////////////////////////////////////////////////////////////////////////////////////////////////////////////


`protected128
P?+)9#"+V.E$ANY.BG)2PC,U'S:"!PR:&P@-%,4ORO>KE-_ER#,[G>X 5&#C5I#RB
P<U&'.)_0]K&.#XQU=.-A)O<:@:9#+M^8=543I+<'AVXC/IAX*1*:M,_E6HZM>#2/
P4XJ"*3QU_">-[] D"$"XB ];3[EZ,W@_8:F#5]JG)Z@\:JZZ^"E5V5I&3J?&Y'I9
P%C^BAK(V1@D"XN=.^#8"%ZN1RZS8S=<D &@^7Y.!RQL'DL(CIM,SIFJT@\63>]-%
P0[S7(W>+@:OIY\LR,D>PF<V>^Q\N3&^T,OQVHU2A>OA+Z)V^T[*?USQ"\[YN.,S.
PS3.!SD58>55^T>?5OH#!R6O]SW4?.HH@1IIUH;C3>/'5I,7C/@_ YNE6QHNPP^MR
PA&+3*[GH=?OC?LZJJLL,B["9X34<"99V\%/JE-Z<F\\6"Y=-=N-OAHY?_>?T8KAO
P2(R0(>3?/-@_]V =J\@4^"356B;9I)^D3VQMD!+RX,F=+&4 ^IB,,TX4*45HU=[V
P75M$%NWB5=5BB33I$.B#HRO4O9FY]F;]?/'SJ36Y,!@EJA99L-9*>,D-E6*U4>MQ
PHVYY%88.-^]0G\,!,!YIOT,/5^]&DNAL3=5W$S6,\]-CI@,^4G;VI+FYU6>\31Y4
P[N>,3D2:J@?*VO *N6[U+C=Q>H=HN"F[I,P<89-TN;LQ5?OHV.<8Y\E@)18I"\D6
P9H@ MY*<T)7UL.)HO)"$4IP5U"C!1YDLGSGVLCD?RLX]8?JP%6(FYU0*K0'SW'L3
P@J[*Z=7CJMF![EUW!DQ,"?]L@\-G!@]>#:+,+2TI@;4(Y'6A&%>[FSWN;/ ?!F&"
PQ%@IL@;_7WH9O"ZK1N2.)&LV,I*7KHAB*V;=ON50@R4[T&B8A=VU@(LLDTCZZE2B
PL*8EECG%75XL8;;)L-4J2ZB3EP&2Q6PG&>Y!^HPGC4CA"@<745(1$5S$8AQ+RB'8
P4,^F?<X57!365U )K0!/GO/:F],DV"]"9AS3PVX6-='I2& =5B]$6>+RA!7#U-)\
PC ")3C*J0&+3)0$X=9EA6]-P\L+I/Y29B6/V%_1%Y LWQ1RKH<$G"5>U(QESO.(F
P04GO"!:,U+%8 0&S(QM!+5<)=9%4[<%ROV":.P-[!%S=XP<@)92-X;D%X>VD>+0T
P<!UU:LPH, BT+\Q4GXYAP/DQ;;2EE*$S'BKHP;AP\11B4F:Q\-"[_TQ%IQRR>R0&
P;M=- !AM6)9B@8$_<)7U7=RKI2N!'WN;1VO,P?B,@.O&<&7U3=:?^W*HSOM:DJDK
P1>KH#FBFT-'18U,%/CVR\P^*.^0":'<XH$JR6?/BMD$6(V!5,N9$OVKCR<"-["C8
P6<E&,:C_#^)9[:C@82'CH9HI?.!5#'3!*DAL'ZO,LLM3\;PJ5[I3*16:) R)S('8
P^(+\QK33L9MOW<&G"H;.0(Q$P(V(3,1HSOIR,8J]&RK6?!,QFO0B-J,:)C7F'?R2
P+D<"[4 5AE=GRU( GLI-;LIF-H0%4=S #(KMN8D_/"U+F!TN&H"NF^=U V<,T4UJ
P2^AB3:OQ71X?<_G@7==/2\C63U<T"VP-]*!T'\!]^ U8CE=HU.*#8!D->Q_T# 85
PN;=V-@GY[4P]Z6]:C6 UWD!7"*5,#/_Y/_R8S&9(->4R*QHQ3A7*/S7&&\RE<I/,
P!VR8W&O'U.W0*<%&"M4""RIK&V=X_#.0C^GW+]>,BIXK5Y+>/SN^T)I.2M68R_JO
P]IB+6X>>.&B38HGS ;[]-FV%E2N8#R"HVO/^\IUZJ(N3+\!(95Y_M%CO/C C^ 2#
P]$N'-:X1.MV:A/[U&T@XDIM:F,@,=V1(C >[&9IP!Z"4&CK(3]O_F-)-77R"DQGS
P.:%HN?KG%Q.[./OGVG;]!J!=2,7YPUR:7NTZ !;-)6$>4E_+U>HJ7Y+%E83QW0,+
PCA3#5%ZDY7B\(IQS#]9VSS2]BKK-8HZS++4ME@KJ=)*3ZT,UBHHS9X:$\Z"VB/??
PXFM$V4V*4&4M;1'=^#Q4SJNWJQ :1[9] YI]I7''RS<<V;>F"JBBI PD5%G_PQ$E
P$9 */+,7]T>Z'8S!9?/S&EI>MTN%EFO<XW@E9*3\C2,R C/%CX*4]5T:S<5ZFV#+
P$**CQKJEX+XO=VS1Z W8G4U39A+^L]I8QLABN(3GYGO(C[,B-9ZF&@9R9SA%-+ F
PMD7.[&BBX,+G"=(*EWS)5S^N@]0J(M$TI:LQ9P.V,J -J]KJ%+,@2>X32'> Y][Y
P$Q.*1M7Y7+-2<^=?88%4,"@SPAV#M ")S1B:5;,(VFCB+S#(5PI4IUP VYSW<4Q6
P((EG-/0-.T+!C;G>H2@M'T$JLCXU/OC6UFJ1"7_&@_G[,_;><263J-TJY5CB1> C
PEHL;SWYZKAQWSQ5F-09\:[OIJT5*#K#6"M^WK"QFU'7HWMEB1L?6)6 /V1_B.)FH
P:$44XJ[!P[@CAVU@D'(E0F7XR>_? WXUCIS7,H;V[ <K8SB0@__X[I4<<DT__NB8
P669&8CQ0H.I@^[KWTL.@#6I-?QQ*\:@X/U8<5F3/'>,="A4FCFIUR\;BQ";/U1?F
P'5@9*)7SSK-(M\.?Y?F"'>U@@0> J .SBQ::ZD8-Y9X25H>93WDP%E)072[2\#HL
PTP%P)GIL+_2GK80(@.PX-T;.:G?77KM 5$<\G*IJ1(2!A5OIW*VE ;,[649+.BD/
P^.ZX+="DD@<CZXMK HT1$O!FBOHA=;ZLZ=S(K<>>>.C#M[FT26BZ-\&]9C8MUG]A
P*EE@,WQ6'XRQ9E%60N^TY>HQ"$I?A&TB'=KTJ/$_(60B2&U-_!@B):RQ+F-72:5Q
PRU1-H#^2B:L9@=4.>Y$5.RO>LN=71VG23DV*!NWF.R!-8',W7,S'-&)6\0\'?SL/
PZ ?X9+RX]2V+^"59G?X)^WU1G317BP+^V_>R7Q,6??JC4J_S.[A5H*! H1U_(3/H
P-^<B%WP6+O]V$8]?"("/N.-R\)$?R_G^)OZ-$T="!&3"6L65,B:LE-1)K/_+IA[O
PYS*C0L9S-J%:Z_=?T=),FQH#5X8)(:%94/MNW>M]68]3(?[%=_,.0DBTKTE88Q>3
P$,#D!SNEX<O76>?(\?(\!TCH#^TQ,)EET,"-HY 6Q;ISQ3<*<*CTB="K,B)VYX9D
P9UM49].M?-BF:BN6F<:@RSG1G+=:6>:'B!8\-:D.Q.]1Z2<^RG -\87("932/_?.
PW@V 6!;M@SC8R4T0O%4>@UG^ \@>^$6H',/NC;=P;-@AS_C5*)77=[KX?7; TI)B
PDY38LU8GMU"YBSZ-3@IY;+NVA:S]DM+EX58]2@!CWGOUVI?RK[3I)-T?)YA9"HP 
PL<NT*HWC=6.E ST$2A.Z(R CF8Z0NJ/CTJ#5-5B*?J(USL8WKTG%T-(>69UVKVN-
PS$=2 U4F\O[2_M^@3;_492@YTCXIR221QX#7F(=C&2O&EL:=!E,' :)_&0:O9 O<
P Z0>I+(-L(CI0_PS5B57NV=>.<QA\TS+>[R6$A["6LCZ0T),UO%T9$WY.*(Q=B@L
P!5Y]MS2X19]FK<>BU<*H01\SR1O#C2#MX5YZU3=WRW/^'2O("R@H3#JR_MYI/.$6
P-_>P3>TH)918,Z)2(^5.2VXM4N4JYX_IMO%*,:/)PN#AS&R>*)19L@^M?'#/,Y>3
P-;"%E5@#B7F7AF ,"-X04,]7S)W= N>LC(:\[1]L8-'Y@+?GWO&QW=0U8Q0/ X_N
P4E<Q&H ;\BUN' TP].N\(\'W:ZTA8742\>Z V?XW.!R^U@]^H1Y;3\]D/D;Y?)9=
P\7+&[%BMO%0%"D=K 2'#3!"02 FYYV."(Z9 W$R _AMV-C,;!4(6S06[0] L2(TM
PH#YZ?D7KC+F;J6*5!_CX*2S7G^&^D#M"90YJI8QYJ#A[N4[LG/5$JC(>Q2@,V&VN
P="&%DIOET)S0XA7ZA%@ JUT=P/T\D+42+)\+D@$E"K',2UP%4;^3$C4%M0IF>?&3
PTH;0")$6"?M5"ZTM-D&PU.TJ2M25IO =F((*KN)"/_3W=5%.H;VG/*J\^#SZZRZ+
P17#MGPRT%-VQDE&"*M6>"HFB:%>'38D3)_Q!02>_D?^SS"9_Y2D'XHEWR(641?G(
P-PA*-.IJU"9[?<>Z%8RE5*M*D[L+K>5/,>D_AZKBB!,V;S7Z@'TZ+ID09CQ"\?*'
P$\&_$O:9H?LG-T+CH^J^>AV<:M+I*P;]E1H&4="R'+3 [*LIMS$K42X!+S[AP^[9
PZ^E/;_$T<8<@D/9.9B 5W^R?1ZA$=;YU6,#M_V&$>W^[ (4%VY;@7:INBGG/WH6O
P_MJQC_S$225%Y39BYO%,91EZ*(S,;2_,X:?#*X*^BMZ$/MT#M0%)\&7#[0J9U'95
POP/MZK4E1O\W/>+=X^6><=ZACOT*>W&>SF0YA,W3#AF-3+VF/=PSR[X2DD$W?5BV
P7#]69Y[85)GFTT)(;Q86CM;YG!=VY!H W1:F5#@0$@4O/Q2("O\:O,8O2NY#?E,O
P"6>P/!0%LIUE_+D<1YW#=YVY574V%<)J$.  +O$*PXC=2[/(#V*'$[G:Q-6QC.B;
P $R<1-00-+-]LZ"/47[)6CS]W^Y./#_W8$.V*$%2OWS>E'%[.0:_K>-?R1AQ"%:[
P8+CV[+JY0'6Y?TO7_!Y>"$(TV;KWQ8"")_#:2-[N4WBG)V:2A7%D9ATU"C7CEU.6
PEVGG2U^*_4%"E11<74;L:"PRH@9Y%;D1HM7,0@L7ZI1+]K)VU\(T;V[Q4YI&A\\$
PBL%9$S:*Q?6SGKIO'>/::G+?;;-RWG## GR:Q"GP0)1/LD%B'H$>+*,019<:\@14
PE20&;G_ADU*OXV4472R7^2CBR\/GV JC%T)8X>[#=\@)'?'U81^<] !(7KP*<*="
P5-'=EMTOX*UP/3+Y[AHK?R<F98XE*E1A5[NB&XD?HDDEBHTMI4J_#*'^:>Q)^KN:
P35=EQ\_"K*><BY%S[75L^+.0-5&]$0XK MP#1!1U6Q"FY]D=&2#!'HL3SA!LXQ@,
P;TYIWX,% ; DC6] >!*,%Q$MDM'D'>3*HEO=OAF5M#Y\*<,")4.NZ6%"-X0\#? I
PBBH47P2$2'T(2[3B25R"] E^G1:S:N$4Y9NU(^5!IY]$JRQH-7;;1C0+'9(4Y3%&
PK-+KL*$)4.HYF=6.7[5UVZ3T<]ME=(AH88GJ15S7$]P0,$HKP;>-U^.OJ?ITG=[!
PS1BZ)8"(K9E"&&Q.32$2(KMAL+!\9JAJ: =0HGU/3L'&,I1,;OW,5=/'Y -!_N,C
PL#P/I-,OR![HOC4/)DG2!3>7C1U;,1FM^2C0Q"5'I0>[BO%.$0G[CB%"'')3G-K>
P2B%R[&,Q?@?V0;B+,H&N1F/NB<KA:Z*(['QA: ;.)F%7EQU8^T"N7C_VW.TU S1@
P-">HV@(('ZV,^@NVN5PEC,?V;X!G+%U/42(/_4_B:=Z.P9F*(9;=6 $FN^K?<?XO
P:7AH<[+O&>BL!+7#*YD.F\_&<X>EARU?[+&LORZ^WU-_,)?7.]H(@;]O#1'$WW6Z
P.M_QB% S*:I/VRPC W96)Y/9PVS2']LF+,'-9+"7,!.R]9(O*3=0$YR#EN3_06-+
PV)QG6>CW&>S[WP;CGW"!*9*/Y3[]2L[Q5IE3E1'" Z.S&B(3MUOKKQSJ,8[\BF>%
PR^7(LC+<+T&V::48I(0I8.]-JE0*,>U^J>",EYWUT:F4+]WB7.\7A$A%@Z\SD'M*
P*VJGM0YF5+6-8?22+J;6($$XHC8 ?R<@WRM&[IP$G$U>XOMW(7BG'F**,#N$I^K:
P/A.>V[/[YM>VQX$+:.L!X\$:^3<K".A:E[OX#AI4EBY?2L&!L+W:LF%9=_]8BHB*
PDL-Y?RM?0-5<>2-G%<&H?,!2U/22*S0ZBTJU?(ZFH#-#.H8RHVZP)%ARL5(@UUAC
P(E9OX"!<7#G9]6&,]I?>7;K/5"5*Q)OEQCN>"6?^G5%$3P*T4A"E%;+IY5V\V.NW
P7O ]QP:T#=#%RK6+VAZ4]R("M)K-JDR^83JG@"[V%B<;52(0?]NK4IF*RLR]3% :
P)I,;ZT.^>_+X>RN>QC#A)>)LLI(T]Z>W ^&>_MJ+SYDL\YU$1()@-5*ZC.<?3:S6
PO-7&R<1KLDQ%"#JSSS!'G%\ -:[%5BB\T8%.*(^QF^7ZM@DXHDI,'I"_1-KZOM*@
PYI=_$7R8F@>8JH'EDG()MZ-)WZCDC!),!QP7N9]*"P1+/+'WP55*Y<LB[5)X#(#\
P4U)) <MWY1J?V/AY9]6'"H$ZV/7]@UKC\5/#6Y"YZJ&Q$SI*CI"+%G\[SC/KO /S
P BFG:U@#<T!38;V"]]=Q&;>%+7F,Y+9T+V3:A ]-WG^R>C<LVI+N%)8D3&?63;9D
PWVRJI7<M#=7=A+.[BG>AS*\&B:H%];G-_.6(BKWH!Z$::Y+1#WP<NOC<%*%B,FU[
PYZ/<$E4!%!4BH='B7[/LHRDVB/J00@6C4Z0Y")\"Q/A4%A4,RI6?WO#,M%=K;>_(
P6E67JR?4S@';H:QMQT ,5YWX"@9.%$1A0^%_)D"K/_)EH=9?!;TL]0Y-3TD-\,;T
P% \2Z&:*U5W#EJP%L]OU%N^K97Q<@^&@,K/-R8CZ#%-QJ@-JP2H2C)LU4RDN"0%C
P5B9^]B,=JY)6A;K#^Z<2 -?;$F986I N S-A931K<Y):V'?9#X26693GCG"C>]@-
P_/(&,GF44/3OX$^8[4T\;>SXC3MD6;^8C6&$=_CN$</._L]1R#)]DIR;M]$/YVO%
PAWV!;21OPOC9AA&)"MK!03S8:_@P1RO#[MT"*X62;?V*\XJ5QDM"-'GQ-+?;^V,C
P34^*4W\]=P<.(P1*A:;BE$]$XGJ4,J5Y0#J_Y'7,B 94&C,&A>/O 6 C8A!)49OB
PGP (WR;PW(LOEJZTIC/2ITR0(A%.5.^.[^8@FD@;QXB4RXQBDW9<.@HR36QI9U)P
P(AKLI:S"OE+TD](<>[E]@METB+@Z4P9B@PJ4QTEXZJWPN7(MT=U.>^.A*-QHI7A[
PV5,!J1@BH0@IB)0.B#O4A[$@-7/S& KO=6BC-WX67-YG]RDY4S04YGS\W),X*W:7
POD$DA@KI'+%@@33XSV$O*VAK#)7KMZQL%UI+@B66/[!=* /?X([:<#S'#[BF>HAS
PHP,+T6=O;X_:S$+/<8U6#25"V0L#@N-US]#>#B] )W/GO?/B+V/AB.%4'Y:62YQL
PN3B)P]2:Z??OCQJWNC2;C41V]1=@IXKYN(DB4ST7B%'@?S)HYN?->/DD/YJ3MY/1
PFZYUP\\ALV_!.2!^,=!SOVA1EZ3-(555DL@OW@P#O? NV^"6*@TQH[[1!,,##'\!
P3F&#YJ<QFW1EY2OG*RDVH0_@?,6>;X))WW,$\7S5TL@"& 25&S(&91?U,::89%4O
P[.\=$W9S2^VJ*D_4M-OP;7,P$0$14##"Q1YW@>D4X:WJ$?2Y-AQD=D5 ?LZ>&K#&
P)KR4X80]V[8.N8 !M@#Z,KSL[60[#>.B+:D:IS!S&%,5,/Q&U7* 2B_D^K;)/BM?
PY,]W0R=; ;B!L:R V$Z.I4#E)IKG7[&V?M%-N#!3$L>]6[A1+$5L@Z4O2#6MG2F:
P\\]I^,'C&M4XU8_0+#AUBH5H9QSN1BN:ZV=BYI,<21'?"1OG"0:"QX NXM_T%6YM
P2#9"E443LI0O6\EW#AMA-U+SV[[86F7;9H;&4GZR[0,FDQ&'\1AU+_;Y)UJT;:-=
P+#/SK "EV=5H5X3,1.?YW/5S.#;]0M%.=S\KP4@I9>=QR +!0@"BWDZK4Q.2#>R<
P:!!@GY;WP"YK*W:L,1SE(3IEO(LW2%6+4SUNASIO0180C1;Q<3L"<HWU*WVH4[ZB
P[3KE#'#L3<UADC)X4(TFGWK 0+3C=^8TQ;W7*3=R0"MZ&G:E:X:Z''_J_E\&EH\"
PPW)25T>#<Q IZ#.>H4E*6X]QQM\5UR[7!6+Q!!2D?N\Q[YF!GWJGNCC+YR VX-8-
P49V>C[)C'(JCOJ<R?VTPMUZD5,Z;S1:3Q C!= X(.4[U5E"J%/83<X'"@M6U+;H%
PSQN$KM\@@3<L_.V;>\B5.HQ)*.MVY:EE#"'2UK.=%Z L<&*0[/U@ZG_86@Q\XSQ<
PHJ)L91LRV240J<.? W> *J6EZ 7C954*I0RR@_KW,H4J4C6A#%&\JX?>T$LQZ.[$
P6CD2KE=5HQ/7[UT(%GJZ0QWD9Z 7G'U@*J")7/1?,:GE0@\!MD8Q2M"'?*6,D,00
PU:KK.<4^)%KO_;ZA?=1?=TS1W)AG4N:D0/V]77<5^9%L33<V=YQT,.A)13):AO3!
P7"O2H1;G#N\7L'"&#&D_6_WX,M@S?W>WEUB4]$6I'-(H7S/1[T+ND-@D[ZEQC:8=
PMFN8OMKT)]IG.[.: (!/9D5Q-;<)U!$QZ4';*KX"Y>&V"JLG.PK,[>&"9ZA4+8WU
PZJ3MD&:@10"(UQ"%@'"N\/?A]D3ZLOYSX_(BL2K8LD8%R 3.9F8)0A-8X)/7Z6HK
P9Q@(#A:P<>YWA;(AI8"!G-,JZY((T(^OD,:\>XO15T74ZR?:HTC!E*5_;IN-%BM3
P0JL:^=>!?]%\7T_9$J^M&)@R5"Q%;'Q7S1!C'#I_^1?7XK70YCKMG:34IV8//MYS
PT2<M&2\K-Q!J1KT5H'>O6'!_^"W@QB\IV39J<V%/<P^Y].K<TQI3AC4ELK$X78@:
P?1;D&950 3E=4D+,R$/2+-P2F8-()(1\T<3ARXHZI#J_<+7*C#??V5.Q#=9_GZU<
P%<'[X,*U*\[?1MDAX%?"\'A0^X;KH:D^'K(<]UB(50<ZP@%_<3$1PJ?)U9WVCZ2'
P>N/K4]KM<[V]7/H21O?G+J+.SL/='M% N:&W6O:1F(5&21#0Q,3G,#-%H-J?:/+A
P.9SX[94BZW?Q]W$0?5BJJ$%T8^IR.R@\>_M ]D !?;57X#2:"<"BLO#NMSRF8%[B
PN1LU.Y SI;$FKDR,Z,CG4ER3VVW].[7;M44Y)/DP"@:S6:N38TAU^RIV]Z,!\2:F
PV.DH6JUB_B0>V!OA:8^9PI40"0?QGJ>NV8-^^V9.W2'F7=GW;8==RQ& MA)]Q('A
P7V>0;.RMI-6)9\U Z:7-=AL-+;GL%LM$067$O6RR$_5+MSY4-6H>H1W8G]S8N[A 
P7+J<L*37W:*_IYW>,K=!#U54SY8O)BBJ8D2DN@K ;%B(;%UKI\5C,[8//AX](G<>
P*S1K"N(\]P_^[D6=LF.,G:$=M*@FI,*\VVS<2/_!"B1;S^ SL32,HW9)FVL1-F:\
PN8AAI]:[YZO-(2BJ\>+2Q%&+5#OX<%@62'ZKK8G8P-G7%3%W=IL S',N7?&OKA\?
PN\,Y Z^RD7#<)QY2$]0_/XSC:$&FZ-/@#?KD0%&L7A"ZS<K;KI[^F^1,.Y>;!YJ^
PQ)!J,C_FNP%5%B(<O]S9SR8!77VM@?O>-G>,6V9G_1*A^5"=0?D-L+]LR6VC50=/
PX^8K>MJLW<'46T^Y(?4+!SP%K"46ZLI8S"*R8GNRAW+1GY 13N,F;E#K':2ZY9A;
PN F0=TJPE"!T7SQ"H9F%14QUB9@&D ,46NHT%4?P!&Q,*4$XWOO?YA*7_0I_@D]'
PJ/K^,.-Z8F(,HGS)5!= T2R9/X!+ZW2P#"])V72<#UZ^VGT5:K$#0G)C5>M4 B5+
P]N%?%O%2$('@=0)Z[NG.RZ:;J@L]TE4B@[PH[(Z9/&B?,\:!7E9A5A>5]\[L=KL^
PAB,0T<1?J_9C91TLV["B&I 0,0NP!RK/9>'G@-Z4,+#8KI>;NCTN>R1T )T> ]MF
P <4FUMH]DGQ3F>L %[G>QK"RII=J@%02X5&#<2?D\6C70YMHJ=L AER$=AA"_D*W
PCD)[Z48)211ML5TMM)^- '$-]-(;NP\(?;(+Y$BJ:F /V.I,XW2*FRB7+BR(SMV_
P9!L%S[7#W7[B^U (/&T<^!;^K$B"+Q<5!'SN/&1C#<[U5P6A[,_^5_469B^4*@J;
PRP?C\^U<%D&_NGY=+H?-FI#&/\VS!0H4&-F.MCI_&M?V$@&( :U(>WA^C8A#([,R
P9)LG;BF)32]XN"G\2E#2M$VU;!_\!6I,-03M>,:\HZE!?I/S1(^_J,"']60=!A[D
PI%T-H"\K_:<^<J4)WP%C(4Z&(4F@4/C "K<YT5>9OD1O3#=K+Q">:]M&,/]^+J@F
P@MX]K/(8$!=X(T=S-6$=>6@F[=TZ$R%W;2R#RGT'7@?*4E;LM]<Z/1/Q-IQ+*=]V
P.L*(U]A^!];AF".D1C/5YQ'99FS_F2M2'YWY?DY4R1<6Q^D8<B6R+Z3I(UV[RQ17
P*@_ST4H[9P.MD<\84B$I3PJOETJ^;EWIM#,H&-QRK2 ).ZL2LHD_M4_1S]+59/?;
PEMMI3,M7[+MJ.HR>\ .SGUN114)0GL%2_Y"#,$-)$I[?N.Z=]L#O"!\QK-U&B(?;
P@C/V3! \Z%@LP/!0 K?;D"LVT1&H.\)ZS6S0TX,4M^4?P'18OX^IE\$*%*-* @[D
PW+K:R<%D))9ZR-A^@4JWU%$%!T_OT,@NJR.^-!0</C)VJDG+]V]QZ=Y5]TO 2S 8
P(5(5K"  M]PU.;C?T:)D;A*)7FTN(X?S ,5FV0WYAN]S[1%ZD!^LUR@%P\RROSN#
P:/.RP;U)!K5YTZN"J7 ;/%+*)G;^4J52WR,^IG-I<^_KW_R#70W,US^,&HX>WE8K
PX <)D,LE$$V^X[QE<<0G!"V]F6;)4]OH">Z? T0H41!N%FGSRP#+>11+*Q$WX)-D
P]PV14?:R@[YVDP!TW;YPH[1OL!X=T,7%H[D>>O!-3F2?[H*#@=]TMY<:HL7=^ISJ
P"$B_#:T-;MZTM7$+I]H!,$?)MR=P ;QR6C=!XC*/^][I4</TKT$S"S4>/=<XL56:
PZ7TRM22IX;-"1?\F.T08SL]W WV>&JL:R;G$J<QMP\T V_DR 99]N$5WT]0V>?H:
P"SP4&B&R^]20 Q@K[Y .^PG.OQI1R[['BYUQ#1;2')?!WWNB_ @T*]$.R^UXODF7
PNP_J&P7YO=$3.<0!!4,N9'.%P.M'IN5% 2GAT%NOP,<:C1_0MZTDEU,?^B4S$,['
PKET0O,I+:9R&;M0:R(/K=\H@D++EK?VJS(DDP!'F:@8N<[UN< R%4-^8>-#@E1>D
P#,W2A6G',SK;533Q]'1O9+L,GV"%$A)WFLOZBU!^'/I3KB/V8G4]F%$O<KAWUP<K
P]DI4&PCL1?]4-L&@8L,)DE1"NTPXW">&)PMDZ69HTV#+2IVP)%7T4:5Z/?OV#$LE
PW@*AWL>#_@^V/XUR(_+9-?ZU62$[VO* 8I04T%19:.$SX3KGT8G[MBCF07!$P5PY
PW\YJIRC:MO&$O1 P TZ$<XWN*$[-Z\3T'F0==HH+^TB\W[3RR U:/7N6GOKOP.):
PD+:X"4%<"W&_\6=S8X%?>O>9 7\.?&PSNE6X!OK0B@(GEUU,LK!_D&H"P3#SZ2RF
PLMKSUCZ)Z'W:0T_R8!L(Q;('Y2KRE5N[EAQ7I*%MA&VBP<0/8)"<J;*&=G)$G4EA
P](+=C/<"GN\7G[F B#+ ''':DV>:PAXAN(R&].:M\,.ZB 'AH@*4(SG7.L:IG7;7
P%W7FLESNNR*P0UE!ET@J-'U#KM<E1C5[\B>GX!U@=X3HC4XP!M93-&N +GSS1==.
P\3\M/&L\3A<;/+_#<N![9LY*\IG(;M%/8LMV@T1C(LA340=HI@A3O,/'BO5$K$,5
PO"&2,[E <45)(4_T['-J6:J8X+":,\:)4S8,\XUH5),N/,AFBK?<\E5T[1K"SVL4
PMM RLWZX8KPZA"^91-)X$B*]2/AR-47^V$.8!A_]#(!)E-O+N2@RWQ:6-+"-Q_=[
PL-]8OS0B\S7^$)S\)OHW*UK__Y7'G<_@U^V_I'UA/2!DO",GPSL@#VBR)/"F.[:<
P#*Z<C^@=*J5I*C1>,N%NO/%R$-';\YJV#[?&0A_/,G944H&(\DT\U2N_2A5<ZU"Y
P)43CN'F^,>*D!.VUS!WX 9C[)LQ:E>+K1+6+T#(P.R>X7UG))P5NI%  PGGF_$6 
P 9S#]C:'*13_:TV*LXDYLL8C++ZJ0<CL:;KC+UK 1'F.,\BFMPXW"Y=\<%M?N+D.
P;)*JEE(9<P9\M]:GX_XO\8K^48+R'J=>9D4CV![>(!P/Z+_.!FIWZB8Y'V_:,5[[
P%(NH*R;4)?Y&U',/R>"!1-(1INIC&9R=U;S^HT?D6U=+^5CLDBB</O)7]Y;KM[%=
PZV=9PZ7R!K_R@C$)HLN@/AG>*';=)*LDIW395,W#_S6&Q'PW_("G3/.Y-&R+O]QZ
P\30!O>YT0FHVP)5'$5,^&YY$B,=_Z<"2BR;;\!_D.DP&V.JL?GV_3PIA1<";;9*[
P=&\&B6P*$PX#!%M!N#2H)D*P3UDMDN<AZJ,O5Z!U'U5X)SGS^ME$/^ZRI(5)KA7O
P1L'X<7O71Q$9#QA<Z9JT.34IXX? 5>Z,' ;AR_AX.'_$A1H2=,,M)_,!9])[6N)&
P+9WL*78OZQM<:VQ!\B7H.V,[VHB[%TF/L!_+(-:.J>D3ID #$:1U52I5S07'I=8\
P[""DI#QWHKN@NT%K-;[M^!?$OL+3 RNBR+,Y_\-#$ H,OSP!9>*A:  B[(#\H!)7
PV&$%T#Z_ 2"Q .:0 *\W:Z-_49():*)MHB!Q)9V^J:C'EC=DS0B)9;[H1 YN90Z?
P1.2ET+FH1$N^@ADN1=5'DQ+'=LV13?_-"P$3%)/HAQ_Z,0'+:'[&/7!QX_D$'Y82
P@E2Z!&'Q3/TX+/W$V?-O(.,RKXAD=>,8"T+R-WF =&F 00,=_U&DT8WX=K:'"*6R
P_IW?:KP?I6*VJIV:ISW5Y*B$VX#0)/BF;.S#Z+RS'9Y"S(3*DOV\XNTM][W2W2 5
PZRT!*?LASH< J=MAAB_C";2;%:Z?<#RKTK.F#JPCGMFX(5QK?7T( R_O=E/P8-W1
P@<]2@0$7FT<\WZC<H/$_68XM5T]L+ 0WNBVP\6"[D@<7X1A&W!&@E?*,C1>SAQ1,
P%?-9".NF/E0TWYM&62'0)CI->N0%KWZA\.4FL,KS6V7W+D7DM<RY0I:K\'GP/UP7
PDP7>OLS:@61I3^&?^[/MZE5341V3C\-'+"3W5""\.H':%#12-&,VJ'%J4KMY&?MQ
PXJDW\T,8>SL6K_PUN-$ZQNI\[6UWRQ[\L)B[EC+*=\'/B<$R #<OGSTF9V9X6GA9
P-: (Y-9Q/QR!=/[4-,?+I(W$,!*5'O#4+BG.]K9M/!9V1'RD8+UWJPN$XKP*"NN/
P0KE4=G(!T.-^:SY26G ),RNQ-C(%A8]10E^V"4KUR?4:@#OI56VM&+:MSB^M#A/2
PM%:JG?3-=8;<9\S DD (D0&$5M^JTH&=EWCJFH2MRZ2NJQH<C>=2DG5W=>A;-VQV
PQ]L[:YG'])L);/9&7!Z9SKXPU6!G9"9+79#\+D1=%+R-3<0]N58)>^F1\ TVQQY?
PXVXO5UH*8#IY>$;+I1<ZV/1P^X"_M638Z E1PU28&O1M"2YPK*4TC[]==I=ICRED
P%9^<"MX9)^1V@[$LP@!5XW"ZX;;8G6\756LOI+N:$R@+)N^B;S\C R2\ZCEW)H*N
P4QW!6=NZ5]@*X*9(%L(8+EI[L^6)UVW %A3W #*2W_!B\:1"Q@H8H.YCNS%)23U.
PV1+S-;%PNHT&\M;=#\#'?.OY%>.$8,'6H.1;_=W/J.AL+HX&G75J""'?VT.GY(VQ
PI?+9M]VA!_DB_##>LV'J_94UQI6*SI;4*(M# >BKSLR:7R0;5QO/F-6D A^,$"7Y
P!M-1Z>B&)VE38EXI-:HMR#WB SSSPE5[I#NK5#2H[4J(NBSD=9&S:NI$53I'.26W
P,2Z!TZCMQFZD49LE/;%U<-M[>W_PS[565Q.F.?#$"!SY28C%_HV)WX*L''HT>?;-
P!PW0;A/V/#)31FK;FH%D:0E(XP>1*/Y@JO*%,"G1$QO[\4*3U-C$%L:D=EWC1)/1
P.EB/EBU:E7482]-T;<8F=D](^":1*)BTQ?LW8D:W3&XH\NL02 P/<<L?SD*'%2AP
PG\40_G:$V]'F2:'=]>FQR$(A91RD>XQ950^CXPJ*Z8Y9<%1D3UJ;\RH#DZ4S[M2B
PG*G<!*]$+Q26%_O]4$=II25= X6C1JL*-()=\0>BS5_]WS;Q>HH*09^47R3I9E8Z
P72E5SF[GEO8L<"YMO'Z81N/*A)NTNCO$E'V_(AG][H^5>DEC]=5 V@O>H^=O^/U^
P/<S,R"*4C">R6AH:XY?CT/$ [$2K);II+&QX(.BK1W#S'[.^/J\8\[%D8E(-#4YM
PB*+#.(.IJ5@ R8>;0,_Q3/#L/RXG\"LX9XW@N:]7J2G'"!+X'*.!61M"=81/N+ZO
P(>5X"9LE0&2]JE-DP^N>QMN&JO[?CAX69"/7/8F+#;D5E>Y ;^O1[X:NL.K(6(G7
P>-=O&%Q(49H]VFE*=41=I-&Y@9>%DT?>@4*X@>#8\XDT(3446;YQ-F3:4EWN](%5
PBCC L/KOYG9NT%9!WTV$H+E,EY.^Z>)33$,/;-E2LM%$W#P^R:$. *&Q/3UL8PR.
PQLR\5\,&&5^&9!F-<=U%B30[%S$"C4K,7"O!D<YN'426BZ?W^0SQ]GK3__;4/(%%
P*=J$"9KJH'R.0B -MNIOKFYYIE1,5CRPE4]P2/GN#_:HE81KYQ^$C,S)T@&!U$,B
PHPV:>I\Q-5&N,K,%3MNX5!XH=\HCW,^R7QFV=9+X7_@I^GC>)-+T(B4&>?&$P;.;
P&*BYMF@%S#S]X&,8%.5OE) ++9/Q-TW,=@4C_(5$-S%>-.#39"<+]. ?A+>4NINZ
PAO.Y/X"*(P 81FY;VGS9F@K@%)(YA\"07O,E:P8--./R3F3'#OD@I,$9M !KDQL#
P.V2G8_]4F9\&Y<IGEW\DGUR(T&"\G[7"G>>F&UON?I=02=E$,*HNG$3DK+A",2,-
P+'BI4,O18>5=D?A4UO(;L2AI4'>CK!]KD+;ASZ*>') FQ)!K2LG86U!D.6^L.S<*
P>L^-!MQ!17[&%C)_RV,BE]]<53@4<" $QOW9V=ZI_2I*&\5H/ 9TT0;9QSYN;A':
P5D)@6_IE/C43OC8Y.Q40Q<Z3F.BKD@X8"40GV9W!ONVLEG('#7QWB'87(O,FB>JY
PR4N3RRMO-&5MBP&,UGV=<9:8^Z7]7H*?#J^!8E41C3$KJZ^0HZNDTEK@HR9*EHT_
P$=(%;(X?1I-.]G!*R\>ILOS\X/G94NA1A'V&!D/0CJ0OTQ&D5BT$C*J2DA]6M@NK
P:4PMS7GQ457HP$XN>/+ Q$N :(.3R9^4^9@Y)"%IW^<-6GU? WI(\T\25]V>R&"Q
P*^D]:A=A:'!?W!]W@!U27L]X+1 QWWZ_ZR>M+Z/HJ$GC=M?:MM^'HR2WC[9]S@CX
P=J/7_YRNLO5]ZNZEYF?8T]S)!G6#\FJ+:=?'B,\HJXB=N&4>R$[%K%'U*G__F4?V
PO[I--EF;YJ^ 14C&%Q9;:=![3)]?1#N@;-8P_6+552@O^?W$S<P8 TB8QMV#4=I+
P_3'8!4&]J]^7F?Z2%VK &IU&DINZ,96/$9R/<&R!%:5_0?*HQ%D4*T3PN^[6GC]K
P#J*50G>;I$!,66CG<2U15C;X504<I,!@J*0_2[]Q!;O',PA8!*0I=! 3BO)+9G']
P HW]RWS#3/8+VA'#UN/?YE"+R/+CTA?#W/FG^QM6*-*=@_=8< !<XD0\'5%,&]\!
PD!#;E".M-FB#*2CWD^6]A_._A7S(PIHHL( 169%N"!?>*K8US$,!4(P ;'PEQ\QZ
P3]\N-HML;O_K6H!U_]"7_[3?U;A:J5B!$S4V#EJ&:6=)39?TS+JQ[Q]ZJ]ZDBN@2
P+?QK30$]/9/S\58TO">\V-VX4!G@@%*/C_E]>3H;.><SZ-E[;??-[KUDO6*++P?_
PQ (A?^\AL%.\+(L%%-:63@[5C\PQZ=[YQ^2%[!I&;C"(CUT:;A,AA%RKK:"?=QAU
P@KSIWM%<"A2IRZ\32PF[.C-"<HI'C92S* #^G6:**F[W/#ARP*BA5?Q?4!XT(7#S
P[9C2359S6(1\J3O<TC /VYDFG2 D9)57:_KEV#+GV0U_I;;G\MNLK4+[H.0V#9M^
P=/)0_4K3X^7, PT.LEPH@4KDLG;C)=%@BM1"RT:4U'"G/>:YB/SEU?N*=;<>+!MD
P0Y2OOD#QK4%-2MH9FNEXT?XTL5*S$1^[Z/8,93"S%F.0*RZUJ!OQ45I8RBP^[>*D
P60D2MH,115V").D7"^<OYJW1#0(2L^ 9V'AK/=>1B\=.Q5J'/H55][.=[I3HS\'-
P!K'UB.<C8.P+P*^$-%B\"K_,!8D4U,P9]9(!:B.CZ5YU(?"NJXCZTW7M/,P ]J/D
P4"?G).%(NW;;']VB0=G][)'^ATN92)VW>U&"OL!3EON,6V[6ETO37\)!CGJN"H*T
PT1IE%.NBY)9+T8D.AYTV6D*=[2\+N5$;XDX:]'5H7'Q+MJSDC?!)"+.EYQJ(3"#:
P]= Z"KBM2_L5BD%&9+#L'*8H)IA^MGWTB[F66"HK\TG8;AC<W<3_$(N5%KC'KH^%
P#!?8#\5:=(MD)!\8- Q8 KB(124T%K130W.LT)-*4KDR@DFA_?["NJ- /86U7OIV
PNH%R[P]$8@_D6 ;!C)J2@94Q3DR.+W"V)8BKU:0G$3<<',&5*'_5W<U1X4F[$*G6
PW=>'L"7I3(*0HP$Q3&"#5IA=@IAUM7]$+*,;4OX*[J"!,2[G*!-I%71AS04GV/J(
P 8I_-2BX:1O%G2* -FZ^^@+;8/1L,>1HFXAC<11&L9R".#QXL[%]]+UY&N@+PJ1H
P^,44H[MWE&$4JD%099SN:^_Y1SCU...S(^*1R]%C&-00L7>K"7D^X$1]^@Z*;ABM
P]O!0<VB<A^;Y2QK=AW@$:1[YG(O8)NO?E'H3<C![[LLG(XTWC<Q\BDR8E_B9'I M
P<2G^"SR]7/XB&7@SD%@B5(EQ812PA=VA5PU9\28.=$U8<O#[RGR-4"F@5R3[1\-T
P.@?N I:T%$C4=Q+54DJF/?QE-Z2#/SCFO"UXLO)FEBZ^Q9"DQO%'%AE/(]H^\FLB
PJ'?>,TI9<X^1W]E ,.? 942RD*(4K(2A+HT7I\)>Q-G#SP3#FC7X&/9OAG0BP)<E
P450,PR)^O:S^G%VV6:7/NB+S\6A3B#L+-7H\=G_UEU!9 ]5S (W[VF)LPRSK/6+P
P&,52% E10L8YHC//;TF-$:'$&O]QVR>QT&H[E*'BV6I@HAAP#4,6+N^?GQB#CV[5
P3^[.A^F+%=H68T\:Y2,@AK*]H!0'P&X9*_Z(SHWS,I?CF_WN[0\PVP4K(M0MM*]T
PRUR!"*)K)&<+"M^*>[LYD!$R5;+U$ PPU6S-@S.7PCT&ZK5#5$_9TN6N'1K] Y,9
P #RQ1)V(U&S68E3B*,$Q\\F\0]GZ^UH%"-[\3*'#42Q32/LM0:,U6YB&$\0)"AH$
P^!2X+S;VU#&P/<Z9\J$K-F%J@]2)/GK "C.^0T>UC;R?_$6T6'/THA@^!X#+:2/_
P-Y&M^]H3^M#H4B#K!;T#-2HE]B1T?Y:NJ)$3?<X<5S.<&4%?^LK3WS8(^X3PTXF#
P.MKV^7^)'<!?:N[?4L0ZY0'K2:CW1(I8* GS5PG<LJ3&&IZ^]M>;#-E,SQ&&"EN<
PV L#\.<_G(,AP:?EEW0MHW=)_"_SJ3/@($+,;@)=L"=1_,69LG"$ ^1/E8;_J61;
PM_^CP-X6:4J]Y=V7P_ [<:81PZOTO4[FLX.T=0W[AD-ZKN]R5C"A%$-O\U57H!M.
P>T[AS<2;?H.R;U=5W3:P6H -V$9O-]3NC1QA7HH+%\FNL'-<";%)">%%@"LQ#A2-
PL ?3:A3LDLN4L[V:\[P"R1')G^4B!WCZ<K</;OPRL:01WY&Q=50:8]H,EEVC3<W_
PT+1AA=@HFO:8]->.G(5YSN>^I%,Z(, VI:M._> AOO7J[-DK=:Y]$O-KI6\JT[U;
P]1'-+=&ELO%4\>?5I]/?IZ?#-4;X8L.G(N_ $\_58YDL3&1?985AT\7MZSZ(X2&E
P+]ZI"+6^5UJ>:F=^$,Q4-K$X:1M^W<MX"",JZ4NV_<6G=,$-C7FMB7MUQZQ*?W8L
P3 \<-$/HB[NF5<-K! !L3=ZZ%)JBY@)A&;],'28II;6C&P_U5>>G\ 3<]$2<,AD;
PZ2.W>>W AP"39 D"F.X#W@_!1A;D$0@A)@\CG>S+>[)U83_K;5O,WS_K%BN@';J,
P@,']SB8"8$CS:9NG7E1N.2)&!1@**U.';GGNUIP'<6N;GS*:'[?@B6>Y 2<<ANJC
P=X3JV9YF&U%+V@I#Y!+*M&0)(#N]3,4%'$*' 5I]EHK,\&O60=IE^VKZ#Z<8,PK@
P?<DE,?#@"D>(C[;PSM-#S4)+^)HCUAQ<.H)AS,)'#=-Z9D4%70XWD;?;NF8A=6IE
PX[R^(,3769 QMFHTF&)"+LY-N%N#S7AF[#U5EQFT)98-9@6_^]#M).A.[? >JMUE
PWR0%X;[8%?1O!TE4Q=V#.""<.#7L[ZE@Q,"B5LBA15J!Y262SRI.QNH>K.0Y9$[P
PK7U>*\Q%3E8<O"!LPSJN@Z2VXQ0]<Q/*TQ3'U&!\79^@?<M5 0D221D=&30[)X?P
PG!$^N(>,?"8[ S20HJ,Y&M F?U#\'M0A<XTX[_Y.J;>P#/DIZLL@OGXJUICR4T<X
P"$%\VPZ^04,[-HQ)2ID.^HU+?SAK*3C'X=!IG/3PX B/N]?4LU@(XOCFZM)@/L: 
P.,*3XXW546E-KT"ZG.#=/R!=@FPQFYVJ9:FQ#:H!H(+@3*@HQS/ \B?Y5@"+L/FO
PN&KO%QC@R;MO(#2.KXVBV$K%?I+=N9*]#4\,^WC8KA K<R3^F?GT'PKN).T?]DK$
PPV\\]^?(:M_IK8]"GT6ROWW5:Q.0%D)X#_*1@OYBEQG@^B R#&0N-47-S<<$0T1"
PG>96+VAQ#=, 1HMV+4+433VIL[GK5=6[-Y=8QPA#JD 5UEBL#4>1_,RC[_>G/?'H
P^"Y\W,! ';HX(1;.1LN"C*4X;L;Q61;@M4(Q28IY".O=N.P+?5_$_.T(Q,:0F:N5
P=3Y!%[$&S;Y8_Z/_<0A6IYAR#I>^Q>,89S458Z3O[9YW *FD5X"H>MC6(EM#4U5-
P;\3%U-,%4HP8J(#P,5/7_C@'N Y]NN;:QQHOBB*)MVCJZLF>"#CI,<Y=/X2?>_I!
P_GO6("ZWSIR[A]OOZ@AY5?=Y#FZ:MZAK/)(%=1?.RIIL&:!6,VKBV8;_IQQ1L;NI
P"FOOX9^B.J>ZHG&6/1JD/<3!<6=PZ+BBOW@'")O&X9:3PQ!_)G1QW@D=A_.RR46Z
P2 5:_Y!M6-/:,/6^DL-V!176Q3!0^\@?!D+9ZT['5N9'%/NIP1(.>@4#_#%=@PB7
P4&:0F618Z^@0.0S9RW?,X'SOB']\3//#.HKEQW.N,6VT\20DGT=5,5BI3:)+AWR-
PF?>PIY<KF:0@0A&'A/@K99I1=QH:&- ,PEOW&+WP&(-L6&1&SL1;/W)C@3QWJ!!#
P.8A?1KVADO&I/=XP/I%&?+I:OY#.Z^[3/DR27(OQ^P@1<A=?_P"_8[ >2@8E;*>*
P*DJZW._(3*CB/=4U+.1J$]:"<PB)%-&75#J(Z:4\)TVP;]+F)X$"3$BO@A&D3PCF
PKE\/^XQ6+7"TI;P0;#[UK3/BKU9_RE08&SA]%9H@<0@8,M).D2QKQV(6<3H16BAK
P8B-J'-*?M45Y.C+BW"Z;UJ\-'5FV(B13X:8"NVTN ]%Y0H L!4D0K6*:MEC%7M&>
P\*%+=V1: /"(]SU9P53?EHJB"7/Z1TCK!D &)7"&1 >]&C(?-O[W8,5KJQ@:P!,)
P:+*#0_)*#KC($]4$%6[L>E!J3#E> ;0I8EXR_;2)W."AJ=^6@@+),_#&\#;:/ON4
PAIUW7:?$.[='TH#I'A=.O9 >AVV@<WH]U#\>8?^HU_$PW!_J@369#.J%O;QJ8<U,
PUR2;F[3LFNBY<>>)OOSP/F 0W#@HGZJR8,S-FD3;02)OE'9N^YIHX/@^I*_R?N_A
PW?,2#!_0I-< #P;B.!WB0*\:T X/0N-[CZYM71T!UTLJWOXKU^FN%I-DKSL>2,EH
P&APCRN7Y/XIGQ,Y'?(!/C1SKS!=3Q%;Z=RG EB2C%O2B%_XF(?80(=^"IGMPWMUM
P(G4Z0#"XIK12:N&,46^$$-NJ87-TC/C%DW^RE0 ,_?4)!087O>YI0SB!B!*05'R9
PQ<6*$24-S4UB&7[L#?+A:[N:S,44!ZRX0QV55+KQ]7DYJ)_3-5=6O(;GF, &:G.D
P\W0\#3'_<1K0WKA$D/ 284")+%YY>\+W7$ZK8/!VOBQI:&I4#]+>-B 124A3U"-F
P&W$7'8Z'(SN_QSN0[!M)UJT<P#0/GB W*X?O=W$2;V'B#0C[%$DQZ/)IK%\=' >V
PQG?3$:1=REOU-&*X9V5ZR@#8/Q$CEA!0WRCT(V^H - ,$.33/PR6O!JD:EW=,D3/
P)(ZS)D2G&\7&+ H(7-F>6FKO]QQ0LGMO\C?G?5ZC1_;OPN8/]&-U#*BBMIH!WE34
P'>N!TF,[4&\1+NW,OT!<S#)-57#'5SUO<NVJ[">4;BCU66_XB5<\!24HLN[#. SO
P@XS+D8''KW(H&J^MI;_NJ&J(E.X/68%)^<7XY+WJI=V6-7S$_LDPNH'>P5T4X>NB
P%0#7"^*MMO[HGJ/>P#"62Z-+Q\5)F H9,D,#XZ;+7.MAR H('SPE>GB\/ '],DRU
P0@M0]V)68[2_&(8C!P):8 :XHU.FM ">UT"R;> +AQQ,>3J)S'%4<;2X._3?9&2O
P>OJK0*U6\N!BRP$?L!NZK[V1O!%@:NOX^GV/*P"9<E)D.QO5__FA="\\6E&PU)1.
PD0:M@_9M)-=D.PNH[05-<Q*#*3437T)>X4Z]BRK.N5K;1<# *$^H5G_/6[+OT\8E
P)R@R_<['T4 +>7KT6EQ2>]FH)(4MRG(TA7W88/@S\#/;YA?E[M%+D0K6ZJM]Z'8K
P'S8")]4 =KQ>'43S*-D1^,(-WU/_X"Q1N\&\GKI<:AK2]7V4'(LPA^_)^?P$1/L/
PL)'S4@(1.WL>0)4POIVU^+.]CW[B2XX^FQM_)?&5R]G8NC8,0E+!) )%U'0_G-B*
PB/)J,[WWJ(9T^+# EM%<G\T-RE2H)V:^D8DX7$2PA;(4$1/$RK7@/2E679?&'9*"
PDU&R]XM.AW_W^H7SE\E["+$[MR&1Q"?/_7)S6)#/58^=G?TYO8\_>53\QVX58%_D
PC?/RWO-U"V?$N8 H,6H)"4BS=LWA IFJ\H+)#R\RI_,"F='WWB$Y**,XT6>?!'@0
P.:?E2CE=B0P*U&>/]MQ1\,%M4*53;#D7F.EC/P"@K0@JSD%,@@>HZ!A?K6!\5EA?
P$_SPN4O.5Q6*MYY>W];!C/"&FLN@/Z(^99EB$,A#"&'2/;Z0":>[\,O_9>O&OJ+=
P[%2(Q"2;-B0Y+JT"F&W3H [)";P,[B)9"66 #S4=S_7WB)8W@7*#?]<DK<;!&33/
P(<]-?VY[+M_\W@Y?9$*$FC^H95?# 3\_UH?$W?CA/N$+ IM&Y(OH_.@7&XSRS6UA
P2<%2R=A!9\<Q>7^Y+^)ZTZ9O;-*=B3"JF >T[_N<M4*R6>H*;7F[N#-784O8ZDHA
PR.AYP&6AX/Q<6;@_!\I3B<4*U2BV:P\BX79$SQ,"F$, J^MFLR*MVV]3/GAPEB@!
P1S3HS]\#;CX.!]/G=-=UA&.>L@F>6T&4OJ3$_DH$QZIM\FT%VZH8#K$USXD%T7E7
P'L6-^5CF^8T; >2VS\@49>[Y''?82Q+))HW_Y;RVZ2F"&^3D)7KK%G K^!S&(!(Z
P5C/'-8D]3@3KH*E&-6+>+K&QN>62$V(^9UO2"A2O$D2;<M69\1X4#@PD@J5_)*+D
PO7/QQO7+^;O#FY#15(.W%HG&#CB%@NSU4+CD)!'FJX'Z38%I:@'\]$ ?^BWIM?SC
PP6X,3#_GM3H?0+/P))(,218_>,7R9*U*I@AZ)OFHP5,NC8 %KX IY7%LR140F\A2
PV#(^9[\XG?DG]+0@_2D$DFOJIJCOI25R4A,@:L>]:],UT-L(EFW56IV\+<)3I8/Q
P:P1ZZ$;HZ2BXU Z\JGF?1CG3%>D4&X)=5V5V=I@U]Y&] F@.*D1&'W6A?(Z/7+M-
P.W/2RF33]"-BO'"IK27T09=<'WC!)I=-LPVGYQT(PV!4J:2]T&W9) W,9JI&X_9?
PBU&CY1VEF^6X(UZ[4[\#W1=TYT^!]'")R[K>--3H?8-*+E6+V_$C9*7G*4'[&"=H
P[80MK$D1(N9 .?\")$G'<B7;*T(>E^$SU>I]M<>YY*7JE9Q6X!N(Y>D["N!Y3DJ:
POR)>T<-*I?K*D/0W/:8#I7 -'3E)3>8$0D8$4^H>/N3@ 2V2@>?UIXQ1;S5)?(>1
P-A!>9BUX-E%%D(MV[J5W*^10Y3,OV=B$3R)+0D(STU.6/:Z<?/@=@],W;8?.==27
PL;Z^?RADWOJ0.QX9; Q/^_.KH0'7J JL#5Y0C1.J1./H0NGKQ,JN#>58O>NZ%+=M
P&?E1AY3W1.*F$:V0=Q=A-U<^,<#2]D@_E !>53^X1H+WK^AE.=_"B$825SSPGIV"
P<[[QN53"1R' W+WDAM\X<CG"G0A9A[Y +WVW+I=1^&91V5=6P5M O39" :<R  9.
P<GC#S2@WDP#X5P"AA2:'[?<VAJWD.IV$K=:='F12>LHOIQ*KZ1'^J,W'6HU:P>]W
P^\I"# BC3V1 ZV0K&+M/0F7!,ZM+7&P^#[/T.42[Y P#@I^0L,S)X10Q?;37_SM@
PLQF2F^T>#-+"RXIKX0G*')67-,K/3#EA8?1DL]E^T9Q=JY_=KG[Q-*P'LAB[]TU1
P;5>-/'$2.=*U:U)ZA&?]\77.E5B:8?[KKH+[(?"@0:]?V?A,<6S!XRQ FV(\9 8+
P:ZHSC\L4)O$-4<%C&Z;@4W8HZ.&PK129)#STR-U'3)Y7NT"7?C^H0M]+N_": TS#
P@'Z/6V(TN>R;GKB,<SNV6G)X%_9;AX^XD=^R#3KNXRL<B^Z"'@8<2A.!<$E5KA>O
P^>BS(Z"<.N F8-[-_.G(R\+H7(%(OZI[+HU.#<T.?S"(;M9991$ <2)G7VA9?MEE
P^4  [GVG:#*(R4$S$9[,HNZ)$YVV[G%$.!B,9G'@"(6^Q.>E;<?O-M+,K.O >&=&
P(BSX:,@JB*?,H"7E&X(F]'+'@E^@(J81P!%G<5@@(@3\.6>=B)7K*24#Q_>LP;7E
PF-C S*L0Q:$/43!)1(P#>9<X2)"[D3(NO,7' 36V5N=@/,0QY('M\<X/0*\!2$(H
P225R(Q5N'H95F:5'M00 O]I%JV"W09RHWB_7C<3A_'62ZZ\)!^31/QIW>E**:9=+
P<J6IYB@*.( C%FPYMO(WDULQ5 4,8<;%C$SDQ+_9(Y=60*73@U.O4/R3J>LFN4.E
P!B"K"EVA'*FJ2P_8J/CGQ/FZS)\ZWH/QA/<K,\RFG:(<TFCZ7]1A>\/\R-[)6KT*
PWIH-?')?G>B99_L>?0K4VR=Y8%$(:C/UB*3:DI2N3%=IYSRB8\9X7)QEUIC=DYG$
P!@:.A@3>20DB)T;!F$U(%IEE.)4C=(A.6PE'ZF,G.E^Q51DX8 ^0[?^H(KE?$;(Z
P/%F0+?)FX8/D@IN5Z6*/)-KJQJTNB%G=!1_SVWA7%Q,H(CQUKT*KP,[=(R$%F1$C
PCW8TX/&<OL27LB_5@0I^(4V)TJ_0RO"JMW*.BN097:(_T?8G%"EY8JQ129PYX_HT
P5PD0H\FCBWC02+MD1":OY'"I0YE$:.ZZ56#)XH8NQ%9*CC=_628<":W15Y;4_)]D
P'M645:?A'-4PN*@AM-2#"PT=V]<^Q1+;GQ&G#F&<3G<^WI+,.\"R\?":!ZG!2,69
PW)3%\@,BT>G&_:V3IL%9D=Q /Q-M-H^)1[6)!&#0Q]M[A3E2L,H*^+VS(UO/=?]+
P#"(I.T0&=7J--L71&[3(WCSQ_M$P&SZGNT,8 1=-!@8'ET#4'R^!WQ:F;F3;-4-X
PGX"Y7F*GH>(%D*U19A)W2+_1%/#Z]<Z,DB+'/-JB_-7"^#6M(EB'&X0X6\@\E,@2
PIORJ$2"Z@!NRKY'!YWW*YN@.6%,)O2S&CG_;8$@ZT)3#_Y/O:OHXQ8DN&$N[C01E
P<_EZ_R#AO:?1S+^$_GPCRM?I)&_&N*]D./1RU6A*TD5$#KKO)%"GYA[&3/6!BSO;
P!C?$X-97^;C".N_&/ =03C7CLT4JSIZ<E8BACO$W [C7D]%^^D"%ZHA .&/D#0)R
P -H65Z51!E%^17Y_:/+*RV)C4?,(($W%$VKJ'B^/T 18C?@/O\RC2A57M#'66D&H
P&JTF>BU\]5L=GTT_NE\\5L,D9.//F /0UB(>[<D'&D7V6Y8,*OGTVYGQSV2WS:6[
P^O=+ H*QI27'<L)B2PVI,U[.9TCF01PN@>IVH>PY"F&47050Q^9N@9)]N#O5^9+A
P6!Y5NO@_UH?U.3%4"JYJMN]0NK&VDF*3C*M=K6:QE% >+A4-XDOQ)%"GZ_B[!7$#
P?>B40/H.[0_VL3P?2YY>XY?0=IA6=* K!XQ*6D2)4S."B=/D:*H8HO[(U<8>G5M_
P<RP5GT&O6]-P_K[#0+P#..<X1_8^/.CP28;6+)'BN/M:)[:,70Q_A^S9U2TG<-A2
P;L1<@JJ"?6=H!"[NS=K"F[_LH54-Y";GQH^4:SF%%0Q'7@Q9<Z70BO%A$S"RH"ZC
P8<)#][TR664Z=7<1,V=<?T,M_7M)PO,S0:5Q!RV&<\9:#1NM)_4I@3YAPF1QWQCD
P.@14OE!7!50ITK>Y:NW, 'H0;X!6R02^"8@FSNBB"4$+<T3M:FE3:.I(;'LLF*@"
P_C(B<NC61L:;.MA*$.(CU,ZDWX"A1U;B,KEUYL(?!YYX:S9D'/S5_\*6&&(1(BU?
P"[\]]HSQWA;LHJM?>+?P9Y-+9EFH>G&O$^+O!%I7=.M;7AXULW&$[#)XXV<5;G3L
PJ4.4- Q(262TU^G9?%D47WERS*3Q\B#-EFC9:#M+WX8H;7VIQXVAW\QU"]>>0DHL
P7BRV=L32K<9)W]&^H:N[+(QT)AZ><]SK,7C-1)>/7KOP)!!OW&L.!]P-84)2=&R3
P/F']F6P)@7ZB&9Q)0M5Z%:OU/B\P@*OL2G.-US5KM!JN+]-A]"3<US-9J@&29[JI
PT-]%RK C7:O7:.3FZ+@#2^/!DQH6^$(>+!VG$L4_E%)\ *G<6B5<F;4-DN24T>8\
P8<2'YC4^;?%H\1KM8W,Z(*PO^OY_P?H^1$%PR\&01X!5_5'LF'H]W9YHL6"M!>C?
PI>=R1&'E7?4^L2;D=PUV(%'1AE(S\GRJ5_,%DC%6W?_H^5].) #U?=F%XE^NQ25!
PP+@MGO:/1*C(3U--1<C&_.; T'/VX(I>J\_C!NAL2!Q.XK6E%X"L^X7P]]Z4\&KJ
P41 %JU04FNZV8I_*GY'-^1"'] U7A3E@HX"S?HO%)#P?,0![2Q:Q[3X![OS $U?4
PNN[I8C*P%"P21K?R= U9OZ!/<5WC#::3Y5]QM+.57M_9B(VYG*%_M"DU\$[+F?E,
P)*NG+UW03R 8HQS]J[(K5OW/G-I'FVR9*I6N=_PU5.K]-U<9-S$H>"1^P2<^!@$V
P#=/E6V?;W-WOY8HC?C+B3+E!4 E'M55H=(0NE$*8"9-FBWNPM;C)]@O;^Z)FMZZ%
P\R&,YNWJJ/R=6A4%^;S631=,?"KP>?X+9QD9=33T?6@L69#/4<4YVI<&^<5M5NC2
PFB@W]H,*VV<Z=/M1WFU7X.JO&5_C<W.8@[Y1@V[EB,+U;&LM;TGK:1J$_11(4Q,%
PB. C8S&7G'U<OLG^CB.<&:LKL71FGX<^4DZM&@HS1JDUZ@YB0F9!T2'(WR"@#CW(
P.YKE>LOG]QP2]PKPUBR,Q]VY[$=BZ;(ESJ$Y_"KRC9>*)&6<;JC.[2!=+1U>H6 1
P>;+0K^H<.PF<6K3@N[=0EE#:@SIA\.4\6,X\A>ESZE'RZ!47QSIDJEH^EYI%F6MY
P2B$2(CU%IRM9_]YE%:_;V;60BO&A(UK)1239 B8(TJIY :X ^E>#$F6LAY])B[&K
PUXNQMY@?,V@4+E\B 6ZU#CSOLN*;@RG:/>U?,PXW.:,!<^3(SC,$R.VQF;3JKMGR
P_I93JY)!Y\[*O]#\#I6/7/OVA)=S.E@N3NX-\7RN;9EU/IO'!3*[?J1S:#%6<^$X
PB*9G)&.-6B5+MDFNN5WLJ789KQ;<SP *:!$U31W&+:4I3=_O:4P($X_30R59/MVZ
PC'EWB0CT_*6;XZF OQ6O"!\P$2S"L1I'BV+JX ;-Q*$$ATK0*PU4T]FQ?T1;<%KN
PUQQLHB]*&ZC!P^[_-..-I%GF]'=,@W7TG=G'3Q8([2)1R4_7'^8'BNV<9>,_?&=Q
PD=?H"D6:X44M6 9;7>&YQ!A)+..Z.V S2"Q]Q\MM&EDTRRGG[I&<9H^C<Q._- J7
PJ5T\U/A#UXSNQ2#E7*BH@WIQD@0;:*\"1\[^$&+(P.JA;6&(D%E0B!MT&J!-5V2+
P'MI)[1O5"5''F&TZ_MS/44B@DCG#I"^QB^*J!#"X,<: WG)(5 <B;:KBUWJ(/ ]0
P>*W8QQ%2JI.88U5%M*!1N\?+RRZ8ST9IA.7^N$RZ]%$^<H#SJJV6J/3 ,V&-CT#C
P7;L<*N8$M785:=7)S.F3HYJ1-WE5\@H"VLU[OS,B)O'ON-&)1:'<FGL298&_@CT3
P/ZH4 1-VU]#<,>L#.Z9&*3WH>NSHF8[R3AN.>'X<W<A;UWCX'6*K1 9:$!)W43FT
P-G:I:E= <]$77?[82SQERL@+HAH:X?+REJ2<K5GSER9AM8;+[PHL??3BZ9"8O.V6
PUWW?RW)FJ'-G9%7[.5S?[ 80A;O_LB7*P+5Z$K-<%-+JO\$]KC'/@7L,.)LUU=?5
P>C@^Y3)2BW4B"YJ<[VV?#U'18EVK89!M8.I/LH>VP$QVO>5W>!)7T55&.LRC500T
P;!FMUT0S^VVS['YOP#I_W!U_LH\;'ZY5]&3RG@S)W-6N4*\GKX&)P?ATAR;")NA+
P<E^.=OS"H]I,KN:9MW=C@0RI5,[9SW-4E4W8 7\H%WOC->^'-9DUM-(::G1/VO%,
PJ P:@0* G#[C?(TPG$R<ENKXW7ZUO>H1&M=,@,-CO2<GQ?EHN$FUYS<,4[>K"A\H
PG8Y!:#[A3L QK0&#HCKBT!F&B@>H[G0!()7S<I[SI.']2"@:N%:-!?4MI]S,S^\:
POZ>!S\N/C'JAP\PVO;$0Q^H*C6TK##Y6JL4T<GX%D.%!J4D03?B.G48S^.Q1N%V7
PIVM Y.D"![,N-[=%C?S&N:D1V)B>",'*!JP.C9L(\6'$='DEW$T$\&63BV?CQS?H
P??TVZ;F]+S%1RXEUHOQ8,^RA-W_->?Z#5)H?E$&3P22\[^/_C6&%.^Z?0.3\BG_%
P;J6SDI?ME7POT%%8O<>@ FB184N#QS:[CMT+N;MC(5X/)/G2;_?\<[$>!!7M&^]2
P?$_)@D:]-S)"W@2LJP1PZ&%=%X;(!D$LQS(61]<N]Y4JC0,>)Q.A)YO;.]N2\,*5
PNJ6*JS:+*5@- /B(\1\_DP?G I#LH(IU,Y.F!H^*YCJ:AK/5!6QP'19[&RE2R*BA
PJ@A#J"+2])'5_X)N]SCT&^>S_DX^NL1?%*:A4'7Q5V#_O5D\2M*6]WY4X0QR6]Y/
PXHL>V;&OP>L@!8.H72^<L 62[P?!5<N#7"/(BW=<P41;-L=6KE,O(N$&HH5_//PN
P0UGG\ERC'>]\I^CD-5M+@D.[V;(:SSY9JKB4_O7#L((Y$/?_W]&CMZZ*$71 ^],X
PH(\"#J0M!RR1\=5\D*T=X6=,,39&'WFAJNT (II]SMM!K9*>L5!;]N^%(1+\Z 6@
P$7K-MHH*0GRISP(@X\M-KE"BL$;G3:O,*ZV??J%(UYZ>B?"HTK=YH^L1TY_!/C\A
P*+<2;)N%J7#B5(^5D;N?S&)W@ZY.Y1,IQ\VF01/[[F=0M834U5K(I"'9O_-I3DEV
P0Z?RQNN++2^7NSW#&<QX_1Q8(GWNPXL;8T@A2X F:B,+9?F^<^LIN5DS=P%7^E3F
P;?V)I<A.PTHJX0G(Q ^I-/'#+_WRX;ZIF=AS/2TW4QMFYF[.NCM[G,:?4J<1H;5 
PF? SQ)I6$8N=O/6?#D^+?0%ZPJ6;=G"M<'>R!BL/5-Z.7,-%"9/'0?L&%7]_(QJC
PXGO*RND&(=<O3!/.6J(0IMIU/;+A,JP?A>^F.Y_#S<>C)WALS=2N[)=S$M99;501
P;UY57#4]=:4$>ZXAN;'@8,DQ7@@RP.K"-.Q-=IKFFE=Y.-MJ@N#ISN[PK(YGMZ^^
PX<<5FME@V.%/08U+[;&AV0)YBP06^YXA <BO$M?MT[L)=S_$GWZSUZ/T>X1BOO8B
P6-<</Q734KZ=^-D.J)-&;K+M;3:[K9M"B[[.^UU@)=:CQJ;!:-S$,2 SV60B*1E1
PY(3MEPSZ/6:GSL666P0B_"X;15X_*?EH%]G'&?MQH1)AP;F>X3#P!!ZFU:JV(R^N
P::Z@VYJ%:.7&NC6_G8\J6R-#,-:#*4@VLSK<"0P(IH2Q0U9W.5D:?&H#V4"HFH8]
P%8_X)Z>$\U<B4^1;XQ5[5;HRE3G_R4 -!6G'=Y@I6P5("J9VOR/;G$%<6$D3N:T>
PXIF2:K2@)K+X0,Z1LP.Q F B5&XRA<;%:W(WLD;&"Y-,[^]/4S'CD,E.[*BLG)^+
P 5R,DRKX6Y3B1Z)Q^WA9@7F^\J7Y?F!A=GM&QW_H/EFG#+,HH/JE)?XXF[S4B&O&
P12)A%WX5GL8&M*F7>M+E@&-J-)RT%;6>4-[/J@P<ST95?+/564P:65R2S-8\?XD-
P/;JUSK"OC3LD:^47?"8??>?$U._CA&$CTD<NWMN"8MC("RBF*#WBV=JD-[3T#&##
PN!+"*<)9OYVW54_R%V+*&)30$%>FHO3_%ZI?+HS,*6NR[]'<;RZ#ER<2.E8Z@-HJ
P1G:'66_^8NPRUE$Z /)@_^+_V6RXAK?%"-S@?QRI2[*%Q$#.>!;/2#)5L<8XE PP
PK[>5LIA4(W JUJ1 :*M%M$F4'!2.(PW<3GB (_WXKH?$(RP][2#7(.'X'"YRKZ;M
P%OX5;J')/KEQ*9(A"H;_@3!/<EU7&=]M;#R6#BS^!">^:]ZG#4.B.C5L<FQ:-\X@
P4NRYV<^*IVP-@7%NUZ9N:!+%D_?!SW-!5D[K=$T!O5,,IY@35=4:-<1=;J%9>ZUM
P]WLT43 %)! 2Y"P:^G0]Z]]&Y_-#T/?8D9H&M)@2;MY&'O<_(^5/$PJHKV-%WI,*
P@9)!>@2%72=PI9>L."WV[@5_HC4_6-.A+%+0D^\;X:6&@$GR(Y5\]8[2*:^U'TSP
P'8AT&&N;E0SQUZ!AY7#0(A!8-Z*8?L*7*<-A6F.09"K<DZWUDP (8 IBBNZIC/3;
P484BPFTY9HO"0/]<*]GB:^>VDOF0(QXG!'Y-@:)!</6>23#J?B_G%D8 9P':T,2^
PA=!1 $&+#VZK.F'K_V^CB8%QRKW;*&Q)+A$I!;8,2M8DQ77_, K6GOA^P.\?47=P
PCF&&F(6!9T?F'',(9$2MGF*QU(&9Y2]%=RH'\Q@/=C$3(]6T8X89-^BT]1V4=3[;
PUC-5B1H:DZ&^Q=/2OYV2O/I5G?<)B]0: G$=%7<+-4CN22$'Y8  :N%Y9OJ;ACN=
P+*]=1_3WJ\87YC4+%,<+*50S 9]T0@?*HLU'/!,Y_5:L/<HGO:B25%V%J1;D3>_Y
P;]Y*US_,+/Z2+,&SH#1L-O^EW(&J%HLE%="C?(=( #\,,G6W!*C2?_!GP\R$==YF
P48&$D&0$6AME5@9$4878X';*$5JO"1!C]U&_J%TUJ8)X?4IZ6&LMC/6_8>$V),=B
PPV[GR%M78 [BJ0J/)/_D5F4XS(9<1$V/ (]>!,O!:74!Y)8%9Z2F8*0V?SPIX"DD
P'FUZT)9["=W\BX -;'1E\K%C_\I:<]964>0!(>;5F'^;D-AAAYFW+Q.M2F.3(MQ/
P?9V1#[IE_S(B %2ER;0#;*]- H6C*)3/92?A6XX_KXJG62FJ("]36RYJ?;?Y+Q"U
PQDU[#/%8'4CS9M (&%#8FGL@ ;?/!-*7$-M3R;7..U-17_Y59,**K98(AZJ%"V,2
P7.<6 KV.F#C/_>)!$R+6E'(]566:0OOIS\,W%< E\+50@>W+Q!'G,&3E*#& /-M,
P4T2GTM'3DMO^0!?K17Q6^A1.8NWD0K.03Q6#A$T_R*R%.[8Q$X)BG"Q[M972\ ^9
PZ6LFD65Z9+/?64AI/RS\!3WH'%#R';*^P>R<.R09AB9UWCDQ1'"4]")CP?5+K(9G
P?<IG:<:CU=AH4*NJS.4 HJ7 723=W10^\3)8^3$H?\]29%(D/R]WOC'& 6'1?\[Q
P_I8G(=KG,4>2TYZ UKD2USF*;@$/ZLG?%>9'V;UMX?99(-HF<3WM,6-N,5!:>W#,
P]O!DZ'.C*TEL VT:8FR^-+XT/UOBG_"XOYQ3[;=0VEP3&NCQ^'[SM"X]<H5 X34*
PCF,^SSSH%K*4*:Z3ZB5REY)2]X7PE:!JT%QNV-.J>]Q58W.9+0_J9 O)\_>A.A$Z
P"O^;&9(%7Y1Z7H1T)8J5P=UB:"0;A;S@C]]-#&?/6+OQ2I[V<0('*\9>=9MJBN@-
P'(1N<P$Q / '_%Q=+EA." 1W[CIFMM%QH[\";BC.;YH9$V,\F^IL""8-TCXO5@3=
P(VJ<:JPRI;BB8P6.6$O&V1)#I/_IZZQ.0/2@]BNF3EOCMD!,!]ZH:DCYJ$Y-Z7P)
P;INZ+H1*.GJLQJ L2=&@I;W2W.F[D/,F[+L[2)1>PEW9?Q5GR-_;QI\NU G*]$G$
PX=7M=*B(9A7AB+M8ZUUM9-+L.%J_^ 8QRD".+76I)2JL!W$FZ$9H04;YE0'J0^&;
PU]6RATW%8(4R4L\-V*0J:+H".HFZG.Q+& HUSUK.0:?1U*O7PX"J23':!'R' B3M
PT7YPB)J?7<__!$D(Z,[4M0UJ-_KYF]C&.N66>N9*-;S$HSJ!-$BHE3#D4C0I8?Y=
PN;T"D&)#:(F489U*VG7_ \(X.;W!TVR*R3#+EGPMF41CZBD(B%WC??BN5#?S =T1
PM-ZAB;+IOPX4@93>4+OX4D63Y9X2L;-C&4'*<9[^[M2AM5.5*V%K5UBOJ81W!Q>>
PE]FXV1H<=*G%9;:IO#ZB3N;@[;_X>8)KE8ARBHH;YCRT#)0KH*'=L6_=C/4_([65
P@5>ECT$F:RI(&UGFA_$@1@W)1>RQO^RH'-14SV\0=O,/Z?"UKK%V39F?6"FR\/CV
P231FFVTJ[L12[XQ[1BUSH@F6Q<EWN&!"UU_Z:%:3_[L]U)$E]?_9C00 M9_\ZY0U
P\83VXN[@V<K'Z&T)AX9?]GAZ 5R+9!E!KJFL4?&[_C'?Q!%E#1FKS@N)FC;TYU^1
P+T;I<MO!RHX-\/Z)4NXT;-.//;VESAQ3!%/@(T9PL^,P$QK+^1SQQJSU0::]7(/V
P@B4,HA)X>^?&1#(W\  =>%H2KPK#<XG%LD/($=0"AU&VI>Y-<ZMY3VUD^:@$3]1#
PE5.UIM*'^(*J\0&;[;=.- !E"W2)FU4GL7<R7<KS$(\ A!'<C!;IHK%/*>"0B!XC
PC+H>DX;=:S>"W;7V 4GNH?R NAMON2(H+).@V+%Y7@,"<<?C=!$8@;F4 WD:!E,D
P%S_JJ OW)R* O !WUW\UTC^3T3=O\5!,S(H:J1)T0^S0*CM!\M1K+T@6!B]@>&,C
P19<?T*:@3^]O2P?*9]2R\.XC5HP#3L,@$Y)J2YVT#7Z+/.F@1FN$A.'RD&)YO1>W
P@B%5^,5H1ZM)@[U)/=KOF=47Y=N;]BR]L/8@B*".PATBNO?@]J^X/FVK,-'/9,EA
P N@UG"(COY/?Z0[_(]MFDW-P+"/W!@K&!6CBT P8EOZXAH-IHU\O6#!MD3N>7DKF
PXT9.\KK?)6V:(.6+@ ;6YOERUV$;NX"[8C1:P-L8\V,N#A*08M1FHUVL^-,M7:/Y
PO7[JL;4331-AIWTV)%9P0<9P?@'<;J=T;N?A%Y+(1,V\7,RU(R6JYC;<SUB@28< 
PH:<F(T'=3W_Z)Q3IZG@=!J:Z<1S6K\'E1SHD8#]120;F/I,W'4V"P;GAQ_:&<:#8
P#*\BE\8&.W4HL^2%F[GJDC1FW(78'&LW9;/E,,[ X-'R:"N"& 1!"_!;$Q6WXBM_
P#%^A*><JA<\>6II6JBZ;QR*_$F<DV@3"KTK"%02"D30)8;^%MSPA54D42BEN[ONZ
POJ$D_3 8(,\)1&_K'-<L%YC#V_)196OG&B(:6)E9F5>7!^0:OIV.O'F9=)F5,@_6
P:8B7,;YH[6#LLZ5W+ Y%O@(RB"A4@[N]HA^Y% ZR18RCI&9&?%FX>?CI0(BZ&^#?
P3<=?>T=)9<K) @X!**Y\E9@X&<QO!\M1$Q9M?HD.0/RV.6 V1WJX407'5-374^QZ
PU^,X/%Y,G$F!>ZL>[F:DJ=IK7RZQS/3$<<HMM3$Z[K8@KKY^5HPZ.F&-D/"PX^]Z
P"!@:P(P0&I7M# N8Z62?,?59YZ:A#I3] G, >^ >N%87B-O_]RM<K TH?'RD&;12
P";N16&>32*_H)$!%*=PH6G?^[@_)4/:CFW%[+X<V'-TA'!?Y1,:K^]RK7K)UG3IM
POY&_YIL,YN53,E 29I?+/VW6>EKI,[L(LTR 77N3K2/:>4UV=8=Y H+5CUI)&K2R
PYO=7[B6'.&FRB 0+#&ZH,JJT9_^EF[:.8A2]91HNX>T^^.OA688:4M\L!%WNT^P'
PD,',#[V<+2=@%W#97>.*M*S4;/F)M0\Z#V907QBBO!"\QZG(B)7H34VI8CLHG3V%
P8IH]I^R=E39ND]EBFRA49QT2Q:6\QD%BRRB0L=]%Q8;:8%"?T SW0QSESZA*;X,Z
PR0%ZEE=*EWNFOY7/F*[FBNVZ,F$AO].+_SKB"1!W#3.PO503]G0/G=^V=4>KXC^O
PXNF_)V"(_S;OC9C97P&VH\3ADF9(VKNCK*B]0KAD@Z[1TG^;9016J3Q/3>)HS*PI
PG?0JYHS 'LE34T<CI $O<1)D;Z8%STEQQR &RR&&K*YR_1..CZQ@B#F2^C%"X27Q
P!G;\9HOHJ(W4T"UB@)\CWV=%=#]45;=^'K*/_*-@6MQXCYO>N@K.-L!LMT[*.S:0
PU'0[G'7.0 @%RMJ+WAZFP$I@SHDU+D#S,]6%4>-?GV)$H5Y>*EJ+@<?5I\PM*PD5
P?;E4CCXV'I6P<T\)[>3& 9UJ.'<K>Q<[@%W0=^L9N ;#G$6[0'P#=BZ@)S"0I&NK
P?Z-&W,ETL^49Y*0_OY0W^;W3BC)>VP8K7UFMZUE#\ +A*5O!1Z;4DD*+G%U.4[NQ
P'>IZWA+3_S[O^VM)<EN\7 %X^GR$=L^4Q%JA!?:(JDF3N<OP<=1[M%]UXZO,S*ZZ
P^T@Y[?R8L2<^#)RU^<5C3W'8+R*,X ]5VM7N *GL0'+ E=>QK/@?9\".61IJ#R9W
PLF])]!W>G8W,Q1..Q=)X+=U"$J)WR9'#84< KNN!N6*ABD@].X\MN4(27,X=P-!+
P(MM VJ.2>IV"HK0NFT$[1V!QL6A/,I\SVB:D_J19(QA!)FG8?\(]?",X@=H+L&PX
P,+ASZKIM;:)3"T4<G3X-C7M)&:T3R)\5!!8ABW*58NR_,<\_M;E%+"9?I,,7N;./
P5;_MT2*HSXZ6R(N@T+PIJ*GE4M )5ZLF(Q3Y/G4')D2;2YS%+J#'P]7$YU99VJIO
PV(RRM.L(0AD0KBV3VA.SI3E]&K@9<SECX&$N/+K(H4FATR7,B_2)>T)]N/;4$[P7
P-+DP+'$'8^(Q;!)#=ZOEQFTN"EXRN_NM66V!A@U3_IOWJDV]_YJW)^).,K' "PI)
P8MW':K;/6+_>-ZC90__$#>I1Q%*WHO.*7UC#".'?PAV_&]F1_LHXJ)2T<*KMPY'6
P^-AM45R;SQ?]U'SW/!'-YS(I61#B"  "+7%Z*49= /^CGHGU[P"K^R*9VL"(Q!\D
P$JCRE1;:FOZD,F.YS4IH?6ADRULB=XD(+'_%PC5G>.!7%G9%+<?;',9L#?_NF9@B
P((V[UU%,STC?<Q4$-PU0Y'EQ^1G?A)@.U9M7!TZ3-FVGF'1A&O:3KCF %<\%8&/7
P7"OFQ!6&>T2,:#G[2.0ML>'2AX:WC<K_/W6'^F\@5RT3I;$@M)T37E1S$#SZO&*I
P)!A(B*^]Q;/3:<T*%Q71U&/@5N&Q=*])=N3Y/ ]C!A#"GYT/'QYQ\-9>A)3=H,4Z
PKOX,LD:7*W!=(^.GPHCZI9F(HP'E2,<&28VK52<8YM?%NJ:]RF'_%J3=GMS0F-ZI
P0=-VP'?+J=,?DOH4PX$Y%':+PS",$D!^@Y:WDQV^@Z91@^I!\/JPH>\N.%2X9BZ@
PDTT2 ";ZBU% 2<?O'Y\L]QJS>+LAFB>?POJ2WFDHV%::>@.==]$>:;9*?8"^(\M#
PB ]K^.0)BGQ Y41-Z1#M]&M31@FYUSSSWZX.]^V&@S96(VA'7RP%-19,R"/]ZO?=
P<3MIX,G_]42@*8 N:#$)I/0,LSIA S?UYVG4492J".P<0\IE!++[$?S=ADO84C??
P&5.II*R[ZXLRP!J.%A?@U\<?S$O-I0D6J\#:I1OMQ-YJ81XYI.3]^( 9VCZF B'P
PH^W$\"PL!UR4<23G+-6->8M(#YQ8I"]DPOOYS6II0.OPYW"]H1%X&#3619K\:R$<
P<>@=^*6Q#O SMN%OX:Y_INML!FJ)H,"&YR2U,@"'D:DOMVAPA )Q,&E*X>UW7'W^
P2$I"S P/\\:W>UIM@9C3U^\/]Y%"9 17;=_$).$F>K5"?'-LG3@<%/.]\4AZESHJ
P"3QWS7MG[==57P<16;)?HV_H\Z&"KP%PHOV:,6TKTWBR,U-&'\F@V>)MO38$:BM,
P-[,_RFO\Z@?UB^]I 2UAG="?C8Z8I]59@JIS*0=,3"##-[F<_PE%6?X=X?:VU!2S
PD:.3DS(HONL3KY9&K\,*\ D1"#)[GZ7#,8$#H>[V0*QAZRA&8TDLV[B0[%AE5&C2
PXQ]+,P?VD$F"#&UP>K<Y0;T!U&'/T\7-SE<#DWF)'HF[)KJ@(&:.R\_Q$99$:8G.
P86!0"0FIB(A615T4?1NW3"L!:*#@HLU&!L=3'W4\=5\^J':Y4(!&^*.#1R\?-=O5
PXO?!)K8^5'T]@+'J>PM4'N-RC2*:T1:,4,GO7N7HR91^\)YE=K2Y0\-[CWH:&@M0
PG.@@VK">ATWJG<<CS5'5R1AQ0G 2)>*Q\>%B!/*[#;LVK6"OMUZ_IU6) 9YIWR9\
PI1W2CM3*(ODIW2W&QEE+*'O'3IE%:JZG,:O9C*U8D_XU_KB<%UM@TH*S'*#?6AJB
P71S+C?%FG8E-/O-E@M$O9_ /FN3V><2 QL5J+R_OUIVS$C":I:-X9,.?>\PA6O:T
P75K\^@13Z'W2-/6HFK1R7>J:1"KY(;&]ZH*YJ_AL@^_H6'2X;2&&4,7.?\D86VQ4
P +JD04@EI47]1N="<R7D3OC5M&U]=S"SUT!@^Q1T37"8^:R!>[]<5.Z:M\3>7KJR
PO6!N )C+R=4Y<7<O8X?N6UX%$@XQ&=#0*?'67;V265CKBGRBC0-'IM (M\R?JM"X
P)_2<NL=5B/>*IL]=#+Z[OK]6\N^7 XFZ/5PFP@0!,=,EH L_1)W,^D ^6;A$_PA,
P0'!?&76>I&#%X6 QQ4LX%3&CZQN, CO;_\=P8"!^]\-V%]R]QE=;@!9I_1$LBKL%
PB0K=1%]BS!CB&-@&9O%ZG)!?C#H7*DP>X"1S+1 'RB;<)I8OEJ@.I*:OG/4$C&$>
P(VY-68VF(1^_$MI]&E"+O1HEEU0UU$>FSI4 XA,795"'+L.@GK+;!TVG:PMRKOD4
PD+TK>1*5]Y1K*,5/P7S/IF9NW)5XI2@'AIH3U0D91Q_BG+6MU#SC01]TQGN=EXW<
P3DD6QOJ.,B-3EPF=H=ATMFFS8 MISNP,D+24ZZ4RU@Z\3Q#FO1ZO*DRO"4Y""<"[
PK!P9X;"4"IFK@I3*ON=,:@V(HG9^<4HZBQSVOIB6\^:=Q(CI84<(E%*3K<\RAM,X
P:U_! 6R"_':ZO1&G^Z)1S:8SX<N,@\Z4HMR,$B -UB?6+NG-8]AN3(0;V2K(U!/"
PUNH[UY@T&ROE7(UYN+F,C^;=.$F7U!.=S;:0;#&X]K:",T20DME4PAB2N<W'<ESS
P3WKK>F8W9K#))= :5B"]UX#=-C4BU*-\%*V+-;-C%QBY3Z1$A?C*?D;!", GA+FG
PFWNV!;Z;Y91K9"@!*32]-!NGN2FP!ET)/B772B&9FJ3CZ$N4E]T43NN?'Y69MPA%
P+W".>HRW#=@5_TH0FG8^10OY*GY.F-RSZLGIGW4+>C6<DG<S,$^&%:]3@*S-E#O2
P"5YTL\V5)S RF(P1X;@9M#^T1#*/+,XXX@O)>=;*>W$%8IC0/;MDGG%&A.)[X ?Q
PT:IM73,2':12Y]/Q"PI4]YWEB0^77E"4)"40C%[LO>*Z^H9P  Q\+2[-DB+[95.\
PH^H<UG_!!X\@S #]A:A=Z'0.Q*)E]B\0(9&./J5WQRF4[&)1FI4MX(/\JD#' ^1"
P -[P&!G9HZ6WD,7/T[#5X)&SZ?_@\["JL;,0<NZ.XLYT&A]WH9[&?#KC?%YM7Z*L
PA/97G6BZA5:ZZB01&^;E>89GAE$AP:8@A:P(UUG0N'I;+TX7H2R=5NGO+N[XO9*D
P+87AJ'DQU]X$(U89OZ]!PMLRF2#\JK% %DR&KVXQF\.,-H($!B@D<KS&G->/EITE
PN]%-119D &$G=:Y5'_L,UJ<%0EJ#U%I:(QFP=$SS)0N>#1@KC/7I_%!;<'+0/K5W
PGH;7I9>.WKW(^KF-:Y6%.;4MP73:GPT74/T<Z5L40=^#N R$JIXRN&U7!\8$_AG5
P3M:_3Y"?L5VH92 M;FF0Y%$3#M_6'K%-<S#2P"GUZP<^??FJ P\L]JPZUBGKM[AI
P/.]H-8?"TU)\E,P#M^BZK*0@$.2C;3!V"^! +GI$9S%VC%A( T:=DJ_BD_73C^"B
PSCC4Y#%Y^!(!V_FB@S3HO3"DZ4IO>.8M&5;^(95#1L+>?GUER!DJ.[\OHFKT":6;
P4+D2#2#K]]-4V[N-(%58@>Q\JA?(#CV<>T^3ZJT)D%V<59P/5,3\P1#+4B6*"%!@
P0Z&611*22>"N48H:P$H\4,-2(GR^P?1@:WZ?^ \AE'-J @%GFJGZJ>>BOX#Q,&K/
PEL[B):<8@F4&<QZ%NWE']6XG"JHU@>R]OAZ +Z^ 3.*+7;9P.9@,64)5*>'6XH-O
P-1I"9>_"S. V>\D/, F4?<1T^K]O.EYG2@]$RTWF>F?Z;@""J;XI0%A/($IHZ,=@
PCZ@PL@WE!KI*;4PQ 1NA'M2.R^?,JA!46U^*?N%>\@2O[CH70QKR,IPC:\[S)K>A
P=C_(VH8WS.)&&U\&F_+D9S/Q^0!F[]LA-PX L@2?V]<%8VGWD]E%!*;YQ !6R*JT
PB68_KHL#DPQZ:[]R&6<--@\P,J 31(1>B.'N^4 &@%\&T<%G/5!ZMU^"B=$Q6WHU
PY^/ELA B!YE,U8HP?61/)NY6"*5!D'"MSP"O=NI)C8\(,7YGM'N=C L4VWF51 [V
P>>Z2P#3[OMJVNZL1ZVIB3/3<_ZPC*XU!5O"'Z9QP(D1ADL5K>T$3[7@NM+F%Z C#
PP\C[-+.14 ^S[B[90^48F'GA3W[&_F(?R"MDXDBUP)_GVP_G1HE?IGP(@UD2UN=2
PFU@_8W]W[6YPA&K64J.VJKV668+,*\H8B-_F&'T>+O0F(N!293NIOTJ.F6E8D^:L
PM3@-4"ZI=V0/Z_W>!V7"MC>6M44YO35/JRNFD]+.X-,DUO<LWD^<(?K($N^>]84Z
P%HP847^%>4HIY"EG.(RTY"65UDYPZ#=3DK#*GEF7)HQ%P6*C>9X[==?=KBN1DJ,<
P>%'M0WH>F8[A;>\:NI&11W:KIZ+,SCP:D(O5#IQ)Z)&/B2HEU,U:G^IW%3.Z?MMM
PJ_-P5F"R!&QQ"WH[+!'P:_-,FT=\&]$EVLZE[XGUZ),%(S.[.)3%8,FFZYX*2>KM
PV':!'/;1JVM9:[,E!RANMW%FK,D4*-2W-?<D>GEQTW+3W8__H@QTJ606:8F*DJ9!
P:OHX(@\$O0Z=DKS3U?,."F2EP@<:GM<P\6O/K+FOCWTX#C?:T%#')5?SXJRSDI/[
P>S&*.!\* OIZL-"UC)!;BK09R^7V[6*%HW#M/?G:UI[+$LQN&%B\FS($E*/AW7ZX
`endprotected128

////////////////////////////////////////////////////////////////////////////////////////////////////////////


`protected128
P?+)9#"+V.E$ANY.BG)2PC,U'S:"!PR:&P@-%,4ORO>KE-_ER#,[G>X 5&#C5I#RB
P<U&'.)_0]K&.#XQU=.-A)O<:@:9#+M^8=543I+<'AVXTH)(F("VI/_HQ?-#)-Q_:
P4$6118A,H'X>*!"A<,G4&4/'#H))R;QOV<)EP2]IUXJ5],33WKX#U;>.'?4VL;:V
P^V/SDH/UGC?=FD53'*&%H5;>Y]TY.KX(U.83ZB@PX-0* N.#370" B36U-SXEC=>
P9M\3+D"HL.@N3W1G6*J7D(W^Q!* --!8!( T[CTT:/AW)XK_S![&Y_:@'IWL.O_#
P0V5(S_E7S27>VO_<=>? [JQH,,#LK]>7)@1S1-D47J@/MVXM+5Z'%Z&U(@.(#@JK
P+/F-(NB]&K -1O2:__8$_VQ3=+1(Y\>&2C9."SPO GKS':A"#"27+C+];(64:<)S
P/.$[T-ID!/>.K7C]8DL^R5S_OU2\+<[Q@49"7RRSD(/*I$F;K+35NOB%C)-T3@+_
PNV:.B[6(  + @R5S*/YJ0=SRU"\657M_H??43]GIYW5_QM)J(N/5ET%4)':Y4RWP
PJFSLW>OJ_=-4=AE'6)_RF\\@;>@<Q&V17=)EO$^\8PY/,9!T0-Z%DH.WUCM"^$<F
PB%BIM\?JN*3OZ'1C4I$+-:ON-[HT3!#CT2?EI'0Y=R(K"[7TBR[->5##WINRJ^B;
PCI?Q;X1ZTD@;0"CLBV7M6Z]HOQ"A]Y5%V04YB@:7%NH%>]5&HFQ2,>!3^8!F8>H9
P0?^X\5_./9>HG]3HY(-MW%U_M=9J&C4#GH$\([P3+F* ;C9U(Y>9"UPG-]?E 'E,
P43V--2Y]6\]9J]KSU_"2&"F!C+L([<W %\GPAY]P*ED#70#I%EX,6L=Y;OJN^YX,
PZISE+U7EBBP2GFM0V/O:;>VDCYO4K5I15><6U+<8RF=#TPC^41+(7GU1M^*\2>7N
P93[NDK?2L9_Y/3)([!F<VEZ%;7+C5=OC86 ."^)R<U*FHG6,X <;ZQ'NGHG1&GG\
PK6U>NC$N14ZO-K$ X9S8=2A3Y@J1]R$MC[W_E4[58:Q%8JZ7AWL%YE$"&@76V[7_
P1O-21<4(N(SOW[#[SH'GIXV5LR.LES:09#E_$5N JCB9!U?LLHM++;)A<!/(PS:W
PX&L8FHW2_V]]0M%52PMOD$C!I5ZIBUX4#8W;=K H?UE/:2H4IKWGN_A88HC5P=_5
P9ZBRB6X_HR3+GHC_N6'ST"66M6>_'%TAC=?HP^NDN@1V=P>@)S5H]1L 1\=:B8H*
P%3_1PQ4!.SI$9O+!16XN85,)?-5XO*E;]4VN):2=Y*(_R13FLK!BQY)B)0WX87Y5
PD KCDY562V8CA %WL^[O2 ;XN*"%/.HO<%ECM0AU4&AF&7RSVH]LCQ(YUUCNLPX=
PT/26KBOI<3U@,MM40:B)ME0)'<MUX(F.3 5.>KJAE"[.:+SY$#$/WWIXIM&=U][3
P=<>NUF3JV<,!ZX2],=KH4"E/X:7N0T/F7\4(=(0)J).5]V@=*'3;5E:CTIB86/0H
PV'^GW-G\50/1EL4G'Q/?DU$QS'9DE6Y?!U.P4\C=N^H6]79@)%T['$C FN;&N), 
PB3$FVCG[&9!6S"6?F!9(JJN=8)%[E^;X<7/$O058ZSU'P[P44ANM9Q'.C'JK'F;%
PU5/$X\FGYOU\7J.8NA(UJC!C!7[(.7.FZ;QH\31Z0MW"&A_.#"@F1O$A0NRY>,X<
PLB9H"*?FVF8%5:U$,YJ<57K^!>DC)BJ"$TP9!1-_VT14Y=;,BA,X]S9($0]4I;0!
P[/3,2^JHXQV:A\XSWJW5P"?GFK1,'!_5NJ'X/9PVX&J.JXW(;]?MY3+M2Q?%(TR>
PCJXC(*/FO*F8@'$#=3LV;/<S$?%E"%Z:Z2M'(A':!EGR(%_OU+>Z.Q\&%O1I7$\8
P3PR2J/47!"F8VXP24"\3A!E/\WHN;2,REOX4UY9<EN?OP@!8:!P2O/K"C' *ZL$K
PG?LACL^:!2R_4H5C/W3 AR17-R]]]<DA/$^WI&9W41K*"O $Q(?X$PNK6YQLSN!L
PPNVJ^"UU"V#J/ ?WDZ[41MY(8AM+!!UTBMJ(?AP:H2!7Y1)RZ;AG2DU>Y)%WCRDK
PJ*,1G6(H$,HA8[D>=GX&"X?W5.H;O:FU6=(=ZYM&85$YN%$@+WB'>G*L=G#% Q/U
PF#*R6.BE"Z8W(7R.+B62P+^&@Y@V?C 6ZV0$"Z I@(YA]H?J:YB*6UDMKC:%$KIJ
PS31]H>U(['>TK8A\@.V]0S&:R5I]LGI8CL!)QL@&BQ+AHY5<%N->TPJS7F@(UL8R
P0M7H*UKMU@G0S$[;RVE+75;I&6>4G+:C_&)H7R8PD1%'Z8"=2Z(KKA-0:)@@JA4 
P1J!FNTF144R[+86*S6X^W("NC+.A0L M$9+3E=5WWN]7QI+C)%,\DD_[TK*VDD/3
P,D$*J! 5:%S\#6'EEPPB(;&=M6_</+.PB>*N38G4OV!+B/7==A=#2>U9B#$31C-7
PTTP4XXKN7&#Z]#=PTOD7]8E\SV*XHQ8L"J3,7QC4[ZI%'Q!!(3UU',OQG5R_W2/!
P6=M;=M3LW$FS;H'U(H&RC/@1HQF8QZ:!W[@+*.&+^[8*K;H,6,=BZBFW5L)\VSTP
P08A6JCQS6EYBE]=#D"NI@S5:9J[?RX1V=^E((51ZV*0WYD\X_WE92F2PT,LF(5=*
PVV1R+#\]R'BC(%=.)WHFM:3,;+OG;2>#'!<FR4Y3LO/JS'_9+:NELK@Q9#M9>]2=
P,BB#C4%V\WWJ;K0L@*^Z<*SV@NY; /I,M.R^SG"!\PQ6%%JBH'&36).D#]8S#I>#
P*]@F]:[-_EB5[)2^ \CNH>2\"M+'HZI32=(PM7K& 7P5V#_UFY!@24[?_:Q^,%10
P?@.A!;FMG%-,*FQOMH>BBLZI>P'=.1XJF%?*"RJ^A!:J3CA9X5_:#:YDF[[Z?8-7
P59S4IHX^A)JEKQF8 %.9 1?ZO-# G)]IPU:,B-4T>DTFP?;;<!=PXPE\%4[.VWZO
PA^%SFX;C1^<U#,IWHFLE?<6NY;.?]FS.R2KV_+R#SK^RCFHD^WW?4#E'X!U"&BRG
P$%06<CX3/.=R?PA?HCL#]^FMSZ%YJT:OD3LQ@;]QA'\CX:BX$Q)#FV*ZTFB%B'<$
P(3-H"L0/K@VLL^"-;L*2WH$-PTUYCKS4L,EWR.0[(IUM[YMT-L^8QP!O[CG4H^&5
P/'_AP^!/L(:)A-!NL\&XQ.@G0'.NM$.#93$_N^ I5?7XM*5-]8@5N;,J$%]6S%64
P1O **4(-<NH5P0K.\34E6"R!7GA:,MYMIG0475ANJD:A7X[#!0]Z.@WX-)(CM7.!
P2V_J4P_C<K=*RPB:O$%TU-0XL(T$-L?%+A#L:2YH5OUX)"^._!ESG16KS'+R)0]8
P;+&_W(].DH^%@B2LULO<71CW8<R"$%I[PC5[S,T-VRPK/PU9^5361?JW12"<#3(#
P0$9U>!,:,/3=,55&<!S,I/>/\5C6I9E9<.<GUALE 7<IVZ'J!T)P1>SLTOV^ NG1
P<FH?_RK/H&, QQ9?I=2E[*)$=7X4]AZGG@Y;J^?T'2JI"V!7 "6RE.+]"I9CAY!%
PH.RN.Q)"#0^\ JOT72^FZ^S2)HZ+81WM ^4&-H3,</D,M=MZ)(<$SB(X5_NXOE$;
P%HD5O< @&P[PO N/-HG]L%EPP>[#W)/37X;LHB4[T(R["URF4Y4A:E!-S3B>H5_=
P;4NZK*;1IPSQT;)N=$P\+R=Q?5'Q]J*,#F4$M*#HP<4="+,5&)VS6^Y'24^WRGK]
PMRPV!>+HE28H@HK>"/!9*1DZ#W^&T?@$0([#TW;91H@& '(T?3?BJ]?<Z)6K_;.E
PU*OD.(<I)2/A_M1$==C.;9NT\T+VGHQ'FGX44DR7(D+8W_6+A_^>&2]"70GN .#!
P\#OG I3FKZN.FJ92/^]*OZOK7*!,-S%1XT)#*O:WXB+A@KT^X$/-)60\#CI/UI 0
P6APT 5PPW]3F^2;!E_@*F2#=+LGSF=T#6_P2:MDNW(S*./_*1F]M7]UH.6#GCP-^
PX/J3G!S]O,B\D)<$S%89)(JPVATZC:6E<^EB2$1A51>D?J>$[SLW 3I</9FB)V+ 
P]0#9PY7<Y&3MI/G4'RSMU+]=>#B8%E-W?:S(RMVF99NK7M=V!H?R]?F1[1IBGMNH
PH B' DV;>P=*2BKA$K7<1O\%@-S7KE&PQ'B*ZEY,'[:^:RA?EUGCL-B)&E?8&UP_
P/L6\$4#3)/(E$=<H(.4 TM"7W[N<33/_3EV,'[<EC6Y*F$["<QJ5XOUP ?45V-.U
P1QN/2D$P8-L$JC)0VPX(7:/<75V,3DI 94\5B/KXU@"[UEZ-Q;<7!ASB3OT4#X=K
P!%GNATMC,#))8TT7#$,"&M2SXXD* ^KL%7JYWT*VZ5=OKO,F@IH_*DDTC:ALCC:G
P0K/XB75)336;O/>Z,6W%4G&\>9_W!T*#Y/X*;6P-RB+II0MS90%,R_;J]:X\J_$:
PHMQPX)AEPJ87MKTNL7526(KU4>4+N5*X:MCJ39\29'YPMWU-?BA6IF9</[T<P,35
PD<\N;Q@1LGEK<J*W%"+2FUZZN1 ! ><"N;YUKMYN# #6$C@Z$_!9'8"+XK3)5R8:
P3Q5)_.$61$( O"=DRTBY< IH^F'$;7$_=>4C8W]$E6: <;7X-)@DF:K#L%I'FM,:
P<7KR)9")4W<STL1*5=D+$TXCZNH6Y==!SR4.Q6(8S$Y\RF-B&]"N0[$$Z]70):8C
P%P9?[R97;4NSCT",>,"&=*D\X:;'C#T_753+S5F1QS:PVDL$=+*>(\U%!$;]D]&]
P5%O\JA[$63AVG'D'F?2RPXC?$@4ILZ5#[>5^V!%ZT&#5D7VT0VAV8\<Q;[LB&6#+
PL@4#9=*,$L=^S>'X7I<AL^,K8%W7F[OWLW?YIBRT1??=<"6/N<%RWHHV^$D'G'<+
P+; ,O8<[M^?"EM#V_D=S;,[<,CR5A/(:/SNVYCE.\9HB(YN'E<X&<CP6^AU_"9V%
PE1P3H)?HW*15S\6M<2BM_@33CK*?Y MH>AO=>8FD%4FMK(#+3YJL6=(K.(&#?]JP
P;);DNU84VKL/Q83)7V=1^,GO:BNP-Z7C4VUD!1V'AJ@YU"DK[:')+'XU45;8Y+45
PUL%S?#"<S)0@NQ21\WF/H)LHPX&F2\FU!2I$"_DSEREH\6PA67.OMZV'1-G,6"EE
PBT1FVO,S)^M;9^C=>ZEL(V*^0+@)3(A:RRTNGK<$50%Q;3F=1KP/SA0#=;G\C6GV
P5:2=F>#3GS69V]$W=VKC(+!_4\36T53@=%X8B#2>-NOOS8_E2CP\9 O_>.'3N$%(
PM@$B[_RE-6PN&2L#X8D6[T#^:&W-I4RLX%A@.%Y2^W!LB-*NQU",BKO)977=8%K#
PT+9:L;Z>V'LQPHXUL!3>@M2-7"+DV5;C3K8T2@2YA@Z,O0RVH45'\"HMJ">KBAMU
PLU#,/F_W_G4Q4+T3Q^=._6]:ERW62"&%L[<KR116=.BFAT-%<A]/PQX\REXH+7C?
P3=[LP(PME,3=6V'8S'5/\K[BFYF>V)WN"G5CG9N)5CLP951J_7\X8=J&:P=$<#1$
PHZ!J(U5+B79F.[:&[:/0 '^L"B6!2!EM7Y! ]",'I>#  <3)BM1LD^X_S91A)S%_
P:G,N D?XUQ]PI$_;).GQC>3:;:^8,Q+KNW2#B!;+RUNRD3#M0_;EWEA BQK'V6&F
P7RD;Z+(_NW%&^]OYI*K J/>3\[P0"U&/KQ2>5.3:4?,AOI1,,!!9OO,;M<>-?BM 
P!#FDC_'B!V8#8XZX^TNMG^2X>EH2( C6*?\R.P?/N,,#PAX[+%Y>CC_?C(-7HFP 
P9-LU*W*X%-,P?$'B=?/6%W"LD<8:X1O(020Q4X>VG#)B(N)!SE%.OI8*TPB@FL\'
P@<!O\B;M9A.QL&Y/<-I4MF4,7$ERD!.=#C;>L(/@DL"0T(!78,(U7+PQ^E#,=<;^
PH'="0YB%DO'4-1WNAVG_!O%1FA-)5+ELR,X;0Q28YBVR^$U2#CF.E?N[Y76K1DNB
P7AUNHL'!L'_*W;1''<__,*<]LX?<E[,#_TMGF=/N$A'2,AZ:9EYU?^ PR? %6V2@
P6K@8<N9:!N,,&+)];R) Z7  :-J ^O)$=9REB*E/B,JYV-_)@56&TJ2\7]=O>S[P
P*SJ)!*.#Z\CJ^H$>-_\ZG;)>9V9$4A+LX^"V+'*N*93W3OR/Q[_2H^224YO1J6\$
P*SCZQ1<@N^>@$_NB=E!SXD[D,R+>3A>G3SM8@>$)(U@4KAVOL"2<M3&ZHQ?>LE-@
P&Q XK*WA7;!G)2M8B.SE'TIAKA$W4>H;$40_&)"Q+!SD\ $5U9GT QBC7#"7]$L;
P<AWNZ%B590?]!5(W42:? 7&0>5RRG@37H^$ZT]FU$<X.]IWHGA-Q<K(UEJ.!RL/7
PK/CYGM %M79]B;X],A=/N/2*/_Y;. 5#693UYYMR6WTJEL*+9\Y/(6)$\G_C1(_<
P&LJ0<2AN"MZ1.MG-6"39? L X%,70X\./X<]81L=FEGLWP/^[HQ+O4II9T;==YKZ
PHC(YJ7[A4!?YV0_#W"-KD(BW<VL1U+;KR_BPI$Y4$9-*0,S66#L8#D9&]@J ;K4_
PO1]N_[4A]5E"&9TKD^I5RA3Q$G<)K+[+ES[.UK V^UPJ.Z]FJ#9(7.H):3D$O+2^
PVE@486M 1JH 5;(LS(0JU#]+!Q-'^,5!_@EE7FH0?)-KFY8H+PGWSD[(B\!BZ=0E
PGK$Q#'Z*"N4]2^N2;..LND2;L?9_? :)N!HP_:S^I7L3+:/B(L]H]E6(RHO"DQ.R
PU(! 5GU<LGB]!'G8[ <+\=P/$R-YGUH1E>;8G5U'V2-F'/3#POX/H&Q SNX"*!_G
PFKAG_DQ E0^Y%# :5(2[QJ@B!8YYGI6L%N33@V,P"".1ET?OOW<W!<ESLA'B!P:)
P,JU/?%,_R\'.C-S1A5]GD0#B$C*,]@*>REY#]QA:8!^26*]R'FGO:>VZNQRY +4_
PA4!@=RE%GKOQ"+!U!5K()P;HY:QQGE'*MJOBMPS<XN\K55]EXE1Y?=UBP5M.)0-.
P#Z"";H.8L?>#0B36_7$Z%\K6$]!,G)LA4L=4E;7S)L'L_>;T^#KQ2G<+XE7!6UR<
P0W6C9 JN\RKBO9 N:$/;J>;WZEICT5/DI]5/H&T @\C',)<C"=Y6T-@G:EN\81AN
P I:.)'ZP&1J4\<4!6BA<-@M?IV!IR/)WMOK(=I_6]<ZO>:YZFE-E6Z/1%QI,^8$*
PO9J5Q'![8/F<KJ BMEB!DT8<$LE2GB7A_!F9*:@+H[HA]7P9?R[NT4A@[9RSBU$Z
PB\Y_*;?][Q=RS9K(]UU;R?*5F2PQSQ=.&%@,*[U>EB=[RBT2G4V[@X4R:]J&AA[-
PTU!M,Q\]C9<GDO ;)THS&*6FCXJ1B "D5;/FTUQ<CED;W^<F<LGXH,!JTFDR1KI3
P ;2-5_>$\Y=+EKN@UB$N(7BMML@$[R7UNVMM@%VM"_,>9"SJT(B7Y9P8,6*C:=3?
P*(/:[F2M+PXVNS2FT3OY+DHBZE8KZ@5"?C[C71-G[8[,12ZYX+GT10<96_3SN6)9
PW$O3,!B)J[,_ZX(A,$11JWEHNX1\O8#W#; )7)Q0$OSE+BED\(Z6F8".?P^1N>.[
P^3SIZP,X#FN29"ZP/9 *0JG2*5L5I,RK/W/[MUW^)B6J8Q>V,K&S(#VSRMH'_N/Z
P]2A_NEP-5,VQ/FS"(AM&KJ+9]3/#XW&^GLW>PC:=V;*U^S#RA'U!_5$(4P>%)0>%
P%?,W-ON6:]V'<)Y2^X-WWBEUTN7J; Z9GN5)@@>)S+ "T!<:L6ZJ3;1X-)X%NGTK
PJM#WQK"9@RD-&^:UD#>Q-'87^]9$*8+)SPD%O/_PI3!,AH)$*P<;<J$ [L[5Z;^F
P<FTN)/X8J]46L\GZRU=NKG@J"N6N4UIMHRH([(0G=C'((<57N7UF&XJFS77Z"K%N
P*?J[MVD)L7P^#(=-D$N=OA+8K9)3H*.$?AN,0.+H3(S0' R=VSJXK3T1S6?UJS4*
P(@")T:MB<D?%G$FJU8C>!HW( H=EZO].P^Z=T4Q[(=DD4<?-AOIG>_!<?);WTIT^
P(8N$#S4.0?$EBQKL82^8?Y3O:$PPM0 J'[S/?G!TJ>\?'UXODG8Z00(3? (#R&.\
P))6WE(""V-<DH&?EC"5'(EY8W=;EC/JOKLC84,G\U8F3)RZ.0V5EJ>-WT%9[8Y"7
`endprotected128

////////////////////////////////////////////////////////////////////////////////////////////////////////////


`protected128
P?+)9#"+V.E$ANY.BG)2PC,U'S:"!PR:&P@-%,4ORO>KE-_ER#,[G>X 5&#C5I#RB
P<U&'.)_0]K&.#XQU=.-A)JE:*]@4C KT6E ])Q@G95=T-MG;L!*X$87OD,MN@@J1
P9Y2UGPU38@[ XCE#YD,R)4!88I.KI>9X-U\7.Z8JZ,1I>JXHN)7KWIF8"E.=RQ"P
P/Y11,!6L0<DKB:5G R&.(<+JW<M(AD6M@R2PH6N&XB@2;!-,O0UX L^V%U@5T*"*
PZJHY_G-#TN]7=?&R>&@C4K[CU":.H:R54*DTL5OQ>;':<Q<O.J52O;:V-?!(T,;B
PC8\C"4/.HJSJ1^T#?OA]%F+W_!-;Z.@G5\X"#!G$I&4(#COWGY!OVGVT)!<3,-B7
PV)MIO>AKB9#_^$>Y#LY$ZL>!/HEDKC)3M[&_#QKH)NDSHW*^8LZ2W36+BAL8Y$B_
P*GH$;"(KCZ.<C?5G*X!P+"Z!Y<[6.:3JY\JG_!GR5\ NBAJ)5<72-<@8G /5=W5^
P?<7]2HSOE_JLSN'5DI>41ZTOO^M)_1N7C97_"20[6=)C]G&1)1/KI=D8X[.\#OYK
PG#JHZWN'/\EMKZ#GTH5)ZQ(ESO>P^JZ"=V55+/SYY/9<SJ4/),"H  &_#I?]Y3?6
P:H\IV6*P:E_4@ &A)@@:04K$^..)I$,#5!&'&PKO1BI4D8B_U2A*9)[N<YDV$-$+
PDC6WI]<G^3,OWKEQ:!?[\O8^B3W@D[D LR0_& 2[V;F^1;H35RZL&1*MSABE:E\[
P13;6\OP@2.TNBH_G>Q'8$ +\#=N/VJBP.0W$42W:SB]]+O[YZENP]"P9Y0L=F]4Y
PE+XH,=;T\<5N!0/?TW:G%M76:\HRU5.J[1K:S)?!2^S. P5&EJL%H#\[EZUS+EXH
PN$=\N>;X'P.=O:_!H]CJ?A\?(O>YC^];#42\"C"?S_>"(X)5SV-?QK.HW0MC0<$>
PJ"$0\5'>&>*("-?S+ X%OB"?N.CI/I12MV<2-9JOO35-G\/Y@\Z1/N#"*BM'"]>H
PE'%WG&M^:3W/P*DHLD! XA/J:T9/BPFB&A.)J]]]*^5Q''!<GRX1RE8### E*( 0
PM'&'\A- FHI51NQV-+V+RB_W#5NT"X:M?F[;0X_RTHRR+<+'K2HSA8Z",U"B\V/^
P$-@!U@(8\HV ES*@'L$PVL3_US^?]*AJ+E<>D,%SWLD"2U%8EML)X@OXR',US,J=
P]G[CQ_#(L1")NI"Q58#'IL)(%GYO,T?U^^2V)T8_\"(?\W<L@MMWJTX6V#7X,9E:
P"L;2L>G!>Y5[QOF 7F9K@$IK4[!L/!4];3$WA503-+D.-Q.5B53LS#H Q]Z'0HFP
P89KIPZT$L>!+PU+7&E)8]JVS4 014TE\'FN%%G.%(-*/3&/+SKOJ@.;40XL]M+F[
P? 2.#3DM%+A;_U>OH;L@7Y)&T7K4\LW;'9PDB@V%,X4M/]X<(QS9XT9#[+%OJH%5
P/49W+M8N0DN9W-KJ<H+62MM"V]-J#F7:8,:J-!Q,1^E&B<B[QO/Y1[VQZPQZ[CBD
P [D\UX);5"O'4KANO$$FV%UIV\RRNN]"_>SV"E_5WJ4;'AOG*( T4HG+#F\4<W1D
PE(SF)C3Z4NK6=3N/FLK&"0B8FGQ&W#_9KPL_65T<_IN2(3=1$Y@%KP7[N( W$;]J
PA9=D-ZBS,,'%O\+R J9TD+><3%V"N<QP5!_KTDP)H+'DZ*5,6!5H/@M5D50^@+6&
P7CNR<\454)>*TT\I2@:/IM&9#]Y5N_08-6?>35TUY?B[, ZK5#.]-L<V2A:E\2IH
P;F%.:S14!GBN?LE&[!H\[EK/N>PB[K-+2;J9#BGV$XH+@L>D#?K:W!W&T;MH!FJ5
PK=AO(4Z9+X$_:;NU6NT0]P4-HWD\9$ZM2>;S3MA^NLC+P[BB08$'M83]0]@<QTW<
P4[S&CA6V,&DR*)Z:*C?F6421GLY<>&D,"R2.CZ&G1N$J;)D[(%%89.5CW9C,&2DL
P4P['_8.OQE4X<:\LF-#-1N8K/Z]'A7/EJ@P3B%H[-R><!P/G+GD!X]%@P.=\3/!O
PFX6.7"Q"7S[&2P#I&;PG8$:.>Z5RYPT_1M=Q K]\D<B:N-,J[,*V2*/5X2&>^VG?
PXK^%V[E4<94/1?GRNVPUU!Z,US'(;B/QL+BM#X8_IB>I )NB"AQ[G=FFP]3+ ^?9
P$F(982%?=0I1OZH2,-]ZFI5-8OH-GF7J[188S(M1MSGTC%)KU$"/J+=+#5ZQR15,
P5/G.VN!O&NQ&Z[6^N49*+4JM<S51$]IL<9)/J_51M&RUZ@:)\4@'HF[NRYCOIT6C
P/D;#[]T\=3YP[MSE@N-*Y'+0PB-&5&^B.;R#/%46<1LOC>G,!%NZHZPSS1#F;)3 
P4J>M>G=4\R"E$#51WTRTG@@4(M/LTC>H*R<8$O;!84?IQT:-0FR';Q24QBDHL@.]
P?H5K@5&B&EA95B/76!8^'0L@,U?XY_KD&N2OXC6]>S4LO3 :>-ER]4O=L*6R*N0;
P!^BUOOQW6D1&]R2WD8L+E-@A?GM=/XX![-LE*7E 1WZ]=[::A,+GN/W6FU[&F7T3
P;#,_N%\KVT0Q=.D&\QFQZFY'TH/HS/\53M@*W[Y,D%["E3ZL2\FMI\@P[T:%REYK
P0&X>*7N! $Y3&/64>"T%I]'1&KZQ=("/?F5N7RGN9H7H5%F,:20N^B_]-V=]?):Z
PG(5=^V/)^,I_O@LZ#4VH[RY6TP89^14\B,DF[+US_<U4< 8\P;H!*C-HHJL0&XJ1
PC<RGOQO7TCZ153B"R"CA;BP?V>-OB4[3XUS+ZZ:6&"944;ORT_B:_D!80WD16Q]#
PI9GC'R'Y[MO\&%H\3WE6G2ZZ@8C:7,+*O0;(9R%L9<[0D#(V_(DVM<%!W=[UP=9E
P2Z^$)&.[-+SF&CK0N"-'1)FN1]V]EI21S  )_J76&<G 1^2;S55O85;U,G3*7D,2
P9##-#VX+6=6K_)FCDUC^&W,1]>N>VH!Y^3"TW:Y"176"=@M@%<D,W_S7NAE0+=<G
PNM37&(?N7?"! " $*BM];&^P#SC/J#*FFC.K?Z;J#X])]^0KY#I6,_V  G]LV8N7
P !F(<J'93C$2Q'3,I55]$%XTA)SKM[5LHI'8F.Y;[]Y3"*6DZZL*C5W&I45S#<=C
P9X!_7UC:<?)K;G:"GVWA_"=R?#-T<2Q8TC,>7X:[[-&'/6TVIO2Z9RF\%,V=+O7"
PB"?.]>?SR;R2-VR2%U6^(^O<*+L39@838U4A\ZXZ$X;C@9N<K\0WRK_&-3MOO+C<
P*>&P:.H21 IP==TTA"I)XJ?F5$,'@E)%F!K-8ZZ+NU%S5Y%=S&G$1?RULFFBEB;+
P['O?>8CL)K9I(""D$=Z9'>M.B@4YF8#(KBD [!R2,9=0WSP5:Y+Z>4:83VD<7$,S
P(?@A4)/Z[,^N)ZDC>KFW;7T!7%8CC8^2:;_5O#\=4QFK>OA!#]*WS 0Y^1_W990:
P54=H;+3,('K3E"\%R%\1VKV?ZDLR'?*+IZT02C=']HO@3^. #93^GZNU%9<H4SE]
P8]HB#D\GM*[$GV<W(\2</@HAF1TJ2<)X:"B)GV+I":7_:$E'-% 5&'SD4"E0U*8G
P1L^P)MM2%FIQW*Y$4\U9VMLO^"I.=#Z\QQ.R.!5%*QEBVAOHSAP&!*+*0K7("^2G
PXDM;A#>J=*,;7^+B",;5Q:-%3/1Q[$8N>B^Q 2/2RSQ@?[]_9\2VFF)X4<R4[(0!
P_G"=]5)-QZJW:YFKLG/3%33\R/'B[@E&[] A0!TFN#8\*09[#V[<_'1 Q-&9?B+D
P'Z1DL1;JWQ7@5/\SU.NR(%L+YBXXRS9R 0NXM[75U]+=OYP<*]2MN2JAFF @$0<^
PC."+RX6O@#8IB51$@0Z*_L#75(^UG "US0IYG3.1TP9_TM[IP\<8<I\^^0N4NBM#
PU\.N!1VY1$+VHL@Q$PZZ2+&&@CL1M]:R?3!P7 %:.\FD3>+^C^7LA'#[KP1E(M[[
PE_FS2OI(0I"N#\T!_<.0H7!8A5A<W=DA.[AXX6YL)@PA;3?P/%-WOPNLO*[*JX?H
P2)C4R ZA65@]D9QN2*(^8BU/HPB>)Y?%P[3J-H2*,&Z3R'N*X2O(IDFZA=5PH./*
P'VLN_;XD+F!/G[25IRJ]R9"NT0V_><Q&;)=G!_=TN#-B/FF27G#X""TX-UX1/#1(
P$HG3&;[<U9'$V1ZDF7_#?5UY*GGD[UE9P/? <AXF>9J'HTDE6C/#\SB-97J)W)D?
PM8(3_HCAFS]'9X\&&C,4LIJSKMV<EU?&>W*?I7*,EM:JZ)YN)NLDHM,=OJ)(2A$D
P!X,GZ;*&&1W,BZ'^7L"R3:$?>LXNW! 3:OY%=I;!MY-JTLLC%5;Z_DM>O:%/*$4Z
P0)F = :CE6W#+7%UKI.FR1:RG\TVFEX,3M'*V?7C:BTV&Q<W*](A>QR,I5.[= Z^
PUM7ZP%AIQ")+..LKP*P%@2Q^/,Q'AP4&VVV%%S'&L,^2UP680>R1_[^->Y6@3,;,
PVD>J+)KUTT9DX=^B7PFMRBSFX>6C_$U>+KB4A]ZR;.;>.CV'-UD&8L]1?9-ZTR#?
P-1^7<DW16?5Z2M63%'Z\T*U.6*$02D#QYE$$4+9LT]T^2#CF,S3UIU[^61<F<4N'
P,74#_J-WM^W/FZ_PLD";#4-A0@%6X";._%>BXX#YF-=GM/,NC7/"'/+ YYKOI"!5
P@]@+K-\"26PWLPGPAX#0BI"*P_&AZ1Y<T.!_EOSE6JF*/CUC=.;\F;FEY+?DSSB#
PW_JA1E*OQ^\FZ%\6"S0,AQ53&LNXFD_?W3V)M:<KE%UJ?8CV5/(354_:3+2PDK?0
P',9GTME93J-_H[UKGPV0_"#X7_X?\I:MT*]RT);\]""!X6;5"CXGBA"I)8W&!%=6
P;NK0Y^E_RB6UZ]HIBCC]@2$RRZD;ST&"4\@(U7Q!@3MJKYJC#NV.VOGV.W):##K^
P<90HG5 34A@>.1?/R!:G62O<G7K4/[GT<$T-V.)EY'Q"6/Q!D_HQZ6:'@WX7IV 8
PNR*+ZP6T:ZADNZ1+;AMEUGFGE$E!C1,B/88_<7@$Y#,;V+"@1X64- @#^4.W],S5
PIPJTN@UIJ(Y;#?-9+6OM'_AXC!\H\P8KQEO"UU[3)7V;B1<%D7M[6X0_/)QQ=+?K
P97SGEU<#IH45#JG,GJODKP9[6?6ZVUF0L3.(!^*@=2DMX[PUM'C<I<0<5R4@=_ %
P\P.')\ 3,+AW#=JCFN90L6(0:.* UH1%'TB'9P)==]=:JKRI3Z?U,!AP+B18'[8A
P,KD'#<9KV.E@_DK"]T-9E%IENZ '!?=5'37"YV5 \UVDIWB'AC$\*[70\F#*SM/)
P*BDA/!==7CAA,+UU@7)?*1#>*4\\*J-3=3"YV?"F=#*CB2& $0_MF2Q\!E>B.0>H
P,/('GLN?CU:'@(88\VLY%]\T&U;HCKS[U!M0OU)"0I57D+W5NV'F^JQCMH'32V^J
PS>%XOS\\9[W27TQ^PYYJZ%$:#/]9;J,NTBC:7Z"O#TYUB5%=IYMQ<@T3FQT#@E(Y
P9+]5>HZX7=#)>S7B[KKZRH<2)=8^?>(DDS,6I)CZ_:)'6;09]MZ7Y4%.A>G=NC&@
P'EXSHS*.YX93_].&@67T1WK/P;9_@>7G@S0Z%!5JHS\DC8!;[(K]U 6T/_Z_K%L&
PA,[P[Z%L_:"CHH:AXA.<"D D<B)OUL0CL,ARD0[Y>$/'[ATS.S/#=*:!B4-8WD0^
P?^!R)LY2PS@4Q Q94Q-5?,I@]V7Z-@305OI?H3.Z<Q[E\'2JZC213&3U.8SQWCC-
P6Z B"V]Z3$DG %_KXE^A,QHXKX!Z^OLSI,F1C0YU?:UX9U!#_@W'I-CO<3+R>%8A
P,,L1+ 3/5!KH-K Q7%S4P?1H!R+4X?85-DDC2FP;C=5VP2&C6!3RZC*&=FH[Z5_"
P^5?3 U"VUN8=X,:CZ(/)\%C'%=TM? T&4PC;+^V*FL3_?$/*#"56S]?[J]X.PL/)
P@B/.J8'SYIE_4%O=KP".?AK&J^NIM56BB.&*<8"ZRNTT6-L6.D+]#;XC!W/1!&J$
P0TURN/J@DJG4U"1]!G:X&UHTN45.$&@LUZKG)\G\MII_J(NM6)_TPDGNKWQQNR8W
PLP'HJI!;JQ-_:"L!QS(*^\S/^?LE-(#MBX(O8.+N&0F3]DHIF2%&U(=IK$H%6T9P
P2L1%(?BB?6[2N,9^XIHBW5JW'GY G*4B.)&#GW33=.O*FUH%9?[4.K_0OL]'HF7"
P-0^Y%^<"O+7C#&O H36@$XB"M4C[I'#04BAA/=:8/%GJ]/A#ZQ7&K=-/19^@@S\P
P9UX9T]-A="1/UXK!NEO)-J-$JG""#0*-9<P-&^%4*;!7WM'QIG]F: 0]L?"2[R73
PQI?S,J7X$VN@L,'Q J2Z*)"@BJ9(8JO>[(8UC[=8ML[UB-4LG;080 =3SNZ:PA;"
PC-]*4_Q]DM =;TW"[?#^0' F+KNJWIKF2SFE$Z4$9U\M6WFR"B[W@Z4)#4?2#@LR
P]C4FOR)V! K,Q%C;DL8AD^W>'[(77VX0*'GEK72H7W?J?P.D#-N]H1# /S$H!R#9
PG091:05[H]('H 1MV:'\=/:O"L$X#*+SKN5SCC**HC;@GD[@:YNK2DW8\/JI*,7Z
PPS R0PL9"DK5[P3DA&>YYO\IAUN%PEE(R(U&U^C%IO+3;!)/#I# \^97F :B*11N
P2!5F+7G*DKK_3\''"5MGKZO0[5+%@8CI*)-C;U-6HC;UML4FJ)'C#AA7L=+GLB$Z
P <7;]*0U)U[8HDEY!F;B>D^WK$F:L$'VD#1M<5##V7X<GJ%.LM!\O_=YKA5_^5#]
PFR56PVVS2N/GW.%]D;VZM/XJA8_LC+D\: T07_^[_816GLTJ=UJ)_RD/VG. ['<>
P)-8VWK.]Y3C4Z%)>XM[=R[S+>.UEG;P-,Y:-R*6=X[7_%C;4OBP1HHL2Q,%-UX+<
P_75EPNMYL<IS-.#\XO\4^,'@KO0K%VU#1R@PBO26@T03E'#J84S:E0._2&P*)(99
PJEOZAH3C>(O@JY;+".>2\ @M,112TJ_9S,P%+L)BKL 10X2HY9OJ[-Q!D='J^HV)
P7EZP$E\P>79K#)LI$'9V]=,4Z-)]/RN) X[^OF"$AA06*5ZAWR]KB"]Y?= 0N9,U
P.+I9$6K2&>Z0IK20&XUQATNF,0CY6YG=\Z\I![N&BL;YDYU\K4A?0 V/:;K]+%"Q
PZH@#J=/.EI7/^.#XP/ 6K&O_3(H3? &>8$D1PX@TJ*)1(=!9># )G8Q7@<@:1VA7
P')1#]MV01I(>=SW!#?VIR"[FH?-82Q'';NK-YWYVBV?*R=[W&I\'24:U',(1*X[M
P[Z7H\QIZ%XI9 VA>8&-EOSMPC"LF66@?,_L/J;??LS).H%C75T^V31[E\R#TJY*G
PPVT?Y^)V,%':@X6SQ\ 7<V%;@06!Q<N  JEH"0?=C'=?PS%^V *[D:2=!ECJ>^?/
P0]W9X42BDSORC<VCM:WA"R#!9'Z])8IVI<9\3O&LEV-CUOSO.Q&21DCHW3W?&J$D
P')FQPD-]T;YWJ&H8G M$-?OK6X"9(I@Y)U0U+?B[D[V)A<%5M7=F?EOI9G52@"/X
P1R^TX0 _9WG(D,:\;6&\Z9\1OL1LY\EXKAEKQEF5@>=(-":J11I;;IX.^[9SJ+P^
P5W<+QN#_4&[F:3E0O3P!4>K\! _9I3]Y0']3/:VSUP.95(.YQ=.4L$_2/:$&K@,@
P,3[3;D0][L5:C4/(,R[T=+U$R.T=JGK5D9J\BB@YLHQJRZIQLL KUGM=]H^32Y&7
P2L+2KA[M[?"H@.68ON6ERLH&!-F#09^K_^CQKN/OS5UZKSY4R13HM,Y<M=6P<\\"
P.OL@B@9MMK2 44BRZY_":OOE_,\!K!GO$H= *E$-8WG%4^I?+M#I5O7-Z:R>X@OI
P'K#+\9L =,)!WW2V"V=)B455N)@W;KYX9F-[)0E8E-DP=6WN9M]A%%M):I53,+[!
PV1AI'T?U_RI(4O.X9'RPHA+S,*1HQ.GD&,MJ%CKI+"*SSI%[2Y83#+9G)\C*^V_]
PF_30!WKB6BX(FYD;-511Z-$,U+^<]@3FI[ H9A+^9] +-%0WD1N' .IELA_?$@^5
P^<L;*C,U8M!$4S&*J_K>KR6+"B+M1<JHZ6;KN0ZKUMYH?UH #'FR._\JD?R\#<87
PEEP!T">(SF+NG>>FHD^0*]<B4S9,)X\BHA2%D[XV2"8ULT3VX(I>C0^7&Y"".9(<
`endprotected128

////////////////////////////////////////////////////////////////////////////////////////////////////////////


`protected128
P?+)9#"+V.E$ANY.BG)2PC,U'S:"!PR:&P@-%,4ORO>KE-_ER#,[G>X 5&#C5I#RB
P<U&'.)_0]K&.#XQU=.-A)OXSUI3BS,P67[EH<Z++18NJK78%]"NP02-^'9PV5QJX
P^B1.EC1+#HW3YJMC$GF=<7J\>X$E"*RZ%4B'T.].=XG)$D44]RDHE=,[.OK5+NHF
P/HT*8>XO2>U9T"("6 J2Q4\V1-X%#;$/2X55F)G$0U6!<$54VJT)H[$BJ?#?S\^C
P #?H]JA1#6"#@QB?QFQH34N>IX:^UWR"P<5CCL;B]U.:Y2MXMTM'A#O(_3L+\Q[ 
PRS']:<GLW#:'$%>V*,;2IB\PS$_5UJSC='FT=?R5)4;/*HX'@X*0F[Z^E6KMC=M.
P\T*:XE(&O 4?=40Q)7<.)6 'DW0)S=! -+Z. >.'[=W.K)J3>T,]B:4H/PNK3;3Q
P_OUE6DIZ&TO I1_XEQ.^OG^R9L>FSHF+?Z]ZBM,M-.\[*XS^GP\23D,+3-V1GPG(
PUJ\"E&8?YW8?]/EWB$M(_8%5P3'E5N,I4=AT W\&*KW9P#:1DH/.+4,K(\E[4T5R
P/Q<ZUG;TOW/&88U#H\$81] _Q83:K%3X?G.#<FU+-NHE0ZE8D_XL/ORT.H!(-Q_L
P0%?8 KAC$8@8C+SH&AO[$/^%7N*9LZ+:N].]T]_ 6U8:O&$IS4=%^AMOS*?Z1XA*
PH746RW-<%>W3LPU-T*(N%,*C/&@X)81)OQ')3@1;YEFRRR:00VB"3<))2*>(E]:!
P*$E*;%F[7,KQR2GU[@[B=& :#X_!V$\(/-W&Y)1?X#$R+1I_8$7\T8H3@.H^F%/S
P[$YD$=*O94N+".[*$8&!#^"PFG]QW+.SZ4^RJNU!RH:V4.F!4@XI&M&[,&J V9A$
P4YQID$-L6KH99]6',&/CG0-NQ/D18,E".3QF1S)PUYE;ME&A$RC]RZ'S#T4!IZ.C
PYDY*6ONKH<4MGC!"[P@A>LR.3W;+Q$/2'MUE7@GA"D8FGMG6'P9K_MP>PGQ$DWV$
P]SLS%+PN@#$%<OT6D_< U@H3%<FAM@% &V##^S'Y+*\^A3)K>/AK>K(!_?E(W W+
P<YJ!#H!1DE=S5M]RFW\OY-AEOAO!,(.V F4*AA#XVQ!$0GC++KOB'N2?"&,\_\$Q
P@.;O02]L3(KM#=1$'FFO>73?!.UP#Z(*VPH*V(.![TAZDYV2E\[@;]5:U[L40WLC
P&@7)5Y43B/UUIS'4?+SA#![^U.%+W0LE_@K5U5\QZ.Y.A+#^GYL=7;N0KN7FMQ1B
P.L:8#%E&209+Q4/L>0\@0\E(.LDEA)U+"(=)E# RBFIG#M=X&5:_;EP%8W:KVKIS
PDYC:\MBGDC66?Y&J]#P2BXHD!>1X%;U+ \]'T@5^#7.)T>OIJSFRZUC5G8H?6RPS
PG6NCO]C8WO.:>AP@Y&4:=5)O(RADS!S&Y:U*T:.^\'85S$\@)"E3=WQ6#)35&Q3I
P_7?Q;%'+LM9F6W<DY?\E7?U':;@@QLP6\RG2BM2*7BK_== EX0>1;>'1RP=']O8R
P$G<0W=<N@HE28__K.6-K B$?1=+S3>Z#G[4]@(&6_A@RG3Q".$C%:.E_VQ^PWW.P
P+SKXE+ 9/!!Y^H[YS+,(*#3F!PF+^<.O#3_@^=Y.4(\-G%K/YA=%#[8@M7CV9.I@
PC3=%?.AY?$-$Z7U>'?I;]3S:/9OB" /$+&GE%L^$055>\<9L=QV&[#FF. #M@NCK
PR@+$$MZLN_I^FQ/=2Z\K90N*^J.Z=!%EFNAC]V;:V36A86#L7C%/M\R;R2=9>)+6
P9^D@X2S+&% <'S"A6T(E9,-(T(18Q ?MJL60#Y@I1')\L\%AI#\FX0$KB"A#[5,]
PO*2%E.PF9L"&5<D;7ZL?I!8+>S7(78$=?@H/(R0$B2IT_)P0/#5[-]<EIK62"%)*
PVGS#-F>XS!>#-)2&Z0FY^;AC5W' Y6P]U$_3[B+7(4K!&_,)_O<>!1K<(2J5,*XH
PK.D#9CC)"S><0I^_3^0>;Q9?N/"M]'SONKQG1L /=/:4?X0]^Z'@]7EC_WKL_C-U
P77YJ;K2[:X6ERON3MA3^KF1)9)R^A&@00+VQZ^$^"ARTQDI'D(/!HUG[)+'T0)UL
PX*$L'2(3D^64V\8*V,I=-U]<K2QN)PFU2BSPV6N0%,>;*=UJ*59#DK]!15C<P ?O
P8!YOZ**?A%KX6EG5M)LH6]I!CC@DO&+R_C]KPBY%0-@H]HJCN#YC>7A$U(8!Q)"_
P4.^+MK/@J7VC(L_MD[FT'O9E?JQDKT=OXC(>B;#M\PM3"D8<8^$7RL!K_;Q>[@JF
P4TGI\*+YI:>37]X=8W:>-3@J;8K#)^9R75OD3J=-7,F;;VY")T.<GRD4TW20+Z$[
PWE'B']];'4?3<E)6KQN$X #*/\ (S?]#/@V_DUHEJL5<3X0OL"*YA=0.*Z<!$++E
P<\)=Q+C'*0*VB)&A@2NG])ER48?!1#,9WY8_MRY?L$2 Y[3KAAW_,E59N]5TP^$I
P [BT(+\D S9+*7:3H@1")CY*%&_G]_ZGEDO^)-'P_*T#0+/ET1&+4GU=^KJ5_>2D
PIMY0A@66D"> *WZ_@(' T>]7UDB )@V?2G3=!$T<P,I7</@\VT@''$?L+.T*M7NC
P3!B2*U]7G5HZ]1(-"$/H69V:B>":TUL>8/OSO;'Z_ZB*@#B@G/U?E_-GI'7R(ZLM
PP<U_$D]K+-2$!Q5/Z0MTF.\@HIS*)]MV@=@_K818K$S#)53Z8^%UOQ2SES?6_?@+
PJ, WC.$"CGR\&V<B#L$VVBP8-563HA))@ZZ27^?3L_8PMDI,*DU2 4R>X:3TIP/?
P@15"<+X:.Z^N3[=40B!U'<1I0^5FFP=[Q2JUKQFM]_?ALSX3=GKBW6S.@F>P;,F=
PWZ1DH=&#M>6J Z>.$B:2,W@]WE3:9I?-3F78I$#<BUNYMH.>&4LVNKX:[5(U B7F
PRZQ;@E%/FE'MZEG1D/QF[4%2U%'Q$=*EOZ4'*O+#5KC+C:8E>:\$U<5/BA<*LXT(
P6_H_/XU=-RMNYA;>"W[\,SO\!$-(.P[*4(XR2G,7$\C,"38X&Z11LT<F0/1'^U=E
P*W(]Z15&V/89&P#>21JPJ+P\)8=MK:+6X#Q[<6$4P: HPGAYFSQ^V],+EJ*J!MI$
PPV]6MR=HTJQA>H=Q2 ,?3LR<0*@/[*%20@74!XW,*3O\.N_%AF:L4R1M:+U#%G06
PUR(EI,G[1?3I8"JG706H"SKYH/'T"C)?GE0,W*S+%+ZZER;T4,2&8V;2#_5GFS<_
PJ765Y0.9PPWUU0K@]5*>A62 !QKZ$W'?G&?S5LE6&(;C/>,X@2X2A' G7K=:09&C
PL/W)PK.T D5GW_D2](GDZ3)DL!%][UR_C4)@%DM'LNV&%,[B@./MK8!#1864J, T
P%$Y:F^Q1K23&3L'3B!)+O!KP+F?]4 S,B7->37['PZR&@2B(4[1DH)TB^6)&XUA+
PW=&!#4NLP'8RI%!*J0GT&N@)4(N!3K\6BTH]6[HRCG6X)(X6G7 9JR1NTF:@SM29
P$AX%W+'V)(7DCVAP?V':&1XMJE*"*29Y+D/:28#O8-*W WT!@BJPEY+J-2NJ 9."
P\VS#2+U/N%+-F#/K'(TL*9U6;S\$KI*,PI4X)9VIBP-<CO74[6@70?3W!%DB]>,O
P@5NDT:UR(). SX7AR]GTW%J&&R9C-C1F$FT]BUG[Q4_)Z;R0,R]E*8"-!OG.E[S*
PG+:&KS=UV_+GF*'1!2V(^7LYO=P24J4N<V%I!<E=<T'%KP>2YN:W[G 8./[CO0F>
P'D$P<+<D 1C=@+D @:TZ./+?U(U68^"K&^15%!JN/>LMO7QBE1D[!.T" 0Q]L_+_
P='V973/;9N_'V&$EGR(D)C<Y;3'Y$TH0Y@,TP3:U&8TQZ@O3$L1Z=I"9IA,-ZQIC
P5!^/3<D9T;>'TW!&]:K87PD\-+?6G]E >+3<1QYOU_ (#J$H%:,I#&80KFL1^1=Q
P#U3,8=:C7F6F0\AMN?]+Q>?,'9;8)&]Z\;/$2M?\T(JL"8]N([58H NCQZD*\QO^
P/W4X>'VT)7DS/R\-J+YMI>73N*4#D $V.XD6(BY2?8T9^,^'Z;[#+Q/@%?S$*Z'Z
P5&M[N+?2)=A'O*[%BJ E@\J41&W+@!;0!L2XRP T0!:-PO(X6ZA7#8?/1DC\D*''
P))"S2>:8PV%Z4'6S:T-M7H<.9$38"S^@.;!>AY+PZ!*9?F+U4M%^'CC(LYF:" 2Z
P\-<:T[LY$[Q>P'^S-SZ"17L#P51#\P56>";O<K?#[$*>"2(\X&&"QE=?8"/>5DR?
PM]7T4,S$LK76P6UC6LYH,FGF0_ZV%N3!<?#9(CV&GGAC1G9)?U/LMF%LC;\-D3SX
P\AV4L,\(VB5I+'D7=8[;PUWW)7\>]7<?,;?^;4)3YST1,Q;'+R+.'0>>QBB#FC&D
P/LOYPG)_?8__9J_Y9$[MF]Z5E'9X[EB<=;@/U]:"TB5FU#5W; F8NP>!#KV"^#GR
PZ,A^A&!=U0RI-2&._*L6@MO MD!>V=11O:Z\MRG&L(:GQ*.*;9X>!J*.5;%842DK
P=TD5U<X<@3 ?(/+!JI(/M6@ZK%*3"B^K-K2*3]CENWZG0&!0.I0DZ%9'[BYZ($7I
PP?5#:2%4@!9 >Q:*,3BY_,!ED91+:_@3:3J2JL>ZQ)E7^S=G_)%2>HBIV-JV!JXY
P [FJS3"D>QN*KU72QSW!U^LW8Y?BP!@L=!).2U*SO\BSL@!_146$708I0J,.YW_,
P-(F 0J?\Y_$4&^H++A>@\\"?.7W62-^C6\IA(B]?R;:9".SI4U:TD0_L+JS/NL2]
P27EE4U17)W_^$ACXH",:N)+1:4KV"(K\/,&C'N;+"R6@:G"*P-3<SIA^;P_ATJ@I
P?5S.;QB+0I46H@F@VM*V/R66_^$NDZ[7J/1XJG7_HP-O1CD#1Y?AV"_@<U0CC-NP
P[R_(O@D(*PL'/[(P<?@&5?Y(X(+D5VDCMNXP)\$+V-.@3MN+V"RD=.**YB[F7(-S
PT9BG^]P>CG;]OK5Z=XHAY<YF4&#_-DP#!5MFMT2F5A.F7Q"?"O(__M>=@YZE?,!&
PNX$P%KD;(0S?BEFA2#[1T!:0C/.!^7?Z?)HWQ "$C\X]R_NG^[,"6?VBXH^&:Q:O
P@/J#AFH/TS>(2%?XE1HQ)*[=N\PWLHAPBDB@(:?TI*&#,S1&)'Y(O4.EJ_F!Y#T2
P!HR>H+@91RF<-L+)BHA&LK% 3]UF/MY[@PD=R"03S),4E^A+9@4@F$FPO4U?R2W0
PJ [,E\[KC4_:"A<GQ \O79Z\,()&O?XPI<UGM((B/F16Z)/'Q]7Y,),? LS?S5P/
P?QW8<7(WYETQS7][O&#O[D)PS!#!'U=X)R284217F*FS6VTU] 1CR>5EZP1O=4MB
P<:P>L][\LTK)1EA;6.&*B.O(!'V*$M/M-K"_RL:X 6T.[',V$H&TW,&@ D$8Z*#[
P/;D6"-FW\%<<F.721WAHUXRI4M,=@W;.;0=86_4,&' *L+47EY"_8;UT89"":A11
PU$3TZ(M]U)B\ ;1 >&AIF> WX-@%:K:&*Y.;7>) >%+4NYM2Q+/2[I/%_!(PCEE[
PH[26KC1R;D.?PSQGI8*4"=(WOE%@F,!*N&NZJPWHE2[&C<F/I0YI;%+Z)8]3VNY3
PQ+Z';IN^!]#U?KD#IG%1/$N9A)T..1=RF)F9:_("KF[K]SUTA$UDLTGK,OIN[ YE
PU2AEC4\;B)"W^2"+\;WX7R'YL=FB'C6T52.1&(YL94>>-$X!O!XTY_P,2+CQ 5X3
P?85Q/CU-8H1V-5<,;%F0YR$R$BS'OU6^WYZ6"%E#MV*4!+@3'G[<\ONS@=.%MF%(
PA#J'&KB/(82&%9VF^XQS%&^-0?0J)7"0\0=>Q/?,;/N>=UN91(?+=/T&+HFLD-TH
PCF>*[0>B&DB'@V0;!]!V0W$P-U>S0<CGM^!4VP721;-]B&32:T!T'#PH\4M+>>!<
PFY91!=AZ)OZ#%F+-N\1JO>UK.ZFYR<AYCU:D[(9]YO5Y4/5I 3@#_=CVVR+31@GW
P959!7P';N6)30_0[_WZ,;D9,Q%>0*8:21#,GDTN&1.:24QQ#4^ $.Q.!P,U1H:T7
PZJ)NSYDH%EQHL=^*?GQ57B?]58?YTX:TRJ*]-GL7N@ORT.YN5TA2(!K<"U"=:;\)
P^ZVV$[UW[OP(D2H.4AIEQZJ"RKBNX>*3KD#N!AQZ52_\OG2J WH07? ORT,:-.]*
P&8:Y] SW&,AMD4R\Q;47D"8C+T\&:ZDF<3-8ILL9\#*0%]GA7L4'2[NE\8BNI.5A
PT:[?' 8C-#3MZ?,_L;\^3A+JL>P4I9%/?1@EGU_\(=ZX)4JMPY0X'["Y8EQ*&8"P
P4N'#^XF.6@O+/JF6-5XZI*T-YEX1_/4;$IX F"_:H@B7/*$"$%VG3.UVH"D^<'Y=
PJ1SH0M53HJZ,2^BQ]1N[YD>W/'!I;J_C4$.:,K_2&^)@G,Z:P#H,'Q"4SS9%;J5>
P,_Q]Z8?12$E[N&C'=>>N@DDRS #Z= 9'*?J?N!&F@=>M2G.I^]S#W%4Q:TJ5KUK)
PW-7,1LQ:[)C^&,K6#O)-:PN:G/*-D=CR ZFO8"&3"\JKQW0 SK4;/%K;OLH!_!W3
PN2(.>TU[$HMX=*GA(2.GW<12__%QS/ 5#:)K+"P&><V:U.U!+$E^_ZMU3>7KJ.>V
PV)0>-T(/_&T>ENT5UR2TW_]P G/0%%Z6G"=;I1XX]CQ/7TNW&3[I8.NFO755 MV;
P%-&8!FW0='>WJMOYG/3[#:.5XD>A-ZW^)MZ0#F41WW++7^<^ZX'?I"J(S2D0E=X&
P1HK[\)%H@Z.C7X[ .7)UE92V*J DN?5OD53U"]IGBC_BJFS./>PS4DM;=5*5&#N:
PK/0(Z\7;8PNL4&&-;$QG"!'R$Z+OH;\')$+)S@S+H5X4@U=97S@/\!NG26[K^?@G
P-#P81N2D<'] S^#A.&8 U=GE==,YFO-*DT^ BL>^'X3\7:>2VQ>4%04(L*['Y6GY
P6;(F^$)T>==>-0,^+/'4"#,D"G3?, %2*3F<T-4/. 4=4Y!19IUU;8+F^&$)X1)F
PKE/!QW%;8&'?UH$$49-"'ON04IUC1/>QG=_T3P5MF*+53>+7S!H,P"+R@Y];ZW(\
P%PR[/EW%#L*F+A*MU+XH3&5GDGHR?W0M^GF#<8C*9\DC2>$-Z4U].QU]U1!'?_5_
P&7WL,]UYF[*07@8?D/Y>7\Y*3T0 ?Y2PK,_HTGU+,KCN^BFRYRM,*8#%%;V[1._Z
PP\&W7*Y1&YB/CEY "AUN_@_AMLM35!L=<A(@&7*OU$ZB_B>E&/7S2&O9Z@E@.%?G
P]Y#3-.K)=Z3'S' ,YP>JE'?(.#!%D/<:6I'Z#LL#HY?\,DU_,>'!C1..'[PEC4AG
PL4*LMB4(\,4W=%_TI$Z*[B\$8E@KKT<<__2-$H\*=EA?20EK=%EZ\4$35$^N+#U4
`endprotected128

////////////////////////////////////////////////////////////////////////////////////////////////////////////


`protected128
P?+)9#"+V.E$ANY.BG)2PC,U'S:"!PR:&P@-%,4ORO>KE-_ER#,[G>X 5&#C5I#RB
P<U&'.)_0]K&.#XQU=.-A)NFY *IV#GK*E4"@X5!Z_QRGQ\ITK*^<WY8EEK2?\6%&
P:;ZU'$N^PW)*QE&H1.RDAQ4U1<G1V@:H\"U%/:(1A_TKN<#;MV 14S5D=8+#)==%
P^[:;+97DA.PMLFT%K!):L/C.NCQ@%^R&8#A,R#J85W([0T\:#9(Z-?AIM4H]I/]0
PVD/I24&,O84" =3[N),S")QP@X''Q-C%;:5)?>.)DP?237_VGBP*K:L"5)J:L[?N
P8,XZ&/-\'2J'_V?3O0)HLZ\&!PJN.FQ/E8X-_,85UG10GE?"HL EW$D*<,9#"D0\
P.<IZJF ]DP!>LOBW<BSEH$E0<N]\$3(P/(A9E,\2WC@G#W7%$&(J #E95?2R"_<4
PWO2PJ==)[<+^,,XTQ3GBE"$ C KY%A^ETY=AO&;UVTW$CHJ4V9J=CLKH=6?8/Z2E
P<%<_36O8JUATSCQ:"#%2TB-3?]DNE2\N__.O] *^0NU!U6.QC!6PL;@>HYHY!#F]
PBG/-J %GFGZ8/905)1$\CI4SA0\Y.R-DN_=BDCPO.M4B7(@ >L4RI[IQ[@]_JFRW
PXR.=\D6FW&KZ!8 *#(O-#/^:RSRL7A X;0"_".1O,KWYV>A*8"EW321"[Q=I324M
P6/+EB5"7N0<R\^K<^[0ZFTQP^@E56K_HV'>AC)R\"-.>GL$CE'2FF&SBO?$/IYWF
PL[PF#Z$\P(?-?C<C\BV+)>+OA:LJ&[5G2Y27RQC/VZ*;XTIJE<#*K85]HQD>=%X&
PQ$_W*V*HH6*(9519VJB;!U44Y4I*;P OD)LZ5K[BQLSI49:G"NT^?&J+_K\4FS?T
PI&R9Q)UF'"&Q>\5@,,L,5NC<"^('FBKN;) <6YA@*,,'#75B<Q&ERV@^$,U< ZK:
P]I=8I2'R@0/L"W#=;PI=LD(T7,#&;$0_,5NEVL9\G[*1W-(734>HDS2>%@2[ ?0R
P"&4IWD4-"=XCWDHX>\QMW,ZKGL!?FX=XW/E34C1P3VH?3PO'8O(^7._=YF5GU"=(
P3VW^4/?I<^B4I4,GR*N5E\RFOV 7%%B2,+M+6HPD"#W"W !%)(^*)-%4DY:-Y*VQ
P8<]DW='.5L#.'&=)PWPSI,!9B47J>,5Q7[GWO^<K;BAA-'"(GO-J>M =)C)]9Z5L
P<]I9=%*+Z<5RM9."<K'/!BAG33@Y*"N!TB5='FH_K_IH.[1'"QL07DK_&\NK6\<5
P.60@5D' APVU1.PGN@#>8(-6BHP(L '<%U_&=C6(@$#%F]"'/F:  WPY= A>[KUG
P),;7IP=:=686>#?L']YST\T="1F]-A/@J&+7#ZGJM@E2VW,X^1ONT5;Z<=9P9]) 
PU=&YT$7!O%6HY7)0)P"=:_&>?F5J53H,HX+G7&%9D>XC&G@B[SN6P?\XF<> 1)$H
P8Q*!U@SUH(*^VJZ7XTS>G'DO$7!+6._\-_2!8;T8)RK8&L:<1S!PD3MC9*"4@,^T
P\4Z'B<-N2[%35H WE^%S=V[0=#Z:0_(*#G)+9(6)VE.TF\3^#PABX-**"*D1H5Z1
P!_8FF#4S9\QD?(E8P'V^0A4=TM0^.TFF=%8S=_ML)4D[A_\*HEGP?_2^JO>V32'C
P3S<O_HYG:""FK*_E(^<M(-1/&?TB[;SS%4@J'G[R%W.7LUZ?P/D9>]OK;CS;4NMH
P"^S!HWNY8V_WA3Y%X_ YM0J''-8OV?E"<:6$I9FFPR*H3CQ@DBP[D5X_1CHCF /6
P^2T")(=LA2OM6#RD[\6(M!B6Y'=;W0G'W7-29CT,9^YJO72^:>3"X=1)38(,81 2
P3[L)>O+SD.'?>5#^GC9)&@DS\N.XJ0&^S&NHZN<F[&A[S:D9LK+9!DRJ#H-2 #;R
PBFXWP%2JXK?2ZT.9&4P@2X.-K]7EC;3)QIC!//45Y.\4(M'6]@_P:/3?0%LZOB;!
P[M!>G^T\24XPXZV"MW&O8(0$B4,6AI_Z!_2N#XMK %RJ"""UU;I_==IGHPMZ.-'L
P[2S>;*JP?I8MOPEXG^ZB9.@O!PC/;5?G(\;O;3[TECNT8-"%WBCB!%H[1?]"%283
P/%6GF"YQU2V:+4&A;DA/ F_X(M,:PH]45CG'N]<IGI &C)\X;F;&>!O)W%.8=TZG
P.Z<<\S>YUK6E_TZ?@6GJZ.CH3J:>X.&+@9E^$AC%H9-SB=RWX?<L2J#)S?H:(EF2
PS_" @Y8E#-X#YMFK$ %(4N;>*@(P;N6E*A[[W<U5RU_)$$<Q4#3Y>U]!Q-P@8]DX
PS!7ODPN.7IEF-S]_4PF(F6_1E-_>PILVW9)F D$>"A&:,%UGH/% I@-_^B5;%-V1
P^C\E9QGH%//."2^+YUU&QIWNTR)C_4D0C"-;;M2<E6'MBI;]N2=.I'HS?F"U_!4!
PH?$MWESB#H\AIWH@;YPAD,V!EKA]18M,R\OSBF]J*DAI&JBZSG$:K_\K*6._A]$+
P/U^;0\)&CM'"U/64:"BE)[G_+U>G>QY.>KE)C#S>M@GZ_EN3O^%1[0H(IM^1?F/0
P6]<3B-H6B',8P1(J9*<A9/2OV7 G-L+='1T+S7;X.8')_.8K:]BP_I0JV1XKT%]6
PW1Q+#4;KKIEB%'NVAX,X;<[0)<G^F#F8U9O)&:N[*DW?3;$1FJC0%@!<(%\S:^IQ
P8S$?7HMH&NV 9H8.S59.'="U&DCI2K([-K2-Y!:^%C83A80%*N.7V)JAT K-R'%7
P#K' D,!OUNA+*7A&*:K.+!&8KZ03E_F>!9,M24F0=RVSS5/D0D@Y\='='%;0-[);
P&'(_S1PS)>I^U@&&2M@;6=))N;_U9IZ25^J[B33>CSN $3;#.AA*1EHSL_(,^G@J
P<)'-+M4F7Z1]H.C;,0M&%*ZRF%*2##O%84*05680>US&S4-61@3U1Z:;*$H!M:CW
PBI4S%2H"@-J6$Q4F=Z<O7IF(:I4J.^XPP(L5OSS$Q%$<Q#0T<$QYGXE5"X(*T]]X
P<S-=(^U&=Y< -9+82J<.EL5QI^\8I9":;Y(C""TF8Z2G_U660]W>?-KH&,+QS&P3
P&(<<E@HY0<,3H$H,J_SQVX;Y2I17F\0.3$&U'DU=X"KL_WD_R._P V8,H;,(D4;0
PIT=59$$%-SQ40'A[P=O8]3.?+2JPQM'UK:.JGBGX_#6EP3N:+Z,77.1JW\KI5Z%!
PO"V@-1K=].DIL.O];9?<&T7V;[G@S&V#!IB(FJTFD&+?0!%569J>L?;UN+<1EQ D
PUQ%:POW0'22!2 *,(81^K<]J<%)&L82P.,X/KZ&5A<R.,%Q+/DN>-HI^L[-6, 0M
P\V)ZCC;V^L#2PFQ?Z#TU<&8D<%VL 7H]"HX8Y7S<>'>.LJ/:!0F5845V#?:6%O[H
PEZY$<>+=\G8((.*U$4)AL\]*!J%XP:K)Z6[6E[;:6.[XGXB]X(W^QJ+T/AD@<8H2
PQ0UTB@3"/,$;P85K754AI;HMZ.KNL"8^TYVG7%_S'(Z"Z^@WH!6[8A_X!9>WT<^D
P(<2XZXKE/[XC/9:T&;P,\YY>W8@4_]_.0G>)LC4:V>%5'(GRH!M_PAI'QI%!YX[#
PL]I1:!Z7-25,XS0ED;*&6F@( )E[KT#O>C<\/4_HB;-D?-\R9%4^XHL$^H4@4#A&
PRPB3(@J)1/#Y\QH%^W@D$Z1C!=T=M2;2V,&JU7\+-5OEZR7QPHQ7@5'$-7Q6/PH]
PDD$!%T<3L@4/:"[$Z3=$<]F3T\BZTJ5H\7*9I2/MU 1R>/$E)PZIQ,F%]VUL(R*6
PE\G2.=+!3T$:7)B&P*$F=Y#+G_,6^Y\))$@1W@31]O=ZW(ZZN4]%BCGTJ<![N5NU
PDRM.G+YG3X]UIE6"JUPQ4U*09SM&B)-Z:*-.A]$9E-38A?K,-MQ?#%QLQ9IA(IFL
P]CI;<CJK!W7/WWPK'5+:;W"5D;F\L'F630<S:;IV$_U<\*3*RTRYU%(TF6!OJ<J&
P(&WX:S1XQ'U/IGJ(I"I%%4WW[[9,NTX[6&#0*=$%=(6#B0[<7=YV!MLR1+=F$ELZ
PM3F^B ;B6,X:Z-6B1))O#\T>CW80&_ QY,7F-5BV9WA%)J-OD K0ZZ?K62 ;\325
PAQ.OYYO7QB'+4@]</9"T&[HF1]&[2=UVXN !8<&K;KB2S/'[26K31TKHWG<K/PE>
P"YUG[H3;NF\>0RK"N$XP H?JUGM.1>P"Z=. MX9T3."-P.>YL9/J+R,"M,8G4Z$4
P*M*,FA%9J:U DYS1&))_]5421QZ2EGWXF.0NS5W.MA5 H $=*"".%#=6:-E4X&]P
P8'[A].:T;E,*B^;3RD22ZKHMNK>=S>=@@M#!I(@A'P*TM+Y6\S.KQ');EQ62;;X 
P;*TD-WCK@>2B;8AI-\6OO $T8(R#/,CY$XSKRB<EXC&Z=O$LP7[Z'C>6T+QY3251
P.EX3C5I)#K%:UJTQS"5F8? 6>"N+ ,'1=BFFZ,2WJ1D[S2%^:,$-]_57)"H]<+I6
P@$S 7/WK$\U*F?Y1Z"M0*(A0T_1X1 (PJ2#,=NO5Q,I.1\_8!>%UF +W'!G0=QZ!
P5^XF1X**R)?GW:L/SL72W^MQCTPYI)8/6Z4('O"_5388M-LV$J6?)!]2("R I9D'
P25@T0.: AMD:_B1M:$&\#FI#1NUVXP!D:2\CFY:XVYJ;]U #W>F]( QOR&A=#DBM
P;;O88SMO.(?Y( ZL@0UN;@+/S'AKDP(=/#VGS[?8#(08G>C+9%)\\*J+4U"360E6
P.9R[Z"UJ1E=*"+^C^X6]=OXD;J?>:%5ZZACR[47+;57I&Q3ODNX).??IY4Q8:3"\
P"HH!M!3,'I+>X$0U"0UZE[@W-22Y#-"7##P$_1_!9%*!>,DG)(M:ZP*1'>,?@DMR
P!71UASQ4MBSH+<GO7$6#D)XB (+<:B8T2V>871^0O44B*Q&]O?X-&_0E2+531\C^
PSF9"5RT>]%PCSW]$O9BMS+?V][M3TFGT=1MCORTC[D*?[!,2P/9V6PVZMJ6_.K3>
PVHSWHT2,D6Z3Y-AMK@ZM :\L7,\A&)XP4[^>(JB^XIZ:57AFAG4*VJ_-38P1ES6:
P-;,J*")C"B*TT'V1UY 2TI*4'U[.[$(41N6]A:$R7*?\\&6+*/9/@KK.V]=AA0U,
PY)H"6N\Q=E*ENR2';XL8DN3_]'^Q__M3D*\Z=]7W?I[<1*(SUL.0B%8K.7!*=4M[
P^F%4<&G@J=Y)VK#=DK/#3]'*^7ZYN&TFU>N VM.=PR4Y-D9<MXEP4V#I>(:\T($B
PF) 9#4'+%*X<V,-)215 4R:P0J:V+QF=*+D(1%\7@,CD/U(BA15'[67W>DUM<V.V
P\D#\"7%9G=./$$N%OM.CXTK!BBS&1#R;-7 5[II +O(!,W.)CF&\Q2N+?/@%#*YZ
PQUFH\7O1@\B%6!K,U)LETW*O+K/&SE8)#*/*&^ZA28TZ,=T(EJ)SEUEHV9QX$UW@
P#P^@5=[3B3J-#AJTLCO)PF=:D%'4$1.)E^'@1>S'N;F%41MWI='/'"$_)S \W%!'
P(X[]ALRG==-&Q;@QYYXN:&*WP*Z>?(++NM*YY1HHPHO2#B\UB9?;?UWMF]AI<\;:
P",&WB)51C\B](#'2S]1B=OT2NRD>L_*4'14Q$CS8C2^EN'T>)P!S<%WZ X\+I6O:
P#[V&\*%AC ,R0M );+IR'3M#_@9F+%Z=-,TBAP-!ZBPN?Y.R;BZYHCB*W JY2NJG
P8QO7BLZG"R=7?CV-<M[59?([)3V[9(K/?'[W20=QB8MC2K0'>N /)\NH>'HF7I$J
P#5D539/;<TW8K#^;JI-Q!OU,#TD_T0IVCMO !"\'[V+_CLD2K8??I9P"/MBB9!RG
PTJY71\S<DD!A*&SU)F:34T%T!G"=I_[&U<YS]AYX6R<TM&OA:W2GF+'AF6KAX%VT
P _@YVV0LKXI9V701=[2X5Y&Y"&:<><%V$D*'W'\:1BJ0KW- AH<J(</%(@-7IC '
P>@D,>T?SY^:G3G,F5^]DTGF(U>_N'C)I=5LC&+Z22'K&8N"]%?#@BKQ$JTYS\2,7
PF2E[)PC=[=3(%JQ%#9OG5GQD6V2=5Q0=D9":#\9@T>C18VZMIO'GVM@1;5 :ZPL5
PY- I#")].2W2!N+/,?L&W)%"XDGPV*4A!N2/;J?)XD5>HMJH\J7EB&TDR4T7AW%=
P\(;-FW;=R24M(QF^PBV=BT.CXJ/OZ2>ANG!'A<NH.-P,<:K@A9[5@7 6#?DJ%/#M
P$VV<-NEGJC07.X)2/ELIO'AX?]#_+E*^G'!?O<@.72$$^2]&S<C0#*R8N:"+*5_6
P3F?-7UB;^6\78EW)B#9&$D^K9:RRSE%"$1@V"K"LOWL--N*L?NM83*]?IIO'I5FO
P7?L*BEK[^N%IABUK_I1W=7H2N2=)K+=;-%%1> (%<82Y:<D@L^6@= D:^U@AYDB'
PLW;CFWT\>K:-5[:1@O_51<0!L\LRD?2^U]2^=E.)L@"$0S.Q@1FF@30K0&FA,>+O
PQ^O\+,Y?9Z-1];^ ?YF-,Q;7A8V50F&*4H_ZC+*N@0\((1Z?U[,E>$]4'^/&V>18
P4'FKO./R8"[:3J;IV=D$MBAU,4*P#)33:SY9,UD/$YTL9Z/F+TN@6Q-IM$<(#3B$
P_]V!$?$L$E#:4\,!!S$,N:8,Z:=['O,RA&I2CL8S[7WH5DE9F#](=&>;LM7<2N91
P[7N9 FHZIJA<<>H43+3%X])+M]3%3.0*!FJ#%=\>G5Q U &BSGFJ7IMY#T_;<(FW
P)=<RV>IH/\V2XG"!/@$&W*TWQ8U?95?:46MY+HQ4-,T6$>$"*^QWHH*#.W1N5:;J
`endprotected128

////////////////////////////////////////////////////////////////////////////////////////////////////////////


`protected128
P?+)9#"+V.E$ANY.BG)2PC,U'S:"!PR:&P@-%,4ORO>KE-_ER#,[G>X 5&#C5I#RB
P<U&'.)_0]K&.#XQU=.-A)NFY *IV#GK*E4"@X5!Z_QRQZN0E,EOLUB4? !?A@M<%
P3%6U^OLS_0*X0A'ZR*T;8.-+R.?>&S]'+GJ)^+W6S4 '!U0L?V.G6X6E_SM&*L.$
PZB^YK1"PHW#CAYWF?56X(]]J/@B6J0X9!;_0.D2K=!-_QXT"!U681D5@(Q8V='8"
P=VSM,PVT#7//L%= !J?0I.C/CV649*6,I8OW(]@^"PN=*(7(/;5B<$@!&\K.N+AD
P(3YH']1,UL=S>JVI7<6%L7VR1\;=HHO1MV.#*]FEHHD2KVIS98P3DYU;^#@WS0B?
PL-12,:\%'<N?61,W03_1C[:H4Z?ZJDDVPK,99YMTBO5!W9S38E'MR*J*"(2KIJO\
PM7/QE$BGHCTH1<:\M\V7ZW$(OT@&JY@HHW(G7CO?;R1O_MK-;O<%ZR.BHN[R*NV7
PND@IZ5P*2B<.09Z?IEP&;(.XS*#\(:Q^ORZ%EK)$G:B<3%Y>W:W@CKM6UB82U.^1
P922&[FG.&;9411"+[;TVBDVE36-:A[9.65INQKI:4VUTTS=F\R.80W!.PE[7V,CC
P$N73K>D0A,**0VNNI!SAWZZJG3VVNLK#8Z*TAG/9BJ$<%ZJ_923*"@C =/;U>**0
PP O(R(72@326!SD"SU O/%P8S_00YG=S%9:W[@0(UPS452@O.?YGXA#*HJTR;/S"
P2O:)GS$5($T1R6H4(\^(L_C .KL&N8,/9@ F=VFUDZ<(XAW-6CW:RT4E /?+3^JO
PK6@4USL-%FL9*J#C^_R_;H%^?Z)J]4N#1"NRE.;'@[O[22936$)X#1!/_:3;"WM=
P+*HMT?YSM2_@ W4.46;,!I$EB-+TQ1G]A1]H).OI)3#FDQU&)85>4TNX[E4H[:Y[
P%]QZB8Q$4P@[FKEN-3C.DY'5J;UR%!0-G7A'ZQR+[I@Q0P/!2;T*/^0+(3AF?F(M
P?200"K938QC,;9B"R]&LWC?5T+>I;SRT)-A4>]D#57P[22Y$6>5Y_GA_5%"2O58Z
P#,L ?&"-V'5V)SG3P/CH"/@QL/^:FRT3VHGT<:0JJ2HE8>Q49)_98J^Q-AHMHIB9
PJ23&D4Q_-8XDTG*8?>+)Y4,2FYR._0WI'_>M)=P%E7]9M<%:\S8>7 ,.:@"N-:A^
PIK^2C3R:!Z]!?D*:6LE(I+79>*KFMY RETSL2C0FS4TS,6PK=>P+6= YD$)\X!-I
PV@(R+&7YAJ:\63TTE2'"Q0^!DFA*#-,*4H1T<K3= '#Z,X9;P6J<OM@"WI5EOG(X
PNJ2>8723K0@!T[5+2;Z<<];?T<S@_035%#EK\=;9>^J@*TE!T^%7 M&U\D+JK8%Z
P+-4J"F'CIY_@?2Y$D;WDX72 38LRSE[$3EN.])%SK?,QAC@37B=[&989!@W-0W7F
PKD-,0F9;_V.0FF#IL!A!N4$VS.W >S7H@61O+C.Y9^NNM=J2^C]SZ:QN@-+95:_#
P"]I1UE5!A'8.%NZ7$^;]$^?*^KJPH#]1A'5%I-2\6/MN/ZTGT:W>0<2OX1L5OP0,
PCCD= 1R*]-)+'M@M9$0BYEQB *]F:4N7U'/LCNC<8>!Q K:>=*NZL&J.VSU0-9EX
P>FMO<S1 ^&G>7,&L3CZVD\]H9Y":X6)[E*4M7EW+1F[=H-//=5F_;]!9!YD699K$
P3N#6N?^NL4NU#@E 4^@FHL'(#&J9(^=V:F3$A2*MAKF<B+-2)%^6G+%+97G>$^2D
PNJR-W_.*(-&X'C!YH,]PM*T@;A.FC&F6!TF5_KR*(WZFF%(D0V+]H*#U<5/*B6VP
P!YF+TL=!'*;5=><SF,>7^L"FP2:4,/(.AI5GLYDMG\1T!]Y::(;5/]W=&YT_P7U_
P5U#1S.<$[^2)[&>0.32]MZRQWJ]S'2U)N &]R1$M.S&]4F%G0I^**]G:-\=$EWF0
PC)8]&>KZFAIXVW&DB.V%/WAIOU@@[5MY,4/."NLW?JN@V<MZVP/R.P6W&:L$QQOH
PULFZ]P8*77E^";ND+/E%YAK W5:&#E3V@;%R0@-D'%1J'K9]PR<JFVT+Z(Q,E+E?
P;D4\W/K#]B#E^/4;,LUL[QR\P!X9;]B5!=2![#[5*+)8G*6<]X=!+S)2---:\TS7
P6%!][C!I+YY$6J6M'E5&ZN8(X:4&9WC^+X:9,VTV(L!G*YCH)_(><&\@TT#>LKH/
PN>E>'/^H.]]0F\((_+A8 _819[:VGD4:>Z0BJS:ILW_E.J9.RW$81*2BY;$,EDF;
P]'VRIZ0IGIW8=:*9#-YD*^O!R%\L\!\KD9JQ<..7HK*];XAFE+"$;7R*3*(&DI?Z
P>EU-]@@*042BAC/OVS/9SREA@N7-"J'-B55Y!@#0I]@[+)\[A-Q$YS[+;L 5Q<3J
PW?\YF)Q 4'8W\S)W<(;0$9H']<C0X:RL$+)M<E:]B703HT-R3)5>OV:BB3'D)4>4
P-5(HNM.N*0RN\^D]5D-N-:.CU\\,"_SILKKBX><+<6SG7X"3.P\H";?BRWV>0J[D
P9K'D2+O_5*TB>E'F#%5FP779D(,ENS5&_(-L!C-_G\RR>>ZDX0?EN#DP2MOD)BZ8
P\.>6WSP%UB_'IHIB P\A,DJUN,8RI-"BK0SEI/IQ!QB7\!O<<-"^[WF-OC%U*DNS
P1NT5X1:ZCG(O?!41DKM8UY<I8;3$Z<D4!>K9&?LP99MF-Y2J>4E1L?>1*L_6G"HI
P-!OXJH/>H24:RYK\W[;N!H6"EWW:T;MR9ZOZ2B.^4UCXZS\!S]-B9DB(.D[\(A@G
P[LWB/B7P]A)R+F/Z\%+Y=4,,3<:ZR6:EQ_(8PB!V[4!RQ+1+E40*X#^DKP(&LCS&
PY<S/$UC"%MOP$W5LWUUYK<($BLY$+N;QK"BFS%^9H#YSB<P5FT\/OM98@T:ZGBE\
P08;#T&"5V6^<K@ARD)Q?T"E5<(5C+.A3U^E?L1ZGYMO*UWA/0_*36_6D;-[6IB$M
PZWYM#?'OK2K ',ND8O6& &(L:_FXU3M+MXMVIJ?_7O*O/=3(7Z(UFJ= P5 2(=&W
`endprotected128

////////////////////////////////////////////////////////////////////////////////////////////////////////////


`protected128
P?+)9#"+V.E$ANY.BG)2PC,U'S:"!PR:&P@-%,4ORO>KE-_ER#,[G>X 5&#C5I#RB
P<U&'.)_0]K&.#XQU=.-A)IW)]]5]3BUW);.#'Q4MA_&)QNOP:XFE"9?&<II?$[>L
PDOV>JEW8<;J;9?7ULGUF06'XM:AC;7O*I9?G#?8G8,59T1I"$Z)XNMD/BXV/!JRZ
P4R!]Y7N+D=W<'5A,A#US(I07YWNL &X7; L7-\UCU089_'&2#NZ3U(CXN&C?QK,4
P:S_BR7X!GF3(M@@,Z=Q16]X)GPBT!>NYWZ;50@"!L;W6[I"HT0W%[)!B.3$5TF0\
P"'J<F&O( ?&"#M,5G":=*=(2Y>[F"5 %LA 9-9M#B%A*8<+[H\9PB8RF?@!^/6+L
P7!6K#OA-X;("!J9D$8/UB%BD8;*7GTJ+,",Y36V?$1P=$]P3!%$2:A[YOBT7;!Q5
P[SGD.WPM1U:Q&;&J,G@WMC.%6)7B6,X.\FWA W&W3:D+2+TKT;I1'V'];EP;Z;\_
PH3W:<'6%']O(AT+-24>9>-$G!I,LA$M_@GK1 :)5I3F*!1?KI\5\CR,FD5-":G>\
P)U"J3#&TTON$FMM&,EOA181]VZY-7/"%RO?[[2%'HX7]!U9C YW,887_T2Z9,C4N
PR&L0,3+,;$Q9&YE/3HQFU?][-]NHCWA'_<\86PDATM%<H'%J-0_2?U%#&#0=$JH'
PF^5#'*0F,P6NFO.JSG(_8PKVHBJMJ2KFUYF:%6(PUGGD\Y-AR$("8>*X'NU*!O*L
P$:EBVA-.?XZK6PTT=CQ4_**_9'CO_:V6Z"L;0?P78QU#/4VI!CWI(VN^)=5:4B5!
P0?* WWY."^"FFM5H:S1#>S<*\>E65EGB7LS3]!E/=K7$P_L!6>'J"_?/# ((#N+&
PZT"X4:) @_.%CX?-_U8/4I>.M&: L[4W+SO%ABM#B<W")X\Y[$_VGH@D)&U!E%EK
P]^WKS>BSM%&B\F"OV(ME<GHL7UMBQ7SR,41K<DVZ@]GW<9GN1A*%H/B&2?VOHEYA
PE\D35?2//HS;L,WK%T HA5P;((19D0<WF\+LI:46+X6_978*RZP),'U8WE)D"J W
P<^:D912OEP_PRT>XSW8Y%V,3\E).7V(2^SE5:"5^<N_AN.N&WVKI&@&YL*G33(NE
PMH0XU<=O+4%2P<Q6<)]_T-FKYX5(#<&^;@7L3:SNZ!-0[PL#C^<K< IVEZ85<=]A
P7N@VL,XN6Y<<O$)T4_W=B04HK,XIKJY[G5WCU]82Z^X=+*[,4YG</'K3[]7U%31#
PXU--##MY5W&9/'D#L/FA5[A,UBR742]TO7G6X+N"_V^I[X@5>CS#$F(@C':_HV0,
P(E3;M$"@RH:?\$HX1Y?7\ Q\5]^9R^+&YTCM\;F]&6\06;:*/#MVEHY\A#Z-39?Z
PFF<JCZ$,0)=KU?TC.X^.#YC,DWN*H2DY&'),&_$(W]9;N_)][%O;Q,9S*^P-1<U5
PL=H\@J4>"."6D=N"SA_\3.#6O^3:>2Y1S(7==-\5Z::5^3]JM"5$&A(ON:OO(UIC
PPG]#T$B-3T=%58P*"]6Z-:7B)2?,X,S?+2A@UVD%LSWTPYG!6N^RFZ;YNS-2!4@^
PEB*VT!<_OU*KI4$$,U-C/@HQ,4#1Q(AZS.=M6X$0?\03IRI?YY7FR;X@<R@RV.&S
PL7[4HY&+C=JGP'ED,+]TNU?0B] =Q(^F\"3^\+*'?/))1CX85HH]Y(6EH?B<7[?8
PI5@4,_7H D5%SG/@$8LX[R"7\_0&XJG!ZN4J4\NR/'=9F/(G<BI'1O>%E1,'MUT+
PD@253MCR9W?0.U/1+ ,72+<,)LPS23E$N<+?]^D85VZUM\ZW&RB@,NG0(R516/IS
P$KGA?%>@VPZ=J&OO2?KM*?126@C?$I$^-4HYF9:5X*-\D=:K50;J//$[V"_GSE+9
P!7184JJ>]E\;^U:-2*\!)[>+4/K< WBC >&8VJZM35<)<D;Y59$3I)L=-P]F8'C*
PR@N",1M<H [SMCH/S+:.IK5:K V[3Y2/D1E8=#6D+N=MSMO:M\'38]H ]N9<NA["
P63V/0N^.U:=3:BQ$7VBJF^Z'*K1)O;= $\4K&]S^;H[-_8'))SWA*D,?.%51ULP!
P-N0F#!,HWL@SG%^=%S0XJYQ_RYFYE;V_R\<LWQ^%)J)8@+P@''N>+:8ZD_VC0:FL
P,_H.9)(<8BYPJ\_"PX9>CC JL35N[UX2;[(6R%LC.>+Z39RQ[I3@MT/4TAYE+Q9P
PFMGBAEF53/SE7A<4-4'5V%#UNK5A1"1)Q7J;M#TRK?D"R#(0WEDU#*[O91 >>DN.
PCT1Z P I"M%'Q@;F]#P( W]P^B9>KV8WM9TI%==6P_J54^AZ1:/@J]_DJP5QWXBP
P&#DA_^B2;J1Q?O(D8\B,1Y:31<"Y6P)P-,ZT!;S[29B/GW"* U0K*#TV0$>< MJL
PCD<Q^5?P_#LC$=;SX2JH,4%G)U!, M@#/W#;,)[/:-8:%@6^LCYR/S7%RBN.?'I[
P/'J5KL8S95I=?2>.\GG]8%,O$#IX*-1[7!OE"Q+$ZURR!G$*,,J)+QQ7>SR!E^=C
P@5IP[*"#I:JL;*8:$T8&$7': NE<^1VA<5;J5-3Q[2 H5;%RBT"2@)J..(">/K3H
P>.(#..AXIJ6A]O,'WRWDS>7!P<%9G3\S"3P3)3D$=XG=CW&QY7XKB<4R9 AU]T=2
P[*E#WD42G4LF6*7/.![N7#OJ)G09V/K-PT#*\W$BPMK9\$'JBQ>?H^S#_-ZG5BZW
P_"83!I9#EW"OVF*6 O)3Q'KRIWU!N2;[!^8-N18]?E>'D]TL0-E@U,7AUDZ-P" '
P!P=Z-+ NL6)&1(BPR"3$0;E):W4#7XL?"N!;@T2IJ4K/#;,T?4$ 6MM_6J,3/0''
PM&Z-J;JE'+85/#]E4@Q'3OZO<^V*OQXQSP@%[)RKKU^I__[__@2&2ZPNNF-9'M]Q
PP,)U4.8TQEK+02B4;DAOT)3 B1E8^SODN*[B'EDGTW%2YB<GH-J+.B^?T$N?<6=+
P6%EK),3/!?;\M])O+ %.J"_:%@N4J%?/@]."\I-4W/!=EMALCZ) 9#3%[PW)Z9.V
PK;.M%CT8F;^(6''>8-B/RT.XC'!-7G;BF@]8F<)+CN?1C@=6K;*BU2_2R^Q"OAF0
P/W3#G)#;[&9>6K:2AZS#LXZ3@^6Z%/#NFFS>)R[6H0](,[T*D9WFLXRJ(\=OS>PZ
PJW.^%=TSLIQEO*OA8;0$VAG$R?D;KB<?*G7W292B 9WX)NTTA0CPOVK;^_"A!"AE
P/\B+(<"LK,XDY!M,()G![G4(,"Q6[6RSGC"AJA??F2+G'0IY^8E7T/N'Y(-_SDI8
P#09 -GMXR= 67JJ=4D8"@5<:(HHP*^Y7XH"N;00+Z*#E>-VJC"H4Y*C(/2V\TSC.
P-GNX(N^_9"OO')E^>RK@-@$67VC0">B/6;:W93T@KU]2JT1#FO&VI@3B135]:KZY
P@'3\>)7]H*HX4,^26H)NTZE2F'].U6Q8'B(GN!/1+]SC+Z5R;EL: /Q[?-HX[].G
P"]:XQRPB7+Y<B 33#*,!(]Q,M=FS/],Z@1 =J>3>!\UQ\%%-0]2VHY.I0,DQZ\MZ
P35."$-_VO YB!R VT45)M-5!]+A1Y%CO=,=F-.6ANQHBD! -Y52]SW8][P@=+LAD
P>E<'QBAH*1N<8R#XC)Y]([#.4RJQ5!K+H/=R1?^<HY=ZP2GW,Q>V<"Y)+AU[LX4>
P@IMHDCFV6#*O&XY;9$+1RE!:F#@=J9>Z434;[.O^E[HRD6%?MVTHOB-)7JY.5Y$[
P#MH<;RI@ " (7/6N*?8.E^HDL]6VS4"1,N[X9CEZR!Z.$"S$X+ 29-=0,\GU'"U4
P7O,H0S \,8(CA0%3QA8Y'JUE5*,8, BM?;(EJQ&X(9N> YGCU_$CMN"U!HWH>!@*
P;W-#UD T%N&Q&#\9[7A8U3& 0IO57+=ZI@&2PYB^>$,^D2#(E46\,V-Z5THG8:/6
P^D^O=G6;;%.+;,1B^%Q$Q667M:7X;<A#NJ-^N%@V[D4G/8SIJIUU9@.R .),IY23
PHT5W.;"-V:BO  AO?AF NO9FBPE1_L.1\\.'+E-+:\YWG^:WP]W)I3\\7<GITVV1
P>_QV8<'[(1@&H$G"R+)PK92RRM[B H&1#LV/D^C&5PD]GCNNHK]^!ND6LJ_:!-W+
P$DR"87P%6*/W&U]JUL@C>N 7 H;  @N+268I_]'MXC'(58-#N^\M.MF-8(MM ?=!
P+\!_C%S'I7=Q#[3=:Q)8V_5FHJ*B@FF/F2XM09/BXJV,7K@R^C$;%W7*LUR"9XL1
P,*P3S.TM3FUN)OKT2U#V:39O;O#7HG:$OXH) L;'$8)>'-O*?AEI>/\V+4%'XQNO
P<>FECH$"W[ENH^\;C&B=899H;<_<(\0/"B_I%LG^8"NB5<:+M<X0# TZ9B*]4K35
P&IJJ',5H);@M?\1W)U<<83)(;:[?^:H4Q4!O.4A=&249LA//SF^FRHCX/(B@+_^$
P.^[Z_S*\LFDN#?@(MV"0'ZHF(^5^SLO\"QZVC8YY+^B_N[@?U% W%8!0"3?&F2O 
PG@85G3*+V^V)F9J$_K-_?WKRM/%QYAFXMGQ,C5S"&V2BN6*ZZ*;RX,^"2UAH;/*W
P,?(&\=@XS#L S0^,XY/!_VPBJQ>[E(H6-NM?3[X=:1_VB;V&.((#R'GV'?5%E=Q*
P3K%W#_-?L,C94U#X) >L%K<JZ :[6$(!<3Q'A.3E(S.6^HG %,F.^#VT'=*SH)"A
PH$WY"8O*/K#X3AK,X,6#M=@,YW6D>/7HD=5-(H&W2P=UX$^ZV)IQCXJN"5*8]4$A
PZN827%]"ZFGO8CK_(@QBS2) !0^M%7[\D'Z&UG-V04QVW5]4DB@!EA9=KMD'QR.Q
P[4Q6(<B/($5KX"J96Q6"X=A5RO-@*E; ]A@]2]'D$,B4F"7@.J7OFR#PNE&IV>G/
PPXDJQS\PE&+\KHR C78PO)^5U5AX2W70>_Z4MO_U*@'"I$2,%*89; 'GQS-?4[JA
P.R-EFL&# K:N__LG6GF:F 6Q CT_LU##ER!Q GX\O(?HUEKZL20H[2&<GM9B5FWY
P3@W9+=E+^'V N/NJ""L%6))]/2 ?>;K>FQ6X;&LP5(NSUS8_FNH*_57?H:#=X5V5
PTYSR%8=>/!IB-^#)%??>T4$R-M\"&6MW@7]86*N9C\ _H6,B@-A,FB@_^V'\2?K[
P'L0.Q/%$8LP^M4.!_17\A:NQQK+=H8[:UTEX3=YV\LTS&Q3&D;M=*Q+7,0PL4Q-4
P6KY.ZK@X*9J T4%$\F]22PE*/W.#XW3SDERG;6_NU?,5_6_*T\26JI-3#1@ 1O T
P&^P^W QOL%2E\?"'K9 *G0?A=HK;,B^PT8(G]/$:@II452/<3_B8M=D\B%L9LQ:&
P0>@5]B:4(/(0QAKPM:1TZZ8I'FO^4/QLJQ[8+L?@6&X&UC.6A>TTAM/&2,G&I+:@
PD)AI7'E:[(P ZCA@OGMVDNT)@* ;TD5)T''JC/.@*XG/?U>BNZ9.I6Q/[]MPB9'C
PB8SM-,&P)+=MHZLFO-2_H!Q-)F.[[ H(I(OSK6+/C(]#XM.L;,RJS(3VB4HE91/H
PG$R\,_55GOVOF+%FP'\=?L[,5*]IN)X@5VYDJ535)P@D;C91Q5LZ "%!#KIMN"8Y
P29$+/JRGH7X0%TJC'3MY:S-GJ</N-">\:*Z&WWQKEDCCF7K]"T-D5'>@;PP_\E[<
PF;;F+K^'SB?17M^*8O0)@;A0(^PS14@&2C7#L<F9JO_D0:D*=9>]!OY-ILU@X6M9
P=J7M!K[8JO-')%%!J?%<W%U\6:'001FM41('_WWGK<ZW_>;Q#NFY,;.AOZ\8E7V+
PVLW4/%_$B9@)&^]G\7Y?R%^O+Y!)"^12(!_7NI"S9N^H=88U'L&!"!4S2BJ/G=):
PJ(Q?&PA;\)-RN8]VJ5<M1:]6HL)W0E+EQW=88VT45S1S D><ODY,&,B2/:PTJ$4Q
P-LTH<M<K=P"-[FJQ.MW!PVL=K[/XNZ<#FVN:9F-V5X%Z5+6 <N:+5!IB*_7['=EM
P%$ABT0Q^$R+NKT/X2RJJG4XY60O+:>3A5GCPE[/[,M/J#WO9.)P+2[-O:[R#GE0C
PG;S-M?G2;0Y$6:(1K@Y=WF_I:)EVP:;BN98T[A4[4/\-_4DSR$\93@?V_>7'S1L$
POZL+P-+?3AA"%-$A2"J+(Z&HP6)LI/!=Y;2?J*7/C%=Q,S/+J1SCGKB^RWX%"Q$4
P"""V_4];"H!YA41^PVC'>'6E$;-Z#@B>YU!M&A8INWA?8Z6#I_W1?P.0(2$7%_+3
P 0D ?9-GXLEA6#+N!](#/60;P87*S^LZV/5_]$ DRBPY^4LO>\#:[:,&Y7-=+P_2
P#*P>-=TR'OPK@7S3HV?]Y'DD/8^* 8!TGQ/1-V0(L/L>U;+4]'Z7X7Q^E][60];#
P^7"W.5*]7']$$\PXN!8#7$'-O>H$OU=D;N54F--9&O#2Q,,ZUS.D).OJ/LX8)==1
P%_LCT$ PT ]EHE9;W_K O'/#O *+IL=Y*9C 4L&F2>]U:2I0AFF?/T-3D01* &,,
PJA2PNDA68=T1'$GV+M4/=*+3(BDO)<DNU39AE.WF><@Y0%J4\AO!DDCA5DB5JH_&
PR$>9B<21TXS/2<9.O-RIA@[W96"4E?5BBCKW0!]^N,^TH.-[5>A&Y&I2L,9&V1 \
PT+R4"),/7E7</3:X(<S;N51>T;L-Q!R=2M031:@G3_IM3%\@" M['D_OZ21)'.3D
P,(9-X5;2YW.6KK97TW%=X^A3\#>'YSEH]D)&/5+7@EB=Y&,V;D1G8XE.:]0;LTH*
P5UM/>ZTQ'7;CUC;)3'#P,'62FNC/#E$JP"@'UH+$< 55\0FW2!*!W4 L(,RLP)EX
P(2RC^6Q[TQ^Y:FI<C7)E"[&7Y/JG7@)7.HY[4\7,"V!NZZDV1>-;.!R:':!"XU,=
P,)%(._5W=(MFQ,!%=_-SML.'9"U;@</FL?+)IHJ+D.!0@]92OQ _E!QV$9>_#X_(
PN$9W=QVUUK/,QDWZ*P?[I8V1X+6YL89&AO024_7"9P_,A6Q)Y+XR<;M5XNOX7QK[
P W6A'QRQGO#D!.0F.!9Q]I#V[W IBOT0?//5J=(C,X+ ];2GFHW[<Y5I)J&(8(-5
PC_-B/QS2UB&_2 ,]:=]?B-VPY<T9 =Q!)A^ 9ZY05J@K_G3ZRE$$@!<@97NQ!ZP9
PC<$\_K389.9)O6!@>+P2@J1("T?Z64D%D:[;+;O&S_&>S- P?4 T?\E?,3DRR\2D
PYI6+MX99\3''RYP,4%\6S /H(J8N'T6?D5H]NS:PE\'*Y;TV\V0ON$V=/RE$YLOH
PM7D" ?)'YS7 ,T]0,^&" WEP/JO'/Z[-( 5IU-2BPN5(+_S;TSJO362D.^)T1S>4
PC\U<=5TLZ3/R_(XW)I4PT9MM^L-OB?.=FV/R(K,5E?5S':42^GK #5^HKF[8P:MM
PODHZ8J5M5+9\/7V-!2K(XGN8K,T=44V<7]WL/ +34?CL&<Q]K/42*WT_4<.E'EV.
PSQ_BG)]&5HG6PA_'0*>\]Q5BI_%N?"7K+3L $P/QNU\!DR-T.-D/!@X3D+#@GL$^
PZ ?:N^U;LRCXN0G\JM&UC3.<X64S!ZIM[17:*I(TS*\Q[LO4%5A;/KQC]=?,7B4M
P1R?,1!G]W[T_028@>[(W'K%[$AW*Z!%"8 6@.ZW"A%(]\7N;XU7S3:8CK0D 6X[Q
P16TK#]_.8M=:VA;FMHW\N+N*B0#6OI6<7)DA;[_!6?K3LT,+K:JTL/.E5"RZ.\!2
P!/X+;P,R-T[I0+?+%Z=0@^KMP66O5V-/A(&?C:2W/BMG>"I'Y]8JC:US&QM,:3#C
PF;%AEJV4D-O.*] XU'"N[3[!7PC&N'YLB4>;U(XNZ=.C42S<YN5BSE,^0W5<>>N8
P+0B_$9<8?:(5E![$?/W&%EPE4"\JQ1:.?A2[K0"&0"MM(?SO(998LYY; 45!7/R]
P)U!;3__BT2U]W@%72V\'5<L4!,Y)VGL,<DEJBLZ-E%NQ= ',@ .?O/D6(/$JQI/J
PN">0]N>^]O]_EK8KP91%?HD<(4@7D<=G$6,XS_6"1:*],+CLY0H ZRYS;T.'Q"95
PNV.',6R./^^?%_7I/\'U>?(RU]64<!ZQ".8\6CX(O?8L25N9GA#LYK?9DV0/Q[W%
P2[-"1%RV]G81(+S H5J6R$\T2#MMZ(E;'8)X]JE@.F/41(ZCS0J1Y[O?87(;\^[0
P!&+\\*YD\1<9?$^E(C, =6R/I!S<M&H</;]92^=8:14)'#SD[YVORRQ(?+/.YH$G
P5#2*+C,8Q[XN?3+BO9L&N $NU*W6 E)MP"N,["SBBWH@"A:UD](X!@X&-0OE'J;H
`endprotected128

////////////////////////////////////////////////////////////////////////////////////////////////////////////


`protected128
P?+)9#"+V.E$ANY.BG)2PC,U'S:"!PR:&P@-%,4ORO>KE-_ER#,[G>X 5&#C5I#RB
P7P%1OW</D*++,<>I>T3^CVG:>&B,YAQ J*H.)CCT@/HU+1Z8F2^-M^ORM&PC<YKQ
PW%<[[_-CMJX$+_&AY%KHR15,4$<]C_T?\;AV[\-V=,H4]_J6* 0!D!UW*>WY'[ <
P)/=JT4 IGN!550LX"U^")JRQ9(K4]MJ'?P4\V8-MSB)=D).M)EVT,C2*O*OW'E0?
PK8-EC5L0BW1JEL.87_OOZZ35F.9G%FFFYID*G!$[Y\T]Y %EO,W$]DWV.T844K)F
PL OJQ0VBJ+)75['.O-.3:@_C+FU-2GSG@OCI)<'?"O\#2E-00;J.+O*@:PCC%*BY
PC-G,R5HRKS[$YXJU "P1SR(4/$?%SN2C/D8/+G8 1U<NN>Y(*[N74J-[!UV:W=#N
PR) ;%?FRU\3CP9%'HL>XDG4781:+K$]8H%%4>P1;2)O*N-/? :>U5#-QA'AR4>)5
P*;RD%;<A[Z9A_X6WC\[BONZ3Q1].$<CCE"\]C2YZM*(2-:_!K$L".@TI55G1P&)X
P81AR/63\B^0&%%G4CW 7SDI#J%4 _/+O%XE*"'OM UVPR&688JUJ/N8B5PAP]2Q@
P0%&GW73]9\UO!0CE,*0N[1TM0+RB>"EDOF<4^1!4%6;MZF;6>F7!:>D&T+;T+E\X
P<U[4_;]9'7_H*.)!PBHPICB6(%#L4=F%!FB8@:SG_?C^]5CL;KG3X!@M@:24+D'9
P5L8@)=7MV]Q&*+$T2]\88%(/5E.(<,K82@>\(97F*O-[E<&+F&AR,,P O>9-D,M4
P(=@MKGMFS8U"WAF3C]2T!>QC0B*,M4"#! 1P&@I\'U"D=LVZI+7968<J<+FT)124
P*[*+!2Z985;.9ZK6TYPU_@$MBH#]V:"^1CHN+^]!,^BQH>ZX74 '#9A@7/QX/7B/
PA@019_F /A_-,.3K+SR0[](*>1/5(X07>)LS.FH3ULM!R%[768&&XSC:96L110\9
PQV%./BL66[[1B?%NX#9GP-+]<\IJU<C#?"7AF[VL]*F0DH\GNZRM: (24(MHU+2[
P)6VS^G4T4L;HI@[/6$:=C.:X%A<OT3W2091J@T7Z!Z_GXWW^'Q2/=SU7L&#KZ8+1
P:3PFF_7BJ/P:5?=>AWO/S+M)L 9%CV=OB G#M $P&)GBP'HLY!-OW2L7P:3T6_:H
P^:A]V/YLK/9O,+PT(FNNI8\0?7/E?C'=IS5#-Y!!I4[;P$N?BPOTJB:.<*@R7JX'
P(,TJZ]0$$+'?ZR0Z*NQ$]X=K@'F!G%,XRJ8NEZ:5JX\P<+\B!_"9XW#?6<^:V* U
PR\7])?@]@MNS8YMRV612. YPF*IE4&M (M$77XHET;N*=0(MNK3UEB6LIW2O'?T[
P_,?Q:X<'/<RIN:KK=P#W);)%/Y*FO9WPN!ST0?K&8N\?7&QXIO4K%U2^O@!A%OTG
P\P=..[.(EPMQ:F,8]>*+0%RQ8?EJL-\-</#]2=LGO;&-&Q!_XEED-ABHZ$H9!M&"
PG%5T5./ 8VNTC2=,V-[Z^FN<\;8PLR/4=7W!N"6N2P6],6^[6&_6!M("K#9K,#K0
PNJ@*>['_*)3@P%=IA!D%5D\=%/H;B09;E38E>(S6I<F$1X9 [%4,BO '9+KBADR+
P2,7L@%0)U0N;7^!ZH3MUINSXF(YU&5A9FO=7O$K@O<SJL2:G_C\7FF#-X-T<RX /
P2[3Y?!($H0+@"?-!C#^AT>]S<6N=P/P9=BX=U_XZAKZ:H?W(["_:_"U]<HMV0:(]
P ZIHDDR+@Z%[3!/:+O O8& CJYH3"F_.:14JW4ERYC^GD7F9,80O/&I)DS4#>+C7
PA+?YGV(,'[(\]%@)A_GLS1/_:ES::;D9$2O]TTDZ<O*9W!*"T*^J=\K@Q(YRY9]O
PX'@U>]]4R,O#U[TZY;I!=]8F6G>XOH_MH6E_";B9,/"=X"R\!_HT4CI7(&49"TNC
P)>R<(RC'&&Q&0"3,S386SRWD$ ]#KB\^I#.@O(R$W ZFUL<?%-NFEH)&:/V[R9BB
P\9A]IRQS=Z#JL_="?;UF.O<_#O18B>UTRK:.X-1\JW(IRM@AJN,,VUOD[HC#]T[L
P>6<+YL>)3*?@/LGW@R:CZ#U6 87H2]MUB<K*WC2ENX]LG!=09D.Y(PVVG_,+:MZ_
P=VS3"Q$]NK6+XPL9.K._Z<^J$5X+=NL%E  H[EO"("=G<J%5*E8S>GU'B?S?%"="
PRF;VX[6YQ #FAFW<Z746;=Z3#]-&91X#2-A%T'K!EEJ]JQDX>U%CB3?1TQ7N;E10
P"A%;-WL.I*LYO?PP].O#]$P]Q4 !-NZ)YBEF(VA<Y-2E2R#8SZ<3%S4W&1$2B]\G
P6@P:7V^55+0L1,T/C(</L";ZB,WV0LB:"74J_%.7EBVSR49%R4-L$JCDTH5@1/ ,
P+>G,+^$20/,^I'!3& $:IU:6?,MA=&G%3Q.K9+JE/(?%,@#"['PH; @;R\-%S6_(
P(38(R^"LL0,3O3_Q'DF[,):+ITF>-O:1#,^2$A<W,P^,+BA.M_*7M_#@ X"]+,8<
P771P_Q[^!!2*I[R54V?M6"PL>\07)/Q]>Q(9::WIV66%'(AZ5B.7DD&4;OIT)<<A
P5*O\ERM)'-C$DQ@5Y-O6:>YK9&#UTN-[N^K-+(MHP_;DB[[!>T #(P]IZI+!. NY
P0^&3OVWC3]L=@1WM$^Q#1H>46OW=EI*TZK<+PZ:6U_BTNZ:YA-?W:J+Y[6V_BD]A
P2$#^6(%9GTT+";&;TG<2B.:XL_-+5M)U70Q!ZY8 3>*8%R)J]%U[P*?XA*H!ZE0&
PHM!4_[YM&IR2FG3)Z-K#O OEQ9_9*3K,T7W*QK49W>"O5?1,3D\0.V(4Y36G[:JD
P;"OK09A10[X921\E6"BE VT(K]<:?M\V1_M4&8!FV I:3\@Q1&8P&5LU_R0FA]FJ
P<"*9(4@NWV&0-XEU';=&?Z$IDT3&*8&>>\).O=RL6$G7:J58A.(-'Y64@ $#VR12
P@$O+1YW("&</Q+G4GJ")%TC4YL[R))\FJZKS*IZN.S+,O-<.3U\QET;& XOX%=^H
P[D+R^H7L'2O,FL>GR^7(VY34?M /H:#>F.=GX'*M$B!'0$N8)9!MC 1KF3*3 Z"+
P%(R/,X"1 ]>3'VJ*ROO7HM$F;'D]*H')8M6K9"Z7#BF:T=W^Y#%W5IB]!CQV(=>O
P%A=)#1ER*'R=3C<)E66YB7"/F(8)+X0.%\$<C>D<S&(TJ7C7(P .FBG8>]ROM7X/
PS:;:T,$-\*YB?Q>Q_ 4,68 H7?V*CD[X,K_<J&6&FP=2MW>[2NTL Q$2O\4]J/J2
P+,$YL:T8*J5_RLSSBK$XY&G'KVIL<DY>#%P>:=1(/M[FCF?[FZ:RSI>#\<?(CM/B
P"NANU6S;<JC+F2#2:S2*!R([\ "# D>_".%E#C/[BI>#SZLT';C"*>.E&W^^,L7V
PZTMN]C1(&F0BQ@8MZ%JL^[H@YD1UW]7(-F*^3;RN':<^ )]&.G 34DNEJI(M+E$X
P/05(Y'W_%WFX$Z?#R;_]&.)H4X[(;)OL/5Y*0O&*'^[9R3N5DQK%,1V9N"&(4E4C
PTND 5+YZEIJZ&\QV'-Z&?0GXMVHH)V%<3(K*,NY[B5\'IN+1,7Q<HZX_^]TJTP4Z
P^"N/D60M^EDMH(T<9*!:-V],+ 6/RP)?B/%%']/GCAB-Q8$\US-6L2$RQ;8>HDF!
P^H!:[W/&_F=M;;$2*WJ.ZVT1V(:LM+4V-)K@I<4+FG1O/O@:D_ZX\!&INU.IBZ4F
P3Z Z?,9)+G0O,:&B1B1U' 0*6\YI(O_'+OB-I,$Q0KBRI:LQ:D/!Q(74?^</DY0$
P#6+0=T]]R^2J= !$D!KNP=']\0-M!NV;EE.<0GRU$7$9M"PO!CLZ-)95O P@HR8;
P,8SA;!MIJK7MG^AYD%X]R'WT.1IX0F6>_I,,::>G IB_6U4NZF I6R.>GP>W4V)$
P'GU7%9\DT["P67M&3PQW',\,(R<@I/0\<[_^_H2-,AB!:D3J@7L9((0E[YF^GL.;
P!V!"))_84]L>5$8)\+Q@1]1 9WJ!@U&=6]_#MQ4S[52&<+,MH#,V%*7*P@!([SU&
PQ+)U&FN)@/[\\1S+AZO""V7R.5U^6L=\%I:!&V;TR+WX%QNS<.?G*TPU\#OUJ>8Q
P%QV_JROET;,&04(=9D \$YH4%]VLK982J57Z"%QKR30]?X'$I>[KD ?-R-WSH(_Y
P3YR"9(T(N;*N\B_GHH\H)6X'89>A9=GNX(TT>17*G>8O[OX2NP,)DA*0^ AEB&FE
P\<!$1 3->AT%8+].-PC*Y4OL-9_KR?XBRC3?]T2W^"SSS,] 5E8XB7P T^SAQ3EP
PB*BQ A<A9D"0RE1;[LZO4?!:&>HXJL13=\GVB:89W#] +9_@]VR:H" A!6&D\-(8
P"(7K+X@Q&F3AXO3^T5E4I]JD TZ+3!,S0G3 IV[()WC66"4!E,S'8%0SZQ\E 09X
PN"-HXB(,;H+I:M2W1L^)K#RG7\-0\:>["7>7T6"*"+\2-S6$,7*C0_/4;Y*<I[MO
P&5]'PKN=<W(K%(VD"?0(!:<-'J<#WSS1',O,Z)MQ4.S&2S^P%:&3<6/&6)5]J'Z5
P:]= $/U2PG*OR0&+_F@0G%VYW5<!ESLT#N(:,JRIEKT8D8[G-[HGC*%X%'=#Z;@*
P(%GGJAK9 "E5NL6/8(9*:L@_VZD#**(L0?3-Y#>JH#1O>V>\W\P[OP<B"+5O!:A>
P)Y^<N7 9%D7UU@O2RZPT22O>,TCNSF=06/\W&T:,Y25NPW4+K9.W=*K=)VR5LIR.
PJ)+=(V.*%01"N>2=9T 'F%1Q2[*^.%(J%R)F@- ? !!:?,Y/O-!=']AG(;-TD($_
PQ,3^T.0'N4"&HI88?O][80MZAT8%_U[9K3XAI-Y4"E1];SZ#"R\V=G']Q0T@47<G
PU[R2HN4Y.I99"['R9NR@/66:Z]SNAW8')61T.YDQ-7\3*DMG.Y5P._O94.48S8C]
PE_M(<8=CPRD)?B V<UB_U"T:Y[C$@QEZT)3=G'%(3%^5Q[IVD/;8C=ZHU"B&*;Z;
PXKG4'_OHKG#N/(9U)?.;6M9$8T[6J@,[K=B/S_C=42^JUG=-_H\@&=66?<CU[; %
PNH-#S%DC3:C'SNG,V'#98R?L6C(2"DO]_6-0  <9/:K:FE8A2D;@+2U?[=/:YP\L
P"TQ!_)15O% ,ZA\L,7B9.!-X]78I6%:\=L4F.A_H?-[#M)!>7(I LF1S$U1IT2Q5
PG2K6U\$0YZ%H)<E\G&I$HP?8R3AO":*CW=FD5\6T&XH6ZHB,%#JK C7U^9:>E54R
P8H7TLY=(HA+6XFFX\GZBXO4<+$7C63L<@:#LA8(FDJY8MNFD7$RA;M=OD$F,P.%>
P$-$ > ,QTB.Z5,3*?H9+N,%C7#IZ/I$U!MR@0J=MJ:>[?VBY<@=HQ4I.$-6^W9-M
P5=DIZL@%D)]6WY7N'3<4J; ?F[3_J;J8^@GZR_P4.N+%%909L:Q !EH0@,0;0]!9
P1F#YZ;)RC #1R8F*[4V'RJ3ASHWLF-379L7L\JGF'32% STH[AH0F<Z&<M!D@Y/#
PTG3VU"#3T'<2C!::9PERG=8\K&'-D$)DO>:DF:/%!?1D\"43T/634!*,B?WVX*91
P+N@K:J.=Y^D87#GLF,FL)I9M7X$UJT%C9*N8=^LCP@'3C4ZVKOCH(;J6WL *[QM"
P/H%R9+A;<',A.2P77I*C&V"U/K">>8S$[KG7WO"3U0*B-IB:3AP7=E &MEO_-7AO
PE]VXRR^;*]^RGAQEJH4RWE"^3#,'(@PJ/L])%]^>\AB0+-;]4IYO1GV/,2)W3W4O
P-G32R[\0@" [)U$?;PD1;Y,'8#UE,T1_P-Q5A$A9>OOB3"&<?U#1\X1X52H\X*).
PVC;NOOXNHQ&#[%(D3VWH:Z:016X/<6:W/M:N7&UGB4.MPL##$A&5Q7N;C9O=>92*
P<\-XWI,&M+=S!X)2WKD(5_LO)5%O_8%"*G$KDS40@9R7S'3Y:<!K)V(5)C:(HM03
PM+%XO)OT+<_C&TGE+]8)K'&L6HJYUCK%VG=MZ_G,J*F==]A06+51D605MA)AM,J%
PU_0N%617F^B+$*F T[B>:N1IV>79W.]Y@[/>'N[(&'P@UCC*(VSB$=(F3WV$3_M:
P,Z#SNFEQ/6@0<7_K.?_"B!YY7ZGVFSB5=[L,7X9)BX$YZEPNO;^G*#ZT,U;!\>?8
PD#XT/#E:*8R1=&>?F$>:O<*/DDF'^\AD1S11^EFM'6KBWAF3_[O^-0LCOG_0(K/E
PF/R_J0L:X+(580@A]/0N9-;/L F0,\H 8>G/ICN%;X/K,S#-BNA<PRBZON)#%<:S
P/N G!<+Z5P;A*.*$Y:",;7WF$:AL8Z$D9CUP"*I-0\5G?!Y+A#^5CVE;8-U;*)NZ
P 32T8$9+K[-_V3XIV9Y6<%[ =':+7*"A&$J0Z,6,PL?LU_^".SA'@#+-Q%[QE%R@
P02 ]TB8 8L7H%.>37*IS <@W57L\YCL26T4X)8U!LBWTV>)70*/!G13L\N=]==N2
P&FF&NANP!@_X%#]E+$8<;C .I"+R7KQ'\^D'V.-K;$'A2UZ:H(OHE9FJT'53^X#X
P+V/;*F)$];NEKV[$2O?*F?\WJ79-]2-+II['E+!"G.T$.KXM"=RNK7%_]3R1D#$J
PSY*\7/%DID%*1"SA!O*4]<1U,WVH5E&/QXT$RIB$'!C0X&F,=;22*!=].%"J='G 
P= ,FF.P^*M)H-N8T1';*F7LTO;'O;!"D>]!.E* Y[4F^!YVL042!(_'E(BZJFB?(
P;Z(;)468^]2K0<LY5^ES_'6O>B])P7I$-C5 RLHY>WP8XM'3X'R!FHNCVO=9$BU7
P3]_C^<<9O,)^*JMN./(-$3L,D=5&K])(A@Y:P8\__DP71(?-FS+!O66= )DZVR5&
P=SYR)9-AN:!)U!8'3"LH-4!J$!L*5M#":F]B*@Y>Z:I/5J$?KZ) O4N;>8WKPF!<
PD4;PX6*6=#N%.G$$IKT30!'?T9B1[D1F?]?A1CTD&3F"I,6+-3V]A+.-,$$:VP0,
PKGG/60:&8IJN6.1]X8 \Q@^'.'W E,HXLH%_6>^Y-7A")U/)G<% <[U$"H^FK4LB
PV99S8)EKQQ^:E&RIF>A9_&F\3T0T(XJQ<*71N]/](=]H"WD:I:[#E]QP"0<FXH?-
PX:$#Z=HX?UZ(5$SBY5ZD6O%8PLK65RIDHH/Z:#<(2! D A3I0-K>JT3XI(*7/IAB
P$DS1\D>C'X?$W*X;)JJ6.LPSJ\F.5TB&"-AH]DDF^-)BN*(WM2>>#E.R7B9U\>C[
P2NR:?5)_E&%R52I'\WQR$;]0X0LHERZ$G:+LVAVQM=N32@;]DTYJ(X-I.L]MT[1O
P\!Q4\?*6G<ELG/YV(/QZ-'*@F$$M2C,XRXLXG/;PJ1X#2=$U2KZY\XDW\M'^_2FK
PLX8L&JOG34K8B60V+,%4#\/42,OQ^US5>C/1Q27*V8Z:79K@U)9G8B:B^&N">N<P
P[1JA\G)1ZXBZMC^<1/:@Z##X)0 :ZU,89R*5><3A_!^Z.8()\*FD_2$]:,=Q%T_!
P#HXL>6$D(:34V;LIY:75Q+@&5G#&*7.K!5:0!>86O6-6V^); L/8EG88Z'&'2LOJ
P YK4[;0@N=8 L@KZW&'^:>EX:_)&N#BL[GI)N@NC14[D'+;N[OZ\?F^)NJO4Z]5@
PF'[0W119CL]$HNN&^(O3MG3TSR37FT-_&B"N%3X_Q Q2XVIMR$6?C!_;[!^#56]<
PTN#*[IA6QQ?#F^AU;O;,',1I,>5U:[_\>;,')<BQ9^]U4@/H30 >SM=%W_2)DMT,
P(X1SN\#(7B$J431N<6$Q \<JO;LD#YKXH\1,#74_G?M?1P4Y?GGNRCH\#G[+JR38
PW<$8Q5K)^,7_W<9$5E-'^BD2%HZ5(;$F'?(I:Z4@K;)8"E-DA7T(R2D1MYE60[J(
PL(LZL&B^1>!3+%GLZYYU= [RL.%2S&+&A.F\MJ01?M[")E*D;FO/HOPJW*-/W]TH
PB=J=_XEB7V@;7S*@&B<QXU)5:^E":1I+8J^%I(N5"7?:DO4JDM--15>)U:H >^8X
P@"G_T$90F>T_)\59L?IW&1C@/&)):%P%'7I3=<3UB@;:/K!.8Q7RCI H3&N8CQU;
PL>;RMIGP3[AKT[I5)/IRBS(B/W&R+9^.#!M9MR8H^E^*/6,/"YH8*1#]8<-!)L;;
P PU9NM-;LQWKK#?.'$!^'>>QIA'&5]C''X=]IDK4Q_WYYZ;QONX6ZG!OX)T#%O):
PO[S[KT#GS"-&J5Q7+16(9B0G1IRVN1*,OP9O!9L-<B>@&RFGEXCD4#;?56!Y:,W(
PYAS="(MY]MQ^,PQ+VA-+ +W4>I(,D!16XV3%F4_2H$<9&%5#H4?:[^G,,OKY>PWD
PP^,P,-IUH QR-NY0,O<:^1OG/=]V)*@1ESUA[K'<[XL2\1A@)L.^8<-[+RB;B7V<
P/W==Y:6D\&X0EE8^^]$X;Y)U.<\E?RMK8-9 @X.H&MM=V_I>#?MNPK6;GU'MV4"I
PM4; TU!PL>P4 Q%$,BN!X>0V:(6&:(/KLB]\6VV6ZS\FH8:D)R;C*'I2TP=2R.3_
PZ=C6L]EQ(1P.P<8Z0NH_!UK\9LN<E;^F$=0?$C5!$#/%9J7>2BS^3DF+2ZNSV&Y-
P@'*G88Z].7=$VO_=^H"6(?J^'E!_?N[WC 5T QO-[%#JH/272"2F1^B?J&@UZ=34
P?'$^P2J*6O\2L&\!R)A@:CN_>7[AS@\VYK4DVF?N,*-Y^VJ*38!$M.;BGL4"%"W<
PJ;\FW>[%7X@+U)G,WY=>5.]R@<_X?N9%S]&4$(+_XTX6_",O&(@78)X(PG_+RB9%
PHQ19YZ.!)0>,,S'E[^Z:I=W 4?L2N>_*F0FF*Y&\ E0H2?!A)UG"6W91._O:_;Z"
PG-<4I.0#JM3WSNB939/-8R2<\8JDB["#%MC.MSP1\B9(([%C1PR) &_P49BRT!0Y
P[$+/R-?SLT<#PZ) 3S!'6_6HE:?J^!I?SWTRRC1!/SWI[I-E[KH&L4*7X\J)/M"*
PDZ(D7?$<049@"ZYXV*5DZ(TT(0I_-<5NF2+4YP%T\ME<>!*[>UR_6DX-R)V9^&(G
PG9:0A6(_"3Z8LAX%B\A#8O/"?+'UOL/+IW]<\%-5AE2GZQVZUI=VM!N !Q%%G1D>
PB YEY"B3$28A-6.1>T<Z37ZXU!:&8X%Q%_VF->(JH#/FD_B1+DVF\GRO2KVCU3Z4
P9<14A:N;^?'1[/O;&&FBKCZ>G&A5?5L5G^^Y9Q8OO6[(*T.$&D^#1O[5%2@Z%1B-
PZY-"HO"\R,J"APY^C,%HG$U%#NF'\GK>-@>'_&UV@] 2TSG"XF!5+ZX]F3T9%GDJ
P?P=B=VWLBIYBM7IR47O+.!-]9M8\T*2Q$WA/.U/I(+P(H$#^$UT]MN%=/5Z_R*K7
PK[K]_ H0%.<<",<V\$80_D!5T+_8:PT[):X5]F%3A_$I!Z*S4C=Q3Q\9QS^0$-Y@
P/X>:AW!_=C%O$:/9Z8K5G\/;3ZV/Z:.@F<C\V:^.ZGGXT?55-Y]RBSJZ!3?O%=LS
P,XC#)E\R:,E-"..17H>JSO^7="IBA\906%?OXDES")LK24;"PM6GF7,U& Q=YPCL
P>3L?(7J6I9I0B.N^TG:[_<99E[_FA?VX?XJY9H7ZD6W#"%0>BKLD[ILHEL@D:UUU
P[KYGB'I 3&UM=0^VCQDWL'RI9S9X123RI1#1+%_#0VQY&7[H84,56MU@7CIZTA-_
PI/$!NN/:M:XT4)-T$YWDQOU$:_O=##1&[R_,&]=3?[5MB3J52Z;'WHE/EY-KB3XE
PXRH1@C(*B&P'\%6KNWVI$_.;CFP.1BY+_6>X5GINS@O*Z#:L21^WPMRZ]<L=)-BG
PV_<&F?69TXK(H(RE#!T/PJ*B$*3?+<+-UR'><871XX%=F)H\5]I(^"K]U/ZJ&BU5
P-[D,[8F/N<ME<.$>=&U]SC1K4>&$_W]G,_$+53_80<"#><%PUR+L-&9YO95?AR_*
PQ6,?!<<X$$\;NP.+,WS1#;1%FUYC*N;&'[*!CSCC8Q=6BM;E#;2Y[#L>/9]&T6+G
P3@6JMN5]8XQ_QI*1GR,K[=C?^C0-TDW5N9,-%O3$!<L55,&%?K::I9[?\-)6E5B/
P>&XP/@_]Z/7&Y,WMX/MV1.UF*M*RQWK&8!2Q-AR/N+8_^-J?WQ$&#NY2R:W9VD5C
PKP(J:85P-[,/DKFS=R.LQXBX6S#JMKA;2L#Z/F!A]X7^]>*'RPW+*C33(2QH(<CB
PP0S+!I[F.(.8+B]_O^9<;C0;UG8$Y(GE0<,6!!]QOG@X+_YV-*HJ,E?3_^6R>G7U
PS+ZG=UKLSS0)&*<F0%_'-[N7#/)1VOWGD_G4'C?EK::+=D:+G&B*ER"@#VW7HN--
P<*6/3$\S"T4%#L'9"7 2L0P";2_V&[[9^K T 5VS8QBQ3"@O5CJ9? 6C17^58_6P
P]>M[$2^M#'8**?&XT7-@ C]FY3&TSI.:!1721/.GEO0/<^S_"^%R%^NHP61;EW6)
PU4*9 (LE8^@P=*=^Q;9'4PR@'BFS'"'65@1+KWRB/CQK>;$[ES(&T^3H -D=_Z<6
P-7TNC'F*;V+B9H8&=(4J0J1<Q@E*5H('/;1:7@W7[L4RAY7G)GSR#:]#"(/T;A?A
PZ8FR9$=\J54%,?:WV?=2^*]J2&I;^^:.4+FM#QU%,-GF V>[O"V9N: M]3QP-MS6
PTNWC,RHI^R5*M:% ,ZU.DPG:R2>4FQD'_9K#\4O4X?0H$7E8@\B?;5B?P9G6$/<@
PBLM%K\;XBJ4!_YS[!R&\"2AO]"0"NX;.DL,C=)2]VO4VV!*E3LZXM[>#5G'#R:Y#
`endprotected128

////////////////////////////////////////////////////////////////////////////////////////////////////////////


`protected128
P?+)9#"+V.E$ANY.BG)2PC,U'S:"!PR:&P@-%,4ORO>KE-_ER#,[G>X 5&#C5I#RB
P<U&'.)_0]K&.#XQU=.-A)LF,]$UFW..]2 $LJ]E=O7T5U41=3U#V2BN@N(E9)D+:
P0KD5N3X<\P,[*9=/R! \?/J1#?,:_GZ%MN>RY7@A]D7-5-Q[H*C@KV,VJW.G14W7
PKS)T3.?#>;/N %>S+U#3>YU[2%@7V-HQI *)1\VI,:,_5!;Z5H.ZE%*TS>!3CZ%E
PX?% F^'5/WI2E[7@$/[V#2N)P3?QY9/EH\F<(,F@H3&1.A*PQUPIK,1]&@@#V@+!
P'3R!#K%%'/K0UN!I6.?BI]:O+[;@DAD>&RN' 1B1T@I7H5[(XWV>($EK?#L[E&HJ
PG0C@;[1R0"PA_-.#H<0UA1<(B!'DJ^9-UZ_ E; A;L34N\D&:5'3-E([2K"&VUS?
P=K/.Y+3/&H\)&<#M[&9+^==",CSTJ]W1QBJOI N .(84JI(R =HN]-%TCB^Y"( \
PHF6,^-&[CF@R?DJ)\>4>^S;U[P/*/[Q,3576_:32E]8(J<]HG?'5LN;E]%*OV@,1
PH\=PYI$=@J2SGX[WTHT>CD"O_-_(7Q&?KW7%XI;.G*Y ><R)F0SM:%HI2V[NAJ9,
PDKCJJ&:O5Q#BY?[/%"+/'?T>_"?YR8%CY*"1NW*X5?$M(.\$80!EO#RFSPX+2H[8
P#[$,/XIH758[/(TR$F"6VK>2'3]+V174REP"#VJW<'$O(XGF],+O,9QZOQYI-=QW
PD=S;"HVHQIK!CS;01Z.9&HE S,O^*_6C?QT>2@'8:A4AG\N)N"BGA(@<XYTBW(S\
PCN/#R?YUY/E=Z08 Y_ZXJ?:YGOY%V]T8E1)G=>\C-V(5%<ATWNI]?^K)A97FE6DH
POP/(=4=>HA82E!X2.9^,P-(;_\4>H8J$U<\H(?UX'?K7)K4XE5TQ]P2@F07$(78U
PVKL^Y-0;>#.;-H*&Y6&V%32\>4X5?LWC:1ZZ&-K,9(G%,ZA2E_ICSI_O^D58[4W:
P+LV-%"T EFW:+YS:NA.A:#J?X4@XK4L7*H A>0VRYREV(3(+3]K(U]CL1C@DF'+K
PJWPOE];EL\1L3?(E#28(00-HOMPZ42(@%]R^&^>-PL/]_88YVE2KRMMY $[%YT:?
PSMJM<!CNA0>@9Z(4W\ 1'/'1@?.Q=9QW9U*C _>Q4YREJNN3!Y[^@MIYJY/QT,P<
P_3.Z<A>QN4VU=M]-9R!NX_M_E>B)>&O/W,9*\I5IKWL?#.<AZ/'N"L&K4N2'R+&*
P"+J-8[J0B1^,^>PWO)7^63F%T*UG(%59G$Z<A@W8XN1FY8P'E48](AR'BB& =*2#
P%A7=:<)??:RGMP*#$RO:%P9*&[U)UMN*<_J6V$CVJ7\#RDPB7:WXAS6@P.*F;SKV
PS<P"(2AS&:ZG I\R'EB^O+[-.9O+NU3AOQ;G/[BW]:8E^;F&,FG5:L*059AS1YPA
P^A6O%W146%C,F<.#J'$Z+B<9]!*\F#IP_;X8UM):-,D*-6&W^Y(XI@/-G6(V7S;O
P9C'!RF7;EJ?QWN788:_#/.IXOD+=TR.0_8$3F'QK0R6>?F%%V)3UOSAL",@LR,>9
P/=>P_0["Q)F)U7+4"I&$Y@SIH1+#^58=PT9M/ ]BQ90)Y^#W\1*?,I+\L",X5^K'
P[5B@(DCKCL-@1<@7$#5[#L(-U#L&4WBWFWJ9N<!-5/5F.H$NK<#7 '20294AG$QN
P*V%:.+RW]/,?N<9:@33."9U]\^XL?)Q-V_-QR$#O0S>C)DM0KRBB_MCH4)\QF6-8
PX,%3A72\<GOBU^TZ?6X20W-W&#:W44(#G@YTOXE^A9$\.M24XRP2SOR)J;WBDA#P
P-S-=1X'K.!=:F^D-Q32)1CU<5*]4_XW!'H1/,=)@0:K238XK\+6)_[G)*]\0E-A.
PUJ\_F@QYI)"<6GM@(PU)CV#C$:O%G@F]";5H/ARQ;V/=V/DVQC<][&5#'AGMN]0=
P[97, H/V_7.SYB+P;$?I0-O;1+@N(7;XW%*SV20TZNOT5_[%(X&/-8O?MK.C_3CU
P-WQH--$ %*'JRMTRM*\GMS(<=&V%,9-I3[-*+TO%$67(0&51*E/"%W?JPMLR& L9
PTM\K6F!A* 2G?Z5*?#3SN]-%MY\;9IGPE@AT?*+8?0N58#+]PG'WTD>>TZTK9+AM
P%56M0'2K?MZT(@KJ8;,.IR4#(W0XA?TYQ5[N% 1RL\-KU44,/0%"0L'H2+.N63, 
P6T]^2V\O^:2%^<G?P*76J38N\!6S#@M@@_3)$66_TZGP:12#X'B:;I?:]H\/)K$5
P]EB";0?MGJL1*10+ 4EES*RK_:MO X)1EA==,,4"&[9\\1O92.(S+4TGG>%,@"NT
P#BUQ@GS3Z_ AS1R#]UQY)-'/N])P#)_RDPQ9M\93@P'KCOFTKU)UZ;1RMYQMN#^2
PT79B<%%L<IZ6_G&^;JW@OM[#RBNN.X$[E7"%O-7CX0'4.1HQ48_ZU(B(C>-&?XU^
PA]&@>#>=KPI=)%)<._IU+N(R/OE]*X^&(O]].CBX!O%\[/V>ZEB 5#-6XB@1H^I6
P<_*Y19\S"&P2L,.'S[-K,835>;E,J_;U^KNRN2D!>!H<AE+QPUC<MTRY1T5*MJ?H
P94I36+#9LW+C77H<3 ;H$M[))J9.Y2RG\H  J$SKJ2XI5!EK):TNO4;U0+==LYH*
P7YOZ<$Q6V27=^)U" #_TXD!E(C[8#??KAS:0^7@[R+ZEY9,-RR9\Z$#:V4\3V.PQ
PSYB!T'ZPD.8R4F>)4<L$_C6/ZIBT&4)'L8]/R#)9PX^86Z4/;NL.T896;WYJ"%9'
P\5*/'EI72)OQ/LD7:LW2]^&;[:<O/]+W_\QS=%OZ]T9(NAW)',7\-L%MZ8L/=3IK
P;)&>M+K1AT]A?"Z6!B@$N/"V=L39&,LPJ!C&/BPT"/7D6&_'Z,:ZPECIK,3MD\(^
P]FG^#T=3O!I"T>!Z*/-8A9U2DTE4* &@W?PKR<]6XO*9T:",F;HE?'..V)_9/SPE
P/B%)[+MJ?.,".7@"E:!^#/VCJWT0,!;KC>#%IS;YU9J@ &3:V+>,HO0T/35K'230
P=8%K_<8,UCKB$=F@XX3SR).BG&ZK+GG\\XE^'GFN)N2^K$K 3.X%<8_T^>K5Y'+V
P-J,.RV7;[X!*1)U<>Q2HEIM;5I4&ZUE,>E6.--$4B=-NB<^G9A37[).1(,.6 8%;
P^7IO,6&P\.)#9N_-=1-^D58J,B%3%F ("-,2W[Y*ZVK;"AQ/F>B@M^8LN.R*V(33
PC'/?I"C:O"P.F=0UE),CCXCZ3V*/0M= 2ERCV[PPILT[R/AGM0K;:_)10UWT*T50
P:1Q65A&G1Z%G5\P]&D%*!OO,;BMQ>9ZCM9ZS:O3\>$IJBQ?QS0"EH9K9;! 3\*PU
P2TNE6K6$+F^I&.6W6"<M\3V!IY"!A,$>-40F[G>@"F_8Y1]#7X]&-,Y8OI=\Z=FQ
P 3GII6$6HM7.R42_!ZO:E"28K>APMV _X:-(A9KV,KT,]UL<W/%,=*UL3+0+,MSR
PF@2.8I*Q WS4,$-C/3J\48%!^*FP8<$(JQ9+NVHGM(>+Q;::_2VEUG-L1$]%N]"J
PQZ^%1S6#?+MTX[7,/<8\ +_'7[<AHQ0L6>PX,GP?4N*G>C)@<2]/KLN&O?L);DH^
PKE!7 +U YZ\ 5Z]WH5D-L>6 ,Z#+#OLCNG;/'YJ$\61L8_\F]U:,'& A!M]-ME7$
PJ#"0$)&%?ZRSWT\C4;8J=L1U)N=^53[F438(7;\HZX1.*'X8?+^,5SSXY([.P% _
P[1?/5R2G=D4\7**;,BNXI<ROJ_/-J2: -=@=<JN)Y?2+024C[B8)O L0+*1Z5Z"?
P>],UXD9P>99<A(/.%^0;WNE ,GV<Y$@@\TFV&4L:>7B\0WZS-)4)=;&G+!7PW%*L
P0I& )9$X[;PTSP;_D/'MXBYG\ZWT-I<DO #=K"+<22E^1D<R)8*S<F<-<K@H]+=N
P!("_(:119 (;7'1TI6 _%"&Y)1FPQCD2+%WU:UD1]MNSBGH>D37;V7+/.9TOU,.R
P_(B=?Z*G"V"U,!$/<8+VJYT0WHVWW12$E=U<@01; F+;U61-HBT08" 3%I1>KF2,
PBI_* *\##,?C1IB+'<"Q0VPGK3(S98@[H+-.)?0BE8T+96]C_8.3Q%/,K$+H+ 4K
P#Y0A.LR7:M0>P48>5_8N62?2VW<8FAMXP%=4<T>*1-,CT7<U%?*RB]>$FYB\J>FK
P#\R7+:!G6OZ\ C1!,Z*R&E=KT*0$A@>+%J6<K=]"+ LT<Y$$)HU'2 YS&Z,5J,X1
P/4<-3V"_WV;O:OQCO=D8.16V;VI\5NG=:G665O!0FB<U]VA:\K;E6O75LVIYNY8Y
P0SJ?;JM*;.IF%L?O"U39 G'PW1 T):N'N1XSRHZS]T\NWCO1<\_5?G[$\8!S3B0,
P;$[L]0DW*]JK1<4U ]OUM JQZLWJPFWQB\.(K;..4"3/MX>8 L/57"=Q_N0:"V3J
P]^7Q@@?1X?$/F.4]@NWW,:9J"&2S:_.9R*08^PNK7WU](AJH\WG??!/,0M@ &^'=
P-079SN"_CU#@;]@HQFU_6!<3$R&"/JDD1_D OF5)TL6]7?,0AS.-Y[*KN81]NAWZ
P"YCKQ$JR@%N6OX,9'D-CD^[>J()3ILDDC-#Q[!D$=]]L,O]*)S?)$@:IE6!'#@=(
P^TVW;. UBLRBI8?7:4]4Y=VH;\;<K>^&#E3S_Y))4ATP%^B/YM(_!+P-POWC-X<U
P:+52>"5<2 34;(9GH!8"VR%=*:C2\LFPL:;W (263Z>U@2K9NO3463Q6R8-IPN<;
P4\92UMS_U0]-@2I-TZ20C<DLV<V>J?]QG]?N[0S@?5L^LNB939:FM+J5!L*(D"[J
P[K L"YHH9!5QYOR22X)B>,E^A_O3\!D&BX<^;K=C>D(VBN4ZZ3:N*3KI_L7CR^4G
P+#?[K><5GAJ[[J[]\_U;,KBNGW,]M+9(/?W:WTIGBS*O1)CN\1DNEE1#0+EO^NW;
PD2QI;28T%@ -#)QC@<L@[%,762[F"X1&I1V_Z![\_,(6\;PO?4,Q@>T_C)RYM I*
PR\YM<#/[K@( <FE+QR0)C[UDS\RQ.1\HVT%E0$V(?8,5A,?Q\D=VO!3]D,<'>6S"
P;%*?%H.MQ73EB"<TN&@$L,<;3JDA7?"VA<A?5C%E_!<,--?AQCA2E+Q?GZ&9=&P.
P)X*,\LL(M"9;,IAZ5!V:S.,PD_^IO&(0VY=+Q5'B);:.:V15K?2X3UUQ>B$!^1.S
P-P0<P?<8*=S[Y[M"\VP_V0TRMS0J=FY?(.U]T6D.G50;N]CL,$JZ#=(7ROPE$<L7
P)XYQAH[2N(KO\>%,</2AA3ZA@SL+]"8FR?5[L?5M=U*8-P^/%T@RH*6>4+]"BV*5
PT]?F$/$LFKZ+%@??!>4&8OZX[ G&-W*EFF)WN/DKL4L $AIN$:+V]VHAD/' L7I1
P<JZ6!.*-@&;CY<=NV_3S!Z(2K]^'^C(I=H^_3(%'HVF7/?2S5\;Z-A3R&FK:Y_EN
P%MK5I]]CP_]07))= K,H<U]U7N)F3B64+)&^89;XO4:>/BU"XS !Q_,"\E-T*<E>
P+%VS<5:H_6GV2'Y+[\0]J&BZG R\Q1R^\#B[R_2##W:8Q0WT-PKN5D8K#1 @0[_%
P<U/R4_V;9[83JG>7SPVJ/RUA0-"VLL#DF4'5:.9 _BR&9+O2/*,%XT?W,%GH[>E>
P?-?J0P*M?R=9?T7%**D[E&RM+87;7K)^9\2#R@#.LPI$4SW?>@D\A:L4;#,$%W[O
P5D63ZE=&1K]TX5Q*@EL@<$T:088 MZ[;\^#$C(8=E5V*UM\\LE(C=YY"VZJ'6,#2
PQQB3W?+-7WSH0V^5203,!41%S9VE N%NILPAB2SG0J%=V8O,>]H54KJ Y5!8E.@@
PX88T,PY>7U,/WXSYB1.,I)@1> [!JK$OM6M )('H600(7+DY1>&1'Y2T4%"D.BP;
P\CHGR5 7>EJUTP.!M_($ XZ[^\7J&C#V6:K9+\/2]6AXN=M=4M'RAL%8 T K"H4M
P^QH]K$"]Z+R#(SYP0(<'-[\)5/L;0/TGDT^LO!W@86B^3F19+L1Y,>Z,B*H*?==X
P*C_>;"*''P$7<X0=#22*YB5/>VQ>@B-&C9,;#Z0KLJV*>A**)"81!X);?1F$D9M3
P!4Z$M@_ARW 8S+>G?<)K6.U>L#('U?5CBEM<P"D/>]J94K<<('/3Y_A0G@6[X&H/
P)';\[AY!U0T;!K)-6[4)"L2"^\QF=R)]>5Z/(]P0X^))ENC.LBHG<^:9BV+]E1AC
P3[Z_!-2XR?%PP_<*3@J8)0YUNI":@Z'VZPE#PRO9JA##,13Q^M65Q&"5:!H3)9?Y
P4YQBDS2&%CV<<6PK0%#%:DSY,):PE@-,QS.;IXH!9!V>8.TW-*9%K/6._L^QQC>.
PY_)I&0(,^@]P\JK[8:Y('P$^JQWO;+%<0:D%9,;=B2;H=H7%F9GP31GZ=R-&Z(,D
P10,>S4Q;3;Q,K+$;CEU&T9S5RX[756.^-):U62>!(<Z?35)PR[_2DHE*/U"^F5A3
P^@3T]4)L:)UTN)$TGIV,.W.=UDF4*'#$DAU<>5*W%![3X37=1.42Y9U63E;U! A3
PYD6;?V2X50-\<CN:Y78\-LQJ36\^NL78I,21X>P:H^3M.DRYS?]BJ ,^V6#80UX8
P='M]&\8 V&D*OP"IJ#/:L6<=$N6.X/98CY#6.E![,F@+ @T62+PQ/C<R 7TUNC>C
PA>=VW^%Y>+_MCQJK(-LJ6_Y\&3:="1TC?^QI@'TL0C,^_V(=$WS@[3%H89>39)Q"
P&8AK\&[8RS0(Q@++C-2=C,3CZ0LZ,KUG5ZORJ48VN+&_(6F<ZK<_.I SEXX2+TGO
PRBYV9*%M=>4:^R::%WQA$?!>P^8^I)PW;X/;I=X-1BDHW5#]%76HZ"*H4\TA:+'3
P70=5MQ[Q45=T413LP&I.]=K<WT%NHZL /\J*-X3N?*?B$&( ![X2YD25N?:OA)L!
P3LQU]P#D0FXO7?7)AN)E%;?+0<^REMEWDPX:B,!#T9T!4_%  =,9Y.LCIR=!C&,+
P_D-]8ZQ,M=1HZ!_!IY=PP,LS);WCVG!?%[OR*%E>0H5$T%L5F>.+1!P/./9Q[/N2
PFH974O2&#<$QUN&%<QN0R.V?LV!M"QK:<>R.0@-:FL$UUE X@'[BC#.?>#.LR+2S
PC)8[SI!<O:@\\CFD?D=[_&A3I/-O.LDS>:BIBWN0T@8V!"!@\KC)+68N0LL;+DT6
P.12]P#(7<8J]:0-?V^BP;)G9!@VX$27FVG^BY<00O#:#&HYKE*$$9"];_OWE(2"-
P@VD;"L@6XB)=DN+MCD 5(N$U)(H7&UXAZ5HO6X8EYU?^\@0EU6M#LR5LM)QH&!32
P^+L"[6*M5J>!&@,]D8H3Q!&]?LIE",TG(]\XI<IA^_/"?_8SE3E[^DM @_RP-N8"
P-70^=M2)@T0D:. 4;78R&GPX=5+72*)8&BF9T/!0MIMY"&=$>U@D1E6&J\_*-)=:
P\"1QI7&ZWU]BK]OJ$B[39?N#6SG)5NOUVN1TMZ#M)$P+V^6D(U^SX% 9QG\VY(X(
P*4*T[U8I@+%%[;CVV"X>%'/+!=&V7N=0OY-LA6]$^"N-[W+YIMNW$"?1A$GQ32L:
PR2JC+:NREU8U8XAO;$M^+>*I;;,WI[?(X6D53H3)DQ Y"F;8F'V$R<]QY<!Y+WC&
PF9MM)[I>VM2)7C@N_ O[5C3*-H:2BY$Z]WTO.H;%5UTW18=2]4/FJQXL;G(%-]28
P"1@,2(N+F*2I55GU4Z=0IN'T@YX$+Y!9'E=C.?'K-1I&*&6 KQ)VP=VR8T!XO)$R
PPD\':TEJ3#\$LTU/1@.&O]^=[!X4NQ+4G3.^M:+>,?EM;K__?K"?$,+*86E2I74D
PX\'=12@*LC5[E^'P'3W[F)=E_;=$^UT T" '5S#&O4+/1W.V3?X3?$W33S,;47.J
PF<:*#UYL15]T1R&(PRFAI6+FK^S548L"0)-S/KLS-MY'RH&0(+19NA-V^C%!54\K
PMXR1^!I2J;.=3?O908_+'!^9=W.5Q(KAE]?7Q7+_@C"AB;5D+H$<Q@M=*%R3V\#U
P4B>U+2BOLIT-6\O_C/E.QZ+5=: O/816K4P1I2XA*RK[S3TA$KX%!'I]%M68LIAT
P=5[R]]876-K6^+<E)?[+2!=<&6UK&$9>N-PU[<5\UUHMJ P@F_CD^!]QGJX)+H&8
P+5.]Q*\7E&?377.X>K-Z.\L.LL6]%9'0H*%1L;!@3K9UL++Y5@WR%3W/_1X",\P]
PPCT+FR ^@9"W'$[-WZLLEU;FA\A12HQ\]_%+.?&EB)'"R9]<_L!/F3S*+(.A8?K=
P;XMT09.I?>I:UD9;&#+JR-2H:E-,^/ XV".'49OE1Y7,[A>_36PHB^H>.3M:8$N 
P.DH*N)F:H]@K^64@!D)E<0/RA!H?";1"4OQ!4T*?:2(=+"&'0D3WMQ)Y&I)_9,<_
P9Q)MJ22DJ.:NH'T93?HM2W.UL]"$J!U^Y$^C:\)Q$WF<"(DC!<]BH]ZN/3]7>)T<
P"WW.BIX\?2_#7>_!20042"RN+E3DGT)=KOZ[GRG;_'4?@RP!G#J<=59(]U[2%95P
PP%[Z)X7=3,0E9<#*!OS:I>K[$/XI*$\_=]YD K61G9_0;,*6@!-N@3B_W:M<U $ 
PDA.R=S=I%-1>&KH18+;*)1ZXB"J7' /^&QA4(G80,,O@.J_@9N/0& DBB<%L[F*9
PK$/S;TL?$1M/[BW"[?#!$:2@P0$G8ZXO,+M5[),DB] ;.4-Q@'4B5V9@#(\1/]OB
PY%HOT'#GW58[68FY9W?$KTS&?;!._)RQ4B5'5P-SCQ-U*8=[,Q'AX"X)'+JQ6AK@
P>GU!J,68*)+&417CFT]ZBZUU(X*XI9,4C>3$6+T%&*Y$8@4QZUJG]1M0;W;_ D7$
P>J8480&@.9O\ SUL-A+9IC)BG9V;M#K+WT!D&>S^M'J3(Z5^K 8Y K!I[!<IE[9:
PA&T)5NJZMHZ2FS#,/:BN3C<@,11^(#LVEJ-QG^2DA_:8[1.:ER8>@*KX1W=R M/E
P!P]-I)8*.<0#>(YV0/2[$&B%6C^2T=OQ@(HD3]?L3M%.P05EEE;A -6=O.N P$G1
P%(KJ5^+7VM4^W3A@W:0D-].-J,3]_7N6=-'\TR4T'#%QCTQRPD&?KQ3?J&_R\IRX
P9=U_ :Y*L<Y)XKOD0"]^%.W$D$Q!@;>*BY]FO?TN'_T$HWV_[5UB\:Y?&Y-%+)]X
PG$J]P790\'>!O*5 [0N&DD3:P/7H=>#SVNVG3A'HV48_V@NI)L4?<>]89H%_!0BI
P"MONB$7.8:OM&+439^O<=0S,GAVOAG$]313>=H-9;(<VZ&&6$ UDA1O-NGU/F= A
P56MD #Z84#\NO^6!=!%7L&TI]GE4VA6?P4ZB7[)(K8'VAD6L)7!9AP7W:VY%J-II
P9+M3]U;D@@L@K=Q%F-NU!3KHQ@"KRGN,'Y\[2KSI<N[N7TQQZ/E!">/!7E5JLW@I
P":L@(*2&8&25+J%1)S=*@;<K%1?_.Y@G,RO6G039;66E\H!LRF8B"*8J>+9TRV]W
P=09N4#_#!J3CD-;PZ^IKUUS3Y,ZJ3<%(0,)I!;7O928YGA2#JMQU('& CJY( K)0
P0)\&9ZGY)+ZMNPW715P_A>Y+YQ2>:&IU'CV.$%C8/:<7%=BOFNW1U0GI4,&-]V\6
P'[LAA"V"NNA)9EP7#F7?PF^.HU;@?+,.GMVWI=(GAN!LJLDYOE41=:=$6[-S>Q$0
PD;'/H:^]KK]PA72X@5<=HML(AM[E&"UT,1R&.AU"K-NO]) I=[UO[;BY[$"L ,-.
P:#]GI#"DL19D7RWO=]?=@P9?T3XCD[.2'_5;[0/JL'N=-HY769FV!7@UX<1US%\)
P/\)H;0"0Y(MH,ON90UDH@;H (T!.]4Q;I:^\R[WW:NX;[[&&\5^ U9RB -*WOMB_
P4;?XLM.\F7A@;E^CO,.SHXG1AFW2I+7Y(Y#W:2_<6:<+I>VE(+@9E$O*0ZWO($)\
PO6/R$:V_-Y,>@3B4D_M[$%)O1);)A _;RJ@ESOC3E+M>(HNU8JE;^T%^65:Q^8RC
P;N43%F#T>1.6RKA=E\\%:)0B/T<V\<5V!VU\@ST#>E<OB!=(TO+,O,.-P<%9.]1Z
PG2WH9<;1"L@<2#0-QU'"QF$H[CL,(SU7-!X+<-KW)^$**@5YYJQ75%UR9>$C1XO@
P9C9QOWXIESPQROS&S]W4S&V:=+D46=(.LS8,)0_Z@*E:4*@&^VPSZ'[%IBOU3)$:
PK =.A:.EPRBAB(T5!*XN L0=8^:DOAC<Y4V"T*<7&$YO3 JN\SX^ZR%'>P1J1=F?
P]<@8)X*AEV_ G*Z6CAX.7CBPOHG%X+IH.I O$*)V10:Q!](]VC!%E7X !6716WFT
P0J<GSC+GFINMDHR?>T?EUR!?T:Z4X^O?SVIB,SBUEAMRBGX7WYF-%2=]EI)?Z@NT
P82B[W^M>48Y.\@GRH23!Q]$S#05JB3'BU>*K NJLTEF A+.@X4[)W1^B49ZWV1"8
P%CJ8SAH=+9^!OCE#M1$Z8.?S"K5?BNMN5]CVP\HW4!_=!TX%]E);8)AJ>(4T(0HN
PEJ'QG?>#_MUD;1&YB==1OLQ-<Q<U.DQJ9C&-.#Z']"X6,?_IRQKR6E*4*JW=)%9L
P)0:C.M'2+/P37T20*I&M8"3>J3OSF<5;H&\/OP, <9;63-/SWF>OY&%9".;0G]TW
PYFB)]RC[H]O >"L%; #>7QI%>D5&S  ^&'9&W59BDAV_&6@Y[.<5T9USFP]6Y36G
P2=WTNO886B(/,[4A!IOX*N$T<B^@TSE4.E@(#3WU<I8Q:N?7=<L^W_."'RE,4.LI
P>CAO3<;8-?_R,Y#1^!5P!]A+2R4<]U9L'<[TXX)!VZ6?5T%FOA1&1NQ\W#*= GF5
`endprotected128

////////////////////////////////////////////////////////////////////////////////////////////////////////////


`protected128
P?+)9#"+V.E$ANY.BG)2PC,U'S:"!PR:&P@-%,4ORO>KE-_ER#,[G>X 5&#C5I#RB
P7P%1OW</D*++,<>I>T3^CVNE?_MW71*8K^<A<8^<&CR&^.!%YJ/*CI2?ZJRO-"H#
PR;EF)?,<2_\;#)-1GB.I1ICC\3Z0G2)C5UV>&55(#%#T*1&M:(]6.R("2D_\!?$J
PQR9"3'>-%;T5AN<#ASL/5=^M)S#)8I;<GTP_R#JYAZXXN2;+)_^N]%>3?.;>1NGI
PUQ\IFG= 2\_\R+QV'Y?HWP%O)J827F>;[E!^%*\])Y%VFFOJ3+Z[:/\XSY%]$8QD
P%_J">2$9%WY,Y14+JW:@2M#7B\G5ES@Y#4^'(OP/_2/.B?M'5YC,2(E/LW^7VOHB
P^ZJ\F80ML,5GJH)G4DJZ+7 V>'P5V9(I7T'!85&GI$QWRS6'\(<03"NY$CL )=/D
PK'\S1Z5,.2\>,A$<:2_!T-V3<R7_]4?-9:K5!GO@%_78RGD,5Z63,].G2(6W.'SA
PVV$40RQIV2Q9[(##!GX%5IN;I>N4<>>KN+:18S7J<\![VU?I'BP#W"SUJ!&H"*.#
PCE\_1#.SW\KP(5@>P@2IWA-OUZ+YV&JG!#@5]QFS0UE2R*-=;\&!&A,8+N ?8;<7
P'C?]5Q.FI.A1>;)*+SV YB<]W)N)(VJ797EC.UC/&4?%_AK=O'(WO)<3L)^I!!2O
P$"KCVIQ4^ (.]G0VCU3PC4S@ ZI*[AJ--GMBK@^6&Y<Y*TR[GEQW/E]Z<X&%ZJB$
PL"9@V;;FOL%\)O:JN+*=*W^FO%'4*)'$#0]R%Z,6M,6>(2&],:EU!(7UC2F:?Y$&
P+BNOZ[;@(;W9B(\)6"[N\_N6;9 /N&:S4"Z<N.(5^[(\2OAI@R91K/9*FC1A7)GY
P6;"I.$2)NZ3<D42JKY0 ZB:!,Z?V(PV,8UD,$&E_/Z/3TZNN)B.WGZPH+!.2:.1:
PG9)V9.]M[/3)K_BA AH)9\T:I17.W*\GG;8/LV>[QV4+?)3F:(UQ@ ,&B_7N3V:<
PB@RD;'C&$V<,#G:-':AXH$P:#,VM]/-HO/%\:W,O40K+9%Z3/MW^;8; RQ MHC&V
PY[-L]IM.0"&2C4"30X=#!]UD,O(<%A>^E),3ET!91;:B A&48&@_253YL(5EFP:_
PJ+P[>I,V<5GF^9'[M01Z^W]WP6DZ\'67WS382,8(F:=9'\FI!6UU3]#+QB*TD9=\
PB$:(%QX?C+?F4)$RYW24+2,/%HJ+-#D/E,522<M3NC1>$E'^9A,!:(UL(1XPR1NK
P_V7&'NCHL.5YQ$GW,B;R=PMSUP\S,.H5G".W[P68"6B832C?:^"3"YWEPO[&6,YM
P0*H6+,]DRF!=RM, Q[22"!G9^V1#+M_\K.D:%'<.:.6AE9'PT.VII[E<PC'DJ=VT
P7WRH<1]YZZK/(-+8$Z6GLF07J]W7EGF5!^P6D@S*H*=M7WO?3^IR&5//:S$C/HW 
P2S2F57$%QXL""ATHI.#R2^^Y2'()\QQB"1&"-2);W9YF>-NED!&0E$(3Y<)5'3OB
PZC5?DP^P-W_<S(=[Z&+(3U+28?K53#@GO=EF[F >9;V+? 8Z6JFJ&5[HN9VTU42Q
P2N DP)WXZ%DU3*3G)TMH>J>O7<(H&&\F>HU8&*FT+G;4PF^9P6?:2KTJL^6#B,(9
P*?V^)4DZWEI,;"_2JI9 J"G0/ =I\IE]".7_V"'6<I%M'81+Q'*=&FHKTB 19)FW
P>F,R.V$[(WE7@#&\-]^D-4\G[Q<W$W;*V=)Y#&@XQ4 4LI$P'N)OV8%U_M7CF.,$
P)"J4(>]ML*\4&$28@M/3U^P7=8)8B>4]HH;3Q]4E(%K1-MS +_UW::B\U) "II2E
P>:W_QKX\$!M-1DQ-Z8_4#&W9%27A1=#1AV-D&="9X7S([C65GH3T]MPO,D_2*G,A
P,B#82KYG3\ %E#9?EU3TAJ]*2^R\OP3-@?((\,"0RW-M)#@0US76&;MK*3<MM?<C
P(Q?PV#AK88.N[ W/3X < RBFEJ$(X4<36E,,"K\/)F*X@-DWU&?%'DD,8VGT1@['
P[&8[AWZW/F*_$^D+1C>BRUS]I3+&R2M@<RQ,)E9"!LY0':'EF<:52(5+H.S.5-&>
PP4Y6]?':\@Y,M&J=6&!U=U5)J.7V%7H7@ =M2D!\T;ZA>B -2!H(JPNY^W[F8^?^
P<A0, Z^H%OQ+7!*$Q+ 0VF9&VYX]J/@75V\FL@311CWX1L6WATGB6?OF@4\89'9Q
P" !]0ZM9#,3.NYR[T<+!?0\@3'60S,&*=!.,%BRVIE>SM#\X.$]$D(_+CO-D9'47
PR3/U'_K#]#G'-/$OJG+ZIDJH@>Q1K:1\KK'F$WV6)!/55;9UY$KGK8CS@N7=C;NQ
P'$SWEF?Q'N6+"R,:F+]@%9+[D;>$#&CKQ(($<MHHB:/($DJWJ3615"'?L[U3_J2X
P_K8CM0:^(S,?\U+N??&(_*.8XUZ!A^) 9]<(!-_3?P96O>V(O):NQ^-,5>5J$>'P
`endprotected128

////////////////////////////////////////////////////////////////////////////////////////////////////////////


`protected128
PDU7H_H3X>>IRR,/N?KT7T<0-(GPPGNX7S)K2O6232&=Z/G(,-RG>ZRZJA ?<O-9I
PT'UJJQ2)\;IC[GIRV=)(O$*N-D?ZHP2>FEQ:VA,.%]"LT\00$=BVW.QQOYU1]JJN
P5H>*Y12CWKCB%"J*UD#<C>>!-JK.1I8!X.8,R7/<CN]ZK1CUA^5 IA" $"R1;IT3
PUG1"2':]"K/&Y=^@-IS6&OYGDM&V>V%I^3+.90Y FC@4:4:6+]+L <TIO\)+6^]J
PV>.USTD#6>RS!"G^[VB2S'<MG2)-*#,/<KL:P !)%6GI58KN2@)!N&Z%[RE_J!@L
P?!,/D9\)\RFU58 DYK'$<Y\!GPPJ[*1)EVB1'T8R[L1(+#Q+BLA>RNYH1!,IEOIH
P:&QFLXI@Y'BNM6"CH17#.&<I5CYSWJNA1TV8_YE@B$Q^E?-@\6L3*. Z0@:]D8F\
PM7XC_RT3GSR!9-<0:7813S<2:<TM5J0X-HB\X2^0"5?0U6?,DPDP:5@B-S>IZ@K5
P=V;A5$4J.Y$ECZ=WA2DL'JZUCQ0"9=*N[.2+GE=1W-*<F)B+M3<"C>F6,1@!V\]B
P3=>1^$JJ?'X:ZA,&_\#6ZK(IP*WG52C4Y<LN">^NK)Y7D@26VI9%Y'S 9-K&9K:*
P1F1)1PA:Z_,AON' 79-",MH?.+1I=K57E8\0H^.ZO.&VB)?_D^R[Z_V],=D*=FF!
PT>7U)%:BK>"_)Q%95'7"X2/0L4KR2J/F+CGF)DBEJN]M3-6OI+#%59+FLY2N*?G_
P"JJON;0+YW)-9HA/=_.CE#1=30*C0THT8M%(AR<:SV-(/H(%C/*B-8WH%DSN!X4;
P&2?-::5PI-]%:<5-B N%UYKHJ$E!-L[6T7^H-8$[G.QW^H)&ZEM?>?[D/$$+W[I"
P((MH" B:<8^..$*US\V\1=<%6M*G\Z&GR/A^3O?064AO;?.\B?Z?.Z:>W0(4I'(L
PM%S_BPH.AF^G= ).4Z@I/ES?7F)DA=M=IKN1YW+H^IME\+-2G0]_'&.0*_(-N/M"
PT2A,*4L$VYK]N"0J"IK(;0$H$LBG!B[X=<OC6*>I]&M%L! >6LG=(>*]6JD7]"*P
P#0>5(FG\==4'5?DK+6Q#U4BQ:4O46<RXI40LQRU6ES\ N:W/_K7U1(\?BDE8"0/B
PYA%>&&:L.:C]A79"N/H$I_G#*^@&,7L,A&>.5.!L2V>(7Q32;UDT,1]KZ7HP.&50
P<^7PR6=5'U4-1JWXO0.%Z$=)6K.XT@ZMD:+HR\" :V (S]T,*9E#),9DNTR$VC)+
P(0G8/3@9+JL,NI4PXSO0?3U7Q/?/':?6CEYP5!JG*!5# D[.!\T+=Z0YDTS-6X:F
P&<4DE@U>8 =0GR!0: (=O\=N<=5+U4^66L H O59Q@LKF6G:+JF"CK+*$V?)%0?^
PWP,69L[8H,^%H4"\^V=E1_!LV?:B+#6G5NZERC,UA;Y4!-<.%,@/"40AWG97X\(2
P1$B1F@?2X;'K(TV.'CU786+K%QF1PP=JD&4IX_KELK$_:Q-GH?WJ..SI:Z=T[85Z
PW0\XTAO,P,"NNF/<2>[JJUX>Y^=H.P14H$M/O,]Q.+4O>&Y9:H7P4)4'(1?UUVQ:
PW< I\@.R$V'M_I,9:]8WG$_K:[S9M8JL'JT2P0R)/#XP!0,G6@61K?AYC!Q<5B#*
P9Z]P,A]"]LLO22E6^$9D$MII_A;IW-0":1G2"QHG4[ZT:-GFK<Y">PPA$(8I*\%R
POC<Q[L#H",*3[JL#+G+FV! 1VXQ(QDI^0IZ?TOX?2QS[OOB:%&CXHX_^P<H-PT=F
P6'['&AN.B)UR2;:@'D*'<F$*3A2P>*JS.9]_9+Z9Q1N7^<Z /LC6$"RMGS05I3&3
P0DSL8C0?4CDR)^6:_@.A2/*?&&.S*UT])KL.!T0I"X8O4Q? K"5+7E)['MLI/5C(
P>XNZ.KEB2\N4GYR:G7-U7[\:$$P4M,SM*DB<05+?06_ ,Y!.+/X][0DP]SZ.:F6C
P;.(^E5*A?D7!<;(MX483Q(8>1NT1+C9VDY-DGKEG:98@%]@+J)M'!=XIP%IZ_I3;
P67D;[/U(/@^8._7;4&DE&VG0DL_^#$E>PFY/2!%TA":)1&F[B/J$3NNWJ[7:O_Y1
PJ71I(V]HQL+52(V^N6%_A31DG_#KQ.QH(%H[=N .UN"):Z0(Y_(Y*?6TIF.B\A^T
POW*A*!U($64]WRSF(L]A,@%O^M/>O!3I5$>XF3N.$(.VQ  >G3HMXV'YDL:"'?B#
P.)_VW_S1OJ<G^5QL;XKG"#&_2W=_YSD>-VNG/P%I752*GB/HVP(R!3I,PLT5PAC7
PT.9+?B.9':PBEW[&4-$T1P3G--:.F"76\,0>RAUV9?K3A6P):"BLV^W$(0#-Y&#Z
P#S#C>[E(F6E.AT0V8A]8'*#C4/1)_K(5+*'GI_+N\5HVCPYOPD@1T"'TM2#D>"#7
PX; )]?R-@%(<\Z]58;_)6*[<Y(U4>#.NV9W$P*=Y<D<; K<>*C3C6(_'3MT53\Y&
P'H> V)*:GB7.SLE)V#]P!U\MT6/.H3/"2X$+U=$(86)N').!^RYO_#$>9GZAPL=#
P\9Z,"Z[$;>:@M170B@Y(38R(*7Y:B]*=DNJ! ,?2CU/B<CND\Y&;;U8B+Z+6;HZE
P#%4NC!ZX!N-4D,?P(J'<LG;C)8A<0'53-VKQ]Y3-(7^BIK5V=2/9K;^GIX<_R)Q;
P-57'9!\;C <1P#6,[,HKD&*O?HCPTSK)U"E=4*Z%S#B >L"V=Z:6@U.@1@62(E;X
P "LW!%+F[,[_I+%S7OTL?Q@.M[RSXT=,PYM %Q[ZA9=)0 )%+OF [?'GZW?P\T+>
PX$LBEAM.C9T-I!:MIS4OK S#OQWV^XH21=?P#I>FXAYN,8.SZ7FL'@;U(CNNQKXP
PXD/)N/LGRZ^<"7L,6BWA^(Q)H?.*7 2[NA16#"> 73[1S1@M;WTS@-+I('B-X\N7
PLQ<C#YTIH7/6_,X2GD'$X_V;R$0#YRFQPCN&A7L[J,/H]& -#<5B1!,H4L."FL=Z
PE?P"?9/#'>>?CH5F"L*[#FX"RLDMO,B<[_H[CIG+CARY,>"C_8%PWHM*)EYT%C82
PK3_?  LR9Y&Y_C'WUH6/2K.EL>TC !Y61Q0^H:KT.+#<_@NOZ.$5/54ZB+I5,_??
P2C0!M\E-E)5@QZ?%QHVG"OLCUO*>/S>!Z$8H>HB%LZ$E_'H-#:/B>_<%K=Z^B\PN
P^L4PA>"FF%QOQ)MS?E=N*]!7M-ZDQJ[B05KJP;M[RE1F]<B6S'&&'^0=MX -6!7O
PLD5X3&=*!XE98=_3+R[YER;@NWU6G'665I$#@OC716BE-W8I_\VDO<A9E'2:E3-[
PRS+H"%2'"G^X2WJ0NURKYN1#G$=;A1^18TO)R"V@91W6K:.O-DLJ#$+.%TG6@\G?
P."-BC*<>J[8Z#VW^753A!3Q)=A2ZEHU(XGZ!9"VX,.._&Z2\XR,AUCA3FLRL6%PO
P;MRM&47W?. ',,'T?'R^SRVNH?Y5(@Z*/;+%TNBUA+9'^9DGQ@DS@NA#Y9%J5SZ"
P9<35%;@HX0+H?^1RHJ%(5IU:P&;:&W4OB='I7.TLW?)8]FVEIHC[HB'T!PA=VK="
PN\X:5Z7IQ6@'0D1\0>V\MZ%'FUS K:;>GA?#2R IBGRN]P?1Q7RPFZD'G>;A8U4\
P-SFP([6)QV99]-66!W,@\5^4%JAZ8@=Z2[D]_6_780:[03@=*@6.;0(5+-7HWND3
P&VR_M0%Z&=[XW2./9- /TH'!3LUB?XC*E?ZWB5U3UAV.N&:N7(,G(HA\_956:R:O
PTMJM?0; ^2<@$-CRO3K0<RP/M];INWG%![\1EY2NQC]1QP-!9B/VBI':$XLR9D=(
P)1'EB N_A2;U.M2AXC!W@(5FWO^V<;RO6H-8-B'T^3.L 2>AN15GJ<)Q,D N7;9>
P@4VVN5?#O="KA)?6:KZ:U<O]*R7JY'&>EX4/G7G4D^_A6RS<^_ )5V73V.A:X-!D
PN P((U&3Y7QJD^"UXVZ:":X9 CL"4L]H[<&BJYU'LU_2XFJM[\AH$ WM3Q-:.($<
PK')RO*+14V,7&>;G^]_7]ZWDVS93[K#/0T>VE2$[D?A94%#C)_KSU,MMJ/(F!/+,
PGZD2IM#43]-M[KO?JV0:-YSB8^ES!]F^Q=V)R.RJ&QV@E1B$;5LKP<I!&SC&*FHW
P/<"]P@VKA*LQ:E^EGV8&^H]#/ WS=)Q,)9ON8P[(1BW>(Y!+@E"#=I 6(>[X0L<Y
PN%>^]G$[#65-C9-@@26]F /I3B@!!/KWO8O,4N07="Y)AAW&BL[+2LPZ;*6YS 6.
P>=[U?A_RF<./[=8\^!4IP84G%.EU4?KM1%3)%Y=B9#SS<4H!_,)\Z A)0>K%4\5T
P_XG4W4I9$9/(ZS;^!?KPC&X1;/$%L&O J:F)&+E$TCIZX#L="%%P)*(S(ZK/N53S
PQ;!/R>YY>?VF; S1%LD?FOCL+>K_B61J]P>5>IU>O.G)[B:X/P&N6];K)B';_6DH
PA\5M,WUHS#<(QRH2LF8.>^Z5MS;WV"88TX^S[@/@7)$\%<#2.5GMI;<G7V*FU,J_
P@JOL;WE_+W&7D\ES"W?/Q%*DN'>-B224_UL\-DK[#GN/6LF]^R5+G0*E#[SF'&EW
PV6%&M^HST+8H&1<Q/9[]Q83$9EP(=T4P4[QFTBH3^2S0H;)[NKZ//A8YQ27(\A 2
PC/B1&@.@V<19E(NVFS]Z>P:_ZWXQK!P6(W6XKL73-R(&U 73+5G6OK%2"/3T?$7^
PA$CN9%:._[OUB86D')NB[]KP^6GHJI,NIR;!\RM&A&'(.;53HMOVZ#')+*SLI^=_
P A*.'D2A@2JN2</[#&/FEO:(\CIDLJ\^/&9"O]:EA9J[@S$+6;C*9#;$_&YKE$QF
P8-^]+_&CF(-Y&.,8=EB.E 32H7LP>A-[/+3'';75LWJ.5PQ:0BWRC!/^!>3T*>O.
P,_0$<1XKQ@SRD6L4@TXM&XRA&$)E,,IN$UW!<_XX\:0Q@(NN:*WUY?!O(H4+@*+V
P*$@YZM48\PN>IX,1BK<$ZL2PU$YW:'T0JY1J+8Y>H22]>Q /T$T,"GV>FT>PY-6_
P\?]6W5#.SP7+)$D"R.RF"$KD;S\T@A:_BU )EL+X30-;-G;"J>Q*>P^&^&/L05 X
PF=:Q%G W?%G#1YF#+"+IU2(GU9"3Z+G4 5WNGATRW>KYWG723M*>>@"GP=9T''0H
PHE(DNDCGQ1>:B:A[$=**IF<ES:!NV ?8#)LMQ(MQ=4!,A8=@?5+F:JL-6A37*9=T
P\8U#4N: #XYE:2UE%8Q\07\V%?SDK405;U ]YXUS-1S7?=**,[2KB,:I!$-P._>R
P^XWTDB:^D;$\[D,/X[.WNPY?Z$2%1,1J$VRN#B(3NB0.ZLLF]Q.9).NZ.IIT%J9E
P4:1V?^GW=,02M@8=\AE>DP;Q8MF]S,>6<;D8NKJI/(<5]@6$LHL_,Y]Z*@U!(:;:
PG,FRTL_8WC2[]?Z@]O%:#B+<U/^Z(MGCYR8.,3=='E[]R99GHBD#N@NXH"9F7KG/
P8\0RYC6=M",;U!-F9^<9_B/=U5P/UQD8)9>:( M<M:]0C4_X!QT';UJ$!M]PQX68
PQ-R]5=':[UTBNLV6QJ%G/PO8R]KIT/ 7'@ P:;8'%&\Q\1Y?^S@BQG+:CV,KF]RM
P_O]FL00X7$5?L+96U.@- 5A5L'[[*[[E^WBQ'N][]%93SD^^$3D>RT8'G_7Z%K^'
P!Y 79SM6XZ4N+[),&,"I_FWCKD-2BGF+&T,5;. WP34<J\8A5$"!)SD#FR=2+ES(
PD":@@-L])338>]C.U;!#D=[V<;WJQ?5F\-XG"6+D1O6< "E2AB3!/:CC56J%]!J7
P"S&(Y#DFR3I,_>P2=_FYH&!1-8BX<!/M %F+U:-M:9+@ITE]3"F_1O(+O;AB8[S*
P3<8135XB17S^2(R1"S!-.\=B2QU0PF<U\WZ[0E$#$#*%L%'0+_CD/$XM@(8%>KQ6
P*..-/2Q^XDNTXMB:03=&7#U_( !<311/N%_/,76OEQ9\K$J2O8\06,1O"  )KLB^
P%6-F$*0;#47-'5$]/B8MU2PT95SH=[^M)>6D-?YHBP2V1#:8_FBJD01KCGT)UZ"-
PV^UH^.'3M%DU?!O<5]G:'VF-WY>'!U-I?!S>9>2 !)_J_U)5M\=3^9RW$"FPXMHT
P/QOM,_"H:3B0 Y!!=%AO\U&W[" D A7G'B&\'QSM#[.T!D\^["PH<,ALL8?LX#X@
PM2RRYF-K;%:Y+Q<8:_).X]>:%-F8(_(7'B]5=>/<!PQJ!EX8>B>49#/F4)@]2*/L
PGX,=FKH?\D??_0(_]3,LF92RO]'M%QHW,JOC$9!&\ _^1;9BIK'J2+<=/0W&WBLS
P$8\UOP,2H%7:5M$V:6V0G8K/V"T2I_\!2#4EDWL^'M0+W98^/;S$?D3+9V^T>W<!
P.([1Z LD![A=4D$%B;# D$)S%C[ZM^BHN-BUH4,@YMX;$Q32QL4-8.CRL3:Z3'!?
P+ H)=\O<@\/D;V5#*ZK*_DRWSC"DN1%OEW<I9WK],+ A83WNW6N@0-3%7@VW.*A%
P0*NF<3;\F+Z\R(C_LYLCYZ$6^M]\60]-@#1J%17^7C3=>@5M"#.T25Y\)!%"JCZS
P5A< HIVF;CNKO09('NN6TGT:^[H7:/:"J:+DR9H%D>): QH@^R*L<AR&3Y1TL0R%
P$,%A,")8; .C3U6+%1=V3F]3QAD*MW4#1@B&:=Z\M0P/R?(K*>9RFQ]+(UJ?ZUGW
P;>KPQ0(!EV_=WTN\!9ZL\\KTVM19>)>7P T,/<^-J)+.0OYJQ6#!A&]UL >_"G(C
PP7K\G*R_3;%?W*1FIAR%BX+1[G?*8L'^)^*6_CL.?05[8R22:BP6>RZ /+XR*"V5
PM:/Z4JLK=K*'.;/@LASTPMO<]$!_D/0XG3Q(.WMT.)SF:+J%#<2FZP/3YSZ!.)C6
PMH;T[!9,G??DI;FE?];!][SVKQJ5\+J<C%Q61\?%XZ!ZAJVXG%E]%^8#)8"PAPNE
P'J>4>/I8$N:S<K2W[C0M!WO:-)6T;6TV27SP :PGY3K8AK UKA^+>B-#!WI3RM?H
P80ED!O?II$?N\L[PA>ZF?::'>_H(1,DMM-S?9%_NEPTAD?Q1[OP(;CHK-=PXO/3T
P7CJ55OQ?/FP+O($:P);7 U%P2=S!3_H@93'<+S,"=67<"'U%LU0I6?]?97DU&_9'
PUL<-;)F&U3*=J+QV]&@<FI2IRV#&2XXMU)1_I5%]K?(:X$%90#$NT.*EC47TOKWC
P?3F,*5:0[4+1&T+QTD/B9<MCGM;7AZE3I2VHJ.11_=B&3&126@%5\-=_WS5V,%_W
P7,X.E1H+)TX"PX"8?S$5GQ\WM'6BGLW)ZLG/Z92MK,W[NI4L_?R>D\[#KR9EJFSE
P(]6:EI1._0'SX)*+@44E,P:??)ZR61::2MP2'CD;'LACK^NN=.*S>4_W5FKNIHK[
PP2'-SX?)^FD<A@@FFOTKXX7Z18&R<?SP4.JCKE(6;XYO/G/JHXWP*U.)-DP5002(
P-IEVAY"9<= OX$5J^+7&#T<L7XXJQ.AU]!'Q4:H]F%R3W"MU?U^6[<>%J$'N=I-4
PQR7\GY*7\B74"!'V9%DRB8B+^=)N8#/);"'O3:R",Q]<L&=^%2@+^DEJ77J\T$M"
P\=?XTX?J83=]@#UX:F _U:7>&@0G))L02O(-993C>S0R#\MV*,3M-BCN64>$5^"S
PU@([IB]Y,X!!00@Y]^0Q&A=58-@+YPFCMJ2LU3@.:\M6ZTL=98]6QU6F47L;WVI/
P;.?Q,%0\L53.;H"%8&_RS9(;XB415MV )%'\2>]I[DT4?'VXJU.A/U?Y1OD3-?I:
P>2^L\ZH[.:5C4.I83N&?C7F15# W]6R].^MB93 FZ<_U#R$5ZG2KQT<W$X**DYSX
P(YU!OH&2*5+@Y)/!3D+_$R$3%P-YZ&,:(:53MX4#=>DO*C/NZ7#Y/3X\00W FURP
PUJ3 <@M^!LIG;,]H*M1)YNZMM[&[5JG)@="2<BQSY5U$BCO")&I(; ; V<8>L^93
P;!>S:"DJC:+;IN:HE+%27_-6'(%-Z2I,!:=0&/#SW=$:G ()0P. (51Z\5+X7 E&
P[K_#O M7R$O$I@;W6B;UW>15X]?N"+<[SO:LJ-KO'2B<!H\JM=)D0ELJ9E!CWW'Z
P8#8/U?I-'2M7C '$Z#YGUK#-\#WU#_H73Y%0:]%(&GA$3N1T)P=BC)\0T:I9-"KF
P5')5:10^_>3E?=#":M@P\N?96OY7>OEZ"G&I%J)+K#A8&'KTYRYC+&(0)X_1R/CR
P+9T7^2)ZU.31;((M2^X>F.&&!3@1CR IN-!LZ(4Z/,=^&YT_1_U45E?&Y?*XF/7U
P22>,XI!^)S-TYJA'R"@,2?6J4.THZ+&A#6,4OHSP,.5+04I3/U$FI&-?OU2;VO-R
P?2YBZV,W06HT)W<GOB. '_-.3\+T4=[^UH / QU7Q%JX\1.OE]%;W'LK*L7Z.S/(
P0^=20MI*=PRB?C<VRJ@N23"W/;QCGPFL$0\KO\FC%<$W:'9[9/^##EA<Y'W*@(KZ
P<UVY")L#GDDT!\[E9SFU=2'3^/?^)T]@U=,8B22:Z^6=<H8= JD*U=,\IYB_$],^
PFL!EL *:U[OY 9)^PV=*=YVG>IH0L%($$N&!5@3#,Y&'0V,+ZXQ%^C%Q:D=H>ZI6
PG-QGLKO\(KS?P7C65(B<"!93"W+33\Z--H/#DBU5]D.D-W]:X[&50E"M=0)'CE/5
P,LD07QB_0E)WT1+D4N1O_HWXGFO9\4S5C@*+-Q &PJ;40%H0_GST2'IYX71';976
PM7OCVP:4&QOMB).3"@V0<1U%7/G'UMZ*46<)N-)$[O'B@\[_*0>4/O$4JLH&J4X\
P;-9>\YS$=?&/4_U^#G#K%^\3%Q2GO;ZL=1"  4EA:%*)?:N;N7K3;F6DJ#-W[%=O
P0(?T+A2I^NCCXNA.!83X# %Z;&&*!  *&[S3$1L-[_\2<F^"42DZ#!A$'KE1;H)*
PM (H]0A!FM&C&;:*CD8CXJ@C'*M+KS*<DW3*-4YL@7S":J$?9DF][L-L-EUF-AJ\
P *3BZ1ID>_),$*6I9.D.1F&0M5A3;[8A<9"C:(DPAXY JATS?7CA0*:U4EA!"T[(
PQ7K2+E*=_!HFZF$2BSU#"-'1OI$E!4P5!9B'IAJRQL^&NECI;4\T/)QXA:R \]>3
P45$8D2$O;WD4 NS^/H^I+)S5C!\A8;G8@^Q)Q&!'#R5!=3> H[18-E8MF$QC4KH!
P$JB+C.(UW08)6KJ)!X<:K/JHZPH?JG/"@<K'A_4\KA>=IQ4S\RJ*CX"UXFV:D".T
P!.\N "67)!ZKAX6FQ:NHSY-AHO_:5]-P[*@QQ:Z%)1U(<EC-814(Z%7-6IY')57G
P4=C+E_&+,_79#!B?7[2Y#B,AQ59K.V[)8+KP. X#2%!'NSIP><E6AE92^@E0%P;4
PXTB>Q&%[28\WWDV::]B9^F$<H&]DU\1?A^ ^B)8(5)\$#]3WHDG$P"@RMMS!9,KO
PIT9%DS$?V6=7A(Q3M5!?E;Z4@.!) \A!GBMK8:INS_*6GO_"^P]LBY#NGJ<K!+S-
P?LKXC;]Z-P?MX>FWR\9RZHHR"X;JM2'$8IQ_YU.RY2&YB4EQ^NW7F.B0.^6^]PE4
P <O04L>^I[J9<N[9ZO%NLRU?=N!R,K7> 6FC)-1)2<SU_!P;*)S71UPI_TB"N2X5
PC:"/(?4WTGW#Q5Z-T"YTG)+)=L?1=@&Q-]X'*O;9.ME*%<\H5>83TE@ZUYU.?L'A
PHAP1K^:61DQL":P2&K[J:)+X)9SLT,6G_([<1Q72ZGIX(@_7',R_-Q.?WIP);=4,
P6EDWH;?(IL*U-H\TZT[,'>DBA!T-4=C7$.Y&;+E5Y-$4.W?"YFMP$6^<^+YEQ>4(
P/%BNQSU##I#\4"GE GHRIF@J2B5&JB'SJI!R+4S;Y5O3HOL6B@,I((?+ U,^*!LC
PE1>6EN.>[.?\QWC%1B6,-$KNH_;D XZ)CL?^-2Y]AQFHI.X8/FS@EY@SF6_(N[(/
P3J!1G=%??ML8M153T.1J4&#N4MB&FDS0_!M!,CS8N#%7MSEYC(;S>89)*A\X3I!T
PP["7<1LP(17*=JU:<&G,UWQ[33O1B%)H-9X#+-WT.Z:I/4)7M8&=S58'(/V-]K8V
P?@2AM//DZ!)F6]:'I#1V=%)4JJ\@EELQV;9UR!FXXX#?/O7Q<(P8("3Z$9RS/P60
P4];$,HD(N#@N]314F^UXH8C/4(E)#?MQ(>[8PB9RX66-MH&:]*0GX+5&;G[X43J+
P _'PK.*Q=6CG*F ]@SQ _T#N7&_+NF(V0R?%E$X!+4B#,6;REPYQXT*FR(0@9[=H
PB3=MU%"BEBB2=>%' "AT9W:BD\ADJO*$$7:'5XK_XKFMT7?2IT=.ZVG!5L1G9>96
PKQBT1P?[&0!:'B@%0X:5T>/:["=ER3>K%3N.4M<FUV7>SXLJ+<XS7_5U_%A\AV3<
P;4@[-&+?8I[:)&\@B^XC>G36F<V=#5W5'8FDPZ$7@2G6?PH:4N.;NY'C1OO!=H_P
P[#3=X^+8F><G=/*%%W[YQNL^JL6XX!Y;_55+V7%-3CYGU8SX,F=I)B)3_+,HJW3F
P=68!Q' 0+ W](<.N)JT<Z"Q0<Q5#)O$4XU*G^%WFPP*18GKEW94P]\XD-3IHK.,N
PXR6W00(/1X2CMHD*"3/E.;8V>5B:_&QH5Q4#J[CO5$=U#<8KM=']J\I0&B20G\#-
PD)SV\E)2MG$ BUT<X_P]H+=P4)R=&UOEH&$H$N1;%F 7^J)XRNMM_HZ<(L#[SQKS
P7,SOU'QI&O/3WKV#%2B&R^Z2_PU?.!1<*7Q-EKGKX<S2#3([H$#,9P9&W81>;[3Q
PF8&N:E,$O)XC>4\ML6#^$ NKU0ND*29)$<VX:K<&^P=)IYY(JCX?\:<(AV.$A>)9
PB+JZ/Z)&VACC&<#NTJBZBK=<%Y0/&;(0_,"-R#?;DSG@*U"L@\#IMI3VS@E".&M"
PW-\=$Y9(9"$(#&@$:WJ]'I8SU?\NHM=R^%'M%N,?>E;HFI9J24']GL> O(W4W$@3
PF5TL#'T3D0)6N!BWF?U(8IOVE2J_>$R]XZEI0WM%<33QZIN\>^J?^(IZ9E)[0:?]
PD+?^BM&63M]O/ \?GM0N^)9A:<9Z/.%@77+/!!XEP"ES9]M)6&RR%0#L.";"Y'10
PN+TD>$N#J07G;!0331[PL/T?_+I(779X9&3IMR.7ZR?$_T2-@&3I )(USIUGA>,S
PO2H6$)#6I ENJ5_JPP2I;]%N;%U5^:L+[:N](PB>Z!TE[]B0R[RO49D[M5#<1YU]
P(JS:"K!/-X,0$H@A3:N*E3%]?M(:R@!,%>G. -CPO%^IX.H,-+F^/7R3QZH\VUX1
P^PF-I:*'@L_[4L/9.Z3$]I'VRSW0-QRDQD-GGW$$D?'93LRB,G'3SOU=J+6RUF,@
PFY#96C>S>G"ECIN$TT9$76Q3N"Y^O(^@++RQ:8$V,[AO^&2J@>]Q%Q*5HUY%I0 .
P0_4G]D2KXY""/N[AELEU:JO/[2I^#;%'5'7^+R$0[6OUK3Z2FLZKAW:8\\;<YAHC
PG:.?T975+K^ #C-1F\,##1O9/*W[\D^QTM:<@+-'K1463_&^F2S8+";$9H2'57X*
P0]-1&8'2@TY!@(Y+]C#+Z'/735LRPT<E*C\+C,FZQK)2)UH/Z^&\R9,]=LQ%IUNO
PEB)] 78KB_(([-*ES,(9+58/9\-XA6%HV2TKQTEV,>2X13)Y=QJ3(=)<B\&Z C&=
P0LRS")2AULBL@?+UHDDCE'5&<J%,/^D-W2$0()1&Z%35^^YD4E>,K1?5<4>@G" Y
P']H4E/*$Z=(U5LH7 IZ^P/5VNI0KXI<H8&;0Y\&3/9';9K4\!L/OA&A0EKC6H@;-
P'56X^GJBZJZL=%?6GD;N\#YI*@;5I[7*UI:+K9<&!4^)M0-93M(<GVW"$YCE/R>=
PG'$M+SK<&$;VP/P74]II3J_Z2F[#_V:IA*U>S34R1*.*PSK[)0R\B$L*^7 (EKE[
P5Z?+UINJSU>T:$RO[-:GFS@BGJGM< 0U'I'=VY:[WD)=76>:#9EBA,P'6!)+647D
PW?Y/DPLC+&.!0LI=D(W[M1]YL+>G9'F8 #I O(4G:XH?8KM"T8M5K.)-^&(S(0C_
P8.-DY5XDN1<>LS_3J!6CK#!1[YH7.M9V1]E,0^?C9F:=^3B[I5.] 8T6I+-ONCYW
PHWE:3S-U<<I09+ #@.J UKD,$4)&CSD?*QXS-?[1YG&_A+[S/G4LO756(>P@7@R,
PNE+@97K>F;K7T\% S7;D2=$9NG?05T34YQXLF,;":+*RZAH\8.2%#]CH48= M N(
PYIL)0GIIN#OTN^#P$P+!#;XG;3-P7(]/NY[F&Z%VP/3-X!;SFL"\5@T?%H*!B97(
PU,I&[+9PQY?O <N<Q7;$"R(QS$R!G99O G,50!55#LFNJWP2,O9+49?LY;ZY*Q.%
PXW.6CL$7]I#)/>_?^C I&SY,_&+H03)#T6=4&]O9NK6V".R#B$?3\5%Q24KZ_0*H
P:A/N,Y2L:@KKVPZ1\]!:EI<FT>1GOGS^^);Y_1KY)-#B#Q;]:+F+JX-Z4S?:HO''
PT?#S 7;OSR/6(_^^MA80\G33T&?%2,-4)E:=S[0:G -9,C':FAC43:P= D2OHMDG
PDGQDJHY$?>A]HLQ[%[KK9J]A1JU9T!1) 2T2@6=5Z%?;G'D[N)J4;\FJ_Z?])1L0
PMIFSO_+948=WEO>"A#<UM)-0*@^I]R,.^(IN]X%*<1<P0JR "NV7/86ZAFB'SB[\
P:C?CH&:4DJ\PT=HBF\AT2]EO?.^&7YR+V:7AU<K(\3TBL.MXZ"(M!YJQ;;\+D99$
PPYX"]_]_&!T2O.3#VJ.5.9B83S[@X)OD"2T;SE"V*4*C!9,<?DK-!;J-\5+$7E\^
PS_E\:Z!LPY4DKJT_/.788<-PX+([+5*NF9:!QG?*< [(FR";LH@2,84MT=\80":8
PP:13&<PK0H;CG?"OBM.;]+JX+(_J[9$HF %TE3 Z ,LE6?;BZX&KR)P>JRFEV@6)
P4_>ZM1"^.,6/09U<PR^P,;N3(2QL!6LH-P[UEF%UA6VIG):JW=/O@<PB@8'*K%WJ
P)L"'GTLN((]9.WNGV%YEXW]C2.5Y[7)N4'38/9 80F;EL-8/V!?_76@+_X>$9:N.
PKM)M;\!P_ATD227<41EC']<:=*FI4_4 -)'T1W>.Z93Y/_4"C\:,?(N*09\K@0P8
P3*I6YIGNS?ZV7=Z@/) <67YSQ1EJC1V:=P^;PEZ3B%2"\#Q&(L_;FC%PF !_K)PS
PA/&7IZ<GEU\96BJVQ,=!GIXX O^&O1GHS#LIY>Q[H6W%1.SDB'(2/J1]H=@4D@ G
PT.M"_Z\@@+X<P]?U,3MW;24Y:UQ"*KWG*N%9/;>(L+6D[ W'4.G+0&@__3S\096Z
P;;G%T[,7XZDJT.A"RNP"F KE?RD+"3"&Z_N36TKG,O;*=8;;[BT[%1;NY1GC?USW
PN*("'7?PHBJNXIF?0!(3,K:BVVI6,]E%ZJ)K.2_?-W;90OG.!&K";&*<!,N(5WT 
POSZ7WFK2:A/46 YWP8H\29;>M6>1=Y$@#H<N\M7=U?LHDFV(UK.A4(<%L68:64Z 
P-/6FN"A1K_E[P> [E; V_]<8CG9D77)&0:?#SQO>7?V"5=DN-T(+B1G<&X#\^%;<
PO<#51]CA.QQ]&423,5W;)C=4V+>2Y'B[U84QQY9IWQK<>.8<:ZG3()5E!$8+)C+S
PU#G9]6H3@N+B:I,Q=B\I%-5S%^-"#!S:\,'[S )CIBJ/O0J2>0F<OW7YF,/P^K:P
P<9+L8RCQ\+1!2^@OLDI0?J ;BMDST@15;7*+X9UC)-A7VNPAJV;B6C [),BI&!Q;
P%+C_.!;9DO8&2)+L.(10"H67')5XNAJ1]#/(-/I>8^74)XT<5&$I\U\CM#BZ*/)2
P81\#].-(X*&KY-91AOX@W<=YCTLW$O!U]&J-W(4(6K@A;QX&A<-+_6 X"+6@=J/8
P3S.-B%FZ[DABFTF6Z6]6O"G2;K3/YRSE#3^"A/I>$6?]XU:8C'=UK;G[9)P >6:8
P92H*)#,SX1=.J?)6L]<AB)"4>36TGZ\0"K..!5CF_ KC/R;=F0=509G](!RXY]^6
P%52$S?!F]18\#=8AL@^F0C&<L:<Y9K)!,Q700[RU;>9.\W^S7BI!=:O D:?QV_&*
PJIHV2?AD^3A7RW6>_Q;US[I&5^]2 @KM=$&0OVEPN>QSBJ8)/RX.2%KI8@5_2JU;
PM 7%7L6T:F$NL_IVB3+Q[TBH DU[1M5S4 <D-Q_+HF(X CZ?+"Y=MEXYAG)SPX4Z
P]GGFBKY/E:47&I,1\VR DU=],PT_4P-FGB%F/"J>O/,_=T*H'P!"WS/T$:-"I8P0
PC"I\(;-=65GX0#,ZW_PY=+P'5-U-D""Q2#;2TXS#<!AVEN:-<6KB=>]KG6R7(4/@
P#<IS:7W^H4O]<E6AY-SG\4I\I%TX"MTIB/X]6)MY(KO^#KY'<,PC3"3K'&LU0D_^
P2,"HF;J:1= ==XJBR5)Z0;.>3A];6FBU5^4CE\5CA?7R& /<) (7Z:1-DLO3YR4 
P7_*N&UT>G_J/]S^=AB>$^2(1,,T98WR79E'WH&MAH*?U..R&LU9U)Q7Y_A=H]@@Q
P0DR@.$T\D)L^[+R;2NZON0[,R$7&K/ ;66SN;0H(NF\GG(MV$._9[/*U K"<Y4,:
P?!NAA)*#M^/,=H*Q9KBF3S^8 XQP!$/JE\96;[G)?RLU8/R.\J4O!XP(H-#+4+U3
P*Q"/#*OGYZHZ65C&A>85VIZ8@WSE7N].-B% HTM T^O[MQ#'2$WS02.^:<_DIGJY
P[$9==@,MDA0'C+"7[;U^F(92V8>P[7)8S?C/I.-@*S<?!'#;\%PCHR<FF7HE$7C0
P"$@<]43Q8(>#-4.\(PX;O)P7.RKI3E&44"K>T8TT.PQ* ,'T@O:>SQQ(BGK1CX$X
P26'R2/Z<E<_X?*47$00^-L!Z%K8G<]I4<.=>7+C5#,IO^CH6:41/QI**<*55;U\8
P4"48>)KX%6_C18X8D<D9-.CU404N0D&'*B-& S$*/.^V!4U(ODJ:BQ&#8B3W+O_M
P*CI/S2@RW&%=/&8),5E>'90HG3B N6O0X_4S9O%9A3*;2AW<TRJQT_%!3AQLTL^9
P%T7_]RBKBV2(>;,HVT"8BU%&W_+(0\1A&'&7)!1(PK<CN?%"VD(S3YFKR9(6 K+?
P88NE61$(&EUZ7;;>47R6$XYY.VJ5C_%-R"]>,"SZ0QN2_6#GBC,]73I\QC A#Z43
P&A7W!+<YG:U#"Z[MB3)TBD.Z=N0V/'[=!<)B[/X*-E4%$<+E50 "2'%L_&K[&9ZP
P@ .%VQ>$+XJS48O,0<H7,:MDQ65E^J^; -)-U;$9+H"@9@*>^'%8_'SQZ]^F#_'Z
P*5$S@3== HHYK)'2'?5#KY^[$7CWD.SCA9(O5AZ"2,%Y.M@?K0EUSG;6:=84>5M^
P<[WX\3=MG,:OTI5I^3%29=$IU'F!'&6$BOXU?R098,QMQOL(-0V!$API99Z:SL-$
P$0%UH+<&BGFDE\QU)YN>\+EWS-IXP8K<EKX-GJ49D7?%)8Y!,*UDM%: 7S?R^QFV
P8NO5?(;!1L)G$H+MJ=R-*XJ=IO7R]@+TTO(@F>!W/-.AZR\@@1'=>KC50AOXFVH5
P-D43=N_2SUT%3*UA\4.Z^.EK0I?>V?5VAL@*+Q@O%6UU!P_3=Q5XA@8)NV01 9B$
P]7*3;PBX!D(&4]LJ8&N$&M6;92KU;(69@K<J5IT/OR2V$LRLQ<]M@SAWIDHG&,+/
P7.<KZWGBZT\W<>3+_.!;_,$C[XWCJ;SCT)18V_(]$<V'<<]'97!Y1F@\+,&I? 15
PDC2MM0_W95$SCV*<*OK&GJM(N_\Y>W[RA:FI%]:<^-:!<\$+M!]*0_J%1A=6H[J/
PW;'YRFDI5QBN8]$Q#RX9DAZ%S"LTOM\L<ED,TLPD4Z?T]?XNX-2^_I0Y2V^_NW;7
P(C$FJ,Q#FX?.WJNK]WM".6OF>56%QA<C/@0#:_N%]2&^[A 9F[+@T)B73?N6,;Q@
P98P%J*$RKCL?2J'IP+:-OR6 (>Y_-;SA4.WI\@)ULS.JAH9>6R+L2YSQ2K)">4*F
P6<R/9]ITP29R<07*IJ9N-^8MVGHEP+?97!;D,:?F)]G#N<!A53[9[HNS'F);OUF*
P@"HBVKFR#,#<F:$8.<1)ZP]W$KQ*;*\YQ+1?B#>;:B3T.R7QYWE#WE^MEF<5>OW?
P^YE=>I,=7WEF8;KIN!UH"6@X+)#,MSJ4IA_:^S.XG-I UR3&M[<$1G5&0K!*6(WN
P38<#0"]X'''Z.J05Y)[* 04S"$'75<)!C?F.W.UK![X8 '9A0R.EP-6(PWU/4'/@
P)7\G)HA0B*MHJMG]VQN6G1^93U)$1CNI8V2F'YOA0<W<)=.PPKDN%9(\D,.&'O^1
P#&N^I]!%_0@W",RD9Z#@(KZZ:N=FMM^+ /-\J!!%+JVY".&C"DLFD8,A55DH2A=A
P3GJ2.F21T$(J[( #(;EB4IT]X*VTGST&:04*!;JG+OV ;R_4&D0CJS<.9:,EX.LB
P\7GPU;(DAR9(Z]F#RLG>XKRG[0[/L^N;0GG,]JR,;YM2P07R]'F/^$-*&G0G;:1#
P-O<AZH>!55:YM/T\/ MLJLG%-@Q\Q&]DH@P0F#D&W8[EFD3)L $7AYHO1R,-4DY5
P=TYQH#2ZBF-K&W^9.=TNS8&AL5] N0# W,H="8M^2JG)]X1>3SN6M8]3W\_LI#\K
P8(,C--1O5;2Y,F1C:J%XK4^IT_>8_"$]N?,@.GAX(MZWK-"\;7J&T"5_EQ!]?[NP
P)\K@WYJ\,HUR=]>$=<N#_^64.JH?@6"I(1(_CK+1GP)+ D_?/M+:4T-<D1];W9O8
PO!MX302N;0(#8)]"CP3=Y"#NX/?]CRXAR9<E41;]YF="665]=I_?F.JS."+H&9+A
P*R2J-R:E\8:UK#&^J'D2U%Q8^6VB(DZ!(YBDGW1)F;78E66FZ*+C4H43<C\<5'XV
P]E[SSZQ;*]ET@$8Q?$W+[/FL:,;PN7>R=/M#B5TO['FNW%X1E= G"4=LI]-MEX2!
P*E6\%AM2Y)+H3Z)\$_3$!'-U#K-&&5$7X8S\A:.KQ2HBT>$]$8S>BI+4F7JDI,P5
PN9HI1\=&[I9H0GQX[1#'<-Z&QC'^QO!9LA^,W\"[3  ADF)$^>'VP*AQ\!I8=)T)
P8]DQ*=5Q69.1-T5 %@C<E\$]D2)K(VR&X"SBFHYY)_K.&+O1?[EMH>+CX+.0]7.F
P,Y7SDZ."G$JSYLJ1?UN:5$IF3X;->,G +W$;JJ>9'V46/2Y.[9H=W6 =EB2S^J:F
PY#G^[!B3W-QS%K6$M*W1&],>*>0GCP-<6G$% Z"51Z2E'<&;[V=,=K>(,G8$4'8O
P1URD_TZGU[OQ,^!G +)/^0['W]L?#0I7L?U*LK"C+3U(XIH5+M:[HH'2VNXO"N 1
P=8D(/:YM?]0:WYRF!# @"8U!8O?5,LDII)/8T<$&@TFMRF97NQ@Y/;QR=]TI86P$
P,58K>LVJ0>4G6S#F'G+8"^^O1C7 3RP]D,KD@[75+XR4H:H5(9_YC2RA9;9!E :&
PP0GCE[ES:,"<O&>ZI6ONA$TX;J4VQ;2=GM)ST7#B$8H49<;^MWJ6UUQ*N/P;FT&%
P6<4L]& =+!=V6VWG-K5%:T&#IM4I]!#YR>N@@'*F8T>.VJ\_;N"8#C;K;%RVLQOT
P0^C5S#R[>R:HG"<WC(WQI=]3.I8)Y\CI5*SE&?(4"S$53LS"FVY)]"0(G#C FHI.
PI>"P^-9W,_"M0PT!^YOE(<R_A$Z[)PSX\[N4!PI=T;?\SJ59;&&]MS4AYD;U*P)4
PWRIQ-DIH6;A^"9*,1HDU2$WO;L]%U' ?(7L^\!K"/KF&/? Y*=VA,2CI12EZ7MH&
P EP,G#_T*22SX%I;:6AM/.YRDBCNK9I="I)>=.K),=3/%HS# @"I"I8M"]U1!,(4
P3U/@S0^WL\==(]=1"-/(1-MLSBEF) [49,@0]#:T<;]25-2L]9G(!\#-5(N,?G C
P7^1N5IY8$TG4S/'E@W28!)I\K;;HF.@]HS)J5A%X)U-\=MG3Z8513+H=2(ZO4A/,
P_.!L,P@V$C!SUUR5Y75L4GCONY,QW@(P3C:=1>38/Y4L7PU1,INM@>UAX:RC2N[K
PE3;(P#-AS2TAR@_23'R1PFZAZ'TK?-["_.V\8P<,5[##L6CYTKO"6)=H1Y4GN'+K
P!V T+U!&):L:,\AD=44_8Z3[='[) O6R-$MJL\'!G=5J:2H +ZNX&3A,)4FBXVT6
P+ BW<]WM86^DM!B8X];.T74 W_/TZ0/14M=@KL@;Z$0/)ELI?T0RIW8(V.62L>F^
PY-5\=*."'X[(+J^N2<]<]&X?")W!W#@T@10 N0*0V?0J+E&O1-VG H<\B9\B&VWW
PWV\:(PA,$ZH,P.97^5+VHVB^OK/*+B0FB'*["_B'VF,;987X^!\PUE[J@7#T([[.
PF2H+53H.ZT[T)9+E1UA5@(@G W93C^/9<HUH0S)?<8R-&(1M+I.0%+2"#!28(?2A
PUOQ(OB'*$RX#=FW_L23^UM3??F\-A40-X+K6N#H*F^S#!P!\'PP'EEZ3+>$]C[J>
PA:'SRSQ<TB(;KU@ZQG42 N8O9#7)6/^P2S!"D,[/G/-23/$M?Y*?BIE547X -E8O
PUO6=2@GAT]I%%UB_0O.=&_0_S0<J%-QRPEI>5(0EG08^C?CYYC+9$".B1:DS9-.Z
P4E4?S0J$=%[V<WK_:",^8E8[3(\7GTJL!S4<JUDV+>D%(5#^<.G;8"E]VR3-$X:@
PSN[&X0%;6L!0/F1'BIFV/[^]GWC!FSC&U7C$?S849@]'R'3.TAU_'VMB8>V'TQL?
`endprotected128

////////////////////////////////////////////////////////////////////////////////////////////////////////////


`protected128
PDU7H_H3X>>IRR,/N?KT7T<0-(GPPGNX7S)K2O6232&=Z/G(,-RG>ZRZJA ?<O-9I
P'(PYU"C>U0.Q;%B>WC6/4B[* @"8B_/X9XNFS>NGG5BSN)N "4RV*E$B!MJ))0<E
PQ_6XEJU3)P0V?DK& :%\'U7W9+O;NU!R@D2.GDA]^;XF.-I/T=WI\D?JAEO9LD06
PWZR'@UFUV+.@ 1'P<2$$@%2Q>14-5[6&D^-:X7.-:M\/D!F8?Q'0$_,YJ 5(9[[;
P$WM^D!\Y1W3G7<VT?H-9@KN6L=]8UH9,XX<E/@!WS+[Q3D?QC)L8V2-)7W;A(:7_
PRKIXFA#%)K11/(QS.N,G&PT*'?3<H Y)$/Z)[_VTSSSJ%@8H*00K.B'=&$\-VE @
P;9>;-AT""L7LV_-:IE0C[^LEKK*1/01Q[BBFHZ.OEML3)S9U6.BN$TH%>M7=(;RW
PJ/UG4J,Q6JR<2PDX':I![/)KDP'S#':6YH2(0S+BM^QER>L?@N?95@"Y&T JE\N=
P0J*'O37WI@!,N=#9)54-GI!%*FD-,H6(#W_W JI^C("UEGD.4 Q(MN+%]@L#@ EL
PHFQZ;GLK.J0'N=M7@<*]3W]//DU$.D[]>?*>V.[H_7HT]>UGB"W5?-?O%QF6CCE.
PT(@S)8[,\'4O$C09C">0ZH!LI=W>,5L7#!U;VRVL'EXWW2]73%11W7.<%64;L",3
P68JEX=!/R,,0'I.MJC*]Y&*8&E^Q*!$,2Z#_&+59,KI"1!.;-M<SR$D#F9W5F<_<
P]56^/)OZ]5I.AV:B +YODW959YV.0MQNK(IOYJ9:]>M.--HM:]=.8FI@0DM!@M^>
PW=F?"X9*LWA[YELAFR^*TL.[8>(NN=?%;!K/-9#YU8;S:IOO'=UP#2C#K [4D06-
PYG,\!Q]V/%%L>BQ^CG/F5:QW!AT5 D2;(!*%C)'+PCU_*"T<'3<?,3?(EYH7)?5D
P(2D#OG=&C&(B(?/MY*=95 E?MCG@\//Z'XB&RWG2"YBL1ABIU:;G)2*X[;Z2NQ(&
PYI-^[I.\G7!J2J"A87O6G(2MCB9,)^@)%<F@(*O;MY">YFHY=&%H4[LJ%Q0N . 4
PK*;CGK$.'7'1:>Y!H(R@:[X/<Z@WO 1P2.0K&L04Q(H\K^ $@IK!QK7_^I]QFF 1
PQ(N[5>:@;03^=EL-OAARF[E*00G!>)W7(\!.!A'EGX$>BF0-"VTXQ&&TC(5E\@+ 
P84R/:D6&M1Q<3V3 #0HV@.>0X"4\P'O+L5J4E%=X%.%VICG,[1)6^H&1'=G&1Q!7
PQCIC<&8#Z, @8HP<2!Z?B:"'NS[9.6.1JRAGFG/3RI")+3\EPBY&]?OL^$OVA"';
P8/1\ P]^[(]PK7P03#?ER2J"TO]NW9=;+-*EL-NY"?7CA(=D@HT5?A: B;PGKC#^
P>X]9'(?""D4@;.6NL3TG#+$%4[@UTS73\!XD@W7#P\W1POULZZT7H4+\%=NTD0 ^
P1UM1<<Z(""I'I3:T'G?M[<"QC;@29%@:]R @N &_$'JMRVUM"KS?,#TT^=X$1E(X
P)MOEL3Q*6G3^+(OKK]4P8Y@SZO(7;)6F-FV,'>-*B%8 71AM",Y ].;="FKPET5D
PLKO._7)8M.46'S;*FIK3$!$5]-] @N.3@4-]@[8V! 4M%!%=:6S*&>K(2H0T]W$;
P8=^Q>>\QJ5&^X[NX@ E6%/T>)2Q\=FZCMU!VXGL"4. 54>I/,>8S0QIM(7V6'*G7
P)B+<JEW@8H 9XDKP8/,>=:M3R<ZWU;X>U=#>6>3RS+A>;9<.QKXBOK&WV912K$F.
PJX 3*P' V"J;,-P=$G[1\XTGT7//F?91@ K72=>*^DU!X%ZI> &F$ VT,@!FD?)*
P.QBV[_B=,T<@QTQ0V@<1^C*F86=Z\&%R\X9:(,##-'Y#7[6S>%*4YT'XYC #WOS_
PG79 <V!0K"X -LN2(U$DK<F")[8&I)1V>YM6YSX6&#EO15"D#&N'1&_@&S#SS+\^
PFM)Q6GH?7_<$^1/9#98\=L6/@PC(V?%][['<IENF<*N]P/9=*G>N$6U>IZ:^F:"I
P2=:IFC ?-ID_'A*?HOLCH2P=(PFH,W'9Y$[\GD_(D\Z H76IC252:* >A8I$-X\2
PRE3=B_#>8FVT[Y1,VM+:LLCXA/K7/O'AM<LI@6&<JU6ZB40<Q=S+M0A&W_]Q(NQ4
P"#1TA!$N]:.2=8I_NEEXD-*%E%G\0/-HC!",D.C1.@!)<P[!_8G6^#R4]].V3+AO
PY4EHO!,S=OJT%@^IYQ4GE(=0)X:I-=X9Z:J[+HH\<3Y>_-#D!=>H<X.-B#L<X>=+
P2G_O?]+7)[ASKST5IL9Y)+EG1KNU;\JXZ1<?;531PF%$]UO[3;W%P)2/IV4JDJZ@
PQ,E8O]E>F<78&@K3BY^XX#..0>0BNZ=Z_[&J6FQM;)](QR%V"R,@?8@P."B]U*A0
P4TE#6\][Y:X SA//U7B=JH^$]55MJQ'^M,6K6.-$T33 E2 S>6!%GPBH;:A]@7-N
P%.YB[2K E!^QP)2AK* !V]UT4;ZU<\+R[)MHL,I2$8GX\3CD0;]:NXQ:5Y92==!$
PMO@U:IO2E0N.#(H\8BJ/MM@R"5\W08D0)UDDU=5R,59\-X;HN"YS8) E\L^=R0UP
PX0F4:4G][!%:(='N>#]&:^"0WS,*/**+CLU\R /!M6OGVL+.-"=X;;NM1#E6L\44
PB 8AS%1+4=H(,I1=*@9__]T7/\%,#//3";IMIR.UTJBX_@=5_A$.&.V [,=3DK0F
P=')2T0*6C<F]YRB3.;#([Z5LU?D9'UZU4<[&XBJI^_+L\\O<<YS<GIG(VRK5-Y$F
P?Y2CQR95?RAV/UJ.-K<#D<^KQ7=@.QI1#Z_.=!K1@K@FJ\NF!O_80D55K5[5U];+
P+R,<@1.'9LI#9X-MC[])UMN/,^'$33DKY'UJ/CDMQ29T+Z1*R@:U,E>CTW#:NS6I
PIR1Q3<Y:*#, %! I)O<X'K7I"&LY$7'?0^-XGY7MX&,3Z+49##O#UZMJ)3-Z\XMC
PX.OKU)%<H^9=T^GG:48P _9MBXO_A8ZBRT6\MK\)EWV$2.9'F>]0%/3>=Q^*3Z9G
P"C(&SLE:MR3$$N>WOH<^?XFD;(DT$6HVP:4 1&$4AS=E=PV-YU?E&R,![NB U7/@
PL31*3M_!NZP!8>TA^"$XN$3M=]Q\PR/8'=>+B$<^<6B@X.>QN,,VP!H.];2;1=SP
PYH\D<A_VXU6 H65LCVL7'$=*Z#_F"]X)HF#DRK;DS_H@Y7+I@L!%7GSN5%M(0W6M
P.$$'FO;\5;EW!(#X(EPVS%@8 ZB9=BK"C_S8)'Z=LV0*79-DS;\NS^H2"83Q\TQ#
P+F[GM4%)BC4:N.8%H^:Q#"CZ=-2\TYKQT&JH7K?ACA=!MD'',FY8:>N![_&;(RIF
PXHU^DML8H[D!&L[+D1-4.CV6>:%=@*33+W3:O&V$HQ;-$CYE+G\/XE@JGT-I'-L@
P'O"I&\T"AS"N<TXY!D.8]*=?%;NR#[+>C>ND9U-#Y5#,R"N![678(YN\*(>8<=UX
PR^0[H7WF3!PUYL JI%]XJ;A>R5&0L'_,"_TZ,\GN;7W&,J'O/I[]F#K&=^T\LTS9
P6C-'H:"FC%YOCEET1L7\78R#R0 S7=SC/UVM+-;=<>':0P;;-92JD<M?TA $_\<U
PF%.?YALJU\:O;;>RHE*?&?IE';B'T7KEY<\/-38N$AL$[UREM?WH4VJ7?)SZ/1R^
P#ZN_ZT5SGB7S="<E9,W9O(MK8B/T,8292Z&8VPSU1MX:J(08]>U3$>YI)\BV'=\M
P'2L/[U,N8:!!DBDU8Y)\R!DW.(,T8@6!9>S,Z$*K-1U83II(SW*D9H20<^S!GFUY
PQ^V16G%$GX/:8:CL36*-Q*K4DJ/D:T*74]Y3T@SLA@FP/'*:2!_H[%A,>C4BY[S.
P;QE!DA"H-N!R'9I<@M!<BDIHK:F[ $H"GE^46-&"BEA>8BY^OD_HO$V,U3'CUC<C
P:2GT2D[;\H35D*T@U&Y_&FYD;L39<F_'1*,PFE5:L@0X^+$*ORWS!Z,$Z!=RU.DL
P#NQ;,$C;7(#=K18RQ/&;#^B@(VB%>X2#[XB6T<5&B^Z",K#]U58BM\W-BW>;FJ*(
PTD73@<U7,(:Q;UWH[(V4D5PHSB=DZ3/C@#>775]Z8\KZW[+RFT=<WQ\E>A?/F4/-
P)$IA(O,L##^^#OEU7PS_J_G\Q$CO SNI?!' !NDYJC791_>1.D 'KL@QCUV45C7"
PG,6#XR2L$,: X)C+D%?<WPU*)#/WY1XE/Z^#9CPTF[E,S[]N>"T45MTH)+6WS^8(
PQ'[UD+TC2%#H0V2@'0J;\U"0:-VER@DK91,CA+:CBBKOD$,))+)#XRLB._+T>PN:
PQ'>8):JK0+:<@9-$>@E$.C#L\NK77P& 44/!&<!K1?W^U1K@RVB30$P,LO$3.$HU
P=[.%NI6]8!<W'/<0W\([PTYJECU XUP1_#M N#TC,#T]YZ,"=8"ECLI-%<6J@^$$
P]!63#(QP",JS(RTI28GDX, +;_?1;H=!O.)W2='4G%[^\J ^ 5]W+D&C:+^P%EJ:
PU/)9\]+&/H!,SI^>.03F3DR^-5W8OQFDT2B_=W![7+IH>L<7(?\2.51$/E$56X&3
P6VCJ .!(ZA8'* E^1H\V]/_8Z%H@;?-CPHQ#WJQ<[Y$NDHQ#IS(3PM7N50)FR@3]
P>-'W('+8"55M;K[[9N3Q:* +F\TE;@6\2T*WDB!TP^"$(J*ECK+$NE!5D\A$7TM5
PIYT*.L\UL2X(_'<;G[OV-L5/W9U>K>&%>CT2O89K0OZ!0>W4\9H P>&K)]TQ)B@Q
PLUU/GVK?KE ?<.JCKTE(-_[="GW=[+*9RII?BOEPRQ<TA;O19>O5A8[K6U=WS$_X
PK(9:5\^VB#K$'QRQ$."O,KR#$D%04#ZLZU'-U&]3<![2S/I'L$FO<"S2<(N5MGS9
P'V_G,O)6QTLNP#I.C@UTMYA B,W3HF2X=H^F<0Q28*Q\N\L,M*YCD.\,:K_&&WZS
PW^*Q#BD9W=AR/E[Z68][:EU^VN&*YCMPRE&M"M #,GB3E>KJR#7:&4G=R8.3D;WO
P'.3[="@*+PY:>J+>,?8_L'^VZ-=>Z'7YYL1KU? []6G!1(Y9#Q)EQCA!\"U&@GF(
PAADI#[*2=N)V&4<F#*4E F*Z8(K<(4NZPH1&G(LHF#+'6:6U]VGTGS6]C5&O*7%?
PXF/R/0W4/S^BB4SH8;T>NH*^HE^RW)?P;+"'/9MG#6^91S75'?NNI ^HU9K*6@,D
PG)0JHRB<2\T_.3(_&R74;'OK"NT.[SG=1Z@5G"DU_)Q.@Q<V:#63NEW?L]WS,\@Q
P<@&,A;91 7]:0RKY0NUT%QD0:6C! [$SCN[]Y?IJ7LR1P7#W #TY?-2*7AG\6,+Z
P9.Z\(<K*)-P4.Z$7I*.Y_2.MM<A"AUH^,]^;L#(NYY@M7.Z9$ZO8<WI?K[:)_+*K
PDS*KK''!8@K)^?&G<[(C8 ) 4+27F^',P(Y=>?9MJ[S)LWSM'%&P,5>P6<>H=%.T
PG9#\S3ZO44R21"Z%MM7)4>&B;&6W3U5/:%&<:H$<Q>2\HUP&;L3=%V) JE^%?_N2
P%]#7<CYE=9H8-@F$18\KBVMJ/N:'3&/.]: 9J<0CL$ &#KTGCU7Z3?*OZC1/?1I8
P&SDTJU831%"\3%S/Z8CD&,IU.B2@ZE/*<=_(!$%.^14FU1??8GN"0_-5"2[4%)V'
PW.%K;Y_2(V*.^WMMG_17<6/H._9[F"!/Z/\3@&*/;BE4&G<]Z=XNT')HX-E(T*/9
P!HSM.BK2G<F%:>FRDSM!/[GVXF\2G< @A1YSD$EYFY ,K,95G#I[G2#EVE<6H452
P,1 :E%J)J&C>UG5N*55>E%RF'UJ!H'RI/&"=M-QK&[JA6;YV!02K(8L[D=,#N.?&
P=>/SX_&UW EDM2;[U 7O;3)\5Z'_MJ/7^.%IR[P6M\G6125N71@QCCAU.XZ.)E*;
P?V2Z.W+3?J5ASW9HG"J0M3]6SNL-)ZH>=<;0PR)$96K) BW+:I\/1N2+6TNV*V>!
PJ@T0>!5M]3V <M>\UE[KXIBW@.<TR]D$Q B*<+*J$C@S(GE55PQ<!)@%A+7%G^K+
P3NH$(F( WWG,F%!+OSSAU0H*-W:D1/WKE2.<8&^-[(>4Q]-O-MPQNCKU3+0"V+T7
PZT$&9);;GY\J;HRMTU(&JGF[6<A>I>0I0.8REA5?U=,Y=;.:'@"Y;4OZZ_T6G,.5
P<NX!5^!Q4=4JPU!)>JO[3 E*2O66._++)T&?P_V0 8)_=X=*&, Z$5$"G^)Z.(<]
P=_3Z)NVOBQL//K-;N_8BK^7&9IFC7,X_ZRX1[)NHAH$<H(=9])LS?+'?"%4\SPZX
PMFTE%;*H!+=KU;U9R_"J+#N<%V=TPKL8U%O1)">'TSPG1G^4XL?OO)$9T\IFV!6W
PM\_4>/&4,4QE.9A($G#L@_KW*1+P X9[F"T\^PH. !.HR.7DPD6E2IJ]@IO3N6-X
P8X9I;"3W;0NW0'&$>>==0D&L6__-FF._:^SQ<ZT9L&AXO=.O3.:@"F7QZ,DZ\NN\
P,N<JE)U!<NSEJTI5TO^^3..7E0!">_FTG0;"(\-\J*<F8[$C;* E&HN?!44X  * 
P\J^/"/TH;[(2Q=\MN.>1%Z5/@QC"U@['U-\Q!-Y+&\1P2,UY(O#8UM5.A*;Z].Y2
P^0$>5!!KV(#?ED*IEH3R*^/;WETR$N&DG4I"NBX_>^/Y[\^WV"\U[*SPOI 5FDN&
P;+^G;\5-&/QW,+2NQF+UP?]]/.=(JM1E#5)K.F9/PWX7\KY>27KIH))_G8Q J5F3
PDG3,XP@JF\4,S#F5')"ZLAR '4<!KUFLCACX;:\/7Q:W946_FWLSPBF!#R(MT]=.
P5#G;!4KO-!65XTHAU M?+# \4N/,_2>5VB+>Z4T5U:1(XMD#.1/GV> X;&AMC87C
PN/^$KQVJYM&*[S!X@+T[/C,')AE,-!TIN6PY'$Y'OE ,-7-YD<TX-P6_WO3PM-TZ
PYLDD3V-I>#&?3XTVUV2UQ7DSIM*;3#UBJ<KRSVIZ6\[F$BYP493Y% !4OWPXV7^#
P+/X]G["  2V/Z Z^OR\#<=S?E)E@<J5$WYN[,^Q7IK^,PL!U1DPU'3;2%C0K&*F'
PJ*PI_T$<6B /0#I.<:^RI]LDB$Y;HEC2]*TJ2^]<MXU8BP[+&#V]GIUL4  &@\+I
P^GT2WCD3M.%8,T^B[3P:3*HV[;$;UGMR'/";.1AL!-0/=2DRH "D7^$)&#RU@SF=
P,%6KG-K2G[3M$/Z"/(79KP;@^+OI)QT^6.L^FH\#DWI4%VOE%;-UH$Q_+_;GKU./
P.;I* 'IA?UNN/!VRA2J?^'3VX$>C_(U]0*/G'6XXJIF2A:8N0$-C'D(F\1Z)J20M
P3M5>32<S3VI]-X*AQM;WC8"UE:R4D*RYI*&#7^"C,@D]3BSL6&?C:-YO",A46_=W
PZS)VM_'/1/8AJ)$9SZR1%!J6QT'4JH>=:5,?T5]=A6=#3.%ZB3Y.42^>[.A-&\+[
P2A])>P'0>?D1OKQ-,J&M1"#IT)+8U*H,ZDZJSDW7\'J%I;F/8%YNT7&D-DMR5)T&
P&8F5X1R00/AERB"]JP=KI8F0T,A$HCX:1<+_.EAI#%P[KA5C912MVP54] X_"##;
P/"WEAT-@W@>9/?)4L?0@4<Y+&/6D6Y+ZTP&,9Z8_[Z>#YIBF$YTO.ZG3CL'P\"./
PZRI@"Q[DBC?_DMJ8ZV($Y-^V8@\RO;,\;X"[96+<X!?11#R/.L(GVC5)%8Z6Z.]U
P4-T>HL?&+)VM/H*7M%?>^9/$?'>RE%'A[/C\13&SI"TL3>PS"KNO?4G86]SP8R R
P8)&'A@$V1-U9-$3(+7=)>/)")&AMJK+GK.&UOK_!B%XF+V>Z,.I %;]B2!?*:"KF
P-3L$CP2;7QWI$IWW OJR>&;47A^?B2GFVAKG8G[EF+^Q^8/X?/23?L%&A HZ? <W
PJBY&!LO[R)C'I"X<E'I'NF@K$M#E):_A/ J>_LZFASE)FJ/QGOK=Y&KP /B7[4.O
PHH+C<9)1F>;A"C$#Z22H%0?P@*$@$(O%YGOC40'$[@V]X;PB3@[=;.!*UY ?&3:F
P;!=&*#&$,?5!^-3EX\"7$<C17OVH7D0W5+,?Z%TK[D3<9I&AI0ZT[YH<O JT5A:G
P#9=6[LXR\@DC[-G?(-3)T-DRU/XY_JXZ,6@BTV)8Q-[=J+,@1UGF%8DG^11@,VTN
PHC@95F3$; /_.7 3R':(&-$"QH9\\1&[/V.(2J=,9_G5F:7N<[E=P!H B?+Q'F"Q
P,3L:T1+DIMLV'>(OB(HIY)$ZH1?_MIH:V[JB<D--(X8*!>WQTS>9/,9W5!&99Q="
P"[%)VX%2>JGHB Y?M;5Q/-Q+%V2RMT#53)Y[Q;VSR1 +A*^PGMT9E!?K )-O'II)
P&.;15<^9*6II0)L[OF*:0E^*M9C)4?QGX.%%]$#!@@3EJ@/*LUD"%?@]J7R! N'Q
P/UH4-<&.)BTXS 59J;D3039A!!/.&'^03_E5*/U7@M>T9<MIV5D4^H:\=3T4QDO>
P+ 92RZT,W%Q56VEKF<4\1%!>@F!JCT^XP@=B'80W7AG"<D8SG&%+PK#Q(4R7!1:8
PN6!6D'+MU4 ^;V@DC[U<0)MJ(UE%=T!-#R MGU=NGJP;0F.9%]0EI#1)2$[Z[P&L
P1T!$:H,8B]81A]<]CT1?HM:"&82TY-)$%>HR,H8F$J]U<C*@B>3/LQTLSN:+>% >
P UK,R82N0LUE1)YG 15-,A0]"WI%[K.8#]RS+7ZMM;BU[S^[X?L(F!)6'-F'8<>U
P,EA8QY&\,Y/&F47X%F "OD$4+>:F[KNM'!29!,94;\,W X:O[\B$2EM8YMJB_;7,
P6=(W4J]KEE9<7G'8:(ZEZXJH5)ID0?T::\:QF_K$9$# (#^G5EHE5T_W9$71CS\*
PX#/T8.@#=X-%IL4UQT^'1TL25"\:"Y,J1<3N)K<A="?C8*N1+GW5D0/O+9_@5Y<R
P[- [1]UDXJ"RG]D+U#DS/AP/6^XP]M:9$=SK]:QTU180/1.(FA:-2(6!Q3<-G#B0
PUO"L&IJJ..AOK:LFWZ.6.+$%).#//TKO6%6BF@\H>-@!$C<2EU:P_DU% 3XPOY.[
PX2&P'GFU0SH3U#?YC2]QF9T#+AE89AF4?<=3!>WB3MAMF#)M:.3AZ+F0W8=F7,8[
P%4^:@U4RM ":+W,(:R*S>)S$XX!SB(@[\E00_HDR4ZI9EE,\QTUNL.X7>>@'R?1W
PBWR:"0::RZE">S:/$6/0?V'VUQH'VCV%)!2^_0YA'#7U0K*PHAZ R:I,R:O?!43*
PA^6ZN(<QWHV]]EF,(*Z.0(<F8B8L<U/:#-EY&\\RZME. 1FXT73F"7R@<4E<31@Q
PWE<3DUG!N6^GSH^Q+)&7.UEM_%?2EE3JL[[S9PGU7'7"C)R@)\4:0OCFB?M#ZV-W
P$QJ5PLSD*>4T'=L"FC"QQ3INQ8&;C;2,R'FK1N6FUV;TV"WE=C&V#\,?0*S*,#Q'
P)_R[X)>0,KIW=!)0]#"UU%5*W(7^6#>^: (PI#L+:1,1+*U(F[2^J%IUO:X^<_6#
PGIT;D).KQ3R5YLL;L'TSUBLL#:2%BV 4X\P5?,(<X8B9=SY9,DCA]%L+^J0NTQMR
PZ#C TBW4L6#"D)>ME /I0^'#"9Y:^4'@@ HFHX3/NFOW8$GKB]0$L:4AMA6TG%<F
P^^CT1T@^,G:GA<9.#932EBF.#X8V9O#W#BIYIJ5<A1:(AD>KO]Y$)MQ&S-YJ,C2K
P@.?BQ>&]4OPDH(;&S$>-75:D )_)U]6?>F ZWUR8"Y%PV8BI'A_PX* HOGNLK[X*
PK?A"^EF>Y>KI%*O\MPY=(^!&(/T)1VIDBA)_B&K."4KZ:BX']$-+=U)/_IU'1<#Q
P#_;]\O<1-QL+U-#*N().N(D)/,=09%;:KF K0>K"\K9](3MZQT%+CJ\RH,W<G!#.
PUPOXGN9&ID7*!>,EUCA*/'_T/Z]0,T;Q.POG#M5P]I3NZ+H5.%I-L.UPCBO&%,RK
PC@1R(NQ&'G4%+ 8A)3%J*T;16,NO6;8$$[3XZ)?BX^;Y[JBE"_46-M.7+>*I<Q,2
P\8^5PT%%-C W>>+.94-D0[3SW;OM]T;!*=OMQ<:PG?<M,0%,]O0S?\1)IR>MWB"/
P)$NYDM>W8?!!@&MGURS4_XJU0!9=:J-5-\)V6&]=2$P]"L>+.LC7G>&_J-YN>3W<
PTSR5,V"%WAU+J4'SF_LTAM%3'_TQ9.I6,Q?.'%/ZLQHQ#PZ3KFAMLM=*][T>6"LG
P'+9@>6RFWF2%$#<>1F'4.V<J ;"(HQE['Y.BKRZZOI-M ;]UHU%+9?+ ORHD_:V&
P94:.#P1I(A+T0K:8BX7=1Z::LT-R%GO1E>HCZ #XO]&3C3U9G4:N(LMGK-;R2702
PH7;A*N&7B4D[L(B9MJ#$1VD?8X6OFJ'$PT, =I:F9="F,(I@>BOVL?QXF*K:\Y*7
PSUHESSB?,Y'Q]$W1'L2<9<I/]K-5X\;)DX17'L9N@.]BQD[JRZ4&:X6-1AB4IQ1K
P5RSWX '9G#N[!H+%+XN7&S^+-G'NC<XZ-XC 9.M7(><#8_5=WOE_./*;EUFOM==4
PI&>9IQYE]*5)Q]C%?8NZQ1$MP<@I3HR0XZR"W(9?O.^+XP+9N"FN\"E_.8V$0HV4
PY.$]/O"NRD4P\*A( 4!,"H3,X[45+0SQV7 OTJ6WI\5P_1)?)^6N52$L3^RLI5$E
PHSK)G@R>V'.R(-V.M'D6\5&?7N6*IHX!JFZ0DJ\^\Y_KN9#$'S&CN/]U[^>RWE3X
PQTY:=.\CKV>8CS<1)UIE0%]*I92[7+%"Y:6[VE#)EM_0'Z?E?=L($>TW\<@B&H2;
P0 D[)[Q/C8'W )A$YL&QO[PP&_+F]V,[6BZ6*R>.7[?%(_#3GI:9EJTR_T9Q/PE6
PPM-9679M\*8$03#_.#:N/PNX^+LVDW@M<!QC&;%8YBL,:NQR,>WC6_P*B+$3 REC
PTV1PR ^CZ[.HMH+QBKUD42AZ5?>X7J$WN!26$GIDTMP&+/4_R=._/7XN</L##MH-
P:>FJ#+.1]Y^]!G;-VHB&_=FWT"E5R1]RK7]WWHZ15'"!X@>Q*GH +<(I/03^6N]O
PO'4WR"03U1/.<Q3LM\LT]66Y[$+*M B,<=":]K276\ 538SF':TC*>$.S"-C6>JH
PBRM*'\KB',0KUI3*9959G^WKM@0YU:EAD]$'"RD5I[F3$;U3E FM#*4]WEZ_S?:P
P'X(%:F]>Z^MW!4!%RIOQ9)',&Q1:D//V+NKL-W_+:>5FL5:?:#N$J^6.@Y)W$=:R
PA+]1^'55T;\'MI2-)E(;GL5Z! K< 3)_.1(!MAV&!#\KE;HZ2^,!*16X;/R)F1FN
PCN,@<_=0^ ?BK)^8C8I." 1MSS 8II@\4QD%U5*!@BVD!SJ(4S;:^Y'#$!+%6?$X
PPG,5S^W<K Z.S[<NB0 5TC#'PN>S%L++-]&XU6F>+NU:;V?GN2E7_R<N#T+*$T5W
PV%*I)2"B8Q,D_4<D3VE^#,RYWN+11-2AY]WWF_[VE:4.$BU8ZZV+^.AA@P'\:?=R
P-RPU ,*&)\:N*@6R3)I3=]^[5N$ QO51K[@0SJ8V]6<17QO?[(T\R,C+]N@=,V(,
P0>4G\"BOV"]8XO!(ZA3* G-0SFV165(.@Q^<SP0C-1>]J%"*+<SR]2Q &A AL&]P
P;& [IM[ 3N VO 80-$'?-%V5#V=^[V)*3C/&O"S-,-<)SW327VTG0( G2]#1.A-E
P06:7=MHSAFM7"^@&SQ01B&7D:L4/I_TI*JKV(PRHK6M;X+2:,*Q*<$"OF#XU)OH2
P[LT=#VOT/@AR/Z[1<.B;1A-R,5/$4.HBQ,])-UK=Q*,1X3M3C??Z4Q\3N0'++?\7
PWT)\".&%L.RWCDJRK-VGFIP[W6X7J)4/!L"L&4+&M(FT3-3:W;!?0T]8<?\]7Q\-
PQE0S4-:\<DBHUZ6]C9?7T5$4W>G5"LG-]X%N"G'#U]GW7"_@FRP%#$?# G"78-D$
P@%_L:M!_N2;ER<])>$<5+=HNQ/*F[NMQC;<;CF!3M\<SO0VLW+&X ;D9F866SJ$L
PRARZ%.4&)C ?/3/./6=H8BK5#H+UR?#0YX)^?M3%G0*')) Y[\!,!>C>:QK:\4^8
P-+[OF-?#(<LZS1&O!NO$LQC#Y?HX4O_61-RKY)<9#654BIG8FVNY1-WD9CV,&JW]
PZ3VZ68T%>-VK*(=BD0M]0W)^3:U2$@B2'P]I/ENG*Y,B*U609QZWE(S+,;1%<3WI
P]T/Z:,Y,J$T*2Y'+<F@E_"AS/?8)4E%!(O1K'OF";E*@<,\H8/-[!'>/&4/MZXEQ
PK8GA*;I>S8C=CE.*K:"N!0,'S,*V7_DTE,1LN&5>2N!%=P^PU\&35@Y/?OY8/ 9S
PR_?DF'13$/>\Q%%T3HNQ/<#VG1R?74D25:BK6Y>!?G3R<88Q '@.4%&9E/A#?Q+H
PIEDGP3S<[H$;!A;#\K_K-"/\DEQV[:#0N0\W86)WD7A.HI^BK*&=-<59HS^26"7D
PO*SMPZY9Q?F;*>G?1.;"O5YS.SW?MU-=O80:!1S? J-0G3WKS3W_!3>$V3X&H.!N
P,"G>GHZX)"I#7\)T/E!HH>)2;+M;$OK[O;7'Z9.*4%$?<.2&,BI;$Z6*;@WN:<GF
PEVVR*A2> U>$U2-$X4-6FE(P2D.K>G=Q;85E;4R'ED+E/U_[2$V7$'<QBE04Q#M&
P3<]AJ*S8B;YHI+63,Y0OGW!-71T9/WSH8FV[XF[7$B$5FVF!)X<#RXT##=<55RR_
P1Z7_T2]XJB;;G16R"GQ:.=OEHBE[24G2A:P'$/*8W.+?5H-$M#75@E2*P/^.&/2R
P;),#,T*)($.[;C$/2ZT4F5B"(X*;:U+Y!Y/CK20#LT\GNT]!)*Q)S$SX;YO5A!AJ
PWD[N71_Q$4D265SAHYATU/(*B^/H$.\5-8,=;I^*)S5O#G97_XRZCYAQ I2FMQ6R
P*8QP%YE8"E48]T]-[81V9 1.@4;)WCP8UTIKC<=J4<NF%R19!>D#H4\+]SFJ)3H$
P5B?9A4=@K-#!EQH6UQ77O])L YL(]?42'0G_A9DC,2+4_OB5%=7@6+<6R6)[<;F$
PR,']%2E^34 =4X/<)7Z=R.+/+4A3!JK<XN';HJX[8/+;1^5;N:YR,/YP/?0A<6J1
PURC:MK6AKP^"L];1.VVC;PXQ\H-,04#N-$U57.VGV@IG4<K<"=F0DPX,NP5YFS@%
P@5:<O)6((!7+<KF*UPF3Z;FPQ ^1BVO!S.FSMI3SZ'J .\6U#$;S53:6?NZV%78.
P ;Z$[*4WC#M#+)TPKII;>R*U"8C_5ZJG=\]OT5:-OZRIB, BPE9"Z:J='ZW><0; 
P)YBY]S"Z"K:+WQS- ,>/JN6^ \ZP11E5L'$ABU*2T#S^O/S69X58L8Z<COPH>^$#
PWJ?X,#:MJ /F4,N_3+C31[YL[159CAET4/D[DD4"  Q->%E34#UL1>T'%NH Q.L 
P3@3J::/+U]V*L\/B%ZA_@URS4^] ^8<I'S<G9^*0CV%#VA\/Q]-8W*1@% RQXL?+
PJBHP$'\VVX8 XG@&>3/8Y?P:M=@-NV5Z33]QC%(S^#C*\PI\&8KQ]S90TK3YE<SZ
P!J7UU2-%D0ZCJ=RR\ZY![DN.3WO-B?7;)EOOJ^4;83B=AJZ'02M):ST+5$@S\!YX
P=NW-K<NJD<5?HV_&ZFN$?::SS1HZ*EV,1* >KOA8>KAMA?NJ\ #Y6Q"]:G,?+U+>
PK"?M$>Y8_TF+T5.-AT$ONF=('D'F?+T"]GR:Z5-K^F9-MHTWP,?E!IUGA8K;:)R6
P%FZZ50%"(=> :=U!E5CRF"I:&:@9$ IO1'&;.<*QZVO;Q>V!F/,G&2TQ:D]8B^N&
P4B2907M-].-<R^+_P^SU>]!\P9PG"G0BGY)M9?L)=W >0ESL)1PVO%!T@=($;:#2
P%7IS)2HG<5H-VRQ_]<D8\.S&P& :%D'V[L<8W0,G;0$GSH$6H,VNUG_4MVJX0$I'
PDT62O?]-\LX4Y:C?K,N,\M:\MV]%_CI'20BNKVG_I$K+P#/R["R.X%=DPF :_U5;
P853'7E/H#SE.,B41X*^+-O['NP[_@!SO?L>[R67OB_EI0P-L04H631R2&:;^%91J
POZJ?(8J12D>T9XI0(_Y+#GJO_V8M$O++>HX9Q.C(+6J$EX5(=Z.,1G(;$AGI.B\]
PBGKEW?*U?EP8Y5I!U0U'K[K$?><QK::7GE<H0\+7< #)FRUOS:0F<U. U[)GW$83
P5TY'H7F+EM9G]$J3E5I7OZB7;3;%Q_! K1WF_(4S^F[?X3><*0-\/K"O%B=+8-!:
P>;;DR3)M#_>1=219,/EM9!VO?R.U;?.V?1Q^Q_*)@5B!E7^1 -;I>_X.XAJ:AI!;
PB%?*"2G#J6\71TD$P6TI$OX14GU K[PX;IB%?#)#4'SM0?KI44Z1I^W]9U+QL??I
PE[1L=$R53/R*R*0O>P:I5SVF "D;K,*2%/=D -B5Q7;V:43Q?1\8=*C"N+T@U(5E
PLR5+$/:G)5P%?R+WLM8#MC=R^8[-@/,@*Q,C,\\),<Y?Q,M,&[89<&;,!EE#8 KJ
P&1\9[!AMLGI-/O$I;,()J1Y->UU4^)&[>5 '_14@EG<G?EB;K;7%#R39@52K=-HY
P]Y!,W-C.@P\#O@>C.FR4,>1<B+@; !@=PU4;AF5 QT#_:W?.[=8J7231WX#\Z/&"
PP94S$OO',-+^C*A\(#NSX"[;QN&4NU,,YN:WI$*RN*&:HD[F:/P/[R_:33)1.9AI
PP@6,\EI^"$JO7G27L%-)YZ ^/(YR7W9Y/,#L\ >:CE'>J&$HBOS$^D4WO]ON%%A8
P>.NB\0^,=^*\AY<UD[)Q>?_516[!=3].3DW/HK;U5=3F\3.WI"Y\,K5>]I+9HWLO
PE.N+D>7U!][D%/XRCT(T;_';&9(HK>(<#]^:(>/6>U:\W2P#,^H8)08F[4\EW5*L
P>#5ER3L\/NU72P?MF@KG[;8S8V0%]H-8^W,<+'4,[*O:!C5243N4Q8Y8ZR9QS-5C
PS>HHT"U^-@[BGJ, 9OZC$P;[UTOQ-J @D+9[SG91B WTO].O-L%KK]6M.$/6A:HP
P\_8=\D?.,'VH/OI9+>XV0G^J<B_XBV8IB0RPW60A^XKY@_*5QK_>."K0L-<Z/""@
P8ZQ%8G2:SXG4@(QE%;F7[:] SR1?J'"K?HZBIM"FAH3&^(FA9#N/;Z0>_8P[WD#L
P?1!!Z?C1E?K&5-*RQ>8V--,+)VS.1474/_>PB[VJY*.RY+F4%/;LIG>!A-QU0]TM
P<9&L!2J/>E-"I+C6E9;,NS*_BJ+'+!Y&W3C_2X4)6D?(0NSZUWP;>PZ;CS1(&Y,)
PFQT]@ YWC@%]A RIX#4H?"ND-U.QD=6?]IBB^R*+P$ASE"H&TI,; GO[J3-6R/^?
PO#=5L()ROW0[!6E[V19GK#'52F1TF@G0=,]4;OHI :#_1>I-KX+*XUO0DO'$4T$9
PKVA<>U5O0IKE*0(UT_&3+(IVG;ZP@+;]0/@W&\9"X]CR%L[IC.AW:2@+,4%?:Y/V
P*50Q)WUL^FB(,?X_[A5(C1;@P().1)<>F&X=])8^1$O''C5N#U8//1\2YHDE,+/8
PS5[JT>:IB@;-EI$7<V2W=;ARN++3'F4@*O]EF6GQ<Q[PH3(H. !TI'YSPNSVJ)UC
P1T"IC<,P_M[A+6)_0GQ@'BB P9)Z_>\ZL%OG/<+F[T0$N+,R[HH.DBU/&OP5FEHV
PBQFF,YHE'8QM%SU_=,>9"I2]5N'I6Y NJ13?\?WX 1RYR69R(LCIBN7!9G>9_].2
PQ=[*N.!ZWTTK$G69YFH6UD=1>TM7!A8[A.T>R/J]3,VJ4[LDPC'Z;CO^HHX?E-FG
PS;L5!!?E9 ,)SVM];.?4,C^=@Q%/XN&ZL00;4/_Y,J(3?:LN?$'M)I$/#W%%7)S\
P8B(3KVWY!@6R'=T9\^R E$J&X&25!7!O=-57_#J4X%[GJ1D16>\_6#/:6S19HC4I
PY^M* -4=W8AIE; <L+R\YN%8$P;=]B+]RUD_"Z$=MTQMJ4L"\-\E\,;CD)^,L#Q^
P#9:LE*PUHQ,V?D%Q0Y)?\5J=#%E?WT1(D /)EC:X;*4AN+7/$4D#U^S*OU [0JZS
PZC5G1IDM?(/;A#MP\$F*@$,QL/D<]3^?B6FR[C-YVO9^"F)R85,2>2G6EPEE^)4C
PH@"WJC0$[,I"%!99JPZ4-=[NV#>+X$)SA8@-B$D5,M06F<W6UOPU YP',9,B#[(Y
P9VCKJO!PE5TC^VP+6)W)+\0#Q2XSS*JK(0'(+/X#^+7DF7-5E/1XC$B#W5M*V^/5
PV,\@OSMP<U"""\6?2&"KU6#JX)A26LB9^X^X0G&]F<KNP*;YF"GX[RI'H&*!8@A@
P0/5-(P#6G>A[G-7ME(/TW*:Y])X%%6)K;P"2/;LZ*1[ZH/STD-SZ4N\YL3V<OZ?(
PFXT ([7/:50(U*W_J:YO_.])<%R4?*FW'^901KRPS[+93<R42+B!:![XW6,:JQVA
PZ_S_KT 4GV8")K"#51[I@1](NW/2H4WE-82F O/AM67IW*<L_W #4;/?0R_(#I0[
PC:9"#$7,1I%XI%@SF3@NP89;>P5L7".X6';VZZ$'HX<ZS"81.HL*)1*XP2$4P5I(
P1!A=;LF1>--+XAK\73%[T\N76%<#BJG8R,S@6% E(LJ^-V%-64!E;2>M*US@SN9Z
P67AQ'3 ^-R/%"6.0XI 44AXL/*[ QNYZ.SE@;> V$JM A+UV4Z)N?D;#HS70X)ZO
P[?O^4X',66B!)LQ2GD;$TTO9VG28_:(3$;HR0+=W,33W5E5-E@-O(?@<VK.^85H+
P+UR4 =C#7NF0U)?%[)DX6TM!ZDDP?EEU_/5*4FGR^TPB!H\)<E1;RL;(V?%Q2 M!
P4>>LR/HB<^ F?:O98X2)DF\B+3?A.4XU\7W)&Y9UF";(]OQ%8(?1]WE@38!1#1*U
PL7/\XANL563!KPY(GU9FDUJ.["XJO35 U/A.*(03M &1/'2G*88>H9[<QD)B,B\3
P8PFSVYV]=)86U@MTK!X.KJDO, -(15 ;928[&S(P-/3;*QYXI25:F=,ZS7+U@+X$
PM[:7\(R'XX%CQ%AR=6S;5OKK-7,D!Y*?2I2]'YABRE6_=UB7QD +$OZ87(^-L7$[
P/IU\'9E1@O<.U;A(V]W'F?IL<E-@5./(#B[W((DB%VC_=45JL:[&BQ>RP]C95J*B
PX2X,#^^N>=(B=0^NR;$MC;(FH&1)DOO34:: / A433/7.BVQOD>22!;_'X>I!\H<
P99_Z*;@SK@I57&PYD!NI68%+.>I?M-J'T,G5J!_L3[S@GLR8&@C7?Z&LBB6G=9]M
PVQL&-G%#$YW%?!H2AG%7)3SRF5,6"NG*."1BC"8-YD>/L[+D0$:HHE1BH^-L?*CS
P+C3%+32I0(S8;T]DJDDH(.DSKH@F?[<#U(3U+D[^0K=9Q[#B(XX:1W>9=?!LU1VZ
P<9MS5(1LA-6%->JI25:FY4*ZG3O@H1!)3RAG>'$TR(S KNNG!IK#PP1]BDQVRPIS
P](+E5T+K]U7#K#Y98Y"^6Y_VY6&/CC/(-R/"'S70*YEYSV#_80L7RE;I E/F2<>W
P W8-$K4=EIC(_JAOR3D8.H-NGN2Y?>&VI2 1P=5,.ERTW[Q#73XPOWBMO-9V.88J
P;+'95-U/4:PI\8Y!$$K%ZHXJQ])Z:^?XH^>-Q8-KEGGF"*NV'"7<-I6C_](4C<T*
P^)!@739>2I<'.QIF3S@XX"1KA%9"BRZSW]0!D2B@8_: '1^3.&@ @4,<&;F*2ZE?
P[@W18ET1FYVAT/J%VKJ)U@C??2@=KIANG&*T^!N?E?*J_()K.?K:^Q1,M.3Z3?B"
P!6_$3HN<M\*,(X)80MDZ-!K,),0<=EL%99C?)+[?^$767U\YO($'(S.ORMP0TZ,[
P'M!S6*6IJ/A) >US+?+G/++].YCP_$>V]5V/[_-@Y07K?#:L(1D)FS%'L6$%(27^
P6XN(!&#Z>/'G/49G108.P\B\5C%VZ;]FO^?!G]B1G_X'<X%VD<SO26(-NEA'8K1_
P!38M@:$.7!K1_/H9G2("/P)Q(8F%Y5>\YE?7(#PA>LAHW58(=CZ_(-$@3IA;>H4S
PD,!]+Z9K19LJ"JNA0>&OK&?]QT3G>#YK;PF1]<34)P?*RY2MB:Q'\/JY$=3%NOA?
P^D_9#;R;/3OW"U4#5A?B^(D8!!8BZ I\./%63D(KI2;MC[I.+:DIDP6Z/::O[\6N
PU0/G)#P0N"([JVC=]C&<!E(O8:2XPIE"&UW7A$SZU?8.?PKU>*'X.Q&3,>!*L6FU
PGDO%R;O YBL;!. [/X OD-016\@)M:T7:G=>N<W(LPJXG^%Q<4H:T,\;^%Z=TC9J
PZNJE4HN+GB%D71T")?^Z<46D!U=HTCSL+"+G)9>JRCT>W8N$'UD$$FY4-\-%BY?A
PZ^L 'W9?9([PQT== 9'1$??]0S&%8?=-G7@/1*"?V'_/\E]Z>#$%7O\::QH@$EG9
P4#D12E>HD\CN$2_M!0:GAL[,T\D@V(B?LTZ4U1=?55:>/2;KB"1]6FKZ[II;/CR/
P^];D*/OQM!=N+*GDK=?VC/[35XK3L#YS*>3<(+$N5O;\@)$TV:5[X-/O6^:L$$LK
P$P'\-(61I65WKDSL8+S,*.+HLQG[J<GT'XT*$P!7RL74SR=UA0C;!%MP8A/HP6HS
P^;33OCMKK'JEKOZ#BL^0,E$3U"J'RA6*CX<H=Z_HNA$1,6WJ*3S%B:2(NDLA0.VG
PIM<6;*0_,0QJN_-9H62_APHI&=B"PF351T]-%;RX;JA&K<6O4FS:<J:0Q+BMZ,Y?
P:%E?A+K]EAQ>F!$KBLMCN 8P)-EW.%RPJ[VSYV6;3W)VXCP[]^9-P32JN@H <K*^
P4/B'U5W]J!?;8YJ$=D0IS"Q2TPJE;_&F>/E?7CVT@&35 @40Q*UQD;8S'0^*#K!#
P+=;WW*2*TP7U. SW_ZROOXL6'"&:!=NWA#ZD0&=(-\B\ _UYM5HB5F]@<Q+U[F=L
PV\S&6#(EN;G_M'0RI1#YWPB#+"1X*^^7(\I;6\PK%JWM< E+U+$H)W3^$#</TZW2
PTXF/50R493G@KM_R=-Z/U^BV#BD=Z:@M;,6$D_'(P5>)%,<PN]95Y'Z!F8/'WE;Q
P#>NV@1J=A UB6Y[=7=\?CF4DY8XW)?,%W3.ZK6?NN1^)FO+G!._:)?<5.8EZNIM?
P77.2BK+#H0PK#C,NHBVKV$$#*;5"R_*\]]P&9/)\J' I::/U_D/+"V5EI$F-;,WD
PS5*L6Z]SJ@6A/ D+)U3T,*4.*;S'(KNP@#,6[:KF)&3R"ZA*>YATL>$M<@VFY/&9
PY;[<R+ ^ZX..72R65X;O&B"<UF:(R=UR#MS)S<-N(9N182ST_6DL+_1!'#,V=Q15
PEJ?Q66*&MUL'GC5=(8E'V6J6A-_, ,:20GR_8ZO6G@T7JAM>M$)IRZN+U><,R9@)
P&WF0TC-@]>Z"-IE/5=/GBP]JU>M1,*ID:D%VU:6FHUN"@QI0]S:AO/N'12C5SP)L
PD_">_K3^W45H0?KS3/<Y,F?+*H]]^E&ME'CV[O#:)IRB7'O)/,M$@!$R6*A3;XEP
P\\('[0]F"JJ0G^/7L"% @LBB@6.9+8*,LV8ZH,5]-]V^?\"( ',:D447'?)H>:OK
PE:*2+(M 3IN,FF?R(RFE&X#HF#><#-?A4!$ &FM9WA+D!FTW%Q.8J5O1&YD'.&AO
P;TH[ZJ+F5)9'EY]5K1-D'@>\@QGP7=:UKKB\^+W_)/RL#._<XS B^A:8# >"#B&C
PD9;G<6 +N/&P7L1Y)-?QSH3*7Y*YO"0>D.4$G12CDU_PP.WT&&K%0Q";OD E-][<
POI]!;QE%!-J/:^;/-8RAYXS'<GL785^/W7<IY*#7I:*]M"!D&W+8-C>\DID9V.(@
P>"_96-K7=J0Z, $8/ZBM:.$6*KM3UPZ\W2(8):.=9WJI C\J,5:WGRP2ZLE<9@7J
P E0SNTYK\U"!, ;1Y@WB2PM>_7XE4I=';Q)WYZBTP%$#OEM/ND^W0JB'VS'S[N(6
P#ED%*M3[IW,1E+7^F> S.!:KW7@QLQ,G@DLN"BM6,W-EBR1=3"-/-*RJH]]]];W<
P* [LV&.$#<O.20F9"VA3,!&Q6R9+^/,<L%*!"+I,F:]0]ZEKTW"<T34WD.(%RA&N
PP6=4G__0'9D/\^G/ZCY+TQ)Z/[+5.<*#?2D(E[M9!=M DVMM$)]L^L4Z!R\\O-L9
P*XI,&_<=@0;/B## O,O+::5T^Z1TUMR5PH2EP$Y29P$OP2BG$S4UVA,&!8KO3B%6
P;A;&9<GGQD;@=#C3KNP#/!OIBV?%U\1AIA>>0$NO^@:[G%QG5><::;L60F4/M R:
P'&G6>N?!XJ*)V>#6G$">%$NTC#40M;F4-#JN.UHC>68N,&VGI#XOJ#?%'CI:([,\
P""XRYM9#4YDKNGG O<$]!M%:D60;@!4?CS 1!$D1@7WTZSHYZK;A,1#8)%J6QBW>
P/[RS//P>1O-+IUU I[>;A$GND%B"::X_8N3E\ZPT\MS*WX.$[*S8@X-L\ZNCN#+?
P,>,Y0%M3'PUF_$QQ.HAF)+&^$E%==$C4,U\I(US $@XPDC46"U\?M7Y4F\Y)RBRH
P0KT9IO..?9Y#!UCFCE0U;NGKTAT[_]NXHM]W[I?]K1M6K C /?_4NQ&E]^S1V =-
PX5M0P$ :?ZZ#.*#%K"5[*%66C=BAG/%3^$2G42OG;8T^Q2(!8V/^DX0G3J$02#R_
P(STC5@(]ZP<%AT1;-5NU7V/JW4K2#Z+@4!)4WR#[/4*,;P%'F 3SH(Y<)?I%ADK^
P;YS9*]8@^7GP"4$C9.;ELN"T72(CPQ2_#V7,*UT924[Q$+3GEXRU5&^8#JTF_JP2
P))^UEG9;J7/JYW;%D8WVQ'VOYM5DU_B0:?HT&&T.(R,#5/M?JR&<%"?L&_5>"*TF
P)V6HEM"U:QR4QA"2GOENJ,2[BQ6RV"T0ZJ8)U.4\QD7="8/YVNC@PSCFVF-\G90!
P+(!8XCJO(5V]>H/ZX?[)*!::C;'B29+C=]-[%O4>>S=;%-,/<78P1E:?V#6;_7[;
P;,34 2$/\I4Z#33-)UV4K]7A-&.(F<RZ%]7(H$4V3(("KBK$ 9VJ&HJ&;4WXC&*1
P+$3MUK8BPZH)&D@U,%E9+%D!W.C_UXHA03ANGAA#O!_$X.9B3</*Q[G9D";(I8$K
PGC)B@Z9?'^20(;N]?I6"+,;9]=()Q%A&K+HJOR#;>(#RGM WFN31$AB16]&NKOK(
PFC)8Z5DL@B^"[PRNK\^U:Z8D77G*+LRI"D!QB-'JBZ*V5Z?P:1DI+92!S6!?$L9"
PT>VPHG):443-8JY<B]E+S%!WB)HRQTV_RLUZF+V%VO5>=?SSH-O>J9H_A[_J>%,0
PX,2%STQGI/GU3)'Z_+Y,8)D60E.U$R.HBQSIQ=S [GLO-S]IN86_J@,\&C5HKKL*
P4<D\Q2-1E7=0$,JL]A5")("/ _J3 3J7MT2W9;!H?JVQMY6;H)HN56$T!5%F-!^_
PB'6_0 G.]$18&&!J*9>\1.?A2,1N-2[5+/PBGVTSO$LN3 %:! /4$O>%@HY83\:M
PI:W[R].HBI:$Q?::& 9JZV=THOMY.TCRG\/U(H4I3:9VM*J5N2;4U/MMI,1-GN_9
PV2;):0R(Y[(\HG)#]@>MRODCH!Z=#C_WYHT"^NMWS3<J%X@)EDL]&!(.V+HL>,VZ
P<G:4O%?Q%A%+.YV?&O^;B,F]E_X*(T<B'F:V9#N$?":1 GQ\"I<\A;8FAA$/YP@4
P1[RFD;\T<W#0ZK0TO/=1$-:LXR;/'#'&Q,$,/.2=$&AL)B<._HP?(Y*)S.YXOKY=
P3:ARU5<C?ZF"*?7RX8M'P%\J(><Z4NI2/"- C_*"+L][F(D&K=:YU:QYHGS/E:*V
PU9-'H!MMFZ]S5;ON;E<'HOQIFGM]#A<.:+G_W0LF<G*P&>0EOK-#%*>9/ADWY1VC
PLOXJYZ!1^#10LE-B3F7#TN]5]]/@<=V%83?^[T[N%[E(NZL[5&]KC7]46X2J/$DT
POUQZ$'3SHZ <'G<.=O+=1JLI+V$75\JPRF;9O="AM-FUNYP1PQ&O \IVIW ?D>*D
PU;EI%Z&&KO!I[@/D7+8QA45+/7>#/MY@M^8BVB<69B5"9PRV=/D/)TPR,V4E3%&8
PJV*%?6WXW_P?AV'1.3HCT*O95@'ZM>,11_VLKZK*ZM+IGOM;N3>>,62>E*8PB/2F
P !Y#5Z\Q$*0>2>'ZB&U%9N+*#+@VJUO#F^CDQ8;\$2:3C2@< /AKX%H_7E(Z3%1$
P8[1<+;*6$PF#Q1OE$+42DB/WV,#S&C&KV8[A4!DA8MTZ7A^9O/W1&3$ST]D[>-J>
P]AE6&60]JZ9KMJ^"))7B_#$W;.FX3 H$WV-6EQ:8X'^&" UZ@2Y&@%'@9)8S5 L0
P+HA!_!SZ5FRGP6]9N6R<9+R *+IDVI$B?I,&+&2"]R3NAWD@("=1J9;@P2CATYRL
PGU+D;?XACLKZ"@&-;-Q]NS-UV7AK^BUQBUF! RYQ:RM6!QC?_M6*COO[;<X^L)H8
P#?)#;&?2]S?<N^\Q>!CW"+W\I;!=<W5G/P!]G^,A?NE],;\07[\A"0QISV\S)/96
P-H(/4]/1[U8]]-X((ET*\7@R^0O'Q*'*M]]4!7):M]?70%1@.:RC!N"+ C<W+,+V
P9&1(8)/!B8NRN.]G+)M7!;/KZ6U[4:'()+Q.*OL58PV8" 7,VC9>J+J/V^_K0K&Y
PT=?N>VR PXUD48*P=._AF_,^ S*]L[_#=MN1#-4,\G-H+:D>,MJ@VV?L4_8&8A%:
PP,4H(L"406,'"-Q<R_QB:OG>4O#K+!O[1-AX>^Q)G7RZ5YX"UPPG3\:'-?6'6[!(
PQRAO-LD+/.O*-Z;_Q.8 SB,%((F]WS:.<_+@UUT)#3JJB80VZ)615'F.B:%  Y8,
PA'(>3\RZG59>/.]!AH'P#=_]+ZLXY27\$+-J>F<EE(I=\Q232Q,X"I=F;7B<<E[L
PS5E%HG6);7ZK1?(I"K+1G)N\P^/6YHE>#F?<7 (O%*C<Z)+:=+R^(+ECB=PYY&TF
PC&=YGRX2[^TXS9'A[Y.MUB/HW& OI*C<,Y]I(A3Y3VO"*\@1CO*(8S+KF9< UP5B
P)U4LD!%HG.'8\:;0@="7R (&\&1G]I7>\9F\]B;QDO#IER>VI45!^@IU7XI?Z$AZ
PMUD_)<2O!D4X(UN65A%71G1FD@?0[TP.\$P4*?F+H D+[=:2)9L:4&^HI(7/'*%>
P0Q]\!@7VLA'R0N#;=9+^S4JQ(F*@I$PGIB5/&"U7JJ^XS<A('\A_KW\=EUD/ 0@]
P A2&C,=#R&4GWVWT+C."/W$[A.LQ[O84@B7 B]G:I?D,O?SH7AR5$XG80/P@@EL>
PQ.+WR*JUC[=9#/<()HGXH!2^<HP/[PO&=KY35X@$*$VTH>T[$HZ[:H@>45X1=U"B
P:3]F4.4.]2@+0'@W[',_A7)_=1@M3'_=TS9[0T: C_,C:MFGH*,D\@?IT\SG*<[)
PS727HF=Z2FSI$5YL2!>BY\ EO?/RM5H#EXB+DA7UX([$SF=KF.;MCXI%?:(_-@V;
PRJM6=(#&"?\'UG*!5OA6<MB1>X^_(Q<,,YK'\0>MV'=39'XY2Y%]=9\=WPC1W?!)
PM.NMFEA'7^+.JZ3H,$*5B'E I,G!ZYYW., _*"@J-F1,E#23:RQ(CN7?NYWN.L7O
P!%IAB,L*&G44PYB@<PP(%HA.O+- 39IY__J)YA(<LNG!H]UV!/?[T>KV@!J2+R9I
PC$28)B_OK%V;ZV-@ZQ+=[QV+NZ*_XSEE-!%'=V:LJ*( MY(;!GYCG %@]?UWY \F
PJ":EL37+/8E=%Z%\6=:+TH9$)4BQFM'>THT1,PO[#:[D/;MW4$LMARJQZZXBYQ6U
P,@=OQ6G-7#N\@@(IM]#GLN7X2HQP.F@DS58!,X,D?$DB!9$D-CO2;8E?2;JJVD=J
P:5D-&[+G?!B?9%O%>5XJ_U6%?RX!QX914ZELP+K%EXWLUQJ"C-M/(\+K=1U"%R 6
PO_<*YKK\S5N>]%"*W\LHV1,"?Q'BO[::/;>G?M0Y,TT4BXZ[+F$)\ZHT^3U)17=W
PHY?,C*!^*6'0%'%MYG-7#V*]95;53BF0F([=BPWJ'3#$FN 7MG]).HK:*'-X>9"5
P5^2/G$2A8DE=W5>+\O[T!H8DF&Y*W'G])Y.R&E@3L:LS-W+BA=%;KCU\,,(,C[]5
P+K)"X5UA)6)=-N#=/:]N])ZIUF+5ZMNK"\-W"IG%Y+U3["WPC7M">9J!WW\'5EOE
PC8+;\T->(/P<MCE+1TG&&>T@<F*9:<2J-A9HFOTK *;:PX(Q>3=R8$J"\C!7[WT,
P/,L621 ]"^SAJ1[,U#JV;I:A'VD4U!41^M6X;'$(.VU69T@PXL;N<.IQ.5^I^39T
P;.A!"6K#!$TYOS/Z"+HY#QRXX<^<Y\2ZZAW$%U2A"FX;3"HP70>RX>2?;.TD4SRW
PUM8%52[@!U5@@[A.\H2R/H_"OJ+C9(6EKP7G9W+EN:R4A3V \4)]S^)+Q@#\J9O9
PZ(O5"G,/=.N/K*V9ZJV*Z'^#246-:I0J.G0F@:U*BA+%&D%$!'W+HY>>U.'@!UH?
PKIAX%3=9.+)V>5P@Q\,HJ$V?=WPXLA<P3\R?7!AZ[A"M$W4450?<'(B+5B7H.[')
P'G,ZXQSNJ2902AXR& %<)L G%QJ;KU]<9E*2::!N)+A":O4@_?9N'H=D-/EGBZ8D
P7LV3LE9:@B19W=\\]YX+$EV,>L :=@WN@";WD6^NCML"D@'JT,>I]L "GYW%$F%]
P>LP4FE_^M^D[GHJ)Z2<?+N_7I?B:Y6$Q$XS !H:DG>*_=2/?=?XT-=ZY,VPO5&Q9
PQ4HN4$:?J9;^P.#?\1R]4(14KB@* O$Y?&YD[%D?5ZX9B6A;I3FY"%K;[739YZ&[
PIG1UU?WHXV^Z,0)\1OJA_G6E'U9FW+B/8"^A>CL"FR/T_T=$H# #XW"<VY!"X^=7
PJ]7.MRA/@Z0ZUPJ9&D&8$\/=%VN425$P::2CW5MN#9NDY;R:M,1==3<^I5EG-"SK
P73F+$=ZRSGUCP7[,X',/[;5R>KY^MG(33Q$7XPO6UO)EHM07PD\$<8?(V2,55ARN
PIR"N9N]X E?[*(L[QO%ZV6<[1@D]T+4W!&%Z$?D.:/[=I^"J?=38HEJ)-A?Z6>AG
PL*5*Y#HK1K!\7\^8+DB=,F%JT\,%U^#TOB=4XO;Q29C<9CK,%-X@\AC8!/V,MQFR
P-!K2BHL$DA^-A"O4P["EH\&R,T-OG26J,]3ST%-+\L)>3+Z)MN71'PS'H6FP)#Z0
P17>>Z][T:\,.?=Z^!=]IL?S%'M;H+"1M"7C7CKE3Z2)M<.IS4:WFX-IGT^$%7C4Z
P\"/97/7Q;_ZS*=\+FL'?<[?5O($OD=XNB@1_]O5=6+O[F?T@N$X=L:01_PA\;+-J
P[)M_#%<GA#ZK)Q)7#!"6G-/DP\AV9'1MW5M(6Z K?1Z9^?F*K*7AA\RC#-L6W#6A
PBF\T'HOLXZ?O_V5>'>Q%M@1"B4:@I!0*P/<Z;Z,6H\6<AI;%8ON^8PLV#\X 1+%W
PF<K<Z\7 -AUI[!VC@*5NS$*Q\JRX%1Q*:R)"LI<8^?N&ZD S:LKPP6JY'2[&4TA]
P,;CTXHJN<0A .YY%IJ=F.]D !W6\#Z:20.0<;#Z6UOZ0DM!O?4DU8O@Z$:2!/VU-
P$T[=;_,6YPC !4L5)W1Y63@QUXK<*?*3A^2 JN^2<5F50>'U&?CU](RF\X:6:UX7
P34GW1"K4C?<".9"?6[VF?:LR3"6;)-R$N,A[T2,"B7$@(VN^1AGL?A&5%JF-%:VH
PDAX;JS$8.JEH6_.VPLP''F>5TR=]P*;=JM;%976B-8H9G?* OL$ X;B2'KTN0!G9
PKGU#].[XNDCR%?)[]W[;BA#0DK2%]H>.]R>7K:K.K43""L)TZY2OA%!#DU/RSW[O
P+Q Z^?5K'#O]3B"[WU4+'Q%VA@AGW $).H@LG_N3Q,MW"4@">ITK?J"*H25>.S/0
P]/$<H79//=!H9%CL6Y[:KJ BQ5^/S,  0!MK<CO*P1P\\7WSUG6-XH9_05X:0F$Y
P1)@OX3*A^PDKAW]1E3X56_/SB2R3TL=P1D=+,(0I+@M5&+_ "P1/-XR<+QEA6UI]
P?+'&W\J8@H&Z22SI?D[O4.HV1%7[3=7?HNJ'P"$1D-MHTBG?@BGE-K5)'<C1Q!#6
PW'5/'+M S =9]JY"&V#4 0 BF/\X2*+-J76O_DN\DZQ97)%SH]C;, I.GHH[Q(XZ
P<EO& Z!]I9$M\Y>&T,(O;==?6X%?4@ _EL @]K2'$UO:%JKJ8W?5 8W8CP'>.)!.
P(2B3HO;D5.P\LX68J8^#4##W1RG]@G<)(&/]8@X.Y<JW.5]","9KS!$8:57K+;&H
P#[30]A/17:N*69F':X.H^#R[L"2N**6TQ]M!S.EN*PU6("F*49G^<",N-XWN48$R
P"?GK5(5B1]<7G4:ZB*^2;O]C#5S6UC@OO5K1XM[M=_?5 7!"7;+,]IN!QF*0+4XH
PB;E85KW:YLJ:92*_^/@FY6J5Y#IS<Y MR0';B\&\#5F9T3H(CE@7&4[WA[F%\=0$
P@8VH[ GFS&$&OP. <C#Z(QH;-)IKHT@+S(!'!$;'*86#L%,QY!,%*EMC+Q.CF@)O
PL'W&&SU55#1,]A0UHK+!\)V&3X7B[F7+S5O'#KY>3_O&LG/(QR(HKXV!!;YH+/+N
PVJW=L/T]1!>)S9>0(B_(M@Y*QJFU4%0#NUHX^#OU=B""^*QY6*M^E/-H>3*EJ"@_
P9S< [&)=+D'1P4N4&3!D7%9*>[0*U\SO2"0(N'ASD57OC;7F;TL3^/6E*-[.]?H4
P<^WJ#9/L.5F"P!VH9CLQKDF"#<3HWN$0,CPW<:V9*@R^__DPF?J3861P>4(XA'T)
P\!=.?]>E[Z-!6LDE#RGYZD[HNQB9V"\R]W &?YC'WOXUR[$/KYDW?UTV?J./;#B&
P,.P^8\9%>/XF;F(-8I5)!'C)O0"9U)<,3GFC4/A(9+$433Z=@#HB;9-7F+]'QC1*
P!(R;63@$HI.=1W^')*=9QSDKZG49'<>SA\I;D.YB XY*_N-*4WXD3*;:8.JP'UC5
P<DV@ZCIYO^*^F.^NW>W].5,S84"$Y>S?"?H6^.T78SR]HR W N*Q80-#O^>!%6C@
PZU.75MK,Z3G?HI#.D[?,?/-MGCP/50[(8F[S'>@QJK% 2PS\4>=8R_.2 ]EPKAY0
P HK,0SMZ!VD (,61"7L>A$X2S_-KW.OS[(O^U4Q9I.<"*NH'-* SRX;C,FJ/R5U:
P[9!C</I\U!&;,PY+>XQI ;'@'H=]:>M1CX_+,RFP#B%R%'RJ<O<=U66J-5L!*O.2
PA\V+X+5)P\;<N&I_/HHPUY27MT!U.:C!N]"'6=+9>=TFQ8#?TM";C>CV/'LH6#?G
P)!OWL/[XFK(](;/L.5%JEC KA$@I*^G&V"L7=NQ3!*D$'F+88[M3(1TH2U=4+YL 
P:NR?<)YL6P9>VZ,SUT"MHOU=H^$#""G[6H_'Y5^HRB5 ."AI53&?Q6H*J"IJ3^0/
PD)+1'OYXF?WCX,<Y9CAID\71*D+XNB4+0!).49LY7.9*?-$2!2/OC3VA7DWTP6#_
P92E>CK0"KH]1;%,VX2(?$<@*[ %C^?KT% E#ZU'TA:?K$C>WAM>R= =FHPTAD<GV
P;3%A;HIT?^N4^Z5BBI^U89NX3AR)6JD>5M$Q=G?]])'/32G/8C9HA0>1""_BY2E+
P"Z8L!RT.C%DG!Q,N&0VV)4E]7:K=.*& M1O]#OFR&?O?H4J0\:OV\!",)#NK7B9Z
P&AIL(1SK@'@)8QA\!J\,O<TQ?)6/K..R#*6\'9O&A^@FQ98RODZVY:?Z\X@&RY%<
P14K;]E4*[M$^G84HK+D7WTZN=OQ9 !*@2,;=R24DP290LH%LS;4<.4E$6.3%OA,O
P@W(YNLK%[9#[N9^!)1C[UZPR$?]9@TPSGR;.53"EN!+H&^4V'Q!Q;9%\]TZ1=W8Z
P"4OGXKJ,N>*F3XJ'+"R-E+,F,*R&Q*Y,W_WW^!F&^=C1<-\0EX';4_4U!HM1](@ 
P009B_ >3RFAK"&;OR_542%>9?V2CJUZ$O(>RPAVH^J<PB+-/1)_WSI]"5<;W>/IB
P"W>;8'#4V#A,47/FT_NM)CXOV8;LML<(A:K"6&GU NIPX3I;.S_@4J15FX5+!WY9
P+9BQEZR:-U.ZQE"E.'D6%MB-C;!('QVV-G,P=A?%ZT/O%77R[F[[74G4&#-&FGA9
P+RUAU+:5+(O6B)ACM>K^DB_3*G:$K<O56_XIDUEH&3S:0,R^()KKH2K&.CC[#%=]
P>:Z/LGSX?\)P#FGU%-@(_^8QIT'43, \V9[4)]Y+,._S,$"L9!A'O][1]D2D9-!"
PS3^'YX1!$-=6UII^YNCXJ+IO=RS %^S]AI%J27GYNI$2G3 :O>YO 9B5C%"#LQC;
PT\4 7G13;8RTJ0CX"*"<@@3PY7[H0LJK!7(+ %8%N(8X^(#7^30WK*(%#5%CEJ[B
P4/?OQ@VGX"JF"M"XP[V105_FLG_PU-9D?^039Q:ZKQ@DKJ 8/' HYX$ZYST,5S:.
P;?"SG<._JSOO0ON>)F(]$""%%FY ON5O3S,"K'7<PE2X"W:H*"+XHM/)9YVG$L3C
P@J%-9*]M,2^P;^-3=!RR,[6UD=.=N/GC]FPYT_HAJ.F_=ND_!"A[:BD=OX EH^MO
PV73N[ACUI# P9D;WR;ER3*VE,T6/(*[)+ZXN8 ;]/$Q[J"EX:8&]?P5)1]KO4"L&
PU%66Y16.92:3^C4CO'1VQ)W--=O_VU/!,/UHXEC>2HLAP+@YM>4-%R;7KZ5W*L5X
PO)_6\:%\/FV+CI(4"_AFA8IT#2P&]"D4(7462T9)6B1Q6PX+VCJ)8.(%HR*R+3O&
P>M\"SP$/?@1.S8?)P%/&/&9G_<*5&T.^ .A"V_5A$6Y@.;YQ[-WI&7MJ"CI#*4:#
P-8):ZQ"4+GR4KTM5TBN,:*?O[I?S=9?PQ^I!=28J)>P],:NI[_1M'+R-,,D!RXI,
P-'Q ^=T=G(TFU)HHSJ,>6@JNDRR+1-GW/([%IUR7G,Y<+?&.)"<83-"-V]D7QV%+
PHP11WO:J*%/)Z[5BD>PX8EL^(!I<A12W>J7P]=WM)0@U- 2L!IRHH>] GY2^ ]?F
P"SUG6Z]HI>>Q0S39GXSI)IARD5X2W\+8C]M_7D0!J+7$\47XVV:^13389319#8N-
P5@/:\EJ]G)I.^<)0,3R,P[ 98>-[]=_QFX?G=IY\6J<Y<WNL .^+_24O)OCB&M")
PG \Q9;YWHA65EKMV Q8E:C"AFS2CN+D8+.OO$PAK$-W%8['I\5&PG=C>U9+14-"?
PI^4#2.A5SZ\(VC,'3":X*ZG<Q3?3V4KY+#D9&?]VZ:GCJM8K.+>-H8>-C_@G,U2G
PBJ._ LI>'NC"G[I"Z"^*3MU2V/E]:LK1\Q;,5$H0)<;9^%>9U.I64Q^U\,\FTA-O
PZ7SS"8A>B0U#^]AFRDOSII.N9&WY4-^%N1-26RQ0(:%4JJU*RI:ZD_>D3_,'XZ %
P.#Y-'7XVOM;X'@0*< 6^N*<<3G09O]L$FIO@C.RU38\5K98%/*/V/%:/;HS2)R30
P]_O^@)6 2PV!$X??L41/XCR3,NW$S*#+CW.T&_!1&@CH9^N4,WG,Q*=TK2[W#7;>
P"Q]M,<YJ"N2B0J'H_3F:ORL0?2REC&3:G'2CN_W%J#2, "IO<.G]LK$PZRZ)PKAF
P.)HW3T%[9#"0SUR&<:_T6/Z)1CKSWO5T,1T%R[U7>"JD:"W72@^Y&W+^&3!5A^FM
P42C-UBK79 R6C\[03%SR4TRTQ_=&ED<@%3@SZ?OG?PS,7-T+?"]?]?;D=U0<69RN
PHT?)859F[-9JC8%9ZO#T3B@B]<+FQ I=5JK:'#D&;N'E1;609!OA.GFH-5/EPQ"Y
P"*%-PMA@7$SCJ\J0KB,RL=OPI60] RDI[B'"CR%+EV"O12+W@HG&YMRWO;C%^YPW
P1*>N[Z,"I8_,E1O,,682PZDG5H%36@T\O%_FXDM=DK$W:[],,-4F%T>Z_MH0HH \
P?4P"Z2TX"6J7>"*8+.=#W*9<B"V$R'\ZL&1\YRCBO;JV<$+DR__2&^6'GSM#'PF$
PI2#9AIYA;/AGKZ)R*Z4?N&-FQ^"/0::5,]?H3+JP[)4EJFN)#%_.2I>>E>A+68+;
P..MF]88@Q27K\+J&Q) RNJ,8S& 1LL;()95IQ:D:$QO$@+/TLDSOB*LXJ:]6#7ZR
P3<8HGC4B 7AU0D?;//T8)(OLEJA26"F0Q*Q!EH'4X'[W@>COR< /?G7FI0S!!/N>
PJF"":1.0C&D^>++S"*L$&,S (D>$.-_&GMDW)SZ_XB\[V$\3\@]W$.>NK>.XYZQR
PZK<^!QF1YR57K8WW&1M&22;6G]+PK+&=?=:^)UI<S2P%E1^9!30KC#EP^9ASA.J>
P6_TQJ,-2NQ>^0+^'7Y:?R^W71'&H"<6@21X 8;)I:J2#=G#W:9U;:MCUW7>3-*0G
P28O%D]6KT4M[@G)%>/I;?0#V==J+(PHP6H,'V7YZ%#1G2S.6D@$]?_*[5CHD,8\C
P)J1+>T##LM5,'QI>E>(NH'GNMWE]%Q%Q)UQ].;-XN3EJHJ(BN)TROA%G6O]RR3YI
PYE^74&H&;J0?07K1FYSYD8CSU @Y1LI"*)X98:15M 0LG22L.;H;A<!/P]:K@FFF
PG+Y7N7_#I:\9&-^\[XL*HHY L/X;+R8;O>VP>7%-@U71HPS)13-?8*G*-K+)\SG<
PB#\+\Y!2<<_%>!"0!.OK;2B%QO,N8(;OCHN_\*Y ..G""9@;4&5=U? S_\9V%?NU
PY2FQ5(]]S9=FZ^%6.Z<OJ42H091!^H06BRZ-LW</?T]= F*?<B.,5^!R;U*H)F7P
PF>5:*39IZ]=$K,JK4'^0L5$KCYL=S/[5TC6-,8%$N#.1Z8&T(]T7&!U-=C2K,BZR
P6;H J=U"ET^CQBQ[?C0'&0VS^L"]2L0,FO8UVS7:B-BZ"-'*(6\X9C53G?2^;"V[
PR$PL0WFYX6)RNR1('-5QH75Q \Y7!"9GE#>75'':)"JA@RZ]ZPMF>+OQ1403!GGJ
PC^=?UO H(@A2L884C3A<QM0M?F @=,I[>>ALE7C+(F_QA[0K'C/,/0 SYMPVF?.:
PD,;3N\W@*IVNZAZ,G5N&$X\AQ0#VHIO;<%GH_5+#R\PRV,[DI@G))(N.VY=:^\VK
P]^1QEJTFV(CCX]9^N(:?P[OZ3+F#^O4V*^1'Y",H\T05*L+17W[J9:MQT YR6G@@
PVDG@KLHZ3 I)6#E0WZ(DP_$*77S :;S'_OG7ZRW4$ZCATS1^F9(,Q?BNO&2&7/6_
P<??$- /41HN]#D=7>61(@]GW6MH!\>>- !;^7^Q('='L9VLHM ?_][.)#Q&JV$04
PJ29*M=-QDB$F0^YU W96JQFE<(C@I@^B@U5#/+8O@"G,8T.(1B#'?L2^D)MQ!? /
P>'DK"2B+*AV8&ONAH"CM_BL;LET#F"][W%F?WO764">K?I)!42;AZ>!%L]V1:.$[
P$?%QURN[5M:#V:CY_S&&A*!&XQW*BR#100>A(*ZJSH(^+=FTG=B<?:13O=;P(I"'
P)O G8 '%58#N^N1X,J]LETH M-M,KQ,&@(6 /7#NG-<."K&KC%!P#]^8 MYU;1_U
P&GXI"0@+B[?W8Q98R_=0\E/7<!QTS]F+(SU<5;6LW"N%73#E4493M/K'6YO+!QZP
P1)Z[S:T["30_'5;%9UTY2;0MQ;FZNX3G>P5BEK()S"F"%._&W&%?B?_LB84(I#2L
P/@0)09K4=XX'@'\F#X''IU*!0+I.TW85[-3T$3F.8<2,!NP#B^ E41IK[ [=+^+P
P<MHM25D-U]U?:@TP^(5PY >$>C.SY;IV^UCV16IG* *G2>=+<8[!@55,3X#$$# !
P._$RL3F%L*AVM80HM;*-! <'9'"2L>&01ZM7L0WB)1%VU!SS=8)2M:VA)W0AP9L%
P%8C_\'JU(L%>$*1">[,!0D"A,8RBFX$S=.JWBO3\:..C0;$2F/6H;G=#M0<SNKL0
P_%;E:A#=)1VI+<X.'(OGU_GA@,:J_<W;;@G>_ZK2R4*B'M()_2W""+!VMG,^ 6DT
P3]2UYX-2[YI_P.0(*Q(8)]M=#<3"*XDVR@$DOU@?6..<P!B&,CPB_;GB#+.3*%\F
P6E/'3#PZI DKB].5+[PB,M)&624S).XI0V_NM]?#%S^'MAFQQ 4P@%<B!;YU84M/
P-?C /FV/0HTU7E@&C+Y-A>C0!=Y$8?$P^P7YW3+D\]XB(*[!&JLFUTEYJQIIQS(Q
PU8 @HX0V>R_ E.E1 @-\>"^+2_#W]EEP2#?4ZF>@7VL%J:'*<M5A$^/]GYSJKK<G
P-]]FJ]L>>=C>AX_XK?VRE'>$X5#?LT1 _N AM^;!CZ68^Z3B7.N+<"(H)N&+9X4:
P?;/PTJ+-<K(<R#"(CW:2,D((]+M X0[%J4YJNG)]<&B6PY$H^=>RTCJV3$-.38F8
PD)^=UB*6=54$$\DVQ6-C!9(Q*W$K6">5LRGG;\.\<I:4%HMX_Y;FZTK,U88U1D58
P O$I4+".Q6C$'!1JIIXQ516_Q%<5>W_!BM3?0!],*W+ #7D[!9/9(!8DX1(?]DT@
PW_O/(YVU*3"M>UVWU+-/\CX>%YTV&#+0&+-2L%CJX<T1N.7--,I4.>T&UVIU&EV/
P1WMDWC1 X^@=;>F'+DG(H&JG'RR_TAXA?3\ @;D:"DQE56L[V4M[?TY==^:BGEVO
PM)*C?@(L2QDDK/,.__";MO;SU2%/Y=N@@*4R<_7#X"/ +M0"CK)"#H!D95R5;#3"
PJY@F,#HBI[^7-MPE'+GXV)TT"%B1&*44@:/-]_UN+WMB">1#E_ ?4\>:#O<V%;W*
P^=O@A0&^/KW3DHFNC/_ QF!VXM QCRQ_M(I>7U$R4Q$Y*BQZ[V%T#U.5ZZ*^9O>I
P0\^ZB?N=?YT"OP'Z@XCD,"P#P2PA8K(Z57NX3 P<N^:E)Q'@83:XP3+;0NZ*=K"R
P*>@^'BA*S,Q""%!"!R,/6C!O*J" #S$Q='M6E_GC/"\>BF[?CA;81&KQKY^3+KH"
PF]\>))7=B91M!1&, 72)-Y5_G6 -P<(RHOT8H#B00L/CW!R33PGEBJO,&STNQ/!]
P*D0G/*G=LB>(@5DZ89V^3[,F-"56UZ2K>>&-XCW8I,7+$ISSKVXXW5F^;?@<V0M*
P\\*F#F[DJY:T@]/4H*1;50:93Y3/1_?2C&0WP*ZH +*L@<(2>^,9=@S*/<9RW[/V
`endprotected128

////////////////////////////////////////////////////////////////////////////////////////////////////////////


`protected128
PDU7H_H3X>>IRR,/N?KT7T<0-(GPPGNX7S)K2O6232&=Z/G(,-RG>ZRZJA ?<O-9I
P)6V2^,?I30Z0UI;:@ -Z?*Z!CS^/3+>IJ7:S9%-P1*EJ-<)XX$9-1.9#9E5^U[W/
PB-4$ )+QO2"V!:33MFA!P0H"[)*B'(,5(B5,GU]A#I^=(. @P&]QW,/I==(M00GU
PCV]?Z5 Y!?6F*MM"#:_9NK^S]4(PFO'KF6++7J01D+-%3'ZNS487BV(L@\8SCFY\
PFIY]\C#F>K;AUDQ2PAUIAK-2^_);?I)_EX"2VE'MI8WG0W]M:FY/KBM1E;."-*[Y
P,HZS/^+QRH^',&PV:S3O>>7_&5Q#OE@SG%*WU;S_>UA)GRG0@M26Y03<[>WY7E:;
PN4>>]#+E"-G3$H&$=L3?BV@GH)&+CP:]H(E)-IU-%;,/DD\ZPBWT#"C<#M8@**"T
PF5%;""K>R# 9"!_Z+#QW(0ZGEG+75&:Q#$#[XBM<82PYH0S&[NGVLWI-NP(10' >
PN&?M[VL-Q6-!+0E41K:>D;%0\]QGL[I>LM1)>++)><A^=@BJJ17C&LM*9GX[X7W"
P-Y/GB/O!S\\4V!+>4H+9N\BT+M,"'QA'16\6&XYT3SY%_CR0:AYFQAORF\X7ZXP8
P4;'L337F_^X#M:$5_UG) DL#.EUBZ6.9=,M"F9ZWJ(][7<3["_KB$=[QR$85KA A
P\S?O>-H,@$&O*X3.'JHBK/S>@>CWH_ED(;4'! WD1W",02/S.Q1/E*5#;IX6^G<M
PAT ?@.K)=R\DYCS7Q[_D]@C;N4VYX7B'RFJZ:XJ<QJK>6.Z(7\P3%PHMHYP +NQ-
P&\:CCPO^ ./Y2=0-E9L*/4N[<!V"]'*QYO%,6N-!IY@4+Q/*A::!"-8(9N+:[ )N
P>OWL-0ZK:*M=X/N-=AHCD>EYVG*C?$V@-\0P,S77(&$@2/-6YU@N=D6"^G*$#WE/
P)H)N>ZX6 U2H0I6(&<\KEKJ28/ )8 (Z,;J0*1)J4PW8.%AEBI.Z?&%X6035 >/K
PD];ZO(LJL<QA7 ,UM'/E][(+)CX\+ 7A/8@/DM<*I]]-*^8Z!R+(>5;!^'7;&X>T
P8'#HI,YJ #FR*J-+Y+P@ZR]Y/$NJXN+(5,D)L'TMK_W ZMQ+/J+C%5]3I5![%"+4
P=7RGE8(PT[6]X";+0'AP3.\4I%7"DI.L&E45U#GKJ,T[9^6T(F??!%JG+_W?_$3!
PS0"9!PW0&"^S(?,C[X8OE24<9JWGKQ/V$T[:B^'<-TV48<0\DLT[F U^YFCN]1'=
P,G)W$+NON\,(7=LE9A"U'R1CO)JO+R'(E[M<-FEU+_3,(6<857R^J$4@K7FVS!^A
P7,_+AH=(5[<6P4U53^AS>G)L=FC(/']2*VU0KL$7;-(LFZG<ODH>I! ,K;=O]$] 
P/;B.9V?N^0R9=<V\!HA8-E8*?@X];T<W97F7/#)O(>/.I6&)2 ;A&WNQ:;C<?=1@
PAM.! WAH1!FESG,P0XY?*A- J/NT7=V/F%A*7[#@RXEJ5GZ'BW?Q,SBVD:8NW0@Z
P.3:MF+5P[[>BE5)CV4SQ (C +,!B4<WA?L""?*@?*EG']&<#;]Q'URD64R <<CQK
PE)&K^?,G4'*4$9Q3WV[5P.79!@8NV)FO?5$\;+#P3*H(S@AU3AD>8"?H<(4*5-*\
P?^CKG0++]S##,_EBIA8$471?TE"'EI2RF>>8/\*W1/Z)BXRBA@UVYYG>@YZJ(]_A
PV;:2WW-KCO70P]ENS>N^+.9WU2,JC^".W]+GF]LA(>*;V8DU@4UO(Z;!<0,,F&O#
PII.>%>F3^KG8*83'WHO[:"0IAB;9'UP$%+V)T:SRY.;*A9J\&JA<%J ^8_H)N /:
P"P&#$.%.#E,$[8C+SFQL@+X,.+%FS+<QX5#/ :N^JXL?M0M5Y#^2"I%*Y\09']A!
P_1#+X_<P7V!TI(?EJMY >U<[OSK3]"374VJJ^XMV0B9V1>MR]RX0B2%1=,&YZ7+-
P?O=\I@HI"$*(D8M.(40*>@@[L:K1NBI%^9!I/IQUT/1PVQBM#ZJJ9E'R]S>*H; )
PPIF<$7>!\'M'R^2CN3*0@Q<^VY!%D^S1/<7Q,G:ZI$0J@T+'(AW_.1A)F#1X_0S 
PS%;(34.6HQVRT[GTBM@EZ:8MKHC^M]O( ML(%N2'>Y7RND<N'7:^Y#:Q/I)C#2 <
P_Z^7XFFKI2PC&^XQGZL,)W$_"7(33$W0+V26^Q[Q!HE\B=+#]5F8\-A/]LLSO1R*
P^CF13'Z$ZM* #TP*MI_WCYJX@,'A1C63[ZBJK'V&2$;A+OZB11YN_,K_A5CW1)YC
PQ*E+=>=^64>&W$;^M.R!P^\#?]J[#!5N\WW,&[0T:W/ZD;+Z$\N%:/S@02QU&<$[
P=L86&KP9%X01N2.!<JH8(3Y# XFDY+_&V>G:S"T!A"&/S%$!1%%U>QYJ(4L2PA/[
P)V>)0E=-?UO^_5E('X1TA3U%S=U:++,HYI$:K1@Z"DAWBO <Y/6P[5H8X,&][QB.
PA9A9<DT10@S[Y_,7S#NE2W]C&DVKX_B,!M,;$FJC[H:7(N0QZ]]$ZK7(,JXR$:59
PNKL@ZXV!_Q>R([0:I[E:H7"P0^R%O>>N]A8'L3/V=4")=<$,PVK+ ?4W^;NDCY>$
P7B#=^=1LFN:--Y9IK!!5T=P'!&.TT%&);H^S8Q(!N)D;8/@O B'T&Z!N+7,SM+2G
P#1O4]A^"RO  +1]" 7XFY-J1,D:AIJ+5P7CNC7".];JI<8+G:>T<[9"(2ZZ),842
P'VH:;K0P B4TJD5<RZT&%MB[*2_5 5JSR"LOQ)SH@D$X#N,J#7U[) )3QIN"F\9O
PY%R>DU#&<28%@XWZ1+S<7_Y9K_)_"OJX1BXWZ4'RP9%"CYKL"OK&+_/N([Y*SYUO
P&:3777HYB"9P2]7EWL-V0A^Y7+$PW;<Q*NL[07,37Y2UL2T4/^<K 7 ]ZE0XP3P"
P'*0R!"GS:(Q=K)WH[QX?9M:<1ICEAM4>L/F +6W9[]@)-G,T$S5'75LEST(:#IKI
PP<K/WIX[Y4S4 XY2690:(U6Q%R[","AL2> 6V@PD'L(1LMV!Z9237E02$I\_PB@J
P_$IKEA>(M,Z[.(](I*G_31Z'[#9F([A=FW%'=7'EJQ S_\<KTS,TSG1L)I3 ]HQP
P1W5<K ^.5UK.UM3<,.O?K+*LV_E3C$,Z:^IHV.G N>PA"I[]<FU91=I38A@L/$[I
P 2 1P@[L)O+ C]LRX:)A]P#JDET1![2:E/%%:;J7B2,(@%14X*H8CZ.5_S.^4Y+D
PLUBZ4D6DWAJ%\]6C7^0;M_1*9#\#'?F@PBXE//ZYA!0^2>;[X=+(M=?6;7N;/))5
PHL,R%;X6R)N2LPFP2E@;Q*")OY36;:X5AH-V+XT;!*"'H$(+_=^!ZE=>DIMG*\$<
PM L^OK&A_VD2.7\\<]K([G0>]UGOB"1PHM)0]AG>N@+[3D8:OS0@#BQ.Y\8 X+=2
P&)6OQ>#P[9Z*%8IKD%HY3YO<RRS99,?4+R%WV \][ Q"4S7QJA&$*H(WA&Q0>8J!
P$&^WW6[_FZ6,Z1X:K!68VQXFV*!7"):B_;-NL=XPBJ/'AF1$#^M"*L9EG!LD >Z.
PHN:F$UUA'R4)UA90+LSB>R>P(FFSDTD4F@@*3[-.A5A!G@\[=8*P&YM%;W'\"56S
P3![0S:/O@HAL1Y"J4@^E-ICV/D/%0!<MI&=L5G:DJ:O<98A_NXSRQ8-.HQ-$DI^*
P01GRU95*,+YJI^-F*3<O(_*;<6I_>MF +AQX>9X7UX5]3?H;YFX U$%/KX@*I#W.
P=&[)A"]:UQ-5@I#"$(A_!CS>4#*2V%IH[I:3/8*/40RT\PNGH&^*;0>IW?0"<'"A
P3*C*""4I9V.)9Z)WP3N TTZ&-8[0(RFEP,;DR-YYU+5OM3ME4T*=2 JVCYJ(2O@M
PXQZ]U=_Z$B=-W'TV64$>8*Y7!/^H/[B(Y7TC"$CN"^ [P+@&#DKF"Y+C#!,4"O#<
P7$Q5WT^3"E>8P17\!>(],V^[F$SF\QD9L4R ZL@WN08\X">Z@Z5$OO\MN*CZGR1#
PS)NQI9>;N)>O$V)$:'SXI_!6+XJVB\B7"3=#9J(X>9JU0<3<JXM(INSJ1]R0[Y> 
P3<D0S"%!F$5+<TT:-JVK"0U%2:^T48?C6=)LTLO("K?%S?/0&_<FYPD-))QAN1GL
P&HI ?R3*X:?WV4*'/Q-8/VR$ 5.0-F&VG]R_U[+=E'*=W#W)//9I24#%1YU:-8/W
P53>@4N 2)=;U<GA+OR<&V7O<K1B<_GW;W]<WF+"7JP>L%>(>WI=0'2Z<G!ST1;J^
PDB02^6)O!'&IZN[!6/Y^7==EU,,J?)?LL\TEM"8%'1YXZ_/R .B@P<1:I5Y6GUO&
PH%=3O 3LT#6:2#"*Z  L'.B=N*-#4U?/((?9L06*A;5L$S4N'&'V%80G1NC)@2_U
P\,_O7WH9*RRT= ] LIIN>?D:::D>!(=@J-B#) ;T?XWN;3',;36L11Z_!WG.*R*H
PG1%L9K#MTR7>A!;:]%*[U(B_@*39H_B<F=A(:F#%HH56CNHI;LOJN30W/R@]Z,8&
PA/BB'<\5SN3E$0^O,UJWCETDB:"M\0M6[#&)5WQKGZ. EF^TE=.E_X CYET5#@Q'
P5,P:,472VG?.Y#;:6MMU#SAMP<UN7V.8RC!W/51FM_E"2?^UE"V*"8 ZSY"S_M^%
P;,!?E4!FM]P+N$@;;^('R([%%-5EYGLVE%JL2W1@C]662FX B_AHY9S@LHSXOR_M
P*(W+"U/L';'!\:@_Y!K[3+?T$:SLD].L\ I]%*E<K!BXT*N#$9FOQM<L$J\)8L9S
PBPZ 4*K,89SN_4WNU28AH;5,8'_<SN#Z>BMLEC<EBQAW2C$/KA@)(.[9PYB?+'U9
P6$ZV\.Q<G]$ ?:JNW3Q#E9[=S^2J8!)O')+T@7\>JV6$8@=J#LW.4=(&,XR99W7<
PIJ"V9>>H*=X@,%HJ-Z1_8EW^^\:S.3M52H*'G;WZ-H+[*8C4W6QBI&7JXKL80886
P[.)D$AJQX.P%QDL/;2ID.R98_,<)79*:CU)"\.AN[K<67;)+J&9AVWIZ1J-89FC9
PPC'N#9*?$>'%K56J.::=6:B/AFC!L_BC*'XR/&A>QI(('LD^LM^09;FR%%?2JX=A
P:9 3.*)O#PA\ Z("K'W=X*4)N%=HFIFQ0L/:KY?N L[N6Y!\$]/F^C[#S87(H@\,
P-$QX6#&XX<!85'%"J<GO[LZTFP\_I4>6<FBV<"ZE[+;#;'ZNI6L\J"+:[\8F *0'
PL4>U'C$,Y=(O@>C]O)8,\)/_X;_A94?$2""8"67$TDC*LGKXC$ VD( ZSB#^0T&W
P =_,B;H_1Q2JH=V1HI+-[_!D#X<GM]JUJ5[%)<O#^-42]>-CI&Z[U]:WUNI>F*$'
P?6ZLIBDF#Y Y?D@=[@Z3^&G#;WX$*JT=AUI79""5@.0J$M]5THI.&,*UQ5"9 C4\
P4X,!D<$(9]<P]!1H/P6GUB=/4^(U7@S@M?$==J-@& /?>+M#0&'>R">\,>"J\R(R
PPOYWL6N/I@PM2Y/]ZV0^!@Z P\O00N=>]B::-,<]"$Z7VSOLH0S-E8CS3%F)\R2P
P(,%TTVFT&>A<Y17O"%K!Z_K1,1%A0FNS #[RRD)51,7^ A)=P@6"I'9*[=L3-=.G
PFSB0WI$<P4//2@OT97<^?3#NF4'8X8[CNJ><M[X7S/75E2&3DX5K^]^VY>O"*5S^
P7HV2."WX0F9\JK^<K*.T5BC+RS@^Z ;LP@/.;:%[D)7B"W>(LP?@(C>Z-&3B&8I4
P;G$Q/R9/^9?6'-(NJPJF,:3[6SHV"0%;^$HFX%NG35QES!&@NW="*9@L+IE[$<J3
PY[S7@(@,-W)^=JM7^N5XNJ@]R-"%*J@A]C%#@5,ZR!6A.?\I:H^";YJC,JBN>+0<
P$?SUB. 4OJ+(':91:(^JG$LC0,X2DH[$-]__4#6T4SH!A<:-!L&MRH1O=I2-A\-!
PG%N36S_'\90*MH26IV F$V67!"NA2)KF]^STCKC/&'@BP^79P1.TUE-QH4[IITW8
P\YJQTX<97",V_WWP!3Y,>VV),R\$[1&:5V  F *]X0DY;0)>1Y?Q%F>A<39/0,=X
PN.-@J-Z']7%"]T.DE>]ODUBO>9RJ6QG](B>QR(C\D&1<((X $"=6R88X"P4->P^O
PP1Z2H_Z<5D3K^,VMR9AC&2!X$\6_>,,KBD$$R?23MO:$G#B\V0]VV^%M97,/5C-Q
PBO1G"&%D_)W93 6%BB[D3QKLFHH>^'7E:RG]"KFD%Q]V7%MV52T7ZA$.INK/03>]
P\?^#34"]L,9 6:1*!O0N':N.8=NN49W?>C0'>RDPO.S['/VJPB9 %7!U&9^*UQ>C
PE0.*5<3>>]8LC2'SEG83>Y=K9%(396(D:$#U:E#>0ZG!14$)3/<"EO&):IL=>$5V
PJW6F"_4/-+^L-H>>8"H N/G"SU;<1ZV'UP9E+*]3K!Z[^[Z$]B@[61[8.H\LOH#:
PS.1;2$V;G-+8AHHDW!NYX09MLK7I]JU3F*!-@CM;M<<]"JE\].);4MXT.,UWA)?H
PV,U"]&Z->2;4@)F]:!#MPJS Z*AF)\Y+\ X6U;R]1Z)Z$UT=W$0GB(W!6HA&QLL>
P)OR_1M$4BPBP#3U6C:-1)KN$++^*FS\4]KP>[$Z]CZ(*T$/S:A97>ERO"JRMC1]3
PFE4E.8_>'BNS[ZKC\-\%1#2!6RFW='K@;1O76^RS-?/%#KN,AO7&Z(RFND-]EP/@
P,BJ$R+=(_?#NZ)BY"_2<7AH8]G-B!X"(S-*,=&+!"8N=K;/[!QQUP<FU?H_9D*.\
POR[0N"C<L1E,/8JFF"/B7M^Y#*]PF0+IG;2PRA9*0FC0S%+6PXP$G(-ADMVU%UDE
PW4C00](:FLG"V['?M7(OG'PP/%L 9@ZE%_KR+$+6.M[5?:O0Z^6<1[JLWCV*KV=X
PZB]\9;[+,Z7'E&JURQ2Y)966+RS5$[-60*B?3\BBLKHN$H4,MD7T.T3*R\_0& V5
P9=BEK7@!T4[NOL=='>WXL0KQ?E^,F>!/M3)W$OZ%ZCM0Z56EE-Z.+Z>9$+\J4/2I
P]"$M@&0758A#<%SYQS1&4T7,<;/QA*V<,P0:24!3)H"R)T!#9RS*>#^2?:_A6!SO
P],><VQ[5*K+_PH]]5Y<U[BK[3Z[[5Q<,C9X .1N_Q=^B,9J!:RT3S(IG7VT?=U^$
PFA;I2B?VV)(WH@2/_ X[,8IC@H%@B =M=30#F.NCFO6:J08")E X_A,[8V/NL2&P
P8Q<"BFS#?]@J#^&VITG]+-7IY$AD."Z+I6#_[1UMUNCG"]5^Y-Y1VSZX!ES*'CN*
P#Q#3]+-505"L6N:<"&&+LH&%#C<B:SGN\#_N46T-QH^#G&P?:B([+EC,-HQF=O><
P#*7IX"H[ +)9XN7%DC)K-&7B1HS7(%!Z,-8O967*4=RZ :;P?\:<\"_RV+DM<&--
P;N4=[E4XY+?%B^KL';:G'8'^WI^(05?Q%^<&9IWL;8M[_J$F'+LJ6H-/((N-S<EE
P@+>QAO)'"3S:,#?9)ES2'F[8>:*<_+6J3<'?2(LOKX Z523?W)BVCV^=C6/@+?)M
P.S>)]R934>&S,YEEB.I/7&NH> A/"S"_Y]:6D4>0!M5J#-D6Z?2!9@PMN^K:Z!P-
P)CO'(>636H+ 7!YFJ_# ]H(+QAUQ!SV]D/;GU!#A6:;1I5":5?RX)_3=KS$K[=!"
P_:PFY7FAL>AKSJB3YI\2UD3_IZVBR57W6@%^R*JHM*3(?GZ /'=N677ARXRAOP)R
P^%\#3FI:GF]G>5X]+'#1$;Z-7:PZJ@YBL  4A#5AVB[1T8$>7NF3<#QM(V- H*,-
P&DN8KWFYL?KN_T:P$X0<7?0BC8*6/8RYDV4V%MTO'ZJW*9%JR*A;,2]8I:21". A
P_7P4X+5LK&B<--Q,4-HPUUUH.I_.MQ?R]U,FF"K?XN0ORZ*HJL#=!CG%9&.PVV1W
PIAB6*PY>U>93596V/G4(A$%F12ZM2*@^A0CJX$70>\2AU1^[E\\8,_=NFC30%!XC
P>!FU6YZ86@KOIX21<#<'. ^QD2"X]#:'B%AA+]Y %86$J^]%7T#03LK>('=!1*D6
PCTP\E]I:J1$C!V$ NOG'(F_"+9#*2I H[OKZ&/6PC==#/J$G0TL$2JVQHI@8Z?RP
P5Q)7-"'P5S88,=YM;O(S\)<BC\95@X8-A+M1K>U1_SP-VT6:U,@* "\Y#AF6%:%>
P5&;9#R.-C@*KA<TQZR_Y"3K"[JTU*5<I9DJ!"Q*-VWXS*FP8ZD6480'9FB8*!<+@
PM624>LDR#TQ.FG8?K_S&03/3;'#^VW#M<>CF$L XTP[7(R=AH,4_^MD1<][\UPR%
P"G(7])W@1K65AW\YY(94[<#+=1".6\E$2Z3=S; 3[.H,VVBBFIP13%]_;H26D>(U
PP,J.Z;M-2&9V/OPDU=@(//1FP9JV"8"'VQNJD3G;\EXO:\#FV- ,)S5/O+'GRHII
P$/ZHGL72U%78!AU5\$);-V%@\7KF?ND=-"805V.P4W'MX0+Z8I'F2+:H0%ZG-Y%[
PA]6= "-!=N)2_S;S9D1-RMRXW!1>'= GY0YQKI!:&9GVGB$T?[WC?!<NW '1;UIK
P**T@(C5!D.;'<J["//#5%T9'NTQAVS;Q=7? ]@ 7?4"4\T7#TXU]Y$\2 V128!K>
PLG]Y8?@ =&Z[N2I]X-W/N2UZR>67+LBR2)R-$2$J4<7RIQ?-45:RJ4?H00@&>CAP
P(:'T0+O\1U!*HZ=!JMQP\D4)#5'GAJ?<9URME6/'\%)N@.<%O]&N[T>O-#\I(EU3
P)4J[,NJT/=LLH:+$C]67$5[*/'&*TC??(2P2PHKB?2& :FNV,%FP[ZWKJS@J=Y>Y
PF2=8EQIOTM]8,8X"ZKHUH,V5M.QQ_=;+T*"*.G$6%C18:^&/45E>2JL].;R[A\MV
P5.>2/&D^$KFF!1YJ:I=7#NY'/\+W;VA4SB?!5!Z@5)"JMD)61<221Z0;*FY/\FC;
PV*<_=S_89U@41M,&93QK.6<%A,Q#G[@_L7*%C2:[,#R*; ZZA62YC.WN5B)NFY4V
P&L4=Z<'=O(_"!#AZ<*BWE/ !M]U)+_^O9>C3)TS6-'><.R71<1G8@PT#9"6__;=X
PTU.A:FG*!]XWFRZ4LSM,,R\/CN(^$<PW*OP+G'<\#?@KYQD4/XGH@;_,+K*ND^,H
P-^M"#T@WDKY)>FZ2<[^0"W@Z9ZHU()7@Y$M9Z,Y&R$;'\IP/3V0,N>&%$U=:_,1O
P899[]*&W3*G^RD$@2F#8]!%SR&B8>( N6A^U[^\INBTC^-7OM!Y7^#%,3=.WL*[K
P,V5K+VJ8\UIPY7N.84X"$Q6*OW#.3M%K2PD[6&"8]UGTWNLT[-;7FBD%PIE8 U?W
P-\\:^_@I[^K*B_0(S4BB40[_82LNMM@9T& &]B_-.\L.M2B>!B'NHKD]?8Y.N]C]
P^Z"<I+Y1V1OL0(J\5_/K..HKJ><'/VADO+RP\%\4SUYD;]0SAH'MOTT.%PXR7Y[R
P8O3Y0?C*;Z@1&=2R"(1E=DP]A$>:$3?;7'+ \</K)$ ;SQC:>C42>PCTC\620>SL
PW-PQH"==+S;&R9=,)2;OCCX[&N^%VA$/MA\IT<SU@J:[K&(]8CC:@W[:+1-:?D=Z
PUB8TMV*F&&-3MASC6JC05/52D!7"Y;7/O*Q@@=(ZPE_ E_HG_)P/"YALDG><HI8&
P#(CX$?0BR<+H9GPX51O:M-*87$2_/'E8:\J6,Z@A$>*)DN 22/0R'1'/LD65;J6U
P+U7X"=9/6(MV'1G ?>TRPS0('$% IF((S$5//T[G:^*/2Y;6.5"^/VY2G4UJ^J- 
P&\P7)>*SBQTUN(M=BEXIS"A51-2\/@H'=ES7AK/,!\X?RS??HCA9!CF-@(8.+6);
PYQK=@Y",^CB<VG7X^\&-M\ 5'-A-?!AM\5^B&&4UJTMG;)@2<=!H^6:]&R\UCJ>A
PWH'(\;>M<<.R#MAHPE].M _S.^6G8SQ4A5>'SMBFM 7QT!@?U&N;97%&,:R#6H>A
P#8T5U]RSO)A00!*E>D0=F&?!.!(#MB E^<=DEDN'L5;MMUID*5_==R3DNOWJA#'Q
P@\2*F<6YPIN%0(T^&.@? ']%2>'K.6NNT<'M.#/F=0#70I6VK4,/R9DQ=\$C($X:
P!]:^*E*?03A=C*8RQ(J]FJEMSV17F$FRUN'XKWY,M#/@+XO.W:# 9RAE,=N[?>E3
PTJEJB=.@DAY40Y0FQ@W<B<[A3L3IGALJ+K8V#B@.Q+N)Z7EV^5I=F_'P*(:!C]"E
PD\WCHO=#,B6,"KCV[E=";*.V .%3, WTWL/N^+>EF529K[1&E8#_>HF6F7)/6!+#
PKP0\E*%I+;':T#T'+S^)3A:-V.C-& JT45Z A9&!")8-:MDPT'IH2?8<XSK6()R?
PTODM?!'-#64GFWB6'K<SZML(T3"'>-=S)](Z>R"!0G7F]FEP^,%?T'7L@-0D NP&
PY8.1<ML#,H0:]4)0???# ^"N.?AWHXO>P/R0X_\- O9CJY\.F4Z%X]6]NVE"5\SN
P<Q<O_>]!J([QTX^/&ZK[,AZ4)?)K7<=P82ITQ4EZ=DJ[KU4?*S%?*G5T!.$84#9^
P_5-,;D_4IV1)%VT'ESRHL5UOBG-WK\"?6D#UL)-$S&./YA+KJ)B[XHXU3(S<8E(H
P9KG8SW]!1Z7X:-C@T)/J0$1:(:E?V2BX^\@1WM5 6,DQD$ 6M(JC LN ?CR_#-N?
PWHY[,4Q%_?MM-:"-?WG';D!.7"M6!?>!%#R%TH'$W_UTF6&OYB"B(>."0:V+H%;H
P:7XCX \H]!\U[]ZCQF?Z[$N]L/_KTZC(*'"8>)5ON<S58T9GR4FE!BOS-ZARGXMQ
PK(A J_7J>"T/QFR7+^D25F 2T2)A]_6$3,8K5_['M'1Q'H)V+ER4&$#P&Q3%U%$+
PHQL>A;@IM1;98-CSL% +K*V ':WV^CF/PX?UMUCGUG 6K>>K5((C9<.C 4:%9N2O
PA6^*ZGH;6;1TA.,KO#/Y$NLY]) J,'G[;6HQ*]U;=3:=5-@&)!ON93-E.IB%0I ?
P7@MN?N7*WT%N)EU,KGT#?#Z'],M0B/U*6 ^0(8[[LZ_*>W;:V??]86.Y1LD=W6D6
PR%'XC6D2)=4-[#7>MW3Y70C+7I>O@W?F4U&K8Q<V8@,\C4M/ZI<*H8_/UVZ#GR7K
PL=N:I?FDI9@@9$ _.X"AJ;5.ZM$1]6XJ4I]CUSZ-_"J32E0!B@]]"L??\:\W_=-3
P-1@1J\*1TD->N4U]4=;BZ5Y_5N\R:J.$3^'@V#/T(>"@O>9(-_9H()++/LAI>MDM
P]SHU4[1CA8!L,170W?89K\C!#A_QYM='S_/Y?AB:D_KFZUVUEC6A%P$\>VAC0)8K
P=92Z?MZ2KE%E+$[Y /83H!G=W%K^](>Y&6IGGCB:8S\R(4M)^/'1BKM#8DDSD@:>
P6<?T(=_$695NO5#1"L/E9"&5<O\\H)KK(*45/,+;B=R!%:KLHU2*2CWK'=W3-8=1
PS>?C!TYX,"K3X'N-45*8OM3^0"L!!1?V9(#UIJ$^$O]=OKJ%)+0]8_A3C^7A=+8[
P6.KW7SO[.AZ'VI>U6*=I8C&AF_9^$'0M=EN];L\\]FOM$4&VG"-SP[AHHI3PL.T[
PL*S&(9<-@4I)I(HIL#E,*"3AD0N31P7%_NI8Z"B@[&]U7K351,5]GA/_"]:5_ULT
PS"_? =BD@:^=T4./TN9)4?FY/Z+V>3J_%8*DR<TX;A4")'>TO :FC-$P\ -E"-/#
P%]8\LS%;!4"8T^73*(.HF:_@9R!$3[Y9\;V$CBP,;V3_&NVB%WX/<%%Z0;'3]Z$[
P<0QW,BM1&,0E+OXMPZ=D7_N![]M/VAGP$1^[+Z"^U:)%3C%Q,0H3ZFPHF-F:T2>+
PY/B3@&WY*7Q=[*G#(U\7/8F%I7DN,L_HWH^EO%=7S'CWBQ<N9C63"D@.*;[N&IA?
PT_3I6.#:0.94R-X;QEGDU=0W%!3W0P+HXX<7CZ*EI\PALM7(8.)J[S>?/2WSOT6^
P(726.FHX^96VS#))$<J'C!%\3+9GM-#+*>.YK<3Y7@[+GF#CMY, *NO)TC;'X<:;
P.<R^IM51393];O1JQ!;'63KPD/@49Z<3<JS]K]D_#ES20@3D8JH;N3ATHQVW2Q]?
P37G1=E3[O\7![^.BI[6T^TDN;!1KN%R #/EJ>XBST;AQ[-IM[+Q#A&[ FN]_#>,"
P?HO*(=D:(PIS75 T;QCC*ZSN)JD,L'9,:4I#8X]2)D5XK;3W,UTD&'?5'02A7 =4
PGE.[Y,?0,;#BLKN.@;=.5A-LNB30$-U!;4+WT-F]Y!QIG#^OMW-1%8XY+Y8*O3!N
PH!XY:$E: Y/+IRCG@H-G$"Z=,TL[40=1C0/NWR\P,RH8N<8B@G,[^[90B.G3TU%T
P.(G6FY:;AH(08W?KW[)7X/%HB"QS;)"9\KJF(:F<DP0?^VI4P.;\0G#E/G-5 _(/
PQ(;]^+77CVCX)T6C$S\,0N:=*LTX+L4-\0F)D!*4!3-'%HMGE5'A&3&.> V0+WJ2
P"H=<@%)B!'UD]C!?E)D6"N:,7OG]H0!OELT]O9;2-?=2XD)M)N9F:F5CL&?!IPU2
PC<! <KUAN$C4-9'X1&#H1(P-AGV)^!*WRS)<Z-;J)@O;,W);Z(CYRQC4RX& =@1%
P0C\YF0U,(]S'I+_B1?1=.*6:(HZ5*JRQ(B%3,&7?*LV?&+[5O)E&JI<Z)%J(\2WL
PH;3#-GJJOF2/0/ &?<8XB:?W6X#_K*NIUEP0=TJO'2UBP+#'#VW'#)^"4B-0V, J
PR#XS[:6(\\)^2 3F)DF%X]9P\0_L5ATB=>MG$H%!$/HSS(!6],O*%2):\3'<P,G:
P?"6F7==HNS85;@JY6Q4@C?(T=QT+K>03%-5URVGAS[,C^8B2<26Z ^25K+JLX=DC
P=*3H@ <^2,O,8,0NLPH*%6V?AM^D[P\.P=;B6U,'I<KZB887=%P('D&M/&=]19J'
PI@I9'$;>28%7H8RL+W_(G9A/__3'T'#H#K4-5Z7.D#Y0L<@O.GN$F(O*O+R-46:%
PM\VJP68Y-IYJ..R/DUB;0LPC C RZ?31GJ1D%&9B$"?AW+O8"UV#2GXT,'B0N*Y7
P$CKNF).P.C.=!P8MX/T ])N4I3K8\8Y+^8$A'<:=E1S^8K.BFQY48K?@2IMP%!WI
P YZ48,C3AC4\,I2)@K):D<]^_HACQ:7]YAPNYBX\T3;8=O@66.%Y:R_UD3H:W9>*
PF1;.7"E 0#;;R![2?5P-B9X_CL\R/+BCUE=<;G!J:JC<QCZ'L*>DXH=Y'7LC2D;&
PQ&1KHI@Y(Y'*4TJU!H[AVNV.ZQ1X#N&1VMDL:TOF)!6P3SS.[<DC>="1'I+%?_G"
P00:]T.IUOND] HS,AO9FPADP,V5FNN&' FND.Y>'U,K<I.N]V<J4=;6KK>NL:#T\
PDE=%*Q@L /-8Q,T^8&A5GQ-/0L09$TO3XM=TM#E'U;NV 8/#X6MBJ?%YG)):X(\"
PGAN>;:!PNR6<ACQ:@_WP.')M/D?U%K'5I/.6;PLJ33(_85I?N)=E/J(6T&KW#E&"
PP=MLCG![=V]ID><1OO'OK4-N "_$6H-;VCZZ>0G,RX((&RKIW1 FH,:X)JS.6KH!
P4#"R$<N]+)T&]:K>6@8&1 D*BQ)_C#(URX,821R"7<%._VD7I:YFD1@!M\JX.M\N
P?31=9OM5HB_*:AKT6-\##71F1-.]?R1SS)S615YC*&'BQ#V,%&$H4*:=\/W;E"L[
P?PM(*F]ANQ1+Q)C&B%X[:%N>+$S!K^=(M)/WUE+#)5PH&"N-LXJCDVXM0F)5./36
PVA56H0"$0R"B#0C_6/4YI:+><VY%,58>,^3^+\O>T2PL"DK9VL:<;<47AUM"[&D/
PAO"N[<-0=\O0HHR*$+2_98209P,V1<-9&J.\?I'$-^C"^P<45?<^]'RYYQWGN61F
P=1ZA-4+5_E)97RJNW0Q:&5#\N^'\5/+I+2S5J3!0%<&M94P8G/ASI+P+$8O[W-F<
PE<9[[H=/U/PMP2T51_I;[+9?'\=]N[.1J*4F?<*Z-T9N<&_MC4Y6PVO!MU&7)0O+
P4?),?ZJ23E%*.MED*Y)"9KIS;MM.9H"'!N5P =\H!G!/;JR9_ "&W*30M4TR;J=U
PMK2DA<9MS>;4:\]>EO!X8;/V6'M%=CRWF ,I\U0Z5UNK1-(;G&+W?+FA)2)4K:C(
P:E=%Q;Z(Z4X$QQK;PUK&N!6-K4DQO(SXZ>S1CZ(UUO+"CS;4)<C]S8)T+XM>Z;["
PT[%RWQ@I[B3FHCL@ ]80&U#WJ&M[\<Z(RW1X@,UT$?,AL%E.P)',75)=OT69]8>)
P=^]O.000X!N[CJ7DWS9^%I1__'\.K=GSE'>M5534!6]HF$-UTWY;/$-?D,&*.'W6
P;)^X6I<8#.\^L\*EW'7Q6#'QOT?I2(CN($>\&! X"Z+7OM7#F@TV8:35BOR09+@X
PUBG%\^7THDZ9,<R&EDI)X2G_]2?S<'LT$476%JJD8[DBIZ0"#(TDZ)+)UMR::9(4
PQ:NFV/1C&:T)$Y8\V]73SU%<_P.48OO_$VMN;9-?(Z=*1<NX*H[$&%F \J.B\HDJ
PG7[$ )5JQ-!W"IVG+@]+>. -+8;!BX+CL3&8BT3K*G;Q&!!PK@C!!FAH>GM$$N2'
P6(,A)\)5V(7R]NC&BCP" D$^V0SU5MOS%&9BM .@Y0*?3:/"OH:(M/UO?6%9R\V-
PGX%ISCFX*[477.BUW,,*BX0_&A=U%H--&3HB6$J]V5$#%KXC(>6CFF,;UKC/<2G\
P(_5 >,MI0.N*V7'[%><EV\8(_LA%PP[B;_,$5H6=^RG$;34S:*5K+7J?TWT4U-H8
PB4$Z#R\=;_:!L/B\^T[$M82F >P +R-SBV*J\#Z0?@BU!\0 R2<YJ6.L9A*1?XT(
P<O8/:!<D\WOR1#VIVM*0(2$M+N?L\G.\<NC4!24:H@LCB'U!L%H^B%WB0(- @Z]E
P)<&-UK2FDVA+V[W2<X',GT'KZ_<0^C+98> *L[4FO>B<.8FG.,',\@U=S>$>O?5C
P1S:MX+&(%'$=L7,O8!Y$;E\8#:]Z 2=[RF-KHI#<CC; UG2N%C<\@VEN(<*:DQ^>
PBY\?+A;P]7/6\7(5YL5U2. F]__\P08S)R,-KRR<BK?\%.Y*#YR\V#Y1[EI!4PT$
PJ*TEE084&&<[N%F;@;<;)C%]19 GWOD+K6NP'NVOB[N\<HOA_.#N3]O#R)*9_34$
P\+A#9J+K+%/$2V9X3G"S0@PV/@TJX;':DN@2:N:R1V ;(GY#M,#]4I_DCJOTENGL
P9(HJ2S%?73 @I;,WD9?J1NIJ6[1LBZ:ZH6%G[+8)PV3DG]=[/R,P*(3WH8 &B^O4
PWL?ZZ0NN]OBI@[1G]]U(SB:?CDUU \O_LYLV0L"_/BP='$&96.@C$%W>=CDY;]]<
P[X&:<&9YZ95R3X9:WI:\.?E(4'\WK[52!Y1AYKW^=354+LZ"MHPRP"@BW(&@VM:I
P4&#5$O^/FV>^A..'XDAPH:8#PYFLD%?NS@LNEY'58]?@R$*VJ.+719KAJ?_ 0!.D
PM M'J19-?_0C-K?0>ECW,I4MIK,*8(_OP0FA05J4Y'S]56(+6*9ZV3/5[8"?8(#G
P]_Z0*V17'14[!Q+\?ID* \X/ORZFM%W(N8;TR;P&?2:1XY':G5=1S7UB?)A#/9(&
PWOQJIYR(L7N^FZ2/6'"AM-W.^-'(<K&N$S")6)+161@!*E>",GIJI[7BVU^$[&F+
P"5?S3:YJFCTO#&YN>X21[ZU9I-8<*L/0-UV-$W"LKW "HL58>)-%-SB!_!ZDI9V<
PTH^&3%ZB\MUWA<A?4[;*, N2HG8+(NR@8??'%YCNFA.+"7[ 9J_'XI8J.#8_X1ZC
P9A(W*)YE@LK)-#;TSF&;1R<U"*6/"8)3^GYJBN:(JFBRF16"L=[5SU%E%NOS:'PS
PU(O,@7C +-HY!PO_-L2F!#*#?GQFY*WK<6P-78F4#G6/5D%FF[9PM11J#[UZ!@&&
P9TOVEX5^>)$(+[7"^]29'2YT:J?F6;+C/K4VR>(!/M&Y<BW'(#\,TEPS:.R!.PB&
P+A!SC5O[JIV8,[(;*CAAG%\\I%S9SNAMHYU12QA9/IS@DP)&S<TLE=EEK1@"T,J)
P?9Z0[!V%9-1]LCE8&V*6OAR6V53R/22'<M  #YJ 0(?\MVZ8D@=P0!^.C0]*,:R@
P@D$4:(X&1%'.S=U '/'\#[[47+?@8=2^+LBE$>QM;4HV/"-^ >]QJF0L%H_+"8%]
PWED M:34L;.@KCG:W[5YIQU6P?@H3PTQ-G95F7?P76,9&37"3 \'H]HG2/ W*Y"O
PWF%&K+S4TWF=>C$T0F#;2['M PW."'IV5#+3\^0[99W\):RJ/<A;,:R*DBLOIZ''
P2I-2]^-P/,,4[@,HJ_P^%$TRD([D1O#0MP7/#,YQ'P.P6X@!RA8(Z)V33H[:N-:8
P,VPUV-6C0+'5&'K<V&URE56ZTA3<Y_Y>S4U37OMFW&V1[N)A?8L_&*:3FY5F*FWM
P)\=T0P6J?0'\(U\VPB,B*?V8&9D!J:R1D0',N_3/J(> 0G7,=@=KA=^J/$-Q13ML
P[-U#R7AC,75V$-NFM2YAN07+>&$0.9CDVF/==7+_-:0:FGAH?+.="#^ I,XAXQ"0
P!\+;_2OU>)%3%A%QKT,+ZEV/(?Y]2EV_#^"P@U!J^L^F0.U,.4@V(Q++4U_(ND3S
P3V<Y>L'J**6F?9#A:).3M<H2VAP=P,JK5*=.+?5H#T#O'?CLT83Q85/)1^4?DMY>
P;99JIMGU*O36C652YBZW%V4-\MZLL5-#1>)'W)7.4U;/W#/3!ZKZUOYAEF5K:ZED
PGC_20+,X]FU""8_:EXVYJ8P5^0U&K.+.4?MM>X*=1033N; '2DH]0].9R,7GQ32Z
P\IRA7%HT[+04,/V-SX$N'!,$B0[_Q@ZDDD<8/\G>C823B8 &KD?<9:=&6X+^3!H7
PE>"%!?E56@:T"-@ P^( #%6S3K/E[Y5:BD,!"-<0LJB,TGI-G!F7C@0:D5(:GV:1
P^?.HX+&-$0@A-N?+OJ]!WQ>U&#-[8N=O&PV XOJ>*!*#@ ULX3 #23,H)=2R7QWL
P"O?;L(1'D$Q?);W%+N%%@I&Y/RCLO55AAN3??B(]>*;!DT?[A$M6+*J3X,;:$""-
P,N-,XCV*$RQ%?SOW\N...=-L\=%O-7KT-LK=PZ]+47@7)Z\/(8UC[.:O?+C7!Z_>
PDY\OJB[IO+=E+$X)87QBH$Z"D$I\:/HA6:/[Z6I5LQ^K)R/^N!..^"Y*$J%+;ZQ:
P-GE$S'??:T8;4Q[D(A!5&O. ]3 U,%BL;\F'G]9,'F;-+FCBYF1,%H3.4?^%OM']
PI&E:EY>Q1^]/]M:]W9&]H4LDQ"@J/Y%>_=^ FN>..-K1.S-N0U*:PJ"-$!)9R"<0
PZ57QIK0[VC)7#%JJ,+:V]78SNJTP.,@LY&*!\E?95R81^5O^<'& OON"90\*J+L\
P4.(,ZX#P13K=!]AXJJG_W]>F36M()_G:V[ &UF6F$P#\B"LPI 2<&5(Y=ZLN<[G0
P\(]\Q!:+NTZJJ'SEYIH!RG.EJ&AH^?Q?M08"/M2TJ+:PJLNNS%%!GJ^EQ,XF9?-1
P/1 1ZSO[J.(:R\UME]LE,5(V;;V+W_5T]'1J/=X3+'59/I7N"DQG&H69[CXV+B3*
P=R@Q7AZ2#%MXA&Z,%&L(-I9'+%R^/\7Z'89Y>2$BZWFD$?IM51^^MJWM\?8))-[/
PHH4<H^>((\@,MC=&"4^=Z,1Z]!2L(:RB5<YV&ZV,H;#)&J7O$H^5A)3N4*%V"O)/
PFW!68(=T2E&<\EKG!-%E:ZWF3K2_AMHCWZV!M#0H61)=&].S&+F<K)-0Q)[W2D4M
P($^Z2 P>'Y!GO<8Y:6*U7VSY?7OWWUS4:KT&-'0]O'[:,-,:G *#;M,_ANE+_BJ.
P9VBERZT&-$EC*&19%/:M#4D1_*$"^AQ7$;E0@>:O^DX8N$SV'?R3+'W8SY2>T&!+
PN=&:"8LV8-SC)K:PM1OWF4X&E<>_3NC/"EIFDURYBCQ(V,AU^*BNP6)YC&F!;])B
P<7H_,\+F$.X83GOU.<"TB^M6DWM-]J/T%(D\V5E;,4&&<HI_-]!'5S.O%,#26&(&
P9:L:C:&TY9.0F0ZFZ!":4;Q/<@5\AS/Q @U&,I;7)7#Y:1U 9&_<W(Z"WLI"5:..
PX8QPF_[R^O)1]:R)I38)NPW]YS$(@O,TU=/+Z11,E.EU+3#?$",#RB1/P0+7 1*E
P)H_>!))IV4]/7M)IY1DZ)KVAIK*ZCC[5I\1G;"5L6\WNW[Z&SYFL5U0M&@>)$N<1
P@<+.62QJ<948,1$QVM14[6WGNO&J@]0\K;I@V.)E&$S67]&"B8UQ;7]A9C@C:=4L
PPH$(6P3CF)Y5@-+4^RJU^VT=*ZJY71:L29*<[A:RW2-\9O=M[N"SA5E/L#AW,Q6^
PSX&90N%P#5.56V-J-XN/?3 ]ITU8:$[:-;2@$FP\7!511/K#9[O5*>;0O7J+4[;5
PS^2S?F=%%LO:X,9Y27J VO_H)C^JCZQY5\ZD;).P^J-NPR,Z$Z]J-]N^ OXQ%L8]
P)VF>MQXFF8:A;)\J)5714 UDDQQ' A9*<08&JHQ6F&3'&[<> R)D$YB3\]=(S]VQ
P^IXCG8>_ELX@Q58?QU ?$#8ID%M0%)2NWZ?6/(W1+W)(%H)O=IE94YJ QU[.&S5?
P*Q -=<[8!-B=;M/=Q&PFM,5Q+W7 IXJFR_%3)DPZL)=(EQ46ESB719I8"LSR"^])
PM9KC*AS!SLTD*0\'O(8\5S'-BQY198>LR-O&0(*GL99;(#IO5LIG="Q7^.%01J9O
P)+;7/U':FUPBR7CRQMY<5D9@@)B:9UTAV>^M*ZA3^Y78ZYMP/V:_;I%A<TW+/Y:E
PO82'1>P@A<RZ6,'(8( ;[(-O^_^SK>47J?!NC[;!EAF?F,TTVH+(08!FKR;:[+:Y
PNS>G[X-Q3EZO[W?B\2FC'1,?$RE$7CM5,5_EKK2Q\?*].RH*!^C4#P70F%@2++#[
P2/DN#ZM)!1V5,5 .F]9VN]B2=\]LY?QLP=&75,8@W]P>:1UUV2=/$";)P&1\1VUV
PM8BF5&,XM;^W#+HC?LEEYAWS.%BA!#5:[I0.,)6U?6^AQT&S52#VS?$,[.-MN&*C
P<H[Z IKL]#@&H.])$U&:MA,M?#/UG:]'56PC,W5N_BCE 4&'N_/]OQCJD#'PVS8 
P2GH"Z_V?P*UZ79=KKW;^&!3X-[/]X*@OUDRV:<X757%<^JO?EF%H48'=GE=!L\OW
PLX3_YK.0)I"=ATWR3CJ"]P2L" PA/4Q)#MMAKFJ7WG7UN03K6?_F4-/ !@R9=;#*
P<;NL+;K(^L0K/V9>/]&#@,;P_:'T)K7%=/Q9)J=N)R82[/]D%17/1A$7,!G2#]=B
P&<@& H@2],INK%?IK0Z*-^"8K2CW;']U 3!F\Y8/N9IQTY0D8*2K)*?T:J?-O";V
P=GXAF+M8\*$9_JI"W[2'299+5.<-?B75<ESDO^VE-XUJ7MRO<,T?X A07P],'M;I
PC7M'P%TG0LK30GW41%/2JP;-Y#J9\*1:PY3]DV%_$@%HL(_6337-CE,EJ_CT_\XV
PS]^!;O9A59>K%:[_M5Z62X;>U[^E(OW,$=R$ZQWH7,6W%\\<G#%6<+R$_VCP<:)!
P4;B![%4B%JI>]30D:<XAFC?854QDKM\>,Q4%Y$O9 Z]/VGMHP2EW\>>Q-K:;)@_>
P[]H"U@3"<^,H&\$A!ICWC,VDSHC!X-U\\-B5JDC4,1&=!M=0#/$/1IS\-THU\&3G
P74(9QHRIDN/+844X51GQN UQQU)A[$]CXU^$]*%MH#8\1BV?(BH$=A7([49.5E0P
PC)O>=J;^XH6,S[NK8-#L//I/;:BV&N$<G2PFAAC8U1P&=R"1XC"2. S0POD>'"[(
PM$K&X:NSV1!UCE$&R%>0ZGOC#OUB=-)>;-;&4]7/MFKI;1-#%JBQ_# D<7<,R]A2
P14!@9?DAUS.U7])G#?;\V66%(3Z5#TRTK;6S\\YP:H[XG/\H.!>9B#!G%J[^3BL4
P%9,87!S!Y:"@_>'H=W"J=6;T=[5V9?.6,1(Y?EP-S50#SV5E0IE>BN_ZAI3OK8-F
`endprotected128

////////////////////////////////////////////////////////////////////////////////////////////////////////////


`protected128
PDU7H_H3X>>IRR,/N?KT7T<0-(GPPGNX7S)K2O6232&=Z/G(,-RG>ZRZJA ?<O-9I
P'(PYU"C>U0.Q;%B>WC6/4N("!WQ+#Y2,0-MG8.LG+%3 /LU2A(GVO&>"+HS]GSYU
PQBQ0J.4BUO$"=7+"Y-!-./AL(=;MC=CZ\EHSB_^R&MYK@&;T*&1C]-S2'Q_VHYMQ
P&G#!0S4:^W\1^9*>:P<(K; %> :Z>+IDM/0\1:EJ!@VEO6DSZ(C!_DK<GVSIO*+Z
P5A=;8*#"YB1M%AH*?=7FM;S)QQL\S4C69IC=EDKO=O>7C3)EF9M:$RV]UQ<#X*MR
P0O=^PF3;4&1YW)FVZT04%$(A. R5E_PL"$OW*"LX+#^])S>#+1& 4'#YG#^&OMD"
PMYZ0E[?N%#*?*D/GI9\/*Q[)40C=$[Y[EA@G3Q<5/^V:&GS#3_A&^1X@UY[/D^;9
PW1=NI/-E+5:JM@,,]:D\,C,H9(Y"PGH^[LOPO$?9I8\MSR[VH%&'.3%WB+VHFYC0
P]]* <O,Q8/^E<6)SZ!O^%B[3(IJRY?Q$GI*YW%,R2<26X*46^.S937_-,\&C->;!
PM$]=):):+Q/B()0NOZ +-1!<_E3)X[0E^[$'W,N+NM+UF$Y$Q2A._[CXZE_19]2_
PI3IN["8!%GX7F?(4MQ<;.PD>H[0DH -B%%'U5/O6!_N+:)7[I%!G/R:3&JSU\ &6
PCO+A(-)\<':VFBCQFX^MN9HI('L'[S)@F'[J8O,#!('6$7-(G1U#&I7]]<>FM-/-
P%O9;67=53JJ:F$TBY_0B;EZ7TM=SMZX%?2LKY2!#[(%1O'T]4]YN2IP_#E9]*,1D
P--,&E3<_-/$^=%>^X"C.$[*D%L@GT,\FI#:*)R&Q %. ,RK;!J$V++A%E;#"T;[9
P.S#&+TQ0KTG.FCMV;>H<(DW3L'.D-.ZN#&BDR"$"KW1V]()Q@ \30-E\[%=VP5TH
PA.-L,A!6Z*OZR<Y_W"(3 X+7YIU#NKI+84S<#^-F_1:?5LM2HB0_<8HM/P*$[5CH
P[IH53VVL)EO#)6V+D>'#LS@I;#:1RWC].'5ARS[B3V ;>$8#L[N(K017GA6";JR5
PD ;$R.XTZYOQGAAG;K]-LD'DR4>*B4UMK\J!7R,T,\>^(:'4> +;ZIVDVU7Z"0 ,
PE?.H/$J<6%2"AU\,S-P9(;DB,\E;\-V.-_(6#)#2ZZH(;6"*KY6]":QTZ/L=-Z\\
PTGC2G8(4"2F4:4P/5M,:2GKY[WH6%,WNYOQ!E2R[_,5DT 7AU*1,5<(SD)SP'__\
P$_EAXB.Y%@378.$RC?&'3[NJWN -G7W'5]^AYM!QJ)51(4@%Y8'E?,])VE? 1(+U
PDGJ;GG/+V,--X3;W"BOU%JI7TUA_8WI91PR:\!'$;M/T5_*6GNUT\= 6[6W@=C*S
P4K?E1ZDL9J;IDC;6&5GWFZGUBJV2?-TZYE%A]D(%J0D027.UUUFJ6,<&3O7Q8AV!
PGHI]J^$[87AR]-.T"NF.>?HMAY P2F1,ZFCY5 H[X%3Z;R4*B^TO#)B6FF'WEYRH
P+OX@!0+NK$S%[F_72B0+ !6/T<B'1D/:%DN;(Z;3R )ILX&!#I;PI7I2^PYDQCK2
P:\]F\?2ECM6WP^]T[>+-(B$>EI.$SA9+/N' )*8YP6_FG>@.A?9A*L",@*?(@J-Y
P+> JC#K1[*2SIQ _#7 [J]KV'?!+@.DY9?5YDSDG5\(IDG6)RW*??3JU>J^ I0/E
P[^Q3;5U2-+6?K+\F'^X!QEE=\I)D0A.L)B,HB3[J,<#<J" @@P!;;\2(-<=& XFZ
PP*' .OM1ZV3/9C7.PN%VR+-?'8EQ5/DHW&NYV#\$67KNR[W.NGZSTZ.+N42AXU0R
POZ5RNCCSZ,A&;H!_.UCC'+-"JCMZWLWIX'[K>S0^[<JTUI^OX/I0)/I/:S5*[(/N
P^4J+\MKS$L0A_RPWR=ZE:W<5!<AVKOUSA6WW=AV)F-4_/OHU(0<$8J9=4)L)S] 5
P>K,)T018T/Z-@DJ!]!L?PYJE1$$4;F45K9)5W(B#_;^!"2*GKK8?L@_Y1CSQ@@=3
PJ/"85/BP+MVH&C:_#E5>CUHD$=(F"K,103)HR^0PVJ)E>9>UX]# :&@7&L;8/<>Y
PO@3F/*!1QYL,W&V\SBBM<+-:A#_BW%!?J.#^VXGS4+V^A<!U/B1<$L-R[&.Z "<+
PB%T]2^/.$/2I6KRQ*1)[OA9OUUOX9%&L];&=]O(#SXQ\Z-)JS">HRN[_CIT78I(=
P#=UQNLI,=)6REXN38RE)U*'%'DKB9CPK<UN @' !+Y4/.S,)L.P)9E<F?JO/3D"+
PX@QK:Z4H%8@@[H^%U0E/VOML&Q9>SIBRVU9)-'L!3F3\LNX:2T,UI3#O*=*Q.F1P
P3(XZ*.UR1-S)(()]^3CU\3@JM]A+I@DQH].L?LK/WLP3-]@'?G!C+E?FM-!:I&N+
PXP=M2ZY4O3!M!Y969:CH!1/^[R7)ZI!X^Y=@<?$0Q';NC7\2"P@QS% 5(@\*D0."
P7Q+G("U9>$P_! ]59E'4;ZQ1=#MEYK44=@4$V</)G&V5D3[P ;6Y\!'=31[RJ >(
PP;V;FC%]1F1"E?[^"4;N6/5ECK#T<-^-O\ZHLA(E,-.^Z]=#84\"]#M;I!"?A"&:
PA7#X46JH^#>UGMJOL>^'_Q+:D% *XQ[,>95'S<B)@SZQ=$UFQUQMDGPN$PK:M_$4
PP)Y-6+^K$GS:?5YER0[/?R_<!-(SYE&WSAXO*64N0>W%09KW2YJ"7\>4.M(JR#HR
P<3D\!U:&EF(B"+ R+N^WK8<JBL,#-P9BU)O?1[I,O.P/+*-@Y W'^D&R_@36YMT 
P 'MNA-[X^TX^^=\Z%5R^72(*72F"&GJN)ZXV\+M8!D>JI:E3M7."RK9$T5*E8R&*
PT@DPPM2I*F%SRR^?2U$KU5WICA?L<I6F"KJ[CG\8E@%10Y_3.$S&G_XT&K)<<EFX
PN#[$^BV--LU2ZH::3X-R-?:-BG-K. 7ZQUS*Z4(2 :=&RT"5>)?8ZNHL=^@BSRA5
PG/ \L'Q]OI*!A[]#W1O1]<$?5!E>[ D<=4(NEUOX7B\A,G$^B>Q'DBB,\8.87N=E
PN&0,H+ +X>I('!!B%\KS&R>./$Q:!HQ5>V#T705[BZ^8IZN+/=4:Z;P(Z^B)37H(
P!2GGL6#^.9'!BAUWUI<I3,;FHG%PG+PBZ;/(GCN>:MN !H0F!GEP:U72X\.H5NZ&
P/:$OHC0*GHBS52V"X\%YO8&Z4LX2-K2>QUVE DNQ^-3(79X0R_O>Y_(U-"-B!I&?
P=S?-2H@,7> (5-W'\P@[-9,@) KOK(!@EQGH;UT\W5JU'H#&JWV^M[NN^(U#?>CA
PD63C0F!9Y9.J5$:64R5E6G5'S6[^(CPZ![8EY\_+11< WQCP T;94+&RLAM"6HX!
P.S6#NU_T5AZ1[8M K?*B9QV=N\,QBQP"^[NV$F%=_RT" ZL)%:R-G98#7 X+,/YQ
PBY.D,B>%I"D0^P8,W!"*\2]PNI=;4"]^@7]79S3F)A?!36/( V %V'5F[4)9-DN<
P>4=<<T[TGK<1[$V'4!;:^\6?]0Q%DMDF&\&E@W#Y!RDMWDN'%!:[%P]=BB7WTELR
P.DE?7KF*35<?B;BGL7T>+NO;3*LBZ+8ZI(PF @VR'=OS"7YU*0#>(G&!D#3QN3SM
P[&Z'@K*8_I;>+JZ64]@I(*[%0:L]JP36S4XA0-=1>]G-S=M?95./'0C08&[N!,;H
P<I83& KV9<*9 Q##6UJ8M<B_;F$)X^>[M8A.L"6<.VT'H33L1'#GV%B^,SMOA[L%
P[1-H,\1=80(N442*,C-P$R<S[Y63/#FDU5E=ISEY.7._/;(6R\1[61" \B'(09E]
P61NFEZA"T,5Y^0KSIN>:ND8#*HX0_:LN>@>$98=?IYC#ZH'CW\=XU=$-M&1<P"M;
P<T>%ZI(;"E5? E<5RNX-6N@,S=-OI4+]FG-OZ"/<YG-,1*F#<<[L=LI)/$1>H7U;
P@00 A$)2Q=5].,9L%[Q!)_=,:_1&$:D0C8-<@N)]2&JD_E'J97WT62K/O=3?C^8:
P@YVHGC[500,UNEZ_B?5*V*"= _?R,%EZ1ZM09/M>QJ__$Z^GZT18+P2F!$J%1J(:
P/&-ZWXPJM:U1N3) VB%O1E?-R=">QQ+'=\PZ&"A(Y6"X;_PJ!RH=77/AVT"_-<ZF
P+:\_FY2*F1YL9P'IWM5RX.C>Z3>+)ZPOS_9$O@&/F)_\/I X1<A@8[E4G9,>P4$+
PUOX_T<Q_>(MF"\J6-M_D^=,JW8'-K]EJ.Z "8%B6:2/60LR0RRTN\L5XYK-)C7%,
P6= & YQP*$"_/<XP1ADZ%O&-.^3MVGUK?'974KK;<:M&B!J8*^/+1IG;MD8F1OK>
PC/$8U4Y93UT)J$,/^&:K9R+J/SD%M:B:U'DN'6OQ@O=O"QU;SZN6FAW7T8"MK#PN
P188WK@YZ5&Z832ZL?8??N]X&3@UXR^B_/N>;^8W9.<V)IU\*Y^LF&GA=K,#+6%95
P95RL=0OPHL'>3]\*T7*8J2->TAUJ)J]/1TD;9'FYS/<\KPX)>6'L>61D4&5XS&+%
PPN@].*1Y0+ XGW[A&S8+,=SMA)IL?B1C]J$[C[/.(RXZ[@%!"7X.1HD8>IUL=P=9
P-XFD@0(ME#$-DVR%0&'3'D>DIL! <TNMJ6=R;/U7^S'? P?>0@E1;$,_!*5=K=H@
P$-YMDYAHV<]Z-@R[X]^<N1&$U4$7'H4WA+FOC!V:$.BSYAHQBU.?<G7@T[GI2M[2
PA^1B";"  IJ60GC$"]W:?$+KVN/0P7]8%_*8;2INS//HM)L%I'N.W?)3\0@VPA-+
P!4 .+X)(.0T@N ZANHL8/2LSHHM>WPO<\!;7^;LIA+W!J2[9[&,_MJYRF$L<FP,R
P"=#30DO.-QWNF*ISV9&CZOEX!W)PQ)93WO)Q[ZR7>#,DE+Q]BC#\1&S?W3Q6$,D9
PPA7E;' ,7@T*-&[#J)RKF2V?D^?<%DH-$K@+<:Y.&*O%:?I-M]I])MG1@!:"6/S7
P<5K!9!,W43)>D>#^<XS7'V$JTO</+>>+HL (0V'*%K',7I]>;F(T!@PEF\P$0*H6
PME,5HYXIC"/5PP[Y< ;8;5'<J/+ABU'_NQ5V+0@L#]C%857^Y#Z+M H:*:9$(3D1
PS1]@?' F@%KUU)E0&MM5:<LNBB"+W4(XO=4*.#)UNW<>Q>WP7!M!0S;?=X,V;+8 
PMR5QU]\8(Z>LO&YP%ZEL^T09+Z\68C.D3&&.D'MAL2X/]+?Z#D"Y^0;'N-TMN[5N
PW08B.@1H(E.)ZKICF^->=S*@<K R5M<SP2I5C.)02*S&M%M'EQ=*[:'N4"!=C[1U
PI6A7N7\?+QG57C@1Z/R'=:!$G3XV&QNF"^?_WO=A?,!48D-1P31/\9@$%>5XC3;%
P66Z[S(Z9..LZ*1M,##2YMSRVHN;^-D&QGE>8@KP9U3S\;SI6Z-IQ[2_.[X077PS.
P,'N]VYD7I/:R52VW/S2_&(Z.>'B$+S.%9ZZKQ+I<*]<-2OK^SH '^C6,JB;10V7A
PDQ\3#"WU*:*F6PSO5&A2R,UX8=LJ@L>1@%C[N.) RVSQ.@_-\+_G<3-[)<N(_H!*
P[^<8F/MF.Z?Y4$'6C+1UK%F!^D]\JN<.Z-/,)S0S\\F4*[RF08IYCH8HI\EKD65:
P/:5:[94A#@S7,SI#'45VF<EE\EJPVH,I)W 5Z#HPD23F:,@2?!X%FI?\KRG?6U\-
P#3@9G/\O(?WQ/%^F)T,2Z>UA(_+[.^*WSS:LE6Q\=Y 5+,$6I'A)1V?2E<N-4(]T
P^,9KLDJVG#T+>QM=S4__E$"+GP[T<5> %-.WAEP>ON/MPI9U)&Y1M\:R+3F+%8:U
P2 4WA46I=5!3J:A6("G+*0)=F/:SA24]+L)3^ TX@^VIK^'$)->KH1ES>(F1QC _
P4SSJFK^4*3+<D<H:.N6Z,_M+<^;47_X C32Y02N[4-PVY\V9J"X+$/0I/_OXR_O;
PGIA]<;IT]V8<ULX[3R:1\-X!5CBDLQDN^CL]9AO]<Z+T&*!G=)Q]$[P5"4Q'=A@-
PJOV[6;OHI&(XWU172A5P* 7I)JU%V<#P=0>^102>EIZ=U5VT+&%(RYYG[D]:!M2+
P$%*O?+0X/8I^L=NP=%#T.U5E@%W$O]\K:KAL>'M*V^!DY(G'$W^N#<;N35 IIDDE
PEP9S!C%:Y,R5HHX3V>8[:KHDM=]!O$@\?@,078H=018=/O5A)([?%_C5!5O$!KT!
PN^/QS.HTNN,6']D=SJ?4K86CJ/6D#F"&=&_1;80V!QYNJ5W3F*GTVLN4&I./-43!
P7BIB5O*?XF7]#1P#M$8\5<6C^G%TS\U9>*8;4V9^#S3?;$\1CW02<)J.QC15()JZ
P7L#%/#@&2F:,+V0\O'B1B.X=DZW+;Q)R35@;TC?U'DEOUDV)IR[DJNX'<MAW F?8
P\:H+(A@A?W5&(=I&%P8+-JU0.V9WD&L[1G:(Y %Z$$I!:**@[(+)KGU>W9I_DR'X
P\W/^528?I7.*:></3$;G['V^/PSYD6H ,#&D+W_AZ)>C?;^T6 [)?%4769NT"Y)_
P\P!E7.-+SUD5 T->+P*8[A9$\&[]N1_HGZC$!A.R.N5%B!@G2')KTEX1B6LQW&@4
P58,Y<&@(9J=%,\.[=YH:)C0J/>_'E%X(NI4*\ZLF)[=_2C/WGT25)87?@55/V8G!
P!O>]H$%_*089-3Q<ZQ"D;Y,R!:_C$>#V7>-JX\F-M@&83"I2IX_W:#%9F-:?,VAS
PWR=?QC+"NU4:C#XCLTXF>8Z:U;8R"L^+QH83JE\B2I*+B*=KWI%[G4SSG@\]0#J*
PSYTRS&&K9N=>R0,79R&!R95DV>,X7ZDD._@Y*#3=(I,7.,2^X0<9DC:)D%?,6N6\
PY5&SG?DJA!Q@6Z0_M$##C)NO/,Y]]46+E=__*:=+OI!&&V3']9*T6PD5!\G6*H7)
PHER0C "60%<0J]I<S7&-R376,U/% ;,'*MS94B[>%Q0E$?7B+G+#KI@R8?U$.?'Q
P]KJE"SM0T9OUA)L_[Z):3I :%DSLUK*0'-A+BQ&9G01/@\R*<V^L)0IQ>A/F;J9<
PO%F$SGOP=)'5JMQO22_:2S4KK+BSQA.#.Z^KUO@/<Q&+WY?!&"G3.^91!OQ*ZO^W
PLLQAE*[A8)/L_W'Z.9:3( W7<D_)B8)1KE7_W?>J!1Q)1&>PKK4>0MR%C#$54)\5
PU)#QQ'I27EM P_<^"?.+W4(_&0Y_I> W?<8_M$U>6)0B_*BV7*\!R-M91V_D#0,K
PAK?+E\=&3%?GC+DEX):XKFO5JGRR)ZS;R1 ($4'EX<5]6D>Y3]?B^V.UY4I9]+$W
P.$D%1C$T0>42AA2BDX,PJM%RZJ<)J?VVKJ*U8#>A@1[*@&";(T@XZE2.L2\W4X=@
PT6?F\8Q_$#3[,QBYC[)21@*AOYD^G046H%<SD$X8L=014\@)2!0^]D)=,3>J_T*R
P"0A\?$2]W*#=HPB[>$*7WVJ:0,AEG4$4RLM%4H@X?1^6''>G]$;S$#/@5,^,!>@O
P")S0Z620ZUFK4P=KYC5PQ5YD?C :N+(WK#>JA'+CZ^WH5(_WG3E4*0#1]W+;@'C\
PR)G@*#)W+.#+?A(%&UZ)B<NRR!FD81%,RYHV?-(O,JB:7[9^#.6Z\7>)VI&+@\/Y
PC5Q&M[K>H>/1N'V1ZR)?C1**T0&-Z;!7[.N04X(4+!9@$DV!JFKRRH=2 UJ)?[+D
PH[2LA**#U$[2%U)X*P)PQD49(.?ZT/FSS5(U'5@V;&$-13C+B;!*$(?HJD:(YH4$
PY<YQ<.?#!]-OQ(U:PCX/0)=>[<@DP*6FG])I\6S1>&Z_;DA%F71^N]9I=C';UA9X
P;)GCDV R3K' 8WQ#2\GF<0&B<PZV)M(>A^5OR4FRO]UT4X*/Z;_*RA-NJV!(DX@*
P<B*L1Z\B59/;F.WS[!7Y-K&>Y2:CI^14@4>NHI@;X;H:F/5XH53^/"5(V*P/(Q^R
P4[DQ;J-*VWOL//;UKL>%;"JQJ+0BXBB0I:[/J3-_N3AWFVZJA+A'?=YI3=X4W'F(
P7W(J$E\/Z:HRU%#G=I!BB\MS/'.O&\.FED[G&B8(DLMSFA&TNOUL@.$)5P:7[MGZ
PLI?P&1W5*Q_]]  PYM7>F-8(T.%RC[).(T+FN$A!>7M[_!PB;:%(#I]7M!:@K_?"
PXADNQ8.95K2[Y4B^BY5T7B>KI:0WI4M"^EFJM9AT,.Y0WT>$.CC;#Z _>%8EXKS]
PU3]0E:]8EY;)G:PV]_GPUP7XNIJT>?;+)W5\/-JFJ/NA9TD-7L$?2=[H/%Q)?==U
P\@7*) 6*W _?N<FNVLQ8DCA.AF[\!LIBXKP##DQ1/,8*OJCZ7:Y\$!OO9CVB^<5E
P0S)$VL)*'[#',B*ZGO0R7N+,BIW>;4;J*R*2%N7\0&37K@G- @- /9!W&@"]%USR
P6DD,*FYQBK.*!\-@C(@&HG"B2O'")RC1AL=D]&QEV8>+7<<PDDX( 9-7>:%'>?M7
PFR(?&<,0LMV;>9X$;:E)$*LFMU$&>JVLK5HSCN['*F1WD%: ]UA^OMHC#T,72YJN
P2;AL*0DW2*7EQ;"+4M1H5'EN9^+"Q<QI\F=W+H=:D1D(;X7RB@^HU5WVN\6K6W30
P 6)*! 8:L6X)SIV6B=3N4=OO)R*MAAVE1O.W.W_& 2K?<F4:P^AT[FKZJH]@(7-%
P''O\/8ML<7\^B.R]OB?2,DO>?0*?7Z&EFK$;B7![V+7^#Q$P@*E( XKOX=HY<M:O
P1.U=O75'M7>)'9H!]Q4#04#8SS\M<\UHZ]XT"8/X,PM&@F[+4;H.687DA2&K?2XR
P#5_)8"X.2]=K?3UJ?GAYT(PMY.HD$B+E,C )/8RM-PU*<\E>OP>F^,(IG1/]DU\2
P&1UOZ:Y?W-#ZS.] M^57FB>\B,AT/9.YJZOL'B%(L7+I6!&6BT&X;((%XP0Y0H2W
PD0F3GPAN\OTI4J GV& '=PB:^UP(T;,J_$VA^.2AVLNBHV4U#*E%- [@^L(G.;>/
PG0ZK[0A>Y8CX.)(KA.2;'?*?;"X'+]A-9J7;'[YIO/L<N*)(^RB*7PMK&(JHIXP]
P* VDLCG]O>/<A_R?@WV- )&@WXO[%O/0<^CY--EJMP(O9,-Y2V4B8: 2L.7@UE'#
PG#]VMO*83-(LB<JJW?P<;Z*1(LP!KS[ ARU@;.'[FA]8*&B04V2^@LG.=K"F:I*=
P0[-*4+D8ECOX#FQ^R;#'^2_R8CFB;;9'\P&'_?2%B784JLI3R?HHCL>E/WBZ+4)8
PO^P][(A\5V,IN+$'A&!M12^=O#Z4=]BCS'$EE:U#F38:4"@.2G\3HB]-KA2T*Z\?
P7SY /A48YL1\:N8"1 CK>AG,E\%\9IP:V)8DO."ETN0@HYK4.T8M[H$^>7^U\*+F
P1CZ5MV$T#;<W8/)JLA.1Y#C.1N*4I*FM?<T6#!M_8;&ZA>7:U@+EF!53\/,A!K_*
P&;NU/2,D!\N=.IHVXA@S+'B7R#/X,5E#]3VOABWJ.<)L$V7BW]M=<$WG48E&;Y(R
P)-^-+/;=9,L+R4"\7$O)5S71H$ 0EB) =T'O.J08<4Y9W6'*CJF\J1'#J09I-Z#O
PQER**,\(%>)(6K#<?%4G+^O2:A J& (.8'&ES5BV'K /F>\3U:_59]J^$PJ6*3:R
P9'MJHG 81N'!%XT3SPU[W"4#)_:F<U3&FLU^[@(:X??97/4^0-XU/-CYJ\WB+$X1
P304XMBZ/E2=POK_TK%-B(%L&3/%$DJ=1*7S,E7K2HF8[7'I,%1D?JW"&R.Y857H;
P/V08W<<D:A7CNDX2S52UF\\ZDK:FS!(ADCJKLUTO+7;MW@]OA@9NW#:)$LW4#[+-
P\+NJ7]Q#@564 :DCCFY57CIVHRZ9OD0RBCW5YJA3+\F-&L&_8;^PH(6N-6HD4B1\
P0S>L6R(J/L8A&N/7TB>&LD36Z!03ZW0H7E;/N[)AFHVAH*<S55$?D0A/:_*LP)X>
P0NRQ<T<'-5\.:"#Y?2^.8)D-\2C@P>E*?4,[3FZ)DZ6FIXH8#(1;/<OIY$(\!'\G
P]E@4+;YH7/EX4<NY9U*J<JT3E247L[N0#V[H4_Q7YJV&B8B[_+@5?'3>9EG..&)1
P>![QB)G_#B_TX4H;E"HFRH 5^&I[VZAJ9S3#9V@$KJ Q/#-34JT'_9C516G6*4"5
P('/&!>[O?:M\K9L6#BF?'7MN"V %X(!F4,'=8!?^ 4)W:?JDK=)E;O;=6SK &*F'
P\I?5?*"0Q\%-N_'TO?TB1%7CH7FZ,$YOU! )Z''0=J?-B:$=7X*G6IQ(]9L4_I-O
PNS+(AA[E 'K]CO77]1Y]((7"W9.KHEZ8?.8OYTMB1L7]^*EO<B>0!+V>#3'XF(<T
PRE^$VX1RSF=L7$TYT>P=OT)R%:2ZOF[@: W+>,&9UFT':+M[#F9JRZ'G&RI.JF60
PXF]$2#@O"\C&G\HM@$278DE/;LRQELE$(+<N[+N+&NP]##!?6&4>)WAUV70_H6?^
P.G\&O"C(.%=+:!D%IMV1IKT?:;U48/!4/*VQG;]Y]MB$.%EJYM2=7&W&[DF[97UX
PF/6NCY+_TF [T8DH!H%O4"+J;IJ RHXQ,Y0+^7:#6S4O^7#^5+TGCF"DDKE3,-T(
P]#_?K<Q<FTK<&Q\,!L0@@<_PIF<19G&Z)O)@'4-?"LX[9-B(MYU9@9?>PGM)90X=
PRH7G+B31UM[>JUXEI8Y:'Y*/61=J__>T63ZPPRSPJ^]H'IVIM&-'\^8M$KVR&Z9(
P"1YS56R0O!EBB18L2Q. /CHVFS'"26^5]25"^BRS>U0<<5931/E#>HBFI]&=L!O+
P ,*D)S&9T7%I._4U>2*DP*GHY6(B8O?E':M%G?U(>_9PL'R"Q1J%\HTEL)WP;M!B
P-M#T%-],MM?7$UM,LHS,S](1RRGO<J/93_WJ7-?=KWH/I@N-P73!?IO88)"F'%0^
P"M'7?O 2G<('#^B5F:>%70L-@?'N2RB1(49'8=E"G])'E)@-\CNJ&[2JZ!=(25\H
P9H*(\0W#,/$+$W_^&!-:F61O_:SW$DNT_\]R50K$ WG*4+=\EO!\,*KTA]J%-#41
P\C$DR.0'/?A'9!L^8#"^@]V'X[4[_[K_< F'=5!,EA@!]31+SX*NQ:G9ME?F0/Z5
P;334<D?V[BV5=2V"G376?@ZP0?'X;($\?2$.J:L[;*-A''^" 2B[9BQUT(>D#NA<
P@L=/7WEK8)OTG/<^"EW0^Q8TMS41#SJ/.4"XN:6@)@J?W(,?#5NI.<2).(G$\W4J
P6^-24=4Q+>V\:7AC#J2T"%:ERZ%G[&U.Y3&\ZF@L1"SB'[[S\C2[]B4SHU<:,&?F
PYT?'DJE)2QEFTS6F$^L+;*3>IV^G5N!BKQW<L<R5$]0?);YH;\,YW6>0WA<BM8RE
P>4T WRW@V&-$+>$DU,4:PS/U0<&3_IO4 >I;1BWLM-=?')]8.X1,$L4@>W.;4 F\
PA&&M@&G!U,Z)T.,(<OQ^ 49=>BL^O<&=7:E#M_/21S%@0I8BR+NG<\!^H#XLXO'U
P'ND?N,* ZK10)Y28>]QKFQXU_6NXJ*/08!H2B>JN"\V,"'9KUY"V/BVKAWS7NA:U
P94A*:-'2,9@I@^RL:(/[YWD".T5]$7??".2 D)_B:Y6[PB2>L0L^$]ES$+)MA3_ 
P%WDO1WUW%0Z4,G.:3G,=\Q4.\)TFY5%&'3V#ZD\;W#(( BQ8,1@"GL[[VG7?UVI7
P==;HIL%^)#G+#(0'KP&JC+9F=L>X1+]B,VASB>/S,QY;P): ?B72,NGW][L,=BQD
P!28P;=O$2;;7#&"4OE\3//(CO*XL/'!KPXA;>.KPP2%9N80VO1"MX4_* @6P1N:;
P^F#[(C=&1AF!.H3APB032D\NR##I+,__]-W;:+<R9HA(TLHF*T#WPA03?V*B%KQ5
P.#^T'C_T2!F[O]/?NTB.*JO)RWNP0_\^A>#R'[57=3 %NZ@JQF!]B-Y]YBC6%Z3#
P5_%H,V<]+AUS+\P033?H0.@*92 :46-Q6>PL*63]62X\^4F0C_/0*L6,K3'_LGCH
P*8P7=%=!H/XHR)#2&>8>LYH)'1CI8D3C1Y-.*=PCNM7H@D2'(9IP!'A&"PGIC5=(
PHUZ;I7#,2)!\0.V)0!+QF[K.=QS;?@D@%KL\RW9[?'>(7&1VMZS$O8C.R7C]2B67
P(2FW4QZEIY>00$V39H;7'&"\@!*E)M  .I^0=B0WAZ[AFM@5SN)/CW&<@[@[9O)'
PIG+"4Y5=]Q"<$Q4TT'T_6-$@\X_&=QMHB\K;##R^JX^+D,#$K/BX?: ')!J/]Y&7
P.]6AX4=>61R0IN,;[V;_H7!!)8Z\W0M4&+/L4T2)ZKA^.VX5..MR!2*8 D"6B4N0
PG?%3^\5ZF_+&"0J82]9K'%CK_9^YDN005X0"UKX57H*+;1F'B?8I%+$[-+FJALHV
P*Y5H.G=RC"AG1) B2]34T'7;8HWW@Z?R/'AZ;C-'#1,L*B1GOS8W%1]JVV.A=4]R
P,6V;9"T!=,%A*JL_2%@<MIG\E&T#%J!.UL'FH0=XHPF&U=X222A3J[:Q5[6ICK6<
PIQ7107P=]* _,T'RR ,CCG4Y/:9\#5QXG:#')C/&\4]L/:VS''D501E,%8EB;Y2K
P-;BE?^!Z_#_G445@^3I5T3H<..$6(0E8!/,)W#3;VCJ&2H3<6ZVB2;A$6B\393[R
P/QHSIZ+;)QMR?[;D @]E#<_^CC7N[L2L8$9YFJ#E.SY$0YT,#XTBX3W).]YKS=FR
P(V_"BR&&DBI+#=H4KJ:H;2'Z;T^2G;C;BE%^BA+JUPY^-0QS^\T6.<*UBQ<KHPL+
PQG%:TJ<87\DWZ.?[!#)W;R9\@?E6>] %;T.YLLKA44SV;G4__6F,) 0"_B!_*F%E
P>E* (N]<I:V8^T2OD[2"LGVMB&8'0H\%H(](9AF![VAY?_WVWM%C1QZSD^'MY*E@
PY25F%[ 0IK\>\)UV44;#-[0I= _#A!D=.8)'KSK*Z.WAKW$12KDUT+K<YX (O<U'
P2 )D"><V5UV,28NC$'H^+#44)XHWKRFWCNH^(.5>X-7=X'UQ_2Q>V</H8)T5LSF1
P1A<T=;/[71F'MIC78C<9XH"N:/K[JSG)2;MH2NI<>F8$[+[S66!!*\1DC",C[29*
PL"WX#/CA7D55(A:GR#4PE1W-HZBW(0N DGE1[=<R+DZ-"&+LI&D"Q)[E]7L0]:AV
P3RD+@H/7=M=8*!CB^1_YU@+Q+<GZ(+TD?1A>'"@=_-**B&<I1U)[>10PV=##F3JD
P.7;@,-M=J@!9EG+,E6-,,>6NU:5@?%2T GMKKU]_J%#CEE;-DSB)I7:,!IEX9;ZW
P/2AS]LB["1124[YI61,F,+H_?)'.CKB#W9V_K$+&$04D:VZ)F\#X.!08B_02Q^PN
P-58.N&HT?AJ\E*:L)H8+P0(C-B/4M(2/3W+D/;^9 "01B"6G<CV K[F6M19YXDP(
P-7YB&)87O)__2BSP\L(:\!(33-<Y.TW ?UIA,4^&%7CU+M7([^5.8]@.'?+0'T%M
P4?ERUO_ # ),KM;_JYS>T,JX:-W)CXZB^Q.GJM-GH>,8_?X:NK7L^3OEH\K94N'!
PMA9(*-(+#:KB1BZ1(?3YA;2P2["Y,DE_^C?$"A(2QD0^2T&I.\R""?@ME*;+;PS<
PZYWE3=LCE>@!  ?O<,)^B;XOO@O"&B>"&%>K_DN#%,&P4/<;X[T16*O<A=._3M5]
P5B4\@GZV!YLZ44;U"I<"H^AED72_Q!H$ (=^PSJ.XHJSJT-B.6^S[/+"G8MTI[YP
P0S+]2>P89O)9Z!D%#"L"%6@_C]>NU0Z]HXJE8GO )<B*)07GN2VJ"TCI?MOH/D\2
P7_&! U0;P.VAIHB<_@0::\L8WB'N/-Y2W8W9&@D$.8<J?]2\'I.C'H@MS4UD:I\C
P9*:'ZLZ3YUV7?!EF">I@_B:NB=HYV,PQX1IPG&NV6_?J:_;WRU_2>EF,0?=J;;3'
P?,7!,"FMX,RP#JD<BU0(8>,-%O_9E+'X*H%E"@^P-J[Q[#+T=99.QG<,@X:W<P'N
PZQLWWY-4-01)J*HC@-6?DH346CI8/)FV-;[0.O#4M&7XY-AQM,G3%"/JXU4JM0P&
P*'<B3MF%@B*@["K64$*1YJY)T[ ]\"V4_R]M(,SFPU(V3/UDPJ1OD350(2IL!??J
P*H:\N'9<",8M4#1/EJ4DPC#[R4^DE>YC'2 WN!G=S5(ZQ+EBHBWYBA2-@$6[O<]J
PYT#4SX1U3L&'V4"RS+:<Z\:)C$U+"EW^9RW+0UBJ]>SC:[D_7OQ5 ]$2MV.TG)]M
P*%.ZWFA<AK,T(=PUR@XVZ@I$8JUS5D*[O7NA#[[[*-1I>2S*'9M,4\="$5FV6KDV
P%QT6_Y*SI@MQ!8KRFE=785)E)5$]+"B;VIZX>C-.];%= / (HJ0/DJI2DP($?/H!
P*;TAHE I$JM[H^+N9# EW:(B3.?8]9*%3)M]M2QR!U*]H0)H5,X1__$T:K3U>T]^
PG$^O_5^=H[[_0I449L]5EG5#;GUQF%P6=B>^P,AM/IW'! S?,)\WGI,U.''1C#5)
P@@JF;&!:3OC/Z1Q>G3^55LF^OD)$#WY_%7@7BPLP2GCT(A9X-(>LCV:L65T7#@+1
P-?H*W[Z+AZ(P'3&RBR"P0:/M%?AOSK[U_?..FWF;8?01^5,0OV6M2M)VEP-M)!7(
PX# &9P-M$ RY,]MHUA*M0#55!,/T* $?I.C/$Q5?3AHY@_Y@XO?ZM=LFQ'*[T=SC
PJ)%-,>8K.@22[>:K4Z2S-3)%$CO/ZQ$)T=ZMZ=J$W:I.RJ2&3W["T,29;X,V6:HY
P#CI]M,V?P]\?^L'KI.:6)IV85M8H X#YPF^)/^+["*Q$6^O(YCJI1N7K:$NMM[+7
P3<BLB+<,SJ2D!DO27^1+O!6G":CK$/-VW8V8^B D_*'O(8K%S.7.;%I]%.V?&!. 
PBFNDQZY(5@XL VGTMW*8 %PQ98DG$OB"3""<;$:MW54-:^F/43]#Q;R-.^7>'/;K
P<5:II6"0<)ZV?H>&;:I9TAJNC6NHD]?NG2,Z$L(QEX<-!8 YIPJ9DLC*Q$0%E,Z!
P2H1VIJDM%'OO_JD(P,+QAVN9;;>B0KHQL@;&@0X/3V;$Y(6>#AM[2KEP2?D7]C!L
P173;F4&8O(;'T4MUPU1+^LXIM1@LJ?HTT@F-"27B7 .1[&'16>[<@(BK(L=._K7.
P!]/.$,5?I+EV B8LHI@KDK>7;>(#B:,(V"A9\%0>*()/MHXTC@2-22;9-U0V/QU'
PZ1_I2F$EH197ATZ\I-D%C@%B;$$@PVH]G!DJJZBK#DR%?<B'[-L?/0U G)++H"=X
P--W.<NI_>FFNQVNC.=MS]P1UM: ?=(E:#4C)>^ T9'U?4#"0QUA2\/.H/8G-JNJ^
P[*7W,J-W4H1!51#>Q_@3VRZ\@U7 +C%Y<]EX!O%N04(M(P8P:0G6"\N8.<W&&0!<
PR%\+"C:AS"F,H]F^0D ;!& <7): ]H%])-$=O-([8ETC7(I+%&7*CB2P=>;2+8?5
PCN7TRHT:IR6IR7O7$"FIX3?-.!,Q#TIE0;HTI6"4E6?O1%?(NS9\ V<:H)P07=#I
P;Z&^JDT94Y,QKL"DT,FKL_6XW)L>O"XSHEU;69:F,X0 0-+FEZ\GM^[ED;\:"YL2
P(@"=Q_4\2$UJ8W29>92G$E>1Z-$)A+=$K7(5)87P=AW<[]IY2Q&'@]J,+NA%*\3.
P-Y;H879*;DK3_3 0LH="S T#_)+2RE$]ZH_ N5D)%#S7V,?JPF;09>+#X/6>ZY,5
PG+LEJMRRRNVN#/;B=W1GWGW/GA'R=H5[+:O0-#>:"T/=CND]!QD%WCX1S>+8]C7U
P&2WYDND;RGC<.T$4X.YY6R2S21<7H28+BJQA0L:88_I%VQOY#D"RA+-FJBZ;>B,.
P-7.E-\A\<<"O>-FV:>_'ML%C\R+\Y<[C=GCFC*!&-C<>Z_UOJ?E7HQW$=F4./48]
P.G+4,C*4K["PWHD;'*(LJ04UC-V7%T+QU[6$,?M^EB^Z^;,[5H,^MH!>737^-+U.
P9,>OOG$&+T2MJ+:F%;*;%Y"<OMQW]HT3Q(G2KV6Z(TQ\HF\S@.!>B-W7<_Z7!*V[
PT&8^NYG;YG.T!:/Y4ET_M$@#8(L_=\#"CJ!;^Z3<I]/&18W<9ZC\ET]E?T%=B@Z=
PHO\L;7-N+ABSK5#0<#LPRW4@#MUH6^_4E$%,RTD!"XF&9PN^L2/'NXS5_UV4NO7X
P1,1VU0.U- AS647Q,!1[2,-Q%FDY@U28MQ'T%0" 7-1_+W494V_.OPH-]"[V6@^T
P)/HW/L;$&CE9#\X@)"\4)\12<>RO4%33UPNQE,YK*<^M&]N,GSB5T<S]4_8BX%[A
P5ESO*D=PEPE*QKX@SG#7S7'#;E/*\.6Q!4L>1R"?I1UEM&GC#*/<+0PTY1]VU15 
P&3!/A0@^G&,2+Y7AY0PBCLT&D(>\O('!U]*9XR7&M^FY-B1&_A]J"DX:B/(GT".@
P'$"K>M0FJL@-L1GD%)+JL.6*N[TI(,RR,$V'E_+)]:,N.]90MF@Q/CPPVK+C)>VT
P/,D3:I%E5N5;37A =F=O]WS<NU,"X5K;<3\,=2YD)6WD^$R,?<^??G+#Q24E*P<6
P+L?  _OY:.0\$K$+NS\NK$/) J:R2D>9R$'P/I6D/]H,-S^:%QDD?,7'K,&+K?ET
P*E3NFTDTV=@FO0X;C)>:S#"?BZ,??9CGY*LM&>J\@69'\X;N4+"$=04I-D.XN! J
P&'DGNY"0/Y=D:O/V;]2DEA8(&UT"-SCWE^\%WQP$X_(X0[&S0T/5Q2 <14*9"5))
P7&^1N_9]!99]LVX*!PZL@^30(+I-(3]O.T_-)!0K:K$5+\XPD5\L0\!3TD2W44*G
PKE'(=44#_=&RVB#(CCV!S>_X-YG5JXF=VZ2_ .DXXJPSED$DOD?5QV!EGV"'S&<I
P2"B>3D<;YH3:- *C:9#<>+GG:F_#[#GR2"?7MHE8.@7WUK!C%H&H.B2)FQH+I&LE
PBZ]7;QV4 O\PY7M3F"16E3JO$(1:8UPS+<6E)]0K-,L<9^@>SFJ43SUYG(V@+J9-
PC*.+[C>E!L'E .0#^'>.V@#2-8Z@$8IN-<1D38C4S !4;"ZE7N/29TU?#D,^%^KG
P6NFZA. $=.S:#SMQNYZ9<4PBF^ $N%\&Z?AN 6GW,HV@(H(.TOA2UY,TCELLZU:)
P.R\*V7H"^I-UTU[ROP+SJ-YI$<,7N,5E$O.90)Z0)??1BVYAZWKS%7M4",+W$L^7
PUKD+>?$DIEATTT%?23+K(]MGDINP/_!,3@@RM#@9RB^5;!:OYK['EEO(9'-ER2LX
PQ=L_+W;(L [?V:6$+O'ZBX KC+TMDDJB.#>;D+H]0J2G1W5859@N8RS8:1^MM'#W
P "F<D+KZP"@_9M2-/KF94<V_\]7)6)Y!A*T-J0P'6OJ[@C]J"K@B5\1BIQ7IOS'M
PJV=]6LH5IF7\)][4^Y^XMP3%%F=<EI9TVT!ACEEE6MVU6$#!K2"78)[U$(J_2OZD
P"?B;)]TIQ8NBH5!L>S%Q9%A:3$J1P0K5I.\54^;L 8/U]@K<U#/"< $F)+6%4"?B
P &(VD7#.FBF,.(>=W@:O+41*3<M!8 1H!;ON$A@8(AE%YF%0VZ!^)43QOQ;X-=/'
PW<$ Q&?%H6V(6=/6LDRK&OI?*&EO8E!O/+O+_3:-P3@,YO!UJ4O-*DOT8&98PD@O
P7^2Y@Q4)JH3*TN_GCQD;*4NAL+\R&;G'O%-(97SASU-!]E=7[NT!XPZTR)]X[TQ!
PE.1T8HSX7/A47<Q9%8.=[=81I5>+Q5625C(AB!(4)ZN[=%V#"O@MHO!*N[%OO!8-
P>[>YYVVATL/RTOL %NOQIT&5-? 5[G!C8VO^!7AV<D?.D5I8<%(T1_OOV^22(N3#
P*20(0]BO9W5\-<MB?2O%YX?LN9_P H%##^%% [O+*3]?,(/+@S8N0;I*4^<2(A1[
P/%<T$=)+<?<M-(W"D$F^8#K*C$(AECRVF28N_Y="CX0B,<J/ZF:#DU.MM&>6FB>Y
PGT+FIB='LPC0@<I(8FIA24<ZK)@7Z\Z3.5^,\=9J46%MAM^LXQV4A>].?=-):(7%
PDE(LR=))VCFG4ZF^_NIK =LC<[##=;1N2B<[6Y?>U@@_2QBB"&#FM#F1X; +G@)E
PW^70ZR!-$CCU&10;E*#71WEGFY'S;[GH1+A%'B_0M]7(#DDX);K(_0(P1SA46,4V
P<G4!+*B%1&^>_EK]+H](/I4ZUCP&9X]C.@M#25%5IW:719$S#$LZ#IAK'DG<K<M:
PR_\*[>SFOZLDG5Y@"P#$V-Z.<]Q-96_J:H<U[,M@FT8 9:!BJ'ET CG?-;P^;M!8
P&C_7U#CFCP&W6L'-4D=ZASP_EWH1@G+$&V-_%WH=7"%V^?^A.0N#: PI7;PE\Y]2
P.2GOM(*"B>(2E"CJ1_#U\F9=-^Y96I/J"W3"((.9&@5V=)%=XN"%6TX9-'Y,3'UE
PGVQ)SI(8 8U,NNSS#"VL4X!L,88=,!=CF1;/\VF@S0G5A72AONT4Q<H38T+B1F.#
P7@D*9U37TP_%?P.]UHIONWHZMSBNSOE''TQ!,O2@C&22KZ^NK]XEV4,Y\5&X[\W(
P8)8H"X$[D!/*O1)69,"PZ3V]F:7M_3B+MX3E*W-%.CEX6?I/C[!:[V;MHIX9\*>/
P3 3NEC.(SD4B&ZG@ ?AL7%'!G\] J^B:/1YJU(A@CS#OZB-:PT2N$MR]?HA@I6+J
PROYMY-A\O*;7AU%HIJ:5_6*;&")HL&O'/EK_L)^Y?A*P)*=J$5,B]2_?0".R7U@"
P(+<;WDD.1\=--\(#;GE[>MS?,-94D*E]Z56,\56?<IM!) ^U+F1*J!U5 ?],S/3(
P5>>F($W&/D-6,=FU6RJ1(4H<"3K#@B45P<-UJ'(-G0?__?0/;+=F='!"@-'5:[,B
PPAC/J,9I?OPE'7@AM!IN+W^;*V'U_B:OA^;=CRR'+W=5ZDR/Z;#;3"7S\P';R]V>
PEF?7R]LR=B?U2QYG]E^L/D^S((E$<_-WP/NARRCYTY&I84*K]0KV] U$@V"/'=MZ
P-/)NJ/0))Z*Q!'W"18E6G8433VI?4 ?LP2X^='3DH7&6.1TOQY0197>8[AI)Q@:C
PMKY0/T(&#TOR1H+4W8V<RP?1_G$F(XB*K()2&C]SHJ?I\N\6O7__S+'5)\(*.JEQ
P),J=HCG1-R!?XS8Z(I@6%W7F1N! 2LQ3*H4G.4R$ZN<4@^\^)A 'K=OU[\B)AH/V
PZ^]\@-'1:F3ZP7B+49[7W24)/+61@05UTHLD7([EO!/P;4S*U!^((0=X[4[+K"=T
P%F!TD'TV8TS,%E@J%P!3P*++GOS#U*J+C/)Q80F$D*%4 *&U);7&Y\3>*-F& B6 
P$?/H'YUUZ_3M1MX8+B3>BW+78L]/("5-ECYN_R0AT?19]R)NME'^*6K?!7U#3S\=
PI(+R+XR"XG9 3\.\%\ ,I+H97JU>[A"EC_DL^WS&.$N&.]^R<8T'-/G" 1;&@@J_
PALY+,V>6SW\J4_1S621:IZ_,S]92X\K2KV&%81Q@.0>:H+D?VHCXAT)J=2MVOCQD
P+6^]%3T(7=7*Q$.K1+\).CEE)0#"!6XTT;&:9JHI36['<L[.0S02 /R8I0(L=?WH
P#4J>9*5H^'8?->:21W4/?,"9BW>M'=*P&3!2;6MU\E'J:\M8P<,&W.E5./,:8Z5:
P',XHRV6.Z'HD?WCM[(I0(QCB14BW0PP+&#8"L1Z*W)67QY';X0\*)H^Y1!Y(=+FC
PI *@+W6U2UY _*.0B<%%M\TO4$=]53_:4"I^%DMJ_Z8%VB^?]#G&O YK.SR''?[?
P8 $@_-GU[W8G0T5O8=$FP5=.4.78\VT=ANMRE\5H8L]O'7H)P4@CU29J"TP?5$*C
P\$+JR]<H0=!7[[OO:.JVQ+RG<V 'TIJ/!G(5PZTQ^?EAG4TG0?S1B+SU0+6[3$I$
PE(J:<?]5S/O5YQ!/\(!1)ZP\WPA_J(,G^UT/TN<56+3]+9\19Z:6>@!1[(F<T;_X
P241NL. M4:SEYY@G@\4G[9Y+84C3>+=<V_3X8'A3?178>S-5=#V"<36\6S#*YYVZ
P3X. SD#[OUI3 /:R%P09&O9CNK]&4*@U1;]*_6@;I$]<VO):F"#[T><@B+>D)LT,
PB%TUCF$Y:J=VS@=DL8@\42QL.8&FH\B@(ZFBY%0D'&C_+XO7C9\5ENAOK.*-082Z
P4K_?".</>P$0]FVBZ@F_-!:$M?XG"V[@?,O]@&I)JM:>Z9 (FY\=#7.Y29PD3_:*
P+/#IQ5A80KHH-%25+C=1:'^H-'(T\B1DV/)V@WGQ$SO)Y<5O.<-H;._"K' \P.!R
P<&(U3#2"V3L 5WJ!@ZARH789\_,#U3BW2FMD;J-1LU_8;9ZLBC,E;9V5PJ!5?&XZ
P%+*UR3HM[IE[L@KQ_>S7 YF0R%W)"UUEULLZV+.^"D+5E8NJ3-MDH !/<#,#BUAQ
P[F2:F_EZTMQ,7_J;D2@4O [EYRT F1$XRRR7QY-&>)_,%2*G@8!*,AYOOYP8.BW5
P=#*G/EB-Y6H$%WKVC1&O=0O^)I??.($8Y.SB=;J-Y9.<%+97-I0^0EM::S:HU.=W
P1 !5>T!=[U[]*';Q.Z>:&6B])?D6B&7_67?9>.12\*'T^_>&PP'H*SX6;ZF[YU22
P4:L;R$F9I-7A&;]LJ%ZL@^&2H)%$1&W(05&#\^"H6!66K/X&XMIZL']&[E=9"U$>
P3&W;=[JK4P!ZCM<=DXBXALXX<3XE$IN"/6Y$ES"POD.=RQ^*;^!WD2/RKO*A^L!%
PN4-=#<UM3;Y2V_)1!G4&]ETH;W.M2X4ZO?E_JS,]/(&>#IT9H4&CWS_!J"\'X!69
P5G27P 8PDJM_='CFB*CZU(>@*/Q2 1$((ZR%GB@;F195:%7!S<<B3[&3F.(N7#9Q
P@LB">$8!'76^N:$^5L^GXL@7;F3R.L3BDI&7FULF^- <QCDQF'I\E,;\%1=)G+5T
P6M62$V .KLA/"-*%D$#=NX Q;.V.+JU8BCZ LS@".B5RHK$$JXZ&,)5[*KU"V>7Q
P<;K^#M8E/QE0;EK 0QC!6^X;8%/$B9ZB>7Q'/S6(A&0+:P4,FG%F"BZ#&-6,!T1L
PH,F#'>IC-2[TY#0S+J\-J._LTC!B1/+%3E+E !-S6OQCT9P'58#$*$"CWG*,;O/N
P@P(<>^,P6:19G>$GGXI$O5I 0> Y^+0^%9AX'!3#-N8HQJ#)W$>"M('.$%#@ME %
P$=%YZ@5.$#)A;_*69HHNO>7.-27<"Y',E?".5_E5>:H8VE''-,%Q_,T+G[![8=AA
P9XSH?#6 6C3V>TOS0<W_MA$1Q7(!P\CDHOW$9Q(0/FECR%#0#TZ=C+:[0$-!KOEQ
PD+:%Z!3C[B?2NU /=AYC)PI-I1S*_9953%*&QA4;OWI%W27']Q5)>T]R<E;P,543
P+^'IQLB?]V@[_?PP"M BV9%H%3#'>8JV]Q"U#Y;[/C))E\G3T#+>"#DY;3V7SK^E
PMWAQGDO\3%(TM'@UN/+KC:7!&">,CAA0^,NQ($EF^=2PPT:3BAW/1>%-EKM>K&=U
PO@E!S30NP,]Q0UV>P.3DOI==\P(>#ID"28=8>]6^#,\H]H^=]J/( 9DY\P(-CGJ2
PTZ*1%9/=<TICRXFO,-NZ[!5^[N>%5*')RA%R_+*5&&/A0<XR$$M9I+0I\1_H.()"
P @7W]3 ,K]*VM)"[$60TIVSTC)Z0PXOMG8SCG$U5M*\L+1#6&*(L9H[;$E75B@(T
P?U;?KR"_:EP !:9N*D+.^AHAB5TKI0/L*"M"5 *&L"43DO=P7DU(H &U=K+:6^;#
PW7(,:9MJERARLU1T[*3!B*0W3R>X4>R5?RY<XOD5N@EC_S-R(68BYA?C$:13BK0*
P:^;$,',[-92_ !C6B<<$254IN)=]^S^0D &\WVE7 ,HI/%M:; @K9RO!0"[GC6-]
P@8Q^;$11S@Q8I$+U\P-O'UC5\)QYQ+Z9&UJ DYTTQN;/354R!,Z.%AR%IZ"[)>#D
P9V7B9NSE,V( M/EYZ563T^YC[D;B.  5*',/8')ZT>+S+/]XMR-2JZP/ ,+9R#4D
P1OQE<;::J!2:CP_X6TE+F0$:777-HCJLZZM< 2M+003\78%>1+!WQO" Z?:Z-2!O
P@QV ;?;5-$';)EZ-G"F@V;8XX/@KCR5;@C<*>8BH>A^? OEZ8G24;H3[#_N I_S>
PIVKUWS[GOQ;5+G*E#RMIU2GVJR;$ZF:-$=FOU0X'G%4B_]Z_W%\@^D=YB>3ZLEF4
PV 8CN>@A!"!KY5>V)6D=C$HX0->3:.2?'Q9!*<.7UB_W=@+^,,4[HGIP+O]P/%&&
P\\I\6 %5W'A@,23]S7'!TN:@1K7%?(NIEKQF=<<G-CH?ZDL'D 0\VO/FTCO1?(+M
P<-YW*:=[*9LR16J3\_Z?()@F^;UJ'D=E_EHNKH4$5MI%B+816P=J%^=;D>HDO>MV
PY1J"&V,+=M*JR.C=A\&6AM:P]6O(&@E:%$/CUSAU!8AUBJ=D:+;#L [X0*J\DV8B
PS*[_Y#O*;;H_1[FOJ8[WZA&Q_ Q"CZ60*3,9]#+]:!5L-FT62>V/P>1?'-=RO,#G
P!,F6T:]TAQF\PTL,P8(#&DI+H=5DH-R@::/H4?F?/C/%I-K!C-"OQ7T<M\HA#><0
PM[X%QJYJMFTHD!+P+JG,7]<H^)V^XEZJ8>:Q]6=?1N)N(#K=:0CT;L9W'?5_\MW'
P[APF!=P7M3>VR<@3#-EBQ0&' I?"',B;Q,_"_PGQ^$<I]V699YY%0)&M]BG+QD"X
P2_$VY!BO2(%H4H01KT9I'ZK?:H/ELNJ&"V3-/G.A.1D7O6$*5*E#*CO8V^_NPD" 
P7QY4%$J<\-3!<CH5;LGP,<P*15,&%:;L2N;P2?SAAW1W>D(V:U5[#PU.<W5UPI6*
P ET>!I:#95!66@)+#35>VC[9J"BZMZYK7JO\N%/#%7(!.-6++>?Q=WRW#RBY 'LE
PZCR,L L'$%.#;L7>O)>$"8VXDH'/B1FS1(AT9PS'\"R7]& 1]Y39M!(U!,GSL$_)
P'\K&AO>?"8MCJLC:>'3,!O/@A$9IN?%@U08H[O8@B8UN;=45CV#0IS- ;AP7'WIW
PJ7)"F:"K/V8("&$510E)61;'2J6E9U_GZD!;1MN3]4 IL-/%+;K\JF,#)]Z-4:M4
P:BM$XKTG=]D*'*NJ :^C?_3O(D?*-8^&J_@$>?X >4<X(DILP3>UK)8Q%#[Y$OR/
P8)G4A^QPXC!C15$?=B'=63F%:'7E9R<Q@[@L*R-7"K7EOP]EC:'%D%#Q1V.2?ZEM
PM+2G%OUGJ&LG-& 5T -&E,Y9(J'$ +9$<9;X+R+2AH^3 #U$+'N'@.Q*8:C:I[K'
P[ %/W+\L-Z#U-"\CE"FZ5NHO%"<\N\ R[8;,+N0@; )UARE9X1QF))0Z)H:ZBO9L
P\4, I)'F']0E\X&,B"23D!CX-NQ^1)*H8CZM$2.T 94\KB&^U?8_/2%-6]UUP'C^
P1K'_6WL[&7+75]P;MZ:($R9*%DIZI1#*/Z'N?]3HFOO:3:I"T]"E:NHS-0-R>GC4
P;WSC]^+(H:QT6@M@RYKFW];3$ZR:S+7?$PQ25B5W48RC](Y7$W_ A@ZBSX7P8Q?E
P3"9CYED7\I;P;B.O( $TYHC:N(6DW6,8)4>F+D_(\FC6.LB[N#);=7+([1O=:[4;
P\<$Q3;3K"2\"T3OI2$ !ZP*4Q'G4"G3$"S8P?L!#Y#F986Q^1HG&:RN$+9 C "YM
PF_%>33955U-^3,7/Y,^*!D1*B3+SLWH!*4;5KRL6!9L6/.HP?Q3B!HOIR+.>GLD8
PO61?%??EG\[Y<0CH(3U@1VPM YBH8W01*WZ[?[P#=C"1UG=4 X?_=_$OKH\D0N/A
P&8:37C5HY11G/35C9#&( $ (IA! -/>5FN="JN'#-]+0%3"TBK'U@D_0G=_,G?K]
P)-7K1F)"U$@9F>*5A]46:*1DB\D D$I8_ E79Z5"H2>L<A >?4H#[F7"R%I+QLI>
PG.<E*J4[,)5\,[:Z4A>[7N^11O_4_;ECHFH;\<?7'IH':M;S@X("4@A3#R]I6\_#
P2 9@'C05LAZI7L]65Y]D__6BAHE=JB+E6I[K&8)P7.#HX0!_W3(BV1G$BEQ+TMI@
P4?STAOS&>0ST,:.8VU.K#E4:I1<T</%1WAQC#:AW6F,:]()"_4IX[6;9Y.0;W2(T
PC<(6T;,:T#O'-736BR6LQG\EKN09A*_ OKNRD)52",)D#3[ASJ:'@;:I;S76YS8N
P,9U;YJ3TN*B1HUO"$9YY3@5D7HHJMX?6J^?A(8N@>MTQ9QI@(V#U_U]*),U=]6=[
PNIUH4\\T# 8UB,5U:F3J%C$"I9DZR+RH@K9UB=-*WE9+;\48O2"NQGH]<;9_RS'6
P^L0:S_@3'>.,-?S*<XQDS7CW^:RU[[H ]")5W!??"ZL9E/J9=,"6PD]!_I=KQB"$
PYE]],+B.^E4&,0#(-SO:*M00^ =X]9L:L""O92)]TU:L2W?Y192^Y5FMV8/RP[[(
P?C2;K3I7:_8<EVH3]Y*741>;#26:*H'0"6J&1T[/Y#S<T)D31R2Y9C6LO:\5>G]3
P9^*6OK8_+0D-1MX MOZTTOFM4)A]@ H?^!PEMRNJXO,ZZE5IBG,>3#0,'EE:\M7 
P#W7HMT?Z/9OYZ$W><Q@]L%8I .>:?\.A!<(^R>$MB$HN^Q-<&NX/'/\_2ZR>>+)S
P?SL.HL#A0LZGQ^H7&(QC J2]%3(1 _>!POQ%VLUN@?F@1-HG9V1*W A(2_A$0\!\
PZ#AXVK4HN=O_ZT/(0X>0AZ4G,QIEIE=_S:S1J(>N0$85J3KT![ 2:^?0PY9DR#56
PV<4L9S/>-[7;';_^Y*UP1X(.Z0&Q:*$"[]^\$*?4(W%>?!8RV]"A6]FPLS XAU(-
P$^6?$PM6A20 0U=]R,72-7!6H(6,38,:;4>5(M[/GE0"W=L2Y0Z3B[KSM*5"'%;C
PKG9F72#5D8CN[MG+SY.!?TT3"_N\+7U780?0G"<YEAG,&24<,A8(LRD*/&:*>=FF
PKK=@A9>OX-@%#[)#Z8AYY8G_3\Q<=O&2"OA>C;6;D=X,8J_R"W3>#>6[Z+ER*N13
PP_%KYWILQ1)"8^WS+>MU9N-^PPG$\FYL?;9:T0SS*?.;DY*A;4V-4F1,;UIF],J"
PN(1#5IM@\GE**CPL!_+X["U3?&1FXU,(? \6QBS'DMOPL4:HEQ"1A3/@@^ 21+1N
PFUEJ>ICZ\*/#Z1\..@:&7 Z$4N2H#N>1$TV<1K1;)!Q:+M=;V"^Z/>S3WP?%DK\/
PTN $^SSDSY-HMV2+G!)D&%"*#$>R]+3JR1WY=ZI9MR8K_[9?+I@73(@50([_)XR0
P#*9%%N#[OT\<.N75>#?^W4(0CY*2;J#'=/B:#>:801B:FW4/5)H2F5H< LDSQ]7<
P,FV!6:IGS@#?VH@K&-7Z79,>=_C>",VU*[R01X=(::R?.U\_.')4((@_1,]$+LX&
P :Y\#5$MZJZWFW@LJGH=:LQ>GRX>>3J_;9;+G?Z2],!#C>:D1E_NWT&QR#PXL*95
P)?9&]_<1:FL.!+TBE=E*;Q9/IHA?5(('Y]0I52U,8"Q0JF<V=F _@2EK1(.P@A];
PMWTC9ZU/R0G[Y6 ^"=-)QL!KETKFT=8YIP=]AU]]>\VV+W5'K^OL=(L447<0D*\&
PQI49SSIH2P-G"I[9/V0"F"<%F(%G'1ZU1RS*\DUH**)VRNK4S$8,QH'PQEPTN3LN
P$I*?J$C44?P$\A@*PW-,R]8^&M7/;!W(?:#&IS2!&ZE$&P[%.P'7!'6R2#:T#IE7
P0.:Z&5:%*EK)-1-M%W=( 9@<XKWIN#:;TL.440$CNI^LR[=>+6(5>W;GW >\8<T^
PE$.4M.C((62@XZ++0$(S\RL4W9VI^+N>IX\GR&69K5OA(&0T-*?P8R.4@ -A[95V
P3?9X][ZYG]56$%W7"*9T(WU46_Z_O2[7]^S&)2ADI.S,2T<8\5XW*>^V'&*QX]F.
PIS"?:)I?NO3TV9CBIS_['/Q!69C1/_7&(]G)B=41L -!_\F7U86:FW*:KHY#XKO.
P;44T276VM;$+.L5QBW?W"!9TF#I>8?8]5VR]!D2(F\ CQT0!8+X"02YK=TXGM@@&
PN\([^%%+!^FI7#V8_1$+U@#Q1VGXXT,PQ*1;5;)1*:-1H2DK8[Q*L*S+B=^A-L?=
PN1\W\IMU/C&O^]BJ(9H"5X!XNIF^HMSGI9LVHRW$===)AX/:Z6AMEYVH %B0VIN3
`endprotected128

////////////////////////////////////////////////////////////////////////////////////////////////////////////


`protected128
PDU7H_H3X>>IRR,/N?KT7T<0-(GPPGNX7S)K2O6232&=Z/G(,-RG>ZRZJA ?<O-9I
P)6V2^,?I30Z0UI;:@ -Z?*1!@'1Y^7&,6RJ-:V4\!H?_G.6)X8;?_62\MDHU0.4;
P[\^3Q.(**[&[[X#""2BH3FT/_0GHTRGM9A5! C/PH-,JPAOSR:[+N2+S+;S)+@J.
P]"RID+UX8P]"I%;%D2,*8OAUE3IDK[E)B#6R[7M"757I63-02"#EXIFL.K]=<)X*
PKWW"@ ?G60^D+:V+&=(E)VB>:?5'(2U/0Z*P'.,]%&,HF_R6*25)ZGN/:'X(./ $
P0R&+U&F;67Y*(IK$0J)@O8^M-N=__E5BE1F? *IP@KY'8Z$3D74H 1W;+F4@)YI]
PPD=M+3*@K7] IR4S!$MD3>UMAD/ULAF;-M28MKFSY3-H'%=9I#"4;8O.O_R\6-MZ
P]^U_P8Z>@?T3NNB&W+\""?52TOW8:TI]\G/RS#_I^UP+4\LY85(_'KF.K!S=\QZZ
P.26.RU22?!_72D6?.ZZX/(?#RPC<LHOU?TP85SZ=@1IY">F),'8+N'D%<7.BOUF8
P;7U$@.+Y8B,4))+%[,?BK9_/EG7(,7[<X1S(:&+\?-$E,(*T'EB_H$.+$U4_L P_
P[IH0?GGM5ARP.WV(/P[- MH*;BK5:2,+J?"Z?5!*@ KL! F#EDYYTA093EP#;[E 
P3RPJQNHE;[_2W6T1#O5)M-+\ 6KY)IN>M^N-PX]]3Q%BE:S1C.YB)-/0.1;7ONWS
PMO8\IW3<E^R>0+1XZ;^3HPWM>U:],VKRQR59A; =")!Q%2IJHE)6.D,O@(BY.*(C
P1B<<Q3M[T*S;$^?Q!Z.R,$9"?+_Y(KRO[\X9EDMESRXJ[E%]3GC+Z_*#(+Q J-TZ
P,71Z+)%QIAJW0]*?7+-ZM;;Y<F>]RF;'7N%9R^E4:NR;_5K@ZV.3D=$@T\D1[[$O
PY.):/#>S5)Y^A)W.I&R>RQGE>@[VT6_VHI=[_&[8$#:47\,3,AP8,:7.+Q$'5HZ 
P4,H$S"K01-[]G6**M8IM_;4_T22"PHN<8ANA/)0>0:S%'>5H5V=;[8&R/?T.O*E:
P)>Y4O:FW_PUB6F<)."[\.^*>B](+C@.R<4\:ZD-2+FG264[ B%4ZKT^LW_48S3VS
PS3P8)KJ@LN5&M#HF:H1CA"?D\+UKB:R4M1;SWRRQR2SUGBQ8 SFHEU\^DQ.C]#IZ
PJ\F1F/P]DDB_)^QP^[53<%R% ]P:TTAVXI_<WN40)6!UT<(1BQZ)5;6Y#:-EP2!T
P=(<$J"89W&[?H@M[SP)?90)]R+=-UO+/W@0G#U),>9>8=K&-W=CDO//UD*K6 CQ9
PSK8IX[QO7&/U# A9<VX*TF7._M1_J86VV_-6UZN+;)\0L=0F+'3-L'N9CH5%K.24
PH/ XX=;:Q/26(IXRK0Q+?S@Z.:OQ6#VIJ+-I4:UD9P _%9B8YL\9-LJE4%*.EI)K
P;K(\SP-ZBW-)]-T.O0^D"_J1&X('UDE+$OWMAC<'8FK*,]4[G_TS6YW2=F"&@!+8
P[:B8'<]2SP9>PDV@ALR@3<%]YG49[>D4G&^VP]SCR)3<RG_Q-(KMO*/PKT4(23!0
P,;%D'";"=)AE"['P2C'Q?R60=+@_IG)%2.8[]#*@TG\HN:ZAG6=#H8OF(L@>E#8+
P^.WJ@95C,<$7,5'IX[-J!;]<>5(T=U? 6&)0TD(-\G;'& 4A22/!I3:)U(;.Y:ZE
P$R%;V%(6RVWBMGV)> )K%HQX<[Q5J 3R<R'?9M5L@I&(Q^:W\7 1.=U_7^R;J^;A
PNQ\6\G:D.^KM=AT</$-FZ/J#],S9ABZ;,T=$*5MA2YK%F89C[B?E'!SB$ST >$B^
PA!\/TN'(P-864&Q?K$:?N!5E3H\F*:$ROZU_RK/.-U+ATSYRNLNNL)]8N[N,.'G$
PB:;<:\;22&:Y5+I7 #*W*3:$'5\R-_A6'M!@*"J-$P+;W<%+VS/<=L@^1[2.:+I:
P!11EURTU]>]6)Y5(J\8S[59=CS$V^_8$K?X=F'_I$*8IE\!Y:C@)2JJ@R]3Z8N08
P6M: $%>V*1JQ/LFCV&PO<,R2C5?5[\\_GY^J?C*J;@>W>3E@#"%SPDFO.5).H+NO
P/C8KZM;_[3(34-X#!&]X.\Y>5X3'0LR=WU#;:ILZ=83+HRKJ;SK<4A(GT@U(FLE.
PD,@!3K0G0Z>#3EEQ<=:U>H/CT![G8_Z^;/++X][I+H!@)E#4T"])0NU(W?;C@?8Q
PI;BMWBU>=(Q 3ZZE/!LAXNAI%EZSIC,-1;5^T&D8E&"E@6Q81,B=EJ*6\R'Z+'SB
P[N4\"5[WM[2HLOM&L65;U0@"S<U/;+^?-LDA?<_E8#BIUGI9?Y!EU[2VL9TQ*MS5
P(6J9W6_,451.*4UN!]:5$8STT*'Z]R&Z.0F.]0I81V5/"'CE9D,G]',A,P'(/C!<
PY@T @\3(J(<MG]:H]B$/173Y!L_CEF4F"Y-;[3V[7WJ/ZB)>>66.7X@+S\Y'J?,A
PO+57B63CW!07[9A!/D1#W 3WCIH"]-T6GK ^$RNU3'49'0(]+%T0-KU0VZ[<TS2O
P)H5K P:HF_:D%L.>_WKTR&]Q%Y,%?NA<QJ.[U *%!\ZHK-AW>M[LR(94_6_.N6/2
P)K(K_NE*4$KG).:B_,3G?A81\.X0,D5;=2['=V79PS2K\_YX<Y1[0\8"\@(EJZ[^
P%['D23$(&NS]]2."WXE<GXK^L@&@R+N#L  SG_B^<O*4Z^('UQ,A:1I/3XMVAJ_W
P5+O,Y1H"E\:K9UW.=<]EX/W&KRSPATXJYAL0CI?M4$C-[S2.L$+NOTFS'E7%.'EY
PENUB4+ED;LEK +=55#"6-]>0#\*\;P4OAN9MGAN%*P-$JXK!7JR=<V\)4;L.V6\L
PB<F]3P8,0D3B"W^'>B_"I$:LL:,)8>P1J1XGVFX'--Q0M6@U &8$"EKH/F'&)Z?^
PO^;K<:C$W!,_%%CBV_O!&97+=EL"V#K\KHF$_29I6X4UD80_0%%0JACA_ &$X>.?
P%M,M7;CFJR>^LW6-H79\ (2+,?6T4!XJ1ASRTG=_>6U=%\0M'CC+J/>W;""C73_%
P.&[M0H")]1+:MVZ>1Q^J/B%2+MJY$7>>_ F/"(M>^$](3E*'\S"U^U>V-D7^_-R(
P2(FJ0L>4P//PYY%76GXH=V+I2D7@Y=:XSK,YJ5'O/4VTT[(BMC3!.>;\],Z7<O__
PGG>NN";1E8*DJ?$EV* VFKV8&L"X#U71\]:*X%$'MWJ.XLHJQN$(-5;^X:I!7/_P
PNXJ;O0_EM I_WJ9";VG>"'8%59L;<?*F&U)?U1%2L",#'QG3- M$V#'?XKHE1T1Q
PQK$@&1P9H"!/TL=UIX1ADK&VW+2>!KD5N>G5'=(*V $4PNN8@EH;SM/ WY/IC[FL
P8T<=Y^Y7R*WZ.MQ77#6_6\-@9";>('.K(*@F>BCI"IL5R"8H.VAT!YN+2LC^X[/X
PLQD+PTK8'', QZ7<N?[*Q.UC\W#BP__E(=XDWWK&"Y$FQV##)[$N<..G*Z0_#29O
P% \)P-9,SK((8#R#7WL)@W2E>2)35Y@UIB/T>P_-2\>=/U>H^+<!DN@'Y/\[\?JF
P.@7&C8KL*0K*I!@2!<F^E*GEHG[VBQ-:B*[R[5!BO%)5<YKE+\FRU9+\%6[\HK)F
P!V#,&'%PC GP)""-4NAM#V^/7;YL^%&02)^#M=R2,I3#H_YI=#7[_,P/?_"*@C)F
P!,V?I71(R=]QOS*I+"U(A<,M6W">@ECP 1*?*E/W/PGH%U12 G\0V=*M$_(^0,HU
PP2=EEBTT3^'"+#UH8FUY.E??+<F:QV9JO^,8'@'ICGV[)S)5.QD!D@6V-FJ+[9BQ
PA;;(3'PH*'_Y#I_&8P5 CU%'0EN<+0JUC+NHM4)-D'8< I&%UF4$?PO7)61(XI$P
P(Z(+7M=_+BT:267FAK,]1;W!RH^X/SGDZKE13UJJ\.H.U O3EKK5^XH9),*-)*>5
P&&/ZJPH*I\QH ]'P:;FQ;+9H%]#_'Y!%%L.CA<CEN\XVMHB\95+?:9"8U7@9+C^5
PSI\M8@''RPHM+)IX6<MXV9&?0@?4] H[^2"DW)GBC!U T[5R])RI<U+I&$<(F::>
P.^<WO7Q8I:)@)QZ+$*89W SC:Q)>W1]V]EL4O2%7 ,6OHDON^DT=1P';<:7N^.6K
P(?C8^'%O':$^@.649E:LZ7]6T%!JT#ET+300U,K(R7[\:773N0 GKX)2%_;ZBZFM
`endprotected128

////////////////////////////////////////////////////////////////////////////////////////////////////////////


`protected128
PDU7H_H3X>>IRR,/N?KT7T<0-(GPPGNX7S)K2O6232&=Z/G(,-RG>ZRZJA ?<O-9I
P)6V2^,?I30Z0UI;:@ -Z?$3XLS,,J0D*2Y<,UBQ,W84;DD5A7_A4(:'08:(&,=OQ
PA/YMX9@X2L$E?!8&C!PF;3->!PS5#C5VL.87D$_ \K<)2]^M4" FCPT?^;4-CK=^
P52C!&]@T/&6?+B,7O(4GE79VU_X&?W,2Q6UY0'HGW!O\[P5HV(T$ /!( BNG\VO.
PAOLY\>UT)<9?N*)H?\'?W(B9@(&IO4\[RW;L)P)W/K_=:D;10/H[V$Y*#S;**^7U
PI(<.4")#3T"T"<<B$@<%U'*4"^0/^$4R]X2L'3  J,1W_Y[58F>YS$P+ 2OA)=JC
P"=>ZE*D &N8DF_9UVI,=OTF]$K,WFG!$J'E;"X$[,DKRI',RH!*\!A7#7T=U69X 
PL)%Q"QT2[B!&3S4HN 6AT-]:K330&+DXR*,3A0S<SXNE<[O=&-2$\[+93V:CU.0Q
P;^8*/*)&W_[LREZ2*$Q^JTUS^(Q^_KIY_KN=%"C(:F1; <NLLX;8XM@V_J?"=I \
PG9_=$/)-NY*4]WI<&]R&OFZ40L1(/!+V7*:7>J;T0;)!U"]"WUY.+'V:S;6,I!V[
P<(.5A< @14]=D<\;0C<BWW]1<:<WB$-'E>9#8/*[=2CD.,\0A,_%_\(HR=^&MO+R
P]0NJ+FBGC>L_ ,]ZM=-17O]-5U?6_W<^2(+6-UCB ], 4"1DW_H #BW@+JYV7MV7
P\,Z9;+ F+O[&%@W1YB2NGL(5%5[ ,Y_:[B$"W>:E3(<<&G9(P8+L2H8QCW*\(OM&
PRD^XS.0R:">R3%0,QU YEDB!?=$WE2&5Y W(>%')=;9&M-W 34!F8YD>;^DH+S[[
PIU)5NRN@Q%YKY?5F-$71@9^G[*,( $H%+&:A7G]N-_/[$8QBQ?WQR)A>.$!$]($3
P5*75ITD!:VH^L$>N4C*C#<V?LJFNYO+1)Y0S^'/,0#5$&C*7V-!$M2C/SP;/"#6Y
P9V/$K[=3'MP+9:NI\+5FWI^VA4912VJ">&-0-L>45P=YWO9U);)F2%>;;V$D03=E
P4)I2&1W&UR'$67G5T.?TKO:2!L]Y*PA3JDJ<YM:V_09C^[WHP$*^4?X&J;<L3\6'
P3N^!P"(&2:Q!4I?@77/O>EC%?QGO I@6/I]T0M0S0?57[YH"JY3%A30^&?K65C*8
P-SX@9D+/$C?+D5W#])%3*HT"*3N>E'AJ [D<Z2_S-RJ7/ L:0M$,JFR'VI/ N24$
P6@44"?+W2R+=!,M.G<'X5%!B!?NV8DAKD7H^VH48F6Y;B$V*:$FF%QQ)WN",KW<V
PHDH;,& J%47&&>+=7=;(N&_G6(2Y&#6[@;%/3%?H">(<Y)0H/X;X9WDO#8,)ZT\=
PS!T?>VY@SM +:"M="C3P#K&:D:@\EN10KB3.-EL(:L-XE'H[J>B@BZ/?/>WK$=@4
P 6$QZ-C]2ONH_MP-?LUWR;?1_3R$#X?LH';!X,&= AK_6V%Q$QJ4=(:+-"&8*6AS
P %7.ZAWN,R8E#@73[*/#5IXD+@O Y-RGZV&O)K\;X&3.F.1YJCE7_(0TC+X=H4#4
P]S+S8^+F6UQY6"&Y58!*4LK)@$@1I'RON%8HHA%A?9]F LFHC^"'M5_V H]4DVOM
PXG4$M0.8>_:A8J-NLPAKMQ X%<40P/2G\DO+!L5+YOJO7X5KI3API4#!"_[:07WT
P0N,;5X#V;W$RI]4J&];*\ADKSU.VT07[1^_#*N72LA)YT-\[9BTK:S<&U5R?"%JD
P(WX;?S<W-"4#M?,-/(].RA*"+/)2IL1F-DZ]X\584;[2A09K=D'YNH73IO#J26 C
P"196Y6]E+PZ<C^X7V-S8@]85NP7BS@P)U 8-@-(TYK]S2R*DKD06KN]1#T&5=TAH
P-6#H:!V.9]Q/[0O;A-TZ>AM-<4LTWV'N: BC;X^D:U+[BZHY_?:LUZD^C+O^,\I7
PJ0;2$!:(*93GM--$SGAS1^<>\CJ;]\^R) 3_Y4X;&PHEZ;4,2W@4)EYEK?>-=VF9
P?(PHL_G3B)&<(&66&U(IZ*E^;%P;-&A-+.]ASC"/F'530I2&Z]S_<M#H6H+N)%F$
P9E$VVB]Z+JUOJ: ?F13<^$4S]<PO)Z/,!-H,^GJ(TF0?R;C2E;O=03HYE*WBT4 Y
P TU!"6%5LM V-#6G3UNN().'OMY?6?[[*B@PQ E0L**VS@CQ5^%VW:+793B84/GP
P-+V19+OF0(_R5P!TM$B%XLNP($4A06(,07)G-JA29(?R""\$F8J$MZ<UA?0YL<+ 
PW]^=#I"WNT(TY(;T0\I; E#Q9LP@6N*H!;\-1J>Z*-BR"A8_3&@6C1P@W4%IKOD'
PPVBJKAZTKF6G-,/;-5FNG(7:578$ (?; QUM&5X@V+'NXIF^?JZHE\QAPT@-V4\<
PA=_J6Y\\'>^I"4^K):K=J@ ,X2,#U1BH<9Y&ISI\IV XCWW';*Q!C&K7:_"4=.[\
PWME_.+,=UP6-NQCNDVO-#H5<NOG$K-1\C#!)F@8<#Q_YJ.)AT,FV77MD EU@'@S%
P*$]+3YY5J-^V#@?#,%!J<PVZ_7^XC L82B5N,'O\#6WB<27^%?RH+^-)J,-/IML#
P;Q- >[2)*B4V.EB@W\"9I6#V?->K-47T-W:YU\M2GUQ35ZA]\C%Y=EB@ &^W;KB*
P[M9"QWI$W-9(E:&]2]\EW.H^AR>>=>C,X(1KVT!.V]?KTI;_T"T'N@X^+#&,$TC8
P@+302U'R';;Q@VS*C__JNR/E>G@?@VYC[%@X(97)V-3C,?M-_1#K&\BI%*INE\93
P8ZQ15IXU^LKO"X%VW]\UKR_Y/EK$B%=GV<=3S^C>_]3[UK2/6O=BW6N=ARSLE1LQ
P'MNC-'U7@9P V[WLMLF+K3&T]%6&*0%*D(OQT[4 UF9;OM"J6*(F3*R_*U[5'&JL
P:2I8*!K/NP'+\J*<13WFK_.GX,OT$>#4__6 P3J^28N,W;BQ*">U]<$PJDLV(NG:
PJ<95T-QAO^8^PI<_TH-T'C;$K;(<JG"Q#&]X _ZE9)3=FOK!XN>KD7WFQFJ12O)7
P_7#$HFC?2Q;^FM4_Y.+A+*WWJU\I9&I?1)0O;@3LE"RV=.AC\K[X)V(@X]S)MM=)
PV;SN;<8( _+YQI:BJ*C3\IKI_[8.""&%C^U]>EFT8KD,XK3W*QE_6%7,07H='9*V
PYQ[@HG/=6M2^'.26;6@B#'*,'IH7'1[JZ=IW>-I75VMUV*$*^X9?H!.9=*T1UGPA
PJ),&82(=)VM&I?I:W_A=)$3V%@O**.?Z)C+2+!5GKX+R]_[VV5UL[$2C1NAS"+WR
P$K@^972.KB:WROOZ+^>IQ*M]#1P1_"<YU@VJ08_@)NRY?B#['E_*=-?1D&2O"V29
PYC06=;FQ"TOH:H35T=8/L2.TSS0O.;*1_0.F9RH9ES/NLO6P4DM^7.\9V&?_ITPZ
P'O@P&,7=''GKA%?/48'N&=972 /A=T^5J3O.SY5L_ ?.QT*F9R#V/%VK0)BSJ\8_
`endprotected128

////////////////////////////////////////////////////////////////////////////////////////////////////////////


`protected128
PDU7H_H3X>>IRR,/N?KT7T<0-(GPPGNX7S)K2O6232&=Z/G(,-RG>ZRZJA ?<O-9I
P)6V2^,?I30Z0UI;:@ -Z?*1!@'1Y^7&,6RJ-:V4\!H>KO4'MHP7SHZ3X7 ?6]I8:
P4R#0X1'4NZF=ISI_+/JD1\@7E6L,ZVM#__7[E O*^!E,(KO@/ZYBW,=.W3CUT1Q\
PZ4X8W'+7$!!NMZ-:[ 9J*@>,YG";UOJ%.3';VU >!(UJD1]C=YVK'@8H=LV@-[.]
P:[)22&FJL. BYZ6V$I]@D-8F>V%A8CTDNV;M<4ZTI06-.#D6)"WPM$G-( B<0!)N
P: D8;RQUJX^;C1F8EY&[ F_^Z6U$C_]T#ZP/&AY0=#IK:M"BJ]Z\.I4ZWV^9$LJY
P(ROIF 6!"NN=I*84YC: J9A2' ^BCB5C$9F,'<B*W/M<%9_MA-M#'$^7[8H?<C#(
P J7&A_UDDQ#V L&\(N6N?%OP(R2V1F<!KV)-!9AK#;7RMVR8=OC;ZI47<JYUE*19
PW#JN;="N$MZ$+:-L,%S5)O"['9C2%"K'N7P\GAM;0=UT_:C%Q,4D1 O5FKORB'")
PFKMQHL.YF'E%GJ-(X?<,'07XO8A4<*BL]C"[MU#CE3+AQ?MK)TY8%3X$]UU6-J(A
P<? D^XYQ= WOYN/O):)AG9R9>2[W;7Z=S+,6^_1K$Y@K%YYTC_FB]XHE>KO3WPS<
P0@'S#2%4J/D;;+'J8Q47SG"AYGGE@]<#Z+T #66PFSN0Y7-O^ 0=:&4;//0VF,,(
PE@XY$V:HM[@5=$?3.6*. WU\\C]2B6=V;KNY6J'166^$Z%9HO#GIT3?4_MU?_'KI
PK&22 &L$[E$']5U:;U=SP48W@U/OM![>VWP'X=,7*@2C4*@\]*G2=7I4KVBP",PB
PG.@+2ACTP3&P4[]<IPAT&<4DH^_WD%<?P[1F\3YU> <XP3I,PW;W25N\4>TL%BVR
POC3 3>3H?.SG8(1(*ZYQC+I+9V-B3HN$<EU@>SMJT^.=CV4H?L5X>E8Y-[<,(L5F
P4QEB#"B(,[ V84 $*"_27*OZA_B,5XYY&>P:OC#N>KFQ,IW@Y-671>>SE?,! %HC
PW_D7 LHZ6^DQ'9TN.2*-/JZ&#)?OI;:'C7_C6=Z,D3+5RT<T-KV5(?%3^_A::JTA
P1CP*%L&0SROP:5ZPHGTJZ+M&6R%\/0RY/]\)*N+X"Q6MJW/R'OPNFF[_?I7J/GP.
P/[]R!KZM4)N*IXP<WBQWCNZ0:BC^,SEP?_ GN^P@W:1-_N@:$LGBH!VL]OX-$'S6
P4$)&YHI9[GX5T?OJUC2,1HKK:JLAJHU^/PAYFK63,\@XHK*Q;F,I/LDWV(TW;:6>
PR&]KSDT^9O,5I0=\XJ$Q,2USVR-:+P\$1Z!A= -9\7B+4(?MO:4K?!X*$ XZ_7T5
P'6.@%Y3/GY?^ ):3_NDM@L=-_8$)/( I#]U]6RS@,^!0RZU^E3"ZM63,PZB^]H4 
PEFV1F2+?#/]J<H&K1+( 77!,6FGI^==.&"!,6P+4=\]\>!W6U7-=?I(82$@F_"82
PAJ22TX@,7M%YEDJG_*:E#74BS:J("((@5>LV,)@;*)BLZYD69W?7&;KEIEYS;O6U
P>WT8?D ?PBYHB[#-AV42](!%P!'74&6W_RA9D+4$N-2EEOGJ3DPIS7WE\Y?P[R@?
P&T1!MV%!:?<0ABVW?,'L8>4HSH@P_W2V00$Z?X2NX>5I6O8%D\8RPN*_]RS_T6>^
P+V,7 CK^UR0LHC6,$;GD=Q5NQ8S;Q<KBI:6"PNZKS7ST%J#8G^(]$;V]G[CF@1LW
P-^GVD+6Z^X(?,4XA:V*ZQ1_1^2I8V<V1T"+Q2=L9W>Q5A.%P-;L%YFRDZCMGM[ZJ
PVTN27K6D5 @]-TLQ(/P>WE[+_O&(4VBG.ZYNJP#*$/C^3S118;U?.^>"U9CFP?=W
PS9I*2#M,[J*AL=6X]8^9&"1M?Q=[7RV7HW=2'&S Q^SXIT979!;-,HL76@]*F^O/
P549++,\D5+F#S55O-U?(4EYX(=LM$TF*0VV_EC#AD?D^]G&9V;]:R3PB6T[M:1-,
PAGC;R6HZHXAG5M^40K>]#0G'OFC)P>;R#9)XTT8)^W,TFV?_$3Y<XBH;\FE@'HE&
PTF H!7I$4-VIK6!6;4[4;$P7*"K^Z@+G:W'N+1A-:4^4:JQ9?V\& VT5_<R/2)T%
P1:YX5QJ6-Z]Q8V7+ O06<KG<JFZD1 5-)4=2I"$F!JSPXG/+M*C@02- Y^ /0[U%
P7<+ZF2+D7T#P# LUZ1KMK)\/N"C]Z9YHTU\-4F6-,37>(NA?V*I//HY[.<D##&!<
PSN=?TSSN9&M5]X]LG>_F?-_?LL83Z]79%8P,OMY=L56!-_GJ+D;#BRJ*<F?@$6)"
P1E2C>GP0_5RJ7*RY$3MC?)G'<U:BG@]9=2DV#-M\WGA$QGY"",A,UG2(;P("R8.H
PJ3A0%ZJ4++<_!98;/R19]F_[/G^3Q RKU*&JI$EU0KMGZ2;0&%KT51<F.%,V+U\ 
P1J%,.LS#+EJV98(2L[Q[.O7U:N=L@_EH>;4&4P1[DM;7#RP#$ =8Q&,\TCF_?@C7
PA4)?'I6-]I;SCKGE\,%]M82=Y=11IUB:R+LP-.L9'9UL]N'RCJ%GWDWWI#'@R].-
P8&:G+O(&E1F;Q43,..$=JSS2MZA[\<7VAFKW<V;4#^H+GO@C>\QT1Z46AII[];$W
PA^0:&H[XA5[&/V!0MRA[AUQ9]T46C,GN4%?QQ^_IY6+E3BJ:M4*F79OZQZ>UIX]H
P'VB*,7/'5F>OT-A([7N_SE">@HH+_TOWJBO*N?4'@]SO\K9+DCI6HK1\.@1F65$_
PTZ^JWLB#]&W<TYZ//G P/R#35!/K1X1,HSPQ]8IS3/($U\0JJC%'B4NC%45G;'K5
PN'I'@[A4VVS)GA\GEVAWJH_S9N))*1XD7OG%A&]+4G7.Q9U44L:LN?P(<RE,D I4
PN;>';0A(RF+O7BNIZ=<*"4V9N859U7J?CB<AML<(4N5?O#[14:IXD...G(&%(:2[
P\#!AKBY#/3&#HA3!A1[TZ7VTP:;[&?1G-6LIU,TK73E"IWP+RDD>B[4<$6)_(AM(
P4UUUQC7>@D;I"T7?X(6-<*#L"F)^T3R?L0'>H-#*!TYY:-Q>X#UFTT&:$($G.$Y*
PU ]LI*7F@N*-6@:G(SO%!CS*OR^YAN3@RD?RS4,Z$U W(<$#7I3,OO7(4++-0GN>
PS382#FP5*H/-FNJW/4_].+!%*:9JN&SFFR #]JBL/A'3EIO-&-UZ$N9R^K--,?H3
PJR94Z4&EO<VQPR_=1-M&3ZI64FQFM$[PL.>J-22M:7V;]QGUBS>GU>>VF^GM,2G[
P)JK" SSA *#[>;MZ0#587A<<_,*L*4^"0D6M-P6N6O@V\1(+9, MY"'-O0]Z5MF1
PG]1>B2,;!L&7-&B=Y1T '7;63Y\@:^J:[%7I@5:8"+O26VAFG:= 8'FJJ=Z=.%:P
PAI]+E<MT*NN50)U\9#(U/1S%5LZB8<<2Z>*/WC(,AGZ,#V+\>PT.$I0C1P"?QES9
P1@/N^Q]4BO2T(,0 4<>DNC_17A#5]HVI';$<K_"[_H.)OK),9HN,H.?:(3M'B,$/
P 9$$:'BJ<3&EZ]O8[5M5.F[%%P#N5@/?$85-]_D4H\[#Y,45@16%HRJO1O1[/[OP
PH-3381:YM?50C[E1P#S'XM#?'RC?J7^"V<0O;1C)ZL_12Y7A0HNKXO:-L)[5=R)D
P'VG."VF:CK4M9X0"O3:[HO<E'4WO!\V]-SY>.B7XY4:8LC! 6"'WNTB:45IS9SSK
PZ GZE)K.U*.I[-@TKRQ;@T[ 4[9%0JK+BLR< IN]C@47UQ3$>F#\I!#HD^(QF8,-
PO_4467O2-]%HBP#.F+SM;!7L233@]3$U)S_09AQL2&7<O#C1Z*'IB5@E!4=1O"YP
PX=0!K@(]-,$5^[1!%P_=O,J?31 K/I%,55EA=5+<M<E7IVDWHY2^!&^,S_IC.9W-
P%Y*-*J3PVEC^F0]MY9PG33O"*KA>"'#HX#TF\<H0XH=R("+"0'U[;8R@"R>8'TB[
PRB(ORHP5*TZ)I=:\W:NX5=<L8BFKN-E#0\Y67V@[6I!;D.4L=GUF?>Q>(X&L44GA
PB3#',@HDY(AH$_;DK+;HDBUKK=#$FB@M/-):K>\;KA3UG1*7CO E'/)%-*'EO%/;
PJ*,N51!WSXP#9 BP,R/T/.0<\&(WHJ G-CQ+8_[0 TS]?4?9RV($<@(=<1A^SE5]
PNR>K@T).^-7#<T\C!"<,4"5T/C#[X!/;&L+X[S?H23FU6-DKJ7F9B:MO"J,E N"B
PWO%9>>X60+=&@D]JA=)/(T![A".L?_V52WK_)6:_M?JYVY1K0_<C-*)W.6AY7/@&
P*;%X!-H<CHI6>B;VHV ,8C%F-<H)VITX4CW8"J#1 /_XYS*VZ$*##46>B#R4!WST
PG;40-B6@]K"FO/+1E5446H< _13@V2+VO]$P0H;4[NA.+A?EBTF^![(:^XNL(2/4
PLTDF0,2Y^)@(A_:-N:D=RLT!"!.X26F9<_ !S6AI>$=?>"H,8;1Q%_RUHS3']:_G
P>&V%INU[Z#SV[AY4:@ ;E\7SD[3>@<N'7("XN\M3V_7E@& EA;68?C>M9Y3JJ]*0
PFTR:4/?OC@*3R(?UB6SU;E<$"@1Z^DGNYTLK,XR!+E79>?BDB)W0_C1%S47!.(C4
P>5\G;N@H:5TKHD*6Z=0^4+ 0%7:,UEQ]X3!R '&ZTIX4,@DM>1A09,V/!@O\?/9R
P'DO:.SV9^?F=$BCZRS0%$1_280\Z[>0]"L&K>:H8G6Y%T[5VID7YC:=5SH_!F"QJ
PNNK-V/>).KT=&Y[I:[B<%E$7J_.MM1.%13^(:CE1M_8Q;4 CI -)0@#;L\$S\]E>
P4ET".YJE,7N($BD3L-K@4&RM)N/\HG1P)2:;P(YH1')!VZ@@1(GU]4*&19A@*%$-
P/G:7#FE6$R/UH(J6PLY(6_A+HG+]##+;S8WS*:2W!8K9K>#;Q@)2Q*P#F4@T+Q4T
P"V^PIE;B]"#. )LBC=@ <Z-N_(?$J(#[X?&. F9[^@:(PD4R#IQW&^%!J09MG@,=
PF$5P$:*N#EOD*2HIT$#E:<TRV$H)YV LH"(?4Q;?:G59QY2<_*VG;H@-VQI)+I";
PC8@;-RT(>GFGDN?"@4##IT 7Y#6 V;VD&DX@M KYNF/Y5JT97_2-XAA8(/KY$ %?
P&M5C@@FRFJ5J ]B8D#,,8=)5R\1/D$C W_B-',-97"0Q(4/2 L"?B_DUH#6\VV7Y
PRVVCD7,+ 40WKF>R7,W1\:3?@7?<*>,ENKA4U_A2K<[_NR&DZ,>-WUM'K,.16"QL
PNY'9PW?O^2>NXU&'YV%9?"&I@Q]6B*SU$,+O]N+5U"&K%&"HZ@8&Q(8X9K\I<QR_
P)5"P'>6N#<6VU_R'Z!6WU,')+$VP1%\%%,H:X&>=_0N>/M=SK";P..XVA[ $^K\!
P6]V?WLLP?BHXU$SN/MB^T/CX_C>W_TRWYV!?_R>=&:N-G7'G<2R1LI1\M<!D<+!X
P@]2ZT^KB!!AKS0%'W6C(*K"(%+]':/'JO+46)+ZG2ENNP?*A[7LS#3\T,$(5,G=;
P/, ;CX:]F4>ACFVK+.NX9.X27M^^O!1W]2N: Y9B4&12UIX.;@3SDJJQY(C(<UP\
P#;[3-_>RY!S6R-?D7[C6(/F<NB]^C(<B9]&_Y;C(4F5.FYBY(^KS:A#W\SD\5'OK
PO_\:@+R^IM/?P8*7%N(_D&!KY+@0'.-S+=A\=I#8X1HDFM"JAXU)*=?IF7!W[.0E
P"UT&OY\N5:X%Z'7CB'29X;9G+ZWP#4;TA2'.3BKVZYAEQ*VL<LGGP<%'QR:ORX+X
P%AI,,,EV>TUO>//M+9.4-8U'Z\A*,6LG@5OJ^O;!N >&2X>"_@9%8-"AZ3564,:'
PN?@.,Z#D!UJ"=;$**PINC! CO:WE$>9JI304LS(H1I6=%:1YX %<YD_E$XX+@_A-
PB?,KWLT\3Q,KCEOVZTQ"$:GU2>C/A#$D9@"Q%'QR)9@18M9('O$G7(4\TQ486L&7
P25E])OO?_!7G/"!ADKWMFC@I64;P^5I71 OKKXD%,GBQRVS?]K3O\EQ?FP-1)/"I
P0>HW+S3,+-#T. W#$/A2#M%-V$3U,Z:=#_["NM\P+.++PG,#7)1Z BIU[0?R@^RX
P;=>21?NJ"0AEL7J&*TO'XY;OLW"+>8PBZ[7'$Y,1QY2\M*F^V,TWMY'X/ H"ST?B
P(3]'6 7X*+*VI00)RB[*[20JI V\VE-HZJ6BC$VYLD0(2O##E0ZVJ3#@ HXX:$_4
P[T;M,0OD@4Q)BG0Y>;*IEUQ.S>7FY$AOL\__53;2+5+8R+RN7SD./VOT/@1.1*![
P@_*'".4T<KDPC[T.,PI?L;<G*ME+TM?*GMP20XF"-PN!-*-#",G2[MV^!X3/[/#"
PF+#IA309TONYD<7.;!%N:.2G/;3.:KUZ=68)H-#\*M1L,S!&KDKBA@-+ $-Z\?',
P75IN+RK],TMW(MGB@_]2_-X1:NP=4;+JWK32!49!>]2U\W@ -<YU$*@;+R,-%4^Q
PQ4X)S.N3_A6FM]-DI0@T_H3 6K< D7^=PN#%*H&(+_YK=75RBIVJA9.+'6ZG0NZ\
PV7A_10OV,B5<&:@NK*&\R5AX^V>V_[8PP <5H#R@O1^\SWFC&LS$ZFN_?KXGE\]N
P@$Q(AF@/5ZG4DL+A,T5!E"]A \CPC@#&:BF8WU ;QVQ%E9ET8+#G()4<_&Z@^?A+
P 3R--0SUN!--?I/ZY:8CC/27NP[8/3'Q#,"4:UJ#I'(C$6<V$/]\!+D:GH;<V4CO
P@]><^B4.I'T"OI#ST^$811J7*+V6G-TFG1J*U:O@;@8J!J%L '_EZKQ@;V\7L^"Z
P%8\?Z.ESPU_YZLBRI(_T45U%ECP(O:Q!;#":+NTF(]4WOSXF+8@%'!LT@L'E0N#2
P^R2/NAEN6HI^'.E2+-403W?/WG#0>D PJUD#Q A/F*O6.Q75<AR4%_FY &D;VZJG
P@BP'UR;F9KAM ?="\>8(T-?)8\I1#8][4\G+8\@I#NR+?,(:0*QLK>W?5NUO58CK
P\7A9^ *&X@YB&Z%KYOW;O<;"";H^>25EG:T&*_/X:I ;4-,KK;(1<'DZW;Z^4EI<
P=3!$A%P8[^GVR#N *_T5NT.MF^"V-H>RBZY;BREJ[>K1O<^1\4@ ;68#UC=\:J6;
PRQQ9T5J:#63>[^+#W+,=]!(3Q5Y<_?B[W\<0",00*HNP=MAIX61M<_P$V%N)M=+#
P'B;I33)GEZG9;!>EE4!N"TOAN=&@&M?.^NH5<LOP$4=:()S[B!,F:Z2:?ZVNL"B^
PPO-GT]NNY-*)GJOIYZO"U[1WWG\!RW",NH^/5,!"9#S9W/N<>8KR$B PQN*-J;-N
P+BO\9$AC@@YDYT;QJ 824QFCBR!]^V=0I?Z2UCLL%S.>FXC:/-<F!U;@0IF(^4/Z
PUL[ #)N#FE>N6?S/G+#F^;"%B9Z*$.<\.$,E&Y[A33^4*)Y9YQHI+;)!;XAT!]QW
PGH.A#G=1ME(-,/<FE$DVH)F?/Q?A2Q)?GBT0<I4N8^>12\G4]"O#I(Z.B\7_B;K0
P"[W(1><Z@%>R9=I"$/9DB# :C?G+$((@SQ%#(M?PK1?7ZV _D.@7&[*;^W;[B);J
P1%%.&@9V3OT3IF<6V)C_-ZTIT5[4X%:"T85X;!CJ[M!(4L M,P_I!4!+<82E 659
P6H0/>>;G^_&*Q7>A'5(#A/,"E5@!2*2!<>2]WJ7;&+I4HQ%++$@"R H1<%X"Q6 Q
P==YQ:)"]IY:X/AV>PM5;I.*@-<)PC89J(1$ @[FZ$E.,!.;SGY(@7F 4TZ<?3S7;
PP6?'V%A2+*PVGN"Z=BZV7OX51O,&8(6FDUZW((/3Z091%>NVQE["VK^FOW0H0BT2
P2VYOL@X*<VA;\N:APG?E%XS!9Q_)NEA."CL\3&HK.8\=EMNC!P"^ :J7U=W;=ZOS
PCX'27:PQ=HN#@PSU$"L!&*-$H/MQQN"#)WZDC\@SDJF,$&C6&\A6]LKB3PLI//1)
PV/QO'5+\'LILX_<(+9!<*9[Q>N-2/0W9$A&33T$GM3-8CY_1OY'YW5S) 0,VCCY6
P+AB_>-,=KBSYL! <\D-:B:-D)W^T)VY,#U #F#*_SK6"8L+(LE1 O]KFS_U=>2G]
PM@H#DI:IR5EM%O2-#?#W?\=MM>4/;P?IP0>J>H_8PO^XG3</._+;[__9.N8OU]BH
P,"LGU-7),YZYX]Q*>? $=(FU?%99==/'3 *PI"%Q!3I6B<( =A[OX%)I: N\ ;]H
PU99NIE%8>V:_\MZ*B\S*?NZX&C*O8\E%M>C9<&A4BXYB^'WXF8 E_#9[86@0" $*
PV=F;($R^A]=[,C;7SXC>A^-#9HE'O][VKR5>FX'#QJIU*S<;0QNIX9Z*H]PZ3SW6
PY/K;/GS,#+><"O\Q0=W&(-G&)5%@8%)#(21R-J!>0G-.MMTB[/\M+V.EFA_B\^L[
P5$(8Y.5C^GZ)=^#5>2FCAA##V*0Y"(\Z<)Y$UL%I;8-X?77\#)K3?L4@\7T8 /6^
P8]3+K?^*ZNEW'5*3W1Z+9N,&*[VIFL =X$,;K3=@0"N/>KJ9[CD#88RO"1&B"#^*
P1,8PNNH9WHUNB"LPW RPF8>961+?6?A55S5^LA_H#]+M)>6N2G-_,E11NAVWXF[V
PKY7+U9-<\AZZ&^]&P[KSIITVS++]@9Q]3"1]!8"U[CPP[QT9)P7TF;XIT+RS'!%*
PKM [X9.3?#HL'[C PS?%G"C1P<_&$TP<G)3)K][ SJLF*_/YW)/(T\V;X3X%7!#!
P+_A9%Z.^':[2RVM 9;@;N'-6+](U8^P6$I7]U !#)QX@28TS;XNWUWLX8988@A9@
P(^P: 24/.R.*_%2,5-MSF'-I7<.2&SFO,HK4(NJ0 #'T,7B &>11(@T8?"]@4;M[
P1']U@]DS7I@<:<6,V;<+<\#&Q<_7 D)S/O4<EU\P@BDX%8RO(\Y^10OZ]UMV&#HN
PK]M8/\,H9^6-)2.AZH,Y,1D4 ?RC9EUG8I-U)?I#[AVO3[QSS\"*&O4EZY)\.!6<
P3YZUF"-=0GJZ'NW #!;].-*E1'#HERS3.IG"6D4:F:A_R-(T#6*;, :Y@7E;-TT&
P#>6 \U)W[$4;9.M(H/+">XZ26[_0DI#;R".UK?'!TX+)N"9X;?D!OO3LO7DD[^Y*
PH*SF\'9VX9=NB_@U)Z=-*4#F$L:]@F]A^7XH/7G/'U-(],5!%NA"%.3>M_*ONQ<2
PTS2KXHEC&4=4$$7(+;\5&,< AJQBD=33+Z4!8OB85GX@50KSEA_S0V2C@"9"5SH'
P46?^,2JHDMJ$= Q7*6K*R1JX/HQ!'4-:D UF>BNC=@)^$V"1X+&PX>4Z"[Z8@(;Y
P%*A53%V].OA;:QA?9V>3:LT=$F8YB,U*'VW"55AL04"))(,PCL#/PU= : S'0^&(
PB=T8&705=+W#EI0_$9\*CW,&N&$PB#'"=_>Z0&P-+C\@< BC[K4O9!BQ1,CXES8A
P:493,M_UR,@0K ])W@%OT5Y7\ I^H*-U 4\OX VM#:'_-_Y^@6  8A-UB:CX']WH
P#\Q3?'3VE1*3UFJ-C"HU@@%+FO2_="\O0K%V"EJH M<./D>@>8#P/R%=[.5RNLO6
P79GQ1PQDBMS=>K_"<)JWU<S&1_-'^BC+6F<3,:DYL19PJ\V,&$T+7>8E.\R4/HR9
PD%AM$DDCM/]%DV:'6PHKHV;> QPAN\MB.R/.C^Q2B.0O!*:[B8N9N'V=FO!/FUGY
P-6XJRS7;MB_[IGK0Y64CJ7$STZADP(LJ&+G(60"I&Y"9.NKV3AO]Q DE%SJND=))
PQ<RYP)?AV@:@P!B'"FRM3S)&0,5*O\."$T<"%(=SSQ7C4\RU<+><-W[HF+M6P/. 
P;!V?J3,#FW+SGO''7=F*IG,RBYB$*(1=+4I;,9\#POW.+\I5JA="*TMAS\Y=^GCH
P&\97:OOE]I[DA6L8U!4C+Q$>$GA$Z>4K-'HMJJM0W&0_UCCAQ%!A80H*D"#PYZ* 
PS^ YO7 )B+ALP"Z\D).V3TW/:,!317.0<]:FV>4B79]"XY ,Z?I/=2[^ITE[9Y:S
PPL+Z<1B6Z_[L6W6_]YG1G#C3">@FELF/3KN"YD)KN<TGZ/8$6$^6^C,=E1M_Q1]+
PICC"(,/F[^,BJT7DC'5[&G<(X1BDX:*9.;.R28V?RO()WREUA4C>*<,-).!]CIYW
PD<[L:TK2))M?15W"K&?.W;@JFVIF>#W\YS3I?O"VQG9-"+))]HA.%;>T[=,9LUV;
P6@E(.MD=?1=U6%;0N_@#X[935AD)F\/(;; )AKKU&6-FH:E*)5)/65@5 Y;)!L[]
PV@U?'GQQI!UB\+Z>JEE$B1ZNNJ^/]XK]E].RT 20FUW-5!=U']M<56[;!,*]#Q%!
PL"#"3ST;1@M?1S%'@ZV^>2,^(5/=$FW' !9*F,9PF!)PM%3XKL4H[$RM$G;Q$UG>
P9\0@=_OS.-YP286FOPJH7;K78(6XX CEU7&7; AVN=KX@3\ ZZ'-AX9A_A'1;((X
PV1:V%;!'B>("LFX"\!2W-12GFU!YU] V@/P#+,+LX#@V"<(EDSJF\H,G/1L=BI5W
P>(PZ6!.,Q/B 6KI_"QOETCV!,W#+ W>,X?IT6P2.7ZEGA;*])>^L"/++=GV7K[WF
PNB_FW*A?Q>;4V3TB$*Y?'IX <LI/<>^RZ\HB+V$4A<3E4\,4T'Y?:<QV*\>:M%>Y
P+2<M%+#**]2?9"-TM=B\ UI&"2WKS]HA.3%(B%R\ZQE;Q4FC:BQR<?KW%F'J T!=
P<FZN94ZC[6V)$ XU!JUXPX^5['U)JU1'% TJ]%"77X#,OHLDM:E'Y?9!#56W!LT8
P^0I?);9ADU1<8+VIOI!73R>N-G:]'2H5@N!BQC&TET].3%),3A)?2+PPW8 ?6!$X
PD]"23[)"*:^[>"8QBA:.C#_ '/K+JF[9T)BJ3I]O_XXE>U& !Y#/0=Y_6"C@5>K&
P9<5_A4^XZ)D-J4"+;%_G!>TQ&FA,2PX? 558J-<XVC.OF$J 2=\(&CU*^H3X!8FJ
P9;>-1J^ H @D!>$+=X<=ZNE;K$0D8?(%\,8BH>SG'VPJ0_U,><(U-^+<27=S5.MK
PC8;DKW(EPLD8&@SDOB"QF:]!YJ?@2OPD-DVAM6(\G',%Q@ER(:TY--!,,[8@<MM#
P_&(@<J+AI1 MDC=HU@.O<?2!KJ'HF&*<EOOB7_*5J)1BW4I56Z;.-^;@Q?RX,'5=
P4W:]J+P(15R/Z^K6D:T+GXNR6!*B7)$NE]Q36"8M2BC3$8\!MTN)G'YWD_3>C89+
P%AUBPW8:CAZRVT%;:8<GS.JTV*SL,\D\1)#H,1J:SR*VWL\LYA52,4!E5]<WPQL^
PMX]<$@VBH_S+7<Q,>IAKFW(O[1JQRV98?^W4._3N#ZOT9858?OG$MZ&VD"JIRQ"Y
P*[B!CVD*495B_ 2]-\<SLUA& TF8C5GTUF#B1@#7)DKB]"SIAN/TSD4ER36.V5&7
P..0ZJ566:,<2$Z]/"4!,24DJ;@BLR)# %J2KB=S;:!8+,'$J3SC>NN*=[99+6+2W
PS8;S(3=_J)C3=5F>*LAX+$U_G&]_R)Q:@++7PDGXHW J2MTR?X)0OJP<3081'U6E
PHTRDOKF6%K'"04GPNW^H7UL49:>3FZN"C8SIU\+4S[.R;8_DB/#HZ!(KRJX'7SG"
PJ9-6>-Q$1Q*JTL1/_L$D7#KGZP!TQL.QWO(*DEBILUP?HKH3]%E(=I)^IZ5$.8:P
PG_E;/+K^5^!)* ?Y#6JLKF"#1C(L:=LF(2%Z<T&<J8P/IW*&Q>QWU%VD K<%X<TL
PU& Y,@?/P)=3UD2 7^E]:C@8DQ09,1,@3?_3M)W-X4E.%MG6]<+=J!P[RA=P,TTF
P0&?##7 K12YLD2<B/T;Q>FS%KC,C8/I)R5\ G2%,GTE7QQFR>.5Q0-D$?!S+L1FZ
P/-BHC-]:&&AS/7PS_I2E'PC]@;C?C\!RV8Y72);MMYLN#.]FRZ__;+K#9^V&X,#[
PO-O5[4?RO"2!-0QPR**H]JNTD[OO,,&)U#G]]C%ZQ=(9J^FB./)PK_RE_>M$G[RG
P%[9V3DV0VY^F;&DH^XX@<JQ *J5K 8<'Y?_02CQF =];S&/EH%8(\3<-+(Z1KIAJ
P4M7YR5VE;Y9FS^V1="F 1L")^*=S3TW)_NE;YTDVM/'<*U%6&=GTQ,U-57V.!SF;
PPXJ;W(<>Y9;P@3B<(FB? M?C(ETGBOK1R[.GJ3T<[$+.SY:"$@B 7"B<7-*YG 5P
P^)@1B3;&T3N35O)I#@+\I(!^)RI^DR7=)J<S)C%:=32./K:G1I_-FO_:>8<I-#S/
P&^U52>_W8#?\(MG,P0SS@N>@Y0E54BORK-WMJJ1-:+WT7NYS%33"[)PG&.7+-9CS
PB:N5CK3'%+\*U?3U:<WZ($@-D'DS0:\]%;:Q2>0D"7AS*R#;%?]8-":L.>.7)1&K
P/K#&+(TAL@+%-[;*)^QU%J*,H.$$M>_^CQ&&PYBW[V&S_&/A=1S[?#5-,L)?-AL/
P#V.-_>&D;*IMZ/=A]"P'A&HG\S*M^>GGG],X,9M'H/CX>-CGQRB+C]M *+7V ^RN
PS/ B)MM97-AR."0OPE/A7GRENKWO$T(L'[N'AL -,Y^EOL+G(],F#6E5X^8I>4+V
P:0YZ.C9J/&^;C@B/]"\:\2CY3F;$OTRW81NY.#S2?Q;C/R A#%KKDL[8@>YQL :D
P3UH>(#O0<M!F"-@/VQ%/.:1-#80 (3RAE#E#O+=*)9OI(]Z50$.8Q C[#6LUQFS\
P0V7C^ K 9%0>CLORL26!D3'E'>;ZYWTQ /D '6[P7CE%C# >(P5VWI#B"D_4.$L&
PEUCJ3NA/7N(%M56\T'6@/GBS[K%0+6AV>^MJIBX; :Q9/^%2AE=6>UQ"(XR(/BRH
P=$F9BVRH_BXHQ??'EP@:>1$;\X6+K#/?C=' O@Y%^<#?M8F3URA'0&A^JZRKY+'(
PT=ZW9POR4.W/3TJC<9?6 A1^#95BG"KVRFDCQ;.1F=17-$RV+^:) 'P@'\3&;/LA
P'AQHZA<<Z%,GW':ZO1)< X#@FV$D_<)8XU]2V#U\,JU%AB;Q-2<[9NNDA!I6):% 
P^65UY<CYXFCUX Y1U#4FF:-=NH;7F&0TG6*]JOT&SR@N\KLUQ ;+L H''Y2^S!%#
P:TGL=B<*R2>1)_PP^R0"FCS $J!?Q!NP$--XK01Y!?YL#:ZRS4H/3H-SU(VNWTMW
P.J==.F-M_YV=]>#-.Q715C55/^^Z/&LQF8\#1_M>3@'0."Z=@"C4\6]!%K30*\3=
P5O<?ST7)-E5W_#C2 <<SID6(UBEZ>M%^4T+[!%,A ]'#:E.&X7PF^ZM8K?Q;] @W
PC>W.B\/G5U^O&-1IH:&=42V=K>N67.2Z9@F/XM0<%8:R3OOX_YB./JSC>V7(>^Z[
PN(@K]RIWS''90I3_/@M\<;'FTM<![@0?(#/B3XP'(@X[EPRP#$+,P0L:2]OW*?BM
PTCM'/4S+FI+4K#KX;<CFL6; G"-MWGV^F=)2R)>0(&AR)(P2)'80L !%R7,X<)4=
P>?U,-E^B2G> 5[V<0Q<T_2XTRVC/(.$)KMOSEM.,-CY<GX373+D_?[OJ7)!KLV-^
P#P\#[Y H=X106_2U!G4C\F5:MCQ &0^RZWM''$,K;,LK6]X+Q#J+R\S@]1&M$FFY
PD[30Z#ART#R\W\\J1WZ"=SSGJ1][61&1/B-X\SLC^J<@P:08=-0&J_=I?NY0P381
P+UZRG=O70IYG1YT*,&;(5@?SR D-3]$>82=AQV2VGC6'U>6)S+![^6NB$:9@94!X
P;7QXH3F6O.9I@@5-;O'A"DO0FI!D?+28@'U'JP)LQH,>/#FU)N^-9;U*6^-4.>5U
P#H7C]D!]]EH_B-D>G"8GT^L^CL.,;)Y+4,P)7V7DM5*UH6(&Y1P76QQO=VX3X=82
P.MR(9UX=NV XMW0'%R7"7&";:_B2#?4CMA[:T.3"N3E+2J3<CS8L3[?'YH1=%Q"O
PQM9-K%98>1-RV1"<?N;!"HA)S@N;S\3B?K60R-VXNM&[6:O9793\*P")S#197OW7
P^$FRG4/S*I"7,]!4#*<]<[5=!UJ>)6$>W9_T5;-^(!J_%T+/<H]IX_B2"8VP]%VB
P80<WLWHY'\!0;7AHM$R3@:],K,:>8YZ\7 8#N^7D#MA+V%JJ]L]\*>L387^^P/UG
P*./<Y4V-<"F+9'CH.)=_D2=!>?KHIR=T\DG7$?$GT6Y1&OGT(L5[ .WB$"9\5E#=
P&@,8</W'EYSF[EJ4;G\OYI5&\0N>1@X?M(WD_2PP5!"@L(&8<TWJ=+9?7@_@IU:-
PYRVM-T$7%U@E9T;9TA2,PRLZ-#10GRH2TTZT,@W*XU(PBI2@VZK"*<!JF!T82L (
P&%3NNL7[#!$V[ R<<9!OT"YK9<!("8&*7Q:&WYDE092?>?J9-Y(('<AVMT9<M7[]
PSK 3-8[50ZPX'[DQ,9!:O671X.UK3\](%;44D=G+#U/S-X\A;_:_@.BL,\A<R<=L
P[]^_CK'W-Y:G;]/R@J*_!+I*?*%0D-XX]2Y<;4F+SD$BX"(_S5"69?:>=[APBN1!
P,'98<&DS4N[#X6"-R[,,$2TD046 CY$IT#'#"MI#MC*I:$R(&>5JSKW[0OESCY:?
PW$G.*0<]T1KG.BZY7EYE$:C5)3_E[?4NI*T^!\A\"']]<,ZS_W>%9]"(?WIEXG+ 
P^]?JM/O[,)V_MB3"*U%\.N"57P5=&Y9UFBU9^MV7=7C&I'$(7G,FITF7@PUED#[U
PG;):%A;8J4"J"S$63  AW?S8_];E<<4W"UZQ&]?MNV!^X&FEDC3O?89\B@ 2OA?P
PZO<HJDPOK_-6L ?H2L! LM(5Z-X+(QN\LL L5W'7F'[#'T*X?*[.=).E<-$4N]@4
P^]9EXOTH49D\#C-L31DVN5NTZ2^>'>H@K>,= K+0I*&:,YPBF9.>#_?-5)(I2R4W
PBRNGH_P1?,H)W(UW3.86O##D\4$BW/"V#T0[.>J3XW0A\'PU%31^E?SYOD1TI1O8
P&^MP*T\N)!3\Y6J;VOY1TA/GIBRWB,G:K0<*^78]W_QMJF4EV'N.[U24/(B:6EA_
P;FKFL<A.YUJ$I*S55)\-?K#<$[QSM[C@(<SWU=3I''5FI1IC6B]$5HI*YCC( XSS
PC7E\9PPF3,2#@9Q&%WT@#2,XZWJ2LA&62QD^U:WD6/5^*O.;DW+CM@YP9&S25K\+
PK4S_AT3&+S!IB<PM<IQ:/CI:NP$JP**S.-^3^3\>:;4/DQU2I[S);FMGH&D.5L0=
PYG+]I\<=+CRGYQ*V:]8O!DH5S0GQ&]!4&G#)3!L&&)C,?_%RP.:PM1Q)EDKE&/@.
P-\ R:O)&"O9385[_JZ-$-4]MH"HZ%KPJCIJ.WGC.G00!Z_QJXZ,U8NZ]7;?&QC )
PS;!-I(+QIK[)IJ@F8MQ,?>7C>ET2H@L?)'!\2%CE4+[UFG5D7M3K,OH:R^9,[\]J
PS-8EPN7:ZU:$"&"Y_ B"^SY_/*AW+P E<;=%1XJSK :D 6;&SZ(!/NCJ;7(#7K]/
PQMU(NU>B8!3WQ_W(^\WV%Q7H1GL\T)4V@.,;_W6C<]\4OS'EGM7XH @9[M*56MTE
P\O+I, [_6NL4P9#X]L3]DUKUB#I%-&[(W]E1P&D:$?T,%0NT?8R(JI!UZ7; :"O[
P&30C%=[W/6_OB8DTXCJ[QWM0=1%E)% ]26Y&'HXGJOWXQV(P4N:;9[#ZX5SF9?FN
PM:NV@EU8M715X+V#2T4*.4R&0F;A LYL[,W#2MKN3DK%CX=D8"K,TA@8=6 /2QQL
PPI)MH](=0BYN^K_0[1J[J)F?WFA#$4U3Y7!Y<$QF%LF GT^"]ZNH#=[^A9.\3/J*
P93O5]V9R%6 L*5[1,7>^ _-EVPE)><>CD87XM_J@XSSK&>3+8'K6BVA#_TJ^8\V@
PX&,YJ;,]F"EM&IR3QX6CJZ[T&NT8U1T=BE:"HH<@=QNKZ3^04K7D/RC DP^F1^?&
PB[J@WHY4*TV!03<$-./(""G*(H#8BD#^_-D \W8)".M(?R<HVEPMFA6!1,O[3,+(
P5]]" *JH-,[*E,-GVG-74O9-B! Q;H+NK807J=\NQAFE[%2K.J/.5CYCY361&3N&
P1#3>J)KLSE%8-JB^Q3D.062Z%[.XUV3O2P-C%"8@"&WYI;PSG)TI-*DJ>P8O@;S.
PKYCM&41H<DX#PJM*Z4Z4<BU%X2'4.Y;) C(1;D([>,73-J/QIQ!5//4^9,D_&WM4
P92H;)+BBP*P4<N>4%FCG<[)]% J9)\GY_,Z7R1RWU,U](A@TQS'!Z$OM\T;?J&/)
PS>D@/WGPYAP?FR;]!!<6EFL6HFFKP^XK(9P.;.L?NBD.&V#W]+SL>O85>O3GH#+7
PAW)^'+.,8*%%';>>;*"4<23$NOW2:Y\I3$L[<24%@[F<:2M_?("SN52SYSFSJ)R*
PNGRG<DR_T\.O@U;+;5S_:EQQ,T?XMV:)1QJHU,1WCI$6,]_JYD9.;L.R)DIFJ2/M
P+;0VDT"GMXX("4M&D -;1:(4H52JM/]@/FAU1AIQU95$PL^+HNL:W6<L"^1UI>WZ
P&,A4-/F^'?//G<,OII@#,ZBJI*<,XDR$JH"'-]MP8H55@-YHN'R;2OZ2H&V>R,V[
P0@:#]KC1O1Z1K!2KK"UD] >C(SO ]+CVW[$L.+2_'2QH'0"%1FO7Z06508(<Q,9Y
PHB$ \.D@9D-.^P-N5R#I@8%-X:@?A6CIOW;?JOFZO-$XXE;; \96Z"D+?(6]2Z/I
P6BBM!6J6,LNWD[I:&8;95.Q?;''ES2?"&TC</SIV+>'W !I,3H!E<!4G.,>9*,ZT
P.502OHO?LP@DE_Z'L>[)/$@%H+P^>ZN#07$]?IM6.26&=F2R'%YT;Z:0FC*OT5RE
PU!H;W'WUH$RG3UY)<&/((=-R>.&_--8Y:$$D)GF@DI-[!,,FP8H^G3*BI*QZV:8%
P8])Z ):T?XQAY\D-<V%! 7&9@' 6@P>W-RNR[9$9O'U&%Q&@AH/R&YLYO(034D&-
PNC[UI !Z**'VH"5I.-VJ?Z(EV<VL7FT2H-B3GRRA6A1%0AW0FH#_YB2M 1[:IJ3S
PUP)C*)1I"4 =@10=T P1A"T5)]!]ZQ3&#&H1=431?+4"7UNZJJF9O\VQ0TF:)-_1
PQ89]GRGG+9S=* ?"6/90]:GPG$QE&>YVI 07/RKHX^UGN'LLV)[\^Q5DKWL6UGFF
P"Z<.3;#+M>O(6X ;>CS^AXBIG[I*F3=/P6?T'P,602L3HSN)& P4AHX&^BA[;U"J
PB(;\?L'P1H?F8K<9N\IJJ\\4+'D4R*^K&WV>8D/7BF-1:_893>2?S!<F8V&_!35K
P ?M:R\V))D'N;VM=1Z<3F2^WB&# $T^##7[W)![R[9D\\*% A?RNV$9>M97$LT9R
PKW+K*\ZQL%$)?Y/RZ#%][P\*T,K(6=*(AD".$QS1P(TYFU3VG"EOHA;8J<&'73 "
P,>M)JK2%ZU@B_Y--0?^LILKSAVE0!&%(L.3D0332:]7Z=2-^4(;_>8G[;P)Q$1!=
P/_]CZ?=4?')M!78/D&O<$(Q"J;$]^8<\2R*OM@R83"_C8G72UQV VRE1Y5!@AH%<
PXL/'$2T%EQ$Y%&10R#V3@RW@_@^?)-1X!00+J@=7Q!ELN:H5L!JZINT3Y?(?"&=A
P);,YJV['!W)#1^W$&&(J3U[_7]XD8%3G->W[:05M)3D$40,"6G@T?L<G-5JVMSHW
P]49NJDI5K]M,[=GO:>F>6_%!0MW@BC&GRTF0@[WM!<P801WE./GVI*'4F_$G/_E6
P@F\HFV^28A 6$C[W)K-%6#>[!_GX]VR1FMCNVW=M6$8)O^A'< LXW!S_,]=Z'/P&
PSK[<#L&]G_[S4)?GGD*$:W"Q2)=T8ZC3!/ OMX6Q/7HT)_P*H?6!/$]'9..<A/$@
PO[ (X<7LGSE![]:$7VYJ6WV;9?";DV>(R1178"![!0Q5JVHJOB>^!:@K<[X+@N_6
PLM<7M,OKY=[>[@*PK=27B@S#0!G]J,0M'LBQ9EYT+3=6D?NOH-"O^HD2XJE_1P=A
P.PY/7Y8_S.B,3I$?R.A:@GUF"[F$\HQBSX',?8/JOFZ0H5^HFSZ8P40WJFH?1PUB
PU6DS*>T,;?2(9#L30[-1"VE65TCL(.6,$-->Z$2P)^"!J!-+*ZP1D9J9][@\74A7
P!&(9<R+X$!H8FKX"<-_283%JD\1M*=PQ'3]NKQSB='!1^9,11KM5X,3:J50NOTTN
P?CPX=,RIAFGSBRY-C@^:[MP0*SA28[C9#'=(X_X#93/L/.P)4QPNK21R4C.>BP14
P.;)IQW]EWSZ_Z]8A$IE:DO1L.>L3!(FHEQ@J[MH<AG)?C,)4*L5EU;=(^ 3+EWSI
P=+5.DE4).=(=AR?]=#$I+3BI9I\(1C?AJI1#MN!68GE"*=>1]DJ:JD/:IS(R1_ES
P+NO"5FI">#WL6T4T\B\"HK(:>$@@0 ;@]^_OEBFLXCNF,IN<AKVM08B+189]62)P
P[Y.D07Y61H'0RG+RP91OYV]H^7QX4YWS2XZC!-IW\AVP3M*]ME=\4I3::CLFG I=
P1RI;,9IAT+A&4.4DU]JC4(CI.&7-<VM(01.FB86,%P_ZW+^RR.E7GR*J-T2/%)*@
PCY I??5:PU3-:4H!;F"?\[BR+;3^@:46L.MU>T'B],I&*:Z?&DX@/E)FM+"UJA-'
P?QRG]AY3%!WQ](KY"J2T1-#L3=0I//J[(H=BQF[3-UQ>(O:'LPZM0;;IK$3&0L$]
PW UJXU+KDS?D@/H,S;,8+I:[*60RK V*@.A+\;GK(PNTV]04(:%(C#&NOVKHM$[P
PECC/I);>Q!$[1GNL<_,<\ST? [ H(_%&9#1"=P>Z9O)SZ]Z[;%]]"6#I;'B<*H<S
P:J!9-I&VNLAX9:61J![PH)=*'4WZ$(>.2S0A=C5=$WIGCO%A)!:D!257/<2H[8,D
P,>M]^FJN5#J)G:A\S_1XFS??VP4N42LC'ODK-E(%IZ?C?Y N#D]<D48HBFTK/A["
PNFQ450OOGGY=%_OK7\D+:CTQ+='[,REN6P/M$W3MVWLCSJ\?&6OMR3/1%/WD-*1B
PM6ROU4*:"M^."J<^&A!YC0>(3O9_)%E,)MV77 3/@'7$C*M 6.44Z*I%;S]FG,28
P.RBL]M2\?&*.$1H9PMIWV5#F,1:&B+R0P@!U:3C;_HJ08PN6RS,7?/7"R&/IVE[S
PL88[&)CI)N:;TC\Z"9FX1IFTI-4TZI:7:T<ZK6B%5H3C_Q*77#IF<;.;)I3R;CS6
P]C][D"XKM-,-;>06!J7;D(BSXRA=$[3&NY&$:U7[>WH!E^.)%8)%!XY,,GSY=]YH
P'Z[/"SQ@BR-K'1_%U1A;X)-YS_@/>J-K).V7Q_;#(I])J(Z2[BNJ>QH^06^H'X/J
PB45*V!251+&@#TZ3%J OX4IX*#6\7KB8SW<"76X63K049'7<% X/S@!<&R%J@& S
`endprotected128

////////////////////////////////////////////////////////////////////////////////////////////////////////////


`protected128
PDU7H_H3X>>IRR,/N?KT7T<0-(GPPGNX7S)K2O6232&=Z/G(,-RG>ZRZJA ?<O-9I
PD!&DT(D#(YO2QL-LJ>1$X6>]N<\'IUB3. !?27BT=8:YBP#L40GHO\+)NG0)+%6Z
PL6=NG3X54/&A:-W;HF=H!Y/YI:1,NFMHZ \3 ?$\F>8<KG-5/JZM#08DY7!4(4+\
P5F%J'JH]J"9N-,A5!_UQUS*HK_"":[U?+,?@I"8^)<^4?+8MN2=0S4+VR'Z) ,+&
PK3L^,JLE>-J@/OJ_%S]U($N;.V+,//.7-Q2>R:=$B64M7_4CHHKRO[7"1(QI:0/R
PCY6'J?6SLQ]/ X^I0V!/9IM&^"7.PL#?N2Q_.*KZM^U+H3[JQ&_KS]=\3Q\6FNOW
P-R$F5+ZO4]@:;A\4-579*^I 5\FZ->V(SQQY@SGA<CR1^EAAH581Q0Y67G%4@,WN
P$) !(.6>Y(O)D)%;&0B?FTW[K:M,95^ ZV2R/-H./<%K0,,:V8 F2=^6G/&+EI ^
P[GX3.#!"+&7*GS%N&4)#VV+\8;Y)N99F_^_08/YK5<"-[UID+71&L<Q,G@A6WGVX
P<3&9>^*!\5 TPUTQ+J;1\ATJ0F8-)SL% 3<@$S'7F?R]\E_SQ8RNM_20UJF@JBC&
P]=EEB\:+"WLDMF01YM;,X$U=PE4:*JI$7+[W,AZV3;!#Y7TL7CC_H1IC)C"Y@IY/
P^,F%;%$=S0@<?:5AV3<]--%O7+@*S0(9$<ER$.C.5 5V9'QBODHQJF[, 05Q(KD:
P:W: =_#I,<'L6 Y)+^'39,Q9G^XARI'0&B041<7KXUTCRD)'T!-7#L59P3I\<P<W
PHS=]8I_"K9PT,LO!R;JB/:YS*W1<<I>151U* 7DJ.XSX.J+3<; #21:(MHKQK672
P*9J6'MH>90X,+S'-WD'V3>5FS,>')W:=!1H<W$6K'I*[8_/Y0"JLFNQL*2,C % <
P8@ SS12P?*RX0OT/=C'RG+>M=H-#(,"8X ^N14GUVFQ><7!&;I%<O7'R^4Q9Z)^'
PIS<3CH]N-@51U;)Y1/"7_/&)&SLQE?O&E4G2*\+ZSP[QOPZG]U3!D]-)!,\VH,Y$
P<.Y\Y1=D_+T0,>!2>"6A*CRZ"9YBTM.3=B.1I&1I>1"HJX":1J9T341X-+Z"F4 A
PY7$_[W-M\[WU'83'%P[G!7PX@Y23>0+NTIE*I,T*./BXWJJ5^>?L*9KW)_YLACX)
P3V@V$G\+S_'0L5:AZO2Y+%R23U3=/8G/G5YEW7H'UIZ_NX=^118[M0<AJGA8B9W+
PN5/Q:#-D2W5EL3PP:;+]\W)Y8HDX&U[7&G%2(IR@,F!W;EJL#^H<'E$@2'7+:?,P
P0^[0@E,^549YE(8S>5-A'WOK 27<EU0FEGV2D"4\"+^$^-+'(DX04O>.Q$$]9A_4
P.[OLF?,*FW1$;.)9A*MG95O-7,*/.S)R \'$^!K&FM8%/^^K^O'LOY_M?:!#R(;]
PEX9F(X1@/WB!-)'6JPD+@VE%A8I),SWI6>'Y_(OF[>5O)%E\G[\YL91FH0B? 5O*
P-#Y!4N "&I>(:+GZW,@;[1::%IP=?*-PS<Q()-WV;EAG.-V%O<*5=)P536Z9\-AH
P9'A\/GQE4JPXM.?L?A1O7&:T/F5[7;[A,1564CS+B=<:I$XE%CNDUV'MTTF ,=K%
PZ* [DKD.KLL7!:'!HZX0,#..0\)CM;-.Q5& DG2!YQ-D[O&O2Y?2G<8PAN94F*#[
P#RV^13:E^L 209^G2'Q1&CS%&UNV]FQN3$ #>P_ND$FVJPCQZQ7-FFU.F,).=ZVI
P$:1!_8G)\+,0KS.2FKEK(8RW@"'K0Z:7?/\G\G!R@9 ;?R<C&\]I4UYIXA6JRZK(
P/\^+/C?JY5PIY0 J\[TDEG [7IZ.9;9(DL]KV8';[:^\U9 AM0/@[QZB9.8L##VN
POQQ"H=_:0I3,M^+(9WAL,8X3&EGJ:T$UU5\2<L;1?R&W#EJ1ZFLM-T/Z8V:[+%P<
PRA  O=I_7T'"KVCN(?FT#DH ]>T,^PJ38A:2'O:MWOF X1%!1O<EWR8<IH&Y3$M%
PY#@LM-E%JS08CAPCX+UFSP$$KRR#[E)_7E&2EO3BT*'27-@;8,3RNCT.#X9H";:M
P3A-*),HCM!GMGV)M)VTL.LCF4"IO:V3T#-E]Q/;"#Y^'.Z]9MLOZ45JLM.WLROD\
P=9\G/WS&KQR2Z-U@VK?<7T*)Z6%B.O,G0D9KL#].GJCI>C@MQ@/HI(S__W1H+ F#
PL+ZUM<EC"\3.>#]Z7_V\?6W9*]D(AD,\%S!*HL@LJQ2+@?Z#H)Y/N/S]M:O==&%:
PMF=="Z(XY)8,F*:'N&-WUB@(?S8^?%B_CD;&W-E_/^8DRQ*BUW(\!E"*\)]0%'AA
P)@T@"L'MO?44"ES'W^H#MGS(+IK_SCM9RO!!#V[1[#X_=!I(JW]0$R!DM@J.WV"8
P_O3P8P!)_%84]&PW2J#L#HR-:ZOF4<\,::C:2P]NB;NJ[@Q1?)>;&GE<JW-[$D[8
PTWC_3F! &/0@'>Z35XS[3W?XYQKJ5\_!A:5J^9N*9MJ]L#XL:;*G:!O6.5P\.L?H
P[&>^@B%!!(KHX03)_<9B$)!SF@DX<3/1N6A SRGX&<+K.^"H6[O,4N&'",P;GZ"Q
PZT!KNX8SI3N!#V;K/)\K&24*3AO)]N47H'IF-F"&0>0,EIZD#8].SY;GJK'I[H.R
P1%W,<(E('4%*1)W8PM[CDNU$!\!@OGY^^B?'6./DF)5-K$-]B&XB7;9T)0U)GK<7
PG"=3_@F.W##(>WH^!9IR <S=D[+:&BE.RHHU[GQ,D0:&+@6N;8&0EBCM341H)_..
PE3!S2@=HXHG'>W;.BT."G<?O,R!J)*,MMR.-)&@M>#<$W.E&"4X%Q<$R[9Y^1D[0
P9[Q\66$4,NRZM6H.'WE;BJ3O4ZA+F/L/VCZ[(7@M:K-4=J&%$:]14ZOJJWHUX\]H
P[%Y]&I)3=@$KM>*/LR' ,T@:""/T\L&+_Y:'_<L+5K*1HCX5I[XK5!I)]?U+9)VN
P_9(>O=B]6V? 0<0D 9_]F,.8L1?8A!%%A8[22S76  D="J5>-<]_>IU$](52K.M$
PJA(F0@7_6&=4.[N=G"0_&'0.',6H,C:3'N5#)38(Q;:!'2A&RNEU6S]"\<JP.N3"
P:!SR&$U#CW-N8T47.CDI7MXR.'G=#53TZ4,T_WK5$$#-MIO$[!S*,ZZWLXUE*^@%
P2>J\=#E!Q_M33I=%OW!D-=OU$8LDR=-(?!\R'WW>T*4;-$Y/F)E=/.=IXJ70_GHQ
P\[X$$FS(""PP@W(O7SXIQ<!7-.7Q6A'IC5<2F+<A>R5_*KU!ZTT_1 51^%PW]2A4
PS#%CYL)\H?J]0PSD^)5G2R-TO954BBRTL<D<W>D5K-M=;'D:NP\!XFS4&5B-)C"G
P02Q VI[Z( YDZ8_]OOUWZPS'ST(A>5.8ACY2V6ZE\JTL-%@*B#/,$J[I=RK'/)5X
PF_L3?KK"^__.WQ@(;C.,6]X.MJC@*'35)P9=Z+_\STE ?DE"9-,TB]"?DN;GGL[A
PUKRO5L'J>)*V>=,P=MI!7\>^OA,4,GZK >A^9'0MPF[&9)H7Y5] @ I^G9B(W*J3
P'A^Y/U@MZ;APOPV"/8#"R+\@@LT3O<\IT&2?>>1+H)\>AE'I$5V1DBSX0M;1/URP
P:>S#K6[787=@/Z%DSB!^72/9\%D"[_,J)-8,QV5T6W01D=+G[:_5<:Q3?030-P]<
PFQ >4CWU>.-!\2^AVHUE$KZ;D?>QY:A3H]BB:(K$:KE#3-D60 >;IN3++[&%7G*6
PKV%W.G.$'H5+UST<K*V6X@U_6#Y071QW0TYEUBZ 2T$G"S06_-!^)5Z1I6W/UMR2
PQ\LY?;VNWGS\]Q?/BZMBG<PY\G:=DGV7'QF4:\Z((Q5F<O*'3+@B:(_BG=WK^<S4
P#@WZ/]"FY;T3"A]!CL/0U0U6!Y@>XLCTS\R\3B$XTT#5K>5"/D]J?S>FF17R*.9I
P&3-OROLL2@@<HN2."#$[$3WT#PGI&IA, LYHI>UHX>%>9=OI(I:=GCG;0Q&TY787
P^*,G9<YCF5@9ZZ TMI690#%\1$\5Y2@7FIUU=_(Z#:S)/1NU:+4APX[_FA9'XEIH
P<2;%0WO%!H'(Z[E><;Y@E>(ZZ[ L(@9) 6-K+7>GZI(.3HR^'?G0(>P,'([A/;0G
PW7R-U#$S>3%QE50G'H*@HVV3NLUJG0#3S]_+=%"-<S>AYIFDC+U.E]0_L[CL4NI;
P?[T&('I2E)/V I]%0!0@Y51(A]Z>Y%Y ]9+X[A(.OG0.@A+CZL5J4-_#,Y3W5/4>
P^1"-/1,7++\R,KH9E1\&VK,:G3NHHJRXDJ@')_"CA+RVI>HF^A?6X:3],\A(,#9G
P0V\7G DNL&S*J7K%=@#&9$,R'Y$)](K+PI7YW%!>LE?.UT>7(&^?N=J@T)*TY8BF
PHY9P!JZ$2#KIX<UFL+P&<8E&VB,6X7G0Y )P(#DJ*/CFW(^"E2&J_8,2;2H?4KY$
PI-C9?OVT!5 L"KHW(O]0(?^7J6<*^DR\UV#@R4EHWD .S[_D7;4?7?9V0TSIAH7K
PW%WV'H$32)/5I2=P_X.SSGR%0;:AN4/.**008P5Y_^A^)"1>>.FIX\=*_#QP5%?(
P39Y8)HZN'$M067(WU$X)G!%YO<U[!5>=@.&)27A^G8Y9MI7A_7CP<[1>D\,JSP-Y
P1F>Z/S>6G]RB2U ;>8@5GT27":Y4V<;V75SN0:C]30,2#X-V>U$(.W,4S>B0M? K
P? PG76/XS!I ]F43Y8I&&62D/)D!8*@#^H'*JF.(BVCUA)LXR>!EPS[^J?]S-[K=
PU2;\ JI-F)V.2)+#YF&%P3B5&&UUOCVD";]3?]-JE@6>&$HLGXT7*.(^*IIGFR*0
PD+^ZM$;3'#5%.@(+TLBL^OAE5,]#1GB$NS:$2O848MN@JI,&[\_7;]-&8L+4PJ+W
P6CXX=S1AM:'RJQ3%ZC=$.=_HKX=9Z*J0J.Q<VB_*N(M3GG^XJ6<BGP4GE49[BM5!
PTDT"R=>23#^V4(:#0ZD_Q_#VQ^J]%^AUX7&PL1"<%@/Y<>=5QL/.2@1:.+I!9!6_
P)9JJE0#?(P_W: F"D%K[-KN^<D_5X,A(#KL,_*RF9M6_ 4SPOT(TZS0$2C^.7;#O
P5J02K/1%ZO/&?28&Y5((F(")#28K&0HX76/S9<?(VL%,?H)\>_F3'Z,(PG6/!:#L
P:1.U\#?&;)S7UVUHAV!5%H):+H-4- 45Y&LIN8D@.]6=48CK]]&$ ZQMP1#HW-_P
P[C[ %Q8 G8L*31HF5.M'.)\&NA%UGD+G&*D.!U"+ "5%31!7FZE^*H/#?L1AZ]I(
P3!BG7@3.80K44VG)M+LUM[:Y("4&-PIR7>QH4:G#Q#21!G]-N?Q),_N@(Z .84YY
P3"<#M@676J+)])GL8)='91TF:PHV^&BCT.8))X70V_9--V:)((4&=\V,EIN;1!YS
PF*KGVC\_2V?W2XJ>(.O_H=N;!'OX:)5>52/@O(W#]Q*N8B!;$18$!O_ MLSG>J%+
PCP,$?A,?/6MPBG'U9>ICS^5_GR[/\_7\CTST$1BGNK*%Q0+[/5:^J^Z2K"*:#K5J
P=94;:L\VZW9>!P9!RON9,8'T"]=E$5O)7?5T!7+#B'EX02S1T9D8HQ=4)X40>[2L
P(?Z/>?X$A?LHDK0*-QJI\Y@N%0.W3Z_AZ8)R\F8HJV_NM#L?N_:1:JD")YRAJ8I_
POX+BB%9\G%W;\<B =M\.@Z\(D?-AU\'DH2_*8N#Q,T1 WJJ\3!MS>/F'41K6D739
P19J5AJ4/_CBSF7@!8K9V?=)V/!=[G(!'JXFWI*NC-7Z9@I4^3-5@T&'>C2L7-[ M
P@U*A2 ;A&39_H1'N:?;YD,CW3["= 7E+;EX\11=!E>,5A-]5:O8\<CRZS+!Q5'J;
P=K>A!JKM^XQK/2>P,"*.0=GEBPH76^F16AKH[5_6;2[IO;:O%WV!6;-C;D_Q3IT@
PQR\+5FR)8NA+%?]'#]KVR2@"_,A1>HEVZ@M"_UH[7CDD]EO7K,+^H-Z.-0Z3XG,F
P3D#A3AOM]OXGE!$"AV'5;O,<W.::I_YV)'CVQ7&RH:/\N?G+<B)^")+X@O_BX\2A
P,[ON,Y+*0/EI,@EA::AZC AFR5R2O5&9$KG2.BW.PPXIS__\NZ[+'18_J;HE-33*
P"8T+' ,"879"ZE<.,%"K1'3$8TR0^(Q1*+,YDC$^!QN)Q+"70IW,4U6,V3D\A0J*
P>\UX&J2[YGRW9F<R0P8+%AIDB))/["ZSB\4C+\D;\=8HX:K6+%O]4XWHY%J^68CT
P/+F!1.HJI^'Q^Y%F7I"@$\XI,#&JWL"R6F3VL4XTF?Z9E;.)NO_)R$VB7_LG@3QN
P# *Z1\7IRXJ/,/4E6G#H^#%:)N*=L/F]FA@J8=E,P+3VN@AHJR!G'6MSMPFE^_33
P&H0-VK+9<<$<61J%)BT^A-8,3=?? 5XB)NL=KU%44]W]L^4N:N]K*>)/\W&4"HS@
P[!.Y-W4;OW"VD&.@4J@"E-]Z2"M@-@>\F38$\$2>7M2'8$="%!XOZX742^V"!H9J
P@M6AFR,(]K'/8 J,6[M>SLLW<Y6-PLW=J8L%U_+5N'X ! G0N>.[GN)1G&40154+
PO0(LY$!QW9[H@D'(!OH [YF#5<H#O;C/";>EZ/!?V+S4KD11I_<SVK3OVW"G8LCO
P>][2,YF$]4&A>@7F/OZCXR-F@=%YK+HHHU;+69;1M78+=GEJ@+]4\50O&_-$13S(
PP$>$00NVUE7$Z/-.;:\8/[-ZX]D-@Z6*5>/0IGDFB=8<<A@,"%;STAQH%OC@&M.E
P!DP4^'@>/I E/:.0,51Y*?R@K@#%>8+N'9J$FQ]^)ON$D[7L(E]:.\./.A0678F2
P4NG9\BZV\(QL:P"I#1FVB,>%N#-6G[TE@*3TUMB7<0+*V"",G#]XB<L4MEDD)A\M
P0AY<<*]U9I[7(L)Y/\&UJ>R/9744]Z<VOO-[W)%&TCH+B)EU&7GQR1T)3"F>L.;T
P4Z$"%WPLZ5HJ L%@T\#Y92@59W 5VQ<LEN$R#8P^Q5E^-P7>=3.?_M6@/E^#I,('
P%CD%Q1"@1=,J@AK%>=36R_$>J1Q7KO\\SQCG'8,OGA^<A;N['JL 48<?7KH]GWW+
P*Z4 Y)CIT$-U,P_>9Z$S"=5/&'?(V$(<@0 [YZ:5_[QF\0<@\\R;HO[TS8_H(2H/
PS5/=$8R;B_MU[6G_'GVLZ'\G\XJO-8C8*4U2EO)T^A1UOLMFAO@XZKT :=DAO^/9
PC'Z)\SMT;(00\@^V2$$RU4K1E7/,F?:Q:?)OB Y90UD23B6&T&\UB5^!)":+'>6R
P<6MVOW &N<=AS5H0AS,;\Z]+;S-<++)5#,ICFR?)>H62.6J/B7R1CYPSTE;+70!B
P+\V ,-?,,X'@UC4F2\(N4 ,7\%*I^<)DR)D#P'FF ,_WHB%Q3-:P:VIW'^F&Y3PD
PD./V"J<5TS*P/3U<+*8O-\#VZ#>D.0)N5WZN5&)(S6]_<$;8B3P\,?2"6CELV5O:
P#=Y;#0GM\D5?<8*<DA#CZ=T9)8B)(CQI81Q?)O&<\23D:R5M7,YC;Y_\% 35:TR2
P[2#CX4QRF$+EF<;7<KGF9-5-/2D>E1L6ILCFB@QM]D!- ,>]6&@A@%A\P[C8D>[<
PXUUC"TEXDY&DXO)1)M1C2*MT>*NK[^0;P^YBT833<S7LJ Z4ZLW<&8W"RAD&CC8&
PE#B9>5Q:.L&^&/'$Y)_*A<DJ@H'+<9D]KA3GQ0> >&:9$7Q80(04ZH7M6!DL6_2W
P#J1N>>Q47S^0'+$".+=DZA$7Z>HK!QN+^68F]-^ZKX*,=]A?51QV':LN<OYF4C7D
P?QX>@U1>VX:I0=MB"7J,^>#)TG4L3_AUUG<XA*T*]&#>Y; 58*@UK'D[;R_(G25K
P[G$<"@ %]A[$5*<[DQGT@&W?'HHT6E#CS=C/I5P%S +_Y,Q)!:3#$1PNQ,=[^$SD
PF.ZL=.FMS@!6.1@^<Y$*B8*>P>_T?)ATJ0F/@C:05<3SKAEQ%_P*WHL&6$W,4GLI
P^?'RK76RU]DR+C+Z;I@.)""&M5N//N=:SJ<<Q5%A.<)59/DPT&=9)="DC)$>?&:_
PWXQGZD"8)_+1]TF,4PA$AI:DN<1>NR?-4;!WP2*/2SU;\HJ3U4);IS6L9[&/,U+C
P<K0Z(_17O;5#M'#>J1WYMH4#4R%@@6Y-P*GP,32D^6D>8.E^&FK7WULP >NR%+ES
P+%&)CN;U'<TQ86(<?6Y261.'5.7#T]XM\N4?@&W>K1K?PH"IJ,CU&H<V"XA^SC[B
PZS=)G'O]YVK'DLWQ1"&C^0HLB,!<;;"O^L0%Q%DB Q56G^A4)3])>.'C8*>6PF#3
PY&JJ_\MY8MKUDZ-";JU<,.W@/&I^+A]EH89/I CJ73K_KZ8ENKW14 +,W%,Z'@/2
P4Z*+AD-@*9!&91Y'AS==CM^F2)JK"):^^Y>8%6 UHD\>!":6W1.AL0O K$5^_1LX
P7Q<MUQ:[7ACFY?E!I$42F:)QZ=D7A*5J<4]*C'NY['FUT+H^P:(]B"AR"(1,=N4 
PE/=B'S@[<3;51^VGJ;O./TF S,]]#'%*.H"9,UY'B8;?-:+S[>5P@!S)NA+DB(<L
P!+YT6#HNL6<8>;7#QP;63U9^^]IJ9.RR4K#06(S]F$BB$)3J2X@I3F]"Z#R@JQ-*
PMR^SXX5^T++XN<5#&2U:?U)M",_+138GQO:9>:+0M4PLFR)18L$></,,91RI@;8J
P?1//M[/&ICY7E>S[FS9<<'P&3-XH/+(*TGS U[UHUV"!<5TQ$[66L5]"Q[V^VA'7
PWD\HRO8)'X,RPK4K9RTV)RC<HH:2>(P!3>_QGME[&)Z'%D\J#8 -.FKR%!-020T*
P+?8DPZP?0.SPF%BX?F,8"T>3*X#=DV3 VG'0>2"A[65::7@\[IG-3+ YQQTUNM>I
P=HK$*%SN_KT<L&&YS*<+(-TZ?VLHZ'KSQ)7@WN+#8L1!!GZF79C,0I*ZQDS%43U#
PDF#EC' A.'7D',UC/NES<54R05;T'"@<I!^C_A%^8]#*J98N>;(?>_].)8M*:,A"
P2+?35A2\3"JS4L*F92YNU^3;2FPED BEE&H4QH0?V-8_*\Q._N-&(,L;ZB3NQ0(=
P[46:K"4&B<*Q>_8L=#Y23ZZBHBH7X9!TR!'/A$^N%XN8B^*6@'QY+^(^Y]W8C=W4
P GXQL<V9DB=1%T\^G3G(*#F-;4!"S!P.49K1H%?V:^1@"2M2)DJ8\OVV$M>9U1?@
P[>^F56W=S96"GY_U*3)^F/T.5XZF?R('+H4GY]>5HK<J0(2&D-\J^-,6Z411A_LW
P'H9"2#(@=*=X40R5&&!W1F3-#]O%H09,"OHQF!)]'O=) A>LRPU[$<$4G,XLXGR_
P)PSH.7S$X\J-W8JP T"TOQ2<XR$:-,.HW;5Q^IO/D-T]L.#Z2.80\;LA(!.^V,P)
PD+E7)+?Q-6/+0?#4%&]F.2LI7+#-Q,4%V9T=X].[CYF'0[2LQF%5< &@UV63SKJH
PBTWU\A*/#0G"Y1;UYG-6SQS 9B;+%:PY!I8XEUJ;/+G,0EHKZ--6<\KUA_Q)/<P!
PMO)">2X3VIT%E7EW?_X/-H4U"*GS>89IN-J&S'R>)4/KC^?F ACB;D?+D.8=<WRM
P*N0JK-QC:BE?KUEP!RC$5AA7P#PBB0$9O&O7SH8O*:K4F=]-;/UE@IA2@U/!IYF?
P>$:$%-$E^,@@1+9P-$FN858#(;8^"MJDN7[L?OR$"^^;RQ[8C1JC(9HHU_VFXGV,
PY855G(G*T1Q<WW@#M_)V7V7"8*+))*K.8ZBVSGXA+EZ*$#JZQD9L9&"@]DI+5514
P5&C_70P5!O-0JC[G'KBK?OGWD6G5$5O8FH%:*@Q[Q&=KN&5]TM8.F052^](MWT8L
P%"K[>#I3N6FRG]W4Y-BB/9),,FPYZ#Z237LHRR'Y$GJC[EU7.P6]AHUL,N*S0M4(
PU=!GZ>'Z1*'3?(Q6R)=I"9VZ03-.97;SMT%^ENZ^85\BL7-()'J"Z :T%6I874)Y
P+Q=$1?#\N&M7";:__VNL$#?N0_@8DS?IZ.)=/'$9::@M^Z9-^ U&*>W_@;WUC%PM
P9V[R9[[3/,QG=@M WFL@;]:I/%I;AU\ 4X\8^$5'1(+UM[XNP6P.<NO(VS?.E4%K
P',+3+!:<:)F#'NBK(U8BB85OF-:?) PYY%[5X*=6&X1/;,=XE^.,#0K\0Y0_2I-L
PG_G=!RLDD>67C?P'!21K#^X%:BDF$3ERI=#:"XSOI+:7RD!!GI2 X9D M;VG8N=F
PL)$54G<:8,6RDY(N9H)M++W?OT1BP^J:];K@%I$>7;Q@!V(Q1Y2]P+[ZW!Y?W7%7
P0'FS@%=3\L8]KCB!^2CJ$U^9?EE=B_\M&8]X/=2@>DN[I/9$VI;4D*)"Q>OAY:&%
PT75E;&P77D8*[?-XU^7BQ5@.&CTN\:/_7T'^D6@6_^W;]P/H4(RJ[(1K=?TY@SU7
PGJL]*K(93E& I<6LZ5>06*P>3S.B^W3!A1.GS8)ZJ;4HL@S6]\:J@K;,[L5\WGIR
P)K*6$N#<'-!7 U]H@K>%%\$<:'T2D$+F54,&?S)&'2H&-K,2D:9!IS),ISH'3Z-K
PC]L[&E9+$6+-M_$]JHX'?3'#G(\P;XB-TLVR0,TMJ4 @*?VN\.BM[,9_K_J\>M\C
P%'D*F0[FYEC9K=&@'7Y)S3><@)N-\TSU.^IW@3.)ML=Q9$!51X#&JU4:5E2P/.#&
P N%H<"#&>TGR53V8DX_'T!G.&0UHH#O^9*QK3.:D@ET9C<8_G5MO-&+8RFG%)SKB
PYN1-?U6Q@/O3"Q/%KD5H+<?%+KB.3A!D-P^LC15/.I:U-I9,!!P'1N=V@TA* IO]
P%3J26V%K"&[/.#KTLZPP@06,L)MW,>UZQB2BG6JBQ#V1+WURGB"02W6M/("R.Z F
`endprotected128

////////////////////////////////////////////////////////////////////////////////////////////////////////////


`protected128
PDU7H_H3X>>IRR,/N?KT7T<0-(GPPGNX7S)K2O6232&=Z/G(,-RG>ZRZJA ?<O-9I
PD!&DT(D#(YO2QL-LJ>1$X8=PIGLX5Y0(/^+8< DY%26N4)54 2J"-[W7K7RD2!12
P3%WY=6!7N,^^[A/IN"VI'^7W\,(H'VG#C16' UR/@"P?<+HY3?_6&N;UK?F93CTD
P&W[?MNT*V!E5DV4@KD:.9K8Z)A0_(VT>8,VQ6/NV<W&<ZLJEF]?.:[*,3X$R-/M.
P1:F)LO;O-B+9L4&@06Z2H4H6C48!HR:FXYFCE.9Y7;#>;5K;!A9&_#@-_M'Q+^E]
P!5T$W@#L\T--37NF\]Y_Z/7\7*E0($32=:R/YF<OSW,'I<'DH"O.VG>^]>J-=>2O
P$<ML2^2@TY(3OQ(4G_&ZB,;,V!8N'L+/NTO3%._T=]L _'5$5:3M-.X1/A5600$\
P$FA/E_:K='.$O=^Z L5P5W7#X<-S'Y'#(8*?AU).$*=BSWY]<.3.:$2./V+2W&_6
PY$.MTIM'F37E!47+=C%R!.$O@.M@W6S8C'*F4]Z^C(>HU.RRB"6]Y[IK;.3&M#2P
P?!?=;7/YML*U02[#R:AFX>HK9UAC5GQI[GQ'EOOQ?ISACG(2M!Z"2BA9&5&M$J_E
PTHG+]QOR>I%G[D(MZ1X>M?G4?'CQA:Q>J0$8%EV8.Y^]"9F?5C"6"AXU(^#'1;LX
P]9[WS_[Z'39Q#)CR2V5@.35_=[/%:< GRA+=:XINS:+?+Y^KN&K(Z\<*1@I5U\L4
PO&'^T@]G/>(A<3T*&PFMA3E/5,.SH(7:<=U>++X0RTH)TM=2F+YR9THBSIHN@0#N
P(;X'#BFMAL;7._R;A2A2!O$X;$M'Z>5E*;2RUF%J @JVFEQJ#3]G&=Z$G>E\7P0T
P"E![IB!27-9H^%)M!D72&.D)OXYF/[95 56TA(;E37G9*Z;Q>?__I826NU@D^3EQ
PBF<RX-<GQ[R+1/=)4VF+4EP.ZW&=!2 K X@F-)XT>^"L)DKJT9411395Y!;D.;G+
PF%/,9\K$)K()YJ$V*")SF.-^RW'Q)BIFN^^D*"A5[D-Z)LY2A:S=1@V],1!3G3&P
P,(IM)<3Q,&PQRABE#.4RQC1J%"W6Q<5@-PW?]]HH(E*-=61Z6KXX]II)Z;,Z&\_$
P,6V.4E?TH.G!D,6J)KEZSB"8>C8_-5 TQMX75Z>D!3(S1V,K9KZ EG>/(>6QHU0I
P/NM#N3'A<#"YD3H;_0Y,3@2\:^&OS[GQBSH*,WHUF^L_#\5G.X-VEZ- [CE4P?5J
PZSV+!M@!K'Z0(HC(?:&XYB8)?4!/,*J:<8Q^:.N-.[1>\('9Z(-VO]/EJY=19Z*P
PQDS,*V;OS]MT0^^H20>V?">\H_>(;Y*0O"@JCY<5!OK.Y9: F![T")]9+$&J_?&B
P.XBIX.M2/&985@NJ4Y0:%.1Q$YW9K&3&NZQ!;JA''$R/ED[C&7K", AT H2"+[ET
P*'&T<1#_169\B(T,-N'W2ID]AXCF[/YVIZ(OSYII+03*?L4B&F&Y$=..1+C8+VBS
P=I/#4,X<M3_#G^LQC6W;.*1BA4+J%VN\\H84S,*'J(Y_,^L Z^,GQ5 (0-[<D!_\
P[[9<;AC2N:2% 5;YJXQ<<C!<*L4A@B/>ZT"*6J"J#ZP+A4_CC5K^YRQU?P9ZNOBL
P2"%K$VPWE%00\Z]AC/(2U\ M$."*;2+-_Z9B*V:/2B^)#>'1'1UQ[NSXS7CH@<S+
P"I;3C(1D^EEN8B5BD[;$;@Q7D@HX3CF,]-@U7O/A-\S5&WH=;E.[%NPC<4=<W"00
P3 ,L7W< 0B?646@L585^1#T-]?CZ_73QKI7+5 S"GR:_B".T]J?X@[3&_#,!X]][
PJW!2&+;/)$!0.!P;:H0?SF;>%B!T&#ZDA@24^/C/\^?1#833X$;)VJ-?*K[;URZ'
PP6PN1V.!SH0D'U05RHQ(<3K*68OW"$T9!7LR9M)DB^45INJ_ZW-H 2,>W0K#2R-"
PA"^,#>]=CV,ADEE7S<<!:S"E?[ NOH;N4B.5Z#&3#;DXZJ)KWL9'&"/'$-I4.9KT
PFK 93>@7 <*L+Q47^N>3?INK<<8-/&*<-TIE7H!2HQCW%<T^V1FUIG 5D.N^!NB:
PM/6?EWU$3:VL./)=3=.&S5;2[6BW$^)T"N8PJ2\:S\YV(!_&DA6);P!5]NNQ/IWH
P8@Q\==E;ZSIE-^Z0)X6XJ?/;F513,3/E0K+]JHHK@[KC?'D(A]!@$^A_(@)+%E"P
PVOC*A/GC! @-[,RAU;K[W8+P1:\D*5<@>JYSP_BR6GRU]2?AN9$*'5J XO(R_EPP
P>L@5*QU ;,9 JD3R+5-""OB8@$Y)-DJ,AG726[6QG(AKX9?)M,>X?___YD@3FOVP
PS\IX(Q'ER* ]?9R5+37"6Y1H+(46R3>S ]9G2U/]8+FU3S&6:6'[E$JI&9EL1\GT
P,Q 0(30S[[@VY#/>-W[L?##9PB<A*P]TPNE;+6/@_.#^V(LO[&A!00QG\\TE'NGX
PLW_<FK9(L52HLW/3R!\![6A9%0;8$+^N2S.,XV/=.;#X9,I$PG^$&II %!.'&W,B
P\:;@'.JO@N:O(%,I6-\Z,=] (_H4IB#2B..\VAW6@\Y#Z7FYA2_5I\,S>;F2?6 +
PSV<IIS\Q["#(,#Y]/>O=^VL#\%%)UH$3[4$ZL\?(&/:._F-48LZD 28-+0<@C0K"
P5Y @7='[8*.2:FQ:7S^&&&(Z)/ZB[XFI [7+9UR6F\3Z#FKRDWFPDTT5OD^V7\S]
P[G/5QOCZ(D&,JKG 0!1*!L=9SFR#,D*%@KYT44RMYFSLKD'2@Y(8,RN,NXT.#.\H
P#5]T;'>M;4(/D=;3W[XIXENPULAGZ:G7A7C4RD=/!F_::LX]XQ^6$W_.BNI'$*3;
P0C@?VH,(E3#";#HY>S>V7(".Z-<!H_^;_DLK2-742MR20B($C)P'<50[F-/A+5ZJ
PM\TBA4X0? UM]Q!"P&-.SW"=]+O;2FT9<95N? MGO?7HBZ72-E,*)!ZTHC,D;556
P<T:3>#>ADX""133=6V2',?XEQ$W]#MZ)[E [5G]]O'3(%"85B%<3L\A/]L,JYPZ!
PB+P.6GSVZ^!'PCDVNND_<E@N5),0DN.]J'^HG.I?4+[PQHGES#+X@9\3E\+ED)CB
P$I@6R"!.F\P;8W I9MZ*,^N(4UQ6SZ5&N.OZ&=%V/[^<WZ'J-MX/RKUXF_8KTXJ^
P+[S(8FS51^CK*$*@DO#HLC$HC;9,B]7'\'&/^&I8YWW%X5&P,X 4U.LP&TNS1 'M
PGX((>%G_4H8'R.$8;7B<0PCO;7\F(7_:G& X>##J#/6RKW'GNB[TW%NIO3H,0H_9
P3,S<N=&#-)W:#&W->*;>RP&H./?G/FYB+\IS^,<?_YV5B^>?L1#61I?B*#L76C?U
PZ\622W36)$")D"UVE[O19,J)?Z;[V?,ERS $=UH%^&B7H4AU''^5[TD074J55;&9
PW% [P4Q3Q=M8A2_#QG6ZOO2/2D<-[G%N) '%>B!RF,L6^&.''RSJ"$!I>T0HA\0+
PZ[V0A%Z[PK-%E7(@-J) KGK.;Z3-&^^3HRM [K@"N$.G^:/Y14\VP%=;I'%'TGZV
P,GMK!-HAYMY)$%U9BLAG>?E6T<I'C^2>LU]4[7R>3_^UFJMNBUNPL0_ CCP1LP>C
P:7_8.:I]DE&F.5;!!O*0CKRWT20T$2Z+RF_]?MFRB%>U=X_],9:485]PWI\?I18C
P=#7T:8+<-(,:8"00L+F*^7YY,?#NIGL]%F_]'5$4$P-)55T&FN S_#/2B1<>ACT?
PLM;<;K]3[TI)_>_@K^PN=\RVVVSK*$"6ER./$>/\1K3_YG)I.OZW<VI@]PO1_2,_
P=M_GM@2BPZ[#@GW/%+U2=@;QP<"SW"F0C/6+SIX"2WJ,@ANN6&[P[F[]:8[[W1_T
PNK[7W9JDQI?J+A@ ^ZQ/12VDHN6G@G<5GVX"/?YI8K>U&43]T9<?@OPN=WPO$%;5
PV;2[>).)B$'+X9EK:7) %KSG*,7"$#SW:=--IY[F<DW4& #WM-O'*^H.9,T=EBK/
PQ/ACE[L!O+;4/[<PE[HB.I,![(E_*7L]4ZR>,3%B);J(ML&^'$1UL"E>XE<U+@10
P5F-S:5#%[>/J\[EN]0'&E8;1BB0K+VF'&LOWT :C3#/!$55Y%RO9N[27)MCK,V3Q
P>N"TL+L_#E51D HX&MEHX_TN&4><"CN:4[$#^D2OU[2JY&+<PS*WY+JW<95&QB7[
P.*PC)LL!2\1S%"QI97M;6I_ /%>V-X*^@!)>DV<LG*TY9E@(_,9 NAHUD^?VKB1;
P+[9WYMIN9[N$A>/G: <L[)('8.<CY2VK[M\B6Q(5G>$M:,!1X0A.R:,^-'+(VK0)
P9&'G8X'FL<XYG'24_3#TBOV-^G0<M/Y?N<I]:VP I"RIKC1PHTHMHS0RS,@V0.%-
PJ0S<<(_$_(W^X+>\21RE98<TXG^V<:Z]!]Q$436^*5"L8K>*E@3D%)95B=']ATRZ
P#;H'>M)%7F+"987!N$SE(&^AE6)<#FXO\-RM#VKFLBUXVBF3FI@2OFV5]M%/[3?5
PTGH^9T0&K]]OV^9M\]V;&;KS-D(3^(;,JED,^)Y9Z,-]T<[&4).TE?TOW :OE5^/
PFGO*ZL C)>Q^;H M*<E&9,A/V=4BYW/%[_Y#;?H.5_^C%V0*<U?-P-)<1HOSN*E&
P6$JL\:)&ZL#KX79$&*W#YMW, >!_6Y:_N.8,XF2=P:U.0;;&V(>(Q2W!4BE0BQKJ
P@P\K1$S17.@[2CE9]2VGB>QQL)/_*([W$G?7][PN09DF XWA@+6GX&NOUI!C-Y:)
PY")>,T5TQ'36)2*["NO>Z(L)2E>JY+L('Z\PE:Z9,A9JUL)-? D\665NJKNHU*>!
P6T5<)BR=K@6?Y&:AIMK-YD)L1@M1+5Q"'IX@PQDC.=2%4&#S=R[" ?(%GV&%,W3Z
PA#="?J V?&0@SRN3I C9.R#PK<X#7D5_%;"88HJ )QD28NDLYJ+JM45A%!XDD8F0
PS1W/OY;%4Q/\?1WNX. 5<HA-/!FZ38FPPA W-M3D&<EHL>YEG"=8J!-Q.3RVU/F2
P4^TNGR%^=O):LQ_:_9\\/2PGNC@3_<U8R*[9MIJ@3NJ9M?439-GY]SQX.Y2Q3W+I
P47?R_?O*LI9M1V38 2 PH;6H4X_T2/S$;'0?55\4G;GKJ@K=&3)RF^N!\J2'Q/70
PNG0=J3 6I_JR&_Z#?8=Z0W_;%"_WQ!8#'?>/5I6U64Y;A9;/ZS> IGY\";:M/[08
P3[44:5];%?!\8)*Q O*R5*@>9@XPC1%**Z4#'&+",YB&QC)I42(K!/JO:'I=1WN+
P&G[D9S;J5W5=I&&P 2D5N*];*0>X7=?ZKL!SW44M,:(&?80=[ZJ!84'<\Z%A8A1.
PX8R#\".><AKWR:(\5@R$]G_T#M)'QZ:J)BMN?W'7K[>TKM_'10.^*EEF#%NV(7[>
P"+#4EQ%/RQ6+Z$]:XDVBZK=1SM3(KMZ>KJW?$.0S3Y=M27X^" B&.+6KKMD,RT#$
P>%)NU=#!_-!)>PMQ!T6:6OUT-,K&C>]TVF8 EIW#VO#=0Y358=M@L!\/6OH%4D)F
P.&$V%OON5M5Z*Q4OZ'GC^SV7^ZV#EB]*2=74?)Z5F+K+-&6JFB)5GSV7GG#4'27M
P8HYQX?S 7O1LS=K9U8R/IM0!%M-=TWY&=ILIUC5TU#G'.N49]GC7PP+0L --X@],
P<9YM';[6]WK^;Y!R ::-*$6":&]F*Z&V\H%F!K.TZ YLW?/(OG^UF1$-H'"SX+[3
P7NIS3V85T]T/$9QG"-.@E.2/I[9)KEXPNRC5>_Z)!+/59L/-IVT+,D[25TQY2HY6
PJX&64"'!>MS5]\;G7T\H]=*0G]8S<PV7EDT.B9B^7WD25)_KT0U(ZP&X!W;:EZ($
P@9Q <54=$D36F>C: \!KI'=MJA5!E;5F:@61F\H(@[>9AW73OXCR0QY[G\H &$*6
P];A@:],W@[L1"[8,&DC]OSM&&$+(2]0^^.?7QY,?F:12; )ZSL'CQ0'0J@ 0E8^S
PC/0!N#X\L2_9O,%Z*>IU&HD.;U$QILE=E%&,H*M/*OU'LK0O*P&-S2AJ5E&I@\C^
P5NW1,])$R);*^7O<*-8]IM8VV%9"^[*L[6 H$<SE9"O@"FB(>^C\;7"D_78;H?QZ
PW_+ON4T@7V@M\>O<7CIIM*-*O/W2K%$]9SV3A\<EE8C,KIETC"3SC!]%Y]P297ZS
PG5();1XD612"WH-Q42L"<" 4# 5@B+OCCO'9.4-DR632BD\Q)&S5IXTX,!#TR%^U
P$"%B F>/<#"DGZ-227\N#1J42*I\MFV6>FE8E\]]Y@,U,;UJK;4+@N+%KA]B!/6G
PFS7G"["#<^$SP-'J2!4[AJ#>^XE!6D-<?1!I[-!/$.[9@F.*;T435$\YOI*T<^PK
PE8-%43ZV^E36V]WT7\G=@2;LNNQMA:7S+?!_%CUI.*6]3V;L!*MJ,"EHL?BEE*A'
P_3M1V@V]\8Q$?RV]G73>F/X"!'65IZD?O-NRCV8/)BLJMZ&A #EGA>5>8&FM./1Y
P<5XM(9".D!U )XQB/S4@'6O%F). NU.R:K3$.&ZZ<\.-K/3RR.^9N^<NK5\=D/5K
PK3TW\VMFNW3K>!PEHLBA?;0CC)CJ\\*@^FE9']L"W1_>HBWEH&23!(]1DD K8 =Q
P]-1^Y8A 9O"DH6Q4BEN5G0ZA^+<1"3"%[4DPXM4$D^X(X=[]FK@ (QB.8V;^_S^H
P_53L9L/)AS/#99-*WB?)/#7LC/#9OO>P=! ^QI!7 1@IUG,?$[%?3KS@V4[])@(0
PK(!"%Z)PBN,$4W8N#X0Q"N&/9  VG09+;_^Q(=6U$EYQ05<[+R<^&1>^O_[D@[O?
P>T[Q;NR7AI^SKZPYH9)CQ^'GI>:$U,[HJ6Q%/$$BX)?-&,SYT!\F'0!]#!4^^I9B
P5X-<01[=F<R_(F<E.C"@A.YRXGO LBN_BY*CDN_"02W^.(>5DX52B-B&3P&_ZZ\]
P!/CL=%ZD)E<"L3%(,DI0K+R8#!-KPKJW(D0.7]XKJ2=5,.?T]'6;PYA6]EUKPK]W
P7[Y>2 %I0[.9NWMBS(Q[9&LS80NO;H.#;:,[%*FAKBOX2#+:#[+9,QAU"?[/^F'B
PG^/!\;X]%_&BC&TQC@>@C/^JP1)SXC+VUUYT[4%,"EM4L1/?_,N##E(=<G+;W)\$
P=2Q@%N^K*CELE3F/WP-H-$ YCZ>K'<H;FHOZR:89_2%($IK6HX)IOX6/8M_<5 0#
P6A^["/BUAW@W3R$/MD]6TB*:H!6T00#+@*#V^-$#Q#]X+8D[KO%CP84$*04:_H^0
PSSDY6DO][*ZC,&2)7G%QRJ"DX)EC@A)S'^_=X3GW.EK+?T6M?#-\/V7.\&L]4AZG
PHMJL-ES5)1L@+[DU=S#1PJ%Y\ZR%@'? 3%K*QW]?M4MPC&(+W3SR1@>@?&4Q?XKI
P?J 3L7GM?S3CA6INSP-WTA]?B?<+H3:[A^CFN<74H(;Y061T894-7S"\;\2_K>-G
P[5D'J*]Y3)VW_XLO=J 81TW/<+7.\/K_'K=O5/=W)-U,%XMZ^&B=9'<*WS=$XI=J
PQ("SF53IT4[8L#>NE%<)<$RNA&O)<PIU\((;P@/A%-85(L-)N'](1FPF@N8>0.S0
P7YI$WQAN)6)JZY2$*D/)NL1@ZC =:3S*L>B!5)A$S2OV-Q:L!M+35B)J[8P[;S!D
P[-X2 $4"-^F$BPI B750]VE]BTYU!@VSW?Z9L>JO^)^]Z]+^=& &B956>QV.96H+
P2*EGHU4E8,J?+%M?[J)QZ$C]X$%)<P^[9*0=GKGAO5Z1+]!%YR"!V1AN,S$RC#IO
P_A_WG;;7&^/GZ!\]XHT%8E*Z:._U^2IX)5CY7(3<[8A]3_J&].M[D)<]7\WNFM61
P!:-:M],EL)X;[Z84C,0,90D(U2!LPGBXTI^TA4$8D@K5^VG.ER4B@>JN17CB@PM=
PNPI$]PT,1\GOQ:3K*]Z+_3TQ0*,;E%!D-[]KSN@=>_:A?1G+A>=[Z6&>KG#;;1GZ
P'Z,Z('DMJ0B%;%T3(>7PC N09)$[AJ3"IJC6I2TO/MYQ3,D>D2<BQ3I&4IE+S)90
PS3'T9_5B&HC6 S3&I[<\MT[_HY):0!H1R,/[,$<OKI='T(\;Y0X5KU)6N/B8#%#,
P>>AF86Q#1FL(B2TBJ)ULS/+Y$PI\351/(8\,>:]?^YWB?3MHH_.>S1:(_'1BB0NY
P6(;P\?QEE^).UJ5C"EQTXK@/'5%W$%/ 8CLP]!]?!>65]4?BR+N' K]0@LM;#YMY
P2]MV7HN<*>/1I$ W"QCG?SE6AII@CT.H4_8! QXPRFN?XX7:XZN1(."),?:&+'K?
PA]#CE6B KFV:P@7W489BBSI!%PWEG*PU9-Y^*'7YA:]XCHXL?M4^FZ$@S%P/55R"
P,E57XI<!&2D\49 %'O#7!K\!MBSXHERTN@L/@:%_(WN.EM<1'M9#D#:F^=AHI&29
P]Q1-(W-0M4Z=4</$BGC;'_+GM->"KD0=\)-A35N3I7M/L_>SI;?*DTS!3NQOX9S>
P\0F<-;^KN7#K :P?M^ A>.7SG[H)C8&D_-AP(OQ3(9>D)-K^HN9.0LERS:E'YMND
P9"\BNG&>LO=AJG!K_I6E43T,'C0$.C"[*=_&WZHYQ^\.HX\2N!ZS+@M[QN5'C/U@
POZJF"2-;:P SFKE&7."0 O[UJ.RO6/NY&@,*HSWJJW&$969J7>75=-.@MD9FW_5R
PT4N)59P"IDT<&17R9?-G,8N=_166=L@_!*0\72MT8&!DIK]],NP4Q3%\:^N5EB__
P_AWOKB< DAMQAIXT%"K8%C?2G>F+BQ*%(\]3B1@OF[N,DN8>-=3R]9BR#L(TR)P 
P)V;>6[+]+_L@/[MJ7@R8^, C>W)/A8N&,DB8%]@4)HW+W7B @EO"EX4MG?$]C)Q0
PO0U8/R$ 3<C:UL8*21VN8(8KAS,I@C#B["W9N=)Z6WF!ZRTN].L>5_P:>PV5;U)Q
P3@\D@>-075@Z^Z1D=M9!TKW73*V5-#P7BP!1! *X4.8H)ZO<0!!COAL;DP:-NPHS
P.ZU!F\N"&CU?JJ=I*%X> LE&A65B.!?Q.$S?/Q:]UM$QS:'Y!F*9B!S?LXSB!8/-
P#R=[O$?3,-0@-5$\U\;IGKII-))E">@IO/FB5Z2%'HTMFL47VERYXEF;/XG",%%#
P,0L:C09PD2C"#(<$$C8#-B_.*<M)-$B3:8'%IVW**R1JC 6+YC0 '!^RI%G8H:5R
PRH?Q@KH=Y??SU&V1Q55U<M,;CDUE[]RJH;R:\\$OQ''PT8GFIX4;&A/K"7,"YAWM
P?4>\:<&9=-7#3UXUQ31C4"E.%!&)B]&=B^^7O@2.(DH+(,.+5D"4C%V".,T*=Q+G
P,:,Q GA;F';MV\!P2A)NGVE>F'J_4#Y7\06QCKA12%K""UMF=,+XS-EORU,1PHNL
P^.3#XXQ>YA&Z6+TQL^P!+Z9@:9723!X6BM7%3S^_C(I&074905.Z)V\+.;WJBRC,
P9IIY*4!JYU@$T%V!4JX<%< 34I%CB6IB"-Q>;V^9GBB>R6$+NHKE@PW3^492]*Z-
PH^#/$K2;._'G9[ZK$QZ0F>SRVG*H7R$QS^/A;4M0?+]^<^6JX7%.%.17NHKQ;:B3
PI+T+$0YM2WQJ7TEU6T,%T4W0&ZXZG(U_=3<NA_X]\I3]N6#M#ZAZY;:+S40E*'PX
PCF?- (G;TG*A8@EW.@(XCSVUR?J*3$6+B92\ ,QZ58,$<^T<Z;;\Z\@LZOSA+>"S
P"<L9N\N<P22:(^TY(H*JE-C@Q- PL)=>=NI. N->VL%/N3+PKWH %U\(Z]^R$RAM
P@1:4)YR9SE+>9U,3H&#_Q;XK,[ 8]A<.KSJE3N4(7?=?A,^4=IDR0:&KWSM/$MKQ
P&/UAR,O[@@;R'RL\%!W+4*L=D0HN-"9@S.UF^$#D)@'F.K7;*WV9XCH&T3MT$(8X
P>2Z]VB:4>F0@9P%8:<#O[O<&$J*1@MI+AER!"(#?H7(ULT'W-VE3ED<H6(B;1$GV
PB UQDQV5:K*,P2W>OH(Q%W,A0T4IL<QAP I3L0CE+4H>#F^4;HQ3[7($P>/.:$RX
PA-5EH"4,^I"=+TC(,Y\U3!_'-/5"4[9/M0.(9E F.([?=;::6D +*;$AU;IWU.&Z
PL=T[%FNULR^FD(@?&Y/:,EOQ8:.GST5=#^' KMU;:*84.5A.(Z5=>*<>Z235;%;F
PQ)*G5</ND5A<95,2MUX&G++[O/ IO( XN3P,A*M(4":W!!YNXS+%+'AEG$"EZ:ZA
PTQ!G\]7%@XF8I>I9-T EP<1Z8IGM]7OC&Z5MKS;K@3,*C5UBKATP^0^&Y#W<BA7J
PLC(^G@>'MO>(V;0#>N!4JWL/,])]*X[#,@D[;^YT&1/J#M_BFP=@KCJZ0*FYQN1@
PN_%9L:#PRMIC5LY3+6 >,YRKOYO0(\.=],*>M1TO[-1Q9=[]XVOXX\;(2:J=87JT
PDUT$UZO6K(#D>ZF"8@!\>:S"1SY?A.]9Z&D0(6DQWF?NOG1T(<WS!?-7F$D':Q "
PC,^.EKFU,JWK@:(;C>$;U [MHX"_;C0J%IWK4Y**%;;?D>&C\7VNL-H*.+T>:2@Z
P5*QP?*L#O)OT68[+T@\;]W'YU[PR+$9,GJM7$(D#[&FR(*UDHER?,630_?"&I:HT
P>G:%K*];?T80^,B3:+"(#F#MAFTMH(V%V@5:%3'0JL1,[U/$G8G Q-;/ME3O0 _1
PG(9=JB=2;3>F1-P%8MZ@$EK^W\@C,!6S0C35E?R9'Y95LI>PO-UFGPS6_<?HU\,-
P.E%\*FHP:GM'::AG]K3-ESVV6AD8G7"_G\38?ND_SFB#JJT)-G%&(.N-;X7.QBB;
P.Z '4D.FT/8=GP9\EE#07P-^#W?]SLZ1WEY/N)V.(3--[/8S"":2+V%,(8U,CB-F
PJ7>DW&H@##VHIW^-?F:D&CZC;FGF-;L](<H_\"ZZK9($_W/-1K=)QOB0B..OEL]I
PQF#SRQC?\ACX!U0V> P9%A7^Z8J_;OI4)-R&E9:MQ-#8EA-KUL6"T5>#A5ULK\\1
PSE2(K^R7?</C!?>_[C%=7X1_6,"I4@G<:+9&$. V[&76XXJ9WE&/Q'GKGE=4<0W$
PW55=?XU%9J0\.OD<G6K$-R$:]A&E!H8WI7/)+0&!@^J<;W)"#N@6]R^K#EQ.%82;
P='5@.CJ#V6AU\\2NMC>/HIYST'J/E24)FWO[YJ0[UW7MM=>3&>SN&R_JT^YY+R-/
P82K?27TE14F3!(VXNO%:LSOAL!E$.&VI03M:"'C?!)NHF?$\$[3J'85@7YO&D1*/
PTGR3:4'@XPX G\Y$"+_NJ*[0$WUF E+.ZDA,YB=*^9 ? #N)XENC2R@Q3:'0"]5O
PT'8#C\:\]"Q0;=LTI3VN=P)]-=36?]Q=7]UUUA)Y2ZNJD)3ZK.%]1O$HP(E2<';Z
PPGKR":6]76J7W&9G*\HRIXA!BN.Z-E&-21VSV*8.B,PG(:QEC#C \5S.=R)1#BV^
P@PVJ??V+4#C'-,GH\Q:L8#)N\887Q7-(/(C!/QXS$EZ$YB,8#3&9];KWV8FN7HM%
P64_@'H2*$/\;O&Q3[H31]D\NW)(8CL7)+^&,_7"V69%Q2P2>E@3YH_'C0U#;YK$X
PB*_'>CG+K%98C,U$41E">I+&_-YND]XN>V$WQD"-M)9R$YYB??8/AJ8Z!X<DBOZC
P+^R/&[VW"82P7_\RB39-*:^0M-CQ6*4SPEW/#.S/;&U'XGAZ_ UKJSZ?Q<S.(I%6
PR^N-\=HH!+<D^J'K;#IF^R'*N6/"HK.GS [.^7[Q+#GV.^X)\:!+\6NP8INF7]VO
P!W4LY+6/!\=W5O)ZBMD.IF3KM@F1-QGRC=M9F6*E&OU'^>_7HW&.3_ES(7B?D1<G
P^8,X8U[AC,TR%YWQTY^OZS&>?A5 [-?, 8M2*"S>Y',6Z8DV0S_ED)1SJZB1Q>OQ
PV+OU)I0'(=.;,>(CT9VQB/:%=%!9T^UVMNE7YV\Z$"=[)YFOJ,?,I4I1,95'Z?ZU
P^WI$ 0U2ALUI9(-1+O=B0[A!AA&@!6AP6/[@O(F&%TQ4\MKM8%O9:,+FAJ^N"HRW
PNK5C](Q3JWY;VZ!),4\2]LUR;0E5*K[AV!&\;>YJQ2TE%3X'UKD(GNUJ/Z;]W6>H
PX;WU?L0QN<(CI8>M(W5;^4X^*AN]:4^5+=N>H"XG3H=0\BCEC.]S;ES9',NJ^V!P
P5BZ\(LI;=<;HCWL,SYYQK,@U(08.^.A%DHNDSUS?-K%)*\1EZ;Q$0F6C__^O74&'
P;:*YWY^.;H1-S)9]FH1H8LJ1YOX;B"G6$-PI6)9$]*N)1Y]E;^H>@04[@[@2SJX+
P9Q0B[]TIF*$S1<LK>])(:P-LFF\(IT]UEGF!C3'@>SPKMB^B#WED%^1W4&8QEL_"
PT,[0&N%VJ5=1&^.&R_IBXP@*D*@LO&Y,9@:NK%@E5R[G7N$TIE-#8(CO.@O^> /I
PN452&O[2V/M &B+".2A]J:/&8--3AGWYN@D+(^:K63XL99PR5!X0*,\Z$QWO?=7 
PZ"&T?'%0]QQ31AMO](/INH]_:"(58!2(A^+%^(C;H75F]Y_E/L&E/@<2; TXOJD2
P[\@H5O4%^X,Y$ZE!,0;>WIM[B&S+&!>Y*4]Q&5[L:<PQ"5%FG$7VCO/'//J=+9MC
PXP*OC4ZAG7K&*\)&CY&'=G3&)6;GK0-^MUI;@,B4Z$>"U>D\!F;N!_J;DJ..\K,E
PFK&M(P@F( CR7#C\+GJ6R34^'7_1>"=&L"$MT]K@JC _2(0UC_ 6K_'ZIT\OLP7C
P[TT-*L&C!%VB^CK>&!RF/=\%SVC+5)XRENI.I1)F-I[W.,N-@Q>(X]I/PD/UV KR
P:0G<S%*.!ATS56=D.#MZT9.K_YP"]K4 07I;A3:]\:0LHS O@8#CJ.M\ W:%T_[A
P-(O.Y 3[!N?4,@N/GWJ=@3X$H+/V#W2\6-> UM;!7 .V-% ?0(<:(4/BU-#!CYD[
PFR$KS3%,DE^*W?DZR\:\VDCGOI3<"B+?[R@#0DQ"$\4:Q;7$T/7BGJBAE\I^NJVV
P*6I^R8LB_F*\ZYZ>5$&K7?T5J>Z FEZH9?P/P$7&'\F1OWEVT>(J2\"^0PX;-%$&
PY09I *&I#U3S)AMHJ?!D%L^>$29EQ*-E\(Y-ZYK:VN]@7^XRCK,SL.<E7D7%PJD8
P)R!_LCK 'Z3B*CV%!I+,SG UAKYWFSU?]B@IA\T%(B;@_79&S)L;@M+N"-#YQE2C
P?YPN#+N0Z?E.RL T.A^I$BXL&DS$B<J([JQC"T'U2S ^B.4]Z6V @_P,2<2%8:JY
P67"^H!&<J,F0-6T=>/0^/2K"JEN'U35V,)E\AQ >.ZJRP-. "9V+W"60:)5B"/R^
P5^$^R\E=7?6*()<N9R%ZD?;CY-Q=<J_N2\:L6^/H?,2O\>OUM^ %PUMRM/<M/#9)
P#UX<AZ.]+6V9#W2"V&9X2H#^2;+'NKKU-3D106>@?1/ "(0C[ /L!YR$F38!.%\,
PM5597':"^9;NAG6U4)^$VN?HA<O'%GULA""#>%MH(,C!AYH?XY61[!2DG4H6,FA-
PIX<^1_]:/GZ9C9S@A">Y'<@_)O1&,$+\:D8W$5R':)!?]K1+:]AB,&&2-=-L,XB.
P#0BZFP0VX1\WU;J?* X[M;44$?W+PNA/:3/&[]+&-M#J\&MA'G E5#GJOJN@JV.#
PIE#=E[XUT@>6QSS,+"\*7.*-K9[3^6#-'012.P;J1PS?2B0N,/#:H/G1GS9L),M4
P[,S:,7U3[@"7ZWW(,W@:!9WRP^Z<<0X7_69&2UZMQF&C!L)AW)6ED'^]-RW;4:2I
PJUJD,D$2D]V8U 3Q;H=I)QG/+8%?0TJ%]9L=Q8K": 4_#[S\C(_0B>JO:]=H')X4
PW"?2AXC*KGG4/FF7*Q@U[U2!QL#*;\EDL\HV6W:+9=EL/%7DRSX&\6NAQ3K'M[WF
PQ;(8UI.^*N?B<65?YKT$GP;Z09&3CQ?6AI6XJN*$-"]T[51>-.NV(O%7-5\;\RJX
P4=IW17JP2IX/^A]KI6V .?90#I!0V,#,U(^V;YG/VD/MHBXP=H5(Q?4T<2"YIR"E
PI'J%W%;J8\@YIIW\+@0&FDE;X2?_Z1:R;O&D[J_(\&JI23%-%@@IX/X5QA'C-&BS
P-I/ %60#/''9EH V6"J0&YH$X SR'>KY]FN;_U] ?0DH]7V)PWMPSHUI$CJ"%S+X
P=@4\:4*!3-M_[8==WW<ZR.3R,L/T=JF-!/*&Y!&! 0%V>HE;4UZO9)_BUN&9CRTK
P+RZI_<+8DD)]3%"%L$^]SVKX=]_*A3EDX!C1LOMP/ZRGUM^@&)ZSH_O[WZ)SGF.Z
P"7*$;G(E+=>SN68'[B<E?3JU:96A)JQQZ/AR6IX LFW+^*3A&U;9"B/NVT4KQ/)L
PG25/+>L<3B)@;JCDT>!S&<DR =Y7,:FJE9"[X1Y_R7Y@-Z0/6EI8"X;=D!L %T-4
P^8IUINWNY)ZD(FV)1SG.>:S:I-VB_PHZ (N>^ >6/%=Q/? E?%V!Z@O5__F2/YWT
PYOB3BF;,S(Z,;)(HYD45Z?5]]ITI7'DK^/C(3KW-)@5,1IA'C1]S_O_,'7ACJ2;8
P9F':9?792P>ZQ> ^AOU_N4X:P HEQ"TS:SW'T#M??V0\[B9M GRN:4/KFI75,.DQ
P2N3:*8ODDBTP",D*W'Z2L>'@XM(I$>B<DQ6PQH(65N65,K\V=P)?&<#N-^M!_]BY
P0(IB&Y&?D,4L[>O\;F8PCT5]9@:@^1+,5LC2,IO^%#TB@7?]S7KJ@D^'E53^*.%3
PAR--0/G7\0%1BB40)4*GGVBN$0E\\X(8E VFK92%JW.<@UE5<C<\Q1%)%2UTBR5C
P7E@F5_UCO.]P3^;,?.)84&X+($R)O! >7:LUD'RSP$/H :@"XFJTI>T;0%V./FRU
P%(C')H6&+G=:=D:VK$$S2+$ 9A2.6QL?6C*^\>\46DO8J5U>$<>HG-=,A ]9M?1>
P*4A^Z!CJ$<?/8O:X[ZB@Z6[\NOO7I]9^K),?4<8/Z-44N5I+1[;=F9,C-\B1&:EK
PG!OIEDP*8@Y<;%,YJ9R.4 >8)V@T.EH0%T(10'>1<W;5RIW"D*J_GB&ILV%*Q,WQ
P^$A;@<G7GI,]5H#X$1UNQ%WV!27&R"HFXD%#HK0A7%DM 4]7L;93_5^N1H4)<1;X
P9R0,4]OM.9!&A+A*W".^AA)GU+1!590._C;D,F*.%2#XLNSI$?*,!6X9#;4YG*WN
PS8C754:N^.2[H?L\X!Q8(W'M:X?PTS0Z-VNH8%_LS>B):P:3,EFE3LFH69P)>G?8
PNMC5 #?\&ZS.P5JP: P^-+DA^4,EJ79'Y=[,](Z?0H3,9-!Y!Q_4)8"B8Y=HB%$]
P:X7Q1"A3!*1D1U*8)'BA T2,LV&S=S:9_E[PIO,_V_MV9O=)%U_&[@.?_-*./,&D
P8(.TXOEN9J]A)'2/E4^#>5WX/)?W)XQ+EZL51\WH4?FG* A.U53-WPI*G2YK.K[D
PYIQY(?@V'YX-.-NY[LP1P*18?#'P9QIOME2 ;M7ARZ@X*9>?[GW25G)*(0$HV@LM
PC(<?+QEE%L!XC^GZ'-A-=)M&^5L1V5Y];\F8LTZ_==YBH4<Y8TP1%I3>%CR6_U8>
P;*%MS%V/&5/9]PQ;V$5U\&L)()*T7ZK_ Y"6BUXL7951CBH3B)U%%] "@._+T^ER
PEM:<AB!_S10>[YG;$O.]_PMA@A\-;YGE[!:DUGN:F(.CL0W06$1&^:*C$'.D7@8'
PDECRO#U)!C3(Y%Y4A.Y4IIE3\&^<J[KL''?,V,9>X4P%3I$^_PD_:^ZF3"DUUC,R
P3IX9E/-TJ1N#+=>'?KPX8TST4WPV:;#$0#]HMZ)\KN-*)L>#RK>NFOV$$]H[I\/*
PL"=UM3NE7XO>%4N!,+A@R%]/1,,B0GE%AL= +Y]FPM,T 7B]@.H49)[ZH,X@G,."
PG.3QHTIGY@J'>@,XT^%-C'^'_Q780Q(JF=XH#U5]^E=ZBYXP_M]0T85EONT)[=NJ
PQTD&IAP8F\9^@')P\9H5PFH;&H<G7;C_#9)NV6@D!AO5@A$NLV\OG3F"D3P>@J2X
P*#\8&@K[/]"N>9?KFLS62BS1.EOO C2$;TZR";_U9-B^*K4+$%6DQTH(66^!$<6W
P* ZDX+._Z]%@ZNX:'AA/[I<B151JWEP -RP++P?/D@'+RD;EH&-1(9IO":8]<.%D
PK=+X/+X9(#AN]TZ_7'(D_2<H.Y@8H7#V:4<8(H1"C#YL1IGF$&8639U'%#5(-+1R
P/;[RJ+34"UQB >7 F^813"?:./LU)-_MK%)SL]T<DMMD0F&3-EA\^KAXCQ6Q10L)
P@EAFXZJ RAU#Y,$K1'<(&YN"1EPMBQ%D6,?6PC,+)74.%I:6_EUZB#%)0VC<,[E3
P]\Y]U_- '8.H)HD_27]<#TQ=M9!4Q?UTHE9_-7<0,P%+B]A3A]3J@/29,.*SK\RF
PUE&B53]=^\6T1FGX&U%)\9'_'G?:#I,C.!V7A2_/9"^W5J)D;)N2/R..#*(0,WW%
P/FPP@P+3YE+GLWX<275UB;EURU;W5UM%3BN>[56\*TLJ"3]!XIE2=S XS)FVV/+D
P</(KW6B 1A;VK_(M;CU<@AR3,<"""V4!-H*JK7?>1JJ6G(\S!7-T]YV/B93FR5G*
PY+^]O\PE3N%T*?QY1<:F>[=5_*I-W]O=A,]^E&U(J*U86@L/]>UF1BY[[95C*$;\
P6.*OU54W1>V[QDI;4#89@I4+71'06Z@H7.))]&O*FPBQQZ0K@5U60=>ES_-!NY1V
P^7"RUHP,7P#$J()<U,P$=>=5UHUH;YW[,W,>6:_,89Y(V3J^$<1YJ!)L'D*F *OU
P99+.:4;'W!E1D#O$@K>K;=GM;Q>3C->/9A*7Q5R(#4K\F_GO= (,*G>E>TB#]3"(
P-RB]>-2\LGREK#> Z88^;;''^!4FOA!W'94(T[5M"A9/XR--  8\E4NL[LTTGQ)_
P@[TW-V R#G_Y]4O$,@"+TE4-2-T?B(7A@7@X["$61?^:>0<[6/)+)9"4,60-K;7N
P,Z)!<G:64B)J9EW2X_S*=*F+;\.'Q]8E7!U <%> ) A^G1JP 9I4J'MV[N07I)IY
PQ)&4O1%N(#3_H1\)1]LXBG,<9ONKA<;)NB=F>@,OEL#+Z3_,(@>%W49;!'XL6=L-
P7.57[2LR-2- @P68'F8^;OXJ<(1U_^4Y7!Z 2*OV%>?S"N2@=02]V \LQ[-7TBGS
P2GBU['B" 8E(2;\ /_.<(6MQ?D74%CMM(UX2;5U9(BB%-GDKI-!:&'5M@*S&\<1J
PUP"BT"XJ?9./0-!Q3;^\01L2(^LW&:4EI1_6C>?3\Q]+U&-@EH[A-^]DQF'HGMP_
P"_2"_V-;7.<REA\F/TX% XJ:O[6-.ZY%DOG#A8>JM4S>[GDD.L1;<V5% Z_#@I<B
P_96C%*[$^E;=AH/;.OC(7$=0ZI?VU@X3F:QPB"I1AIB:HO-[,.]NB8FB?*08*75C
P].^9&U)X/%T(@:!R=-+FTDTZ<O?:1J':WW2>NUX6>K:4R;!JX=-G/H2O1%-L+DX&
P^U"'RRB]UB5$'(L-#))4[OTR!-^,V,CAS09Q)*I2TDJV7/]9,_P/P#(!UV)5@V3O
P-H2IB^#])A*7/)A5:5?Q76O4D-IY'=?FACJOWNK=5PUT=*#7[_-?SN$U56LV[(T*
PGV;4*_:ZL&@VULZ<7U'8A@02"@W!&&6^5M$V$?U,DS_-U^:DF3]!D1B4*D#,SQ U
P%!DU]/UUT*[RE(<Y/[?K!W4D\X+_3(IDEY]: R)=(U<7I4Q3<?[W72UM-KXRV3RZ
P(?VP=S0W6[: HLVP-#QLYVF$K>B,HI%G'$$LY/4TQC/#%IA?T"3W%Y2!R$#T7,9[
P$*VD-JLINI]T SN!4FL,'9KN?;@$=136P 3*Z_M=X"C%SD9=:+"P>,7V:BW]J0=3
P9NWNZ<@>^:M/C&N^.Y-\*6?^2P'UB-0KWP-<OKA)_X/C^:!G?@7:?,5)%%F0ZD4F
PZ=.43R1R"UHD5IPJKP?1HP^1F)+R_*FK]2*1O$3[):4PD+*(&H#VQ! E/"0"_[]V
PDAQ+V*V,P-+@8BRQS>[/)Q$/<^F%D)P+$1,_4[H7T.9I=F2HSB92*8B[(*U;*K:+
PK%.\P\'GBUI*)Z>'/ +">2O"&FX^?Y [4<9*1MH3UG!+#0D8YHCQFG^"@G_PDJL?
P,8UMVJ.&9^:564ME+P(U"QW(35(-N#]F&464CS4(HMVMC82F@&Z6G:I(3$A-C^&1
P?P7P]0J!Y.D>L@#IX!SNH K^IMF;1!,N #JQ?LTD<Z3_2Z5DT?>Q+O'(Q$]!KLAK
PV@/7A>841+^GPQG%"TSH0'9\2X02QA4-]YE8H##'',#832GR>@,9'K.YQN./5]_V
P>  +@F0YR#Q[9WKX>"T)/C#1>E'6=B@GD+(4CJ8T))6/_GP\N8[=:N^)H3;9_"L^
P6JI)-#(T7ZILFV,=[3A*7[R?NB^DL+M 3/\6@4@JC$%/_+%&4RM7.6%X&.+.&"9<
PRK;="#7M'$"_()?>)0 ;<';LZW5<R!H  [9\< W"J:\&_.6/\!T6(4""42_=4IXS
P/*9?[2\N('DDS?!-21K3?I\>5OX+(+S2?77U DD+DH]_55D'O8N$(IN,LQ!*:%A#
P]%$! 4 \T.QA1>]/H0MO\&^,O%1SI\P6!&=U)XW!]#)?%^Z$MV-YV*AC^\PVSGX$
PP(5CNT45!0Z;E4,GW1SKE@>3K\2B>C/]XQ8=3WG\7[#?G!BZ9\(0%&.0YW5)[FHF
P@B&,*UJ&7-/S&5>@B^W2MC>#[:?=L*>50K(3?N+5\7'5L$MS$.?#@N$?)O-I2_.<
PG>O2=]?]DLV(6]89\;..3T)X.A #$IJ4;QV.E3M=9Y&=6B)]ZX%-:QUU\0J]BA1F
PY.UTI,ZY=C 3^JE;QC"M(PP0&D#_=TF?W5M4UL858?J2PMZ H)\U4]:#[(\)&I2;
PHG2+C5PLF'"W78'<?3J\+@L,[XV1<&A?5W]1&!:L,9/.J .8-JN^3J_19H?MVIH7
PA>.,J>AB9EY TP;>^:PK0YXWXQ63L0!YQ!P22#_C-TT_UA)!2,L[)>XTC5MLBM,C
P[ ?CJ("M/'?=P^E#M.ZD*RKSL):HMIG7;[4@;-,6%C#IQE3Z=YO2RCLF.[SK6^/J
PKRUFQ_\ZI.OT*N>;MZ]%VMEV& XH8 LGIZO1 <ZC^DCG:^=TA!'<<;0\Z$EB0F![
PZY"?[E8:=XTA<1-=6^7)V+KE<Q%G#9+UT/A1IS&N=!BLX+2&<>%B+Y_ U<)2A!LF
P18U:+N6D;+).D-MVB.#LWL3%.^2"Z/BCB>ESF)="S^0VD^N\*15[43L&ZN4#F1%X
P+%U+X>=O>KENX=3F9=4JPFLZN1>0+G "ZI8:HC CFAC&R,1TM\^ZY7=DJ?SXVY()
PTL(<5H6O1^\58O7Y9([NXH>OM\-LZ-"Z_O%E#%S^8:*CC?L#4W'-_WY^6\GBOX 7
P!(A@"JR7M%?]S73_NKN%36C(X+"O8!-E,72+2_Q.2V7GJ%8 )Q'],"I@43$58BK)
PMN].ILP5RYE">X_:SE$.1A:OU2H2(A";9TB9/5)3SI"A8\9';Q#@#,AZ,F<Z4929
PLKL0DX'R@O +81+$7S9$)AG6EWBAZ]KX42J@C^^NJ^Q4]G[_]:"$RK1IUSHF:P,L
PF;&T98QS.;"!0QY3AX 7@WQZ.)OTJ""O O<..'UXVR%_-^B81]4(%-"G[W0JE*]-
P7:EKPA?0:5G!Z[DWP;Q]S-KL^JBLDJOE"@],DI0V3O N 0>F[LI-(*]6PBM]J*@ 
P.CJ6)HRBG%V)U#)R/VD_WYCW%_&KJ[)R.=;\@.9C<*=;!9;BHU]V]W% DR[VF\S.
PT(F.1VZ]WF35Y<&7K]CI-NMQQDP-OZE[M?M )X)KN[WZ''J*FV8A1"<V$2/S<U3\
PQ\[34G9'4KW.ATQQ?<_XFUIPD^RX"!@GA4[IFIC:H.#1-R*RA$/5?-L])'6"&63[
PIMS;^?%_40V"F<J?CP"NMKI,692' *(9J<]I6B!@Q(<AG_'>0-4'U]+XN,*>OF7S
P@$QS#;/<C7K8Q.+8N9$X<=L57 <NUEX\$+S,E!C<OU 1H6^)-ZB.<'Q9:IS';/@>
PNY-7>/5AZ0@_S@"FY?V7$H*LWQ-@FL+1\/@# XDU-E3TRD7'!'.SEMFG.NO0M&O 
PK%"Z6IAQ-*A.IMX/]3P'0_'\PE2=:VV*NDH1*XYFR\9K6D2PCSV0)B""%B^/AMO1
P7G7]HX\"R<#$5PXZ*H/Q,554*X%RB ,&5$]N#M]ERD,4!]]./\7<6LPP090HU];Q
P:'_>#KF _!X>%H)]O\'*XJ.LEY AD_#W;%!CA#=LM!T7#LP2^VO*%L]@LV#"'RL5
P1YF:F9D3<!4%F["2F.@SPJ()2HYO""9F,;VN'[U$K*.LD_6\W$KPE ?6PU<JG5-G
P[6C<OKG<:.$%1$':@JF<$L83^5L%]C._8Y\@H^)O-O-_S:Q6D'=@-,RKS*L\V1$#
PV,@I'EZ[RX7)_&UR1E927)/VY09/ _G7!,JTH/2; N8B'C@\:M3D\^&T#X)=M2@R
PAW=M@\KM^('-&F9-QRS5;E-LP_1J(KTOW79)G&.='1,4D#23BX+4;T[EM;W+W*ZH
P_66F8T%\2C0[13SFZO>HJKFY>H TG1;>HH4C9$^.L6H<@SP 1#4;?[YZE-<O[&%1
P6=5QU@RVLB> S-!6D *NE$B#?"^0Z>FN& E3N2?!89=?'-MC)9:3?E"F62J6>!\D
P97'GZS8 X/GHKT9&!$M2_<D LA87%A,_XIK_IRS\!]ZHHZB06HWB?\_&#J?.I/_$
PE6I 73=1X,.$6K7>1:V* E4F'N4^?$+K9?2,Z-- LW];<Y56"%9]DTD8I_D^3N^.
P(O=)_\;P74J!O=C?M7!QA$Y1LU]M7IWL]9S/UU'I 6HU-)C!LH3.ONJ9D"(,FUI&
P_?LJ45G"H[%OYKD@),14S^S%X6;+U;OMTXHC^V4!?-@3N*:2RU[8+;_*T["1X(0"
PU5DP!9,4\P]2!:7O(T;N8IF%BC2=D5A(#U@1_J3,D&SE8]=U3OVN_/-DG[2C&&X?
P(QTDL-I3W!8(SFI>##Q9IN_!+7I=XYRK-+Q&(U2T1 MW!(^<I:!)LG_*T@7'U2^U
PT33ULN$4;+7I]9KVG@@>RZ.PREH$S0\U:5?<:?WS!3U?- R< -[."BFC@U.8378P
PUTB4TO#&\0D$@:7<V\ZMUXE;T3Z@5QJN_M![>RI95Y(4^BD+?&QD^%.I2A")1'&:
P4W/,U(*+WTEK;JD3!O="<<C-41/[]B]";6?B4,9/M'97_VMGIKFXYG4Z4=S!V&W?
P:R^2,:%540J*>'=!OI0T3%B<)F#X^RKAA*D)&*<'X<W.]*)7IJP2H<<M3_^L7]!<
PS]#7X%8V\4&&^)V==^+WKL-TR<7E4-<.B@^965O#X6)?'7XUOYD8Z%_J^TP9J!,+
P_.57"/_MD4[RYS@1Z)27D0H;+4=M.+,O>H'\I68W03-O,+IHW-_[\>"]V'0EN%CP
P?I_<C[22/ENO]=7:,G5_=N:QGXDZ(VB_N2.]$,A45;D-)8@S]2CA]?90;I&>3Q20
P(-(+@.'9JH>O:I<?/O8N&]>R]<U(_R'IV"U=1.\YPS?JXR]Y$, R54/:^JF(;,@-
PF6_7F=\,KHFJ74B4"[-]B?ASRN-OC-;8<(=OFVF,AYZ6_$_\GV[A6K=V]G<_/>1P
P8$B/6Q8^E.H'K+:!!,9LI3C\"MI*5DEV_#ZTYGH)-BS:(4<)HDE+",&>/%23RE46
P$QJ*,C@BJ/(%V 7%%9A]U+N^XKD%$-XG7<[*_N"J<3\X._>[UV)(1!VTDP'9U191
P.JZ/")BDNW_[7*7ML8A(PF4UFX+U.\9'T"G2Q9]W]Y,GK3(*$%Z<36[78.;6B1&"
PL4LHDT4/]UU_U?=C"MEG5<>W!;AV*H6Y>N%"E]Z5CF4A8 @RZ$4O139SNA%@.0-J
P,2JX?,;>_/):7+_F]V4)WE9OLA15V0OYH^Y,RT@:TO>S'&R]S+SG#2 ,\)J-D=40
P+:G[B#%VEICC6"3Y<E-.-P 5>WM.=7<^GGVML^SZ\)(41V6I)[,:==IEJ,=HID)N
PB>_\G2]85QP%/J\8*@LE'0V^7!L'*[=(YA:IJ3@Z"^^:>8B%7TV(':NW'"\W)+8)
P!0,\N[^JW>Q^C03'QCVE2$ *"?-VZ%YS]H=.[&R0DHS7EX\]@^QBBC&M RK@_5?9
PKZY-23AR7%H_JO9[#O8-KX8H.T^[6LZ:M$D.IF V5;'P7WHONYLYG0IN$@B$H/<Z
PO?'9#>T*:CXZPJ+OJ50HY)E5E@V*59Y:N_X_19;SLX"&(!9>L,5:?#CY9V[8>;>!
P5ZZ2]@?<K'&Y8%4+.0R.=<!;&4_NNOQ<L\H">"^U&QO/$&V8^J>PTEYCSI1508^%
PO!)Q_B(/JXYG]]*V7F/:+$STR]&I!?[$=QGOHA2E)),)WD\(VVKBA0= ]L+@[29F
P5YP'K@7@)<4FXHM=:XD]DAFTYV+2LXV+>_ Z9[BHG\3%<NOZ/!N)1Q!(YHS'3HMB
PZE[)\62;<NSPH+(D*5,M15LB2"+;43,M8T-I_P,(]I/<FD-4 N#R!U+VD-;K'YI$
P[3@*:4XZE8LWH/U)SL7, "));I6$Y!RFII+6D43VN?7['^WDK1#7V@%F5"Z0^O_3
PVE>P SZ^W_HIG0*MO(#@@ V$X$8P8^TL(>$(- UM/A>>/ YP2\<#45Q[+<12@AY+
P5(7LJN6_X/KY8'X=<<4Y%; ')^OF$J"!,?YOMRY;A2T&HNG:&@>B3*'56K\:VL^6
PMT7%1YI\FKR]<+<T8Q33VRQPV6QG ?PHNN.#45S5UL=Y1NX/V%!N3,[N.>;];'\G
PV$05D^.M<S(!GA_Y$;Q'5DW^5&]+ 0?X]UA1$7T\\&K5$,N_V;.<1]?*ME_"&Y2J
P-6CT#&><1.9W2#WH_UPG=*.+1Y(X$QM41)MOEW)P'6T^DB6#,'!1EA9;-E%%O;F\
P ?MT%[/=1;=1FHP"4X),Z_,B0_PSIJZ:=+N/L$I*X<CT7BQ+A:PEC^?^MC>39#U=
P#$GX)K-XA]Z2@O98C)4@_X\*/[]PD^]<$%\R)A:CB!/2:XDQO3;?[AXJ$54E)64/
P9H0<O5X^%N'KMC15A?!48#C_/D$P5Y@]=48?'&W^V4E:\0_8_)KGH3;'%Y"?Y%?(
P>^X:S1<6+X0N:&0LEG,_<<-4XD-8W8<BTEZ188SG.YO&)"JLOP^I/O+-,#T.80L 
PG2O>J'VI'JG%WR([6UK9PSL1B77C!-XTGL1,F4C'O,KKIL/'XP#788QTL.^+!)ZO
P*2F0T'(MO'!*NJ6MJ6OL.[JD@S[MD"X0W &QO);3R\&UP82J]X7"7=\^U\"O=9D0
PGK!2G^C #=YS1H7B= 7[*Y]'_]IE//\17-=#N8DRD04(416H-/1^ZIP\\W$CMF*N
PJ#(!YI.4+  >:WY7GT0EW?YARQ%>GX?!.&.*CE=9F^D#0(.^N'J7NI[52TOP^,.2
P 6:)-GVN<Z';Z3)Z;$.%E,I7-O G<8=(>[D S<^G]&0 5(<?EG@6I+:J3<I?<O:2
P;E6F=GK&^.0-#Q.D7+/R_G<@@:4W](E3H<6_/(9%"/1U$>K_BGSM![OK5N_AIH1^
P0F(W<=JKDM!R2+>WL C7A5" [OXL-KXH^%!Z"1>$F9L)FS&XFO#A/FXSBC[S]T6%
PY_E'D=^VW8DVR50&^-U!"H9O\947H61FKBM3Q+(#R^"NG $Z56%I]8Q2*X 60J,\
P+8;2I8[4P.JXRZ5=#6RGR32OJB,@%^'O"X#CCR;QQ1<SI+F9>.B%:/?D9S20<%;6
P4KCMBZ_?9,EIAA,D-.<698&TD[\O^A!C%YWU E[?0^VW<D<X.#ETW",BCDJ"5(^;
P5N,BE4%.IQ5X7:DL4"O0QTU<MTK$\?H)(Q-*_5OHWGXU)4!?Z[HO@B%K5Q+D9EVV
P!J#F&^SJ)N;Z#57"!1&J*TH]HH98II3G7_MK["_.$#I;,Q;NO5L;2#P!SJ 7O&Y]
P]+_A_']Q6U,[P<0U?;>V)\D%@30XYUGJ9IX&W0;/^^N2Q@/X4$VD<C:<:>.+!P8D
P>TN,,G[]KW BL:.[[KT,Y0+Y=:?%-J]!B30BA-N7(;4M#[>R2->I_A H3N07+W',
PZ16ZH$RH)J\)=N1US"3TDJ'.'YNL2&*3LM4/K^<7N=$.Y,Y A[AWE3"LAMF>B]4V
PL5P#LJ=\POU':8AP)D0*#])JR4],I= ]%,/EU@\))/^D.V(UGR/3)MI7/G%Z[&>.
PQ6GA5<X[2@_N\2_Y86FY=.:6F W U;W#2A"L-6\*H\!8F6(\<U6:#KYV^K0-W31!
P9V4\(I8*^>[F:?S 1"NEIW^,@?RLQ<=\-B99?@K=+.:4GH1VBJJ5F5$;F4EY=(QW
PG1\F5,Q9P?'+(O.5%4,)WW6V'_[??[K<R@1!N&,EFI$WT? #,\/L<Y_MR]B4NH88
P%;4TG]B$#F$6&SS>N2S1M;<$K\@0/TYI?XM>-9J*$K.%2$8H$25AQ^:<$^G6B!4_
P#E'!-3R=]CB'<W*MUYW/EKN'X+:9X#J"&X>"WB2:_4:W*_.3D-I'I'=@#PY0R0=:
PG684\Q)K 'IM,>Y)I5?PT\),&R (YF]0SOH.R1,>\2E.CW%&SO8!@_8GP%>Q)TJ;
PS9>4_ZC(K,A4%0#BT0U3>!80\CM<7V53MK#@+)0*-Z=%9&L0BG$H&5HM_EL<</ZN
PA+]&!:AS%R[/T4?#/ ?Z^(M>#F5!D:IJ5%5#:/T!X+FRAC-ES(4ZO'QE[9-MN3%W
P.O5#[X9F8H_Z4[/7R!; GPPH(UD/>!!%SE>8?_FX2(5SS7^OS(("#W>!'F@4N>I<
PRB9^A;!9.R+#YEE;)F*&!W(;I;3&@?I?*WDNC37SI:8JV05$WD2@6V^?D;F\&]49
PRW_TAB,9'L0D5^!1@B-O87?]:8RX2<8_P *AQRC\+6+_2!8'*=P\KW'DZAW:PIMD
PZ'P:&JT4U8:#WLI/FM7H[^.0ZV;P L@ARM(CUPEI]RR =,;F1M5$5=. XTV1BS*5
P>A8T-EF%JD^PY-AL*-B!(6@B(]E575'[\"H*>\9F:<V*RTT4."9=ZA2_N"UQGRIH
P>'TM85HJZD5\FMY*.WZ#"10>6YG$")Y 3N:'C:@AK908K4@,MV2:#'^VYZ_,5:F3
P^'9%9U;/)4T/@7]9%5_XD%L6]P&O$I[YRS?4OV0L33<2+73DP32:A]M"^6KY>MMT
P" I.PYB,?4D<K)2N_HCN3Y[ [=B?3[!QB!N6-!%7<A!C1B,KN*]+P&U1V]7%-I%P
PBS9Q?=?AS@I/70C8TP^KKOL?PJ_0&3"V5]#^;:<(?'-SS.(AJSQ+'()NIER*91V;
PTM/)RV\$G8YS-Q1MY\@7[N :;*!OCW?;[#U497OF,",??B_N,$,$5AIZU(?3Q>?\
P %L5-1 T^SR/>W.WG@)FFPVU.?;TVV\"@,"IA1B*U6J!1'G?)S5I[8]I6+3RU1(.
P4LK[W>Z@KCUE6X?N*,-+U+ HK=^PH#.4PU*DFS.2(J<Z"[=A,/' +)Q$P<IUERDI
P7H+=P?.V >^<Y7\10W*MHWZ(FN8?DY4NPMSH%[D 04WF6PYGW5N9Q38&Y32XQ)H1
PW-FPQJ&N#O\1>&O66SQY;1Q8V7JFF*YT))M!1?0$%6HX;,&Z!,LE_0J28#TS#DTU
P#R+[%-@$BN#94[O%3 Y<R.M%0WFG76R'J&Z[[[DW_*N1'JL2(8K SSC8 Y856KMN
P&87*Q)DEXAVJWB&E'E". 3B52!7@0<&@V-)1T8GT7=SSMKC&+P<"NGVYG%RJ<R:$
PZB;M%GN;0,+@M\8<U"E@:$2DNRTYEV8G"]FLB("<F\:5/E+5QWE-( @?40I58UZ&
P+!%#64H?&@Q&@(FK W4@JP7',6OUCW H#%]A;@Z_W4PI^B=DI*RL 8KF>Z+I:*3"
P(B(D'=P%8GM9U=;Y3G1XFDR?$#O'>6EQP(8@G+KW-!<'FS"D4R);:(XY($T,6C*P
PY8MQ["T&S1L[W3+*KNV$ARUA0IU)\G3C5J \AK5919V: B #9!L>WWPVFABQHB?J
P=PR6TPPV11J!4>WNHFME9:+^CMI*<Z, <L!=^O-18]4\NH?$0S%SR%<*U8 W !%)
PO0,9#%%3F)#EREWN!;&$BV\MA:JA\]-T"NB W$**M^NKFD'@^*5\&>;PN_/%-6O9
P@^6=Z6'6=Q\U?3%4TKB[1,;YW1 'ZO)&J/T2R38PB[G1EAW J/IV:V-F?H5:5SQ.
PI_QSSP"DU=,.O9JFVB?18$FH\&<'/<JM'F94;=!BTDM8*ZLE,,RHGM]&TL&9"*CO
P60(H<%,A*4?U^BNP@E$PZPY8FR&*0(["OV2UN1GI!I#@?\LZ->Q+-$[1=QFS3<T*
P!9E-5V&B3/-C2W3NQ"\Q-K\IH,96N?3C0&;21V2;E)EWNUU$6K;*<QG/DQX>9!=(
P=IY(0DK0%CM'J-E+7ZVDU\P/&T+!,Q&FZ3?:,/KZK>.#(+/@1/R?(>]&(\=1SYJ?
PV]%,A5NV\%6&I]N0[J#6^]#@<=)6D#+?)+Y,4F6[& 1=P9-F@SOK9(05<L_8$Y(N
PDS.M&?X5)F%B A+F"!$_AK$X(@RI:7AG:.A]&\FV6J'JY;MW:NI*;@O['Z;;Q12=
P]+?4Q&D',YWG^M#I;WR6&&+*4N ON^M_K>35D=3VG_?7!,ZF*D54"C@!Y7+-]-'_
PN=<+>4N]:ZLHWJJJ'.J>N 8H<.F-.:JBRGK?3/]O>:F1Y2:818AE2922 \^__Q(U
P?0[)5T=*5=00A@/6P'!)O[ =7)C^#:\V411KYUNAOC]3F7A%R*8LD-Z/;Q)V"_7"
P_/V^O\VG4BIU;%C-*%B-0A!2=X3,L'4$O:V,T."G'I;@KX+*KCLWNA7H^LM6_CJ*
P6VZB2-4NW ]B"F&<8?24'SM5X8W7_".=CHDVJ#-F$ @'T?M;_[P]GAY?]N*>T)'2
PU\P=WSW[L,+^6: .>E/<->ZEDV+ATB*T%WB@),#)+7AFIV^7$NX D*1^#S\^OH1S
P>S:U3:.1&+51+#$1W<FYFE'UH&R\V/RQY."DVH+P8'<9,8\Z0@''XL:QOT4[6*^'
P^[0*F4)#$A7\2#P2K(QBO.%['DH2*],#T&F\NAB.IPJI<"RDD-PYZZCHN5<@>4#K
P>ZW5 3Z.0M2PW_BV6OY,R_-D6<A8*._:=@BV[[=P?\?A4Z>T$[=%A(3KM<RB2#1?
P40& V;DM2MQ_!!ZXJ]DQ@NDGL6X%J5NQ,"FLZ"W2<;Y\S.%41,DB+2R/E]6("PW>
P:Y):L]FR"B \Z:54OTIFCLLB"5^('36A5^W%3YE-!:DR+T/&K1,#:?AN DII,>11
PC#C/HA%7I1\W?X*WZ. U.RU]Q@>-C'?-7I<WT93?:)1&3-W,[H(BP)#JTR20_#9$
P&3YKM\JT!N!AL=JI0V#CQ4H4@R!!.PUU*V1HV_1%V^QC^K#P7MC'Y83LR 9P$J.W
P0]4$^-,R68689PD2L',-::QODT$81AUDI[<&^V]M\6TW#)O//2/["^RT VR1NTY7
PC_)<IT4QX1T\7 M- T*S==S;TGS"SDPPI1_I(T.?5HO1<GQ(4_.P3T>LJ\ORT_V9
PCZ^ KZA_]ZN6>Y G(KWRPK-%7P<-0#M3^C^+44J/S+0X^M' C'Z(=(1PQFLDZ6P,
PE[GL^<B!@D@1$[97"2QRDDU'?]Q]!2-UE"[&66WQ6T$6NF5(>RLLKTN3'S]43-UF
P&#F6VC8^C&_4UB@V>LD/H0M]P!O@BE"[\<4JMR4CV02(\=CPVP3W<?4/&TI(9KB>
P5MGY[C&4"6BBOKT*'H@THPB9Q.#-/4W=9M9. H[5MBE3%L_>AU)+W+%IUY,,"/Y2
P&@0U(TN7GN_;MQ>5K7B=<US;G6N3XFCIAB;8:YKB"T8V6SX0V)8;PKXUKDQX/BE6
PAYD'&*:!QLT:]]K$CL[(\*3/8;DV^:Q%*EBRF2:5M[@MOU1H_!&EB7>N/TC&SIYR
PM-JGGZ7WVI8$TR-1:0UQ::E9?4JR\%["X!H]F_>O*%W,$I@'EW$]%KV<JK;P^^=+
P[83]_JP\]P6DU'C<XRMYXJ5UW=F\''PXUG\>%!O5DF-_YW74?]6G Y/V?PX#@N5Y
PW-QXD(2#*"-S#H5V,7W0>-*WO8A63*81- ;+'_A#=-=WGQ(B7(A 9*[U>S,CR276
PHJYO8]GN3X&(,+R]P7GBCY-H^H^ROR1U;-QOGLK[NHVV>H,VJYW#DP,P+ YAL;8"
P5HMR5Y4(0-OW).(5O(]6S9W8*7W%.(+6#DKA1QK\35&_*#2N+OBEN[3LCCN5 ,0@
P<5+2<KPU?3]'"6?(QX#G02P+9H$X2^(]CL@%;FGCR+;/#Z>5#$9Q(M!]+/MI2$,H
P$6;:B:3W->,*&:O-W67_ZKM'=8)$Z;+J@*W&X&GQ5R2DFXWHNT0AK6#E/R/M4*P9
P)SK.76E$[ A[&#/YC68U&I9(SI?V<Y0GQN,?%=^Q_0KV( V*QTQ.YN+[.VNH2%ST
P4(+J1E&VD-E2QYYA^']!44GSF'7&P'TJFD.>O%+L5%6H!JY54E^="U?'J7Z (=EB
PX&X'/:3;$"$&C"0V(>5LK.#&4,G7.[3]GUL<K&+J:I-M(.6L529!CD 5(BT#*[[]
P&0.*&3?D5NDU5B1R'JUW7&.53L0:?V,7J"TN8"C%!*G:>WF\ZSXG$EEF/A4AR=7^
PT^>^\WC 3<-7HU=:&'23UWSH83^UVEM_9,3;E9O6ZE'"BQM8M9D9%"D+#A@>@K#Y
P'#-#\9*_)VG[;+.CP+UGR2F$'O_GM=M^6>C9:71%_^DFDA8\AP73D-J_S__[G/UB
P>D/SX39-6.,O@-8J-08U)@"@T.(Z;5!EP^D,9+$ V_ ;G:9M,X&4VU;;SOF*) ,]
PX"\#C>W('T[H]M5</7_70_4HS\*Q<-YUU+U2TZC"'DGHFH+0X)+PBM5F;&5;\FX4
PE"#^'&$6(0K:H3L$'Z:C)^;&=PU_$W,SO!Y"WZCB3PMOCRQ,(K*016Z^L%CS1QZV
P^>B\@G?]X5G0&_^"!^,'(E\;5[\J:8EI2_P&]H-()<*1!+KMN\>N>RYY:BI3A>4M
PQN2UGVT(S7DVA6T=:/VSD]S.@ QTMRN,GCYQ%[#*>7Q;PG'RR#9J=N1%?XRR@G@C
P6<PKC:'0'CAF1S5V'XW-JG^ 37"2A4#I:)/P.]Y=>:Q1YN*,23]3VM')N:[22:45
P7:/ SLX4MC%$P]3UYR=ROR8J,HXW#5UX^Y]VL!I)]CGV2J!1Z:/8(QDEC0[I %2:
P0R6)_B6C1=4;<:@81)2JY3R8,QBQ'&CF>52O;*$D\EJF#PX98'NQ3_K+0P^#FDAG
P0P<F?K1?O@JYS6TIPN:_?@U/<N;R;?7S=^3*ZU4B33=H.7F2YE[;K#R"]TR!-)TO
PX?[VTS1C!+T0+M)5M(-Q$H92\JCDI/WV CFGC6?WPST/QC7N5BT=?8]Q[JB8ET]Q
PS1>CQU'EY(Q'VN/!8HL69!="<]&#V'ES$/1#^X_H@0:B6AFT%&H"PD"=%3Q_@")N
P /*  ,S*<=SSCU#;3!TAD-%6>M[G*X"L!=QO\B<R \TS;\S"U%=0)H[WEB)89M7E
P_LA4UT/,08W"H=M[L9XELE10JXKL)KO0.']=PS<!M=5'H'A']=*YHU#;ZZ5M\%P#
P7N14RR7S=EOL+\VHE.K;)8<+FUWE40+N1P,F\13-R_? 3)A:]F;V4V4CL^ 2VC+#
PQ 7,IJMGX?$LDV)B7L7DT\(DPWT;?NAW::F5:G-!AP89O< ';LQ&'?_7;G^2FMS&
P-Z",5H&Q!J SMLIB-./B?7S0\R<O5@JHPFL1L:NU--(O5;4F?OR=Q6,J2%8)8%Y/
PW9QS<"]DMD_\GE968BCHV(@DN: 19!1&A6CIOJ,J[:\M8^2&D%MT5F:XVD*I%WS3
P-M69HS&@=X$X3&P)"74XN4L[7@A*8_9_]U%;9X+Y?#UFD>PH\RX+V$2!I.L3*7K*
P:JU:N$GE%X2&JF9[#[%;D]=?,M!*!Q&7+["*9KE)U64F/>+0@/[H^B??L,N *_5%
P>\/6RN:UIGO\ZG;M O:/X%LV,\B\I/=*[SA@0+XCB'*\]M-Y#.U+4V=\/=S'S_%?
P!R[2MZ_]47,J =\ HR*(3,/1=1;7)8")?>6.I9DLEC:=?0%77[?HU>/B]SFHUWP,
PS+B%ZFP$/9+C!5 ,47\(3I%1BM$#V,)G\8OAX1JE16L5%,@1GZ,K%P$VC!)NC:Z4
PDBV[I%7'2I(A-W/F";:+:AU<.ZX*<#:50O+.1>VP:C=VGJ&#:825'W=[X,VC)5([
P6P);*9N(I7]8'2C$6WT^M0R*#?9=W)D" $N36R#PE++./ DD$XKN;:(TAK<2?*1K
P:1$]%_PT!=^U#TL:O[&'#K?];('S-ZU<"?B9/L%1-^C(\9B('V18SH@&J[J\8O/ 
P+W WP_NQ_,O22/E- T5U3E>*=YX'F8U3*!?/U\QA\4@1/I%4D5T9'K-F6J^VP.\9
P&9D.6XQPLY$6M^ZF9A2L$WPI>U'!.IED:;_\V86OF,,L5;Z4SAV%973[C^!<]Q8\
PTQBO^&H\4%)^^:+AG*.28G?F<Q),9:A0)3DJ-;U_64-$.DI6$D+?W@Z1987$=A(L
P_ "!A[,J\6$+K:1]/+ <G^'%M>%BDY-'_,\IUK5Z3KZE8GSX5U&,A$4@2+?RWY/"
PL?:4E:O<(@DDCF^/RX8\8NHBOC8SL?NVK*@>_9ZM<KPGTX.(\ VB!@7. "N93-'1
PU)"K]*_1"H8VM D3CGCC!#IEES !ININ@'.:RBB%N&'^!Z4O("0\;!ZG0:7C'K$A
P68=KIXQ3_9*5U'\CPRV&T9=.OQ(<V&CA%!79>)9'SF4$*">B"W@I\8^@&"WI<(!4
P^! N^) Y+"^6@QX"9(\ZI=CBS$0BR,]I'%D$%@[UXY[R!\$L4M#J9JKBV-0JN4[8
P)-P!BN.N"6S>U8=.AL/$$@M4UNV??Y@"7MG5*_#D,R_/.E)R(+;)H?YIS42%U74I
PWM.[:(_ R><J+9W;O"0YR5SFDG/8?)N.R/KKC@EF?/SM3AM JA7'R#!T-Z>,!G>E
PU4F5X#L@)QH]2^#B4J8=%<PI38P;9]9M12][3^PME'%5 1:-%N.D4#/['343^?'-
P8I(&O7!S\D/@[@O1_7S#?P<SDZ<2!GQ'.X-YO:^HQ% \ +GO;D/WDIB0,N:PQ1QF
PJ7.[1%[@&TVQ$(@+P1)(!()6.\[/6K!QA==3X:,F=D)+K^%/:]X3\B3C6 />IZ3F
PH+]6A9<B2AD@>Y>H@+LQH V\J(<YF]0'1>)Z4H3/USG@G_5%R3 7$L>O/^P4Y$0F
PG)WTV.CIZ/%K==^300M9'N11LD^Q.?QC1N=Z:M.,F.JQ!(_+T1;!GR)^A?,%DUX[
PI3GY"H,Y#X;RDZ67;+B6=,2"4XX/F@@#'?KK"<TQEDN]VQ=\H423Z'[2@M;\8^>*
PE#W@;R!^,(QC'.9;"J$0R="IK1#'YZ'U@"?$(G/DZP^..E!)*Q79.\69KFE<OU?0
P.P@N[O2@\.JY^YV;\O2>29 YY,=$+X<K(18+6D7,GW0ST& "CQ\-4GX,^A(][6AP
PI=D\NV8.,-VK1%UGL1/3[&E][[G6RER>&Y73;++GT@_B\4G2#GBC5)+;BI%5KY\=
P+J[&S&CTBNFRQP#V/A"DNK;<-N2D.QAAZE<6^/J_OTXJ8?H;WV+7J;+1KTS0VW_G
P3LUF0XV <?+!-\U:6"LP=W/H\"!M/U<ZH'>"B:UCF*IA?>HA/?>:SZ[FQ8KZ2%^&
P[[MU()V%T!T#;8F 3M;:E)#B)3>I4?UD/&DAR1AX4F2_&(<&3DZ:HL:9U?JR[W#R
PTL;.(?BI9)"D,FU.JR>MEMD4#52?(5V/CH=JS9_4>?\IDN8(P_ 8DT_M@2*@$7@5
P0\I?@HW9?SR$4M!,*$F_37@*V/"6U,/H?P"QC9(J_4'6XB659SHDY04Z@$@7,1B-
P4)BN%*>@N,L&'/@V*!'H8-:!,)*T."YR/@A/R$L_A[[.$#>]I\MS%(&SPE#MT/F&
P?/8+\CI7/EM4K2,[ZR?/W2?^=PWAU\1X1^#GF.X6V-1^T@>_Q=+X8?RA=</7)*+,
P/ :@J\'JZN!7HX%UP$1I1%3^:%[]=!Q)[K&F3.6Q!O<F95H$X5#R8)I]+?'WW_?#
PO;9M9SOS:UGDZ:9.*:B.J]Z486U,EPA(QZ7EQQP'2W\PO.D?_Y1VE+P49K^YK#\ 
P2W7W(Q:<J)7EI9F*^IF1)%3P$@]4EUE7%FZERJ*6X0J6SW2"WGKP(U7/4.Y)L(6M
P+[.%Q.@SW@"4*&M7L%"#+A#NN*W,UNC]XU6=HI&0!CBWUO*&%S#5GVR)#E"@+$I8
P]<9-?9XL(D_,\C!2@Y*8:!N#!+ZJ%^CRI7<DER9L*6(.E!D]FW7^JI;GS-3RZCQ9
PZ3JF.+EAWH-K/,>G0ZT%&(TQ5\5\$::NC"4O;J^:+C'8%=C@@FB2'7N/8GA;;XB_
P 8U9T]^+V5\;@M>NT3YJHS#FLQ=7I<_4OP-]J9))=[XGOW &;K?]J%:_#FK:]@$J
PF0YZAQO>E.[Q2C;=2.TE+YO"5R!UA$CW*"_[DVB\[:[$WXLWJ=._&#<-EHXIKP]E
P3;XOUX9'I+VG*LC,M;-7WF3J+@TOHR^HWHHL7Q3P+B?3J0#55'WLD(?GT5"V8!28
PF I@E$1G4:^9![M=AZ91N39BGA]LPY$DT*>0'./7D6#^[@TY0)U!EN/W,DTFT DU
P/!'L$R$!\N&]P9@/-*N+(^-U])?Z= RD,Q:Y:F\94YN_Y[.+'EY?%1@.6O7^X;4-
P]:".XM/!GK I]IM9##XG6>0?6>6A01IE3N5<X=2H&_-6.0S)^?VH&T9MA<Y=[?\C
P+?4S4*47M;5!?D3HU/9D):[@>&7^ E*]')I+M/AU_?#/?_%/Y%%(?>KLDA. [AGL
PG*Q@(GG'43_@$_?9J;8LBJ 49A06CF V_BU6%H3)NCQ:B*Q)BU X'0%.3A#@8JS,
PL6J&P?;^P6A._L4 ZH3#[V6V&)@H&[H0VLX,6/'Y8O[3PE&/(KX;STQ0,L.A'@CO
PTQ4^]+08+K06&,!UC7+F+=\1NIX2GL:DN,4#PM\]=&0Z*'\?@2Z1Y*^\16=XD19&
PT36,PJQ&?]!I'N&YH86+WLL9C46W3".>KNI7T[B7IN?6 T;,D0N;9%^%(1</1,XV
P]]$)" @B8.T 8KOC8^DFWIHKOWB=>U*TDIF"G/_K$@P*0Z!'E8>T/GM]FH!^7:\V
P1;)'V&_O 2EWJ\B^OPYO$<_AC8*QP1H@"YN^]5D 7AN>W>0E(ZHVBC]"96@4S9-V
P-\R> (-57M>QA;K[HZ'N,P2-!ICH5\1M76><DU<Q/-XA"*>%%' >+[]948IYWU_?
P?K^\FR[&[RIV[<*FST4P#PDB#NRPDVV35J)3UW=O;\?30+K8[XPPLG.>2XUB%)9:
PHRE#[H&H 4^WP:"80IQ%*?:+%H#$*/CE\\]J*0\#KJO3;F/-V0"1TJT1B':(MD9$
P-J+(U>6>N<('_YB-OK1Q3.!,T2#.EM8(D9+G,Z=,-B-^GTQ%A:=,(TH]V>&==X8I
PT).H]2E/T[%::=$0Q<@22 _SD9-$M<Z\]@Y>(@V(Y1H6K\CS7^0!0P6H_MNSRN(A
PG9D@H!]/H60;^NZW-1Y(UJ9!-)0C^9.01&N)YJ"NC2G%URA\@<23TU_"H?YZQ/+V
P_%B/% _+014BLLD!X@+A^>K=2]LZR:V^-&MI.JQC3+G1$0'%D"T3VV+,F2??)(&$
P[:H.N/_;-IS76V3'R$VH%L66-/IUD3I=,JH]-YU*LD5IFZ4\UV-KIH="*F O.F3\
PA4A!U"5-+U1GE)C$@>.YO5#4)  !P"K'VT"D5AF2HZ!>85NOJ%IN,1 ?-.P6S.!#
P5>>).#BA-52,HUZ:#A-PU@:Q:5VB*\SUBH!.@X7HID<O4<40J?>VA?'N@DD>_XUU
PL1P/%C>2-@M:VZ@JPPB2GW,_MC<ZRX U$W'U.V=F!ZP344U27& +MM>ZE B0N8I&
PN'_KNH"L;%A5_[9HWQ.@I U/,?,%-D!5TT%(<\;E%#C>1;>G[!Q+X&,I%!X7!S&9
P=9[H)0V(%11QN]S]MCXHWO$9_'KE(2(EP<(ZLG">6_;K3Z>#N[D]BWY9#PM$WT+W
PX\MO2_9D1.!5<,5CD,06(\3)>C'#YA?O^,I-D2\I+ .K'D#.+JQL5?I'CHLP.)6 
PXE;S>2&Q%=B2:*.[^O8Y,*KD);+F1!SSH_3!,EP 3Z1?E5"O>@L7:_2XY/MQH5((
P]/B-'GP\.OC6>>Q9_]+!UF!=PR((,[I/3TUI.&>(97>4;M<X=65_7U^]E:VHM\N>
P8RTSL"T.BDH?,/=\^IO>">S;D  ? LQWG9B"@HQ9IK'RLA>:?.>6P/B-9G,A_!N]
P0N2JG4C_PZFW+QW+4.^(O<B;=.'ZB^T(&Q_B8Y-5?5[\.MY+G8P);C-7M%AO,ID+
P"37=\F,8O"U LXAW+<8DL!T)/13XD 055B%/XC(#DJ@(IMEI/&.J_/%N,.2]A[R,
PEI+W]J9*XHOWG?7_:(8!!3DC2<$([9)D&P7=@_M\H1,J:U^_H^Q 12555-='Q.HM
P2ZZR:?\)_247.A\^ 5C$W<YXK!;)25,;C*]"3G';@Y49M<IO&<RXC=>2@<P>H'GN
P5K?76X0T6X.X&/0@6N,+7NGDK7LTB#B;3"\%@J..4]AO_NIWFP(G3H@5F\9 7+Q1
P"I)^L[W0*%$]D*??Q&K*?$F8PQ>^3NS*B1^ $^G[U,E/8C%-.X@')%,1R6;'$A:2
PI^H4%W?F":>@,*1*?[/DS0"57XZ*L50=IHGA3[EE,(;)CV1VQ7=&,T/CS93QS$,X
P#^-MYVF8^Y[B/PB8$#^$(A5P>X9J/ -MU>;^31!M3SJ/0961M$SBE5# 0_9ZZ/\,
P[K#W%R[U\O%4 "M;ADM<0;JI_9P7!Y=Z$WVF)B5,A##^2P$.O?Q%S@<6DR4E0W!.
P6'10/7ZFK!P#P=Z],*!GGQ'- 'H)<@EKO8WL>D.-:U\.QUD\(!8T\UXL4DI,']PD
P>JLR65.M.*#PV0Y3/PTP=<2_DOLM???A[*6Q;DHWUYO[%XYW-P0<'W+G%AUS0P04
P1();PCC".<.'P/TQ"O3L:LDT_EN>5E^RI_,__7T:\._1KK[&+G.#I"CE&_N9=)*+
PCW"E_B.Z[CD)2 4,\^9UY@&V,H'-U' CI:5.14O,IT$_7Q-%J.6QAK7TB;L=0;0=
P?TK?/WYX_?Y/(<+0G):QR7GD?PJYBPWOMK./TK8>& G5Z%^4@5K#V0-F-Q>[= 0A
PI",)YVXX+*HNWVUPEP0#89G!L&AV[_BAB&U>8'4(BEIH8=V+.^"XJKVETU9]7LPC
P1U$@/I)'EYZ1LX=M9]&-?26KJZV?&JA2,EFU4=3[5,[#B_C,72+%< :D&:$'/IK"
PM,)Z3T'T1;:Y!WL(%P'4R,P*JHVY#3\!Z8E:;I31IG:T\BP3';KQ=H]\/MP,M6?K
PI<1Z5$6'HDF>2#HBW#,2(T["=?Y5[V_H;2%R,^[29PZO21QG.6[(6Z'/_9#(\+@S
P6-X4G6ME-<*U5VLOISHU&G3VI#*EWRO(8MQAK28I"9L\%GM#'<-Z:2D[J%8?UBY)
P?Z>ZF#&IRNR]155(NGV37Y!5!CL$,FMGN%L!.OD[E1UE*T_4-8_^K$_8;'UR--&Q
PJ72"D3<'-&@Z0MHV%]+VZ9E_U\6T(32FCJ,[WOO*!I'Q:^^<6='1S]UU/#G\&9 R
P>T3^C6NIOJ5TMP1WIR7"Q20-RK0C]4)GOUK]^*M18;]_JUO-O:@_XJ@WO4%%";! 
PV'@R"V[D+ V*[#DA"U?BYG,R*) D%<UJ%\0D0Z87J?0*<_>0@VI$M%B&_T4RWIO7
PY_!$*Q0'+.HV5FT@S)5WHV@^&D<\P&5$"F@%GF9Y3\U=F,*JW\!K4LP-MC<W_)>0
P3#:U\2S] J6=[']=].&#X?+)H^MIUQ'T+[ =!F4]FU-U(HIT</ECT6?\W75^HG7G
P8;A></ WI)I(WKPBXV\LB")1+;E"L,)^;7?RO-P*)N=1A?7#2\CJ8JKOZ.LDV0*V
P#G@RQ4T':8O[_$S\"+C,GM4M)L(L:,K[%+W78P>>3<Y+OE6L9@[W:E5$&&$WW$H-
P7H=V>FMBML<5/AQ[^7:$@=L(JL%08'(/#_9VS\JPW!M>4N5:P#P?J]5,Y_2O]YQS
PG'J;>&P,E9JHS8RL1]]SF^D+$XY1688SH'J_.[&B!XR/PK*1#9.IP-] 0/3!MT(_
P12GD6))Q(0O9PJ%V+FH&)OUN(H8UK&HGQ!HBT^N5W4,D7HM74O$@M5L@6' +6LG*
PNC;YHTR(P3O_4VV <D55-*Z!/&RE_YT1>@$IW0^M4X#H^P5TZPP-O88ZB+JC$D%M
PGS='Z>#-FAJLM\__$9??,&>HTRP!/06%W<KCG67G#Z]=R,&')/ V\'WMEO9V26F)
P=FM%U'B%I0U",\L_I8!8_7L2[[G?K,;GI3\V$$[(2X$OJ$R<ITO$WG2J4BOY<6']
PD 7O[:*#Y;+H!9>F#HJOA;?YC-G=KYX%(D-&+;L!JMK32A&AU2WKF?4]QM)51ME!
P(=4AKGRY8@S-'F-.XR[6A2[AX>$%Q5A*ES(^0SPJK:C><5O$(,.M3$(5]FFR-^;,
PN0DN5=HV4(>^V(J)HNA]?1F*?V!4F&LO! @_T0RT9 FHM#MHZWWM![";,&9RX9D!
PO K+P,<JD:2W(S,RI$F_[ 3#OZSN=')T6+1.0B&+.RT)V#'%0UF@_,0:E)<!L\BJ
P N$\LL]'G5\7(IS[UNBV_$4)!5'\TK.T-@VL"<S0UO8"1R,&8H2X.FW]CWV4&=Q/
P(2=Z\TMRZ,)A'4<>:<QYZK5.QE3T/BF!FHH32YU?+[OJ]" XDR5 OJ@1J[\R1AY;
P2VB6U,1#G<?CPH@&8B9;QG\L//=DP5F".3GF5^3-X/5#X.O"SM<4W.JUA6_>5)QS
P6V4/.^=3;R<Z%E_+*)MHDP(&@%$EN?F#79ODY:80B&._+">1\Y/2F"*'X\U$L*D9
P@HE-Z9BH CB!M;&6W>?!1GL93O1U5*!)YJ^66IK$B+&,7^X63[]R M:![,;FF,0;
P&@J7 >Z# <20QF#S]G'?62@AH]F1$$WI-W:0DN$^@BC/1Y3SK2THZCCR!\"$/!&#
P;C32&>/^"C!9HOO\!F!&HX@96%H')*_1[AK%"DTW. U/A-/) _E?9=ISA@LYPZ'7
P?8L,/9BCH'29QTG&UC#C*Z.(7SV</]6=>S2@-^J'5+UG*U+&:B5^+VSR,LPN1>R9
P=#.E[U^[=([P6[V<-O_I*'Q,"_@M:'\\J+A.:-/N-=LOAE5(K(2=5A'B5>D17@K#
P%!A=T+%LPF-&*L\,IN5]'SZ-5J#@T!KKNDUQJX)0B W4)(I[-1@XS-?7[8>6B0TU
PH089W(?.<6TX5Y)8E5--=' -/-<01"]$D [6Z03;:^!J6^VD#7.YPWY+>4U;SAAU
P'NG1G*\3W*(+C3R-@-%VO-N5@</78<,BL/\JWAL_4$Q-3&*<K&G!>>0:]P-3)G4A
P-&_-M:;59CUDJ%N1 =_1"G]IP;:?>OW1DW*;:JRH^$NZ2'5+VO=[OHSH71KRHI*\
PY?ORK5"@5& US2]"D'>)X^AKBH1,NB;?TVUGPECJ\=Y\P=*B+?DW U]>MI*%U!(:
P@"E=X]Q]_<\&WND57Z_/[\FOPM#<.KJ_Z N%/4>HK=T&O/H#RJ(P4KVK[&<A.OA1
PS@<'.*1L3-U__$BVW5JDGA4R/].ZK@GDGCATN(O!F9\A\7V[&@J:BL:\[+?HKP["
P" 2MNR'43G"D.U(?!2<5.3N0.[DJ'1^B/A(P8P_Z&$_:] "Q*)MS1HXAMCB&0/:>
P)FG+L;63;U9G2)FXK9D0TLH3=ZZCA:B"Y&1AKS1I;!G.[- ;*S "<C@@N5;6.GIQ
P,<'%8&PRL[MRA9K7:Q0G=]].]P"_ (O<M[!B:6'<M.+HV@>8.@N:W?LD'OI(Q*KY
PNV7)TOJ;M'SA1]E2UA7)O7L^6?>-D_X1R\@:WR/]B;;%[R9@.B=;V?84QC\W6H8:
P8> >\[WJ'4*>NSKBC7-X8:LC=J:G@TCU;=?"0,15M$H>AC^ N=VILW(B\*ZZZ(8/
P]Q*)N [BUV]#[/ QI!Y@GQ.ZQC(3T]WK%P^C1M'9%:B 9KL,[E=FE^=5U6.%@ X?
PU:N;"Y?[5:<NH%>/X8SGE_?1VMS-VGT78=/ZGR 5T(J3]R1'Z6(O2!RJN*BNV5:4
P<BK*"S^'"VDJ89DGS3X ^83@T/>3Z4]G;]8YIHB0-&V/FUUH<)G/]46NL^;C-98=
P7\NNA%"YW(G!O4PR/0*B\+E&RZL-P)0B/:;A[OJ9\9,&CSH1N99:U8<_ ;'D4@9Q
P2!+_3?&;"IJ]0 V@\=BGDPU=F,+@=\'\#;4MOX\N;=37%1,VDTBJ6Q4?M(I/HAQC
P@0]G?>+#3=^8-[]P,8Y [YCP=_"#JFG4'N_(]LJ[US&U+9R+V$9-KPOT9&K%( Y=
P;!1SF+.)TSP!26JP]7VZ@ND*< NLPC=U,OF:;_Z%J 1UTZ^_5EP8P=Q1ZQ(XV.=-
PNUG]+[8_O0O4$IL$^I.NB!B/'$A]+1??LAH%7BQ4>F;^PP5_CBZ-'(].DF,[M]G(
P=@ <TAM&+FLBS"M+R7T1!S5MU#FN:;.D $#_:!-3"DEG'4:[QM;FU76:"81)9N%"
PHPPA3F8\&#JR6'AL/ [3U#=&XR)<QJ\P&^OBI#W7PC@U>[M?ZS%_@[X&CZ'+6;>=
P.GXE0.VAB9,L:?6O3?N \:8!@\+\MD-IKWXE#,_MR4A#>6@%$3 N]HW*(FLS:R(W
PA1+<4Z-Y@\%)(KW+O?PX.1:F; >N]R(W*FKD;BO27/X$E]=S?5X-C)F?_#$9]"KW
PK@6.+/@I+Q#<RP[>_-:^3]!&#PM50KUH<8?0C@@E$9;F+^UX_#U:!&MD3\8#OZNX
P6N^R-MP#&+9/:5M*K?9L^NGS+6*$.-$%V1(O"&53[!89&2VP'R(=O5NTUUR0ALLW
P@"@R<RU]J(74>K9.CG*?I%C@)/;&0:CL..OODUF\<4''L9"MV3""+,FU;9]:3)TT
P3VYFC,W+ B?<!3J  EO^V<QN8*IZ,G"?<6HR83;XEPHHIY3<9]B<EM6!: FAY=[-
P1L*W+PH>."U_=<-<*O+V:%$YZ5^G\;R\*,Q%D]>5E:S&7O0\]UA6S*<<V/&-40L;
P"2J%1=:C:,=.USYD1L68,O3+CU6VI_C$1?);_ZX>+C,S7HQA756A@^A](D'/6/?;
PL,$L9KJ<9+.OH>>_D3U\1M:!NEH_9]G8YK[ FTW.3,58!76X[!AS;7*M_7<SBB/+
P"9-%G_E82],3$&&">(>8D:J\7;_\P8:OBH2%A][BO$<72?=T@)YG!_!]^L\WKP2H
P/NZ&L6ESUFPV ,&G]T6+.T*TFX!L6$ 'J7:$A]ILT6D"E:"[2J $9))C-P/J/:6<
P?8(.4E?J[6=Z$6 ;65LL^W2+>PLVF?%?[CZZS*?.A9)T. I!B,SD$K(OU0(&A4@J
POMYU/E0-7+*?#C1B:$X.*0$R-!1RR8WC#88%Y&O<=JI#%>$3#1PX+L9@$AZR-2],
PR[3.FB4A WY-<74QF?=L]?$$Y/.;M3X UO!H3!_#I4YFX@O,V,\5M<VTC5?H)Q-'
P0X61V"V^YQ%LCHOSW%>G1)-3&YF\\'*3ZR_';^]F)5!^5&,-VB&!C"S+?7-+\U"6
PF?D>>YZ3'U_)Z*NAN^;J'24Z0*^3KTVF#")$(#4$]/?-'UM.VV@UX-S4UD-?MY(M
P^LN[\Y9UI'DK$70Z\U-^?H0# ==[<^$K^<9L%;Z:"9F]Z[WT8-7T-Z]P4%K4Q'UF
P* ,"=$7NM8UJC:!#\5L^M35$:.USKUZQLZKG*%*,8BWFWX9V>SK(IO>FI#"Q= %N
PL-IW3@M3J(K,^H\*<&\)_$]-DP.QU2!6,9/HLR2R@CC:?DZ[(I^[-9K3-0&>SI/J
PO@PG#Q\Q12VC:7&[<BLT,Z[Z_UX#.":F]7<GE:!70I$7<!?8&/+D,ZXF\MRNBJ/8
PO.ZZ[+B8T1W2\NR#=*/0A,IH'(L")U=6-_V;XO#!H[4_?>Q6/JN1C&P O:P;=POE
P'0P+A-P0YU&TY-M).845G:H@7'"V9QM?J=$I$EX$8$%SO0OLT]**7<KF6[4BQS,@
P@AIZOIOM=4NT6Z=4(Y6D):&3G#DG@JL>%W\8XTE2AVY7 "P'#";,0]$SBRK#+4LP
P"*!+GRH(. !9VE0*;M-6W [C'YPH=A,9A$SZYKRI7V@J96 ;ZN10"6@S&,%LI&T_
P<8(GDH=/-E\R5A4/ *TF/E[3-8% (0=77S'5R8J[2?=/];(XJ"&)\4[\M- QW\G!
PEX'F&(E9R&X<.K@HSWS2C# Y'J(V[#>;9KB^DB>4_=8_I)=N['','>]'J3B1@D&J
P3"<#JYA8N+C6#?6%5^;&+^E@'1=(D?:6FHIX_/YT<%PLW/8,5 ^]P@V!73GR@WG3
P(-'K'ROTTD0P#+6GT38WYVC41Y.L96H]O!\"'_2^W(@+16>#P4$\?64?FE?QF,-N
PW5Q.(V5AWK,[ZV$<5^00J#[=\ES,1K!(&ZP$L[!1ZH%MUZ:">"D#CKHPY,8P,.[B
P2AE4I,<GSM^A%2@WPCOFUR1^L*\'FE@O[_,^$)2GS'!XWE'G*J-*33QE.@6I&UN]
P*;+UYH;L)8$SO?F;]?L<9'B/5ORP_%:N8#JO:Q&&D-'NE;U+R0UE0R3G+&3"&U'C
P>AF'DHZ^)E_G1:=_22#\X6D?J$*2B\#/[-27[HZHKDLF;;D%,P ]L3#S;@Z._, >
P+G?81$4DL,?'=LM*)!2O)JTUG/'Y/#>V!]11G$&JT1V;X'C?(#(<VT?>O3!099OB
P-='D@*Z,E6.YN:WC$WIS-^2XFD1A-ZX\DKNW_L>41>=0GVV#]F7S]43VRPW:G[+D
P9K^:^(7KT!@3S9'M^;D(Y?6#"QM! DD@7@*-?-_(,X[>-S [XL=Y0^["*. =2T/F
PO,>"=D,+QWK!)V9D3W3VP<FM#</!U\FVQ1;W9 IS8-(&T5%ZLHYG$#=3-L Y:N2]
P_@ZLDR_(#Z[N\W2"LA6A_G#["&2=N%]@HMH;05JRA#[\">.6J#276Q6\% ZFT,J?
P!^?Z_F.G+_QM]ATY#GM?1F"834<'O=2E=Z)@5O+YK7B"*"[#HF=HV//8(0P_(ED$
P->/ 'N]X"0^?@B)X^(%W+MS\0;H&FU"XM>1,2A=KPT:^?5CWV6DNF\,6()B=Q]3P
PD<*4+M(,_H%C2N.^QF.&PHSU7>5 V6!+SSSS9EGV?\OFSU.(8V*XY5:V7'*'-&YH
PY+JSP)54H'B*^K-)**_1<OX^+M'@S?EJ-_C5)![\_IS<7&;@LZ9I#64]4D5,AQ._
P$T?9A9'D<,^V%73C=/XNS<'6XW<J2\900^W"XR2]?_7>V\BHE*48G(*=M!18Y@U:
P/"?"/6)7:+-:Q@;]6>T::K[9H9_,?U"+,!IWR\-.K5HR=*DT3?Y1R8&TL60(* 7O
P#61B;O"O?P*)KE#W$R!*@"=U*-07U>4<Q.;G"ZZE#DO(9%K<2[F_RD:2H;=6_B85
P)5(Z*)YSI9VK.S,\'GEK1R>22#9%&>^$\33$$I%PXQ&U=DT\2JHM6D(-'1X"0J5C
PF-OIS*^.)\IB=+5G8_GEXZ4 @J]2%ORRA+.PBU._5A R<D)H'M<XUFF)8N23F8JY
P8GH U."X8SJ60*\?Y%"UP45><@Q4["H<6L=6DG,4TBDQ2E;:>QO ESMCM5+RD%1%
P[I],*[=*,!!'@A?5ZL(_-<<Z!.DKF>Y^S@04X)-DFY,F67#>6BLW\R)NU&H,UJO=
P+ARSM<WLQ+\S1(D,/0&>%^"$@4I7VL9@N,3I:_K9[=Y"VMU@O@8*3U,1O_B>)^!B
P( ]:#E ZD&X7[A",/R XRLZ=@25YVP%\F2.2:HW2UG2-ZTQP6YWMKH?WB=FG?!$P
P"A7DR;'_W6A>RYT/4IWSWXIGPGK%N" TL&+OF3<)X$%=AE.:U9E:@BW>)C62)*LV
PD0909]G#K73TOM1X.1[I,87T+1:]9 'R)C&CU7T7&G'3S6O)&!)>6B=H1<Y47"<]
PT>5=+#TO<?B$;\2V:,1#]PA[5G,I$L#9_K7SQ"FP7(QOLT#;*#L0Z%8YAB3ZPP;H
PT.8BXG,PCV_Y47@RD,O>#OLV+$?6*XZN\;K#UOJ63/W#7+#?873@(L&SG>OG=Q97
P,=;&?ZSXM'.%GI."X(NXO"'<S ;U'(/O>H5IV<QRE4GN3=[__"&N3YQ,6.G6:#;"
P@1[1;G,R-<G@UR^$5?P%D])Q?#$9X1@,8AKMU7).XS4C(B.7'HUZ&">A<91\=4Z[
P5T+E%#;:KS!NH3+'1A0+B 1KLTKPF+@R_DX[Y8J=TF8.0_]H!7B"WZ#[6Q*!&Z/>
PEHZ\V-WJE77!AB,>378O$KO#B#BME#RT8] @@Z5PK+TP2C/I5+G0[NYZ_ZY]*B2&
PR&R.'.&1;._KVYJ^R_3D#%:9YK5ZK*,UO9;%98*$5_2P!=DV G$&W.6=U=/N/06\
PI#!]I8KA&\8]VIW5\N,A.1#K. >5&AQ)H.8?]H>I@>N^C8)YFB$URYCI=*-X\*B7
P182\]P>[/[,BXT7L9OV('T?4#!A^"^OG*9L[2MWYO1?IM"'JP<N1HIK8"LIS>(#$
P K_F*XZ/XK3^&JZD5Y:^$?4R&9B4HM8P!ON='U2<!K?X+TT#UVAK3?@&\Z8\+'^)
P?:1^._H>W6Z<TW6+9\4\@.\F^:+C?<K\N"F<JY:@%S1;T=;*[RQ*W6,&#3\%$]M5
P -;9YDTZ<[+NPUW#QR^-L9R!.?UR%Y4O?M&#S"![R1L38<84V7$8[\NJN-98-QK,
P$UL)XO9].LGD<PQC[(VU:MO-.M]0(5*"!EGI0SX)5.]'*4;+%6=3( >V1JV]G7]T
P9ZE[.MH6!!EV$,OG5M3,U,@V+W,Z>]?+-V2'O&L,^R- 5'GUBKNAG*7,(3]P3XT]
PO,EZ^_W0^PL=1<.N^]R3 U-_A<?\?TS=QAP06A"?%@'5"2%G"?R>8W;\PD<K-=%=
P2G)*7.F4[+ID%H-:9K0\!A0&) )M!/BN$[8!R"4O9M] F1UAY,^.F-.;Y-6.%N3@
P(I["$&3?[>4]4M;9IO$LBI-O^<!,>UA"3O.+9S5E_V72X3 [4/I/#T6\ZJ[C@807
P'TI0DP/0=>5^3/J1JZO".;_:C:O[3YBPOSR316'6B*Q2Y;2;2P5\96%7/3,O!M.$
P?QST]QF'3Z4OM)5$U4S,RI*7#O>3M]@#+>4JA:#\OP8$%M=?;%UP6X[^7>]?HF["
PP[4\[VWW[F+P!.5!P#0C+EV)7S$G[46V=2\/_D_:&[F9<G?&L.%[R1.>(3"Y=<0X
PM2$"BEAEG(Q&BA\*1E.XY\/=G<'*-$[\E2HKY/'X#Y'E)Z6>Y[0?W/5R>Z/Q?*Z2
P(R[$J=O/ R<\U&O\GM9U]$*Q12U[.ZI'!A9@G*T,T*73B3S(S%7RYMV5D6F4].%#
PSB/(/A0TZ+XNVT5&1PLQ]5)H,(9FB2-]1YW="WB4-Y"J\'^N9_8,,@TRNWWU.B@(
P-<FL/SH;4E7) ::F\Z(TE1*/JC_:C(KSC9'VZ(2<X>.@>!0$E!Y_]:*QCW(.'?XV
P(^V<6;!*G"LDZG&\7P_WB2"(B9Y&I 'W6_Y'M;CHH1!/RA.BZ\ 0'?1RRWH2D&UD
PW:K_/L#B3_0-5S "0!_8P8FGM?P<5\ZU)IU$BDS]\5:5W=A]?T=U5D#)#*EAC]##
PWHYO'9<%&\F>6F5(3!9%SPC1SJ5M0+<E(/"F2/:"C51UU@B%2CRX(.#\2>U^[\&0
P4( 1"7^GVD$:;I-MUCZFUXZUK#WY:_:>M&)9\D1M4N9R-MN6QIV=G-C?*$=:(0TC
P?ES!!Z1W0RM2JQ:,\32B7GL;5,80X9_%^7P1]]#SQ?N.D'<0F1BYM1<IKAB089&?
P+;#8^.[I+<#9=J0(:BJ3*QP)5Y!B;$3F!% _E4X]+RC5_IG&M&K?&W/UGVO(^ --
P5AF-6MQX!<V2SN'7!!JCRX[O%UR?^6NUFMKQV4'@&%@DK?]VZ5J"1/V=<M[9I=Z\
P"0MUASR"5H)F;SY$R4\I27?U$^O=Y.1PDX,!?&G*:<469/1;VM3N6T+ ^E],02"/
P&R=Y'?EO^$)%3OP%*.&B_WCC<-!HP)#=G=<F?PR^PI Q5@#)U\ M5O/<LKVK !\2
PU-FGVD.K&;[_E=3^?%RD$::\PNUY+0N%.VMA5B&/?<UE]WQTE$](U_00A4+I9.0<
PSV;\WY+YS,&#P=H/H3-N(3%8O7M&18#P@? I%A,$S&H4P;0XR5BDR)[4!8<X<G]R
P93(N/5J548_GZI.1J\(U'28=90&5"C@$9^'<5HCF-=6CW1VMB[?CU:)G6DDJ:'GZ
P]L1J<&U*V 2Z]' 52U\X/\N\W)H)I)?EK)KXEOY <X#6_E!$&%C8?3UZ>X+\;?J:
P8CP20=ZAR*N.3D^,N>$6XR4T!'-:Q$W7Y?VG7BCD0M*MX02<2$H=*0+YT%/<O667
PPN+ 1OB5U2H+3GIZ7#+-S=2L.JZD-/IU'&4&$:M5.A-&7O"6(CQ0^H-U-XKKL+NO
P-1TY[N?#$;D%UK$A^UC8>V;6Q\YJB44OOHKJLT!NN+O+,@ I=&;R?WG$!/Y[)=7\
P9%TQRM(,"?OD>.[6H>K)3D]]I:D$<X02%70N"JU&ZYG)?/+;PX*OJO;=(TMQ HLJ
P,Z S]/?VH<)YNS[S^^W=)MASV)I_<B([++TD%&8"2>V;]\2"Z[<MU3C3PF)?;@C$
PD:JSBH*INL,3%9Y=4XO/_0N^L/EDH/$3*2/([^N3)KXR@0&'S2GO^@&L^8.P6S]6
P8)3O6QX;^#?3#L1TG3S[=PH&B G\3ZB$;3L,7B/;H_G0A3/@G;S$DO4M;K#0C^RL
P2V,.=Q.P@L[D6UJ;JJ 4LW33M*!O[(;V\499:^!)!PIO-_ "2 (%VG-0^JI5@+F*
P#98D.]BIE%PBD/"BP\ M"NA(%FZ4QH1M484.G/=S;5T- 9JZY.-[Z^J%E,TXP!%*
P*;"8Q6N)QW=%X1GK:'DP4A:%/,N\B+"UEJ)5E;W1K@\,6$VOR#T%X&\;?<H48.#N
P .V?N*'[S5E;Z1\CV6&RKL'\)QUKOM_MWYQ(Y4QXUP!*)+YN@P\9)7S(CAH4NK;4
PJK2'61SX8/2[H":4FYK(-8!FM.]=*U(&& 'B:I?)LC2TIJ9[D96&I>FZ1!.DP =R
PF5X\.^$)B?/Q*W_32B:O=J&1 U"YKC_^U[0(O8IV:--NB]U)",V8JE"@_ZJO--!K
P[?F979OC$80(@X\'-UA/")L8ZCD"NB$RZ)-,<[8$/G2=J*E8KV0-M;? @F+'&/@_
P&::EYC ,!:$U7-5)8*P>$+9 -#PEL\67%X0U%V_,OTEH>[=1H4=3"L0"6&M3A*RG
P46;A(( W?S&0)1AO)C$&R_P5K*5SY&[B>* MY=#F@HS"(K)YE(\V[=<T5I\SX3= 
P&&D[:WS];C+ZYJX4)#A-D@*MCBI.OY>P?6;JI&7A-@.-Z0P=@=(0I_9.'@Y?I@$\
PC*^&A(CY<..4<*XB3I!JM(51*W(>OD8CNUJJM$G#7XYJ1_IX8642W"@NQ'!W>QX*
P[%3&5C6$Z.7?MDW')RAF\$$HX[-M6IFZPL.^5I=@;A;4P6E;]/]ZSD-ZZ+GEOY-$
P-9#IL^&>3B+&U./77$QDM-\P@/2-2?\VT]O,.D!4CQSP&I25%QX@:Z$6'Q3!B>,'
PIP;Z4UI=BIB(XSSR^@ D K?3@0)?>L?0]SMDG8ZAD]\S@'!27+M26"Q^CZ'00OCV
P:QT&Q8I< <^ ZMNL'%35_=Z(3G%,J1,5P6)L' EO.Z2EH9ZLN=4DMH9^J@5,K&B(
P;8[28Q +>F_Y@&Q&^S%&%K_V6>/U(8Y#YJ1+%#HM$_>K^8,NK/:TP<UC>XZ?3G>P
PC5_?'BV54R8[W_HS[O?VD!?=J< ;L$@I-@7,A4[UC"E2L$\PX&:G\1DL@A8-PP-6
P##+$<X\L^2$ 23\_,)M89\ GXXH$HEEGIAHY,NCN3;TSYJ',OG&;0T?E9+ZJI5Y'
P90&_3I'9U520?7%U4KDJ5\SL+G0=X(UT%:-\\(@Y.R-]3 OHL0ZE^'YVVH[S'#70
PZ7YMNW0D"GM&XG<RY]\#U#LX4!T:2GHSH@"M<)Z<=UM*&,S6A,VQR"R\G=AEN, @
P5S9T__9[2B)]:XTDM3Z^A]\CT#1Q7#7@^]8&NI.QOK1C^"8O?D2=5''1T?"0MK.?
P78-PIB?UVEI?W19TE4>BIL'(1]*++?L[!QD= G)\;:D'^:GLBP!5^T^A:V1XRX"^
PU<5]:TSF!D>+T\*N2]#,2S*IKRWR3>2?G[ VXM_/ORU<42Q3B10J[Z8EUSS(^6M(
P$ G5IPQVJ/'R\M58JZC+$[=R;M&-U[7#,J88Z#X C_?T#<-I7$*#1$VKQB)RJ<=(
P.B]A-$*^,WCBPT&R7B*(]=%3B!O+/;3X.$OZ>\A4(.IJ)020-1\RMEXDHTYYQ&"T
P)6Z9\_WN;'%'V5N7JL0#P'"Q/(<AU-.GLB^AK2B.%B#<B3OD:JT^BO$!!N1"E*6/
P2"5/)GB<95Q*;\)!QWGPHD23N?6VB2$OO:;1,<7FDR5EJD)$Q'/NX&#LX;6JB\%;
P4EP8W_KDJE\V[K%&L#PW=;U#&1R]8R-_7U%-QU>^;CYV1%Q:W4?/\S-%1VS7U>8%
P,.E*[T1"[;YEZ#K^Z<0&WH.-9!Q':B+,]GUDK/+Y12M*\MX[=[N7LZX5GTD,HA"&
P@^CG6N,3LE%X)DM,%39= B%TC$"6'MVWT![/>%_01H_M#.F"F.!Y_:"M@"A7P0WW
P?DAOR\CL>\CU<EZ/837M434DPRL!^]\L4S6OOB,<\F?N2O(K[C&)AWK'V(,K!YW.
P4W;7O@DYZB3ZLP^6/8>0;JF[TGH/7,.;((_2U=^#&!^("BS2 "<(Z/=4%39F_UK1
P?^U^?8D]PU=Y4)U(M<J>E\ Y0!,!TYC7I+<3.NV3]+<^C=*F?GTY XL1F.";;/3;
P;_/,CG%#O*V<8KA>)71. ;,O_R=U=D,=P09TMAXNH:,3E;APS+^>H8[/*TJ &@"K
PQ]77#E<;]/G/CUN>VN$L#%OSZ5EJC9 %0POV"MT@]&.^3_<0N3/%;J>I#K>-V2'6
P@=QB)!NV2<%\'8.B\0DT#TTGH<![M6Q1SS8[E]J='\C(/'6:/#_"HF8J4P@"F"/%
P/$-0N[Y)89:M2E9=U4VVA%3^<A(UCR3(M13+]>\%<3.U'1XX9A7GK09;AZ&'HIP@
P07B_%1RZ<6 ,#-&F3<[<&?&AG+8N:V,\40?*\(A+;W0 >3]9OJ.2*'^!UU_?P3\3
P!33V\7+MBGD#L?D*Y0/^8*C24"841$[+(-SVGU>:VVLFK8W:GMD\G9\W'M(-A]"W
P^L/:VD<O^FEH3QR'V\P#7)[KD 5M!ES'-M'NG\TCC<HH,'N5J5)2V?V?@ZM6"S9O
PFQ_O6"C+)6"*437Z^NYXG\WL$_C"7>=Q F-Q__G2J8"X677N^=9CW\Y5^ZWTU#E1
PGFP'<C+)E?D'2*X!3EB<J8>)1_F)<31#MZTGJ\NB7;;>PU/BY0(M^XC$IA2_!DT9
PDTU5T300-B0ML'/@]Q_BHY\!*[@+T)+5@J0K@)S4E.QRJ"#A7TT)HSXMSG7MG=?:
P7].TX/"+HU"J),%\6;5.F FD8,KF*33,B.<N!<W_]MK:.?+/#B>.N=H&45&D]HQ'
P@MAOI([NJ26'?_<"JC2F#:=2C<CY^JJGQ.KQ%(04%)9<3Z>&HQ1_(*J$_.33.@)B
PE.E<8:\P4+;Z_=P>>NV3."%2MSV%;YR&ZX^^A*,,D$FFQIMM2B:X:>]M8:G314VH
P8CD"@!3=?YHH5 5'#LUJ&L]+&]J_AE0F,%+JPNUCMP#R3/-7]M1(P!GJM8G/,P#N
P6A22 '5I/QL;L#NE+)&%(M;9?M'R-J6O,JVI5F2T\,EN/'2J]8!_JNF,%;3Q+!WT
PJ\H(@N3L^R7 Z$[ ?-U"<(N6F$(?-IZR..C' 13V@?X@1$]>/1;(^KSU!Y'\I&"U
P1H6RKD?/U=5BPX*?)S6B:7^7[>)K6/-)""IR*<K&\(T>F3@7*)T.P(Q@K;H 090H
PQ1YI<(Z;B@ D*RRJEC/ H4H/_/+NLI0?X_-(FN0E<Q[&,R.')D756!7#0(#?$77 
P^V$X1F**LD/^'\_EC* &87\Q4XY07DQ<4$&&7:J7V'P314]Z^90__3+1'W5'N25I
PB[M[T  >*9M _1:[)32#,]4GY #!/9 /]6@$N46P_# (<M?;0,KQ9ZFR'B>[#]2O
P16W;XJ]6"1=!I4;YOZ:PX'#/^BGX&LJ!^!(6'\H>2,:&W-9P2+2O$FNB8D;]PP(9
PR!THD5F9LU:^--^=NX+R ";GBMT5.6#G3<]H^[7]JF8%KSD&," .4 EB^"->\Z+(
P&*# "^4TQ#V6U(L[F>8K0.5\++Y'L+H]Z*B'&_=)54Y0,8;H3D1TGN#*FXD(-R!;
P4=M@02VHTJGG#J2Q;05R6.QC>#DF8XG##%HPOX\[UMQW(, NZDH1W^)^Z6J@HJ._
PO[DN+I<F$X:X4';*^B77F1$RKP!ZW*:HA^O6'R7TC!IST4YAZK(TQS)B"YZ=1_HZ
P_*TG9XMVYZ_WFP^W5.\CGUN*C/H$H6<X/HJGF/4JW#G4(831E-\:[*,(<,V"6&0K
PB?7K)O#[;T[-/XE %B26%UJ8O2"-3;&*!-.'7^)ZD^C7QS@($ZQQPXQHQ'M0,E00
PJ&8TN>U=0/K6\/.]/C7F/8_]PHR!R4@@ A6  &EG!BRQ#%A7PCH%^7B-V?; LL%C
PA?C&I]%XHW@Y3L:FUS4FXX^Y=,$L>T#@X?NIWTA=%W):-T(Y[1R ?L2.!^6_5%RR
P"^QB@$-4I?XL3C5+*M5"64KH;4-:GF__Z5_=.D0L-!F!@=&]47IXT+1D-)Y1D[,]
P^U&*H].EL>1>H])C].;MJ/'1LBM +.K_.--NYK5;4/:S6Z&YKARG4<*91=FJU@;V
PBFFP4U)P[Y+LS+9Y8+FC"7!V*21TQ1W*]+E:1>Q16;Y]8Q<\Y9MN&]"N)-?!VT;U
P+C2,50\@<12IB,](G#70;%5 _:S);,BR%J_*2($98$Y@E'@.&-0+8+3T(-;J@Z$L
P-=+B&?"8#<DNH>+UZ>YFGQ=^^E,&)^:<FTZIA)6>V@8Q3:9)^V(_4<9[=DO422BK
PCX8)F>1N]W'KM3)(FDPMU__;^.+HX2!T9QZH:"KJD<*[3%AM8<#NHY=E0M2.*&<=
PDH%[M_?8D1;\&S]S%*U>*I, / VZ*)'$DR,@6< 8O=7+P'2CSQ<+Y3X#"/.0[<;G
PKA.JDV?34+//O9[2S>RDT3HIDE[ 37E$I?"QZ+/^4#<"##_9G^$#$#^;F75EP[0N
P_^K*7 E9-RRU<5<^I;S55+V1OJ#L78MKA+81+W-B1T&DCNN,'CB8A'TZ@-9(B'.!
P=)CZ)G):, T.2K90-S8GSK=4/T8Z@6&,OX ,!&W^!T[/OM<K< 738':BZ29&Y+9U
P45$F+#+%KKEA%)$<++; (JQV'AQ;ZD<5V4:=%>\OU!I$9ON!:45K!BBVPP7Q]E1-
PMLUN?)XDY2L>NQ)BJR4/\T<@%HS!S7V>C2VB3&Y8P#FLGD4C]YE.9N*>JVUVA-;:
P#GFZPW3N!D9RSSUL)GT2)OOSAOS*:368GB;"PCL7NNZP]TJL<-NNI>O@?/>"*%('
P)"C)_!W;CI?] &C9YEV/NWA4-^T<G9&XE&'XPA4[7%)+4+LO[5?JVO18<ROL45\T
P+;6KI6MM-[G1[5AC"GLL[48T&K72%DZD9M.E!=>%D5)AXQT,;+4,M\&.'^?*RY)H
P.VSXO!/2Z05C#!=7D??G)D-R/U+19CVE;X&$C7]>XBN>=/-U/K>C<5ZZ&I["$R=/
P&@?]A*X;Y/NC$V2+;BZ[Y1G!,(!&^]N=#:+?)X[5]LAGAEX0#* ,M#_4 .EMJKQ?
PWO5Y6BA)/^C9^8EL+3_KO5++C9<!D=QD*=GV0DZ<!6>>M7XKCM*J&HV%IF1!^[8S
P$F*S?_OLRD"$SS9#UU#@TX+G7A2O[*5R4/\;8R-I(I8T0+ F94BS.[;E.=T;Y,;.
PE)\(YKG.MNZ2?AY]8GJG"*+B\T&KM_ 7>T2#<LT5&8_H=W$RLAUD2+7"DN(-X+WN
P2NPWYP+&S70B&PUD-9 .U:W6K;@5KWO"C0+-H"U$LSWDT83E0!%-X6_Z>RE@ "<]
P@=YFP+R5Y9ZH0EH#:0H,)(5MJKV;S4$%>FTMXO$F<P@ SUJ20XQ#6^&P&H>7>3EO
PJ^7 3&QXMQY3<(V8 X*&)RKSYSQ_4S:UV16-4TN*G[\LY4P4:9RW*P8#L7L"WAZL
PDE($_)GC"E/O3$K=+OL+IGS:T5VD2/[Z:N#S>CH"8*BC+!%*SW"=*'!47J3*&I\I
P5^=!% .]1I<(3/C^:8S[A]$Y#(EG_5.X@G>PW$&G;",'T2_(3X*%Z,AAY#Y_]$'3
PRRC;_;RBF$(S!8I_%*$=HCFW1<TG5,K<P^J6A-&67$:]0DH^8/J:YSPOSUX#G*+H
PHW!"\OBYI9Y1QM:B<PIT<V/"'G3W6Z*IJ[SYU9"0>3$&LO._**B=2&0TS/#]NR^H
P<:R:7V;H@?EA?.>"X7?O-SJJDY8'(K8'%\!W+IG(YL8R$J )VZC_7\8.CUZ\1"UU
P.C,L6(D:#BTHEA".JE0LNR;JUROXT$X3AK<[V?HVG7:=1:Y3%*/JO+*=JM/T\[BD
P);%$=3]F?VYG\0*^4BP '=!<)'/5M#VZVV'0*XTW'/$R E7]TM\GV+?P#S%-#8RL
PP$=SJL45\^MRI)\=DY]M1S2\IH8A?^8@S>UD^'DU' 6+9CVA2_NB6F)E:PB["07$
PO$5XZG%TN7&8LCG!UPE.:[E^T;)T6F8,=@-Y@2(#"28T0EA/<J*(;ZW\F0*P*^LG
PE J-/Q;'2C7%!2EU'^#04Z3&5!Y"3C% ]\-A1#@,^DX_4O(E:-Q7;_P:\2)[:VJ(
P"<DZ>$ :;?3)1!P!;2]FNJ)1Q'2Q3 D;5@:(_8R30(@#U/+Y9RJAZ)6A8/:NN?E)
PI(*MWKZ^+#C^@Q B&OPNO'WP9L,9%5#\TPIY-MS=11L$. @NBC',4%EJ_5L^5HVL
PMU?N5[FU&+9<9*<[J,YHLIT&<<86(SP&P>VJ:*X8@Q</%#?P"9<R32Y]HY$?)ZA(
P1:VQ@UAKA-)0ZZ4%']7USP"Y*2)8XOD\2Y\7[#61 A$JB>1RXFGGHUYRBY?$=[7Q
P][:#U=#C5H5:^SZPY%B5H/ZZZL-%&:OWW-JRY />SY;G10,1H<7#M^EF_($0<M8+
P,DZ9T0G2!S#YYO\RC%8U,:4&NHBCDBQY%N#4/$!T&'X/& _;+BD&U"5&G<SN3W%*
PB1<[TJZ,1Q5Y:7%W:9R"=[:60$,V."O%<<-"/F1HL&D=)D3K0_=<,+)6*/1#]2K,
PY\:^9JY;19):+(<8=I;*-30]LLE;H,C& :+435X.!]KXFR=6XC V)"FYL>;^?HE%
P9JE/S07@ESDEYNIG*<[Z$D[IQ9T[@YA[, ;G;JR4L[;-IP_MZH^=BUK<C=_BX09Y
P-&*M(5&L"G)W/2M*8^9B;=2O4N[L[UY'6^GR? U^(<A)"^""3)ER/^JT?'MV0W*,
PLW*BPJ[]XX.Z**P[Y<R9RC4_H/^X.F@V8L(>TZ<(+AUZ/'><,HT,]/2[Y+3_#BB,
P"(4I&.#?[H/.2P4O<^!W[S92GC"!B;X.?&R*HUFL8>/AF07F3P3U)\6A7J6A:?PT
P1>[PZ\K<ZR.[U>5^=2\YL68D1M@07K)MOU  >EQ\2KM'/21A1!-T_,+A='4@X.LG
PAI]4*(G94,;.1MY8;FG/:N% \L_6@;9S*D=2MXF@'8/P!A5X56V#'#.A-3&(QRM_
P6KM7ZV[LUO3]!W>,8&>G,L=JA#/-M?,=V1I)[.SU)I593S ?B;8/1M0&@8<#F/2K
P6)7%)K<7_ME#9N^UY*FE7(NQ[D#)N!>:T81!5QR?F]E^[Y#"KCVDS>=/:?[&M2MD
P2+KY,N]E[W.-?DBM]-']\!V[O:[;9 QA?SU.+ZF./)$W)25CXJ=3.C@/O/N"@N>1
PP5"#N)1%Q2L\T27R@OS.[&2M#B&_4KZ@-I^SK2\,"Z;K"S',!&P\E'Z1[F;O-*TW
PUP_I?-EF"7/M[KO_RE&82<.?@3M6J[0N ]A3)V0 4_JNO/(IN5[6\R==7.@"+,P"
P==R_>?+ "@ >'GB.6;Q_4UGNW'@<<KP94_B2 9)'L/!SE:J,_/%2CJ/WTN0,,HEA
P5S3/.$16:,+1,0N4Z(O0!8A(%?/U!2T7O"[C)4\0HX.M!N$ N+.1AWLT_RK_>UT[
P5P?N4@Y2:Q/6)KJ=^MQ@R8[05J*A*(=BR7 239/B1K,W"45)[)N41)QI=+!CB#FU
PQ$\\4Y';2)YA2L$D[GBH98I7:R8#=KWZ20Y[18N/4"I=2E>XR/0W*\0@C13O!<XD
PZ9UHG?P,2<I /;@@^V^E8J&U;#;W.X$=8Q=#>@OS;4':"^1&&X+3B[AA2#E8LC:8
P6PKI88L"M,XF$_=@0??_@L=Y)P42QP/"W7,Q,W!.!/F5_'SS9(Y&P$%\3*I[,2:$
P1ZI#TN.UT8M@/-E]1\:%DR\%%4BC-@XJ"Z;Y)Y,(<Z\8MJ/[>*(6IPW-8SZUA517
PE2D(N@@A>>NG:D(MZ--'+,QUD6B+A\]HK *+8DM=H16#ZX^"DP7ONF0%;WWFU;C!
PS*6&GAMQEUDH(@6R%(#A[1A?23<<Y]4(M9N:*0E?X^IDW5V,*\],F.A4"7KV6?[L
P]5"!-3-W&?,KJ996AD?J+L#P NB1129.&]L*@5M-3&,Q UPHQ,B"(=X9-,)<91-_
PC]I"2W\8FWI$Q>$R+B28)K-65\+A7G8P,&+-LFD9+F"HXLWI#3H32N'(();"9LN1
P#,W<8F=#C=]K&ZD6^V]: )[5$+JG_>G.F'\I6>(68K/KO5^C>]AMN<-W4SL'[1$*
PK#AEZ#F$BZ*'^9J\QO4\08OQ\KG@EG5]US1GUL@3"1[8R1QN%G <MU<\6@0*JZCD
P+.!65&;B3&35&Q:OB"]@RE0E'B@^&])WL2-Q'.\$"/1?;LR71[[,-'@,6F8O<W<S
P^D.1U3,Z:=C%Y:?A-T8DJRA5NFO>:YML4V 9B78+PF0/%U1^S64L4A+,I0 CSM9@
P6%9BPADO0&4'H>>;JI@F[):'G#AI/7:,[O2F-:HE+"-T"E^*0\>%[]UFW6,AV'N?
PMVUP]@=]V[]!&YK9/8.$MYOH0U'/.8<C%IAXH8"^ME[>LB+$#>C5?1L5/8SX@"^[
P[],[B UH-D]_F*< UDR@3/"HAC= $2(M[!9$]N'O>[_./[MV^H5T0.R41^ 1JZ_O
P$7'V%FL!RV\<_%C2ET(NH$KCK U.<@$2PCFR\\4JX(@8URQ^GU 30'';V31))?;W
P7?,+T9P=MHN"+.74=PZ)EQR$-H%F\)IRTD!TF;"Y@V-&5RT)OMS?L*7(;5WB)J[I
P6[CQB\5CQ1SV_"-"%PZ"<-%: ?)RV>6'6Z=O2\41"D"*TD)# NPPI;]S8,[)N)HQ
P2A49<;J3B6!P@MB!I]*P6'6">!RJ!WR%V0O5;8T:>35(6SD9Y*]DYB\#Q[)]J^DC
P_D#)PII<GCXFAK^(C0*4[N@N_W.K!=5RY>USYQDJ]0'5LA#+)&$\N+@(J;'F5=^^
PVYG/7]S.#WG&R(14#:!JH!FRCRQ]#,S$$K)&_&YFG0KWB(&XDN[I\EB33@$<,;I2
PVK^@, LJDC,)JI*;XF$/I;2Q?1H&AI)Y(@;QRX8/LE.VE!$$G6C1S&<7$+NI-&)R
P#2A];9F)!:L.,-HV9&H#36;<NA-RP9: ]=KB/=%0E0BJO$W,2;3"XJ1LI<,6(6K>
PN(8_J*(<Z>/ X2Y#/(7W2V04MPYICZ5RBU^@\;>C>!+Z.)MA1LFZ'N(96(%*&1+4
P/(Y2YQM04KN)V_^TY(3N09[FM O$2!L'73;@OA*Y0W.>CPV2$\A8?3T>ANSZP,7T
P?HSZN/W&U2@,9"\]R M%=+[8!2VK&\,6S>M),;P-A<0R^D,E>L5S);EW#/>ZN/#E
P\S,_/>\:J(+I @V;[8K]\CV;NJP(Y8H3G9<)%K1CHO/C>64L5D(*K!+V,O!/+K8K
P5\TKL1\7@S<BY+CL/&7,%*.$ <A60]%IZX%TPZ003-O'  +9C7G)"Z)*'27A!NXD
PT;!)5WU_5<?:4/33M6\G:IL +8$LSKWPXUP><(O#^J^ A!#J]@P[^V2CI <<_)@,
P,@P-ODB5@2.?TPR[I.R3:ZWW QY/E0.]UY"KV$']O_2)C+PI8PZ/(6JC@"8(GL3,
P;UZ]F-=BL!B?%4/*RAD[<(SL.($!61%>MJ)'VJ'^=!G!=*']"7%,N7)N,0&\S)'H
P\I<_.]A/Y9CGU6+O].#   U\>>%-O* RPL!,E3:0X[ 6:^HY!@R.7^"OKUSO[<4;
PM>P:E IJPDSU "I##0,1,Z@E,9[ 0G9Z/8X):!E9=A U:O+YISSVE9J.'<_-,_Y(
PKC";T8Y1!4S8T,1\ID=SIBC_%]DP\70O.(6_$8,2GXKNCUE=G6\#)+)FR?!(6XN@
P;)'D/JEPU3'#,AXB)3)S0HWB,V*5R>M5 #;_I81;-;X0WNL?%6(PV1@EA:^<W-2$
PWIB47%B1434+8G_/,=_>B(^:'=*;A]\Z^Y[VYWDM_[>SI+;>\47$"BUX<$R:(BZ;
P;:J'JSU975=Q/U'555_A0^EQ/G8Y=@CED('_HJG"[ZQ-JX^AO_7!66A?8M.SS?OU
P$CJ]-$%:*A. [Q]PN7$&I+8?<PUA-W=&(K9I9@>\&Q#0SJIU#V-IBF_K?[OA0]5C
P6\:526;?R*I-;2(SJ1[K7.S</Q_NO,*ZD=X,<K?W5I'CH:QRG*"+%S\XF"P#8^['
P5QV]OT"I5;3:ZU*!9"U%U@2A6Z0^A=_,)6E(5KJ?[?G=2SDDIR1U'II]J1-"_VI+
PL[/7C/3#QYOXJ:7C41>(0@M2LAN4H8C#M)XW>*]>R27K4KX7[7O+75^++_"L.B6T
PI6 F\,DY:6L%6S8F[:YZ1OV*R/F1(HN!Q2KTWY)1RWO5IX.SB'+4U4$-8BPR5O_(
PS("$_#<1?&LD=I.1,,I(+='A[Q;$ ]=O&NB*#3#.2/=L=*%@S32T+ZPN'51/9*.K
P*ZZ]4!4,H;LOG2!00_D*&(KV>%HRMXH-\]\SI%@_=P%B#HJ\*^77KAWJ2?LJ5/(M
PBF.8?D!QF6GU"K.8E*5 B$Z7E& M1!=3:I891-F[ZMNH+550JRM+O=;/L.#KB)Z%
PYTF:V9;;I6, (@$ VSD"K[/B[A#Y63=<TOH!$VP#UT@OVW4G!Z$A'1,?JVL"7P8)
P+?IG*3DL ?+SI7%*)JV.I,T!DY@K58)^E,W .+]Y1J98Q:Q6 \X$YL9.>>P#*9M9
P(:"U+:0BG>FH/P7!N;N=J6>.=%@C,:[\B:R@TG4@]G<VE4%?S(6.LE^V#0?UN)(Z
PEP=EU9K,Q0Q3<>GX77!NBE@+QK&0"R;=4,P/E8]LTLQ8?';OFC&(#V"."W7P\-70
PJ[=4_5"H-\I5#9J=/FYW:PHDBI=:Y7(KV^GW=77:2)H_RD3%5/KXAWAGW;=Y39)A
P:*U!@I-2TH1Z+_VRTL(#AH-K5_)"=X*.ZH;[EQK;D9VI>U=C^P8EK<>8>>(_GY, 
P)PAB:#8"#)%@J/OLS".MTV3 RC8')8XBYE>D\C9/;,0"I.?BKWQ&<W<VQ()BR^VV
PN0N8UOM/&A'V11 7SX$@;A!9LZTU3P02SKB#HI?FV'&Y0Z^Q5@S^F0N(,C0O[95C
PGZF^CL8/=K _].4;),;(VO:;B-1UJNDFB(^'B$$BG.+UR/!!7.X_*E_4A1B\]^0F
PX#B%XPCV,\I&VM<BX&C(#(935!6Q/JF()5.2-5C#;$-EN:\>C6UK:BQF+(M>X8P9
PKGCBG?V4XBJ'48//M#00 1*=%] ]I4YY=^$?T+]A'._P[!"D4A5P[6(_^T8!LJK.
PYWBG<=",4'P_,7""<!HVJYB.Z5"N\ZADUQ857Q?N#0C#M5 S-/N0RJP;2BQ)F:IY
PH391-6_KM4S_ :"#,Z@545;MY[>LL(1OXL*OR2Q+":W#LR\V!H\F+-_Y1:O6KB>D
PY3E6!]#R[5R#7L/(^Q^K8),*7-?IW5-<5PP,;!LT"EPU-MO\0K.!C@=I7H!.*C6>
P#FY6=OOQ#/0K4W. QP.\V^>0:-H=V#_*9Z:BHWV?[%47>6E.1_.XS8-Y>CA!?&.*
P. $;NQ*;6,P(1I2N+LU+/TEM4+8[C_GW,1<X4QH3;=K^00;)7R,^ A"$RZ\@(T,"
PDB>ES'A2]'[[JM8;OM)[]3U3M  %>3/JR/0"$8MEUW5OF%.&V?B&)&&H=#T<?L>'
P=]$>C0:W.(;#YQ>9EOM4OOK*'(U6>!3YR:Z-NSLVEIX)P..PKKRN%8.H2?0;DF81
P.TXF3!1W[@UJ[&=1*FA-P>B DJ-619JGZ/^.)^773;#O^#OFXC_C$JLZ0Z:#>N--
PEM!0?9_-?SK+VV._CI>F%49/D7>;11_YA4&1O-'[QH2S1=#E^@0;AE0;L@ 094L>
P:'\VK3HMC15G[_S:+$14=JRSJ4^'+H9YW:;*+$#!Z]@&K '4\Z8N!\18L$S2'8 E
P\'])SNF18'1'8HXC:OXB%-(#<NEK.I<YQ1M]4?!M8APDK;N_JKA+I44=51P>77Y>
P]9/<@,8?/K\S<.8V Q&&?NCUZR$<XYGED7Z\,2<\Q-G^E$_X*S*Y:BB!F''HGOF 
PSO _AU<7IMT5]F!+?5DS*^7P'W&79E&,,N"]%;('\^'QOQ))]UIVY-U7C)AA:X(B
PR 6' ((.?N8"Q*X0.*</T*QU&,W/NA9OU 2(!LA+I7U]!5JINZZ$?9]E1Y#2B!&P
P #LU^3#K7Z &S7@E@'G%2ZH^A6X84XKRZ6Y*FOP5C<GJWV*=KA=?T^97]U%3L+_M
PARZM!=C4T:ASGZ3HFMI^D5*QF';#WEM=)XRC!7);KQM"DP8&,LA1KMHOU*;WB!:K
P@2S,1UM7W/8V?>\_N0T3H8Z^9_P;:SPB6FI&MP/1WM]$YO)\:L\SHVMV2/HW:SEZ
PZ\M0%4"L._6.I>?DAI6-[5\X5RI&Y>D^_,$(K) *)#.5L@-JK6S/M5J!MP.=][ D
P)!.0=S>Y^U:T %>DF';L1@2U_]>Q?G<GS?L&HA:G4,?CCP2(0J*R?^]XLC6,< [E
PYD%9CXZ][S)3CO9(1EB@V.I!]L=-E3 +MC.E4R!X<JDQ!, ]/NDPS8-[T$[R&[7E
P%(O+PJ,-[\#ANQ22BR;\:_+/-9CLC)-O$W%+ZVLKD:VZ]^8L <Z^HQ*/Q#[[F?WC
P"W-C_8BYM7$BQ/\G'$;VME\!UY9SV.Q 3&-DI?/[?J\'1'OV9]-GRWAPBQDD>RR*
P\$V+-C<EZFX^,YO;L#%M9*>"Z9\ZF&C^^C*\5>X'L2EOE*FUP$LOK2D-:=@O(QCQ
PHWGMI)($DYR)NWI"[&+O6EAIS"Y:R?N$O@<ROH,R7.IHJUUK.=\^CG!L>?NF#!7;
P(]6A_#+0=V\_I'J<EQYTB+2#Y%L+$>M4!=,25**.\87)9\;K"DY+:QI8J;X:A)>@
PQS=?8L>F^(%</MRD \VN JPVR<[B\?2(-'$B0M3 J>WW7<K6(O//6)>.>CXM6,R(
P83"T\QA@138X6\X[>6:YB%$Z-.5*QP30(S_.'  J"^$)BSJQ&-BQ[@R9<XN/XC*%
P%783JF#.-)M3_6FT6>*8#J8IK;1. EMY\&:TQUM\Q90DC:(69JVL_I8?E\%J6U]G
P7*;@(E3EOG,_Z.H4%?+VE6-D=#\KJ-L\(21(Z;5NOAM:Q/ B[E&UZI1V7>0AI![J
P$H*0$W=,("S3=X:+ 7>3]61V_=E!U:#+*N>Q3AK3IG)/(=CDZ,JB+".,$Y0DL')T
P*/O:!B[>6VC=+SUBPXKBB)S/5/G#R;;/*\1A5#!/8U8HQ:US#CMK03S[^[W*! [C
P8X?&81C5I3<].L]2H&X$)GM0#:,X&'HKV4]7W 3PC!+I_L-<96C3)N4!UI++!8E\
P7,<BV#5P2-B.\(@A_"1.D7Q"CH@/W1.TFE[ /P8#+S8>ZXZQUUL7A:47P81P)"@S
P:AI/0H+CY\T.NKB*B(L#[\I\D%^J@F;T>_MYA4X%,E29&%<CU?RV'K#I,WP?ALB-
PM$<&9[+EYF9"-,)\5B.YEX+@+QF>^![VYH>PJ=4 5A?V]/I0!L,"WGW*;W;62FC8
P"^J7AP=-9?"NMN9D43.]AUTLZQ);A/HOKAJ/AL,6RLF08$^^^Y*,P+$]3".Z)W*!
P.<X8[O!'EA2F</)72C8'/4Q[?>L<)DV&>M"^YNG02P1=F[/9Z'PMS32?G:-G^33$
P>D"BX%XSWZ2:!DMI]<UOM1@5_NI6&'Z_R]464;7+W>LFG/I'[;PK;"4 8038MA3)
PYC2$_" &!J2_XXQW%W;S+FIQAD&-@?_P'/LG!DN<N=3&59%U(SR$P[=5]SOQG1VN
PR4@U9V2FN?IYIK&+M\+%M/U,/MGD1<$85DD12*Q@FI]2N[U )&N#,6WG=S;C*^S*
P7#N5'N)I$A=7%,QN]U/0EB#.*1'/)FF0_ -" N0B"%KJMTD0QG/? KDP,'#%AK6$
P*%P5-W#-NLZ1Q$ /LM0I&YJ*L%&[=9%76K M+>:^3%8IM>!O-*(B^?Q7)<M4;^SH
PTV)=T,S" H<4,2=G)'2'*2YE>+<!>@*2R%YPGV875654OFS,IR O+BVH+"HE$@[]
P_2I>8 H/X=$C]3Y5),C3['TH\", 4$"BD>)A1',I"F*6*B5(3)0YA?Y%WT^-IV]U
PQ-%^8N]*(3U$85%N(L%CF[]K36KM]F"'N6.Q;-[[UP$-I6=]I&WSD2B%3 L/LY8G
P](_@L.I,LBG@3X,6"=BIA<)-0#Y0Y1-K Z5[T.L"@4H9]J\6OWE.-%LPFY]+2>9)
P!7MH6AVKT)]-KA9RJD]X,4RM?WF-@%[8MD56.:=.XCH")*H4T-F*%]+HA+7OQ[,V
PVA=A"7O1HGX_6M<'! _!)2<=<-T?CNC"EJL_P$6:\)-I/Y,RSM;&,^U^N5@6R;O!
P!++,7DD^%$[T]FNE,\'61R2;N_(DI50/&\\A^ZK^.!FG3O/^[S&A-(HMU?4T-[6T
P*LK<&30+QL43+PWYI 061"SC+U*X<6',E@?;E@Z.K3%0[O5(DN<B%YBZ+X.RR.+*
PVO#U.BB#>K5G'F1W[\4F9NU<JO_,7YUE[8(X!Z%//9M)6#[=G'V@N>#E688C]@,*
P6M<J@3]Q:=."?&I57+V+S6%[).*:(36HJEW[<=.U7S/C$^6^1+K4\H]%ORFGI692
PBKS^V)(KX0.\&<9V1IP#U*0]CVJ/<XV;*(&) ^2>,#"!J\'^:V5+(K-N*4N=!V>1
P&V2<MT))?D]AL8S9CNKJ41N/'<!'_I_C'\FAZUTR_RX,/CX9'%*!;/"1B)ND]18,
PCY_X-X)$P\-'R4>VC>79Z4&2;/(+RJ9&%NOR0&EMU.3X8XO+0^E2Z5F&G>ZZ$X5;
PTQXYV]K>NZO WKKK157?'U?>?I/2R.>^",P"]RU-C4YD4XZ.8*^K1I"0:%C"\)R$
P2J0')1UG%]*C8DN2^";,(-I"KC^7%;QZ1_'4F57J6U216PWY'4*D#99[;K;-7JK2
P;;;NGV+93Z1?&!<EI"@.*+;[Z-U-_I]>WFL612?5G!VN425/%I&I4.VM#]X>R* @
PK(MHP"J&8O!41DCF^K IH+'?C(8=O1T'*+4&'V"AH1)7PD1D"/2R48RMDARX!Y<T
P7-4DG"M4L-H:3@LZ'?'5GYTRA)$8)/;QW/*,MV8ZR^%>N@ILP]*-1NUQ%6$>D0\A
P!D5JJB3_W<MBP517D@K+=T1P(NQ/()M-DHS+JW?LW 9A474)^Q)4,NFPAXS"?+!F
P2?MF'9\*+_[:C!DHI0;2T2*_!/EK3#ZV,QO(-:L29CL^^,,CBC?%>^<IX"A<0G$(
PLP'%TJA$^#))V[.+STB#DBVJ9T:"_,NI=03!VO!L:N $FV>!,<HGM%6:O(^%-$MQ
P8 :7S/D<DU/?]Z9YM%>"93Y%58#&VOT1&\^O/-M\WA+"L4T;4Z,ND<'A/Q3["YM/
PW 5-$.D^:DG"!S45-S*R=T&I^39"+WA>Y.0%NMA/Y(8\+T%>[ ?5E\PX/W0\5K/U
P^6;C.[G._09<$+_'8 "E571@L=:F(D8NVY"010_8A; -K):HJ"(Z1Q$)T?8&AUBW
PY0>"$%.%3U+V)E'=U11R%=(65QG#7TI39(P/Y32@"L0$>:P*HDUM +V1' HR:W)V
PAKP.*^'LI@\XW0&T01E@7C*1YI2OG$8B2;U/-,Y07IO(>RG'XAO_DL2?'MQ/F<:V
P*UNMB\Y;U#FB@W"N#0YS([1 +82N2M+%Q7*@4RS\ZHSKJ5=)O3%X?<V,^.XBQ854
P8UJP@$]AZ0.[-L_.LLN^A6 *J83+ S?'K=29Q\[9CB4E1Q9E+H@VD\/"D[9MA1L:
P!X\G8*R*Q(IK @)@)7:,S$-3.*(DGG8^HQ7!CHJ?-^V,+FY=#^>39>>'.V$+O@BZ
P+9J<!'-<?J/^]/ZZ$A$<,-BKV[SPR=2S_#E]9]4ANM!%GM=_1'$%Q4XZ#".$GPQ?
PS+WF C"@E!/*>J5VY)!KX[]G>S,3RO.J[!*EXLPL6$I1Q69D]XX+QZL*KVKBQ^=7
PR+Z PY'I@B]-"LCD,C]J4.H-5Z)H$:[N&D224C 3^?,2<Y9B+,(T<W%![^JUXM]>
PTN.V.O@ZNJ'W8Y"/,PFF< @,Q8M\=]B]J7#Q-B\2+&1>OY]3*.G)RA?& +[$B9]Q
PHR<%\/@;C%I>55&(!9'R4TS]!=ZBSU/@OIZ(/CF$LS5V"K?KC+Q<$(1 Y@RL;'"'
PGR9W@!K2OV[N]TORP9<^N?D>R'ZSJOKJT6AFV-PD)5<OL%<(5^&H_AX7O< SRE5E
P_-U/-+XLW06&\@+'13I$OJD67WL?9@G+P15L#S(J??QA><DGG%M8CWRD\$S]1>22
PUP84(:XH4I.U-.P.\ZU(8^!K*S-"UIK[XX'3Y5B6GAO#,FH._4]XP-9M%Y1I%&7&
P:V&*B3;%E@2JI2/=4%JL80\@&7ZJ4)]^+P<%8MM=U-35&^M_%D1.5;AIGQUN#:II
P"DY#TP HR3< V4.[4_W$ILFQ$CS4D,,-KWI? [:(M!&$2B+&"Z#8B9^3"[2MZ&L-
P@3E':*UT=+=K]K MC3%?0Q)LS1LJC4L'0;-O=TBW:"6?W/Q2*Y=,_J=T1,'_U2-O
P=K9 @4'<0W/"XL(%7C:;*ZO%=ADU?A^3WFM@7*KPV&%86Q*.\*45-@24C2_4DYEZ
P,I<XWLT^$): ]+J?>+<9IV%K1F.#Y'DA&^;(DG]#8:=]Z"EQPZ9U-CP"@.^_/S9G
P1L *[QVYWX6&Z'PF@^MF/86IA""F-*+MM@(/AN,&:;O!3[J2P4_7VC%-PBC[ ]*B
PK/)JC-HD;P:A6Y/!M&B,9<Z4L A,.<$-<M9R3;+ '9%I5N,I^(&E5 =L&A@$GT5=
PD"?7U<<S<#LT%V[%Z&;5BJI0#T^43M&3M5[GTZ&IO?L=R&4RUR!0E/R3H#3H68Q]
PVH48RZ63'F4.*QP)W=HJ#^0^417I(;@?P@E8[? OWD@"J<A)<#1J2%\CF>2.1"M.
P^N988=]*H"H.BN*\<1_A7H>$W#@[7\=\7OF+L <3TXRT/LA RRQVNRW[D?N?B7S=
P%ZG]#^IM@B<A973L)'1W'Q%9#:]=?GO;GH./>!$M6([GBQ"#G^E&O$9E7C\]/T,Q
P*KTC@0CR&.&!LC2E8GJO*VCI0'GD5MP_J).I L8218P@D:A.;B[/(B5O)+M)XTA!
P(/L\^^T%/M9HZJOK>\DY2F.D^+XU )>RVEPO MV#W]4LOG7 V,JH;XR?@;-)MM0J
PS]G4!4W@G#I+V>J4!Z>O7?MMX9T(OWD.+0/ QOCJ>L7^<DNSFSSO;Y8B88\BUXMZ
P0F@GK 4 2D=H2.9]D&S\+3CD%$@(>/(IDL9>B"L+8AH%N? *LA,\(!-IPZ[S6#+^
PM(K:HG-CVG>MBN7(,OALXY3BW-6+I':E,O O?H'Q3U"KT^LO,NZWJ$/XDJFG$=S=
PU$;#WCG1 -2]X#RP?DWMM4TGH?_>"]9G,QH7MS[=H0.![$[@H J_YA6RR1FQ((H+
P+EIT8JX+6QV9O=.2V=^C;B1(#$V\89*C,RB[I#_ZV_YH*[H.KFP5S#!( .K9I%Q>
P&)"QGN8*5#:7$-31XK56-G)Y%X2-V*-E%IV.,.JB,W\RIWYYJ*+FV/RX"XYC96QY
P;(Z&R7)]K')/-9#S_%48+?0D^?%L?8M9$PL.:\/!@(R'(WA>I3)1U6L(=Q)V=,>0
PV^;KOX W&C4 S &^TZAI=&-O$15J7M81+_ZU'.^M.!QEIYBGGOY.ZZO8OQ&0XR0^
P5.=G'/.E F*=.#W78+&(?(H.?$%G:,JTG. L8_:X>?.[IKY2R_P1AU=>#LT?HA*G
PA@+(+IN_@HN7K_L=*?%$A+^X>Q#X+@-#=ATJZ_>$O7782;=+>Z<"%U3('U]<V@"P
P0&GBZ!7>Y/SM]&N9BBPUKO]"9$TUG"(&"7R4?2DQ.*=>V8I3?O4H8AAA&- @ PPB
PP3*ZFJE@COK(=<K3=0>9U>15%Y4&]2ZURGSKYYO2+ M0.>YNU.FWG'.CF/C<U$D^
P*B^B$1SAR.W7@'I/RD"JYN&'&=\[)[UL@"^&CBE- +C_FP%>2I&.RMQ$L?GW&1<2
P!AL;>E(C,RBLBGVBX7)R&X='BPD']0:S6'<AGX=6N/ WI_K]CY8\&-E\]D^ETW%N
P+\W[N\Z+/ /&EKU<N\'P<F^"N5""V"X;A[A9I8T_*NM6EH9W;8B>_%6?D981,<N/
P'IDA)@+Y+U,0OMD$586M0%1J.++:O,)<LHKOWLX06\5L$6+80G/)(=%Y"T%:2G/_
P<2]K>WB<=_SDU4.C8P$7L< +I(XD)E.YL@WJT[$UXK K[7IV&3E/":OB;LDPYHP/
PU,WW@_C_1?C?^!XYNPF#D0M?KHO/\QV_HTL)>N85DP<(><"[32F"U*H_=S"*02J7
P \'_?V6F[%S^NO0LD)&%/Z-UNKWOC),@Z4MZAS)+Z<8-(3+]=*CH#;9HB1XZ<H(Y
P W96>G787 3@2R5ZY_,8BR!E86;6T+K.I0#(X+C?G,R7J.>*24 8<]/<N1AH9:7-
PIF.L/#Q<JFB-9W%7YE$56600KQ _N8Z#AG1,XC2P8M5C5$)5V:92$LYVM"8! Q(?
P[]P.?R-5F;=LLVKH?TX?IG,WBR9:YS!*70-1BVS)WE:7Z/5<?\IKPP#Y:;>AZNN#
PM=4XO5"T8^E/@9C B?BB7(TMFZ8/1B=7 KIJ:V\;D5LT/OQE,>NN[%1'LDY3= ''
P*=3M??K3&QV-L73%E0&H OQDQFZ\_:[2R]K<XYVJ1ME_.3]K82L@H*F];R228]6R
PHM3<6$^L+KV_,UKT=OHBT"_#.L&V.V]CJP7_9VMB#0)Z.+,/%;2X47D210>NRE[S
P5RM)?GF%H"6TY?AQ B0$MSB>]DN'"MGE[JQ*+,I&_<5=Q2DG_HO5?C>AT6+;ZR(B
P3B)V](.\AB>CL.MX:4$ _6UJG"1]I>XOOS+*X4S-!'Z8H2!5:6C.A^WB?F 6E6L_
P&O< 2MIZ8!HG&696EM)*D0+\,B],(1\E1U=H;TU;<IJ:>!V$0&>TWL*8$DM_QF]-
P_A!@CRIXF>T$?]C#Y^ V<?_X;?]>,>C^JK:WNK\W%E=P(%Q('8]*:^:&O_PQ@S5"
PWS@:01W+-E37I+#?:MX-UP-.=%RR]HIR$<@3VV0K=JA<J<*MHT\$6NS-/SC4BQKY
PG,Q"9$,5):@1'<>\#NF;!/P 9FSKG5NY:?I?GS1.M;5P>G$3R )USHJN>G.FN3\&
P,CTV&>V><6D?2@^X>+N85C70;%\OV16^[?.A"NM4@"Y4^&9<;[_9O::H #-TS:(=
P5HC.\@<HW0-G%6=70@AO=O&Z@1"8IT:S_Y=%0-*63L<MB8(R" @)'DJ>L66@C=XE
P4.S,G_BA$1XF-Y/[)DDYDBU 4WP?^5XFN@:F])V[0)<F.E69@B?E@BK^\E%2.%:Y
PB@Z$VT"I?R*OVY7X->7]O_'C%D?A_E[#+,[F!+/&RF!ME5]">.-8^6? V1W.\)JC
P+7%C(;L7TY]I[XA@H1T3CCI*M><VH4>Y5MIWD[I/6(S\;G.L]Y9NV6>5?P1K14>_
PV8;-LNT@,G7/7X1#YZ3'^?5=W/#8K0S)$J7B"%>50^^O#F#'\-QM+%-#LC).&)DP
P0+S@WV;$W^:!>X>#F)0!38;M*"P'(6>(-7MS_PV-H3BNP6I?Z>?LDWGC\,7)_6)3
P%K9*(+5Q! ')#P\ DW2#V=MJF&G"B&+BJ#7Y^TYF2&^@GFFN6CJ<K-IMEKUI3E #
P^IF?/+Y/DQYAP6K&?G59D3;C-X.Z%QR/R#:(A&5T>BYQ+(';K+>4F8M9[:6,!V>L
POV1TY ?NJ KX#YMT=<N+D<:O;,,18E7NR>P:30+.J%<1<;,0A*BSC#$T''.8"=X!
PJ:OS6?L1J\&QH@-^UF/15OYD&"B,(8M!QS';)E:"6'VIH>,L-V)5$TOQDDC\34$T
P9\##ELD-4NV%5LC-FYP2HT,*'IQ0X$.O>N>ZXNQM'O-HXZK;)'BN7^[8#T,RTG6G
PL:DKC:CT#I]Q\G!V0%NA=;.&TVR'PLAU]#]IB";3%U1JH0:H4)V,O?W%,B@\56Z2
P."%G#68-$N,%.%J'6]\0?_575N"0Z+X(^/D'DP:-_@)4Q2-!J##^+G,]E?MR'9)D
PEY\L27',R8FM>9_+\'L-Y_0C2(["&@.ISZA%8XKHBH!%'V,3>VV-$U_Y8D_%,<0?
P'%+L"2/=,(%F$2F]^_?%,3TEA70QQ78VQ[:<5U8QUZX3"T]"&!SUT26S9WZ!Y8->
P>O]C=]K,02V"ZUFLSR3R/QEWUA?>9 +T%$8CWJX57<J@/W">.B"?@.+;10HRKL<4
PGO)J+95D2*JUGJ0K.SK>[W"\V.,27)\;$5B%-P6 <K![8Z8E89QM#$E6^HJE$9"X
P-$U'Y40JO"GK,%7YM;@2\JV=(V)-<E@3MV 5ZIC5\9=!-D4=I0>II?<EY"[ZY$Z)
PEYZV9[*VAOK6^%J&RIQ)+T*I-HU1>'M"" GUM+C,Z>&M7%FDDV+I(]8%V!6M]/@$
P5,;T+&=^/ /FA18'OC2:U)2;<O%JH!EL *6RK\$B;R \>)GA!-V]JFW!K'E$'7E+
PSJIP4=<OX+66M?I;+/"[,NW?X:3]FH4);IX1L!J !F;69ZH%:\J5"<E_0]]=WD5U
P39E77*O^4QJ74)#/I107'J_GA.+9VA V)IC[BML9!M]&44#12A599W41_:!X*KQH
P_J],CSR7,(?)YGMAMCMI8BS1I8P^W565@04\>-YU3R\%JP&LU?>/%0.6]9VNWL$)
PR+':S_FUR,04K9(E"$ZU4D=9<4<K='-&WLYQ +M.)]3@8E[(B&RMS:23N(EONE9-
P?IA9GPYZYR=3QI-&#4UG2,>^DB CIOQC44PCH$%<4:79#.G"4[$8K)VYBO*J6L[U
PGKR7QRZJFN(P[.UR-Y1DP(OB?[-<F]7Z\ADU/_Z%3@@7>%<JM9?IQ>LZYN/H6<UD
P('K,GS^>*RA)U4U\:2\@8IVI?A6^4TV"(?)#L"=L.<M<$'V1SGR\W&"HFOC&=,.=
PW3CDF#1(3EB:%&.-"MEH=F2/T2B3]\X=SL)XOG6ZIWEBW;2$>>4_I;\"7!Y2KXOT
PHR?,'!"T+O/N*["(CC)70A3R7O0]8%P%.NP IC*T3FI="-2%=_0G=86?>9G8L4=3
P=A[Y@<L<5LX"P>G%!8\>6!/5Y.B!4E4%KTH26KF_D9H2DSQQT6<@SW&4\2U&W<\%
P+9"A(-E>+I#&F2"^G@FM2*LEC]&YN3F/"S$:JL&*RDB^VB&P>N6%ZB(ZE=027H"K
P,WS?YX92,]8)V]3Y.^[S!*;EY-,7%/?XN:10+X )8IQ:&9X_P)&8O[:I/>_$7Y*:
P##&W^8S^5R?*U^(M$>U@90??=K%5HH#_L$-FWO#XQ72Z#-79QZV$ADXOF4Y0@:AD
P<1]!]D PN0G$#R>QDFW2T 739DKM#C #(JX*/W5#W= TQ_72U"M(7O#]MO+$/#):
PS-,/Y%Q09EV)['@CN^MS&*H28BOJ%<@%9LWP%A=XWE.JK.?_X8^51*["R*<^X%YU
P K/M07K]SN%(R(#LQH>P_:>4MH(P&OG(Q+.]E ?H%U_EL+F./95#+R0.](^XF=C,
P94C.&SD&DW52?M!<,BY$\+%C&4#-8WX\3D*JI,>PXVZT^U+R07AF;1=18<3S#!K.
PVF7<@+$(IZK?2PWY[2D!YH;Q')B,PDW3+N/KJD&?3)[3QJR$:=J$,Y9#:'SD9'2[
PDTD%*C4ESB'_-*XH>TPS&H*,2DFJ-!1):"-J.Y<0D>.KNRZ=GJBP\K)K+1JD2R5>
PTP!*@*P?MW$B?CELDJKB*CZ]=+)H_V/6X[:P,:( /YUB1 %C;X'"560,*,85=OFM
PM++#X&375DS2+IY+DE%/9,L8'OB+=.S-7P+(J"R(6\[VOX$J,:K<1,=9WU\]C8N$
P^ SJ>F"QK5,[L._10*4BWPEM-?<:_L2A+5X-SA-*5)PG3F0X6->2.+EL$IZ=73*-
P_?S$**T.'=?TR'5!Y3UD90L=QQZ332S%*?JC^\R5EXEZ5VNU;6>F&+K[5'ZUI/EA
PQ&<P.)0,(:&KBB*0A8YOO[A.F_J8/4)SL?FP&)PA!OQ6 SM3HFYJ+)BT-_/>L'MG
PZK3S,KOEK@*!A+05N""Q)H..:MTK9Q<H,SAG8TVI'7D]1=@GQ/(@N C3_XWYP"T+
P'T%B7B=SNAN67:G^@1GCVHGY7N&*CVZJ!Z/,DOYR%0B/[)'^G!'V^0YCCE0)4P=(
PQ'-PH1FHE%"='K?^.,O7^:HM>YNODSCM(>3*@O0>+&DA7T/-HJ81#)K@7!=T+WOF
PN8'PR KN2JD*G%JZEE?AN:D#(/T-^'".F/C4(83M=A[]QJ%VS"[O5AYI\"<]R['H
PN%H=*H$]AT/?L.9@>(T;WG-^C=9Q$U8+53[>4J*%MM$SIFU(Y)0 PHL(W@N5S!-.
P\?<I',)'!YH+N8IKJ'-SXCF15/^85WP5.^B'A6/+3^1AO1>"[>EZ#0JCOK_&RUJJ
P_+/EC7=S.'%QZ1S,(8...<>-"\&I4P ]#"];&A"8C19'PDMUF49X8B9VD'#CGKD[
P>DC.G8GGZI"4Y"#Y^LGL#G%(8M@9)./QLJ"(/W93NU'>H1YE(,JUORM5.G_5!!V 
PK29KUEKWV4=U (Q$QZC0N5HWK<W;5O$ (IL)?R47U$K[/#6%:*'"WMH )V$!/L;L
PIO.U;'#KC(3J3RQB/++*:ADGXHF*EQS14GXD-MVCUQ-CJ44;B^>1*U2<4HOT0*R-
PPVH]X BK44&AH7?NPKS\7H --Z6RW^3^#AQ+&DY5UV^TE@=E;75MOH9GH5VZ#U*(
P\<K\6 4GE;A?% H^R;N=[BB;>U4:=91K)]:KM5A='&,.N3@/O'@2P=CR(_G(4PV7
P.;[7;^WIM'AE%A<,IM!Q>@,ZRP/WZIOBRBR$.=97I'"JH*FQA+U&VJXI7^I:LQ13
P,E05U \W3,%*BY_UP%X\A>,;6^,3:E:-^3(%(K@L77R ,%C;XT.Q<0_N6Y2UIA1H
PSYF;J*M'U@+-@5VB%0I'U<TQ/WE:Y#Z#K&AU>S!X+;6KD/LRBGLD4IG%."^H<=F2
PH:_Z_5324PG39Y"5V99V9V$4MJ.[1N,*?_,6Q?%./%E_ID61QJ1*)JE%ZYX)V@J&
P3.IBM(@C>W''G&RJI,LS<,<\7C&  EP+\_J#56WU@]ITV; 1PS1+H ZL6039CQ_B
P)SGU$")L,B//2!(O-_7D4!0OGB8-RA-Q)I8P&IBPG'3542-F@=;'CX!I!.#5U-\=
P\_#HCK&&3#^_/-RZ(0O/70/[! =S=\55:2K#<HXY("X0,=KB+=,A[;/"#-VZFQ)'
PJD*":T Q\+Z$\ M%: ^<Z+X;J7Z$CHP>7OISLLQ?-3.^[\+Y;G?>O+@KKVEHQZ&T
P--L&?D"[P^\<&')V19IB&GA8[YG;#]L8H-'R$WD].Z,[)^>&"S]D@X/1#N#1 XH_
PGCD+QKBF*Z#M'99,Q"_>.^[[$4"@47B;7,**U1?I7+@EEPA5K:@NKOLJ<#BEY8NP
P*G]]\!C:VOE(E,(,W08LT\_#4:G8AX "N*._0STJ?Q[#J"2#)Y>NT(?"0MMNYT<N
PJ^UC"R.H;)K88*6VRZD0*"-"$+IN4H)4^3++FB>L"N)T,]NJ"T\=?<D9:>%83CJR
P4Q%W8CAY#_ZG3ZLU['?^IM G[47\W/^:O'!A'@:$] 8O"16OB(+[PBHH(NMG'X&Y
P<<U2WMV\]+U[=:/Z+. *%+6^Q5%[\(F8[@]*[#AD)\A2%N_0CUQ&-Y;6U_3-'=8H
PHH28EP;':<.DN!^VT397T#$S<WCXM$*S90QM-F\C(+6%P\2V.I\U'CYH&08'X4#=
P.Y+'0GXBCG#!=59I6UF6=47GU2;]*)OQ'SU%WLD$,0T00@>X7/!)BI8>7XM/5_O4
`endprotected128

////////////////////////////////////////////////////////////////////////////////////////////////////////////


`protected128
PDU7H_H3X>>IRR,/N?KT7T<0-(GPPGNX7S)K2O6232&=Z/G(,-RG>ZRZJA ?<O-9I
PD!&DT(D#(YO2QL-LJ>1$X<%&MO@^+6%XNO#N516ME]N-_.3:092 V2^,I3\SG,"F
PBLH!WUU]>XD<"@6 0(FOGP=2[L(7<96^GX3.RYJ)V&'NL#)1OV^9[@FAL39@"G!M
P5+]_#;^0JE,; I':[>O.&FSU*1#>@42-^DYC<I!%$!0\-_GEPVT-T701"HCJTK^H
PRO$&'#FMHEW%327F;_)97)*9E18R755 "YDLL>9/2")'>?N1.A7KP*\.*;Z?,CUE
P>._1,>$BT7YL2$C4UX\;JVANO?M(E\.5M\5_0^(_F6%/;;T:!*KLKF:DK XC[IGZ
PSG;'42'4M,^+2[6<]0?]P-QS5C1I%J#U^U_/@7]B'3+P\B]%;RY;V+R!V4V>#7IH
PB7?"@:9<1X2%@6/@!;.Q0(*->A.:K'+7(E+<ZF?0JRT1"0;18%Z*8;W)@^S$KYP'
P*/-#C+]Z_PJX'-8.Y,:A!*?AN7+%P6]2/LK?.ERF,1G9_\UK)4$Y:A#I'2['5HPB
PTJ*M&*VO&F_ T>^;47NDZI#'QLCXO!"E(_)J7JT[9 ;?6&+^&5'68U3Q3*7;MU@V
P&]O1M^"W39ZW\Y\7#)I<#7N_[1%8Y,EX@QA7=7>69G/)Z"GUX S=M9%UMW0):VH-
PAT[R9[M31Q&8>784P5 5F"^2S)U+>'#'C[WUZXW"+[H0_-QS.PO+; ]8(IK5=H;:
P1E+SRI-<?TKYP':K=$15&S,O6PKM6X3M/B_:U^N+IL,8: #852QT=)I@^N,]@T1#
PM,_-T*&?0NFV)5#W"4/+T7<741N_TZ\JY5EMGGIFH& )& !-1/2Q&",#/ <_7/8\
PP<RJ0=_^Q<B4)C>(,NL0UC'Y  CZR&U6LNOHWE6O^"0>2?>E@.P;-C9E0+K^$8\+
P,,F-TE%+<;XE$CYM^@@<^11PJFB(BX"_'ISNJ<XE]89S&S3E\TF,:+4]BVB\<U/#
P\U&.[I5VD:'N+3<Z3+I*\:KT$K38_5U892@\  "<U;)H>OR]>&%(XCM=EX'O;6KQ
PU8@D#'C,%X3HE> W*D?2A*^,DOE^)L%E/X?D??2@XS"_DTQ"'C8(/^@G<T=(@;"1
PE(Y0)5N%NJ(<-Z#O>3%[?!0]I@#06N"_-"A1OO1A76SIM.<T.T$&0X.WCC,]2V;/
PTTL47OFXZ+5;LK1G%W$LL#'>O\S0ZK\#5M@%Q,_$Z=+XG>N_]#XW(="B)!;TZX)K
P/I'.DRG'!X[ ^D4,@B9[!*GN=C+"N.B#!FU([[><'6R6G]V;IRT13]FREX?+ '(?
P;'D"4J(\;X WR F=(PTMG:!N]*>>?0$"S=!A(0 P?=(E$[3)%]'@..?Y!ETSS/$3
P_:3!S?N=M!.*F[I@NE./M!?"V$)@C$WQN7#.0F6TQ9#;]T'V+KG\8==5]Y=ZV63_
P9N1"9G;9_+GX[G0I#B9@9AQU4&"K-]R\00'OD]A%\B8GZ/8$O#3FMF[_#9NQCV=!
P7:4<\7)#X%O_Y(2-<)]A<NA[!M38Q$NO3<L*Y=B(+]^6H@0QYFV&O+#Q>8$4L2?G
PK8J$"D$M!I@.AY82AH _82(N,O[5!^QRU/PY__>H"!QM2)AO>>2"8X .DA48!\2F
P&%>,9PYA$!$OP$./J:#C33-N92B82-/ITB5UDY<@2YNJ+FCBT;Q9^!<POJTBQVQI
P1/5<7_Z; T;):Z46C@G$B=2N?JS/?A+H2%\#?A.4]G[JTXSA%,U\U4UQ1?U[3V1M
P[MF>5'?J&'_NG^.Q5<[Y:"VJ)JPYMO%KULH+/:2++Q\J30E]P;K8@#B+'*R!3.8J
PI#O>\TB3Q :U41T!NC^:O=!A,H(X)(MZ4/U7H.DI.U;V%XCY]L$7T).B%HTHW;25
P;./A,#'A_\QD,@1UF8\Z[A07F^,3[T:IK$C4=KLZ@79^46JKVPC*C]+%T1R!<]6X
P 31+4K QJK<2H%&.1^(Y_0PXTD_R!O4\ "KDG)B,_YG[IX=!G%NX[_NF7A^JD]G4
PF-LQK;@)'10*HQL\@>OY8#XFM'>!\YA]2;6)/\\3*2I&*$KJ4<9,7]09:)=U"DNB
P.UGZ<E&*9Y%#O)=B0!H)9GK'\X,1Y/Z.W583N0)WKY):CD#O1L.<"A,V'J0$SH7U
P+X"QW F-X@NB\8R+"A+],&VY>]&43%P<:_E2Q\P(K/JY=.9L5_]PHT*#E.MG]139
PKG)\1AD_#2U&%:0<);WO TZ(]C%+9M9V\;'I33_^<\>0/S;7[X+1-#^[:.55YQA'
P(:5^R\&=&\<;KPKEN.(#0:&9\6E_^3@4^%8=,P_^SF-WP<HK^M64D'(&!.T07</Q
P="F:& "/PLI^)&&FCVF*;D :7O\"M4O,0W@=&M>U'3_%PLQXLA]#PA_)=N].83,C
PXOTF\M G[*9'9;]WT&N2^8\CA-$Y<R*RT6\+DA0L*(GK>")4%/M1UR>8R93Q0P)O
PWM!SUHZ--Y&E%WBU7&IT8AJ? 159HVE0R@>^/[K\<GEM!'5:9?4%-\>?43<S!$C&
PHW<:SXTMEKW%/G"4#V;QG,_/IZ[V&*:&Y,R*RXBMYP"V>25V2FCSD/2F))*2QY"R
PN$>RUPV@8,90,G;6V]8+=\Z4H>BF1XT2%D?,#-;,M%/$7<SCWW%BK2?34^/G=O9G
P<3!ZJQ<X]@89_SD)FZ?XA!&L+46 G^]1GX1!PV?R#GDOB<VD\K-$\:BY3TI)C@:3
P+NZ4> 5?F @-)-_'IK:4,_^I/GSVOM8@>@>('.+?*U^_%J'E JM-R[,:Z\Q!JRXI
PIZ3$N;Y"IV:SCMS87Q/2W&A8S##QOB?&,E$+L8.G634)5$M,)'2G)C*%<AVHO]C#
P?ZAI?Q1!$"8TQH@]7YM@OVZ@CN V1.QQK:A>72/'?='&5_O5 '9INQ;<O:4H!#\ 
P:8%6\6/&K.+O<\C+L66>@KVWP#';QPB1C:'1&TEP+8#S7 Y,-*T'M NPEV)U0N1:
PQ%WT\#1FU^EXX>M_K#/;1G/9V7Q\=XK#?Q?QLTRJ@G+8>3K,1N=]-8V^F>J%L2<4
P&&YFD-QN3!VB;+!22&!F)3QR,+1 ON7C6_I(_5[5#8HO#EYS8S?5>JF X@[7(Z=-
PUMJ YDJWS7@;"%Y:AZJ\Z?%;<FSU[BB ),WN@Z/#\Y8G6532DL#R_RVK6VT"Q#H[
PBLD1MUYE]%B>N]3>Q"%S 63:C7EJ!"?F@K[D*PMDI=Y'S"<8E^O*V?(_XOYW^FAE
PYE\PD/G:%CCME[V5:&:'.'H5T^#P6*1JL+)ZO3-1O&PU8 PMF@TX*^)()I<,7#5$
P8Y%*< 80>.N9CNLHH81K3FZYF,"2##P@9^#'"%/67CJY.:(FR(-IA8^<N-A^<&<*
P1AHWVRU_4*-+$E)S)OG6%J6U'SI^4K!&YK7#$" ,F1#!JT-]I*4-3Q.^R\?>-[O2
PS%^Z+][5;NR2PX$@LF0H%Z$;7$Y4R-/+@]LSF57^W\$D1?T P25X;9PD8V/^3*M.
P3OMNN)T.YQ&<2E<IGA2E; !I3;,%3,=E0'VBN>6-VFH\J,[O*&W:=MH2$<(%-A4N
P,C>!3Q\(_N%F6! ]=1*<@F&,T;>Q_$%Q.F Z'_O>JX< +<D5)\RJRH FJ=, .@=*
P:(T.7/06J_GU().]T0 >&B%X'PP]VRUVLFKD6=P4I_,4%P)0%3C"A6(9YU8]/X64
P"^F "ST,,+K'984%/DS/(F_H=PK+-I;R:T%W%LZ.Q_<#])1* J[NI0=X2LVC@BZM
PIPHWLY\(6F8R/TV=:_.UL$&4$K2]IG!A9$4P-C^'(K7YDDP_?^=>FXK&_4TX9G@>
P+W9&"1(P*-6*_%,*^G9L3P7]$@3K0!#0%DS-Y='PBJ@9T^:.)YU=9K??VU_KS"*$
P'*24WF6500I--,Y>PRAQ;HQU'"-;TK$8"'S/79QMZVJN+S ?"[!H-*?["LQ&'PI>
P2C@]V;<S+TF3*!/ .BM%_A\(&S1^. 2T!\/>P3-SH5@KG^&DT;?#:#S$O8&&^Y+H
PPP0ELJ*L%2!3D(*%&$8*G:;\?X"7!A)/T)WRX@%40J6!<? MP=A"#S.KMM/BEK(/
P0[.^B94T;C<!)ZE QAATVF/X:9Q"=ZB8>2S'?_0-K4K2BV7_3E08_24@SKTXT YY
P-3D$#1S2Y.%S]2!G-['EZ);@:XY+"!;F*?.XW!3FV"QUK5G,R.A$<J5V%LW-H-!S
P!"B>/[CZDGDAFP[,;UT(\&T#]2Q7@(['*%".I?[%#F[:RH'RAB ]$_U<#6/,,1-V
PZ%$(B5EGFFT'H,B)<XL$/4<P;AIH<3YBA6@W]\BZ*R\%2K+L$],Y$&ZO"*);U"-J
P1,\#ME5;4=7:7_[M['V0&/ELE8):Y /8*/T2T_+WW\?XX GP%M%ASM>",X:$0%+1
P%0P39J$L0_'$U0*PLSE)NU@5$$MPBD@[DV1D!Q! I9?^\8YC:57GNCG@G>CD !?2
P,?*PU;<EP2)3M:?\K@FFY?M8R';WA(/'P%4DF<=><BO368IY@9)DN5Q/=8]/JE6;
PVQZQJ\2K#-'!Y$-D25@4?:B'D,\$42P9KT?@]\))M8._$>P\Q++^Y,EPI^4@3IHU
PYVYUS"09T#/R;2<@!1_]LU]D]G.:04Z!R7#)<6MP'CEE1*> A2S:;??#*)0;A#Q_
PJRZ=0E?*TEJ['37[D_I8DJ6+D,Y@O7[MQ2\V%]*:%D8CZQ_-I>:6P^^T?%G_<.P^
P('HI97J5,/;OZY,*+5'002-"9#I&+-UKF+LPG&L#R_U2]='.Y!&O6Y//\OGM-\2_
PA5,1DW[[@4)DZBYB[A8'CZF0M>,/B6=P";!W[7$/&MP_8<E*]0*) RL@R@SH&7N?
P7M[S:15K9Z_Z2OD,8"'%?RA_I3 S/"# ;FYARO$0A*]HKZL55N$>2OY]C?\/M;JK
P\L@7FP;L3W#;=N#=26N3X\\+Z>M" +8)+.'NBWZ<1*_?SS_<^[?C\\?00!:28T3*
P-!S9S!08P#;[# I?X*W, 9/4YXS'''T+"L3P[H/Z'<T ;?N_Y9@/%95"7PX-'7Q#
P#BGTG@/;RSGZ!+Q$[2OTW>"[J_[9V?^QA $4Y7D&#M-!V,SV/&0&P2O*?ZCL(="W
P8_X;?R?BUO/YO 2QPR7VD C55K/];G\FAW'#8[;#LRHV"_-GVH<<3Y%9J!<L,R1C
PX+=<*&:=Y[)8I6 2K7ROY>:H:GG)VYM,\,0@M\6 L";FB3'\GI8)OT@6RXW^BQG/
P:\3JRDN-I>&5SG[JR7S%D(<M*:Z(U 69_HD$:)$9/S+.Z&PGX^:>'TMFY-1] (8E
P"1^S!,2AK]6#3QNC+S-?'=EH7NC8MYUY#48_'<YIJ)_7[DL^+*0$WU.[;11N$WE5
P=P?'LZ&)IP:F_%B_4OXNP-X9Z'&T\FXA[G#5U5H:PV<WGFSZ-11Z,Q6\!_ZP @M%
P&:-E$09)7RU'(G!_LC7>IQA0&4+$FGSR6R(!K-_S3VBD/%!PR"I3O'KA<WY]6/9I
PMY1>5G0]B]-;\)#0)A(Y=XRX^@K<6/PP7XM(2A;3HZ_E9E$XR:ZK#P\*"P](I>;\
PF>C*/<"WN%CH5M9:XEU>/N&#&O2HW>1)#EYP2)"HIK72H()<Y<D#B^/#-X9_*'BK
PJ%4:&1B7U 5?A!8)5-GC% $%VCVTC,WC+&[0 6B963!LY(8 GYB5T?\,*%UN-$D1
P]N'R0P)QVN8%Q)6D5?AE27@45S&BZID564XH/B8!!=EAB?HDE!*UA+T'\RHX$ZZI
P;:EW"(D59$8BYIR%ANY$G1:2@=$X?W;EEYM?+9?'C\@M3_\AC%ZJP'&IY?% 4Q1W
P$   <6/!.3ZBOV(?MS49(ZG&J733U_@I.9&1@AWZ)R1:;I(D.?5PZ<[[HP,G0,.K
P,1YPPS?K%/9JZ&#8WQ[P$8R8]YH/#+L*7T\5D%_7 )UVR"&>9S1T-:+NDAJRIRJ4
PZM[25X*R<>'JP[L"1();1*SY<9!N%HIC9_+"L554R4!_CYVK8JO^]O]IQKE?GET'
P9P1GN.BSAJ-M+5P=53RIA4[_"@LB'_5!HO\/*UT $?VO667SK!+&*?V^7M>*S3[[
PI1]/_%K%+/">B)=K'8[W4&+#\$J,]L3Q]=Z_3$C>&1^8'-"B=%=6Y7K>]5PTO(1"
P/-FQH>8^'%^<;"*:!9ZL)AG@HJ9#MK"9^\&"Q+C]YS]7PZ=\?*S2\VHW0UY63J 0
P=X?>QPVX'+*$NB.X%L==$[(@*RR)<=!8\(T:W7V"+W0I7PY4'GMH^0O8<ZRRQ0=&
PY+#>D9BN@:%?1>D>7.D#62^Q>=9EM+^J\4-+<0X<=Q BM\# S"E 5@\?8.QZ>CG%
P6T,SOKMKR=5"]#IC^[)2+ \3 8H-;XKL+M_!$([GEU=V@E2\%IU7+'S-:B9$HJ,=
PF;! 7A2@\6*&8&RI5I7+%I4^3AG^Q,/^6D;HZZA^YSPSVG6T)X4DWL/%PF5[T4YX
P%Z>;QH@%J;T621AE.?$(48=M"DG<7K8AQBZE&L4G'55NZ9IH9MQ@X]W'MTRUXB*^
P.3C!('TFQX[> 91$*I:>=Q@!9F^'X21=6O9U1EZ)&Z.'.AV.(7+3PT>O$.=I8&I.
PID_H_)OS3B-Z3(>CVO);0[6;>(Y9#,,N3>3I$+7-]_&)6)+IX/0M(E98G8=C,LMV
PB0+$%@*S$1WSI@SW&(]88N/O]@\1 H8?K_M@JY18Z[KD:GK"[[T]N'C>FP@GI>5,
P9@E1BS D%&*:R[2]9OWK)#[G\+@EKY8W0*N:&P16U=;(\8*\_(NSKT$6&2&7OFOK
PX2KP>J?BD4B51\,--$'HFFO ^J?(=ZFLZA6G.*P[Y(]<6UG%,57N$&?C]P7<_EG"
P\-637'XR-#GO0T.-OJ*67F#'@D,O[F6MJ[3\VBO'F(*L&'IS4<T$PY8TUZL*L/9.
PI56<QTDP5\YW*<UT3>;K"8;9XFL?Y<N4"JM,+N:SH'QWF]]T%#JO%J;FD@PH?:2M
PQUX JP DX7SI&V]'9+O\J_ A+.]#?X^I&$Z,BKWG\9Q];(&%Z[L^DTL%I>RK[.<;
PZX57GG7J*N_QY2R7R4B,J-EHKE@AW!:EM %^3AO&&+Y2V0&:#XJ +5,IP7U9+_1V
PS\X117/;^9*)[&BBYI<T82+&Q:?WW[,U2E4H<T_Z2!C+D@X!L:NN_6(_V P _K%A
P..G!/BD1>!(P\^1]+$EKVH[MZS?V8P==B"X(VL+=N7F<2]#]8]T%4@+7JY3[RGJ5
P"#\O#W*S(OJ!<HL(C&FF6.CR1B0!,OX"SIU.,?F[##NZ8AN6%"ZO,@'LXURO0N6<
P:G4L:T<%C7E2#5*74E;JO?6Y9SIDG9".1]W,NO[$=T\WZ@,B' B7E>2N4";28X>6
P'\\;)'Q=NTFO*FH;XT=:46O%?\]L#X*3M3XP4EQI?V4Z&_[S4*ZF<T=8'?F?FT;L
P-K"C>30!()IX!M0B%M1K=K3\;ZXN0OB -\ 6R-$@390 F;)B9K2YF*<Z0CUB]UQ@
P)*AIGS!%_AF%Z/58HHJ<SXG@ IZ$(#"7K4T=(@U_W4_2W.6F3<Y0<N2O>'-51MU3
PR%KS;@\',SUTG0IHK,Y$!.)?QB21CS!>D3ZDL)88(=B3<[[S!T A?<-50I1]>Y>=
P-!!B5NOKI)J240X_]21QMM7=3B31J@"12:/B.4[IMNO2#S\J"+U665C_6D/@PL-M
P$>5[K29)\G1C:/<&,@H.5K8Y^%=[!WH!R).U<^AM=-QD%/&*?E29O(4T$W &KR7I
P]PX^:SO%OT1U^^W(X^MO-^C-.@/&QYFS27G %'($>[@(TX+5O!--?NRB3-$L3KPK
PD!A_18;IO.H+D(S1^39&(4X-47&CVJ7.U7X:Y@Q?<%(B/TR-_9@'+>DQUQ*YD3YP
P$)6C^-XS.@_7Q)[OVP"_W"SYWGS$@"Q>ES@>RPN3$*8RAPX6T7?@A)^A "9H24D?
P V&J1\OLW$"I'U%_-,0(D SSH*W 1O4KIL96A-\K>?>P;VYBOO'(2H3@?'7%?+7+
P;/,/-WWWFII:3\L'J]^HMV+#9Z$J+$X9S3UQ<:X-A&#NA#V&69%%E88B-Q6J*^##
P4AVG9^^^M;F"<J9T:T*=)_#8+[=:#;AE0^8#WY^B%C.^#CXL-OK$:&>][5^PR&'_
P=4"D":DQW]P]]<J8-X173'-_F\Y==*RWHV7EBCZFO,ZZC4>5(S<N^URBTJ%&.%/*
PNFRF7*-#'5B5IQ?"*P'G'[\(!XOQ#JO#U&7>#4%^#M8BQR^,R/PGD/V6UU:(';: 
PI2N/H @P\_P)UL.1>)UW[]6.:ZD:="\Q&KE]^\KQP72>NB!:7$1[*ZK!F#Q=BVQ$
PQW7AC*8'!Z[3L*O<#;1_*TSHI[3/L.2-B%-8S2&7"92(M)X)'ULT*Q.:Y"KR6,&V
PBWRW#MM=/M9;964$OTW$MH]'W^DH7<?9IGHA$-_S3R"#6,RX"3+ A8M $8)P5AX=
PGN49MEX(J&.;7YZ[IA#(I>6PK2 8L$5M+'Q):6S1Z"_[Z!(MX$V_7D:RO,U:Y414
PN!0:U@I<3C45GA_4W8[E:<'SNOL!ENB3[B4VK\+.&-:''/ T\C _NOTT^LK&M.'4
P2<J@4H+[,PI6*9GG=<O07),=+IE)7@J6B^MAUR?NO$E]FZ;$UBOJ2F7GZO5.?#L>
P,8QQ- B.=<X&(F2P_X+<G4-G0ZB)<BTLV8K*'.V)PZ J\[(2AI(,.G<*03%/$!%D
PR87#@G%= ^4]NA/?W#?Z1[6]>>;8PNOG'HDLB#@-4-9=' ],@*+S6Q8>-]=!]&N;
P"*"VJ*>YUVD4V,4PG>?!R>L<&4N!#7 !>K(H6/!8HE)KJJ]8$!C97*L!9W2'[)=Y
P>_N\8]IZ<(&\W98>9]G #8X7O0*F^B>!@J9-?%N&)C/'3&Q*[T9G_=!)8?Z2E TE
P'B.&F.7^[O=Z?VCB\ZBK_RUY&>'43XF!,"T0#F:KS1"%,4T*XJPAZ//LVD.O'?D\
P K[Y>]![8\IB6>%N_\^5$R@24P"9'VTZ/ 4Y? AHI TTFS0!X^"\+U5%'/-J3T*T
P1VP+ %?-Y3'E@WY'1S?;)0LAT[F&VD*?$@H"-0U_F'?-7%ZCRPZG@=@RCC])3LY-
PRR^3N$+K$X\A"@;&3B609?/OS3@>VE',BN%\H*;8L2#$$?8%[89"00UT1!O\3,OW
PPYN./@P<P&8>))NTZPA]D)88M(JG.86*/5ADY<ACC],15FO/20IMHO#RVXRHI/-*
PN.-?5AY4H?+,2>%G_@\ZZ9]@/A=1U.5\'$M<L=$VKSQCY_;U->25H1*Q@&N)!DJI
PQ 58+6QBY>7IX=2!.57<O3$N805W?>&JQ0;USC-(P-G_EO W _K81 +>6ZSQCC[R
P:V7DL7]13BZ$]LU0N>' )!):^M2(NQ=1KF4_L<.""E/S&6M[IJ9U52[/5I^##LR.
P^CFX0-L&73X[(AE2:1 #3KQ%B:Z4LW/OB.E#PX9D6F#Z)QV:NL0+[&U3G$TN@-BE
P8&\R"ZI2)(:\9]W$]UL"4>"!5[5M;OR=23A7]6MF CZR@L*>IS2J1_. 6W$R?;!,
P5Z**]&^\OE^0 V5M!0->Y?@.2=V%,(_S_Q=E!^:07^\GBR(Z0XU/\:?STO#"^D1V
P%SK$TVA;4)PKOF&'/-%.=@BNE61#H)^04"84H,G$7!VP'RA]GOKHYCX>,M(&4K+ 
P@Z_,VEAZ9JDSUWMFU+6RM6 O;LOU"I>(Z;U&E%]HRF(@=13+"XR?,]G&.F&6I5_Q
P"4P!D5VEYTUPSW59[5%?>EQYQS- >)=/)M^D,U5/-56G/[<B_XOXM_P.9()>?J2*
P4Z1$CX]:II',O'ZKO^L9%_]\+6QIX5:%?GI=01=][*#IJQ<B0 P<[.FXN$. NSO)
PDITA;1'*,59X+D.\1IO68K56\B6!;IZY"TKB!S3=XZ<1^ZIZ^0'@G9UX[FQ% +(7
P,OI63-%QE89/0".T,2_FQO5;#;0EQ D+OV:O?RC)[BB&T/"?&K-Z)4UH,4-FJ(SC
P?-%0G*%;9-6\N4,@;B2! 6.NY6K U8V074T,Z/<T#VODR?V$Y'B]LNJM''+*,76(
PM%6G- U;;0%E3W#1,O)'./CF1R+A@VSL?3#>67+@ #K*7#:*W-KS SL"(:WOVNWI
P&U!$!L#C& S[W2H$C*E@X\@M;DN*:RY:XU[X$K38%W3B89>G!^?^4':QJ<O@N)!1
P,MB+Y85,DJ"?[NXCY9&35:QZL!4315>DCW?TB-"046MY*(82?-/A5-+ LO,#SDYQ
P T0[E2I!Z+GL-TWPR%9T;&(+4]PN!IOR\\^\2AZ4,\SGTVW3FT V8DQ67H;I:[:6
PY$@J]APY' 5(_E%7#D.%OZHP%I(//E88J6UX5,N>JM<'-U*?7[<*YF_@Y);CR")<
PKT5.YD7V2T=ABS-F"8!CJ!'(E!PQYHC8;8KJ*?+%#%*41*LFEG,Y5>P8>I._?JQ&
P_#ZQO2H0""Q=FAGIN"#LKT)8"/4O<7%Y972YAEJ">PH6U7UN1BE\H>\MVM[&/B4F
P49DYK"P&U&?LD_?5SA0;ASYP>2%BPFPYH8[(BN^9#N74@S;KF/526&;^]YJ6+@4X
P,XR4I5+B_M_[BVD;:>?@?X_.8&,RE49YHK'HR+*'? M+7@VJT.[\O6_IB'2U&\4R
PP-\/V0BJCNJIVVG.MO%\,#K<7-UG$OB<FH=M,SUVJ1?$U=-GBPWJ;Y1L,K[81O@3
PG.4UC>SID3LE@H=\-G">_XP;?G3!*H,$=%%?Z@+AY]*IT/S)UT3?ZI\XVYD1(&1&
P.,RZYLU!#3F 2^2]5""6V##%=\J/5E5].=8&9$(QVI@<IL3"'OF&55043TWQ"FB7
P&FRYBL;W38#)<'Z<<^U6(IF#["YBZLBH4RPI!Q[JGYN2A],^/9Q.E^!2-[^\^+20
P@RPT;RJ5^@$]ITA400!^,NW"KC_4\!F5([0'=.V>!I&2.B5)ZH^QGU18<8=89Z*<
P./GCO-C>8(:6@VK)XVE&D_CDO;)_0N8>?K,1<.E,TC:K(]W]57M +B4N),#A,E-J
PCY,0$]- L24I'^Z_<-/A94U]>OZX6_C[4>AVQKS2V(A!\/.*(43/57GM6%CVT]!F
P(WUM@)@08U9MH;3%V,<G>>@8<>BIUS#+M9J.A3JL+^9"974LPDEB&WJ7%49NA.D2
PV.^2Y>6*3#T2K>Y40D77,I?^2V.96.JX4-6_2Z@%JA"@%4,=0#X5=NMP;R&*Z2F.
P:<K!E")W[27\Z MBXG^6]'QP_$KR?(,!3&'&TX,%[@<@94:2+3./JUZ%_:I.SOSF
P2U *0.5.V#JPKO$/K8T^%KEM[Q'0(2_12&_)+=E;MU";Z%;*'GXPK]'/@0IRU">Z
P:3?INEN@+B;DD-I@QR3),3OLL$+@G\CI/=67@37D9'_Y5A2=H;F/O]5T4L/,3S[V
PG@IRK5[LP,K*<II>,D+2^CTE]SYT8T5%Q=\;<&-*/3E+S,'S"QDZV9DJ>,0):I6$
P K(?V- 5:2,,?Z*/5)U(O@G,TO*&:!_4;#.X[+(!QJ7DWI 1%?X+\)64A(2%'KE!
P[S,,01$S"-1SHX&YLA__[FK(:#CB0Y<V4:V!">%_I!\/6BA[WF?YT3D=DN@VO?*B
P!M/E_[0)([(.O!;\"@SP"1XK@ZJZ%9/QWK60B5L,JAQZV--#.-E$,R=2E%URL(ZJ
P_ZA+@D\NI-)AKRM8(]6O9VJ,/$\F/B63!%6Z"V#;=.M]D7JJF(H10MS"L@4OU@O 
PL?R%(T94'KD$M&^)V$RD$ \.5YG3A#1I:P5('D7ZSG_ ]VY1T+;5E!2(=RM64XWV
P3#2<"A_R9$TZ#L=SJS@$O3I77;.?&CUQ06PJH7QT:UM"7@^D]"=DMU&(BI5(C0'_
P"8HAB%\U%M\X20+A_-N'" M%KQ$007E,*)UEP1<"[B#?^RT:.(1M4)W>'OAZ^%/%
PW5['F^@+J9/AVT]("(P8)S@AFIK//DE"D<W\/4_+D,=)6I2+)39[Y<##G U0A7TA
PQ/)X7( DD4;Q)_XFGO&C[9]-[-;,A5-6C37,.#=B1,O(.S^:0:M'-.V/[VHVTG^%
PX-[U3]_T8(89[_\NJ+:@_$X>NZCPW8?P]_\L^I?0&&!J66OZ<0DHT77:-<RUDCR!
P,>YJ6;>B%A:'$U,EM^WG/:[7)MER4_@A$6L)(JB2 90*R45TSL(;ME<M"?)R8?Y>
P@6\D*<'^CM^V^E9\W)BHILJTW]2B>@L)MK)]PH75MU<9'<"W,&3\'&=O](^,:7)5
P8"@=D_L._NV\J%*86)3[1."! =YZ%;]1*8G\,5AF\'1<K4-9^K;IX%UM:6@-TM:L
P6YU6^LB4QKBG[WQVI^9AD]#K/]?4EJ%51QR4)<+^O)ZOVYGOAG:<0<FE/S_("3GR
PVW/GXK3R0.+@A9Q:**YC_0OSF8("0/@NF\KO$6O17\NF=-)LNJ4A'UYX$(EN$>_=
PL\#@@+JO1O]25^H&_E?'DJ;Y><DF+^^, %)O3IC_PS_*)C!RI7,*:JPP#DDT9$_J
PL<F/&DR%$DZ)N&8?[I!*'>1%<&=SA2.R58\S=0R4F68T2KU"YM$UH[^V6%G0=7G7
PZ*F^FWX:+V1]$/O4*0S->]I=],4)65\N@@YP38"J*@42?*W3._<@1@0!CVU4'/U5
PR+?10O%/XR1X*TBV=P32&XZ5EG/SDZVK0L@>5N\">H@AU98=YO(1:'R3B)]W4N!Q
PU\&C<[_LMZ*BTUU8ST\NHP*\L,?BUL9[?7#*^]>%R43-8EO?N_9Y*Q4#N0?CBY0%
P%E?/[M;1+ VH. 2I[A-L.'/%.7>Z^RXX*PWSKXUDS^@PZ,U(+!E#R)?Z\:GL_K+A
PTB6B,BCG=8,S1Y3QGU"C?Y9 D.=<4'D8_$=A*LB"3_8]'(S!+H"/P7*O@5M$,["U
P=,ZP\$:=_<8,+1@]*TI_GD!DG'B7X:R ]I/ ED\8$,4@>E)+NG"]/"%[9\Z^JE^Z
PK/<LKY41C;M5G,9A+=>'!L;MSO0R&_-N;5+&MD]:3=UY25DA5^U^I4S<<=EHJHG=
P.4'NAIW$AM?!3I/ ^CN',[55EH10"Q/J]V$7=-L/'2#,82  B<QYO;I#_H/PQ.V$
PYK\8!^;-_P2VET_!6><2I)V6P>'H(TBJ  O^!Q\1%E[(H(?MVO^;][OXT]9(5?'X
PDGC_Y0.T?RMB;X"QQOORKK@L7C;SE0"$7C_,HVN(?N*.%:IL.XPP;88@+U+=',#X
P]*G._2I/,W!^,4MR]7 K*C;.'I#B$@D)XD2-1C\+[I7(+EY:]=>?#?W[ZTKUMC/T
P%[WE@.5<5E&DQO8@E1&M0V;6<+C.I)4P-N%/3\K7+KM%/OZ8W"/\8!:SQLQ!R&C^
P?'<,%H>W$@QL[R9U ,JP3&4+A&VW9(.5 %NY>HHWA?.NP+0BCP\\SNX+I-O@I@I=
PVD:)E 6MAVIHDL:<EY5)^]9-DU9/&M></)&MA:D:8!"*?E5)S/D$&&YV@QL'$"#3
PN0-=@ ),_SQ1B<5VMB%]O53$7:(9Z-9MU/.-#(YF9US%/(LD X9YQ^I[170^)8GT
PZF?5%*J5DYE)S\&&PM-[/)UO9G O_?/UPXD$MAOU(9H<1:]HB3=<9KZ$%YO(/Q!%
P_51I 9M(ROP!NOD _WX$8\Y]>$0$C$*570&'GYR\'Q^2[UA*T'1)P9CSQG*)@5(B
P$KIVNG[S-;%>C+&5MDC]7 D<(\X\<LECKMNP " C_4HV!%82PT@GHZLY%A5)X^J7
P-.N1*;;+JYY$J)\P>XF,QM4>6+4ES_R%=O8)8O$3B*KLI.]IHXN:(MYP <RX+_HZ
PO9ERW'0*]^"\T\P:W>1_>"H&?6E$S;@AVGLL;MB=UA]5<@PT#OB2](809%ICK%O'
P*#OY&D5=UV1P\"K$@C0O+AK"H#>RM+(.)!HM4KK^V+F'ES+K,4!V$H+8;+2<,>TQ
PU&@1&-])NS?C)YME<!?[2*?QL ,V[M.X]1VA6Y,-#>D)+24H^*I*E@7%\;?"(8JM
P].N94\+^D2.C<M73-3>K2PGETFJE$3$LD$O$H2L!N$E8OH+D ,!YPGRS30O=XG,0
P$8?O:3#GJ28%6-PF>=?DJEV48$Z:'[V $@)7 &%(P47@X?-9/D@@-'GO.-\8':(.
P/LXX*+>\ZC0@8VE^D"YY;CWSYN1@OXETO.CCY]]&D?^>Z=T\B><"J(2"+"P4%<!N
P[Y(3*$]IUMW7,.G)(HFS#J1 -E9D\_97VVNUJQKV1M$%^QK&R[Z-9$?;TN(U9\ST
P<QMJNC.$;#;#M9J]%)YK2PP0(&. 4#[>#O13 C4M,XHAY(TU+N9<%YM?5IA1)18@
P"_RM$!1>]\R*5#&R#_UY>P02S80ONJ6,\?$RX:>7"H4BN?%2)%PQR8Y&X# 1ACZ 
PAX&*RQ,;PD0&HW\[R_"07;)1<G'X)]X,N9<#*GF[S;]D*7:6V.GH6CXES=/3?"["
PNNKRELZGC$ R>1>E_'!O:/F!A>^W&RVLR![Q?.7 J7:FT@\JG^6I4LA6^?^]H=_Y
P_@RUTHHZH933R\N\:2*TPZW/7FACX0:DA0[-$EM.#D'!#S,PQ)Y@9O7,2>CS1#>S
P\J'GF:W3!17^].;3&%LN_7+N9GX_#D7,WN5V?@WWNVVM3 V1F$4=P25-T8I"'@BG
P(JKW#%D#A#4Q27Y %S&.QYHMB3AS#;>3;7M3CF/  <MN<)RU&CM9&K$00H"]914B
PE6>R)W2Y*X=0A8AOP+)&D3J=TUY6%^<Y:)&%PDYNE4O9T),2_PS9,8(&/M\G&F)+
PS&C'H EN7EJ_V2/D6!85K 1TO8)DO*F&](D<W0Q&5+EJ@CMYSF6XXM/4.'\$\C5S
POP.LQ!*TPRG:J$R8%5;54T2H@,?+_(O,NJUU;WZM#_7?+D%1[+R!BC^=,Q5/1\49
PB*TKTO"U,8@6G'3[/N4MOGC5YWT+O)Q/0']Z\XBEC0I&@]UP7"::L$'?:B/:FE4G
P4+P+F;AC3*:X!5WOAM:^(!#]K^_";88XA)1\Z>KI9I(HJ";RGK-\84Q,*%F\,?$T
P^/PJ8B"'=.6SA7@.ZGEE;H#<,M0<(!6[_::KK>'(1A!:A4[B_+JWG_AE6V%Z8<M)
P#2,),Z&."BV'O P*ZK*Y<?I)7C <B;Y3M-/0N+QJ\)!>]E:BQOK'"3!3O7%,,1LG
PT?%QS<B^&9.%NE$X<I_8'P\IAJE(#JU-NJL\+ ),#*P+#EN#ILP&"'^XE%-QIATP
P,\D_)"'Q&1X*E?^UC!F^?K+A>.Y("#O5$TZ: 19MWBFE:ZY#;44:\)/(M678/Z!L
PI,*_L#8;LM3ZKU3P)O15JWL1UXPCDU2Y3HKL<KA?QG!VSIW,6?G%@IHF/3]X*L3K
PN3T5UBM66$+&EB1"D.X +.P-B.DP(3KLRDJQ$)2FE;N?TX;\W<\GRK+Q@R._(#\]
PU(_FW/EY3/!<BT0T\+06<_DNQ0#-NEY_-7?&^WL)K)()NC(4JP[)3&0@!&N[0OJ/
P80$>@N,\W_'2!4LGV@D=Y$+8!)1Z"SU0JX)<BR/$PQLJOGJ,"ZPGM,+[=W92&N*K
PW/Q'');7%'!,PKUT.?4U9=\-L6L%UFFOB#P#1\929N2 *?8K?U)N+O(J0OW*V# @
P .9%87".(2[W+,F1<)$]=)M7<=UC__;%A& Y/AU\9W'Y(9)53Y*=\,K3;0D>Y0P_
P$COI3O[+7RBK"7_5373G_L"!$B4!B-S!HK2#<_,FP<W\["R!U7 !0GY=^GGTOTM%
PH)1N^NFV)C#^GL-PM.'$V9]CMQ'\LIC_.!Q^'O*\OY,4F]?17QN@ZJB505=S>L(%
PXN/N$I@K@(4<Z0VNCRR-Z^]CV4[@-6PB&+F7 <]B\FK",1C-!&Z'.=&8*,> A.E^
P#.3'2MAYK4$1^+XO=H#PT=Z<_9P]2TL\ :G^PH6A+U%;AUC>H2/UGR=:.X3;H35 
PCA3Z)S7MA3\*A?(I?MXKB00&$8*&U#/\[C"WLA1V H=Y*XYRKLC5R.5^G&#VO\[E
P*>0?J?3BUS*8#4E_J.E]J+O7>M_,D'66<8%95"#>QA5QUI4PK&\;)H4S- VG@[F;
P0:F)FU(7%ZI\#0:&W" ,T<W.5*GI7D]A:,<A7V*#BP]'N&#;9=[+\W-&QY<-:(L"
PU&Q=10TR>R!.C?^MTPF<^C?/Z*["EF@?L4;.'BP"DW=T=*9K7,.]1USN9)M]T]V^
P4!VMTC L05)!MOGG(3-]=S.(9&4.C%W90B1U-[(_*^;T]XA/%.(C7Q> 0 =M#8L[
P='R-YF;UX:%[_SF!,*W*PFC_GL K#6F5.H=JZ7C#D9YZ]J6JAO[#\UTZB @[?U[=
P4L[!0:#S(%H6RTX+D64YDICK.\I'IMWZNU\' -DAX-3.YTKW EMWP Z$,>)[&P:(
P\CCVX%$Y\B';;A^[O1EOS3(_6;G9.Z?,$5*3D[RN4XWK[ )0Q.7A)?H"NI9(W[2S
P:>OE%:(8AL4=+$@+ HVR, V6Z:.W&_I%8B+'!>@U R#X0=J3R5J*JY)R^.$Q'?X<
PY,F^7=]4^1<EB64.>%#8J+&TI_D]3- JZ^%X2A>4IE*F<UJ(!@P N#XTU3@Z/R?H
P0"K@<6@ _'*$1XC?'4!$U:C42BOM/S@-7ES0E;/FA 5DQ>7<GK2N,0!#WO P\WV$
PYI,":E>T5)OJ.>:3\;.O"Z;*BL*>]-R^N4"##H(](]Q#\S YQZ._"$Z0@":*<GHF
PX[YE:BH72\?(VT_-;_.1?-D%'45+$B)KHP"T2<TXHZS. /JZMG&]D\JAFU6;[X2Q
PXB<=-+OTZH&*_;NKJ.91N&+UDET.%K[$G8)/4UXA<6\+\E72SK"42T9ZKB\JM'ZL
P(\(M35FL<UN_+?Q<-#^SZ!C E,HELVEV>WLOENK41."ZS4*I$SY5&ZB_%#OQL?U6
PI&:VTAB4BWC95IFXLE]JZ$RCQ@6<R>4\<.-GP653!&"T:-YLF]Y=CW'*<\KL;3J]
P%Z@Q\H'[0-0Q;HXQT+]6MX05A(+*5+4PV8).(LHE#A(#YSA\1;?^8 A/7-39GR/;
PVKNE2_L7WD!.:,!:&^>W/<>?X;X@^K&VM-$U5(M'2S1H'[^!6=*R+V\Z<^3XG599
PFW6$:)2A39J!_>AE8QA@3X+S:X*VT0VZSO,JPD6JF!/GH2\,JQ_+H;[U75\(U 5-
P.5.G@J7V2WB(V)U'QY7\*#*"17S Y$DZZOK*9[.%<+.=8<T:1W9YV@9)S.(_*4D@
P/F,6Z V.3"Y1'M6B:)"2/CJVIL,AZCV'1<X=.^^M91D \P"UVQE?^.WBG Z:<Z/G
P,"CY'I4\G:.$I==:L"\8\D#&4=C;XPEMN@N$/AG'#+?!];5DA)U\4=38DP.>;"#7
P!H@;'AJ%J?(>CCS4*QDH'HU\0W(2U0$ W8^G%L]DPIJ;C$F^C<Z<2 (W0H3\;T;D
PLSS^\F(E$MF(K[8Z6DZS^&QNVQ,$*/BSN-K)-F8/VF+=$$&02+7>6=%GQ44#P/!E
PML_-"GM<X:#&AWS>HL43JT..#(N'UWBM=C2.TU5]*A8C8V8M>;1A\)[NW'O19R)^
P#ZM]32L^W1T;%Y14;!KTFU'>J=O"*/!JQF\)E601?5<IN,Q.>]J9.)O)8+0-JJLG
P() ^EF)\0C2R\ESQEN%'H[*#HY;TZ8;77;I_QPI:'C /6)U) PE,Z,95E\[1;$V_
PY '( [[Q4E,.Y=2KX[^<1!(CYU8/H;R'R5NYM-[:&-H3MS5 =I*@<7F1'UI)%+'%
PKW\GRMIIV/]:LK*G8WD7O#30#),V8;-0/L#V!"XS@N6IU"Z*7ICM,9O7S%V[\@;.
P+'EK1CJ+HOZQDB01D[Y-69S7F69[TGP* 0=__LXGGX&WL9'0M'9J:LD9\_Q?LWWV
P"S[1_.6H)^N(%YG(DTO[.P$DJ$OB2$!$5.?-9]11QW<//TG;$49&*C&'QA+'-DYZ
PDY+O\:/MSAU]F#0+JS@-196A9 W/7YCE&:M"W03HBN)<0S /#?VGB[$V)=[H4R"X
P*CW+!C4EN/Z[C#Z=,BB[8XLGN<YL;8AD_<_V!MMK7^?/UU.*.ZC;D$)A86-^T8)7
PK#MVR*$O X1[&@,2Y>G2M&<NT.8Y2,/ /ZDJWWYSMYFP?:RZZ%3Y%+$= +TTHB0.
PD$[\..,ICZ#WE,!DOA=4G[*0YJ+!$.>\-E6HE_-IZ;/-OEVX=WU=T41)?Y:=&L>'
P>V8!)W/1W)F(X&5]=Y6L5?,_4FDKBNR/^D4X!_J1NN&7)YF/6R!L$V-%6U3#R-Q>
P+AT0/,?_7BD8MEXDB*L1;2DX!:/J [G")]$JQ-;5O/6%B34(!'#T['6-'/E:P*E[
P;:XV'F0T@<</_.0GKG3F0XR*6<'<(A'2Y#KJS4A>N5)1%:IIP;<4?N X,&&W>+(N
PTU>@I?S&X"=6XKJ/AXIIT3JP@M';)ZD-3!%"/XM6\IFJ45@#5CRVKF?G#"1L&B=F
PA@ZYJ3@J&947& 8$E]]P%QT8"U\/%%'K<%>U;C.%W__)(N4H@JFT<Z*A'DI;AKO@
P'Y;_47 EMFD\_+Z')RPM,M#M(YZ\(I00+ZPF#D4&Z@HS> X6BZ_I^Y%![Y^& GOE
P4D'+.X-O@R>1V?>X?N8R/BE&G8$O!@$^@(.#?2XXXI3\CKZ]R/#]3D;8AQQ9AQ;]
PA'%'_\&]*.)XZ4'0954ACS#B=Y8SR+.-11Q?MB,LSL#"'--IF:@&*<BMOM/@._M6
PD261'I4(E9'&A*6PD\/B;@,8KPA6QGI5J-;5+=D$G NL.U!N B1!+##ST,T&R/]"
P3G5=84H#R!6R-M9R\:FT-5&6(^W+X:&S9$H5FD+I,><OMI+--E#LUBW6> F8?%4 
P%D?PUV_XA/;L=RJ&2S2E^;VC3GYX)@6%Q=\,SI]=DM;9OTX162==,[(_*R*6#0K5
P-DMN.9];9MUG%PMPY\O)>OB R3$!0@\RAT\I,8"*;8KY$ @3S+-/>Q!O$4?9D86M
P]/PI),W,EF!IWE/6)P:DH^:K*2VL\?$68U-2FD>@AMTAW@D)KOU.8"6@-9RX98ZW
P#?Z)UB;C2'*G:&MQ51\?V#Y<@BWF_UOL"UN TDFK$7ZT22!Z4@T@'YJ)JZ+? <[N
P:">,=EB;MPEJPXC-T%I1E>?;8[\2ZE;2NHHII \\-G$%YCON[EV1!5^,]65]6R28
P*,H@B.0H.$XOU:\5.S*:0B)]^8Y/2^Z_T>,4)](/VSFKL &B2B[^T@M('363PW<0
PP\IHEFDZ*J N0:#*S/ZF^XZ )61@7HU7B4"U\$!F<.KX$[_%UFI7Y81::IF5*KK(
P,XOZ)E=[@5.>1[7-M[\ Q4;W,A:>+F(7:F@W7%'BPQ6"F$RGWK^)E?P.^T.^%"NO
PQA4DZ_2R*.P+<-T>;$?LL;O@>U[(HD,%%-BB*P89X[Y_V^.T'5+%F--?'N<,B&_!
PK/[*D(!MNC<R7?0!O@<E3,5KY93 _6'D8YTIK0H/V;+S4>&,XAU*C93Q?J#KMQ-6
PGHA>210^)HA[:?5Z=H84\_ K[[LA[N/^V;&X,UKH%[@K OIBQ75\FHVP]#7(A(*W
PPYL14*$XYB(\TG2!Q)5<6I9Y;69$Z,68H,5:@^D>2Q47ECZMEA$UR?QN/\/%/R\8
PF=B?UY<&Z%IL(%3.K+];C9PIRA;]1_0<B/%\^BXU<C[ZS9&'IH/:620O_RB+H.%5
P:0H]@IG@.5(W\_C&^2L=HE\$@.2E5=!-RP!6RE?/.ZDL'GQ5]MK<5 I5^G@1=>98
PJGDH%<J69I$@RG;U7+.H0!\=T6]R+#2<1F!SK##7#-/P-.:T-J@>CPS>RP;<[=K,
PVX3GG1::,B_"3_/9T69I!0!O0O"4VS9F\ YM2!^3M;+H1QG&6>D<;VD2T/&GM^(8
P[?NPN_:I;1$3:75I0,55G%W>V+.98J"<](:)I?O7S<CBYY#^W&I")USZFJH@%+(6
P[ST.,1, >K[;RWJ1N-^U0Q1FZA3 <X?.FF!O83'"$[^P"^0H2X!'>-=112USKQR,
P.'!KVOG@1U(#4OP7ER?^^R?H=_>C2$_EN6]!.!_,S)T3Z2_T-(Y,*?S[;=/08C 1
P3N%H !3S_I"<?@&Y! .)''FO;HNUX5H5*H&C6Y[U6YWV&1NI[&'&KUBFS:]7!5QA
P.ZI1RXIOI+[V!"U5.N?+?<:%Q&5]DOK U:-G-)I=#3 (C"*@"1!AE#:\"(FP0?'G
PK30Y']SK (N%V_QAP5(#SX8'_QTSL"> WE3GXCV.8S9@7-$09A19_0GC,ZKV?*!Y
PD)8))FR\%DT7@[KWL[/D)CKASS(^,#AX>K'M$8#!O>O=?P2M+L7>"R(J>1VK[Y?M
PQ$*[=70+E0\\9S)-!EPC1*9,J_A\FC LZ#L2' U:!1P&M>MM\5QIX8?.),E6YQ%W
PNG?;_9VNU]'WMWB5[A*@"<N*J/CL#9J;M2@]P_L, URTYE:,,EH!#M+NQ.,G@[.B
PN@4MP$ME(RZQ:L>MS*" :+!99FS>OKFE(?(3MTT"@K.J=W34D?TV@8%S4L=#PRYI
PUUWZWMN96BPU7-VVI_3\-CMT_8O_%= Y '-6V'+'&=M.4RJIIA";\%".MARL")I8
P[%-TQTP+0U)\VCWBD.(3/F+2)1)3C"<P*;#X&N;Z1H8PF<U#GM?,I_W!&.(UHCC(
PF3L58+)6HQ#6)"1RL?NQS^%%1%X;BRI$!ERIP];[E_WW'E5VF-FQWM-T]6C:\/52
P9I[W/J?5V"*QV[5#M8UP'HE@#);J,/%I/ =[*I"3K>,A>K=%Z_/;'PNX'74P:KE4
PN3KX@Q- 5:>Q/L(E?CUD]I<;^S3@^HK+H]-?F6;TBRZB@%S,/FA+L3[2BD:CGCOJ
PX+;=1 @ZUGT[[=.:[#-<!7 \$A.D;//?S3WF^Y)75'P(K78>DGAN/CQ-,8>4&!6G
P\T]W901=+AG=_'")QH9/IWQ!QK)]HBASN7DA%'2@C7A"B/0[9\E@*SYPY%PEX5@I
P/GNO^ RSNI FW_13DH M43:UZ.=''WYR]KD?4?>ITSKA*,TYGT*_$='0X2B"53;M
P\5WE@L!H"[PV2)_3L #'X<_77(!*)MP"_OTCIG?LGCR;3%BUYQ/EW+R(64F(J[XP
PK\4=%[#[** ID@D@ADF^Z3>R*PV =4?U8KD, %I@SDLI@A*4GT!]]\J^<:CX97J5
PCGS( 32*2#/=WZGTE06H-"B]?_.<$-U\P\Y]X9&AW,6EK8!=HA#5^,\5K&&LKNK0
PJB[O:<<$9+ EXDLI7=)YO\P)FX,V@H>\,ICVF)XE4GL0YH;U_X5CQ.T5,4Z/7L4%
PY<I3(R)/<7"J:$7!)>9L8P\+\ZM[!3%J Y*(F0./<FC9VU]18Y;$IT7=7.ZI1+M9
P2XYB*%WPW!3)*KD,#(S"QQG?P/>C$Y*BBPCKT=[S#O6T9N>?@%5N#%/X@KZ <UXQ
P ZPH%@-H[W27OYX#8W$\^R"DA\T9"X[!S;"NW(KDN,JORHQSE9!T)R_(0X)82H%'
P$:W$=;I!)3MBK;K6-J?95?^E2$'<MC8F0>%.*U1Q"Q$BL38K!R9!'Z,'0I!Z!>Z'
P\/B$IO?R<BP8E:RK!Y.=Y:"[<-\\9X262>V&2X3ES:;>DCU;Q[?4FX7Y^(M<XQ;]
PP47E:A-8K#L3PT\FL9DDC966NC.>&C9U&B(">'H'7[4K9HY>X\]BG PRRX.LL+.Q
P9)(6! XBAR96>"BV?V<PAMN6NE8$4_XNSL/:Z+4I?%CU,_W*#7GRVVLH08A;H#5;
PG;JD7]/GEU4UFB6-T'0'G!TQ;7@#;_4^LQ<^0'-G:#'LF<>9BIEBX6!'>'2N7HU!
PU)E@!)U [;H,(S&$P/C*[>-@TW2WMN8SE%CKR_(9<#YK&$PFNYYMU'_S3&BE:O1B
PJ)PW2LHIV,=;\P9T3B6_@"\;89W788JE:XDRA\7NH4G1X*0D=6&BFHC:#K< SO&P
P+3H\LL]D,F<%N TU,"-<Y")PD<[^]9H>"'I#SD+MY82'6]UKN_!>4P-<-P.8:$>=
P?%^1P#Y^@=7_ D=8BC>@& &U"Z 43>-+XEGW"F%FXE?C3(#XB0_K#0J0<S)=</7[
P?1)J(!>,-8P5F@9UCM[D#+^W=Z:ABXP&]MMQ*H2CMQ)13XBEF9Z'+;%+,E-[%15[
PV:-:<\/#4G%!>[M'XT79'WW>L7- #O9K90UE#&#5MI;/5L,G2X'W]H</:*_C4=4R
P;SK9"5J0KY&Q!5+FAH[$>"$\0R[V(CKCF[>;DE>$P6I4JA.Y9-]@-G1J5:<G[TNX
P92=:*+C'.LU<%M/,$^3+)\B:$$&@S7=M$]9ST):)[_"XQP6P;ZYQ7:X@W"0##Y,)
P>;')8A=;PUX".%#6:+!);HB!23#JN]4C*6I2I-LO_5JT8=AMQPOWS7L[KP)EL"GP
P)I6+JQR7 .T<5;# P4N]T:#H602UV5WJ+<6WXYHI_=VFIC:L5*ZXY%Z80N88Q$I&
PZB<6E]8]A9#Q''<\!T ==\U.!C]_W*OHAN$%( ODWN(Y$1*X!O^42. 9_2^T\4*-
P7#!\ 3%++#F3: ,Y83'8(@0)['NE/2I.2#AW8-(8<3%<WE3'SP'0E5OP/5JM8?1R
PD84N=U.I5'U@ XA2RL%!^5:->Q->P"(I?#1K F]6:$UG9;N5&/AR[ (,YH 6)<^V
P+54;0$.B<@N"4.>DS$I=H1?M4 Y*>&/Z?YP\"S86GN^\V]G-C$XD]+[_<1RA1&,D
P]5J&48F\7Q"J< F!PR9PWRA,@F+:63J*P<1HX%F>S;;NF0VO&@]I1(ZB0N ">X?T
P0])7#(3LE5.TVM:[Z$A?D LQ,;(-)H5@S=O%?Y8_DZU#88_GZ@UHNJ%'T,P$ME?,
P,=R:WA,==3$%O;SXUQ4=93]LFPBD/F= [NN<!&2<E7=07?R^H$$1"-DX",]<$SFW
PJGK.HN2.(G\E1*H&HO'4FH.T8.R*=$V%;V?&,TZGH-SBJ08*A7^-YU#<!KUT]G^2
P&$<SYM[HU%$S@02[ST,$H@MYXZ1+ZFE8[8-DO_P@X ?57YY/%[M *[OT8DK1NU8D
PE*#1,P@:S$AH>"R/&>AWMEYI>99%P#U((T-&,XW9-^K.GU /)ZJWR0YP:'4G1F_<
P3&-,/MP-UE1O5^IDN9(>PUM&]ZI:5D(RW[A&9FFVULL'3XR[3,J*\3#_)GWKK,!O
PVJVZ2S%!D  ;]+S=;4WT>88HBES65;("$&H58,F-0-R<_G9R<Z"_B1S;5VB?,1^[
P=0&YX@RTL:S/<KE-/I;5Q%.;'V3/BG.'1-H7MBX$H!$D="#$_)[/><?J!T;C$C5N
PA&>(/;Y#^ P@K9^193Q,$)X:XN25^=1B)=@H4E?:C#7N0'_MB0\@<*YBY:&MZ/@<
PP$@S-MGD6)ST5T"%:C&_5#%!64E";U6R:4#D<-7]*-5'(A6^!$U!NU7>TM#*5K=-
P#<CIJ1"N>0##?L+HG(J1/=X*F153S6,RB:GAU4>_9>B]\&*<4!J#T"#P'M$'<5@4
P2[;HJ4P5\URZJC<.>#]OT^[W!F]JK_IC5UMXIM5<,0P+I64S7=XDJ@96:L1A,8\)
PB:8QTL)>13.S2J>',U<TS&<2=C\,?\0G&XXBJVG1L='H*1(DI3AX-14+9IB/TM2:
P4C6^/7.;I1X%FM%(JTL?BI,J?XF6:D*MM<RI["9.CV.1T,2]9!DGO*NVA*6Q7,W.
PZ#[P1N)9:QE0A.\I  RDV@2(;/V;U4+\$K:AS$0IE=K+]:^N9X./^M>Y2M>O+P3H
PB5B]I4E/"<(78P4^*D@R]W8X."2*B$VV'J24QR_+&)T4@9E]4'5.K%?*S.IX-Y5Y
PIZ,(:G9F'&VS*5NF9CG=.<G5#R_5: HJ2*N:.,D,#Y9$4?2!TQ7^772[*>Z@8B:@
PJQJEQR3"/P8*NG(@1P4'1MJZ?M3'\Y:O(X-78](YLQ#68TL$F\N!<?L-HB03)^";
P$PG(V#ZU?BA!L/PJVI]+CK^#IGM\BPFMS$[CX#SZ 6ZE-1\G*"5X*:87PP5N=<[R
PRB&8;TH .8?*"2?>P=%?N Y+KRZ">EL@SG#B'*+YK63G2G8=UXOM (;:CT4(O,[/
P?F/0WV'85;C>UIX<GV[\A](#?KJ=(57J:<&P\+D1]6<0:NGM[7S)Z9I7VEL&Z"(A
PU$*.".GCHW*NS]B"M;MO-S67I%">E01FCS&R[2<^S ["OVAF=)0B4>9B&[D8_66:
PHV!M;_:CM1.-+-*P_MF8!8S/&28I0UBF<T5>1"6[7.9C=;M=^(XFEU#TE65<BRME
PT"_)@GY'WL6;>!=X[7QN>_*F)BM%E8FVU6**25*K2 >-('.WT7IIFM##NJY#RSI[
P45CYD14"HNMFS+DRY"3* Q=Z^L#OZ@VJ*XX+3M*H;8U&>G;:2H*%9+BB%@8,/GJ#
POL-=J>LZ1HYEUO$I?2"%_:6J&H>XR*YLU/6V7^*WI]Z8463\1'5UTUNVS3<'&_-+
P'RNO^"S8RZTHZ8T$WG/"7R+VHU7\%\R* EFHECC/^A>.9# /0-8:=YY93N4-VU-J
P,[(\1G4/"XX _M%HK[W_48$%R_N@R%VH;UR%7=2*-$CM@E0S>)H:I"QF<R9@K(SN
PWL4."W'[P'/9/? D.,E/B+OG3./DU;PN0#\ZAZ4;+8B]QST]7^HI00HRTU.ZYX;]
PCBIF=BSHYFQ0%O'6/'9;U[#^(1#V@:*A&1:#@QVQ;L],DKH0\/Z5CI&/BED;^IR2
PL7U%QA@,=&?K]BU?DOJ=AL#' 2T>V0M/%0:$2"&DJ=G7LMMZEX4(LEK]WXUC(D_3
PG%3UL,=O@4@KV<,9!^G&W"ZDSS&BB[ <896X^+=V3J1/#>WQ@1R"I$&@0?)VFWK8
PI%59/BK3<[.2+ O^&AC4WX6US;H/@7'^=Q\(H\0[MT\ZB<CXI6G%M(7I'3Y:Z3X9
POJL7]LB19PRB(M[E2<-!DW?3MK#SKHS5_&9+I:<UDS"@3]"G=-H5(F2Q(6O*;ZE(
PW&QPWL)GG^/S?S0%J@*?\@4U#.@*MNX*-;T*K8N%#"54?,3>:68P2'":7@AW%?)Z
PAW%CW"+GUFFD< NEI5F>.+29O<93@)AC8,F/-/T9LHQ""(FB:W$Q;WT(P3(0465"
`endprotected128

////////////////////////////////////////////////////////////////////////////////////////////////////////////


`protected128
PDU7H_H3X>>IRR,/N?KT7T<0-(GPPGNX7S)K2O6232&=Z/G(,-RG>ZRZJA ?<O-9I
P)6V2^,?I30Z0UI;:@ -Z?*1!@'1Y^7&,6RJ-:V4\!H?[Q#:S3XF;L)<'.>',2@=%
PQ/"/!05,54/&&N9D43H#D!\K\J3.0M7L[PFY+NDGXEFQN@OGWRY<*&.AID./DN=#
PU1[ZS7*1BSJ>@IN\N+@=^["T>QV1(U,R)_ _.MZ)1ASS-KT35&Z#O-_Q870!F #^
PVQ WT!=)&TQ!D4!MCA[I*VT* 6]R&!S9US1#R935$3!>>:#]BQH7:_O9I#_!_)P<
P_0)U^B'96S.%TY9>"6*C5;=6T900S%VY_5ZT3]M4PCWLMCD\D[WY>X;P&C:.4Y9Q
PSXBKYKJDFJ#^#HC$;A).D?7O]Z^5HR,Q?-N4U]@SHV8]_6TJB^^N[6C2J"GG)BAK
PWB6/68HIRYEJ5@VR<S?.N?#"54]9F=DS+KO72Z+]Y$!_J=&B4T?#G"FD&2N[[0"#
P[1684<QE2C$*$%NI"[2V$WS^].<<'ZC5T),\1P3XL'O[][AO)S%:.<2@"YRGS!HR
PM5D^\LO-')KVBJ@?]!BA]!V+]#5?*;WILF][^N ]<JBO_-\O4"F;5%0EHB@F? )0
P3TQ]V;>\MOW>=[>IBL:F_QEWR=(EUOG#%B)-&L-JEK_ T7!)8_STK4=+R)J)#LPS
PABI%CK?"2.>6Q7A>_@\?D'5L/R#;0E%VED.OPXID?V[2JKM.U"6-;1CKV-)J;Z 0
P7," B5_?>0>KL68)W,>2(<"F]WBW^9"!V6Z^@/8R\8%+":LM$!9-CE'-K6=\=1W/
P31YLE-'Q7\1RNW/5"O\ ),4<10:=.ZZ_-3NK<(J-!3 N)A$)T^E80&F.U%%IKB-V
PO(4\)!;C[P8RSY2S")HD3G2< %W9"6U0>4N$>;7UW@UQQIN#T4+AMV?I"$9KGNCN
P _(=)]3\T;*Z1^7[I%M<)W4=AA+\OJL<M.]OQ_,&62-^WDUE4PJ[1/\2G$V-/R38
P-71UN +(><9*>J:''LF_:WB6<_EHL(@4D8],KTE<(4!(NHN_1%^$>Z(99_\Q#A1>
P9(0>JAX-N);WA5NN(I^[2N!\.J&\>HYQ"U_%-Y46[BJ8=#C14ZXK^LP-T7K+\KZX
P6K(*3X]U<V/C- /"U3*V@<S??XZL7M,3C&U1ATW Y6*1J>HU2U7 WMZ,;U/A[>X-
PH7Z^+-"[TTC+!,&/2"EF)A)P6KJE@<;AIRM9#H25A1]6J 8U%1)34TG23S#N,.8;
P!'>%!DL3(=A9&[B72\Y5;GY\N097YW6>F#?N?Z7C=-@_FLO/T*TPDR5XJ7.+X_A'
P06YK[&G: >?_'CU7;_6*693L%36A50&%#0]?R23CCQ2?3;>1E.>TPZ; A=FFG\%$
PY"B9C)J!.OKY;'.^H/STB7>:^--L,%4J<35;=M*C*EYQ<>88UOM4.6YU?D0))YJP
P/.LV[%5?I3NG,],QLA\FLGRE],4S<9T]_PS;K/4+T<-=-E0UW6GL<'._)57#M/BA
PU6(!YK3]E8MN:J"=P/M]#,#-"6?/*"[)O)<[(8V"?N79I#];_V".9_TJ#HUU9#O^
PN>7G(?Q:6;QMEA/6KR@:+Y/="@[Q)(*ZE$\GD+(RC&S7ZU[%&\)\T?.1 &);ZA&"
PF$U8CQ'?"A1_[8O-5BN6<DQ&(T3(*P7RWAR^4E:3\&*',7H7364PV#8VB\W6:GE.
P0P=^ .RVLY/+N@Y@'/4_P0B?.P) >*&^4[>(4>%(RW%UYMZ.*T0X?09&>7M<9SZ/
P/R+YUS^DL$QGVR+PSJ,%G9)O)E@$_-E]]O3A!_:$JKM8'_]SV,J!+MTC4SP8-? (
P',.I*[6XSHTOWABSE6S[M]G?VK3P3BC6BJ/KJ!0#SD PXR?EWES__80Q,U2ZQ?AI
PO=9O'ZU:M#&P\*AVX]DY5(!TKL:97@P@;CVN34#[[1DP[D.BQQ%SNOD[D6&KW"$+
P/LD*D_S_7MZ</6@WUUXK[JBFCAOW'UTS!TVS0<?AD-]'+)9 XL6,'/>=*+TTL-3Z
P,^).*P<4'=BP>R!H.:[J\L#+SLG.NK0*?QX3Y'5]2H07N%C)=$@6*U#?R)8<@[24
P7L(MP:A8E'D6CE=^T!P/X2&@K@PLDZUT(E,,+GFO3E%M :#U?MO<UV0R K-DL?ZW
PK@1O>BD8B):!G/8(3>Z *]PK4P%2&TPW9HOO4=40(%%(?=[VS&G58":1'W70\$9>
PQ*[UI.\U177*!!Z@"J* 5'H"J^W:J>%TJC[XS!4[T$:QM53 8J]9L,% H><,HTD&
P4/*'KE#:$*5<J!T'IZ^JO[X=W798@\F$V[O+;;$BHHF8)^\^(_0Q)ETDH\5SD>5X
PRP^;F<^U'?B<J\(2GP.,OMEBRAB\TMBF!6A+]6/>5U2T%IF;MHV*Q\VBQ=[Z%1-L
P'&[&E7IXX_+;,XKRUM:%+_96=UBP[@ /#$:Y%I9?D7E9ZH%Y(>?08W%X4_ ;E0,_
P=J\ E<1X"[M$44J*WYJQ\$NPQXDGA/2QY!-3T#0P3[UF,2^98[!F*?UM#C+_D[Y/
PQ%"\-^EF (6^- F#2AVGT)I.>W(IEWOBIF5';(KN('7R"5)/#,_)ZM,L="X*R41^
PT6%[1=H,$+Y-GH<TPV4%6RMUM&N@G,4ZR)Z)<]]QR!1.(1V EKMA?3I\MH()O$3O
PHNT_I;('OXLA7<CS3^EO9BFVL:Q&(=._)4 W]OF='AYX!_@J5K5)FLX$;I'B1)YP
P*3/Z!/_XNNA>@%=R/8&$IKLV%!W4I&RED:R4A@--[4=OBTQ%N\=@I)J0F^LW/(HA
P+-G=XR)_Y<M\V[1L_V<;:Z4)ZROB]#Y4NI9'A#76>).8B\6^VGK",Q_X9X%)OU6A
PM%)K_^^+Q\D%-YE]S-(-(>ZKJK^* *W)%1\^M"8P.[ [,E5<T;CR)F[:D1JOG6M8
P+<GQWD- >!UD"UKY9:I8.O''&R"_Q)<%)KR-SN&H$P\U5RM4^(V<CODN7)IVUXJ3
PC?-3'3.-U(QK:9"F'Q(E0I#E2Z906"&+%9=95EN75J7"24^Q$D0U#8Y@Z?,+G!@L
PI/\73AOH8CV\+MV$_-U<'#KLM[3W+:[)+*;7H1<N!>M!U1".:,,E&ZA4A 3N,572
PCJYEZ]2?1@9.B;/?$\Y\?YPFJ<E+Z:4:CR[<$JV(P69-/2&F4>=Q[WNR"AA*^Q,@
PB*H"^-^IA]8A- [.J0[9 PJ>7>4>2GC .Y%S4IC&?1)+)_DW<A&*]Z!F2L=69E.5
PG=1E8("FYYS?&7N,ZX/;OWNQ+V?DK$0<[]4I.!JC0F9&QWR>G$I.W/X7S*EAV#M]
PY3@!'8U +2$-\FDM1&EIK9;2,LSR)W#H[+'M$AZ9E+;,.1NR\<?9&RW;XMQK!*^2
P"=Y!@WY6W"R5Y%+3#(V(%?6XC]W>93.Z@KV3_PGSL:]+VXX=N0ATY)J4T0<DD'=6
P"LWU;#JL@X5T;(QS8FO;9SHNNI)K"@ICNZ-YY"Q 6O]B^)]^QDGA1Y;RTNB-ZM%2
P'WD;=<5:\2U6A40(W;X2R_B<%W,BA-1B89?9CL,J(.2MVD2W&D$3MDS6+!ZD>I9C
P% )7S5 I=,,*%D[+ )4E?6T(($1,V?%)2M$5-NX8*19]/=#ER\%D*Q?8?2_)I0K2
P?D9'%_H-V]Y.$I_U:U*:*4>7+J+?QVCQ,PM7C$\==$TOVG=,K8%C2_EN4Q0"02.>
P0;]3'8#0ZCLN?ROK#)EJH[,O15AITE # Q$-R3Z=Y8AIYN#9:W=/2T)QH0' W0^&
PON@7F+7-C,*QWZE@?^>>9J];Z>J/OD_T!WU0+=XY@2NAMS)CPWFL) DU/,C@/[6S
PS($E$U7E?+@0.^F*WN2,[Y;VL40Q878Y.O$HWM[B+&6,F4$1R^ =AY87V#\3,K4U
P* W386;9ZIJV+/NZ"+YQ> :SIF1#@: @?51YQ/X>&K6A","1;(QN; (.4P3XZZ\4
P'7.R)L;6!HG5 E'5QT(*L(I;[BT7@]TMLLSC$QM$X^IY$\D*+1 @M]I*U511I9JA
P4]!R,1%2]^<[2T"9'O! PI!A1&[O=2$,):VKB\Q*,B%&>O=@=<_Y=^)_B[H34B/<
PHVQ=-%UF06%-EVMY#E"QQ>^/0UME?-;=!4H:M47^ Z$RM-LC07T%R&%5V4E1R>A<
PMV?=UNM=H\W>TH']YZ-T7#QHR3LV"T* 8]U1VR* 6!M6T$C5X[/+:>;GZK-V)U;?
PI($MJ=HL7V>K9!0!U7"HG6J:914"<0<-?3 )B$H_EHUO5 _@R6UB2RY5X5;U%+,/
P.^<1)OG.]KDLLJQZOJBY]_]C?,WAH %:6 OW!#V[<GRL9=R(@W"4_8"O\7M+LDE,
P =UHPMENM8+)62B)4'R.A243LABKM$(-!OGLD+OG#C,PJ*D2?"T%+P2>L%\>>/P!
PN(1*B; G&'024'1.<GHH5%UD"9PT]S/!'-I1<.TCN!XSPD^*9=J_X]Y3O/U)7@&B
P4LAW&@AQ P1N"?J.T$CN$+2,RB7RM2$4O*G5Q?GM3$[*H<B:@A^"CI5\>5$"IDW^
P49R6L@KR\GQ2H(0/H L!+VHJC,+$0'"4"]0:3Y'#&;N8$=WBH]/[)ATKS,Z"60MD
P'4]@O:^^'<.XQ_E*30_G$H:>W. A2JQZ7LG@*:"X73Y_K"]I7_F!R"3I*F//#\&X
P3=\2V$'DMU1'R6*S2--\+-D=TL1RUA#E2))_U!0@C$Z^WL*>[3@<2:R($Q*H9W2H
PFT5$2*C!F:]Q3"Y#B^/W3RAR.T@[]K?KX:$/BNW#B_2UUV>URZ:P'2YQ(,%3Y$P@
PXQQ*IA'+1 V6SP!JE+HNQ*2V791&]&J'J>[@F4O@QN$MS1"T7,;>0\L;T+A]%"G#
P4:<J8]I93Q;LJUW&0_V(GA1 7O5LBN53X-!%1)==_Y%N/\^Z9(#F(D1RVF.O0^2)
PRUEV0]/AG$V]$L0=-PQO _VBCEW1B52M;6W^I.R&6R<M+CQY > D.*(,&5G0;[J&
P&?Z.A23PR:+9]<@XUZQW M1Z2)*+S\Q1J$.^<//T"UDW2N=XAD1S\E4K$Q(,6:X*
P?!M^+:'\[<UV?'3BC/XU/N8C]$</H?*7+^,R$@MV!&(FB[X@B)>RR"$G'K'QJGY!
P>.(,58S47CO)\:]Z8I^3+O,IN6.!4^^@DH9+IGA1R JJ<&ZP8OBF4:[7D+/!2]$6
P[U?@GS@O\E_DY^#^2-2@@-J)[P_IR8%IDV%/-M9:<Y2@TMBPMXS?@\P:FLQ#J%]/
PDD@E+A$4297>.6!$K&S9.2RPEPH9V7DAKUW[6LD?09;375LAKTR3VY^AOMU3$7S@
PE)U 2G1L8B 2/?>;MCC$<^XUNYD'OH/'EY\[<PM;&H@GU7>"@<!1M9<."&3W#>QO
P *Z<$)O.<E<8,L7Z=CZM!"\'ZVX[TEZ Y;^-&%1;01(Y3Z]=LS.P0P^MZ3NR@T0H
PH36GQ[][Z6FG4W9$RX;3#4-@X.*;O>$O(SCNMDS+'#H9.XQ"S6($"[OHD $@N#<.
P@S>>BGPR1"6HO2F("8-PM9X; 28/ H5:?:(_:U>T)S=&CXU:+GT,\O*(!MS-6\:L
PTV[/.^42HX PU-&<, N&#$GC$Y,.]]4@AX$1T<098+#EACB_5">4K[B5*AKT=(<M
P F>1)HN^%=D@4HH;@+JHO-A[$M,9!"D-1S[4]Q0M#<U81^I!KP5';@7[#[5_H"TH
PE.GFOU^L]DB&S><07=&I2@BN#$[M558A1$ F)L>JLAN 3DV=UPF>^72DE!=LN4G,
P%@Z^B7^5,\ O'X8&_)>D9)$F3/=*8;LD&%/WS\@QG"7CS79NMAW EM$!GKF8Y/LW
P210]!.VX>OL0NO<ES9<\;"4=W&A/3Z442G@_$^(/G$9L&'-+&G%=+LAU*?J;0[$<
P,8I-W8)(XW;X^36T-PHU.4,[1UY%)H$XFI4R4":8_^ED/=7M<>C,KMEA;W&OB)"W
P[]4<J#')/KP)FK4G9F\./WP42>"%,/_4<*HP8ZQ0)SY%+4,.+2-O_I%D=YA%E3S#
PXV[3GB]UL/J)M4JB#9ZC*C!DE-T.EIK!B1DKW 'TW'2Y$F:=*.@(8+D_)3Y'C:65
P]J4'KIB90]$%G,M+B0EMS($I=8;T[^CW,OJF<]-Z(:A22+.2K\BDKUA$2/>$4Y<)
P0\#E]M?'=6A1/,O$-@)*HKV3F#Y>#"_H%BN8ZH<5[HZQ:Y7X]&S\%?]47JI.SERG
P'B-E6K NU'56L \VMTA<^U#W/BK6/&,_(^EAPO7K/N/^?RCT]QWRVZ.(VH7Y]"2?
P2NJ4@U*I2"SD$8^JZ2N8\TJ'RFZ!R!M@O>V%4WP+80Q,)+L1G5./VJV#6P&5 2R%
P?&,<)%])GQ&!Q^9Q:!UY$:]R1A6:%)D@TE%/C@(KN_:WJ8'7VA'#&JZ;DDI9$$WT
P+0$,<QW*G!1ET:=\WR-QY 0'7&\!T,B CW(!:1&,XQB?/26H<TLI%:[*1T-]_01;
P9%3R4J\$+M=.;#W2N0Z7B!U0T%&O+$@AV!E;#[SS@H(^9.7OL8%JX/]H9;><)<)>
P-H-"#30,&0RJ4]0K:+]7 R6;60FS3I2S^LWJX%BR'7XPME]\WVN>%9"[ONN09[V.
P!S?W$VRNL2=G.Z-S"O.:)?8/YFW+-)!6*.[KIV5]SX%YKH<LF=.Z?++SBM#'.DOJ
P##!Z3#4K<ZF;.DE(#^5WI'>8,V0K\W,X);Y%B\SCCU0>Q@E#X9@LH&1)%)3433_%
PYTB<ML#4*.D5U_\4;Q;TX[6G 9L[WZWB1).DA*>?_#*)0F]53G&' ,44VDA2V>_3
P!WB_!B*"EJ)\QGAX#VNA&?S!BBPVX$;;\F?11WI@F66CQB$J1HK'DXM8KPUA<]*5
P<_"S$4$6: 4P+$')3S]I\ 7=K=(V9RCQHDRD;>V<*)]).V"0T*2^!%';"_YWE7AW
PIE+RR&[=R=R'^YTN!P5D_OC/2H_Q@=@ L0M+& T^Z98<#TL+C5S1QO2T,E]*;4E#
PKMV$CX$IG3A_';%B@[5XN_%FAR<T1<\O7&S9,'HYJT#*\2C8O19"O@VX,'O7UYN=
P4D@RDQ]N.DAK@ I#*9:WIG3 $#T>E,ZNY<J0/]EW:A9'$/5.(9M0PM(#DAIB>R^<
PX5"2T9;L%9=9GS5.*8(Q(-=&'/"S_]OR)0]PS??S5OR&7D*4ISQ7"X"%UQ5TD<:7
P1J^5PX]4K.EY]&FJ&*09KF%\!U#'[^&&8< IHP2I !-(C*&^A_S@UM-\:]4T^,!J
P[38-!Q:JB^;TNEZKK,PIWH@I9Y95+:RP:\AU_#A(%4Q.['JFV@'2D30/*1#)-O0#
P70.1<V40 Q@:.:>MBC;',M&UXC<IVKI*I$9&L2@B%>=!G5^F4A(#/H<^3?-DK%[4
P@<)Q8'AJ7JM&.OUP\V;$B##\Y;A]?$K.>7@XK(O-/HX\Q%\HLH[QA]&^'7H8@WET
PS%]V#E:RG4410B0W+\$(&")SA6CHZ_ZA7$2V<<Q2F85AEB^1XYUD),$$<D$T:^S>
PC*QAK@ W?J_FCZV6W'T=J&#DC)'[)6-#>OO>%[0%G K6,13!$?I[K5_6IVX>K0%J
PWARRTR+OX4OP*::1X1K<J>'V!J0Y3:$"G7 #A;,&M6839&XSK)G+V-'UAI%Z.- [
P:(@.W#T"?C3F;=XT"LPH&IFH14CPEY<HUVY$7*;TPOW,;]BY/6U3*K7)#]I*T>]/
PQUX%V-L\]X;^+D$2 I'7.TR^L>! MJP4IAV8GKOC&J:'F10A]CDK#AHC;):7',',
P>),:4PK?1P<'BTV<+,['S_<<U;+[7C>:ZZ^5,PG.3\H-5<\IU_$@C,0Z>C,A ^@!
P2#E;&.D&\-K20S@73C\\VSPA5;R.1R]=]Y62!^\-2=+O\3I$IX6=P&3AQ>B2G_(1
P;)"90:F=W,4)B2#&WR?D'N>8U6,XZ9QS_X(!IQ3*6< ,^ FZ[#>UX&;?&Y0Z@S"M
PU'_SS7IWP2&A;.:\K.(#;F@M?_X"L ](Y?=NV]KNUB[S(ZXR)$J[Q!;:2PL?U0B9
PQMTBE.[#=J?GY2N775[M@#W0=Z2(XHT+)"P:1B,'EZ65<[S>HPQ$J=46.X#.X-:0
PK>-7QY)W?@7,\@#"3'SE9Y"1U.:I7?7F??W#]&E[_5]O,[OJ*:*E[QM\U+6\;%^:
PX<] ]B7]Q$7@$F07LMGZ3\O!3OMJD&EI"H<@)+&#-67$_SC+G9)B+Z(1Z*+'4X$6
PO<A]Q)04BLC*!(L:*I-L7=JS%<=-9MH'E ]%I^^&%T]HVK)K J@TAE6.</Y[W= "
P"@2G+C$0(.FYYQ/QS'LS@LL>E"#'\'P'4K5-* 2.O"_P]*K-KUJA\13I;S-I0P9,
P&3T7>W"S7H:DPZ2*90][ 69L. B4=8^-*.)F+*G-3\AV'?49=4'5ROR;>41J%9;^
P(3G/>.3=$LF&6!PR1AHJI6Y2@_-.$]S(L@#?:K*T:JCN\]H=Q/O<IO0E?V/^>JD@
P<+4=AMVH]0P%,HKVU$OO"W[Y=KELI+D<#><:?&6>**$[E'4WP(4<@R;,4 !8/DY[
P%A*P*R1AU&S* &SOKP)9'"6_^LJ@:M"/;0.Q0($5J\3P%ZW@CGE8@^B!9OZ$R/OR
P3 +Y5H1%S ,L %6HJOZK<&31<!AC+=3V?9NR'3"77KQYR]LJ0=V6Y<APZ,A&YO_6
PKH>8@620F\0'X 4G5K:NRU_;;'QH?,Z\BRR8FF-@YJ[4BG1N<7Y5#SD8#,2GF8Y"
P9#*V;0A)02>QBJJ,,2>Y3@R2\&F3.J:I'FW4:UK\@O:@HN5)">*X,*2#,7XJTA<(
PZH': 8/&%2J>GJ<TG@5L_K55>)@+'?CD98^UBS/R30N@&$@]%*0;BEQJVLD&II<<
PD@EN;%&DSHI@>.Z:P^2)G*T8C7D2R584^B8)S&D6F$.C+[I?'7O6G^/I=*W<7QRU
P$F=M>&**BOBQ#O9C N%^.?/:4J9/.C-D"_)_W$7*+3><]F&<;9P%+$ )C!PX[3I&
P=IU,I2[-SY7R!/A*SCQ.M <<7"W3 )0E!A6AP'XS.?LP"71L5O6)BB6XU_D!/#5$
PL#!AE89*7]C1T!YT!;% _ZD&0H%E:Y6 5,VFQ>P]Q ,L3VMKSM6'1*?Z"0*P6;.#
P@SYH)6S*51[2,7GC8&4YI_/]W[NP^C4J-S P.W4U'=44$A?YSD869*_ \I&\D[(^
PRK&*!6_"A]@DSQ_K.7'?[%^_,ZH05O>S7!Z;9K;NUJC5!&JB$SWQV2]]M0_EMIY<
P*_];^AT1[,:4^**1\DO+'T9TC-R<,J6EJ!O5!7IA RW9[!/GZF8:),!LIZZ!\(7_
P/4_L%J VDX<=/Y,4+X"]J:5[55'] *+F30$V7CL]H&[O8M<!(=,C<!7&[>>V%A4M
P2*U.)JGGB2=$I%8C7]#@7)=TLM)UX7-IIF'[:0M8E+Y67$S-BJ:5#C7H*#H*[$>+
PN\&%N8Z+-WB>R^_@^&.'XBY<GF'<^CR@D^]Z5F1,Z"<KYG0*4UCZOFM%Y[M7ZN5W
P!"0EJ4MO%/',.CFA[G-4P!LBD; (!2&!P 3Q3'*O;*@E</:';X9*1<E<-(?MB18-
PV5D+S"W)-_,KFF>QG]X4'"6OGJ;D4P_Y4S*2ZIW08?K5XHN<.H=HLE,JK'(EW^*(
PDUP6(7L,XCIQT_@S! ^O05.]!#G/D/?)=W7;H]D][MV1A$BZ.#K^GC3ZV_5ZHL./
P7O;#U[-0:D4,4O/^@.E]W^J0P7H1%K5B-DO&5%N$G)0_K,FME5_5N,FTS._K:/#G
P5<UY#/ AH[^9;F_O/JOUV/EU[DE9R2T_DAUG+MJG2%+Y61*%5@LA3LZ 0)AA8F*U
PGK"Q?&"+$ZH/U/@RVTB%!X8SP]XH!^.J81?RU8W W>Y["IK15O^5YMDX^I%#30$-
PEF>]%N5TE;DK,)6;U8F_\(#54O&HJ$+'P5,(ZZYR.\#V#[ 9.%]PCE@=L> VD!15
PC**@_KTK"/N!S#+N;;=YB7*ZC/1I6$8$M\UZN)S22^ZT A6BF ]!Z[GZDUA5OA%J
P'->-6/J]TK"7? <,..@>*4V\%*- QH,U[601V0;7)G?F7J7-JR8+D[#\:AS<FE0W
P\!\]\R?QM,%%YH?#6/(C4UFOIK_TQF&S.P"42)YV<XBY>B26#VVA2*_%U7:E9S=K
PZ<,!-6/4M,U$$:Q&("O(3'$B&ABIUV")4)6G\PM,>GAR_V/060^L#<;6BYC=0LO-
P&8NCL5GO33$7?W$<;QE$>_\Q+ !+*5XMVE^-U_)+_\+';>:M.$0%Z QJ;4:D)AD<
P6X^BYZ^N&224OHP#U$/AN/+6">Y=FN!IT6@/IE(YUTCNHN;VFJ^1J+62FUB^T!1W
PYNJ(#K))2]:+->MEM8JM=_)O\G)'I"<DZ86(H[U,,-TA ,K'[V<C.3ATWVRD]M0F
P&"MUG5-8768YV+DYB8?N[5 \=, 2\[LJW5I1NYF1VA\GG^_0$,.&T0[RKS1-'#Q+
P=8(O!V@LA"HIF#Y8.DA>IGD0AFX1(V;]32,?"W0?%A1GL^"_VYCE:O+%AAST,W?;
P(>DLK6.(R;$!_V9H_=*61?<NYF[("9_9I=6]B]\+_$2TN),X<N9C1D1S@]<JBZ<<
P)< \W7MR0NQST6,RAR=^VP^AV%_&'>M8#I-MSXU*:PZ(6"N^.0\P/GCS+P<M\5<)
P>'\;H+<#PJE!WMW-<7YCS/1'6]3/]*&V2&F28ENH4HJ+]OD1VF<_X4!60V%_TF 9
P>BHR<$O)KZ_F/7%K6$4[@Z7+?S-ZLK^LV\WM^Y$%;'CR\?2A)PZ/\\ \C">+?H1%
PT*_6U@Y!*BFVH4M+/!*AO*2NPLWME83B&7./M1QHR(*<D*/P/1T3/ZCN7;\J/ R8
PH[[K_[Z[7X/SP9??ZH->@["9-W:HZ,L;;@;2I)"7> %%TY?+QN]O_[.GM*W$XOI*
P2H,6T(;<E-K7(_VODNK<3(B]QK$H_'T*Z'1,R.07_?VE&/3B9#< 6:!)J88IL@LL
PQZ^O6FKO=FSD4C1Q-2/J(7"VW4XT+#UR,#=<RXS31+R^9H$:)AQ).^X#UDD!9GA$
P";GN#^['!"2=,0?SBLTRB[WP.3V/YT-GX-AE*>M[9G\0-COJ)$E E0G$S+OC0;;.
P#=\=O+3;6;YH090*LI##9I]ZFS.9(+OA8^]GYT2$>X?)<U=:;)&DV&W/A@/2W(G6
P0VKDIT0D7K6;14F[I.- W:S%;],9<=$G:BV,LO0J&VS64<P[0=I8J4@W0JEP/+3J
PR0F8=!HIPSUO3/@%D3S%^4]&.B;#AD8A[D86:F514X\]N]<O2FLV]AFH"5W]@%-W
P0 P\PL,!U1J3;^H;.6%[':Q*ISE1ZGQ1(T753+W?,DVIS7F.C%$Z?'[1=BS(/G]Z
PKGW+N<W&(%G%$B/6,<C_E7/5#W0LJ1'W)S8#0^UOO,YG[&4]E=,GJNL'N/&*V _S
P $ZMY?+-KW:2?1B-JMXU\0Q^6@CI$^#,4JW<-!(2]H#-[TNF@ELX_94KT#JK;80"
PF9,Z\FTV66?XQ,L ='T]HY;.,(Y6I3 !#&M-6K<IRM43<!\5_'3&4(RDZ8&-H(B$
PP[ C""'Q41FR\^:5_ G24^93/=$/>]*W2-\ C:*[1@.$U6J^O-DJSM_OHWP89!]Y
P@57+,Q<#/S1\<Y6X-+QH56^8,@U_UD:"UYQ_]:]PXI)@M/VT;U9I<M.X/'*G>-MA
`endprotected128

////////////////////////////////////////////////////////////////////////////////////////////////////////////


`protected128
PDU7H_H3X>>IRR,/N?KT7T<0-(GPPGNX7S)K2O6232&=Z/G(,-RG>ZRZJA ?<O-9I
P'(PYU"C>U0.Q;%B>WC6/4HC.[V1,^)A"QOFL2+GS#V&0 O/LF@$&+0H:O]+<784#
P5JED%HG$(9>&ZVBN;D+.!TY6TX4\EQM:7I3QU0Y-TRKPH4I1#?_/#EDX8X1]J'E)
PR@!+B\[KC.HU&Y.^(8*U*]'K0I0L0[J)O1#)&.>,"H?=1_CIWCQ*I<TPA:,#<6"_
PIHRK"",*NN4N)9,L<*]ILHIW/4Y9S\73-B^^XW8IN=JW-$KCMN=F,;@"?A\".A%W
PY2%#5> 2$2JKTPLD(5L?7.X7F\9N\*H*X;[(D_J^3,,&(M)T6&2EZS!G!$$JW,7U
P8.G#POEY!?=)UL'9/J;_0@6Y\U@7_**U3#*C#_<H+KKO*\<BIJ2L-&IVO^"5M/5G
P$H:J21A3$ I9'?,41$2*\98GS*IQ0\JT>U_N8-L>=7$?6"X7OT//+XT[%5'"*=[2
PP-E@6;5UJ@ZE!L")-[ IU+Y*DPH,"6)*Q>!XW!A"'L>SWP%"@+R_](]I.VL[]?^,
P4-%(YK16BJD]A1ZC@@]"R*-(\>H*ZKYC.AV 8%:F4;)-)"4EXB%A35HXC[0VD6'1
P^\L@3PHHM;U=V.>GPX#@@#5$6=5X61OZCL4S4*8+/9!?&;4SRO&2;N(90NNUCHX:
P$QLJ$%KT[.0O#FDI8XPV >"T&PN:/),8<(.IG/C =D]&%2299C'\+8W8=I+KG5P7
P@+L.*Y%U+(!9WI&WZZST/>90$I?[</2*09AW!&<OT5RP]&J.,@F&ES@*VY8/:>NP
P4F@O?):-AY^PU\!M:90(&<_YLDQ8P#U"/HJB;'@/KH+J"GT]0+>HJV\X& J(I]M)
PT?/?I7NIN2]9U<GL9SL2EDXYHY>>!4H[@5TH-$V7AOF6R+?W4B.'=0J2#@L_+.IF
P0Q&R[BN*:D^\7FU,F1R4PT&RL3U":.\F9]R;(=.@\5KIQ^J!6)##VJ.2,ER.WVTG
PQ8HNY!EC_Y,T(F:+/ILJI2_Z\I>[D.:?X%E<E:*F IX7,M4_TVIW(SIV3.PW>Z38
P5V5&WK#G%YMXV/MM4-T##%41QH86%UO=D[]J-K/WLRY=XXJ_Z$&TK74-/O-D'3;P
P*:B+7[[@-+S:]8/]';*'5H2WQ@=,Z+2<FOB 3"PD=M:&JBS)W-B4S[8V$@!7RD!"
P_%96-R3!,>_?LR+L:"8X:4DFUW*IB9._@2RK\+KNK-0TD-;H@]?<Z(<QUE[>)OSI
P'</;AB<F?;A=<WR@4:\!(^,9-[UB,0_S;0(.W#9PF\&EK"2X5+;8%+Z(" PLY\2[
P.LN/<R3ST+U1,[V3;25[R#:"91IWK^9MR:IY\(4RX,^]C@=2#,)M;1PVF+[^!(M!
PZ8@[+NYWDV"CIG+Z*$&1S>S!8U 4&VJF+^&,-S\@GGU.#B<&QA>8XQ5A'\LNWV)L
PI&REGP0J)J>_+O5:B!L$'G7QATST-7;*(5QF[HO9[9632-;<\)<6'VU- &(#/H*;
P.2KE9M<9F3*7,_>0*DM\2IY)<]DTN#G]]GM@G:PU!=3*31LN]^2#M$ET\=D*3HK?
P^IY$JK9D5"H]?.P&37G#2+Q$DA.3-YB2[V:81.Q$#K%Q$-E'_)2^1M,-*5',, I\
P0>\R=NY$N<A%F)R ,$O"QD)#\)*FZN:D%&5;NKQW(SS78,IC^#KK041HD71U7T/Q
PA%^8/J**XHG,N>>KY+NN)F'M<-J!7;C!7>O+5U$D6 AP:55Y:W&^M/,=?B79U726
P"AYF0+Z[ G[MB_ELCY_:(G7HA C#9DBB]*5:',U&TL4J!UX5/7:0_'3=&WKFUL $
P3R\K+X0L \),'*3&A$9'>#I-D1@?\/(Z4WZ9H/F@#PHN$-0M%?ZJ;;-,- -<;[\S
P81N%Z!]U^/!.6;-U.7&UQF5]7$YQ$Y*!&&'U$KI8:/TE649R4[,9!SFZ%R6>ZZC 
P9OKCHMEWPU!WLCHPSO24Z*/<MM<,^"5"4NPV(^DLXYDN\Z((9S(ZV#6D*/X)>,'V
P?BBE1B02%;\(';"\=(#"PB_6'8-["2M9T7RR6">ZJQML1.I5?EX6S\OF)IR#_M/ 
PV5=OI,:T@9TK7.LX1U,3CT7_MO-$\>"H649L=FOC=*0(+V104N7-C>^S([B?8E[%
PV!3C8J ^F$A/6*MA:N$ER4YFC(8B>RQ,II\9[^L!.M.*1DLKI20=/ZC$1-WH=I!E
P&KA42G.!AO'F! -UK@B,2'P^G8L=.6VXN W0(30I^9\!F:J=-UXN?'U:E.E^$J7'
P3>C:KL0'OD]$,?!9&S*2(ED1ZBG.9$.L+=11=#K@]G<*GF55BO"&UA,M^NABXTXL
P!$(=AP8O0&JNRZ$F@(8V6DTH/F'*\&>2TG-F8>-%I9[IU8<$-L_IQ]JF%Y,!7!OA
P(O^G]D$V&"V[<;>^&D:-]"2/Q!CAC[%@[/B$" /LVK]&[?4B2<=N_@JG-IVQ*9@W
P:I2N-Q!LSI<LA; S.4D7!LGD@"?53T.V"J%FO=D=D7@&(NUE: G7RM[%?9\3=O(L
P(9NI=_RVUV0?-WM _YT94$BTD6"HD3>C]J!$@MM\4NCF&'^N@S%,3"%9GX8*XE-I
PG)+D'<4QNQ@,DYHT*'C"A$HPGJ&UV>P1+TJ@EU;F+-"#%5YM"_W^S5X97Z-FXUS+
P+WF!?\'PR-1S0A+[K$CRR(>?ODY-*8 H,S+FKX,4G-!K69]/"*9:O1[O Y3,^$-+
P?&+#"8)V[%[>VSAK?"'DQ8$SH0/[Y\;M><A<I:]YH*RW) Y_[^]C50%<,["J-A$!
PN*'WT3!^B_:-E5"5&];_5O=<U60F<S,LJ<M#DA5V4\+"%\W[;JJTX3XI=E!ZM&L9
P232@"=L@]9[*DJY4X]X_6#]) G*S+6O NH*S0HU-.3;41_9,L5<GW\^M&=0V+GKG
PB'AO=-9"U'5@!4!?<X9+:?QE"W0OH95 \4R0WO:O:0HS*43X5VA;A!GY*/N5$;$R
P"!N*4/Z;#B?((-@1=4\=+.R:@_0$G4,Z'-)@Q/,Y(:V%YTR3D>$B9ZJP8FUF5?B5
P8"/!P/=;>IX.QHNZJ":]ACL@VH;=B7YMP/JF>-4BS$:#/[*?G=.S1DF8__;WO'(P
PV56!]AOSB?@4Y%GU2&GJUNJJL=MW 9Q&/=B_$UA'9L!<'>HGAX.C[A;Q)B1^)@\8
PC*E_P)!B@MC9/^)[/8)P <R6BXGD.7O7?>O=HB9VE2! B=<:^"2MHQ:>+FUS,B1]
P]6=8B>-QOOU6>WXPV]CQE9!!][&X@JM1[///+X:VV:-;+_[EW1=C6W='5X<D':DS
P8H^/&>A[6%H=W\B,!+'L'<P2R!L?HJM#JJ J&I:-'4<!NN(P L[%1#\T03H)'GX 
PUOUFA!:FE8!'4$JD6:Q7!@WX#P99QZ.H)=)B[Q+5;FI(*.EV[RG_1<*F"L51/O:3
POY^=/Q%8G)!=N8(BE.XDRFXXEJR]H%/@N,IS.L_%IT"OA\V"4T@G'_@\>C+NRDZ*
PSX^'%],O_2F/6S4@P< N;[M)>SA$\>8;84J5=97&HFBI]H=E,@ \AF&9IV#8H% 1
P7/N*_WBCR3UU7XJB?XW_%]H!!\+7 QVU!:&2U"'I+XY##\O:>WCLKRQF'=NGB3F/
PDOQ6L4B>$<6N_$.8X_C$*QKHE\]2P *YO5IHU7Y21RG.(J&>?U78_['ZI.UC:%UK
PM$[S')NPRK^:8;-_MM.SPEZOQKISXX-RBJO5XMG)F-MD +32BOP7:Z^EF*QR#V1,
PW3!72%82LG8TPKPDXN!!J-TU+PV^Z.U"->=M1KC..X'K)AE>QQI>F[V@W>B59_.Q
P7@""K$O20:A<'_?@AY5'$."BGO.&("IC[,%DSS?@B95E9>G!4J#(>C4NHH?S.32G
P>>U<@G:ZVBXA,3+Y7 <AJ"YFO;+#!\-24%]+-ESM#^]2@0O&>0_)O\GVXK_3RP+=
PCU2^2]G'DFLW4W#%_>!HG:&2@QTU.#U5YD, FW^D(U-/-WKJ>6;)6\7PA]W)PV"R
P2^].!(J;@=Z%?7:#=UL.>?,3#@]L3U$'BE7EA@N6?V[1YG8R^P$I5$NF56!\>M0M
P];Z+63-/)^+FLY# XD:K(E W@$J@Z"$X-*8 8LLTO68[^34YKJRE_8T^GX=YEJ(+
P#S#[_SKDK8A2"8LZZ^HY["%4DIR9=5\3?DT*%K1F%5JW\A_&]LNL>XHSYAR7]7$#
PET\FY7C,DJMF_F.!,2$*9N!_0;(;KW\ EIZ(B=K":PWF=*^WYF$T8Y(+P0220QT0
PY$>]W(.0J8030CL[&9>UHS;RQ[']7)LLNG\#*IPWBCC**QNV78U?M4F:Z9-XNHY*
PFN7W8@V*4A$"U_ C:6YV$('SL*RXQQU!&5W+$LX*6Y);I3OMS9=RQ&"=)"(3W8#C
P&CIQ$X^CI3$ '[TBYF*,W0-':3H;0H7*XL?9,I[#47NE-J/K\(/L4V%+X]<JINVE
PN>,(_=ERJTOH[$ZAC[[CX1I2RJYVHE;ZD(]HA"TF;UBEYL- P4C?7%C4X'WZ7$A:
PTA==3_+&F1FLIJ=# -/<!M[R2'?!I0O"<7$/(OV>)-,H.3.?4'*9)%V[@P-E7&5_
P#;9/K  ^^_D4&1'/3 V-V3RQ!YU[B,!^N?3),H&<\*;/N8FMLC&Y2S+I(%4TXJ>L
P7^OQO:'3NAF*N7\^3AO L:)>O:M",A[-^DS_# 47,#S[4F%E#?F8+VO\6'3X(E_M
P'8UGRJX',IE9 :O)\,_HY\W4R753_@]X5LG>U*[?:%8I-"?/>D?<ZJ* ?X :4U>U
PV]*\][X=M-(2YOU/3+MX1H#=]0G!7NVGANPH-3<7AS<7:C5LRQHA>S&HFLYZD 9&
P@#"EM&^N3)F Q)3MR*!'< *9JL:4DE)%5Q6U*WD[38H$ */E12(06[SYL\*A$?33
P%::7%S:/@N*\#?WM9 2#8?V"7= _UA/<="' DVP$?D!>R' 9OEU:&I_1PWM1?I*;
PHPX;_RR(+$.&F*LI4ND54&$6TCX+DT0\\O1!SL0#BNJJ -+&?CQ]6BVEQK\W#R3S
PJ+CHB <=\>,9_@NBE@FR/J1XU#VVO B4O(L3#B9&<!Q'^#'1&ZQW^O3@9<00P6C3
P)#9(Q^9TG8U;)I4*/EU\TO;0D3@60W1 YXS^3<,XH"%.E9>3>\A!F=PCK[\HA-59
P8;2':RE51F^-P7>VQ.QX5U9$O_Q8U'";/S,U\.YG#%G0P+J&4;BX$@P^F!4D>R!1
PZNZ9Z!PT*AWN6&GR)NIM29>RX7)"NF,XO [EN0P5.&4LQK'67<?&% D#I8N)1#Q>
P,,PQ*V(&Y#8",C#S@<2NYY1;<>G> NFW@DD^2H[$8ZY#&^ C;+4BO\=F;N79B91"
P#(?ZS.L> QJ)_*9Q2N)B6_'>\H=<)))X: K-.V1RR"((T\>RDTKG?)+N%]S5K-[G
PKD4N1FEB=)DTL9CJ6#6!"VN[ 9 LRSKBJ!HG2 1.+)Q@.(PX.8),1I%3@Z\?',?6
PYH"6X[@1X/QARB.8X8OSH@C)2( %U08))L[]$P2HIB$^$\1ZJ_!'VH5E5[N%CR\X
P' -S;8;Y!;X!N(OR)=,]*MO@/I/1?0!%8\RFJ7X#K(> ,:[DGU'((<TA=@@EGO$B
P*%SF :L8J_+4->?9V#EU7-LQF3PN&-8Y/P?8;2I>;*#ASUSJN5-@U_/(!DM5C6]+
P9+>MP@WD41><8+7XVN/W$;K3[ 8>;\QRA!%IB^^ER*+$?$9Z-7 73\>*G1PQ!E>_
P[@H%"0RO:IA:T[5._1DU*O<>6J(1Z!M%CG%C](OML2;;IQ#$1$Z)E2\Y>D82403$
PZ":QER#_/U-I@(X[@(*O)\&,+_LO+.SJZKJH KHQ=ZG B'>*M%9O<%\<H6#KOXF;
PIP9YM\4MUP),GF>&A[D 'N\X"E[OI ?) [Y1Z](_K=P*JR.FA*+N)A<'$"0-YY>V
PS6ROQM'?[P 3."-]ZKB<%[\"37)-[^%^(*42]<+CZ?,K#+<W$#>(EZA5[#UZ4GN0
PYWA8NQD6%3"L$BK37<0YE?&#;JYFJ"4?/?X'@Z>7CZ?):@N)Z],5?^4HGZ$NJ@AM
P;0(Q2;RUB =MIF=/ ^O2J<:H3_#'9D(([SJF*@S!=.DALZM\-D6PKTD:G72)"+L8
P,)GS\S_LX?=&;&IISK%@H:+LJ<A#/8G!2]BMJHC=LG@STB\<EO-^RZ8*^Y0,^!SC
PT30&?33EJ8']CX*+0G>8;K(>AXIM5&_ N=8M8?@L.SFAS^/S+;/  ]:,AVT4<:YA
P_NTJD:7UKL*/YUM$2T@-W(J\QBD#Q%$,A'5^R;&,_)%%*9MG8WE&*,4:2XD$(W58
PS0H%/9RFJ?J@B3^/.:5$&Q??T;OC-,W KG_NZK>*\00?!<!;3A/?_V["(5(,G^[>
P%2 Q%\.P$W$PR%%DAGO?*P'2BAO@#ZY0EF@ZKT_&QJM@SU7/Z0.R:9_@><NX\'5$
P/A)5B8D7[,4*D?)9/HDA\$YTPW>=7Q)&?!8H5@]6.\373XBE&&32W<I1"'?Q[U$M
P6.;?,7K&TX]I.J U,F/JU]*+-WPQO7J=7OB4<QH/%4138$\*[&X*%W)*!7OX=-@!
PSZ_O]8_TS[&@A([3==!_3#A#;65!GXRJAG(]][:=*5K;"<RL<$B7),F_3B-&HD4H
PD!R^@]1I%WSC&&R!_"E^G=9[:<>A%L9PVJ8H']"Z2XIXNW340Y*$@:>GD9X^<#_&
PI;U5F,7G/6>#MFFBG.V'1-_D#X1BFYFG>)H5#^"Q$NXZG&+^..5\I4**S5#PY-FO
PXG%TS\*JI+G[65/$:&7HM]>*XEAP%L4!>NAXY?O<T:?_NO\.':)NI/G8ZFW4Q&7L
P,_DBE4&0ARZ6R"H&GF:?^[+NMR"T]%A.B1O\N_#7+&B3U2S@!C?PC6DT@'V9!GJ(
P#ND("T[A&N[0;N/JS',C!&DQ TNGITXI2+URI;9JGA:\Y G?O>]\'[ 2A)[J/I@Q
P E7M$6;!E#:-Z^T)0RHHK30<;- 0=3(JB?X8G4NHL+<M[D\(I]^E,3N'W^ 1ZKJ2
PD#JA-MR4V+/&0(+3",%!Q4^HV\(V0V3WLEK>D"R'4R0JEH=YG]UMY4A"N]0=2A"=
PV=*<]Z*Q)>2K("$6X<\\LA 5="OBYPGJ.(ZPTS@*?7$G5;P6 4 ]Y NJE=N^3T:'
PI/EL<->""%@'\1@'Y*5V?7NH9U;$*X,4O6K)';13IC@N8I?:?\8MO;<[!@/ZABF>
P1C+=IA.ZF:Q"1<&NPJHTO6K2B<\3J%\3J2#JIY]+W'D?<%Y]3?%EAIT>9^! -L3/
PT*C_*PNK'4A#-<5H(SSU2\!<X&^\,4R;L"F=!$3S)F5!.=1S]E(<N!2#MH,9,[,H
PB3#UZP-+QA8\1Z6^P41)ORX/'H\L8:FG@DXIS3V'Y:H)54H.W#1%#8+9H.CY"8E.
P#-^08/ 75?PVR+/_K'A4\G4Z:W;D*?>< 6ZDHKVM #*".[&G=5B 03]#T&8R_^50
P&>BIN-0LXR$9H%TQ%T]?0EM%Q[20;HJIY!UL?%E.FTA#1-QLEWJH4?+\1*"1;#*:
P6X5G-G!4P1^QZ7:EN,7E 0(41)"-\CL$WECLE)N680[OWXD7=Z..UYO'OB&&67B"
P8NY/_0;2PY ^_;)YV.+P]Q A4,8W6AS\G3('LW3=<^+J]CGV&SBR9I@=W;9XNWA4
P1#*F_%VKLS,%CP?,7IGZZA6IA118&,2M:_EIIK\M<$JH";"T@T.@<@@LNXNM<TFE
PA6QW'#<2C_;<-^?C?ZJ>?KKD6+TNXM:_\_E!DHD:E ##2V5USZA!8#M$_1N<HCS3
P#S'(*=^[(X:)N.R>]98EY1*"]Q&NYB8ISA9>EU"I&C-0GW4[Q@ZH?YZA(@Y/?D,R
PUIG7A;]T=Z##MVA&ISQ<4Q/L T\8?5]Q=T.@_3)+&^C,BG/3L7G%6F8VTAQ<0IQ6
PYG*Z<O*9L"9*0=\+@S/DG\[BV!-KH4M;0/1Z8Z^6='<JC?Y8+_ DN[?FF."YJ5=1
PG*Y,<Q'B7D.QS &^3C&CM9K8Y>L#18O[HH88"HL?["O!!N9)*H -S%OC4TW00$4R
PTT1G&K[*,GP_"J3*[]]/_B,I(WR[Q?-<4:VXK8_ Z:!A"YO/R_E[H@AH&OY&T<[9
P HK;'N]#9P$JU\$:G*QZ>E*+\>S"!.@_&&"^A_]LM7U!T K/HQY,=IJ1&4IK4B,]
PB@K#1#9W@1;_<U:;4=F:)L_^HDC8ZY9*8DKL6"AH\ZF"^S\#'M8[ZW=DYT4B/ET@
PZ_Y:[N%N0(%!'__FAZ^O4S3IH6I%<8,!I#Z%(]SZ>/H+ES%9+.">A*Z _9^R^Z!4
PG /Q1&>A>NR)6M!TCL*Q =*M*F$< KU7/^EH6R#LV.A!R5DG_[D"Y.Z=(;HL-*9'
P&=VQ2?$M-=MHYDV14-'8"!6O4A3'6?P38:!*/+(K8DA3U#-ZATA$/E4+D:VEM5_G
P]>CEUDC5';8H)>54?;,1+OSO;HEY8FY/:!8!13G](UU]0=V!!GTK UA6;8P:8Y?4
P8VD 8[75 =YOU#I]E[5)Z8O$A^KA]K?G2Z;QNXD,S?9&ZT-;%9?N<=63' 7$11?Q
P5,-GGB<EC2J7*SRMR\T(\!$'+/)O02&P(!<!F>#W=RXO*,E.@(3K5 >(:SF[[XSD
P+8C((:)T>1BR#,DA.OBB?Z$8X5XB$$2N]7U!4=?28 LI:PD!K!(D\1JV ]$P[PAH
P9P8%1C"V<:BRE^N&DC TOS'RF81YS%I5_PS1HA8'$_V@MYKA%=SP:@H,/.^<#.>,
P>(33W//\B3.T  5+?E@I3M+4P94(5PR!EF2"*H#\5$$M^;Q]?Y4RY/K P/21U8]]
PFEFWOOI+R9?XJ_GJE=D_B)+@ Z=8%AP1H7&%R8>-VI:9.JG2C\"_BE<5EFF7D$F9
PSO)4 F%Y6C5RQK[+7D:\4-E$7I%Z8Z5/DPSA >+;@;%+3R8$>KOP^>FQ1SKCFV^]
P#@R-1@G^+GT::*S"9$S_^*O6WX5%I!M-%VOE#!'30, 7= N6N'JAW=0(DDP'CRP/
P+&%^#(^2,OI'@M"'(H^I*<.\A*3/BWD^GE_=L16[K9%J[72I%+8<"'4(R'E)B<9O
`endprotected128

////////////////////////////////////////////////////////////////////////////////////////////////////////////


`protected128
PDU7H_H3X>>IRR,/N?KT7T<0-(GPPGNX7S)K2O6232&=Z/G(,-RG>ZRZJA ?<O-9I
PD!&DT(D#(YO2QL-LJ>1$X7*R+2B9;)0XH%QGFK\;"/: %S#\1 ;$PB[OX-[AM]YK
P/3;K/?,: ((Y^J\B,D1CXD8P6SCF>,'? ONUL[W!"GA O3!A0=2P!JC@O.N'Q=L;
PN?IA()CX<V,@6K *(1KO793SK78^LZH<WA6'-(C[0]$(*D#D+C3R@V .5HF1F\-;
P!UVHP#O6K2(]-?S %CN":8]Y_?7Z9F)H^/%V)776)B>^VI@4Y4!U P2<]'T^(;^*
PT^3O)W91><I/71>F^2*2 Y;BYP9:<LQ@M&AW]U=B_'R+^>PO@6KD4QPS07)I"$E=
P3#C'+25&3P8VP:G*$>/OV3(EGFCD:?I&P"/+PX;!%R7&9J2]]-X<2[XA)4YVN+,#
P7,L1L0XQ?'$^M5@,=D*)$U[0S@ '=-_)8:AG$G!5<6S)H84"S[/_"NK+#S9(I=AB
P.Q \I7!M4+3".E<'+7Y5+F?"'":SEQ[UNR_WVG+M HMPNA]D9ZFAV']DS')GTZ&G
P0L1>?6>UFECO./.U29%E66[:@A#M&,,WS4=EV S(0K?1!;J(S&$W\0;?Q#BL?>JU
P/A@J:K(-+P@Y&D"%B*<_W4>%KF]U#IK37L04SD=J4Y1D/CD%MMN884HJ)HBR @<7
P5#QQM6%S%\YX+9EK@3\&U\, EL3RW,<*8#UF,*=BDJ_:<:+A[/2Z>?S8;6&V"9$;
P7O=141F_:;KYZLI&_9;= R/=,?/-N;"C)=^:@IU86%&&FU9?5._B>O1CR?>AO7N"
PPZQA)%P87@?QF=]VT,!1W,3W U"]#?9F'@?FS5]>WQ8]&QL(A<<_[:2P= 0S3Y(D
PL!.P)3N4J'E#FS3G4XA PM+ 1;KRV;2^1!V*!^$>G6>?4]XNW/T9KMP^'*A6=46M
PAGR&I@#0/T;TM-OZ@TS.; N@$]HT9J_HC!A?@1;>KVJUW]^;6.M/C=':JX=@Y"_G
P+)UQ\"V()']OC-3<O@VX7+8;7IF$.79V][LS^)<E-)+;J*-S-!4H1B'U;J$+?8*_
PMU_.Z[&3)MA<+BNK_K:1DC%)6 ;NCL*M$UL)5W[S+0K(@_TMIY^+*O*/<TP>^S#M
PTGNT&4_![J&:W LWFVC0DHS+\LR:-A#QX)9U;*,L_3]$'51)&C!<!KB-6;"<_5[H
P4;.'Z.>;5ZX[^]P_H$>:6#+!N['HB1U. @_3W'=A4@+U!IY8O<U.[D$80L!87?0.
POZIW-(0<EVIV&DW56GN]#<>!);\$8"3,[LQM)F#S-?-,OL]Y#52,8U9R@RWC;FQT
P0;$J5F_YQWKKI^B!6$GWM_'BB(5@4E\F2KK^^?Z(!?^/.Z>R\:B"#1W7XBQM9&'1
P5?D<AYAE%J@35T3K#S]9+*<'E7F2Q48032G/XX7#:KX>?";'F>T#(ID:)#"<8;?U
PT ^1FIQ1.UMQ1I9^\\H1^/>^NYJWP B'3,'63G+<HUA2]NI)9\K5'&>TWZ5_0]7#
PM"[2!\J*C\!6!YUAF>-76&I1&=@<?-O,FS ;'H H$]?N#U>!X?-41QE&CGF=I,1C
PLFZB9ED!T@E;;@ER +W6V,/3KBN&W*\HZSS7F.'LH&+F@Q#YXI,:8L+Z8%NG5%8>
P#^#,6.=$J:GN@1/+1\=$+"'UMZX0N6;4K6Y"?8BPMY<>250')W';++H^! ,33KA,
PLJ7\S:%1JB1IL\-:*3()87MB2F5_Y7>;%^Y4'?!6JGQ*U?MXNB^;QE&136???,14
P:@ ]OLE.NHT!>QXHK3<YFHLJ^M.]SMY:4\5TO+WC-7W4$:IH^/*2;F9[JF9MZ"?L
P$#'C]9^E[B-"B4Q1H0KHS 0P-D=1%S*;$[E4Y3$L'"2-[4_3@&H=]LTL4].<&/]Y
P?W1)7#PJ9H:7V)Q ]_T/D9F+%%SN;=^:Y-M& J=Z5NX12CE?@_+JUD/'@6?,\DNT
P@1CMZ>$87+O&?HEXN["S@XXJ05X+:)D2+KEO!)9A[: #M$RU #PZNQ4=1)IQ,M2+
P(#TQ-)"88E\.,?P9 64[]_JGS0<:H&:_UW!H*457\TR-H]B_IT4K0X39E=*?'!$U
P35I,K5\-.6"VG<JJ@T#X<WO]M[&VZ>KK?EC&"T_(\KC$M1WB&WS!.&IM3TC4W;2=
PH#96(D[U";HGE.2P 8[9P(+32^!A&_^ZA=7[Z72VT#E;76VNH$B@L(VH69UZ$A*$
P,]I/:)?ZUB%HMZ1']N&M?^C()F@?T_6IS:H^ORXSQW9&9MHGVNIM,5__,I!M%CH:
P>3\3#A+5(.=A(@ZV(.D8LOG*HUJX8R*JM*W^Z:CHXA;NJL@ (^XF>JE _SO>W\7%
P*'O[7W<Z$:8IYNN'=5@'(8#06-]O@Z1Y1U1/8(QBF-@(.LPQJ\.S4 73H^.&Z&8F
PA%HY"G=B%1('4+G5H[LPR6T4DH]BJEU=%!4686BC]&6^A"046_'V"R&H\A_FQW;R
PBN=V/3\,%\.$V5 WPG/<+[>(EPU,-A3L A:_3J-!LK>+7[](_<;_#8OX[3-<H;#0
P'.&'AO4XXFG+%$L^)@]1.CEYV]X^IBD"+\SKF)SJ;6H\@4"]U =&'(-=*HROH3V*
P@>D.@JV^SH>J/N C35</+6H=S)%!W&J\B21PUO[^"[LQKJLG7JC),C55%*0P/:C\
PFL0-QZ_#.7X-X:;@C-73'L"A+CL9%M2P4U>[@_(7%[@>Q,&@'A7/<7$5I5TMA%2C
P?A'4%62H7 6MHB0C5<,=7<Q5:RZ3F80V_U5.,*I2:H'AN1W)PQN/(M7\,O(^;I!D
`endprotected128

////////////////////////////////////////////////////////////////////////////////////////////////////////////


`protected128
PDU7H_H3X>>IRR,/N?KT7T<0-(GPPGNX7S)K2O6232&=Z/G(,-RG>ZRZJA ?<O-9I
P)6V2^,?I30Z0UI;:@ -Z?*Z!CS^/3+>IJ7:S9%-P1*EJ-<)XX$9-1.9#9E5^U[W/
PB-4$ )+QO2"V!:33MFA!P0H"[)*B'(,5(B5,GU]A#I]C$V7"@8P! E/B85^)UP[/
P-B2M@UP37NPM*74Z&&Q*#^.QA&#W0DMP1^I ],VNUEJK%XE.&IO>KXMCF-'"Y .Q
PC/[USJQEE:MH9SSTN<D*_G(LY<XN-P8O<&ZO^6H6T<,1(OX!'2;GPE:VZK9C;(!;
P(DTM^"BN0/_,>I99C[%G^($:7\TY-E([;3Z20,C@XA1R^:9YF=(NQ(B\4 )Q73"X
PYX2O)."?BGE'L&W$ARI#LQ<?K+A"[T>('&#2O/F?!OGXF>U)M=B$_>$XS!B*-=@Y
P$/GN"7!>*XP,#6<T<U2S<'Q997]")( ="X\=RZ08>&7I8OS[,->O%]+-*&*/BIS!
P(4STQN?NW 1YJ@HD7O Z"[XF@4/'N1/ L(3M/[XZ[BL?S.,:L-%YX5;(#S([CGPC
P@MP@7RC^/S#!\RQW.,9V5V@WRS<,RF'L0I= .)=EW%*GKZIOJ(-$66FS^F]M#N>F
P/*C.=N(P5EIWFRD4J<&+9_DM$<PRH7BG47*$@>AOLH>[Z_O*M0R:1Z?.&, ODQ3S
P9N4P=R5DP1=0#'SBV8E1"H(AS1*^:$\5KRM8--R7_3K!*99CB\7"F8NFO.YS)J\0
PH]-L;61WV-9=T>FNU697.G9$+SPQ+<LW=O/]LX!+K$%*O\* 0OB^X."'K^JU4(*X
PHDH&R1UP"U2 *ER7TY1YS2-]744W&$>GXHH^1;>EQ!8KD9+QBLJN1;VEXRICX0/,
PV)B2Q(FKNUP!6W"[Z<:_VTEA18@(T>XHNS%^?:R_ZN# 5@>?,7,\P?]2QM5M" -8
PS0IQW>E-J+3:Q)80+SY4RI-Y6J8_0OVRX*@2@GZ<=!$/ 21:LPWO[MRYN[XR&7M$
P8],:L^+U#*X<2S1]ZUGYOG:!;XJNH9^ZUVO.D,X<-VY5[YW'4GJY:K&C2KTY4K"G
P0&OO<P3HN(XVCTY\-@2R^/F[YBY\(S3=(L/]_AI^R3*9%\6U0SQ(%6X&:UK>7S<'
P[>X0>[.*%D^OPL@?L?C<F!UE'6@O?-^JYK0(!T2_<!GGGZ!&(3K/ZS5<[RCR7@][
P 8;);QEOUNJ?P[=;>-*(#\]5TX(34]RSKAPZLY/Y@.BVFK_6ZXM8.\>W*7$;1= 5
P%EC@H>T)[KR+1,!RA;B9@8(+/$N-WC&LDIEZ]:Q?/NJF(9(3;1IDB.;=$GVMX=0R
P,HK;=H#U8&9#W_ <0.BT2UK%+"BLE$)545&A%31J*BB*UCJT<7.U?)J\&[<O7M^@
P7T]_2Y2R\"#FJG<;$%#TA=+^5&P!NP%'WZF6Q2=,376:9%N!KMGITC3LW"177T)U
PM*92C,OSIBZ!P1"&IHNSNO]?V)NH0Y*)>^V<Y^B=:/ FCH^F=#SPO+0&Z2]CPYZ@
PIOG-W&O40D#.4D)3'.W0J:/P("IO^*552_#G/8.UD'OP-C"8"-NBD1Y%2KD"&!H<
P5<OQ"W CM(!AM>7:GSNJ_VJ+^-KBC1W8$D&2I-%PN0'O%</(JZ+)M.9I >H+_O13
PD*Q_-C71<D3IF!H@2H@B0O4U] V<5+* @DG=*MC+?-I//FNH,N_V.W=/;*J A\>[
P]/!L$0>)C_#%2Z&L4G'B(-4C\OM5U?_9X?CFZ6OV*R&GR&]U@L72D7:A8&XNK1QG
PE2-3\\4U-H6:AD#;W'JG)9(E!BPRJ530B/<FA(D0?&>[25)I%Z&HJ$XN1XC<*FM3
P!.)X]7O@!3$8V2BA!3 DB?=9X>&4DP:I*MWNVIQ&CFR3C .8K'PRU+MK@7Q!;GS3
P<(L2E\=UFPL/ *&-L%<:L_T!/0! 2)//&."=+X!?FJ\P>:6=$[V,LW Q;:1-9=M5
P9EO?+"N6%TXK1ML&3SV8=VU ^NU*3Q@/%GMUXPW[M^\L*P&MJ1V/*T.R_2K;O_X4
P9NM9K_2 :;+9=DKMA7AQ\LI&G@B/F8!@Q BQ8+6%12[*O>A[M>$KHXQ#_K@2'I_6
P'1&U^)W+PX$<(K&%K_02M.TUFM.8W&.,^KJ3@_Q/<,\@;&5>0VMN-VG#JFTIP#S&
P(E(P3R(69X/<;35*K=YA3%:5V2N:8E1M?_51ON8/\O</H6WUJ.-S&:(&O95<"F$6
P8%"O%'W&4@;=*P=%ANQ4A8Z@;BC.B^)!<IP!"G5GECV4T\-S%LU9I&_)^,E(X6K"
P.X'$!NZ/Z5/)DV5E3)JEDF1,?M5V1R-1:?L5-LIR)76LX6EU?,.Y3W 8Q:M-4ZP,
P!L>"Y>WY^@(&YMQ@B&\>"O]:M[>TH"PQ=Z97" [UZ=FCL.!A8C *X** \C]O7Z ?
PQGVFR;#3Y, ."/\2:KJMDWFI^O:[]:,/[2Q6]P1;U"S=A$7_8WM@B1]HFP9;Y,UV
P\R!7-N]$")WG;J#YJN?;_$?R;*XI^NI4;:$3U2C)]Q-- XGZ'&A!NSY8T!6RXUD,
P)HIEW?^A=ACH&^!W/)BA.\Q;T>QRAO3U+ FEK.6/4?R\#N ^NF+@9S&!X6]*FJ,_
PLBS( ^BV.M7;W5L%UI(6N_.!IQ UV-0 [ITN:.D4$X.&C=-5_C%A5%<R)\$4UWE]
PACW+(N7MY?'.V]'&(,%#CUX<>I:G)&),FHL)>@+@0.--WJ\EBX-HLEFU/&#_9&\\
P7CN&I!TL,C3=X(H(2"YN^9^*+NO/6VWMIZ/9WI':KM4G*:"CJ2CE@]&#)EZI2"T4
P(.<*5#887>>NL_7HX:E7U4.U+)JAL-:$JTP/7W1;"G^LC>T40E9CD-LC4Q\RM?R^
P$>L%_6X3;C&LX'VI5U/S]3,'$20_+E4\):F6!H4(,#'8:\*0L WUR%W)C7R#PD^6
PBL'Y6CC>85D5.KP C.\%*.9GDY"39YY]H(-VS2&%V!G;LTZ<"@4&Q8]NLJ"E%VJS
P!5$R:%,8[R16[AIP]L  12^+%O3 >U09O-*%)K)+$*L]M9K,.H,86%>_P0H+2J-(
PCSE>)S6[_2MUUK,%L9Y"MP97[T\V9$WWQ*]V5[]K,)UP4QH%#A$R(%I4\JLHR7MF
PG@)O :_5<N;S=##5H,M:7"DG+4XV6Z_9<<%'Y]EKFIQ[\]1>\^&M;I2,"P^W7RI#
P(O_?$1=*@1!70.2F?GO]903GWB6#O9-E6WRS;3V4-\6T[?MBLPA<C-Z@><[PZQ^/
P2CU7K4_10J$#2J<_)DX*^?_F<3S%(,%?9KPR!=C$/%]"EU^C8.:NDG]*T$L'.-Z,
P<*D3&+37FL'I.[<]TI@#NJ+K6\2K6XL-W]5Y3LAT0#.[;Z1&3]=@S)NR>$076T87
PTB#H\2R2UJ"*Q47L0P6'_"6B=RT <TSCQ,;2<FX<W58L+O4KNMH<5'DEZ#N6,<%/
PDXQ8XB7"/U%GF55LW(]%$]%F+B,!1,$'%$L-+NOU\7W2T561]535!_R$D+2HJLX%
P1#BA;C+1RRYFX<3ON("C6@T4F5).E?%L >FW&.OQVOA0)F<V[A,OD:%[T-TR8";E
PS!V]!(:0GBAFG!5Y,U)R7P]23HZ.<5Q4HAZW[Z19Z4U H4+,;((#KRD@;Z' S8SZ
P<!ZJ\#$J$#;X4KA9X,#4EQK<; )8W%O\X9&(%%>>1TJN*RP]S> &%8ZHYJC'IBT=
P,CK][^:EJNN..95DY"Z XP?:/<LIZI"2;66)*VZ6.L,U#C86?4**ZF$$*?4B*95F
PR)970;?'JQE FT?3=!'@F,+RXF27*57!(: PRK>LJX9V&.33Z "-]UN\&(UJB',"
PCMC81U*@ YQ!.[A6(HA6KF.>LLR@Z(2SCQU'C^$;Y]Z:;_@WP$1"C.99[I1ENX\3
P<WG&-E^WJ, 'PL<C54)K+(?Z.O#M@CXA#T]\Z(-"5%?G@C_:=8UW+BC]W'V6LJP]
P0H ^M#8 "X$!AUGZ/ 2,?S!=^#\ZNVP-R3@PLIW?WQJ(5&.5*7IYO(QAB3#1LM-H
P=DOS$X9*IX/999,- S!M@*?-I9;%VK)R$[!:5>"N?QNZ;K_TU*#[S#"7O7;X\G5=
PEZN+NZSO"9>54K30E QI=)()!-(F*(PQ)<CW%JTMJU8%$&T0H37*JLM>O=(=>Q^@
P@?0,OKA=CXOT5AW2AI8N*YL%I<3E*'R_<87O]47HS)/4%"6Q(;;SY;&MZ/=QM_K1
P*'=[9+4 ]T%W+5TU@ RXI?G9YM6C\KI*]]1]P#Y=-7XGQY4'S;C<@>=,C92)_L*0
P:K3T7U^@]IIWMFFU$J=O1YKA;Z91O"J<%_= ;93^=Z2P>>$W_Z%L#\YL@6PGF,RJ
`endprotected128

////////////////////////////////////////////////////////////////////////////////////////////////////////////


`protected128
PW%6N-7SP_SO_TK,3>DL!DT-1M\7DG![]> 4:6,=?0!8.J\K]2J55I<2N=C=&Z<7U
P1HXYKU)%WM"&=D>44HQZ H7T5$?C]OT8_VY&]$08S%Z^N] GYI.=&9YAZQ:@>08 
P,ZHR A,T(3AUG#.]>\9U,S)H#T&@9QA^&Y@Z 9YY7:=Z>'6\$C_M^\1OKBBL*Z"R
PYW<M%/.3'R.<T+>TR"-V%!Q+9>+)X&;PKQZL"Z(R%7K[([_%D14YGN(N3OEQ%6=.
P::$AF^ EG*!+\TY2.M5\ V NMQ);/ A["K]-(IS"Y7V89'$B\#05YNN.<,&FBL:(
PV$?PR6+T85-&SV(^USJGF(EPC(>D*>74^I\).?ZX*++F1=^AMF^DX(@T)1B.V\H=
P[6H%C_'1JP$3HO3+3467^0Z=Z@C.=0NHTIT(U" N&]E#V#6P4IH_7?85=0)$1N#(
PZ(91DGN<ZYL6\S ]+:Y^P+[D<R8&JY@D020O;$E:%B'5.E[S[BXDZ4B)2.2=92V:
PTTNU6)LOAV7.PV#ZN23-;7,[WCU4\(EA3,S&CEOUP13"Y\6-.IN0[<*Y9T$\5C:N
P!3L/!62$68BG\04P=\]PZ&8R4/:!>P,]CVDOF/F7CQWO-175%B8J:A$2*;>GY)PB
P.Y.8A+_8P1'=X]FF2)V[P:XRH GZ"\RP WULFQ<?/6+0,+DQN:P$R7F]D326#SGN
P^/)+R>P'I,%C#3[$'_:J-TO_(8=5RV'EN&*+#.T_7;_:/'._WRYUZ,3SE"<U:NEN
P6AX0^D8A:Q*>//,KH;W-Z/)%1'!7I_NZ1KZ]1,I%:?X:(BUB]LGO(#ZCQD,5*G::
P5LX4N9-I:W+P:Z[=YF!/AL,C;-'27(CJ."(KV0A\/\!'2BG#;B?M7E*UE@*EGW21
P DM_MOX;G_?7!QI95#AR1Z1R^8. 00"< V7 6!A(?/LNQ]7/<C)O@>3L:E3#B34[
P\U'D%EG),\5S.-<?QF]>(:HW2XJ.49J&RM3$]3"C40T("+XE.4V0@K7D7!9O_E%.
PO"$BN:GJ-<_-; ]--AJ&Y,P.;CM-J26Z [2[8Z":/EPKBTUR^1U\OE@XM"=R^DPL
PF:K6JT6]%;,1:5FW+^T9^J_>I'UC0:MP<6"D)4"1WF' >'(!TSB.Y-T$K9!K'$:P
P5 MD;[=27OH60%;C,460]G.O)IS@=^H_.(K2TXE=L^;E&D&[13I@CIL,A=5Y;?<<
PRT3UXXQQ<A1S?*>EQ=ZFM---P10O@4-W"M:J/5'/+U__:6<V[ 2L-CS-!&F,9?W:
PQ]M4;G[$9&3J(TJ)N3EO&XZ?8%!5-H:O1H/GZT>7O$TB__@=4>G-+-,NA5$"C:$]
P51J'X+?Y:0I*54O6[32%)1U8VIG*9(@4/+M2D(.[_',PZ.Y"6(=D?*.@4=M!..V;
PU)=>Z>-'E="KD^*1!TK(1)4(!]!N4KJU_ OD]39VC@LW[QC[W)Z;(R1^<SGO$TDG
P)H]T1;>Z+(N^?.IPZW[[_8M'_>$1\=BD'L,M( (2<[(JUI!<5;Y'\(?UA8%,W;5R
PQ(1#%;PX:(.HRBOH7\GYQ,^,.JW(Z^(H7\;,%@4T@A=?&/=D'[VVPX]68IL*2K=G
P*U(G7,' %Z. (8)I]3)EQ&KC$8?/WX1\:I"WU,R1V#QTC:!_D<'%SUV"(D('YD^C
P[)2X]Q\:O8C41B816-C'9)-=F((55 .2P @,9R GO%W:"C%+=1_Z-:E!6T6L#Q'W
PY4/#.ZJ \&5TQH$?8OD**<XU0O3:=X*924<UN,][AS=;OL"HPH6H67W/LPVO#HBK
PJN]FQ*MC*R35#7:G8=UP$FV3OME3T7O+90*G^JQN^;%ED6^76DLQ*<T/1C6@;R?!
PXCD H-E>#W?VVF[&;5N!FK15D2%'8;(RR7'B:,]$W.K0H;<VI\#CU]U^RY9%$XZN
P'Q4G=NZ>*FY5+TX-G$C?"&22DGK,4#D?;'1#OJX%9,BP!JW(.HM>7&XJ%,KK:O)M
P9M(+ZN1=+&"+:E[&FJ1,LFRW^N X(Y#$;A\OBMIJ?2;Z0AO>L\TWBTA*SJ\NB=UL
PII/HBZ#J2]I*SUY>Y%P"J]R&S;>*<<:&B(YNJ9J']=*Y*8NMV# =D<2;(!V*Z^-F
PH/S_[?E]JP>X(1M/M#NT:R2,'"LTR#UFH WDLX\HB]?8%SC.M*WUL27,O@L E*\?
P@GL!NXA?'3]5Y%K<?>:Z !(6E"0IB/H"<_OXF2]*;14SZI\43095:M5*=K[Z,.<-
P*QCSKB:Q8-;Q:6EH,!+XRU<:#IAE?2ES%%U#M$21X#I\EKRF;33Y:[F#=V&F0E7W
P):P/3WXDBP:G"D."B-3D5PQYX* OJ//9[J')]].8LF6EF)]0!Y)JM:63[MI?,0SF
P;B__C2ZC]%TZ_J+1-KM!?2@KP6RA<^9\.<X5]G+U6A%.F@9Y&9(S0[81%%V3-*,\
PZ5AR)#%;;+V>WF\3PLI4M+$#+PW/#]5VT^0T.HMIMXT-BKK<U4C[2J_U%G8%BV"?
P;?7F9\3& BS/T)*W5V?_T.L@Q-)D2MRBKS,$>EM@P^#X1F+K<-1=0K /Z'%$5#,J
P^ O>3TL2R#4Q.K=SF]+GB.N^<D<BAG^V"5GUZB=1R\<LV6FM6$OV).Y1#=V(,[G#
P:VS=,<M %RAXIKE9H3@YS"7CZ1DJ3ZR%]2@QET O&4LW8+V7OZ+#D(*V(GVT[>KQ
P!OY%ZE9[E^76@?H>IS8VB&M*(^!'PO#]ZNB8/2UQ[52F[[C59&N*]IQ#E[,]_L,<
P'?_3*"B-_77.$HC$2YZ@%QX7C=)_3CRJU"D='UC2.$_,E>H"WF1HKWZ-S8?L[S)'
P(?7>!O34N+5,O7F I<TYXZ(ZE[K$_[@DBG<;_UIH9G[?\A;E)DE7\0%?W+9H_WJ0
P99YF75PN1%^I9![NI*B[JR/RU14)^5E\W*ZR#^>UGQ"4E<38)@JZAY<DB;9KHV!I
P1*$<;1R"RTW&S$Y69Z4/O$;^I+D$^%QZ'I?X9&V [JG0"9^?*40OT?S5TSSL+#6G
P^OQV$+I0Q4$;^NN9V#B#Z_]_UGG03D\(?FHZIAO:HRP:-4B&L0UMBIHAY+'\.=JN
P+\77?G-@643;*EWH@N8\0,YI'M804%[EUZVM%OZ(*F[@=GI\G&?:=M.VC#!%W/<A
P=H"YYW&;7]T7GFU05_>_LB2W8WB%".^^X73P3L<HQ0X0Q@R E@-6VJFG'1MP=VG]
P2B7S";'J@"#4WDR8LJ!7$LTG-]K8.UX_?!OLK#N="\N8B?XO4&W9FC_W;P*]60&<
PAX@$.$@SA6]<(:6$F^!'RN)JW>0+2[*!*+O H<=]F]/,)["J8XU9Y+61K-H-0ZM:
PBMB0L 7:$@HZ>=E5TJJ)%8_[Z$C 0X^*'\:Z2G;2 $'(W1)@W2#+@9VHO;]K=50B
P#$R:9W!8:[M\JZ %(P4#K1YE#4A:)DEO+')B%.YH3+HR30<55/-;@\N 4DO!L4X#
PFPOM;5/$;A[5]RZ\WI-2B^<!0K4HFDOQ%EZ$T@WSA ;Q\X> QOZ>^#RP*!]1L*'8
P)SPC)=(.3O0",6NOPON.YF5AYD5BO$)QIHFUY=SA>WA/W.]SQV#8:(^O;ITW#T0A
PF?0_>U#8"^;Y]\-\^:E\Q%QA]0>C=9Z+_6(,F/FKI*#VZ,LE$Q*!7UL>NG&8)3YU
PXDDSCA/%8[#A,I$86=Q6IL;DQEA4>.T7=QFISV/+Y+90N,!?GCK-XEK#QDR+:-S6
P=3'0Z'Q)[S%(D]/20R<]"U8O6I];PCC-34H"K;?%'Y49VWF.KWR? )Y,9&V.__RV
PR+Q;.^XK,0F?3PUK(\C8C&T[0V_0MW(]19CD;;BAK>^])$+XBL3-)T'F,WN4EKO;
P#DP!-_!O?EC']>VX"=@WGLG??#$.<VNE)S8V%<M9P#*>[ &.+I Z('>&PQ3SF!CS
PZO!V5+L]-S<ZR*:F'E9'$&E)W3&C(I55R]_)W8 4UR%%BY%=!7)2SE3=5?>[PSY,
POLD;_8R#YZ2G'^R_G<92;>3D=/$FQ7#M#<G&><V@W]XMA#^;@73R\-AW2M8?KH#O
P[:XPU%O<3YAI-0%[D2Z$L]U12?:.?=-;K_RPRL"1LQX9%S ,'/;C6T QO,*TW$"N
PW0RI>SJBMB4@BH1F'VXTGCXGB(VKTF4 QG.,"C;!1A5\9_UC[=,*+67RT^9U0G7_
PAN!HF(R;$-_/:)"OQ5/WXR4D3> @E3F4.T9&HD* V(C%M\**RR?R_4W+G(WHO$X"
P9CW]ZAXDB5J.C401@4'A8F308ZB<-I0[PH_D6N%.\O.IQ;*E+H;#.?H.346US4*.
`endprotected128

////////////////////////////////////////////////////////////////////////////////////////////////////////////


`protected128
PW%6N-7SP_SO_TK,3>DL!DT-1M\7DG![]> 4:6,=?0!8.J\K]2J55I<2N=C=&Z<7U
P1HXYKU)%WM"&=D>44HQZ L^1*;-_5<27\?IN07254^>:(YO*WMC%8QSN#JD-_).R
P,IA9V19?C^1[;_B9C?V%R\SM;OU09JZ3'K,J??B^;YFIJ&B'7'$Q5Y/7NHM*L7-S
PDPZ\8+=F&&[KC\TNE!?6ZO'^45-YTQC"%BL%[R,<&&;V=B1B4X 4+9_D7_R%F#O5
P\ ?00Y^.I?M0P5J!BJ!"_@!O D=_5OC[965;Q0?'JUKC1.N*F\(QXQ%+NC8>C'O*
P&"'5L: C"7TAH^F\CYNS#!7A] 7;Y"=_D)R'20JL1[TPN7O#^3ZB+@FTT4ME[BX8
PJ4O>2#(U51[G8X#L]JKL+-HAYK:7^0\WP0$W3D@[OS,/ 8.QFI:(]$7>O/G&#.B"
P+/@@8^_-HU_O;MHB?UBNJ#=)9,0.=(C^3G(!Y9Y;69L;UR!I5LDM8#S2B%=<3M/O
PH=EL'_8E=5^?UO@,1>NNOB,>'CC/W;]"#W^D-ARXX&%O<1'H=>4#SPC\S8ZV-8BW
P0^=1FH/E%+S6@S-$VZ)R.A=UG08R7775C68D[V_.Q15<X)S+5WZ,Z\+I*1K DL("
PTA]6='[?LS3"7?06<)#VATWN^;?LK3GDFO4AIPH9[SVO?#4Q!U61:8KB)L*!J *9
PP<N'PLLW.I:^CA\[(A:2,EV9DS?.$ZXT]MW=R:'/FUH0='O?PAM H&X=)CC7SQ>"
P3CHC;O/9Y')G1CUP8$</H?(:'7RNV1*JL#^$94,8DPH6AN, B%Q#;^7IG-OY4.$T
PN))SBSX[HYV[$UD&\$J%%=P=&<H$P< $U"@HVD'KX@%O_\QM=)1:=D@0LW%OK0;L
P#<&K^^B42$<CGBT3PXJTJ=#+[O^5E;/EF3)ZO"X6Y*2CAY]$CQ!J=)K-DI&]Z-[I
P2'&^KC27*)IO2JA;F\EYIKX*.V_%6<-EHF.]>WLILY-J>' 1R$93%]&**SZ^M$)Y
P\3:%5$.]\94]F0$1M\9O_XM)O(+3K#"YD:Z6#4\5,'@\^'L\7S<_.@S'U7ZSG1OI
PZ5G'U.09IN[:Z@23QCTI(5-5R<=RZ2"5/"7$K3P2C>\X+F3??6-0?2X@JL,Q??.N
`endprotected128

////////////////////////////////////////////////////////////////////////////////////////////////////////////


`protected128
PW%6N-7SP_SO_TK,3>DL!DT-1M\7DG![]> 4:6,=?0!8.J\K]2J55I<2N=C=&Z<7U
P1HXYKU)%WM"&=D>44HQZ A=7/S=:]6_U@,_UP\X!!G#L =LX?#WOP7=^AI^K,W:G
P1'BU1++[6*XK\0E0D"_G49@JH,4P87EI>UR^=NW++%_2QI.9#MMB+OWN"P=4XOB=
P+LJCO:PV$W<W[-@ L7D3."C3&M,EQJB(0[#^1(OK!BO,$ME'SVY\75I>TU!$!_KJ
P0\Q$*F_P,U5H8UYZTN?Q;ZCG)$>BR:O_$@9_VCL8K9#QFGU1_!DX[ N7SVGW*?84
P,:#!2>&2^;BHY<PH)]QS(M^0>1210KROM=7J.;;'W3\5_8"@4&AVC)J"U[!T%9W[
P-\=VE""#RK1&^"\:+J$)>.55+]4O3VG>^^19&+(,[Y"@=NX9N!EF/X(TH8PEZRVP
P,0WB<W4C- :/&:MR(H:!BI=RB-I_\Y!@V,'VC=KBALMPM?U 1FAG'QJ<DE'*Y^53
P[!?/X?.=N)]2"H"!/LVUB=L/>'4<D+$:MO7GEDOP83F6UQXE[,;,$ 1_F9<34\ E
PR(F2*=.3R3)RUQ!.$ >/Y\3U51-,9*9*;P;AHIRO%>7J3@2$D#G: D4WF>*8F<(!
P&33@VR?*X.Q%+181+/AUWJ!@.W:E,03UD)5\61$='1-OX'(!?F;/W<WOOBG=(^]S
P*#W_&VPR;!<V2R/%)'Q7TLX)N-,CT?I/$M*#DWZ7YY&;\/A>%*X&BJ!@I*^PI!V;
P*<D1RVJS0D;RHH_ROSIKM(9%J.C8D=F>E2ML 5?1+>W%:/TCUG:9(I5WC"9"(T[9
P V^.%[V"^HODI7)2Q'7004KA[^H[L40U#2^WM-D%9/?SUKS"6JSH4)5^'ANQ6M"G
PP"M,Z!T)?QAQAK##\/;;CR-7<#!>%'CY&6$5^BHXT!JNR06/B_O@)[KD2]G$5!76
P\>S?/E#0NBP)"NU_8O7];NFT) C!#E=4'U,I'OH'[OMQH6&\(=)X;Z!0)A0BA\+2
P_>&[.>K"(?DP__;FGI(RUX?@='B C,8.(G<UC'H#/97K42A7RU"A_9$-\6A.-=\*
PDNDNY9!PQ(1SFS:R3*G+0FP)41Y8O@1O=0H46.EA1UQH/9=)7^9H;,;I=?Y8*15,
P+&H^#.?5))SY!HXJETE#^2=J$:5'<=+0G(:L J(UID,;L[=4H8._&2M "%0+@-9Y
P  :;QR;T_KM&4XJ$2D\UXUEQ@%4N#,UA3%;!QED/W1BKJQ(IK/D'-;DZ!T!R32H7
P!19MD^+D1U>>>2T(%? X-&\GA3+_A3"):AM5GHN 73-[OF+"1YE?RT<AO<>,K?J@
P[U-^\M:R*D(%%]*[0*?R)M-I@)>>/GGM#MRG)Q>JNWS >S_[@_,8@P/8#P^C?9'!
P2]%;3J1R86'8;Y-V&EPGX68 GH/\]^4G2\@@Z8\6Y*JO*Y .Z%RR_BNQ>FFY+1?&
PS)F<5C;!C?Y/EOG@P@\:O-*;J)R\DLV6SG7;>7>#E*0ZGW3%16!IT6:%I "L(%*]
PE89O2]Z40@Z;Q-N4 W$@#1+)AT:' HUN:S[$FMEJB/6RAV_%E3U1E/(+NB21$QB[
PEP9$!BT'Q]@$P:C6J>$KJ&%R=?>\V:)\YY\>>R;BV 2BIS/>K@86@#VF_?9?(12U
P3[CVPSNJ"_=.#W.M)ZF"'*W-6*P4 9+\MJKUF],5))GVE'1_8MQ^>&%+\!X&'4Z]
PY>"3N?=76OJ3>2/><T3R0"/KDF=29?BOO!A*JVSP#9'-_W-!V2SD#$*ZS\@[:-P,
PJIZQJ/SVB.>E%?V\DC4TK@2]Z%$@\Q)FU*-!PNP3X%5K[\#+T9?YS?X#J+K0V+$(
P[7;(M D7C*H2*5 *G"^AYX9O1(4BUI"7RPI9-9D!+## #GK+KPQ?-LW1=%#%/]J^
P!7&-JWOW=[0U:MFJT"0'CWL\R2HLV[XFP.P-Q-WTU6A\N21RWCSWX:WI=P4USXK'
P<<9 @EH1 QG)!3HR6 2U.NW(4;?S=&.<W]6?<L75G*K6L#+6Z-D>)"N20:GQ7(8!
P**Q(75K5[4];Q+.H1=A\!$"D_/B$P](..O6GGAVZS:@R+!L3& Q0DD)7_?OEKL-=
P1J*3*D?RVE&ZD&M63SC]27K3M__!8]EA))Q7\YGIBG'.*&8Y89<*"5NNZGK\N?#V
P^]FCG6U>TR5:KA#O"IRNH*V0-F\O;K$N!<H4ATB^_ #:*8<(O8/\\!3C"42Q_K4W
P83666_7$X(#FQZ8V_$Z^P-7!NW#&VQSBA*D*C*&_A(.UW+7+C5\/-#8B+YBE>DQ$
P1/U03M9](N5"7,W@A]%O45ELFY7_5!$'XJ5C=I</ R=@S5L+7'387D:IS\TL7-IT
PX8Y*:Z6V]W:C->%4Q^YEWA1A<L=UR.W$[GQA,X0!#?U#9U"L#@5===P0O35+V[! 
P#;FAX2.QP!9?7M(\DE#*<S0$RE^<US/MYSQ:VE87?=N.(RKJ[GL0X3(^RKJJ5R2*
PH8Q6)?D;NPV%OIWE-N:0\=Y]"N5N508(29IE@3&G_KCE-VY Y0Q[BP4QL8?3CUR#
P$2IC8PF?AL==L6Q<>6A/4O01@"]MT-,?&$M.1I:&^$!][$,Q#:Y%>4:7WZH^!.80
PGK):HJBSCZ/86KUO*-:!PT;P[ /TG7W4TEB]D_R=2?H6C,WE(<F-97@_OK1-5(1M
PSS5S)\+Y,29GK2L4SX.)%.#BV;/']?/AVKL,@J'4YF2E6FU3X59R1Q(RNN,>)4#'
P@.VZ!9&P*E A=4"J7JLL9*<[4Z!H8ADWIK6N.M XL93+_STH]U6A#)W?ZG0O@),\
PQ<<\.U*4%0X"I\-Z"# #2S+'D[3VZ.HW*=]%</,G$9"YGKRO*LE(A]HX(J1_.:\L
P>RI66??+(>!L42VXICU19$VV?Z"X-^PUI"<43%%@!(&4M7'(FHG+:97 G?XV3$+Q
P94Q'I0D==U4;*3LDFY7ID<$![KD>P3=S4&(XR&F>2D>^0L[E>ZX>L>ED5HZLT3TL
P@XIH7B]3/Y8.88+@13'7WR8=+NX);,7*T0&Z *#_>+8RG$=T;R2>)V0XHQ7B*.HI
P^\>!@62904N+9BT;<,2HU^<\M3AS>=Y"EU/4P'_UWQ#W917:\N)7J@^>?  -ZI8>
PRIALN-&4=WA=!P/FPG@1P'YS?Z*F'KI\)=1K<X<:99.>%8"WE.?M*"$'_%U&*3TB
PFV-58<TQN&6K%/YX<9K2K!8A84[ODC[W;LT(6+?+<J^SM1>@*-(HHK2>O?$R]*?;
P7'8_U\;W0IH3)B?ES\7DD9G@5[MJ":SR(,#$HEJE5OOG.F+6@X:P0+RIKI&[FX;;
P_ L=<B'@=>O"'*?NXN75;@H5;MT#]0-98*V;*?#K+;*H%TQ],^8,QEMO0C+EF;_%
P89?)SQKZDTKJ!7/@2E-;Z4W5H\+HX2R$=ZY1RT[3AO0?$%DI&V Y:3I];?NZQD&0
P.!OSB=:#A(Z5ETN#2=(Z*X-;_8Y>DW0Y6)0P/RF#IH?1$8M4YY\C<ACABDMD@9_A
PM^_ *$[5,P,7YL#6[>>L6?+(/B!2_]U)A#UD:>\&;-=1[.<!KV'G)++K:2245'8Y
PBAC,3-$FW0IH*%9(EDD_ N"&ZLV_[!\Z\FG%.F+UKY^M:E[=XGZ$O3%6GF."Z-#8
PNVX]\KR!TPP)6QV"@K@JM16TG"5$ 2%E6LF:&>)K02FCD2K.P>@@VN!F9\3VFGP-
PP^HX%)J;FP8@P!&3 DAH\M2!#Y$B=GEB>\ 51\8I1U;$*]J%J?==6/W3W&J<]J.-
P()(,V\Q2.W=W:?#HHPJ4S3MK*5>6.KP+%]NRO6?H;-H:Z/_?06 #!&WH\%@_$D;(
PXFX64HK'9>3*:V 2Q*J52=X?>I_Q4;9%7;@O-M-0R6>^O/;O)?$$V$*(,[:K=YHN
P9CK<(=.'D)CL,8TV I6N-[5\$&2ORPD/MKKI.M&L4U2-TB(M"!C%M=?J"4T&C[*:
PYAEN?>QG[X G;;Z346H)6,;OJ#<%&G\@NV_95\'848E+0^8-]!:3*P0WKBZH.8EC
PTDW94M?9N86$!AQ2SE!E%"^/BUC?PGAPK>I,_\<\)ST.G(<+1JGI=+RU+39?I3J;
PF#[J*@3R;4'8Y:$',?D#N::IT*<55%T4,%3*X5+4?_!D;+%$3C_5K>"!"&-@$I"#
PO?U>#PKK"*MICWPK1[!1I-K18&'3TI:%3^!= J8.LN\@D;R_*V4%@U9E5K9#67AO
PW:S"AVP-YN+8#.[LNB\%Q'>:1WC/A-PG,JLYHZR?97&\ 4U=Y.%XYE&N:E@&8N)L
P\U](^% OA,6LZA?*8BT:576V81L#HQHS1ANP^Q?=_=) )Q*4N?[@P@1*?W@<YR3)
P>%1961Z+8VT9?=_D:T_0ENN:D^JH6S._X)&7@X;F@-$F:0YW[HP];>?9[L,=^N0E
P[ ^ZV 3OKM*K#F/8V9K?I%YCD@G)\Y%+\"A@L+IARD_!G=G-9C\R Z.1*Z#N?0]!
PU<CT1]=3@J$&39,HA0WJ&'6$5S=:/D] >.<P.EK'G/H,G"WZ;/T0F48J ^"!1)0A
P^,\??SP-/4YIIK &Z!JRK07=*7!@:Z%PV:T?#&A*'/] ]7%Z#\7,1$45G&<)*&PG
PP:]E)4++(<7/+^.PG'-'N:LVI_0K^*^*YN%7JV:/U'??+?& @@P7C45_*BN!BI][
PBE\"X: "4N,4UO]J ! T>&E:0[L:'3[40HS!23*3B8,2Y$%UXQYUN?RQ:S%3V*Y.
P+T<9S)T"QH G^@1+_#=UK1CX;];R+&0,B#1%U/'LG=#_1\N=*P:6F3S&12"5T*MQ
PT_?(N9)500?QZR=VUN$W,$Z"ZY%W(6U<Q3M!S919EU%[0!L#OQ6YK$E-($:@;UW_
P-8.)X]!Z_I<;N'82ON3[NPILFIV'R8FA444ZWJ2NP'K+V8#_H/%RS>U=;+MS-=.[
PP+>\K0!R!%URNY:45!O65)]Q/R,O@_,*5P#9=J+RDCP>OH:BF94.OF8T#4.DX%1Z
P[1L_V&4JN@@>J8'X@R8MK!!1S$RRRJ6*=XJ^D9(CM(!$#)KL$1E,<HK+S3_F&O=D
P*VMGS_( -?_C!%8/I@ A92-1O1W0>_+RZP?E .V> ':K?Y*-]*"*(H4JNK>^HSFA
PU)(H&6K;KO-R&S)38ISJYEC';B7>,Z6HS@]BR;7SE&PC^<5+5.A AH;3(N0E\&RN
P=Q;1.*XRY'GO:,]C;DT%#3K('!-S$'0"//&7I+N3J,-*"<2#7C]ZI_5-N-_MX)D<
PK*9+_1#8?9)1 WN$#\N]63NK?G(8/!RZ%0>5\<*SW0Y>G.AV'V$BPFK+6F_3?^5O
PYP0I? =#  &(%W,6DYS]?UNT/38*MSS[+=C/Q)]._<4]P0?%+_6>EP^.X1ZK$ECM
PFIW359P+&7<&G(= I8FMR4-_O ^I6BM1SQOOV-,T2AK;.(82MG$79TCZ2)D(?.+R
P(BWC)K^/^;#;]244'Y(ZX7H/7)DZ*I]NB1=:CY+\]!\]1]T>]-S_ >8PD"L-@O'>
P>1C9.JS378<?F=#7YZX1H)5I4]&T?.[*<Q@9#G,+#VH.Z4/B*QGS4W:0SJF/EJ%:
P5DI4#^?R/(*.<1BD[Y?0=2>!HJW>8"%MHD\WIL+X91]='HYJ32\ 2MI?N@>T+X)X
P2FYX(1T+^50EW8KA>--UTGRS1BE#V2<.LI %+Y;%[)V0W#'S<R<,Q#[.>IT:/L$!
PVH_L0T/ E"'64P4X' ]/X71NMVX(4W_8.WP@T:0:_VT[V;@.'EQ\L"5+FG>@'T?X
P<,W1G:,D/IC"(&EPJ%$3*3BT8M4\-+-I0=J 6)RR/9W;8$>47I @K@C*+ ,^$LU#
P!=%8=  D$#Z><<6W JFX\"B;Y 56J&;XD&,D!QSG;?UG/G7N%\D2/8W/9?SVNG)D
PDN T+60!MYJ)SRM6[6]+SOD>0>8D5))L">NL2(/NI_I1]A()>O3_B[9KAI%1SYF,
PY(#T%)19;M^@XU89D0U#T_*D4ZY(XY%:F9>E)OA+,^1)9)L3KAP8&XZM+'(+A.PV
PN>FAITE[U"%MT>[ R,3&XD5^A]$!' ^A,WQ\:J/%>30T/B1Q*HFB^8=XY-J#U>EB
P.[)-)YCO2=:F=)"&4DT?DF5!=(ORO.0XS=60ZLB4]^3SJ/,\BJBAP]Z=5>;]]YG6
`endprotected128

////////////////////////////////////////////////////////////////////////////////////////////////////////////


`protected128
PW%6N-7SP_SO_TK,3>DL!DT-1M\7DG![]> 4:6,=?0!8.J\K]2J55I<2N=C=&Z<7U
P1HXYKU)%WM"&=D>44HQZ A=7/S=:]6_U@,_UP\X!!G#L =LX?#WOP7=^AI^K,W:G
P S=J-\@R)9XYIU4]13R@]/A:H\DY52,;\DL>@ :6$=2JX*#%L7FHL@\D/[A0B7S:
PY2L)6(_]Y+H*1SRN6P@H D[8N:RGA8^&_!A\D9*R>42O%0P+:A1:!#JUM$XBFZWG
P?<+20<S+L7<(D6Y(7SVCTEJQZ"J)%+?F$K1"7ZHCHV]/;G;BKA@YY3/1N?"[?,JX
PG3MK9I5 6&R>&Q8P:I]W.?=Y1)#"D\\ZD;JOTNK@^;C;7+]\8D8P4:PVF8ID  XU
P!$JR8G2K;C5-]5$TH=29S2 2+]EP8S 4:M@UP(;8_0#$(*V(@[3MAGDJ9M3! V?K
P,YT<X<\O"1!#X(.>Q58H\ 8^$W'\FOG)]%1MYW-P.( 2?*&T1PQ;M3EN".S7'6=Q
P$8B/$'$_/)I(NG,\7W,T"'!"$>530$O>[Y.J@ ;B&+A<]GV]_Z'>UAA8] P%N'QB
P*I2S79YWP#DE<" A!S+%XH/^W68C<UODNVN<VP5A<KW0*#Y15S]7[?T]1):5,K :
PH-JO[/;">2G-TV.()H1DHRWX_!=4AH%?#^J*A!<T!/+N9BLL4C85KTRC/;J4@L$=
P%M\]9WK^H7+CBM1R=.3E"52<QS-1Q^1A5Q_3PDYM-B!&+HV!2IPJ2/4/5T=3//!Q
P3Q1!CVSC6?S>Y-)'LK)0IY./0)_3BU?L6-LP\S7S4_:9%O.B3'U%1NN83]XR+S'@
P/)/VE?14B%]KA*4!!?]WG7 WK!;8K/74;T$Q^[P71=T0G5^%6?244'GMKBN6L4WY
P_EE]-+C@MW'ZU(8>6DH/$G+>ZJ^N/,)E.\Z28JNL?;$[J=>/K.0=).;$+[DP/BOB
P)"%"<HSC'"<+;7^A*YPB&/JMZOH-"G%QV;+->3>M(&5N:,6+F)HE;8;I;L4K5R9U
PC,XX+#)%)_+37\,54=11 5RFP"6KS9Q,@@T$"G3YHJ<@,SZN+_S2-0CY:+CX5>'$
PQPZ6WJB>^_SZZ3$DZ_K X"M&KAL3P.#H%P ALO.CJ+>"^6?TK-O??H%PT+05N;%S
P\)EI!!9^ 19VQ"@<<BJ"H\.Y]/9ZY;O #XZHY)S*GXJG4Z?X4D?'0-9N8)(G1GBZ
PXW%O/5W@BF(,ZZ<9)=(*C+=-MSORHAX>)78%1V5V0D #IZ22%2@9H3CF](Z&!",X
P3NEJ?,7,TT 5Y]"*3]E+!@4&FF!_AX>/1I&4(62$C!.D3FTY(2XAKHJHAOR=$VW!
PC5W(_VKNI)DM\8)X@?W-@WG D-@D*W1/Q>_^X1(;'!B"_W<P=%8^]<4F&0]\,H2@
PHH*[GK'97%[PA'F6=(#IS]Q)V*O8W^48P6Q(S[59@^ZEH9#J+(4XWG3U]])01:A;
P]V]6&0!L"/WO !;]:^3]#',%XMV84O F=&$EKP^E_"ONXPS88"L]GLK1.VL"VC'1
P*ZW !"-'1UK%K04>Z,&_)LH L4Z">3.59F<1>6@BZ(#I*R" @Q%?Z2E;E55>[&0Z
P9''=$M<*RW=ML+7?79="_.=*)F&;@*[OW6!G_4BFO0HFL^@X8]%?A?B#E;@FAO*Y
P''KR^/R(;Q@!TRA(@ BZF9X*M^H8#P;[U3B0..$WFC(#4B@N94.@PE/-&PG^D5W2
P;&>TJR8*"X5#+'SXFFG'=,0WO!&KI!D9.?:V5(L#<',?0[4R?B60![H'6+ 2H[PC
P3B"&%';%0)>/"'_$T 0"JG.:?MYX[KZE33X.2%1NMYF'+V@J=%5:(RO*2W*%\9I&
P$_.!D3.'8F'(85:D!_(+*\"IW-35X<X#7 W8^U/<2T'H@07'9TX+/NES'. JL29M
P&SY=S@T$*#% [:-:*8=8J.%@=Z:D33<@H: WH.0X\<VSB01-SHZ5H)U*>7R@@[8.
PZKP5V&L9Q@J9+;<)I8L(CPB_("EJSMMDO(Z;=UP] 9QN+F<]M2"9\FU!T 1M[H0C
P75[^O)V!V)O)KH"..?EDCR]0)EU5=9QVC:0UP$$V\[EC1F055;;<# A[2=EHF9MG
`endprotected128

////////////////////////////////////////////////////////////////////////////////////////////////////////////


`protected128
PW%6N-7SP_SO_TK,3>DL!DT-1M\7DG![]> 4:6,=?0!8.J\K]2J55I<2N=C=&Z<7U
PF>S#:'*-QNR%<^)6=#&>ZJ&AFN_C&J5A/56B++R;YT#1@(X=2&7#SN(>!-CO_JK&
P\GCII$(MEP]2@M0J#!4()KD1Z ";,,MMH1KJRO]1FBC)8QFNZISMY4$6BA]DKS7*
PEM:6T#,9-@ZQ#^N(=_^@# [=\&N0,Z.(!"?^J 9,6JH)$XQIC'W(5G/PV_&8/7HF
P=C0]7X!4AXK5OY];R$'!YTI+7R,T%L8S,D&I2?6\''H#L@_0F33Z&L<L,F%1UNTT
PKDR+;< +LJR47)K#=N!/\Q[5?O+@R%9%DM;%QN.D\O+(>Z_YN(4</ V2M&#9\(Z(
P0DZIHR_LC7ET]1R,8+*.P:H$T&![IR'IHY@*@^J+>?-J+VA&3']PAF7=X =9,X1A
PJ'4Z)7L6:VX?9W0HVQ3D2-OMWF9EO3^4GJU!/V-$%9A0S-?* 7A$Y(1!YW??.*%#
P A'?P$F/,BWS>"Y"=7%U9-93?0@#3K+R7W]'%9S! 4:PVJ9LH':@/83%W'B1GRQB
PY.T>U)N3(#1/U\HU6--@VD]F9)7V5.O:<%N"2%'%2 QSH /N"N0@0)S$WICN(;Y/
PBC2^5-(R\J77*H!&1<+6MQ"'3XTA=K^V%@T]LQ/:$=&6B+7R92=<"6,[$]S:;H7<
P^HQ3+9E$]0@:[^9,+($;#+!P2+\OIUDX\ETKUH/W'!@IZQJ"H3NJ:V0[903*S, S
PCA+]KDVN*K$1J#6OCTV?F(+YR_QGTS(VO(!O;5(/>^C&2S(J@B@9Y:XZX("1&Z0\
PU/E9CJ0"#&E?PP73FF!K(9O\EE]HFJWVH]+C5,@#VVL+U-$A^*9?@^J2K: E.)$)
P1O7OGGY0JN6,/(?JA8; \ZP/J3 VYJN.'8(J;X>HM\WP4?=.:>$M7 >Z5<1!<HYF
PTB[#P;>8+&&3%FE4A 45V9?B,NP7FD0^KVD2-1E[?MLW48B1V[LDX42CG.]5]3M%
P!P/]D-0TNC.8TB$12GDLCPC49GV76]L#0/SA-]@#RC '$L@%("2'1Z)J^EAV_BAE
P-Y7Q)N+&F@W*MFM^\O/(J^;-/S/"61Z!=!\Z6BSF!9:E^7 W2F>I^_1D*:[=BA+N
PIF27],)\1-_@JP=)0T63T.@IU'DDF-96V9W,PZF[]7VCB'F]_!>1'NP@'B UZQ2=
P)+EO[S&.M.(?Y#I9($.T[:41CU6 GKF(.;P @T*97:'#[0S1_\)8,9#S-U^>.R@0
PQ"(TO1A,*P^HV[F1!GH-K67C[FWC&[.F/W;W7IV?'TU4QRE3Q(&_*.<5%C8=+.*7
P?4T_.)SDGJ&F3J20,NYMP[G[&*@G,E8E$56C.Y*]6T?-VB=H0T16QF+7(U E/F:U
PR3 Q?=QUJ#QB8>R>J;W-$CYOH6*%_+I@I7[,,6?7T82<EQ:L! ^RHVY;TWB+HXID
P8(!6ZK#_H1Y8;GT,Z]B#Y+A.;6PA:8CY),\&_&SCY1SDQ^^'(="/XYKV:[OLVT1H
P*$TS5<AV"4X?8=[F*P"V5<9=)?1JQ]O8_>ZN<?WVIH>6F;V9-+&(1NONP_1V.)2:
P8\:1!N4$:6XEVQ<386$#4T&KBD?"VN,15W$>'VL"</0ND4MH1?O6^8Q]/&>7H 6'
PC37/@^AOVQP_!9!^&)VRR!!1H=&KQ OG^UM/T2Y.IWBKH&!8J2<G1RNG=%N)H;D*
PWBP()ZG1Y4)- VPDRJ^/UK *P =3K45Z;/-"7T8?#YX8JV.3?]-_WL63()G4;BV(
PO>=T5T"K"L/% ?:1.&&B$AMI;:6P/QJ"A<'V:J_6G*)R<P;%-L<NVQ33W&#HG0YG
PEW>/BP/O>]D5,2^PY-0MFEZCZ'A \/1F/G7F286V5SW@N)#WO^$WF*PX: *66A>$
PS*9LF,B682^XYNQP?PH!'*%+05'F2K;:'QJ"F AF3J]0]VM#5I"K3@W,YW4%!8OI
P9U/HW/&\ 9B=C-A +GV)F0'Q()RDZ&.NF7>@<'!&-WH0K;1;6%,WGNAZEC^%^5E_
P+%#NH5A@$0?2_3>)11$9/5#^?I,RK@XB.2;]Y.(EQ@6=OB0R'_M#[B*%7T@T:?/Q
PS\U#NTHDK!0;_1Q+9!;2&$4J5]F!6(C%([PN)*D#FZ4'%B S<C[6#)<P#E0L&R"R
P_9*_5/IKA-W(<^$FWN&:K<X5SB;P6(^N\3]6;)X/ X\K66S?P@4: FL7 DN3#L?0
P+ 6<][<O#!]5IC/PC!UMO-P,-F".E_)WT3+QA$LI#8*SZK##9;,  +O'[4K2+D06
P@>-]?BBRXGZ6U:8%LPV: 2B4=W'L@!YS9"+B/MCE+3/B'XDL/7PT#MH\4MZV4W*7
PA I8%UCH<:2!9==>[]VA;=$%%'735X$^^O/A.%VF^8$WI48O(.*<]NO2S++5"'/0
P.#P50(G%K77A<28VOLFPZY.4N]8:47RV1A]O*UFA%><P=O&KH[BL3+$%5@AT&R'!
P9AOFU8/%:I3:LUK)^8Q&[%0HJ,+$N9]U Y/%")10FVB2OXUC4>["+O]^-3K!\?27
P5E=-=$7==R"W@#TV'4F-.'S=JDW771)#]K??>C2:^7AAW"F!SK0FM GJ+*D[_:?V
PZ_9\OBO#EK[J6_%'K*'W4KX8/@X9P305<7QKOP\&6G*BUE\&8S>N@"]3.$8!'\K#
PPD-KZ$**6$?9$,L>^:4O)'[_4LDO?F>LMK>A3YOOY9[^'*-.<O)1O'7-%"DSMK8@
P^03TJW50KE0]SI]-91O_*YQALA@9QSI0] :PE=(X+[UL!Q2S5]FWGT3-@.B!"U2-
P_WX^>RLTC2DM@_JPC1#V\:C!W7%D.3^"L.FHHI7JH$SW/FM(PTA\3,>=/ZJ9!@:J
P&<MSMBM!SN5/FD'8.JE<$ 9H(V,"A'I<2N 8()$H5[F$6G[B<VN86S+@J+HHIK,&
P?"ZK2R??RMVX5%C#/V=%U?)Y+PSIQ(3GO4.$R($)%4_Y8_,SGL3ZB.'-(/+$O>3B
P 5I//3>FJR*7N9W^$%)%[PS<@DH^F]R(MRR@'E"<"*DL<4"][3[:"@7OX=ZA;KTR
PN5J#[<_ A-W\4U8#FM#1G-JVN2GSHJVT\H8=E&OT"62\OL7O\0;.#)G?_&D)OUW:
PQHFWC\HT?J3VZCD4[.A]SZ7QA$3105PC%/.UM!!?4G+"\$HJ7=<.1.)2U4V!@@XR
P0IZ3,.%]&F_"FYGAOIWQO';C_%BV&G#/?@D(R!H13EV&W7>3;!4PQ9%\*I+]2#2 
P;:XF)4 )LP_3O![AU7C-$$WW2U8[=PEX)X?'$^N%?1PKJ7$CA]3!-)"7.I.<2%U3
P(E3&XRC3ZB["? E8@\#<]W: =\PRK8=(D8HDO1-X29SZS?#(+I'+5^B,Y?/?((X#
P1IVF5 9QK\,PI"IC,H3*AI00(]($U&?3);5GD#DXFTA/.SJQ1Y*^S"1J&.7,#Q.#
PU\[.+17G6[1=TT3:/%>:/Z@,N+"Z/Q3Q.IE%&#,\-?)M:_>QB.@BW93C9M--%CF"
P$5OFV>*2CFX?C\ K_]E&$<^.[ZZ DC/)]ZSF-!KLY <&4WX @-%X(^QE5^WF)36^
PR>51_D[\V,<_,6T_3&@#J[ (K5,-$EH+UT=:S64%P2:_E!(EV]&_=XA-!1'#]F6.
P%0-@]7&W->H=7!I8T'@\%@B=F93N6*P06\W$+H ![/$3L5^:HQIO2(UW\:9F$*@8
P=>B/JL!$HT !K&<YWT\/%O/&U9IM.."YW D35ULU<"T3>O!_+<TMW4&@;Y=C&J:G
PZ$6%=\JC5S0\B34,C@93R]Q+.!?7$3F/XJL?$G+_,>(V0N(_B_N^A2VIUINEO!5!
PD 69SYG:=!]\@4_1 @AG?/_KK^>\#TCP@W@S635-"P+ ;:7-9]6AU!2HMV</:6_J
PA<A$IVB^#'9&2ZQ#EWABT;8IIGL<J/B\^'V_0Q< ]]B7L@#A'#%?ASCDVF,,)Y*"
PUN3[Z3>]ITKMP:NM:7$&L#V4EQ(QA[/F8 !'^#:Z1N??U$J(4^/7=\OD7^,3HY#F
P_:Z:-<F$3]]-J9)EBV/K'*T!!",MW.I5D26+C.9_?^BJU&+/L1J0"R]2'3RW'ZV%
P@TFY"*TNA,DD]G'FD"$$&<FU\0N"(B._ \'B2DDN\TZ#JQ&T=JLDSBO,J]_F9S-Y
P_K26+1DL0Q/9GEBJJFNJ0/WU],FW9A<%13"G=@8Q\Q*].[8O%<%\T:8Y0K6_='G+
PY/:E*BGB)%ZBP9PB2>:6 3QZV#+7[0K2!'F%XP-'Y [?2QP(+0W4O08 MC)$>7#>
P>(;"Q_F/DOI/=A3RO,-M7S)@:=\\W=LIEMWX6D+A6IL>"TI1^+4C3ZY7+DML??K.
P@]3Z*3-(HM ^B7^6JQ_.5^Z;7N4F9/3-XWE7(7RIB3_'&A>2B)RI3S@JDD 'P9,8
P1V8Q&RS.PK./Z5X,O,7*/?@,*A0VO.:;^>#A/SO+8UX;W(QKBPFM'#IFB.^:B,.Q
P04S(\'0E:W\#Q<$ :XP[%L3SU%)MAUR0?IS=NC/J/.;XP+R4+"%\]L&JGO*015W9
P8S-7M?L9H>F-DHF-S"(T3X/W>QC+$XG:>S,S%HIH?NKM/11E) JVM+URJ"VR^_F\
P;;W]$@W-!L.DV^UU4,5MO#JD"O8"NH+T#VQJK@@=WQS7ET(>,3V5O]+GE$ZX+^/6
P(:'N0*GF6-D6$$%9#(9FRIFF5?;M=@+QR#]LS4ISYRE1K"8(67_&M%](HWE,%'F4
P0,:*5L(8*;FVIGL%.)_K1FV5-81DIL>2]XX1E.;BIV!JPEIC%2<\VU&I 22J-)4.
P5,C]K06[H1>QU[&LO$*@;D,!:&@<X6=Z0#S$:#U$F=FD0Q4X+Y+E\H) >VN]R)9C
PG,S00)#_M,<]O[IP W33SE>F YD3U+-<D<R# 01X;J<[$E%7PUP,QAAT;K?L.PVM
P-_\?)<4JF>*N (ZF^>.),?')ML:],X/SO<H%-^>/I5%'6+[CI!(3;=^=_4J#*$5D
PD$B/>L[/R"N<O?%[F,X8'Z)$*QA/9WR-N3 Q[Q1;<>S4V$1"=X 7>WF@$7^&34,X
PACL2,ASKD^O$L &!*G@?DMY:,437_6W+\#1HN[I[F&K*%3\4T42VY,L)P2@Q?GI&
P%ABP&M=1MFSWCY=XP):6Y]'DZAD&&HH@J'/N 3^=I"QYA<WS2LWZ]FJ6JSR:4+>Y
PYT$?Z\/ F;6.:C&!L4]<\3QQAX6L^'XU46Q%>&Z^,<;3.\\MKJ8@4I-IOC!>@2/6
PH(*C0L=3&""=P?S?O*1867#V96ID4'6)<G,1+;A-+. 8[#.8\7J,/U29L!1U$]RG
P*C+=-!.%S2;CT$1RL!.'JBYG4QL-,%,L6_A"-8R)8T2=RV2<46DQ-;*BJ-FSKE;X
P>#\;SBW5LV<<,I?6K/1YG14-[65^CF%0O: %B;<NE\<1(<<2@_<9T@7*F2X3O\"'
P8Y_@,Y,MNGCK3UBS@9 /0N5;K1U+2G'8)UPT<!0T_7 7*>1D (7ZMO31(HZ!8OX>
P8P189ZW $\RQBH^&GSD=[DG$WN!&(M//?$3=!OMPGOG"9(ZFX8NC_;GDE*K5N,'J
PDT\*,:F[/(=-,6UDW"RL,P/OH?!?DNZ./X$ .RI;DT, F9O7^PC^TIPYKHV8V3B9
P>-(B6*3GE"FL2OR[Z>\F</@G^2Q,<FM(0<ANFWE/N9-G*5 2X)BA"8RW&5?JE\_P
P$N;Q&L*%Y-^>I ZR=%KF2O$I1#A,VX*+#H+S"PL?W\H<"]$YDF2D^RS\:*J3)J$&
P>*U8G C;H(4V-,RN?+N1+SRO%#^$T(6$QJMHOW-,.?L"5KN?61$!!C!%V!L*-<LN
PL)\[T8SN5>T!/7"!E>E.F5_?;8Y1ED)WF<=:&0!&)1/J\^W5BVFV:O=R<M)T;,KC
PC;N$Z/U@#RDV[C-&@!#??AY%9$@+>* )7%%R<G')\TV)I]4[XWB2$Y8I4();&>T-
P\E^"=YFW8QZW]65*QPC:COE%1U! ##'-6K*0! QT@\IQ0VES0N/Z322>#8^',[O&
P-)L_3_L^FAST+I:8MVHG:-TTY*Y33[Q++$H-_&Y;3+[ IG[NPZI=4_D/ZIEJ>U4.
PH$,J!,7/1&*'0GJ=U1-A;M#<P25 'TB 7V4D)*"*ZP<P;8O<8$JX0N8M2-D!^C!S
P"Q3>(!E+'\QC>S:=Q*FT<R %H':(4M5;W1!M ;T76UL(-*5+<F-A6SP<DP+[1G4 
P*>-?C HSQKY\WHMW*(6C"1&<\2KC$.I\11\K@DGK,?PO( O_)( ER$UAGRFM&NJ6
P#%?_U<O4JG)84'8J(KX%32[3YFFMKW@6B#&".](!2N!@G6JRB8H2AG@9Z_Q2UK<4
P1#E(Q<U!Q5N[2: IP6?U3IIK&)[<E#TO4/T>M=I6("C #Y]._,VVU[7KR2>S#VJN
P!Z-:[,:[(AWMB9',A36.]< LWTQEZ<UE8YE=(A'2ESO?NR^T66%^'9NVWQ10R1[E
P]+%K[_F J<:)H  ?^NW5SE 38CYU3A+P\#\%* RV1^Q(K<!XNM,7T XJH%3'97D\
P@*.UL;S0W?XCQY@X& &GZ6. !V@Q-'KT ?\D=JI" E\Y5LR3-04*[.K8!EC2#SMM
PR^N$]3V6_T2RM;/F%6>5FP+?O2H#,^>S^!!O8TAP"25?5K/G68P]?9=CM-(VZ$6R
P*AD0<=7/TM;5#VA^!7&358K'1[&<'$ FIB+,G>VB1J*@@VM3?QZA*29W0+)@5MR6
PG6I2&:6/?89S;JY6(?;%I_ \\@'HDF5-P U8=V>1#]E=1V)\\FE:,JY<.0B9J-2"
P2HFN)S=ZH8,:BW1NSA($LR(?6QX3%"3_(8 *@,MH_4Z/MUP:R:+^%[_$>?MZ5 :W
PN2.-^4XS^F%*4A?B%G2*/H#3W]%6F36.T?R8[A<.?4NZ ABG=MD1@UC?PL6F0@$.
P^\@?]""\&K*_8/LC8R9!V9- N)4 UBY!,)=!LRS0-1[9W[( UZM84>$(\R%@#",L
PCO%FYF!R]=4<[-3-LC3'MNKO(C4G0 W%7E'K\-4@$E+DYAF<X97CY< -K>FT5V0[
P9MJM*= *0^Z(Z-$YI_\8\TIEF/-\H+(YYSF5:T$BKJ>R!9>9M8!:R(F+>U[Q[>DU
P(((4T6C+A6A8:6M/'6L7(S\&1CUY\X.XBHP4%F9/UOQAEN7BC_6JDG55<X26%/+=
PNN>L/O?BPT*@PDE':E UJ*[R%EN4]_?R+L*_+R@EKCBC&7\U%,1Q),&.(D#B!5BB
P/M5*Y;"D(9TD@9N*9K78UF@AR$F2:"W@K?]&GOMF(G^6T(O_-UFG4%@C )&%<.4!
PR6IC0*OQ4CB#8,=N8I)[S"]8K<[F%O%<X58T.0Q.@\11: $',KD8BW&_TU[ESH>D
PYAD6DTV6P!BF!L(U^2+6!0W[,+#(%A1*7)/Y0PA]763M(L1NA-1B,MA3K^4"ARN;
PY,IL#OFFJV64^S.LUC;Z 55):DAHC::J^%NLR'D).A]"$5[8X:=\MG-KB:I;%#6^
P1N!B\01!8[*^(F'!M6!$T\%9]:2H2'';3"6>(MC)SUC<ICA812-CJ_V[P3HWTQ]Y
P/?&'-7R9FIB('\>E2A[NQ!$R76RLQ@PB=:N"17J_(&=7=QP\T=F,:5AR$-D97$_E
P" $K>CFQ^]PXG6#%1;"LP<:L^"N$R<6ZTO=$^E55@F#3X5TA8E35)-)-)90&: 9D
P9.71B'IM*MCJ(C]U1Z;5AC%K-1,5+RX+DT4&"LS1>=DKJ=SS49?0%#&L9NY0)KYE
P4GG-^\.NAVV4U?6+1)&9[LA1@3?51LT?12)M]')U;P_X)1#]-0B'O/*OND\O9R@L
P'>VGH319EEE2<8+3>K.N#GXHTPV*K+KG,@AV?H>BC(E.(R^:>9VWC#G:FJD[E8]7
P3DPX6DY8W))T:DO9*PFW,A\YJ-]0A>79>.<Q13=8E]W2A/J2!'?&_L_>:#EL@2;9
P%0/H;6M7;S LF;QN)]WO-AXGCX]*UUHXU]J$MR#91M6?# G30H84 !:B$C'F+?LH
PP'4:!<([G4M*X.D2[>C&/# <Z7.1A%5C'<\I9^ -)1N2O'<PC/V!0CG4L'CJH5]5
P-[6R8!>2&EK;&FR_R6U)0[6&W8\;H*-M;/N &C<7$]-"RAL'X/LGP 0PB@I*K0HK
P6>>K1ZS4&TJ^R^R>ZFN->]$V)&1C2$%I"YA^HL.5W<4M5F?QG*T,7@O<6Z($110=
P6J+:G.;SFM4UE?V<^8!/@907(N1OH5?39B'9JH6*_#S'2W;,@VMD1.F_F(&2/R8M
PR>!00(1W/(GIF79XPOR5V.9>/_X" ( =MEP7&$',>KY!U"O>7]*+_2X*@"P_2%#,
PSPM?YTRK-.VS"<!*%Q#%TNHNDT@ NFKK0]\.CX%3MUHW%;XSY$:V4I?YONRX-.VG
P$JRGO5JN."J2-0"QMCA-QJ,&&I=5U$.1C.2?2-SO%'@_, $B;$ .;:..@RW.)W]J
P'SOAJ[;LLQJ[P@'@(]>U/=$[WB>>QM_0EN5Y4JQ<$;?ZC_1\*.03&5K^H&-I+'T\
P(YTA?$52_H 5:V[5%^'!]L:QJ1JR] 79EWK!_HR76.<E#\BI>LP6"E[";:1XE'\J
P'X4$D2267]U,9)X?PD =Y/?'V@J4WNM,WU':0B<"6#PM@SI8=4R0=*M7JF"XF/0E
P N8ZCL#X47AU40WJH1^KA+GWE5H:G12@@["?!XY:F(SW!HCL+T3]U"! HG2X>F<&
PPRSUH"/:P9(#4_TJO.63"D+-07@F<V%81F&7+!R"G&Y, ;]WG67 AIQ:5;M$XPJ<
PON"S5\NAV%L>K#< J:(:DR,4W(/<#>;&-LB'?^RA>\X;4CK+EFU++:<JQST26AVP
P>:_@10WG.!<WB,YA89W>U:I<-I[=O/E+72TX.WZVK*VG%!3^7$$A36PY1.W/0=T1
P!30)X(D4-6IH.93Y&^1W\3X8HTF>D G#Z]&':*KHBF9DCNRJF;4<JG,;=/:)'<;"
PB0UKSWUB/?;"LD2R:46ZT:PCS[>J7D;F7-FL+J7*266;IG_ I#*5XF/A'$7]-9XF
PH54$GU,J M'V#]7YWI:P$R:O^ ,=[ML/&#U4+.$FC\J72YF3.+7<WX)H[P.8W8"H
P2@*V.E^ 0+"L5$6A?=9C^IA:*&L68$)$(XM'><PK]'CM+P ^!S.]'AYY=JQ+[*F\
PJ8C(>VEGA1A:2$*#2+-5W6&\NV4DCD%UQ1TH&98F6O0E$9J-\ (KA #;M>LQ>'?.
P2:;#22P.7!UKXE)&_\N$&1C5LS#*GPSLS-O N-?;Z[.HS.VCM'(4:EO20\D;6GW:
PEO(KP5KIP?ENRDXG+K73E-R"]]C^7K_RC&[2:?>M(6=;)Y3:T+ K+3F61%G*+'W9
P >@T4M_D_1YX_J.*#TJV'$QSA,PB%8.^L&D=BQ2D&#>'S%FFHHQ2_B..&&4C12KC
P 0T3*KB_7O"C<.NK*UL?8;ZEO?O>2(A$\$=YY1_Y@W/3Z3Y[F&;5Q/-XLQ5H5JQV
PZA/-*Z;I7I=HOU0L"==VH=J&QJ#3+V.A/U#"=)X]'98JJ$-%+<YQDT;O .2()3SO
P6.!L'Q^$C[M!AUH;WF0V(-K:U]5^VW"&DS#]I%[N0X!LE#K*ASXJBCF_3$FV"QTF
P(\>9*M-U_"[KZ2W:%:6, M</]"!R&B2#U2*.=V_1DC7^FO/=2_M>[.#-<O41LD J
P'>6H0W3A5T.)[[+=".JC3E])X]57S"BM&G=:-YYAG#>J2+@J6]" 6DT=F-P+F"M?
P#'ZGW!CC_JF<EM6:3_CM)?^HHXQH(4/GC4"L-G $$3C;_R.&4C]\PO!0]'UB@S[K
P_XYTOTB[>^5%(AU-DN;8:"9)*G:1IP:JNVA"MQOGE*]4JP.D16P&M(^"3W2RY0EH
PNY=;[XRJVPQ7>9@_ @>[B",BE&;JE'&U-.;()13OQUQ;&[E:!2U[=YP/I NY=QGX
PL_=<H"12$L4=/V0M.C!\Q1K;4RMLS%HQ:4ZI$'G>B0\\2)HV4I?*7$$'J-!UW)LC
PA!M\3J&99X-6 ?"UY/#]>"8]KW5"9<3&[$895:)XU<69X#YR(0GVH?Z4#ON^Y[2M
P ?K^QY/1S;JIN4BLXG!XN8)@4#NX!J'J%WS)B2^<@L;HN[$'3Q@;C^HAIO/F!<4C
P_!8<=7A:#2A9<4;&?NJAOA[S9$33)A-PVO#C?T=_?Y!EZ@*;%N'G:&]ZC2<TV<+7
PZ@+Q\!> K!\_6BZ[;GZ(E4CU-+WIECP>@:9Z*69& 0?S!&F-&(+W77#ZF6BLB:#A
P0=-$3>EKO#![OYQ9N<O*_-B-;&=1-Z[T102'_L0(*<>GG"R/RUL?4OYPF8APC(UL
P?'TD63 C--K4HL=NJOV>+=<",+&L_+0+^WK91K3RM37G+=IZ.6'[,XB3"?AB/I'V
PZCI00J?\ X!JXJ6=V5SIL7]ESL;R+TQ!*-[B#?W_P0BD[ ."1#]54I#$Q)55]'4%
P6HJ) U<D0'3.+]^*LO@G*%:[XGOIKY6^X/?!0PE.=XKD/X4$U-T&2DSW,203T!R;
PI\1PIX M$W;O+;RQIZ^(%#NLD# 3QR24[C+G=W)]Q[VLQ;];P:1M&WAE4H2JZ8[0
PW7]0'H>T$Z ]%N>A"RUM5VLR6[AD33E@,M#\4I&Y"D#S8;^_O GJ(1+DB89V '^L
P^%Z3WD3AFXP@^/?#%L]GG1U^*QH#U!\BVC=IQ5;)@J;"I@@GI9M$,X7QO!AJ%$S;
P6^T!>HK',8O&E=:9PQ$<1'Z-ZA90G5< QRK0U^[U1<:UD,,X )BHOP<8 O0/G"\7
PS&7J-MXFS(O# +&<2DDJ=IG/+I?C$S?QA%MYUABU2<?T8@W#[09 MHE3H)&FZ,:6
P/H9^%)6R$V<M"5\8(QN[1,UNK"3R#N#B6\B/''%_;LC(+<[$L-XN%J!G540.234J
P>G9\M'ZOJ =%Q@=?>V"7(M"\[LCQV;?</ILZ9\69U9XAD1C) ",[E9RTP0*]\?:=
P,^%'\T=$+H6^;G_- !6KQR?&>C5]82B!%--GW)MT7/5 +E0(?2?_07@S5^R;:,ZW
PYJA>UJXUCI\ZH*%HM$2A\"B<]Z 1VLHK/73U)3K0PW%$@["M39CT,;-F+VQ]ZP?5
P:8]D"^#2K4??(_CF#5P.V9INGZB5PHC\[7ZK535R&(2JN[*?C@^A-N@U*.'.]99&
PU((!W]X>(SG1_T9']FE4[[UCB2\:S-]\;G7/Z?-M:,%!7N_O<A0U#29=[Y(:5Y'0
P B1@8,;<8NP:\EV9Q.@$/R<.BX,J<=HBUF+^?;Q9DRR?O99]>GM-WG?,GR5N:70P
P2]CA#%/=1=B9T>IG*([1,>AG_-+9K+Y"Z<1S@8V"%7_.0F2HU8"%0?@__C;ES]P?
P,BP3APZIYYBPRI5.X8+4W\TE<@=6??F)UFPWR]<P"@#5+P&7G_1$CDGW"#^L3!1>
`endprotected128

////////////////////////////////////////////////////////////////////////////////////////////////////////////


`protected128
PW%6N-7SP_SO_TK,3>DL!DT-1M\7DG![]> 4:6,=?0!8.J\K]2J55I<2N=C=&Z<7U
P1HXYKU)%WM"&=D>44HQZ A=7/S=:]6_U@,_UP\X!!G#L =LX?#WOP7=^AI^K,W:G
P1'BU1++[6*XK\0E0D"_G49@JH,4P87EI>UR^=NW++%_2QI.9#MMB+OWN"P=4XOB=
P+LJCO:PV$W<W[-@ L7D3.'(6XY-*W2((1GPZ7^=!O&Y-%R._5*OJ6/L,^F5RU1D1
PD+!])J.)(: Z\%5*R,DE.??HP6@+N+M3(TF.%&"Q2U@7!=2N6FNXESZKE),.L,:%
PS?X#H* YLK%M$8#$#C0%_,$5?Q:8BL-8N,4Y)6MV]X$LEQVTTO0'<Y7#[!5 ,6EI
P;,!=5^7"L213UR99HK[=DRE$+U'Y%*+K]F';A<[BY90F9Q:897$JW_WO"+U,HM\9
PP9J^"G&S=U4$!($U.]]85QPC"@.Q+:",+4%;_F8Q4R*.I@E:<Q%YBKUJ&G"CFPZJ
PDER:E%9$[L$TN$6%+6!I960R*\!K2XN \169F7A=>)1+5]+JU4%+9073Q'!:BR+S
P&!#3D6A*F'_,AT61A*VGB8Y(' =V_XU&+E]\;)H*H0">2\UE;@;(23-)7*7%;;<<
P[EDQ'CC7&#6K@FYP0'V^DD49*79H(9<J%3FZ'1^%T&PNW-QD7'>Q^.84_AGGHA;6
P[,TPBS(TB!]4?'R;,I+Z)RI2WH"+*0B3GP.QCRBK1'T]'?LMW726%V5\>542_EW=
P=!TAF0B/K>?D?8ANZC9<5:JAX10<RRH6)_,%;"Y2@$(2<P:OY0:Q77#A# @B+M2&
P7;O?=_UE'M_6%'P#S+"<NU5I4.FWEX)X_NTJE\"\$RK4:KWO%HB,R<$SV66.]P.T
PHSP3!_G8T=Y-H>:..'MBCOR'0V"(,)7)3?\@\7G[Q+]TIO<*Z=TNJ^6[Y)R/+],V
P^/)])'ND^=0FAFP7T9 -TIK1SN4>;S=<KEAU%$36?7'N?Y4RMXB9HM#6L1ZBP;86
PO"&>[?O=;_49D)JB3X@"VYV&CD0)U-UC+<MTM?Y4[6ZG/20T(I WI$3BH? K2.F]
P//FG7DK?"%2UH+B,HD0^BXV6GUN/]O-ZYL#>DT_!WY9Y[%IAY;!#U^<YO#JI4DZB
P=8A ,R77OA/6FI@PV\C((D5-PEX3+<%<.Y4Y#PU[MLY2N^O97G+@1KC(L;D@Y!H^
PPH;R=71DKT<CDZSF9#Z&?M&07RL"* <+*_ >)BJQSX?"-&E+1@F((^#UHJW-8VOB
P">N#;-F;5<.>[%R2:E^JTK#I-F_2V](53J*:V3 7FR8/+/Z/\X, >*0/?(H:N-&K
P/ZF_T/"#+[8#/9:]XJT?H:CWO-FW:B1 ..R-/LEI@CB^:ZB0L_5:TDG]J@B%]!L:
P#>C*;WLJ_9!=T*\4#]7,_; AW+3/4SHV5# ?BSHA2WB?IG?=>-.YG3)E&?Y9U_9W
P4MN/Z@6;23E\&B:4]T58BH:LE*T:2UWD8WW.P7;]8KE=7N5%M"C\E]@WV.B#),M#
P06_/M3,_>_ 7$BPM>LKM(P5:0)> )Q^)!F^8ZZ=7*>W'P?^TP3;J%8>6K37. !L7
PW=9V"Z$N]VJQ9TP;(,D@I7S">W1MYF6B%QULL[WY,]W/X&7X%29PWZ#_$"AVY)N_
P_41N>ZLK/7J]24.'9VI_:_N(60=!C?%:O*MU,#EJTS]Y\K*ZL:<0T6LY5=HU:[+ 
PX4!-V :'E[01'T\0F9W^'#;*X=!9ND@A,O4[FN)C.,.)@,<W+*^+$N8+5#0W>/]?
PL1RS%Z/N1PA_@CIZ>7].BGQGG:).39"81=4;JJHAP=9K\)LUW0X"9Y=S,_. 32!\
P*\>AP\:21Z<U=U>:5NU!LI_O7K*O\0S!/ZG=;#F^BGOO--60EQ#=45IM\$/0H.0>
PT-:9NYE*R;OX;7+71%D(10O6B!*4*)ZRQ%&_.<EFX:]Y[$*S132XMP MY\Q.3S!4
P=OQF@4&G;?S6!85Q5\T5#QV4^0NJ"NZ[E=P.%/-P"^DRD$KGVD9]]#Z!5TD^YC#*
PA',?98S,=U:K8MOMJV\$<9B]@HHM3VLA+E2)EE\:6EE)U9Q )L$/IEBWV.L)9]:A
P6&]\B:BG##<-G;>,*>N%H/R*$#,T$? JN+.!EPYYN#,NI@]()/O_V6."Q2R0'X]3
PZXQZ%][A@5]Y?-6S*4"7LF8'HEHNAM%]*L5,.O79[??Q[_VNGS6/0"8:'6!/?!I3
P8[C]][6W$@;Q@5M,E%\8#DQ=SM<9^6U\@FNM0G@7U&Z%)PJ*"[Z/]O+O5\)4S*]%
PYF4?)U[2 \PFT@NO,/C)$;%CC@6#.,&H7!%8]V78:2\.OI,R)AK>C7D2L9TE9?,G
P=7)EW_U&'Z-&^;-O-J%]OID%.W/KDU(V3= ,2G[2"FF:AZF3+70!_;!",<RO$J??
PH3=D5S(?I)O%@_>R'_+8JG$'YUH 787A,-1>KK*UF,X)<LB?TJH$0W$#&8#)J;;*
PNSRN%"GOYLX#437'G'?=J[T5WMV=Z<X"3"U(E0/'-"-.D&4_S45TOAT6(S&2Y"]Q
P6@1Q!P_$.3V)H&GY0]9CGV6;V1F(,&P A%;NQ@9M 060O^QT)1+(3QEM6:#</G5T
P.[3%X0?*=]4),3PY(U1Q ^YINO?],@!0[C$6BIIZT5^Q;KG?*G#2- :D9D\T)(D6
PW,!XDLH" HZ2/-21@ GBY[(&5C7<^O';J? /.'NC-C/U5#B1ZJ#Z_&<@(&M6IH^_
P7<JJ#YB B T^7Y+:*^PQE"26-'I2_&S;B_Z0"F3!6&?E/&;G]O#-+4D,W'V$HUN5
P'C2"54X#I>MI!TU=V)V=?HMPUZFYJP?V.;T 5]W-289*0_#Q0'6VG#8H.Q,*!K0-
P2^$;=?;W"7R(60XX;92OL5S"+&RSWB-.@&]--2XQ[#YI/7D<%I [":E[?[%"(?59
P^3'*&M++9=;YAW*G5)EQZS=GEG*W@D=JT^/=EP7T+DS"1OMQYG*-/R$()PA;D[D)
PQ+O3*@5=O8R[-@JF^K%]V@^$G=(/T-ZHA,0;"]/\2JU!/%H];SWXO<U!FER9[4 9
P&< P6068!G<)XCV6^PD;0J\N6S$S<\+&%.N\ <!,S3>E=/7Q[G7*'8=H<;:10SS'
P5.EG@CU.GPRUBL:-([[TPPKC&HZM7D"+1&RH).6=C*C]09O*44B%K]81*C97+]C0
P0W>8LJ4"B%G06/)J_*I# Z@NH^^@JRG4GVK])ER#Z&757%).VO*"\>?5N-)*=&U5
PI9U#KRR685$J0="\3FJ="WV'[O]VU3(!S<,.RR)G W=?KT!AZ-.);&RSK05ZVU2$
P07@>%,I,R)>;9CF3#(+#@\2RPQ(K!2>E%0P7X)H0_L0^OZ('C>3N!H*Q(@R%JZ6H
P-DRVC_7[[^,3IW2^>/XU7C09>E$(HT6;GU9P5,?!OC0_##H:\$IT<M/&HXRW#*L;
P'FP/\*6%9H7BCGY$!EBPF$ !3'2^G[/7S6G$^A>KEK!H)TV1WK"Z64YF+T[!O1N3
PD,)H0.F!;*\$\6SZ5%:"G&/,>@DR.N:N@K+1CM)9-!83IS:'00)1$&13!?U-/65#
PYD%I!0M0;C+<\"W6D*N8OQ_>Z3;%A7SFD&[D$%)INQ;HS">I;[^'S2S[\GR!%)\F
PP47(KI=-+6U?HX8N5629SU,1W; J);6-:WXH5>JW[\!)J;C<=QN+O)0*%L0UP(;/
P-'(P^8J1LPR9D Z-E'>L3Z:9COLYP="6%[X=F AC>>)ELZZ,9W^E.:^NN8TAY$UQ
P>D',6OLZM DFB+T6E4HHC]"C7V[\*K# U7B1;-?S[@J^)0.5Z8(.?^ 7WX:]JA*;
P(WL=DX^-]#&:Z@T_"L <$OR5=\WU66[OO<0.71:-UO[V(<^PT;G?AU0AJA>!&U%&
P1\(%]4,IGNW^9J]F;4^[A7OSZEJD'/_(E73-R;EVZ5"+RKJI*J<*BPRNH98:^-A0
P)XG-GEIVI->WX&,3E/F\084I;U.A B= 'VJ5/3WJN%X@JT;_M'.0IF11K6D7^IX 
PIO^1)OG:IDLDRC*2J-2;:$K7L5\>X;M.!.V],.,<@C]LCO3:;.J*0_=SW$ZYQ\#V
PNO:%$"85EF RLP1TC9%=+=F*:W37&((@RV7(8(.+>9NF& .=N*"U2[J$]#RQ6%!J
P'JY\Q"#@5Y0^&;JWK\*AF\P>O]_L#\5UL@WTDDOY')XRS_\+9XQ^_MX%5$U$^P[C
P/FR*VY41!@Z@N++C<[3W.#JQPH)CE5FUZ$SO=)4#HB H;"(-X$0?S8T0<D1=A5X'
P*>(3.GGMD3J,&1O9O 7)%?.5(S['"H%QC'9E;>9FE/-O6&7WY-J#5F2(#Z&N'43*
P70;66WN9)#*<A9U;A0FZ!UAZS"6]O#ZHO^'+NE##CEB\/ONV8QLABG!K46W:^3=&
P499YYGZ;QJK07S.EE%CQJSF_%=6#_G5M]4]5<X '?3I"8Q0UWX^F9M@ C--.RA)/
PVE$%*V=:@/$AIQ>3N?HJ]R9<YW?#0X=AG!.-C[*U2J&18[U_S(:#)HN\"@11IZ/W
PDQF(?EJN\6>HRG!J%=.'C\+XLG;$&I!: D%!NWHP20%:)6HQ&*I:1OWUW"]UA'5]
P_NWX1R E(=3V)D.4N)#C7;,21/U2L<8,N=^8$QUNE$9]"5T^D\Z.R"\], 6<K'*\
PBH("$?UNJQBS%$J10+L#[X7($6B,6@JG;R?TZT5AFU2!*6=TAIA\F@$U).-3#S&8
P8EG].WIXPL:(TR7Q3-'$ 5+[[D2Y,_$P-V;@(NG2QNM\4W[L_APRV_A+]N=7C8Y+
P]/Q$\Q1<Q_89UT*_U$2IS+_90(3AQB*LV(FZ]=H#+.8TI6O@5N"5YR^^HFK]M?Z]
PQ.P<P.@NH),8#7RPHLJ*@6'UNH]?O,:6UA.PVU],M[&KJU-;(VOYG\8L07:7V%I[
PFSXK"D[=6S>=H\)@P^U\S_ YM$H0<K*7%'[Y,C_05AI:#FU>U'-I85LSS/)="IZG
PH;JK%;_E_IQ&&Y4%D^9=M4IX^UX'W:\^60>[_++L+^*F9*/=K!PX@H!?G]>KB\X=
P:XM4 FGCV;"@IC9PT-WX_@4F'5^P\P+=WI8%;AQGAL_W-;L824%?2MC8&D<(S7Y6
P:U\L A]ZJ48'K\8!?U'.QN$9S@4HS (EDYUKZN2)+'FRX)6!A/#+1RFYE-EO1F&M
P/'B4MKU(+J/QH9R"=P">?_$D"9UZ*AKG@<U$FEZ4+R):JK*$QQANXAH;_>LM@M5_
P0]S"D^C%7[:TA8J9YAMP</R/,*7R>7-TR4]\R72'! ,XWES#S:$DM(5+/LKY;+V0
PQN<!]*QJ;;:A0[QHQUSZ"H!9+UL'2TQ=0'T!;LB.UHKN--K+.=U%-I[CT3S"EM@2
P@7,ZJ"I,T!Q6$5T:D341R#IKJ<[0)>0I>C("A1ZBDTBM[IJQ7P'^#9DI/+K:W]]N
PF&=L2^:3 A07G 3)$S)Q(B)D^[A<QL9.0GEVSA]M!4T:)$@F7:<RWH%WK(V@@__"
P-9'_P*>$1PZ7-ZV7XZJ.M4",$N+"#K"KS*MN+S]!Y1EWMY=0: D_Z!#(3??LVZ+D
PV]G=YKW=AF,W>)C1\,U)#W)Y3"N34?:&]P_LZP2"!ZH4A.3U?O^#9C/UGLF(^=, 
P*8D=]!,?]B_8$A=1ZJ+LWNL0 L]8BR3G&\=CK81G&8I-_TR%N]?[<$>DN> &DJJY
PVR0>(B@=.K__2)00,)'4S-8#4;(@0^P04II1&@ZN;B-4A?F#D9>:+3^\["K.$]]G
PE:#9:K.WXOL=JBGA3*+N',Y.:C-VU8#O#&U'*+JG^Y]0%]&6LMYZ_2.*&T=:YGA:
P,1UPT3I^?_4I.3,:[8VUY(/?X0M@N9OC&:(1J]F^CE\^,"-"KKFC=R.JS<&B*V.B
PEH59I^BY!JIE#_%:A\^4#W,7QI<2B408Y[\WF9Q&FZ'*HVIQL<M=$\R(NMT=05]L
P(KQQ^-&>45/.AYHT"-JF  7ZB.=#P'GK7?6UY/:\<5+9E OP(7)-R<=QB@FIY,BH
P;6,A@-E1-]%>L&U<.L_PL,I&AFE8>4-]3OD?IKZ@KS(H+%<F$Q8*N7X&O< (E4U_
P+X!.V)LM .T[,:A&W!+G4W>/M=[:3.AOOQ.0?DCN.)K ?>JF](-%WS& ]8P%*2D-
P#1G'"H,^J1"[EA[Y>-M7OF1X($-A,S8-JH^>5TGG8;F23&^]]39V/&$M27U<Q>5M
P[HAS#J3M#_>L=#P^0,4.=]%)F(7K]?!"C%#\XMU'-9Z@\=]R-5G_]EV+-(CK>!KN
PC^>\@;#Y$L?*Z1-^124)TOM/::+O+.!O8,MA)A@%[7;\/,O>$"D_MV@Q/*4/*U,:
PPN^4YYHJ1PJ!S<3Q15Z6G5.PY"7]V1M 2YE*>0X\A3(U_#\]V0 ,)$^3+<&3V"1#
PZ&EZ0<(0+PPM#U^MU4NK1L/H FH H\LH)+Y>T5 ?\<<TT\KD&.^WHQ)<DS<V'#7I
P%.?;7=N&!).SBO\X[87(FGI*C&'8/3J&P^UF7H!3;H8CX/(J8-IAV3&XUZ9X@-.9
P+4(6%58SC&OUGYY0-*O*[;\KR6C!4!=9EJDM#T;IP-J%2TJ&JM]\AY7WJ3Q[ST(!
PE9*_DL 06 &P,$^*T00,9S*]+%0$$(T+TU<AN>5F!VSFCN/59C1X+TLW'B%J[5VI
PL_O6;2YVPF4V]VNB=;D&**\6UNUZ/E[ZS56;8IG!Y/@1.O.-J*GH_>R1E9<'6&N 
PWB%M.%**)HZ'QO=0-53<Z\6I,5[+%1,_7%."E&7K;#*$,QGFE]5%/B!%V$G+@<-R
P>G1JR^R-BXIHOV8:;9>2O)\1PU?"ZH16P1&9?6\<KQ=UWVQ=JBL&I.W'"K74DV<L
PPP.VBCJM?E?_LD-Y!S2?5(2*<UA6W:_#IMQ'GUT]F605]C5SGB'=(A2.ONE>80ZP
P/T[@#2VW'H"Z8X6(9'RBK/'2?=/?IZ_E1P.P;HR>$[B@*I=5<DQU=]9!-7@3APB;
PP+0VH0]3)D7\OVKTJ/4 FHPF!NZ"WGSAM\9^'FS" Z[(1+__]T.J&H:6Y6,#6G%L
PT(<)K#<M!:?I(+<9>G[WQS^9^H&T/A2XEQOGE!];;O2\S)K$Z]E)AR[;^S7$^I'?
P?/%[C['RC,H!0'JX?7/$$OA^%%3_(WW52SD&>=NO<.HYEN*OTR7S<1Y3*?*6*HGA
P0;;QQZ'*5DO:@=!9ADP5>FDMTD7LM@?Z?K;2ZK5!>7H>/_\#9N_A/ 3KFP@;6IZ\
P'7$AFJHEAKTY>%E_4S5MM(-P\[TG](^O-]>XSX@]J';4N[#OT9Q<QVU?88[GB;W 
PD)KXP:R"3[RIE?P]!GB:S K541VZT?>^UBS,BG)8(;A%[Z[%D'""%'VV4(1,LJ37
P/(];QJ/OVQS(*1&)<.(:[\]8'+8>YAEE)_T%RC(=L_PG(W*&-S3TQ)DLX>:B]15\
`endprotected128

////////////////////////////////////////////////////////////////////////////////////////////////////////////


`protected128
PW%6N-7SP_SO_TK,3>DL!DT-1M\7DG![]> 4:6,=?0!8.J\K]2J55I<2N=C=&Z<7U
PF>S#:'*-QNR%<^)6=#&>ZE')M\Z%;FR13T(<YE5'8(*YENN 9KJ_M?M84AFMY4**
P23\K$DZA2TI^M.F8<5=$),E.+X*]&3@G39VL]B3NH8R/UH9V=G]T13JYA'!+(L'N
P_PDF_E[RZ%A;O P#Y.[]%J%HVR^:;$R"R"<?:F;1P]VOP7=!R S%3H#U%*$A8X8N
P'&DZT>BU#XM7K]@;UG&4JSEMH^/^]3Q[ J88 QK<GL2YD25(7*4.+X-L740QX!?S
P"9$( A%7 NWCEQQJ]4"0R(N(/T4Y&=4;Y:0-;6B($9/V!N3@:SQ?K0)%<)]%;J7)
PTQW?@&40B[*>5'7WLKFTRB_[T\]*=7^"T',C&2D'!I8)@=#-/_MVA/+D[(%)RP[L
P+E(X,QN$]OTO5$PG954W"A+S3GT,V?;4%4?AR# V[MG_E9_W08,=KM^LGVTDT"U-
P56:)AZ#O"EVM&>TJ#EWN_^(KEFE5=#@H" 3V12]Z?S";'.J((Y3K%1G"E!FWK'@6
P2/&[ZE/E #B"GGDWY10N[$/#^U1JH\L)4@^GHBTO;[A[$@%?=X5P^J00_+ZQ;<QP
PP*A#:BO.*?A -T45)X)/]L?X-R%XPR)R:1IBJ:L#<.#X&C\H0 %=?-GETV6,#&H0
P/7?[W2CY.//0%9GI6Z1JGEU:!>)8)5H*$M@BK 3T*4&.D7]F0SP(65<T< 471">!
P!'!+?XW?>763")JCTU(<U"B5\0J!=8]25W:8EZ?0%#$^4KD=H" ,2/A(#\CWHZSO
PM1IXN!3$N+ 6)15/_))/SLBJ'C[=\1RJ/O.<8C&A\1RK1:W 0(&0E\H9<SV74IKZ
P!K.VM!8JB]%!+3AT17G3YWY+<';&M(%^CZSX.>C ZI8@L% .APW'Z"D>& MOZ ..
PK&VA9@6I]*#(]BA^8DTZ=FJXM))%0*Q)E!HG\#5Q8S7JMJ77)ZM=78.FGH BQTG#
P,B[QV0"<Y[79QZD[:W_PHFI9;_T*YT'-J &*Q[-&@+X4HQ4FY:."!4^%TT.D:M'>
PQ+A#U:R1>L-DO,4- O7<S\,  I7'=8[@+GNY& ]NWL&;.LDI "2>0KP9*^=!OTX6
P6S9S\C.F6O_.%(U=:^H?9S9F+>P?<4:5]0.WB>0<PJ=W34R-^'>XL@3%^.]W$*8N
P>V[>5-4\L/72AV(,<V-> HG:.Z&&^59"D6G8*&_BR4S\&&T9>)=VY73,!2CVST '
P"+ZFR2.?R+_3?N*JW;K_4>!X<(BU=3 ^L-R%/^9X?S.5R2KQE!81!=]$FOI_4<^<
P1%N0II1.OL?-('&]2=3Z8EDLWR8IL;JW.<>#U;ZQSM1HU# ==0@9D8Q"<')_+!6?
P^5$C>>%;IY^D?OQ(YJE8_G1Z.ID-#027?8,\#\Q6I"_UA=QV'IRTC?)O/FX3+OI\
P"Z0RPC2NR<\2W_I=R%5&3Z!).\D6IOGVQ@^'J[!H*D"]^\E8@Y'I^N<QYI$/<V.F
P+;V;&DCE0Q0Y#,58YXE$?E&34?>)9?Y,Y]TLJKA9GFDG%0DKB'O;Z)*5C4M-36R6
P6V&?3?E-O^"!0=B7@-FA# CV6%@;GAH !\'B'#O@3$O\ >CM3'1KF)@JY4$[VA9N
P7T5@>:7C@FM&VL$4Z*#!%]?ERXZE$0!+B<Q7%W#4.S'9ECF=CLI4\VVP5]'7M1_4
PBA]^!H/#+2"593^F),.S*G0\I+I<CCI<K>ETD-Y-H)/IR]O!SKGJP2IR,U>S=3>X
P6T)A]5/DL565,;D\U7R-]F5TX5>Q)I;>V#$*DA-B&7T8I\P!NB[_.W>\H)MV0<YK
PBPV1OAA@">A56R#&_SO;%'TR"9]#NB+D74[U?<F23_7_!^,G+T^;&B+"0"._45Q3
PJ?+(#9( 0A=%92,WTDNX,U9.M7MV+XY4!G& RCF\_&@Y6]O7(ZKAW.R)2^DI7;^I
P89N\5L6X4,FE047P(J($OAC<F_HAVTCS_<A8!CJZUAV]BL\(L$K>A\PO*^[NWYPW
PNG9759_R']08A ]455<L+DIV_S@;I"?H8O30IISBDB)#_H>=J:NY57]*9Y-V7O;,
P'BUA%B20"4$;050\,)3G[D<G'OJZU@\F$OBUIC646"W]L,@-WR&&L21#*O_3%:-)
P:8Z;DX*-9VE>IM8,7*%B%\8#BA'9A#0]RPJ:ZZ EOAF<OK#Q(W:=1C2P(IM40'?[
PZ](MD1X?XN3-%@*IP-$]A&7Q8G1"3K6&)90E.UR83>)-ST_*I$!*ZBJ[^_<)ZUHV
PR:< YO0LU5@SUO,*9!"]=+*N4L8I@G^Z:HA]0UF]-J*X-2O@1*UX'WRQTXQYYT)X
PHR"SG%@RL4VM0E%WIXL ?IF \X DS.I&RD4,H7C+N%P]Y;?>4GD*H<1XU;BY-_HJ
PN.A4T3>#D+CU) @!7$+/E-'TP<_?1K"1"9]YI/\(3PQ'ZT'B^LD(2>VS8?.L+R$C
P84Z\X?J<)*T]+;XB,.[=":R22EF0/UPH%.SM.=]M5(]/US&)$/G#W?-1&S-]RZM&
P5X*G%_@8MS_-YC8I7_;>%)P';4N:+K.H).#'>2O:@X-/<80C( 2(7?H80CM1)OEM
P[XQAW"(OK&>%"@;GD 1EQ>&=:\ E9_W@;TVYJ>JM'[NK*OS$]-.[/^H]?@LJ\?C<
P\5G)0;:\? 3TO>DWE=%O4*',I')"K.BZ:I9=AX_8UV8Y^ADQN'CB6!7,F(ZKV^0V
PE02S[LU*'C+JD0@^CZU&0$VJ=1@$91*?;H[45 8*:YC/8HZ>< X_H[NHZ(U3*C.V
P<2AXQKOUHEI,B::F<?$X+@R<M,>9]:0T4Y'M9K0^8D=>CO[5UU'!AM.4(C=L\_Z,
P"R?826IL>%"/+A495\_%'/J!K[P<0U=X!:T6I:C=K>$_@6_MCW([,X@1[?>2QNME
P*KM7FI=UR1!FKN6PQN!T YY"=\^>V1O]8._S;/V+_&04#ZA2JZ/?I'EF*KR<3V<?
P6,H0AKE*7>(FGK:S\9S7\BP0,.[=0>^L&"4\CO>JNZ\&DUM#5)7/(;ZT7?T?6K[L
PNI5Y&4(EZ**^889/DFJNV/?VI#"8!S0#0G^B+836<!%N &*UE4 EVA)@ T^&N)47
P[(&)PI6[<:^?P%G\%%=HD1\#K#$WK_\@N/MM7H05;38HR)('WZ:DOMW#ZGB:NA.\
PG;%IMH9L08O34@\QEG6:$]$X%((YCOZU\0*47(3-4AY7[A$-OD,^Y='(Q%W80[3L
P&2AO487]:<1M>0B+4>O\*?-\;N]N._8++^(H3!!5E7F*0W"D-O0#*;9<LWT/1^KP
P"JKE7JYY3_(NQEDFH SN;?F8UQ[]\:3AKYXN#T&U1X<@JENSX.0';$\),Z[_H^)>
P3_<XJZ7?U]3WFF/A^;6E.='<Y;/),MX=*5YL/S2U*-2J'Z9!:<4-*\@7\OM4T#_"
PEU!8L^.""M7:&]_>Q@INECLDNJC6BV8N"LIDQ"-ERF;S\,<OH8<L0GSY =1[^(\Y
PHUV=#C6OC4[K2920*G>M+)(O)IC#OA#GF\+T:ZD* _( )7J%4,$HL-W.MF+/6+])
P9(%A5]?R;$K,V-C4*-X@/ .W-TP&M7XR43+')8#Q]B 52*U!FA1VTUDMVXK#)<N@
P-6,$5:'F'[]/D<8G9#D%_:;GQ.A2'XEVZDB=-1,Y4]_=>.GMXA:5E=/ _&",H7QJ
PBBX=IJ0K%I[U@IV;$">0+E8\#V'W[8+7AOLD?WU"ND-\7@?C4-TR_W=?\]Q34*SV
P5"&Z<)QZQHRO(SYZ1(62A*;3. (,ZTH^JE:._B\E"I69^=+L(5D7=>D?F?_.E5/X
P-Q0C/\X@=ULWCGOY.H9*KB:OJCB&6T-#;5()JO5@]4#25IO9UZ$<X$W397>MU7NF
P27,NJ(,$ >H:)N>T58]CWR8AEUG1#BQ[W5TC"* "]*QS[%&A3Q1$$WB>-;4'L>=+
P36S!KBQ?3R0P7)\*1(H]$S3B@1"JTCI,I14535>EKY[S9V)9RJBO9O>2-B5H'P[^
PY7=O8.JJ"=F],FV\P?_,3T&W?3A)[AZ+X\%1#+]>?FH#;]>DL1"X549V66HGWCG8
P6C21*\!P&H#+X11S@Z9\^2MKZT:QF<)8]'ALPMGXFUSL[XVQ6X=LEF3#[#@+EA^\
`endprotected128

////////////////////////////////////////////////////////////////////////////////////////////////////////////


`protected128
PW%6N-7SP_SO_TK,3>DL!DT-1M\7DG![]> 4:6,=?0!8.J\K]2J55I<2N=C=&Z<7U
PF>S#:'*-QNR%<^)6=#&>ZH9R2*YLR[&9O#;?I2IJ#P/'8\XIA^##\FZNJAQ;)OH 
P7& /&EE<QV;_<;DRF,"'>=]PL!=.&'.Q^,\1/>8P\XK34.HEOVT#/B $\MT<+<:[
PO;EADQBT+I83X)3.U<XP+C.P&66!!DMS0U9OF*]@N^L&2PS!. =N3\P4T\0;O)B2
PY: L.]).6%<1[+^$92LW_^+H4& W$2RP;KI"R/5-!@PH7C,8@CT1?#$%+6^Z1K63
P]N(OM\@T]FX5$OK ?B6MTW<\:0XB[SI\,S,&IX",7R#!9#1F:29WF.8Z?$;4E_],
P7W1)7+A7VQ@S?11)_(4WC6 JDN*)E_T&B8&^6^*O<F"6RX[!-.@4JFX'FEP33T%[
PP.;RFDAZ^$H&"<?0/J.7>E:K)GM((':(O!9,$G#M2MQ@/2VWKRI^$O54UF:I_JX6
P&QG\?*S!Q84G%_/S1Q"E^?*\ R'[>IS4H]UZQ AQ!$31N94(!6$Q8W_P[" M/Q/*
PYX!6AE05%>44>4N"YJ\\4'LY4U2,AEK\J"\0$BB*T$J==7TL(1"R+V!Q,DRZTB7O
P>'%S\@)JG8)=LR.="%N_S1I:GF;SI4VXS)0#'L1;H'_\>57.1>V4W(6,\0P=X67;
P46QB&]:+!9^=2[3M,)T7H3H<*NZY48['%K5?[5KLY_=99\Y>4DTG<U\0W?7!E_#=
PD3Y$\T@_\:&I:,G9 P&6=3R00_4AG0.()035 X@'"O?Y@^8&.D"(.7]Q@;0![(RM
P-F-MW2S6UT&&,%[#1$"Q]2WCANQGIT..[8;5JG#>[9L$2XC!:X] ,A"]0#[*KR%1
P'J&Z4?EW\=E0YEE7$GDH<R.YE9:NHHB[Q=YWQ@)(PSW&AI%\/'^KYZ52$4[PR:?J
P[/ZVUD5T)S@Z/QP_O'#-.="7)YGQ".".<4#[[$?N9^U-65,%;<^"RP9>R;("0V/<
P+DNV/@0Q!6V[#0."PCL"JS@7_4W7(7J5L3@>"8NOANKX-IKHK+N8:K38=.XG.%'D
P6[Q0,'A27ID5.N^WW2;7!WXM"AMAH:(<T$99LT9QC?3V%':GEM#OZ 5J/MU:6B/F
P(9TTI3T1HD0\;:,YS V^;0% 4H'#F,,4D:7>)"^NS-QC6WW[ 8W] 5*5""N8T1"%
P7P@/36OF2[F/@4D#<3.S>7RZ12/#2$>HEF(L4#.8:-&?SN8+ C)2-!E/%4F:<#EE
PO C'P_]N%GZX4#JT.PL*W\J/ZG1E4<%"[F ?-1%*[O?*5[X!E^LA%'F1S;GT#==.
P.]M);R*(5TEJK]*&<*(KYX27,@40ARV.6/.M7]#3E=9!]>I<<PSYNDVQW08J,G*2
PA74XU5'F!HKG2V0,FBK#K"O1"\D4 <D[OJ/]9SS%)8JO__4P;R^) @47]_PRSZ'5
P95;$1G0<KK+M6IR+^]TUJN+80LS;W!NL2QWJ%HN/8PU,FZE]:.)K3+&&JY)^8*4,
`endprotected128

////////////////////////////////////////////////////////////////////////////////////////////////////////////


`protected128
PW%6N-7SP_SO_TK,3>DL!DT-1M\7DG![]> 4:6,=?0!8.J\K]2J55I<2N=C=&Z<7U
PF>S#:'*-QNR%<^)6=#&>ZHI_88*_N+!/7M.2$=39I4#70&:ZHM =:WN>')9-LKQI
PD@8I*?XZY!< EE?L\4!8C3'W<"JAKAF,>_R:4BFLPXPM\.++RB(-1 ^+UR/Q>B0&
PY ZSK[S8^TJJZ9G&MN&%)/<%& , Q@IU'RGW^1:J^[H@ZA(37M@$>C(_IVWBSL:@
P6 U2W+'"%@4"Y7[8@P@%A^8!Z4A#IYQ+O\RJW?R)4G4/ NQ\5('(.0TDQ/T)GX7&
PK*4EI(.^NL!?$CI:(YR>:-6.\X9/B(*F 1;P1YLW,NH6M6"0[JRX\_FF&N3./UE!
P5U)7!(*2Y/Z$/BO,++51;14HR86"JKKB,1SC(]<J4I-DV. !.3.CU^79KEE"[1_,
P%XQ0H?W_&BS7"OW]6O[-YD'M8EQYF:D;A2^[B46?[MVA;9)R%QZ0T\6>K/9.%V=X
P9/JF$@%Z1 ?S(8 2]Q,-9LQ!-*@E8[$U_PT5M5.W([/O%4.K>7*'E/]%:;4MSKS4
PDV8S;7LZ)%QNB%Q14>[IGX+HC=8"EP='?77'^S*IK8]@I.)*J@4;TL+U#\3RC$S]
P>5D5IVF7:#SQN$8-]T$%K(\1.=6$-QG7Y?O=^H6&UU?VX9KC92%T]/1OR:*BJCZY
PO[D\N'Y<_?3PC:<4#%<JF1D$T]3=51OH5)C" MC C9CJRAW/+6$!-K$7/KE1RBF-
PZ8S*)F2>6./!9./BE'ZU;MO(3.RE.<\C?Z9 >=!A2(%Y>!M2'^+,1UD'VKF,IVGS
P/@<3W+(T?T7K+Y\M U[[53MJ-7Q]9K@E9+Z4MO*(U<.!D>E/3=#WS#WENU(T57,G
P#<[99CVZQGV%&XX(,TA>Z(N[KE,EUPUUC\+'FA/);:=>"D]#7RZ;AU-8NR((CN)\
PO8XD6C:=D2E>&VC4WP1MQ_B'2C'FG#+?%ABM4<?\+M4A?/PGWV"UD)]V@D,YIYIP
P$154@N*2DY?OZAU[*1JXR$V-,E??LD&:LAS _L@VQ[9R4EJ49Y7;]@5O6;2*K_^H
P0O2@.G&)^]NE%6CGZ6L<6*+3M#&F;S8<>!8ZOK+&2.^-MY<1X=5_7&KTG$ O]+<)
P>UY"(^L@J-@T!L:YO%X.<I0"R[U83\I2TRK$)J)3226BFT>UX'W7UXP?SR]289YC
PP?GTH<'8R)V]F'-Y)&H%PWZ .3>NE>=1#>!-%$ DY$>6JNL.G&QZZSUK6SRB69UR
PXG":6B/\%^+#'7SKS>6PD_=R+<RH\NU3\3^M42W*EWP>]K W])Y)"9H2 *7$G$=]
PR&;X\&GPDH/;)N$C&S&_8577DN-*<GOHC?!T=(++NE<4 T>C94;WC=%_M:KX3HI^
P)5^E*]EHP\_Y703(HHUV%<^)G +/Y!&YCCRJ+1P]<^<KZ*W)EZY.9U1".M[4\C#/
P6%2'^WJL0V..NBN E\+E $NQ"3[[JL3P>T(T98HXU@I$SK%6Y9X3VD6?F7 5#HG;
P @#]ZG[8@3BWEF-^+#F]:D?NE!5RJ L!AHX@KJ\G.JY$$3"OGOSN\Q 3D@L< ZV"
P3GB 1F;/#5)@W?_05<]Y=PZUK/9G2"X]M)S0>+&/N#WU/Z'Q+:P%3/%#1:V@(+'(
P$-M!9T7.0ZDE"IR(L><I^@3ZP:VV2=D,[@T8D=RD8G?@_=[#*V;'! 1LX4E\'A3:
PHVG>D1V5@F@['#X2F# L?1V''5-UBP5\8^;N-5OV3(*OC?,_Q';).*.*_]+A[RKX
PH:O]\Q:JO=#6E 10"U.]MTP\63"70FS8>J($:!P!7TE;R)G\E"A5)'_G1\.UB@ O
P![Y<8.W[DBQ;-RK^#<O EHM*SCB2FBXM[M87X055;LO>EKGR,MERN"TN_5,A%<_G
P3+E) ^SKA0Q8BS#[ %&]1N]I#*'D"-7V,8@D&11?JAP,9,T43C&I70):EVLJE2U&
P+VD0]!4L-7L?O[E0U "???4K)@*U5N#,C"^BLZ.U2LYZ",8E2V=)2I$ S_P3+0IM
P474(9C$XXQ'] $8O_&P"[<J)@TA./&;,I-MB%^T8YES"+%$G?X=F/89Z0Q&[I<4=
PU8[$3H>%A?SH&5'S+VK[JW^-)+[1?H8C_!7 K/],3(K'+=@-[7K<CMT%M@\WKK2=
P-\%4KVJ2V^"%V[A1@$'=6AXR^%>#E5B)PVYSRR3'/OX'_GT+*,IQS%+_J9*W'BT@
P")5/I)X/HI&.O <)UBX!@+#-Y/J :A-FO<'[B"(Q[-,2H904&,:7;G!,&;=R&""&
P[(3JC(A4%BZ4HCJ>%,Z3R)G^=?&=4H>5NL9];_13!VH83V9-+57W':3I,F2,(JN^
PNNW5*:"0&M&9#DV]Z;FW;?&U8'@6JE'D+&'2^LHLM&)&91<*TKP?Y%\*#HKMC.W+
P_?G1%58]F D^12,03ND$SQ^6G"U?MBXJ*"Z'5.-WWG47'P'*C&E[O\X7Z^2?K?R$
PIYB7VR-KWZ8I]$ >7V*T5@4/RZ\JME&OD6))*%@!*2/"3^0H($)_V]N"!W+':$\'
PFX\<ZGT_J,OQE.,KR%EI]*EHH,F2(L!-: !?>))Y5Q)>],G?PN.+>[%P6"K0>P7O
P*U\1<]'R3C 'FF>W8GS9?7?Z'G*#!*[A6^O1B@(I6]H$Z/QV8%;*J$<R'XOG3Q?$
PIK@Z85(;(4^-S]R'#,HWB0'"F,:V"P>[NF+OQ9&[@(2CXGA!D4A1:<AK1T?+:GA4
PR?LVH-F88,G7Q2N;Z7C7D>QR&/P].R40=].D.LXU<GJ(T@CUST4YG&#%OI'NWM]N
P+&1^^ @0'?:R5$U]73,0 Z'$^=;-GD] N D<U+!!JSJ[&#=Z^." ^14!-UA/Z'!#
P<>-5_%%2^BWLSMV9Q4E-E_$;8>9I9V](2.L_Q=0E)HT+]'Z%+F6JPT$&XX4A+3U%
P!527P?N()&1W=U5/T1C3*,MSKP;\"SA$HG49\Q 4J:F!;-VU*<GQ=(0Z^RB*F1>1
`endprotected128

////////////////////////////////////////////////////////////////////////////////////////////////////////////


`protected128
PW%6N-7SP_SO_TK,3>DL!DT-1M\7DG![]> 4:6,=?0!8.J\K]2J55I<2N=C=&Z<7U
PF>S#:'*-QNR%<^)6=#&>ZH9R2*YLR[&9O#;?I2IJ#P.9TE<N[GR)2K]'*?^QF^-"
P8,I8^FMIJ^_@9F-S'J7V U(8OPB2!NN;3I9*RB'[::QN_N:>T[:,-45('[ 1_+XR
PND_''#7[94?>V=N@)0Z20G\!1O$TTC0?K10\P?L4A3N<>]95I((K= Q<[<S*2?SK
P)+/K284(S!=8%*05<01IEHY=&:O87I#U/>,62C=Z@5@$+'XJBN%XTV,,3:#O^(RH
P"\N0,*M*98=Z-$/NF P8A2^<#L9E^34,74('9S&ZSCCD!<_NVVLWFCV:/:<NCNB5
PR&H-L00<^$MVY=KI2E79\\:F'C7!5"7MO((9AFR1!2>I4@Q@&Q_(.6W2*ZV7A1@U
PC="_#3 JV[PLV8(Q3X=,RC]=1-:/])1JUV3ZU$-H=..<^B'DGUM.BEPK+R= SZ['
P?P"0U!CZ*7+9.&1B7Y$REX74'@.1G8@MML)>5?;.40=JS!%<ENXJSL!""29-\_[T
P6T/K1S#5 8KH'W%&9<P%-=1P30!7T6YU%OR&M-NU+![]4E<UF<RD51D%0!2K68BN
P^?>Z.0>G=#B-"UWS[K/0+.]"_ ;T5!"<5A1_L66^&"Z1U#E0Z6KG*VCLE2Y73.M>
P&(T00YA3-*=[N@%R'!VX8NK4YOSMC*R?A<@ZF3U%I@J+?_;]$=BOJIY%VWF <7?T
P3IF*R@A]'DXCE7V-B8)HATNG2 O75=+2?SNHC>.T==$/G1W+$Q&K0+T%I=A@:U=Q
PGLC3='JW<D7+6=X-$0@C_N.^7%N@UHN-C@4)!NU3/_,04(Y'ERP=MVV#T+9% [0$
P3$B61%JF)F1WM0!UB:^!H0V<?E#I4H@ZIP_U^,8/E9O2;N'%:;#2:")BW^;AS*8^
P!E.[T7[CL7'@NWQ7F^=3+>I@>AL&LPR);1=:_4-<FQ^KS1&V1"I=X8>#J50%O&@Z
P.?.!GX*C*:US1BJRA![ARE2%6=)=&YB83J[]\"5V5$0L[4J#I':#QE8NE MO-J"^
P!73;"#^RKFQMA\)M"53[$4<^]50$BO5'<LOPB@T,OAPA4RC5-O8TW<R1D@K"H:GB
P<K7>5YP<(BV'\37[CG56TT!AEU9B@RXCHC?^4XJF$NA&,M ^^#*DZS XASL[!VMZ
P=(K5Q80O:1UF:(^]7P^&520VZO(\_/(*P,H(]/<"H;BDE=9$3H)W0[8JIW4S(,6B
PUH%)T97G2SZ9&^9)$IKDD09B$I<*#^Y2KYBM@&>-&^V+#?$E9D<=CY2TB UJDR/-
PG(#?RO"' T>7^8!F!>K=0FM*Z^J/=$Q94FY6>'=0?63@%*^\+J"@*DF45_HSE::9
P)+FQ-);OBA$[F%1*TO+8<.=Q\L[6$L[ <K@RY-ZIDX)%0ZDU[ L!Z>6XW*_!-@@8
P$%.">] -8C/H[WJ2P@/Q9[\,%$J/J*@&"&X44"##=)_3=MURZ1E,XF27 ^0W=V_7
PN6%O)8MZD"$M,P RWW8?MB,\ZBU!SS+3X+%EI68A1X5%1"V)@5XEB^Q_OB[%(E6$
P)X\%Q/-7>\KZT][!F'"GK'B#G'YT>J?.F3*<U!*"["H\HP,^G&9S>F9@N)^4FMLF
P<\QGCSV _YXA)# (0R4C#<C"5-&5EQO$*+>?59Z3IG%Y[]->:HFC]WM$<@SO<SR2
P,Z4E@XC#4+,K'\Y-H;>4(7>$&DX5*/KWBN<IKX=H!&&WWP<IZ'( L+B*7P(^X6EN
P)QGT<$ADF,*PK!T#>8$O-70!TXAUC@S(VOK+$X.'G0A73/0)GG1W@C 5[5#)*R\M
P4@5V)_0%Z=$50EM.[4O-.7[;AQI^^PB,4,7")GQ&1\LKVP<6GZ5#8%"9P$DCV(JC
PXPZ"-OPZ'66+F"$@+M8B>8:]DF<="N];8^D@#^IV;B0)/,JI'@JLJG?[/S%_Y O^
PT![%8\V=6+JZLG;I#&U':U2[L8[J/SBW)W$Q^<2 X5<R?^(<'$R?Y$%B%0H2[Z%"
P&S9<@(Q$8^6!(./@MKIY!IBS*!2^MSV1%+FKDJ\NQ_DA), G6%UBE%%81\+^;VIA
P!I3.;)M%]$+DV!FC3(HD%>D93M\DH8@BKB^AK#/[&;TJO2&6K_]0YM?:U(_V?-(H
P'DXK)_%;2Q>7JAW)1TX=>"*AH_5K=-[N26)J^9*S5+OA!W+?#F^_\-Y(\RQH+8J 
PW4>_*CS_.KA6QRB.DAJ%RJ-O5!'BW?NCWW]M!*D"[3S_U6[?+,D2RI7''8]@[W[*
PXMJ]4:%)]4/$+YY1NA3I>4J^D'B:TONQB/ 7ELPTB*\GO'Y\3*]C&\[44Z_:>;/(
P+6V6-FR.2WTF%<0$R7!R;HW-,X.YZQ+E/G*?(&.T04_(UN*">RB(&>SH#@=KM.7 
P_B\VYQ=HB[T7-#WDTIFWM'N"1Z!UIC<*@%B/H(J&*,_OL6'Y]'*"]8PA (>>9OTA
P^I.!4OL3.[5"UK=DH+ $-H^F7N!BI@4)H=>#<W( %Z B*&J:SP*C$I\TI?JX1IB1
P>I (LQ2BSX&3U?.*UKBB,>"S5_FL2H.3%N+^Q"W'*) .3R[]'U:G&DM?N8[V,2(K
P+D+/HV+'ZD'%@=9AYN#T%0 %[I=/#?W:.ZW$07\[&\7S7Y-PK;9X(&]7I5_*',U+
P\.YQGL&DV>3B'"T+_>N0F-CQV/CV/W/L<')'MES8(9."-7L_*"EGD955YID!ZXZ?
P84Q'Y\C_9@]F\&13R%FM\TN:(&R"U7\[VKM%[1O+4&8YZX-L?62R]15+WN8<U5OC
P1%RK@G.L-*U6?I\#X(WX*)=K#83Y5%_CL"V4W:-I<P!;(?7]VGGOY+U.P?+E#U3>
PVZP93$=E"ACRE2#J%GH(61,]E:*G\?PX;4/7T/;#+6)X7[!7FR._+4=_Q1_O%2R3
P,V%[OFNA=GP7U7(([16J>_(\I042U<";(ZU9FXR')U>W#"T3+]5B2C"S:%P*Q[BE
P[WW-QC&[T_"!=X/#,0.<T,'FG,="1IVI62?,!O5N$RMY?K\F;TAH=G7TG%'QYH-K
PT6\#>W(F#F-^#&2']LIQ"$.)B-4CBQ7*,XQ-)NBF;@]^ '[RM!+#!E<+872(:)%Z
P^[BEPPA Z[F!<7FA^0(=<?#$Z+LP]IR3B VFC49O.&27R]1^?%_12^ RY.7R'GE&
PZ$<]%*6[N!>44=N4<BUNVBUJR*,>O@T>FTQ]6^($@$^ 7*FWCQ+,?2VS]3WG'9-#
PL^VY3A:KZ9K-B#'CX+^%KO^:A1_P5:@E\2W2[F!35JTM'Y'PR$9H3IL4+&)7+8!D
PRON_7D<CY H?/C:X)RLJN_\[4..3+NM5J0X%$@K!P0HR[5OH'E3MND@8]!O/W%'W
P J6;OV@4F$=XL6V4BO="(ET5(4%@Y2WIU>PO6L0P!R@D"0 ^/P*&?26A:C(?@H!L
P[7-.-Z,#GG"E."7]%(7;@AAYD(+CN3O 4,#'9DU(!=ZQ;T_4YNL'.(R.Y+/3\\F!
P"[P9?*]$&2"%"9>N7S$D@L\64L[?6]^Z>"%<IEC:X-?K+68G&:G=->R?S-;9]7DO
POJ[JSN&_51!6R 6NS25::['WG#ILU1],DB<^]6>.>T;.\1;K@H%3*3?]\QCHF[]4
PFOD3!6L_BAS=48DO$<76 '& -;]7+O>N@[$(&2I&(ZRJ>PHWJ:0VY*,D7#;'BTW\
P@53E%_%'[O!$UX)X#H5KOP1K6C0S^)>T"I]SL3#;9&"V#IQ1\Z#OJ7/^*L2656@;
PHXM>MS,I8V2L<TOKJOKO4Q@^>:GTT%'<++T:7D4]8?1-'](5"KFUX=4QC4^'$M&F
PW)DA4)_5<1+%=VF>6T7Y$ZF>1\9$V<+QE XFR1!%]%FX4#?1IIN!Y=X3>5X_2H@W
PFW>]^5J] :%*XZ/@7B^]CN%#TP#Z'^;U)$"S\:"JZ'0;K5[<%%/+0Q: ;$"E9)E=
P^ AIT;9)I*=:Y81YNMJ&2&*R)0B[#GLV^7RU-:C/7J#%NIUHO"/$"1]=OO<-:"[X
PTM3R7D9.%!D[</AE5/T4VJM(WK"N%U]ZSUT_H/)T++M8!9U7?._BH=VO&L'A6F0'
PY?(Y(F,\E\%833$(C[ 2V2?1<-L_8A_G_+5**!B+RDJ]' MS JM%RZ)9D/T!+_KQ
PI C@ZRYZ+?>9>T>E$'GU2A\=9_37F?Y.TIL-5$7BM%?%^@'3-=A2$!Q$K@3O-EY7
PS>;A3)U'W[\X_*S<74.V[@8WB9&-Y=2S7:X/-"O];"9Q3@&,O)>JP(Y!$=8D%/>R
PHETXH.4.@T O+*B<:=!FV >/FYF__""_M%2^<?_,. >6<>9D[GWN<_&,/@J+JQKX
P\KQ+OJV+F[6U[?_OGK#!VF=<K[GN-.T2UOA2\5;EUE!)S[A*\VZ GE-():U"*-0T
P0!Z+SYT462-N'R:KO321"MRG1UB$(]&IUES*JG#TZWR(V1V_%I^4,R-V&#OM:$.-
P"M8V.KK:GB<([HO'IGW\B.*[DMKB>*5]B!@G;F_.PNHV5"2TM^5G[C3>02N6/XMV
PY#(D^IU;[#1_A!GQM,S8"P#0.\^/&;C/ @\61(N'A<APJEB-[R&V^<3"8!M>IR[X
P/A2#VHTX( WKR"4QZVB=S3;H $V;)\QMF>,-T/93">K HT3*RI@4#?^S<1)?\<A2
P4#+@G9 $U:I2^1DR#F56L#1OWVQY_R!OP[08.Q"!=ELF,_Q*47%-6;:DA(_8J$<C
PEP]N(6J&NCJF[#:+MZ-X9[_1$W W^[N :[0QB2\1VE+@Z_-!)G4P*0*<_/>4(N]+
P[X[[C".F"E%48?3P_*+:&UT>;KW3VG+;X_-,;Y6^D3=8?^&0"@CDV<#Z;=OC"R\C
`endprotected128

////////////////////////////////////////////////////////////////////////////////////////////////////////////


`protected128
PW%6N-7SP_SO_TK,3>DL!DT-1M\7DG![]> 4:6,=?0!8.J\K]2J55I<2N=C=&Z<7U
PF>S#:'*-QNR%<^)6=#&>ZJ&AFN_C&J5A/56B++R;YT T]Y/VCZK6\QPIZ?H"RQ!\
P!5*R6\(,5/5YV_LH7!. 9=4=8J1UN^2[!SNM64421FK\RGN^<_]'L&=L"RVB<_9R
P?FF.+Z@A.:,2XNG@"8Z (9M$O-0S$TOW^J1MR]' VBU1^BCT*]8_'MPRBJ!XUM2I
P&A/ 4.,RLP 0A4G;2SM-I4;X6G3ZC52!K]J+:(>Y6&BE2AP;B))=O,^+LC@.5I(N
PZ VLA$?#^IS<#4T5_P@-7PB\2C/;U8D6&=UT"U&:LZV*B7:_-$E=RYM12)R&C;2N
P\?J!$MP+,E94*F>50,XM%R^#-A6<;\O]Z":NGJ5(S++WW2MA9SCXZT*C"[A?FE-_
PKME31-+5G;J"/F6JY"DE]D"?&!+]]AN1[=:GJ-0O>:>_+! #)KG:=\_GT<YC$>/%
PF8G0PFESQA_0TH$4TZ59GR7V1&-7>'"_H/MC?D9$,E _GC?+UNPT5Y>=FTBVM-WE
P;L%YF#I.#'95BG^;FT? ROVX%O&TZ9D-*2W='D@%J$VRP[06MZKY-Z+!$ +AOO.E
P2AW-;0W&W?<;+*Q2%$#I )*6G),?Z3025K,+M59RN2L41?BV"\+UY#H/-Y,<F6PQ
P YN*?RU(]E 9%N6%C\<O]P\J_CX\"Y%+<M_6%$[B*,U:+\1C]H2D=VF N(8R:MT1
P?1:6CB?-(XJ\:<>F/!**\AA%V"?.+S0XO  '#O6$<@(A_/++@Y_B1J%#PS"UR>7I
PVGYKRZ&J[6ZRJ$PWL.$JK@<M6L.84["PS=S(+@!$>>=V3WVMV-]&T&XU=Q<WD+$Y
P%@$QBZ@B.*UTOY#E;"5T,0W-PX\_! =W0* FB@OL]')R<WG%' J=%_ AC,\]A(_\
PI#OY*0+!BZ,X:1?I#,D<V5@IN#C@W,0W>+&R9IV^&Y7RO%Q_7?2B-V_EBPW^=\O-
PZ^?Q]=,F\KM8G%705)3ZB+M%:(AMF=K@\#1%EOH4YY4(S\P;'S=US)8QZE<6>C,N
PV7R=F8#.G@I@S$A'!,>"_.CED23M49&.].!93$5[/W$CJ0) S'.XPURJ?;4W[@("
PO.-U(Z?/U40'>3@%.> GISP<XD.@#>R#LXV%;U/X%4BXSLZD/SL@J<OJ6FQ0OVGT
P*!7B/'?0[Z04Y%LA?JKLH]RL-]YY O*3_>R]P@ZI/$X%9-L]0TW1\\A&6(.0YO"+
PS91BAY#8^6<WXC(>()(\X,<BU'(A"LVAT+B[.35"&\/!R"NVPH"@VJ_ZO">9L1,V
PZ=I$:T@<1/.1*!&<Z^V2<5@%P^F]QD!_8:G-,UMP57<(UI!46/%Z&:6CS#!A7;=N
P43Y&GQ,I@'UF"?RF>R,#R5E.J^(35/OWG]2U^M$.RB2<-_1O#.1;QQ-UJ[3.ZD#>
PL#0];"Y^@A[W+AS?CLE+W^.J4E>=+@1#A&V61:P8XS?XS;8(T"I?&"S26N.?&P#8
P_D=@,&($W3VW*33L??3NXYJ>WSJZCM\/,W]83I([Z8!L+M](6]I;$6BI[!2:\M+9
P]T.564D]LU="/43/81%F([(\\K$OM]=GXKBI42 ^J7<X<&&!(W5.\M_T2!6;7E[3
`endprotected128

////////////////////////////////////////////////////////////////////////////////////////////////////////////


`protected128
PW%6N-7SP_SO_TK,3>DL!DT-1M\7DG![]> 4:6,=?0!8.J\K]2J55I<2N=C=&Z<7U
PF>S#:'*-QNR%<^)6=#&>ZH9R2*YLR[&9O#;?I2IJ#P.9TE<N[GR)2K]'*?^QF^-"
P8,I8^FMIJ^_@9F-S'J7V U(8OPB2!NN;3I9*RB'[::RIW1SR7Z[YP@$%XJ+HF8SX
P*]'O/*H'R-7@^(:N^43)*>;)CR7)INUA?\?%\]K20U3*U=<LXDP+X#NRS751DV+1
P9>J[KY1+5NR@/_=YGDUA+TS<S^2BQ?,>,H2%MG^_])P6ZKL  .CR#4A: (,[C11C
PVK%VBZJ&[)WH=-0\YGJ@R@N>!4$I> ZCTEU01QU+'CW?9(="Z-5.I? &\B>7"$TR
PH$<(PX<3[$>=X@ UA9X;'YI 9,JZ%SZ]=[R)_K?]#31.= H#2<.AD5%/_)QF0@RA
P+P];;[#H6EV%SW.C);W$(^PE)%$1OV^LH:Z]%[8?OK &CMS@BXR".^_.5-6$4N6&
PAU96FPF&FCRC/R=3H_V0JL75F,%88S.>Q4*]7T^(R)"<*.V1UM]UR5I,LLZ3:.N]
P\:=EVK39^.]YR] _LIU-1RA-.CDN<@<FP-AXI<@G]_W,^=8J:0KB1$\!&TN5$L;?
P!O):EMMNTOAG;$XETSSY=GPG[[/Z:&;4_VQA07L4TE/$0Y01$4P#=/N2/4O/M)X$
PXOA_@AZ'_7D+Z?.D4A$WP34"=JH8._9?=QE1,Z9P7*EB7TRI*LFGX#P[?[AY%%^X
PA/M81[TH6?T<P^VA?I,NOH/W]JEN'U!/N(<+2@IM@S.D&NOMOQ]?=<<2)C6%6VC\
P? TC1,)03SZ5DQAF(,IDOV*ICWFVTP1EY@M\&?J!+7$;_I*[\!R7PJ9"*=<L0WD7
P&*3G=-]SHI4O$#S*NL#7@'<.521-RPB!!QC!/.8Q:^%-6ENC65"6.!-;'E!]RJB!
P>5-R=^W$-3]F;J<S.4CLI% NQ9](A]>\KC3U.:H[ 84]8!*;-'JE_R'9;V+YFR]/
P:H<]H7J<PX ^EQU#T?9,N5*X?O:!4>&V;GT!^%+O%S(Q3^=3%0ETKE]Y5>13MSJO
P# +_C/"J^?J+>7F::)'/VF%WI"SLN8^YE@;;)*&I+SW4F?P"_61]EFE"JA>6DWK$
P \YE85-,%@L# [>O,KM.6,4#VT(3S-YPW"K:2$@*>XYP;NJFZCF>RY47^#R!MQL,
PDLZ1P5C+T\![]U1\S)4CH$(<1>C-TN6<:Y3?A78)JQL9XF3']3+CO3#1$'#\TY*0
P4,^AHKB=SFQULQ;?>RVPSW)+6<BBY/$K5]_07^95"+2 8J(,FXN2=#N^JP?[)6+'
P1EF_5=&=X].)3A'P)CUE7HJQ5J:.IT_#HZC<+,-G!QU:7?@/]9*#K L"./44O"\D
P)\1#M"^4YE,S&*-.U7\(DHZLD62.$0#/@RU>ECY2V)'E;'X0H@V$:55B)P>"&O7.
PZQ"?>3Y1IRK5G2!@&LO+-*FJM#$W#QQY4\]$8G3 0H%CE@5N6MN3WOQ!JB#@LU#;
PDF]MB3T K\/6_;<FF>3.SN(6^$KJV'YPGDIURUF2;4FA"GY@-*S$6C\WY>::>*2X
P3-JA98.;IUI>3HO3$;R3CD,R<#N0$!^4;C,:-_5;W*WDV,=+X!D?P3(T'.SO!XTB
P^7F5W&I6=SAQA?7][Q7,&I,?2.]X$Y_G-0L4/#YM1I4K*\/+P_)P 6&>.=Q%(,GO
P_E:R%C0Q!H'N^9^)N\\ OG*P5#<B'<TOB<?HPR\JDZK56T0RF]K*D9I#RQ;%Q2<1
P("GG&@T>/IZ>M-&YAMZ.C2G(P:+?17BVO":[#>5$Z#*(QPR)E 0QZ5B'G63!&+0)
P0OB:R8(1^_+RI_WDOCBME0(S)3+&?"<Z(R"X:X#@2LR':]W-DDI[C^V,(/4['('0
P/F^Z5E_T0P"%;P]"??ZV$QR4<I I=89ITK-0 4G'L[YFO'_3M6MKDK)T5N&6=-61
PL+O,$J"?9MY2D2O<^VZL9H#D[,KP8<>0&=@]6]>C;::50-M9H:BF-]7Z?W[2:NX\
PB*3H7O%>$[SM4,0M7SMQL.T>GZH5! IX3N?8+W*_%V51'DH_FEF>V1N#$D;:0TC3
P99%"6%M7JXKW.^S=/K_%_QRQ,5;996CR/I=$0L^G*U2FI[\D@5BSRNR_2185FG\K
PW>*90$B\,1=$[!=WT3-4>1X3)OZ&/^J@#0FV4[\ HQR&WWUI+!B+?&OX<(/8@B8(
PTAB1@*4:VDV!35:(N0?6D"/.X^4TCQ8@EO^W%K0_ '@6F+T!!</I3CIPP9X<FSB5
P:\'_F:")8")L(Q];]9P-8FJ_$:Z,@$+2A;>)I^XXY=1<K)Y]B'@R&VL4"V5,=F4K
P>K4E^QCE=S7@PXPH"\]D!3O,\G72*N'*P;Z 6K773Q<1LM83E?-_8!1U\'&WGZ 5
P]"XRSB5P-K-)*VUQ7ZEE4N1H=Y<8Y;$W7"$"9,EA.A 53HDF.8'NX$Y3JRVT2(Y,
P!N ;PL:I:6?:L4EXH7V&,;G 3F[/OV[U%0.V4_%XIQ 5&9.^OS(QQ6X\8'"<TPD>
PADX">%R=F^D*(-)6N_S:%X98]O2@,A_?+[/'&75\%USWC_@5Y+R'OV>>CE)/%&?Y
P[]6:B\P_W6N'Y^#>+M!R/TI16<DUU&X2]<49H_O.C<WO^EI#B]^(DC6!Y#M<SM*F
P&Z_63B%+G>3V)GNFP:9X$@/8.$'&=(*QV^Q0>FU_I$8F^%1REM=WK4WSHR(T\:W=
PPBH<S#&4*N0<-DC%$=X5:@NYQ$.\T8LO6*U(+/#(CL$*G1;@\$]S(ZZ,:*IA'L-@
P'NJA2>J>PD\)3AQZ)#E"+<[55G#MMEH ]&RL;3F.KYPX:*LB7$7XKXD>L6(7*^?G
PV]=ZNB7*QLX"R&CBG?4>B,$DRWID3\A4^,W%T5G5<NOT1NVW^\UT]*@+-0 =:%))
PF#:V5A-V M?@)U^8):ZTM6R4:MG+=#N"MCX]4./,IC?3'*1NKL*PR./?]AL$TVD=
P?Y3,Z_:N7&GM*'/,KI&4G3/:_?<),6,&W>YP9]3]/#B@"PZJIV4%:*KWYTE\[M*%
P<7=>U>+$7Z0MR?B!UCSQ_L94-$J"360QTI+HJ#IK;?8)E^Y+*F[M8C3^"YB3-CS@
P(*V3PYI(+T7BR6&6RX)+L3QR7+CO_6>V7:#L)QK1%)?:Z";_+UD0LO_+"N57#DQ(
PYQS[I;-VDK#-+YV>WH<E2X4NX=[(K#@)IDMV/"E7I?\<S>?]FBUE@B/Y$Z3&Q3]^
P>,+_XEP=(U1KCMVMVAL>K1YZ5[VR*CYE>NPS9'(RH/'9ASPD[QH*X\&8]^A7 O= 
P:+UE@B@Q[;>H[6:34"<'5E]VJ^AFF*7574SQ2K)&>9:1H$]BAPF#X*GG,F0G 8C?
P,I<>'"-DC<" ,DE%B6A?X#RSK63@W8-HF%W.JIO6/X!?WR/R0H)K2X# S[/-9;YF
P++'?+@,(\':RN#SO%$NRJ9HR2AXYA &<M<3,<,;_QG_?R['('H3<T8"R@J!^R\>%
PD-^O[TP&BD)/VU4";.?\7];Q'!"#OM]'*V1E.48\207X88X?Z>6P)9^S08I&A)5"
PC;OQ>N-!!Q>15FA!<UUY8]!(?(X2*LG]GO>0^Q%S:P$Z6-NOZL).3P3 5$Q7"!0X
PT0Z6:0WLB/@/ZV5CDU01LN_J4_5W:)G(0OY3&RY(JQ.A&->ZE3-*+E',MK)'V!2B
P[T?6(MY:;W=A$E\=OV#49*?^7X\1%5&,3<RR)]IJFM]K\J=N/6:O!%1SJZYGIU&H
P; 'A%A4)*C0^YI"+:Z,+1&!J=/YW+EI<IR^?HTR&M%"(D#_)[]QV+'%_<!E?GI8>
PV_^V%/#YY@O^DR(W;EZ,]D!DW!MHMF-LVP]X*VB7G.<7/,Z)T=7PX\ILSY)6^_Y)
P>4T2>*+ "^HTV3:V"4)U&%NS:@R]RB%=#0X_1V SK2F,Q[F>J\:3Z>WC:L ]C,)*
P),<#6H^98!):SI]41L@A"!XU,[EZ6X@I@Z&I\(#-W,=GK/JZF^$SI?R_ C;R/Q\<
PHWZ=;UF%*'^2[+W.L2\87\B_AX\:6);Z23='$EFNA^IGXBX]%]^#WGD68FU[?%%U
P,2D-M3.U"3]NCCZ*FO;4_6%+?;TY>+W[4O_'!<<Q^VT_L8:49S^(G4K\.77A(X=U
P?7]<W_E(Q[S(ORS;MR^*DBQ0(55[^M_7@=;'#3C>%*P9@EG2+T& +"%:@@"E06)R
P4PTL\]2S-%P=1P<_A7<AF"]8@ZRGN,"&0]?ZUL_@9#BG>"[%G5@=;8*AZH>;V3P%
P^A%Q"S84?;VRP9"VVL'I\[ NVG;?@/+]$I 8$3H,P,'X>D4HBZU=CZ4Y'&\%=L;+
P\V(=H=P$HM&8H2>N1U1..61^;;$RP2Q_H-"),[0/<QM*57DY). DKH *5T3'G[/Y
PXH>L>E[8(F[J_&D4>^.EK0B&4S%-Y>%?Y/[XI:0AJ,T&0WG!*3+H(S43^5$K-F V
P&&_]?^*CK$0ZL2?SL__\)6N=!>.]PF9NWGCB-3QH(W=O]<KD$\L&EX(;BF)D9/#-
P4LFK1O0R4%H?)$?_(B,_1F2DCX1'[^I.9V97;F"%5R.N/VL;0!;,U9Z],I7'Y9CF
P<^6")+LL'JOU;H64U/2?N/*2F*L=@ED\+5F$,O<[AANI1;4Q:W8?P_"HHOT\.=+)
PSK"M_)]]G4&#M:VI8AB2U#&-%ODJVA1)0#6M'-B-:?8VA66D%]@:4,(+.%PCE&=Z
P4%62SXTRS^5^> I&CV8]A)T@^ ?,3=MCCG"/[FCM)7!3XK+?J3P_7QD"AWAR5Y)]
P@/"3K*0"]J=4++4#$D6.GE\RN$F-_;A_C\%Q!8OH)E JSY_B;UNS@NU#H!KJ%0_C
P$SEY*00FL9399]B_U29#,I<1\'P8+8&=,A-B4N!,E_IC"DMYUSDH4KU;Z_0>ON13
P(W9_]2<A] KQCRIAXQ*IGEQ^;3F&.R&/U>NAO^HXHDR:E'7Z,C#2&4H?]E.9!MC.
PNL5PLF4L501J[XQ? IEZ_A$UAPVI+L&Z4E9TNB8]"QSTR(3IF"YMZ.,H@"U6)E&&
PO<O#+*!^W6]$NS)<9DL(A>IK0!O?-4\/Y1GID@WC4M&:++UB#I=\?B8,'/$G_[HK
P]>=LE3?B (G) 8\><;)K+O&J]$"B27>55W=FE1/9\N<UFGAQWGTB@X<HY!BJV%>,
P@',A!](ND0]O*?%9T9@GKZDV6XV+P:=XE08 =B;L^0Y']TK\LN3T.1M=>X#"@Z5X
`endprotected128

////////////////////////////////////////////////////////////////////////////////////////////////////////////


`protected128
PW%6N-7SP_SO_TK,3>DL!DT-1M\7DG![]> 4:6,=?0!8.J\K]2J55I<2N=C=&Z<7U
PF>S#:'*-QNR%<^)6=#&>ZH9R2*YLR[&9O#;?I2IJ#P.9TE<N[GR)2K]'*?^QF^-"
P8,I8^FMIJ^_@9F-S'J7V U(8OPB2!NN;3I9*RB'[::RLK,\JXR#>P-.O5ZI(<*)9
PWR74S#9F+YC!C4DA:$14AW>>*.GWZ9X_S%?0LMB0Q&!X5,-+QJ&I% !2")N-!%^ 
PNYBK*B!,0\>@9 CT(J)9W,GKSFU9,F%[(]1_J""U29R6]+<[=(+#@0CNJO2G^S:\
PJQ?5<7^GQR\\7NRA)</9<=,NK6C\:$:;E\0-7D (63!>27@$BI5?C4'AYJ^<E9CA
P(D!M\Q+4$9 %AL&O$[I2I-OJ(2\!'[6_W,QE&0B8"*KMLJV5VED#RX<7H=C2."^W
PU,Z3"+<$[TS?A;*RG\R6N70LH+:%G,.@@(]E=$J<O("NIO.(>/JI_RN$T$6Z^"Q!
PK,W6*,&#?PWH?0J>'):5F(.MUS[>$]!H\YZV*ZZ@2E:A@@6Y]CVLJ98U;?\2W.,.
PO,CGN\0^]?  *Y5+_"(;)PQ6:#4E$6];#A4EP768Q]0Y]G#A(O89+0+)DK=1XQ=S
P/U^<;$ +W#SJ+*S)]9A$:G69]<^&!P,W2?@L2:X#@46T4*&($2KK%DOJ,6M\YBKI
P@$GC*V=VO</:S5:W]V)'0KHQ0/YH:4'!\9MU"'4PM;56E<RV>9%:F'@&6<'E&%>$
PN> =,+$E?&L A-JOO?1RJAP673ID69/V[$M@B4.\YV)WAH+6LC?2F$A@EL$^L9,#
PET\$BXR4$R.7*&Y$P<^;6HSSK192JR\&4*1'8JH)&J/I'EO3/0O6Y,J7][WE&JI 
P <J=9N$6C_/J/7U#(U1J.T<S)$&0'#**>ODJW(:73"N7+:0Q^H2,,<<835Z%.<S7
P1?Y<A<I64TG/H)-'$M;67[0NW7L(_4VTB&:E["PP4/\O]._NWR<M.YREA0+53Q<#
P*BH_'+;Z/3\3"5&TM*0?O5/&OF$6SNB=V[1C^;9/VHM\*E[YCTPBA[C&$M8[.,#D
P%5K&.%X,A/].TZU4M;WR.X(=^4(VDHL!&P.5J*;GF9 45& ^+%-$[T%%@%R)(VI0
PDZ=PRL*H0SC(*=*T3^(8TSLH_?S7_2KQ<L[D:4\J[%DB.0-_THR^1DXCE^?!0E1V
PMY>LJH>2WCQHETAK'P@J#KW]-5PG9OGOTTF,2SP55;1JD4DK+;G5U+: "./PB7V8
PZ :!-ZB>V[LW?FQP3K:B_DU6X@EF.Z0?W3*2?ZI6MLQ<:!#0WEZSE:Y 1!1@CM*0
P;(/\XQQ^*I6QG\MS*D]U??N>>]J8196GJU1X$,@-ZM9Y;V?,"! W'#=B'"XJY,AI
P:1#O HMY<UOSW+Q(S]1OV?^-J17(5"?GVA,YP%Q"LS$O7A2=P [F4@T./9<NS6V&
P+X'4@/^"NC;@?1YY9VYN"DZ'&)==FE^)C(K@A]K-]L WZOR-7"U(O!8I/FV()9CB
P.,@F[C!RW+^DP#'R(8)-XT21C4VG%)=UNLQ6ET%EF'$,*Y+XI:0".]<G"UQJ&[LT
P=PI=S)-@9P#1D=KIF!=N^Y4<Z5WS\;"HL6CHJ_F(67LVIG92MJS@,RTW $=585-*
PGWI);?68>'>CW(K#N*ANFJ)T,H ,>6M3H OIZB<8YV4@I+D "WC,!/B'M]VIO;:[
P[D X2*KR*96,<[8=]6*$KD9@=771U-J'O!2P!2E*CF1.AX%#Z:AM1)39CN*FX?0;
PM["%O_;6Y[UPZYBT F4TDLF[HR"8*049<&-V]8A57C<TC7\;)O<#$KJA:U>1Z <Z
P_63="GDI#&5I&O@FC=D#Z&9G!]7T54XDHXU]9%KR61.5R7WV/LS,:(6E7D"EJ5Z8
P5<I@DH#]V,JJ\L"\?S$U^9D#IL%YR/5Y+^>AJP%='_K^2OHA_>D0\\*!&VAWU=[X
P1NQDT,\!Y2WDCRM9(KJ'@F8U9B6)V)7_V*[HB3':P>J6.Q05O4@SSZ]0Q]!4TVK;
PZ$^6>*X:E4EOZ/)J#V@7/\(_+WDK4'L/E-;_ 1F/1Q/$-E[E0',LFCWYN()SG10#
P"8OD'.-)]Q8@<@A%G7.W=Z40?+CDQ1S$1]%PAR^#,5BVEX?F[L*2F4N]7,NT%\W'
`endprotected128

////////////////////////////////////////////////////////////////////////////////////////////////////////////


`protected128
PNV'1>,0;%GI:;0X(%41WOFORDK9R#+1*>>CJM^55G/+4W?PE D_54W6?8@B'6WH5
PNZPY:,HC8VI B%_I?%H*,G4$BR"VCTB6>0X, ^MNZ$O:W-MFJ!%AS#3Z8;-&*]$A
P96$6]S[)=] 2L4XP>QEDA,*!UB*<OJT<7&$%/K*L+_ 7ONNLG42B_VQPJV0]]*M@
P:*HK>U#KTY'<"EY=L)U:41.9'W2+T95# 0XNU$7D)A#WCX-EDH2!@H80=<">' U4
PM!+X)79?"8 P)W<+<ZT*3'%8W@M+OC'OZ<3W\V7;]?I:,F4]H ,A'E-LN>(>T;C8
P==H_]+N$-$4Q46%E8\=*EY9WV_/1(\$/.]\-X!ZOVLS'ABJ5[[FT,+IH8[SC<+-@
P[(5L*%(J>"T>/HD#D$H59H1P"%PT,4E=F@4K>U1Q0'HH[UP&T1RTF(@/A>J3[(8+
P>L,OU'=6&8 QJOZ7;AJH"Q"$G.HUA&KA^SR8&C5N5?R'8 H?5"=Y:+OOY/"@W:_)
P;#I]JCAV^NSPH8Y)/P$F>_RGQ)VL6R'@DN3]6[]@^"T5@/):HW%)89+79.^9;+G^
P^3T:2?E0^E*"-657$DVIB*;SOV3L/ZE2:9>#5$[ :Y5P+$U#]CZ\FFDJ9\C>3C>5
P>8GJ51DT%^X*(?7U<==-5AJC^KJ2&\+; N,;8^O^QBDU=D?.+3S?&1_3R6;+?/UL
P3=KI;(E^7?(VA7A";78RLWP3@!FUD+O@CF]M[LJ/PN&H]P5\"C5J:_D(M)G7BL4@
PP3/P")'OWO*AN\$)"5"J76+'P0"V!__*&G25+>/GSLCE_R]Q/ -S72RO(S N!7 ]
PB5H"6^F1']#&O7_5UPO# VZ:ZVMTB5.GN(C]099KKI\P0QD:]9*:5 %>*I;X=\55
PS2@*Z;.MO*\(>?S+]USKGO,U1=?>"21P$1*&,%\^B$J5MI;OPCU=B\V-(% $@EY5
PS!<<9Y(?!AE?$"1<#$7)/%\Y0+'-X=LW[2Q5;@#:I4F7L'F4'H^_C/,3B#YNDP3G
P[0 ]/C!7\Z0U;6!16+.LJ2FG-U88I.SJ"W_7@)3[S%*WZ6IS7F6B,&?MN($5O>A.
PC!/OE"1"(F+.W66K!'(^CUHGI&O/0HB;A2C0CNL!:+4<BD:2D<HP(XD_6)F L^-&
P,?R(KL4GZ!F'%; B/\.WK[:C]O7O[S)@4+M-OG^746!)X,K]R--4M+^H\?+S'.*(
P:QZW\#F.1F\8JU9K]E87=EQ:>VPB "K(4[=1)K(AC *\_+]]&YVC<Y7Z7,/P0W7Y
P?,A&QW5W$N&XCGFR5! GZZ(Z<G*^PW%)"(Z=4<)#[3/:>5(1%W#_659([8].*<.0
PN4EH-J@F1&0=$^3)LQWS'=?$C)E07+ E?GW1.S2(@:!H1F++ZZ-GH^22 8KW<.]5
PW?+,S,C)JE>Y4,!>P[E3VD:BOQQVIA;5AO<E):<N627@S1=+EFLN6O?AV?IYT&5#
PKXYN#4S6.@[4[$Z'.:,Y5844$!WI B,1N_H\ I<NO:.PM(Y2666^-<B=VPOS;9XX
P"ENU>X0;@.6&^*8QP*8 3"<-H<3J1CA->OY]2V=)+&FG+ ,,$(4D9K'4#Q(SF$M8
P42Y4[#K@-CM((E5ZLU87EMM-\MT3T@W-C[X+?07S(PX9ZY ((J^[UKYG/#ZK$5.0
P<"P<"N=B$E[@TB[^Y/>&--^!2]$/_,(4!W,1WR$Q&9-(/REYM9[R:C<U/SR3%_,"
P]'K#9L]*/IB@_16Y@"44>Y6X+2'Q0'/6UF&$RZ4DV+E3K72YG2;/G?RR@*\)-YEI
P8,GTK_/-L!IKWF[1:A< ]?$E?5JZXG=F#0]S7&!=.$DT)MS4H=IAEJ^^Z+412L(;
PKL)9,)Y>0Z#[ZNY'\[N'-C(/HIL@[R86RCX4+D-TJ)I*- "?W(F5@F7T1BNRF;4,
P%6=M=TEZX*S\U/$VPDP:NP^3LWZ5/[+C^J7$3"HO$H?92[3BFP&:Z[8:3/GW755(
PB2?/*!RN#;9XHJ13)L(/**HN=)3J2?ZK$7\3='WIYL3U./(K*0(!VI3^(:N'"6T5
PK@A*R-FT:;2':8N!X2ZZ3=YTUUGS!=5RU;T!\]DNW4F]&(YG]@#91!6@XV.5M=C%
PBG70TL-V.Y(@M;X'1BWK(DM;/!7T/J"/G&J&"8PQ.;>-A%H)8  8Q,H#GAB2@.&/
PA4K+4H'(S!TM1,0 2+8A61D(,/VS\,U]69LL GZPQRDY\W*QS]]?D7UX9^EQ5.+N
P+J%8*IP>R3> WED6YM@6A(8M.8]BL;*])!@]845X%^6.HN^J)"A(*\JK D6J9+5G
P+I+TJO1\.&N'3.9? B3=>#E@-W]*W(972@L])W%'T_N_DYTD6!@PI]1MB3/?!RU:
P+$P-Z+$5O"2 @3?X&FQ]ZA5Q'?:&YF&EH($;X5BA8ZWK;&+5JSP;DOV57?W2N1UG
P/@D=_BQ?MY@S\Y5]3A/Z5HC,5C8@ "=7JN:IN$<G^MDH9%L+V1*M(+KIX5X2)0G5
P]#SH*)<\1:X8 E@_WQJ9U(,T,*!&A\^-#UC@</''"\W)[[S+^S'W<JF5;V Q$4]A
PY>QQ@=!GU0,+K9/:%U].!3UF)3N4RKQ%XRLS.I92S#>SC.TN<<!9<9HBNR2<-M-A
P0M5671I.6L7VM#+W<0+L DM,:LG[;5BX"%LBYP3/' @#_ S"*^Y^)IM /=K3 GX<
PTY:/<1,TPYUZ??=P1K!,?5A6.MCZ,H8%/K16DQ(YR02<DA?^S:4'P%.ZP':^RZ=+
PMMGX;R1/0N(<E.! OBW&[XGIP[U=M*XKZJ\IP&2M^[4J-<O]&'C_*_<;7IV)^#CG
PX^M<'1.-7A]DU8<L<W8#+L4!/%J85":I(2&QWI(C++I5\R%_/ O0H7+5'L#E-"=T
PEVI&RZ"YB*)\S.;BM_63E'H@4H3"T(S^0^P9F^>/DT_66(L7@^NMD%NO$[Y&-%ME
P(Y7$+RK)JJ'7<KP!$1[BJ3FOLX2:&(.\8\Q2&8TH<AS<-W2+70S)J82QJJ3O3<7\
PZL*F?88;6Y  Y#W!OKTL0F5"JV%!T0VG5*PI,9Z!9]W-#^&(A;R'QL-=W#_I:/PO
P-?>D67GW6(>B ;H7NEZM@56&<"D>J1?D5!GC!O.=W:]]P@F_HALRZ8,9_(@7GY&A
PU8E#<W]4H(:7DMKX9FQQ'>":"B;X*W10XV8C8EK!K? 34=Y/:AR/3#-8&CIOA1R6
P6X\<HSBJ-RZOG/1(04* *77I(R/C<?,C1[=#<$ ?A"T/<:_?]>_VZ(N_]FYR@'1;
P4RM)+&50^IERP>-^D:F M>M 92BH<M9&><8$2VI7?%5B=BUCHT[?( (M0S)FP=\W
PL>J_KIF].>)] \IU2C!(W"NVFLYCP<_G?BMS^S&5?1OJ(T44$&TC/XO4JKX; S.=
P0P(*HS+:O@/4Y\_PC#IF+J-%R8T!#" <>ZN1=*!FG']<XZQOC^>1ESS:]*=,<+P*
P%/L+;S,D88M.V.4P"30M?F=#"?%5>2AJFKJJCUO:X^ (C D]F:QG?)CLY;RP;G_R
PH$WM2*WN,.3H5C=@RYI$57C8CA9WZ*%Y3!VL#)2:4,<SX>2,(#_#T7_F@%9M-5=C
P%(&Q5,\7SGF^1@2?C./ ]E?+-LY=&?^0)?25NKFLP4Z5#QZEQ0\LNXQX$/69IY2M
P$'L\8WK_:Q^.QK)NPV#("IC(AZH"!KLI%()8;HS<GQLCPQP?1^Y%1)7K,IOU/7PD
PD6U[>'7M02BV#EXWTIHH"YSA2/Q9Z$8\[&V%8]>O>+_RC SA-I%S (,A'T9^>/9(
P?P-K*53+Q(!--C%[4;FD3"RR(1TCC/O(&RM"EI*Y,JS+"O1*_6'2GYW3J[.9\C'F
P@BZ]YDI(I<=4=W&)#/( D/H%;9Y64&1R9(,!%>_VUZB6Y)P(=(LA:ZF:4*+29 O.
PX$-+HO.TJ1.40,0#(];?V@4>7-P74_B?<SB!4YC@C_ (SCH LW89#:U#/QXN4Z8"
PFE^C+L^6]1$K<*#52?W:L;*5&UVJA,WL80UNV!\[CR8D?T^-T-#K^6'>DT2NM+H>
PJC@[211!E>)R$)#PJ*XJR0K 4.A'0J2=/4A4]93%6XK[) 0Q$%P<U!'>OK85TRD3
PT.; U98_%DI92,4% :*76X9JRVXEMJ>9O%B?!3$I']F2M^#>8+C[Z4*W&O@#L1_F
P$<:\_GE_DP C/OH^))!;H*B:&;5*K@2I7*QIRA[EJ] L([VRZI+H%^XB7EXZ?^+R
PG<J?J/6PS)MQN:]L[4+,>>BKGPJ3C'4RGXN;278Q5QOM568*(!X5T+K[G^Z6Q[YK
PZW[K3&5Y(@E:T^V$.O!H<X.@V0N^LWD<CEE);J+;+&DQ"=[W M3,>=:];A4H4>QW
PHG(O#CF>:N(K<79/#)PJ8QU&+5,,,U\/(Y(H?IW$%&9,RX04VK\8T9% DO"*2+-N
P'_380:($1VCZ>L&8@ZA,)/1'-JJZAU%HJZ.G:#<LYG#T*?U6$@OM@@[%X,. !%",
P+SSP(';A==RP]# SYIG>2?/0]B>B<3K!4AL3[)"X$Q]I$0.3E#ROO!9LR14>6]RC
PH#\2K[%Y;<[H.R?#1>T$M6).H(27&PA2^2Q2F"VK,&Q#N2(Z<!G70=5@$BQLKX;M
PRZ",7A1KQ4*(6 8KU8&T4DRS.&VRS(LNONJ1%$K-LV4YLM*U\'K/HUT? E#)<X2'
P:,[MS!:+K5I,HL05.5V).8@Y[J(GU)-[F:BC?845;JBL]GHN+HZ86K/BMJ,R3="P
P!1-C-+XSM9D%WR(9T%TV,R1RRU7Z/+R7<OX<D.+$DK-2N$BQS[,\@(G;!4Z![1C=
P[<_9&*'#I%/^RN:8+)<LV25H75'&!7?%!N8H\;J6;$C]C=<>19"F&8$!&2/YN X[
PO:^5T0#+2CUT65G&YXI(XJD^)!5AW51F2L;\6O5>\?6>=CQ>[SN"6^D.0+;:!T#I
PL$E&(F0:L)GNN.I664#TH6_F_B<(1F?S)993Q/'8!TY'4A[+=5O^&FHA-W$<QSW!
PR,'5:5P^HW5D>!W3"Q7J'!G%\1B,'(P902#2:SD*1\M!4YPV:LI%KB=\V" ^ C>5
P^?80_W8Z 3(1&,"-TQ]64+Z(?B;7C\4DWREQ$4WVKYL</^'<S^3 S)!ZSY!OW54 
P2*+&$@'Y C>!>R"OL%LK^OC'+@ZY_C8:8-[UJ,9%T:PA_0AN@EO 0%I];9#=WRA.
P8Q/069][Y;?T,Z,T[]2+YO:5A>J<D<?2J>8:O0H0!I+D(80WK3_.ETEG% ,6H?<;
P0M8S0]!*3-O)TP7KIK0&>F&'&Y:M=>A*'2(3GVDMI 'L]$4J=H%YQXXE*Y+5^A >
PX[!%/B'<B(Q<6R.$ZW$T-G2YG5[%. [CINTL91[5B7.$::/_N,O*:L[*%F0&#LXT
P4[.M[E1.1\_X33&NIA70_E@V54=V[DIQL!^ \8<UEP'GZ@KIK:36V.@;;]>G$%UO
PF'Q)-A1J>/=XF:R;J5==)H.J+S1I38]:M \ZY"]D = 0S%E6#2I&OD5;RS+L3_JP
P:9> Q&']R3Y1V+XZ%(0^HU9?MT[IO 'V_*%7B2(B:XFC/Z?@R2]8=MU+33,!KKZ9
PDX N-;]0LN/8#M$]3_&84ZG?-HK#^"R[AVV4K;]Y6$IPYP&XZ7V,^HYS3AC:NQ0F
P( L#)A0HM\.+^?]N3Q3V>L% :S[W!5O,\95@Z@A"'RW8L R)A9'M0?7N/1F6Q$0N
PFI1&N WWJ0T]6V=&7,Y6O'IG+$X6J[!^@BV\:*'T:;E!=A0?BD.O$V:(RG*BW.;+
P<?^<1=C&MH8#OU6DN  VZCJ_;#,0#HB(]LQ,'YT3U489>PR8V6++GUP]@BV:&?JN
`endprotected128

////////////////////////////////////////////////////////////////////////////////////////////////////////////


`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-1", key_method="rsa"
`pragma protect key_block
Gc4kT4jn8BUnIl4Ym+JaJCsODNGjyZqHwkCgJ+iXNiXD6lZCjHOKBp16fisekpgu8UWOFFtBm1PW
5vRuziaNadYj5TnK/JgVqm+aBaYqVsBRl3O6Vjv4eAPjygBiJruQktdVJS5hkynZk3N39IQTEVDg
dt+9afULg6Mvu9TEZII=

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Synopsys", key_keyname="SNPS-VCS-RSA-1", key_method="rsa"
`pragma protect key_block
u1S2R32S8Y72zGic2JBmZTg257Omg7mmiFteDYIMPU0+gNwVgAQPozhJOikc0DjF1BuC3Z06vGeu
OEgPftmywkA76YxGQwVIQQX4FwIWbMgx1GUJV9FT5h+b9jFpToyT/h8CbfG1rZcBWuupWZD4aWCD
8j4iZ0PYpmNbok6rXA4=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=13376)
`pragma protect data_block
1qROTVpef2PjSHx4YM0ueXwb8DKxJnksOGeJFeOuXkd3eWBBjrZTwlNhzf0ymi/2jm6Wj6Ty0Tjm
W8K7hPBxgdarQgbWG/I5tran7w3m1987HitlvTh56dPqylfUuKLo25oIRvaIZPJmgeTnzR38hfPo
dDzlHN4M2vs7dnTQt3iHEorVjgwzU5maJeojWw6DeIVq2mgbdbbC06+MgMKwekqyXE6guRaW9DeA
PZNdhNe1JUtO6VyBIR0Xx9Mv5LxDhDMR8HN+9FzjXeqaBLTV4aY/pwRK6iRBIbs9OKB/kMDdmUWT
TOSzhOaIu5q34cQJoqB/8hsvKIJCLEOj2TgXNMqt+Ghr/9Ev85F/nAfMXZO5ApGbOQSf3NkuLyyT
yOllcPGonHb/RT9VMR62s1vr0XDmvPkYdP3I3hwNPtEvO7xCJpeITT4ylRMheVzGjpUSGg67MgdO
fQ5kYjH2zdMh0AAfZBKSLn0i9VspUrQoJJ8XWGj1cMVS0aE+gNVjFTUrfAe3F3/WV15bAEK713P/
ows2TEj4VTwvQTFEtyXPn27QSW26Gf3CpYkaRmtk04HjxhMl7G7So4JiV6iup0OGnMhLQgNwANxN
yg05b10cZE74Vnagpo4dlhFyLQOVcmc3UTsprzptndWovP/wMVzjJh2J8fXWLEdmpF6waWk12fIL
yexlT+xYIPoTU2byVQZfzsKnvZ+sq7a6QD/A62Etd5+M2OS1g5jT5AbQaFdrfaNarsmdX9jZwhGV
xgfiBHFBZEtC3+RaJRrKb4SpITXFTLDLVUX50A3qWTGM3LnIv8FvQhSpBcSlbHwEZrC2k2DMXbhe
CmYRgNqmA7YXXs3X2YaT+Y32w4t1ou4UA4uaoi36nKG0NXpxh96NlTJHfNR1PJ/PE5+fxbs078Ok
g3ycn1bFgvE4hBpgvW2+yhjPmzRJyUK3TUFRgETMRKI9tgpIo5CVh/lVHuInpraJYD7eUtHYCyhe
0FPYiBzttr9GOFZ0SA60Qtuu375Zm6Is0XEd4CQrVLWGyaVYEXjQxL6IcFpnXRfy9nY5VyKVjIK0
eMec593UOdv+9YJ4KPD8aGdXPJYJTbEz/WW27Dg4pbAV3eYP/N6olV8D2pSbIONgAAHc6WDrPFzU
PcWvX8LM21WvvCGOOGI0Q4aHbDC5ITgVhzR8pSokzRE1qKnIeVbCRZbrQ1tj94ymbv8pZs1dL8Zy
GULrefdKUzB4zutmMxIBMW1t2QC6KKiHH1wkuz3hjCVQUs7k19K2EharLNEaqJrSMqhxJr6Ny7oA
RLw+c3yPtouhE0KWqqLc2fx9kl2wEmU3du1E97XAMVr2wJ5UwKtvl3sX39GMuiCURYbi1/YrbdwF
JNTl/2CZh/jCHZB9d6GuvxBgQAUK2bmZH3fE3csvGtk/8Xfk8iLAuAeZAd/OpCU3U0G7nY6N7iuN
jK0H9P5jKrb+4Ef10Ls+3HWHJTDbPuQkG4OcXH2tpKaCJg/3h3JDi5O1sjegLakTEMt1u8+rOd5m
PPTc+gHx409j39roEU50bHCWtxum10aSciElAo2OTfk1ed5ui+5eIZ6M/BtngS+Z8JczstcVJ7gJ
WeR7lDvQPtVHLgQdK8gNavjojUwy7Mg3d23K5ClYZR3suY5nJg/DDQqevDHveaDrwvXJczDOdeLq
8xi0M33mYQ5zdsA8Woybg9UZxdD1HRIgEvGeXIMY+QBHjPZnWGDRv3UFrHDbWCSsNP7hgtEQEojC
5cvNuQtEPdp8Un3WDUELpqgbK6W2kbHGS5ULGEuwRdGe6Ey3BzyYf0CMZ42NQbLE/mnOk36ygR29
o7T+y842WRqdRETqQVcbIgEX2Z7QIXISCWuxAjMLiye0Yy4YGvr9FQtaMazWFXrkEzXFlLwsfP7n
5uCtmq/nyEZrP27e/9lknFRxJ3tcuclHnljHYTUTgVVVRQr61QIRBUu2E4zGeapK0ydEIHCAZPNV
215cU1IFAhTrU3l6OIam5o9hIKDNuiCS9i1tpNPA3TGw5ohAxYlL2F/r+ZF9qRpedZwjjOVcW2Q1
alPHkQ6LeL48wNxK8nX6kJPyCzqkH7H7gpW+iFYQuVpAX8+L7+0/beEk74iu7amqWwJ8tIB1Fws/
xHweqlP1kfa8EO5IqJBymv2I7nfDOi/5EPac8a78w7vQ7t6Y/bq8+04A2QoxLvKP35H5MD2hdCvu
vSIGJuT1Y2TPkJMZYcLi2Oq92hZ0N1ArMxOFhkq2jq1ZOPkvlM+kITm2F3dVMABW7lz6aoY9oAZp
e9gBNPvGOLS5u61Mo0zoY3fyEw1xbnvZJWV5Mn5eo6CtMut47TqvWW+UdSCNH4vfYnJeKkgLQriU
2r/V7obzzoVIAmpBZ4xeATAU7bv1+IGbAJATGqFTURfXTsZce8ESxx2VJPK6CgAZv8AqWAt68xXD
TeAEDdTDFJ2JGJ4a4fTML6+dPCeN0Fj+5IPUUbRBXYljnLjWke0be+b1sMCKC3X5V69KZfL1fxuo
nMuC2a0fQv9c0U906HNTVrZHwzuBBfrHsyxE1jOluZ54xpV21vsNVKiA0adyvCMSXUyYQ5SCrMea
aOHZIiddAFlA/2gB1+TxLaNKD/dnv9ECiUJvyEwvQPXPJDPcIhi46bbfoIlxd8kUn7G02cezah/t
kcGDL6ATc6pe6lS72vu0uYd9uDaUtZJcRhbGDItRfOu3jck6HHy4r0obAF3BVGyr18ayMOHm+CsS
yjwvSjqC7JNjO0Z37+ioYzECY7+C7ezjSIJ2p0GvYQ13Sjuy+GpVzUNkFB9wEUZbJCyjbZ1FRlUB
FQm8KN5mWYooFY7a43/F30/FsVqSAbm5srkAMIpci/kRsDBamNHbMdEUj2CTFEtCIvLedw8uQlIS
uK0Y+cZWHFuacVykDo4n5GXxyTKjs2bx8CSWtcLzN0bHGBAXvWba2wlT7o4AAwoK9povWIDOWECl
EK6hG3C8WYrUtyaTm72b1N62DCXC9rGVJlkRpWwzRoi7Nc7OpjDnnsSI8fVLVZQkdbdLWGtwZUWh
cwJlLgo8YpH1o7ny9e0YL+XFJw/hOCYyxXDE+iaSDHpDgS4Db6RuNOQHZjBMQOheeZtWAvMKmAeT
idUZSnuXDRJ2F6geP+3lZAXyme605WU43EX1E/HIrSlwPP6PE1+AMv81Rzp7J1cCr4DJAQP7+kBP
YtCDFfhLJsS55xz4FZHRbcLJyq0xyCaKNiFH5nkIEx9bH38r2IIK6lyXKGV/YkLmmmbS9SyM/xT/
uh6vlIkxgG8qLbO1/xZ9rhEASngd1lHHEHZat4nfqmoQk3TrNI9RzQqsioYBeAGZn+hTRat0q+Q/
m1NSlG0hOpaicEAJ/nhLacGb7UZ68wUo7qCtLfUYAqEGqwIUEFuKUkES/QmDoAdVcwJtCzI9VL0x
dwX7coOg+uTQad6ikAM+BMXn9FkuLrBL5hEFRoAP5ThDQPF1YBLHhGe3HjWsd709CZ//6mmsPp1k
vc1DILluEPpJZV9JM3ZV9DVUdTn3TUgL5QEg2uucXy6FMzqgOEDaxU/P0m+f6+Gb9aMI01RfKPjS
vOS/f3XlNDHegk2FdQ0f3Anaqb5Q4q+QV0rU37ap/4+t+XS5YvqHLzcFxfOTRhgRg/rSsP1yVinA
H/12jG1LoIvLqXCf8uDA4+LhVepgalCmt20E+4ukYRrbDK4Ci59wS1nFdlarEwVZBo4nd+CuOAuk
nHQnAveqbHa5e1BcJur+ItI+NBCcSgWrGGyGXbL9QVvnX5cZqfMDGYD/e1Qj2JoojBpT5iXdy6Gm
qlVkJsAhH4h67d6lMYbzKcvd87Dl022pnmai9NVqgHY24ot7MYVdZyw8iS7QsCZf90IkgVmnkGRp
QWB8d6dA2akvtyyjzImr13DEklF3hs4vNHFw4Rn5AW7x3rJLYfhW7NrLl8Ro798dTlKeJCmjos/7
sTv/c+9WY86PqbnWDboHs2jVPi/VaF1s9eb+AeIGg3P7LgbWCpNBEa2aVWfCKneqmSSr/KC/UrLx
OyP/jdI2NeetyD9kNZFLDjq2CKOYj3FPzf3nrcbYKS7ofLk6laP3Qhbjuc1jq9NQ4Xdn0rM3jufe
mjP/jyP1fiTX/I73nBr54XZUnqhYD/durpf1GWsUtWYZiF0eWsrJA5I1kL8ExRc6Y/3yRd61k41D
ewYKQMrFGWo409N0mWZV/JetahxtPYT0uenRcRhXfXk7hWAN8aK0QUsDSTi1h8yp11VKsRKp52UC
QDK23RqlDQ1NjwgBImmNw9OjQIRrIMGhVfFmXp6mW1+2RovOeuFd8Amn2tjBmR4WGZZG2mbZWpOM
JVc3HxZPV2iABBoOIBOBBVilLdqpHoLdpX/1ZMZFKoIfinx2hH9UU/yPdMXra3/rV+eGX3vFLyZB
DA0P317lFm9M7MxGA18snhDZZOzO/26fV5rpDxTrsjgcIwik0UK/ZE7+CVsR3xJSFGAnJMEOfrjp
sbmklUp1uHZWe0zn7dXowY0ip2tTyQwi+RE2NcgpC+N4/V/0OUsyUgmNjNfV5+2NQSUxbpunEbBk
rzUMjL+nuyQmyxQn995uz2BWbqqRv8bdTCJ+u9M9gOWIkWoMfAhgZ2iHSc47nLCI/mS/1cMNFwq2
9CtTvUToAANWEqdi7VApYsbSuvISr77fNGb1/n9WnAnNNe7CYkJTHsgIk7QmxkgvKXMviRMaOqzV
HRCQ2cYhFf0xds+mJfmlG+ReGHr3FdhL7OoWc7wo2zJ9LsLbydcRBaCETdjSbKp1BwebvwZhOtBA
CxQXYdDfqahEjjKO26NiTgj4zVAzywD2s598IpjZPS5t5jVVXIRacPIfUxQfcYlSCkqTI3pq3V6i
it5oIFoUFd7kwwTfD7BRQ6lai/tBSFI+NNQ081BiLy2Y39+nAQbjy41smXw7vmzr0pf1JVK4N6QX
ZIdyZxb4tDYJtTLLg08yGf2Rb9Fqxg6u2Le9Ra8atUIe+ow/aMGrB/qpdiFfA9WdN6I/gjtxxagQ
ApExVlG2LvMK41huUo/j6jiYHgq1ZKAFARrBwTdsgLhtIjIwHTFpFk0QgMc3nlWxK0zJJxrhvFOl
ZZ+0VbMrmr6UTCX054UN4XFp66VBTqyi+OmdalM8gf81Gbvlu/0EIgg76+uuFTAwZ2TCtRu1m2o3
IiBTjsnzd2ByQmvZtf1d2laNVuyXvbRCSX1pt8AkldIbSSKnODtMENGOfIY0w5hw/ty13TeaIkH1
IdZTEBxd1x3FeTboCEbrudFOoN9FuCwib9E//WjPYgoOTeAxWUkT860lV5q6Y49KgAct8aLl42RW
VdrnXA+dHHIFilgcB+Z73yIlb1cN/aZAW16Q/5aELr6drbzdeX8hXpWC1VcY4yr+5kjHO+nPsuAh
nvtcT2LORSvsdv5KNRee2fsn+qAbyprow1QSYulnxX1f9vPvdRXHUi7Cgqh9+1dh8pfqJXORxQ2w
BCYvihGDW7OWdt+ORo4h7vj0VWygb+scuVo13yA17bRl/5ZSIO1UroJ1VCyQHG/eOU5DI7PWtOnQ
g91U4Wok80atJHEu8gBKEFjkclkVsTD47Tcr2UuboiYsSg6JyXcD6A5+TOiXdKXE5dIchzwRLztB
NjSsz2rk/1VpH9fzrMgzss4pg8VwkjqoF+yR1QnCDFW12gpaOLsY6I3nWfg0QCNC3UdIfBJDkY7I
exlz2EVvkl4+VbeFNLnaSPyZSRxR2A4aueN30D2+FnkD4y9LOtOaK/M+oW24HfAMPPCfCRT8Q+Ht
WigEgGWJnib0RbsEKMqGWGI8+KVg1rG3fNElM1elmEL6Gxcwa8FPrqUxVdoaWo6vYH+Q64jymD6o
cvPFJqbY8f73fpgMvVhN6LXaKp6rY5unxMKwbEqsvdJk6e3SouuVPkrQVrY3ttZcCWk1MJhl+9M+
CKQJahJm/ZVv1T8TzbF7uoJI7q/AaeTfaczHlwjBmlpwKEllVZ8/nYAT1NVVQZBMxMZTHwhufmWx
n6X1tRZIm51NQusHhlLTcyaOcyb0wFWNvZXSciuEUV5Jl33SFVa0E5zTfCtf05pkj+jEc7d6S28g
pRfI2NaRHgN6S2ZL9JL/XpE5J+06gezu4WjyNDH4e5GWSzkHp/SkVSc8Ehq8sngMkklo/GJid6pm
C14+imQsnl9fqvEjudjH+GSjZbeOtoXIbmKI9ZUXlsX+o7O/5Cz8tkxHe0SO5TdJohASB2h37LF0
WB54SRvNJ5+kabdpGTPfqsBmNhYCZuyoOvcjpacpr2IitfegPAWDfgec/p/JgLvRedCSXMujS8Kl
GxRUAfG2Ay7dWe8QtKUW+cGEnhS39a+UxCvzwikCLfHxFCW0x/d6kPpGdLgQfpO4ZIg9caGsWxun
AKswg//Ja8fpvtpSSQSDk7Ri2QF5kInUTwYvSf/3VuuZOTCedB5ewAULHUmB0/XO0jIcAfA8T+MS
IhwGuBHTFewVtleNKmN4SZiR/QePwcUdoaTyofD/7vJ2VT/1ydVe71zUVzOezHFnWbk8UD2yQ+7J
MmswSNjWVbU19E8/p3BMhu8KLe6Q55C6mx/jVGsBp/EMqn6+BL1pWv0GJqx5RogIkjdqtqdrV///
bGIrHDnNmBe2Hs+/FoTOHdVzjmPWxd8uHRbOmQFWY6TEHRJbo9BUphstvPAMBLNaEEikhj0cN/Zq
PZyu/6N3DcF1lGQnYgsIYT79gOT9M3JNkkDU/QcVWXG5UmmWbyVDtJon9B07sbyZ6zhZwbIt/zbS
Dwmd+7YCFqeydsSxUbL6Hx6jvqqhBGJn4/5k6VdXo/6N1k0AlPzglVgoQJAmFlzvdgYeHXCuKn25
Yb56IxBf5hdclQ/+fgYu27hu5su5Aw7rSQvs9Z96YNIIZQt7lo4nVYmiaKVlVEbgXuj45mPbMLA9
4TBTb9HaEfw0+cpsexb6cwi/o0IoEVT02N6doXnhJdmxgBEAQffXjspChqd4ttO/mROJYyuaB/pS
85tFuJzxeBim1QJ2H18TqcnXT3dZMBEvdaxISevvRIptnW4VyLQoj+s4Gw2bFtfuCa1n0Z1Q3+zs
CYPhXDUzCaWwBEgf7Ln0s804S72ygVct2BNbRCWw7BOiM0bg/BCKBrMv2UM7QerwW8EANx6A1PVF
vQ0O3gzxwEXnzZC+vNSYVgC/wJs92+swPUn+VzXxFCGuCc3bdl3a23CouUkSWgMsTPDuR8ODpeNT
cr1nllPeqkboI1bCBi3nMOK/MDBJRgP+HFwW7CbiMdRYKUEegtQHhXVppJw7ttBALn/aUKlhptA3
ntiDzasVwbVU8JZBCk3XPR+V5E2tHsrI3d2Jt5aUFinqNVzGph/4+AwZaYyuoO0jCmPAXWZdDhON
89Tu/gUoZ9Lpg85+kIC43wEq/dfi0P02Jhx/UGsfw/eqZ9/OpinoZ7FPQWXH9SOsY0yTXa2jGYvg
syGk/bODJKRG8YLYHFta9FdWHXMyuHxeR0H/DnfkOFKlRXkQUDq7qZygPm5DEHmbDMNEidAa53ku
U7FcP3ZNBohEEiAgirX1zCCeHmguQISeLgXrKCCuyZ2Jvilcr9rNz+GZA4gFrF82Llf0ZW7shI9q
4WwuYqCw97xMKtzx4vmkFhjUNoLtMEbHL1UxI8FRuQ5hSC2NfOFrVSpZoeFUH1JRA3WCZXahHuOX
83arEeUzRGd8dQ0SEAWD+Q9nKQ95EalgdU9cyuQPXy6fhCElG34+BfFY/xCfH7Z5pGlqe5W2IFkz
L6nOVh9cVbkPyG634daFmwzN6yAN16R3wHGznKSDYp7VcZPTef0zw/hbj83CdwtRheqnSH76Z9FA
+8YCfeWleUSTO1Sti9EJNg7rLVHFsFLqqFCnUz4bhd38zsEqQXqBS3V0BiBUIe3QKqxcyBneKNta
Ra/8qBu8AAhN//rhSUgoMyBwTRUfQpp3pPV500tsQcKJ+2DohNdpC7sMHvkjdu9ppyx1tLGoPlfB
Erjkwj08GIQOEAQnofVNpePd7PJzsYkv4CegXp9Ym/NLRRs8KldEd8YhUirVMRNmMQCkzneo5anb
KO0qpl+Okf2QIvYnqn28awZvxoh4h2JjvoXmdDY9TcHxhRdqhW/w+KObZhuPGJ7ph8+OT3mwqQ6F
k0iVw735PnpL3tw1hNLm3kYa+Pavz0t32QFIRy+pI1HTowQeGV6p6qMu6mt6Z7iYOS+WGJ6V7qeD
8nFcV8jcY5shBMsexbTEUS4jp4Gvy4eY79K61S+EwOatRUl0dRTSzvspMHiG4w89mpjenlUefSOK
nzsaJyoV/gc8GqEdNKYt1p2cdO9B6iee3jCeH7zyvWaIzRQYD5G/YfyT7nRs7HOg8+bxbXt9N+HM
SI0b2AJOu7dO3qQY7s0WulnsFAdstinlqA28IBKUKoTU/cUlLUdyMlww634SQadOEomNPktDSzgX
xRiixJGKqLTc9biWbvv6a4hh7XgNjIlTG/NYn3UqwGc4awqzFP/qXV1xQd0AH/n2J2kCaK63M3e6
+LSQ5a3nBZ22zVgwVpTdV6/hez9EYEpTqzPz4ivOof3VWWZsG3ilFzPXTKTWURPl6ftNmrHqdtes
O4Q/FSRXVMoEERG5MkBC6RFibpbVGpLneTP4zZ743CFqAvtFheJLnccZXz2w9BCx6qc2NEk2tekY
H4YsSp43wzUK0mhFAd9QHkAunkRrU/GsJMT896XM0msbjBvX+9j7CpLUFE5bXYz6CxnTilVFHxAZ
kBRryP5h/LGA2zv1EKQsRHnmapwgI1ydU12PttZBTfSOJ7NQO9Mw9mdtLoMhNoqSQOrHPROuVfsJ
FsvG8SMxKT2RtOtSyem14WXhOQACFZYFLMZFKaja2Cgjm6MTVxdXV3zSfiWw7BI9T0g2Lu7MpFdr
UpcC5o/H3xAMlCAJ1EFHpzH7c1OyTa7nXo+1sDLHV+Hsbm7NzNI51vp6svUFfJXMDd5cCzAbT0uU
DyqvtbpYf8cFyJPqml6cfz5H7QOvPRHaycjQ80xGf/mMEeS7wOoUbkpIyQCixhWd4NzNpKIOLErs
1aWcdn5uYf/vSdqrvKGfBEPQ+VU9MVgKGyoXa+FMw27iEdHI4hh0qU8pLNs6ULxTZVKlEPHR5L7o
alF692U7v8ERRrRHdKwOBxrMwDpOLHsGREObLcDr2kPa88zY1E7xb6uBw2CD+henPj9zJZrGSlE/
j2IbBs8eS+TE+sc9VYVQ2XYF+zAitWHOLpZ4ZxDBoQEeTCstKaCTIOkIrYNOeLs6tgcd+I1klXVR
340DQ6nHXTpOtdkDSwZAgz2skJzztA9724j89OH2lG0E2SARpHynyW0Jcun4/ofcJ4HrwV4rH/Ko
ny+OjEjHscChdcHhbDoif3S2D5IC9MV4H0hgKLVLUI3P0m+RVpCW246RlmvZsYETXOQgZ2NVaZ7e
kVpiNS579ZKSJyzD/hdggIBE5tQ6wcx46/XxmmaCS0LJMDN2LwA3gDX+oBx8qSGDeMxq0y/DDE/5
UCTbCTPcTnuyVeMcIIsf64JYbkURLzC9UJ0Idyp6xnwSF+OY1+CmTE3oKNCGxfXq5I6RuhjWnldv
RqJs0JEZwZB80xCsAykXCUxKJumJd/xe5CnYWdfA9Sd8jn6MO9mH73PWG1pMyRHdB/M90LIG7G4H
5MZDxd1EktBpy1WGu0a8+uma/16YnYr6GG1Eqfe2CBcq7OV3hk2JbSXwmP3LEh1M3fTjIya6xNKo
ijXGJ2OPuSIvp5z4zgPvVu6FLuMhnOcPT6lMFLtN6qafndnjFSqDqoRzuIgwQCok6ZQb+f94Z0fi
vNWgD5jmWP3EWadGge1RFK0kzR6m32tJIrvClQ+E1NxqJoPLH+UmV/UrXIAyQfICoWUbiAmFvCqj
GAOdncDiehvpzCg+zqw6b7j4Nehaxw2C+40rShyZYYIZfQdnUrUJmNnHXvsCb6QFmn4NABxSvdKn
4QHv+LahuEa3IBFBLyhaKBSAcDZK+uDR2smQhOoqeqokL8xOLWpuDKupxSFM1CKN6oBW7qOkizQw
GlvhFGkKI/tESVXAjJW63TESIk3Zmm5Q1ecOMm52W8KQ0ZXmHl1OsM4KiJpUSU41DDhuew9pBLDj
TbhmykIXsAHwOWtsNJZ+/3N1pjxthMQPSoB5sym+BBLYYRCARctn2nGpjk6g4ljqqvz3fpVGATBz
BlNlEWplMDe1Nni38IirK/FoRFWXqsG7nizXsPJUhukybi/IoTo1K3N/2Wbp3Wt6Bo6GxhykXOfO
pxTwyNVtqxDE9MIxm+TOkRjoULra9exnwG3gSn+tAf9DzsJnMTyQ1VxP2be3IqsjFyUX3vB210fk
U7Y5K0xOf/Y7Q/1mjYa0uje2EZCqYkeJJ1ZMuEjxi9tOhTq5dOXywLU2JdmtoDPhWoEynA64/7KT
1LFz3SRjUGKnbRKvxU79RStIHftCUkhct11gBcd6dKpcFQPkqWcrC+hhU3Ms8j83U7SoWg86/3/2
BmuCJALlUV2yiF85/FCYQugeOSTX297KZH4qJMB+suAzQuX22TQj6grf1dPbrXCY0HLzGeR01Kng
vE+y3T1iEaxaghBQMgMddfXHP63uz/BaYkvdXoLwgc6+mqhGG7uLyXxFwmAvyRkXl+Vm4lDG87Jr
5b1yTo4FA38AwbgHETfBrFalBO/Ge2VeH5COslMj41ZgjllPFg6lQukmPsY3kvqJwe7mciZt9VlM
A0PB5FvIkDS0zgLv93+vGzrJX1uFfsJALH4tyW8yShH+3jPTYRYSIrhufw+oFytzu5uKJQMsCpAd
kPrhY3KK/2J30Yld5OsGeC4K5Q9ru+QQRulSFOtyK4oThWnGx4NDWJJAQmvJWpwbg5Qv4HG6rBky
TQZVpu1VJ04Xbrqb9ViMf2/dv9Y2RxNJppve3Vg4wQQML+a02mZh4K3jFnbHXDqFZXoW41TWMWLy
HsWPrb/qaR6MXxHeqOwohW2Xs7zXD178/u5qOFIFrdb9ATP1AS18ZT0pbEnguJohcDk7THuEFfq4
STwKfiHYSc/BhLFLz+swkXLrVXn2LR5ffw9pX8xNQrMkyf09mSVjwrnVsCQ3p+mifJoZ22VwYjKw
zqvpaNA5yo2h29QdGmriBlXFhdbSPFO8xoDwtHzF2Gymxj3OQsfM0H+vI4PX5aAqTavuytvT5PFV
yn2iR4no+SZIbde++gnk0MtkEZTrxlm8geIWDFRuDnH3DQDoMwoCvJpo1kYUuZ/eUaT67moSFxcO
ohffe61M1Jza3jsQgVSLTPWJ1cwpIpeOHh+wAbtWRvlRp9D4nk5Y7q2yHxBxEFDn9fqc/vY0DgM8
X46TSvoP9MD1LgJ254Cr40VQ0lhBdlnTw/Q5InQA2WkD+rAY+rmQ7y1rl/vRhCWomEc9NCLG0vss
rgCD4UFkIddiIkZK9rvXuCCqNtsFA9Tf7mhAcRPlmfQVtS5XCNSCPnsbC8dz9ovIBpDgVpU3gOyJ
JL1n+PN+gveZy/5fsuenZuPqTuDvWBfy9uAjmaCGdFDCOpUG0wMGby5dM2/4rewQEQfhFwZub1C9
kpaMnSt3Z1R9h0qPP2YDA2x/KakGTnyaEzjS1Wl6E5ytUedapfxsmjkBlC0CHWEvgOwIjjcISLhE
+w4+hT40neGMHva1iL3Qy6dVu95FugUxe561RSWG1tdyeRXRW1DVTzWYpZpVDOQeS7Z2gKwU/I6t
bzbKQSMVQILh4WtMy94YrAs8qO2dBe9FwO+eTmC5dyuKXvnB1LTXkym9xtK0X/D9SScXqHvx2qGh
44U67lFdy7WjWFz/DedLUDZ8lBCLsQ7ZLpGmu1kXroC/tyKJeqp1ronIxAuzI4GNdictmUqPoBe3
4pdl6tHpZKv+vwNCwe6p5quWJTFE8HLw7tZF5i2LPNxD7Ic3SJbi0rKD77RiLdO/SNzSjqrngVMc
R9ohhS42cbOGy+yMGFZ9fvQ4oInFWwvnBN0UE4ReRAohAFbZ9bbfPanRLaCJt5pBj64z4juhK3Y7
AGiWxmOyyXMBUfw5N1X9ydSV3FM+wOBs61ZcGQWF/II+10lsXJrSeD/WHj3bAO4Y4JHOLkkF3fwF
VBSCdUIECBBCgkzj2206zk8Eup5tlOJT0Zs8GM1XKaawvSr3AVhVqdSLD7zmXmH3H3prJMr57pYt
qmWsHyLrxGfBnT4BPLcdYQI2Oj6FBSXTI8rY4cOK7P62e4m3+KCZio4o+QbX2R35qfSPGEfXR7fA
RgqmBfwTZphAPSBta6D+5NSPTK6yYGYgrMlFcnIQBA5T49mxH0nGteZfV/04cBoOp3SL7+fb0anT
lEzxI9BGRyIaT3uTleborpcMaoFF0BxI2EvgaeN6WCv6It1umqHpfMYUjI/G7VkJEGoSkCQcfpDy
IeaX9A7/UXTPEK+Y4E01TWERnc4CoEg/kjIxrpcL0zObYxiJF70usTvmFmbV7fP3IQoDFFgNj82g
HQjj5wfimnahjeFkftzgNKoIbwk5lUYERItNVAnDWvALhxzEF06mF+H/wcAWdHlpC61EudNG36e0
7UV2MgvhxFTOzxiM1LPa8yCxT/m9V7MsQBBGSElzshPyRv5irhI9B/E/0hEQJpJPMHJHsTLGBYZw
PJr9Wyt97XcwZmLwYmO2Rdm09JVy3lJS5gM4+KluJwotftlmFOWMvFMPD7QRrhNBgobdKIAd6Itb
VDYGsoJHmLWDNhShlxi+HuxaF9tIcdLk25MYvslnNnPfvKawxkpMok0zCHvs0igVi9EYOx/eyA8r
xJLbsne5DSGtQ536Q+XYlEDi3K+yGP+tbk/ZoLk2jn7l9O8HEvo3Htbe/bbbJ/lzZLzVbTciCcug
RqFemUXhqcDnpHBiqemSq+13ISIw2XEIkjWoqUAskGfkhV6ZxPi5XlnC0WlPa6OJvjFVEX5SIcis
2148wvOoDJWc2XFnEy/jhOxyOkIi0FlWE3IQGND6iAzv1gQ13P8xqzCLOih8+iZGy/dKDNHiwfah
6K+GBV/9mVCFj87pFHXKkfrP4S70UoGUwNo1sRqTeSfdExmhf1tpH+BrFqPuV7bcWPrKs/C9b3Oz
XYyU9NWGsqPJA3WOtp9y/Qk40JW7zKSq/EcyyPkNgIb4tMDlTbRhV8GkFgMXpcDwpKd7jHRig4Wh
PUXuz17yS3o2UMRCSfaLlBSfvrMjOxvFGpoGZo4FMAKtlJBmQPambe7NQnidEJWRYBS3xCOsOO7L
JSWB/6bwKbhLDS+aWpuAMzMagOz9y0+BmJC8Nu+KyNC6+zSO5UiR5hV2D/r1VEY5LCk7fDnb9FaB
6NJDcDkLzJlWEj3IMpz68kIxZ6oTUYXPmvNCc/BSPctLkVWDtRooE2VHOCrLVNVjzqV9b1VWUcwt
VKOhYtxHvFgW8Nzo1jpxiME3B7EQvY7mzYZGT6ZFN/2gMbGdYS3JcsZ0SZN3KItjlEenfQ2WzJHC
JLdVS5McU9gFv6/pOlne1cypBg6JFGYeMlSCeX/KcL6VFdddmkrLLogqmJDratgiY4yhCMNY8z1j
NtL8yOtsa4C36jZRUMOPeYLyL2et3dWwDwFrhpOL3/eIGaDTFz+yUz62Ea5dETUcHgF0JHLQVxQt
QHQxEgzk4go6MPQ+pVDoU7D3a70Ee9XoGuT1c6qKTULA6PKc4BpE2Z2uS3M4+9LeMyK61RgZxWOY
LF5IBuQoeAXa+TNZTyJDqYrsABEzZlfnlYbTjLwo6zT8dAurzTxBYQqR5vFvJSYCOXfe/KZ24/Jo
tRimO3Z7Z1SfgJgoZ0reL8AnYJzjKjMC/uSCJ+7+H9TQCtCtB5KnP6dxLE2JcaB7YcRz6BPf6nLt
oqN9K2ONiyr3Ae+09TNhe1oI+uI+KmXDLyC/0NR6EebgUmjF7+WijkfULx0pWavB/7qmCYtFMan7
NNoRbK7Cn15V63HCtDJRS6/qH1neW3BBt+JedgpzKGHMW+FOyo/YJ6/uB8vK5J5Ji0BVCINS6bjM
ntzyDrpt/wqGadZCD2KyV4ujVdRko9cBVu1MrDmQxlhtOt0AbztEGGuCSz//ZyGZw0xwsUrcGez7
WkCNNVe3p/F9kKcMhPKyeCJ9zqGQ3sG2+Ah9L4RKvwdvFRxIAepn7Li1f9efYJUNfWNaPVboKWP/
WaMfjR1y+aEANEudLX7Diz3K7fkAR4MsB4nX2INCAxV2+52P9ZnXxBPqFHxjbx1Jdn8eg/921WOc
srY0Ydd9SaiyJNiVlNdSx4FFEin/uf5ZssCvogqLWFO5MWEnRSR0KkycuQ5bh1nsHLTQqxL2ExAI
Djy2Xoy3W6dnwjCfN2WexKmAIbuVvAw7FeJ7jn+IZBrhVPMMRTr5PB+/fAG8vllL7IPrLgyPv+Pc
B9PXKambi72reQhMv4oASXcxS7TYbhEytCy+5+xhNKCBwBujKZX0ztFGAhzR3cXjkRx3cJpmEoWP
TQeXM4/rGU69gWuEELhvZS+VnBXIY3XN960fXdHvouOFTHbvLLdx1q0fUW84zCSX9HxVBxVRrRlz
7eED5Tr+VIF9H7zKR9SXOLviBkc3BdEE96Axajk9Eac2ZK432aNvFXeOE+4oOWakHdkzxtB7ungu
+kU5kvw/uvo28rK1UqksCpg7E1+of8edtEfhY0V5tmYkD/I/wmzUH28AbrZ4DlOn4Uo1PAat4aQL
UwjqnGCWLMiuxu++ap3I3LvtaZIlhFV5zO8LVpbrAGcYGfUh/kRihFRhm7wkmu4NNfKUy860pjUP
57l4Z9uamayF2d5Hd5gKu/35NCZPtO2WPnBilhttbDiWqI8S3EKq+H5hYvtSoxZttUfJ/xCiAkxb
F9D+VrSQXgQGdJeFGmgjxFDPUZcD/RW5rffis2WaTUN0NiovpesAcDwakCuMoHcg92O7xGDHAUMy
hKG5lX+aCWd9G6rTYw/1Ifipw+lkjIcaVYuR9HoN/dyvwdiEXkcWPW2Rvyadgdw3m/3jEAfnTdlF
fAO78c+PPqKQZHDSY/FEJdLJrTfmLO1kLhdNts4zWDU/G5173La4MWmVcjls/kX/wPx32ayjRCXL
KVaLr4fdUlkqqDcof/JpohoWapFx0mqjxz9XysB8mM8676yhWjs2CBUOHNjpJGGciPceT/ejp0vx
sxzuoNkwukSvfqnoPIK6F2oERWe3THgqj9y0xsgewXJ986RKdt9/F8rq/mFf23b9nKcSjbNYNDqX
tjH7MzTSUpKa6b1zpBH9ulOE1OXlmRvZowU8xHHXD0FjMXGEit7FmjGdUYkz8aRam7qfms0YpQ+2
x2DXhfviFV10yQ/i9SGwMrWq7uqwNbiiAdajILeBggqHz3FSHt6tdEhvrwlG8C0pnQj4iizCDvwk
hwPes8hssla5NTSnmGPVYtuT1qZgYmMKgd6F1ntfLeSkA4cPH1oMBSBj5X8Ku5Q69vOfusnqvuFV
ZtdTUUcidlMV/4Y8z97hMZpqnYGRV2tCknzLL8L3pUAF5iuEZ6v85LuOAWst6Iwecfh15vPsTaVu
+0hPELxfZSH6f9mZGMvWOmji6ZeeyWpF5j8JqeMI2WQ65ts3J8palJJJd8ygJqKcfZnIRjpDCIg8
5Mw5svvEMZONEEj6vdgdXns2rGSG0aj8a/wr48L0zBYjSK36J2hTx+1/OxZ5PNdCWcSvtUXYWVTu
2JCX1Jx5W+l34R3J7IH6jXPSzbzxEjvoNfjZfqxq3Q9vzUiA0PDk8yCz7zBOAIaQIJ1MtqM5hNX7
8MJtFhiR5bYEHXf4NPyBmmmCvYrbpbIXgMAXH8McEUuFZV6E04fJafKf0mmlH98h1sS6c0/PhPIb
GuW/EtjP6G3MywFCY4em9OMFRFnyIUerGj7ud1IayQvigQLpi4o6sRXoEyDloN4d/tHCEybzOmm3
GIEOodpyj2S2w3bThosXqREe3Mvgvnok3dVRoXO47q+pFz5qUUKmNDjtg98IfE2X9Gcj945sGKce
954VQOuOgNyoZNrkOweVX9zv+Rm6YJGaemKYRESTj+8r7zkYOFda+8kIrwzvv1WZEV7qgf6S1xj8
u+09qHlX3fwtNx2roSNtnBHpqQJV8syRfJRsoD5dCnWLA5h7apXPsgGu+HpE0wDWAJtsWwoTw0So
q1Wh9+jWv5nJXnsLVvPMGgYfhnUOwpSdCzcI9moSqpOZ2YSxu+PHg2SOz+2bFExcM0ph9VZNBzqK
e70vWPfAMpzC+ZQrBD5A6Y9qFa9NjuEdMvt/S1AIeWm1TRKyLDDT65hLbZYUliNkL1Vbf6fD8M9C
9tKkB4AiwOdSAO02Ki+seN0aNZ3XcyhJebS/3kVVCJ8VME/zZXYRV8R+d1oVB/GhFxnO/cbNLJs7
3Ht2xTz8Uiqz+E9IYSEqPU+C9mtbOZUsDVsBrkH5hBsw9qigfnKzsG2YzU1tkdpGWroH+s1wTf7C
xAJ+jO5yMnGBQCGC+yCOJL8oZW3XhdsTxZgWAFlm2eowqAu3NgougOvs4za0dkWIwkBKhBYZTuT5
Lgo5FVhspDyEEU2jvkeA24tCp3eFJdB3qxHqhZYP0ad3yfjMItA8jxTIA/svlvE3zIigiXYMLCnU
r6IGjp27VxaaticqeZirORvNwSePbRljYoCSqkJsznpru8ZcvXhwAfwHPn/up2HbbMydTog7njbd
WBX19RnqfCDZJPpl+mfsFA+zeJ1sJzM4gRlqRgYySHSKhTzjLSLjQwYvQEkzaoBhlr1edcmmStmM
XgBPl4kRpfVXY3TBqBlKNLH+JlONmfn0pk8tuGABzIq2XWV4t6mySWTjV6sA54RGQSqmE5N+ymH8
lPOi91EAOS+atdizESNqFHH4uuBXzVk3LN8IPNqEhzZ3LFmUgfR/Py3SLvn2tx/24FMC4JrEn/Mb
BOcUExDR1vn89l7lf/fk1NN1d24oG6hXirUtEAH46G8oRxzoZpC8y9DS9/q0QGO6Pa0xGcB51H0H
3kTIw9jY/Y7KzqmK7kp2fVXUaVf2vvQ2DEffIiV+ZWrZK137idxc2yy5IlsIHDkqim/FePgX6aBk
3OUFje5ZkzO5PqBHQt+6hQmInGhDpyquGDflIKqg9QbbcpZCex+MK2DPhbDqqfDFCDih+BesF2Tw
bpYj70HbzsVc+m/kdvE/Cm6ylSenB8Plb2844aal0e0Hzd48w12W0Z+xyj/wQNhUjieDBMKyz32b
VQBTUTaiffDmlyC0uYy6rUAYZ7AhQ4yBAfoEJDpvcnTRWqyV1FuCEdgxeNtGpHeK0UtV3cJkmJat
SX9bX6mEqd4mz/0Dj+fijAhAvL8oNpFPofdOEOoIv7OGtACQNkWdrMYPB6g+jIWwvbYdFcn33623
O8KMiq5jklLHAfsgn9QmnjJqxlyPOD9BWu4sEuKIA8Vrbv9rCaNGrtq4MeT4ugU2B03IQJjAoJP7
N1WNpu3tAjlkCGxcStZMoVLSCMezm3hhpPIU5vB2XoHRpX/SbOtjSvnBzdxHm97DkzTkYo72gCkO
Abj+xG2KapaO82KVuX26c8qYTdyaEClnxhkYxVhAPk6FstVjVsKONc5i2187XqmY02A+F/TL4FBw
rt0TuUVbzvlzhtIgS7YGbPh+k7NO3uQF3gLYAsDC/AOz2ubCcCgWdpIdEI/ltUQWyEiO7KM/8Nj6
/y6e++lODth9h046cYSSzSVd5fwaFYnjm3r1iEUA4qj1O8emQLvEQNN+J4m8bg2AqFGp6r+LUuyN
nU56D9S00MQbkz8HHJUjTJEfZhde9SkFRn47bUSj7JDuhvYlIp/f56gLrCg4uruNwj0nVX047cLV
mJpDP8+hiXFaVy17Wl8Q2wj55Orx6zI7b7Rwuzp/pawO46mxbws=

`pragma protect end_protected
////////////////////////////////////////////////////////////////////////////////////////////////////////////


`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-1", key_method="rsa"
`pragma protect key_block
a9MZXZYJRwI74tgXoaPCfXdj8JcqUCSmI73DZuv4kFK3BRSPa8izvu0dXvputLqQ3BsI/M7Dz/Pm
d4pXY5wTW6ObFt0+1z4npqX14LN9DxmwUk+B2KCgsL9THPecRq9NM6Kb2t9hx/utDoGDGogIOma3
4fw5O41SrkGxxB8Gt98=

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Synopsys", key_keyname="SNPS-VCS-RSA-1", key_method="rsa"
`pragma protect key_block
bPMM2R6tsueN6tkWOE8/mTmic26hxf1/CjFVzVzPJSY9l/o2evEHW/7PfEYEN8NeoIVaHsEKJtsp
lA82u/medk4+7NiBv0nNBRSxSSTtHP/XSk05ojDSI8hS1VmVlIkH3tF7kaHcMdm9sqvTKTFNDwQh
kvMMub6ezus5CmNsBzA=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=1712)
`pragma protect data_block
p/Z8pPqxfSDOByVmXZNyNZjgIKlc/EXmwxFpfinoq3mC/nr+XHQ993P05fGxHpYVNv4R6RIS6abP
euiLyfwHYgnM8u8sjUC/TX7EJRHtFDC7FGtnwypAaV5Xk511Wj74OgYFwhlrFyEWmJ6BqqG0WUFA
PT4MMyFtc06CUUbvyrmPtxdEqkA9tY4sunjzDaCwcY2X+Cn4ezqdVFF66SwVtEcHzAGJBEoeIHj2
IMz0AsNxyh2s+83Lt3rqhOfs7xcFZX2HNJrpOMdocBnTn+5CNtcoAl9QzNvu1YH7/E1Vc4w0TK8h
m2r3/Od9SY+QMdKHfl2mx5WE+a6bTNZW5OoYiByQsgL/KW5pPUKa3XTf/wuqZLpYd9rRq8B1dvWQ
+0z6yJiCa4gXwhX3eHEkjLNmEnQddHqPdoDRPXdW/GAZIrdHj8+fuZ20lIp4XcoAsJmLcT5RBU5H
jS1TsXWElWxwmXVPyOY/PJgnJoctq5qqVkY+xBLSzk+n80JfYKFJPgQyvuEBblDZLcofrl/0UhLB
mnc8XnIQ0S2pixMU7De29t57TsOoKnpk4PPvb7T/lBBwN6mOBNve3iTk4h+sk6XyCO5/z7m3Re0b
YoXBoD9LY3MaEZYv8FC81iwkUBozHW1IFYw19gcAGLkYwkTSnFuYlpcKliQTHwXsw5g1u4YooFf2
PrUnvHCR+bi0ZsGgUlARV4kAz4uwGWmbvCEVMbIE2515YYjOicHCaLJ4tu1mIX2CzNMjbYInH806
sFN9jaVA9Kwudcxlxh0FhhpU2zrjVg6BwUqQk2u/quEyVqBriYcdVhtAUF85aT2qhL4FQx7aiPDA
tZkgGAjKcqB+ymndCD4Xi3p8b6mXXbrde71ppIDjDE2/VLljd+ORMHeJwYKhSvy5n5dX83fqsyU8
DvGmjj4QNvXoX+rmN0Ka9Pnix+skSi6+Btt+38wPf4znofEuzyrveoE2Y3435owMFJPaOeQ2DpE9
CDbXO7aB6NocBrk6NnhyCfMlbQOx99oCSZuLisRZrh06nq9TOPrjwWEgMvqVmATj8k4kI4BREWKP
rC5dVtD6HwAelQRtyU12dP2p4/vTAog5bgfEovrAKeYKf1dkXV4cFf33NQA+ABQBNRhuOPdlGRl3
/IG8GKl+BA3S6dnuIN00ap+amwxxOLqQB8frpK8NB0ONsy6v4qJ2ps1oy5H1Pvk88mftluTyNv4H
raGjVd+jdHqIpmIvNux6puY6D9z87K17zd4AGDEZgyclp86puX1WH/GU1HCZs7Ca34vxkzl+1ZMF
W+GK2ddueyC0N6NdZ0y6hRJSGOS1iDtQq2RR72ZAM6RlS60nLxFJpDwMhTPwQNf1UumMCXuuM1mm
4Syc2BClUweQ82RttWRcXpAVR/Fx1s9frMLjQL4Dbwb9ttwpasOAwGnsp1QnJZtKE9DKfyJqJoa0
lfTpK8RI7pfG8wgEvos54FOoO7LnIVOlBholmVQqvlhTUDus92NFRr5mepNSGqq8e7DbN3v/sT2i
nRbnxwpi8S0upyYa9ahWfpeMOxz8GkkhxQyASwU/Ovl8oM+7XN3jaB0w0D29il/8azlpjybpCVR4
jJScwZ9PQoNlFS2u48iDt3D4BNxXls6E6kNHm1qh5R0ArtmzoIIO0ahVVvRrbZjptq57QvVNSvK6
y9u29yYBX6Z0iGnQEaNKJ6rq7ShASROY7AjphhtzywPH2rILj+F4MtwU3ivHHry0s8bZ/2Td3Rb4
lfk8hDSe+NtWxvhnyiNk6ULhfxC9Xld0qgluEg2Ba3R9gjVwwatuBxEtHLexDd/UHx5bvvGguMGX
wBHs/l4HbH1rAvUHgQJdEVH4mPZfVGWADf3a2OhWEtzepsfIvf4+1duCHI33HVDBEOTk1ACB8SlH
D2um+mx8FiIywkS1DcZyTbOBgF9dJvqz/iZ0340c817jgdpmO/V19L3Pkm5UvFbgxTQLUK4Lu+rS
P26sRCusbvJxSe5/apM7oxfYGTPKuvI3JDWjIHKhYZLG6AR0cEffvKQaIUF/v3J5BjWj8XDgguzZ
k54MvrJ//pQYwZD+NvbLtbVhdoxNk+V/15wUrWoGR1NxcGdT9gQs8gVTGqalCOtMCTlaTg4ENisO
ibnHrKSx1dZTtrD8QPHbllCKXjWnz3r0kufTAt1gRoDEov/wRsWSBOYqo6D1R65RgURUg4QBYFCI
nnkTQRJFsG3mAcr4++0QQzfLisTps30ikzOgjr0bs7oRlT3ektN7014z8CsoyCwqexPO/fgEz+11
Zsc=

`pragma protect end_protected
////////////////////////////////////////////////////////////////////////////////////////////////////////////


`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-1", key_method="rsa"
`pragma protect key_block
G8S5bs/nmfTg+XZFFeS7vhO7uSBgxNl2N3tH1ifIJ8E0LBBZjm13Fn4k/oaiC7JjqysmJR/cO0Y8
wGSZfYqBnQubHbODw+IUNOPVxb0tNR/yYhhrk/A5D5L4cPXwwDiA6xqCbnTkvVwWQutBYsobGIUz
wEPLEetp6Az2041s+WY=

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Synopsys", key_keyname="SNPS-VCS-RSA-1", key_method="rsa"
`pragma protect key_block
QfWFqGrg75J8XwLPC+EZL1SfmPl2pCUbNxJttxvHg7T2BBndRplsKIbE/I52KxvYWt6cx/oehzvd
WlSxwp3fcRQmVPtuq1ZEQ4OcPvALvGYLT+Xtg6lCJbn5DUVdVep9S/sZJPgzw/a+wZdWlbYCAx4e
Wg9ajLBHD9YAOJ8G4yE=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=17984)
`pragma protect data_block
TiulAyL22vnSRjlv6WIgM8YRvmylxWMtUGmldYGs/WYVLLn1B07zr27CGRcY8IZpFpWEM44/jl4X
dc70Mfk93Wn0sL/2uInwh7xP/19uJNs6T/59LQGRFIkbAU4WpctIVDmkl8CyJIE7BGa7Bf7/KZ7o
5si/s/VRL+5RLAPCiEkdviuEZu61fUtoEflHe9mBPNTTcaOtcvnZ98RW8g520k9SfU31tdmiRGjg
6fN1IkP7r/QiHa8Jva0dKzgelAKNyZgwobfw7YKIurrRPKli1HFgMi5kizwdfEY/0SxCikRmqIRW
MPRbTjRhlZH1GIyKTsb9EPWmwfZ9ubZgIyTWuDDQ5OJ2+9UWpRPt5hHIYj9/JGcmvkS/QRk9YOlu
l9yzdvgRZhwQzntdsGHn1M/qGNXSQroHF3iNmB+VnOOsCYrDVHCyaL+6cU6LZehROEkxTOsYy3+A
wKQGiUbSy+F/ywLJUHt+VgQ73fdJeiKSd+A9hLIF3FD6BHlGFsdEwyQnQJH5s2m3Q4ZiaWIDDFrN
T0UTgqYhgVwpTKWdqJYLCMM9tfhP50dIWz7097WTc1tAztuxWnob/+WpcbXWKvKnSOLRISaEmEHD
OxHJSU1VJgnWYCMHB03D71IMwnanNCTYII5sm2LFShQUYzXq8PpuTni5wUuxogJATDzYqF7pweqz
bDj2K6J8GWiZnalXe3T8pAPMoAvNiXRKYbv6yfC4JqXxAwV6DQltg+6mmOw79GBNQR8F95mHZMtu
jA2zioNHWrP4VA24P4NIJ8gj1gTttpT3EAN4r/2MqPoTTf02/IGM0xPnTom9dTDzcAPoID12nOr8
T/lcT4BJKHCEXQsQSSW9VAgBd/a2CuV6FzeRUFHqkN057f7PFaiSNK+6b+UelMbKyrTNmCkyXpLV
+uxGbKrp5x94+h6qHBx1jO88CofedxPQrBqH5+0i5EnUtLKG0Nj75lkF4dl8Jqdi4uAYkpRBkMnv
xoLyyAN3NB58KVHXzZgdIIfo4d+IwAfWpokusRCMUhlIUIOa+s0fPUv+OmLAj2uvRfl5qnUGvmmh
IwgL03kPc8M8SupBmUgSAgYM3CcyCEPIJUVbd3bDR+hybI+dnncJRwPRYdtd3uJflFYGrtXLwHQH
gKwJeLiCbKsdwc8+BpJ2qZC8vFwKMhVtLT44gbHMc+6JMmiD9wahaGWLi6LtdyJRVpBK1S5lcITS
6u+Tq8bY920ewfJC0HSMqtpPSk6AzoM1mtIFAVAK/B/u2snDiX0mWTRFA1zlrNp+aC6ZkhT+/mKY
fEP4Rt72AqerEHiylwNAIlQarAcpRaJdYi1o6JtdQT9zWmTclXSVW/2mIRQ0LjXY79YsOIq3qgbW
iWXYFJ4S33hwPbpz1EMIPygVIRbNWbbUnkCLLKTSi7EWT5y0mw8Meyp46aK6pu5gYdBcVc6hsV8v
F4KPxNjxplhYSL+uHuXHX2nyIaI3JRKh5gMDFDo7boXGp5RMZVs0whXF4BoZFvwMJrgn0T/8QGHw
b0wW4PZrvgT1R2GLk6rGpj8+UdfYG1+ZUTeFxPFY7zdlfxupeumUOfn3p4zmFMANtUJHbQqsgT0G
1V5H8gZArCECkNOujX+JVJYDLU7N/h7aeIk5Xfg3qJeJSH/1DMvwMu1Pb9/beoeskl5FFcwwMYrt
zlV70iGQAHwv6O46g7V0IQWkSVUxPYTqp8KP6qEucKI9CygfPIFzkZVCYiVouDMz4bvKlgN5TMNM
zsHVp+a4jzbvkj6NaqyAJiTGnBI3W4KmkM66zdvSkg2x3GD9fgA0Ox07WRSWvMsVSw3UXKtXpDXO
Cp9G8pZCUfRLypjRNnFxV5siuYDQq5pswoptWpdtjDUNm/mZotgShAI5s8evP04kyH44l17xd2TF
oIOvS67moJamZi+xaXEuEXEeejkosm9+OioA3UInYTF9g7VnObB7I0V7xapTAflbjWBnMMp2osIZ
AI5lnvmq6Az2+1xs6YbsGrMdwMiniYsxzMsmiRmeJWim24VEH/imMfYx/9farAKNTxHAExymotVm
5s17ndI5n7PH0OdLV2SoM6tLIF0znR+mVuqCRvdYMSAeNHpsDnQX8sCj8m9h5sFt5L/fGHHRUE5j
uD8MBUm9D2k1K2eRaktXyodSq7sZhtu4tyEpk7qjw5zw7TRj7+tBvjLAtP9cWJwE1oqnmrSRPmhB
7de7/x+THRQ9P0+5nTy8ZuzCMRI5bJpRCTqa17xZ/8EoTDJkXqm6ZdwkwSwP1xa1fCI0T+jXcURg
lc6M8FdWeKQeuAldHdey62a7v1/edhVARY3rbHQ9lkx16j3pw957C2SU2pG4+RsTGnTyJ+IGQ432
Vc5VkWKvUA9gVOKfZbDoSKci2fm62mw4Iw1rx8+ewjutkzYii5zEl3DhLHPbiCrIyypXTBoUMx7u
8gKSN1gSvekYazlACKWGSrGF6mYd9c3Xu3r9IvN3oyy0/So7xRAx1FUb2wLhgL2OCB7ySD4Fq0pm
Kun/AkxcQ3Cy6uJ6m9Z29X0bQbvHPz3YitKXE65uq0ZduCJ/CDFjvYTqqLhtODjVfOfrLWvxVymT
jp2NZ/DZl2hf4qfaeAROvBoawJIpb+EFZT21aWGBGw5NfPP5EbSiriYPUFtxX8ZQVJVzRjD1lc5x
dDUai4SeCDvV8m1fTJEVAaEXTTKQ2FJKi5RbZiwVmDkAQ08d+ZTA5Wopk54qcvQ6vueIm/kXxO/D
6/mRsCDbkzvepMjigbEMy1X8ZqzoDu6N/MeuUALUe+Awdz4NuGMvDeAh9CmUYCPTIDY1Busa46Xh
tJt5uxRp+4joYvVkcID7ne5QhAEcHjOreL3ixkNsJL0zTElDm9FDG1M+ypyhODyJKoBzb7X06Cdl
H0Q3xrD3BJZrYYzpxdqHTfY8LsoeW35D+tS98rxaArDj9qq0CVkxsE/xoRiluRkH0qoxoQw1Rzo4
tpRQRDWekDFPMMT5IHF6aP5Xrbcnfkqj6s0U8hHmksFBND6gJNFlKEUguipCymntRKE8Ex7qCVMg
25GAKZ1D15X0TG4S33/f0CBlRab2riUp3+nWGMRdOc9NUdOQpiqVLcVamqboJ4VtLP0QSglzYHFa
mbJS5MCxEYbJCy/3094a8KHFi9et60HMgQ5J9zJ9x1IZODXDszVQp+zRteY2jWBjLoG5lF+3Lwe+
yHzZxVR274E5U3sxOejugIZwV8GNrrr3SCwNZ6l1arvYEvm5bk5U+Cc1kYYAr5ndrHt9YZg+cXop
nF6NtMLj7HDTpRoXQXo+BhVQTBthYX1NNZNx9CH9aZrcDUQkqF1Si+k48QZdxEnn9CwQDZ7+z6NI
gRx1jp0CVKVWezTijwRi6hnI9OsetviVCxYuk9n9OZGPfVy7BN5QHrAfczhhlBx6KY6e3NTYz7FE
yrRuy/QE9ar6R9p5iGi5rs/AlHj7tNK2jfGUXffPZn77S/1yBjelt1bunq/9UudTbiXjbTMyYj0U
xj6bIzRQkWzvFp/FEO7EDD+LtdCvuyF7MMoFAClCwfUN7Tv5QoLwRcd00Kn/QIiEPVXLQh192azA
IHCMqd/vsOYO+IrSqu9q+kbf9k5mTu7VotZFZpQ9zGGYGT5e1eAhhQ5mbgwRpwobgivtCVFoAsNj
D5gMgIA95isBUFnmkAXlwZDvPN2Ny49UbPw9W1ou+pmL/hI7oxwD2wJ/fFYgNAoC/73u+zpd4uGe
UvjJtZIOKwjcK5ZMh+bRDnaZK67VRROb6KFsKotecsI79P4U4iSzChxlQHx5+VrijOL/RAublpob
1jSwJX7bQmAJX9JwyPVg2xjzv/nL6Z0ht5lH86xEBWMRNQzT/xKJfVK5oWurF5RzujCOZ6lr72WR
HSgTn6Z41rOPaNUdbRXtA2k27XKWGH9wz0dD371z+XGwPhtxvaR1cPXaeX+KphuU/ewGuXLrqY5W
o9AYXUaWeaI3l8e5o5pXJyJEuxHPIwvMsPAQmLjRFOmTMLAc/le9Z+nem/7EpeTVhVVRKQukeYwL
/hVHo9kbgTXatBwf08BNtOj5IV87KrNRy4y6GWZHMoS/oKWmgppF6WhxCAkkiYtwcCN9cFKCKAS5
Trh1XEaOodAImFX180oLsVdWz2MLJI/TI3xOuRyCty8YF6u0Pu+EhHzbIOoE+C1TQuMU724qh9Zq
B4BFLsX3PU6ShO08J7/Heep8hUR2A/7Uv0GI/qianLmh6Y7Rcm6uJBbWKLnmOho9VTuReU5XIoh7
VkANR4xTiNooG7epYqToZXlE9qCRWh8x6UfurlbGOm0vpYppTYTen1lDOmNFB+wiCPnX/KCEoV8h
hqUmUj086hiwIpDH4GLjW5V0IxPriPVLBotyfzlo1OoONIRkkm7SFJiz4utphT23Yhaf3fDlB7uB
bfzpC0tucFHtQuKJVMMIwnlJOqbxXhoYU8fftANISzudupPGKrMQApPKRRAfb1yCoBoobwpvxkzS
arUtCAMtTDDuYOKK1fCd+WulXdCvMpFn/f2DQ9P83A1/9B3w7++VZfkHYta8Nx7SkBRthI2iGgTw
tEvwzGewFTxbWV3pzGJwJo1je8TP0yAxAi52CnmHpBuzGLI8eKntGoFtnAupoJUFYNcXES5bmaZs
b2PrOcQ6OGqLZJKxLazSTGVH4gW/xDHPQgN/5aUXeokL0B7XoTgfbzWWRYX+/TOwa47mj/HvtPD9
YWBVektl73F5FVa47J7d/JAqCVG6G1hXMI8Hq0ASfIcMwx8/qsswjpyYN8A4UcM2u5505JFeiotJ
X4nwsUEwyoCPe0iRDGOgDVHXwnLdHe+TAhHT7NWAoUVIwem6w80ZfzkfEdFjIob34X6IhhWxYB7V
u0CuH8L8Ju5d6lO+pFN7PN4S7/BCDyYvgPuhOYyea21d6N78Jn58Ogl5yLiP479eK6RqcCrWGodm
+Ky/Y3LhUvsvjq7dpNwXKsa3/oPsrm14GQ1wIsxdG17InrVp6Q+aOqKjX9TPH0WYKp8mPty1jz6M
kG2JzcbLEmPeMwo0De/4W0QwbDpkhxIHWSbNtHWDRO6zCMVFnFEu+V3OlVTLlNBcKGNplpbXgjF9
8LSu59W1tdhqD2Tnwws2e2AxxJGK+lh31Q418bJXgsX19CtueOnUoGF3/ku/GYj4CAS9ShYFM4+o
mESPuiL7diVMAunSCS+npnBNb3+42Ehmszk3kJymz4HVSmHlTTiGRgChxci3hNolurTXQGlAr19G
np/3aoE74jBdyk62W2i5k3rgQsgoBXB0E4SAjVRb2ZxUuDUnn/KF3Ss1OerXxf45zno4DPIob7/o
1aOQ1wju1WEC7GA1LiIzgs7ibK5X8lo+ERn0DphtVbm964S8eLgAnFgfrea9Qn1ES7Xld5cLP1/L
1iSg+b2QxSx8AZSR62AbXUP2LQhQJ7+MWvjLrkpfbvzU8bwrtNgU06Jj2nr4c9WgMfGNsTBWSeYx
KtJGn+SvBXQOLvkJ6yg/FFLxsZvjEGrmiq/JIMZkQqmQ7SXWpN9GqAWjBWCX+kOe/ZJ6uCkwTVUw
Gdw6V64yc61gDFygDGaTgSRY0b76a/xjlNNwyNN0680NVtK10dlchzeHLcZ6S3eJlS/+GkaH5Mr2
7sMsJWZ33Z5/xjexVwjyzrg/3Bi5+P177dND/qj1c8jCaLhFqZRN50gO6OqC2HGSWHtMTBE+tOaN
xM6YBkAkPCO43aGbMdbGI6w6s8d7ioxoRzOC+7j5Nu7kfI7TNmyhZa/wI4FZ1hGYtAGOqUcje5rt
QVJNgxst60/TXvbHl1tF4PaqgCHOCglswQFKL2u4R3ZBzTvndVw0G20OJz6vPYjFmGnu6A+eVlnd
FdjOeZZWt7DPh5ewvdjY7NuPQGw9mJCu8+ZwRR1yb50B4ItIEL3KgGQ18DFZWMR9k7EwAl6sVgas
s2u6yjMyvTGDNp388kckjHYmFm7B2LEKIYjPozhESwQK6XV5z+VHDGgaxlg7SPombP4aJhfzt0Jq
mJ+B4ffnTv0k1ZNTn3oB9K4PUAtq/X/jcS6X5bXjZaRbnb0E0jqtr/d8ELvx2V7sLbxqAGNinBuo
Lq6ZSiZnq9pqXp1lPj8sxi/GQXLKBfFMkX4sL9Q6KAEp9tcYtBOgiHmYDK2a9fP79Ye/SWv7XiRB
YkfUeFxz+2+txBI05giUYWARJnaGcTueVdkXQ4A4lR4IW+0kuP32cJjtJa2+cBKGUFRcEVVbtUDR
PpvO/LMYPyD+IsTYCv1oxX0W83goR3vtIsMDo5vW/ABodYatR7hWWcBXrV4/mkBTfVZ74SsxPFX1
Mh7Pt2qCO3XlPJWgBATFkttXu8m8KWomZiNsgfemvCal5Hsa+aW3pI81at6anj3nmIZafYO+YJgK
wSP7BYNsK1SOZwQlZpesfsuYB7yAWrfrRHtkqRiVnenWhfRCDlgnyfcsMmua8QhVso0NQ0BUvUR6
SRZZNB7trLnpfjj03pKc3n2mWNtus8IUBGIw7HdNhAKz2IbN4YbBUv+gishP17oAHUL0IIJW7xY1
4btuojLIIkIovFyuPGfKSCJIbLM/njGA7Y+8Y+ZtMd2NCxDb0xyG7BQeHN5mT0fvUIut50eBMzAX
Du/MnOSeOK2C6Fguhv2lTGeoTLBto6Sh6M1ETI6Sr2MSiCw9q0ByGSpDjwNZRMr43WQppqhkmGp8
q/xe3KJ97PrPPx0u/fksnzCBAeQG3BwB+JalCOPaOjciBe5O3fqSIyGxLTIGCQB06zjiST+xAlN3
E48gpfyDpieEu48RxyXAgjOB4IPn1IlaxED9f7yU1IOINOyaUEygOnEagmb+8fdNF8C6/uqMpwfp
GXPlQhER0qWwiV1teZOwfxTOpHbO7nzqlNULsoY4nYzStBYhO0S41HpB33j5CJGPBeuO7OeqNURx
lF1NfCOmvJL+2mKvs8NKgCYkpmQaFv8eQRsejHGmAn0uiWx0oahv+VaJ2pc8S7vv23dVO8i4GNLR
rKMCaiAiOoxYsmaMuXqMLX9wiBl9Bkycd9uP+iuodURT7njdHrFUakt+MSIVZfOL7mTX3pLC+9dB
fQBk/fhCvnLbyBye1A0f2jHrwFGYNSvg4wwiMbe9bPx2Pu+JtDgArb7mY0/daWSnM9rwZ0AZfTnM
k/vyMPuJovVzgFia/yoo85Q0PkLTD4ky0CacaQOcY0Yfv7wXkKoR4885KauBrm3ysiiKJidoMlaK
tvaph3dJGLO3VlMEzVp/aIW1ILUU6Z0v0JwwMNG4XSYjHdkh6q/oXLiCYou2rtmuqVU1VioLxogA
vhjDx6wLaM9KMQhEt+bSYtHwDo2+XnxEDBvklz01Y5vNpO3gnpA7hC99NVI9Ch52Khl0RePlB4kY
2dIQTBp7XhWhaUTK9nLz+Sh24WjfszuSb8hf3TVs8hVwgPYdQsur5Oy5cziTtDFp8CANfVU8/Gw/
WY2Q15rc9paccgzEG+8EAmWyT9aH4c2puiceNF8o984DdrKUlJy+fjZpzDYJLDGzaXNE+JfzH9gY
mWDVDqZDiH2p4rInsyyUJ9AYRxjVqaa+okrxiZT1RSSmN7jTYjlXVUhZ2zwjSfrpnGiYZ9aNXzLc
HYIQEreEVm8QjrzrdoCc0BdZYl39iFFsq5kYroj3o9+IYXLjBOzrEE67o7H+LwVVvBfCB9YW1/ox
t4tvLpMmL2GAhw4z6RVYjq9u/zNVBfo6dnFddxHo16JtmOk7S1/SIvrYY9uuzik6dBWHVD4KrN55
ytiF8M8MR25LmRlXQ24HTNmn1ClCga3lackxyOQcVo1mpTF86lJzQhsRi3CeGlFdhk8jg3AMBHVX
1PlO3WKWEWv7ftplFsIJn8AUzQcjKbRyPozodHEFgr63Z6iFmUdrhfCfTO0ukbWMWlYZ0ZbNSabh
SCDTVxbNUZee9MaNraJ45Rm1Y04pfvxwbkQwQ6ubBa02NubZlWgyizHVxOwC4fjyiO3IsdJISmw5
AD7R1LI+DUv1JFt9jbJZbZxYcmNgXYMAy1BClU/R8MFa9+0cYMe6Q5w/BBYKXscNQ5ZHRsWINyGN
TO37SSNBsjR7eJCacAfhlr7ct2YtrnVE9fKpaLdwRzWmrDdMta4wrO2YJIB7pbLUGK54rWUubzLu
JWJnA82n1FOUGhVJxu9gK9mDDYvsjNIAhuOGuA6LjL224fHjXp41TfhuODFcRK47C87PytIgQZm8
b5ODO0HxnliNK98LJIJfMBLz4P9Yt/XFY/OuFihayTePdUVio85KPhYzjKcR7RVU8vRuHcXJY0Tt
WyZu68Y5OozqDkpJnZVY8Mtky8IaiWcep7lWhrzBIWqnikt5bBiZl56IebWIWGPiRJPenllC4TCV
SKsNAJf4cIE2Xby8kvn6CqMzPSiZRExxRSMAtA0VIDu2FslNjRwrTO9nFxHyrSI+xkgIqzzG/I6x
aaqAlDew9WENUYqT8wXSB0TcU2dW2lS3gK14PwlwAWzTM5InSWAccIJ5x0cppB++i8g/QZ+nmAdG
ZSGt4suePe2YfHGfij5klFeXKA17cmvv3du+IZ/imwSTMGjx69L3WKH1mN5sZCLpflqKERKEZ7wH
DvSi0XrwuFb3tF6kTZTF5Ucyngg2AOADpfEhkdUkMePO5/ibT3+Z/RQCmhkDYBSLUFsYpVrasz/j
nf4d82TCn1WGfTXRkXK775XP+Yoc1JbWpGCbvkPHl6MxJZWiU790qeeYM/hSEoRqZQuWKkgMhzqq
SEasFuI6d4QP3DII9BiGuIY6U7iNPjuoJnjjcNzPRrwdGtwMAvryUDkniDJCg5EHWj79oc64FQL7
+VbeNUOwKx508VvlcDGFeTb2CehQHmBs34SAR+5S3WiYisQ/Y9SNBkUu0TB+ILMIFY4BlnGPgsCc
jGH4zijqQF+RD3RU4NnUgSNJRwnaBw/s34LcLo1lIvIx9/GhgWqEK0KB4M6Ct6ht27Db5yTNES9d
Xs3512A3PE9oiCjN558H5Wo9VwO4xzHHtZVYODLEdSpp7eoT7ExtFnuEMTxQi7WYdii7v5YKWY2I
21HTa8OUFt63gCWnH908Epp9nuFyHbJOePPa3a4qH3ePDzBX+Ozw51k4jz4WOxQE8aorB7EEvVKV
15KA3L2qCeoEiK5ZG7cnzgWf+JH1vc5PLlJ7qeSpp+yyg4IYAL3/70gZLcJKaQv+FJImFPlkz7Du
9p2b6LvEVntD8o+KKhifutJz4r/Y5lWFY6mMoqj7EFPWxP3+vBvKoR6HoOrqW4US/Kt1e/FINT2z
w1D/YT8ii0iV9jVVV7gbDjaAL9Axm8yII9vK4jDxyRT60mOVr5HjV3nd81FxCbUXn2EiP3cole8S
8sXldy0Pg0jAlPDJgGpyoWu1cJjCWgRQ5EZ+4Hm+UoWY9/FHkroSV+tf6gxSCRZkMNDwXwnkC7Ng
QkJ9CPX9x8Rx7bgrOdqOgbgCKk1SkY3iiFBbpjMhdULsBid4cJ1iFhiZbwTtWq+zqDim3Ksm/iDq
+DvSR+cVpKH6J34r6wGm5CnYp0Iq05tR7fxR3kuUodqKmTc17cECQN41KRUh+XGM9NJ+/UemQcVb
+WdqwVPTdQIkbSZ9bRevBTsjJER8JFXRC1/PYQz2qW8NviP8fAcW6zOAAy0A0ELPUGCzGkJ7OksO
QOeb7ljPQBXdhtxsNn1F8SwNu5+IqWZhsXE7pkZ+YBwhqG33FPbMRcY9lzBgdul05aQAafzt414f
P9Vd3/8gik0zItx/iNszqYViTwI4MM3xlxb0eEqmUj6I0cTjtcVpRk3MFppgS3dGMwxCR6Y/M4l0
dxO9VCYBvgmK7tjOlzfPJ1RPw4bF3qdQWrM5IB4y8WN+BRv0Yw1exk9FRjQ8gD7QTiZ5Ra9uHdLV
ehlu7VWGFprTSEajvPlGVcH38j2EbaAOGJEkF7DeNKRf5rp/ZVOeGw00nPfFQAjfeTfdJzpRRpO/
RDNaCZbnx5dOUsgucLLe66KXz9j65MPXmrasescMA9lsjGzDj5OKVOGxArEA3Y4zJzjjGwVC87nV
SuI8QITw5wH8X1CCM6+BnNHo75Pz7Yrpvg0RM8Ct1rw2FSuIqUSbr5XGzanESq3uzg1WuYCDuuxY
pq6JVn5K57kTutNB1zqPTgvwnbfg6/eHD+PvXpxsvzg5X8PdbVRrgljZ9XAcsWZWY8BboBG1ljgX
dO0W2KOfkR9QgbggMw2WltWzY62FGml87qiH1+gg0MOyxB7Z2gyhZPRZaWqWKVyAa4m3tJvaT5ap
tHyXb82fE99UANoHnotuGC2S/BGD95kyzaqJjkD/lEmES0hAfwnRvHhypmlubbcYVlEieEVkOWWX
D5B1RdjQCmmRXGO0Eg65Tx0E5AQ0yadY8Z1y215M9MYYa8bzdu9n0oRMCt/RTOOIaIdSJ3onLp0B
a7vTxKcJ77CEsxtWYSv19WX45Gi1Aj+g6RndZPZuTmYHgGeEo1Hv4T/V/ZBv3kFbOZPlDtA9Kzs2
GE0CuSllk/U1hRCc97bfU7QlesM27Z2na2sIFUYsNQnn1LQMgBdEIsV3uHEGcKJCd/LZFdzGCI11
78xCEZ5E5y/MtBomCSKsik2tNAKP29tdWpgjRlMOqTwm9uCk/K2ivavPdo/h4W7WttAAUEGMwMIu
Qu3/DznbdW6m+auUr1Wc7GUkuB50SfWKmrTVHVy4jUxPYEfMHcY9rE1sw0RU8vJu/MGX3tz3WTrZ
43McabqaxbHNdbfWDe8LjcWfhqCx3n3NyDyjfCqeLQcNxvkm6j9t+VHoJH/Szw9IpQ8xn5RMXeqp
abO4aHDeam2ap1eH3IHurmpV1YLlwYAbsFcABXcWaAXy7f1Aqxvr6jIs1vx2Kow+UFSlseqhppqU
ctFNCAFQA94o8lr9Z/MSGPjS1r1yOAgjlzqkWwwlTz+W9SRAbG3nFzKa/bY9cszz8r9gi9DuxhL8
uxJuo7cWIiZehUk40G2igeQ1bNf+Tyi2SGLzVEer78QWkC6eur70A7O4HxaD05FT8ulc3IHkmcv/
R0dAknJCw9rWtmQDdMmukf0v/oc6e2YG5cNwmYS+uagr2OJ/aKtnQRejgxpyUZxGQeT+np8eUrgA
FM3jpLpBrYeu4TTQqLwGcKJsqcP+6CeLSFwUjC4AwIyttHGy6H2kNYFp9uEoJOZ0ZLe5c5cADyQh
bkK8E0SYwNiYE0yy6rIOdwePz2fAV3GncaX77x9FYFW6bDBYZDEjbQihtvBbSGY3LbQC0hlaOgs3
8OYAkf4WqOV8j+2W1/A91BV+KYLAR1bVZPTc0doLMDw5PMOqLK3pa+IStLFQr54/NJeQpQS23pSL
TinXUyuex2Bk3CCfzzKkbhBNvnkukJGif17nRCDORM7IVCI2fHWDh0Y9YO27XqVRCp8+Q4AjAEvL
8BFbUW0IU1EMvzP4i3Juw7Cknlw0WzC8qbxXQpQ7IDKQf8LVo6EWylvNPiGxQkXqQw1phWgRpPPI
tm1Ddd4KanoILjFYjN/nCKQ1w1dy7L98aWtklT8wZ/WI9sYvdC+xGu8E0mflm83Ay1le4ClK2QBH
l1y7tq/lyLduwUYXBdYiXxn1mELIk3q199pJ0oZ3/InNzzk9ru3aMV8FtI4S0EzyhH5f6uvsTj5A
CDqROiY+ctx2ZEr2oPCcMN2A5GU6poP0vgSE88dfn9octbc0lQLgv1wsnLZUseZhJSy8vnEY280u
x4/nv3TLGESP73st3l0NyQae0xlng6rgTcq1Sn3olzc5w7TPSR8gBBBZeJlF53OxsSq1uLmPrfND
8UXHUiAfoqc4bA84udIL9jMLLCPx/M1ZDP+CJGoIXOaAwyMmrOtFecW/CXRY1s6w4zwPQBUgIwH1
BwwoDosw7KJYl3xXC1aDqBpCHx39VbvI44uAnuwNR5sGiYCjxQFSZrLUpapM5XK/9qm6kUZiIAxy
j6XMlkgi/yH4YzlvjmFXg+14C+8p5fEti132PBqprFBnvA5acei4hHsOglO7I32/FHhPGksHuM+T
pdGOqGq+3ddponID4CmFgugniwzjxTNzBqu+A9boEQl/ScDsF911dn18Efc0DMN4+0+0o3tmfSxQ
NbHa/S5ZM9pPRP26NVpr0IdY2hGWHwCjs+OzIKfuFVwp1TOTBzZM0BD3yKzaaEJcWU+A0rPJcmWt
X0ABBgq7xN6+dNB4tJRQN/zNUpDVK+EFO9+uHUvjp0lhFkkVNeIXIcWGJ85R494Bj9mfsS+p3Ay8
8MUSJC411Fx1DbapJnNtCqftYRHVviTCbOhx7RwITYW9BPoy0idp7wxk2cGRRAasvDnafjYSPs2V
RlrCrf0RqkRJDw/F+718ld0iO7mzSE3bnb38Us+PxUdtaM4xomgQna72Rc9+picOM4GYbd29+pzF
tTl9FbifzzEcs23P0wLvVlkGNvy6RLLOI5/xJOSfvVrBsyCzzRKH4GY8v3tjMPTHLzyVWFoqjwR5
jmHP0ADhxSHZZxPPx7FPXt7LZTfkdGUImoyG2fNXLmPcm9I+E81noOJCqOgGsU5NOzuSdxmGs636
kOWBBFqQHe5P2fnHUtBDE/m2GDG4cjNVDeMUI1U/vRlGMvUIBa3xs4nkOPajw/hcAD9Vkfpam7GY
ehOXiO6c03Eqa3ySM96SJlZyh09RPpI2F81fsSfxQDeSOcneHNeiNpjXcQ877PvgfqjuZtU9UBTs
BWwQU3PqMdcbVL0WDobeEbMc9qfXk84qN665y8DDdoPEYCfMuzSdPSZb+4ssiQRBzNVO6LuZF6sK
sR5edOc0ISQkm5U0B/VGYCAHBpWru9IYzAwaWHKzwdRs+BcHNvDUELkxYIX6AeVjHqRj75SI3+X0
cAvg9cTCYMTMwsHGjp+FC07nBOupWzQPkysu6mx90pYSF2aqrTWJsIu+ft2S/LwZeUZI08kuwa9F
1r0xjN4jnpde7+4dv7Q14HUWVB3ghikAromUoIGarxAxSDLgL21FUtNAqcNpdUhBXTNyR/ZSm+oV
shBkXbMMTsyuM2RBmLSf9bR3stGDpPZtqGjfH+XYQLInoLeJK+m1PsUHvg4g3OWs5H4HTkJWAZJ9
Kas1W9rXTLYCPA2FeGVCV1oL587XZstidiuyaXSvjJpkh2PO4te6k+3Cj8e3Cj0oVhUJ3l7JcV08
qO6g+DjAsNHcWvDX3YLQWTfEMlPZx57fkBOgEWkM7ySp+rpo+4C3lis4z7qrVhZGa8fb49rocj9G
DczytGxmEAMRlStl68pUKbAzrFxNsgVmZl0uCSLjevIJz6OlteZDvRLv4N1DayGG70fwng+3ZfYB
PiU5PeWMJTOJusBclel2Vj4/vzRXpyolAYiO6xNtCQjaAQkkivw+Xd1U2Y/ChUKv30OneHjHw52I
O1suGGdjYxPp9a7svXtt69XHbL1WN0DBnD58ae/LcHBp8O2lvNiLZZXYPAxZon7QXRCvacAOymXh
baRpK3k4NxCIVl5+mJtlck39j2BcNXrmnSGKaMNV+/QmAK0at7ZhuYhkNgLBui/3ZsaMpoAp9pHi
E5pUW1V+UCB2Gc2MiBq+CpwWuMqIf5yD9hA69UgkQAPXGuW9FqQqgAF8HXytaoB5eAJ3uMErkEQj
OH5DphbyrsGcgOG8fO+vgs9yYUfY05lbAvKHf0uKH4DzgR9kI2gjC17O1aD7J7LumyGWXo0DbEET
j+r5eU2xZdXkm0QiDd6PkgJQ7rfMqnescrxEdVNiml7ypkIrXB75X/Mj2Ci1PjXrLMZ8DPpJAb7j
s6jw4W4mszNVO1VMiTlonBA0TxtnFaqKdO74mdEvRJ8FKsdOocJ+x6Pcdwz2kOFkAZRCvLTtnIL2
drNHSwOe3lsv9F7UujQ9D57ZzW0Nebqs+3wiHgjVpml/Eq4RUTBLMhNCwta8rYm3eEAnlddQxuon
QEhq2t7ZHmKETCUgfVIq9mX5CTaM5nXjU+S5v9Jdoz0XTMXwZ92At8gVjzUyYKiVU0B8IcIt7S6a
Dr2q7b3BPmOPCh/P80yhNxQm/d2WNdKZVUlyRUEo4ffWZkm7+8eDz+ohVKGu+9W9mFTFCTSMWFVE
3QgLww/hmEFEE+QDifGIyOn3qnuOOmSCS0m+bV3s2S/PWmF63YNSrgVoBRUGx51t5d7NUmbd8wmI
k6PZf7QCfXpKvyjijZMjp6BNjDyGPoh0Z2suxc5m2pr80LHHEhWMFWqiwrrBELSzvbmSKhJsol9c
vPFpWkbtktjTPYOQlpi42lEHQ3lNkkmf2YXCIfCbFzE6NLH35hzTPG1Pl9By5GASi1gaJLYwORgK
XIBxWwBt25CJWoxDSXq0uptF6xY8GwZ78S1CvAltX2aPn4ba2C6Q5BknsHtNheVaFmwTMQxfWpgj
GITJPzX7+w94kI9kfRsWikoY0Xrwr+OHiJhpsaGXQuMxkLdWmGyNE3h//H6MDNvsDyxGxv59Mf3h
TB3/+hVfLHn7fyxgGtFxrOtjm6c/Jc6FzEFpBKhkf7uW6FxFtbEZy6CI//mkc8cSTvAQhu+e5B+p
HXRk22NjyKcwsV6UaaeOiLaGu0f13a1e14gWXkD99R8+qxNSP/S8ArkWKJ38Ri0dYnoFOtxg7gpa
cSltIrzCES0p7+j44cd88Vqb0CVj7m/jcaZIoE0RwbgZMFMM2BIxnIG9NRlA3oZKFWef5V6veopf
qDJMmYYECJ8KXudiKluZCLB1pIC8cMzCfi8239nmmBXE8tvAQbrPdSkEKAfiBZC2U0FdSxyE/Q9P
gnHCgs9E3Y8bvNtBUyWClkmwj7NpLvyAqO6qoFTJXLPlg4z+l8k2bUwooKyARxR7Dn3oUrSNaodw
4r1tyaWGyfH/3TTbx0PZFMxKxvn9Jcnj3mChnEne5LyWm2uWywr6EVFy+jr5/UIxTAWVv8SYEQ7O
pr37RoGQhoQ1+EnpsRt6xRC6MaQPUP2CAY19Fk6731hfBoowYsmSS4iMLxDkGRgvE4zkVtOQbNcY
B0cTUVwpF9nJGFVAxhsrd63gNdpCpoGlEroEo/EjYHQeWfM7bJTH7bUXMOuPchTFqOlAY5hAFsqb
pYT2SzjQ56XqkVdCCVAQCUOssXecTzh3WXcqEoNS4gieuO3+wE70ljJZQC4zuYjA1wXif3eFIJrL
NWqS4UEP3fkhkq9OS5s6ZV7/w/Q4PgZdEaxldyZphUpGHb54Pb7nPBr7Hk7XlqoMnv0hva8HNOD2
XJ3h954tS/40VHkta6N2EYW/H9DEuDRp9//lfVTW2jLPS1KRyi2znQOVeOEpRpORoBorOseXjz/5
3g3B2fyyb1+q4ajKwl1sUEEOTozSs2+sjJCk6bO+FH6KcckhSR8yL+3x+SRU7M/mIIMOLL/1ID61
OO93+QSdTjf6nUPT30vKd/RYRoiHPxF8KL7zWW8I/WMYazfUqdOKKy7YEknpJKKxVRLZfLRLvvn7
g15xMYXbv8+5c+ZFv/Dvay23lt7RsmFW5QQ71OZqgx6jI/20AtwfqAam/uKGoNnWhj5FPcd61Jfc
qOH7uMWYDEHgxmQE3UhclCfRNYHQvg4KKfWwi/X/HWH+G4vlQuE9CtGumcQo4m5nrW6dnHiAYPwp
oa4nNLL0LzUYmPl4G+uFmaUYC/yAgEWO7tuRgBxVpVdo9v4xCFsgW/V0oV/2oEZxb7G/zTyb38cB
fJCJj/h6rMSOjd4ULS/VeHIHb4UDw6LHrWhQPrVc3ZzMTtetmH0dJ4gIoDs6bmi3KacibBnbU1vN
6Bb+jy1p1cdi3YpibmniB/cds0UZW+ZmVCBNWE8z425MYDFf+co6Gkc+S+SMUrwoAz4+wwIUevhB
ZfPtDv7T7fNGPEbD9hllPA3MDDQ+IpEyj/IvYnfote2AvGahcSAvwSJH7xhh41qOyI87SJlMaqmV
Qon6L4IIydJ61cZotLCbA4CoFXS4fBiBH6PbReNUJYiKB3n1hhoDuAkf9pk6bjyphnq7ZDUFGJNp
Q1M6hOLtZ86cdNujSNmxQNpjvMBNOywYVwL9PeVZjXlhO5IO15v2bxm5avENz115QMR4pg7YqQwJ
zApGnASVfezLkkGhk6hCqZjp+Kow+6HDR9EA6iwTaXy8rbaHtIO7R2YCaPF2LEdCW1mvtnJ1kVY5
GeknJQkXTXAOfbi85Qkyi9VTAm7vOjuaFO8rouEjY+mxkiLDLyApNK71W5aRlnWBqJvIs4DkVsS3
dbLT3HBSpt4PsqgZVecxbdq4dDoZEzL1FB7hhkQhq3VwtKj/UFlEC6BhlXkDYZ9mDHHup+tMT7Go
3w8XOGqVApNwYSEz0wnJ8Q6ImxsZeDOjOSRRfueviIG4p/bhi0LqyaZDclU1oGoOhH2d+IUUCv98
RW8UppUl98a0S3LpLjIb65vFBwxqG4ddrwLlpUeYUQ/VJ+7CI5kowG3mHvW+9Xay3zRmu/N/QEb3
x+KkIhvKLhFgyXsv8nZrcTV8Eq8DO0n8w5eqkH/Cp+jhgb0c3O89PjjPolVTfnnVwXCUdJlfuAAG
pPdEuObS2097e0KkoIK3r3mr8UyR9erNuxFRY7TXmbJtx2KXl+BHRZFNTJyRM1Dh7cXnZNE3KV++
dorfv0MDknZnpY/lhu9cVxzbdOSWfBEvOnEIrWpyulIkOmuVOrbfqXTa5PdDBDuCcNgn0mt0zglm
GbFEePzAqpBAHSg6/B0nKQVaAo9ZYHfAkYqndBNQsDt82EkRkeSSDU1Z8GAWkfAWJoGSbje+KvDo
bcpsNf/TZk8awLjVT/uxRgfBFfE5Acxdea+S5uFAa51DqaTv7Sho5jzwf9NCJmcIWw4zJEMc+6i6
Tb67W1kMAT2GlqRLiGc4p37Or6Y5CBFlP9yu52157Vx53yk5yBzK9SGs4LxaUmc35OU+CgZvtv+Y
C9jQQ18voG27dKVhjTC8v1q1SPeLc1o4MPnMtbjg8tDzHb1x4vcZiDLh39GwHrap6ap0FZfNQPDq
DDWJdE49kbtYqqrESG9JP3KZWwqbO04B7stQdpAQUd/5ipyJKzihQZAgAk4yZXeYEknjg+VL2p8y
81/dwJJIKDIS7enJtDMMtHQoH6NIMuwNfJpcjMHOTpObtTrPB8cmWnXdyqbJYH83dDECGwkQY47i
XaI1W1FzJf6f23aCO5eCcTxM/hM6mm/Kybqpabm4Wz4bPD5PWvQeD41srRWbUChXPTJOR2NA2knC
SG5PZ55ptbLaEKVIIymnuCZH9FNIADAdarNWwlYyXxezPXQV8kD1OGUS0mIT7SN+yMRzD49KRldX
OzZ00xzsNKs6sS//hZeIfSAX+fepYlu3+NaSjM3yostS6pce5A0tbutzYgz+6EWBRHoEVHqILQ2p
ZWOPgAt+9mx6viKlPQnRTHSYcfqxKHsG0QPxg/1zpsM1xIr3dBn7StyNvuLEmWTACgTqyuMB1atY
zDPmZeI/BFaMy+xz01JAkjVKuyQ6GfIfSgSA0NGxDuUjjJdlg2qCxwWGkXPKZPa7o8S5kSNj5zWZ
8BUm3nH6+pWSRPTrtLc0VJxI+MUcpqKBXCOyyN5JCIVnRNvy6mIAU9x+14CMdvrPFxXXav5nPWNT
fGKCStL+vfJkC33URuw5eovB4jilP0suLxKIW+YHphcWinAX7um9ug79c7HFOeoaA+aOVO6G3PoO
zvlXvLjrzIxuz9IaVeN94p97706Qb15ZSCrl2U+s3NA2weezGenA6XLByTLcDJKDjXIs3tmAAwaz
q79DLwKOKCF69yFS7i1lvcHMuaWR5BqQJaOUGOee5H+rcpStBpHNo/a6cMsmwqe20Ib5Q8N2YBwX
HEhnlfWY9t9EJ4SYgGUuB2zDomYmWTtkMgrc/SwvLrqKKAeOvTXzhB3DE63OC7ZIgM+HfiVkDZk5
ioFyeBt8WCnsLR3BPTf2kHABRjm6dz9BqsT1rPje2HVNH5pHnaXrhQULBtLn0g7dNzP40in4TaWb
J0p1oN3p3MGq8YXtw1eZ3uqpkBHRQaeqjDFBYyXH3CkKyzFjQmilUj283xqay7Nr1/qE6J+QFS2h
iSrpxX0pvSlbT6OHl6wOp9YUSXsbPbBaQ75R8PaKhtI69g+0KH8ILr0SQHjzIA6NgPsB07X3wgqD
TZqafLTvMMmT91v7BXVRAP632KrmzaRNfqN1lfIgustxalE0oFLd/UNO+t9CP3ESFSlpbSXjEQ8U
XAkBhl549qt/id51Dy4JWx1D9TdRu5+aZCTfy5VXNGaU+4zu+aZUC1uskSDOl47c6ATg4Aylvcd4
eod4V4sFMwIZW30okcEJt6u2/Hj4GoZLknSO7QfcROeAo1Ep56UHorMPzEgdeFKcfRJEkBK8kwbC
GguVetql+eQSoGkSA49QzSY6fm6EsXlebV5O7+bMGKVB8gSBxCYhOdk92u3W6KHegdRoj1hV2ei7
eC3qL4UUnqxJ4C73lyEyIodE7Rj2aAInUhI6BsAhy/IpkOoTKkpbNZ3baZXDV0QcLq15X3+WLs/6
FRIlf9VBiuKJBqRZKwSCUVRDofe5lfVbCKHs0nX895DW2RW0SOQWYRc0u0xPgvu51J91T4dnBUm0
RWi/umZ0OA7LOh3xoSz7EGscydFliS3kAL5us5X+PryjBBzKtDePNFnG9Fv72pYoWgDOwHa5Fup9
a1VkjpPaZfaFaPLWV1uax8edbLgk98364Rn7JcAwvApejZtYmOXg3VIicd314NTOT5M8P3inzoWD
YmDCHs9pzXPvvYlTOuUVmzWpuNqvqDhSSNIXZkCGn2Jn8GoFOiGCsHz+sKi8APUbrIkvztqoTeR6
xYz4I7QT12m1bP2n/6jC5I3dNOFk0wVpR1JisYj/Tqs89ZHEdArlmzX09x4R3HKDjCHlaO5WS/iz
HYLwIF7cr9GNM8B+B9C5d9FxyLC60Rj42kt2lb4eaDZCsssS6o5FNJiKVd6IRTVlpAuDp/Qp/L4I
EQdRWwDzgqx3sagbCVNaZXTcqNUeBsynE9kQSiRR+71ZsdMIQHgM0RwWVPWww4xK+mLptNfy5I2Q
4vkfPdulsYGtUVe5lz+93CFR29R5yc+U6lFIpNhBYAPvPCtjVZzVtQ+Vp9k7Hwj2e+itizzEy1J9
8Q+j5piP1QjAFy4OOCaAE55of6bFMakFLSNvdqYJJsmqIaoxSl8KB5txn0F8bdzrtvEQckhagOeS
VOXn75V2PcExvgZIW36Hdo4I17pLML8CNNs2u08AlMhZRHf09eVy1ZXw70Ok/0pl3+Lj76fAeTRb
iSVUNXO0wHVcUTUYE54autkW4HhuHILMLyZBaVLL+iaiHGQVF4hH4+trdNa+/b6DFoLkRnb9ZXUT
aALDcLPfVfmhYRyB9JaCrZz/VtpRi9Ilcts092yElNypCtlW430JnACU14TcIErUpRcqj5F3roBt
sK5l/MTaF8voClun07dApc+QcJv7361M49El9V7e20JVZQ9pxcOaSjD9Ob3iyyfT1jEdTmoyS6zi
qLetV6Tw9Nvvfv2bERz6jpScG5oE2/w1O7ZGUA/eIdGbM+/QIsBR1czUKN1vp9GYi7OR3xfVlyZ0
dXixakFkKW4ff135UDM0/i8qWJ3ghDFjo39J8cZD5CgO/h3zgtfdHaQPNAVTFWubXh9kLQhkeUUT
bcUvl+gjRD5d5LhSgDWI0k1wwh/z0jxMLKCmPRZ1QpkGrPR3KpNk3EOxi9jnDm7UdwUDeSjEe2Vo
DUxWMbc5JZBVFq+e/UdubkSXb1Sp9I4rp4Fy+pl+CHmOjWiek3vIMr7+B0STveDI7rmQb1qW3bNC
qlcpO91FpCso0l6l450nuDCqfzDUxTZrjfFfAOmA3L89R8K6bXoihbtyjax95YlmZHe6oedVas10
P8N9RSNHH7BrEH9WqxIa6/mh3wKpxmO6+JyHfT4Rffpuc+M2sWr887ajIWQG2fzk0v4j2IjAn4uX
vHRIIzFCouozuRwUEt1CJbSlyjTNKOZ9T478IixRC4+XO0yNy20xOvqDpND6v4wLNJVvDK6x568x
nQmKznJxPfOY+v8N73/AqCsXigyJnMHrIi0IT8NWHE8OlEKxopZ3lwm9isQp2alxqFZuyHg4JhmV
+433XY9P5iuI/IIqHTNqDwoxa+aAoBlkwDn+t9YfK/4AyiInC1gdZAXOrbo/fXLif0PrZ7mnyDiy
afvpMpw0JJA4y34SDh+US/Mya+ppfWRrQ0abyym63chNwxKY/GDCiKD0x2s+oCDNdpXBXBp8pMv/
oQ2NcPV+JrZuTtfzPFyl0jYwSqRwUGcvBfi1U1qjwlyx1Oj3Sn74S/NU9mXb1r8P3a7AlWy9RQNH
prydknSBPDufE3yD8TcdvU41z7FsECBObxIVlJoakinJkEVKD6b62+8HO2z2Nok1F/h7DB6Sz9C9
JEMZIlT+dO3toyNPz2vCkgpEsgxVAArAketA5dVFO7l3GR+INbObYGS+odKbiPYex14+YHgr0WSs
Vlq9wTaPUJ7KjmcJYky0BeQIRqEmFCpOnPL6hl9LNHKUm1zFsRgoRpq1Xm+GSo3se7J/bZhfWsR3
yo//L/DjZ33sYNGj7SIPAW+a3t4dqarNnWLAwVQ6pWkeFIAh4xRSLDQdEv1FVygDgXj8yDmYjEBf
2Stl8L4WWKDSOD6ROV0VI3FmAVneCWKdboZWyA2aVvx844gVnHeuBui9+gv6k5Pt29mQSX0Cm0Gs
4NwnhiYVR/PGUj4589fAYo1lYmetnkCFm8An/N4JD4aKcOu/Thv+2CaHKjOG3JfS8f7yNuQ7elPr
v1A7JjGsn01Z7pXAXkBHlxCKwPJC3tNYCVeO1Q8tRIJRXpIMImvvbFZpA2uFx8g4K06agflaRMlD
EJ/3IA6puwFR+tuFOngo25V4tuKNbHtBMewwSi4n8GdFuhEQuBgkK2meBj8RkC0UhaNnU36rrU3P
skJWMx8+f3oN7ipA3yUvkKuU49EpIc+5KAyOU1CVS2m7Nn86T3lnNxUkvT4xpqHtQcqK3ljV3e/1
H7rRcDMhJwqxKvVrtqJTDfeF6u6nC437YcIZ/y7nn5ufIwuWcVJYOSCDEcHauP+SSr3cLgr3pAxi
zkSkQtoEH4xUS4/Bsma06duznHmb+BaT5oedLqWmko3mAK93s2/2wRrnT6ciZsx4ClvFR8yx5tcV
IvCAvjwFLfRVFsuC4QTDSqvzfffHdwZnzEbrU5/+x0OuRTdKW7fxhzm0Pt9iAMKbEvBvb6C0vi7U
06yVQEKo13tbWWl0Kjqin2fDegEd0nKND9E3o4svrvODOKyhiGrp0IUUomcWhzBzgkxAz4O0ZAu9
4mmSUiUGKnGK5Ias2N/6WvJN4k+VKHAzCaz/Awja6IQEH7TCq0jgtRa7Q6feLn7R1Al6hdFbnDvI
ZL8wyG724LZN7c1larTW6GotuLV2RMMWFvsnZST4T+i7HwvB1rq81n/Dewvl6Qr/Eh/AfCplsIQG
8zZnciwexgdtkEdl3WbHtZjZO+kg+n5kpcZ3ShEBzKbzTk+gQL6r1XPn9jT73eHwTgMnXnnvc2TX
wwoINv2rmfMSKNuWJtmxycgOXf+uXwOR7wz9tRykWuiXhddO7NcstEy/35x9CmJD2zzmvdqN/F+i
VYPpUT/kk1BVC5iqHRW9WOezNKbs5wvoKg54TUF95v3gyw/0oFZTH8zIW9lSGV0REKjFvm2r9B6j
rwUoybQokpEf0gy/Dr8V7tWV0VQQ6taisNIUc3FSlWXNr6EkLf6/26HgSyafFZ9bYfA+16c/Sc02
wrDbeEOZQI7BMtMNUiB56qcwewuOgNV+7Kui30/RsmALrZMUxfIlONRAXQuER9yDcm0bTJihmg7S
gb+7Q8reD07+prv3Kj//8ufEWBz15ansOM1+SXHnmBJqp7FZM/VPaOxs1Iph9dERbcKfu73nTSCq
kIAYti6TE3SglpeWybTYSEhVJlGD4yvC3q/YHaldDBYSi34Ybi6EjAVQv9Wbj4xqKMuoeD6YALcf
O+Sx7w6jSlf44moiPBicF0wSegVWwQSKDASTzYG1p4u4BHydZr2CfM265XEcfGIZO1GW5DdH97Mu
iCzYKlxM0wLWYKKJiYLTvQ7LzRSByCG2nT1V0EHGQ2jA5vmFpt+L1RZv7gXqzEVceMD8ewcslzDq
ffzBU/jOgOeG/taq/kJ9RSC1eQvtRd/Tqi4X67Ql2KUiE9HFQ1y1pznXd13Nbgqc3mdZ+HzJ7bq5
4a4yD2I8vq9EIt7q1O4FazOfpiS80YflDQxfSHph4LA+QC2CQCLIaA/TNyqnznHJeXLJ1P9oZUqY
JBAtCrmjuGn5Yn8LAKn7qBagW4YoEPRBGZlXWiyXKpKCjtTh+rnJ4i1CNofFMuN180ZPwRkeoRA/
5BG2y4YSytRxACUE2nWDwEg61EBc9hGNCqyhinw/L2vZxpPdjUIx8LtE/F4hdF+yoUY1Aq6pk1Af
Ty+EsZpBN5jPRv32+YCOEczVyoOD6TsU2roeCGexgW8Lor80xjLFNkxROhKEGo+wLT5Bv/5zNtvD
RtdE5laVWG3L3HreXaOGHPw/uHk9DRu6c4509U6NYAFoCbi0V1ngIdtLLxDApCY0RNT+/h2dRGxP
CWDncj6qPYM5yMP5K823SyqyUljUNfT5Xx60AvJsgqo/MnRBWk1aZFHaoIQGWinW4378TO4IFlKy
SJ32s5sqlXVOzEInVqG7LTgfG9k9y3zITIFD62J7mwx+YkkE2GEGchf/iM8U/wwzWkXjQuaOjWC0
ABfIJtwhwPBzVnqsZqPJ/Yn+m/kdt5/XwfJ6bdPeR400TcArVGWMuMqYUz28kcTlXEIEA5HfT/QW
B/YC/M9yWTAfiGalEGIcRLHxb+An87uMP6Ss/0vUWOBVy7EjebpJ0yy27QpTNWfTcahr0pKH6gJx
Lx/nAVFoI7QtGpcfWRrycv7KsPzP7l5MCrTZcCjDCRKSY7rUhbLSloa8HlSyZXUQOpPx/pR77veh
eRpwEnswqtjGgfmosE/6hnTmJpLgOqGs/M8LCQRmxSt+7NPvMtkbf3WITqjsDe/PvVaJTUg1/QrH
mQvBI2gUeFtwRWzBFbwjtUqK5izqHP+q94zT/mYiD7WVdgVHMNEQBJaTr9R1ZrVZzPwQEUEu779W
iCxYYhiB5MqgwUnYWFP1g1w3NmuSGRKYcImiKH1wmOUVyHK9bP7bOoUxZQt7alnHmbe52zsMLqNc
J81Cl25SUeAS6x12d+BrW/+VB4qV55WnWEpsdjwvcIJG4ju6J7HSWuGo2FyF6YchU8LmVZKbkHa3
KD2/MsMYjSL74mLRJ+FZbeq48T6oFcqDi+mDVvRDDmYtCKwkQap7CwO+5x2THvqNgj2srDd0gCcG
PVQKsP4J4a3vIPebBnYHVpHPxMKkAjjDiz5kXqLPWThMk3ZULJzd2aK/NPpMRf29d5plsSIKfqA2
xjkyL1uRxe3Pdn1ehPnb11It0IS3R/L9zoYRbkDMbG39tKOoDoRJaWBvEs52qcAjtNi1ssjcIOHq
PE1sSfJ4C/WYW82GB02FdFP0YYTIbgYLXFW1zihEkVGIA35Afi7VyFkjUzkbmP4uhV5veSMw4KIk
QEIF/1mimRybPaglj0J1CPOLBvqH+zYyzKAnG/0gSYxV1lX6jcoWv74LOsj+tbifYIUFS2vC0tBi
o3HRHxa9QnrmGpCbGeoSyTSt1oF04BdsKJk5F42q+slMZ2uZHMYIEfkAFQSSXpYD6+72OBCLeTee
kIQMZaWC5WRMAJ+4vE3fNjilUH8t5bf/HFesSrRqdiWOHWx8EHj8suHpAVHFnZvGQcbs3mcMko1+
9a8SLhtFdLrMIZOrJsg7O0VazpI3/vJ068WTdjLHKdgiqvMke3MjfgiGc/yhZqh7TGRq/6W6Y4lK
3CxJBTjJpnkaD/oacEUGoGoXRX43WBSTRgVYNk909RxVPfORSCeDQCsHjl8hmYjh3FDIMxzhJ3Yt
9xub1MU7VvLDzJidxtmv3cK2Sak+3bqXyWNGWgI=

`pragma protect end_protected
////////////////////////////////////////////////////////////////////////////////////////////////////////////


`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-1", key_method="rsa"
`pragma protect key_block
Ic8VH1PcaXxI81s2U9fd9K0aHxHrF8Rk9kRTk/sdhr2INU+B9/2cr7Y+uWIPyux6FgaBbN6HJ1T2
Yr0Hq4UddM9bU7wjWAFUkaBdFPHgf63BKYjsULv6j4L56KaX6bvf8PYItlamiA6lx7f4gpOSSjgq
tsMa/KepTozCEqjfqYM=

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Synopsys", key_keyname="SNPS-VCS-RSA-1", key_method="rsa"
`pragma protect key_block
q1APcYx/QgKVzUxsXjhV53FbibM64sgE6ThQiKryhPzL5OX6IW8f09T25WS06KDAUeKDmjOp7ans
hnuJOncOeBh05MNxpypX0m7WbPtXs5vPXk9Hq/Sxj3ShXoVWugktyYm7XBWPPVfhr2ZjrD6tPk6R
tk6J8bvcP9yRDNtAnOs=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=1040)
`pragma protect data_block
MutUfOw83xprhbG24EwCmq5FlEGdhDOqDw0wcnTTszQMmhr9/FRUUbGD1SKcAMsqkbeuiUW0oZ7Y
MxecCiE+RkGjGx7FX0VPG7pmEh4X1/sHrZ7/REoo0vg+Ks9EGJyeP/DlBJqSMt9ALrF0gax9Kp+4
EWIKeGPxZjGSzQMyihQI4pBBfkHqmPVgFSYLeDc89KFkiKDXj73WgYxWUuavrhjjxm+GI6FmYGfT
PkwlJexBPQENChuXmimeHBgmMhOLnfcgjk2oNnOMYwXGCtCjRHJdTsMllB1Eo9KCUEUzYI7xRI5I
ExBVkM+0KwPSDhQJVAL/fjPIJUBrY8D43xBFeO7e5m5OxR4cbP5HbYBQRPKWAzkvQM4yrvKdT+4P
6VAAuCzlVl8+zuSAZkvZsSfMKdy636RJWvSxOnlaRUasuKk58oUm4ea+OVX05vNHVgIphcCFIri3
AGGY6eQouYoUGU6kgKwq+W6DcwtosGT9y9cnFNYsAstD3NNB2S3ot56g0LBR3ddSjxM6u10B9V28
sH9zhQhLYkwpQvf1228BRj4KLcm+mqhShXpM1hNZ1/LYh5wkIMfV0nVgfkWP0bbI3JGGQDMgGdbb
HM/KO6pzvQobYWwzBBB7jGKtjyrm6HGcnziWL5w8T4n8bDUfv0psv4QPonsal9YzZ4DzYw+FVGsk
oTD//yWMDaHocNFX9hayPvue2Qavl6TulR3+bAvDSTc9Y1AwcLZ7Ema9+s6ss2nBEZ6A8L2h9Q7C
NKKoKyq30nstyudAFyxkwqZ00ET+FY1hY0aNvCYffZIuz1F27Cao+SVLdIcgv+O9b9mMTyeU0aqA
xWhD7VLbEk/EzprLJw7qyOjlhrOkgAmT/5H/R+2eW6hNw4LfHv0rCJlQNSGrB7VEkOTG/xaVcYyr
UJ3DVthvi3kHmk0nNJsU1LEeMNIYteefQA3IR9/ocaDRYLTBBoUyTI/eWWQ7FvCNVWilk8CNhZ0R
TfAOyQj206nWcHYd0djINWAnCSkCA7q6MECfd4bQS7sOeZr+pWWLqmIuSjoGW34C+tDz0ctw4cd3
hhDre9YVc8OLWMjmjkwZgi6OwHKWFrIrzbmh2WjhkrO2QkVuG2rQmigbbAE8iJDpQ/FZYcbazoE1
7QU6XJ8lW0mQQ7zQRDn0PROeryMtwIUZZt24shHS9nVyE3xPeac2Be7iZ0XDvtdpWqP5hltXJs+y
ByfayaKZ2z6MCH/wJiiyiQdPC0scLimv3tgnww0niFy4PeEx3YztrXyWZeiLFWixLSHvg/YrzYU+
M/073hHEU1OSA+gHFKPAdnKx6FtbpCQm5xrjchBjllQrsJQEqFZ3gx1R97Vgid72sAEVJQafrNdS
1aTGGQVLmWODKuCbwMI=

`pragma protect end_protected
////////////////////////////////////////////////////////////////////////////////////////////////////////////


`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-1", key_method="rsa"
`pragma protect key_block
L4yiNGDl0Is0ICXT53kha8kCkv4zINp+EDY8Q1Ohl2eGayeFxDxF0VyiJE7Iec8hrXqVMxcQbEY2
dVn529h9bWkTStZxCoDYxJPQYCB0f4xSNW9GcF512aPG+CzLSVNypR5aK4DgEu+V64pPOuNRt5/7
EozP90gdoWVS19HCIag=

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Synopsys", key_keyname="SNPS-VCS-RSA-1", key_method="rsa"
`pragma protect key_block
nwYSkwPHYP6P/L2yaedugfAUNa/bdjK9PHq4kX+wn9AwFIvtJxQPJxryfMLMfmuBENKRhZFwxMSy
vsnvbaY+KGQmfPpLSThXBkC2g8YrA6b4EkekLaj5g/wUCtK11MU+5NruUGCEL4H/ovLlWKUCD+nm
cvQpb/MCbx8PwPXFJK4=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=656)
`pragma protect data_block
zpzBsSmcRLERDfyuwTKknk23mPMmi5uEdAuHBGF1YFgZ4NSPMUXUZOn0chO243VwrdX8na9rv6aF
bPli8yoKZ7hwLZma0nvMQn9E+JACnrT4RNWYgrkIuwV2OUhU1w3VqnGP8i6/OSqjtVeB5LLDNpba
9BA/3trKxDo/lGGvxsvhhQb+AHkYHsOUmB3kHNhV2GDHFZjUWPNvxONBI6WJV6c1P9P6C4bGi6tR
ex6y2UZQcGQ8N5MxvyDzUAV3xGuM4hsjGGDoB9exX7yCn9Z1hfz0u8URb5g07z11HhT+ozsAi4tD
6qgkxtiIujRpAkiMIANdejWYpZpP2teydbmIryrT3lAcwSnKQXQpJbJv8LGpSzAyNcZLMknkUoRD
n4k+ENOyZBAZEO57N8KXTt/0yH4LCYRcG+4CrAf6KXa88y/MGDie+mTHYGfceDo+gXmdIupZ1B6C
Uuaq0UlKI2rduJr8YxJV0pyITWL3Z48RtQI1l6uo42aeWftSJSecj/ESUt1wdbdA394GpPKmRUVe
8HeHody66NhmnnjHz6tBXwvEStBi9lxdj0H0QKf4L3HWDciMTVQQGzXJhXqLb12T2u3UJcULkAjw
ZJ7oSVtrRxARBaj1o9fatS7FkgmOph7Qc77xkFF8hsIPXHvsT91NLa1/azl7n6w5u9R5p0YB0Bsl
EezyQsxJcMrbK+dUwQMW2p/aMCHNJAnd/KFQypdEKhD4Iu53vn8Nys3q8q2YDqWmxq/PNNdBLbaw
oWky8H1i7G+el/4tUsCRQ/m52JW9n/X2CRYjvUMbcSyHKY96LT3wmtCVixydy20VwXrALeolX4Ee
eedl7cK0AlSKWGlgq5VrkDT2+HlxneqRrzEhUuk=

`pragma protect end_protected
////////////////////////////////////////////////////////////////////////////////////////////////////////////


`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-1", key_method="rsa"
`pragma protect key_block
PwaGx8hkz2M4CB8UuwTpFxmiyBx5yC416umgjwAUk6mjlgyZXh1xdekXKZQ6qT7GfocRo0wKZPMo
V/5wWMcSIndd7YUaRe/v/D5f/bPj7B/ODnCD7G/DR+1lG8TnkQIxo4cb51l9Juw/5DxwIc5s8HO/
hMnBTOATVrTpm22DKi8=

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Synopsys", key_keyname="SNPS-VCS-RSA-1", key_method="rsa"
`pragma protect key_block
0RKdt6q6xIe6m9rJntrRDt4JoICguPEulGfk4afxAboWXoOG73yoz+dWBNYZRtNDMONLdMH+pTN4
uSMx1QutXPjFImgcX5X2EdF3t/jxEexzadlZr6mZ/Hssnmt3+TtxXzCjt+SzBH2a7cLVkO0ZAwts
VHcfKuoC56QqXq6qlsA=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=704)
`pragma protect data_block
Z1vQNhvJIJidkfbbvMBlq2/aQEtaIJZoRHfq6RrXg9w9n9XYyYLmZPWzXZJCSQDf4PbBQyaEFFc0
hqiVYk11136JOAYhJBIMZpFDjhju1jpn7A8QgW3htj0fv0yxlOuurSmsHmRSdYReYhFKtyaCmhoy
yLSCPW10iyiVem2zImnZYn6607CiCjCvwt00xl8KrpZY6ekMqUYb64ATWoWBf6anWNyyJFagtunS
ni+LpFqVXxcYatTbABHp5xonzTrAP5OJsXSjIn9RU77LBzukixXP2zxIqPN2ZoFJcwWbV2Z+yhd6
BpqzyULA7q9uNmRWsfuA2IO0ndqzFcFGQK785dUYFy4hnLMTvh37BWOw4EqCBU391uOIEAG0sOCR
+UTFDDUit/iIhsslOW95dZXytSMSDKFkT7F999EhAOVMr0G3VabHm7SqqvcSS4xhUjNP5n/Pv/W3
xK3JwSBZRHWeiF1R6JbhgfT5jnkLfoGyaygABouKcw9RlPGFtq20y5x2BhYxhknfbJnNNUcyzmJP
YenO9shv6vufMh78XfwjSeX833dzTc+euXuw6j5vO/6ut8ZzC7y7RonofPu6BrVGYCuzVhNjlXQD
zcMMQGy31bfH9kp2gfgvvAhTiwbj8h1tjEYsgiVzPFu5Q/PLOmCIMyFWOjPLEG1Tps/UTwaTE/BV
TEP4awCibAWsroMCEBZqHqBmkgTudUtVL6lDdhLEhjF8RNBOlmm1dO4O4zkxrby0E9IlSn++aH94
qLuxRpZ6KxKqJWxgBfHVmf/Y+IGrbAHF4rz91vPKfG7cYOpdtsi3HgiMyTtDdQFLiOcxNq775ksV
tmKGU3IqEsLVKgGoXC1ezKN2aIVium7sohWwrYvi1JcD1K/9gPP/jJH3A4ZfXSn+pSv6/QvAZJ+s
uY+5nK5BUAG+HYnThczb099dapE=

`pragma protect end_protected
////////////////////////////////////////////////////////////////////////////////////////////////////////////


`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-1", key_method="rsa"
`pragma protect key_block
e4E12ROGT1v2s6+O68BD2nuEC4HU2RZlkkrq3in+C9uCnfGwbBPRrtQWH/uqk28mpQZ6f4PeUkAi
NASYRrV9IIhc2kVfLX5q0lJiWhBglKDS4KvGgD3MP/lJRE8BWDrBOnmq2fbd3U6TJopW5+LMHImx
7V6Q7yNYm2ONcHxaDl8=

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Synopsys", key_keyname="SNPS-VCS-RSA-1", key_method="rsa"
`pragma protect key_block
wgn20OjDEElsjSoDSv+LmIWsbaegh0B3iEvFzA+SC6DJFz5/pmV5BuOlII0v5rHMbhfP53nL5BOG
As87Rk0Jovk4b4PnuY7S/gA6zWHJHrSPMmCqZnW83AC6lS5sGY5PxcxxVdkYJnzsyF0WN7orvYwq
Y2B8OsRBFliqaDyUSz0=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=126576)
`pragma protect data_block
O4xBEDiNocrZemKiXomaeNFBre/TatEEoQgCX6fowt99gBWrYlmMzVaQluKisgTkdgYGMHfTmbss
WtUERDNSKHts1mV+TzHirg0nfuXLB/+9JrHHulREeFwJuDvZmlVvIFEpGrwGcDKAZuEmLTJa4Aq5
r92YYAlfVKMFS5tzyMMSuWyK325mHRwdSX0eOwL4HYk9/G0FwYmTzIERVaHSSXDQPnRmrQtDVE1z
Joa23CIGwOA7YPZeJ15wEPVyv/0ISSwsmqZ/xFWL39bwqk4pUqicPvOytKUV4R908hZBEOA+A13A
tL6zsrItUoLFyV9lCaPdsyJ9+6U20tPD1O6xLIzwI8Vs8ZeFQaKN86Dlx7qOWZiezUJXA9RFHyRj
UC9D2vsIXpTBu7yM5eYicZdDCNm0BMvp9eV8P02uw5N+oANRqioad5jaOmBbgrfq4rn7C0CVeOa0
gJOFMTjwTtTX01czdc5hmsQTGJAVSMXgWdPi8rmYxlZS6qbi1mNEqHeSyyRXG7LEQuviTE+XEmeZ
KqxOWS3XB/BHgEATShyKu37IFjOvRmClCPJqWujXA/Jl3tD4QhgAKYjWvQUR37eBiRGibzWv9JCT
Ql5c6mdn1XH3Ze6MAEzsi/ELsL9u8taLUPMO4CGJZY3ESNGCKvNGYrnYL41hPWs7UN9zA+RgDvwX
jeQIM1TQ97J9WZSsJ5fFMpznbTIX55Z+sv+TLdrybwKlNNaKu4LBROopZ/81ZMTVMKCOVvrOODfA
wryN6vzNWNsk1Bcia60ecL/Zlpi5qPhUbyPZoPByMilVHE/SwU3CIPKzq1NLhWgLXkYh5lU7NX9v
7zHd0an1pYmuGft9cQ6Fn4vsaJzGOAjzt6rfhEcxBZLv/CrgKfusR11ORLPBtrPu+Y62TrL8ExMI
QF0oRjSHvy9iQYVofvnK9aqPl1oB79c1JRXlMIP7eTSoWAWTmq897iyiQ575g5eyQ87rtPZW4POd
HR+gH3ZuQLZjx2WSi7oz6PLfmfxANbaHvriOnP2kU6RDMUlhc/7Ja8HlyaSWWgdpsQdXSEYzxJ76
3C5i/7SMJ1sOfo0c4lh2N/6pTRd19pAH6snm1ITm+dtzdjzh7JjVGDH/n+8vXoFwLrr9NAcRnupy
EIZBwBYnHqJir2Vn3pr7WzxRnavAzAhbvh0kQ1P0BQZZ5mZP0LxSZkumDhnF6FJwbUZDr6iNXiiI
QcLAktHfIzaTO0zSNhKix/qkTKheSmyktehu9dpTJfK5o7aeVGFon/BrYv+9mmtpmlOVcsQBE6hP
g6G5Gn2y8CuxCc4pWb/LfDHNp1oGuh/GONMPUprGkyQ0/0D/owKDhLZW3cPXflFmYHS33/5Tw3Dy
V8taO67Rk4MYvWNlB7DnlDRHSUBKMZ+p0cf3l0JnFYkEEQ2IjmHAF0a0DSN11dBbtXeCtKF/c1qi
h+hReVA1uk5nssB9/ZNfSd+CpVPr/7mDQDX1f+0Mmc1yi4A9Yc+dNtPgss1IGz8p6S5JahkhXgR2
QB7HeoNbGvSD4ya+cMusCONkzq/hjRpcbMs3H86TEy1IUg1VOT9bsgz8M/xEaxUg6At7LoYNC4Mu
CCltkk8FPKUF7CGO628ksr3KdzFJxBXLe3c0//h9iZMYYp1B+FE2GVBobavGrAueqxJFmr+j2P+D
Mvcl+xQxccdmg7DieZswjl5O6BfGoUfEB3AYQq3i5ByM8TPbWAmjDvstomBCnOgqY3g3Ra68FaxG
27zBOtQGXvj+cEcUzeD4bvLQhBZw87kSYvM7nZpcVglHT6OPCWAprv3dulPrUFOMwR7sUp0uLvST
FaVjin4qr/otGwX4mSD8rQ62BPqQvJBWgywBQgXhnBJP5YEQ4faM9HCQjQFqRd66GY+CP6aatKmm
zt3kxFx6ZE0bekrzwKJZSN4a53ycVEzz9cH1ZlpDYR8D53wKlJ90d4Dk3B1FmU7CZ1uKFFK3CB/n
qJIJU4ciFm7HGM961ZpSw/4J6uBzCp+PBN9DYnB5ecmmEDfvZfCebktH14abKXKRLfxfQLJRBC9U
GAGNkK1QOj+r5Y9DdytaGOgkAqxThClaoBc9TX4f4tE1MlKbExJhFcqZba0+M4sJs2O40Dveqsde
vm0rJPE/jks+nK/othQ+oM2aBo5uBQj+aqvu/Wjd2kdQLttN8BPf/1h63sV4BcyPNUkDCxIXTheP
KGolUHwe0rQaIXLhh29nt0+Bdp+kjsfx17TW4raLB3yGvY7VCHgO1/GxDqUpJ/mw91j7Q9HXjE9m
Ye0UeG82ZwRB3YIniCCzL93m7FnFIFwCpPZujtri2Av8zM9vHCiGywdrFU+cCz/iBIc2LQ5cnv35
kxJVHzALRnEL+vwL2sdy9U6urBtJHj8E57UYwn5yKKFRK/mjTH1ajJ7oF3Qs9HFSIbeT84rcfhRf
JIpxUgQKvrZMOauykGwXTjn8h5B8EhxvQdDuewpXlwVGxxrS7fDdYnNMthDwkQ4HyrXLJLefEz3z
QR+cqbSVTbUhhrNgUpKZkoDmVASS0/YQNob0v6HDc4aGb3D2HhzGt1EOGdREn0qVBShht8410Vm6
vE13q0yvh3kOBvBN5KSIC+CnLIJft0I2P3QH6W8Et9erV/DRBZQGdnaNUTgBhE6DXCjHpSkUPUQB
A/wUS73pgJSVeDNb7yv54LgkM9GPayljivgEZ8p7O7L2OazbYEA62p5Qf78g1qkzsCKcHhYgdxo9
C9hPswp2V9S1zD/XCXJ/wiKet8kqzAKeV2Eh6RWu8GeTH8VfOZ1+9ZBDMBTfTcqTGTV+rCT+7jZ5
0WrB45LHFeuXyst9PUAMmiR5wHnvLkVrucxslybFDh81txR5v2B9iD2Kr6ieKcya7R/TGBZzzoG4
SvWnPvQrgnG7KN1KJniat8uSL/FZcgJUbzkI8nWiCDBRgJ/utugDD4VBcv7a5H6hBjh7FTDlyCHh
+B0hxZ92BREZ/A9GJqHCNz5XopDdvHzzMmoYyyOeb6t1Cf0HrL8JIKMmDuqJCzWsuN8Xtniy3Rh0
9eTyMxJWa1bEHjp31Mh5yiOA1oXTi9nXMifgRfhRF1tqcm+e1cQORWaDoV67B3rCltciO2I2kllS
kBZAojHrIs9KqB8vlWZhdr6UvVDr59551W8q0PdsrNVgf/RjlSVYYM5aW4GI/o8cYJRswKZsZ7ou
UnzVuJN/2r1AdUZjK8Q1yjroEa/SIrqFY3RWAInq9FbqH1Eq4JUghhh4wDU0SRQbt1xGPiUkc2xS
94eAimtC13AkJT3WtkmHnHQdJ3pxF2wxuUxU0eMB7iF4H7QpQRv9cTNrAzppW2fYOtybrTO/sAG0
fc0x3gJxN8sgOSepopzsYT4YoOKIi+sGIEHpwHu3xFggZr+Gl26C9jvQNGGRbCjFuXg50iBJqR6Q
CcYbvZIYhOBV1RxSZrzM5NsIQDFntG4ajJpSRXQgeQt9JEUcgyFZeJgw+t5TNO6F2Jj2f2GqTsaw
nitNlqhwwYXYNm+N56pcCt24m+3A4R4S8iVSvA3ngUxH6wZU2BWTWzbqjm3FnCsxwjz53+/HUiyz
c5gS02uka2fBgmf3c+bcV2AZTSP545ojMm18pxYuq0Y1R/9zihuNyLZJi6MLlP/2mpK6pHF1nOBp
mjjJDFbEFsOJTVpwsBHG6I4jCQp+zmSzBT7iQM5POZ/7f6x8ytq4+2Pg9zuCiRJfETLBtj548XK2
x1by9HuqVJ2xQUUxJfblbA3Uv6VBpsWS4Vwgc6jpLryZnLY/rVFz7ghW9XXNfO/pvJYyeWjs3as8
ZtehFuPPlK5+dgfbqzLEV+Pq9aqDtnFvqVnmUsnwJB1M8RF5gVd18rxnE7ybdV1mUbrAnI6lYdOj
15Jn7z5D4vUYT98xdXSMgVwRrY8XrSDyZnBfYS436gc3Jf9bg1XsFIkhVwU1BQHITTHttv1r9Euw
ny+O0NMVvwLS5jDCOj2QB0wxJo7oEvvL8B5/WgrclElDyxWFrUXQI4ONJh4cFLKxvhKrjJOIb49Y
mVWQoblsgksbaAqr62HTe/jo6dBgqVegBZbFKfi7oWS8uNzQgf6A7H++wEWriTVhEBMTlLHaLLn/
Ts4pbu193twf5ChljA+S3tSCeCod+nANWEQV6zwX4GG8A/gMBymjLOjP0sivdptOJalzsWoNltRy
8jpdnOVYtfZPZSRKFpK9kc9t+dcJLYpnP7aNXbEbsiwCYzCzGpouM3BlGQA/1FaeLp3AYWmL2+Jr
RKxeEws5iEtzJZ1UzBzNNL4qCBG2sMkXvd4vccX/DMUhM3mnNBlzuzq+aqyntL/PhXosZ3EgaM6H
svMW8lXunqzO7/EJTfd3b+oCdO+1ZnFPJX7scVLAN58vd3nFUCkRPw7V4F7od9MvIQmKeqERkfxE
g3VFIhurBhN4sQNUYL5LQRf4z/81POgwzK2uufhTrMqK7NdCHOplEOUPHWm8pO5YtB1gDNaVCaig
DljGr4NVmLY9QdGCF4uU7Dcasuoa3HkIZrIq2e1bBfPJZWTIHruAlPjzhyYe9VtO/y3T/x1eSf9W
BIdgSyJxMOATLX+EASLBRSN8kmKxbSKfmH46xm/eA/giQTGTgaLdSqrrTFp9jB0t9xYmdiRyuU6S
x5f1Ie1kJzF7wJ34Mvb6+dBaIuYvjx//QGxoDbPOv2bGDzF6kRjXcOlYeQiAVTD7IBJ1dLs8X9Ow
UYt+fWgO24dqvooqQhjek8/WGA+/CBrIjF69Xlsx7wBrTrHz6bJQlLiDvi62OWyEqaNPiHivHEPv
8LihutVspHOCpqQ7nL65TF0VH22/xVgGLrGpOhP9221WOp6c8q7w0vCX8+a8iQ5knWMQj0rcF5PE
uzf3BgXaJGQ9FiQWtjEZi7WUkSvSvaVwI1s8UBu2TVH29KTMeEBNWpIHsrhnySLkXVXLrOfvpBLq
tpJuXrqy7gzdoyOXDc3zHljOKJTmKbR7kezwtNsPBpTjyN0Q3e6R+FgXzo7BfAStQI2uYpjxEVlX
usLKgN1NRZcCEfktGLVygplSJ2ySB3itFyiMVY+iY0eOZvk4eHlrlzGj5tzopBFZTGoSh1c7m/MQ
O8uevfxvM3DtdK5Ulhc13r2t0ZcnaNRCEyxjx+MdItX3e4x8imTMfQWT0rICm4p2Zwp0JSSEvO/B
QwNzD5arV+ttlhTUMM3UsV2CIhyfpQglc3EYDVdEnn/mkj6neZ0zt18fIz9EMopQsEmqC7eCZRlx
NSdLJf6bjw48zzJ4mUJmf79Qg5WrPUj2x+k+OU4FONPO6rA0icKptOTTw1lLXarm0OBf2g8uVVeV
mcEZRAIARY7bEqHvmtW6thimcV70fzooysXeeCIXZcSXD3r4J7p19uqPAkhFDBlIDI60vVr7sRfV
Zhledsh24Jr9wkHWacaSODMqeIBrOaGvwkLeHdY/YGLKzy1sSsok2/tvsRj8ejnuVbYmazWbKjYJ
Kn0cNMOlz6DxmJs/zAdlCIHWZPFAgggIE4iPXK51Qv6QOoVH+VEBskZWxKBB4iMDwHeiskU0QRa1
GcQ03X1ckaSzfibRMg1gaMvpLCUSp4gclsGitJCIheTGL96HljfJfwevyFUOcT37C8xg7P7lp5ly
/0hk0w6GVctH0RgqZgMpMansb5FjmOh9fsHUTBBogz7PL1iI3wspe3CId6ABVAgZkfikCH6YfarJ
2dG3gDAhu1WwkVjG7fjsrai29KGMjbv5JMClyu1zcdkaweK3YJbJ1gOlXf43BrkGnu9f1ZALuxkL
4JVE71ZgKxlRepx+D+AoIxIwllFP3dcrYG3EZoUgbe1J4DorFrP9FXGWsN4A73SNP7Ima4khCyug
zKSF9LRJ3Q7ON4C8Oh7jHE3QIXX2ked6t07D3P7au0H1ocOI5JxbwQLlHca0wtd+NhNOcQU2dIZD
ITQjydWo21FvFHVAlxrxHR000AmDhtHeXmzjeR7rSs1uqeDy0s78qr1hIwaM4CRU/bMup19DnMWS
muhbRNbAWQUFmRcHSSQCNnTfGme+lnh9T8fMhxu1e+cc7TG+1Ltp3ZNXYBq+ZKpSnItU/tgK8+Yu
jYcWftn/Oue5Wtp/J8CU9sxbLyyoSuD3xlfmDDZ4aV/JB1E9iT3yMfS4G9+1czeiqGidjXh/HfXv
i7AIUjeYhMPLYj069121km6uPtEJxtNT3DWdh/8N+VLATZ+njV58I8fpdgOivd/9pGTJuq0bYpCS
TGgsDQ2tpHMDg3kbh726d5uaPiGNeT4Um+TWiFY4N5aasCkcbNXFPpBMcohHm7gLvaequDKORMSY
QG5pWzKQXS8+Kkzjzb2A1nNin1V48BKukqC9myercrJIA1MZpN1udLbychxNp+jsakLn2xX3j1UC
uJePkLSaWItP9rNEjWrwwbml7jEDY2GTwkJnDoYCXOFzDqOXJAsuKnbrSCN65aQG2HMd8RlFFpz7
3RFP/JEbLhboxra7fkC1KbjEd3kCoGqbxciYtYHuKZ/mcYjJoTxMviNEGRmwJUNKLgxvSdp7N2ku
wfWN38289p1wh928BXLU6koYL6RWEa5a6IwjTEG+IQSSt0fMZhX7A+QI+YUXnXygVSvcTZH93jMg
4ZH5k/Qa4Ikqw1wa0vUmNcloDe7uVZ7O+OG2Iyt7ieAsB8YE8dHr7W4L+1vnYYwDCY/vdBQ/eCXP
l0WkXJQoj0twpWoV4clX/cJK1k4XElllpJ9lxnP/P7SWGxpGWbaAZUlHssj5ubQk7//ehffXoyoa
lQQlxxVavfYgLDqsXN1GYmjJq2b+q1zAEmBXXRB7D2YUrUMaci+0u4ig/y+xhgNb4TtJlMKDYhpJ
wM+8SWzdrQvCki3IJk5DVOLSDEmYxRtVcr3nLjEm9NxCZpThC6sExDayiyTk+sB781liAmiJI010
mxqSXfW8YuNDSmJvsIFRWXzEU+cEIaZz+Wr4ti2xy/L8FznhLHr6g24mVYfrDXXXPRTWSxLtiRE4
GrRESMqw5dDDs0RgUKTZi5l7+EL9IQCuXGYs7p1J4ABF/SVQDqwoGVTExAxdjqe60A0Av3txQagk
nVPo2H6uuWDgCS65qEIdddhMYwgWoAIIKbds79OqTNgKqxvBBsWuBRecg7ljoUp5zQQRhMKyuxNZ
EosorMIBdMEfgGIgJN2nhpMU+guQnJVY5dPlfoK/sLlFAV2dFcCav6RLzQZEjl3nWJ4SWStfFyj7
ZKraBOQM2cRaHhxsaLMLBlxrIi/9VXbTQhPGWK0w6n/Td8109VgTIoBhLY4c6gM3yV1bRC8ylOua
mAs/Uw0KDHY2UNWQbjY6LYQ4naENJfeKWg70hAM66tM9wlFpdDheASxooaf2myZLNwCn78c956MI
KijrwIBbtlLB+FxqwGwZ/5pzJzTBh6RX06qyThc8aCOZKDevClrK0xxwTWlAlWmlNycIauzEMN1G
SJY7Q/bofg5rrl/k5X2nX6bFQUDwRLMKjLbBUZkcKDZ9P6UfMPDjXspbPg+tn7/BViL2L9RdX8p9
WX7NqAHBxDK/cCPNF0RoUNeNhracwIXwI6Cc/okz2Mbt+1ATJwpHWzKxEQxH/X9UuvPXe7OqhxE2
r+falKj1tK6JmtxPrU9gnYK/4CQLZcmEhmZVVUt4dhF2v81EF46i026TbVhUeUH2ot815SYSh6gS
Wgyih9mh1Ech8j8Uoxa+9JudsJa255BxKQ3FKNp9nMh7yFk5RIq61pg0lUgODy9drbTh8OLepXkL
wBr+Qxew85BMeXh+VX/+Ld1mgkQPBRvK/kRrVEdpf2Gu+4im/wDsIKuv3GNIGxHQzheNUrvorpUs
LcVvCXfQHU0Tyj4dPZIzv6FxMvyYetJV/+EZVGgI3bw3GcJlVGtlc8tBmgVF7rWWGeWfAzSMV67o
gJUqV7QVxtiwzVrLCmdtt68fgbb5VBf6wPRpkBlYAr2sBB9Gf1d5z8OgH26iOxfea0hg3qPmrdV+
Dzm6Gz8DbYSo/0+RSpQSp3djo6ZdHNwnGAta0TZCyw3TivZ8gmQJAl/sLKafKP6QrWNGcatdWlGu
h1/Q7DLO7nHUhs9+GQpLZH9cILl5f2W1MujUAVvHxzrt7eSv/LNMnwRZcY2h9NxxW0i7KQbHQlZT
wJMOq5L4JIHf3dkZbctc7vctORLeoipeCFfHfvUUI4wuy8vc857kN4likPF9x9gPiJtKnBE2Cg22
OV6AKHEuZTM1/mQ8+kbPnwOkwLv+RRStqQUpxxgiXRCFgQslf00Blv+6OnpyQnNujW7QK7Guz5x5
hq9PRnYSxP3WTxmy0+2KC54qMH9RQiZT5wsmJiDPawbTrCDdcNqZOkZNHHRfAVpdeC1OP/Oxlgi7
NnKmCno+CD6hEwf98u6CtHg2j1zoZ1ABBTBJEOYffdU58trEpkCPDbo/In8KCuqLNOdmVUj3eWlD
RbSGyUuAQMykxdsSwVKqFxlhwNY6bSvy21tQ2Gd+dsUKR66Q+qJeHNPELyLS8tX442YcxqZNXeXE
LmSS1+ngfsLALtiFcLvEU/0YqbVz70WpPVDhFn2ya5hySb93A7TgVGFNzJwfDhJiTq3QJwvu/XdH
870uEOl7Jt/z+ZCpUiQ/FSJopHM6kKJ8VLMUXdrKro+U6xqN/9JkjbFKmkMn4P6buVcvS/Qb+yU7
JuSZwQoBQDH45fs9C6xDMyvYiuV8MF9Pxdx6jTP0J0q9izuBdQVBUdPEs5/28j1Wut+iGGcJvJsa
Dfyk8m5IgRiF9xt+9nDfbaTZBilrZB1GOEmI0iifa+n1HKGv7I/rrPm5D98jlhjKrFztijCLJlbV
qtTyLpjnFD8uTSOX0/MgPxYP6bMZ+p1+IAaJJ1/F/Nk2ACj7UZEZvIFzLrwRNA/DnyE5K6uWKjfD
mysFUFUf30DAtjuFbHwkVprsNRIEbmebkN8IhV9U9AIOE74ji1HmHMrevsYk+G8VyENCnkxWM2Z6
pbg/qeTNpnHy+LpCKCPGiSYmXKCOryIUu/14b+drR3x+wz35ppIDFL5B6GgWpGixeQU2CfSAhryI
UdZfVJ9L7julIb02k+FKHgdpwjbO/3X7hMG7ulC8BrVNEc6ap9DRDeqs5J+loYhz173lJJ1eGP3O
n44zT4ZxmsBo4J23tzlvkYU6yIhSUP05EWu4nMz5Wer4SJ7jB9qDKJvZFlVWHTKdYd9e2uSbk5H2
qhT0vpMb2qWOlV8tVpI7Ge3d4bSRh0ASHlHzM/vS9WSa6nD/HXOWJ8XZ6awVlT6u/KFBrytan56u
ETzVBDSuMVpOH6A7BGkX+SIVA0BTO4e3Sdr7lwGZklZ1glYcYOefILk88HAFdJ2Wdl4QcDCDa/MM
AGyCBcIy7TyabHbfcTNIJdb34OWOGvXYofYCL6ur58d9VA+sPjAIjC2fQaeTaAH1ivrS5Hnr5Prf
gR1acpHm1RK/1LB0pXpM9LytK1YiVQAr3f62QJB/6IuyGqa7swHuPDg9Fg/fxi5M+G4jKMA6hRnG
9ln4kWQBFt/CO2wr9GcULOlQvFkn6H48JZuqBkT05tnxYARPw3K8FUNZG2SJkR0shn33T6B1xYVO
gD1GIR0Ox3r64VLLGeKuRZlM34S68nQpTPdh2z++DjN1m5dvCph3Y08U9JYxl8wKw25C6ZPcry3B
4Y7sVsViwswHYMjgBfWQgHDDlNIZNyiehM394iG3R7RqP8rEUu2oYU3WEq21SjAKe9SLBr2wGwPU
2LoJC96bk16XmfySAek6meovvuDA7uYUS52RjvRWy0nhjcn6ETVXcVcjq4H5oeayTQm1KyPEfLHG
Ro0UU0Aiy7WfeLaDqdWd8FlXJ1xBdnctFOelBVCbrQeoJANbuTNpdfrnhZU6OIddE2wN04YlJ/tR
+DUf4XiTivR8arg1yLcgFAp+nOVgqVMH4GZ7II+V5g6wLSfgf377tRGDZNpqF0VL5ycNQQee27GL
4ZXY/NgT0Rkumd5wDuyaj5iICe64qWDtvWf6E6WgubQ335zq9S6PrSBqMWrpTq3ExI0VFNLBib6R
LFLTf8IXV6VdGksNX80Pr16ofegsWxAMNZ2iO7ad94TRWSNIV1PNlHhu0tYb2Bc88KEDOq0+wsIv
YjSnyx+SZOifTl1OvpNjQGgV8qapC12HbkviVVjv+t+p30od0ZIE2Zq55eyp5Z6g+0sPprsCCioO
aDystPz+2KmKGnwMxQmpVRA1OliyRP2MMtmvETTS8ItotPJizcPte5Es3mag8N8cpWpBkzV6R0pu
/4blKwC4TXbGUxKbB0s58feOofpCTL+Ybg6iqd6THk1gW6sA8t3sk0xdFyitfCgVjLcCz8wHN5Ov
n+cZM1QyejflF5oi/oqKHH4fdgcdG3/V8Pi68LQa741UWPM0ZHWCSYwbXHFT6ptRRN5QwfL0+nJA
TcWPhqyh5z5gnMT5e4NuLu/0ifx9WgtnPg9gF8cpDk6AY7hUWZEerBZrB9GWYSzbIwND9q61uwkM
UCRpnJAqC0JWvHPPchvDRp6kD1UpWbs1nEY7lCLyCFovyU7qrw8J/W23YPq1lVj+kIxdnaRBlOYl
1Jkv/HvJTEO3n9C+YKYNFgq+XfbPr+NusK+lFMtLEBEmaSx0fVXrz0BgGcZR0M+zTgbXXXl1cVQ0
1J9667AtCebOB1fzcrIOBhxW9gA0/qE5kIa4G3+rURYLZIQ+4nnelf1bYfkBAhtshi7HD8Mmf0SE
r48WUoCKTdJ6Y27yXUZrdY1IkwxpYf2L5sJSN5yrqhkp02GArd3m+1jPm3Ib3nfyQ2G+uNsnJhv3
H+wFIlmjMFQebwwBg20Qk7aL+nuLj81W6FaUrrTOgUqk/am8bBvtw1KL+/UWma9UP1spoC7Fhgnz
oVMQBZqq18eGA4kQJ1cqTaSFDAhNNon7G/H2LJIs+FAsjZNTrcuDtOHULAa7KXAKFwO0JTsPvF+N
OqW+ReeGH4lBeH5NT2LV7M8PyMPzt2I6x2mYw3ZATe0VLoup5pWYZgSp098BMwM+oa5MDAElJfY0
RvA9J2F6b1HxA1K3ImQBihVQr6LvXvi1Y9p/SXltVZZd1TNoMKaO9xFIVT1eGf6CbUs6LD9Qjtqf
Vw9ovGQ+UOu01KoA0pqfR3J4D3obXMI8jQLjsB6/L0cMSSO/ArwlKA10/4dE5l27yuUnpJoiHF5Z
8sefIkURrShty6s+5mbIHuC3ht85seVjBa+kG067+RLce6TZUnE/AeqYROvS4vhy58MJU0j3ndUY
wRpN6T2yIVTDwfW0Xf156/pqI203jf1Gvy+RGcx+uCirX7cn7pXqHHeaFvXiRVvdakQeODelQmJt
VZ+Eh6IPRnbFbILB4IjHV5SQ4NYMJ0K2M3L1F6qFtNZ1Al0AFqd+lR2w/N3Oft4+RjoZh5JbZcnR
Cw0pjbvVnpQa7TzHCsI7l3cPNAYwdZbWf5x9hYos8E4nRr8TmgzDBGqPopgv7GORPFwjvTdxRio9
akTBzEYcqG6lL5cKqdKBRwVxmFFspqDfFxljMtEtWIdMBDu60E23Pq0ZxjVR4G908IU0m0TCNOQx
SsDtinxfCZorda3/ERMv1v6YA8Fd7L6rSD94xNvR61uNby0M89hZMH3cX9kbK17/O2p5UL0nBFcU
qYPMdf+z84mYqWgIKck3MYuIxuuwSBhfX8v6uJTRVfwcjjWGjUxSJa0eUQZ54YPlCASfCeaNrp5G
MQ5CaBlXadp6RIY+c1+ChYytfmw/lku2nVQq5p/PjNHUQyIOulWxbG6kmLoFI6i/niuNk5zSdKnh
ILwW+5Djg1rBKLObUGvN8FkVksQh4vvepSOhfRUqgkRYxWLWOxljKvLa2537Zh7u0cwU2A9DJ39l
s7kriXoVmFvGuewBAAKUk4uNuhQJct+HTxIF7LP9BdUEkoRxB4ClVILtDVQWoik8XE4SO3Eq3hn+
PXpNn+xoNwaYkSTpZR6uz+pt+RfFuPo25Gsy8emHtvEg1gFwE0IE4b1TbWxRaIBWbNkVFZWLAaaE
mw5G3vw+UjpB3c7SlUojFY/LrZ4n6GZJZ9/s+oT6AKJnyVWGv1ukIlKoubKfKAx5abKHSa0SBrPg
mdC3n6CNFzsOTRaw2KppoE/j0D9O449N8I1qvzgnSg6gQVMzYsGmCQaXro2y2CCUkZmhbcd6i1+6
JHGPmnK7lZ0mKZNGiR1G9CEn8Xf3ZetN2P1w1rdJvfSKWFMaWFdUqUCID425w/3Z5Thudvkf5MRW
39P5UulvgZgP0dQDkROVrQhodQI5QOgPfPKbxmam/j/65tfWY8h26gTnS5UiT3HezHjSuixMbv+B
lrNMCjcTfwIB4LZu+YaJLuE933SZZn818B/Gs7HZdvPRzVWtsAvEondVK6fXP7cJAlS8nYpJddOs
nC5Cwz76ExONLHM9x9PuJx932aYFv0TpWk6BJWt35ZvXIfMJBHboD9PRAWInLU4jmC5GV/ABvgE2
17aVcBtkbyFWg2axG4DFJwE+++ZM2qsmuSTrFMLUWvjXVyAcqmSbpvTbAlM/SDw2djS7DQvnRbRS
q9j/LkpqSytr7ZFxgQdVeQXBJ3YF7clXDaSmygxYdfJDDAq5NHWkkdk0BhfErcnzgr8KRvuJtXqX
VNIhlfrTKde1gL59RlifC2+fBvZINFwB91lFFpF8GIwJrkoJ0BIfyOXT33KHBTnIaFr/YeoJtLzA
x0ZdyCo6CRCdxDxX8WSHB8hbzyJ9of330LZ7axccTmnMFU75pa4wZhKhtGmecogMpYAQOMqW2DSA
No0WL2+Dhs8SOHo0uxVinxZ9oUOqtIUW2Rax1YNA6asoM28ItzAXrv8gjhCvDBZYQmgXdV8qKoT0
wCcdqPDr1osxpV81UF31bU/VZEpRhTRVl9XRMpX+u1tgahL5yxtJABLzlnnABN2rVoiNVX/7kWnE
CzKMjJ8k79+acX+SAR2/11AafuDFZzvSHxySytDhodcJdBA3doMBlHv9GrJyOhvKznlJ2FsKDBuh
nq2kn7O2cDrhCaUZAa0fJKeiZpxAal5edNslT7cbGp3dd4N9A5G9xboqHCdvVnWFZhxxKhsUshoN
oI0HIpdYkPhfqnhuUBMFsugtHcPTql5zRnP5Yk9nKRi07Ae8NHyi7qiuIVQR4bfQiXKrmNbN1IAr
FtUGnRDN02/7llLlYRIWC5VbLktqf6W1X+6aNvig+AIXN/Y2grLAGRbNC77B0Lm0Z97MtgBxShs/
wEU5Rro262XatpJbofaQ3ctQO3vzviFYeoHk+4tfgi2cxRPDJN9X3kLozOc93W7d4fcoJf6qVq1W
hnv10EznEFK17522V2u9/zUzUrGOg87/pDx5zQoo6FK0Lg07CREcb9CPlDFiw5gzUqP00jElJOpA
V8SKkor7mVTeMJFK1gmBPrv3DTwbqaNiXARoTl75cJntnK8EfwcN4ldFHqh/hSgVmDPC3rOCoAnY
UESewiSV1NvBeFMFxuTv8wayLux0RhR/eUEC+FXkSaYoMhy8Z1uu4IRutsbT7ZunEM+8Rc3B6UcC
Rk7y7yFxkNTdVNdjpVqq3bAT9/ay+OZ2nMd55C9saxKxLpd5SBZgLFnjT7nE/g1+7dWuVdON9JNY
HInxLpoDW/DiCwBtAPXQzlzhnPp7oQh1vDEY3xQgMugApP7xGJv/SrT/u1N2xliiIMFf9IgYnXWR
mDyVmBHynjKY/0VVD4Rgrxcrzm4Ka/1GOH7F9B6J8OVXfllBNfC1PFHGYxlw2hL1qRk8wOKE+NFH
4GHFugyVnMV6sYWhhbAT0A3AUBuZ/6EgnjY9r8S/yrn0aoWQRip39hx2x2ZE2Cm2CuRhwMPWAFsE
u8Ntzddr2i9NLKzMoHnBpd6vr7KdSTt1dK4WGiHOrNcoabyTac1czFH7LUxpafkVN6s3suzgOT87
LUbh1nKtMBuLOrpi7GR1K9kYvWGaKmfH2lw2RSdRGiNOdTSythdgafcUQYQnnG1rv82oMkc7UY3r
hqt9J8Iv3UGTGWU9Hu+39M7127iMY+HpcHvOt4qm+pzTuZvV3CdEZYV9eX3lmq8Rq1y36Z0uL1DI
VbloCH7EHRyIBMTsGwRGJu7DVZcAzC1CcFxxRpS7oCcBXlND4BUTKEMP9uBkLex0AxWnHgaDSjsz
pvkDRwuZJWlCHFZBbgPcAGpvBlYufavbQHLFxshA1K+esXKGelPUWR4wkXyXzd2Km8+f8/rRjW54
W6Mp+0w25R7Sz3XAsxxswD0jQOcaK+KTHc0VDatgU54aOxffeEPQcKmlst46YW4lo1mWAUXZf0Am
4hs5F2D747a6MfGngxCTZgxfd451blrVUlFZ2oQBLO0ebfmp63nHK/62qEPntNyaLzfBwh/TNt5w
dfNWp26tKZzFg1g7kJYnuWva6Gr0tRLazOgY65eSz3VTo/5vcA0JSyyMo3CPNxV5xJjiYl5NdV4n
8zz5HJie2FphTGLBusqJ9jo8NdfgYyun1txzSNzLBOKHcd3k49srdOFdm+Qea5kiqEpXKlUsMWBm
OQdRx7q4OgT8FfP6kZXX+o/Bfct2qEUSQPcteyYjFRW/vXFfG8xxJcd8RPpx7hipChAg3gyDlHT7
enN8MXqfuQu4ujWi8k34kIHRZBDL2gYBUDHFbmZaQiAE/PMFFxMDgNfHafDq3evJKSzlha2sm9Kv
8sSVANudNIEseDU8ks4pofO6nVc0yJ8EDMXoLmdEBuVVNNhue/kGuE/lw2sYeoJupc0L1cNInWQR
YOli6tMD25mzdEOJIJ7aS8Lk3E6PkmiuSpCEO5UpPX/6Ddj6WZ4LKgZkzcXuHwC6w61efOzuFf1V
3aTA+WJ91wNo9V0I3X3u0SmD2AyjJ+M62P692CAKayKNJTaiTUuT3i1nTHRaiRK1zNiq/k+zW6it
X3N3J0zo5O+xvN9+m4DPWoiT64IOrymldUa/yNEvFnVbTyDBBNrpGX2CTy8/LOT2/NVTq5yr5KwE
aY1J06vfz5vij6ptqFcKEqKedSjgZJnxrRt2H7J/YgJQTABoNkLf5+LHGhV6XdCqK3XhHMYo0VNt
GFb2kM838s+Ey2dVDSyTEGtvZhGeH+DqwywMlbtaLvtdjDW/CQ0SWCt8+ErzvkA2afnwWKXZwL51
FKdcxIC/B0kXBb79lqWofi3Veu+XJOpzHoYjBjA5D3jUV/YunRD4x010YMHv+7dYSojoLkfb/rLD
gVoS3wUt5OHCfan7lPe/STb+/vvVw9Idb77W6peVVsxnoD9B7y/h3pO3yz224bki7IovQ5szkjw9
rEIcerl/6Cfi5E2JzvIsN3bwOrOhoHADQrTAWYFgrxzvKFvpB4oO3lQILuWOjbgaD3+Q+QnHxnPA
CA6v3FbcBxGKi3IL/MEsRcuuWYJrVkZ6srAToXb11koya4nrm7SEPQUmRI1uLmGprnzeFsVaSBPT
bOvRBu41qrfbpvhqy1FsJM+amORVIripUB03YMu2b8ANcb6K4VmY5GZHiV6omm7ootcK6/Gi+QPP
hJ18u8f1BRXQ5dKWTP5ZRVB6Afqxg3B5M3VSjpD74fGtVyinpOjqFrgrb7j0MiKPyS2oJJt3VscO
GEVAzHh/rZ+MIGH564uWAFC87asCvUs4CkYl45VJ1JooV1rsNTRAKnRZc8FNquem0KJOYG/YUhKM
ZTrVwZhB+YPz/jUJ6/Ey2CCI9Cf2LgZ+srOJ0CQtGpDL0ymPmhIJM7COWk0imDZGGogT2KwqmQQi
+HMsqyt81uofWulhV505/y9zHr8t2K8kbzNaEeupWbU0GUqG9hlDtQAkyC+PjOTvet/Iv5nyx/l8
gaWr7eOXN3xUYFkgqtqq9tJBJ77YCeoTU5PmNpUHyBvvgXl2hANQw3n/mP01LXbQbrNVXXzEFjvm
x8JIvxjtthO/S2gEua2D1Ef7qJ9a5ZhiB5kG7PvQmz8T2P71GmCr0YlXYts2kno7ZdAMMIaOZsyc
5QbkqmCGQM4JpHqUZZmRJk6LQhvOHnO//p3p11A0KbCu+3tFV8MjRBtIlip9IU008xne+tSZBd7N
O3HFFlq5WVVZGMm+EysEWqshTvEVw5WbNUD5V0zgdqQ1PBr/B0m+KfSp5RirjInpm8O8lUVYXdV4
EmE5sCDCW3O6Jaloedi/9EGY4PmokekI2TkttX7V8eywSTvLtE8gcSaVaLTzDw9wU3bwh3U2ICXv
QZFMS6z3mQ2Qf4mQ7Uufik4I+WrN6iTki2UNgliWhZh0Cl7FMCrPKQl646Vgir42c4ITrP85c0FB
sQRwa5dIIWfHwr17sFzg/JVj8iOOzZAjvmFtDVW1cx8TDdbin6oFPrO3yXH1w3STgXSgsUbEZxC0
Qkfa2jSaJremGCTSsjqBktYedImxJ8EJcsSj8uaLW72CLhRP2uD/dQH624T+bnsokIp7cbIBqL7C
iNvxu06xs5pTmikAFzLBtatc/w6lnUSvEyHktuMiG/cU18XNeUPPmMoL196IObwXy3nOq+xBJ6GW
C3ZeU1VgL71W1NdzzFq9WZUJix78sutuTeecqOlW1r/IA07Lg+Iqs6ZbLCVCCJB6FHP6YP1PZK0E
swnnCYRyzbu+EyFbbYzjLk6U5Pb7MFOR1PewYaLwBtNF0gLgmQpggMGReXBCP7+ilRyxt5UatZ1B
fa0gJtkNd+lD4Y4m2rC1tNha/sqcDHP7SW57G/o0XljgmCx1lpM/iuVmn/AdeFs+8XJ3QCzQzZPe
2lITGyWArwfREqNwQxvop7fCIVla5XNCleJSo7yhpyt27Gp9ffNGlSWzOSWl37Wjob2wOcyKfN8D
T0vursYmKrpS3RIyv7Qfp3L2zZU0WKv+t1rC1Ua4+C5B7jk6XARXPuEX6OYIe+v90txqpx6bBdBD
m+eHW87dlt3dDak9e2PFJ78mu2QQ5p8yywg4M40wuwp6O+MfBGjKujpAJdKjtdi+yWLA1ToxOZ9H
xMQCFoUPO3gJi27kMqWPLjII64wd7JCnvMwJaD8mQgpDTYbViJ7xL6L30DEwgOTBU6VvYFPGgkfM
Ge2pAyYG6oZEAY4E3YuLTaoz8qkPGvg5pjPvdq29HX+/cQe+Huu84I7vi43nLDPDuMV3ZfoNun1I
aT9nT9lgsA9ZbAA7ouZJ2Zbt9lzIFCSbdDqYao5RINKDifMf72sSuh4LW4ksHYPqEJp+W5TjC2/Y
K1nwh9kgQz71NMCRgIv2idkS/df+BqU7TgCXRXEDocFWSXSsvLBLAfHlTr7iZ6wg9LC+VtOMX8et
fGwdSPOOnxmEDgYLpbGvhU6iedYLZS7jQE864asF0oq+qO0WnpRrkl0zNFNn8eJGbzSrj7zI9/Dg
Ucb/JDwmvzHzjozVlJvatGjrCCTdOSNTGJjDpNt3LW0Tt9luCScgNRXPqNzNBNq7LZlURsF8gXg9
06wauSVbcLG2CnbzHpbwEQ1yY3CqR4GM1ZafGsk7it+U6yu7JY9YAMh9zlGCyzhCIe39/Wj05aiU
55a+gszEMBiIAAC/8zlcN6m9TfXnX8QfsHXvTCyzleaJWw60bMTHWWnjH/iYRHFOEM8o0jUYX756
zG2OWkj5nCmopSYZIPUopFm+h3I1AXJzxaadf8NA2dwmKM1aeZS5rsaBC4JOnEMshOdzTRRmbVze
Dw6qQEMQD+E1tWzereKwyfT0IIXtfNEqt40y7XBHHIA3oP0FvA2k9Hsfq01GQc1oXG8+QlM/tldO
2eECOh7xF43kS147FYBy/ULDUcU2NqPOzhBYJWO3ubB4lFfWGvPvrEFUfhvXcXnmg4OOmVoEBugq
4sW7ceh9DanOKgowQQpn/YOEUbXDZ5kZqM/Ke+aOpTtBSWRQwLZpkND0yWWpVzY4p/ZvD313sYKl
z4FWtOInwivOMP8OJtveXjcevRZxFJvG04rCUb5d0+Y9VofmNeNy4MIPuL3/nJVTSbryfj3jI0+u
joXUf54lBABG0Tw70EFrdzrLtp/jJVG9C9yYWHowgQ+7SNwAJSNkid7hr4J6CP0UGcXIDkAA4Lf6
1TPmvJaEORO58gdQyD1fxCx+kSp3Sl8aV8SreuqeKnlqeyuP35nhwGN8Ib8ZzoVgQLDcsSG6HXh4
vhuEJ4ZOPhHFG/xjZ1qk6p11VsvDINqs22YA1PUGJZNtf1VaFhGg6doo+RvLPs+ruh0yEd0fRdVe
sABmTV6aYZnQWNl052Mcz2r0KJ1UqWDr/Uj/bqCnqptCvCTsW5RFyXFCLz8TP8hPE/cB8fTlIF8D
aoSf6WiLG+ZLsaBG76x7iWRyJbGc6VRUzEh3/CWbFR2+LU04cfxnGro+9lAVYEqp6rMEO8E/5dmy
ou1UGWgc75QI0dJr1C/qP83BZWXHTx9xBSmNRFZ+yXU5AIXAxd+hitRXr54L/tso8qCoW/FgTs2z
JWQT+/tzh8YnLQnJuxLyHMXVogI66WFwPl/rehP/12GvUCJVXia/4xRa1sq96y6dl7jlfJeEbzaH
1PTbAI4ddlv8BAlWVdCL/9LYtLDrW18MLwzu5S1J6O+OUiKS/77L6zjtYUiI1eaqwso0fdkKMhdA
aLQ9deeGVTOiwPvam782toijNMP1Rzc0x7QxTmEM7E+lALaYvsWSi9jDgJh6Yk9w1QQ8bzZNNtKo
lKTBf900j6fxQXMTN8P9A7KNZp5GtYRQSa+Af0zf33Ug6LFdaZ5SH4WxSJh6dM4mrFcoFzrP0DRJ
CeQ5ucVsp23z4+kb9eIc3dp17x+jgfAnPMonl8I/bc6Kf3vs2smiYn6GSJ2J02Tjs5VuSbHbE1v6
0XN31Pf6SBJZcF8s1+d8HCCZxpVJpYN0UCp+xemdT+vG9oON5Prw+4fg0RrH4xFImo4knZDFkkvD
BK9Pp00cVPn61jfXPv7dr0IcHdV57MGcZzJCS0E581X+8F/nvCS6tssSLQ30OCS24dBY+KUH0wOY
TmPNpExNsfJ2b29k6IjaZGSwB60Gzhk3/AvWV4jLB/5Pg9gyHYH5zdXuh24R72iwTx1S5y3HVdmb
u+ScEJn2xMkIBwV00b1V2bOmU98pIXpJvGYYnGUhVCXbPiFiGWKqOy3K5LDb8ymygz5z+/z1vp8J
dcBpwtiQPIkSZD5vSuV4x74g+mVBder3C/YSXxroHBMeltBdKEpLz5Q03dy7S2mtIwI1e1enCYAa
5PjnVw6OFCA6vWmqUegqu1k8TrRbWdZ2c78cJWud76DYoFVp3mLA3tEfb7GKi2jRgdi5hUV9+A7U
G/BhDUMtOaU9py5l6mS0YbttJuALh5XIdKH6L6hSkTW+q61pi/4ofCJVU5aVr57SJaGdbiQoYcD9
29y/mqEbxQqCaXZxw9qww9hlg/hOgYANOxHQeeZo/5BRAqfN8VWvZKJAu1XSWKb8XwvIskle76sn
sllZAjAP8/P6tLk+Kx7M25yVlnlNnSYx7ROzl7bJdXo9IGKifWlzOFJKW0Z7W71JjzVWiYKFjgEE
TOlXLu1G5gubxaG1oeCGWH80i0RrHXiUP0Xd97hNth898inYGnGeFssDVquixkqpToHjg/l37L/W
Bx7MIECiZK1KY/9Lbr6Xw+NNM1jRv/0MvjA9VrrScYc5Lmu9B7kEL7lYKGIKuZFK18hQSd1REssJ
miLmzk0XYyNKKNFaZ3IrySiAPKJVmdwcRe3ux0TMXSL1FVOwdDctgSOs4F/NGKuKx+p5U2MIG9dM
3PPykjvpvhQ89rB5nFMqpR8Ly438ZEBeAFNknXg3El6Lkaaqdx5tdDVcV1M/9eIcBG1iqXfBMDgD
6gcQjypBXqPJP5FNjaIIYApGwLiWTCjdiDmk4jE9rKn7mrTP32nZJm2ekMwW50JvvN+//ojumv8h
OubTuzZ2yr1ufE5KTzYq/245ikE4v53aSNorXzZmWHS0MxcceBiR4VSPGFs/dqv+YrQCg17XqoBK
Bu/LT5Tisj1iq2ji0N3kfK/pOCPq432Reyp6EbETuUoGVeawzev0QhTx1qAc06ms1X1YXED966Gm
7YRfiaSMZXS3RMIQJg4JPExIPOcCaH3QKTRM+mV62rnXR2fQXySdH5Ga8+ExE3Y3t4xIOyq5HoUE
aSRC6Ao09+CePLuHxbug+er7OqCvP5A5OjgJXmd8qPTU2l2gcgvRI+eSFrQHl7xnzNciC//Q1CV0
2x4sYBg1DZIBma6NWoxl9vzzDRpPGeO1sUQf94n8mjiyIIaWQ6/DPeOg52qSHu+Mrrg9OZoQJY1R
gfEDxCoriWapItvv3snduh9fHFCEW/PRmix9HFfyiBszp1obzvOKRn3SrYk3j2UTIqwh57/E1wfl
27p59OU7ERER/T4rTkqorMchbAxKVsnwXCVvNXyoiitgrtskY+VYnjiAXl4efBx4X0f+6hOy84WN
QB2m1kTOpAg/6pG0n6Z+Aix2M3Q8lUrTPwoKD3YecgI2E0ePfTxQmL0+lUFR8vUdbcxdAtX9gb0O
VXNem5oPeBcSEUpoKMODegqbDanW54owShsircoGOGGhMpCI67dQg4rJm3t1jHS4tN2Mcroo0fYs
AVlNLLtrzPjOWG5YYCRqkRdKJwUsPn3JdqmPuVv0eiPZNa8CQJ/HBYrLL/ni1jDbWVyy7wRTio/I
b4wRzZee0/8cpjCT4KP7dpF2iHVqqBKCUPGdY7d7CIDLFazGcNe5KeYwy0YFCGIk+e98Kjh+63Qv
NSOEr5j+VBviolBCkBWo6bNSdOvbjb/Y2mi6x/HCdGZ5JVgF11TTlmpRSkQ997FArbSIG/VSvn/V
ATEd8b+EZbt+einKOEUSyBX1A120ZyXjP9cW+xh7ZMtxkBNIncO1kdt+HrF4zZeDEbWOyvcxCBI9
kPAN9t+jteg9dyUe+5FbS8NY6Ee12T5QCzOBNfBS1t5R5bPMYhMKo/iEYwnUw5l1CijyEMBkCbSD
4oALYa023VbVkNXt4R21Z9btpuZRgQalZ4ci5jvdBiFqbu6z4dMGqnjVp/MaUTVNcF5gOyWkXrws
ocp39wPK5xPiCjmMvpiZnhAtv5Bku4quqOMtV9D1c2tw2uVTl+Nopzu+njcbZfd6KpMEBFbWpe/h
i89OgW7xo7ATgCbZTOgHHOIb1QrC0B/YJd6V5K/F7JeenkdU14jR6m/kM/6dY3BD84MRMUNK2nPJ
DW447CSmIw1ik1Vd5sWryQEMQ8S5rGMC3CKkzEv1mTuU5LV99nmKMLkePpI4rnjbgQ2rHv+q4SpX
KLNQL0LRQSQIxD/9MhxUWS3ljDce6Pp1+0kB2xTWoStNlfcip2diBXXwf7A5TeKCNW8c9XtkHIjs
S0WfqRkQj9XFhsBe5/b964VN4m4hPfviJBVOldFj63J3Nz/6BdmKC2PB48yfqb7hig9JFcD8y7Aj
zaNEl2Ld2ARMGRRp57upZbfnyv7QFgfhHL/PBWoGn5cnevgSzihsXSpeUmcydgtreRlS6Y4u1vYd
aKcGL6Poz06SuvcBPaosbiAeWrImAnZ2dKrpVM3upatrmrFnQTt8pe+41XWC0VOb+YQb9pyL5u69
i/6+ePznfNL7gc7MXvqWhBT/VViMrfnNjh3qAX90cP/ENQI8HBAQEk/rlBCUa0zPIi/SvX/KTCFj
J1pM2g6EToIGVy8VDuuIMPVik58W2hLvFCtQDYS94PlbFkq9+9suZ7lR5BaazXGDi+DsSrtdNXby
607j5UiCnIntJfvfrncPVwe6MfgEU3fbDiYmIEy6DZm3bL/T6I0HPrBn81S6HOAOdWRAEjP/K2nX
8HYFUuNiMrhhwEVEkTDrnXxgBrbk18fMCM84fSVShz7LPQkvKg2Gjm8KkX7SUXXGFdSwNUcVLPYM
a7tO+28a3OJc4Eg1AMqqAVREyk3x0uPRZAmS5Wqq0fyrRuVC9CLHQ26wKhpVSRqsZTQhTSu4RXvi
qFmCQqxhPdD3ig9twPD089r1pHZJuI+uvqqI4mHLZHUSTQachCqnZsXEeDCXUnk17opzEf5NvoWP
NATM+4cJYxybsKhel+7im3e1oOKTsDv9rNEdbkk9ZiCQT+7PlbQdO+yMocbkKDC/rG3o2nJEuxz6
i03pUDZaOvM43A/NPBhMyHfNS/roSWCWy4lZlvrGh7qCq/BgIPpkuywntYh1NhYi8yahprSizxop
mywUi/k1rmUkXau72lBgQYG7UJnbevrd5flE2QpInOK7tnCGGUGyKmEYlZw9jmr1vWlQNjtff6Y9
a/vgLP4VxGtd0cI7k17/2kMhCj/8VQ89WfElBkY+s8U62N1gtH5Hvdj6uofPvIGswnPJmLOMfx/q
LKyP4ybZYR642Dgo5hxyvQdQ0ZYX+tIJu66i3SllsNTApj9NvkBPftGsvGGP3f6fDWYMyuwm2+1r
3U+QJzZEahbP+3wlLsA5gXb8gihRMFyp4tt/5/nXwrph27ExrSc2HqHhiMIdRkCeKUf3tEjJr152
FJzQt+MpmjeQbK+bXxfxF01Go1evG8taBQqa8pwi+lw8NLXuK1t0WT81rW9hhlz5gZMmp0P38p8J
tL5tEosKm3L6XrUrrPx17hoCQZHeSUb9cj+TSSOtVt1tQRJxihVC0ZfdrC6mM0SS9UrrnCJxP4e6
/gxWt5Vsm7eVqWNPrhD7jV8BkD9emv0IbP8QlmiLVWku02RLAp/NYUkEDJ1MWHIsnobqLXs5wU0P
JzGopmBZHFc/CBqLzpybBYRbckcmrmYqKjn2Dkfqzv8iaVzk7F52K2PVrrNwlCbAHW+SUosVFwPR
o1xt33l8Nu9oLWxTBUwopDfTNecUH7morul4M0cwx4PxLQTRLLWydcqEsfdQNqLph4OPTpoapfdK
WRaC7mVHhcXHm1tr4F1cnzwp9tYD5aGUyu57I4Cq0IuW8Q+W8fXseZibPekfrI3CZNJGOH1WAJuO
k3qY3GWZTtsYXxU3wHbErgYNvgorN42M0L5jPOEYZpKY5pvcNJwwbGbFhy6wlz55SBK+6+W7JIrQ
RdM8D2P/AzBb9netyVADe4PmVBJ3yPAN1HKt0U9ohhyeAT9EZU0Pv0X/ZlOswKHulPq62hRKCJvO
dGCk2nUeBMrB71PjI/sx1f5CPaqxytVUJkm+TmpV8ChRQsvbpQN4GgFppoUOBjkIgzpfrG9hZqNj
YLovf12yp+PvtcnA5/LhiyjUZNr1jW8YhYn0C6sfC2BmH9lW+6jfcJSLkHx7/Bbv6S8fgZhOIJhn
toLeM7ZGOhnzNtnUT2unLbyscXP5uOWTquk1GiLET3j1El9We6sG9H9OobiPBOst7wNbCCtUHQs2
GK+xH2NrUfiP4KvofUYwdS1C9y64vF5F+Ay1eUz+gP/Umd9bPmSgD6NlWjjkUJ+oeVg8nqRQw5g7
kSKDCOhHSmI4OSK9AJTV2d+DRVHmnXk91ILAg4EdI+HEwiU33AH4db5n7wAXpazS5E1db2+NmX1V
o2TgmXwezCAvhc9eM1hq1Q2CIXPNepJyPPwjaKoaBbXGOCiO9FsqXkt6zECVKCZB/KFgPuigrezE
5hl2duvq7UAHKw6Wwi3XC0yXfnBdvW8yMVxvUjS0k10oqjpuBR8FS6WvYcxDFc/eLu9qCHKTPVih
CC+d3W7m6mQcX93asqjcdNUBoijdeWjWA701WrUcWu70hTPoPmNtaBkN8ndIwLVrSU3Qau375UZC
0xI/7S7TvdIe7lyn577eOUPGQ6YOk7Fkk+EFnYpvFRiEK9pWpTayRh+ymGuPpPNak7jEK2iX5n0M
BxpD7XCI8QOpT3iakdELpoLD/0hx73k1I0bWfgNpjusfA++9FYoZh/FU5wqs6goukNOoZ9lhe5PT
+gB2JXNmCb84XemnHNF+so8Qq8i/YY2jQEXuWsTsOq68SdhPhKMhvxKy3kb/d4a+OSem5w9B04iw
eXmtkhes6TEeE5+gKTBMUIo/P1gRSaAj40WM9AECEaaaPWXqHqAfV6DRXoDNTMpjKYtArEHBQ0N8
QaWZd5Ro2VZqCcmnqUyT4t1IJTWTCVSraTkXRWCsxPs50dTVFnGdkN8Ofe1EONF68i+on3BeGvSe
U9/BD+RHM7u9OqYpHvYMXHoP8ivMvR/BCu99I6l81VgDiUi0ZIq6KGi/cygtw53Y4r/n8u7FqsrO
Ttp4/YgSXPCwlGnAg8GIAlUfX0CZJxXVDU2sJCDvMfSgP7clOilHTFGAF4rSWVSMpm3srn5aBHqR
y46+5OAYtYTu5X7oGOSaEDYniXrWRV9UO8YY1eRFkO5WnFLAxYDRdDFqQD8x/9URMY1kf5kNDNfd
P6186NBlPbyBFC6/hdMqF3PI956bRhj+ZLdMkUw66Dsb16ch/dY9kMP+9wrB5lvId4gacJ6Yf3q5
yijv+pClVPfUQrKG34iZYl8TAmTn0eiiIOqe1ORqq5HPnrMWYh2ylYHYncoEGmH2NBtnlPIwkeGn
8axEGxkJhnUM6GgJpS8eze2LDBR5G7RDJa+opsn5p8f3UFC0Xc8cbc9oXg/PWAo8rQcHE0YSpKQs
qDNM+O6CHsG8BaIzIp6ZvNwpCss4SGRuwMy6rp1Sn5EEKnlWmO5d9opWzi1DknCCDSR6I82xgB2G
NQvnseW2mxMub4Ejjp9twXLu+Mll/aGnsHjft/A4XfvBbZE7MN5e2Utpu7IlOrBNjJjCbzHcazTM
CbhxOiKRfVBC0HtbU/OGey9j1Nl1Jw9ouhjX9410CpJojlnPUC5JLefKefJ08ipv875SAVCCZt/0
2KcmqccDCM232sYKVPw1+z1LWNNu3kLIptmMHZcu0BET9P+SraqvqdxPsmO59EUsy0ZhhjBEpqwI
rzry7ygjQ6cXiHIIv6f//mRDHrOddPZYhnTncFvTJ77S4YkHSMUrPcNfYIiJKEOhxYA450U8AMkz
C+dxFfKho9YOFCsjTTdNqH370akjMX3yEebfQLz81kU94xTZ7v1sJbTtZl0WwK0sara9lx5SlnBp
iMRQcO9TqmAxgz7vWCkdwe6P3bhNCRCb15R79ohEiU49U3wWq5jMqeNovr58BB1SjWu8Ak3QtvIn
4L+n6v4otU0Cy2IGPM8ccE/MwPjLVST69jQ/xNKCqEMTVCKuDwEpqQoaDbYPujwIHQMi8wWZGg5J
YcClH0iglM1Ttvr8pNkyRiI9tSIJfM7D16B+viot9TiqeCGSteGtrdPxIveTjJgiHk1jQW+fv3iu
2rSBFuiAl7VV4MlThK6cErKDPVGxCjN/xAfKN2+Pn8HBz8IqvYfw4U9352QwpyqxyeNA46oPITCw
8cbUH+UGWRKwgs4k2IBLRIW5HI4hR8/m6qercNU+PGXkSMeJQn+JX5N77uPiW6INFZQafmqHSNhI
ogcmVwGidIVcrolmWwgvWID7e6vu5ml8+SWMjGx+vl5TgHEsStpmgJ6IVNh2qBhcfGQLdg24pIJ9
zbeCW5eO99erz1LM8VbsH10xKpa3Y+Gasb5ZQlM1PQCVlWI3kA9rqr8GstiGS+fZSQLeHzmzEzxc
bdpi9TO4w/GJElMvy3VM2lB50M9Iz0oheeONhGd5RCma0KtGerpEIZikojDXNKdWP0ZTBdgL+ucB
heIrKDaY2mJEPuVLWJcxIln2qyzDWbBbE1vamUhwCanZ0kqHgySvz9nxG5TtY0HpTAMqsGL1ifPO
w9N6heyqJWzm1shJaoODSpL1P210ZFaiT5yR07i2escXm5YWLXbQqQ7gn+ZXkfhUZue+/iGR2JqN
sNygs2rEEjIeF75jK2dua3Oi1+jVZWOy5FG+scoT65rVKzRYP1+52deSIgF2KtPVWQuWnlgjdK16
WP1zLUmLR6eOv3VPxU6QIOp8B7uSXKmPv6p3NWkfWVj4T+pG/1ALPIeD594Ikx6GP3G0cGz0pQtr
CnjuHrtvAr3NEvY1sUu+XnhoC26FpOaAzMt/07WSXm+a93OxJni/ySMXAncM2YL4PQ8ASDgLo5jD
YVk82iVIXkIl+SoqrHmn+5nuwCHn2Ur0NDyWlctqUnTgSaXdJMs5COeqVd8oWu6z3AlffRjNxIiE
WIxm14Z8hZHzcQz/kCKAKj1dZDtia362vBoRAAhjzvWy3AcVrmdLH1I8GjWaWNrnIH4WJnhDhDZj
7UrdkvhyZl3l2LNeavSFj/2Fi75EKW80kCXH6puTpWTbVEMeXOTJGuaS7H0n92HkIN4048KflpSO
qu5i+RHeEAA6k3JuGAuO/QuatOfWB9+5dXSqdJAUsIoX3t0sIasF0ZaHF1aVswk31EJsjSihm81N
SU39enY9m6uz6arUCoBbeznsdAqQOxfqPfsVN9E8D5qLT5A4k+DWuwq9fzdboa2vwDGizCgVP0oQ
/L4GQwzO83cwsokTThEsG272qUYCzJlJDpmI2UCxZbNqhoLJQMG25ZBPy7n0UMFB+Sz+z+VehoVL
/Z7yykez2TeYOHV+dcGJjykh9AmJD4ZzryoS3QGeQbT9g8OAhOAYAbOHHh7psoKC5rwBjWt426gV
rrEqMOFWmC+MFOyEMMfB+N/sEEXxxCnCkPZWxpRUKO+/vyvdj2OfoiThugKPoL0EWV99c/aDS92Z
o4QK2Eb4T47DemTLJNf0XQfL9HYD/RfX6KRWBLrPCrjH7/gTpsgFCSh3SNtK/31W/mlQLgJDCGc7
23I569vtiUjrCUzWPudFPuZgRr+dZGlQOkuDMrQO9rAeA+p+2FYc9O79qDOvjxu060rSobLCHFsy
2ubu68KJP/zAHjyWiT+Jjvm0+hPHh13IVlPxQRjyc7K9g+IMSgyDz/BmndCE/SdGfShxvP5iJinN
q1TpVk0OgIIjaJt9apYsHwsZF5NCVQA85yFheXvUWzdOJXnQnc3LSWIvCzqcfarCy70iV0kWulBe
TrbBwbDrbvYf00nMorZSknE1VrWBmAs9fWjbJqFxh6aPHH1G7iNmyx50jG4zF1raLDpfWOWd2oE2
keH40S7TP0Jbqw14QjlI8E87+mKLINVi6dO/cEOenrZKQD1O4ol9sPnfvX5QNl/s35+ClO7Ai8Dx
exipjQmoLDk9/mPNGz8IEuZSN/9lu0qpDnqpmBpYmxX4g2zG5qVu8hT72CA6j9HDutkf5kk1+Jo4
rwqiZh8BG+XnV7/lqBWh4k5l44B8nc82Z0rVsXKBoCudQqsIF7Z0CmRapJsXwY2uY6fFexXlxT6/
2VKDs6+6yLhnllx+fX/o6aMxWAsSIA7n0bmInldnCr2xhQvvowLBXM7T5pZmZ3VYQ1NiCRCoeTSH
6C23V1ZNWpofcA6kR2VNXkUE+z17+oPQLnf0OI8+gbKfxDtjCk1Wb+wbmfV82w4HiotURSQKQ5kj
1tXrToHtsbBD6X0iSyRULL+R9c9+8pgvbzGpwQ4E8uOotb3224H5qTEtSV3/tDgzHACq6F2cmnAV
/X+zK9O7xE5n1Xq5HVOqPvVQHC8/o4CceI9edW8X6YlR9BsfYwID9p4EeOwnquFVEG8Bh0B9WJZR
pSNuZArYIfnkwpJmsUMLLOHxlTbGyfbVaCk9JvVK18YXeKbUKfKEfsTi4spuxwtzCZzulPTq0i0e
pXXc725ud8HiwwK7LUPBMx4O78bGSizASWmQmnNDJ+aEltYYYVeUBuQ3Tk/RVisfNOHAYq3yihuj
b06/dvJANi7mwLhu+v/oUKpxIGgyhfKrKNncJ3WadwRDgJoGOliisVbLyul29IsReeHLS0qPfiCY
EPe6OWvtg504QPbDDcudHQ0mMjm3paxVpDTBx5tRY/8Xf19iwHemuSTgQjX8xcAYK49s36V7M5j4
OiMgHswUbk6a6QtcgQusDpjaoE8M23zqbhrmTbE0jQxDc1VTpvwN3kNdsa1zSPARJsXaAyMmmtbP
/85vBcuQXy/Kk4n09a7UJSqVGMDRyrIaGNqOOQ+yiDPeazzM5ZfD7uX4BCLH0LUh6pvHySQF5OVb
76h7gZwfnWufs2LF66iH/6K6+T61gboX7JVBfQN5Es+LjHYtOpMUqRTwbSTCE2yGUD6M7+BQXwM/
ohJ80X+ibwwYCeubGACotKeqYkZ/orjHnXuacr3owKPZmmlbmFV59lQ72WKKEPYIqxdRA+f7E21V
xM4tphol002TlEmL1gBJNwQNB1z+u0ijVv0wmQetZOaVcpNz+EBbfiVb3ySBWrbcCNPcLUH3Rb8c
hugypvBs1sBPZ7HC1lURvSD5Wn/fdx9nRdltxEgC95fZqggUArNeSlZApm2arffjltPHlloZc61S
DKhB2n366lTjIqKuHzfovNpC282VWungBnFOSuBMA47Q/ZTGkFIIg/h4nwHg5+u1AG/5g3NcT/G7
KMpy5WIMIiXUlfAg5AyVILzsN2BxuhLbdD4/90eZh4nivyFZaSTgptbTKoQngtmN9UPWuvQ4nrLL
7FzGm7jwN0EWS7sCVaNzNcsSH/bFWooFsvlJjRfPH5amfdv2wVQC9lvomuGHGoLQvrxWh/3Ihvzk
a5xEAQ4AnWeFY/Fh6EisE+2aPq7QX63QBmaN5TCp3QpyeApdb1nUj9OKyLr/Za19IFDzzXlDQKtu
QeVcPeMug6Vm7UX3T0xiNipK55MRWN9seetzRnEhyzSMWNcYmztWkLG8hR6nsA64loR9o7br9asd
dVqWG2e3qxERQjy3ARwmrTa7jJDTBj4pcyRR6Npdpi6vhPIVO5exlUNn46mfwJy3tSJlvleSPq/4
DxNblErSVmQNz6QeEMh3NaSYt1RBP+GgK0I7j6X9oIR48i3odMRklEx51j/FTsT7S5NIhhHQSxZp
YAeMpJtvKMzprO8Sa2ISGL6lrozcTPFBFfYuwqoh53kocO//g4D81YhTdfcV45CbL1jIRtH39mkO
p2qGqJYspK4vsInOGymg/rJG3SiO7qLpmoLYKKcaZW4B7Uvt8LNQgprCUQyYA7vahPPaKqYCkP2q
+6FC1XBDd41QpiCeH9RXVkMa844cfKTJhhZt0Be1wcHtohejpGChkx2VRA0PwDqgy8DFMSb7+LcS
z9PkgwmZBX0x5Qc2geHmu9m7qXEoMdM0nzKleRv2KfamU2NVyIs5OJKkQmJ6+gEEpTOqdJAh0/Kb
JRRnAcs9r/VUu0lu2unEM5qBgyX3ajAdiY6udVb/Axd/ibaIKTHlwA2PnHSJPaVcU2SbI1DS4lUG
hkIk1zepmV0JoyMPuA5UkUQM8rOuY8PfUc6xzk5bVDwtxpoSy2PVrS7wEXW7R3H4ZUdBemDsarWy
umrQ4JjQcZbETBuozD3qjhoIdSDQrjq02DDP+yn81HJykup4V8lgXPLXqLO2qFCiZtx6wAkvpgUm
NRDOF2byIg9B4Dt9mxP9I34UXGOzBZIF3Jhr0DJiGJ/1pLm7GFVCA2Dkc6O/1PqzNmdw1nraP73o
BQoKAnM+7kv8GmhjKU3dKML19Y73S9gmzwjCqT6HG0n2JDqUOLQF6cYkOPDZgMsKX38ewqhOUkCl
vNTyM12CkaL1KVODPy11M3PCbVhdzXDSJ5UII6BTFqLFnq6oNngyFVkB89xE1HIF2q8Fo/5QpeYu
SxhHRRDUrACRBYtF9v+g9WfS9+/J0lMTlvQUtP6bX6zMmJ7AiM40J4lBGZnL70s0um3/G+iY+iys
54tB/W4e4P9+E3FnUjLZjn4n6GCTLK2zUNp/O79ksO/ru57+5Brl3gQvPOAe252dBJwsdvq3lewD
OuiSesOUT9OwV7JLVq5RoW+Ghg1qamWIfz51LHJJyMipCnDHd6lkCtcJVkcIy0L5tmpaQRNsY+wq
hqSBZ5uQdMNZwMvjeQGh0YEqQg74eBbeTcNAKKewhY8dES66BNcpM8QMJrF7x+qmFPyvTBZ7TkQQ
xkVqN9hE5rHbe7BeTlb0I/4CIVjPlqZiAa9TEL7TNLYZzuKAju6gpWieQOvJ35ME9DFNLwF/fym4
3qDo/2qvCUa8AILMukTQ7gb38OP8xkmGc/qRgYZN7Pr4nGUG+4W9qQoBoz/jvHoxCdnbCpoAzKty
aLMLSa+EJyTIgR9Db2SVnkg53K2KN/40P5mUjM8txlNtLjb+Jo/u2PiejLffJ+a3wQ9a/twXNlif
3h7N8nkExiLXexcHTytk35YbdJeDkyJCvguoNN6Igzwa6YwoOVwYDkqiZN1CMrCgdyz0MfHwzevv
PiJ0WfZwrIBybidd1ysA+fe5Yk4GuQ5U0E4+5XxaT/4Mw8DeiVQ8F8Ccgo0xMLXzQ7p4/B+WojqB
nI/XPjTDsnzJ+TjsuPjKueUZRefsPcHKvw3JofVR+n8AhpSLCVcWVmT6dNg/Huq21fbJGn+D/moi
SmqEdMz5Yswtw98ibLug/DBW1L/4YzbV+zNUgMFyojsf2BlxcdIYUo6TO1AKu+b/TTS0pAusiLVA
3yhUa6ShzTTGA3+BJ2haxW/3bTqHhmI5Dr6vw2ThT2O+eYA6mUALIvtvwPnPj4prR2tLgVP/xjR0
4cMS5P8xlKfmZMHXSgFQ7x/2E1jR8W1DFED9dc5IwQd2vvofnguQFaNg9ITkpmAyHcQypDvU3vMX
O37AVIcVYRed0pScMhX0c9QwiQThLwqdQB6smmM1DD6rzuTxpmTFGc3R5tI3ElobPfpOK4KN1if3
wgBWWKaXOgeyDPlbAOLSAEDRRUmR8qiVyCJGu+24GF0+L+gPUiDNoiQiZQHd1K8JbTyC9gsMfW9S
LzRIw4dVjIfvIhh79oHzG1QQ8Ll4tWVdMUKkbcCZVQcyrLxZUqFjD9ufKhhmTafdKc0HWI/sLWXj
vgvRv6Hb8eYzpmrEKtaeJEUdxb+kZvv0pMZWiZt1g0pIGykgFmzkpBia0I3UaLo3ItIvSpSLZmL4
QTZlQ8XPD1Np9j/xmtIPaC3Tn9OJjfKSENB8ccdCZU/jBj14YgCOfirF8LXPmKa/2QBs9lnmDVZw
Zewk/ECpCq8CPS+2TLIzZyCbwVU7c7FY82Y0LQXOqO77BApoQO1rNPohev/zWsjnhu715dxrQBzs
S0X2v137hbZaa+2jGxqgA3Yr0lc/42tmlyOUCkYM0auvMI7WB7HhQuW2hWbBmCnYpjXzy24qcxlx
zs9v6CBmIlHkfoxN96kLdF+1y9gOWPRl7XbBdlAawvDzI4jE/dzmkOdsU8xOGvtk/JO7+cx8Pa3C
S7K+F+zrOzxju0EM57ioa3XlBobDY+9yM40b+sIKC3I+RUd1Q8Xk+YKjbcYE6eXl++X6IJ/sHjdP
nuuf/TRE6y1SrnwkTX7tKafWchUqhr6k8DwFN4c3rGmMxVIKTeNpBthv5wOKIGerhd2FKD5mhdxd
7efTLGk7YsXObi8yKEmmevArnxDHfIcM6Qe0xHZ35vgkJGruGmzkhnZ5P19q8bo8Lk4WTxmJJAPF
Gf9gvhpeb/ChfHHYwmHqaNilJNkW1XT7ZiMAeKJjUMQDhgMth/PB4TFKMXtGncRtTdf3u7yAcZgD
wtslnewLBlLeNxs1iWjR92qnC6mwlScfo4dxlDXmtCKFSHnr1ABNr/34p5TO9PcCHMesYSgyIQod
whCBncW0aP+41T6PtwuG2DkB1roCg2633X2v+FdiLVaEaAZAMvlPzu94wwb75zZGciIPoBvp4q+G
yUKBltJkYD4z4a+lbNrUTC691Yxnk4DM49wGy27RmJLARvENA2igNKtj+OqkZtc+pFDTZ7Ty/oBd
TxdpgLqyQr4pDXMDUvma5sL0YZChWnF/sCA/Ir8uAkLUFANCXVC9Sc9PBA6uAX+iH8RUfTJgViW+
p9tMpnxzIPTlkSFewa3PQTLqdKtoi5wWlVw/4TXga34T6eT4zX3n/wNH4ZIpNgPId/5vrqAEQGTM
4SMzREgQED5TbM9z4sGlyYYc86T9lkgJh07bTm9ZTUTt2lMCqyRqUIt2El4ryqVzM22fT+1WGEEp
UAxoZ+gyl7PC90DhhUI8lgSdktsr9v+4GTIumli0VcaS77vZDwXYqf2eiiEcE/dTi3MjxXMUUNWq
gPE4CUa8o/np73qEqb2YHoshQPqn8SLjVzJXy/FbrpQdjXGHi+K9Tvclu/Y1pjN4J4Ul9WyeRUHM
a+6MRuNig22A5sb3TemsnYA/YndcTK5NNpkW4K4Sur5hNL8XQslY2vJK/zf/hPcjnExS8/yFuNFE
N4gyinFY0ppOjLl88C1lJ2wK77Uy0XLmxX7CGS7uUslpRuk9w06aHQ/0laYBX4k6hWkKGZTX4/o4
aEpYNhl2DrI1IOj0RUZEw/1WC/9RFcDufgiHmCpJsW8HaVJ+OJIQykmWej7PODe2tDW/1F6GA4Q0
Mjgh7TM7CSWWfJUt1qbY7MUAsgQw+KKoLsMXMI1KdL4V6M9Yf8tJ7upcu7D1UqPz51NA/KkXwkgM
VRE5jqx7lVkLgIm2A/arevybL1EYk7cP+RhMbVIZQ+jEUpI7SM5xfw0Nguf5KO9jIckgtXq27n5Z
qSsWZGOb7c9ouFyIWq6ukna4wvjkuRZ17jHfKPsBiy6bwMhJBFa2d1VA/XeGty+ev2Xi5NoeeP/M
gQty/5KMLLUOhqaIcqVMH9dQsVylXenLCLbh6nED5xgHkKgdbi4/yf6Knkc/Lm+7vl7P9ab0EqWH
j5i6RCbTFDVkxrceefJ41SYCUiHuhyHvepJ4bZUW+lHspxYbMhzUtKZh1qmLMqB/G5ry8yVi7xHt
KoVne6FLhJ9JdDXG+vmZRl3z0vMCfChs7oe1UdTdJVKLzjGUUlG6EJ2/e5f3iU/wdZykkr7XBvI4
pH7W6Bc0qL4hSbK0FeYV1KenCEhCPd31XjUbx2zQlH0gxpIjNO/Dsv/RwjR7NIqEg6xhkm92FQMi
BHXzW3LpZwFY28XZ37GotZLTAzkeOjvkrAylb31VGQnLYtiuBDnMi9VGWfdu+Tjdjz/tc+YUsUuO
wXhiUagUGvt64XUjUYRLVtzv7n9WoGp4vpuTtHABOhg/QRcmV/BRsLQKkF6/9bAoLDQtj7CsnbtH
fHhazfOYNuud6UX0ytKhBm2O9wkh77PVetlyTFfu2CoG+W+kRGZ6q9pXrtSKnyozef4I/ZlaAUc1
OHLYMzc6z2zaf6WUYd8xOeOeSxu9oW/kP1nb9fK8uh5xbR1MRFyNWezHJ2rcON3tln/66EIeTjlN
ca4bkMs8fCCC+oiFWktGu/Wen5/cC3uvqwg+/6iKCVaEgjv6C+DBWf5mwrIbx9GQwJ6/AuQeRcLz
f0yZwTk9a7YkyPbWIGxDptMJK20C8hXmFZfYcMvHF2upgsvHCvZbFyIz9xJxXzxzL/I4iReF9Wfr
or7UlkKHjHnV3cp3vs6h9nE/yGtLc0QxY/OI6KWN+RMQPm0TIqnoSmy9vO1eXbsd6eDwD8lGcSUd
IZeKNbllPQcglr+QzGVTocKE/XraWNn9FnfvHhpb6WCoFUJDRvRoiRWdB4oIRD5OY47CxxbIhbji
vSH8XxixvBk2c+t9UamFaXNyt88z/0i/Jj05EC70InKmElLwDY2VUt+SGJnC8onGjZhUH6IhgsDf
p9Mn0BmQXll0ai0KxuYBDEAqsUcQ81gNAlj7hxu7fBgk1Gu01T1wLnPvgSdbbkM/Y0xX6hZkvLJH
qW9GYrB+tDxTlXHN4xyxzLg3NFQuvxMRQR5l/C1X/hdr/usA2hjt6a2FKfC0GgB7Mnx/A5akdk50
Hv+PCK7wjTtqrx4yoYYBhsww20r60hAiCmVMkipxi0bgHi5juWLrk5pvmtQGuUYBOapTymLd0ZnS
CcUn78kO11DW0jkIUT06zVydSGKB94If7TPsdagii8jgnIjexOSzh1rsusC1FHgyjG4OtxLO3eA3
+JaEnYFDu84FNz4bxM1y63aPywGoL2ILMD6rmVx20V25f7H3xho098v8gKU06PeM8Qr/LLLTP0Wg
0tqY0MOtjavrnoqebFul1JJP3gVBEzA2+vtAJiTlcmHPya2AYUDIqCoERlCI6zxDhdy7RjvmWqZE
ipmdByQjipv+jyx7v5fcYtrWMSwrBwYpzeIcwJkWkESViZYX660APpiSWzi99QJtaUf+/Te4VUU/
dWBfKRDQgSyuxvcqSRURa4bU+449AnNynxLxUFEHdArAzQQXlLBN0239E+Tq2V6w375mQqn+el8Q
v7CjEBc1O6mskyqM2q0MukrKX1k+vFD1jObJZXXqsgE/+GRY3A8lvnhjhM4pW55j7A4I1LVcxDSy
uUXCyfC0nrAj8Rzq0W9RC+yN/T+Wb8XipBOuiKKvtrJ5cEr2aXK+f3tHvOtgednrkEiPK7rixpBW
kS6ORjjKC2znwm/8cR8qVmU/O77JRhLqJqSCdHYKwoE9IibnbHTl8YCnra11dxyJo7iFMztRuCQU
CIXUivEhCuteDW5IF4lDyhXm3L3G8fLgy8BWAZK+jz56t2DfrOjZXXINNjc+PUB0H0VnMBXfldpt
3oMGq/sYoBWZjFR1YWZ4wx1gS2SBl7upuxA1WAv4dXeUuplxGzvBYxuqsHdEID5Nt59itCcfI0wm
S0shPeuXK8YQsVi+XztHvo4iuemzoIP/VOp0EM6gZFmTagxDdQFP6lpPTywrsBrskm2EUSAAY6/L
8peCI13VxW1fvMS4asl9gM3lxudGMarTdZQ9JRr+32v2GK63/86E5o+/YILYE6WGuu8Vr07ymJ+M
s9OnYu0G+cORp01yPZpc24c7F4OT2KybAwUP9SvVsshYwpvAPObYlaXvk7cXsxugoWX/dNlnRJ6q
6Pw7nMTVlqANIpJecIhjnyLp9D37FWLz64ZPwSoGWA9Acq9MqezlRkZAR2Ji/PGz4Vxi+iEHyh2H
Cv0hDs4v77FJCIYBYy28isxyCM9nqVnv4gjv9J6gmrRGeS7xgFjax+VRHbmwESL4+ekKwJ5Mniko
SCPILt0mmPsy0aaADg++E73ZGrJBFdLftWO9MEnC+oOTU5Jda9SY9ksghEjqX4MMA9YvSJyrz7Sc
wpoMVyGpL6mQURg21QMT6oRC2cFDIS6iXgNfLvceZzicw/HRCXvJpSO0/qhMqPlhvCcz/tIOJV2j
eTWjeVuUuwMNYuezL7DB4hqhtblcJ8o4h5IWGBlpEjVXo+52+OcV75+y4e4v4OmuSZrJz8lplE/A
a+1mjJw+XDJ7Bp/tgkjHFRCH/FX3ttyHmkYKrz8eXAW/L5sHC3ZYYlF6pbypxvlD2PZYk2zhDc92
YRsB8MHYjoY09SuK08w4ZeJ2WREv9gPQ+jXN5x/O2D/FTa4iT5ubl5LsZ5JEVCZ/qxaZmBhp76e5
zL5XPqzCr9KkXpyl/XagTjKEboUMAgGv+ggHMDFcBH6JhW0HoLN5PchFVVUgmGKvn4JBJ/UFniF2
Dtmi2aZaHovxrAUrUAnRS32YZyS0bqMkKfUc9TzyxvMAXQ5hoB3AvPBqTqgNSmLx2ex9ChMzRpN5
Ko6Flp6/hFu0jE9CKqjc41tMSnEAkrwZ8BV4uQrzcHQ+Nr8EpFl1BkhgI7Jd7JzrBm6MJqdsjKgS
KEHjDrjX66aiMMAcjSF8QA3V7qYgLCRhGqtv5l6UyXEjSJhdL0IGX7QVHs5NYnFdHryAcIXNDd1i
L1wXO/pOJYJwKZvpIslxYsCmnJPEuamMoI9QUlrbQi2NMTkL+MC5L7UBaZIQZ3m1npEwe+3DLTa/
hag6uL/QVDfuxBZgeK6kuNrEmJlpacXIDS75dtxxN9/h8r+um7I7rONXWuVqzzTTInCXkT86Vcky
kNxRxkc7KK6WlGLQ8Id+yM3i+k4WnTUEe1tt1a2lPFfxcBHinkVfrkHAggnFe8AIvQCa+4mnqe5M
5A0/LoSXz67a4Uqntz1ozJE8EcRY8JDDtG6CQKKjkJjT1ROHZCElM132E/now271Gk2Im+Q3Ojj5
yAY9Mfi9k/COfVz4+1pNO4Lh02PycXI9K4T9HKYP9uM+eQ1tQOhJz0rGqeY4RkvrgjmTDkF377n1
p0isW0f3rKf7ZZp90EWZEYRvdAJaqksbncp34Bd4GS/NSGON2mDf8g45fB7GV17yTdFALHTBC+lD
Osl6n5LdnxRFohNRxc7vmbe8VFVjbrz4JaetXtp/Wnu4LWmXKkFfGAynARsxH1/eGib391r1D8sp
tELTxOmW4ufwaMVaMKdZJUpwS5INRto3/ahh0D2l9A/vY6m+nkd6cXbaQ89D+XEsNYSo809aTS16
h1mJHdAl6VBMgqLcfEVW8mgARcejRB57z1OU2A3hbjhxtClES/6is3PPT+9gKXLqh/5mVVwBNmeL
P74lValMlWrmds8Fk0q1EaF+ZtaM55JsCtwXTqXykTb9Q7+TS6mx0oaomREGZmDBs4yOUbAjv0vX
T9yqK05IL36TZJ1A13asrEFyIs7O4sTJUPXpzAcaiWdauRSqygie80MJGDRuwPbcw0lYS39fMoJ0
PGisu5V28dMeAB+UWuJ6KYwnCi5r1Fk2yJIWLy+m6NEB8iRup52XND9oX2/jVs44zZf7XN/ifZBL
b7bDrZz/0NzFxaSCuQeZSRG5MA+3fX5o66M7HwPWO/40cpVkx3B8U80uaKq234cvvAZJpc8I7Ie/
U9wVxpN2PW6/4T/igjh+NhXA3zN6EL4aLPqd+2uHqeobpUii6np8MhCu4cimDPTSYmUaA7ySq35T
v7ItV004K0PtcEtYUC15C+8TiLnB7Zo6isBODrSs1q5el521KNdS3DHMiryFM6o3li2aH8xbCQl0
FT3UCNc3kGnLlisUagCjica+rRUYQ+024OKm+LzBPbUWitaDJ7vXCty8kTh+0nYqkoIa0343mlGD
UQvVnXfrkFuf8s6CNV68vPKGqyAT2xmMBXDqsbOCBjrK/tPJavqj4ofpv0dhoryvx/XyjpVnoLwu
f7Bw87U0kVv9Hx+U8B9qCncvX7UcpMnpb5J6ALW3K65MyMyGAMcm+EMuyNREnQAxa7DNPwxGHVou
DNQRWMLXCp3KFTCIo10YdzKnjbeDaJIVkxJAV2PLKRISQLF9LprkllxXdqLkByXyV34ZTP7f2yk2
JK/yXzGYvvo0n0ccXkS/U0Obg82i3M6u0J2KfwgUsMGpbP3eVzCgkiQ6jfloq+uKkTcFABp6Qu1P
y/NHAwzpK9pptH6gZEFCycBg1XK2FVXIpWWTn7sbIBVw9YkbY+zVkb4/yID/Dqg/VPHzLoZyn4x/
Uip3H7bp7o/VdeCRN5nTukkj7GzXzuzogHkbYuOZXl4xm6rUslWF1/NKC99vpK4IZLa3y1xgDtgc
hyj4AfxXem+OIMg/oWDgKYQlU2Zh6Mmd8gs2cjX8IgEgg/EKDI/54wNgM5/von85fV7eTyzOQakh
R2uwbyzaxjfKesMokvxitwC+YitzXjwAKPo0w2ETlbkKuZvkgQGKqLNrVTq+Q4snpe9ErHFgMAHa
NcUToaSAGqD3j+UgWiPvVWtZCq4HuyZ7O8i7qme1dtiMUPM5lGVZVwxsWDY1w1RNVB68JwZeJMp5
xG1is/HBiCz4e/Yt0AH2TPCKHdYU1Fa2YJkYgvjSdQ5mIegobuB72oAEhtlnG70YKYksxHE5igCQ
uYflKZGG9P+Uc/P13k73uR1jL8gSZKC9AIBTJUZRG4bRStzgXZ7xN0fQcaDTeifb8MKLHpyXhURp
7SMjmKEAp2/QPy3hAmXLeD+PwurK7ZGgqrVb50U6Tpa33BB3yhs5eyrMV4j+oLfNAVBOoi4w7+/o
zuJDikFjSdV85HAaysgoSKfWp4CbY5Pu9ovbYZxl7nYyg+rqke5xN0DdtRiQ2n1sgiHP3NKrrwsl
bsWLDliiO1TSiD4DNIDNC997Aab/mtW9qO3Csx+1VXaASHxVCeshrnPAS19oh5bS2LbhDHUx+QfZ
4qjWd8Q/BVQUWaDRAYB6dYe+CaoOYEywSP2y1RbSGQ401rYi1RN+5dJ976Yzakjzg9c0KrUd+nQG
HzDx+8tWHnKoTSCDTu5ttQgwxsnHp9a3QJ6Xoc6A9LGH3w4EWLxdnnM3kRfKc3xlZXx8ecE1qEID
KK3YBl8XLfZUqRF65wMvht/0zCe04DAnxL+Fwkr3lGeJ26DAeADQrCISfhk+GDkuC8uIymPjpCUl
H0mfvIeUifThTAoQ7//Q+VQAb2rqEfDbt+Rei1P7fcBLN9kvPVaS1Yp+kEkRBolcweZiFUI2JiEm
FNcLE2Gs5WOeN5LZvBDnmA6FJ2b1ftbWbIxSTqNoHIDUx26fLZQnIa/Nm+C/+SHzaf9vTXjGA/o3
QjlxjpPkC17e+Ju5dZvaYuTrvXMJq708Qo1O5LhG+Dww7YG9JcJZtniXsryeAUM/7Nh8bF1zgz/E
LCHMAsJlLvv07HZI7HrRhp7GGzUSrsXTS5q5ILRi1qf9/yx6FnQ99XsXiu1Zx/7IB0hSdQL0Yw+a
wWCtXHiVgfbQHWgbZfYrwZc9SZr4+o6juBzvZBr3UWwZ0KjQZearW2hl2GpcpZJgKRCTCeNHPYmb
10h9egaeVDPlNJASynSBBXasXtn4uZFLpg05yARxfA+goEMPboWyWVg1ZDg3NkTDoV2WszhvGMwK
3iQAgyOaO4jzx1JK6TlIz2EoyK32yEFnuRngVFjeSWYpHS/QUC7O6o57tJSZFABn+hjUysB0T7YF
VW+kHzCGvEepb8daMk+0ciTMQTOZmrBZVgHODcupEAiwOE6pFZfFr1NhiIE+vySeGWxjUyvcuvtS
w99JpVUcMOE3ilbMAFfBX2rQq4yovBmbYdfLPOwBlNFE6t1Qwgk7vnXyJ/Nv/Nm+RtnGiemDPth3
gbbFYFWyDJ1BEPLRMdRIjDdIpebKDIDt6InWeJfQD0HtfQqlLtbjqG1Nue9SemXw8b0wYTpWd8KF
1H0wCIZNh646ApBJXwKcR4nDDNbG/Cl8jR5AbBME6z1MXy3mHXrpq/Qof6+2jWD6IsBaKl0bs8ZR
ySl0cHUtD1OzyfwIxTXORY5GFib1QSzyDE25Ypf6b/noCRsD6DAqi1gxMSQuh8YzRLsvTDAxZzTR
UJcVfQvX4z09Oj7pBGpZS+QNpnWN53X5qYtj/qpaFmAGyeF68qOI9KhYtsOz8b0sMZ+XJtdstL9C
x0IoJ/4MiWjxgGhcZypZTqtwInmA7Jju77er/87PPDNcaucJcsa8AkgAKh72P0kvPw9hbRn4LZL0
EtpL0IylVRMDJ9HfB7w+GzRk+st/3g1ATlQ1mXVSNmYKUzETY4jrBRx5edeUd6s+3WEivrE0gxZ1
Lx7BbeGY6FacAIAWlgmbK7vIV1z5J/01bO5P7zCTzpvggekL7D3T9ctI6ZEsZI4lfl1bQEuJuXC/
uslE1N/i7La14S6i/ZTVXui8Igx21+BGDVc3EM3dr3WdG1M/uo3GtPSbSg6VEa82LULktBFBpumv
HRAbDdPKcHz02+2qTE+ThuX1fIwaWyzKWVg0RXZKmQdqlM4sM5se0DlpVwZ4t0eIONgCfIHkdOT/
St07ijySIbxpYanxp8EsozTw760TFqMVreZIlSeU6GVogxGWW+eEsVH7DffBiECrfFMJdlgEzQ2z
P19Kq6eckVVBCqQR4OUyK6Q0gZ6EqoehmhTfGgy6bHi+RqEV1L1xJ08nepA5aQHDkJq6AjfgxyF6
nQrQ8sFonBFIKlDWpgYBLbVzlwtD/XayJGaYHIs2a4RM9RMCJvFDYyPsmvWrJ6TyQuDFLt/TiQIN
oXqDeKGU569Jadbmlg8c7N6u9Ho+YvUR1KunQeBbSmfj1LA/fG5KfA9jfq3mXNc4inBehGzvVapN
48X2Txovqrq7irPIuXh/admlOROvSPWEjij7KXuiUjTljmx4PLSHXSU8IlwQhbKe3wH4rkgBA0zE
0JllVc7/CLEz/lFxRbbVf7t/bOv2E6iLZ8UW6tGCbVqJVXOatGo+p8kelV13oqG+rAaRrs8UiyGH
5eDBobdqwwqX4FTUkVJ9jchHM4kLbOX5cK2GKUFrFjL0spM7fbJQhiPceOtCPYYRjbVSCoriZeaw
h7yJPcH24aNl0MsZJceimdcizoYk4o9sZ1l3XBmccQhSEvaRkUNSAoOoPMf4XqMeO/caLY4OoGiJ
eyR/qCDA4vRb2T5DL4S5Ct8k5WZq5tIP8wq8J8OoT2J2Rh/MVS8GFLeGMxfLlGl/F2ivotT6S+sl
TzqsaDSg3Il+cu9NPhjn0aH3J/jlAEzg7xf8/diEDvNkkjWu/IyFQk6Uos3w+whFH05OYkVc4MNR
v/cHIYCsPTS0fdrZe2Qmh5xcb3kfSea/O4LCzjiP1f64/vXP0gWAArwXUmaXA0+v1NKeiODI7K7Y
n008SCTgCPzxjpttBaDU7sv544dVxWsAoc9PlF6Q1lu+3ZejBoYFHJOXAt1yqg0MKAnm8wqnsgp+
KABxdO3f/meoB/1FGrwYvt7kg7HstPR13NN3o9Qs/OaOIt/va/+R11tMyCtSQvad6yrFW6+jPsib
mkDDQb1GiZcBubBepNuIM0bW3Ixh+AFCDFhBNUezq1bX2OUANfJ3DO3+fPZy37+vWELWWIEj+8J7
OTIzyt19F4OJxfU+hbyo/DXtgE7FnLcjzp8cE54LsVBeGbFRktxbmZS1YPO7HEc6V1JIQ1hfYP66
YzRWf6gL7hol/XsWizkcZFpNw2PIuHsviIbzwXarHyHdELels+IA6/nFziZC2eIJ1wDKCiTG6Rrf
2e+xGPgyxUIfGWAY8GyGHPv3pIsu56yfhU73WOGnTpVl3dLWOpSMcJZ9gAfq9iDqD4FelAZYR8JR
Nciwa7lf66ua13LHAzw/5rgug72+tWLAhr3lQiWPwcBEx0X2toMtk/VUvScNwOkRu4m+VjScSJIt
xhj+EzweVXIUw6+VxQL0OsOAJK+HLGOYQj6fx7cD8P0cnzNu1+2FkKCnUXo83ErNWZSgLmaAcBSk
sKmMjUDSdPO4XdPOJ2Gh9KF5lwQiTT7yVIP8DDkGV5Dl9sYM2B44GGKpiu+k9NSNf88ROIMb0tfS
GnOemlmxg/7aQCsmkoY0u2A3uPELHH2RyDQAqeWu2kKPaVRArydiQS50OvgUjQADKz9z9LSGfQ6+
k/g6cz4l792W3Xl3FRKEmlRFYrVyAP94HqZv5BP2FAveVrLcel4EClqROhteiP5YsF+Dznp+aG1G
BmjYO8DjQy6P7JcqPYh7jz+SykwBRLCJHSMpGyoUwh+D8okxI1JY/OahUqyVam3kbtmCjmPPCc1w
aDCUv8itWqBYRv3gfU1RN03sVSQFnvz8vkrSwm6K1RbglFN8uJelkKs2xQu8OYnKev3n8YWu6bS2
G6eR2E/vMpUDV2ghq2NJkD/JSjHigpkZq9CaPt26Owy7QwK5R4gXfQXBTqhQUKywz1/hZASfrhlY
FQmHtXeeYZs7Kp2xJwjkyvP6C7ShMSkbM2sdaqBHHkENcvCokRw/qLOA7jacIYkmN/Sp4/BwlF8W
Jeq0hKCk+ismS0IY9Lkhdii085NYEP5gS3Gwnt64tfiB2c4Fj12YYsLMZsqs1aNws69hdeLlfjNe
udo1sJOXIlLfM9AkSD6OWa9S6N1UclDqGw14THlWZyx+qtz81W26xGJKOcF9j/T3hgkjBrNShar1
XAkRXJS2DQW4tnuG/y8uMHIKoDWJqic2gljisSRDCTFm4eOPfXogSEvZnSpRHx4tJq8KpALrWL0E
tSYfpBDpIFrXdjg3O9nscgjLAcrYFUdImO9jT2EU8p84pIkKiDpZdbUAg/inWI9+M6Wj7JZtS0GK
TAhqGUsAcmC3OeJOmYEkx9AEsTaPz7/FJCo/wCGUy3H4+73eXdA/QLNVoAQfD7ykqhorg7MXXWRk
z9Oeo9y7bdaBUyLt/R4vb6yAB0ET3N2rlZMkezssIirDiB0EdH/7DFvrqP1pxnmCRFcJPV7nO3RF
WSSEjtF95D/+6iMheVsjvI0OHq8V8Tk/QAIrwOPJl9U7r0HB9vQmilxOoxt56zLe86UeQIGMKlDB
+VyJ4vBltdzI+UG5VSDkVZw5xPPOHLxwFY4K5mjgcRqt+YZ991UUxA8hc7A0bJRhTypN8R6flEhI
sbZkqY25cyhd5iL/0HJu9Qdl624G3Wz8xXj8+b3bF/d7yZyenQotkQZfGsN6MvmpqFFjNvYJlSDI
B0cDT9/bc2lw9cz7bhcKenPYMGUFLDb0ByYrdhgDVdKuixuRc2efLAJTgG2AzE7weAIZr8U4j2i3
xESGW1k5D5XMSK+jbrwNVeNyCa1A1oeIcVrWxE6bKAWKnHkSik3AE8YoBaMpIkc6ChDrcL+xiEiU
jgZzQPdZjFONNq0UAGv5ykz58xkJm6QJ9LmyFRxxkRyDeu31rZ6vDbiSP9eX31LFoHV7TzF1ftnY
N6FzwfDnuUcXGmaLuQqpV4ohW5on7jn27DNnHvJ5kmtutZ03X3SwMr2PoiWK04nOyR09uNkw5Ijy
Z320q8Fvf5G/9S45gLn8nbyi04s59BzQV5ajsXGFk0xzXUId3EniLgsk5uE/EbWSnijJCIIputNq
DxiCcP68tztrKspNQYwCiuVF4ye1i7AkcNvI6H1Cnf+JByPYdd2alqJagbmDWlU07ZJtQHTV8ekg
fvZ6UkMrwVoyhn9ZshFCRh61OM/VZHo6syWg/DAMdrCMmVBb/ZqmbB+cGljcIWglwxHXJgYDhchN
C2EjLz6zwY5I6nIjfO9HP6R9dpw7v4ssNU1QcrgYHVAXiH7Ni3PqWOPsu7Re3Jmo3+WKzv3HQwT/
5bdgln8GHE5UTKyjHjphfGnCYd3hmvIIKKfr0nuLjviXiEustH8TGQJicvWU2yObsV1v/+vRein3
lH8uoU3/bM0w9AiOlN53QrWjGV5y5f4jI8q0gjZCkC4tFIxCcfZKpaU9tnmPGwIuh54hMEgDzju6
TuKbohPRPCEU0JEWKkic380Qr38AeX/qpY4e7aGOfHJ4HJmeiu3F3pzSv3aXyIEnbHtrxRVjkOj6
jxQN4kfvnxsTWR5OTwOP4rK6fxHyEPVVYUnQT/Xxk0pJb89k77lI981PX9eh1UbopzMZoCUhOjZo
GL13ZV4IqrQcAXwBuQmDDqeBoJJOxYqrZTsklT/X3dEdh03POdrf2Mp59cfGhtJLNYDHhud41e7V
spPaOP117q8QtodK+aDt8ZO0199DL/BAS5J0ldjoNads5Of9KBH/PLarLipAwhxDWmZoaU3uaFHW
+INFH8+aCHv1dZQEx94ZHX2TQZi5kGQ4XXRFvJ7jKcj1noK1B0+9fPGaRY33K9rZQzjAj88pnMQQ
sTmStYW1qr3PzUR/pPx+cBiAPE2NPguNzHv36e4GIRuWKm5ORjkxB0gOojhYNHPnVf0YIhw0zi9W
R6pGZp5RDSeLafzbvSXlUD/VKaNCGor+aN8KQjJFPO4K8ufYCebv1UpeQc8QLvhIni9H2QkU6h5f
SlGmpgiq4OG5Hu9sO6Io9xrMNL46rr9ePAuswJ6otfcaGwvKuevoU+1p4+beB65fPZikCrOmaB2k
9pRW6S30gSYU1HMK7dhyDc9yzKVgSwTbemxfpQsG1spux86qTZCOzUrMXHQigRKk8FqxPgGIMDl8
Vvu0AgUGesOw6265ue2L5b4+fexR9DgJEpgq6KmJkla3S/mG8rf/RsUl8sVhzDzdCY1Hcp4VlXMq
EpC+4AfrNI0tAMSnPjfuPVby9fUEsYuyz4KdJQifVJlL+v8JoRcGxsf+2icSTBiJtu2tWAfhEX5u
bo46FBgj3IAZsFhEetnYvI/gsB2rwIQ4fPfFIE/3eLxm0/HSVFf6aXnN0BB0jVCEEpgfIHmPCU1w
Z9HtB/ocPJcBYiFTg0ylJhnoavPrHcmJ845rnbzGgGfauWdX3HXLwCN/dIndzMJhasXtSFtNUOwI
Fmhd3u7wWzUErykV9f7DmZ52eHHR6vFq8zSRNQF2rMh8oOlcyJSIaG1INLL3xVhvgoKTv3FgBKSc
MvvjY34NIMmYT0kFhc5k58hDloVHkeS5nyABHuLYU10oGB15Eo4NOA+82HXytuufL1WPpU/6asav
Typ4//OA1RKNMrVVSuod7y89VgfDCv1CSVaD7v/7X4PMOvakpBnh+CVJrT71Q7YqQiESdttgYz7o
0fEBud1IWhTp/RvhLfuyY4Rrm3Nwm+pruCXuDbxU/9kuvaaXWGs7HTfxLGxsST0OkVk2ftyLuoBE
ZmnJrdUwGvQFyv+KQfzZjC5qJua68+6raxzdwlb1ZYF/kT0cOWH8Vec8zWZ2iFG627uaCstzQV+Q
rIsWgcByRfqGGuppATdoHVHVStxiWg75Y3/G4oE9UM9RnZwjwrMvd/ZEp9ViuNk6n62pKQDLStrZ
o1VxQD3hrolm3SV50AV7QbnKGjMkW3YwHXL+p19xw/tuE/zTIMddJOypGATDISBSkgEir5ueh08V
tNFmKhKzHGNPTbVIKjKC+canTs4XA3k6gVvAFcd7SIhDacbrRRQdOs00mADxs/sQI1E86Sbks1BU
uiEkT3uc9J+FQ6rxE+ALNhmTJheYXcqorglxNG4cCOirgvf3UOfgOmjYNgFioBxs6WqOecVnYve1
cG12aDMUbjNfZyxSHcwbNt7HOV3scY3xvMOtioEGEeDDfPY97AaN3wGGUr6SePKgIgTbe3/2IhbU
YAHS5bFi2SlzyRmlK9KvRnd6on9fU0nWTVUov8PiX+8WY+2+2hPawf4l8YYHT2NfcbyqyQI6A/hu
npHA0zigP9M4YIF96Ael+NHxsVL++QNxY+l/K3QbeYrEglEu7wwPQFZaTHXo4U9Kx/9AOFxnw1EA
1aCL3lUK1IRStdtubW+q6D41VIBsgO9VRXdVeRxZF63ZJyvghT01rVrSNQRfPTEPLI2F2jSYHol8
7N2pCL0RMnOejOUmvklbE9ECusDcgaWNxwMs9sHRXf8zsLttvwAbDDi7A+u/yCBjpXLO9pPe2mRt
PbI22xVtnphXP0HGFnvdSwu1JeNbqwwiLc0zrv9vBoNFnduzp8jIlGiKks3tXn4yRl5xJnD8Hq9f
8m6X63ttzlV+v8WLbN38aQJ63mu5Q0wcfPmrs2+mkGGVyuhBpGqFyPIxdyJ7PqpEk9A80s3CGO8H
zWdKo90sxfss0X+2TtaelFoDCVyefesJp4A21PpLtQLWLRCjJWfgGaiPajbxt6bXrtd6rh7ctFuf
sPFovtMSPxwYoFgNaM0iL1Bst53V9mNmqFQfeHXLwsVlJnc7if80BK2iRfsAPPvQCj35HTcEaekB
i2L6QAXe5hAVg3G3YJdiVZi7yUPOzIR01N47EIld5csZlTQEI/m3l/isEpr3R4jpzSONqHWK48w5
LCGSegaL/rfV8tyV72nOZdc9FF5EgkOztJXfnZOSrJE9n6eM5ftLDIGUXt/8U4jbuWrUkij3Hcvl
fvA+3aBPVDBUKl0SJ+MBWkjBA5mI1aQPte4wuAvfZLyzTXK2p/qOtO9VdVeAB3wxhEwfv2KA+Jvf
zh12tuerhjbOEGo3MDCIjY9q2dVssp5Y+5JCqF6o8shUo8RaMKa8vGZ6ejLPSx6eSzOKAjPZGArb
HXowziGQE4cq7ktkOlWUBhJOAwAXb+GTE2/jJXB0zfrsHC57ZQ6uE0CSWFANjjvXJTdlyK4zDNty
l0mpEBIhrQqACG/+QcBFioiL7uGgSqmMUxWr5Abucsou9KtufV++HT5I/K7vGMpIbk3yKeMlndDS
GpWqYx+2Yl4gUfXTEaHTqXkiuyAC+UZ6wQr+YuCVd3Ir7elTDjKmG9gywa6e8pR8nx0hnBhmpm9W
jNcXn1th7Y8Am4ReAZkK6RXqs3afq84/bmG+4UlvKmZ712MCACS+91eBxqVLvGjfeak3quI0syZt
/HXEgx/5pZYgVuvdQJ/dZL19ggUq6ShAgWILAZY7yzhumKPXoNZpkxy423DSdbubdnwPhpN4TlPP
U0HplJuwRaSmX3qt0pKB/80qKQTe83OTtSJ2XT3mVoHd4kPEWf6zvnVYFL2/pdQ1IuyBuCJtNXia
YWKaDP0KxZCibpfkr2AN0tLvRU/OesRf4iBSCPY/5/gYrT4+2BLnMVC3UfnlUDMTmCGR3b6Ksq4g
HYdtoXYs/it03HW8wqd3l7H6K9ZZzflqiJiwCvRf32BHXYKxnLv3DPNJ6IFjkYJFXB6SXbFaw2oN
zUJr0I0P57H7fnWcGOhO8F22jJpdOd3S+4d2lFTcF4rz09YQiTP40+lkZ1Dvjs9Rvklu/ZWYoDTX
9GNZMVNt2Rc+McOlNky6r/D09QqvhKCOZbzwJtn6Rc4Ka5H1+/0NbfMgtsH2yjfzmqQiYYZ7H3k8
4ptEPdcSXTzotUBdSgBzlIR3iIN7pgJ2fEzF5yt58yIT9KkEdvTUODFYdD4CX7Q4lLoBY8a8i+sX
U+A6CERElFjBJI8mEC61bpejOq26eCK9jfno7BlbLtv1V1RxhwY/LAulpWYzg0DN6+u0d3rwrhoU
v4lr/hTkktuhZsm8nVGuT137E3v73e1A1HfSuRr2LCHr+TrRKHRLKIBLOCSFytboZFgFdrSO7Ojf
iKVSbKfrG0HrvFqN0EDbsUN5ZOCknUnm1ooPdTcZf7cKnTUSMwbK8awO3sWQ7F5NzfudL2QizCsR
WefykSde7JsDfadgUEBpBQm3JQRS8auaoXfsC+Jj4tgOw7eSicP4QbzJlZRFQfvng5WW8nf7PHjP
zANcNJ/wPVTNhHsGTQmIMZOTAo0I3aoZ+BATHf0j8mIgFeIfWi+LDif+H/DzZgnCiGw7MmXTxXyN
gHuOk2FDzLhmBqzuEQPd0bxNMLApu/L0ansOc+GlxFdCAH9U+E7lEVKSwwxmp63ZmRhRyj34898L
d/iba04FI83Zi2SaWi4C2BImfviXBW18X0lmSy9GoKWkkJDkTSYrPDFtGIMAdBsU+/uc09aoEA7Y
uIl+DsPPJootLCuQnqrSrYWRm+lTpSQjkeQBJgQfGGlfu4lMlSUCawwuGJGT8JbgqmSPQFAi/owC
JtYpZMurii2NKU8A7fPWCohZ4PK6orWR9/1H1OR+xIlJrKD2JtOs4zo0NaPlDjJ68h77avyLo5B2
B7Clwsxj8Iy3XP9x/TaOpQgjOgXw+zL6DFLKXF/1ghFAnsI/6TYqvox7eySr5CqHPg7KDi65BOkh
/FLT6Y1PBR/9C6H2wU+C5Qn+wwHCEZNBhTaHis9DXK57av0c+BrAkH87KJ70Nq7EBiqmXLdBHkBs
7xPxGkZqwMlaBWJ6aRucsBPUkLvEjLVbTYqDL27sGAMN/i5yPNAsBvkN0ca8iuCuln+QI20th2Rg
ApYpz49ZpzxBqaQ0Q7jneBaQ35LulxM6GSiY1h4X7GpwFqRU/UWpY098dbrR93Lgnu3aSrtnJ9BT
0c1PQomFhjPp241EK+PI8idOaDknXp6EbAabLNk/fqIPIqlk9ckmNk4ujR9Kl5gaTV6vfKiApX/h
sP8KbF+CVC4IfMcyw9t/M7NQOsBqALJR6btjIiF8u0J8/eKyTXIOPY9GQomJQaU+Pp/f2RJmfKtV
NhrfJ5YEweHsJbhLGkQPGEnXcvUT3OrY4Xm0UcUndusyBvl5ewk3rhm6DKCJ/sCcBsPl/R+wC9r9
BgHwS7Cz8c4KME+R2tymYd7+wK14n3x7XWp2gUAhY6opMJXOJWuItBI6FVhxsR14sxGnELVVVhFf
Z+QFziU5XYEYEcgMogJsp5s+PQeEdYTiOLS2wvt93Ci0gpH+EXfOj9H4eRwoW7DQAzR6cj20FbDi
egqIAd3mSEUI196mKC6m0PzswAUUb+on9UBPqEZheWpVxdscaRvN8LjTw0oQSl4SDjW0QqfqFoKA
UuFEuZ7vYRujgb1HkkhW8g7Bzcshyh00qC2IBCJZG37pwviIenziHQToSSdNZNq3aFkAOFr6WXzj
4IzXI13qXFdapVzesKLyPF/ovyj7bleomUOcWCACmzhQ+4PeMDazXCZv2cImwNwwyVfcswl0LsWT
F7Bg12oXet7uuvgOSXl2Nftu4GFqN2NemwI/wpqRKnBC+XdFTD6I5bPzWEKizssJu5XOhphyVZj9
QrFMeDVq/lQBm8N3KBC//E39+1Z5F0sIwGkZ93dbgiP4lPsnkALxQPgPptJeqHrTPghaCjRruUO+
tmhG4BN3Cr6bjlYzBlSWoWfGTQKvp+ZAdOyFjcV+y9XtGdSujtPnHPKTe71Td+1u5bI2M7wYw1Q2
2nj2ZNZbLyLJW/HDFhQp8wusyIfk5XD4MIAEKqu7A/WShTioegZIh/eMgDWrWPrvX0lCaSWeWp1s
4S53aS3YJ44S+YXQw10PZIzweoRKOZlC/nzu7I/Ramwsk4nH+QjXSpOb8aNlSkFSp7Q8s6qh4bPM
ElCU17s8ox0J5/4xbx2OQqLaaiS/0ogQkRnjP2tkJjCnYd9NI3Try5RJxCUjZoSbkwh/lp8vdTHI
UmxTc6NF8mIX0OrDBtmFWm8oXXf/i309nheM2X7Dty1HuZxptBO11Cl/p/QZ2tWO5zJRkr5mmUPD
YKtgYm8kNiK3XEgSWyxU0jCMu7p7G+MloE/XJ0LX45qVhfGPR3zfd380O0Ajuc/yaWSqyM3jyONS
IPUJz90WIzSrIG9aZ0EBlGCRk3qfeGcr0yZNs9FDwqAtgSMM+qUA4fusZzaZh8xry7G59OSP+/Rb
rMbUa/d2unty/gAbLUcZZsgZ0MRV3cqc7VwjSjeu/vYsUpnxB1bow3fPCYE2ewEAFF632L3Mryim
lxXH9TZkkvMYZ8dDLL0z826CaNixlOtZSabfPWs1sag+kn4k2k4tzxzXNkIKC3iXevnP8DkgwO6O
zdAvoTnZB6iba1PgzpAlzWCzBNdbaMYoR/5M77VnnyBVFX4cBZ8wH+SrY5JTN6Kcn/bWkJSm1j6e
IPdXoRcAaHOZfIq2+CPsquWH35oyHtITynTAiNlVq/9QBz1gyh7BWCJKLMoP4TATfTGBK2x/ygTX
jYaS2+j2KzI+CVXzAHSa22nd+5vX+xz7ZD1aEJXzJX38CxCKskcn38lgYQ2uZQZmtu9L2YbU1NEA
QwOzZ0b2Qbv+NbMYO5dztqIWfLCv1WkAaA76SIFU9zRRc/SS6OIH6ey1npidg8ecSneecOxI8y6D
t113SYcvShWXuqR+XD5C5p2thuttB259xE7iTTXUS+EN9JIqQBuqCy7RsvBTB8lw8918SU1TEyn8
voh3GycYRbxV+CzXMt2pErCJN8rMqfqAtrKqfNABfdRQu90zI5o8n29aftWI04Mpr8T5TjQw4Dgy
yOm/s02e95e8uyGlHAOyO7WPkxzlls9FJU8I631hpjvhhKbjz0LbZkP91onmyOGScgDrXkLTmeQL
vq8CdOb4M2NuyTQeiFx8dgqPtuRurQu+G0kWhQDrjssTJJITMTIF3CGfqSSvla1p3/hpidkPMBbw
PP5FRRrsYzSl8ziz9BQQq1YUCJ8lFA9tu1e77JP5ZvUkpBG1QAKTwjI+52e6WCkcFdTrYLu87Dtc
rdgRjSQQF8ZcTRK8b4BqWm88MvkwrLo9MwDx1lVfeLfrp2UiyPB1hqlYC90cIRRXaCHNTpVXQGic
tk4gK9DwiqHQfZxNq1ciP2LGb9XmpQdiunUDDNs6kz5OoSyryyOdJrgkQAZmeOo84Ad766ZTYFPU
SzJpRkJ+0O3XEik09Kszq4HzAriz9cTBFcuSfDcxjDwnsID+j0QoN7j3+sN34X1DJcw5S+EiDdYZ
Ed/+pcj9/84hvAutOuVVJjEauS+/44B5ZwLpuFt5KqJ5egjoWBBY2ms2E4PudCvLMfEz7G1H3UJE
GDxlKYfuwoevYm6Yec1dmoq44ksn8ceSZKSXkho4zqC/6J60Nw301VOFsmlxJ21DQqBjk78W4r/w
zl42NWzeROpsMmyMRkckx27Fsn/GRWC96hbmq/sfyS60WybPJbUF0Z9BNjcgka1B9dnQ70gW/91w
GO7tx85mPyETVMqzwloO0VnzvMUFU0o5apXiF/16TEXxVuNhWwpp/7KT7NRfWkM/lyQv+wOMJ9AH
rPjgOgSSzctWOKBMRl+Gu/2qSnrIlj8GNYZ9gjaYfHeyf3uxyAvWcJzLak+cDaMpyomhZldw3+6u
CYOfh6FUXmpbV36UGwzta0l7XhZdMt+pcK//EBVtE0iEz7OHeTDv2MO3G6bfpdIF2wflcyA5Hmfz
53Rjb2H+zESv0SwqxFsFPiUSjNlukrhuYX5y1s22xfLfinmCit3kM+OEsV0RAydOsWMGwcLMy1jL
VmQqG7n7FzftquXW7uvnxgBi/V933qtxS/r50B0A4KXIloI8Iw9qtOefW9FLkpWy6yJ2bwrzbKJ5
j/n3R70yL1ug2vHFVKuIYcZ3JZvkRSxLmoXJABaWSCJgfCVQlh9tu2s01ffmvtwbcNXeI47H3AbR
NKZnyFLgLfd9WNpS4mqb9RfQYP50Bd42pBAtZLkuwS+mfGAlg2TqR5q1kx6mIqfFl7hGeREWH2Bi
LE0taA9XOHb+BmrgruCQQkCYwR6LQzxeDfVDA7PjnjFno03CgdrKxf+oWYVMw7EYA9CEeD6XeBV0
XrlwWzwbT73V/fxQvApM55zl4wbo7RWMJr2LNjpZi2hi5+KWEDWSCm0oSENSRh/vWUtXzltcbEJj
1fUNHc05erh3fQYKrTxur2102cxa1Hkw8uc0wGi6XzWtSzrFAqdfK524SCmp4WsYYSG8KogWkip6
vnokbkPftI2OTCXjbOmJk+ur3WaYIPqRMqbbkDdqGRH4J2xj8qSTVUkXwFPN8q9/rbEtUBfMcxI5
0PAvfeZhkWrbK7AmiPBFY+j34feJ2byVF19aJpcZJqc0PtqnougnIv+k7dFA51I4ZFBfgmkz2TQ5
wU+GzOdU+9QX+jgmHkM/+7dAUPszBo7N2vs62SGu2KphGnYzCk4lgDj+vjQ7c+anNzpBeAh9XYL5
oT7WAktYBFYPKEnqytGT5DxXCeUkm8JmMRPgaleqep88YVkGzePFPjsBfiH0iXAFDkLkmdCbXC+F
yU44043SiEWVpbP3JfNcmfvjy9WRpZGiu96CaZMbDHeq8tNke+lr3VDZlppyT9T+OBY+DsEtYuos
g7UPhIjQdKPLv8qbVaYDhsdTwWVCB8HEk2MaAe8t7m1VPhs/CW4WlhDci9VUM1qF1a/KJ14wI2Rx
uvC1gbicnqs+qYzudX9M59hq1vM2SiUcMjeHqCnhtgXrsMB6HK+Wdu6NCDR793Ghs8PsmysEcl15
fl7HHGUKIo/HYENuBswDUneVK9Q48z5C/YAIXfe4S5zWhGms8GJ9Zd+MSyzugJ0DyQU4dx7jyftV
oWSyPvsjAxN4kDQwjT+2sA/mz/anLibG6FiWqXzYqMiza4DgxRtWVEyVKttqWnvvOjDu/EX4iH8a
cyox6b/YGnZ5EbbMT670CaiXh0LrcJxwdgCiDfHN8vJuSjqrtM+1BlsxKCBpJV9j1G3PFYE/Vr5k
BV7/1e5E8VJcJ3mvO/pH+YUrdI9vsyEvVd3exl2slM8erYJzHzE82fJABkUDTl7unAcjfgZiFfnC
GMimz5ChSDPWF8ZaABPtOOvk6eJ6F8nStj5IA5/rVCAXsTfgkWlBi9h2pfDmrpXA8ZN1StuBnEKQ
WD1IwLfG1QjQi2VnTdRon4JpgT7AMQ/Lk855EI4rngkdWZ9w9mrHV3dlLTRpItCcijTvVxdWPxvW
29keR2C72cvParIxAIotgYVT1kfUUICRgkAsRrVQWCL9TBM6iM9NoRDUdYlIzvxqXUi7ll6Ugut1
qUHnD1kwsH/H/4eWkwij1MqGuJ1jW1Ioq7qP+nLa0ZEyIyJvEvrVJ5HF3fiUZrAWuLqv2A8URKsb
vzCba6aZyIuBPS/QQA0mZ0wxOecR4XbvozixPiX15C8shLYImNZj5prf2XgadCYvp+tMhPN8rxka
ZlOvWmN74xsZS4hhaUQZgeqioDcGFPsjB3e8NPSSygVP9YmyeaNuldlouJyTpvvyiAjN3+bH5M/l
hO8TUN8urPmSdua5RThz1tOoKu8p/qUloGGwvrJC2rEFJOuTiuBps7Z59YpYoWIYS/1z+FjeVdmE
RuxBtOIFZQWhrW3f2EbIGt05ziTmayIRSRRk89iOksDuytvtEQsyJ+ZDuTADjlNgY5dUfuMs/bZi
0vTLrxeAr1ZkjVltE659ibtLHDAVN+LRs809jiZAiAgvuIOVfKaatoMpa2LEB9paouXO2CoXc2Lg
uBQ07x/YviyzTItwtjW3TSF46LQ3GkM7f9GWKUaV/Rfma/ksD2tGL4vxeCd8t+ZMfNQFXQMRD8aD
SHW+1vYAQAm/wtiFv6eia0+Bbp3crIDygvHMMtP/cYozctdu0Y4YEVEz5c2PnpvuaI3pfBTvIVje
tGl71rZOmdIt3lGy4PohVMaJ1KY58JZG3YjEZzyQzBJeIwOC4UQb6HPnCO5RkSPuRu4zBFlRtJX0
RyWhf4rHBPu+8yZTCZSlaNUArVMmAOiwXx1fO5Q1cn0ttXSH+NpK60QX1UYnjLrk6cPL6NIHEafa
JAdAm4YbTxz0bLkvw4UGLOBWpRSSrOJUJ9D9udnK4d93cTRyH20JW+Qg04OZKqtQcKxL0KLu5AzR
Bj53Rd0XL575DGHOVVRkHYsgjx3tbSjYN2a+tcJvmPmZJagZ8DxEg0KKdl62+GioIYhQaGijYHl3
MeVUZhUxr155xZbk+miNmGO+rfB3FaYSDRKnKrxoJdwVJuvPeqQU6k0Z64X41iUPPoIY9CFMKqeD
zVK8QyNn3W0WqP4jtN6ahdyr7ISwQqr14yrtl8teVffTdBaEsraCjrpAx5ElsPEdVEy6TyAzB4RU
d9i+me5RJCE9gA06YNlOVhtNP1VaTxnxC0YLabzA4yjq9zFvJfaIQPLX00/D4NRd7IoGUvUmk5W4
GamVycX1Vn1xtDsrq9r+ZUxUS439hIhk4Bw9yiyICfwKtHHoP45mjhySLCStOqWUx+d1dA9q35BB
lFVf4tNJ01fIxYDdxfRYyIVx4PFU3//7t+24cQYSYLMUKhZwb+p3qIEnHXIUlqW0ehrPzncpkzBt
O2lRqjLVlQwq8Q1/m20c3EfffMw6/F+pLtq/2Eivt0hAnSAjpoYX/Lj+7UwQ3e94a7SND2GQr0y1
jGHVwoYjxZJDDHNkAf94dA2OlIc7RU2dMEGY2RBtJ/JgbSnI5n0Osnq45iZGuRnrVt60Uyt3o4So
UvRDsagradlih+nuwOkgaK0TKxV9qGlQesZPfmsWW9bG8JXIcB/Pqt9fMBEM8HVmdgLmaao5JT1u
Do9bjSnjZ87Ey0kwIFU5kWXujaXB+JI2IqYlryZcYQ2AK4zaOB9ryj/D4283XlB+RQ+wIm7gtYEs
xqUm/f6KyiQ+mpr93NqZloHXhg2m5GNBSx4wUL3GNYur+9lJEODOlOdr6OYSwSpdZqNAZPzWO9Ke
+w0OkGxa2UU6P6gXiiEovNgd7ax7wUbwMqEoBuXvb0d962mxz3zdr5fm5VBrpZz3ygTLu5Xx0udM
4FBbfsenlOpdWoRAhPjKc5sdDcTI74Ny8FWYvaIn8T+4AYqEpibMkacvZ61ytVhZdzdnscPIEiMc
5Eaalby8TmGuzmN6su7H8sMs1yu7FblEedF1j2+EgWvSps0NIe0mmuf/yUOqOOcQz8f+jI0X3qpn
4m13Qwky7RmeMnLSB9dWWqqoRHUe14J6npdVOrIoq/Kegyas99sq3toOAZXj0JikLAkizMjaE78p
rlMvczhNI0F6GnDjzKMtBzyiqsZK6haIWs4EsY6aLauOO2a/iF8pzgRvmoEAdMoyXPezCyVsDIkU
fvgzD4DZ8FgqZjDrJS1i9Pov7GVyEVnXAp8OWKM1k2hwTKzCTmOacu9p99Z0x2YDIqmjOx/Q7kPv
l/9PXDneK43mwrU9ItJ0kIAV5ifn0zR0JxXPFaQ0oZxMVzAl6f3gqeQ7I0sImiyG6PA8KP+yaICU
ZUo4nN7vAE5+CPA3gUR+8Rqm17rPHNub8PnAkr4iM84wL/JzOXw7+jT+1WplovRHcZtRhUfTi0QH
1CwOKonZRyiF7sILxJ3QwscF9ctu4EauyJ316BMIZn9wFBTmBtxAjJot3DRB5yWiyYCVEwZjwzS8
UPpEvODvNOj4vqx5uOo5cCXTCkvp7ajS4fu+GVQLUNGLKuLaTZdlebkLGL3KaLSWD+ShH70H71mA
yk+WlSVx4/g/XzrIjGXnZUSkdETqj4muCZHEFAvn700XA/or+LjQ+4ta2CGHV/2YqjdsGyFFleqo
3PFJ8/QdxvjDMkjFp/pZDvKBUi1qXXYHJFmSyegDRIEjxUgCgECI6B6xnZm5jvNYNF/TEnptJ8BE
SRdwOvGxTVnp3kZMx/3pYsdWa+MvAJhH4yfAJJJ9JduQr0Q/zjob2TBAbFed5voXxL0LDVMrmUzw
+STHA0wFPgoR+G9zk6KspPnAkntQBKOuvTftBTcDWCLRg7io9SV04HK1CjmGPyJ2voaR0ThtMlf4
m3ux0P07KXmD5kkMI/9oIebsJxlh6Zp50ljaajWwXX+ZR+tQqxFYDEwJ0gXic4AzeiC8XIWc3mGn
bzw9gcJ2ipnWwzM3f8m4XYO5LaOcqmM7auDGZ030fIrTmHJwnzH76fTNiWf18CGSwGzEjHuWktpG
FiX4jHXXO9cEKvC0VaPFLaI/Re/4W39vTj1LJZTJEAo8eXpDi3qkoDZcaUTNWlzOkDFQa8GEL9Az
2OXX6mnYawcWL//ADULj0IEohOAQzs4FvEGQeXRCAv79q0JqOPveR5MAkguE3JUpNHqTQT+Nrwwc
IEtGFNtvT5gHEY/LA86WMe3De59Gfe2gq1lp2TtXGrEQUpgthffgLkQZCXuHvD7bBqCIVDHnTRLs
k5qY7f6u+Cde5v+/lnJg/jzxPHDZXIScyTkns1OLIH08ynmBiu2oF2m90BlYn/LYx3MjTi61ttSI
HNqENUTBXbb1Zu77uHSWXU7pqp2rd7lWJ573qXcDjURAq46WT/5kItltCdSniYgC5tNDPvbGy6Yx
B9G5bJOoIVbLnTkPYclPm7mu4TKujKQ1PUzpOJMNjh4pMOAf5d6ArzeMPqSrDQS6UrSO+TXgipK/
TqH5vhtKMT84TyA1vo5LEyl5/M8N/o6wPM9RgveuiHPgfYFH71JkXwSvL3OjiCvVbbre4nsn1EU9
tj8+Nch1+6Q/1Z0lVIgc0S9xfimp1a+apUa2fWAmg0ZEkaVrwTv8lFEnRYybYHpiQyiUzM08DtZF
4vS7s9Uiae02Up65wZ9rsWsIWfk9Xmf/wEcwerDKDsIrH1KNeVxbKJl0EvP9pCqwkK++63iubu58
nkEWK92RKD+zqbpguceHViXTUdyGg64rUgzUWRJ035FOnP8MhD9Lapx2Ygc4J2+xnLiH7WZwy41n
lmVKLIqfar07CzGEUNnkSkeacAM7DANkuYur9MMVfWm+/tNv/WLUJKw3IKOsVSs5X/Q7zVnssTZH
cB0subyEAp1t5HsSLNGRhrchSDFnqfK22XLNgw6CKFGc5zYRE4E7jVu+csWW64SiJ+fhphwZHkpr
Tpfo9F+77SsC+3vUaZOCR9/DFi/wl98BU7aDe1HsRck0IqQCzsJXF4+/UYXYHIsC4vstWEI5zVf0
rXBZ7ayDrburnhClR/P4VZPB+DdsRsERyuH/I4KFikYXztzDFUShTxf5RXYpUe7VJ+kIc8le9R4s
CwaqSVP/9nniUtiYotPp06foFrNa4DdKHPA2ULVVbht2xn2Ywx+lJr8k6Xh39r8McRLDyj4hjZ57
9+JBPG6+Dy1Zbhw9xGYl7H1dHZPx+wKn+1pfQtBHcsoVsm7kxHNunowkElrJmxIa91hFi44Lsqum
iWXoAJXWGRTJRq2lltqNmGNTi5thkRckcBouzVX8/vbo4eMujJ0rcEqs+en/xVGUk/NLqEyJB2RT
0SNT4sFQxpPt/QZXv3gAulGsVlNNoQlUPOuwtjYemKBQFbANcmZz5fAWp0sLZyysRT0yJv8eAYkk
fusOn+Xg8Cv3GADMI27l4IlEt9kS83X8mKPHEPACXZe077y7HIVnyQtQXKss/rU5LE2+sFBvBRu1
vKr6dSbDESAm+aLbna0XvMMpm0p8WSq0BzgcFGBa2jht+BsniThOWB29J9LuAVOgc4Yy6cH2/4ep
AOxvAhfJyH0E6HaSbGcF7YJeUHwnKNrc5mnfBhD4Vt00uxpBbJY4WsOm1jvIWip2EEHwpTGKHrYF
Fjq3eiCq93uH+YtwLvAzULi4ZNKFFYZDhYUPdPHafnvt851rb1m6DGeg4iG9rpa8zksd9YBaREA0
hmrObhvJYto7K3/C10s2lca6Gr9npsLb8a7PyD7vTZmjgUszFXbOqDwHJ2ELVoFHrQUijVw9lGcO
dLjkcHZWHVTSeg2oBxS7Zw2M5KsyNdr+EGYcMIuy5PBtBeQpaJ24t1x0Ipz0Hj8qHsgGylLmXlEo
e+IEqhXaYbgM/AiyD0s7Ghr+FgE04xCfnlmeNAjTnFnrW1fCLM+ONkhGKtnz0jYmR4oi3TUQEE9S
2R1bowyAjrVcOArSrsGMJMT4FBV7bPqcCwaJH4LAcMFTMRIkchU+qMBnCCKps6RnHIeHGeFyFgjY
ypJUcnagSOrJI7WILImS0QS1OgIiT7f+1To7d8EPzy55/FSbidrCsDQNcZg8JdgC7ygaN9jwpGXa
4hW4oIeseja7hlR8f7s6OwQwFPVNmjul8ILX1Od9lGtEEgSvuC2VUwpJ1tjzIGnfArVWGqm2fEEt
b5/in8xsbJDtk+kO19Tk6FggpgvV9Wt5K9UxxYH8ccDC4emkuStRJ+TDqzVFyGBNEoefjFYItb9S
++mQKvgeRr4vG/7Lb0XCCt4669WyihhlUcG+dI06PjgvtEaOgYNeLzjNMTxjS08GGsJk8RjFgGBT
efrzyEfn0F8RRGKxZGOpTy+A25wWqrX/Wlw8l30JloSGSG+8P9Kl8O7Gxe4SrNsSj2ArpIc3ri8u
Wc3+NMXy26Pr5iL7z+7hDGKeph26mrBppyHQS7NvcGne7VFcRH9326sDADeJYS8R4JWje/N9BNMl
0EIQSxxVgYiwii9lfgwgeItfgB5vT0YmxDshAGysc/RWMs/q5NELLrcDeJlw+HPyc8FM5qCiDJOu
+iCAA3SyykZGkSc/6nS+MXE6pU9/2VgaAeyba8soRRAGOqW+sjDFRYJ7utulZxdAE5osXVS+Us2/
RP+b3DqDdEAfD3QWGW6Vp0EH4pLncuwY4ONSTJNHL0PauTjAW+K2Zcppdf5/LUErm6g2XYIt2xgt
muo7ZDLp4NKvBnZqOlTvKOuTpDnoBmA9NPQqUjVvNS6823KgwlFBvU7raMNSWNkCsg9SMUg2QU86
9xf6caU0u2ptOq2iv12tRP+55OsNUfoFH+JuhEHNF2L6slb453khkBv4BjdQrG8hHSLYEhrxL9N1
8YEC1fGIf68PfQhOZcF9l/fJM0Ih/SRY0GzYKdhE/1QkVq5HsoCU/0tn8IN/3E0D7NPz6xPgUbUA
WGPkDTcYYgfDkbv5K2/xTjhmRko1XOBApu3TrdPii0VthNamLlhAoBUn9zsPvDyH7JFqeXjOdcew
Cp8vOFcZjwGNk8/Duhb7zstx+R3yDVGG4Z7j5qVZ74e91bjXp4nMvLrFT7fOQT/Bg1krh36Rq/hN
aQYG5/ewj98pUBKk5XmLmTW7bIvdxmIitm7jkyAc6ICF3jkjgqbzGdX9Fj1x2au/5KceLGf2ruzA
+Yj2srPBkoJMsoya7QFGHR26yFQPBzL922ZVCCE9478UbS4+xB9q9essKhhxFHeUNH+7RbHsiQrm
REPBA+I9FoNOQOmZM01xnh2YVk7AfYqQcE29A2V/J8+mKQn9Ovcp7Fm9LHOemIoLOGmjDNKr9WXx
zUq1SGUMXzrPxO4PccrNgPcl7QLcQCGPUtuarEIj3DU5PtWhg2yPnIH4JRC8GUV4b6yW5HC1RZg5
OeczIUopJrDa8ft64SPzIsB2LBEmsovlV1fNtosnChOIWQB2rXUdiVfTObMA7czgbTTZtEsNEsxI
t6jK6ehvF+Zze5kaTPXtwZEyVqCM8jkBBVHR7OcV7lC5dUhVN4K7fENpNCxZS6lVn6/aWOnbfSdj
hoRlBzSTDYF8O/zXPnm5viC6lNJ2278bXmV0nhjyzFDvcJBaqYIA4+oO4gb4MMaJAIQcocSdra0w
HzBuxq3FvlgZyxnQkT9xEFYN1ruapQ3bg9Cs/z7BIp4+tClrE+IvPgRORIqftfP/+JXNMMZCxhyS
UVDandFgbaEVdZofOIuGmfu/AaG6vi5basY92QpGXsbJF4nOtKg0D47bxbreChfHwuIZYdD5mMUe
eWOxj53u9WIwU0bIuVG7X0qB6modYC04DyTKLNOjGHqxVYneUEpBbsJNl19ZQA4DOHHz6sZNXP8F
G5rOlJh0xY01Imu5w9LXXt4Oc9YeKxFoQiGzVWTgicJekOEfu4westuo7PIfBvUk643MuXlQ5jqp
Cd0y7ApdOMPfKPaZW2ekaLGCdSPnhAhf9OxPqYxPOq8b+RyrPT8AOEHkHVQMB6TW0hLKizfn9lll
f0aE394Zrv8AM1wqvtCEXHXFn/iwGR1bbDlg4ZFlcNbmL6/9zD12RrX5eDlTAabN5vI3rJMtYMNF
9jD9wAJLfHOdFdyrdHLBhu0snMSrImnveS/S9XBPVWWpdJcCybJ+LFFByND+9JXZp2Rrp+OGeNs9
MFMY/wXXbTuWYzQ8MabUGyA6lQlrZ57+wqqcVY2jlKgQXR19EfNx7k2ORnZJnPBQQgstLdE2C70d
HaT8J7Ey3dKIV3JFd8k7BwCt6m4WpFfOyL2hRfETqEDEsnTw8J7ifSJpOSXJFp0bqthAkPFgJxXt
Y9zoMTvXl07n01+4u6qJ9iCfDnbH9YPUX/LGbOd9nMf50FHPYGqy51rhgWFFHzh2MDMhbhuRs3T1
vrW3VhI60vg7RTsfEBMHwcOn6Iaa8DyOdWwi3gWpwU7qc5+up5xTVy5EayQdOvAHJOjmf+zwEWXR
albk7ZrOpm8a49NRvdkLqQiGTaEwWJY8FQsxafsOM1cHy25nfSVhNqbAabr5ww1Kt4maSavP9Egi
K/1oegtvf9iBaST2ajHoNQaWCf7pAMKKg/zTNR8qjEJyNsLU2uzuh2VbH7wC3VFzHRm9sr9O6B9W
eRueCys6uxbsZiptR6QMz3ZGYyBoFys41OoZ3gTIC7VR7JZbGOY44v3EOI8D2BbBf/qKMVA2No1x
vPzXIht7h5dOZZXkC5zKJ7XMpr4YwLo7zjYP5OHfVxV5HHuZbeTlZyEveUpfAQUDxLTLE5w+2csz
JucLfYYsrH0OMqBb6qd1cD88OeMqp0NtJRd3BwEAA5qLs3IC8QxYZPmEP/nl/zwGx046hR9RQVL8
KknweH2ogzzOiiq2xSwmGepoEbJLq1gZVE/3uQqiSR50VtTCjVsiQ013ED4LvTIozxijAV4Om5Ka
T+A0obA8yD3giLB/HDa8ykZU14gcgLJNQHO5xB/xu+tbuAifYyWT1P3PiCZAD0LTHFIRlDeHF6PD
ZcUsgpZuJIX/jb4yXXdkmPHm2bMt5LxcjRgpmmryl1M2AXzfnStUu3hXMcHIuOiMm+3FkIpDNOxD
Y/J51xgllphjwC7CiTegg4HKMgnnk/1APp+jpUXic9JvoodaHls01id0iXkVK9c48Lt71HDyiY64
hPt3Uh29ZE1O76Pw7f4DkIKlLg4jVU9FYvNzJWoVS/tssiq4dN9km4shZ/kQ3e2kfqxUDEuh+xCU
dLKRRYX6uf19udNbOBHlGEUksYR/R1BpHZZtDz6M3QW+rFMl1RXbsT1eEZs0/AMHD1P7mpC0F1f2
Qtt8ugNFz2srQoVdW1iz/0t4PAv7P9DydfaTYEykOf873CXSERzu2TDkQbSOxqSlHOd3NWipF7rg
qmMbdJ8tQ/WzKF+XjO69KXKk3iXXkidLQCTEa3YTy9BUHImEptfRAcoFkBEVio6HJScV+wRiXI2W
cl+iLIuVLx0Wg2epo7tWsqncbwGpQad01o3zlUIo1wwCivg0bm0lZQ+TII1A25Bdg9/WPd14HtBU
2Yb85W30ugaA1cN5KKFddQ58u7PRDW+xfySZljVY7m2CGJFbUNjErR8rWEbuSrFMCf8kX1loXECf
WXbPHQTWwSHYQzRAqbRZtQN/MzOSa8Mk/wKA3WEwN+BkML+Pk0IY7h7sDdhZUOmfQMK3lDd73eZa
1486Z1tvXnMbrNz0wnyTLi8TdT6aLUW90C9V1h64qn5elrW8k0pv803mbyJc00HiWdPh4Zvg6qeq
u233vximJnP1Ox4peXweXrdIoc8ikfE8HJE1XyJfaa4JmzS7zvEeHyAuhSKMBGISToytBQbkYYRY
p32WivqlwPplt1Kn1FDOEzEmvD8lrik0qTETEm5veaXpTmhlZn9cNx3Upk+4x0hYtFaN86+erSyD
2yas5fcDuK0Y9yrQKnNT/BFYE9+Yz/gZEOjO0vAcQiLDMvs5hGKwsLBMAk+S6ihitwbvks+jlmiS
RSwp9iH5hWKi1bi1Yjvryl+yL0RB2KwLG1+JlfRED9EggWJTOTE3tS7H9xEjgIS6YssOnBRHJNcx
1al5pY2/piCZ3J9LRDm+CZyY3ob+n4A0RlGtdFgUIDHWOM6x7irfi7zU936PTgussXA1pKBnJ+6t
S6H8aVzXc3AkhTYS+AITV6GPEWRGt9MH86gEsV2FI1O0JSsK6Dbwwn5TKHVZVJDMrEzlO7viEtBr
A6xOKqDQLVkqZIRcnCPa0vsTWWz/RakwZ2Y+7q/AQZiyeErtjYio1DczCJ9rUv0xH2xAPBcm9tpG
WmKKxZV8ArsBVjgiRm551WT0j9OwyUxnfvedd4STsdDUjTJxJQ4a+ZwoQDrG4YIDpvdvAQnt7fzC
pebq64dh9MC1GLT9b1yFl8tHexwwuYlWFkliebKIvRO+mt+i8ePGAbAM3tz3fOKDxbAGbqv6Mlkz
MQ9W02QiU9hDFRh9YRvd6CREaOoKN7/I6Vcbp/+r/wa0SHT7ZlrjdwHnoVnE16DZatx9x2O+Qs/f
gSB8Yy3jd3j+0aQg/IgjTGnqLoIFWt6iGlN3VwmJ3FCCdhun3o4DEGxH3Fpq+eG9YQLAFGMFI0f1
lPu7al8gGgHCOY1orfEAGSu25poHQanD6nBzuC84+5oyrHCh7kSGMaz1P1PUl7v5/rNXaw3NN6ho
5HXgULPTI/7z57AVVPabNNMbKWTErqsuWNUUAED9kL98b0h/vl7F0oL6pVpYAzfgmZjAM63YdPtN
XhkHTh6fzdgqORBuK7x+3zSSAo1QKEQzfT9VGxoBHzOC9qWtnp0Cl1JMIJl1AUvgE8HAy9EcYio9
iltBdb67fbMg3vQW+p58uv7lrFj1YOtKGnv+9CmupjHB0xwG21pyf93g+ghh0ncWw73L90pXHPpR
+ggdSaxblAol48jKX1jDaamoVeP+imF6s2EMrGW6luN3neTrGJEPcp4dCNgB6aQDUaiZgslhHnof
CbbRiV+RNUU8sO85HBYkz2lowBJek+1xZjXChTIb+i1uozPYdEgZYMi0yIMUwT2hxCVTMMO0DVY5
UFSwR7/Z2+sk76FbHMeLb812sT7VCvzLl+ifc9KNo5qJB8o8MuFLBJJmntot0w0zyfZMRaLxtpMF
9mWMjQW84deacnqXChqmqmE2JwyV5jnT+OZMMtFeIUzh5v2H/TlStURP9vI4KsFiYevLgLuZQUnX
6SSyGPoZhY8XGhzdvNZMm4ltcXf2sdfBk1bYxnAOTYxNsM7sQ0rKgRdPWzZM3KpJVZGN4rZKCSdm
WEOhqo/CsOvNDO/96Shs9A+JAKxXCx7+6jaUPtk0H6MlqBU0Fkzr4J4c4oUKjAvt+G6VAAiaTBOu
6WOHoRXX5XANjAjvymdatGQYBH651xjof5PXh8WJyFlALf+oat+5EsI2hWxNqx9XztMdB48aci3N
9QxsYk+2Nm51uAkVZu/FrBdLuvMv96UtbsuGcBiASDDoYHdwoPQu3koHRvZIuwd8pwvMramtCNR6
J08cEyjN9vfA6jCzywMRi+N7wHAiEgGnMtHRE5LhytYayczl1oTj7/fPAwdjPU3s2a3GSUwjgOMX
8+O/yDr5dwefEhe3KX0jbvcOqP2jQqi5rNy/Pub0mZ2dEWTKnBn3FxRDQpf5cwsbVmkElPwTbcJ8
HNHi3ZbVn6ytMHQNzq7+I8DEChobALmLNEmutRB9PBbu3oNT/PmvD2bSqgqhrwKa4mw4LuIqaNNL
H27X1F7kndiafTrw38DC14AghXlU5HHuMNPXYs4rzufvoaSriq9RiWS83fZXFaFPMU5krOyf8TnC
ZJWuh7u73nkhdTBKCMlHglNDtIdRpibCm+cgiaRW0MYa7m9pFaxkkwAoishlphDyaUDS7hoHIn0g
1r3f3KIy4xlHNVy4ekd0XERdDvbrIhci8xEhYl+Z1iZF2NjVlqZkLVYGYY0KRU7AhhBZiCMU+2lA
JI5z8Xb84A0GhJ9BqsiAEOav6c6RB7+JIrk+qDfA+sVoni3nAHc9IlYzDkpi+/dZSt8QahCSiJJa
tHwyCpZ8JcMLNJBeh8VjbekGBK3UEPqTD1hMx8r+QgvBHdr1wtp4LVdgBOOP5GVL8N1XvmBBbvKX
aZlZtWmhU6T1OhcFY4TY0UvnmuH8E0EG3NLzJaKa4eaNBZf8hGa4FBf7Xi7Tj/hklW/ZQT0JkaMS
ibpKbWEP6jkhCyy8SzTean8VS9sWsOWPdfg8rWNKqpRbiJAuy1qeLpOfvpHYThpmont18iciZGUB
lIFml84ApqkNNMct+IXjuw1eHTSR5IyUZPJaC1tcroxEIdUV/suJqVgDMv+JV0h6ozyEIkljQHgC
dqVqt8zbhzjlH9bnsQCvrojI3kQtWd1eUF3mNr0z5iu3Zkm7IH3oTWYlQ7Pwe2GmpJNx1LnSVyCj
dHx7hR+zZf7pbk9ZdZaxrbABnedT6/KP121aRlpzLezBZxL3RkhBwX6AbGngs/UkL+vZcnvsZbTV
hOuQnPXIpWKf5nr6Fy6WUjWc4F5xrSfOBlH9666EMXR2GTbyCg/0fkB7P5tmMZkepL5wXuY6JlGZ
zSrDvORxEWcvg5m1L0WYTzZOPKunUrZQfc9TDGyL4bWfDTM+DizHIJdWTGE3ywcaNeIG99BXyETO
a50UAWMrccSRTjeHVt0kYBbQ5ameB//lHpxjGWGouOeIrMKB7tHP5qDRqQykipEsZd2CdHTPSxVI
Ad7RFQ+91BMQtCvj8BCsFtHVQTNsHENOWcAOS9sekVys/1Czxf0Zx/dGiCqTSk+WolJfFBts4AGy
lR9K2cg3zccelQm+5P2+PD6/Uxj+os/D3s7up5auXN6MiDZ0VWySE2ycWzfAQpSaArloe+vJ/dug
1iATpfzUOfPXFgjaTtM0l24we7mqYzcy88x5DZmgJwlunLx/CRo72PMa9f0IdybsviKlecoxgrW4
0JNe2m+lKvdpYESXbfpyqR6htn73Z6PDRJNRqVyjdSDrqXW07jKgvytDKLIu4RsBFap01PRwbgfK
zRdgv8pJ7pE07PyrXPNmcDXbCsnjxm792Lqc/YKebclOXxDWfBOhtB49aNdhnyVhIrU+pn0sN+yy
h1hZzXCdhwkmUDHfDt6g971hiyXpWM/rHr4u0PZHW5A8YT6sqAb3HSCq7bpZ9h1C28zG+x9r7kvJ
03zr90qnkC4W7UZfwaDCRiU66JVhI3br0CEdtg8SkfIpwKQQ5NIyo4vhdyYG/NYHEfyH8wCPvrQ9
0BtCcfGSJDmdwNw7BnR9DNrPNga5Ft46qgoOWyfnq4feGwOFHK6+pPBrAtFF6BCDr8/lvRXOgvgq
aP8Y8jguaHJ9TlNJaKzpUBXaO0zKlkcrnkgUpiL/RxeefrKapJiylaseGg5MN2n3G/XXYTylB9wp
bwksxmq7CmddLeNjIEwTitZsyxIyeRE6MqDWnbix0MWW9JkDt0w11ES1/2EYUxnfDJHtGt2Ns8Wu
lxgxOpMnl9U9H5Y9yz4d0HD1Vyp3OB21uj8zKDq726o2DtxEtWaCuYSQ3+WJxjhOsimFiOpeVKTk
kixX6RbIBXCQKaMsrGMitdiLdcEDEGQKVAjMc4w1nZdo/5rDUJG3sckSWjUhqiGqDIY+NCsPTB63
soZwxaYNQankeR6ZRBtcpkyO6N5V0Wf81Ngu5MkyPmCKCmE3eZfsw9Wd4syz4LHzJ2dn0lw0YORG
eOdKxe/5VsVt1SfXGXBGmBOqTcLZw0jkarWzbd6eGNdm+9JO/VmpOjYwq6P61lX7dZV9Fvrv/clO
0Z8YPeJYT+sexQub0AVadQaD1kkRIeXCG7HLT1aCte+r4MbRUhwiQTS4bBRyvTLuiRV72Uv1y/sU
5ww7FVouPULJMOvO0j0buGPHZ3NgFW9DlllBAuXXz7KFAQ193Pr5HawJQVfRk8CLPeW0M5lsqTLu
Gi+8C0JInuNGd/u8fKzqwLLghsjflNGhmhwdk/pUpWVyAJjHg7tCZoZk5eFKGoB7BVBnKCVhF/tR
diowwcK2pO+eiXBcaHBb8sPsbCRff6knBuJtMhX72T1bwYt8v29JRXyxPB1U9z87blqcuTnVrunU
aetUSHUCRzXp1j9zM/Z4Pi4AEywJ3fGFw1DYRTHGYFfxksr7YS96AQEyxd6RCOOV2W5yyQW64vD5
litK2P7Gj/W/GTDvjRDAW4wF2M442lsEvHfVedhTtAIAd6wFciItLflfYTjz+vy1x27D3+cZDlEl
moXSRxxSb+K+hl/RIHQLBUg3Ffd8+rt6dTK+iItbLxVoZL0Drb8QL5XdCBpNrXxshwJz6EnR/sg9
CyOIvHBl2xQXf2usg5Sq0bKn+2laJUuHtYiz4a4UayEGSXE+O20XP+pi3fqyiP6H/ntm1kWS2IWW
FyGJTsb/3/rpNdq/XsJifqP/wyeRmKAZt4qC7eK3GGCuolv5cY/nJadTNSEM2hC5UhBy55GE474t
eNPJB5KxHTx3ojjPZY5Ar5FOIJtwUP5L6+tDC7lY5IQ4JKL4KmqzlMRfTN9hR6S/BEDavPtnEPdL
8MGMjAChy3SxqvnT/4DbHaQT3xfHBZ4muPpXz9gii0enzOY/S8pKQvJWMtMxExKMKwAZ9Ieyl0e6
uS485YYB0ZcXk0Dh129IZKKbLUNuVS4SKHlb/ZFBFkmGJ/KqoqPYIkGao5LN7HJlnRwrl3v7QGJc
vBOtL7I4Z28vGZS7VOI9HUy3cRW1V8+8XI/Pldoz8QOjsOpWzVlGRY0IBxiSWJWSRkmKcDRtcFwB
eL+U08VTUb4Qse6xVLdymkKOOG5BWXQ5CuNfFmLpaoF4VEi5KPwl+8lQJySoSQ9BdzqRejZpeAQO
kjAWvyAs3VGfxvIWrpO94DmIpmOKCC4Qzg5fpVZ5nRtPzmAkFTU0IsEusBOHbl5zVI6wrgIYYFjn
pCucBNvQ8hTGrlIKb9NyMMtDg6/FZJH7W462G//7hg0ESbE6I1gyYZJKwfmVh6BwIX/55h0lFfRW
oP6KEtoivEbIu1yRhR/Gqqzs5x6UzLWDDubDYao+pYheDSY1O+13gnsOEAAX3sL/bLLVE57jhbhl
/w8biRFY+Frq+2sH3EktRtrn9hdFZvzV2ua7ybTrUD7H65EXhs+dlogbhEV76LCi6ohiN8IYE8rG
WZLIds2OT+o87I28Ebu789liRRYDNjLoGiMLZ0Dumvka1/pQpfxJomG600CVD4TIWM31FufgRhSu
ubulLq3ux0hjWwbhUpL98M/gtMhpIemgBcE3U1b53iYXFKkGXf2FqO4mL3myx4EZT/TonWirmUB4
X+aSB6rMu+CYDF+tcOD3LfBlUFE9C9E9XUF65fQmAErJyby+3KAhdF13QjtUY/ClAiN7fVSj7k/B
s4/wOjtMgQLHGVt5zrsmbn6dM37HwKKXWd26oGNA9/ioCX1PMH8hGUuX10o5r2ZnXHibiIrChV1F
etJlF5DAfaQNHXXvjP5KOGMba0YZ8wRdm4mH8XQ3kPWumL5W7EXClLe3fWknvmyx4/D8TRX9+LL3
/+KZ8fh89J/YEC+Kvsh9bY+nn5AGo4ER4sVf6PdY75K/97ivwgyoDvbsPAUixuKdmeUMrdAEq8yv
o5jyV6HScOeu+L6Phc9OVJvks7iLseWNLgveFsK+AtUv41WuZfslMmSIXXItBLn4Ez0aK8ijeuYQ
nsQ07ifSedKVYk/ATtu8VF9WG9c2i04fYOlSKOKuIVOhG0lcS3qoFdFMlvgpKJG+seEhmEzcR5Zg
ZrYwHX0SJAUm6M9q2sQw/xsmm/ro0li+PB2c6/6dSOUvT/NKGv+/BecKkkJO9q2bY0M3d0vVk+ve
NH0dGeF6Q+JuaVph++lijOxICMnuQlGZchmX70/FhsAOwSbEU3qiEWDf4qD43ZXCTrV3dLAxero8
OyYD0ywZlsS8cS4KwnzXXrsbZH9NnqdVSjCnq/9LZMfUjxz5MAdJEhY33pnzPJJBNw/MIdOxW9P7
gVchORSZE3TMACrJDWDBC/+74dcwUImahnavELydDFnrBu4gS+nA7Z90dzb65Gx/85GMK8OSI7EJ
NImxmKZ72w5te/wsihg3zGqiOBRuIAm9xWng0+Ewfgvc/fLs9l9DJqQrhl4cr67qtu89lIRj+HDi
DGDLeipEec+z7SNzQ0ZWEdNykCa13cDCR6/bkgrgufe/L4d5km9dtP0oSITva2QHaDOZqqhw9R/J
rc0s6fUaFOyjHsY+3qEOqdAxPVcilGgDdO30TX32c/DzLdU7ja8lPmZeXCih9G3SR/wZWQJhCcxy
ZQ7sKlmiYJ3K9H3I+i3Qzg/UUq3NwIOhFyqhEl+9ddKhnb/EqcGc6s2BcAsun077H86dvNhbqZFA
Iw2fcpIgHrehJ5OI59LPMeGbV9q3UWzolRAURDcocX/ydv7mSN7w9HqfucuSF6BmXjWmXLFxDtw5
2gsenUTyv7DEZgxJO8mIDzPCgSQeul2SctyKuP+HZxBDJ0hwbUqRXAUL5oGY8Z9vhTcQFH0R2ZEr
qhGQumOHeMSHm/XdBCByWjw248olCFaf5aSKaag7+mwFoNOOR7TEQCOxZo9nWFINKPtRbamKrEEc
eqtJm3lT1EQS8ZSmRHx6lt1qQifilvbwaePBG0u5RlW8P0315muWFG5CTxIJL8J5DFo8DOsJ5iaW
vMeIzEaw69ovuPMI5ECMdvxBUzX3lN/P8qcDso9svCSRzVeIdTOOIjUEazUZjv3j1kAnzweEvZtT
cR66j/Dbn9RL/jeBaxTigRjfKpeVGAenI6HYLJr1BDo4xjNKw0ZQ4a8txA10f9LT+d9daIovo/7O
cZooKN850en5ni+AkKukwwjcvrzrGqEtlY+RS6L6IWKg87GeV/UBX/wIi2Y6QBE0Cpbbskx4IGV9
5IRNBd2PWLxPCBs3eAnOVL6rzJkcQJdr/fqaHtdQhnLOVlp47pYx6EtwkFLOSeGjd3aPRZLspii3
icUKGYsISfOxEhuT5vlwFOWEk2vIs6L0t/Wmu+OYgP5tlUxb/EGyr82ZejKX8TJIYEMBP0D8q7Pv
ozr6ulrABHxsDkkZeMNgGJS1IDLAyGrsUv9Ewh6gdyIbL3PJ5+EtV910IizGEHbjtv9znlXR38d6
CYHjAUj/Euh/42tLGgb89Th0NU4xoLvtcFGQ/EtgvNG6hjrww8zE99tQfrRnln9TopVJQX6/wK4a
l1Ik94LpKQBjaGaEVEaMl3EwYlK/WweiSNo3Ll08Q4fOCUBdEXb9zbA8lC75rKelMlGYlCWMaOxs
P7HIG3iz2iAjEaURZoFpJO1/bODd1/Cnm2Telcj5SRhqeTQFOD8e/6t9BqgUypwIDkb42ccD94VJ
UBXXjqaT+6FQa/2UuNUP0cn1nTHVyHlkTjXV1NrKTUbC4naET2ZzW/resgpYITWJA3zVqYa4OTe3
yPf1Tb2rJ3LI3qi3PGlF8y7r8VFd1d2Zo/XrJgiVW3C//vwO761UDt22Py3UTraUuesCLioma10A
npsYAY2U046Vzn5frKLGcnRc5r+MMr/QVpCX8hiIz1QqLZyDDr2OR+07JwUXJzuBL/vfU5D3NSPW
IRqQk/oChJ4R5eC7251Fr8QLZDppbfTSlhNOWif3aQHV7z/LzL/10h1ZjOnUym2FzuBz7KtiXNyd
SNO1fb/Sgy2wETFLyufIqwtSflqss0X2VKH2nAb7YP5NLZG8evttZP8hlsX/N4DjUepBTX7/b2hr
kEEnl0sfqMNVE/qCWjX1STeeqiW45s9eKYUL1tdS7hiaWDxHYrXX4/B5hRG8yNDVSZWN26LVWbkg
8E4RcpYVcQrn5wipSU1DKkzrPbo/szVZTGpqiy6RJL23ch6XUiIfCE4r0+DZlRPH7OSLKQfcHsh/
MPKLNm6iGqJgyu5JcuCFgD0JfBNyIWSdGApa8jvMH8ArAHqb2ax57ySMH65ZX0VXeUfO/m8YClIx
IurTKFasztYUeyNbpmMr7P+g1WHtM6hOJjXe6wTcXiuuIZYnj9JDRCqaowlHUFf8yRmTTu50JiVL
2QzQiakMEkvpuKC+6yU5OEh/EcA4B2Uov6i5amML9qZ/5CcCVRjWJ5HW7oyYmCuThfhDW/G49dgA
Thhp4ZES3KM7rebgFmMLgZtKnplsMK2RScjNfcK1a8owflRxiqSNoYofZJZMbDn3eSmS5N3L40Ng
ayj+ODTnBQZxNFiRRVnIPir+q8//dQPrTLhW9QsN7DHo0oUTOMvs48bTHPX52EVOSvwh3nxkkv/Y
1IJKzdNH1kXw6nIviL/rX7jlTp/Z8J/sVErXSaK9SsTe1rAAPG6SNxRIr9QL3mOZ3UZpNs911E+r
zRp1gHcjwhrfjcCa+/w/kJiqrnTBTPbHJKzu3kor4cGV/NDRUZg3Bsg+YpGrblJpnRfWnJBHuulI
CUdSVhtyQSCZxCZepdsSLUdYA5781KoBZfMuIVQ2dfd6iQWvv/RsjLC5Ar9L5VqRSbi/fNio8Ytr
K/AXo7FRM3Ncku3B7Z0cAkDTHLa0/JjgQrUStT8+oURqyQPbKnkCj32FTw89C2mFR9Qi23OF3HWB
bsQR1ZVCBwnImhQ6GnoeN51x3ObNKN+bxkrHFa+3fMxvV87a0aEcLfCOAkjCbJWGa42l0MvNLO3X
mb6Hh5ardaL6ObbOcOzdFiMqQYf2+BwuVPKkvxo4D2lCn6M38kY2RjmK+YQJkt1RYEHZKbya8m5H
Q67ogRiK8lqrF+gLIYHvoQbZvp953rPp8vwO1zfdNIWhcoHl/nXHHzAg8lbzhdcdqNRIFpSRHyGs
/Qlie1oD9bm1dG0fvCnlbu8FZUwIkj8MKdrw8F3lBYN8mzlJZVW7xpkhO0WQNrLmN5C9rP9NaDiZ
s5834BEPUstoWa+LM4fIRKIGdVKKv9it1kViRA68Hc1a/LkrOE/VhfDCji7Q5Dt0wmNfpAizh50+
D1BWCooPCZy+q7+2Qg/erJ7G01K7A0NzudPebJyruDzmaKKxkaaC43kfPOEmfXCOgsWbXzco4I/L
jjLnBWTPf9qKiVFMq5jTCVvdLzXjlen4jeVhFAbMZo1dkqcno+/LsAAas1R2dm7sLIYLmlIDY3Ms
p1Cnc7Ow8g6bR7lwXjsCZ8tCr0xAhMqINj+jLVW1xe9SP2/fKUnwRA7pphrza+QDYcREAnzIJ0pI
+0TeRsBm3OkYGQNWLpBiJrFfv5OGWz+BBw5f/8h53G5SwRUPthkvxau6Blv83oirhjkLnaOalrXn
S1sJNjPt2rsHg69f+u/cpQUFqOm2L99AFK1CfeuVJm+B11f57flw/RNNtFFbZPE9dV3mu0BqkOoD
f6K8IOddJOPMGxclgKkxJV0mb57LML7urxqel71otc8wxm29FbhzmLbkgaRyOKEn6r5SXbsm5BUb
Sff+h1Glus7bGbk8TJeOK74nCpYXB5xeGSVI9t0hvO1S0aOnKz3aosl/Cx+mqtHJJrnQYDF3+omh
El8FH8V2/v2Cs9MFwSPw4lJ3u304JB4wK9Ob4JIgFWQkskRU139KZZnYT8iHvD6SLcwuZ2ESOfcw
CHEIi3tEzm871/BSDhtYTALgJhWInKKnxTEIiRCoC4U3sTE8qq9FqMOEGizQkgYLr6+UJ+pO3ksk
S8WbEl4NfT8mX93nKgGooe2ZgklD/c/k7F//Eo1rCTXBNQvHscEXea5nGHXlECAGTtM9PtLytoDT
adBRM8fgnltVZZrjHlxQt16pTvNzv8ywc4XQp8+N2CNX0pDiFmEeYic8u4OLg9Hbw2D6oFCVPGDu
UF7oKVoaDXKgXnuWlxkxtuq/7I4kUzXPvWwcD/GUl+2xt6upjhO7g24N7QmkpIsgyTh/E9nIR6oX
7fTLDPuENJ9gfn/XjTBl4fVQuQ7ZFvAHT+Foy/vUtIqKiKWmB8lB4XDifjQAk+KTAZxqt2XQgESI
L8S9N3/4FFT+d+/6BKUs9i1O5DIFFgHsk00RL7l+aNMEPKWS7l2UAJjeqUqG+YSpXqn/ws6EDjY0
G16hYsqprq3sFT8UmGA32qDcc53jz+JoN/qqnrzAhEGu9ncJozYhpUpZwWtDT30mf1LlqHWcUDYL
RyYg/DXEZTI0O4ppBuGyDEZR+rPjgmXyEL9SwHibu8qq+e0jP4VsJm3t/HjrrSyc+oV1ZBr1p2WP
T4oYXOcY6RWnewlpzbaw/RQQhjsSqalsHhLXTijsR8Vum68NFrKHMcUVyYsQEK485D5Thp3FopdB
tt0eHJAuxXJEg+eilGHC193EHZxbqMXYjGW8x5C1Z425iBsHvMsiBxgTxXvBnvbvFf8UaIVpO0Gk
s2toImn43KpjR/xMzQHCaI10ke8C/ISv+0x6qywiDN30qHvUWQtmt8siyj0pu+Chbf3N/EZgRttj
xo1Eo60tr/tWNQjwSx24eSyWwqwqwpAJElmXbKRsUT7ezx0Hs+jJsNjitmDf1ZWMIOce8iS9+/or
Wt2+4DE3cmgf4XFfEzp1B+0sLhpMrB2pvZAxfe2+Ui4uxXIRgQ9KaOQjP581mkzxOb/BCaeZt61f
z4SGLKKQ3hpzLCVlrelUyg2DeRJX9pZ9hEqDHhyDnoq4w8fcBQuAt2R0RBSpcmWi/1qNP7FiK0CP
/gUo1rwTr+YrJUHDqcThMyy7KnAV7+7x9BfE2CyCYGQ2k4lnDZm/u4BP67KTh5zKUEX4zqKBi3xa
GG+nsLMkmfDWYV97iMKhUQqaU/EzYfRuh8MV6n17P8n7qKuY10wnsUHhC4IzesTRLTzVBQ6ugZLQ
PlfkmbIXOTmntqUssvgZ4M6km1+6bhRso1h76/HQiVNtfzCwGejMX0mNklBxjgWVpFL8ZB7AMkgr
vr6ZH4Bcm6hjj6njWWNrs0jruIWMIZ4pK75dZam/7zKxU4JhC+ufLM5KNVewfIW5gn0RThGiKPx2
9bpyoMoVI6CPqGfMQ16qeM8k04Jq7brZ10a5tuEpSprCl586B7fKLIELUyGcU+3kNGMpa5eQYVSP
/vOE4MBByhhBgtOmnaEJjaGDcs1LV6K3o/D8hWuBTkW2y4gmIMbpqND+cafgLkNw5/x7fq8+u8dE
ucGv18NyUJXCWjaRy3DPYKWo6OfGJHzM7IovPp4KwGooeBd5rbNdoJUEQ4hklPunXJxLz/XeoiYU
iSLgH6CKV20OsSRz/1DEYx4wW98oxoplGfFoH/CrFPeUekyN+GpiDB6wNADXy4Iv7bBr3Fav2f4Z
eKrSm8tfprIBXz+H/kxd45++bC6kUhwhCXf3olPOSLSePUs5Kd54T4w2B2JMAb52J+DR0Te2kn55
5zokuGeXaS8xMfXVxMFbc2Vx1euGxkDA4ZdLil5R8x4IIxq6DTSZBg0jI3W0K/LJcxiI1h26O/oc
q/Px2zkOmqITimpdnS9+XShTe/karzBJ4NTNVc1d3ttYN3hOYzt6BbsED1oUXIpQv7La+BgNnDbR
LbZckNXSSlWSRnWBvboJawu8Y5SImMOU0fUYii4PnVIUa7YZo16KNtDoTNiC25s3N3q9yiJBynEt
s8pIzy+9ou4rZ1wxXlMjnZ5b+Dy8YSDWoMw7DKyNJ/R3/9XihYMqVGeWHXrT70IJkfzSnP1uqS6V
ID55Ru6DQ5h8oZrTjqhbl6Y8Wukz9cZNPUVpJMHm0oq0WB0s2mGZzcbV6+ZTLjDjgE976pG9Mcm2
04+TUIxmo/Gi09fRSzmMCySyTs21HkiPDcYd85JrfnrYl5fzb9lRRx6Y0FAuADTTVkHlMpW7eRj8
joFWL9rFIzQi1CpzJpNYLJ6Yy8tcEFsXB7v6JSb4BBYNbW2OoAY2dUB0vj0cOMNaYRi5ufNCEP10
V3I64N2z4FTLcMSArnakT2MKcHNseEzY32US8NoaUyx+dOgy1aJ9o48Shhv/oXqR/QJGDmm+010A
TJ4cI+Oq7lLjt7HOncghJxxSqqUMlenSVzGMu8UE5kL1RFnka3ImNcZMhY4DGyLaC60G/gyYGeeH
mpsTccWDID0eqqqnQbX/jJuRk/KPKcInbJpGGiLExRHvuK+Een5AE4KoavSx+NiC1TgB1Hcgp3dm
29hsIJLEuoyx1AMWRwPwAXABB+lzMxPu+saQ+SlhZbP3AN6PRCXRVSItA76PqwoJQ1SLlW98CyAH
28AkaY0KSsce4TocfTrnANGHZ2SVmiNgoyvMCM9C5+KHiBGQRoWUe1Ngaa4nsVEoEX8fvi7KCR5s
PWmJe+Z79Qr3y4g/XMlRIYgUd1THMDbPNbGjbUewz2zWn0J17ZCpZ5u8OEdayOy5cPv9TvY/fk+b
iOy5vTUR+RjFXxgqwzpUG9hdjjcchq+jIo2B/2ecJwv1hdprz3k0WsRmTzeYcNVBUy7GoxWahbj0
bYb9WW9pZ3psJcgzx/ljz960OEJXTBxC1z1st7v4oThvDeC94hiujxx6FQJxRzow+6LDf2SrQSy4
8LGaxelivoY8xMJAcvrYpXW1sBDKdbKO89BSefUDKXT9yHLsgKUSYqc+2GHu3ZLABiCAONMHteV6
McCGHvJALpDCaMYvJKlis5Vv5I2O9B0HyzhyM0n3ISBW6sM1ET5m0LwAE/sAotBI3Y5EltssqPme
Ka8K3Uk6JcTZm32nY2mrysbn6Oa9rpINBTXZ0pyPbvQ1clstpzyyfBYaktYHSVd6nJhZsmFZZLtv
+sSxNanIQ/h1Z9ZHa0w6If4R5GDC88FItq0urDyUEcswlMoVia0B0XbVo2VpFIFiZZ46nS2VvOdZ
f066YMLkXleSOMYPkF/vECJYXEjbHw7m7zH9+HxSDdQyKMrp4dPQXiqRqbbSBxNUlLSxQO+D6LnO
KsDIXzayYG5e82XXBxI8obFCOuXFbJ9HUmzgO6YuNy1+9/7jvDhynOxrhkMQgc05k/qkLeWzqk9m
T/mprCQRP6BfbChdhi92CdCfgwm1Zs+g5k3F67GkRARlG9hS9lgKMbhKFSq8TIXMdk7ISrj4BHFp
owDuKR/oQB0SzLsL814clOdu+5/lfcE4w0g1OQIA1eC1hQ99jC8G2SfuhMa2qCNmNX3L+dojsPSa
8lu6x9/pD459DB9vEnQ6XrmTIH+3fk8xaumztgZ1LaeY5lM9wzntJ5Yoeh7sZq7b5LcDj+fP2K0v
CvWJKtoIjN7QGBAyZeldi4EOItMFLqffIDS5vIW5fGCvo58typ+1etCBQ39lSVppCLjrnde9wx5/
sJrrIVgALrRgaK39W28binruftt3TGQMvDiUr2XidEZ7aKP+TUPn9p2PpY4NuJTh9eRjEwD/QznX
nfyDnifrl741FQ7AW/srRnuHTau6LaGSth5KmUOhcbFUqHrILcmlTYYk86j8U/VSYyrQQOJWFOQg
oV9k2HFswjscaUoA4TE2c+w/GqIT+FLelXKAPxYDqKkSDDFx53+d6Vduwces3OHsh7E1YPLL4T2m
jJaE0nQCnPRLc2Wys+oELiamR5dTwoSV1cW0hbUOod2Dr9DDUwXqZeSYopBMA3D5JNhRNBSR1dpE
tl60yrkYHkFDoL3BLrjhZmB/GELsDNSseWCOg4Gz3ufyhpFcBm42oEoyh9mkJrmaZCE5IzTu5rQp
KeT3IiwcekWIq8MjeHaZ7u+gKyvEZvMVGT9WbsHgNi2dpCBsVC1cRYHjR+ecg4gbtey3ytGcCeZr
3K/0Z8j+e3uo9lIk/ima4OacCUDlszhnnepRRBRmZ2wIdLnO5S6YBjsc19A0FhvIrvbhUVe3OMED
/YrqMu/NPurG2CF343DbyNlHyZlIQM8d1E0OyMnl8dtlY1pduo2V3xD7isQpYajt3eJj8TxcQyJj
7hd6x/84vCyitr6QwtkMXP83A4fe/yOvh64asCtuiS9pDMxZSw2Y4TA7RWBlTtT6Z1x7ccuoD9KK
x3OBLlBWz2zURCrMCAqLDkOaMzQXyQFjFiWjncQAKPD5VN4KBWHmp0q/L8JStdCSsyuibeclA68H
FSsKioEQhiSNl4b027ZnAH9AiqS0XXbYrfVXCcPcYdmONR7DkCFd0NVnLVA4XdgwcqvkpG9UtVbF
amdT+8OdyJ2x5FvWk7bNuzO6k+k3MT2uCBmozl3ZO6HGiXSHTjolOZWbkff5rerlybbbSgC67ON0
k5VpYXR5AJOhqJ47B8cvjWcyez7AjNl4PKSvHeftqUSeWg4jXVnr8O3dOy60GmR6C1MDRjBMh9na
ebHYr4ZecZ1bxLB5xdTuV06t13qgcyZs21bn2iBv1+LpMr033SLihIUdiIqMuT7nWFEkRp1hTpvl
KNJzMBw6P7pybMek00St7LBpRH53ciJ44R9MQickaOVT9kOPwjDZ7edkD8ThXPfhBQTk2nJ4jx6x
FOmBr2TIGu5i8C7msNU6+ds6errqGguXgSAC5O97PsdwoQfuZk0zIdohnz2adBlwUPn/a1eUNFtx
fsoUFgO0gJ+tY7HM6ppVTEgw2F88zg44IQSiXjoWkKhiFtiJ/jU0XFyvBSpF41Eci5ETJmXo1NPE
Lf5fjO8ZosbY/zgWDUpdylpdnvarPdGesgAJ49CUzI/JxsntNkbUMmBMtF7LFgNv9qIYbM5PTaSe
Gyi5gqCA7oVUZ9aswC1dYHAZBElxYuii5RzvLej+wGsFQ/ZR7DMWYGL+3Cro/ZbacnhxKHnxtvna
DJiWXFP5kNZQJ3aJz4FpAzN9lt1Szf1ep3rQR75VhSm6upxzWksegmUdQiGHGBlowwgCTDYWdnR3
14egsrFx/6+7wiho5bSm5UGbLx8405A9yJF/5C2xuPj/PrfcO32FQKZpD44A/tXYxlApKpH5gFFA
dTiE1I2MENtUcFro3vtPTSmXpw27XRlVEpM1IFzDMo6V/0wvKJQIg49Uy+aKwTG7GSiRNTFLivKZ
F/jATvH4f8/z//ITYcDks0iL3GE6CiJxG1l6pLHHVL5EORYMKbx0Hh5fasZacOVBOdpSuSHwYj8C
NTmB1mEQic9CGa7jPIfqcNlGNJmOf9522LMcOI0e/rBguhiXq93xNs7GMM7sKG/xaYCiS8S8nEFt
Ra4ZWYLzTO7PS0FU+8slaWI6JcWHKHq0Qf2Iic4yshQ3G/u//Ov7TgRJT2buYFQxH3KFYtwSfV/j
6qdpdh/a4crKXQUbBntrLgehbDUabhHGHHcfYxumBIIGegNZGM7bvj/wEiVmrWImJf6h36FoB+Lt
ziZ7ZB6lVxjLvXBzoWsA/AZzXDc35X+KmRVwi2hsffpSJJRAVXpZAZetV9DMV26Z4N4l8C29Njua
m87TuwLaQvgD8puYOIEBtz0EZUFCZuZoZjz/3YvBcnq4CvCsOsNteDy8gyFhApUp3LgdGD1w3Jrs
YWRPeqHXsU44ksz2PPdSg2sXH1FYh7Tz4qTzPf99XyQFrSH8kzYmx1zayb7+clYVaVOyXj3PmheL
ZLS1/hwHkjab7+WPsizAikMqUDFq1G9S9UrJ1eyduSSxU9Y2eJIb9WIaL7nRLEHS4iZz4kGr3XeC
8mP5ryRDVh9R+CQWWxWXf4FnHh2qzOykg2TdGeHd0p4PyqmZz1kUL6+eEeRPNJbmKhljc4Z0zV0D
8ENJKT1bcNHbkrl2JBdWsSSDe6BSalRYXtyj9TeQ8mWWLKnjkVAs+uC4JL3IHONAudToetOh2kJV
BO2/F7NT+3WX7UeWhShguoozn8H+OIV0eeqQoGgjUVPFY1VOaFW6c5+BhT6FMRKJKRpgIG7RkIHI
F5h/EVWDQmqdN9larGI8vIxNNaCHsTC438Vley0372jUxZ33qMNIfxYaLibRHO9uLSC6pQ6yVSB4
oG0T6s3i34hYMhRnhyPltcXz+h4JTAyU7IEwyEzPhv/AYptRnNlWWINkOvGw/jKH4ph6/g7zhDaV
6/bP+v7tExLZ0AwKcISdqY1l3pGABKFs3QET0N8paLJDEKz8AzNHEw4OT87N8kVhnTBTvTv1WI18
aM04L/ysO4SBYCzYAmbEjdWYErGMYJZVGlAPI8j2rK2QbX1CRIwX6RdSGomiy3a6THpVKB9bilC2
o69ZLasmsZy8D6NuPnggNk+2FMoYw+/o3wTHsS8UfZWTuq1eT4QgJYrf1U1H70g+24GO+UeTuGRa
a9TuSC0mDDspTXkA6q9RXm+AnrCZ1dn/JC+YRRvQeX44gXJGHLrufmC7Ghe7Ta3/NrdAjetwtCrd
NJO9cL+KY80VayS1siYH48Wm7xQs1TUI3poXm2vMNSLPcAmEQEMqMetvnjAyJ15cDcSRSDKGAWyJ
p06p88uTOEJSwkWZCzXAYtEn7PTkiazVskWqFCwTFCgMNZnB565fK8Ev5R2lFpDSwzd3vyl4IuNY
171d03/d4qwnzHFxKHI+TkOfXaIEqtTftqhq+ovwLCA9y2QwKbWEQKkXgPK08bmf04wtTHjQKbC/
TJUnRaE6645gArXzhnTEixMZe6Ck8a1+u5R0XS+IDzH23KKHB18kXOv7bZl6OWRhSahQQYibMCE1
u3vddcqTTQ0ccUkiQOx/3hKb9kyABuUtKEWpEwjoKKDCgTgFJypJjgsUjn0GTaUEJqjLDV72B1tD
TuZVXUEoumLJZQNHUIstEZD+HyzUdUiuyUQNztnP5ykrCJMRTTfNq86uTp0lkhoz1Xu5OJN3j/g/
hy+hNP5VFd/KjpJh00B+Nng6N6AWQKTQB+i05O5QS2m7bhGyuvxdo9bp5IDitXtQmGnm6J/FMaCm
cUHY62kCxS0kBRIWg5e3zan4xg9YB64vpw4RnUGCscNYmr+6xIcKJz7tuvKA41xShCz5/e9ZIZ1v
12TxlIlzTcbFAc1XfVeHtPsoHs48OZ5Zkewa/yz/izeJRVZg+uAmmHQcJNNzVzyNogNmtD4aRxIC
knyqbykfbqqUL9CKUMQjqTyLf+GPAUEqpagDbyOEGP7qA3U0XOBJZYCJteyYBWw/824MteQe7gWB
Sef9MALo8jsK5x7lz1631hSSlPE4G/+mr0orsiuNZkgIBQDUOtJiAhx0NlPnBfXqZWM+aSzQSIMW
XE+I5uxmkriq9aIkpTZbJCJZMTAuveysnWVKn9JEbGVqC0VbkrdbihUBCWZ4wwjBfzOdsmOKXIoP
QfLwspX7jMRK7TnHkP5Y2swv5WeZd/jjikt5foyDKsYeC2XnJipbMWXRYEqmwsOk/HI5IdwU9RoU
RXjM6dxe+vqXZXEvineSwxws18U4BdQQ7qfxQXYdIe2HGWLiDdnPqLMwyg0+rH9ErWBXN+su9jPG
2dTjr+J0FHtpC7AF40T/tlwKAzkNP8YEDIWoLyuFViqzexKvWqo8ulWKGhbtdF1DVNaf0wCG6QpF
JkMdMUpoYPKUZy6+56ma/y+BKTuQzwEwGjWuQGP51bfnU7mFrah0ZNcLDE4Nizlnmn9LB1pMDUzH
0CKtcKhKncqifqqLTzZurUUnczQ094Ls+TI3yLnBfr3YLQ2RB4t5atFMT5B213/e2van3B2/w1tr
srUImh+Og/jvC6CfIo0crXYZ3Bf1L7V61rIckUAhA8WS58PCOhIMaU96+MtPpJiac0PcJ1rmkVuP
H3DUIVgwnEXTsS8n/QtVeqCAp7LPouCq903QET66A9ukYVSue+mO4KuzcvNDGkRdV82jef94P6AK
PzXKYDP+Fh6aUmKYg+eQvOcXU4KBTTc9KN3l73rBXaTpAGIh7rIDEM0xnHwM9hwp1Z7NVm37ntqA
C3gP292kIFR/CfE9TwfpegG0hl7Q2LVwST1BWJWmpGANJiT0637wq7gEAytdel2Fp7uYtOXiup/e
b43y4Aj6rYnDL+RqfiNByadfH0/bGJXI8xd2sRzA9R/TtWwFzYQRxqK2I2sNR/I6P8TpPJU6H2RI
wsmu1TvJORhjzf657VQyf+ItPsc2JWQjzNMiPfI4+WNd79OcF5p0SATyadt2MlEivE3O7qTriOCu
wjegnLfK2HoqGXeGq8Qx3TwLWHPZu2g4tNa+3BLRoYATm2+rfveCoBMUOTwTnSkbrKdBz8Boha0H
K7Iqnk5FMPT87wV4qGwgdGi51+Swz5P2FWmd2yG3bdPTpPuK5cI8qQYctkMfcuaB4mQZ8ASlj1qZ
rELTR+xxLs88AddUTfx1yC7neCW6WO2zYFYo55k0XXTPkgFmnsJUqVnkQvFojjSbO17E2OTx9B9p
7abEh8DDE6msgUCUIYqhv/7RoJwLRH31P5XdZdrNLsJcosHB/0IwH6CHqYOU0aloDH/Qox1rYcK+
wb1iV8tIjhn51W7fo0xo5xieo57tKCo5MjJVXHAcOXX1i3+kBI36dY9Ce3I014bgS3SLzfE0sV6D
u3JmTZ51I22mZsX4ia0QySiSGGv1PvgSkNwEWE/cUterbOWUWNXvIpyox6aoHX6HiO2fWdHzq6m9
8snmSJYnsb/0e0Cejo+GNGbhBVxyZ17MVtZqCOktgC0quK8vTeFixgSqT9WewiYIU/IkuhxfVWP4
I0VBXkwUyPDQVVLWr2BnMx2mVhPqa9UqdRJLCR1P/ldngocr5H4n4nifp8muHzBQtgtreinqsAPI
6bvK7z1WxgZyBd6OefRlOfY4txmXnpDT6nuww6b5nfa7YUJSY1jPPzsA9xiqduY3HE55wxib9OHU
gjCvU8tuUC8D31RHQuKbdFxjYzWhrfS1Xv3nkk4X0KJ7J9FWGAKZ0I0KCy6fMk6K6Mp0FBsvoBAN
hlcT3zZSxLLTvr0Svzjcqbea1pl/tbBtuDDP3MPE0O/tfsgIkTDxEkNzaJYNt5UOZpTAABDXAO+u
dgQqPLNnhvctfprAMs+i0xrPoRWndM9x0wfTzxBrBByNPIqxoBbYh2vq65QeicdMzwbjd6RGJvmC
PQ95aOmDHzjIeyNj3mQ1inV+atAmmBJ+tqJaO2UDJ8I+a2dZNmj/4TLX4HzQdxBJWlR17ks2Sylt
WLLsagGFKOzGrfzQh6qehEO2d2KVNGp3miydNqOE0+l+CA3eOoHz+EZ06BLbFCYEdp2EwvXzvjlh
WRh3ZlCm9EOp94dVYI6XpzX/hqoH5l2/G74LVPz8oCVEA4svJTcCUxNes7qRYUnoTEji6TrVhaPW
K+CHpzUVnRG5Wts2AoEPYo9EeNhtxt+kAoMtEYw1AtzV377yhmW4/5zO0B/+KDM9tiXVBEp8u5Pa
lTQw/uZV/QNODHeSHcHmTkOlL8Y1yq6dzdU6jg+M9uxfpvKZnursy260hvlKrsHZHcr7xewbl5iJ
pOLUlTKcA6KwD8/p2cyZtwqV7wRF9bfLJUXNjfaskLQq7kcJZz4DikrUNFVirc+5ZHQIDgXJcZe8
Xuf5spo8VpxOotRAxu/HHJ+uPWF8gmiKLKBOcTDwFDjH5Iq5834Dy8DRRFBIxVi3FvlfcZ92JAbV
r7lpnqaDSrEgoNpLNYArAmbf6Eop3YJecb2sUPUKNuYyrGgVFpD3o1Ug+aGwabsudxOLfqRIdZaT
aMIH+fLldFoH/fLhsrksd641WW4wEXbprAiBLE2dqMiKO+GCfqDYYCRZYPA6IbzS8+wMcPKAyH6w
kQNUPROe9oJon2susGZdUz1Wrj/zPnIXquLYsrFBnGGHERURqMnK2PmT4l0hcBF4NHhPXZ9ZYu7k
NLrx1m1fuiQGWuk8dlu6WobFZ9LsA6KHj10jSPq1wyvvZa594reSl+M0+DnGExRF5Sx5ryaKZFoK
9BwKussObWdvovFFFekdTnPL+QcxHmFfR32DZ8e0mqK7Zorqp/Hfa6yagFENF04I955XjWSk6WtW
qLia2LL+U8pROTVtwq9KjV+IDdUXz/Z995j3hWf9UGbv9ULcpCeWmmhsj0T8aRExOfAg+1jrTmo0
rxLVUX3ZlYOUUo4YY/zfrYEj3U48lhK/077BpABXP+ooiLDLt3ZsUsEcXjvXn0CyQBulTGWWgGRr
MMEKhMPoMau/2yv7y5EgLqm48VhF9u6NIC1kJ/QNRw2EJSQQzfsljiXhVegYwVNEBUERDzkag0jW
IFFmycYRiDba3NqBSrPCLycxn6YbqihxR5riKk5ezykj6jhGLdnDYCCNAm9zcdhQQs3JCE2k64Tu
884nE4RQf+vp/jZS8SFdZvoVKQ+efbFY2uvio3zn2EGInmgBnYCnQU2wnqZsDqAX9FOWqcG2/gxR
uuDUqMA7MsxVRfxLPoJTSXNU4SGrsJv+mqDv4u39upJF4J/iHdwtvMkf/rJNObljutJ7iabObVvp
Ixsb0CHGgwMuFtbZzDLyNmqYPadb+DnQzYY2YEyUzlpABpItViuY8ufeGq24zwTNUDW/nOdyVOUI
3gtGyoDQnGVHL4lH6SWwYfAbJZ0UTefnnUEJVnF2Vhchj4LAiLFjdLy7KzIWq8zM4HicxweogP8u
bM8YW8UPr3dboTetJvQhCyFjCb/WPYiZ7gRUK8KupKTjwDsTNDMMvmFDvMHP2O6qkEZ6Xep0+WPl
c1rpI8dg3Xba0/yGibuyFU8Mm1WtmpVzAZ7yd7EcNyH3rzogzQA6gSWOwuFYW9US3unuOwN3W5aV
/1hu7IX3Kqlg7F7+ekn+MzxJEMXaraxO6aSzRoodpWUki6dbidbsV0rMD6L/W09rq1WjLR1xjVwr
a2SMRnUR14XlD3lE0ZTN+n8bbIzC1PitzHQeGs9lCav7pSnCWCYyshE9u06Z+PDsunkFUPa2j4Ai
jGLnMpbxJ7Snundm8yPSoQQWpnpCMFw1Aygk0IyNveDBX0dQUa/zzClOl7g8QwV4O5fz8BtCdIKk
gscbquZL2/nrnkxaq7zMA0demnpEyyYnPx2/1Sr/r/wn5iRlEMZA/5IEXDDnOaVZldETteAf4FSd
9ipc8cTsWcLXKiD1kWRsNgTw727ZLBJqHgq1tztyO5Uvt38OSSX1nCh+CIyYP/czjSPAl44fuiX2
IALbMBCXJSMa35nw3iv1v51JmLf+gGgFb+I9kRfago3QwUSiHIZ+JDbnfS6tqxVclEdePUHCGqQF
KouLavNObzUZp5SzlL0EMA1RDsbzO5Dd1A263JCf5z7SQTqLx7FqNiEFv5LQvBMADdyjFOzRBRYO
EcI1I4AvM8KN1BEAbLDGJlXBbqvLEIDUOAKaME30ZtG3vF+81+ALf/wBZKDoy0unqK8cOZt4ve0h
U0k4U1VsjrvDpfe3WAqbNAGjTNgJET1ITsXYQJkFe0L6WPIkzkG3FTMN7oI/Bte2E6YNS3up80gQ
jfyYq/CyZ5zEarTEDoUnw442MzxITWrLFplgItKHFgNpKnBJGv+O2EyS9xuecm1t5Kd6gM8bbwX5
tIFapxco+Vkyl9kT+hifq6kWAfWJmwu9UlWOKdVdM9nVerqP0R85vvzqKFSJK3TiW++K0bNYLXDa
fFynj+BGHDmKKWPKOndCS2xHgF2i+QuUQd0b9zC8aJXIuHBy1JFSg0yd+I+8ALjqpH6J9j6KsP8H
/3mz3yHk4HKRUIfcI958mUSij+w76xg2vOm0aFEgFRSwVn/6lD/WAhpN2/we7+oIIwjS/dpRB75G
vUWZfKmlu0GYP/vhVMpbgj5FjASFKkdZSNrsi7opB/INjno5Mc41kqGv0yhZRV1KdwH55gwIKgF9
SXsIDDO+U2NuLrf7AH4KSxX+jQ8Tony9REpCtDSOEg5buJlG94+FGXGzwap5ljd3zGTucng7QkGZ
WuYhu7R3tBYwK6TD0cnGmSoSQatFLmY+YDqdRnVJopQ9wX48aUFdNQF28jpJ+LcF7Hn7C/o1tWi2
ejBcUpN/czh4a6yLYLygV2HM3eavQrVYEamELtJdGINe8Abp9lfWAOrOwL5RnIjZJUngxv7+ncSU
SQegnZLpVKQfCXk2r35HEtkhpswW3bAP1wIWk3zKy2Ul2pHw3TWntS9eeOff2HuhbIYT+N2op2lX
/uSUoaFlJ8TgFFxkyMY7N6Zs4X0K04kS/7x9d0bdAveR4PQzvl+V6C3Jug9OCIy+fP7Q7KpaPk+U
jyVbb/mBgA7g/8XPE/EUHOu1ZbELRxu0YT6hwBzFr8AjO2wF189b40YCxKxnmPV+bdEGMtoCbd6w
NooiegM9VlDwe04AP74RuBIftob0hr3HnQIXG7Mj25Y3lfNWlm/xZTlEh6TqrfUuo1LZcy1bMt0k
4uIuLbBO0xYBNI+hpYrR7e8Q/Mf79MK0obvLtjimzJJmcpce6RFQALzDnIOtDrbM5IXHohrtVXTU
jnmvxtboB0SEuf8Ws0k20e5ZqhV8Q3tmRo1sMF7p6uMOsjKeDU38RY1uV4GgCH99Qw4zV/yz2XvE
Ae6PjdY0EVHJVPvhnGJKw5JfEjJJ/8mm5BcqO8pUbNVZYcRiXtxHXGYFiY79yqBqLqqsxNpgzEvq
mjQ3MHpdPihOdxy7b55uj7Obsp9nIts8on7xHnr6W66QjF3SKqikXN0W9fNDIxegJ3+wz7ECaMlz
n2hy8wngjmrOeXuAF3Gg4ezWs4TtiVZgw7Wa9N1JmTzmDupfbBAFwOblQtQU1vTrSoB7Zg0Rh9PQ
t2m73w6yZG+ugHv5UaphgTAaFGAW9G/+Dll5lG8ZLG+tqovv109rd2s4pl6IQv3CoTR18h3bTBUU
IcPfHEDW2lPc07z1la3/R8ZPg99vR6wWP3nLfpG3FmAqi4TS69y+aGKw8EmFJ/NG5rIneXuzUJNY
LnwgCnWJJGWoCYOJ1YiLtrNVk3o+68taWLLdiYY4SkxkVpjKq842Q2AI6s6SwqUygDgjR3/X8Jux
qQYmws5rlA0ehlNv3d9Ib1g9NH4DSzTti1U9iexW3CI+d7ylVbPYKHohT0pOVw7Yb5Cfak4XEqOJ
DKQTG+SGPM/dT/Y+GJvYVMoe+CATe3fj2limURuW/mQ+xwN4OmT91Q5JrJXC64/0V20NthYywJtb
V56QnJp1WXKaYQvC7jxwFfwQ9Zy7g8Bsl2k3GDCF8fc/DafFoayE/XnrzXASHn/Q9DpxRNGgHwgp
6AA2M9rrUP427x0Pp9VSu2QaiS9GT5NIpQpYb7vQnaclWtteCMQXDiRrGXDl8cSS2/hpff9jtjfP
6Lg5hReQ21cvDP42myR4oKlpovSYWSRPxxFoeD5D6F7Ey0WVcgzeB6vVA6Bu/r8H0994N/Uq6mEg
QJn+yW7NTZ+nbltkdZsF6QSBYZ5Rtv6S9/GhO22WPL+LCuVo6TY/74LYDIU6S2gQUeZn4eVOTcFT
sgzU9qg5Jyt3ue5ZHTBiuDkGUubfcWOfFHVGZWsknZVRlAil/aUwMrFg54CWZy858f3PHt1aqPJb
GKWsb0HVfp8VOsIfgR45s3RGKwGfxKmGBpzmEnE+AZ6Tet9I0eXTVsMJs3BQebU4gqlE9AeMM3QY
Oraw2AI/pfeuvVkzmu3CdWtC9VSadkQdoFUrxmoQ1M2ANuvpK3w5QeSln7B6PqQaXctlncJuTI0a
N2+lUhiJ0ockb5n9vjPda6JolwLF7yk5uI0NPNW1OSlMutiJoob52Lvdt2ONGNzPCwbriJ05A9bj
Tw84374OhK1ScxFYxrMBbwQrslrnWjamK7hyxrNvQw0R38+pd64s10CEh4L6Tjpu/HdErsyCiIK5
z2tZ7cPtZjKTu2wMj3SzWidxP7QrA1fjaTXB9x8eMnGLMz8SJWKTD6B4qFubaXt9JBUbrHWl4FbW
TWmWciTp8aGoRtOGAlCzWRRWmZZc+8d74dEwpuvSpbRj74yhll/m5ucyGXVwUYEVUjDIla/u5iKc
kGwfmShMOKkTWT4mwYc0HlhL3SUY1m9PhnZa/etZAleoW0AogaQ4eXRYxxmdqPz/Q61elmrYQl5T
DR6z2g2kQXUUM+NpWAxGSouY+qSiVoYhKOD1w0taqXZY2/cSrjGY68sSSK83b5FuWuoCXRBqxnxQ
FEfEXjfPzWL2tRwyBsaVRLMWWxbm1AO/hbxceLm5GuyWZDVpWnijfhlnUtZktOe5VulgIGUmETof
nxGF0H0dDZbbNwNWpzXgalH2R+8qpDRthwG//1V6arbEqYCg/S8zNojskfQkAmF5iHxpBVzPHk/A
/poap5S+UOXa2T93MWOaj+62lTVNeOLJYNAY2SfmOk77dCNZFNQGOQEiKi6tyb986s7QWWiFp1PC
yuAW6YcETv1VX+XSWwkiCH0lMzOHhx6Wr3BKN8/banADUYl9euR1PsnfunRMjAK4MKJumXeLpelm
VVyX1VicIzQBd9yw3dTw4cX/v/EwMO/FdnnwITS5QzHhtVmXtNTVrmdZ8Hi2/dFE/K30CeCZx8Gq
vuAoTP/cDvJDh72nwYB0eLQlntRNJfItExp+0IBcmHnU75L5YdnLUEAzIaOFQKI8dKGiCZDKh5NU
WiEafCp+xxoy9m+6+POQvypyFEtcuS4M32bBrJcWCm3epZPIUpDMKeZGmSa/IdN7S+1gyBpUujfV
26A2hVGqh0Xfym86uGwtbRLP8WLi0sIvEzMUgXM2h/+N46YQLwcx5LO1SbePq2IAU/lrrYp+EzDH
9Itbn/ek0tqp7Ck+Aki3lBRpbUkmhQXz800mDkX6vnG2/aYc8Q4UnuEtFXKp3aA7Tu3tw7tT8A5I
lCHyeqAXnnzZdas0ye89InhZoZyvxlcTMpEzPtAODLBo0RCY4v9FVOhbiuDvWmhE6bstTr/WtA5n
o1LWJB49O383qXx6hxh+ngyJmO9a3k4iloIVbeuAH+BHTSKSNQ7aGDQpDidtizSMUP58bQPlql05
gdZC7gU1MvuXh1G7A+XitxQ933blT61E66lk/mcVC3oWzsZ/RTTGJ7SzxWmsOPCNyh6gTbjEvADX
rdliVucNCQGssFcWA66f6/SC4/9W8NrRiMcrIqyZkt/ATDb8Hc+FeWOQnuz1RCk2Bf9ZCnhBrHia
rRjVm19pfNhppL62scfZlEfys8GlvksHsOOhWn+I273bEf0gqUbiQKTWluexrpMltcCuRZLA2Zn1
7NmGN9XtPCpYOlz0SGRPTdD9cezjYRqwfQh3i6x9cGzCjuVZW4Ac/jkIvPYs4Zoz16LH0dcPP9N7
3ft2e+zzehbjk9TjR8o7lATain/M61jOf90HIEj7r0vukk3ofj3alw7qh5tTaSegdyU7q2GjcJT+
MoPS7F9AbtynCFtnBjKBIyUHgIDVK/S3GAPrCSKKgJsNx5JBeeyvRk9NUBgqNp0GpV+UpKsdy1S7
HMuSyvsXZjI4AU1j53WLzq9ILCyjGlH5AzXECxjSx4x+UloxYkXxalxb7xh21n6fLq624wI60fv/
0MRbMkGYkE8zaJbCp0TKPfrDfK8rjfeuSNxV7rYM2swjGV/rdb6fQozuV2gzoLCwqUVf+PlXpWZX
cNz2wQRdQdd/xmVSxbUJBZ/hsZNPKjvqxudyzqS6A7406lP7soMDMSzdgB0aLrnH0oQOMCIaG5G0
fEKwQiqk9I0vhtiY8uaCS2SLs5SqhrFCljdyTUaoBPwedk8ZJiJnIRQb9tJtbuL3PT7qtt5wXCbZ
6ceBoHF+JjUmXyX84z7cVItJTxoGA1ypKscQ572F0BoPk8KZlTEIXyr1liUjWPKodktqCBeG5/x8
sNavyJb9sqxnf6AO9VeI3WAQv12jgEEhXagRS7xj9WI3sfCo8QjzbouGb/q+lPN2TGPriYaQcD24
3QnEShdiFnxoZwBQ5c8GQzX+uBgpk2pGt5SId08R5ED2QiyiAz4BUzOPB1SaFXlb7hhN9EdKwY5y
9YRbW/nyaTkV5+WXmNjpZ+B2Ar0EOCem5wWuZAbOxhtqN0xItWQKamjrB1LZ4LSgVBKIhVEffW9b
8Qgy7/fMVD5Zv4MKy2Yt/i4USF5URKqVXTckAm2+OeVt426KBMg8qvWXO0EU/p1AIRlajp6aVXoT
dMpYO+ghPKEfScbb/UuEItxYCUuZGZGUKoJQyxawVEAKf9MHrWdojVsJSbhCzWNszm1TMEwD78SS
6tB8PoircGdR+pHYlE6wy5bUSGWvT5lhDuShqc5dbooqwqKKt4Uwa+/0mGB33u4ZwJ9UOnttcXp/
iGOmbRQF0c8qNC6gvqd56JsumwpnRISUvL2r7f0HI16zVJDDbqEI/GIMk4WI1OrLAqvd5G6KiOa8
hqGqrFyAWBm+0hcVlFaRa5NZUnzwM3OxP/zRI39gq9RCBVO/kfdO8l0BIBBtN4pFzAYbm7M3xoA2
iKg6JkvMtyzieI9uKyTva2qBSdi15DCu5qWrJuapY4Uh/D5w7yXdc96EARxmjLX0HaDejN6Rgcsi
lD5QFJL01RxctupsVtN6o2F4rxEhHK/V69g08nu1ZE+lApDKJ+8mIcsObLhwFbHz9CqvD97U58os
9vT3G87XV2p7iOmTR9CIHBFGKzY+z5TS48wSeGAKA5/tiiXHAO4POwtQarV9QTAaJ9hQRLG+UY14
PZkFKfA7AChvE48cN8wTiEJhia+xZZ/uzOL4WdRYO0D3+8XmR36ABYmWDLtXH+dhAQJfSJQOX3kI
v/takk+Wj0XYJdkMEe8vQmdLJveJJAuVkxyWkPbKIkPgHdrAU3AA9P3sB5761dljFfx0bwQxkZf8
ya6ukVdBxATbsV/fw9FdReCdNEqusW1uBwUWJO/0+9wXCO5sD59IO7vaANahjx9a0ubNtFiqDYR1
YzB9h38Y8hj5IKKmgVCMq7939PmciXg9ai439pYMk5T4pBJx7ALeaOsw23ivezQboaudMFN1N6Fv
O+vvUZ/NIwqXNhNS3TsUccds1Lu3tKol8akAgAnQZ143UIJHhl+qOeCTvMr6o5e6+K/3L2+wxMjy
OdFLPI+RPIyMZD8tkcWDAU1NtIRmwuWw2q55TBp610bsd5cL7OFqw+9rhEzk/NlK438A6dDeGdDB
sVm1zNpb9jng/pF/UqBfz+0tY2v50eXfFrrWw6HReR3syiB2sjfxTEyjRV1QjaqOna3zad0zDO2s
CtTBuuQ0aVXszcI8UgOYTBjDfDbtvnxlmajxJA2EK6JEL07/W56xNs5L+r8MxFRJLQOnv0QEOk3I
UOEatvJ7yLJ1FT9VeoqqntM6TFA7aaNbEpPFNYGYirE/iYP1a1ZAw+CgOHridH8A51s+4u/0yg/y
t9NBTMm7PMufZnZAJZKh4ilMiXWEImdrcjUWs3GQtQQQ74oJrWivfImZ12RtJyOFENJXJ30lfdfR
WJzWcqsDB8gZaqNTSX6iBI4XBtpBLhPe0s6VZt4Twwa2xOfNU8E0rT7D1liEV8hOyli2HqqCe0io
WoRw/R7hmlvu9BUrLx4MapAEFTVzF0xH5kgD+btsC5mjJv+oEb+l/6aeE5/XY+5yW8yFFzT4Nv6i
NRHkDLIovXRXJr5VhaWTp96ISI68eMnp6j5yKn/V9zqOOPFjE5Eqln1mhrDsQiGGGJFT1fET3Lu0
B3UrzNg5YJz2ZvcCnFay9GjZ0uxeot/IpcTyWnyX0NDPu2lfsDCuZ6OBRWTea1AdoDWvnJsVpMYt
eFRXfd3VBK+iExPqVQaEp59huB9PO3x7fz82kYbs1ktDstdxm7RJcuDAPYhUa9ljstI/6IpT4DHo
MSYez5qP2uRClzeqdrET3msKsnqzS8pTp5mLoulOTx2LgI/DBtJsLOhylOwDlMiG7k9vXGlSzeWf
T0k0ZQFGn1orNRYi6o4MR+pjuBsQmLpoJeWiDoYyqkKn6dF7LjoI6nfh5568IwTTE3tZvJFkrXQ8
aOwi9beQcAWl+Q36/UqtUWpXx1TOtG35MDmvlUsdVILPF/MMToAwJRpR1lVS5bEhh5JMVb+m0PAG
AoyIAzW8WyLBbdhfZv9E+5qyXUa8DvIvIwDQ029/bsaVv17jeHlOpqo4yfwiAHrQDWMA5ddUf6B5
WfCH73PrGfzPOSUBqjZT1TWyKL6rD0Bm5yUGV27TcAJtvEEk605cOhBjiBhj1QQHt6f7shM60qCo
tRedECn3oM+qmlHt+2dIGUQiERxOvXhKWa0Cxp19BKrs83fDD0wljGBm/nshrOf++8kga2QDXgi/
ryEVRWhA5jHJH9Q0pEXpl6fEYb209T2M1LNCTz3Cu+SYJP2IONTa3P2HJBDimi5JBA+qL/lDtuQl
b2io1VD41PumWS0/LZ5IicE8Y9waeUTSz9PpIJMfVWwaMTj6mDgRPfFwZbXAYoIl5U4mOjpW4G1N
c7SEdHtk8KZWxzSPDBxspVTKo+FR1yyj43+fmN7xQ05i4nvFa5zfUvNMrOPnp58iD6yAl3n9phNg
pcSpOUcChLdxa9mVYARq3AAPchFyHxnnsc43zStspdo99kTV1S6ueKQC73pEBURi+L8rJg/afO5v
u7RqxQIdzc+DsHK4IJtY0JWlZgEQvqsiTVpSC7m5mL7oHJNzsiBOh+47E9JcGhfliThUlHaL9UvM
0xAa00Iu+a+Q/OAUQseTCU0iz4j+lVX6VRrg87oM0LsCOepUlh8WZroRZFctq4ogAjtO/3renmR6
MMqQj5KRLLOkSjRrVrtLEP2KrFBFzGxGUvIDQKE1+v+/S6vkNbwP5fQLhmA3wa+WoCkUDXxphZ63
2TFTdPm83dbUSXJx/hS6HVEQ3xGpJ2YvPuoD52iHuCrJKpoQKhjhfOmiurpe4T7u/DqV5AoeW2Ld
7sjvBZBpRanqcryjdW0UtNQkQTHARBwO882vmj/+4DAil0qmJNSRRefcQbK6j0I2WRdhu99O/TWm
q/tEmCmcFu/LAd8vUnW+rGrCOnZB7q7CZwSb/Y5kVHX+G4C/UolBPwYk7VCpP+ZbZoX+eYczxqyU
IMaWmort0Jh7h5vvk5QFWo8II0AaHtFW7Ezr9uowlF7gK3LaAeypvkIvE3mtzzTj0J3QopYKl/dE
u8+MwrOAoU0sP+ZaVd23fTEjQg5piaqeJAsAkxUH57hpuk8D3jPQMD+1y+xpKmDLq6XTrpFwuIN4
HVVljapCvWYtuciCl/IQILZDjPjlSNpT1LcoscV0xiPp/NuD0RUBpdkZ2BTQi7h0437I4AlhSBs3
2Il/JAG9cnuMRYP841FFj1Y83bwewr1eAl+LF8yotoXMwVHcXM8ubOkIedWqGG+lluiEAa86RMNM
TIcQuXHNprqe2LtqxDkY4bEOZDJjfE+XZDcLW/UnNeEyEJTv1Tz3pGdk8i1sPBPbGh484VKNA502
Un52wry/zbBaaRqndseqJugEQ0Jb5A/OFPmsq6iP3oY+Bwx9gJNRtsnBW4mBucLcUWr084yrXCWf
4m8DqJSpgtiEhw8PZ1yx+6EL3ad3FsFZlrU4W7Tk41iTdLBsbqSkQ8K0+eU6ZkbO6xvh0vk2trG7
O3hdl/Kx0E2qW0mloJ6dBssYZscG2hxZr3h46fBHAnCaNttkm5yzfkFIS04pTaA/eN6D1QD50K0l
pDrcUpWKIEwz79g3VzaZx+ac+J+Ab7J6G0IkjkankffoUn52ummaovX2Noay3GkgTkQTQQ7Mwlue
p0nPxtIO0iMwxPDyYWWe1PoaJz1ZWOgt21yBnaXc3xW4BVc6htniE5doPK4weecahDDln92CTrB1
M8cFgZpaYTe2VyXbM9duot18qAuB4KrNCu9AOhmO539HKU5BCsP0IA5OC/LAmGB9UKPz0tL7bDXj
A99hlywCUmZPLYVJACOwf0LpQL4096KpTxtbzOOJp5wTyojFK5Z5/prvVqWh9IegXnM09Rno6OwK
gVp1uAlhS2RVUocqsgYsYc11DO6B0MSOXXLnovQjPW+rU2rJ6KmApR1r7BzHs5MjYw/cr+zVegRC
jjlBep7wxwUJ4eeiblJ4lIHxbblpWv1yKb/iFygDd4i1qS5EirR5NF0IYDyCgUEshQqb4sWJNo66
JRpZfMXXzrirOIsCdSBEcb8gmCZ6wKUeqDRIcpqVEf8sU/siGKFiwVO5j7FvVNNXhkeHx7SbbrIb
wZDAffvQRQTupqhlo+0huFb5vPvXtt0UcTzIzrr22KCtTD9if5hAWZwwd+9stKI1TDtdz9rPEtPA
wAl1jamMNCy94FpNwYvxgg8rrVfYVdNUHYOS+jIlFRVL0BzNFi4C/pDQ2kGSYOOmri/r0MfikBva
E3qylj1M2b/H9LyMb5TXIlFmOTTBtzNsbSfGLkFMFE4/SNeoEy6SmVRwCkGCc5/5/bjVAs3Dg968
qmWDl2D+F0TAMPad48C6BAhm/8RFRKUYJNvJB4J3yR0HDmQrHlZRcUshsV8F63alfafpEM7leZ9a
w/XPIQkpXFWuyAWoUCw6mxldwssAjIS5CzfB79xx3XUbmcRNL6g8+MrEDSTk72D33/f/5aGxWsTK
B6EuYhaxaNYJYnW1U0YL/uIyNURVQ9hVj9OZco7Om7WCtH6mQqPTbu6RlqIeGBYN2FIOOj6wy6y5
P/819Dc3q+Q5tq03cHweIeO9+sfZEOxBgNBzXjYSpFWpsZW6a8+bnq6jT7+NKOCk9Q8H7j7gozBg
So3zZPWLGUEk3m9zU890IyKAH0Bgh5K9/jnTCxIAVnK3CmdiXuJDetx1dWxEpt9BiiJK/l+aY41B
KbStX6UEi0dfH00cqnC7jtKSiVWo6FRc6czhz10qBhkA+4REDhaL8rN/Ke6775jlddTRRudoRJon
/1C/dJVDmLEc7B0QKF318EkVH43BYt5PaMyaygj8v+K3yEr57GcWtavGk9qWdciU2hAjkFxdS+P7
AhF3Xhzocvr14bKMXpIccGEPWSKviwM1PVlFinrHDwO7HgBbtlHPoP2MS1I5FLKJe7gmdKC58hpn
Sezguh1dxC+kbJpEiEp8XNe41VDYpe4RzOHqgmTfIsxO6TveEoTOAwKX2R8m5JZxzP0ZtjCQXo3s
nS8dYahsa4arc1GkYUuL0++Hn0Sqe4bpOPCdpx82FFh1nFXyuif35o2mXmUYgUhkXGIcEKWmeJjX
KbXl0my9E3y9W7WGXahTffzUU6kR1rsWhr1VCQ+6ci/j+SltaXNTJQ0cbo2KycGv7vj6IIzZF9L0
HPVrwsW42oN7xyQJjypCgiw7BflFqicF5E9imQGDwav1ygTQRnfJd9CUk5oMzj3G8U/yPa8Y/nEq
zJfQtfzJCDltE+CJ2yV7vCphpNAu4tlxVE8vco7KJUvkUkBkoufEliH1mSRmOvJkbuMoyD1SA0Ro
w5GuITzHPyMWTbpeOtOyvnAFovbvjHtn8QHeUknm1wFAbZUwKz8PZQxgx16doUwbxy/sJG8lS3cL
2tegLVdsI+4VoVHt7RYx34BGWQTewdEXTgUvT2HWyyzejCFW6GhrKbeYmRwNFBNfuTkTgM3TU/zb
/jGKqL/bgAeGUzioPyA7i3uMEC0tUku5U6enCiubuJ1lX3Xe8GFrpU6nbKgJO0ihXIl05yivQX2c
R8GzuJa7KHvMQ8hoHTCjTUPl0yHcoLhx9fFKuW1tsG68Gs2XiXB5hsCAdcYNd0HRAVWnkW9aeJab
6sJJbYVsQqI6O9Jf9dtrOH2Z3AgOWgj3sPBROL6xWaXwwd/Ec/5wa1w24CwMi1HP3LLCgxryAIng
0AQ2yrdUW3LTD1I+W7c51A4/c2G2YUeCU665+sFDt2jXP5TBdDytb+BtTf8trfZVcBrMylUx9Zqq
gSGziDy/rL9EjFDAQHsPqEQpXlSRIWEyJn4pDUxlQXtIxLSdmTjw39Qn5iccAQlHXWDuTxXZHV3E
Nn5wCJD80rikpRLqaVIBN3cLPtwltgbzywdn+FOxADV/YDmKZP6JmPUEyEuk9KrnXd3chu1UAdTA
8E+8Ri4IQAGM7x6U0ys1rCOJnkGrk5BXhH/krLqXaxAe2SZzHgS+3VRTqA3nQCZcNzJskpcSawz/
WS+8AF3fc8mKyqX5N7g4piRcotbxsLU2Qm1wi1iHrt9lJLFnXAznwCtP85Xa82XuttpClHGZM9v9
QSzbTdq0BkHfEKLyZLbCwF+GYsLK+YcRZbru4vPz3LbdgBe0OUtHheqn6k/8Tphv4hJ7iuwxiImu
I6lPgFeJXquNsaTeXg1VPvHBxA0HmlV2OitQ7dcEuwBFg3r41bi7Mt0jMTjClqIECy5WRBhtFX8F
cDN4n0jl4nOT4a8bCwiIrfRcU1ktKsB57fxNkr7p247nsID8BHIUKaa/OuuliHQtkdOVkhGp/2/P
u2mcjTCGSGpyZevA1RUa39R+KaMa6tVEjVFwTHpENNXQgT4nCesBRkFUYS4gMKWItVADVAeTUM7M
IlBSTQ973UueXcRdh+WAR+cUPankzZbT7DUsavrhiEBVvkTiGVDhx5huiW0DlLMB3MMlWbJwkkUZ
fPkBCxWFHdJVt5TnDHXdqbeN2QFsuGzIk01QVlXdVvivBouUXeN4XjtcAmuIbD8lSPmqkWKRsIYq
e2PAohhM0YHvgiClFV8zSRX1t7uYn/LA5wcRBDeB8h448AufWQhZIMe7/Na3XsYgOLgeYyvFd+z0
3SxztjSGiYXqQoLb9xSr9OnCDWNYNHDLV6wO3/ridJILt7Tj65Y53/OPKmXLPpBIRa2P1VjRecCK
TXeu9+bgpWkQyM6hFvADFoLS+hick5Ngy1RbytZFxB/LO0BYxCGjPS9jhSaeRJ81XxfzBjPMchlc
HGAkJw1ZUnQpW6fT8ZrXAnA0YqQYT6wBDIIy/ZUduzgmPzWRekCwx+siVhAgpkwOLgbwQBWyxXrZ
0yX/h2RE1w0vlh/InYQjCpxXrS4KwdCehePlHPC0FoJ6wxM9vh2fcVQrS2K+AeGRkXG5CeVZ7wYl
+7bqPDH20vB7Fe2uGBs/0pXEuA/a6Vh5AGHKPPUFxCH45ZhzzvFskTN8Ws/+E/nfichg9tJfkaxN
mS5IgoXck5ZQN4sF4lbObRO20c5qCFNYZJQHSwbsB6vDIedPqqe0AKe+VIgLHEimwHXjOPo3RYWa
9r+G1l4BVeQFz3jAXDk61AtYZmReAgYZttAf+jYzUwT14yWeMz4aB0OILHoSYVlEjRHpRgDRiH5z
zkyiQL1JH9Gji2VLyFECGwWD6XBtdJDJhZb/p7HliqCd0GYWuE9L0Hj8R/4lE0jyfQFbhpe2axvm
q+4ejy+h89+Vvv3UedKSUBLJufROt0QCpTwAPJkOvPOSxa5epP2mj2BfgCRsga2CBWU67EXw2hRL
Ydpq3JYrnSof/+XBwIOBWLJzVnzgefwpW6fr4roLrty0QPEjoxu0Ll/QeimwR56cQ1aH900w0yTp
IRVGFH+RzAnw12MTvCiiRpTfkb/I3jz8HMTjklf/EUurXNReCYb4Aesxa6RGaD/tLQEWlkKPHNs1
Z5l+yoxi36WpHUoCal5ajlr3VFPtgJdIWtsFeQCa924iiqN5DM6GbFaUdk6CquH1KbwoQOy2xqvy
cftVs6ME1y3bBaKJy75w3q9tymqw+jQArS9bgzCGl2JaiNcTTaP/o1md3470flEkAdkmTC7g4bmH
/Yf90gqS3MdBi/R0XmzO1o+xWcbL4rUTiooNicv3Gq0FqBVqsdvWuBEt19qh1d+X0YPukLkcgEil
NlKMYphXkXZwdwT0HonPVKw+xTrQz8AQk+AwjQNCOo/tiWCuR2oOvm9sFyRHoNKLC47wCVuUkxJK
9jqAiX1fU5BJyA4f2rw8alHBA3lvhbXBjkLLCnQJwldQ2iHtNXuqmfGzwFojyh01iwXlDUwyCsnu
spxDopRfVzEXVTLul2Jb68S9fmGeat8HvAx2d1l5xQBdbj72DOhlvmCWHskAOI9sRVLw6xHHFGay
Nm5W0M+R9+crB1evP16eeu1XEmXhrLxp80z0hPMqD48PC59/KHc4L8aJ+GVh2KfCtgiEwWgt6ZH9
6J9LN6GgofFZkVBTrQlkH/TJKcqly/ZIesrQWEDLgZByAYX/4UhZxEUxTeDKwWO+H1lorOrsEECI
ClkHLAQwLwCWYrTLgG7/HMMsVHNz0SPG1n1iAS2ZeCbtF0LVP1JrcXv0B1fOucY+jdT65nDZTM8n
LHER8QA9DSdwFJhpgAztbVv4YCxeX3KOzIFopFEZ0zH/sIGX3eCmF8eyHB+xhvRkPmNQywjyTHSO
NW453FeDzELnwB2MVQ7heq6y7kt09uZpDE/jAU2I/cjsKyycoAUgEpWyP8BSCAIfIuQr+N5inL21
Vjxu0BMuPCp311jxka3XUlzJGbeIz1hp+Rw0ggnNkBs6iuiMf/7e19sp+HqhVd994cXZB4HyihTm
q978EFVhmxO5lYseWeINUmO+NBStmdeOn4RpTDpicWIF9vvTL/24b1v6JsHBXZ8sFWW5N1t4GwAX
rIkWIYsWoNz9oWU+ON28U2yYIrWkYxz2sLo91mc/EHBC4jlE+dK/cQqCsb3FaTH2LvkpfnGUtkJ0
uak4ImoYnRN9rO/LktPVqT3Nh0rT3TJG352Nfk62Mr1n2v4BTQQmOviM8BGbjiwku6xmeoY3LTNo
2NvbbQb2o6Wz165mU5YnuU48D7bNdp1qxcTqCDhX88oePfHl699DuQiVVVy5JzVHv9gtsDv/kiGS
lLT2ALmKj4HKFeekKsFPcNbcXa2m1ckuD1V2GerW15eQRobeKTcGr709HTkZsINSOHWKXPry7GbW
3fjeI+CECPBqIS7VQSnCSAxjTcnVxlyPQx/qjQwt2+p2IImlj805K92R6egzfliSUIxYCTgSIMdm
kBALUcGyIUjd3kSuXk2EAEcqCVrNaLluzYcRh4HZTtEl40cvI26Fm94DMB1ZxlmDetmCJh+8tanR
xRT+yGbr7C2nGay3Qp8e4Ievuft/IM/oEtkLVPpSLzSw3QDgIeFTjbDh07X5raxZt5M2G88WHOos
DriGPfSnSO0gqOhQC91I1vxlLLfpRpmeuVxwRs0sVs4avUP337irZLIs1+omrWQACGD4XyCYVnC1
FtHWiw2qlTifLax6Jd6TaVi/CAWkBKDIoMn1cpQAjOEe1JHzfAosLC5QHBPd8X0mpVeq2hVIc883
aqdamJQX11MIFNNjJDDdpB/MlN+J3AxRc6HOFOIufRlODnwotDJCIR2QRK37SfJ3cxgAJUQkNIsh
JGJM2T+GSzfvtHG2hetJmbkzaxNqclxxik3fVwkge1Sms+4F9cIPY/0gxOLWs/Cu8tzigOBT+k+A
dz7YhbmwvDL2wk0wuwIbExf4QJU0c5UqCpmsSWAU2DhCo9XE1fblLLO0syW6JI6F+WcZvXCv5zgs
a5UPgAt3U72GguUacyci5NWUsVjdBSHKd58yZkrcBYoKJSFg4sPwd5mFAH5+hacclpnL5EKp+wSa
MMY4Y+wYVblAtQINIG1M4lw8VvaEIFFM3pdOwDWFkuwwMreBSuzOhoYViRsTwJ22bpZ6DB/IRlPh
rIR+o9RwMwjFnAzSz6POY0kC3t4u2B69ulVviZu920e+93WgAAdID97qNR8sAdbUz4Ynh7/yTWHh
CgsllXGPXZoldQ9lMIQM/kO48SvxigtUeqQBEp5Sln8lohHo8vV791RW69YdzCedElYou4RydmXS
xaWzJhhRL/d1+0vjW9aGDeNklIsGlCG1PByMA4hnHVg5hB/EAAN2cFyJz26GrlHtqsMeoUv/u01n
R1/KRUOqM8gvGR/9AN+pUYs3o5BeHiPHJyIVGQf+ZpksAOXsv7CF/6yxE4eavIrpOUGO1Kn7LRdE
6+M2OiCPOvn4PurfST8WAALVL4ENPRcUvsoRPdg8qA3gmuKf7pJxEOGt5w9evegNcXy49FxNyCBy
1H1ZmxOPU9V9WICZMBYz2aPkKGoow5UYy2HG2O5fj1Avk4g4hibBpwkModZnE5HnSCom5w6s4LmO
nhpeEzw2dengiocFbXjiojUu/0EgtgElX0a5kn/FJ7frQLc8hSoni9K1CeTQNnLjHzaLukfG1sZM
UZ/lsTl3sqHbG1gKf8iasMqMpdaFjtGrHPkm+1mjvrisAM680kmkiT2x2qg1AiqnYeh92xPFUtc6
XK/ZuuOtTW5hhlbNVvoCvjE97YrRG4foAf8aqqabMMuKU+5FRcXPcmvmYWtX/kyIr7FA/Xv5vLiz
CNm36U1LHHJ1dcRQeN7Erj2xWP8Kwy6nrOsWpPltBeRWKCMlJdlA7oYPZ04+MuCkzDLM7+3QgvX0
YFFTQ3WbZk3fYDoXMHpzVgXto/w5zEPzmYwyknvLJMqxspfhOzXiDtc3/WK1KOd/s2OCrLhGesx7
hQwTPa/Xtw7ti17BVLz+aR3mqM930+aaQB73Lp85jR6lxAkk1iYt9aShxcpqeMstLJ7zx9YVDBt4
hYhGuIaKgHfSkAelRkRIpN2h/nJfH9d8O+5ghKX7ar3w0o9DfE04rcS4sptYpevZbTjqUrVHRU7k
+nt37q+YgzG3I7Q9ZrYCB35IrxtPT/q6Xkg2L5gqX42LSdnjXUPe2LqEK+aEXZbXHEKlPEz6/3fO
0byyDblXHprj9Q6xY3q9zYWrUIgq+Q9OOjhdMGgWHGEtwekZ1f8SpWAWsP7P65P+6Wrt8hRvJDg/
icfEf+HO8MHun5tu/M80ZJBpy9f5jleKh+AEB7T+e/8D0F0Ih7mbN74PpuZup8V/0lv/YrC/sxeV
wuTGyEBJ6dQGof5qdRKbEDcg8bTA5uM4lIlXLO+A4NIzTsYsxK3sK6aRsOBDk7nGNc1ulUxHjobP
PGTUB+eFsB1l97xzix6mIh6f2YkdmtHGwfC04aWODUaXZJJu1MyrocOCDLWrlYugJqJ1SFoHGfVa
rEv1/SJvvhp+Zxp+QkkOQ8UW5oLA8bqbgN2bn1Bfks3IjEpsDs/lb1UTKu8ZNODu36kiI7Wt9MNq
REW5p4e5FVGQYsPLpId/D+NN9HFASJA5l9xNoyGy4hBzWjh7sBqIRk4AOn/vho0JJDfbvI81Nsny
f21j12mOmV03+N97Eb4k125gZEUeJ3hHpgoMdt/GpFTOzFDEN6xIff6lYHnh1mlrFiJQPoNukugS
y4i90kfl/R94ar9WV4iAM9UgUmZfIw25nWH+pY7ykewuHPMaKNC1yzHEtYDtxDbvMHvUcreG4Mp+
W/7sXcIhbAG9o8fqnUeIyyiyeFssYGMtjeRyvhIhNwz/ClPNWqQRvycXBFn1rwpxCic+jYkJtJDw
NhDzWLmZ3KxCTdh5tiYF/t5VRukNVtz9q7JaIhnGwK8KD5tXdc6Ou9Ean6A1zg0LgXwcIPVLUIrs
uJ7sdaBJMs1fn0ZXhSwXrJB58CugUD742hQDQ0A4HuAcqWj4TsLni3ERzkXDmOxm0emL+Vj+t8Ft
UNoCqZ1OTdupFSqRUILgDH2EtXzyqmh/tsMKuKC4eAP7gx7twXWRuFBNdQT9hGlDyU2nWlxEg8ZW
y0zcfu16c5YBtYHHal+6hzK/0fHXFXUkVogFoUbSaP6D67H8ZYVOsUDxgmyfkYfSZ+V/phJzFV8a
HXEE5b95kZp33M7IlmYvfKXbKA0IxUBZV02OXMaZ0euRNRY+fAxTxNw422ztImEi2BKJU3G3IsrI
QLKSIMuZRGTZcj30Xkeevb1WsAQsFIq9Fqe1XMKFTNnbYUQ/O7Xr3IFPuIv46UX9BdAb6j1YAQBN
HztbLHd2NhSCjeAGSBeste79WUgaFZFvugE3vyO9xmaoa2yyE46d4VzPrQk26mrXrCJYHZPuedzE
ppIK3j7BuiIPEjalLb2KXCEbOTHb4ZdPV009Bu1R8a8rmwcxNjRIMr8L2HTUy8JIboJrplFGjYR/
6zkTgMRXrmNu+kD+Gua0dBv23u3nVVd1KJ2o+/hDsUSlQFjyW13z1iSRux8zvx12nIe1FEzozuD+
vMNcsY/IXxIHPE5JPsUQ07/9b6Unyo94SRCnsCZXWfGSP3/qrMQOBlf77gUQhLogN7y+w6mj/m9Y
gPyM754xvrmd+C007UseEn2SiZrfj7Y4r3aDEfq/Fy8GJLpQDdRKaDiSep1mkm6ozQQ3213cLlan
ZJbUelGu+06WHisBNnrRBpZoFCHrRHRlzj4SQRyHH+ymKo2bFQ0uwpFj4kZnY/h5Yx++tHAvRHwi
CAy28tAQ9Q3OEonPNtr15etZis6kYbuQPZZ3my/5qWxEkNa0oembv1ppOH8oIg20dKYerrRYsKGo
x+9xeHVB5PnwKzKfqm3zKSEH4AaH+L4XUt8b+F6jcjcCDcHq4M0VKDjlF0f+GofH8kkS0FTTob2l
zZMGdYjlFlBS463ElY+wvS8gLOMEWr6CmayY24aFECu08/3MkSNhs/2tS/9juGe/D5Uz/n1XgUWN
1CCIJUyaFoZkHqWvJyDpQabhU9qNrIn44e87Lkhf9CSnwuQuSAE40pP7MP70kndix3/36YCUCi4D
6IiPJg0bXTuII+OCWn2qC4AmpfTwpuIkP8QgXVvI3bvvJao0VtGrQZoq0a1bMBxkeVFJUvdiE8Hk
j+eUe5fH/EwhSQNAA7Hm2AzlJmey9GS9eDbL+v0SkJPcSHvo51NBLJq4Uqiw7wdYbfkjaprBFiVE
iQ0RUSgyL3FWY58m4rialNzQEMVT7xh6OZA/R0fezCuxZ9JbfStJ6IonPjzikW8JaWK5QH3N9iP6
a9QbP68z3C15gER2ZwFvuvdGBJlkDOrl03ISEorCQJIptM8RyUNAIPJpIenFNoM3JGXQWocw0jdu
1zyhq6XCeL+V/4VZk8Uo0QiIp+3kjR2ybmskvYblXcaybkSp/UdvyI/rSuWMtfe9Ld07yqxBa+v9
u4krSx0/5/z/WYR75M0eeCFScjA2uVccNtPw4gHjN2uuNdISYQp9KP6FtRXKRfkH+QFTLpmNuCF1
wHIGLP/0Hph43rbJwtRvDgeVjf6L9E8plWuARFYH7Tz5vezZ1BRkxvLgY3Uv/9HyU73HgandzAAM
ULEswQ7ZDGwYO4hIgrLCFIGByNbRdGKWkY5oyItG8PzySmGwdpOHhNL7Yf802H672uhRhDM7QPi5
OF/xhiLlrZ51wqaqMjdct6i36miKrSbZtNhesLKn7ldmd1Y8kpWLv9VsevNXLJePA2yh34F4ogDJ
fLZlyzWiA71GPX7KlYdRwFo9GuPYnabtOhJAVKGJGzgdCq7N/FugMLB+WRQNp7Z9LgkVBdsgjlTe
zkqO80RC1e3xqcik5n+mcCA5BYbvOfQM/qm9K67jwTFBFAUMxJr92IwIIc66sCv1WzWG+JPxJyZZ
Z3O07ajZzEGT1JFuAUmffWeBXX6m6uQQIUxce1ma5YCvg3LnOVWsOdrNe2i2AK4nHieoFYUyJlCn
hlJjQmJO6Z3zHAsl9tsL48ND3nZrZBpFG8XCr5k/P9TyTi82f628urANRFWk/1dDWgi2SUPoCTW3
AeGiHMao7lphrA2W1FTI9UznuC1SNeaYS1zcVIZfxUw10V4oR1qXrqNGnoJVNswOn/fnSb9qzT0w
bgzKcEC/A/oBA4js57EzMHt++JzvIgkoZm0XhDJePncjhNqfSPM76QQQH+VhFco06SMYWKVSUOXr
/zgn4hyoqTD/ZRbnk1DKQmFTMr3K6wE3A2yLGjO1umZ1JrF1S4KyDdXj40qIVNxngK89kDDorwJ8
WcqXco6j1zuOT8SzFOYb3LaMacmBM2nNeRcYn/SDiD9TijeZTVq72p5fOaB2AXLIQ95p5kudv5qa
rZRyl70F+cRKxlTBIfIU9BRmAQ4k7ZmYJFrSHsoHFpHbf6k/Nm55jh4FRm0p4iPQR3NINAklKLcd
tL9kb4CmfQteUXa/p/w8FIt+ueVyqXrDFSBEoMe/sLgiUCtgGnyoxWn0fAfJQBD0yMGl9kCw3T5c
e+Oo5ZjvEPOByTnyPR6r+cjxQ8Aq6kL2vjrFLu23emeAi0nkxKYkJQD3JIuBe+WltLeWKPEUTFyE
isNZTvwySREr8OUa26LJccSGkLjoleg1NFSRuFw9XF6A5KlXrUlqhFrNpVc2WYq9E/hChtFjXMGn
U34Xk831Wfn05E+WUuqrmTTBe1g3ShwrfT9RYIxDw3KcBfkprA3C7myfjXEFzRFJbgozAYMH32Hm
3pT2enqCb5VeOChzPUZApJZ+T9gLrzFG1+1M3OV7uxpVnsThL0wKUZV7nQAScOMyFEGp3W3ipNxX
GO2vI5SX1/JEjbCR4sZWjAqLDnZwO39M/o5osFxlNyKpV9HaHy/45KoT5X7uSNA5/uiu/SNbjcxL
V43Q3RmRgZTnhVDPYPQsdQBGg2XzbC0wlpOPV0uIW8jIRB/vSrsLMiKtV+jAHMxSD4B/TYqPjRsE
0UgCq/Tf4C8PNDy6iSDlgRAmT2CFtx1vDGs0cHVPiCsuPvDuahi3r0ITdvijjCSzJ+/q7UpTLiVC
ex8upSfTqvYKwFC0ZVaDXI27tGsHYsfqPPiszqNfTuSDDFmP41AsDeVu+Mdbyht4oyF6zAeteRFf
yW14WYZyuLso6nxBl7POaAU9MeTrIrOyDUgOIzcxSYpvONz9jKWqN+hPHyufuU7KzvFcDipTZ6VC
y2TWtvMX33/Ar6mzwkQ4pVOX5frGWzXSbIXfuyusgb0Le1XACBCH+13KZjQZXpzGUqDGIsFIjzOT
BHNbbXwzC96z/9svVxUvS7l/aSaxu2OS0YvfPLNE5wctrggd4vpjoPIvM3yMV4eibfX2Wkdsg8SJ
vuwxMeyhB7QGzU1NN9clB9cZw+ZPxvG+tV9AwyOva05tFbrGrJ7p39EnmTYLv00i9B6PZb0Y/4Vt
pmdqTacbGBedx8ormkzQ5Yn8MGHUe9COAWSP1zdk/Cf5uBH3cFOnTJtkCG0ZDkO2r9W2AOKIVstW
Bo5pf5CIYYtZmm6nTkSesJM7kIa+f3uc5CI+8Gnz5ptJddi3LMyE7bSR4A5fyn/VL1qpy3P7g/2K
uhRt0oW5NFnFcNyMrwSy/f0vOOgirhf/UK884mA34QMPJFTV4Kj0OeZ2uIafRyWhuFewwg6yDGOe
HVSY0sQ0gmFyHgx1l9A83xRwP3uF5ZoRQwzeypj8nX2moSqaWFhc2u3YUvx6OFV3GnEXjyb5cpZa
aDWnG0MRDcYuFnun19VrFb91ZnhxxFTIRjuSD4tmnFgrDqN3HmjmidyjeJlhc5VdO3sjF7m/q14X
3hn+/HODWEnWYjjWbHG+1zbgktnqvaAbzRq3E9x181j3iQtt2VtjM7H6azg6oYXtXfhtjHe5BsSd
UTysmlgYPxAogUcXKG4WN5BoBGIMDTO+Vr31oKhF0AEOQhINYWemVrVHGlEzaZk7YfWtkbK7DQ5+
UKdNK6yVcGk7/yPQufIM2fRc7h1QhQmzV4cL7iPSVbdQ/oGiNvhX1rriodK1jZ5PQW+3PxarGO42
K1zP7/TvF3sIJBfgao4Uq30c3zrxScMYnU06njGvHmTwYZ6Y4zVdfh4JjaKrMTQeifyJFkOxG1Vv
w9ShWdmDfXlXrH8HDzbYzKdgeOH8Yczditi8FH/YY2kOOLqeW9oSgBLkXj96C+P3ESNlK0BqrXjE
SSFfvTIUD2bvBX/k6nZTnxppqZZA+Oz19tWXhF0aIcW9yy12t9F+vrLjWXoMwXSYbXDrgr5jej58
GuZ9MKwiixL+kd61s/2MKxoQH0eI3l9JhE9M/MBNvXfGHM5BUTDdiV8mV1u62dDm14LHqw3PUMNt
zL/uxic6GRVyh0PYhVo6YGvvQwjGVmiMKFfvvELcNj1KEgqcyvCJvjGQh+RhXKJniAXn37Fekrw+
PjlLUh5Tib4yhesUuRB6dpJ8ymNgDPQqbmYtzDQeb4r1OAR1yAk4c5+ROHwkbZzaTMSpa7ksHHja
vQrHuY/6oQCBYGEQIuh5uJ6ulgjw7FuiVE7UztOEBR6fY8H/ENGcHlRv3XJq/uHzLEaIMuhLRlWv
m4oWbRXouE2Q1oV7OVFF3Pxc42KH7ucLKBqOGcbFsA4O/q3Agdz2fSnibZ7+iCcNGYnogf865Io/
50tS3VuT2n7JKYgwV04lfUElQPwIfq/bFzAdiTHQ1k3k5Zl9nLOwt3rzX5gvP1MV2Ycih+l7uia6
94iJkKH2P9qJN650LK8Fe0ZKyKy12LoUC1g9dprt+baBVpwqbc9Gg5o4/0WxZKXmD/m+LnxuCz+j
UYiIkZUW0rWopsnTiNH6j4cu6jb7m93OK9tH+QNLaTKjLvh1nnmfMRHEl7H4iPCtjc+6EZvi6OMN
+xZO84Ri8C16GqTnEwaNR6mcWbWduX0i8rYCmBRSVA1stdvSLpR8Wn8ABsa8NR2Ac+prdCAFbWJp
ncMBQ982Cy9sattiwiZBp4HpEwlsbFnzmj7yT9xPJjT+N3/H66fr1vyog+nKoJHQKFehfH7sA2Hp
VvCb3WaYoGNxXgFpMepdcgIb8b07Ka/mkNhcJoKYwtDSh7rH9E3T64RM57pgfdMBlQ5qMQv78IYJ
hUqyfiMTtdswjmLDHBltzBYyB5qj85bf2129q/E9LXptI4AsGO2TGgiV9SUOeVCYvIUx8G9+b8xp
5L2CBhkmBNDwmill0dNXlxuTo8c/nnTiHrAdBPrcFsNUJCT8iFSG9ngcAImnj6q2EBTIem54aEuP
OLxZ2B6Ggm7eaRsd8sWnD47tdoB/49O3VcH72QYi9KBTHXWaOkM8tbtshLGI14nQgi2U3kkXw8Tl
Kw1S+XlmF0S/CnBTDEUMSINV6lCRbyFUEsiB6dh6rapVzsZqr/Y5jj93dEtDnSZj2S/bOKPkL3Oe
OIMc09bud6O3FhulG7iGxuoB1DcTPLKlTZ4tZToeCua/Xc129r4SlYgs+OxDaqLO9kv53yOmSOsh
BCdUNQXhpbBHoCiuT3tHQDzv3zGnKFw4DBYV0jjw/JydWhH01P4dZJWVlEP1u1OVjMCKschbjuNl
ra+5tp1vvEktde0nR+sxZsfMQy4ZsHkAPIbN+Pxm7eY6JaRwiBuDgxF4k05s95hFbc1goouHh9+g
GU91pOwOO+lVixPvkZP74Eo0U++bvVifXFEHyY+mYchBZq2hZoeA/YGludXA389lryg8NQIqDBGm
JQzgwYIc2Y8UhamB9KHPPM00KcyVcWxHz9hmJG3rtOhDYJ3uo/ktTF8c3nX2B6uQW/ZdyY+TASY5
v22Hu56zIXxemZn+ZmcCpIU5KzVSKFhDvpBY/p8WK2dTmemu43FRcWwha+MhxsrpWQ2FtgcajHq7
V2bDwa/Ckjni0GbdKgFBvt28iTNVRPhROJks9f19ow9bojQoorXBgigXwkg0N7mO+WbdWrZGVm5f
JuCgeuibzaRvSbq695fUfUjPx54xDQzctiThGrGZdtBkin6i1P8/pqCcUZ1SmErwK4nuftQLhm5W
DMx88nwaNjDVj2tm/R44Fd45JjNMstYqdUcRQ50KkcmGxlYtje2o5gAsbjXsVedUR7oeaHliXQ0a
n3nWhV8UOwNSgbxuCagsua+o3qPZ6SyWpAXgFcsV0/lz4qBeb5XNVntE/3F7NN5icjttFmGzBrpo
PCo1krrUHB6nk0p8Mh+eF9KjcZvHfe/7IfoJfZLhUJGNqL8w3c0JUWUBJts0Qk1yVyj+IPZcNWvd
Wm3u3NGkPE4iz/kBHeMXGs6HmjJQErUj5eechRMW4+3+mswbC37A9Tth3cHCehiWaKZJX1cF9rXg
wrUengMSDEVectXGnG0tQmmbhtMTiy5e/mMCmMuRMq4iF6d60xUwcu4cQ+HQ/BMoWFPyAnPIn9KI
Gm7fowTaDssxb2zKriVdkTuXg9Zblk6XxZuG18n8fUjLdO3Hol9Ap6HcDDW6J9l72oll2kH+4Vvb
abFESJ1h09yeIjknOsx3mhu+PfS7K9VOJKIf9ELhrinIF6LG8mwgYkERapRaIYcAvE9I3Se4AcvE
1IwCufOsmASHdvC5bzq1vF9AiexnXAuhQ/sZfHNJ96pvhHQvoi/jeDapud1SK4wH82gFqP6TEEop
cB4PksPz2T5BSrnNA0e7JcO9DoVpMDmM15wmdoAFYzUB2h7ubooH7OFCmnrTh6DoKPh0XjEtPqrB
gMLSFSBtSAhalTPPFrG7Asg+Mp+m2TlJ03XODxKA0GzNO7b1LkVuQ7lOlTIM+Mh4eanLsBZEAGNc
K0FySman2rCrIhzLs7BT2SbeqGER1cADTxayBMFBX8zY4sEpSRiwN7Kc8V8zYYviMO+oYJfgA9aO
m72MgAcmD69uiv7ZHM+ffXL4LpD7vBGnKR7emSkwnyFV3/Yusrgrf9O0uyP3VTYIZsTVAn7H5+PJ
u+MuaoSI3/gwsa7Q5aM7sl1nVgjAgpt6G9MEdUVUMbes4N8tQmBwlabsD7DrGbBO7eXszKtgjHV4
UP3FZQ8AsVuF6zii3rO6QM2aoebxmtUhx0mCRmnl+xR2xWuF3CZt/4Yo3Ckql9v8k5hjbTW4IdwQ
JSlAtK4q3OGkkEPWn6SAeZZ5sgCqpascEC6ZEKe7ki1+HpyG7TsFhoPPYbZH3QqULCz4i7FJ27U7
WUpSBH/KKLF8DY8TnKHGYRV9XiLRFcOwOrVIajvj1U+Zqplezxp5neCTs8jdEtlxQYAI0Pu+kNkC
azc9wAQGcRGM7VysfyWXZgYZVJ0te0Vy5jHxxsb5S63ABwC2Cyhbjsinys3yRyIL1ogWizzjMLCh
w+B2RvzKqH0jS8qnIbLyt8ij7A/VUGpzPCvBuLvzgsJvGve0/s2kbmk2sWoT/J9j4vzxA8Cmlt9g
OFmGAkx2lEJEWRdaICXqO5rABFHGEWUGtq+bY7nXL4oYcnRaLn49TBnNHIIWm4t+ivYo4VkMPFIx
ldZnsPBIod+MmbX4TG/VShb13fPcHkAAMh3+eleo69oQyDqcq1suekrqblsyidMBPg6LFMYFTNkM
1Zas0CKiuT/57sD3/M6+73adGwoq0yXEJ9lqc0WAS3qk0aD+F35NxIu18HPBDMXfUiae44FpUgsK
qw8fR/1agcvRARhm81cwPqMBNicCjTVRH4nm4qIocSDV61TaaSONmG7jH3JVrrpAeiblB92W03eA
Z0HlaZhH4J3WU8q3hdcoktUYPCrPN6/fuTT4RnBh5Dn3G/PF0qbDg/aWkfjTIfVxGhmi3Bi3AVgX
IYTbNp5k6q9KcUIuww3N3gEWjbmaDBGwAEeUZYRMK4fodCCj6lzScVvVhXew7XGi7iPZl4GFTzqZ
/3DUTT/0NCzyAjF4su0g0dztorKgJAcoLOrqko7mB+E4K2Rj73Kg+iNuhULMDv1FEiAQH40stfY1
JtbSOYhWnDbd0OpoGbD4Qa9qbBz1yhdsUJbkKeWTb5nyn3+V0iZLukd/k+dkrO2WEgHFBnKylowm
31DxanNzc7lAxA520sB6vs7KJ0YFO7hTIPPuwT13FxhJZ4UcXZYjfqVh6+i8RKIimol5Lqq7Nq4C
8o4vGuuWbw9Bdn5+EON3cgXRhpJMIuUvDRG/AuCcuLE3kXSRc9vVK+fm6IhDyXJ9v89MLAKVyc4m
jx/Hkle8fl6xPCTij6fanRovZI876NX+ZRWROqSvXO3WEJe7r3SbW8fjCNEWtlHkK9IUijUsERFO
nhwjmgGprEheLxIFZh+lW6UPzVll5p23O911aYF6T1cz/8l1Ohi6bbd9rcdkXzJlxoCXKVj/FfAJ
mY7aMFGTE5Wh8FZu9QUIAiCK46P9JY2bt23lw9fsXwbUocXmgwLUgg7XOdOu+yXpBJC0np1lz03k
/LT5khTmKCC03cYQeSk9iQLKZ+VPHmmOFSJHtJuzIfRcp/iFca207eNyLaORgJMytcl8A4rSUXGa
jBiFB5ToNvzuFqqwcWhDkU30311Q5klkvPnuegRSOlUBbHsbg2kWNUxEomBbx/K/+Qujqst6mLGb
RCKlmcRt2VlVzfZd/8tMwJqWk142nanBkKt9I8dVrtIgnZiY9aNSi6TZmhwU5jt6W2/dIHnTNpbV
P3H5SHL3uPFdMsRGY2TGvOnBm+hAoYgIpBwy0cx8teJoqkuav0upNtiwBUyM036bdxhG2yY0gP87
So+G0SGMe7bLYAEGxvdlcCANQOxqvqOJkKM+6FrROiGWrKCSHG4pW0wVy9ty+YetHhu+s3imHNbh
hB7Gq9pAPIbhhv8CY2JSrCXI1qCFiNakOVHwZCVmyYJepMgKImF/8EEbfb14nNbhW95S4rNdM5m5
FQSEQGfyHWzDvCMaJvH8gjVIEz5Fxa/pT+qIE740C3oluOScuRI4+XAtTAOFFbVW3S4muaMekiB7
lxzdJ8luux1C/KQ93GgdIP0UH5Fgkq/9U5vtoe5JZQkrDuYLQb2UCWOQpn0zY8DKflcZeKQ6ngUw
UYK4zkY/96BjpdK+PbmZWhWfhsMYoQVrStV+d6FM7hFtn8nP1pW+wPEbI4Y5PqTOSWhbHU25aVZo
Lu4dwtCXhLolVxWMqIUQeQrUIqJQ8X4+3VhXPbQdiqMHdLYHJ1FPgL1Kpu5tP/D9BT0BbnraegWM
rjA88++UntPRczgfDLSBrwj2LjW/jjpqJyv8YWGzN2wtwNKjsNX3DfQ9xQ/vQ/pzz5MUpoeQbONT
BYYpqojmkyU3ROkv+5ksTtjkhutIKEnknPHH4rFQstq564fSPQMdWuBL/aZqvkloT4wokuVClRHs
Cd7Ip1l3W0aaYqnla/+YrIzGvVjMePnSiozIIYJjkT4+9on0s4jcY8SVXeaYiV3LfCX1/483shtP
DyyJR8BQK5cvZrN6HjfEX6HPJ7NiVIo85EbBz7MNuMgvcvb9AuHSYeprMJ+O8jnKRZFHpWDSiQrf
LwVmOwGzzzflu71Lu2A4AIq1HDi0ybSx7EBK2hRlRjomDJ6sc/DvbvNaQYn0KylqcYLUhMQpHN/p
y+WSTAjTtd9nRjAjUegIVsHXsjjEHmsWof4pwmzRxjj0ZVkWXGKoQxlYUBuj+6Hjw5pAStJp0Rod
1iv+0XgdJmCe9O+rjO71qqs0ZGeoq8aklb0rNcwkSad/DPuOOTOJGntJWfDaEwzd/uRQm1mOdrlF
dw7q2CxeXRO3NrB1Bzf3oDZTatqmjvG3yh+9s2Yw36sPI/TaP/0izPFVAgSkqK9XAxtcS38pKBfx
Jwja0gc7rqtt0bYE2ctaHDQQBcdcRANkwNfLDz4hAkZrXLfOQur3S2skGypUcX7czPunE3R0lNos
k7lt1j/WoKhOBJwQy7cpd6+/FIA5YmHJ0EJ8CFsoye/rkpsB6BXd7Z53JAQJgSc2hljOGDrAXf3B
0X78LFiWzAsxXKVCwJxPxHonmKqbB/72b1KXwcnZqII+MxWkaTb8E/yrP/twDmLENKKCc7BxciLy
FDnMMMIE1HTrP2xIPwIbF1rylt1IE9yXCksOn/zVrTeETOiJGj0bt9DqJ6gXiTEMND0RNIowAtqu
b5ydzW7CiPwZLq//sChy7QMT1UTUqksmQnNCXrvI8TVLxd9O8tsu99JTfSYzFje+Y0acbJBlj6t/
EUkZoB1glhgbCPCMmH5yrp1bbhqB3qmOT+VwGQYLDZ9Iz0XSdzKlfek5uzg0jyUbXoU6N4Zqv0QK
0Wxw8EI/kBUbqROAlhJiukU/Ve29eV9MNB9BHwiP8FrgoraAxPsh+JPz6RDi97Y11j6/0Al4oTTU
jx/xyI0qPWrJRVNIDv1Vu7ye11gFk6eSgi9aERQEtUdM6Qvc3hJKCM8JznvY6EIvNpfAGdGCjBCB
4kdVzMsTG5M/w7lOVpNjXc5ZLeFtV5xrbfFDwpNBCkk18XWOkCmchwUPg06blEcpqk5zXwNuQoW4
kdVSKiPhNq++LMkEAUDVWsg9+T910EyKIHsp3JraYrMGDQ237lcP6T8Xyx8FuFezmxDMTYo9pW2W
kBmWrtB9aOuaYiXx8x/iYhPBV9gU90I6NBBICsT2zeg9QKnBwyG11nl47WOtxRNDjhpYgOxYuaIu
+DJZTPrnoCau7nrUD/sWFP93cKTTcjx4AS3GSAss0ttzuedvDWKExiUOKDF4wUhwMe8ux/5r25qS
l+L2q5WJUXwZhKxUpyNahhSJgxaX6qxZxBqFGCcS4FMjEZDiaMvWx1nyc1RiqhMzlgJJAddcoYbg
Mgw516ceXEJ5/t+K8c0+2l32HBPemAvurRKl4RyYjg6pW4WCXy3Pe0IsPNla/ziyc4W+O029pigA
5bdE9NhhJBYzdvEKwa1S32sKhFfzd4jPCR14iktValCvqSKSoevQZwEPea1UWIdcQYOopTdczElt
a4SilHu8IGLfyKgUeqHL2+nF0wUO1+EavfhU/hoibxGcRva0XwkJzS1BrM5oJ/l64Livwpe4+jzl
oC0smyDGmjDC1l4ruPATxQZzuDXpZtJbFUAFzX/GfL68E5mopD2WY79J18wODUq0JM3n7a1sr+7m
A5Q06UTM6BwQcEBDo6Cl8KyIRfMSjFVtzK/D9UJeTRyoRq7dggtRZWPUI7ms5iW4rBPhf4sSlUlt
Et0hrU1NEDDg1oSdOVldr3ZflbfDUaGvhpbYFiekED/ICD+zdcPASJGTRjv9qaWXoy0+mhf0OknN
4nx5ST2Q+NXo6Jb3ZEOVLfCvdC01e9zklRQ/4I/jHq95oFHx/RAzv73fm3ghodXUOA/5uNgWCuoO
7bTfLK+DYZa2I92B4X5QWXlyawMLKpCkWpGBRZpjhEAqCB7IAtJYL8W97MUHcPy8dea/RRnVQmtN
nQqUiuUNR+CSQoFcTb+raB8yI16mtl9ZiA0YeWvuRdPXLaodTYMEqCRXEP1WKsHR4QJFS5ztBuoE
RYoFHDCTSwTSOXbSlcdI4SC5egSJyzO00ungVt2Ukm0wxm5KC5GPVBrCuJf/RKm18u04nlh6uruv
zSw51N0YdJscWqhhYjt+5J5w6sX9aSi5kiI1sIjULxhJO0IRFhIx1v83g0+lakIZXSRra1cHGX88
kq/IBXQYyD9/kO1aLXnVFfaBWNcu/8y7Bh3j6LLSW6vmtQc3Hk9E/w8ADjHfTsV6kOd0Ct1y1/L0
lJM9Ckef3pKiRDOytmNph6/qfyNgaorCYAe+VRwLuc/zyd3gcYkCtOz0oFutVnkYdDoOojgKZj6d
C7hKvkfduvGWcWC4L9F5DHJy+rmvySPJ0ac/Y44DisH20B7h6ZTXimGrQfC6BGrw2oUe/I5k98m9
1DaKTsNyr/FiyWyLmDhTMiyrJ2bgHc3uvHGyorXR1HzQ52LBbGK1dOfSfs/5CN6nsJY4ET8QsZTV
fw6wv+kUo2rtIiDnmrEVFRi7ESP7Zn+Qf6gwNAYZIRWvfkPdZN4FIWAenUOLiSr8WenTa7FgfeWu
+FBLYIUIWM3JyY/bCe9uzSbpRQjdeJaclAlEqgWRwADgba9CQorRNt1LPSUCSedCkwTbd8zMB9w2
4WVLDPEVGb1XGTmegCmiWuIIihm9w8nHGvKVa4NuD4dPXUkivwaN9etmutxS/96G7py+FqRBFyMW
KyTZTMcm2IMDTQdGEx95dShD+DvYAPs454nCNdHY7oXjnGaXA0eTE/HoMewReA0sBljXPKmvpet8
tUCUh+yrNZIpcVVR1+5tAcXcSiI+UKWKrrE0AtTblv9MPhqBQ6LSbbhB0x5kuYh9ClKpj+6hSw4l
hcSm9z80264fg4wtdoFwfgFITrzO9iWuo3gHJgjtifLPTxrFr13zlH2KbIYkEuygKZ6MZd+QzxNt
u9myj2O6QnCLOSBhZdwiB+73HhCXIPc8hRFgjpdyVSKHXjZTyu/69OEPB9GflSZZrchH5tYrRvCJ
/8MNY6IrJ1cIjLyYhNlwLXsQbur1n1cv+0MRTEd0rPTBvTZHhNslZ6JMLiNm5AKXYhJW1Y1VYlOt
sSt6SQGI2xx2vJhoSHwPwsPYnn1zGmc08UBv6s+ow3N5/1TO20zFiMtEux4YhgDQphUOmJsiaH7c
QzWp5YrjCgfV0yaFN5IcqZ37jgtuntsjfyPqL98H3kQ7yCmnT8RYjHq1bN49hovBOohXZb2SxNyT
2ujhPsrREG3groipg7FjtheXOT6kwbSRqxx5RzwWrQDZ3X7y5rg0X4dn1xyRXn/5g+kHhTmlNxw1
6Mw/3di6SCjZ6d9Rr8hiw6U6f79mV69gFrMhESoejakorApJPF7YVG24azCWXNnVLYQeneNKrWRp
itsz9sqax3uko/3OAKVFWpHyxXArgiaM9fhGVVrzH0rYB4p255BJCLfgmAlJjzUX1Q8IcgbSCo48
TlQFuS4bdhuQN1pko+72fmUQ5sl73SQ9T3rk7yemQV0oOFtMaW+6+QDolc5f3JeRB/SjBfgp9X3w
huDvyBgs2RM7Y5qZpq/HEithETYxtI0oIupG6uPyhoVoRmTyZwDXJsWCliuocrV59NBU8ILyZkgK
ZSKsj/dz/YoqJOhdjAABY1uvPu9dRWR7fCMG6aDvcFVeEvqj0yP5b13Xa9Q1KCA1ZoMaM5H74ptw
CCrvYvu0NMA660LOyiEyK5Epb53apVl9r7/OUSKzZeyjARR3IE9n09EMEuo15/2kiaw9FHzajP8S
j0FGPknb+vyU5KVf55HjDSu6zBTzD4EEkxrnNYDSDkdwSaZidp0m7rVfBvyvgbuP1sFu8aG27+Gn
CMQmj82CDy/RTlFtN8DJ3Qx0yCyeVklsMeao9yjkWKSwLYgL+DmxkuBUQ4gb5deiBXnjqc4tv5RY
srlWOZg5MPuk9kuy4DPbduAoQHwtJetZ3y2KpbV7tbe2c8UbnnMvfGqxeemwNsEP5IypKOcpN9Dz
6PVjurPZrQNK8q25iysSecALQBXAMJZmqPWEPm+oEy3kfhIQAkLQugiWARhj0V+oLzpGu78Gqy/c
PgmccWWgT2LuP+22il2WuTM3a313aQompilSsbjZ9i03ITXO+3N9KbJLTva3WEhvrOqZe1WqbV56
w5JKYgpqCweMZ4TSpAvoePvSmvgOO6A16o1c5yhr1Qkz+aWZMl9mG/w9mlF+UviWwv2BABcbhymX
kyzlbU046/75Dh7VliK8l3W0TUea8AiF57aGlK+roXWVUxtJ1gk7tsFccraL9IikoQUe7YN2wDSU
W7tusrxJ3tjNMtgWe83kXiKEtW3H56kMcp5NfEZV9b5aNZtPzJRnj4XRv7mpGhQHdNVzpCTAJRoy
RCpRArKNsKW6Xx0DtpcmNaWu95Md3JoKByXewFZK80RDBiyUHOXSbm+h7Kht1AS63T21wcX7Fg/+
YJ1n/xaX61Od8drnjufk/G8VIIY5/H5D5yiMyf1xvtmX+8EdBW5iOHDnVsRceFjsp0f52E7HZGvZ
9wAGRi/CAtJosHKhS+nNUofYhfUwUsl17hxpBhBcGWvEaYfsRPF7iHFeUq4awfw/gN12Qu8lwJAq
8hz47zBJ8jlIMiLNmZO91tWIKP+5aKs7LXf+rj4I7AJlD3POa/1Aoo8Ix1KMMqhNqvN5IOzvCgdF
Idp3FO2cHBWqBbFQUPxThS2QfqRCDW4KcpJd/h1XXBtkGjbjcSP6m9Jd2WW76QnyqioEc8moYV5u
91ZbeZZOvce2hhN+2jhicb4ezanN6r/88kDq8i/xN8gVTe/D12VfFRf0l6brUgGFfPYK3JC9cAdU
anbErxbFxWvp3lNenu2Jr2hUcLOcu10mblj9HTLz3QpAzUT353BFLRMXu3Jixq5tKjJoVU1ByZyZ
XSP7QW6Z7e2toWWwQHMD8hNWGJOQPN4F/xMhOwAvQFbqxaXP737hNgHnNkIDVEmnJlrgY6w51O+C
MAdsRTWTlT/I3um+o3XTUzDOakLzoUBQTKa8ca4XnAXNnfCQCV70E0VP2H2KyEY2pmV/9G7U8Q+3
pwN9fdIUijB8LTazXVECi+tbhwkbIOTwLgJMveGlxsidI/6rsLwkzRLzksspNDDBnBqvSpktLwib
rUK1JVnason+jBawXrvDxBl9338mwAXB6TCMj7vDrleto8Qsx9fFje2+tpo5SX4Ou15JAbuTFdzs
zdIvIDPfv39QczHfU5kDidDDW/0h/yeJWu9S/oliifnOOlRj5EM5M74qCCbWo20zu9PoSgYyA0aY
DduJnNLxJJ9ez88IJ3Go0s7Yczp+rB9g6+2zrohPgFCr+VqgpIpA3FVSE4aifM9auy3gNIGJWJpa
WN7j9eCawSTJaeXDsqMTrnwu4QU7OeXviEkFhvatMFmnizta1xkVdLK18wSsl9POs66b1/BLv4sO
rUcqPaCHxcpHqvyfp3X5qg/lMKo2GCuuB2J4T90wUIv/kJEDf5eubAldLY2tnA5B1TPGru8T59ix
gUzKWe09F4YWsoSbnEzPWWpxANmSkkj5AF50X78WQHrKClAxmultafS1Bf2Ox/idEWZUcWi1h26X
LYNDCQwLPt4M0GsbqdPdFnOwwRtFAiQKr1BjMFfHH28V5H7ZaDyNtp2DhMcAmBFR9c2xVDh6Pxfv
r89xq1MsDuzUiT3RKaicCiInuWMhqX/nIUmEkxcUaKqUEG2ldsuU0Pb2YEW3e92czL5zcF0D6ALu
F8dDbt4mgASUwFPyIg2EQ8PrGqY5UQhajlheS+AOjaCP+7EVTSOaK2tIKUkGPEIH79PpJZnysLAa
WyMmaSdom3XsR/voN+BHk3W3i7dITJyzH2HehKSHMcDedl6F4lSmuDdqVwc6TSr2Io5wY8sXPJL+
DH+khV7EawSEiTPe/FVxRAstxAVhOesL0hAT/U21iuk+J+GhLzRXXGJQcpD2/6YkhgkO1Lhcg/qR
RJCzp0WQcWgvqItfzdyE8MHn5i8ev5WqzKwialpz7cKyILpNg6NjltzK+jtiuRHl0XFdrxIlwJPQ
Za4Bx4ktfTi4cBJAA1hk/UTeoohvsF2U0HTVD5KDXFD0UAnp3AfpNUKl3KZZpNlL0WH2msrPKh7n
NyuFno0dH3lMm5PPxEI3pRNsmuzny/xlosoYnPUTYIBiVQZ1NHBb1YA0i08HWiXRkJOKtLpIF5Iy
XIR3bfiCi5KqU2RITXlfuCMnU9lJOTzUWaC6SIHNqTV9tFa470pehfbvDV9R/aElXcT1aJ7W8gAs
+tU7J/lh48epFMGgGrb24/NqPEuYDR5uJG0/4PnkcrWZOBOYAuVdh3rrTCUYN05SdFNsdULbjLT2
wVWdz8PiQZ3a+ce8C2fR/3efb6W0KRPaXCLi+ksVW42y63Pe+5Uo8q1ZM5CmH34RIQFubCeSsF0J
20DfR0HRuV+N2cSuujaE4IXesTifHVhTXYXyQ6sCpTteQiXM1UtIl+nXzMpMWtSq/5CjCpEb47fw
U0t+V13dDnHdU/Mm+8cjDbCrJSTcAubc2j3JIhu+qqzqMc4LYLgTP1sxshU77pWpzo0AfKRz2BKt
UDg/PctZYZu0sQJGzZ2HhXZ1aBgh1IdInpn3Z/W8upoA6D4+pbbasqa+fMw8dq7UxNV+q1TpnQ+T
esa7imCOmK7+P6Zi34q0205xV2ECIupnNxFJLgBvqHpVozvEXeoi4VxuQjek2Lh/Kw5lbMVNTh2s
W4/b0V0iZSPYj+wBZQm/iy41uM9PYZY2STzJ5odQ54ABcOMvvK4tJj0urtOGMGtdb9zzlZFLGq2e
J23AUY/R0LiPS2xoXi1B1a3cO+DAJw4ujCO/3mWbUKi2T5cqM6mbVoxDViMDREwIPKB2lNlXy6wt
5CWiTXFKQA00GcZYYOtzdr+nfJ+86LPeAkeyKmwvu7g94sMYJwbuFr10HnqCF3O1glKmJWgmBvio
/ZrYr4ekdN+QSmN5PwFKrqIEHvWcq4jLLJUPHb/JWmShfzILZsTHwkw8wUtQ8l/YYSVolm2TZAOu
8T+1AZUBnWhQHrffLjUnRA72jJ5262sJnnQaeuJ57CunvwjveQYPTska++OW1l6WivFSG7A8WMMU
NglKgxuNxtL6bSLA3AvyH5L5de9bG/8f4vUEvnYT9wCs4MPA4dOQt+NMKPOKjIFSeJ/v+ZbRw3rV
9fnXcRh3IHjAy2p4ieu+gNA2kBss5t+qSZFR1dIjDt0vnhGWID6bN69xf9rlXozIvkmYj+5fDDrs
Mf1NaDTeHT3qG89Qq+O/cN78Ll7IotRVmwD4L30WxF0qq9H5x1+JPlJThW5fvJOKNLwUmJ0s7Uyq
mc/fHJjAYXNlrzz3L2/jGHQzG8G6SC/6YMTsGzIWY64l/HKB1QaVta+Tx6o2ygo0jLm7F/EQesLw
Rf3dVCaDbPE4tNJhKvrjs00rnaUvIgPfkTXWWFiuPMrXSmlDtvUP0EZubpqk6huhweqdmZk1+yvm
B07K5W7e5Kq8OWV8wAapJKkpHJVZcXjcMz8anmCi4OIGZdaZz3N81AuBWirmQUjKJOd81tp9wb10
4gojBlGwkm1b0YcJFRALk2uymdYJDIuJiyL4YABRt2FqkhIiSls/CUwHJlefxa1h7jF4Q99DfFgn
xZdOYdekzXp0t9wkcY69fbmDE/HzjIiTUkg1nmKGqiCKmXMN/k3DONc2LOPJkIfAg0f8v4FwMq58
LUu3Flhz6XP9WnUv7UIjsQxBIrWQm+ql09rgWYUsbr+JYvVw5R5TxsJrhvHHLi2+PVNFcuwozDZZ
zJnVQRQ2e3RAXrQMbQ4NBSTtSMAaDxI2Wo0ydluF/mDklK5nna2Mtohh2wjfb6JaZiPl6wr/Uvm5
zWOcyQb8uVHojW7cjmTEHTz/DFn7kS8AY286kimLPlJVvB4yHaLQ3YEF5BMUPP3295UT4GqKZ638
da76qx2MbY/LXKmXcKkH0zHHgRWR4XPssUePlRT/GFJx0hPNzPKceaKFlV726V8F9ldA501rq1Y1
f/R123V/4Eq6xYuCKW7lD+CKpX0D/7tu17HaWD4o3fHvnm4KRWkkMUipnPgiWh6dTe4TsvzVNoOo
hg0lqIvKsBQPPz1U5PXU2V6pqvueKfcpUGbVBzWZcdOR0FaVLV3iYDyH7wFW/d3/2gDErPh/2isD
LDJC0dU7/AALMkZgYJF10AmNggGtwR54L1wG77lDwHDyqEvGNPW5Gy9hiz9rRUxY5A5zB54XKtq7
nDZjCKgO+ZwtCIPMlA3G8Ww1zza0vo9Xzok1JvT3buCyODj+2gM0ZQS5G8r4LBZRCvwvWYdedbKJ
4OcE3iO2Qy0tV+prITnt33iTzPtKL7/aWqiZLvuTjOHRARbY+0d9loLUhst3pIKIN8AohXmADIiR
j5HGAgpnHGz6T5A+Le5Yq4PQ0oa6SgWvIQM80j0JgLaCk7z+ZfQ3pHfcPIrHxy0Ee/+0S4wWEi1m
/xwHtOVWB9NbaYwP9OPjAJ9ywel0gAKGNV5LMNxsyzhWgrmf73V+qxHGD765/2Lov2uqnAgA/Tom
tG9AVMBUQDR6wWQzVw81Hc2506MJI1PwF6V5DWnov9mPSEVmuwU3s5obGx1dFNkCKvvlNbOyfiVu
enBFVYuuu0L+eJAAfLhw/O3ADHaXbAgRXaWen55yiBFIZsQUBdpZPLFAEWzRkhMiz7+iJXV5ktOY
16jdxaP1zI8MFD+nOgndInV8mfOD1vPFxI2y+uIg+K40kIPtRlLT+nHK0RK+Ye55T2Ve4akGwCYi
Fok6S954jZWXgxdCJyWnZUGy0YkWiQA7WBzoBv+IfqSIZHCvwoszNGh2/aQmfAyWFJP+wjZfu8xk
x1hh/eJjeF6Cyw/Hhwx8wjj8m0Sf0sJtukBBNhDXPs8KraB3O60DIBiO+lOqP+1Z34TXzRwn2njk
iBaFEFAZydhrJx1aZI8X9gZifuLHsNYt/qfxylQ4adLrLsevoFPAiRJT4Z1oRbYjnHe7B1+iK927
BGs8u2iZ8rbXX0+oCpnb0D9Zm0miLPeJI1ajN6PJolz6lFnOgGVQ56RvX6xyXFJvZP7vwTqctqcE
KGHYQL82zmr2cperC1RJLwP/7vKNTw+5a2aBlGZFFDRv0E4jWlnF9rYokZttT5EmSZIpQprjrvad
KXgN5s0OEpXfOUQABnpWrvABgZOcT6h+5qnq+DKxrK6dyvPTM8+V67TnY+0KRhYywWGixTCyU2Hy
jePbfXzfFYpMp3w0ayeLmKnFCvKGZViAYgxJxzPMItB1wU70N4nWRvmDRI9mLSdgTw74rZ2lZ+mf
felIGwFviNcPTNGcpc2thGCUruenqZYMjhBvOcC8Om9WSl9aIP+KzP9SusKifM0iwT5ArMsrA3ul
hQUoKwCKyDjCYPamPBILibMy4Hzi7H5k0kyHmNQSmAhtKKcu6UnQTUTixLSOQA5ghPctxbrxaQZD
WkXsIunOteXHqBM8qy804Ii2xmhadPHKLwFUA30bgwdLZtZ0IeUIsqHtAwgg9bLkEA/Ac/vL/mMx
YvAu2+A5m8EYJjFEtcqBRYsMh6o8oenk8Ktw01zAvABQilDjQZGOSf7BKlc4bt3dMzFUkKYbzr64
sT3keCoKo3Sugh3AWmNSo0YzknLuXosuimDPsKNhDBWrZsODjU9Q9JBV3aKEAkmGU2LtPARP86VV
mIr4MsTmWfVR6ZyHzM+d03APq/HUGKlhGiLtAQd1Okt8qjwU9ZWWV1hcYjPlJR4L/to/9eNU6zr1
uWJd4R6A28MgN+KG8pR/3T6wvNnHDsomumSBu4tb9s9eFHxoH90qRP5L4psy4WCbv1db9beajhbt
b1wxVVJzHCuuo5TdEe9JNjfqCWJoIHtMTI43Y69H+nwWYIIQMJCsOaJU5E3JWbo2YSK4oVXtpexh
x1H+4V9dvL5IzsBISFfqNpZvsahugrfzOskOuFCef6xpI3f7FN0iPsDITEhpaU1t7uT0hABRhkZb
YqVLx0TYIc0Pd8x+keYoY8Ryb2YoX/Xsi+mrnuxEH6RcIRp35ldWTaNvYNBGSwX1jHG+XGdTslAv
umzedf39Vu7PGr3JiuagffAy85xt64zFgiz32BKY09Q21uMxNEzF7G1g5yIY6R6211OUdqsA+BwP
ShfNCYy26mkNEO+MJX+Ia2wiM+3xpDovK/LFzaIdUyZ79nOtCSYGEz19Cs/+9MMjQt0fXisd7KDA
vZgHhZkVXj+vEwczaPv1JyGq9keRLoBOHjadfRl8iQLMZB1ZDjwh+gIkKmDpZHY74kke99iX/iuz
XbQBVQy1LTHSC5w60/cVaG4bu7Is8ZZKrbONu6rcLbt58QTOS7xmShOcr6JRjcTbEc8DJQM3XFrW
g3ZJoNqkDX9Ch0HMp2CZum0ZRiTnSc0CwILPQo+Vkg/k2rfaRr+IWlI5H22LbbTHt0q6PsCD39mX
Z5QTv2iQ92AsxFI3cCotS7g6FLO1RieiqVIU5vD9d8DBQq7tkvNAJbcJksfg9w5uNNmf3rR1h4HM
rNn5oNMlhivHHDuWc7AH1Ery79tpdKEoNJR4pVCDlMOgvGqMRl6uhMGE/Tqr56zAhmcKNIL3rjpl
/tQl63TFq8YNu4EV9DDxNwZiKdAu6cfpmBCVmeFW0mP5wFS9RyRvEU/vJTa9F5YG5/4r2N7/k3Vr
4bhUWmSpmnhJvTabxTe6TwCOOsVY8nmv37aYjkiLUvjepTUVCwm6RJPE1s8v0FmWGUN6oxAC5yt9
uay0BH1V6Arvo6jjZ9dok9jktY8iLHWHClxuiUMffnrMez5sRxk8ZPtZ8w8PuNicgq/u3xlls5Dd
gscVdTvAK+wUTa122mV7pQ8svs5U4pUrycpgNeeVa/x44a+9JpyOwLRS9zXlDf20em4PC7vewABe
KtreabIoAK2WRdJeiB0MEuXZgrXJnAzydIctxENtJLKQrSQsaoJ/+iLo6kzzQSIav1/za5Af+oGI
Mu2Vy3dOeEsQFvJ7uYN9tc1n9aw2ci/3JDOkR1eptN0UV5RjdWKPRT9hdZ86AZyWxlTLfIZ3ftwF
rV4baAvHUIU/MAubkCARpmgSXSZz+LdGx9IjKMS51pbPni2cm974fOk90AJnpGXrtJ/gx3FXAnap
evEXXu9Z0OdQVA1pOCnzX9/YsGPQ3Hm1jr0FEmCEsd9KB6H4/nPxbN84ugCmAgDGPAriUUDsEMcq
nn2A9aZ1bcPw8BYmUsyZG6/OmCw/zPDzB4rsgEvwB/0KWFx0feENbADHabTCYGUyp6fHgyiXz+xE
CMX657WNj6/cux08mbhRjvSK7LEpHNb97o5apvNEpYsA5KelaTCSEZjQ/HSd/sjw02g+8EA90a1l
4jGAUCi2Kfn0hhfGQwz1LC8+tkHN1lP7bfQk4Y5Dtgoc6zxF6grW0qIeWA4tTL8zQlj0/I+e8n8I
5qKDUQ7QZyYwdEPxUFSTuu+M4AJqiNb0Kyj3gLclwYgJMCQeQ8NJAxYzRTV9NUTLi26OjhEH2KzZ
XlAq1nMAw11+q7CndQMk3hQjZHM8E3UIOkI5CYhn55HsyOOA5iAjKlwC9IJQfAI/2YLccSBMyvXi
uLpgb+nhJ3lG4CAWEfcV4SaOIZV8DrR+pz2X+HIFPcqoTHcDYvhiw/hI++3MJdsWvO55RvGqPY3H
S/phiwNZxziUKvvdDqNJ7hREjoaH8vLWbPVb3fP3YbeJMhUxGAxjv6TBhWOKcBOJZrcIJN+G/wdx
ZZtOogSRRle4kctdPs9PLc6/B3wyxLgxTPkt4meNv+724aTPVNBylBHcFXmqT8dA3+yFFsSULfPa
58p01mWFZCnbDBwUxMULtQcYMS9J99redbFAP8JWHmhJa4YS0B4rjufqCooLQ9AVHXzLxeBkqK2i
DFk0ys8vghfs8QYoWqydI3GHQm4+kqQImZbo9WNYo0dG8lUaFYp95ZoAlnPBvH1qOefZXtykLIGs
X64XQpkey1lByrIC3Abxge/HrPEMox5En6cSIbau0+4Wi9oU0apUZYU1crtoAGTZ6EzrpMCmsJ7t
dTFgyeKuTTKztjBckPmOa4zf05VENg3t8S/vZU7gryhAYy/ymA8XRrAcVpB3oSlHzLbNO6MJYaMh
mAaKz+FqR0XJxlcPirquh1VAt6Z9hIajkavysYw7MuFFsQt6Fs9XUepkSYQ9JceAHaZ1iwBLl/a7
TimYmnqT9UfGpX2Z9F6ITBlZn3SpFLhBdRg6ML9N+sJkp9GW4IUZ+SiyresjP8srhv+5sAmW9Xf2
na7kwBbF+5E/JAZ6mtompA2yqoKqT1zLnu1xb7yneaVxrlrnl9oproJ28BRuemVNau8HhUwS51sC
5Jl7CZ3cnQBoQnJeLjlz7QEimzH7DczLukJK5FpNK8RHGfgwXaIAXHkZI0Sj5me6q7A7RL7rqfBa
7Cw5kmZ0YR/hSEid7aVLUc2rTNCUeWsJ7wc8ptFCwJrtJWw/Nj4Wo5XH+5hgIZlxX3MlSx/BPE1S
917l1VI0cVEQYhvFR1lORgm1azSnv16Iluyicg6es2gIC4Y3i/1fOTpZpnzVRc3S9YCtYzuufTcD
D2fxyROzxCxi2zV8nUwCDyez0UOI9QrlMiaNOI9rakZkYt3SWQLg+EAQ/XsP117PNgYVyyXSGr/F
NL/3TXg3nVseOAQKzV9a5BNhUHEMwHU96OWkktiM12Bmgicjb5eGhOZlmRdGt1H05MpGowUTjzQv
24Zo0RLp4hwOL1cuaobqttG9ZKmcdNGRJODguoKfaK2WTC3APWDuIKkfQN8WtDX9PcuSwfSzsTGO
AeiuqVjtruR8EVyN9V6y6rUHlVgPBOH3WoAecnbmv7D55nyQ4cb5MhvtGQxf+r7io2hUVgrZ1mTP
Zzni9cvOuqxFaUf/8o/aHsinnBPC8eh3x52DgZzkw5YB8Cp3vSM/aePfxjK4oLewzl/ohfBbGV/w
g0xMIM2pTbQAv33bf03tbIvoB5oxmYVxQRnS9TjM0bnvKvfC2MCnisfWtHxLaGORhuKctHu4m00i
4QpL+gov2X0kXOYm+2vTdkIkCuk8o8ZCwLS0m32UFrbXjeT0LRbyqAsJ1aHlUgPoZfiQp9405ur6
q4G2lZwEcMKtNv6VMraMMB4WcYFoZfUqSMwU+ZD3tNP7Yv4MxwEufInjdgXRBuQki7Tb8mH/3yYY
CSBCJD6GQtegJbAu36AAKcD0MyDepAYLnG/LU289NDVoNs0nRRoQSIZw30IPiR5T8a29te+um13G
JnqT++K0C/Kn+d1mRaXKNHDyR0OTv5NTcOevycbOsX4c0+VurH+o7bx9YLVGnxXU5hosFpBg/Uct
ClvFF538RvkcSpqf4oZ5x3kBq2E6oYRPmmjVrKT6IwCyeyggCiEMza/s/HmFtwN15wSnGw0tXDr/
bSZF3Cg+ykg8KRBD/+nHV/Qp3sNWBHqfiU692NWnBuWz8SdxOsDzP8JKwjT5Qww5XC7ULIF+Ukpw
UnDmPAGkDJMs6U3GNUuRf+qNCEvxO7zLqjBBO/2VYMHZt4DirE/jEPCC26bbiFfXKP2OnATWkBR7
QR14mbX3CysUp3Q4iQPz7Ce/1N9EzeRauS7paojLsZXNsTMFL+yAKWz83kAQECuocdtz8i7cyF68
fb9sCnRAEFnQYVHmk4tdcsc541oD38HslbWXJvTOiuC6uhrVbVqZr3uugAyucBusUJKMSJb3R53u
xbH/tMe11QHQ4sKWN56Dspr7wb5MCN3OSWBfbxUToFGM6ViCI5+88MQrmKrwiy91dfEzxN5NB++t
31WORrcp/olsCLO92fYuJvwsOPp66gpUNMQdkr+T/quR41QvOeE+mla/Yg44bqeMH020elNAb0g4
tMYYm7AhxkImoIDTgOVGf6DdU1o169oI89vFJb/B+b00gC/+N/Sn8WBtTCJMx/SGzzsni6jjq4TL
13gGNCNMEru3YS7VEjHBB3FY1R0jr8JztqFE8KwelYqBecYSiV5lC55xx5TPAJqZowlzIKJ1hNlF
RY9Lsa2FDA59SW92bSYmbyT9ewkwXycLN37m+mHr6yos51ApHiwCSZ8ymVA+JoFkKltKlYiAip2K
TX4RwWzAJfgUWAX4Ka3FHLJWkftI8vHoSPlctvuRmJ5I4rEpj9ojAXQdLJYwmfDCNLFAxfY1Vcw5
iDG23EIFJSW0K214fWhNenICZ69Dyou8rVklmWUW+L2NaQ+lVFGus8BbGFPeIAqhc727SFC/ef2L
YnH0MCFuRpVXjYkyrQ2D5B7vlbZcdBPilFNwLjGxmc9Hv5Z7VPNEJrWiuUV7RnkIhpu8M89RD+5A
c9p/GyRe8qyMTKRuXMyPtkAjeUo5dDJZko8IGsuYyeRl5UADUMfoe9KzDctOwApZhOTn7rl/fDNS
STg5+lfeBuNV7AobrbfbT8/vvFnk17tggTANKB3pWpjbHpdZIP3WvNTgUBH9/7b7twOiNFSJKXZv
p3KGVUMX7dVYhKZbe2bvsgiuxuJnurTe8TZHRxdrB3lg0t1gsGcZCDxEnhZAmXa+fWDuFirfaUQ5
5XRG7rIe27zfF3x4E2MSK+XDa5xs2mJLNxKYaffILsQQ9pTbceWUwfqmN9p67pJ+oK/jkik9MrIj
2B4HJOka50vKarzKwVPPtfVmqTqg0eAtD+2o+oz/IqoX1uutxP2pD04h7LczPBoTvaE+wl2HsMrH
sVg/e9I35+UrC6Iqt+Stw3JujarwYVVZOo9AKrn8P0/4bc1lNfmEhc1TXg/RldJBso9CrixbJto1
l37pSaHUuL5ce9UqNDku+hZfbbDFl4cGTAEvGo0tz9hep/1QBbjwz1+VLDrmqPKUx2PnPEejp4fj
DtEdxM/GCf+lhi37fabTD7SSHUUjQOzcD1Ug5geVe6DUErZjJiEyZXJ1628U2nTRU2K7Dbkp9jxU
JbX4Od+CAKgQVlLzPpJIWLA8YpmWye+74syBb4O9IafovHE99bHg0d7DrFOQQWCMAPFtJdf/77u/
SAoU82bTwVdvHChtxaFGJPeom3nshpo/8oTmbLBuuz+8iqxOIXk8hzRQ/6dDoUHbytVtZLV3b/m8
Ql8Q+JwX6yT5ZtIjrLcHqC8M6vnAVZHBwDShT6PsoDRLdhQs4KDe8wDDv5Dk4eqnrK+9xWNkqDKw
kgxh5He+yKIw8VSOECWZWE3S9Qg/h915tdD1DWPJyQg4a9pf4EjfZdPiwcXxuGtj2Tmj/rqre+7u
6baeiFTpjAQZxrdK4j7T1cEBVuBrDoBuW9XiBaCL9eivsnwBW4itEXt39sNu4MJ70ffEtVgoTbJv
I+2PMblhWzavbP8iLWeW+Z6yxq+r6RNczUBz1UGcDWGALTOel5f0nP3+ttGf6pnscLD3q0+3x8DC
hZelHTkqUh7mnNWLhjh+vNvteasZMmQBcT/4heH2UBvF7cE7A8Z80nRdHbWccr8X2aGM7JP11lN1
GB8HLB7oSPoyacX/GyB80iFS0/EAaScRCrlyLFRt5v+iPVsY5lZSvaVDnMkpF8i7W2Sdj/YvVoG+
mdmPm3brmHtwPKiCVtFlH0MK700yuAmarvS8GCLlF3Q+0Q+RfR4/uyfD9YULmvzXGnpAsBcVY6lC
qK2JzYmp91F1K5jSo8MGkwm0HHQZvXM6h6cKzAMqrF8xliXKUOkZTmNMX9pHi5/vdsDzFKFuDnhC
NPZOrJWOpSjgAXyDJnE6fl+lSBQvpr9pVxhOIthsxnbHkmfs8V1LkAVHsugHSoH/YOOiRXj2b+Ts
XZmgwjqKh4mzrEOy4YwgsIdGdOrfEv8/AdOQ61llkGB/a0rMRbRCmN9YaVTyR/5as4IevFvFLjr2
jhPIDeO5GFtnanV9si4XTNuhW5isEQYV//+6W0OKx+ve+qIEQjZmsseqAbtn3TIGEZuUB308cds6
IS8Eisw85Kw4rL8KzDjnLcVpQ96Eay6kYyHxIqdcA7FwAtWo9I/YpUiFBfsO9Is5WpIqSewzEPQI
zmln/fZHIX6BTrgtGo88cpMVEdyy8yYmMvJMRcORStc7iplBIwQKQ/7wer6zid3JAcjr5tLwIQMo
Z4X0eFWq3bKASfr+0v+Zaue9XdXmteUfiIWc5tHrWlA+XLUSIaKw5rWYFOz7B7jt8Nv8W4e+Pwlp
UxP39e/iWUWjJgQfU54Cghgq7jwKHjWrRgNsOAsQpXnkbKNnGWcW0QTJiUP3l5d3m5s40qUto8/5
YWKfwBR8V7tCqKw/o1cANu1BZObiPHM34/2CAE/bEghG1r2x3SPHS6q2zu7H7dRuUHRLl78tH6NI
Ny8nSMPz0LSWkfEaipSqWQ/cVrM4QN8ISHx4rBRCQDld1s4nCnKF6oZHp24fOOJJULm9dJcNPxRx
BZceMno+s9suJBJKNn26CleGztVj3isYX0oEYMNtYT5A9gN2toaD8/Bk1SoKcRNnDhfTiBfHS8v7
VDAME6O1Wtos0ROPXOPXCnKm2L69z4SoqD1dUnY5BOtUZSbrsfkRTLd+9M7gBJTNWriIhkJIbviX
26P6n9L1Md2eBuGdHriApGPOFH8DAqt3Dg0BhXmAs/SjBTXCTw0wsLSz93k/EC+DNltJOua9iUpq
QZq+TEFn5+rz5Eqj4tJ9wSK/mUZDfXSBhA8yH124A6S+uGVByToMBA+fJMgCn1gTAwZEJyHOjawS
qly1vaq7fph/9tleqmChRpwysB//kKB3AWZOYMMvcClIRTipTKtlMTyG+URdvYB04K5ZJKo5vv2l
GCCgv+CwTi7ZWMUKQcNfK4slKI7TPCnr1TYe1bVevIJfAywMVQz6Iq6H0qo7yo4Q9vou4eFGUWm7
z+5NNoGuqmEMzaYoIV3wHaMknGDDD1PBiCqmA31s5de+lEKh+BDllTHErQ3yYrK9RBpY12e/U7kt
uLBqw7SG2gn2Fvum2bnERQoNEmxE3JktGPCgFjNmAyFG1ZuaUNww+SUEtpKctzQGFZCrnDJ00hHD
+ZCnsTO3IrPeNzS8RtTDT1Fhd3CmZaXjq5tNilaM1GkKeJjpiUnNAup4xr2HTexffL1Jpn6zvLRw
3kc3VxSbrp1uYnQGiHz3NdRje0HNylsiBN06CO3ZF3vOvGGhQPG8q2iOgEPqBVRTlZ4C2n4nQY1V
zeODj2IfIr264+zZzMxSTWS+7CXVdivkOZqv3o3FRiEelwNgYsL4gsenxPJPO2pr58/shdeHiTKS
l7vg7fnBsXQa2zEltSEqBw4i5MCJ5F1UXS8jNBOmk60dIdfA7w45/wzbHKhXPF0R4GN2FoVX4Iol
sIJGcHs/IamwcW86MkmTMMLD+0e/oLZDE+fgqUoI5qCM7tC4uYpFJbNkY7B+eSFeksEAYNrxVzFy
fXkYWCPq4VHuuGGn/II3Xit0qqluLDXs81Num3KZjJj5NkOLnqpWq+w9lgzt7wtDQhqGQcqyovEs
qx+IgM2zJu5biaKAtEEaB2HLmjzKTI5fwdjkx2LE0/WJ+D+aIBOYk9/bJBSVihV0Scp8VH5PbkzO
NoaAkC9wNYnA/moNVlsc2VkmyG2z0rLQOaPWljbu0spTgFExl5vkSW0B8Y/ovN3XltCIlFBVijj1
5Oj92hNBYz6RDC0gPBIbWNrl79Shn6psDGwOniqwQHk6794gJoRF1b/D7ITT8duaiEBUU6S+VTBb
S5kAYr2LVKQRsnH3ltBcIt+cW+KwbIYS3/+7kGJOH/TDZYp6SwwYAT6efWTQ9K5BavoH9rmleRC3
a42YYO2WcGv5rEinLWwqkCSw4aXZMaCMzz9d4s2KNz4tl9GUVtxVI8FsxZdoC7GbTIxzZBLwC7Q9
CGUu7diAjtaE4S2JBoLBa3I61QduyDuAe5aqyIwH+hjHomGkV/dcqCMcsR8oFZcdlYxOoxc4QLf7
1d4U1Fj2Jx7PUNjbEr5YSi8wQQNk2lNZTuEnClR8bRVvxE/omDDt5mE9l1c4YeuhQKhbUUJs9OmV
yuu+gGZqrzLxBe0XdhvT6kgXeWCD8arKBtJFEq5PnkJxpwnDQmvWnwYDg4hYo3896Rjr7X+BBnXK
89/hQhG0njn/26ahYBzI7TsjgPNmmoudP8Aq3RjOAbNGzQ4tlV8l3evoq+yo5RNCyHnPsFxp2KTl
tZXydfkpt5ojRdrh3DdpuG8kTh4mKhzd2ReLmYgUa0YwxfjTqok6ObnJiR9ziHo4lROdycCn9CXe
k+mi5oMztbd8/oOfAvJ9pKgcoESdBXQw8gDgDS01eHPpzEeLTY7/ssP8XbAYKPqj5Vz8E9HmUZMs
pFGiTH2p2khboVB/y4+SSPa/eW7+bSFpq48W70xrPQh2y3q1hYPrrec8rBDw7N12jEXOZDe5vuMu
BmOBkzeFFUXImf0oNvzOg9eG3pwSzEO36NrQma3LsbtPv+uILIeZiOh1uYQWjf+ejcpNGHm32+62
1ZBZsy9xmJFbZZDgcBGEsR9B1QT2ibx2Oc59U7/UNOXm7o8Km077Ivw2ch5jnqj+pnZ3Vouworyc
UE7Zuj9S+2h1ZvfJezza8r7xhnzlWGhbmHpladO5CbS53fbCCfGNDCeICgiYWnKVtRPWNUMwQ0WY
LaH/CdyWJmWnVNibbjTF5uKrQiDYolIA4R/NrDX2MX72VB9xcRorlzQVCIAPeEo9wQ8dIOsQOzHA
f5+MJcaJXjbrbg9so8zrnm2CNcHJ9yzaB5trHwm/JGK2yFMFudQsNyBhg57boxHdeNFqvT8aMPEQ
gQtziRgquDjD6aLBUOfHx3KKCK0YEXG7RyThdwGYx8RqClTHH3DDd6S0DhSxEcPZO0P/vXRVANtg
ToJ1vmr94jQ3/a8LV+gbtlmDy5pkq9039j6OCFFoDminyzlZNSN9kR4LYA4+6cISAfPHoqw+EE5M
1HYsroQyA65iFc5UY3CWBxLKq7XEfs9XUhyUE9HJ6RfcTNTIpbKE+8WhghGVBXrF4Pgw4dcBHFh1
tSoqxPgUk7dHj6ngx+Wz9sIIA12hwylDFNbR9AjmE2YWQ4N7RA0MUT0L3OU2HgcmeWrxrMdL3mMM
oEc/uZSF076QOiOS56+iqMmsKTBhhsxQ59dI/0eVIytW8YtJbszE1C1oHHGyGPhOonPyzH4arPqd
KYZuXUoQ4HuMd2nVR4/DfZSXV/6fhQFGmhH+qz0JnbkL6Mo8iwhNTbCo/DxJIkGVTx3MlQgPlqiY
KL8lIU31WbYOyC3E8SL62kvNaHqNlzS+Abr5bkp13xD+DbEhjkcVaoQbvcbW/XgkNaqRynivpRTO
FGxk6hvAD9yH7kgdfpi1rgutDpUyqQSwNyU2rBOLQsh6d0TfGkev7+JdVCUgSk4IPobnkgMeqgyO
lSNqLN2q8Tf/NFYpzYfGl4Gva+xsvM0lPa4+agR3NiMNtoSo3nvfolNn0G9UPNadJ2UyfX1lkGdZ
KzjYGo78FrLXis62SfkV0QH5OBIUxcECs3o08dG+3sTckP+6I7IrtYTJbYcY8jsmKHnR2X+yJByD
NkBQF7nRrijVDDY4WPY/yvHRSYWIrmnCAhIcYshUCGgWsmWzJfJSEmIgjjuQvNOxbjvnnkdRBMSU
vRqaP/sdZ2KN8N3aEGCQ2dnNziD/9IYwsLegRVyt84aI4PEPhC8aodoHycZLrYnxLLUS/IXwnbKC
t7OcdDJTc6q9cV+ow6yPf/M02vZ50eE+yfww3VqU3krTQL5khU+tmCTJ40KnMSGn+yTfMk8ubbLL
LPK/8tnAmw2B/EhH5j34uMoGGYkJRF+FX26eswUYFwEkV9QE3S8wOreLs9q54X4wHGjvK83HFPzQ
FVgIFOF6mGayyUCQv1hJcVrtXV6WjFWGRcrA+l+cr/A2IKFXAG9thzUvqVNubBzzXgTmdMi/tDZu
ckT1oCVorEJCTRc/AJcjJqkwv9aYT1REEirG2gwMyTdLrVsaQ0wxrZA0TDeiTWiv5N1Fq416nssl
2T2aOOEX56ALAVcDzR8OOh5RMKjUayyfaONqqh/ycRtqVlG+n/ZoUkaIyTKqI/UEPT6gXD/5phwy
miAakN3FBq5zs6o3MMWXaPngckZg8b7Z11zSZ0cKVMIO+5uc2Xl4WCc3L6TlhyoBelycpPe8/IJW
KpDJkx7pkpdQrpuqXwWg7rEutlcbEnzFISS/kGqzooFXD3conlJFKQFehU8EyWgqo7zRuSzW4mZd
Nm9Z54R9i/Tv0kA3a/WH2cbEvGmyGotXdK0BNm0Wp2kbpcZUEMjaTWpKrepMwANlK2D112nRiYne
XftT3CSleF0Gr6vN8A9t52zC5c3mkeX5MC/W7DsNAYX2tpI8xri/JQC+EBHni65mSvgN7q1OmUuc
0vzJ07OTqlwXyHp8iv0R8rC5GHPNiDTihFjvZeWTQPVUlOX+M3q6s90leZU3orYcP4NjcePCI1+n
fGPD+hMFbqBgc7kgOzYe9pvXi1iYG1wXNp/tipnpYOEzhpVZZbgDnQWdCBehNmeer47/hd7TV3mF
XnHEmDRx4LWDj+HSMib+xuQ3aAH5R7i82xPmX3cQRVZpumqwsk8MfIwPHIEMPQSHCEJILJSfKkAD
uTfd8WPxLduhW1mo/K8vbZXJRkcdPqhhFM9ABm14I/VCZDH2Rcm5wyQqWVgRanfzjkbPbFBzxN1O
n4uqydHnxpX1KLwV8jJE1vq577lGwcAAmuXPK1nPBr06VAedkG/ae6LMuWtt2UKore4957uGSMdL
ZaO9e51yWESX06S65ICf1rI0W4U3WsDuKI7eq8yZR4ja6QbwgCvnM0EOVXKVqtrcn3h+HRFFZery
eppS/OxOqWZfOdXzy97FhrLQ1vmko3w4AywJ9pGyaSqFGGpLXM5Ob9n9zsHYAgbN2NqRL9JehcA8
oSxhc1UzcUIw9JAkKWGOJy53A/bUBG+LAy4+OGaPuYDSRChxMJf1r/nPPI4JaI6rNHFUiIddjMg9
XZWwrRR1DAC1Cqc1QrBw0RORRtC4qgqKChPWnnPNwEYME7sf1vV3R0dyqEMGMNY5bFPAXl5TfDaF
UyUcldqx0yVGpAXnxB8aiI3qy+pgPupn5zN7C0pfTCeeLaqvi5IFf28JCUXnOON4eP1Y1hlWeMky
hXKMud6f5MGCu5LnsnorayzDlK/tEQDngE+KILD404hxXyxZB3ew1XLTe2Y2CXy7cAwEVbyZQC3r
WmkHOlPMEWU0OHNDsB6nv5/o0xCwO3kBn5Vz0zZlim4TWC2omdV8IMSR+YCDYJATR5VCO2cr2U5d
Jb4vnKWSlFY5Qcnk4ow0S9JqFM1YF7vEwH7aC5a86pL6MO4e/Z17gjUSgKE8DAD1HKZjHEflnKAR
OwsHiRnX2iuvhgMG3RgKkst+8Vl7ZO5L/Zs7mL0/QeV2AIRsNbu9K3xYHwC3aZhzqo0zi6C8fKkO
tkAOTsT051jdfNENrP7uL7E8Xtp/T+SmQR2zzpMBOOtJxH2KXbr4gai2ahIn+Y+rV71Ulpt4LiCl
ywlspEijxGbNkw8u67veEGlVLwO5VQlkJuJUpnSKSe4PscgdFE553sfgk0Qa3cipUWzxz8jg0rPl
Zgv3EEvxg+6EeaEkfx28a3085pYsQzjVBitPc6T+Jq4hSUK4dMWph1WQIqWdsby1oVaEL6iLKRK8
rup76HxS/K6qHShhsMGtBaFVDrT4Rl0pB/gicx0KM7goc2q6enJTrpqsvaT+DqNWliT4vNybE6Gv
OTaMv8tra7Z1u3AR3x56JUFpSLjNHqsegOesGagNFesvNYhMmKp6F3fwUp30kHeAy6ibpaDl86D1
mMtR6EEd8ZeQMiyZQZYFxiVpQuKsWlwNiv656xsllakKZkoS1svHkOij73/vaIxoFm6z5z9CWkpd
igS571hSTxkGr63YvC5vpOAHMlNJU89MwiYQKxB6HcHY7gh+LWomoWapn/REsEuerl3Q/HLtlq4c
rnE6askc4BQJ6J/EFwDSQflXKqEcz/f1Z7KkZ8ZSXWhvuDSRH9JKnT+2mrjH0b1pB0cvcOZKIUNH
A2GqM1kaxyFhshBI1Ysz16lYMyNbviXLuaK9RL8i+cYf5HhxUtbN0ojXFSlj25wm0z0sx7Eo5R29
1507UjZy+XuA7FJ/+7OEwSQcZYWuJOeEnqjCYUTIXuUACzs3RPreSXPcg0D/J/JqFDpbCpa8LZyE
Uq2/sJVPlAhivH0eEDQyi8v9Or0mVME8SPGQxkSA/dW6PB9ukpazMxqhvRykJa4wZpRgYSfOLKjG
Psl9Z6w0GePtkIfSSfazwaC1/3w/1zdeil55lPb3PUsfwVlEcWkrZSXhWx/OrsNfljFlYWmkviOS
GmiZ6ZGYAJGPFCPdYqOK400bHcCaNoihM/J6lA8i7gNzhMk9h92F8WT1TtzTCf+Y+fQJ8fwQyb8s
+dK4cJZWaBTIcsNaAZ0kQyVoS2CtDLxefMqrbDAXakSXp96Ybi+OWIEGEdFHd+0yCn8Qnr6g9jQp
SdlnrfoiW5KwGn/CWNUJB7Vtw2Zr+SeXkHsnhsaVLf+QqZJBvjfOZm5x4Ncn4vmSDTqnbsYx8AOL
dVVADssmkWip0MK9i1icTu88RE1G9w29+XEyvR7bXHdlGbBKqhMIAgNwfo6kpZ19dXY+jNLWgt1i
bYYr02ioBCopjq7RJtQHliTmHutB4cLUvX/STVS6wpjKJ23C8qCVYg6iTznQN4uCFBbRZ6L9KC1Y
/6YUWxKZw1ICC//qpMfcC1tnxudhJIpdsKk1orQNQjC1RTdnyvEhqlGzDQ5Rm7VCxZpkgfSz2nze
nND6JNpdOLKEkFIZMBviaG2s0rhb5shzJzwymkE7cLrRypzg91HCKZfyvQIrAqs0BP9bu2o/NQWD
bEsVAJy1lRsUTOqYrWgwfMD5QywUiFT2YFlDgm1H61jC9b3hpesZOQX1dElxfXU3MvXRuIHMTzpG
v1afkFbC6vuY59mlHNFSyRs0wqPrQ8vwvnIMF/ql4jCL0zXa9vEi8QNpj4Yb7M8kCoGMeiptGm7p
/ed75VxuYt9r6qy5cvLns0LxQoJ2+ZDnA8jXLAQlARdE1wDS1/JhEKwSCdCSPj+di3QVKgPnq4N6
+XGqUeg18f2A2su+j1d4oAQRqlRhVzIWNQKSDSEFzD7X8IuW0TXzkB72TQlkK4/2qAL+jLylULSr
oO/n8WlWWtP4DC1cvLRx94//d8ulzg8msWLt+aaPNeea18ujhkvbLMnk3F9xvkNX087c1hLicfUk
b7gwCsIiYQAeNuVH03GKtqgRw9yv5YoAlC3C2AJ7hDxqVoNogGoephwU3YMXwL3sRfxi/ursxyV2
eKf5Ef/rC5Cy8aoh1HvqK4PhPrVaTD42sPJnrB7kyUQSursifVrlCsneJGbeKLewhNZ0cyE4WYvS
MY7zBI/Lzoc3znZmXT5i7Ysv40woOzVET40C4lPYQtfObhOG6JYa6BBEm44UIs9kuNDagG4/WTKS
L/gcavdLMNMlieBNfP/X3REq9G+Y2r8nPPXO/kVHx89La1kPJPqJbiOS8wv8RbbmaZslS7z2pYLK
yLRSSfjICBK7694vVg5gw9R4jivZmK+OkOE20AfB6W7bpzGl+xWXy4UhEzMSygDRAZ/XM9ADxJm9
TiYIHo5XTzSodR9Yin5vxQOGNx4JMPVKol7fr2LYXKOKGX4NQxdjBMlmyPq2C6FWbwlqfNkTAE6q
8BapDLOkiqR5AxaLPMTHemcahQAQTul8phiG0wDr9XOUtTVCIG0YJLLiVQw3u4XCW+OAl8/nGe65
L0gOpSRKk6BERgnIy9EWGqnGuXzhoRm23x5sljO4HD8YfKu1w/t+4yIbPkzIAQ7umZcnCvhlyAcM
VwLBeeJdkr/lhRxX/Fy3P3E6C78tLnqPWmyEXMTfnBNb5OhOZiAy2z1lbGbfIeqa5w0j1JKulcCV
NCxyJn+SXRl9RsMzc9Yo32lfcUF23kEXth+GCsn6osNqsR86mlALNmg4YTKbltOKZf0IIrLTawd/
a9iy7EkrKEiM3D1mb/TDIy5abFJefZPjiY3gsXDgVi7tQ9Fa25ZSblw4SfwQO2guSjh9odUB9RXv
dY2VpOGCkelyajHsP0VtLkdGnaJZuQTDeokEqenwlYLuINHMmoNtSvyIHpT5MYiu+z4Y68Mt0Y1U
GNYaHsxrhDTWpy2TmLsHt/XZadpcGrtipiyQNhJowCeAmBZgykpoU63SUDgKqvh3PBO9aEy9GdkA
EMi2rbXy17NYDAdWA3aFQNKvszxrHK/YKcYjK/Panr4bOOT4e1rZEi67h5tTUOTcTY4lguLpKJ3x
eopY7h8WJdcDD+HB+M7gtxl90vEsZawXe9ReBFgChmBIIF67RHfeT9RmXarjGF/rk3icVdnhC4JY
/CX8XZrmZAVQLsVcltyAE+NXvv+kmcwiDkRbEw4HbUARKWFdNif4TqLpXse9tLtnDZjvy9EeCjrW
DwQnFHDmHiF5IuDfj5N4aodbloN7d1gcSAiBa5vHjZjJ6830nkoserB+SF+0A//V4N7mgUeTUNJa
rNdTgmcaeulCdQI8boaSLNWIhPu9ePkZH8niVk80JpPGXo8eOfd/SuQ761Atr4i6SD2lmggP66rk
MvamE0A/W3WHIztMhfNGP4Yd8/7/GQV6E/lpN6WOfNUlm4Qm75UgEwm5IRxs3bhFVRGL2S6vgqKI
lvKYkHV5vwA7SYa7gl6tINA4khdzdyu/cBd+evh+9YzjmdoJQ9/UAfRvo/zKNOPmR5lox+7HlWRC
vPTIXT5R3kbzuJ2L+vyKf7L2K2FMiLvUV9o8kQX6cldgRsJ+oDgC3o7bdYfPMODt3CFZFjJ8oJrH
mdIElmIW5YNDPTPl7q1fSFJAtxwTZ2AGcfMiclG3C+L0BFSBDgmpze7+jxeFbbDJlF4c76L2OTkP
YTpp0gT1z1zIKAkEocBYxz67F91A9enmyV1qqpgExA+VYLr65sNni5v/VA76NTvGlzPwwexo9Qme
xQkvmqb1yuXAdzV6kKj2XQK2+Y3znHSBjrh2urJCyJBnlvya//Sied+SIA5IcS02dbcNmPpOayfT
+gCLApFWQSl9kRjgyeITm8Id/7vsgDEM9ue1dzLLKXd4Q4H+PhiJpZlLA/ygUEttLJpPBwOeig/W
zUsSs8L1VczbFGw+Zxgic1dDn+EXXlaS41PR+H2lsF+43GxsDaWZ/YFANDr8T1YAIgDG9bfPU1yw
rtvObxJ7AKlgHFcHuMQLH1u7Ce00wcMwpAVVptB4nK7tlTBDeJJM/dIUNPsEiTC/JNebKe91BCa2
tInWbHzfBXpNm/D6sidNOe/ocTj1QgUm2NFGQc44gMLWEdOqcPJjlWFTAePoVlkSaqZ88OWXJZkf
awAxvXr6+xftR54f+JGZRzLTe1Ih6Mh1/CXIVfk7V+Ua9aOeubNO/+s7SbYTTJlwE8pE5DasROBt
iDUHMJqgOd5T2UiYaPDR9a8vCfUUMvXE3o2vtC5hBeQ0R2H6GcfUPIp54+y7/0JiVsBfa8gFdp2S
GDB8R6v1wr0IGndz99tBymDwN9Uv0a7p7SnBs7q2w0s8SOQbgJeVa44p4tUsHSM7D2zN3Z4zupBg
3pUEgjPKzsbQNzA/0QvJcADrXhs6AaDPTiP4/WZxXqaez5A+zi5u53j6sq2odS/1zHSUHO+IKEqz
pkBWHXbLPf7ZfKNNvgC7GvjaMyRtBqr0J6Wo1mcsq84ufTNdftOdiTLtl0BQo3UcvlN/mbMNzVpV
qTuueHaRsYTGav2BqaPkiyFuorfsIZgNfD1M+cpI1hu6LvovHIqN5KrPP9glT1mdCdXOMvKMY1oU
u8bnRBInvrzHWnFlpBvg3M75Flnv5a5CNI7urTa4EY3+CZu30GkkKmC4Fg7p+qGioX7q4OUFB7wD
/R6kSlSxS7TSyYhvVdRVeLsfP83Iepc2cet2tkENBBaHpPNIbtCcTbM5z6wMnPxuBvACMsQ4gQP6
uGFPfFYVMHTwWrV2HfPXUADUmP+NFTL27g1u/dGm758mjtDH8nUqqwV8dxJjZ696+c6+9FuDRmv2
QdD7jxeslUvrxWpiSrgDoTWbO92YH3fFbNpdz5AuAQ7j8HMsnk2Q/a8G7c7b4wvCrM6dqzpW9GPQ
SxlaOTeMEVzI/ichQb25G/r2vUXGDwSDYS07S4FcFZPZg9YdFTPwI1T0bFmxK/YNgLK2owwUO9B7
EaWlRNMydGz0FsAJwLn+l2nAOB06mUNMQwpc8QMRl/jZJvBSH4gWDMmJV4u0teFOD/jFKNKHqd9Q
+BDhQsybCvO5rxEkSlaFpJjmeM1mW3Du2qeNZlPDLJE1+JFHHj+F9nqcoZrmnU3srERosqhtpJ/v
cxQADQHAtrsrto12KAr7Jongkb//6dmELXCMXsvOu5xwiY2YqIyZtV2kkV4PRVNiAkDun8cKraDz
gjH30+n7ZRMwWOwrdfeEHQCpF3/EuiufjeinJOnoXKdDIelrO5kGBdOj6pQVFOKOl+TQyVIfXbyX
4BVEY16eEe6yKZ0icx1lVJjMKGxPFESqIz1X53R+/XQOwoKJse217ny53W7hBE7MZ6rt+7OGeTNd
SNFPrGwMZ4QfH8A4IXhCpy1atSBq0/GO0fXdpmutpIudpZQIMbZJE3edKaboRg3UCy3l0ybQ4D7T
rI+uQRFXCJmMuH5ff5ZovSYwieEhWOGllYxR1iqtTHjC6PgXEWD3plbRUOqNat8bMkeXc3d1bEoW
N9lI8vyX4KXCg/A221mYQ9fpnSAQ6z7/l97dyEPGn+AHq83X0Nygrn6lfzTp0Zv1A+2llaavqprH
ITtx6HESQFik+daFkeQas5r74pbRKC/qiiwTKPdVDz7HIkdAcTBjfPtQGqozy3qpH3Dd0rKzJ4rC
u6LHER1zHLiyKo1/e2XTC+R7CSuXqRNUyiu1Cc2pRJDw1IeCpnnwirKuQBMVIOqGvS5VXbzezCXx
blKasWaE7UX0NrPoTOynQgwoEODdNb4qt7GAvstIztBKhjp0GHfWQUlkT7HxTHXTtEP3tqEKJ0/E
W7aDrXC67lKDXurC4whgdMUk1593OEuy0l5ioPTgXEDWXc3PyInzObHoDOM0TMqGtw+x0cD4bEN4
kiMjDPF8afmv8K1WIP0y6VAWQjyAqPF8XDqTv2InABoicIDtD6XfUANeYy76puKzsYfkk2YhV9Cg
dgZ+7fzY93eJE15An79Yr8K6letFvVDxP2/ILjm7kose1SlTCf1nKhPj+4zxrjfh6TJ1qoUvbB56
86S97Dz8JfL5B6bpUSzlm5CQHNHwvhvPq8OZyEr3aQ6LKSJ+C/ydrOReE6k4iN49WILy+bFvR4ze
oLKmjJSgG8xNt77TOzJ5xta3FCx+LDWa87oIAawtAkZ/fkWX6V7TEqA8By+TlpTPJsPZkidr1euQ
wuqRSzAtF95B3QpW9vz9czOz4TqkKWRgeCRsPdGzoWsPhe6mFD8jziJjwZjGWqPsMFulYOAAvlW0
TaNJmU+h3ZZopRJ5yPTrX8wH8Lx+nTTPbedax+RO4Xr7bjnrZOKEUBWlBFDqOFxf6dvgxfVNKE/p
TvCca13RmFYubYfg9PYJuZJvf6HK1j9hORF7RUSE+snk3lLF9kCA0W5NimOB5MpwCS3zs9ScwH/8
7tZI8oZEoLjpw7eb8Zigh/zI6LLYRSlnaaF9trsgW8ZXfyH6f0nxqzHUE4gm8sYRBunswOpKGU53
nI3Gxs5FVdDBfPcYg09/mrdM0l4NwQwV+WW30JcdrYIOrUnEJhyqbscGjdq+boJbrJE8vnI3Mrtp
OpDLiaCXJ2jSgZzFIi1apgX01WAs9HOAJ+SNg2NpcwkJZZKD7CVuB2d9wWO9BrtY9wvD+QovXtkv
p5pZIhSj0BrrOLuYIR1Q9cjkJervLEPWy21bAFlnIavOfmyO8gpOoEp/qbravorniE/lnku9wNnu
SFyXjAohvhrpX7lmk2vfl6APFcygil6GC0Nk09P+ZGDbKhTs61VA8Ep8Dfgz4JAFmo6fs9g15Tvo
EGInRv08J4G6JZXhaBFHtYUNJPkyAzQ3EH4YPSY/EGBpLXpiZWdvGP+sPgUivGyIjw74N5454iia
PVL2mpboT3/vLn6D8ljxpAZB+l+Zi+Nws5QJu6fp6GE8W9mygw6w4TmnD8oGs2CiivkxPDteEGD3
ut9dnYEruHmluLknsJ07DbzUfc8rr4wXMO1UOXaHCcolaaUzl918mP0HniK+CI7UzBFH2fpT0OGN
6Bmvtw7uOeloFuTrTYYQR4R64y+RQ94cuDTxaqNPl+h6FHbpbDvSlwD5k6MEeIvj1v1E5fGBUv4A
iXtL/DZ1VUiVV7k0AMjsowmneM7TIc5d4TsnFL+bVWsRQ0NkPWpPZdY93IOmfKExE02HBxH+6ZqC
eA+IMAee+DbyrTKp1rw3mB1h5uPeafLRG0uhuqpdCU1z78aqoInNebaas5ipCPkmg06BVfl+smHy
7anlsLOm0UakRaE9qvXhvneYFE22Jhk7LCADEWJII2uNZ48IOJGSX65SLrPyzaO5doSHAWa9oI/T
zRJIt9amvi2iwY4UNCDoy7xJBj+oz+AnkRsv199jLvipDAm99aZS5EWH3DbbDb71rqgYu4iA5i8z
XJBlM/UnJhmJmewVl5nXysyAUAnb2stDHPoS3vVUVRwISElhob/0YaDgcJGPT0N9UivR/uZHUOgp
WAFGp99RLQZVzx+NLj9Xt14WeTOp4YHWQ7/GfzpCnWIAwKvJ+rq2uxN+HGJ8Yf31mJeOgdX7MFtV
DhHR+rmOmL3TFT3fCu1DYycORlnbyKHACJP1K6S+cR4YjlEIObpynOWqtHs0qM3PT+ENcAuEH0JO
9YvtYEm7z3p6uXdhp8/UU6/bsVqN+Oz79+bstfS67UVFcWZ9I4yg5jj/UcHSuflE4h53ZpZc2qSA
ICzDo/6zc2m4qWlfKGgIdbWExeRtiAWTUcyC5MQEcbeRqoQNlaIK8/sruJGA96IKYqK6itH/TU5m
dXkGskX8MXx8iWPYHaz+G5EELs2Sgr7uBIvUHDtxaaehoQMlPza6t7mvQyYDaPKs/UtJXqnK8MJG
SkYydKW68Z6mvzNxNOgZzd7tCUxQxE0NE0M9AA14aY3AseVXvoGN6nEvJV9L3AOy4GE8wIM7GpgZ
5Rvioyb2okxFLoqmbf9c3OVr+cJ8cdin5RH1qZGHiHdhp/L3sOogmqKFQVQ1hb1hqEeoZPCPnZqK
9gv4U9m6sRewmxhrL+VooPMpX7pQOz4h91rg34YmqYstvKxnf9jNI3ppNVOkV991B1NqH3CWg43W
EJzQta4KWSGbh5kjhTNMGEGUtTHHnf6e0iP7ho+7JXuJsJlCszBD+sozGzWBjYTtNizQQ3RhHGlF
bEFTgzM1uakCMdtjfKCunwSW4DAu8R7UckFxlPsN6M01SFfmtKWYCO+lJK+u28aqwBtnchbn70Fm
AQkIBT0IWOSXxofvCgpbnFcLDeeQQ3VsvLorgiNmMYAZdjWC417t14ZFYT2I2+6ifQp6SNEZYhJf
BIO6F0/8fNf3QkvA00fF3vU4Df5L+bwcU1JiDztp6bU1RTegWi3P4tQSNqZlU2KvxXIPVEuFj/5L
Km9ajeiQmUucTwKWbJnzJV7jGFauvF7fD4DJvg8Nq5sB2xApAy30VoFxveOvIYtgk4/pCIaHDKHK
H/Q7kzesFNZFICglB3I6FghkNgOstPmd5NgdB9J+xVKKxl/wXPHbonIITP2dBPmuedY12rU91MWf
KAeiTYFkresapvSiUf4ksi+MgEZbv1OdqovrBw1nmjbHtDSS6763NH0yuIZ+2gvX5QSUq3izoRUu
GLHLFzql8EEQUb9MCjS1V2eCJhMe2WseGB4X8KRXDlrPM1x8nnrtrkowOjB+a3zt8X5fO26HVC+v
rR00zHlfIkPyIqrUXI/zGUb1GrF9oaVNGm19RDeh/6oOF47LZ6iA26h4RCFMfWgQm1O0U8BuqtyK
at7/gX0A4KJyfSfImxnbgyMO6ZBayWeVb5EruHARDxOLjusr8Rwmv4grqLN39I9Ph+5AE1er2+9S
Y9pBQQFkCAZv8JXbWEZiXMRr4jFcErpSfClZspnKoSP9Vrlyu/i1iepT7n7fdfKFPgqI8x0luK1v
MkzF73jeL2OTjoMAvg5r5XGlPIWZP+GkjIaximlZvkEsOFkLAB0QgH1ZPIjbUeoyXNjeQ3Lud4yT
0W98kXwt57gfmgPCYImbzM/PTQ4CbV3sCn5lD8NOsbMTO1duNb6MZ5TxL+55ydivELsZfJAaz1Po
xMIBEpVmHvZOR17D9Gcq99VMT/p02yFUrIBjXsromKe9KWCuRfhL6lltamz6hcCtOhrWlki3DnWZ
m1El6ouRMeh4p6xiWQC+15tSvXLbaAicTEjTDRLceWizwKsmHfMU3Nyys/O7MhP4sCu1sCg7gV+r
go6tOsHV1x4/7B6RG4SMdCEpM9/dDSQaVvWJp6DezDR7hl/Kjfcgk1VIEGtffIcqiWO78rmvLvzW
fJO0ytZhXowvidiuPscvHJPGp+L6rSlr7v3gCnBkfYN35rOQmP5/gYl1oSi6TFhnG4NKcJHnjdUB
vyvW0+BxKl5XsJohB8gvfLwtSCt4P6fCEEA6hd+v6jXyk/E0lXBXs9+pzoAX2HSeyLnZJmfzGYYq
vx1xXs2m6iLbKiColo7unj+WdbPd8GE/PtcW5TVWHITEqh21q8NhcOnRlebCvWLDvMcgQsEQEO5U
+EZXIOaB+G/IGbPOukWBnudzRf81yHea9YPsV2j3NRmeBdhcePxj2e2FujoqdM6u22YZZLi0Ur+P
NW05yg3Tnswb0I1vMYU4OQyQU8FgE1Gcjp7U6e5fVHjugLyGTXstLfLTGiQrPbmGZcsO7QWCE27L
V18/oo5q6YC0vhulgXNUCWULJwj3sz4Dqu/7ZeJv08h7qNZhXL/blZwbIKFtQ3s/6VEh6AbeZ4Jj
TJPYpV876BXkJO0Wp7jdZ2gKvCAVbE3aur0nb9392yjajSpFmW7V29zgHTsoVQDlf3gBZAkICsHU
h/6u/X8UpyAc6MiQvPIVGrbuSf8akQNOVufZ3aSbCxOuGkNroCbkdjIS3Hu4IP7u+ifmRa/zIot2
Qia3mBfw0USu4B1ydh7EVU2vv7fi3kyY5xfEPHXCA7dSZY6mFN9OtBTiXjHHekBR6+QES7PlA4+q
L5zvjk9zYB5bXG1gbmdW7Ngs/jrIpPz1kToSLW0WalVB3p6HacfMpwGtdxyZQaUeQq7zqrAs9Lsw
FLl5qakzOUYNTlXPG0/IMnpoD7PGkTQkrb6GUcjdQJ83Oop4Ua7hSNpQSknEDHERwXrgXNRegFg7
RazDIKaVh3SHJHpmRpk/aNFInVCpffLOz1Ki9BdR76fDVaVIYYRcNFF8F0NrQebWxYCan0zb08B5
dygUF9EWzEbflsCBqqxX/qWu1TobPT0LunH6u6bwAQhfcgP23hSCmEicspVh/YliDjfSVt42v5H5
dseiaHWXlVK3tpNxtlWpt+kKhoOge97X8O9LJkg3MFfx83XXUlP8amevwxsxbl7h7S8v2RSz9Q9u
75Hi7VNNGg/FNm9bxi8gvwn22HLAv3hLuO8xcDF/tBUOMagkAO3tTSLCHPXMfMH6POhIS6bvJ4T8
RllrUQmRCoTcjw99N6cqw5XM1q4RY4qkAgbgs/csXg6tYgaO+WwB3mybQWzc4oxo7ZfPj5XFCL+J
oGxSPPFGlDz0GlHMK9og0nkK6+qfCPgRFR6jSx9BDZQH3VI2EP3pHX5d3Ms9RkUEie+hNPdERQrP
uTXL53unDRXf7a14RU4RQqrCMIwpYMFskRGE/rOtAUSIXAXLQDopEitiN+4ZDKSgab2AwNPQUaMQ
jD4rKyCC1OweOWolywABTJsqXjU9EzO/Goyzl3nHpVjeX0nE4R8J0B0Dpkaxf4yHcw/83N32BUY5
U3eSO9cZ9STUj0FxN+BAn7YphwbOW8rjP633IHAeKIBgFEtDvy4MNt21SmwHAD7n6DQljMMXWx8i
N7oKVAwSjY6HMXqmegZcos64w3yOWxO9Xflufwy1QH3K+vU6uGTTGSMwF/ABRry39Pjq/0dYDXWK
PJ+DjslAmTZeEZbFMN5azEx8X7ElWgqblabdr9sWw9sqTQ1HYEh+YrO1r/bIJe5zSPwPH04hruEa
8ty2xZzmmVssfz1WH8r94MfZoo5CKLQ92YhQ2eFd44QFPzitwfzhrLjCjh5WHQBxSKdCYlNHNMsl
RjriLqUdhDTed3+VJn5B1E7+4GOHXtj1sEFytWVUfS0qcpNh5EO0zZL2rV/3oHvenfZ0X2mI/Jne
741iS0OOoXZ6pe08OPwDBhG7d/0+DPLuXcYaujiKd9AMG9OWi1QmHAMVKSWVX2413AEFHG4EJOsB
KkTMPJiam4HPT5rSvaXvcaR4ttpbowNdUwkFqiIAsOzQpOwFRldCidxOYs7YWJcQtx5khH7SxMY7
RnAYqFSQsDwccQLTGr1+cTOMrGSYOIEd705Reo/25dbdMdbe+jDcoUpBAK1R+Mlv6scihMJURGOy
X/EjpJb0UVyK6LVxTRyf1FezBybMaICLLr95mColGHqfpAZgdwVDSydQJ22nlJTjOrVRxcceIBrs
5YvlFfKnBpXUKKNA+5NYbJxD2h3LmXGYvF8hBJGkj8KU39RS32vSSGeZw2Ec0G8B+P+h9V+ZtqEB
JxeIDdYYr7p420aAZcYqFgxm12Aid/v8KRxsb/pS2tDwGJaCiOh9MkLBVo3YNlFUIgLMhYut3ya2
oMu7b6O0R+HaCJ3g0HgIUuLdiCgoSffmW9oJVV8j89hokx5+Ulmxoz/7mFvwo1tVVRUWF4YnG/xD
E4ouue94aOFMKRbZj15OMI/EASotatxGhYSAJ4976crE/BosuIMhoBkRP1FSlx2SzfV7qoXnXe0V
5yWF2EonN3YHIZJXYjkr5TggN/CJd9rBoS3qexJVKFcMDONL3ZPgpIWoXjoI4pTR6bbR7WvcHtH1
cXDnQKj3sj7Ym7QwxkCotrNQF+f3J7x0SfwPCKyqnqGe0YGY17KqsdoPYyubCU/3zwMmSH4f8GeJ
ToBn6Pvrd7zMFNJeqlsRsAFbSjkcHpz2dXZXkfNYmj8kmUfc1wftdP01Er30cY82FV73HuwPdTq9
YnD4WgI1hWCmRj4G0D/6/q+VkJLJ65RMzTKqLbcfyTo6KMG37opGVwsvFH1Je7biBWxZlZIcAt2o
1S6h0O975BeCrQk9aUmKmfQlyCBrZOSde4XkDlLTk/kZUWAl4zewGXKxu+QbYdeSvSsS6vTKrj6b
pm1KXQBfUN1LHxcnuv+RG/gUkgaftNpXznql931HqQGY1Ji6vbpwz2g96xgmBWpfQSQTmVblp3+S
CsYqk6ooWu59lagYzGysu3CE+KLkzf9FdQozOODB62iskDp8U76+hShPklFnAv72qUcRPH5FyLCE
ADbc5C+G84UBGX9ogs/deocTK+VdmtakQATn/GqOPRtO+iQ3mqcnaxkNR9GeHDagVGtMu0xjRhHe
9qoPz9ULTWVAzfMVjspGR057aYia8LAaQbvn9HHiNIgJ5ItUNg8s3IYwo5tX/dh4I8hdMINntB8F
KcfjUvgp49kwH4GT6FG80o0TmNJXI9LXbxGQuy3O6oOZD4zWNf3I/UG6d/ELhUwJqvgXpfJs/f1w
Y+x23vZ8J0alB5D5AgsxQztgFHFqqX/uAUmDj1p0d9oWiiVHlVT6V5ELHK9NpeWlI7W90/tGj5AK
u1gyks91Ra34qhRgALfKBQH9I83K6tZDUzkyWOX2/9gd1EbSE+OqZNSpR4vr97eSSLhMedp8odUL
vq7y++QoqlSg70S/iaap27P4dp872SFf4dXHfwjh1g1s5voJ0icC+oh2St1rzUm3Qzo5LyhmIMzk
ym86pDzKPTUhrX0oHgMrsnh5DP6e2Pr/lPSlPSYXsjA8KS1MUvmNDr4a8Ej8Zb8KmCxRNrwnhZIo
T0xRA8soEKvdI7MNrRSBRdN9TloQsemBQR3/xZjLKDbg0d5FL3G79uA0YAZzSwF42ILCrVKL9b09
a1pDV17taiK1sx5sMWAc1kF0YiOfBNA4seLp6y6ZOzwD1NsUPlFTcwbbsi6vIDarXldCcH7C+Ybq
6Ar3U0WRoyLmDD9hnqfhkW59Fa4o6itPaki7h4M/u3UUSwfiNjivkzRanBKrejf+MhEsUxgxNxVb
GXi6q0Ww+4SkXDTYZy/q74NkuZnrseMToj5ZeNTmwqmR9Bb2VZYrMeZWmU+qqW7Yk0y8nDVdDgaz
lL9HG2Beg4QMwF3fvziuE6+pCgUdNxcq0Wj7MeoAlIn+E71Ya4HG1v6MHuKhcnP8KfjXMVRkDTix
ZRUwxkAYiliAtWpppz2fyPBiz3rGeRasAW4zT3Z93AAoHH6y3WwcTJf27fQriJotfp5xWzJhOyiB
dR8J7juH64qLq8/8tHZRySk6m9AntNmNA/bnUMbtL+Q1zISDWr9LARU+xTmu8NIjeWvmrEURj5QK
bH92gqbVGi39Ej0/z4VmTV64GqDHMxPt0JB85mkJrwO2Va6rwatE3tMOwmsYgyY4fjbOR8FcdEZu
ffyB7Z0F85tXJ30jLp4wJHvo9kmHDHRBvsWDyRde0uQ7o35xK9IGv7JmpmCxXoaWB0tIo08AIcz6
uSoncHWxbLxmMSBi/97RoDdyO6VcD+roNjHuRyHBO44LjO19Plu6tVNX0hfixmAJfMZ6VZAsivht
R9vUyv6kh1j0hdHoMMrkjf+3wrQ1EGoVFnHYZvJyhFKWTRhZ/LFQpfASaOnmR00bS7gJ0XSYbzMc
jAcy27RjZ7p9XrqXKYHJ5C5a6QHPB94HJ+OaUfpmOyP7h72kVeACV6wg/+nv7z0qUfiuPZ5WTuaP
b4hNqJQ0aXKCbtHegNFuLPTai1+BxDXgBkxDI1U18Gd0y7kjpR202cXD0Bqv3lfA5XTVfje5AL+I
EDq5N6mttZ9YOFqsDXceB/rtcIsmYvEZPtWJPBgGVw5j75FdR8NDU8SuyY1FBfOwaJhJTIbD0HXg
+zBCv04dV54WQePsrl/rKrKSoYH3qDa7cXED80FSMrHFI2/WPRGLMjPQeyj+dfoyYWDAKm/kITqn
V4uz4ZCVtqePueusR9BDTFTQ611n140+7OnKbdVrNfUgENGSrhKKQDiA+ymZZn8q91TEezvEnV7P
uoNnnW/o45Hb9D4hr3zpEdUwGDfir28JU4AhMeSRnpVewLKaokRqX3zxYxpam4aqkuCeG1OYrNSs
eKCeVSQTM9IIdY14rJirZfYwfHVNDCA8m3vLZJqRoTYt++A1s6A1dXzOkJybQ8oLC34SZQpEq2Vn
HN7vZUjC2u9lN1vS16VoJfLjevG5MzS4i1rGeG+uSGfJTc45IoqIKV91Q6MlPjidxTti/ZxUFQ8/
hSQLJDwUchKrV2ADoQNsMLKN/8exmHJcFi3leM8b1gnFt7Qyoty4psF5bxM02OFaFq4LKHLMOf+L
VgTcZUhxFgkaqwZ6RGhNzJ4VnXBscKInspuEYeqKgsoibYETzu/6STcN8YVb7DxLgu7O/cjQ4Ioh
FSRhB/LvUG6Dp6EciIcJ43QkVQfeFff0VfIE+eBljwyYLD6XDYYSm7ALAcRMRE3tSAROx87bLZpF
yvJdU5hzmqFESMoCJwzx0Z8/Je/0CTvP5zDh5hgm1Wn471Kw9JHwTslqQLJ+L8kCur5pnalhF1Im
XnJ1HGqzi6GZMt4n9RKYyYbWC90vgh8HmmO4P5XdMgN4FNI/G1ix8sh8PJPQxaZph5+F/b/IEAhD
ReIDEXwI9AEigbov+DzmDkucUDzxTy7l8ScGmDghLIMGDGMGddMmS1f21yuHY9m7UhltdwBNR9AQ
YrSFqeNasrp/lUQ1vJbgdNRzEYLnaQZirFL33eNhQBYBU3VFspfVzlkM/1Dw+KPcL6g5tt9zKrGk
daQrF15GzCTTAX2moZErNijW+xW+iDyLNeaYyNi1+TmiwP+dAlIUzuWMksdG7Z3rdwkkVMrZ8X8d
p+bWdh8lyR97nEu30YHzV+b/n5KGRWX3WhN/H6fGddeSWLcEAR9EntKZF4b6P9ZB/9inhYaxRYTt
6/9niuq7D3SPCo/lWaYtWag/WN9V3DOXgpgpaooJ1wz8J3nahoufvx2ukWtvkL1Qva1TJw7+I5q3
fUJ3UXhNiRNAWHD6HNmbTqmJxRZAuKo4FezQwX5qzXE5nOGmFx0ay7yf5xMQ5cs43NifqP65JQYA
m/VjNPcuZPW8HkMTV4xq+rK2t+vuGUY9bcD8o+W4MwaZfp4OdV2kA40wsqWwwd/OeXQ6z+ezRcNY
hAFIZ7uICBdnBUY88MAELbWLVeC4rFzlt7urRkvronyHWzyHrjVn8eXnSpD8CUzvvqKAWLj3pfpi
E6cJ8YPbzElVJs77LP3JJkyhlmSI1A+pTbVzwnULkLunZP4mWaXBrh8pFh4iTUTb1n2NQQDSadGa
JQJ073OF9wkVw1EycjH8WOUvpX9VIwPRGLYn4UkiSj3BI+4T2uaymIIw1IUecUrmm2hd3m3GS53V
WbLx9fi7S521uZNJxG36eXrpgXkmuHdVkrOzyr7TPg0p//MiK+ivxghSAd03AiASoWk/V0MhAjZI
EW6W1+5Ya3w0mTVDevopKxHsggEBxYXDDj8im94EdyJTt2nlY/bDq8kO4YkAkuRRyQtDTdYRIPJW
Bg0pyOEKWGyA/tiQ9iDpjMg0WMg242Xqq01Lx33tAhO2A+jtfuSXN9H1aYikAtKm7ro7Q/PeCTgW
TY3dkLpSVRz2i2f0R5AClQEeODT5v2scq10sN7A3o0EWfs1D1lr8kR/vm/NhCc7WNmqOkKKjQu+4
PljmRFwCnGp4snDMdIM4wgA+UUErT3S08QPiCrqaPaTtpfPxql+NxZ9Os/uZh0HiHw+27/p8fT9b
gLiw6UKhMFhQvqLLrQwfrcjNO86VD+j4jfCuuIJXT9urjZ88FRsJYphZYIt5JVTHYleSOWIK4i+0
MflA1QKPXwIDk02+7UViXIBYYZf6LDkOUojki6PhbIwFm4HTs22NmX/uDrAqVZXC8ZhSytfhiPig
u22Ljpp5m2k8o8FIllf2h0eVnB9qEvOkmSb1IKRT5KqkRZRp+w2RAjoPw+23wCGsVeBVz7aZG8jf
GVp+dzjnNMqVzmFFrTI+rH4V6C//zd76m1qPL9eYSDlt50XhTjRV8mrC7VPrvkkYoHWQB16soXBx
LwodPxb4lEO3ISMZ0zXjcB0feawFyN08Gya08m8+k8VHT2VqNfkAPQFW98Q1SGiGKuON3rVLr6K+
lb0coZmAKjwtfkhyYm4mz5l/zOrMuv//Y3Qzt+9/I2Q7g5OX3W2WCnVAvfhdMMlEV+tpfAZ4Krt9
+05KA1QYR7kB3Zbdb3KR1OR3zeK1TXG96KxPNlh4bEsk9yD5HexC6Ii0J6lMzLPktVhDSicuXKBr
HATpyCZjWP4ZeQUHno4FFY3jP/oazGI2Q8FCs09o/odv5/kKnTBH75VzgyaHrZG9iRC7cIBu0vCW
lNvDjUnx84oQhY3pSGrFzW4Mybf60D8H9ExcmOtCqE5r/Ydi7Cfdb2KN5uqCimfXkCuUfuzJzKUX
YKplxAp1kQjhBVvI3Zj9ZiCoLklLvueleu3f52vBVIR4IYDAgH0zB/xnyxO8WGFZ1Q3NCfuizXmq
5lcQNRr4oXl/gNdnZR5Ztl5jz5Dw0M++n5iJy1KoXaDOBIdGuhXqurTiLl02nxe1herGQy8/CUsK
UPPFRrQG0PMW3rXKovCVZou0K2gNfI7Hf67YeDMF4yiS1nToksvGVgK/+KFwrS5NRmtgNzdaIllf
J8DzInnR/ZIIcn7THuKhgImhwQ8EaS52VjFuSQ3IoDb+D8KEpFZsDdGn8MiHwQ18jD5+ury9tRin
xWV3SI20oRy6q7Snlyn2WYwy7bBG1SOtTMjamayFgliTxOE2fnkUpfFn+C3SqluuHFLxAQH6pg5x
L5tO1eolFgdA4wxrjath3mnIXjDOJro2Fr80Y9Xy7YXfxm9JHy+IXIcjp4bFtJN+wJ4xrL5KTW74
uCjk1i91wWxs6AkCh+JwqCe4VUkD37gIiO6iVFa8EyztgM0zxdtTM6sF9bFWz5YBqQeMjFqsgLVS
QXmPbE8IBOD0AOYtdq1z4NYer6GtLZkD8633fEUJ2944B9NTDuTqHhxXYO030M+fvLyN9p8+GTLZ
NyrQ7/4MUcHt+JEPFNGHdzQ5hAPRjVGAF1FeTXQPzcqPhaKkqjuScPsVwrRH/gyHlCkqLycOveRD
Bar4+IWFDMhFkuho3d+bNbMlbXIDPyA63TX1FnRouXqYswc4ZN/tB2XI2R53ISmtigLcG9XePvrz
aUxSsB96TLvahTQ+aBpp+ZIV0jjnGFhn3sBosa614ho9Ldy1NpeyMhTREUp/GzwQQN1TaPBscmaz
po84116ypJ2ZXE6yW+t200tWUdhO2jFxY8Bp1a9hrs32dneHVRRWThV9Wm25w5JsE9ihcjDyBF6d
SJIXanSnxKXKqxQCa5g1sQO3/BOAU2DMVL/xUbJ5AIuJR5PiElgk9MaAwHDExOBsPN92OFh0LKzp
MsgX0Xqv1uTWHw4YJZ/FOqyFq+Kxel//mzpfWDAWEb3nTT/K8sgf2yW9INsXA38IlO+5/sBvYaOr
D/Vf/u0WeW+CDEULggzUh7IVwCm8AgJw6ChFe4M/X8YkCFnbpuYQ3PmROavMZIXYHGM2Z03Lmk4M
dIWEmxpYPzyfQE16XWh6zrsdqo/7t8UXYV9bcLq61B3yuC4zdu0eBeucmJ+OQQkUG86MXZcEbo7E
1SoHkbOkMaZS962osWv8DUzQHvIpbBxTHayUqPl2AH/ym6rBsId/YjdESdeNsxIjlEETyf5Yelgz
TeJQEcI/Ww0rpQexjp4Knz8hbNOOg9iswUcl4tGRbNdVwgo3RhAiU6bIH/k8FMPKchMhQAFP4gVu
poTq90uduPO/6BWlW89eeg0Rkz6O2HD2qDrOLXFiWQP/senusgdZs44+2qjER7vDO0+e7tMtGUkm
7AInokfNCxPCOqIt0xc/9vIt5sNzcRf5sxjcg/CD9EncS7CDDZJxHi2H/qWo1x4vnT5IJcct7Wgf
PKK/ZSdLUzqcEROtzLbzqnJJ0G6+Hs18eCvhnDlsjbHAxqljwD+cUXBDsJMgD+67+a5AYVL3KCVM
5BMf4Zk4fYtxUWK1SiT4wYlZtO4aAOy35WCHBzLLPU4qpdv4UbYLtyorqDmrIGDxUBhzsNAkraYc
WrfgYxfJc23EipxqlOZPSVdHjPSuH7mgOax1/gFql+Pz9IfJFTpUQ+RMNfOZRTpavkwVAwbgvwau
kcWRO1kVkLtA1iyrUfHN4e4Urb8zIciXGYGqKdTkk14hIE5KFsM0Qd+hGkj2NxO0QdkSiX6j754x
4693QNg75HW7jkfjwHXP/+5jzIJ5JcMTWoUa5di1/b4gYs4fKZLCKavyw9YORS/yWTIBiyYiySAp
dDe5Kv868APyc7XDFDnadzUaOloagnDMD/YBOHZErc3/seKBPlGP8nN1OcHxZ3d+qkjy1bW1fctx
bhAFlBYI1CFqj4AuEj53MFnpC3Evttu92+42M7zJBmOBIzkjTN0NmskO8kWbn4wBW1KUUdI9BZ+K
HV5wum6W/YkPoKLxNivxh9kzhJGB/ueNH3/YiJEmaz5mUmLzelIBtflHXh9jZgyZ4DLww381E1Fc
8lmQ3JZ19hEC+TQwabJTz/oBnm2NNMFTrfIRyXPVAe8fN4uqCVk+WYuA5HH0oGdamd+u2S78NLyk
fTdhmN6MBfOOnWWmN7YEiVRFtSgDXOsZQeZH7a6AMEql3vZcGEd2XitstkNuxShnvRwtIZyl+yZ4
v6L8pZd18512o7VZMRdnoPVahuCaX8HrL7BGGSp4DyVEEiOztR5ZMBhzc9l9sVLhSb61Ie/0Woy3
r+ojP9ivEEp3OkKxvE7Z3zzcwR4pocZqV62JDYhIUs4IEu4iowAjp61IlX8oHr9oangxwA3yBB0x
I7SXS56mH4agA9mLjOq4uA9PSyrTw0fr1JxhW98lrlqE5OBItvv6jjoefTVXvmGHauRtRIzADSD1
HecsDrSWjO82Wr55c5ESGdEYaZhaIk9cgAEL203Mfup2TTJscVpXvsNFbz1EwhjU1WrrGOTT/ndS
LhDbOBKREaDTjz60zE8XwS59zAYplSfgkvMw0z7h05lA8yZsMm/cpGii+w5OpXBG9H+2frHJVKlg
dC4rrSp1LfyPNwF2NlIb+EM4Vt8VZdeJRqElyosQ3lRR9W8zQ/wUX2awWMcbchLdWhN2TJnW6nep
E2azzhwtkRc8FMmg+PYJMe7LYdRVFrZqmXtTBcAI1SijJEu57dRjG1hIxu5KSeVcVcfGFMZf4CAe
thLfoD0kv2/alr2r2h/Sg+H2Mt8++p3Q55AUNmwbyoed5Xu5UbBog9SxwSUNP3Gv/3h9GKdhpa5K
K7ut8isux/wjhqnjVhDYytjapjJPPTC2eSDpPE3TSKIQ7lqXutsklEGzWBOLLrQipNfuMDPnkkh5
075EjqWG7E81uDxnXn/DDz6ODvXxp5TerXvUdUSyjOv10rodaa3eI9UYEWlbHnZM6EwaO+5Vq6+g
iUJDDmJqOD+kAn267SBztJOrJwaoTsG0/VuiERISLLImRnRMUwMVQRR8k9l0i1sEd79BeFvDlq+1
QasHtpOoH35CWmpfQEHqf/JH6d0T2qonbhgVkCHKF2RGtK73LyDSjaxuZ3drhoeADspQkn5Wkwxi
2sPJmpeWzYyVp8vtdTqb9t3sHPStgshW/j+RdI2iFBM1KEkO+a0fVOLPPfTX2s99D/gXPDwy6mz9
FX/OVlp4RhoSGpOJCENWA6AMjav9HImanHsgQaYxT8E9Bdt412vQCDzwtxBfnr1mS0C2rEF2AK3P
WovQWF4jlCvzSEjMlW44dIbuqbV9g+Qcj3DRDV8JQ8fYy+8xNIiY6y1zdslrP6UQAgN2348X8/mF
yeUJQfxJ1xQcANWOSSSY69r6q1YWgGfuunKW5eR8gwRGFWKKN1DrHaiQ5UslXArfzEnBgUBM1wya
r1xhmF+oQuSMWuWtnhwwpgd16G1weHKZzDRs6zuwZEhZdBsnJ9TLHd4UwgpQTOHedlQ1zKOCoGbt
1cGGuuQs4jo+2HZSS3HtNsDqQNs1rjzk0KgMwrfPfF+By+3aSuu7+n0pIBX26WjCsemDyHGhxTcA
BE+bksU5ZjGnRVWh4aUVSJI6pJlrEY9HVTEgJAk/BlS9CbJwv4FBE9wsd5fgWSoQCHZ0HjVEzsss
E9ZRaZ07OrNcHMak9vhAMX8jGM7HpXs6xkvlue0AnZq9joJ0ULNKgj67dReGnlYek3SmnLUyRIE9
eO3FeS9aMPKPYB1eYiRupILdNG61MNaRG2cJUzZdJg6yezQo4fsP1vz56zFGV54CHAbH4EagqjrH
EIbJvOj6YldQCBvfrn+/sKUDQ4lRO5J01tlk5lqQVU1nhok3/lXtWnCayKZvLFfz4KeixDslPUoo
b/M7E5/NNbLyi1dqAaQGRt3VSIAFiEQ3nEwqrJjscJWMEZGJ9lywK/A6maPxOQk07gPqZ7DOty78
ee64lDqd/LRzrUViUnmS5XONlRm+s+78clcrPSzRw7WrELpp0ukMg/hMvr+Oe2L6G3FdHWJUmwol
cmQfDd8RBo10ORKyqqlJwyPUgi20mb9HOKG6HF1WIqEvyJZM0ncMmhv3iIkVWZkr1xRBRyNjQUKU
8K93rhhQE8P3v8efItvHgQDAPdWJuLXyDxVWK3nxe3r+LanNIFQa8NjpXvhwVhATyedBxb3AWJxg
Lpd9Np6r7/ZUb9x2wtfs+6DIwj/i++ekZSt5KA2mc+Nl3nxfzxdwqmFm8yqWCydbu2au9Pn9DKQf
QQ1cpKA2jfQLUFQ6CoIv4MQJ3ihtOttcKiLSy2ON4PaCSnz/JqhoN+GKT6Um0pi/5+ynfWVTDzUK
7UYH/Rt67rBj8fgay7KxCTi0j53FGGAAUv69Gb1sScJZ5bgxYGkVxvcxmLISHIFbBg2lUcHHC1l0
DO14O5LDWUSrLyatxO0eOJ7uA4m029VYLei0uO8cz7sD+VumhYi2/vxrGE5G++/0W5FDGNgBPzL7
8vXnjLaaxGQ7MF15dnVaj2Rz94MSmiMeSt3/iYFwKaTybcyjgFUJAk2fkc/IYl0swEiHlH/gPrGM
uhukusPvP0IEigLvn5GvvNSHwQDvnSDnIz3ZXXglScyQuN8PAN8wjOePRytil9JgyECyMWMCXnd3
BPNdQVDmGX7LZZnxF0YI7Y1+tQySY8Amzp5SBPVNxyGXEcT8qj2uaDNqBvLrQsJrlq9dXbusSg4k
PyzK993YFpyezlcs/ENc9k/k9Dey7gkS5FbFz1LHzflpPaa69aK1IVycLehHYvnXHww6L5VS1j5V
udmzX33ihZRI/0VjdgYfhxKN5nPEvuEwGjf6r+9Y3t7o+22R1fTZPxGdYm+l/3neLn30gwgsc/rB
/QR1Kj4PLFJDraiFdaxPfqx8HrN9GLKtYY4hVxxj06Q5MyEkLyLCSb6eQH7NNbWTmMMla2sIT5uS
4HOskOJLerY4Hus6qz+iEVNQPtZiIy4TryfsyllHq7ss1sRL7+bOS2RNmo56T4injyfMBuOjqRcl
X6I+sgpN0JXdOwJ9JB/s53kHwqAdtb9IVKyi/s8vuZ+RomThZbyd+mVEP4xWhJbGBcbYJNsxrl6z
fsicj4zwU7PNPRWtQyhZVj1glRhU9ZPd5sF2PPPVj8QyHUO4OJ07v49jc8l6D6j7ufMoiWoiZPt4
S/SVFHp1VU9NRhzO3Xb2edCNHeH7r0tfAvU7uHmgOYFUky8xT1T/KVom6Pr4+T6mqaUCfGWX+82y
uD4p4A6mBLC9VQBz77+bCsfCVpi4qD7z4LiMA7Li8hJ1wEaqI7AXZJ4oXTYTYayrkf/V8XlMPdoU
lBu4UopFR+ArO0m6OCs+3Oxif4P0PcwkL1R3wHy/6IQgMu6k1ixSu2YbDG7E61472JQ64he2EBCS
PwNdbitGcvxEqkls+MnwJmYwnZuKjnKfMN6v1+2gPnaHwenggV76noWU90VutzuEqoTTAgmH/hqQ
QhgaIhsnuA8J4pj4UogwGvQu+JmkgYCHv+sWhcIw16URs3/pFfphXKSLJpTXH3cnNfR/WeikcU81
SEuo6j7vw8Xm5Iz9icB8DaLjBD1HBjFC+JJDpKkUU8NHglTiG4bTvNreRga3K0+MgiqFLCSe8QJU
ejRi1FSx6Vv1NL7M3QaM/ZaNIm7KiMGlJy5p61PhCA3lN9j8JJG389hRmUCodcxpenPOT2h0dGQb
Hk4tp6+k6W2jPhRkXej4ThGVv49si2NKXZbsiV66xanUHJ1QJirIo/cRU/68e2NRuTdCPe1a5hw9
QuuGpg0+SQFrBhFg6/F/ECTjSvT7aIU/OPBtVls/xJbRCqXoWZCEM9qIbDHMugXbbgQ1/akFAzn5
THAeeBniGjVfBC4YPuTo+8UTM1+dY7NNAha3ruqDDdpNxgnXkckM9yKFK4wOuPH9SmwdXAb4Rvl7
gsnlqTgri6flxvc/qmOsVu8D2wNUQHocu8GmpqSU6l/ZdOdlmAvANVSAphjIoV4BT2dCi6nwL+l9
3bRvD7aUHCgnMFz+XxvW8SVjlYUnk1xu1HpSkzUguM4ITWZdyDXbLENaM2vNscm41vxoMex47Xk4
xKCwKZUkLQ2kkbKiydN3m4J9zdMQh0odXnGvOwA84yWsj2rzGLh+WDTce9W76fMo7Sk5xTTBdQGQ
zUp474a3twvlYT6OVMQ/VgDU55BhqF8RPz1MTSqHtnrQGJaBtIXmaUuBB0wGhBpEO5J9kvwcLjC7
ghzNsTXS/ehQsV2geVWkiW2YLxahdvQgUfVi6PW8drprs77CguIsyS1Qitip2JHjMJ0y0AxGXCMb
T0SHML8lETopgjYbfPxh5MJl9udGyATvIBYYAEooyMpLQ/ex9sVnoi6RpQw6J3hffrhdLtbPw/Kh
cYD0y9MxdbHQAw3op+7Sg9MNLPFvVkcz+LE5PIROV9QtNt5a+0F0nzb25KLre4ixe3FRB/wlMsA6
GLEGwXkqNtU+StaBVyZ+4ep+BHwMbshtsPSyy7tWK+TtVFzPQGlT9MSgVaNJNs1A8HsWXcJ0kh1l
w0Tpvu/E8zW5bmxza0JtQyB50PbIYBearO/tfr27hewpa9RraHqgvSbA130M3jSKLPbqe5MK6AN2
KauTn99fj0JF5c7N7JK5jiJgRbbaWuNXCTXueUuJ4SBKB4oVTz8QDmBOVy66drmEzllWfIhC+hhh
gcgNVQJxkAOvhHN3VPmWbVxsTO4UTCbcO+EH/d+ZtUtJ0se5WBWLInr5mhIJH6X9hE8EpZitAGPO
m52ghI2P/hwN2l2AuikqZ86UK7REIj7TGX3GsuNhFNzAW4MeTDscxryhIX0fPIZdHXaA7+qq/YCT
J/GV3QF3m9sQwgdjZqVMY9NUVZug4nYpGAI1MZWUNGDLbn4W9dp7I7CVSAxklnGTWtDzaqxRYqiT
wifGl/GednZT2jjrmg0OfUDT4yXxvy95JcL++szWk4jHDi3lgcVWGi6fCJjYdDyoMfGUzBi4/cz2
kZcsDdAstroeM1pX/UKjQjIW3werry5T9Krnc9hvmw42acl8P8MCtBibaRq5esXsuJeN5W+1BhtN
6l28xQhMQA4KJghj+5mX8UJ3unaNRLDCGjSyLKAFB/HzRqTImhmYnFYqA3Ovo21+qw0s1hPp7CFf
6BEjzeHziEcvwRKRSMgWVCceOoVHZcdSUCOWuF8Sn9Eyvjk9ZIiFTqtAA+6qqLOSPUGwTTB1X2n+
Al20vSlY/tbJdMkJ99XaTKzIMdJiOvYq8uKSBizSv1IbOOS/Md6f1y2krvs1fzmDHynUTrirD/w8
eCtiEPjhlIbQf3ZSsqBT6EFO3AmILFvTx0xjmaw5mKAl4oj4v8lR4Nuy57qjhvhCPtWFs3cN1Nvs
xQp6+ZaigxOIBeVxgcm9bt56O+f/z8ijvTlJC79Ul8zRuuQa601PEzZnwmTlN5n3beZ7Qb9fVMRn
ywTAtJ1m50tjunk9yrpneYk57C6Qk0WCUkiEUrKiUpQRJxq2K5FzB2W7M4gjP96dT/Z0G1WVy9Kg
5xviL9gG373vMsrY0xAcP4wxhQYkpZxzoNRjYMtLOTEFML8F/G76D9BvZAhvVEPyS6I4V/7aERZt
hmxgTBDCNfuYl5leCE1PqDs3ALvSA9/YMlhTlV1qN+9ovtNO7KHbVlKTSOcg+M+zuh/X5Aizc6Hb
8tNZkk0SfHP6W2F7OxdxkBCft5YNNSKlzc8OYAg52yuUIUwklHv1jEUUXMZY+ZcrS7jfawbSK7GC
jSY80p9k5pFjYsy91ELdVHQaplgwRYOUEmNxE2MCAHhE/boKOW+9s2Ypty/dDl1qjygoGNbgv6Ic
4h0H+0iKDYInbnDmdPlll5yAGWFm8dm/nDyJQy7a5cv9jdHd66C983woxhm6ahegJ8/aqGnx4iea
bohojnKpF6BPbBGYQMKEFxBA0XOcJhqcJsXtvu2kvLLLOI2Y6EPmsVLNlSEgMa5EKp1H0r0vUIx8
HLGN3Cnm+ShAKvfoURf4YO1+yrD+WkCvoweWVullkPwY9yiRJrnC9ZHousnt+95Jto9yardJWSah
CRhXCWyrr3ec0JVpstd9exS3mT32OI6z/I1FJCKlWuoDgDb5B/wj/upGmgwhx56pw8MEtkYc83LC
2RaOVJMs4v4bqjwn2FQZcKA8aYTOSRMVgj05EhlJYv9qkO/qEFX3kpqRahnACUt1IbM/bH5/Mj2D
kdhqM8DyTgoT2q7i5SDbjjCcA9sPMTInWavo4x6rjmGKevwdaRR7DQhLWdJuzKaKjOHufzF/++Zk
Hip7aI8mOLcgdD9/eFx5zg+3CuZCjdmhiTS+4X4O8OuDjJrW9VjXwdiJD5XUDB7UQ4eHmuIL6q/o
kbgHcSPgJ3tD2Kr9R0hx7ZWYPhdBrHEkIVIkD+zwYmM2m9mXin3AoniOjf+7X9cuap541oWx6qIl
bxnfI+gJbY9GH2g4J1rJjkkbWB/YGZb9bz1Q22nkLxuMlfy3k4yVObtJcR4qCS3hEMRB67Q5ZwHf
HBYW2zP6p4Lik/10Ad+vZH75B6u1J/QqudQnunCEtcbnJhwQwKAGJGyyHzRqxWqt46aA9EgLk/I+
WZDmx9Bd+4iY9Sk0Li1nL4zNCJ0EPTHuhYKmMrACUKPs4Y9CcgtnVOP6mkTVlvX7nTSKRhTC64k+
l7XuNaBIi3L8jdhudyQw0H+eXuZVFyX66eAG76M+oymSUM3cqF4AUmTZwKHQ6itPVdOe4myC2us7
GDZzvxge9+2VGkl6WuPw/EJ/mg69zVjCwLZlGEYgoqmOPDFZoOU4BJ1zhg0sqJTZf0Es1pKGuWE3
GG5qvqS3yKbTvnCCB5Ri2XxE+zpXfbWv0Jyt8y9nCzfhiRHHFNm0EW4j7IxlRtt8jqo8UUjwEJHU
TsXe5k42CVpQgKdIFHQywqZ3JX5u7HJnqq867oHHDc1I5dc5Sh5mjRCqYvaMt1QoOBiGoZAmZPOk
lf9lr0H98FUYKnfOiKBWsaiQaZM2XbQDnCGg4BHl6jq5JLa+xJqDDlUAPJ/9VYA4YopWWeVwewtL
YlSJY8Wq8ee6wa0Vwqje55ettjv4xfUq3WjGTt1vhqmrtI2P4CmmDm3V0rD0EnjujMG/cdswblHB
wEK//fIDpabggSt96GuNoDiuWLIHQxXaCvAOdeBwKEbiFa/W8D8feEDaFy6IHPb9jO0w3Zk9u2G6
03+bEOYfcwQdfjrI65GKGiQZddg/xmaE7gt/4otABxnU7dp6iufc8H9tbv+mNhrjVgsU3qNEB3GL
TxzJv2nF+TAd/bKqBc2VGLiWVZhnat/FMKSW3nqXhMbSHMgbmVIsDbWZU62TgLWzLrqWVqengP92
tQU1nbG5nnDjnp2COhX7Pwk5F7h0HUNrFFEIzxFcPO3uXRo00quRUzw75VMjtMlYz6d8AWQeTFqj
7pKdM4aX+ph9vOfIQAyJPRFWox+KKH6MGV+/HhNbOCxxMWMVWFBO1FMo0MyqEoNW79egGzhj2JNT
4y6vAZDbZ3ShYn2qMyjTc7fihtExyqJn7af9T2KK31/0Sju4gIG+hJVvNgk/wXjnN+TPUjnsp3k7
MvI29x99Tt2IhE2VDHiaLtG986D2USPjVDnaxdNJ+sEiCHNqEqqUaCumLs4vIgZ9/h2hI+VehXYY
ZfhYn1LVU8cVsoirccWqZAbvGaMJXgmbA6TOvAj5tpVFmkQdb7TF1vrDq1xE0RX4CjxjMc0kbQtg
6uUdMkY5oRcWuW48N37qYUibbZDmZb9nQrvAkRpXqm5m15Jje8b3lnyMwhAL2Srt0061xWLDR//U
+nKdghT9o6Hxy50kuBDadQR/aGNL3oaHt5qY6CF9RQa2tro/7Ptp9Godp7htGSnwJ00iRPqGnpJH
SbjwKJWLIyBNUDxuIPGVqwRlIEZrV0c32D87sICeHubKkhKXY3BZxE2ZWMuUchFPMvITadZOk74l
k3N3Y3h9KnwY7nMQGytTUahGKmKyO7KM1f9bO9AeyscXEppUY9KfVrEAhoLd0iabTO7GCRd5P+bT
eViRK65/ghB3yIY4dWEwwd0m3FkXkm3uHjYnthVzzHQaiQHm+io33R8yQTj8ASOO4xCzSnAe4LO6
oV6lldsea+68phDfd+74zSMjnjTUTTZml/gBNqYC/6NCbbQ7q8GD2oKz/sJ26zDYg7ZP4iToU+DQ
eCok+MMEwHO57So+NILlRzLzJEbHKn960rKZpSL7cN2VYfD4HaBeO/gMOy4k4tMOUuaSFtU7C6Vv
x/+c2H29KcuctzRAbmD6YsV/Lk4rbaO2tQTrX+aOhArTbyI3F/ZHG8VkXMcP+GvxWu2GsWHlRplv
0fOHDakL061s+Zrbk6jmKjRsCZK/7Q2E18z++QSnHNcyeqCpNPhPGJsePKVgd/ROlUDuYGyul14O
+q4m73QNSVLPaR18YGVKE2uYuGMP2VdsLYT5nEVGXb4dIF1SnrOyt2cDYnGloYgtOzMsvZREngWs
k7LgH0vl+2E7vCzKccUI+MXxR3LLomvPHwJXSpO6nEYsA6Xwy/VllnGndM6a7zeeyYkLMiXDM76A
JqCABPu/0UGfipN1lP8cA/zXDfi9thznejGfwWllsAANVHCrOt1L4qGaWZlVTqwWiqvhjVc3eqSU
ze4Xg5tDpt1Kv03L2uEoG/sDP2g1U68fUlBq9MYIsUXa6JaOPHKeUYZS+mt9r10LWHNfqCP6qv1s
yyJZmxD3Qz3mH8yoQRegTOTQNjeKAv5K8x9e3SODqFYrLRyukhS7YKcKQU5Ab6GMwTj6Yz0vXGa+
ushzmTkU+xzv4srFJW1myU4OuBCsS0r+B/pGXo5tp/2UsKywh8ySnRtBZjy7yxmBEtISCxubBWtL
SKkDe1jEy2OXGggCAvuQj932gr51+rTQ+GedwVNj50ihfd5YUGi1Yoq7P/CeOm+AZHRMW73HIoJr
jo6coZkohQzh8sCST772NJtoPoD0PHc9QkJrwm1Uk3E2mlCCKfe6ZqjJAiNGD2GHO4adOB01TQJB
gpyYVbss4TC+NIYmeBLEuGDpF1mXxvIQa3Uv0x2D9OQfJnZmLvF2rJa763sNbRjjqru0cGrqAr+7
ZNa3+LO1GgAggTRMlDsVWyebyzk5cxrQVFd2Ag0cTCDz6CwG/WyA1bj1WsTN0rzF64aG21Mw+KhB
JdxsRqplLM9JfVow8DC/e1tDhEfS8VACUnEC17fGJCTosigXRPDBZpaU7yNk0VM5+IuK577uTK2k
t6o3A7onkXdRdMOtHT/5YSH7ypjsO2/Y8GhMIWPN2qPn8C/+scCdNajBTilYIvX82YjjpDi7rShT
aLkIbqVco/oJT77wIFNZvxzkRU1syMx1viQDUBIUKLKtOoWMDHHkmB0phYQRr9MnXoGl4Bilmk94
sSQiuCykj+xOZl1KdysxIj72c/uVhPk3Je01KD8BHivUgq1Gi4h1K7hpBcx4jOABMf4uRKot97En
SD1hZPFHNUmgQ9f+bwqhw3ArE4d/ZcuVramh3q8D8e7dVCC0M1Ec2xBfJFj3clOoBTDI0JaFqkhJ
pi1KYgTtoxTdOV07PdhgfEtOdQqLJ3554XxNOxE0rPa/43mADQCtotvXa2Eyyh7JPezjbE9K6Wsn
gfOhE5WozHvA9iwpptWlXKKUrCmqtvJZYaTXaKwy5Xb3+/TKzUZsj4q4+RkdNiXqoR23bkqQ3Uh2
JJuStJKs7WMw23PWd/+aLbErUg/vZFZa3l4PAwLi9A/QOT+Z5w4FLx59eubHELPqUpG8uBjDaJjN
sjheqhHYhpaDw9vNZMTUFOY+0SUYueTbmCvvZPam50PPFQrPHlzhvg0IhxCImnwmfTovcx+p1Cfp
i/vcfFZy7/p5kYBhpRUTi40GULLA2kvYD/cDa/IYPsmQyK10pyOO1URJ3d1hA7WGTCU6Ym67/hlL
bfErNi4S5WxSY6uGUOCuvMv3kclCW5zM4Rfm5dmVDsb8O68jUUunjXnPGlW+7xx0MvsKroIIjY2T
7KFnGeuECJDWDRqohEoVVBrpRl6GBy6x3VcE00WImwqPuNHpH8wyjyeN3zjkhO/ZlSs3JdxZH/UH
nrdpSZk7/jb2NcXj95r2/7EuD4nQu4rU1qeer9qQqVEIKwyOKJ8cPDwGBH95xIZJjFl7lld9KsFB
qVgshdRZvIFbOAKl/o2F9J75YRnzTTWd4UD/f7ap1ItoMBNyVTaVDiGl83UP1l/JasvKnDKiitBK
ZXJYLk+bXEs+kd67Qxc1I1aBkTgdYZ9DFKIiun1A2R45kV520LbIva9VEuPEWS19fwYNoVRpo5GB
EnbtPMs1NznXZbQ0ttXxTqvLq8sad5SPw9Bt1pS3ncwAy/2p8Ov36XFEACQeUuaXEm8Pb/P1LeM5
ocJAlWtyfqoWVIbpwYgZ4W2n3irQg1wFMDgwcv90XPpBHbzlzm3Bcq5VIra9bZxYftpZADO21YHe
f5RVwE3P+vila702Ec0Yna3+yTCDa3iKoLGZThmZtfQFoxVinou4wFwq1t+5dZzSvCkLnYfT6WxB
UE8/WwPxV6axE2Dip/XXWtvSsK+rSM9or0/GCdSpq+3pJLyk6YK1dBQgjabX5A7eFPB5P4h21BIY
D4gwl13i2L4/C5+agNtCJ8bK0CPZUNQMK1L5qvHmZRZueBoZpOgpFH3m6R+mvKezdOcwGdiQSvdS
l2MFb8Yh1yTE8D9gX3pAh04zqNHta9iOntwXNazt23fHcqrH4aQP4Osrh2/EJa1KfU/HAM2L0L/W
4ubWHBPAkbsp+a0jQ9mcGQwcmdVJIi73sD0uc1rmrsiH6k30wOwdy+UzF4dMctqaCFloZOxKnr9+
o8QVriEJ4k/OTH+k+tLL8LEndrC2NsvwNQBNl6GLl5IcfvVdI0VrKPQG7PvQf39YPBedXZg/OUCi
Ae3DejwjtNvrNNnyUTBqSc1r0cldqnGlxD2M9W0fwrMDGn55DPPzNyZzZmtv+GM3Ng1mKffcD3Xe
BwpQGG7Y2TB4jwAWuhunsI+DeFbBi4HgoLM6rT1mUE3Ygpfk68k+UvTguCEy8gJ3wmppKBaZxIRw
cVcBX6K3u4k7387F3zylHCYlyM75JZEG7ZdpoAl1IoXUw7p8cBsqV3QsWhCZelUPvTbmgbI3Sm8k
WTZrD+6Exity9dFmOY1eEQ9PJc0YFc85429n6isn+2IZZSMPgtrVSaLHq6CQ37nEJe8vu+Bs50oR
YwjFrbdLXB0ZJGWdxaMOBbY7RRZMvQEfSHX0z5G7dA1nUhUperuE1jLKb3VoCoheMhd49kwDiaTn
VbuLefYCnykrQOVqHM4BzohVOdhjprQ6rXsHESb+CimHw1fRUu6QDzBmvggzl67u8iB245kwNaIl
Gj0f+DOgV2nd3yQSpYTUFyRD5mNV5EzpmP56W8E/6sVTfiSzQ/ouw/4WPuMGZcBMKgU0o3yq9Bve
x6zeGEFbIPjDJE8ls83wvvyoUhcZFs//Etbm+ZOvaE6luN/NsbcT9OR3HzUWYizWMRm52M9Wkdx9
dEdim/mlRtDRjNJpvP3v0WUTX5xOYZiEMm+vgneQwD9j3MU8nPqLKTpUhhEdc7rWVcQsDwdOd6pt
KQOnEyyxS0vHp0KsqsGA6MloBXGQUb8F242L+hO29SGOU3N/bIfx7EWIW0Cyn+s82JSwGYCLdLbe
NRgidwy2eBlyeO/gNSdkxsrG93oDq5qHcv0VQnyqGnsmVEFtVL3lE8xiMWV6iiEN6JkjsubMTAvu
onTCLLS3KjpYcC2Sp4cZpiXocnE4osQmtlHDj39nSdJtvATZHHRs17nGHGyPtYsliEWDoeSf6n76
YVCZ78mP70dwujHw+hnR/G2CoXNakSMKN6H9+SDuerq+uwqkhK56SeABTZTB1YwoE1jO1Au2xkDB
qr21Nhg5Wb+dCCTvwXY0p6tiqKAlgD4YKG4QkMP54rg5PZPRDwYJFbPRWKJpcw6Jx0967WKWs3ea
11yunGmT9RwW2YXtTdpKiTOxcSU57wnQW15QbyyK9w3wfxDzti5YeEzAYPxWUwwxOM11uLybZX3G
GAdpDhPSgc0+iV4j6CiWgLuKD9tyFrxN8a0o1H4zo3xam4+jWXif111xopoLPnZlJaADSelVJaUU
pi/1SmDl8kuX1jW+SjOllXGJBhkKxPhZLBXFAhjXy3ncepxm2uE5GMG65iBD3qt5OV1lYxrmDXcD
5uUA0SVCJs6tumy5Kfj0astxXmqx+toXbE57fL3T2gz4ZarTMrLVfEQJmFujxdMZ3SiVw2W+sGqn
LJqEe66tpmzXnmxwpMR276J69lwrsg/KzD7nTgcLsdQWKAaFqw2tlYS+ijSvpRjQ+M1QX7y2tRGz
V5+GyYeiFsl0zU7G7c3wladaYrIAT7uTg8dPbVExjj/qIjDeUm5RNv/anR1FbEg4FetG8Icp6CRG
cvg2DyRnq5I8f/NP3A8uV4NcajLkcaq49vs81S/7386YCOq4Jf9POgp8nE2L/CdWaycOIbcamz2V
ZxkULzXqfrFMaxnwiItcjsDuShreHOI9f022zy1612yHGqnEVQghCnnseCbfPhkD61JqaCOdUKs8
d5WeAlAh1rN8zVSRW9nHqLBnWRs7X1C/4tKaPblEyiQruRYdQl0SYiJB2cQi5KG1iRkoQE8/s7aV
U8O3G2P8oYg1VBamJopu6/FSoGQnOMX0knBQ7M4c5skBxT4sLJ+4WsW1tMdXbJas8+W+oWqtpzZf
j2FOdOgdp89Yg0v35OqHm4v/+hYVUWL8jEAqcCUJLDt9ICnChMsLTNXdemAT2CRpy4QEjVK6gYy3
hetO9/fmlJ/udelriDZuI+hDUdCNm1o3ebUpwQQx8cfJJXhO4IHh5u1bRuEpqWCRG2ctCCiSwJ1n
RDh12MU4QBOLo6K6UjZOCCU/6DFV6NsCjb5ceQW7Gbj/zjqoYKOPVp9a64ldGAt4jXEMsuQoCvTB
o7jaBbDOKMCSrDYrybwE3QIMFHcOE6Bmci/UijnQiF/f2FUfkA655m/kTQDXVRlCq3ARQWNP6p2z
EMfIs15NJSX7v4rdqHRlBBeec8EMSb0QEmdQ/nuknJZB48yild2IDffJ646aTrsNwVNV4IWD4whb
XnMDeqWCF4QI6w3akTKz2V64yijjaPNA2xberpgCgzEdNaO8cXgQV9IW6vTuxGxy4ItmlT+mH95e
+o4rv8Xkj1w1PoveYPCN4dPQnz5H8Xz079kONeF86N3V0VPd1SqPNo4TDJ93rYY2+4suH0oMx5QE
oTZp6DBiF+ik50Te/UeT9w2E7SmeJXt3un8lis1bV9Aor/k4aNcM6sjVXOcnxwBFguoJFvuE2gMP
1m/WGUHLeadIaQmNnnPqTQC6Vmnpe7GjaYr76iKmeWfe4QBqFIkpPf7Dbni6XWiVHkBXsiSa044z
9W/L4FgdLLX2QSsVstv8QTgvNT933DCzFL4wZOaIpaF3TuDwvhTAziw16glNlF5o5vfRRcNnco2m
HksJAHEhWTqQeQwhgYS8j+Lhil8kya/PFiBmCh8opiZTV+Ze8QzWXxuvjHnKAXPAZTr1yFUVegzu
8GBrsll4UwJtSA8To39PGa0PeDgH9Uc+jCEIccYFJNYTky/yeJ10oMtSKcXEEfBskF2yVY7q9kLz
i+KV6UrgLcuF4zLYt24uCMh/tibu58a4I85JUZvg2YX9DP8kqohLLyurWDl/NREg0x4Na2aA2RIH
Nci/rnow1us5svztSpOZ8CfT2ANBlDN5crExUN1c1zIhP/DNJRszGhIXJlowXpnccYSFbLSNCSsY
7LvxJ+Oa+nt20vddLWSE1Cv7BZZpWpSIIgBiVzBho+we1Fkx8CHoe5ejyU1vwQMNu/Xf1MTDSkEx
3Oja39QCG/+THumjJEaTGEb8uD5H0nDiBh+Ph3Wj/i0AApaBuxsiq9/wTZ05Nuya4OsiaMLlB6TU
zLCfcnxTz6q0hJtpZZbcWhkmpQfYyWhd2XQlum9Edze+tblOHQkTFYaGfkbOFkPkUAx6/IoO8UmK
A6fTV8o978zDlnrxdPveDAPKk02d2mSO6x/OXknNrNradDSxtVLqhdirZvqVHlzYMbdSQLc66YOC
gzJKDKZKpbre+n2H275J6/bQcQXRQb8gjxa74vBDkydMKcw2ssnfApBxA3FHdEy0BwCV8v9sTg8R
DjAhJ1nogKMOG4ADtVIE8uthcRIWDQXlKntnJsjvc3fnHsPZJ6Hk996F6ak7bWDoLYBG3GDKz45q
ncM/wcMFi5U1LW/aWmRMnY2Nmv9evbspqq/SlTiGXYcLY4I1dx7AlxQwcpLn1mLHG5D7NrZ6fiaT
2SwbeqIFcqrdL+tk/+RoplXX2Le3+FHkzQKAqEtF6EZtqtoJx9WBawoKc/ol57Qdp75+PRCeY6Bg
fM3PtuJa8AiSqeB/pacdSrsvB9vyPxqm0zErPfyGFgMqwr2OgvWluZgjamCCc1ZwnesKXt16VGoQ
7yPoOt1EoGjaUBtHZtqrk5E3oQGfeRBnFb6SDtPKgXjHdom26IQF9bPnorO7PgEy9oxwQarRFmtp
srE3oWqE+C6pSFiMSRxnX6G0ihOv+RpuA4xwgoTEfiPANLchW7CapW4T2tKzhg11qmqwwBo2Yrs8
nYGEvqDhI0+hx78bIUFyfquXrHpWZc/V85xgpZgRK4wkIGS5IoSpxwXCWsW/QrN70saK/dEqJJLW
7/7YkP08OxKC1Mrlmw40xIclSya13NbZ3+x9lr6cYxSIMsTLNLxGu2jdVHp7Swpe9CX2oYn56L3I
7IFBt1spgXEXXIzV6yJHIPmcLncM88On5bUUGrKIPRAuj8IEeD5YVB6qSEP3enOioC/nfnMvJH0k
jCxh4Y1TVCIwK+6tUrmtSQOqtKJkF9Tj51NdoCSn89cdG3xjAwy2X7ykkjAGUIUx70xqOpRMzU6Z
0qQ2LxyzNmseIKFkXCgt59ZJBYqy5nfc8SJQx5qz8Sc2j51CXXhp6l3MfpC7kDDoYRcXIVIOxfWm
5ZITDGoaMuHxLEGOW9VJQOKZ5zwfNPGUNCH+PQiaVhHJtKjSmmOfDygVhJaPiQKd+F6cw2m4nxu3
sk6tIShPbeGW/NBkxBlLKGRKaheRqHtT9/ML6UJY4KzfCfP89UQvXaMEKbN3p58ZO0UpA6eD5+Q6
6Tnp9NjcjdHOcB//nAmPkjsjVjgEKQN8rleuebSgugN214c47NG/YrEgalpWPq+TtxKx1gxal7R8
2Cp5LoJP/TbpsvO5Xqmqpvf9eLfAIc7B+yiA1fK09NwpFbUp5zTTP+nZ6PUEvZPMKuuiqUmei273
9OHzqN9xqFeBtUzaJQ9eWiNMnTT0VF8nhFOvyyDrSmzYSaihWZsKYh6OGfJ8KtQ2fF6Z6w52RkCp
SrauGl9/hPUA/HHPAIyL7iZCsvgaH7i19JFEFh06hV8xTrBr5y4VzcyAeG/pPdiY8B1Xml+b1uQY
ZQUujiYnGvOmoK6SxoC+eQWS3CZyNtrb0LRd/I7+gDvBzEm4e4yYURKuIHq2c3W2vxpTRvilF2LO
JISyD4rmiZdJN1Suf/tDh9lpHNmT6AI1yhsNsMefWVUXlj7fiDEuyPqp2QjpPc45+Wb1VFZTqi+s
0cEk+T/59LeFfpMbbPxYVh/UAF6JCYVZz3EHLZeWhhGo47WMrCvzRj4y5SIIh7fF0y6AiwuODXB2
FV2cM2DBOHopqBjApPi/f7bgEJlaekOkzcpHYi01QENhYSi8+4lA6rrTzOkn5KVJGF+FkXaRArjT
gPXIHaQYXAAKedfApDoVXrWg+mBh664heokCBnmho5BC/fBG2HFNK1r7j/iGRksmujc7hqGcKvNM
3EcNc4xSrhMYRo4e8x/MUnGpRAJG4Jsp5TILduUNElvHj74R7TRK62X9e7fyTU+W/6cYr8Q5DGC2
AzV722LWYoTVdDxkkFgWOJ+xfJ7TT93kxvMqOgFXSZ3U3SYQC8nABPvnbaqxj4m+g1ZnaXWAHxGt
D1IyWI61rSFcGuzHduO0krMpeAWaiWIyOsIxBfmb4z8eWSR6XSpRZQnoJ4yl8PCITqMatm7MzoMJ
zSNGZmjnvN2QZ3QyIbPx6xytTlfHUQTWpXFJnRipk0fw+m72xvNS4gf59tTr45AXjccQg20Wzpcd
2PnuhN9UnILarp2RY+2vSoh8hKhkrnrdYZdSWiDyH5SftD/wy5n0xQeZJbNkwFxsQeHFFa695ij2
SoqOHN+Dk71bI83Z3XPNErvxkjONm+QJy5fRdyRLl23rol5A44Mqig/SSaoPlYapTIlFzw8TrWbu
8tEfi7CITA8ARv3t+TRRPseJZUE96z12CetxAY7LPbxbj7wgnfPBkgIEQKBYurW0GWg2uetz9A6E
2LGHhyC7QsnneJvea8xJUt9SOAQqYlnF/Qdhz7olQOS2Rpm6HWO3qjUEm9INzBosb+uFEdLoF1yL
dw7u0stfhxyvd9AjdTEIjMUpZHrO36lOuRCifISI2Pask0wyrhq0saqxMBMBsm5sq+5e5i4ptRal
/tas63S61J7vD7drED+JUYhQhNYfCxi8y6V1lj0DWy9jEXZMDrXieir8byvhNmRj8OQDfwNeXJoF
RZ6Wq4FNqLFM99VSvzIg69TQFpaTItEx79JfOcIwrqn6rXfTKHeBvfTPZyac5Bi+GUaYnUu/AOAV
IOQNg/FNk2PStCwI3rZVkwhNeptX+4I2ZQTeBaYx+VOEvg7qQxJtRaKS6JP9VdY/0BL4GfIRddH7
TfkpLSZomVcmFEYb+4xHJx3ut3IDVMcvqn09Mw2UiXWiaMdms+DznovhBhC2jhqb4yi/tDHmm4OG
JH50hxBV5ytttUpK7HDl5tJqDwBHSlVN1C2caZmrT6AldnS0n3e20MFQsB7GzTMHQPpvNmwgwLdg
Lp+TJRVZAVDvTygDVLDpcK5TtlDILZNqw80nOnFjqVWis9hGr6tESO07uk/hwmha86Nt+STMpETb
LyA8bttgy8nKam6jNfzDCAQ5nBa8F10nMHs7L+2QTom9xwPl79EaJ4dhNzutpBfRKlVIT8Bn7Nn1
bBvQte0/pRDY7pm1z5sAoqLjlcOIW8gBgfuXcRSoTVzOrOahb2/4gGmLRxyEEFFHfUEF8Prgpfzl
98rdcz1hPicChyGXYZLighEzgysUu7GkDnmVL1/40raiz4njKAhya0/howH1ukLgE8qXa7puIF+k
30xEPHiGDI3NQPqHldx5fG+mXtwTl/qGOjQH26AionvoTrjQVb+bQXhWem5oIeVdeRUQfWAPZgLJ
oQD2PQR96lfT+pXABDVl+I2kdrTtJ8Ue55clJzDZbcI0MXFwlKvaVhEX9IrwevPV/DNZF/GMgmXj
UMb0cZepl/pMc1II4nPbNT/bErVJCDEUXCeGAjHVkcDxjh+traL2QDKYmEuF+rLEjY/I4vNENUgc
HROKzZ/4U2UWU/M2EMij9PQw9GCuINaugssXCJKVkyCBn9ZlTOh4J/3ZpGBbRpkv7LNLog5RyPDv
eXNnZU25vIRV3WInFL25sN1gKu/4uCYbeO8AVSMZIbr4cfTJ2YUDonPauaXoHqffmRqjHx/fgW7M
vypl8kB8HZ8ecg0/hzno7+1+dMmsIOnPLbUoEU+TsK6jzdNqBr8bKRDuVk2tBURJtNoRn5qg8+Os
cVd8ECddZi22oNFpX8OTG8/YNEwWRUEpeXlYx+yFf0t0ZWYrQ37B74GgOTUPoLFeToRkiLQpWXDh
BE6Sff2InaXF87OS17A2gDag77BOcES3m+FcK9fjZIiX3TXLA/Cy/J/inKtMRhh1cfsNlXAmyqOW
YbCUteJ1Xmkr5F1EFzOPdL8GU6Wfl1bj3r6XE7r993YfYlMr4BBKInQNwCE/cRywTlhSt1nsII73
lWU5mGMwnvh5rqEYrGB2LFqvPh8338dE6gA0Zv5PFAnz0D2I3xDG1YO62jYtKgHMD9TZQSHFwhyc
IYct5t8L5arZExqYYjMuSNzKydcqxPeYa39PEiiDj5n1XBtWrx8o1RpptTYN+gJziA+MnFuF/kyX
c99KncrDsTJLuxfj2cekpyqMFPDI7prC6mmjMpyZ2ibru1nu3hIUbwCDwYHSf2F4PbcXhT0B5xol
j/z62QsIJVMRvI2+nYxnFqjxDubyDpBlqr8NxdPNMOQxegG52uk2TagG6bKHoliTdupa3ioT3U8l
mp+V91Zc7ehCZOedsyIXJJBV9kZ4wXpExpo7igYrxIQeQJ+Egjy9Nwo+0/TZeQKoj3Gf4IEKYZx4
W3w+nUEpf4tX4UYvFWv2YBJeUogSzemK7Pqeb0Qk6RnBCjslfJ0+zoGrOndhLqQawPBaHV5/Fz3p
z3sbdd9dREOmCbVlCMOPz2PAxK1S1xj4MdzTr9N1Nw4Qphdt8e9S7A02iauwjeqDxK+lyl60zMwG
WnZ3Yd3jTyYO7LRw0+6DtBeY3Sf1gKSdwsDyB3o8aEa0B+TKaE3xeCXa5m5VWil1QklQr8TkjluS
+Vu8eoiGURli9QR2x1lZi82h3vQ6iDml+sUpqTi5LHkjPPDVyVQ3DKgm461FWEf1qtUZ8iFUnfUU
YE9/mYi7ojqbLNWYikH2nfESPRldGkFuSTE7bNo3RdVIm+czRmaYPKGbRYKtM4X7SZvS8oWjv+6y
47KQ422nxJEH0sIJxNLMeY+jBOjQ5/qgiDiiH0hGJMDJCuQxNgHuw5WNaNUFKj/YEkuf3PAUAIqJ
n1X5cmqUOwTrkSkchLAaw09zkRtYlUZVkdb7mmK9gFVBp1ZexBaMtXN2MS976IethYuIFledwxx9
Okd0DjMUkhPjM1/uNQpo0udssO+1U1VWkfsoc1PW7AMPXRgO0BwXRm1OxBOCsKObhjR+vT63o2Xf
QO0HKBq5Htr4UciCckQiYmhhTntZLK3SYXQClL8TYndSiZgQzTExwdXNtkdEDTxEPqOCXNHRcVP/
0hCTXr6bCJ9CyZcbs38KMiB/bZL1Y93PMm0qvY11LJHng+16Ilm0NFBQBbNyUK3494a4MAKGT0sA
TP3V6iGqOozb0YcO5k6U5dvqGStVPyvEQVJxaMa0+kQRhPoR5gsc/y78roMkNWMjc8bAJBa7jAm/
0Qz1MBpEuEu/eFmTVyBN5Nhui1xHzOPuQn+zpOWi/hixxo8LHwCAr5Jqw5/lq8kyjaTzcqcRK9/D
jBhXsulEcxe229FQVK0qU9L427pe0XQuVVBS9uDIAE8vE2b/tcfnLkCIoAcUuJRFgLN/r/A1eXqt
HcFP13bLR3bobXSN5Onxt01rpXtEKFm2Gj+1+dDOee26p4TfoHz4oBC7O+6eBsLbZ170bSMjniYJ
MFIgWFTfrCA9i2vgCvF66H3zGnNBekght1xwj3yoHHyOBD3FWijtFFtecOIKzJop5x3pHfQ5gMUe
J52XrJt9QirF9WxQ6gjaojM+XSTLzGk3l2XhoX3lokOzhGJeJxbhkfTuCLz4NwZIDPAOh+cSxVxq
BlbJAQcVnqieKvR2v+aLn3E/dX54VEjJ530vk3X3Q1W9W6RQ4K9p83kV+hcAUuy5hYO6rnomdAbG
CG3pln99sCZE+nIk+sTJF0X+c3+kZkpkJNubyNEk+4JvfO7/Qqbv+6RiMGhemLAk37YQ3Tuynw0l
K9KHsjDJkQdMtda502CCDyKd884fQzzNmSPb7R/AqlJ5hlPjkrnzziln53GoKH1HVq5ii70Utj97
CtSeO+LBrYAvfVnfTix6jlDg8yyxvVoudfE+Ct1PCWMqeIangJFrMnRFYCW5yQ533NjNFEHCUtD4
sWDQUOVvCayyvtGyHPmJxPHK6lHg6aGBAmq3mKBozY5P+88dXoAeGJOJfLf9QT96A+Hj2C/yg+WL
oPs0h7KsJlB06hl8dFSNg/LoatPixetIQ0hqCRoQt2qxTANIIKzIlX466yZ3FF2Q8z6+VDHBYbTa
tfLKXwl2f2DTSL3vVllhtEP3f8R5uxC+Dmm6nQXTHv7drU1Ikjjd897I36RQ6guTP8GSOv2ZxS0/
3lj5ilDZwoNtPw3velgGhMdg3Y1lJabRgpcEiUEzcpeLBmzlCX91wqp8pm5ELGu4gk5twQSQVdNf
xAe/zT6k43lYx2dz+G+m7lfszGKGhMJZj6vl9LXuIkQniFzkbVp+rKDI+vjvXk6PUvgMJ36I0Tu5
/cm3M1g8FGpuHQwHoA2x28sus1bcEy06ENJmMCeJjQ3vuoDnn60fjSa8g/qafX2gVJ2nxkjla9TB
OU9yhb6J14byKJBiWpylBkRxUNXCtm44NsP/F1+fPncyyxsA/KBs8PmwLNEsle8oQV/mgmh7I+t3
91l+w+2qSBPw+bC+Q3eZfbyiGSBDSEmOU3MOTWZlmC4LO3TmMKyxoohletzt6W8IQTjA2UnT52pF
GEjL3ZIXty6VoAE4t2G5qt7dEqhP4tEcvBFsLTSvkfGZgKCI9J2kW2QElTf8TYQTBWqRffX/Cm7J
X1k3p7hmbnxCE1mKE+rBEzed4+UB9qD7qP7lN4IqOTR9QCiI5EXAlCR1jd+OxSNw4hGg6bWnMwia
l6Al43faGArsImVAqBo/hX5q0SIU/lS+pVtZ0o9Vx1T4rb1ouOdUvITFhGCYQrzmdK+EXZgp3hRU
qRbDR/+iUoVcz6k/g1C+DhJiEqAnq2iB+5W2akLD2VaDJOwFsIM3KAJCrULdxpejGGTABJoFpRir
ZA7ye4TZ8cXLkRI3YaLN/qSEljzPBPuc3FEf8OrrvPFRJtg/hgr2v1GsJoPtnJwbHxTbQqKyxbNv
VtVmHD4GDIKfMwT2EoaQh03thDN4MlaiZ75geBlhIB+lhuCdaOlpc+zqow78/Rcpav5rv80ru38J
smM1Uu2FDeIj29MBqLZq7xKtQ9VXbhLaECOgXzbzibz0ceFnr2Lwv29x7QThQ0LOEPtAgYmG462A
qNV52MQ6C1dCXoLJlLsMfyC/ASjBV3UUY4aJWPTIfZFjoeKDpySc3yAF66YoiPuJvEO3r9NP6guk
XBPkol/UQLXVv3MK2oe7O0M3133y2lTSDrsmTYiSiYqq9rWko2YfBpPKNDbbglHL3hsA0v4d05Or
9qoBIYFrIv8G87nRV/vclRpEEkR3EKPPU4dMACbkMJxTC/vuAxgXmjZY8oLwimSY8g1g0gEoMr28
77Quqyn43z3Z/tPTwJEiiS93Q4ao6iE0fjcBwYsBnc1Bo68HxG6VX26bin0NGSvh2aIMPm4QBGcE
RGwqOnBGtu4nhOW32vVCWhYUe/c8j/llLcXbMmahHRfKNcCkp9YuwbuOEweaT2TTkr1QxoAL6yhC
PHCnPVoyHtM81lCXIDx3svr9rooz7FPcSq10cFv1uDwBmif7WAYprjzspiB4F60OLGDenQQl8niu
isRp4vmBtLbhMMD2vJPg04Ur5mB37Zfin5bv8vcjKcaKWfklpub/PcizCoewLWmui388gsIgh074
Vy2IJ6FawNUhZ4aRX5kby2OWURV/eSjot2KLSucKnu+EyhBjnN0pmebRZNmSsahHxce4/LTluGZK
ZLQTcDdl+D0WhYpL1PcxcWL2VkHe2mioGr6QBa9B6PV3K5JVYRARGX6/zE1/RAeGrohr/ArPoosv
EDU0DvSbNC4fsSAWnbZPk2WM8tP9ZfhhVu6XILjl9s7aPOU4FI13pK8EY1HhVx8AC5z5ovgce9br
mrvEfnLzpEg8ilf8QHQhl0u6J+ZWEX7uTHDS5qRV9I+TuFJBsP39v3Vx+hx+oDypUvDebhCNgBCV
wLZd+yhdwIRynWzCZ5xx6GlqtKS+2lob+6U9PXaIWM+INe1L+qM81CiEuWQOWWf+qYqRAvXxC1YR
FIbYCC+NWbkz9+e+hUJ5S+pL0tt2G7EV1XdsuC3Q8V63MgDCPMA4fnHXagrYLmpeM7HHO7Ldbo28
BiH5scdhHJtn12ySD8LBpOrfEsydX7YRwxEqFW09bid5/lVd

`pragma protect end_protected
////////////////////////////////////////////////////////////////////////////////////////////////////////////


`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-1", key_method="rsa"
`pragma protect key_block
AT73zx2OVs3NmmZnzAKyecvV1h0J76lrbNfkA1UWrpCdQ5ZofgTAKanclRablHNcVYnKzPBua7lX
leajL2rXBfnD84OkGiwLeTA3jCLiAEiHh1OLM0tCIUGkGHAtpaCcuM1qF3NKPUjivZjbpSMLrsWm
W1DTVh0KppRT6OAqZoE=

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Synopsys", key_keyname="SNPS-VCS-RSA-1", key_method="rsa"
`pragma protect key_block
otAx89ru1ytbxx2RS6w0k/OQF/wDfWkZC5Mk6USsCnWwJ/xbV0xGZ52qKlSHw18TO28ow+eeNd9b
jhNoSHalknJtvN8Mb5viMfNDXxdvtRT9QQNfFC2xT6aOd656Ks/qoxChFRBUnYcbRtIDkosqZvcH
bIqfuyWrymWOXodnW8o=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=3232)
`pragma protect data_block
m+/PL+VnogwTyX6X+BYCH6eK0gpScGia8cj09TUjM+hpfM8w9W7Dt1n+jfsuxxqfrOL5r0fZ3yMA
u/v4/ek55spYdaNJNhembq51ywjYeyPNFb0ntbVSPvFXnpBH2yfj52lyfVwm4vD7vLiY6YAvlKQc
QQe0Ap+k1zXUolEIYjzcQdBAMeuezGxIkGyO9iYRuZbyrW5KHLxwjwN58frokxJu0lToAOSUoC0O
TCtSTBv9c7KeEIOMWNEpf593BR546Jm+U/980DkFQ1K+SDyLr0XWav0B7lf45esBkowPYW/oUKn6
xvn656OzhuhhpzvyVC/WAgVyozhqme1LWfPjo/SA8rqT96WKeuKe3Ekt0Jm1slAlT3EQyw+F2Gqy
tShcYND+yWjE2E7jo24tg2HxTQnC9bPfXIMa5VVYty//Wk4N6O//BW/yT3AwbTICPHkVBo2hQSdX
l4B2tWeNHYh9gD7pEMEnz1fFqnjqG3GE1ZaNwvNpEmIouJI61trRrjTVeZ5xR10R8XdTirgm4kXa
/dETBc7giARWy79PE0GTgfEHCo8s4iN9CTwTYUf0/fSklls4E6VxnpGUmpQiQsmTBpHbQklXjOMI
J+4/RbZai8eCRZvlLpvd6IxDdTuBAwINiSTMcWCA2x+4ictRZAfpzjf/TaDUhjxMCHUYu9BsITwu
KWni89Dezz24B7QQpTAS263VSn+a2ATpW79l5gDZd9ItHSiqNj1B9YDv9pZm0jId+qvuMS4sYu5I
7Nt2ZXO6w0mSD3aIzYQ/dkdlONdrUgzoOnt/zJhNj8b0I5KoIV6cc7Oaj8GfUxAk5oq/kLOXC5Tz
diDOsRBCzAnH+L5SDNtFgNLvJGZligvasUYWYJTF+pxr/ULoXHZc0dGiB/vPkngW+IwmMJZymZxo
P9rz9gHMEQyrngtFLKEno6uPvW8NL8WaeTIF/hqK5MwT2prAZzQG2RK0EYQtWLS07KvaQnRsT6Nr
eM8QZ25UQjVEexB6uFB5cXQz0bMdJ+Mdy5b7a7vLTDnTQjC87dHpdwRA2yRMuY0+i7CwGQUvCNHk
VqwueGjG1BVdM3cvZH5ow9dHbHHY4AmIAo15MHkDrbbvPBlOSkVmImN1K7URRC3vCRlpg6oR1Ywi
6c2TArJhYbNLPFBiprRAnqqUhbpN9mIL+5h1/oV5zjG0GWm4BkSyZeQ5gCD1gEdR/yKl3kE9ENGc
8D04mj0NyphOKOE8hJTwgm5nLDAa3ue8sVgD8jerBeWKebP3dvc1LX7jMszxzXy0Ai85w6EuCeKZ
fmxR+rSIZll/nKl9Bh0MHVnS7ZOTPcloygifTwr/7Gp23pPLfnFRvo+VFvd0F7n7urmskAMajoNm
oraamF3Ru1yhpN/Azl6YX8jQ8PugsuDHrIQcGYJtunAc3k6Lz3cZRhbRtWfB9YJUNyjEPoj+P+Bw
HNqL0BZSXLgdn8NHejx0sdsM3622nmYJPKL2wLQ01s+/M9QZ03QZFXVTFPpcuiSDbEvPsZ+mBsyS
1MA+VjU/zlPfp1HL+9la/yfKGCYD37K9En+kcsaS57XJ1+8wqriULIoOhbIoNR7+Hhl2QkddKmKh
A6im+VPqYIMtg4OFclZp3ztMMN1bidajbn3qeKKWApk++DNVhUqs1RI0hmjjUV58we01pYCArg66
CQ0wX2BvmSoVHIwDr1siz9DTzfLBxbxZJw/nqNwO15s1fYE4k68ndHekDPi203iOyBFx3pGVOtWn
pwLbDT7OW4D8jWedMhyKjgKGFQgKqyJUYuj2Vs1G7/cjtS4i9kE6NL4FjXYRmVvDN381ggyrL2BF
Kv27a8LyFIuFFqPQchmIjcM39dZKs1cfaeh+9E0SV1xqbpGrhOiNpfGewZroeRinBRG4EZp9ibpy
VMkgaT8+oNNmewMTgghJ+UtrtjbcIKa6gt0+ydWvIR9RRqbHg8qxpRKOGvp5e/dp1kIjyGfmiAip
wHHt5qScw2pSqB8MwgA01SMC4xMmRVQNfolPUR0bN8wiZsQo/Hx4lAoCBz1TcAi/oC824yRm3Hes
9EChcXTLakXWcMsN2jmBMXC3CxlEqVfnqzVMxWiEWxtWPNrjorqR+CKhw9Cs9MRW1QWjXx/T3+1d
x2klYU6n/HbujkMhbiYvAI7Znf+D1EjneWcl3yojz5gYflvaFLZvyJMPNGMkRrBIOIg6v1G2i0rE
QUkKtfExbQLIAtz9q975sX4yy1RNK7f04oz8PayoRpQRKskIUNuTAhvJCMOGYqnb5ju4RVlZY2fz
TjHLVBCi7MlOl1ECV+M0jpE1t2sGptOYVw2Q5KUaaixBSy71odhhtWYrjJg0GQuhXWcKZoOi4/Ij
a8Pq4Mwh+A+CJ0U4WkEKSvn6kswfdsrTktvpO0pD/7Ug5MlxjhXtkOIfRrQNZyDNP3U2bmcIRl4E
y3LCNiiloxKMQjXpfTdFbum+lVNXCQ3aJw7QgwRL13jeRTSfI9prjbqEEoWQHduHPryi/pqzQgwp
NszXond5N5BA86h9CwBUiwc+57M25umxSw/4YfsYsgyg/m9Mdzmi8fhh5g0YV7Ekxtj1eu5tjZZ4
fFr1eKac7kDUqq001gNRyQAAVKoCrZ94v7fXCC8K3erEEI5zEz1c91i19iYYs5DRU4llQZ7RecPc
1ltjfC6aYVa/PQuzpdt1ZXFW+i897mlCsZwAueA2FmusBHvzKhPY1uBB5b7BlN5U3c/1/6qclvHn
nK3bPoojn8/aYmoE73zGdt8ZJPhpSrSw2wzvjWUYw0eWM20XZXQO15ybBQNbsTX70l77/1ZAIfXz
eDNHWngA/56mT7cEnGQPwo5Sv1seUYKZhFJHutZ8/cil9S8zjTDKeWtHXxWWnyDo8grJHTKJ3JPG
VhNVXVM/wymkfnreE02ETqB4RYrpkjhSfDLnqO5th6VnSaYkjLAdlIFDB6SrVOMYY4fTSFoO6ukq
IGft79XmkaiglOQ5j3W1dZsk0olx6JxDukE3qeIZugfL8hCpLHMGFy0ouoPr6UuqCVXhVQo6LrcR
mMRMZEWuboHkxIkmlhkesHutPeNUUXD2g/UWLyb3K7owjOcXkW+uJG0NsY/kgQ/aHAqwI0mEwqrR
t+VmjFWsMrMvV5r0QRmLI4eMbBVmOrhy3CuYio8kRhLkDjBZi4ZYlTaplTEETwlzysWpMQ7cB1kw
aN7CWr8RMPKTGoZhUazUmWvpWMf7mbvUTZCdRXvBPMYQI38IVEcb6cj4riVbwVrVZnrYW7PCPjmI
+fu17k/H0SY1XECYPF+Y3O2PjNgUUqmqi1SLQUW7KOkyasB4WDKpjT/K4wo6GnsksDCSXox3Q5O0
4m1sdEZvKBEJge9T+RZ73qG+T37DXkMw83dT0doaocPlyJEqe2f9bQkto+HhfGn0yP8HJ/LMrtJM
miNhRsFYO1rACK1Nw5ENPef+RBwXhWsXLXeE+w3pP54XEOva429EPReirVhFGFakceGf2yxk5rSM
CnbLM+tHeU3cnqOBqnZ5mekhRll94PcbicrRT++ZcuF1uectQYpHiNNSzqA1hwtZo4/r5vFKXv0X
PdddlgQ25s2W7dtNuksaEoM6FTVTys3/VeHchtMOspAYBwcWIDmnZfGlKyd3wWGDBphxNLDR2ppG
IcND2qb+hsFhXM9GdrYIoraru1r+Z8MIZ/e/wouqLIBTiqPe8UaqJUmzFzFBR6gRkYHULQJCAvTT
9yC118BBPONk1KE3VwFRLlq6d2GdlopvzHLQUeVffUaS3av/WxbNdaWWgYpCjYDR3mhv9YipBx7G
PPSq53FNK7EktCkc3Py4ZKCWjiO5MjMA5nMiM1v8c085t4ECP6Efc7NJhFQNEljnvfz1bHxt1U+q
rcjqbTrYYycaL+wXjqu9AifhTBYirQCRlRVciuXifpNUPJGozIaK+QiEmnlPvWRZncEMd+oOhltn
2+hOFVgdu0Cz0DFZj9XELjlBn6Ges5dR76k1aX2Q01ounDZILFbFYDlYwEReP4X1C2Q0Yoh+hHw1
ZP9fOcUVouDkLuF9HfaSbvc88r0XNIymJWapFqG6FtD8+E2vuQxhyjCJ1tta127WotINm6RTIUGd
ewG+XZ4RMmUti1Hu7VUNo4XNzFPwGUe55HPPpDSW/sddmabGQyK4SxXLCpFGsQlxB7nvd+3MARbE
CEvTcRFMomahej5TOBSSBFZNnPsFyn8gm4nAsAXH/1yDdYO6gUeJShz2IVBZ92ELHV6Xi704sLio
mCt+V6NjT/QeTydIdxVxGQoZlTbrzkX6ovT4udR4QItS96azQZdZiQ==

`pragma protect end_protected
////////////////////////////////////////////////////////////////////////////////////////////////////////////


`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-1", key_method="rsa"
`pragma protect key_block
OD4cYVm2EjkkAZb4djt9JS5anhwI2dsaO7OT9f2uRxQUTIhnQ2R9DHIci8ldX3yuNylJmjjJLPvx
VL0KVWigerEwRejJKOYO/M/rOcJXRUxBetPNT6ipPnZ2iJTMzQ1ddOxI3hrtzVN1B2SKVd81l+Pv
y/QYvoVoob8WtquRUZs=

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Synopsys", key_keyname="SNPS-VCS-RSA-1", key_method="rsa"
`pragma protect key_block
r6I0kOXtWnO8EPvprvPdEsjWLFI/PfB05M4eG2Jx+T2x7TVBVJ3CZLjhh5Gm9oJa6w6dGuitgB6z
G7XqKgDMgHJ9ohde05ZCPkUGRJXDAfp0VQX5ZnE4PisNa0R2ikdIHUVj+fqyQzmOLeZaUVvXxaI2
eBAhEPRuDDRwUUyADeM=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=3712)
`pragma protect data_block
PXHPJrC6dkHUQQyR9bs0A9SQ2NJVQ8GrIt335pR8k/BJB5opisVB8yK71x48u+flMbzKff6uIVA+
qKGBZpnODxHa3h2LFLDN2G3tuI09pBr4q/+Q3nHUkC1n4648nngK2k6pjDE1uIldAHGhpuZnkgi6
nkL6OuNDzr0KriXyi1RvNq3kkbM0ROfkrEqA2n7ZnB76A0su/OoBi8UVHNJES4nYF5dco0dF/JJH
311zxUcxRzTtimk3Cr8cMtRVvJj7TN5Xil5vQCws7rRQxPOtU+jkasn+gS0kTLlSJoBbbWiP7rFM
YDT2BQF4SZbtQsbeWwUv6H52mJfSjRIFXdxJjAnTHIOBb82h1esq2eIVqIZZVHLAF0ymsTeqhSdf
/ben5jLiZof+KolMI5W2hHkcPIHfvnc0Qop7vLLijK+jZ7zE70WHNQ7y/CkgAYnYhdqzwdJOHkPm
BBPf4Sx4EBVkfots/ixD7okI7LktFfuF/v/GA8MfuGPZ9wA3SBQvrEDYFJyQ70k7Qg3I1QAnzjq8
2F7IVp84fkKneBcVnu14R60oLrm/NIzOAmu1zAtxuCPp43m3ffarmAgolx5lWO8wLoxQpMjkpPFc
ga2sAhnm+U0/ZlMfpORorOsw5Ict5naFB4IclmDbeGwZUIYumj0BKpzNJOoI0S2kY3FYiScKivue
RLndKwa1jTUWfXZMsGcg7DCuNgcjYeBOXoL6EUBRntoGk6XAqpNGzQOrCoL4BvbZCaH/ItsSg4RD
svrvtsp4k6ALR2YRMWnCTj/aRIjydKanCtcBlde89FVfFlTgmJyhg+omcHh8qVIeZTSTDeXp7vPA
A9P/YLSRMZvS6f59MEX2kvEVeJF2l4SmsyPaP+gMiNxy8kZiZx/VJSTpWPAnCUY4c4jp/PgzhM85
KoJf0W54bKVzGeROHx0t1+mQBs9WF1JuwC85zh7YMMtJIWhfieg9ssA+Wbk/pU9DIRfgs7lIG3p8
Q49RwUCObT8QnSX8wzejUW8McWtldSeY5fCULSEDKnaFqDPD4t+ZJXv553KIeIwbGnop9DJDMv6C
S7/CxEZqzkWIY4+KwpN853fGnEaESQvA51UqvLAahGxr7zxWe0giJD1U9hWKyWNxTSEZRiQYhg5M
g7067BxCfGAxsUqeTEoh3H3Lt+Eiq1GtEceTlq7paWfS+NJskZwZzqyuBfClea3XKuM3I664Fr6J
O8bOTGeleUGj9nzmxVANBNo0o55Z7pUsU9jyz/hnyv7n6Sgvk0pXbos3Vw057zGKm1tG4/LUkObr
ti5ONwAnwj8chyd5S2Aw9zlQYZAwIPp+Vjoa+HGhlka54JT3q3cx9jKqlZ2h0F0KIPYvod1ncNNw
6QhHHzrH3KHXxmxtF+Mx3qWMY8jPUF1lS2hKKyFLzk3SLuHmCSNqkCkMcdyvef8BtusjYpVSkWRy
GD43UrfXP7/adYd5gaBP15v7QogNmHXSXO3oGV6//269xSb0vrfD6vvQdfnZ7QzKsp/rryfjY6ye
ctYhF9BaGSR4RnM6THs/iEA93GHaHKIk1ao1k0XJm+1VUyFxqjoRH2N68JJK8sabYpx+TPt+TUf7
cdy/O0C59yOCjl+I+h6MmY7BcYJYlYkpBOWeo6UDsXlSRV4qx/uo2YFYB6uYCsgal3+Zng4tb4+m
oanPogprFxFRWroGSOObVR4auJDGUAn+SdT+uglgECR/OOXX5BMJkvZWoFonIimeq09Z7VrrZyoI
rskuryCgP3K8FVi5AlzEpyC5zkR1swUugTz2jhQnha2kI50Nt9X5jeY3dtOoSXOsMwsmUiv6gzb7
ZWvrkUvXr/eZyyRRnFUORZdmDkzw2ZljKeiis9NH/nWBZTwRkhm9CUPhj6rrE/+asAd2gXERcgJ0
F+klxkC7s6y8bAmjB8TBctTZbR1+FyDBca8mBLkm/L8FOPiD4CUJjsyl4in+a+dgQufSF2g4MtfO
5SwLHFdX4C2galp78RF/22Acnbxw49QBoCSX21h1LZ4BMATvH8+6/SiHBnBxMorxuJ3SmthMf9Ls
CL/hYOjmLjk+IF4WHUP+9OApcceYZw8RNfM5AX4x6/s89uHqpzY70i0ZSyBBC/8P+Fnu+MtTatmA
QK6QSvVWwgcQABgQx3tIzjNcqJ9ejgN/PVekuTAiABYVweS8T8vNDqzwy4ukGP+Gg9OnVUcr9OKY
niKO1PAYKzRrOaW1WFd2/PRT2drEPVI+QFWtEttKYQGvivEKuOc7CjGua8Jti1LKx99TsLd7HRYx
G2Ohg5/ABfTt6SpA3dS/YUdcDebWBdeMpWnWyOHlQtoQbT2U0aLDEsZuQdDXCCDwbdeKa0SUWy+C
1hQmAjD29tP6VIV6EEV/bvVI0Q2udhx2eW9uph49jCtr8RjcRChmj4cwfsnCMuqkfS91C7GzhMeg
ZJ8OKSkIkJixtck2+8mEopptN+PmHuu09aWBOkVonVG9nhrvEveFnCG4zXzuYzNjW2+R14aQK2JJ
MzFqV4u7XfP3gybUFjM/4DZhRX1qTG1sa5pnn1HflPHOqiKNY+vliGkEcMCALPV21GTvOfamWyZA
4KxVqFM6vLGc1A+yzESyk1e4RLE5AEXRa9036UmF4FdMKGAWe3LngJvm0FuxSQApw/OqzheTCoi+
c29YY7lApxscHkXAoJV65TdRLRB5RVeXwJylcvG4cHazZRvqWBi+xiSH9C49FA/Psd5GgxUVtdMo
jnEN9tHSj900Vt9WKbe9rT/O4qCCnnS4ijAWEnOF7h50DQFavzzPiaM87ocCSq7Z31G5vIpPVxLq
Ur/yJCjud/y1RqSl1JPiTmbn1uKNAaVyqdD6EGAXVGBBY/EoAodhDu/nFK5G8W8biXEdLB0tXuWP
fQOGMvR5/CMDkLjITFtgS2iEiEn6Oxyn7kqeX/3B8i9tbNUNI9Q27p2xu3mgdBTn9M1NqSJzFfXr
HbB+FQfXkRcND/Mjqb1NzbfsM5ocdGbLKGjinGT3uXk/mKjG7HTamyVJGCVP3q2A8kHQpTyfp0Ft
7j8s+tM3tWRxVtW7WaFi/wCt7yJIJaTmUFt7ZrZYxVRsVKs829DvItdsr0ywrdQxpZYMW0n9nWZX
2cBMBk9/Y8PwPt0Y2XKPM9kpXJ4mYUik/WDKFko+zqQgQaRHhwJ6qzNcQZ3hKU0udRypy0b3vDF8
iOwX77hFHMZGdvvK/1c0IF8oQxAobkDjAke97pqhCIZvApmgsKHw3LsZNmbLUcZvSzpk0Hx4bjJu
GVOHmhWG3fm5jS6cSngSuqHG0fmZxmgpqIOEruDYOo21oYbNOfoIu/B2lMNgIGLJ9jqv1CTobEBY
MYsjEhWzODfefmgvQZi/rEv5+cPOt40ELMscDhR60kM6j/bxO5fYyLpSe6fbgyb/9XXRmjX6Crin
LcM/Aw1JnVcThy6jTYI/uoSFy2vLwpS73Vo34Bjdfl8b8Fv9cyHd68szTL9nkyWAsTRsXSzxGXTb
IH7xR8McIkBkkry9YP5FuT3FtMI2EwBGZDnzYN/pLgBtbgNxWVyNDfjXTKJBZpvEZ1VUZaBStW0B
c32irJ9qL2ifsr5ukULmZJUcLqQ3Qc60uzerASvcBqDhEh/LfQ94dNEfNweyCjqFwy/B16O6kjrz
EfddSoCq68DECC8opoKD7tcOv/yr/RHfuei4EdN/MewHQe1mZoa2ef0u7WlI1GY9lRLzBOvxWWLt
9Mo2jDu1gAy/NMGDobqQDVeHylYQabkW+DzQ14LhcmOHSYe3rhlLhhSxobJLSu8oZhtSV2WHu9v9
Jl09KUTKslBPnRdrftMEvWCuti0gjwp53CtFCT8NhGkgT3QPJnr+U4LaOpUpvpevYopQkZpDnTkv
wn8uPx0GySegp00soMoUVEvvGqaaX/DQ+YEtzggdVLDaGvOYZRmJLlFrm/qUJwt1nFKVN+nJ2JjQ
EP6ZODVc8JCmRhxgdOFs8/SdPNnUUABWGsxoeHSFs0VOoEAvlMnG6Dc0vSpWihtcj7F5a8yzMzDb
zCNnFstIafpM9NdnlWVENGl9pTSLCRNsZDczQVYEbWensk5ceFtRHq3yQvvK5PyDZ9ivTj+oRxEN
WzVTbytDd/i+hK2AUdxU70q+5geiq6XFsX4C1pXKGh03Etl63Pn3j6MxPCx82BVqbzHUVPNNMA6N
z8zahJaaD9RPAq5pbo5arYUMUzfLXQbbYGrzeqO6NqmwQo5QKwHSQH3EeLiFa4p1kRwFL0drCJ1q
5izVilDlEwjj/86nUni5E1u+yCF0bdKax/3m/IVV15vv2isy/I15RvkIBBqFw+ebojkHsrNrjk1E
EIHuZiOkevQWoNcWMhN1Zp56t6WqikTCD376dZ09XKzhjvKLO7QfFJQ5YNHS9S6yLIZY+RJ8odlU
IZchR986aP+Pf40OIxuTW1ZFMuCxDv5TUiUmedhvhaNHCfi0CsfC4ezZZZCi1lZFCD/pl87Gkam+
DdxxSaKybLhqwLl3/sC5Nob//5K4BI/e0+YBtsy4pWgpvG1YWlztxXuruUNye6h5PGwWKHVuI1D8
9ux3GBoc67rGjc5kJt53QIZ8XtTu3CQOp3XiL4tlLmbnIvZm5/AKgB6THMDsPlK3Vah6ltQyEqV7
5ncTPHjavL1e3wqdmIqVcn0yWue6kScuu82MFsVMOJbuNhH5uJKw4x1cXmo9AfrPF+wK2UUSYs2C
KCMHzp0uEfLmEqmb007241GsMyi97khf+YxjNY934KKe8KYn5r87LAnMu046G0a3gmh/fhUFHLdM
PO+9ZrgtJ+MY3g5WRlR7dzei4tYjZ8jUaDra4h70jCb063FCXKUJ69nsVwuUwni6JtN4iIPKX9Eo
BWfFSQtFkNGJ4DkYjlmyndDFZf/VKM2IXq4YhxKe1TgvkZDSeygMEpMnA2GzugcuIOTIE4D0sFaw
Ar7J2FrtbA==

`pragma protect end_protected
////////////////////////////////////////////////////////////////////////////////////////////////////////////


`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-1", key_method="rsa"
`pragma protect key_block
RNPBUXgikxhy5tFZnJCoCWH8zGPbcFauWixrpQqM1eyVTbBVSvhoos/wleaUXB8dTFZjxW8CfI+Q
wE4G+eFRqYA9h+jmNh4CEXPkWwVLCapeW+E3ADmBGJEfr/KuJKkAvrkqIEffA5sRUHsGs9YvTdxD
BH73UiqXYa922NR58XY=

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Synopsys", key_keyname="SNPS-VCS-RSA-1", key_method="rsa"
`pragma protect key_block
2CbdWSNt+q8neZErCPnuR6EHBQL0X4VwdzZpQYx3PAVaTBDFxVuWsp/0FiGl0aeA7ivc270NfM6H
CSsnTi8+vj2XC79e9J1CB0r/E5BZegtqA7jq6LUDoXZ8H9RXeR9YPmKrB2y2HgYSmBTj4OHwh/JY
+HmaiC6YPTkmS+rx7Ak=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=7744)
`pragma protect data_block
F3qFfcD1wtXAon/QgkOw2r8ah8UQhix3uVhDjNDjZJfR2rv/9zee5FyED8fZTyklOF05GKFUvWGP
52r1eHQExN8avusyqJOIotLXBp9FtFoQcE3OFyrViGAUZx2EX/AQUBMvKj0fogFcjNsSTtT/jTdn
Ju7IKaS1OXo2xLtvlk9zynclVtPD4oegI/bBINvaTKQbBZBnr/8YUS3amXe2EMsMsLgmP9BeUu2X
pFxcgWeRSK4IY9HsLFuyljrxztCIYHz7Pb/FEJ1hl8PoNF/Pi6T6cDqYzfVgd4wc6jrVZYr6tMQU
rZs221K4PDh6YPAvdpSlDjzrVdUyZ5u0n7ZdmY/h3uxcuNq0OcAcPgTI+85gUJR3mRTSP37UeR0A
sMniUC3neriBMW5Pz4wu67wpJ+MQqMFq0HCwZEJfKqBsO5oC+lvgaDmMXaKkh0BDRF9/AEZWY1Ld
j9t93OuVq9fcLjhD7W8wpyi3qG8GZ/LzQux3185vy1xS+DjuQyHYkXlaHNpP7eZRor3eymxNMsdw
v8EbOs9Apt6TkbGa/llJSSE1k7DZqgZGQqt9gS0NY7a/EeGIlFL7Gb6dxwCZeg4/OMjo+gjQqmrU
97gyC+gsGlnf5Q71QBCyGL3zlFj20dQyrkMOXi0uJptgVozN6xogwW0ARP+ySZNqTbtHCweTcLK9
xnsavoQqcB0Y5H8XuTEUETUU169ALVTDM/PfwR5+k0+qfqY9rnXbzNGe/iCEMHWLXJDyozDKEX9j
nApbT6BVi3xfCkeKzUuPurGEI2PK9WWL7I/3L4QeLZ0jCrHEKpIA+9Wvj8oJ7n2KdnuiYELho8Py
4IinIcG6qBtUV6gVzIGT2udmbhWCaYYyz+SUT9VxH77AtpTRxd82bOww30MNP3z2DrALMPQMgaop
G2pRUfA7v9L2oA//NxLUvENUeFol0trUb2ak/NwfjE8alJ7xRQLsV83v9neRwf/mj+JqX7OW/GRn
ZJ7oMkVqNxfSk/Y6KdrhjqlYZBmtYpcrqSPdRqckar29sIDcL6dDyz9VDE7ZidhbxE3rseG2YXOz
8rjKhYUwM3+yEY6et2NmaQSCgX3/yxjxlupBp/JJlXmMSZcm/bseMzv8tvhZ1lXjslb47GjRbG8A
r+KTdpPkBEh4zw7uDMz9DNqR1y+DJorXgGP/sieHp2OvoTypDi8gH8pZqxzVI4avHfTEdshUynrO
80e8EB/mf9o0OMPIuEg8vdkJJhz2ooSBPM0B2ollYjARZMDsjJJTIm3AAsu4msmKn2UPT6nezkKg
LYpNmEXK5xY0wbkML8LUWxAeTby0S4CDCjl9woEwwr30Bo83m6K8ZhQO3RArDipbg0gaAjxwlfFd
mbt6GzKHpeYuZ4xjKXR3JjwpxQeRa38goJIXCqc3JqnPDQ1uOgrjZk8gw6Vyf0JFg516ts2HRrid
S3khFub0EO4INSIGFfUC/GNKd+8Fsd7nF0ie0ntxxO3pKNL3IU5+1xDXJ8gnc86NX2hnMo/PAaky
Q85OPUZ1n8FvX2hMJNS12ECfYKSzPXoYu9lDjnCRGwL3PGGy8StpI8a28moV4bArSYVAy5lkUiJs
jxencVQWKUnOVGhkCFGk/Dy8K/V3d7Ey0ZSUWiBYBnyjqtM4WuPEEOJG6R0P2/IygTTPH+98nQ6M
nxwKgdAhntBQ6rTw2KDGUAbfpf+tjmq79ejSJ3mEAxWSOux43h+m5LJRt+3CxKVuzRJcP545EUHG
JUWqyXleYl7g9kutaj5pBDoWE+UB081u1x2mgBAOR3m7RiDqMLON5AzWukmfzvkXQTG+L+vxO7VZ
FA6Kp0k3+0E1b+mpSF6QRazzgL4JVi9+yd0Y8HJx7Xb6M2mzCl219n5d9YZ/OFnM7uHAiY8VUBuu
LBAD6Ky5XKaYFTNl2NyiP7ktRQIlXI1RivORRgDoDY4pxDB3YhAECYTo5ViX5unBxmBS7yMnshWY
ceX/8VXgInqKi4/EpKVbMdBpIp5j/eToRz5yrMX9GU7LNdQ7GOD1xACxWYlJXez7JaPJXZvqKQUI
x43EsA+m7TXqHXmGDc/KpmTSmAN0dL/20+K/VCBUGACT+c+zQpj6+xj0qnZdFBMOd+DhHS3CxWPY
P8PNTb0nsAv/bFeERJvH5sUewgCotADZ47uEWrU9uxHkGTzXJTXHUkli6NxcNngk9bvP2CBa3EA0
k/PCM5Q5/4JDP6vLKY5jnpv1IDy0Lkg2VhkzWiMTXKOhNJm+0BfPJr1Cw7ic0YwgBxkUh+eMGqMd
p6PF8QoImGnLmCgaFJtE93w2YKS584z1mWzdvOfCkLrBK70zNf+h3R4bNhW8LdF1mGv8iECcum9T
m6tWGRfB+QILvIr0sMFugIJ+gG2bxlb12a6v3TBnvb7NMGPgwZ/YcqjdKaMjDx80cdoHWY8RF2Nt
qUuwO0hPfuRN0qjZ0wL+coH01xU7vyAP3j41Zo4eugA3X2G5TvmNx1G1ybr1gq55Bjkcatc4eNzF
HOTpSrnuZOnttbXuGB2ZeMXtWCxhFL5SPMMAU1Ares1crgMAxafyEPyEMvCOaGKj6oiS5iiztakj
uL/+Z6OqhMy6Lq1LAodCXo56WUbBuqjp1oKDiCFdIGoAPkMejZJmRqVh3lzmyUrLwPyoksMngdIb
QKsnfzSk0SOw+TgXQ2tWaNEDhaeP7h9w8m59U7YtoUZYp6ilNQoPVsySy6fIJhLgcmPgMrTu1ooT
ST6XeW3qYsRp1IGpoQtC0OMlfAovNIooI3rbQePLd7j2jBNxuuLMFt52HlhPvPe5KScuVXMq83HZ
rg6Djt8wDMwu2SNNCXxVmTtwGtRtETBSl6svaDlBhTrLKIXHRriuv8WllQUmB9k4Ec1445klls+a
t4t50gTr30g6Ix9IhiQeUXvRIwV0xTuNN737+CvjMaUWYlikid7WMcwg8atzB65oALawLg2JOIbL
zs/yJtrbxOzpkTmx29WKdkfUxxMUmfUsz7XgMr/s0XfvgilP+sXjSelH8XJtpmqBeumhlUZ7Rbva
xJcXbajx/L7hj6LicHlnygtEgD87Kdb5dNSA/0VjCjqodLDAqxm4TPaS2QlNH/bzp0NK9IdGmoya
eeIREddmr+VChICaibchGtkqTkJp1gRV/0oIh9Uk2zbU45gSSHdO2MK2qmVkQLLLPtZW0Hw9ukyF
Ief9prElx4X7yZtmf4RtEG7o1wzCer77lwECfEw6gQOnXJVIcC5ou6CjFvEm0bxVhZjZWgdv0sLC
NEzAFCFw5Zo28frY+omXdC7vtKIvLdHQ3BAL9MvlxHryKdigCOtzOirVkMHqE/4lb1sggYURxO+2
BLXj9Mni48KhQ1tG1Nj8sT0m1cPzm5qh9aoZVbH8GU1r5vOZlJxA1WuJ5rzce+QipoYHBJXz+KNt
LVKma/9iH2pcQ6nZwGWJ3/K5xeiJ94PyBfbE94Nh9YJ4lYc1WGp/2YLS2Mj8rmuOIyQr/qTpipwd
8VmoUWU5lcAo3+pstrAQV8WppJE75D2tjT7LXJNRAljeQvvEvyj0dkkFr8fgPUv+luUX+BF8fOzt
wsDmygNqYrW+6HNBgegt9dfAiMJDgPqB4JePKGpaAT6runVpnQkKWnjXP/JGT4J5BLREQvmjOaVU
nHld/ebB/mjvFeW404VFxHEnmnuZfot32UviU9c/IZZ8E3P8o27YEkcr6VI+qR0byiDL5wnpHN2d
SJGMehyrplM3BZyVaxz/NK5iZk4LWl9vjo+O2Au86lvzYs5cSruv45zpxCFYDUsbHdNne1gbqjAX
pzy5670cDDMhK9qzts1SZUblFuGzu7awK5XDTqQDT5yQqvuNmDz8VHWJtlGNC/mgBdgIdebKF1GY
0CWEO3lPMBKnHm86NmsexT9NgB0plENOSqfgAWyQpzMhMKv8FaXkJLIJR0hjOh2osTxQlCJqphpf
Oeoz5eRZ6FsZhM0f4XMCUkP+7iTZchJ2bY5qZscjhzHqpFNoItxVzuuv3287imrkLOlmGlAGy9tH
3dz8wlLqibgAx+k8n+eBWcJg0aOq17ioGmUVMqfkVmOVJcbXJfQgUt2vto6DOHLJt7r/aujXKRJu
rkAf4c9Q0Hsht6U/tzfTRwiFss9T5jJksBRJ8rNBCNWNAndv5Z8rkafxd6iiQEnG9G/YjIfrmjdC
HV+/mszRw+IF/teObsDm7kiQvkftd7pdxiPM7OAf4RiMcoYG9puWma5o8tWCzr3yMTr4Tgbb5Vjq
sp5HFcIf7DOesM8FAoP6adnXRrs0N886ETyzavhdI6b1QrBJ9ExRikD5lNGUDhaP/OCI5doykf4+
e5NGo01/Rl0VuWUdKETSgebyPdVWiFJwK713O3TRSJ5iw3JY3Hx7xbr+hQh4GABRiuQ+Rou/6q4o
YizlZ1SrIvJX6Pl0iPnZEo6Mv0BRX4GUynecR0cus1CFHmR4uvtZk5hJ7Eho8I+ed/Rixc0w149a
zyHIYHRgYRW3HMKWXXHckWGnsZFC74KksNR6K3+XK5FdwwIhAQYzkhFA2Iu4GUAjeB2eXAERe3t7
rv8GeC8ncxTxiXscwV5bAWeGQKUGs0zihD5y6sXe92Q6bOjOrBi7AfaLxZd5XvHbXvwr5N6n3s4b
L2Va4DfSfctaE1MGlA+Y/x4OXu6IxPMlR/ShtdOe91nK1aaXFnezS+XASxHfSoc7SLhLGq1Zcdbr
M6j+MDQXCNjBilzfbcNKJtepbLJEtihSkqEG+CCJ65tZJ7v0taFrZuf+sy7PKuH7fV0TLObh/dDy
mRdBAyMmkd/2lpIawDyrEU1x0AAR7tvdM3pYd+X5JvirOyPfgaXVfui9etDmBmQNkEe+tdfKlwX3
bGXoU1TcZ3sBpdHJ+5nCpHSyKW0BRaSWe3MOM/haBnbRtXHcgIl0D89UJLw/Zs2YceNSrgZ+Byvj
scw7uIt55IkubCfDn8mUqqT5Vh860Wf0E4Vo6JtUWfrVkT5el4f6NpnxfcLacQAASZsol94Jo+g0
2D0YqgCr98ZflQ5l6PtRxnhcflo6PGni7nnEWdUkMVLEQ5WmjZtwELnIkkgPftZWZvkjHvjdXs4z
VBA7iALhsniS9K9NPuPmwucnKzCLCcujWrJJOoLSALQNpNwfGzrMFvjuUq/yHcrPOXA+60X4l3D0
nu3SAJqaFGswcwqrdmfngmMCT6ZVkpq+DscGIzC+vkD/8309w0V/FiKdayevrrq2Lo8j8XyGesie
fodlzk6JrZSBuNGBAcxM9gCIw2oVz8JkRJKCRIn/zCAuhqMURYyvTnbd0uqb9zsG1njSUL7kZ85L
kxpy8dlE5cKYEzL2+K8BGAgcCBff5MshZS0hiRbsG2QRUvt6hhW1ygnzd+Gn7f0u3bJRrz5UvZ/2
GizRILFSjSgWebi1cQVA8rpt2fym80YArwDA60idHFS/+fFg5FSRm/FCGbeRZ9uqjcoZteE7dXcf
2JJZgSgfIqnAykpkALnVuSSar5WUVnmu87bpOPJrawdYrEM+Vt7TnC+LcaEU2zAEr11r0wWot4YD
7pdQ6PM6xeADc7MpBCK1hG/VSeOefMTeYJG7XYGFp6mJli19O25LXONSL6/hIda0ywoQSwwfmck6
wrDkyurDMRnlMIIRspWogpQvhgwoRJyaWbQO9TfyVqNZ5dsrODLQk3UeWrN3ag+uyp46Y0kBXAcl
yV0ax4mFfS59wTS1+u6yRSNv5G4wEtdVS4iz2WLot+rc7zr3+I/tX5cScmOvkT56OuGC76EuLFjd
ianiiSWHarXw+swIIM3vH3WABB6+UWepeGD0vsBnjKrbDqWcbQOyqcNktMs00e2z9nao1urP1SKd
F93oaaAhQkmgzGxslkBC+bihVX/eeonYcITzrjx4G7ZtTfSM5ZgWEMyOv43d9YNPgnvSTMwRqCJF
KVGf4Z4wUVYy0u3zLgX6otcjcDG+ywj0MtaWfyNhR9fppztDZ0EcWzyGwzxFf6/BtC8PcbETP4GU
Z1Q+Eq6hkRR7T5x6fg0GZG5MtWA3FIn1YbZpwd74fifj7p/CE/XhUO5EbUY2a5F4H9oTQFqD4kG9
cc4iSIPOaHL0Xt2I/hRaIh91BfKfSl8cOHa2NVddyyxRt3C3lEj5xVI/ocZzOHWiN7IoOieo5TDj
GLjrMRWdqlMU/Bs+zBnb43oDawgnA6w9zk0BPJr+1UQoKDASDUCAzOteKOGFKfXox2kf48rsnKM4
uii2bGJc4CwUMyUlHSt5xc/JdZ/GrpCEZtUSycRhiLAeNe22t9dOOBu+yotO9Qa6st4m1gEJb0NA
Efp1DDxuZehbOu+hLTiyOhrPjpwCuRcgFdxULrPomVGeOex99xQngRzU0XaGrJDo5MXCKf8XLkD3
mcg1vSmxUTgYzQ83GnwKsSEYDhaqsuqmQI9wBieKDaSNeYedwFQDuFejb1wma5cUru8tmWwfLz1H
W0akVp/ZlNaPNhAt5hVASN5C52/SJY9ZXjTqX2Xe7ljiMo+XCHeKfK4/ubxidJckvAlgRnZ8bUPx
mXz0Qh1WgLaSAFdq4HDh/CDZevdk7C3WhXxzjOXOWOXf08xtP1SRLAHzAyUTCoDNxFZwqPaUNKoD
HbTcTt5k831UHzwwukfDvWT0xpQTXgOQWNY+WiJZfCMV39BlCPO6Q/6Eb3MKlrIeXe8ljBKPGmu7
08w8aAeZLmu0YIW4Zp9imk5h79qCtHLDznbv9cnzmyk7iCyZKd2UhrTTKZErwtrLD9FqC0XSFCSp
GIQHMb86YXsUNzyrL9/V7LHi6BkaKWMp8tO332UnZF8tdtkjJdt4ks69mFyC/O2FB1OYSYbJHJhv
az+vxoACsGfRcEHaf3mEhIOeH3vkrSyDs8cMOrjtfPRUfwuPbaUBpR7m48lda/VHLIU2W1hlLZW2
62qcCdZaIrZGj0dVM/dvrHYB5fH46wzz7A2AeTj4d2lHrhbEUZuWH2MmvmBBvGt8y4p1RqdpdVkM
oxNftq44MEL0v4gmWRVvbN0KJs9b/Pj9a+mPwV70GkF3rWtO9yDE7+5cRrCPPUClQWvFEZGjHOF+
KOPPgl6lOwasH6GuEQBLfKPqwF6Eq08Yt0CqJ3BfHGCsDuktj8/sHJzu9jYDCWkM7At1DIknZcXH
vYX5uQdt33XqqWdFJixZsbjmQqqZXxfUAymjroEAz6UsdCfBfO7mRn7M9cyKfW8N38LV8i2W5lYV
dJvzYs03J3mAkZ+jTt1grEx/8GMz7GIhlg2EtJQ10S+2VcRvluxkPLF+5kMS33pYw5DlXQYtN7Oy
qt4wxcigr6z/ZADx54BzQE5WJV14GThy+1dxs6sQzA9jO4fCVeh7tL/aOgR4pg4JlRjV9WYxu/Cg
AbVMfEM6NkkFaAcVi8ksQQhalcLov57Ey7Cd+uTgLgUQ97PMrRNkAuLJKgaEcFtAG+Vg9dpnPBb8
VuuZ/O1JRB/90slR8Ph7Aus4spsej9PBbQwiY8VK5jVMyWjsZ36ZtvvTMREIvzzqdQ82PLFsoXqb
B0EWFic1if18szjuZTykIvmT9xMcfjclWOyrWNhsFKEqkOfKnsrRvyoEb8EwW3KfWrh9zXejdAD8
jXYP7WLbPuhCYLJCw2vDDBX0bB4IkKvYuC+tz/YAMsXGCc8bwZkS9mzEPr5e+q9S0Pl+GE/rVudf
EisaNoocAQ4FIPWNgA5oHxuQeXUqKwfzCffX39//5sPdcSQYs6Zxm/1SLH+sdXuWyvwqsIa1wXJ3
W5a6jrkaKvdOWPKN/tcHxbLj22B8ZwfNvhOQK7NqcARosyfRdbFnlBZFcDYtuXWcgYKD4OiWk6GD
wE6luzH2H3FPP0RkukRzpQsJ1Pb6a8LH5DfbfAgC5tKUdmz6JuUCcR3iMPt4oVuqJqSHrNwdLhhU
eAo2bu9cHjlQLrZBz9wgz2EVc5e55vrPHe4ss2J27mABCTfLu4Zn/TcGpur/TAneLMyOOxlocnzC
C8h9VWDDw17IiAHjsYZWayaeUlvU80ywTSa7Xu0bnUZ0qwfaAttwwilnVRTuMASF/+56cKh2pTyC
7dEZIgWdfPH89BOoB91lvrnGnnOysSZ5Cg0tX/y3/Olh7B8GoBssYc51IjBbFUE1pYYw6ozspXSx
LS0syJsVWyxlXawzrDRJ4YjZQmAJaM530RYwhWwmIRjT6LORYXhYQI4Hg2YbDBERIqSlvOUPRCeF
9ycdaapSElcgZQinRw12xRlJLpnjYZ9cauEzlkmdUzn3O1HKkkDKqhtF/NEEzKdkxX+P0Z0KyYyX
JodMvmQ85INqDpc9p050ZtWvXgAuG8SQpUuVANpfjSSC7/5sEKBHsLQA1Ea46QwotKenqEuKrnQB
rwTHtks/JsxpZP3rAyv8dRzNAc8tW0N9BpeuxFuiRln5Tv2IufjDTgBBu2AKXRwDiGV28WOhKH54
xik7wUCnmDoTTB/K/W9QHog9RvcDH8LBE5fmCxdMk1LCzAEzjCofQld4lNg4Ez6T0FaJxFHP/CdP
PZ6ciVO/iI9fh8Roy/A/+HWV3pK6oCrU54qQ3c2j2HHMVs3Od0iCZ5/JTOVND/AtLwvXIv+uV8YI
yeJHoqd26Y6NMeMBT04eUCaRYmbdNNGuIhUTmPL23auSWxnIKPYKuVYAPCptruzUTlq3whHYnDZJ
tCVIXpk4iu0yTiRF21DLRdv93e7u0SCdLjxmZwGTSX/H93JAhzC5lC0Pb0TBzILcSVb3QZjLFHvq
32QYkVxRADOSJsxc7ewy9+j/r1/y+6nPkHPyKyiLMO1/YXAfjz2E4vEA4vie00Ovfg42upcHxxK0
yv4hCiXtogMDzhsVCdSDDvxz38QVVBfImlKyW6XhNQazP1Nw460Qqqe9R1+EdZvLB/7xM9AZ36QX
oCEn4z0GjQFdjQEo3jgnI72eObeiSt+Sci4Zz++Ca6PsrNHFZkNvFiJzLqMdfw404WaQK3WDCLUI
bBoIJMYkNiHcw2sYxO02eubjJqt0kM+n6Zk9wI9gZGKprRlgQaVeQB9vwB+O/ZrYN7anoOR3M6cD
5spzVSe/luWBheump964IGJfv6Z9YBkFbbTFr5D5sE5VMOOWL4WhaJRX1GAHUn9cWHHHyX5gjt9r
kgl3yjztPFJQ5fpuTknL4+5+DxNCQzBTr1kEVdF79t6VO2dY0h3x8Iy0t7Qx5sG3IW9zpB8J4ZXj
RQIkg/Ae9QWpYTCCXTEbYm3NJeyqg6+FqVTO+PRRJsGfHixN0Dkdm5TBgQ0dVGYMAqNVdsKiyzZk
OOC1fhSFTd7o6AfAKAXGACg+GXYAJsgCzBv2I7u9djZ8DOpbm9fTEpHhqoE9LF5wsOPU1ZAJEHFW
M0x0eg/HMWGYt0rBMYe3hMR1IVqUbUt+f/f3L3zGwF5EIbXiFDYgMFXcSJGx6jkiRvAai8R9JiO8
tR8dgiqCxjxiVjTPdK6ldFXz+b6sqbbUtihVjqKLgpKpIJUWfgGk9ENNvypNnabSPA8b+3zoiWrm
IgJkqD0Pn/sQoKjtFiHlGrBNlnhYb7uoEp2PpXg94J/TeluA7ba8yrvGs3LCFQ8eBZ1Wq5zDNJk4
ZNEB//veyAd6HhNupJivyubAmo98gjR+MQMPsvRX7SPVGyahP9E+rDM45nWrTLW5nrnnhewtsNw5
pbe8Z9v2AWagTy0me6DsdDfHOo/HMnW5sJ1fujG4KtqVaZaWpouyTqF0JUW3qQ+Dqc3j90PMs65n
IseqUgllzNRt3+SHQ634dWhAIwhmVPHW1j7LrpPpfKnHCbSoq8ocTxxHmkggo3jlyY5/HHTzZB7u
YEp4u9BfW4pD+96aEvWiJExTfC3NgnjYrOAup+8k/ISbuZaRweGsLxB0ppf/oG8JXYKNYtxJ+7BU
nQZfPbdGR5PuxpmywgcFCJ9Tx4zo2iy9u0RIh79fl4QqRJp1r4sh2DkZqTehCNw+A7mWQBpwbDOF
LCullfQQP2EIaWecjqYClt7L1eWouAl8KpvCyx7dQ8nhjUbe0t865WYOyEq1oMIcDeg49aeg296z
hs/LmCgw6WVvba4/MPNOrEWyH/eiYXKX4wfjHYXqH1rxdn6/JAMKVniilVOr8bJix1AMa5MLZNbo
riQ4D3kvPKF4MkCge6k2a8BWPx2JdkVFIHxmYIc51xGs+TEiJhu8DE6PfaFbRDJ1UgrNwDE5v+qQ
XQ6QHQwPUZSfNG5q3mOQyIZf50WUoMnNQBH4uV8ydI/1pLfeBpJNXYtjQKqccEzYbhIxAEEXpf7b
/ZkwiSCEpHW7zXLrsVG2qVso5n+Zf0APLrITki7RYhMqDf0JGTumRAC3Z9K+f91L1Q==

`pragma protect end_protected
////////////////////////////////////////////////////////////////////////////////////////////////////////////


`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-1", key_method="rsa"
`pragma protect key_block
PWcRi0OI/wvi8XI8tqHJjp9nN1rli26F3cqVhhMY1noAFKAHaxIY1cKWerAlCkRTiZ7arEd36vZ3
7eOIQA0vs5zhGZnUH0uSELUAUBN8bAEbpzGVw2yyQttLRPdt+lQodZJesFcYvzxj/nQ2dbZnht30
UvXVw7lNXJZP4RbTKvY=

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Synopsys", key_keyname="SNPS-VCS-RSA-1", key_method="rsa"
`pragma protect key_block
pY5fbqP8o53Gzv1hJpa5lrp9YeMwKYV9AzMpRyfbwqXcM3nZG49+chGPcdJ3UN0jzrNS2u1kpvuh
Yca+NwZPscKSLX4b6NqokbV4eV5PwFsL+yo+VN5ruFyZ5Tsv9js3Su19NzBmT+orwuplIrsLbdnU
UATYRM4ftEsbbRZhU2c=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=1632)
`pragma protect data_block
ZFiwJwfwJYkWMLYxszLCw2l51YqsYqTMLATzct8r5iCYGUHVAmEe4FCgWhunG0yAwDkjPANLztVx
ql4Zs2Mu9Z71vh8YoqlcjHYlZox48W4n6AJpkbUtEMvnj7SThV7ducXPv1WXkN/mbhu4QbNp18iB
KN7rEAYKohAJbeB+//1Yk1XjudIFU/wvMiCUrTqlZCjklpr3faiV5zsknn7fLShu9f2/hFYkmAWE
bvpiazAPWnek8vP8XMDBXtdpuB0QmuGDYd+ERtaznbucyM8X1SXLwTRNH5AasgIImdiwY9J1+JyT
SRqd1TWFZlyCwmObxyWgEnHpNrYNZjCQBJ4LuHuPb5zgU9/rD0L/imrwaXBcxk+ru5PhlLvshd2D
qRHwEhqTiaaauZUyzW/rTSVJAPekOuDhXKnLiqZN94E8TNFXKINDVJXvCMW6kdgRqmP/3TcOCzl5
xDJInLlA9XHZitw/NOJCDxLEaIpxbKoWKcPP9S8Bs/idPw8y/eEdQ99qdFamYvQvRYNf+mcnV/EB
Myvd5ZrR3B2I9tNIwoXpKyAUC8Zzrbge8BizA8AUfO0qXSzvzAHl9UMHZEi7y7yZAUzH74xGkUi+
GFG4aPgiznzq67B78y8XAiUom1d3liF5XBFV+CjH3El5NgDTkZwnFGZ6vPEFL10O6vwu/4k4ZJWe
tofqYIwmC03d2eObjgpYRllGqUxfE/WbYWeCXPjWbI3Ewc2niSOSS1GT0Tpyf562aJC70rZiOavq
bkZQ2j4fJBIHglPIKCQtPvjrEtuKAD7wuZj82Q55+NXHstl40Xi+J7FNLMkogAeKv3dZhSHVfLLE
47JXOilIOLruVABsBwq4NfIWGWXwUfdseod/2lysYowoXICS1JdeN5K5esC8Tyk4Pn0lhIJ1Dxll
lvKidxmmKAMq9Nve1Rj4+fTFUjhORnX2AQGgkLdO4HcWWzCgPAHPL08ZGzqKcLv71zYL7Zesr/hP
veOv21Ba4BP8Z6TJPxGnKTAwLqVrHZvA56gdr/QAz78qUYZ4b5DSyxEZhNy7V9zdck5barzTCHUB
LzPNKcpVlFgtiWvN3dIurWz1h5QGDr8P6xBgQX6QpH60ydernswaiaxDqMdHTKjvtwwNS77BPYUl
1ZDJfqL9U7pU2JIZPxJOAAwMnDJC8XZSb7wRbl2SNQ4W3rjyz/YXPGWtI2WeygcB7yGlRyPpfjY4
Sibn+hopPNiKZazrSAK5EP0rsH5virFYL8lzDGBs+wPh478fANC5PNKS4d1T1kT1Qd+epj/xwLEH
40ZPn3HAhYuwds9lppkoktAYm+WVDsaKnIq2wOUWVW3TN0Lm9HqakxyFfEgIy/t64dJSs40zD0IR
ohbovo8vkE6RrRBNsbZVHxFR695RGbcYclP3aowt/WDX0uajcfooJwRbOoYhudzW/upRCGWLj122
C0kU+lQ4DsUdqxm7ucVj0ZFbxgxZVClPmp2dcTzK0gM6X/HhIgAym2FTwmuL98LiIKxVPTE5a7qE
4eq8YZm0Lyv028rDbUHESpVmeXW2045IrM5/TmR+gxb7qCjesqQV22PB1rtZVcagXGA2jiXMPyly
4G+GODkz8GChkY5+ayD1SL+YwCGZwwZQBHZq7Z/aaJ5AvMtfdaCBhJOFFP8Pjvau0cmUjDb5LBJ2
sx1P+kEpca40kr2RtD2mKIx/DLouYaUtNZTnqhC0TKg+gvshe2CToS173/h7UgeknlC4fo2S92IK
iOaIAwSLAT2hvUCqgWw2aLoLLwGJx/q2gZsi0hWM1jLzbPnjSVgfMmk/m8uSvV96cVdaVJdei/UZ
3dPs23k7lyvuPeSlXbw09c9ekBa+EptuwciYDEq6UT6h5WSgCvvc2YC0giAvZGP8VYuEk3s+1ZE2
jc1GlbbsfyTGADuto7G5TrYi3exUg7w2WzjfhcYZoG17N9yFoj3y+8UKL2ggDi2GnkXV+lXKjGJm
bIX8AeH9UPAQijyJ6Dm8+E6y08I9jg+a56wLEQuJg1Of+8+uigAkWOtizsaB6w5pNEmP2iqjXsN2
Z4m7N7xIZS0EWm8gP2UNW0f2EdMpoel+MFsYgMwypCVT47sLLkXgJzD0TIzHShsEMNTUgHMdhQWQ
DBrZKf5pjUBTJCWqQ4lcVO1WmZc64d2Vqj8HZd6kFvR02P8Y

`pragma protect end_protected
////////////////////////////////////////////////////////////////////////////////////////////////////////////


`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-1", key_method="rsa"
`pragma protect key_block
RAN2FBw8mrB3/N5y9K/D9FuoKzVCQKFxcxeK451UBy3qdPW+MPiJsb4QiDZS7pKDe95ZVa8a3Sia
oPRSqLGQgQth6ZmXeioQs/zxP+JSHXFkmRt+Qo3RKf0Zh1ZEMS3vKgcBDPF3EPBBTTLuOIOU0fu5
vIymhs3obqDd78xtrqg=

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Synopsys", key_keyname="SNPS-VCS-RSA-1", key_method="rsa"
`pragma protect key_block
hQebkjhERSu4ZCYkgwRdzLm7zg2bl6u3moucCqHjaZPLBlggPEtzu1mPMHcH186RUGO30NPTva5i
BnXA6Wm1Poq6oHC2yoHscs55vj/NEu7BueG7f2mlbQ3tV3kIESDTmLsQtk4VdI4PNme8mX2Wo+KY
QzroE8MKLzB6TawMgrU=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=9552)
`pragma protect data_block
AuYXlHx+nr80NSIJOZbi1IxmIgAhg1/a+p8uV1DZHsziZ1gd3yX7gy+JUUFGQbBtJ6aFWwMQsvvu
/B5iaZQUtgZoFbMpOFvzFnP3UQOz5EsAg4DkrDubffPn1mFqTofrxNYJmIVmqz3TPcy1L1HcRXev
o7CbozHWa/QrPeOeW0tKqJFvPB2pxtTm9OLPhGqWtXwgH/gFV88M89yzr7WxAsKCq0J76XmiVVY5
zA4M0lQdmRlJDrE4CDpDKtZcgcWmGu0W6zQfyp/L82ksCj6xVk3GzWvrysPU/RcryN588+C0wSt7
T2pCs3ni6y9ktv0Hb69VjptfND/nM4Whx1Iji2x3Ek5DO8UxyWYlFCN/prJhuUIglh4plPLfNcTj
2AB7/X+zcXoFXtK4yWgO6q9Xbjuo0Aa8C62hW8u680A9Hrk2NF3hmPZWiUv/f+G6aYZuK0CWP19h
OK/gwIDnqvEFxdoc53hPC9EtIkKWTBnXV3CuYQIkQ/XCLyQ1D3NoLsy7vSQBymyUAOIsXU6PzEuL
8khByzG3qukIugK6JdipkA7NsuUhiq+0smkANBmFuXgmTAdWZE15P9tOR2sC/h5e1VpNiAVcB/Yk
iOFyCHULcteLzDLi+PSd1Qvqo+7wExk8VrcZdERPLf6PnXW/Xlx+eFzWtfgVIlSr8gDd+ZV36VC8
tDAR6WgYGR/2bJ/BA0TcCZaUwRKHGJmHsAJskFIAvKv+cO6+Da8KA7sMFzflGGBPqzSsQ/F4ni9/
EyDlXZjsbvh6Lo6QuYu7rNumUKeGI2LdfvVNkr/rea1tce0FFmo1aqVmramq1mUjOLItvLsNSeQl
/r0+k+Jzo0jRTuMkWmftvg507wtE9U750SJ9UCC5PGW6AKIYxkFc81mdIcun4xBFibRgT6vpQH7z
KZ1IoePCDnek7njsOXRbylFUO8dpY4idufMT7ZEu8l5MRKVaC4zU1cdSDXxwbphBPRYXcsZm31yK
qy3+g12uVKbKD1mg2Nyx4uChVThVAWgoTn9HU4v7y3tlmahA1eXEEQTsPaKZAr9zo2EgPX3ncCcO
4EK9PY5bAazmPmqy6ij+BGgtKixsnnOaGpXL0iQaAsK/yCsLeKae8lsLxlM7YSKCXuBYG9p6e+E5
nfCHvvGfaoPxSO6WA0mAMws899xufbI8kUAbtlH6L+w9z5CLgO4IAF3WVvkrE0dxGKxETEKg5DGN
l7LbJtmpSZ+QxU8ELCDB+zHjg55/eahpD8tRNZpXys1Yr0YoXReTmY+HEce/cp2YUISwHuNBlm63
l6KZEmBvTpsfr4T7yewD7F/qQXwJ75wNLejmJaR4/Fh/xAoweeD+bSCRNHa7u7mMZ7+GqJurs6Ly
5sxZo1A46cQ9pi4EfmWsOlAfK2iYOls8yUtl3bwVMlmeStTNDKI8869yE8+RTa2AjUuHdmS6/KE7
IX6Od84ov8WqOTuGUCpsACUlVUjpMw94fR5w4Gew1zTKg7w+VlA1w7MSfbmB0Wd5onjZlzaVP0Ay
ixY7EI+gircUHk3n+EhDXFPUGnSlX+Mh2WTQKf617tQlPsYvWp+lfLN+y8F6xa6S9w9GyQqhzfsS
mzOmHAWFSFL+u1Q1l2d5tBxOfssMr2/CDmMkAjOUlsSibdLbH8dSlS0Ju2C1HKRG1HYrjcGvamuj
kDqS0JTVa53op6YaUXoK2af0FKw5QIf4XI//NkEqVL/B/7DweKkfDDw+fKVoDix6FXvvI8fSRQM3
dU5NKFtAJ2bHfiCzdabLi1WiYT8HNWGsYvFuNFO7rdIOxcwjRd9JkRZ9n6amuBubO5/oBnK+FxlH
kFU6wp9/VtOVDBACO2sWa909vH3IYAQxMUE3qN8IhBDhB+DTr4gEPeuiB8Z2KmEmCHeBjUp0JrYI
d6YRjURl6Y05KhR+HOMuffIyf4Gfc0lsEQ4PGUAtPuxdVvqdSwNfH6LKQ1tM5iyvVeIO6ocMDcW3
cUdZSjZQtIZM72oeJLCxpegxb6JSGjDOsnabo+pTphsFloswwlbcLgBAFzluPCyx0Bew9Uk2MZPY
WBNqftHfyomde1LsfcMo4kiBe+e72OsVur5y3khsV11j1g2TCCPPRVsdUcpfXJza8SC0erSnglJW
hChiLUoUubBrbAuYmFNqLukpOy+Oz+MCTyMfzXLJDb6pqKvF4vIe4ZsjzpQA93UDrE1/GXIxWWQd
T7cyhlGuodihm+OxI4hKpsbs0kTualt7SGtbevDzZQWZLl9urBhorQC+Rn/qoS5T52oLyoEWr1Ev
fT6uWPIn/slJZ71/Wcr0+sHRUTKKzT8VJKdNx3NBt2LoTC399sgp4C8bYDulMYzqB65hYqOqT6Ka
ElNjfkTKdoXLio0L2WpcfpLmpfpVFKs4dgx/cg7D8caRvnS4Sr53BjXaqIHLJ9PEUJcU+YNmh2T4
5jEH+UVt5p7EjyIbylz7Ccs8c0VMff8Y94jRYJm/L0cmu7gx0CD3K3hbimQZH2SgSnXB8i2mWTvB
f+gSlsWlIu6olbUkC6TO6rvqTUkdxrRIwnnWPNI93vCdXTpBHGz111tfuRK1vlqYetE9y5HY0+lX
cXvmuIvTHY64LaxqyaFF/9RNQffWWyJ7fPfSWsyqnLoll4WgGlKsllswv/LUgBFAhsIoElxj/0FC
a7uj+sSlEk4eIrEcFsnhGoSVBNOudWgLOw0sY8MKlBDWpPoXruC0kjeON0BLz8wmucSbyE1bPCdm
Lce1lKTKgfIiUt2fTWaasL+LVI+lndAXm2MGTnT5ALNic+pMWZHBPP5WLdJCeJf3SsS3sb8HxBue
XlWCrn1htBrOMQyJVZxjMsQpw/w18+KP7j/WwQTSFnUAIB7cvo+Bm2LV9PBsyv/GxXXfWRFr/1CI
CtHY3HwJJF6WmWaim7XSZpqjas5rFiuRz47ZrzBMTKHZVn6o7FT2nweC4v5yrzfF6BCBb1H0zOGk
/y4rXQs6+ogAEf8MZG5J3/rj8b/3rOGzKN7IMN4se6bM/fzxegLc9/E7v797u7wCD4JMWh97sKuS
1OeEKtUZWFj2r0m+6BWORgVZJSFX4EiGURGuP+8ddU6m9JQTa4lP/HPpqKW9saT9eKuPWBnhZX4k
GQfr6QGCgy74JNmyHc4XVhyM2qdJJZLv+8W5WdgWmqSVqYtXJaKnfsDTj/Fe3h8QloQwacDsmLbv
+Vc9fS6wlz+mCzTMN1pSuP/D/uxBZM/2JIjbPz4Bioj/3R6tbT3c/iVqBb82HX5NJld2iAAbxv8b
R9gLKV03+EIFAdJRIaqNlLZtwHxcl91XN1oQZ0d+KnI9vZzcF1Rm4uWNVvtPbEFPBZNIaEsCaj1q
ZPk71NBQcycqIlPVt2XB47M8DNNdzo1XClL/JKjAydOo+d8voUzmhdu24XtNg6l2EFJmDVp46hFK
YJtI4danYFTzJfIzsiZG3ThQMAktNxQUj87qHq9MJ9qsTMm4jxOhOQBL3EIvH3C21S/6YegggAz8
9KvhXqQw5CYDA/cajLaFWZZoWS1vPEvTx2XVuNW8RA19yd4jXqGJiajx9qOp1cC+XxSxbF1q+1Zo
0EessD2cuxezcENWHBbq+/tLGcqF0zR0itnG5LLak4AYKkZG+E3GGyiQ6TaDq5z+9eayCTdftoBt
c1tDkVKpG+E9Pzo7RFI9qnubnckQ4/7/QtWN7uGfEy3FkXTdZ+etE5+34hCRLjQjvU4faVEULPNc
Eo1vXK+jCWE4MRLqTPWvS0oSaN/FFnh40iZyP7IZJ/ezB0NlpumJb4otauSnDRpZISXU/xDo3W4w
9cRWuDRzNLgyiSYsini62/mPpWKECIMIUsUTXQFhX/KB97jaoapM8k1vFrJOMXPefcwHnl0qvMEV
5KM3TyzBRlC9UhdT/MPnrDKgeHuS9IhkXoYPr32hm1x8hA1tcuk3C551+VHO7nrcHS5O3Pzwoqiw
UoKmiRx+Fbc5BsAhVLMJ1rXLgECi8k1uxKWYYrR4vxIOXa5dY2Q+URr9W892lCCZ592O0muVALq7
Yqs9XN4YBiLeO0EhnaMLV9Irq0Hi69SCcFoMsMWrid65REkltnn85/yI91jeYOy1xR/YpBkMG8RD
HFVxSFuBD/FAqSSZxuqmTK9Dt5wHOwv1KM4vG6ZQfEmb6aZhhwm0K8+sor070lyAObTEGT4bB9OJ
tmpOYgX7WnG+XEdFlTOyJPuKxo0u2AoZQ7ZVhRs7tS56+LISdRaiZ15/K7lMeeK6z1kSYPwzu4NP
1kkYWzuByCV5tOuIRlL6Ge2PZtY41mffhkYY+qBHBSo3VdF25bSnOvytDNLWR+ZOqSTwkZT/RvIF
xdnw5YkM1LRxoRcfmZYfoNqbiy2Ocets0xODWNba1btWBhIlhaTOzGDaYhB8tbeC4s/kh4W+F4dB
ROlzzvHAGsQtFHZbBO/dc8Oj+ACT6ZNpHwlNg/eoc7vHXNIY/6paweMkFDrrGZEOMKizcsQVLzAi
evVkpohi+U/Mk7gFTMq27vc6zMOzCLRShfOjZgWiequsOM9fZlaXUAG3z7dDgxHizgFjlHjriRH8
QAlaBGjffrR0qHiODqTycLZ91YVZKD57GH572AOD08PR46SuJJJRNVPomfL2qni8rNEWQtqS/I2j
jccCYmka+Og9Ts7R0fVdcQjG5wz69CZ0LkJXh4gG9gwj7FMgnoxC6axuUouteWpGebS1KjUXMV+s
imNUFaBbcYKie8qjDOuTz5mg32xSBTJfsdfbPFR49+w9yUbd/TW0hgBU0yPkOgOE88fixKMyLC+8
bsZUtNdvwtyebCzYJQOHEVMKjvjijOGuHAErT0MBkZvwXGdI6sP5wTQTbZCMX3fACLTZKfwbq6s9
+aVUoOig5z2OwM8dkZUKGPv//RCD6I3rMWp9108uP0XWVt0RfSooQIviAK5/ViO3mxIis/DQe8FB
NPTK44DiWEdWTtv6Gs+pAJpydjtQhDuWSPVHLyDcN1IoUnvSCt03J+06n0vZDbjwaStFwmRtxrOM
G2GeOe6ayeZQzWRWSbHbVNnP/Zm+4Ywlrrk59jlPWvpRnr/IdGkWFq4s8qwhEO+l6viRXBbk6V5w
tXm1E4xRHkbSCwxyz3FMUBHQCSDkdY1L8OWPLPInOJh+7QH8yTV40sD3GfG2XCqAf331Wm4DEFKp
sd1poodBhbAKxHBv9GatjrKVrDHVI7hdDt3erKQwshmIq5P1iFTwULF5Kr8oVaRYOAFrT/B4YCUv
iOkkNYxyHIPgV10PumIiUC+53a5CAxY79dWEmS/DhtQdeZ6WsnEVEkNbKq5+JyaZbxLYRlKVcl0/
YUGmfG2xAduI1C4Ysb0emWDEXs+BiAMERPtKGkDnvXRvbAXFAvfh/q7Uj7aLLMVUXQvmDJdqPcPk
NuIlydByONdlRFUwvai775F2LPZRMoptjVJn2A6yjAbKAfD/aso0O4KL2JeR9yFCweeQRTXSszna
rc5a7SYtv1uDoi2dB2v05l3PyJk5qb8DOtV6hC6Ychequ/JBxVtgb27LKilLugj4ig0v/qKvoX+B
Ra1tf0g5j24RBYhmiJdKj/cvcOe3Mn/Jfu50DfYScY9m7qhZXcOQ/xY9OaWA7HzvRHpeqqyKasbv
OzOSem9a3CLVPMZBbDSUdvgiAiBpEYD6Ibf2BWT735MQ+yMoQaTfsroxioDM1wGCz1N9Fah4KH9m
MGSqimTaMfDcBVI4/ChQmEkp432rNfCin7HEoBH/zSMlgVZ1aWtDimJklzNW+779YDCOqn74628T
/XEb2zQVOV4e3cwQ12eeHv7BylPPg+cgRgGDn3uiuFF1XijVSQ28ccKMEuIpXyDE4Z637oMr6aUj
uhrK2qKMZje+FiYxSE+2DMnR0y267XTQ/lWyMwbCE3MxnNGBJbBTmM5297Ef7VkufKLgPl4ImGv8
yLE14ZmVDUHmnvd1cxktY57UtSaJdCbM3+kgywdRZ9VgHhfJxphpYPfyFYw0uxQkx/vgdajaVkiy
wSj5lP+bhqH6vslhyu8aVZsPlndX4W+2Rn3G1tOjMLC56xw28VYOLAZfiviiH4pJSMg4k2eHFkei
t0YHAbz5LDq1UwQfUrtGOne94noXTkXHM8psFi1WGKpnE/+r9EbUel/KnDQnyoK+eEDrwO+tWZfW
BJTD42z7Xxay8MEhHjlg85WpkzOCCQ+rEhdPtvmGrEo0hlte80OXEl6uH+SdkDOUnHLd7Ypau9Px
eL3TF9sjR7JM77YQ6tYpv9Xb9IW6kUzzcXQA3dzbe7MTkz9Zw3k8EY47i4tRqyJO08bTZuF4tyGR
+ZpBQnGpVi6YodxOvziBNCgC4oPu+aJAQmflRjFIAEMcgCVmEn9Pr5c7Ov9sE3Vet/y6jD+HRXXm
760hDNVG1QiFrqqlAVFaLh3047Gv2EgpEFxuvQJY2k0VgzV0jBY1k1yOY8TbHUJJ9AuyFgljz9aP
iMQnDVpkDiSpbWZ1ZakiS/NAdDyudGcgUI93R6oU/dWZ0ten5RCoLyVg1ZR/8wbE3eOayaxGoC4R
vPnI20zdWQIhFhjRUA4e67ToLlyJKxg0NOxxII/qGdpZ7bgcMdR3rU2LZIdZR6IpKbsZ38RJzRZb
2RP3gWSjfnv/mUFgKQKWl5D47qnYvsc2Fh8fLO3yzHnwsMl2zJwHbEtrYYwQDmcZ+ROT0SrD+u9X
qeYQGojP69jqRxxLTB84pQEVTcs28I2t4fLWDbfwmBgiEZoLcqgzGsY39e9AqgwI6YXPtl+Imi3c
Aqe6EXt1RRgr7+4EJUI/mhKf+OPjNtDEnI20OHEo8NSGLvVc2cnQjVRWWbs1T3RmmZLgG3W9VPtK
VBpWfkzxFMSNUBVGPLmQTNqBKacFYxhiLi5ZBTJQTdiVnZbd7pJeW/F38Txze4ssnuDkwU39zG8Y
GmoI5SQOQnOdFHMHvNh1/F6HPyiFS4B/x51BRwGnhEiVnxCx1ArCNd/zOFQB/gpxMXIQQZE/asQW
bquVWWjAVeL1q7TaUrZGj/Su+g0y3kiQgzCK7LRh8+T63ZtWc2/C/fhSD3lZYbTiUnq8UEx7ytA3
SPIqEt+9bUU0Sz/Gd2vb8Cfj0vWPzV903yJ1x/LGYqukg91EdmmCXkWHBuH1bNMFNCkdXsUdOaqB
dcX8I4qk6m7B2TFW7l20xcCRTG44P/wuGEp/fBz2W/WUvtVxbCcc4AA1Z2wQvy0Usm1Tg32O15rg
hIeKmzHPjbp7QbyIed6m1YZxh3vc9E8gL88rE5LSKzj7yV+5hOW3XCBwgWNN6U94O4KxX8mUuipH
Poz4Ok0vAPBC+EqtAsP6xVPhcJBOiFiy9Rzow7GNVYmyAEOSjlXMYIZfPkY7uGnyvBschPe0T86b
1tejE1apAb3WhVYfIGrD7YQc2G8+1rCv6bTdio8Wwb7LuvItB8eAKQ2BxC51Tkjq2qiEZ6oHe+h/
uYv7sDUxA7lW0SxwYxiSqet02TACPTGu1ubMKC+CefgQKjqn/9bJX0hEi2VQcmQOEHJ/6+/5Kax6
mh+rgnCseOepcHtRrErD00QXC/nXM/UAMyI0zuhYlW3O20emFPkGEY/Hks64U5V1/tU9raoejDZu
DtgC6u3Stcn0ixT4K7di7dCtJo1QHJCS8v2ydppeTapjoSfr59b8aUB89w8pL+pB0edIgIqXSkLr
t7xyaGNhpqzko1p6fbGOl02peNlqWwMurtu8nPlZPg8b63Lip9FqItPkaMeAPjAiRcok7/4bIEZQ
N6V4OFXuwCBGf0VqX6AIhO4NVTCYFFl7/H+6Gefr53RsqMzk/Lpmd38aW2E8j7BybuD/VBD5ly64
ZP9kNK5PBgiSyIL4Z1A0dtPUE1sNm1Y+ByYNlXLmY/zjBeeruFelyxAHBW7i9rMT2F0Bor302Rmo
Lc7u2E/MzPk+i+e4ekNfXfkP4T8V9rplr63hmjry9eKpqoKCyvJUhrrkW15xXBU5iRdiBkorPiDf
De/d3kR89W1lNcaKZ9/wFccHY6JDaTmXTiyjQfDEtc2Wd6k+uSQCNg0cJRMZcL6w3O2FluQkESz3
Cj2ZPBLiPuet22j8dhOMSuA9XUKuLJUtfYE3nAUq8u/tAzDBP/VJIOmE9ONUjAdNJgkQQJDbxD4J
AH9dEnGANkC51oqq295g2djhfBKvd0V7uVwGRpqXbaNALTTA+mNYuCMmpmti+xm8WIQtJf2INDyb
CFQNGBl83YqZ7hsUvqaipT9YhqaGC69jAYhrb9fSPc3EDXquox8FyORNAAnvnjdRsJQ1uL0zgaM9
/2joWAbl0iY27WpDzI91BlHFzgYE1Dtv0CHUqcxjob9aNe0jQuPnAA+rd9DgBRBmfCvS+i24pR/W
ZfaovN1fJC8dF8PTuUohH7NaEcMOUUXMScuFoH+yzJAWNI7fNn+268p1Lr6t+jMdEvm7IBlhmj9f
nUXPL8FDpsvkAI6QGg/tLamlIT+Esg5VNOSy5DCPm2UCbRlJt39JR13UL4SI+Z9ex4Dnyg5GGXGP
aKou68Nk4NLHzrB5ZhG7TjG2aG97XTLFplQtWO3tXI+3hcVCbKvPUMccobiwyYhksLWASFPU3EIH
OklxazXKrfz+SUrgUh50jYUddeoKr4yCKXsebDpfr675uW3blTcgl2F5tgdeB5/utDDs3JOjHN5d
YTgwdUia2hPwkPPS3orx3vztgBbtMmBu1I3w9vnXFlUEho9bhUGaYnmwWLgZaA57CmOgVftlmdYy
4xvqpZeV9HpuNsSow5pWBTEFfuTm9bSbgDu5wLGjw4Ui2Ez8wP+aJMiY9b5gigKhfmid9x12T5fE
akjM4qBClT3SLZxZADV6udfgnXVKVHUcyakj+sDZgDDymV4b/YWvEeK3m0hP6bN+JuQMi7cE+fGk
QIDGAdqK7zChK28Gb2kuNGYbm0Ik9RTnGIPg+M8G5ggVDI4jtrHS3FU1xncSvk6++ergEc/aHcq2
z17SHj2Aka6J+jYJikscbBYTB3UT7y6VXhrrMxx1NAY4FAPO6r/uBJiCfNzuOi0ak3P1cp/WyI4A
Wzy2oL+ZYBQezrKZv2cnBXyZJBJ3r9wp0p+OOHMVOfmF+0Uu/XxpryHz3bv6ZP+CGcSNuvSTPEO3
DsldW7silmLTrDMOXs4hqD6MDII6xjn2j0uewWy3luTqab/qyu7uhzSjHwLhOeHFAdMAcuqPN3Ip
GwwOYG44euKSAb0qpp+fLalVSGIxjVkdawbvLn0fgUZuBxpN61nv0I5aEi8Jh0Qu3UFTm86enkoU
w+BwWq1zIwFOuETXcGEg51jQ8EpL/ZfO+oT8xsB0oCL0suJKh81E7fCwBwbIqSdOl442Y/GZQIlJ
c/dGqu2izOo/J/iRkWy0Si/zOar8sHUNcY7tbQRed7KVAx4kKthbys2Bd9MT+Q5X3uZwdS3PHUZR
mGPsNshlnCnL2IRCeV6eas9foyXHGHO8Lbyto3mNi26czxPXqUMd0yGdEzvKM9ecjZXsge9SXzog
pVdZWy2uSQO50of9fRDYWkhyl9/pDKye4YbfDkwVWoUW2mIb6NHk6wBE4w9Wj3K68rXWkNu4R5Sx
VExbCqITdP2NmV+l2uuVITQjYr+iELWvI1VvFiU/i2qVBoclcyxWlPSQAeFYqq/RZc8RNYIoA73+
uSM8J2D0UZ+Q4RTbNEyY7PK2LFhiyDnsSXS1YlOH3Y4tQigQEn2QavgZviRh2k41okfr64rf0u0j
3/IVeB6aFG7gp8lJii6EL9OmVYF2K3Qj8oh7YfRPMUP6GlO3iaHArmla1+VZDwbRF6Q2fC/mxxCw
x7hnFwJM/PgcDgIIEjRe8P3m6giAsCoAFrJS3XJiis/tjpxje2y//ujA5IQ3IJk7rQqcsRaHKqkn
baAdpnDBHzbIVk0isfbEJeM5ynqJbunrOBI/F+xFTh6RxN6CcCoIgXwhCEO4ORmKof0bU7MXcr3Q
GSojIdLeg6l87YeOh4bDPPZUjJ5Hd9t3JoWvEmp1a/xgdI5zWdPrK/AO8G+Ps+LkJg4cD0RWdZn2
dEDe9zJVefltjZSHPosPaPRmmY+Le+Gu2HLLQ1LW6Ure24wqlrJip0juiXQ1ucVX6gbA02uQjEhF
Qso6X+LBgYMPMBsyzpJatl8V7dFbmE2LX34M2ne8tOv4I/Mqwpod/9/CZiqKBMfOydS/T5Anx2LD
gXhlxgYygkjaog71hFRzZ6AyPGWYXMQXsrtXzFnO/R2/Ab2oBVYxDDB1jTV8SRS1nSKLYNRbghqv
qKc/lo99mgI80aFN4vNXPw4OvflD8j5icXwqxq6j/Ns/De5+t/Ffs172TtTix0FMHVpLhhKeh1gx
L9TG5xV5MIvJEsYMB4y/+tH1JJ6k78u3yg80Yu0gXUv4gGvXf+dqxzo6oIvz8YWGqSaTY/SBWcbU
YZcDmupMn5R1wWCFtXqyCR3U9vXl372pzfdsvEGyRzhU38jh/hC5J9oNch4ModDGXZekzuK75iHq
9XXj2GNM+KZxkF6IgIF1arcNLEXnvNKy6cMdko8EaXT3dplACobmhGtjoThFfdVcl0xZsZI46meU
z8rhIvbxMil9sjzxO5VOwhRnh6uEYAXr6p42G0WsqvNLMI/ygtQR29tUp4qxLh/qMxErdoZILriA
eSbUqNIOsoEysXi9hXJnchrfzbNJf8+oxx+27zp/3dUUgyU6CozCdu0G8rmI0V/urisuWCJZeDn5
0iflvXtfGMhY+bC7CjGahMDwOVxyii5T6f27pvh5GWFDkHpxSZ57u6lT3clKLJqH4adDEE4IBi0I
oSqJJKAbl+deojybFAwLngp+U0pfqxqZeTiuFk7TbMiNwlcB2ugHZRgiZBwNX08F/ufW/bbkCE0K
0fOaggM3cALjT5uExhPi1LHEKBrc0nAdJ9GGrApCvwp9hN5S2ru1obI5BBVcTqhgUlj04+xsuGkZ
Cej2kiDl83rqd3EcJr6MpiOAacis4Bqo1QNCdMmH+C1VMxRf+anjjbqZHot9r4RKaD7n7EU2hbyv
zJwPCOLOIcWJ8c3dA8S3+cm+/OCXnp1jxUIKamVbxOXUVCbiwWn0Zx0FmuB8FPGQISJGTpi1wYvc
yK+y+zLmR9lZc4PyTVkHvOaD2uuW6+wwuexRROigWpW7+SrxC+6iJ1JPfKokG0D7tdmamA4tZRHN
gw+8/rhhQ/d9OgA6/DLMr4mv5HlTutE9f154EfumEVQkGQMfHte1meHNeDM21eOgCDEH8+RnDCEK
Kxe8RIFk7CSiU0k8ZPdfY8CJptATsSF1SINo/p0C+yk+cjLtc27scr/UcqtBafe751i+o4CemKJq
AJeVebmfNiSzytoqbIugGV3JFLD9DNACy9IzTGs4LkxFQglsTya2aTjPz0or31hLXtXjwBs4CnW6
7vWEOn5bV8EIa5VWg53nYSf4581GeHTHkpc6Vgm0kKd/S8Zt1Y6SVwZlSKMVT5u51ViYN1D1ujU1
oeLJ98e4i43Hxapr+tj0JtX9B8y0mnzA1rbsjRkhGdoazSasXi4gov09nY9tBDo1kJJprVbZHGNS
YqpkOqBqSA4nVgHNx41cb+vFu8ti64PjCVwHhoQyqWLdx1e1hdVlfVx+bcxJPKCLp8SEEo+yvJ9F
iyNeW9Mkbd89u/rWOlpurPI3jVBzHwjHoE7+JNgzpxLktcloFlRXgPtSUecFaHvnGZLd2uWAcSSj
JIcKKU2gwPj1f8PJ4gyHhdsOnvpkEvNIS9jbpnQBzSWfNp6fLVLbwLAtW3YAzs+aeewKOQ6QBcYg
VM0Mf0+QBS+E7b0isOo4pgoG3H9nhQMm/m8x0VoY5zViIjZJgFITaNjo31qy7XWYrVX58AdCMgO1
4vkxUkkOCyJBByLvCqVwx1ph4EKDtozxfSsndE6RDY6eMI4nfkRFDdo65g9nuugBp11vWirse8rY
B2Vs/6Ewq/n62bbrQpQ5Uh4iuGknxzBvkhngsr4i2Sw2V6wbWi4cqf+SLDwboK3+ShU6SSABvTAt
50TIOtN9ZnoNqcDJC88uCxlL99dqcyK+9dDl/2BR0dOe5VG9mez/W1SS046nSvqklKLvHlxeI+ai
1Z/qK4andvShnYZ4UI/LqvVrS8k6PTNCR6QS6iqZC1rm/tPqqckdRehNpbzMwFXV9rN8ONebvXkf
hO762IY24wxVy9HBEm9b7lwBeglL14yTnuClN5KcqU2pvx47ocwZNMo9vN+Q7w/aHw1Qr+y4be8x
/EhEroWVEUYJrzIrS//sWzFbI4zkcQGFwHIFI+tkCO7I0mLFszqigLMvgqSPfMQYpEAMJO9EU1Lr
5AJ7jhrGTJVZ9cPYBrU3s41yaXNdJTFrax5wAkPzgsQZl8DPBCp8lAgsB6F3QYFmD6IOXtywoeqV
ApFL0LukKSqXW385JmFpISH/cuj5NBjsJUXNboKUhiDipysgBqQz8OmB1/oQ/o0h7ot1lbSv1kDG
NoyqWJjtVd+UqeEcHqm8EQbQBHAZmkZPsCtw90MJRQpr+/msQaG7NFkSnhWtjKSlrJv74BRXeAF9
EhWO8SSWKitxT2f5ON70hX/97oHf3TgE/NVSf1Ncyu75mgg95oCq6e0xClRtq7tvNmhRZPVXQxxc
zxyIs4ku2ZFE91zgNYkBV8g+Za68vGYigaEovl3ZldqYLaz90iA3BR0aFKfV1qWWNUvGhzu5UU9s
CGVi+kB31NffTMP+qkAL0/mrqVK+uFLpldSZge+Cn2le

`pragma protect end_protected
////////////////////////////////////////////////////////////////////////////////////////////////////////////


`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-1", key_method="rsa"
`pragma protect key_block
gNFcUfwKF9Uj5q4dBL0ugDdl/ETLXdHHRjt/zNH0rC/dEkg3vie1jZFVP81er1Q4DGNnrgRSYsZC
RqTTtZ5rK9527gZ90nmVszufYsre+FmLbof40BMurZ/wXBRchf+bVzIRzjuzWg/UQptfnulVyReR
+QXQ2WgFRxAlfH1mq2U=

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Synopsys", key_keyname="SNPS-VCS-RSA-1", key_method="rsa"
`pragma protect key_block
NhwooTBnjqhfmvK4qgvLkOK+6r6Vlo3SJ6/cI3jIyjxDI3NpuiGTNHR+QowNZ9iKg2gcgAibPl1m
M3zPcR+JGrHeTR+jHZATovBKTQvJ8IJxoolJh44DUDfj6hBbVqqdtQuIMoLeJ/5AuSVGOAH5Wlna
5Kvbo7BLcS04jGqn6IY=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=1120)
`pragma protect data_block
sYnl1uha9e5XiQsdx6VPkDKmz/dDaEtQnWbtKJDYa8yS1uMJRItjD2Y88e82601FCUsBxXU57V7H
JlQQLrE2ZooZs/NcYEHaeXhEl8+ig1ISxmTqO6MGTJ4WPi3kIkDGuFjMI4QHLIagHHHMRz0NEgs9
rrRe7RrNkKCnFGzP51QviSOnU3Bv9vQqZBnrbb2xs2F/r5AXJXAheOBBOOMhqXeKauY8Dzi5Aqxq
nwSTPhK23PX56oLKcVY3Hh5J3aZxg2Mys9H9dEbQFIKqQWsF7xbduR/Q/T0sImFfPB4RZe/BCnOL
3C+n41Bj9NdhyFRE3IOsh61gGP0aAon54tPPBwo34TOg4NB/eau9ZP8AVvS/7U0RlpsklEYISX3P
ekUkv7u1/6/VyCxGtL7eLK8rUVHpzF81H6YR/9ss8kY0u0YpfMHO7ZjAzVn2A7o1zcYEf/txvpm7
c8yg5SgGTxjiI9KuMNMjGoZpZ2Ix2mrYlOS+PH0PXZ7SzKU8KvtSFha+fdrOAmxxUuEPd5yXWU1t
16zY786UExeHKVvMXGVhfA2sRjYj7433Tddc3+Now/zdNKX1kMmtXidscIZkkiwJLhp+F7Es54IC
2RRSeRSvLVSugdC+1nYukPk9WVkokm19aOT3/MCRxzE5sEBOIRaVkX00wFOpTMkmLat7ZWOIFLjj
TLymbg1HBbOt5vkeQRdJVxjLcjQnepN/xb6/XMUA3U6aQ542gzK+7DPRITmO9BC4SXcEIY5FR42H
/CtBQuKJmpIQwPCjdd9SMc3TADKACQvpoGLytHjGHJRcDGmP3ZhapgZ3VCM5oIHh/XQNprhkdN6e
VJ7aGCl3uFFF0p3tIn8yAYP7wxePvCYZsXrN7zVYX2QUpMmtgE/ZV5kdlZ1x6BKlDaZhlCxrxZzK
j6E6RFySMj5oS76Mix8n8K5aBf7IYdK37DErQT44BE2b9iEXECFPZ6M9+u3xEBwhXiIUMS6UbGvW
mc5llZy10ehr+q2Q3RQsmYNvadJuMQD8R3IHERdkcM1kpxreYudDPEmnFmg8S9yGel6f9PDaUGM5
N5uTG7JfbWAMqKYWft2+7iBaPgPFBkqjC9aNONGeZJIilLpR+PTVIwhN+KG+9PM7Xzz2njwEzszN
zF07brwtUNtIxO8S8rAlApeuhppwLZ7WZxwgAWAKv4/J0MPP5guBkYx3tpRt1+oH9pz4LJUGrxC8
D1ux+1UBUnBj+4nr2IMUfvOzVTO7fKROQuCc2GKj6kT/VTTIw6jpoDaECzRpOTzR343yBHuSwjE/
DdsWtDjqEke1I/Hx03vQhoZmca/emPwp+F1PGSsuOv4dfPYyXxss+K7M2U4jD8osMVQR5jAX/tcR
0IB8vIwnmzMEqArZCJODEY/0xa7gsFv0+i4c3gQvU5lSclrOqVEdiVPiQZ+bIhCwVCRvNuJ89q5k
bPVosKsa/Rs7WASgb2LSobcaqCGAc/1MTcdFaRMvpZBLADUo1Q==

`pragma protect end_protected
////////////////////////////////////////////////////////////////////////////////////////////////////////////


`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-1", key_method="rsa"
`pragma protect key_block
noHXjRraXdNLvzuRwcwm7xCPM69deLAm6Sp3PR2eUwwboh0r5hGA8k1EcfIzvTWDmA2UuQwsfU84
SNdSAEGeIvmdk4vpLQH7tMBa7MfnOmgcJ8jEknnjth2RgKJgRVZTeOObF4vF66hhFqKSRnJWENJ+
YWYPbVIHMLtlHypBQdA=

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Synopsys", key_keyname="SNPS-VCS-RSA-1", key_method="rsa"
`pragma protect key_block
O2CEe1aqv6eaSqPXuT+89h8kTkWKNt29RD7ZkO/s5YaKPF45XOIXF+gMXhx9RtzbNnJ4aAaYf0Vl
QvWr9+2Qv128fi5W4iq6k3Kl79vN7T42THyDKK4l7iea57Arl6+ZpRqd/YUZUGsR1/AgNFSoNbCC
kNeZuUc3mjwu+SnBAtQ=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=6208)
`pragma protect data_block
pDIA5MhAgmyhkHdWCMGoRPck6LT1QvGCTAg5CpUVOcNojKwlRDZ7PrVP3AOdT0+rztRJdY3MwHAx
UZtr8kKyeegbHAcqYQiZqnqxFsk+QbPnbsByitu0xNSkqtaScglyU6yAgAOef9BI09x7OMJgcCc/
zkU9wkPxWJqyI9MTGM374RQRlfd/axwx4DJsbvuESN0QWZXijX4r4NTUpXO3VbQCNmy+5KrLMziX
bfpZO57z6LtNNmv//O8GJ4jfTOUlD80mCu29wwJsNuOOWMITG2jniZjhBOuMo9hIFDyqntzIzG9z
70sTFvXuu41qL6w1RntHN/iLoZTMTJZtwM6HjaGPlg1OSLnv75BJuY9Wxcgep1fe74pAWGRH5N1i
Im6jHaUQ8amUqr6YKA3pKvKDJvVhkSS02pBFfWb9VPhEK8PRXxIUWKjGuBd6VYKmKWSup3+c+JnD
M1rlgakQQ01VRPZUGNLt5y5UxizeqQDPaG4aLC5RcGJ8rJvpEJ95gwu5t9S7iw+XF4681NrB01UX
hVSneBx5GIRCPnrE+yn+hI3AsXFvTZ5KwSP3ckGGs38a/SaSfJYmOFZkBnwZRTRNs73P16pkuMB4
URsA0bTzk3Q1f1ERbdkviEwniORnXJy7TqzcDjGG9ir9PH+MHE8P9hTF+h8lEOWuwdQFQ3BGD8VG
cntHUX4rt4he2GqyaoHrdBlytNf1M3tr9pszFo8jTTWM8hjZREcZKCqGkGCRgBZSFNDfODauCK2o
ulpQd0D7SzDE8u7LGL9oPX1ENp0vGALoJY22krMxfgqSHa8kj7msuO/mMsaFNJrsBeKKaifhk1iy
TnjKxZeEpRNdLQNtaB77KFX6mMxQGuJ4MvhaQRbEtU4fCTCbfD9+YuvLzp+UYhKso4vOvPMe63w8
wkIRF1w6IXgVX8CpKgP53FmgfrBsqpy4ozZ6BJ21fEIdyzCsmuSKVSJBrRXWMxMq3Ui9J2kksH5v
Te+fpg8Z6WkJ2jMBpm8m147Lv5FSuZY/0SuOCk5Pie6GPDRfxdRZthCMmYVksLLsjV5Fn+EQiHzE
so+7YuislsCnuuomwHInJhhQIRlhDKUga6Xaoi+VdJJzf8Jn0PujUKF+BkjsGfh8rJxV8ym0Sx2w
uLiP4Wbdm00T/ttQ3KKD46+HxtgQdMCwFSG3KYqnw5/OqYdCCz7mfY5OzhMDVaIPRWSgcLGGGmYe
eaQSrhLbVOEsa8+NMLM9KwFWFgNxeIUCO0lW0Ot3nv3jtiF9+4f80nOm8Up2KqWl9LBPmT8Dci3o
zr3uIR1SYH5t9SxPs4g4P4NnhuN2M+cW/Wy0XpKzCSoOVcBdnRYAxILxPUoAxH9EBGMi9QJ0fWwW
SM2Ji+e+iyLwb6VEPpS2agSeYiqIvVoz9aRzsYLOLglYYhi5wuBwH683E+xk1BSSkQh8UXC2c8cr
O3+oD9v3uXQGzZOB9eP8WU5PfIXlfUbzdxz/MOtfDdlmGdxuN3B5+CqhVkum4PptLhHOnefVo4tL
ZZSTZdvRUtYQx3vlGyTLeRrZWBs0oXuBwhRuL5g2HUELML76JPNLSmt+g6tLlTKPyaak3P3yOOQW
go4RzeYyWNqxpQVAZt5IqVmdk2FD3M3WH0QSvBeNphXrZoLhmL/3RAuxYMQBfcaDDofIl++i0/AQ
avNwEX5b6KNpg0vLHSdF/+tniIjwCZQ3dv8nB0fUXrSVMSLJWxyblWV2jVE/VvhYvqzzRQR0hKPk
AAdm6M6UliOWUwrUSlFrgwKKGNPkLqpmpOtplc3gKev5NUHQrZzfFiYSk60spK6+GRV5YQ1eemVS
/T+kSShjt6ZH7NIXD9u1eal1hoYG4w8XbaVEtJCHG95oVjw2Kw8sMf8egH5iHEwXY7xVbCNBa+Mk
hOyeQkoF/6hKymXcXNRuojTdyYY2ySWookMpu5RXpyK9mNN6X2AyCWuI9kwoNXifw4uHHPX7264d
rLPi9Fp1Wx94H1m/iPeXhhxmnOznaQE5o38sVFwkUbStrnz6z8QguJ2uhxymnoeKErDgAkI6LOpr
zgAKZI2qiQyT7liK6BLRA6dg8ejygPmTlBCOnot38jdIALQMbakV+zr+APUy3slEQxx0SGdDZmoH
fY9+wTyh0uCBuclVzPtmFyz2MmNuBojrExDSFoEJ8ndAVbz1QBf69xSD90aDITUdRp0DqanktY+f
1It3l83Wir5098/K5kMykkPX0EtvR+BcIezXcPAYToAgvZMZxOkwiyndbXdwCycCxYiLwI9kgUpq
gzz3GdvSG1negnjin8FmDqX1k2aMhNUaygFKUkMjayMa5HdeMEhTDhSlkjB+X/LGa4BAiQy8S+cw
3MAZyQevDi6OFwtaqnMuGweOTlXltKnE+uZogxQp4BgpebTtOKPPje2ayklpFyuUW51LpinkUIj1
Zt9+jXnims9GbRYbHX2SYyCzFkGN6V1klr0p5JswwjooI3jXhGOEiH26nGjL2ZqCmx5TDf7LqtS3
VwkPxZat/MNFE24pVEZG0x4DwWQr5M3z3Zs7zN/6fudd10k5T7d5Erfiv56cFaWOoxwzuo62JnnC
7jcaRulimCM8qIPOoYAQjBYOYrKntK9BB/e4qsoE24gRKVDiyF3GkP7xFyxXe6a9hafOIjEpsx3B
9dsXBWvUCg38dLeB66aQHSLAIJGbj/kTX8nSVYqCbIZDhgaumtjP5wPmvmuIL+281dPMvZHPp1r0
8DHsNdU7FqgrxFfgLr+pKieQIuNqD7nmifHy/mVdURVzFpB8RMHylWrhPnGSWREU/qEVyQzHvqEK
MvlvGLmzN03IUn0Ys+H4gpVAh3J8aCJ2QHAbB9kjlZzdy40phkiwVB27eIXCYrFrFx4TBayot2nC
yXXo6rAFbRbCUGED6VQvEmNL0COoVFeYzPY0ISs4dJt6TNvoy0dSW2yEydn6X2j9nFdUANYYu/MS
URi3m1MMhDOtqR8wr1PQVMODzmtw491D8vSFzYcE9qLZFv5bl+9GRrZcT/+8GzRzaBVwkA7G+NW5
QRu3mak/SbP+3gxW3W8wmyzxZbkh4Sr8nMtQrY4ls8Qtr5CFChwZuhiltP0ooULdSnEaVD4BxZb1
0cC0i73ejfFzAMxxDGMuX2L2S5vpTOaL8+AoUBBQqB19kr+YGI1Cc2F9U9AbYly+Vc3VNOXP84zp
PLLSYSY0VaycNRQldlz21P6VERXpUnt5z1emZK1h5uVXILmx97P69Kk6Hy+t+jBxw/b3kRUCKEsA
1we/8IhSUJK+MZyYFvbcTkgby/yJtYjJStZWkgamcABkZroyWKBCrVaJ9QRuY5YII0jPYroDApN9
dJTlOWO9JnkliH9EUGVBk7aH0hd8T3fLwDOAjdx3xpapWIJ8icAsNiypjyTA00RT+QvLz2iQPZh4
XJYEHgxyGqDTRTVV9mA9I5/MCBG10vZUy0SNgokIna/CVs8VattvvvirA8xr/xui6csXwpGSkvua
wwRlba5ARHps8VKgxLDw7Yy/tEXGyvG/Ha6StSMfZDBFKiZD+ng1WdhS8k0nhlyL7UqCKTrA9AnF
Se757/Tmy410MqNXmABSWp0Wwe5n5LG8wxZ657lKVMlge6sC9W1Ql+b8mcpwuPYpJ14gvgR+76mE
kXAYuqt2s8FjlV3wwq45QbC0efjh+kX/hD9xvbUqPQ/BeCNCHVdiQN+KtRJ2oueZNdVjet5rwdk+
mBeHEWQ4jH8oxgur+6eRZaYJHS1CoNkwQH2vH5VzHgaEtkxC727G0wQEv4LAEchdMxTfFKlKyutg
DKxNoLQpzOK4g7MTPWaMw8vJSxQNIGditpkgtFqfP3coXG9wNSYiLPOqg/S4zO2zUHpzuQ0ZG06m
uj5j0zrU57pSK0x3K7y3X3bf/uGqFK3wfAIbT4N9z0J6DsJEADdS/5DdrNlBQsQBJARvJunceRjD
7N+yTAX+jZlt18af5FM42wHbnoMSm89SymbaQN5MQhd5lh9RvljkJj6OnrjGAiDNq5bavknqryu7
P2yv9pZHzRmu+V0vLWYCYqTjMbkjVqueOq8scKskE7qSHNVgbGG1YKQtPZ9LO/2sxiMYF7r+Hsww
Q5C0IjOOJ5Z1KTOjUNoQSiR5KsWcpyF8ve6R3ndxT3VzGL0pqarfbRu2K1WKHdCv+8r02sFxCGa7
dyrRA1SfHg/tTUb+yMMT/Ir9pdliSyZS1ncXc5EcNxAXCD5NWZV0Z//kPNa+LkhUg1CEF0cLzkhI
Kn453Ei+c0Mar0UyHOWGH3HAqVj1i1quLXRiS2xS6Bi9U1JZ+9gf9QE4I3IazN5axcug1v8+25xO
3Aqht09B3EfAF3nVhFH0qavooWiix0Zti0QHJQvkmFeQXnqEfPygd5INj+JmByfJQBor/60qo6g9
plHjN9YBz7xEal5HSnqbi329ftLep7wqq+P9uSJEr28wVUOXZN2mo+8MSUsyek00+imy95VrwQe9
0n5ACzW/RmCf7W1CAMlyzgvXZmv3+ygSZBhCWufdv0JUGT3Z5B9yYAV3h+B9QcFcyB3xSTilSjQV
Rc/K4z6jNb247kc4BPnWKgxI+G38gUrlVwSFqYGC4aj2TVTGbTmTtXofhf8t8+Vw/p+w3F4uOWRp
OaB03JoYS1DP20ODuEjoKh4gZxIWLiTfEYfa5XwdQ4z6k87ZO6vLI2zY4wQThQPKNUybaQ8uJtT3
FO206ypJqVniDLkqrYbsp6zsAVBwtwBgwmGMgkkoYCkUSUfQZGNmRIICW6Yr7VoX2A0RFCPAlm3d
/lGmXR97G0eST6woSUxfagXwHbocNW16UEleb+jBH4CuX1ri1AtYOwcGWqDoNtD3Pm0xI6M7CMO5
BP5EjbTDdov+VQbLmpHMjpabdb8u7NlscfZs1bTliZNNGouIE0u0U5RUmaqJpc95XLD6OfloREXN
iy3/kQIIt+uG7AUX+/89kBdb59C1uawbH0Tg+FSk57DjiTNh1NgvRrsH6rzXWJjVxn49L5+2ONZc
y957VhlU5aobJlRMtcFzehF+hHoO/U5puG80yB1Dvy7usuqVBcPMu5SHCXvO6AYH9+NmFFlmHvRA
1UNAUh9t07ZmbJwb8n1Jw0gXvtf+Nxg/Rv2vHemOxKPv3iDOS4IW+R6KMIFRSzdLSQrXCudCknxu
qCLROdVsS6tZNTcXuFHssufuRMdxjVJ5fBMo4Pw4LLhpSI2mR84ADhcqnm8U5Fz9oQFkJOOK9g6c
vQWrx5iGrHPeeoXXE7oRzD8IyD4oZD/fx4fYKsjnSPorT00IZMMivmd/VccdNT8+ktWbBEE/DhjD
zxUDMen6MbaVk07fsMLl6qTn5GAtx8Bg45UVzfdRpAcJwiecnGOzrZxiK4vthQeK64fa6gbprKeX
rLKiL6+XpfSeIerFYwG9CJhRbc5L7UqBNjufqQrKMGVXJSyapKpARIRxjq4o+vvYdONHCfw/7yRr
cDwdGIXbW6vlMgjEyBMLmTjR0M23ls70I2W3hGxHwjlJo7uwqxuvj9E+fH0F7aNzWP75L86jg9B9
bHSwwL6FHv9Y0TY7kTIrtxTLbpGikst00hsDsaWp6x7uDz2ZtTCPAL2flXPr+6cXKOEDBgNUmIjR
YqBGdnBRt5qg2vK4O/JKyB0bMH2UyaG3LEie//sgDHXVS5qo6JQuXDhgAMQlPYRrSsxkMJK1sZJ5
pNknwDVFX0rzk2qhMr6XVBEDmGBFQuZUcamqujohkG1bMu+n/8ge4D/IWgByuQof9F2NdCAzrAUA
fc/SvHVd/xBMV9dAxaJUQ7RHlczO/88n6ZCNVVZkDraK3fihghd+EoLqDEsP2TQFZAJ1vwozIPXd
HCv1QBwHkjmxjoNNnpiNOf7O3s1KQCuKZpuzoz5PcMhrOHPJ0Kr6EhNvgklK1Dd3c6GRlVN96TR2
Pt401r3pIbT+xyQ66HV8DXPB6k7VKXwROjBB/NoUS1nQPbdUDPRALwGbJChCNtkXm6ExcmtgNxa9
DYvdedY+AeRI24QdqTni/U/kKn+p5uoB/Pyhent7BoVi2vJktRVmYKS7NJ+LtvisZJeIgahV6nSP
hej36YivXHn05AqY1NmdkWF5dveKNgwxC7AG7wRsth9HB+a3SJLOn2KB5liWkbtbJ/uL3kZNOR+x
8nfDgdUQDNYU/79EZMFX6eKWyS3JSOeue5UHI3+7B92SBVQ36gvVuPg+GocA8sOBLRn4iyg815Gh
i4qqQuSnu9kpa/5jOzK8hge7qekVw80yJFVsAVF+urSu6UMYAZAMt29JQLZKzUekAn6+/ZgyX2Z6
0GQ9l7n1yrZqnh2n0aZJA8xmr4ZGIHkpgzAFo5s9cCmyBuuTxKmOAWB/OC3se+aAZgaAO1W7UwvW
FLDPsH5A8PJDnfkHtpck5ZOkOYl76xEXZat/ioJkbO8fKcVO3q1p225fj2z7vAsLwTyyJlbfMryg
/LwqgALbPizn6Xr6LXqrdQbXFUbjuAxOm5v/Afggj3+hriN8lMFv8TcT5YELUsFOnyYZsx9+ODbT
KH4f9JRhk9QFj0oySXUgA0QLYksWtL4DGShtvn7KaTmxSSyjOLITE41Z6U646rmkD2pNzci1P6XZ
i83FQ2DORgWduVgTkyEMlIaUbvyn+7JaTZt+gRXEGy79yCqMSrtc7j3V+hrAeveRkK7xIfi1zAPB
0kGB6do4DAV9jPrI8HH38kiJvNFjxa7N4x9lQAfw3uMQT/vEzBlyb6sBgNsiDMRWLxtabY8V+Eq0
fGFKZOZnP0v1UVD0p4+RkyOLIhMvKiYUUSed+O5W3+HOgukd/TYzLHAsQDy5TWpTnaWujShDA0FL
zrhmdKsSaKUU0i1P4bz87WZyDkFIXQqHtwTNyzIwTiNNqN52T+gRxfEjvvGqaUUHZZlcZ5YrzFcz
f0bGH2T6FjFuNgrfGj3oqnt5iB9Kf/KvWdFkkfzOTeB1rIYpXE4NMmwVC6mvh8VXZRMNR/b3QWb8
FvEA5UvnW0JdONmlPlL3yfQdMM/S4iRmN13/IGTmvzfT/sPWHdclm65xpbqfAsF6x4HZKFjikNLh
IC+nrAAEMqtyy6tY363MOo5SOJcVXftVgzqi8w5ECtwfe7ttpi+gUcp303goGYnt7TGjkI6XQR3X
RT5/b0VjYxZsjk6DQmR99XnKM1tfYU633V32jKtVIGTB8GjMGHqqHvw9saR9C4/rOiV3hE7uvi4P
Eg+kohWLnUBXXhYLDVFRYbsfrxqxHV88grFhhD1tR4gT4nOFj3kHK3oX6uPeLXOdUbTxN93RcRMk
XLgyWp87E3jA1wfAUksmCPUcI02iPbA3VwzptVWXIybYiZL/16ZP6HtDa3V+XMigheoVGyMyWo+C
8KpKmIVknHc9uXUF9+/UIoC6z20aSGanaKwt7qfZxFZyPN088EgoPXRLDHVHy4jSUp5goL0IvyWd
HMaIc5XhG6kggjBghBQqRCWUfQGfX/eqU5TqZH7RmvP3cfoq2dt1FGmnYLkRXk/Kt8wuYM1MoTFG
I+a6GcOBkz7BsTIiXPEd5KSZpd+BNu0UpNpEg6bafaAcfb2onuXF4DBH8yKEGTRsiAp8gxZ/kZfF
DZB7mRZnhDYPyhF2hgoBCthU+Ns72u7Eq6ZKccEW6gH6Os9cwaibOYjYet62C3TO4NDuq1j5qXIG
VN5ufRNfXZfJl9IrAJ3YeArlKV1+HXLzcgkTOtnUxUkTgQbu1CwuEvXKPcBuyAyFncK68kc0P668
rci8vANhYz1KOlgwaxgfrphuXTetjVvL8pNB0GCoEXBhV8YZ9XETQftH4CUMVOFht/MOGHdfvlY1
U4awi70PknapBUYZzdZEdSeGhgObKbnQe+VZOl0vpL28985h2a7h3I0ZznR6c/vmDaGAOyqltiJe
rDaZ+AXXvgx+/uXv2suu8kcvzX/zoDob1tzAwfay9xLHBF18a8rypJzNjqf+TSLn7xphowIXXico
8H+CXSnlos7ZBoZ/RlkNGu4XtpMelIaVETXmhyeRbd8s9jZ+MUbKnaqH419Ws3QN4ZDOKVMyUMYE
YU2EqlPjlAne/Wai//ppfXk6+u8x6oX1LxcbveBtU3kVtEop/sfv3O0RJUt/tqUORuyVeUjx0tW0
e26/uZ3M+6vXmY4X7ArUK/PbqhC6t5xIDVnvxacDU7yEHFEgM69lTGHWpDNLQKnFaAIc+Fgu3fXJ
tS5HtGv0lvTCOXelddNpqLjx0w4mQKiRmMekbjb5BB1F1Kgnr/VNFZYDvri/gpg3scdDbQ==

`pragma protect end_protected
////////////////////////////////////////////////////////////////////////////////////////////////////////////


`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-1", key_method="rsa"
`pragma protect key_block
owhyHhj9UjF8lNunSUQOJ8mkD5a6djknvtmibnIE+VhIWQVHagHzUHo/BMNKP4ftN+YTajf38k7e
mbto/oI0mG+3dLWdkv2bvRrEWs0b4ffqwnRyzcKC9Vwfm4Ja68zPHZ4YkqbNdb5HbsP7ihp6BQkk
c7kO/cFOM3vbMDnvtrQ=

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Synopsys", key_keyname="SNPS-VCS-RSA-1", key_method="rsa"
`pragma protect key_block
Z5hhG1D+FLEiA0fbWVg6WkVMLnMQdT4xdwkEJvK6ufaDebOgXPBgWtwsQjiYWq015j2+j14p/kUV
ZM3uhdiwv9n3ab+NdARFere2uoEzAR7SbShgjMVzP8RnYlhenLWVzDUs5k8DpMvSmajYj+NP+Vil
kMZkYEZkDvv1wlLmhS4=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=1952)
`pragma protect data_block
NSqhYI6n07AD2h/38LPwsHZ8Na7kb9XfLzn91Orng7Vjxr5wp52pv2HoEwnopr53HaNipInwDjLD
cUFWT+iMk9FXn9MxPQDq/Oqtu5WnCF9ZwZH2gsk6r/kaxXWDV+1SuSGsd8A+AbpqqO6offf1KFMl
PXt4MJw3mVnX0W8t29NSMJlfhndnkcS/vd4d9key9WtDNIxET1AQewK4+s3X6fsLwnbSbKM0nUj0
HpCsbU33kDoiz7Srn1NWPOPSiojTbbH6T99ip4eF4F0vTnwWu56FfrunsTNL95xe1fJdtlpjmuBo
4YTTt9XP+tIliVr7jPgkIpa674/H+cuimuIuVss+y1P53LTARqkLZXV+iyNsy/JRBFI1X47yi3Jy
SIUfaIGLqPubdod4O0crzp+5q1j5NFFaWgp9HF0Qxu0+Bkq6T9AjvykFqSIvR2vPgEFHsAFzAIoP
GO3NXAY4JwNZMD45DQeK53JmKcWXzLmVu4kgs539WthdOKVOod0z+8JU9dviDEfuWvg2qZLzz02x
sR14VhLyClJ+wpcPuJvhs7AzSniPS3BQGVhpGQeMqTOIYVXmR6kRV7CLaqiJSWLtsDdDja89Bvla
N0Tc0R7pFtZmHXYGRJsoww48EfP66078UOymLNlRZ/BXVhXj8xFnCuWiK1tolfD8Y+YmPqXD/occ
yUo+aJOU47Tuz7vnNvJsrSNOIU7my90V6vyOvoww2u8UKq2I3/n2gP8mpy9w1si2PzAfHskS2snC
ednzYfJu+oHyOAh8ZVOGw8ZtQElqV5mGCn1NfPg/l2GIwcfIIz/09MPF8M9pUTHBAa/Q7Avk0CGp
zF4KYvkRwpxfv9NF4a9rdSZKxbYU+TdcyniOWs2ekEQVZ7G39RAg0EYOuXQ5ipQUiT3pOFkYX5Ep
mDxawk1R19Xa+miJ0xrrRTZchYXvoOxzTYt7FkuVZJBzoBLz2vIkwW9eHF69oBYTVJFcxYR1XPUd
2/WhXBYHnonTiiCaSlkz9i4w62c/hfqzhnqPBXbT1UlYqBQzx3LVgP8ertsRkWAzwpGhhXvfE2ZP
bk7H0l+3+vw4AZaC6x+R7no5P7+oQ1jvJmWhM7tVBNhhFVrRFPJhBs8jo8CRSA2tY15MAzBHU8YQ
RtEwKiHUriHjUHS+dJU7wxYHVim6z/Fhx2GbqSTyMx2vRvTljMDtCqVbA4AzvOm1qtq9PbMWBRL9
XNZiI0PpGeGPBB+ZjJb2hwBm9V/ZYk4jvTbmoey/jwEWPerjvyrp1Cz/u3yJI1aHUOT41F+UFohw
SPppoUKwiYF+//WMwQTjO43ptB0JkyH2c4xc7cxBuoMiPONxwrHb0vPi2dPXnTYiEJr9+bqJXOb5
XSDnVX5QL8go63sJzRambqkgUpjDe1OkVksx0AmAU1IvkS0xmqsfWzRBLxUvS+RE010D03TjUJvs
Hea8GGEJiorIJPoLqihlZ+zmmt0nFYyRLcdiwKX/BOEufvjRNIrqFXssHQ1l+yzRnVIDyNK4WeEC
7OOYmQvD05SSClk3STjFJgzw0k6UnOVuQxe8xrWb7cXNAyEC88VrvHokmp/TAB6rMNv1mBgAuza2
ZmeReAajjxG0Z2cNpL6hRUYOoap7Q7mfYf0vg7t7BbQnxKcHwi636Bof0FFf29IVb1zA/ys2NQtG
YgByCljLqMh5dfFri/T9HTXOjxvoMkDwSFQk9/Pyni4CAH7hz/lxV5oyLJnCgA9A/3uWXYegZ4eF
0WkG69dw1CR4zLGc2GY5l0jB2bjGMRecRPXm2ZuWI6IW+vzYq9G+TxEuRJABIoRCRnONvmMadd0s
7kjY0LL9uzZqw8Crw5ZrO0PikQ8U9YnX5QBJZ2EiscYWGjMDbs4n4nwJ9HVLzQglHgfaPcPn5puX
AwCttKZ/zXfrjdBhu7Xw4ntOWmzdPi1rSak7VyTutNfq/WUgoGeUiUIL4GukYMYj2T8sqAOWVmX9
mC+Fn79dE4a5q2gIYfjxJQTUKIgwaBoxPTMqXldiFW+TpzUI9YgPPWatIp46WSykb2il3A16mxx9
V1Qmpxd/DYCADko0MU4PNAVkU7KiRdmQ4XDkUNk1Hr1mztB4kUGtKo1xnIZiAhcrpb/jcrY/Ll5I
GXiM5u8kf9QsgUjMfazFKBb7LQkVKvwiMK68r57rlU95rmuMDqS0kpgPn7ZdDExzXbArKohd9ZtZ
Ws0olpMgV9AxqkJ0c3nmNHPMUQ766ztUuRxQlRDgZV3qMvxAdQVcuJ5XQOfG0goFVL557gmI3axS
sBDSwmaQ7xUrTDYrRcZU3+oLBjGxgI6GzdrgGMXcOBzud2BuGW2PxiVVm3ZmS5ugDNbCfA2jhX9l
LP0iRnqrliUHQgEno01z4J8z+J9Ejtj9EKMKcaytw+XUqNv++9w94+MxBZiprvYbWpeeoMTqXxxG
JIDgPOsE20KRZxIT34u5tcUeB463dIarHrTbAMpwbL87gD2p5XcEE9LkLHyUaMzgFS+EwhNeZTEb
gHROnhPpO9KVq+HsatZSgNk0jy7OBKkuMQnPKyRjf+Vur2Y4LsSTDOKX/si8lPLeU96sV0XfYqSH
45GPZX9SG8D/b12RIbw=

`pragma protect end_protected
////////////////////////////////////////////////////////////////////////////////////////////////////////////


`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-1", key_method="rsa"
`pragma protect key_block
JxHN0T5s+0/BKaJDjHicLw//nI98Y+AcG3uHeH2YdS6CKOH9l39AKONUUyUyEPskoRF9KplgBtoy
SAaNz+5A6JUC6rdp0v78vLQ3aSNZ8SN/wwY3t6K2GtW5RH98UPvUSTzsD5LP9q0QQJT8q8XQZrrK
WQcCFmv3CEAXy9kcacU=

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Synopsys", key_keyname="SNPS-VCS-RSA-1", key_method="rsa"
`pragma protect key_block
jI8RYE96InG0tqLdvHxG+vIo7EuCy0I+UklUhxgmdsr/x+ANOdc4lSggaUcZSBqfFjriAb4Td/rk
Y5NQUIAq9iobdLs/W7S0r2RFcVKixxjbu9uZlv+fHBxmBtUIEiU2LK++PcxjEA0ackXdp4NHQ1YW
Bkz5h64ELxwX26B+aOQ=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=3968)
`pragma protect data_block
Za9Rx2udmcT1S0BjReYHl6HB8z5YVp3z1TvbAraxQdwGWr7IgjHXWAm5SzkuLf63QRlpcyt7Kw3y
sIHSEWPIzHv7N3wFilza6gOJQnTf4AO1SLL36xxPzxcUV8z5w7WPayftVig83j+ki+aJKMMORAiB
T3D3d4Tbj8XSiQ83sKm1asX387dsx1tWSzupZlOFM3WD3eGv+bQCneOyTcNX9BQeAOXNgS2s6NOJ
DASeHbdZ74CWLInTF0KL9M7Cy0Ls3ewjhNvya5bfarANl7Oc6htpn3gY9HbnQ0WC+Z4m4mQks0iq
4MH77akWgt0gGoj53IN8h+ZkZNS5CTZulx72v1XkvBsuXnIuSmwqSOLiaxu8XrcSZmWHpR/5DX4V
1+2PqwDcoUtEP5Gaw9fogTQp7hL5jYX3Ykps33zJK/W+r43kpiyHNiAIDTVVucgOwCF0pc2x4Edb
rOW457ldDY4P911d+P36pEgQuTYtdpxGNw6cOkGXLJnAwxARiZ5TLJPCHDIfOfipyGkYtvc+TZiy
84Fa9og+ZLsLbCYffFfby8kF0GH0vgThcI0Jz83Q8FJOA5SAThwtzVnLIUO0xLCttQfvePEQ2Wik
8MxWxcb7D5naSAGe53tcVrySiVSLX5JZ5ybCz0uaYcpYhEieKHsUs8G3A6iQJVRvicQKjRHBCpky
Ubju2QiCbJvNS9qBdDnV6fw6HCnxqcC0CZzQPc21TJz/0fCrk0+YwzNwrjqTGF6bHy1+XIUo5AQ5
GTFbg82/wy+jnpRITn86VJdPER3nPRZNV0m/vHPF2nP5oOJSlDYXxoYkYm6rTCyr33QEfps4ehsh
OL6CWf2JvKkV/M73ABX+HKsXm3Pgy8RpteeLMs+avRzFx+YyoG3CDilFDuue8f99N23JN+CoYHAQ
grZkAZRxSswm/IMDlqCuq5ZV48TKP0QN6ZDW8VVMC0yq4oPHNvmNxNsMOW3ul1z7Wfh0IumGmpU2
206c8f06rFYs8cE6dNgvGjdXhiY2Z+wX6r6HNK8jPKoTDIPVEFx8y/PoRhXCmD+EXu/UK/BjKUmv
JWCVaoezv/Gx3bslsYenUARRpt1LPyXiu5trYRKA3tqB00Aa5cbYE8DpGBKwKm5a0UBF3hgDCBSt
RMlMyjbhmsuJjgbvZmukFQYETuB8T427Jb52m9KZugAMRPTCgp2XwLeOoP20pq0f4JfbHrIsGD5r
az/sh0nkny5/2iJIFxVht4gnk7OZmz6yncsgHQnrLJ8aI5HLBfCG2uD/KQmpqLObricxZVusf3rD
esSJv0iYN7BTk6upDqyVkgq7cwq2QSP9i9wmVBwBftOHkNiQkP0eHuKgAXuiLdxUVJ3jUTZJ1m67
kIPWYoFpf6rhTNNn+cqsjenG3CsWhn9tldebCfCB3nG5bNXCRTvo2uJvhf05Wie/68nqD0UJr6Ox
LSq8Odb7wbKb5IhRq8DoDOEgDGs2ZrTbGn77g4XaCECnHfHH9puck7wRi7OV+530Y+6t01R32um1
iA5dmqD9FwY6NEf3Jp8JoEQG1rM38y6TD37bG65TLZvR+2kRy3vxNmFkgd3OpowIibdOdMZTXapk
rUGe9JcIQGSPP//xGAQTp4gcVgj0HcLxCGZypM6ZMc8t5IF6gvuiJ1C1A5dpgej6gH+5R83gVdiT
ZLyiOWMjMDU1OypqulkzDuLkzOKbfAdKa/QzrswvSiTvboCleDeu84rKlgm2zn9K2hPbBX268DtM
nIcHYZMddxR1u62R1d1bRZ99c4kK3AsRSCD91LF8JnkLkI8nMDTh6tJ9rxLbOJ3QQaFzpQ8DrQYb
KycfiPh6g4//RjpBwhaMxC/1HbFEjUAmz4RbdPu36L/L43Dfjp/vc/DWWjTFHx+E1QcO4NOly69C
URReCirCYmQgl0S7bFbqrpCSL0+NlarH0FkbLo9OguXQ3tVzZxqw/5n8xraEJYpZeew0kaQ/RFqz
Iyv4umtsJkhD3xc4W4kCj3mzxyhXGmTDK6Tg/0kCPJEgkhPIb+r1olt/YvHoSwKFMftu6+daDeMF
Hoktn0CNyJ/W37yD3O3qU61LSuo5ZZgZ+13mW3hTg+QcYVDcKNqQpE2B/iOYaQ3zkQE07XAztedD
2Ch7NwCvpF2EHTovaeaiLYFkPbYTNJRtwc8n1s84iOg1+pwu/i6+yUAxikcAh86tFm9NWDeZCyzH
BWk5X0xlueAyJgHwftFSV9l2H/ChWbHF1l6gU7dyyCg0bgZskZw9YV4rEFw4ifTloCmjUzZeax9N
hh3QzdhAgr6GvWawvu8Wrb5pOO1JFnOyn0l+/qVNHlWCCDzEdOtCZtOFE2BhbcAXuAypN3g7FboH
Ry30KAdmtW97JLWsMPhBFX/w0YlI/+1IDDHABs8xrzDFTLMjci/ZOC6VYF7ZaIsFkf86q6/CafjI
3WAnWdh3kcS23LdilLecBUyfa+3+Eu1Ds93UdLDL1TvIzjQo9Yojf4t2a29HH7y3UMAWShwF9v83
1aEHF4bY+YZfLhleT/4r/GrW0CXmC5izrsdQPQz0SStQArYHsFfJQ0xopO1WovFkIjOw6IRHBDjc
rRb5pwhtXPq1UkIN1z/5Dzb2GQJZluzRDBwAKIXPOlf1R7FVw7wQKWNp9hKBLwzPDVOKPB86jiVC
BJ3wyybZ1LW6TU4QT7/Akpu9pGNAWZ5/laNot4Ko6sJtH+/zl5A8Tqs9M9emcGkUFqpR1+xZTNCZ
KmVxq1+Klnxif4+tFyn5C7LRE4vkZyA8JidBHW+JymfciBMvountK6RxZktO1mI+ta+oUMcP/x/C
uueGc9Rqseb7LmI3ya+hB8F4E6UOxRQxh3CsbfoC4uH6gJPv+3hAVyE3sSuZFhrN2mz2m0++r0xG
i9GlTyG2vYrtoPpqnSGS/lvg4XdUoQkEYIvex9Mb7P5t3U7IZqOIZGR+E4nD1tTZcC6xE8Ev07gF
nEJsXgiCLYam8NToVUYf7Rp5UINuqmewPa13qgPGySYS3/1pV893IdHVdLtzktFmXNEhxU++d7Bb
Unmbp6lK0rlQxQjsuqyQ/hJQkLi05G5MKlTbxoXcBf7re8yn/RLr1PyahCEuDHSXW0dbfTV9mmBM
wFYQj4z4cLnOVotqzshZIeuQfxXAwmufwzPMS3opH+QRazuTFiI9BOKbBPIfFzOgV4bnQZ+uK5KE
WVcGAAB87W0d/lXWAx/qy9j0qVhk5jZ1+ccHXz7Iv1JBmY6ykyX6EvPD1Z3QwiIaDtwre6efIVP4
yM/80QN9P7sAKfGd6BcX4zZ6fpFG29NMp77fvH35y72P4grEnVY1kLkkf3pRi59RMoRI3WOAnMCq
uGGQjORrRpEzQr9wtRNb/ko2ByQ5dTtCxBKHUxXIlrY6UTYQiyDLUKNDtkFvXW5C45lCJKkwbM0+
yfZkrbJ68VEQUJPCeQu+eBG18Q8+DHslQz7IYpmEFu67BUwdQ9g0Y6grPFPAF25cIgWW1xw6onCe
EzQJ7k9+QDxS+X+lB6Oi+rIxEF4fro7ZxAWjoiHEN4xC+6VMWmjQQpl970FqQ4jNr+FAcEGJrinX
OWI1zYK4olLWJAKuryAW3D1tMdPGhXDu7UtES5zIZjUV3a8w/zcoiffqNC7lYMFEANHmAx+sAaPk
9LzkEeps+GjC3+nonZFFAXOWhA3vcL4Iy6IZHDTCiBEOqglKRpOp1tAztFnJpFExOQeDZuoXnZ/N
Tc4sjIfrB02c1PFBuWqOAkgQkYQ61vF6mHQALsn21c8DYFIPBlXM32LIqbajXowcEa9B36hLEiIm
mIK9yugMk7UcIv7S+pbUm1Wmd39cPgt/pvO/A/MQ2RZoeyDcbxzWmv2l5aR1S0Anx+jmnu2sbVCy
wefzFYK+xBoV81vOsaoPkd4rQfigWVM5BfgTEy42V9BLs07N9YKDRtecZ0r2JkI2XSuUwaSmnkeR
kYXndB6Qhys+XLLRDy15O6hvVslHz5qNs4BoMpbh4Qn/yP4QOqEhMxyYCaNi9MWZaOglXa3trnfW
SXR3261jvrcOBKCOIDyKusPNfSDllidPFp+hMp0rDtc9fSPn9PCTYpwOoIra9yLlCKByfM7qswTh
QS0/fAvZ5s3y+cE/eZnzJqjaAdSvbW7nl+MuO5seZV9ykG1ApqF7zkc+hb5X9gXiFyWSGbGwkEd0
6Aw8XA8WtTJs5j1zTovATnnkjsVAIAj7UKQVSApKgzIOOwz0PKLzAa7ngx0pd6FIIS7s6+Ah4yYz
pUXKc8sCUbkU8Utc/wo7fKEOwvh92IJSCH/HRPVyMFcLFafedMxOH0cIqa44vCegzr8sg3hT2Jgu
Kna2PR1KFDv3pA+Zzxgvfb8OEJlpDJLEw7NYIMXNVsFI+aLrel9avnA0ahvQGn8KT/4r+bi93Jt4
bcYKgcx5Nl/RzK9I/YdvH2RNHm/Yw4qCzYMblLYErd2883YkccCA4cFvNlxMmEka/YlfAx9vQVhS
LCKOrmGt3LwIP9+IeK4EIqsWScNES/A2B0lMP92+NfueFkaujPkX62rl9JOBSKQm8AfG7+FutLXa
C2XXUPOBeEEfKD904v46mKA/i8/boaROMKjzeA4dyRch6gupyFybWA/cPJpA3pMiq7o+P7iewAcM
4YqBP5lGdYLxr8Ojwrpc9p8/QWpURxsC0iDPI8716HP62OelRxBflvBT/aVFiidmwjkz7k7Ao913
+dfBZqDlSEk+fO20567EQ2AiXHY8rC3+q/nuvd/g44Wgef3czWdjDbTGwxrz5GJluHvw2F9jcQSS
ov4egJV36RrhVbwyb1Cd4KrEKAUEFGTIvknZgxTzlIlLjGC6MfTHbLPzSvV+sX99MRr5CGMlWnDR
9HUE8+imLTEv1ApLE+j+YBZZLZYMAtBasKHvH3wD7W/Guk170g3Pw/f48G/gVk4E6DxoLCpbbWsc
tIeYXBNcDAe5cxOgXTE9njauLO6PHWXf2+dzmS9q30By1yB5M+P8KrK0vk3/0rHzzaBbaoQMeWp0
FkqdGncfLp+zrgaEq71ac9FOQah9v83d7VuYXXggu9Z8oBDWB2IohP5PdDkBeIfpuyGqS0d3zhij
SmkKQMMQcexnaHbxiGJkss/49Hfy+vV36KuJnBe9GQ9bRiyVwNUi4ZvoE1stDoLXDydtCvfFlH//
0wJMI1NkXC3vzaAx/c94RudCHtc912wT/MDQJPgY4YnhMwuBWBvqNtoe7B9vbEx01hHntMZkxOQm
CBa+SNfrxrkzpKdDDKbegav4FjBeJA0zL06UcsAxrSeSUTk=

`pragma protect end_protected
////////////////////////////////////////////////////////////////////////////////////////////////////////////


`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-1", key_method="rsa"
`pragma protect key_block
AcTcXnssstMoR5NRd47KJt+DGCTTjHqu9UEpcwvBw21RdesJBDTInROqJrlETbDz+fk9/sfYc5sz
es8alTGKzL4C1LjbVSMlwCyd4ZR2uCNZ8c80C6X6uP+E9TJQ7TvOON1BY5mgw3oC4/qVHsrNhKR7
MzJNGHY6LHESpxwK5ds=

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Synopsys", key_keyname="SNPS-VCS-RSA-1", key_method="rsa"
`pragma protect key_block
lp0pepvv9xL6KbrFKBm/zEoHOQFzj4TreHr0xq4ZJ0pQtcs/JRb1CSVTtLcyqfiLBdGvFo6o6FnL
dPK/BEGDUb6c6FZm297xSXeqXt3YiNrq3i66JLnW+zhtGRtHhPKosNq1YqTyIQZ4rFneTikxMvGb
7SSEb0/0QDL+VDbJdME=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=11024)
`pragma protect data_block
ag4WdKEynI2kXlkARzbVA92QUM8MQvY0wjYcd6j4Bo18ysviOCBvNE8fQ/jw2RTEgvfFDzTZQkmx
u4qhGgpr2KxGcY10AS2qyKMThKWKBpbBGOLLAvVH0SwxpOF2F5bu3wcrTfd2SbSmF5URdkKRr45Z
q+Chv44sEYi9PLV1KjfMstxqWSoVD9OAIJiwLfKvSF6biOJiZ0tXgLLqBQgVahtdrIpDmcPPR4KU
eXdRKPiG8xMbT+oomT3/NoERDKl8ROBoobEGIeRbzm8GysT7axzE/HTJQkR/c+CO5g0k8m3vobLH
YwBowAHZpF3RXb9oAB4yKoxZ4XENY3MJVQFI8zfu2iTD0I0ZagRlqD3w4k4blhbBtvam1ri4M3gQ
s4zcmxCw1mGK9prat+VQ7gffv1Qx5JhM9/tOW20jGMnq8MH6lDvPGUrhZwUajZge/LHJKL5gwhM9
1cDtdrah3Akr1C9oy9MZCrzxkOphi12QSNW+T79s5mFtt9nsUXShteFdneuAE7WR5mFXIq4OTHw3
/PdPNz5+ZU3svYGu/7giqaBa2Jt4ZV2ELUpgyNBhkx9esi8UDQSvuYnW4/RCoqd1gQ8W2PpYKcpb
nxU4OV3lddfiEgRQEKXboBIPXqqmoImGz6meGkKxDRqJ8Lt4kTnVUqYPoY87gFalk530p+kSp1SY
N+ZH58XIXLB+xKCUXykB4rj2ooXwL4GJN5x840G9xFIVXaoxd7MzlUsw9ozzgRpfREhwPGcDt3Vp
+4SyL247zGBWcnXDjBYKTZWvmD+ulWsz0rPAhDnKWY4PgxmdNUWtd61Fb+PtYJ+16dcWthDrqFl2
uX2btIkMRhPG7Oq4Yunzuu/j2aMczubVMRB6b+6irpftlLV2xLRhnurcXpZcrVQU+VORL9VMI7ZA
2Rdr+x0sBbf0R0bTuIxlqIZGd7NGR8Vyov2eHV8hbLM6v71P6pXHqVvXSFdxQp45XpjXp3e6eBJT
rbg5wExVoapaGi/ZNtxGpodHBf1+hnwd8qjQ05r1CuAgGwwV2SaNAASHYms+7JYLJ7v6rH/8cqrf
xWQhGsU0F7Hi0Z2vaEt+9724sfxQhNxZ50mEzv5WGebp87zy1pWmEJj1ygROXbtlk066/vTMNWMH
XkiZN4AQ00onK3KOhs4ExSq0iTCxBmBQOAivVZJvpnsb3SZGsB5rECL6IGuILQFQX0deAYBU3npa
CF9yP9sD/4eCuHR5lhM2IL8AJFaCi8zgN4KoxZc+FwzSc9CJ736Pd2HwZxxBzbcyDpfuCIM+wBXv
A3Rwg9JYKCiWNo3k4jFhM+boSJRCiJDh7Pa2Cj2Ela/i41XoDVw+1dC+0xGrtcOaUnwEFJ77LJuo
j5FcXRI9f3SRKdBbaAMohR/Q8Awvq4+M6AcR3LGogXLWLM+zQsL+zduRQmOnNRvJCU1Rvf6M1KVH
KYWrJ0B8142KdZzsUGSeixCmMXnOzMNjm/WPvjq/vvTMHRIRSjqXbkaXc8fzSGmmJIy7iphpkYrw
qWBhYg1Co4/479wQdR9HPt4zS6xYkZsCcre4RjXK3HYeFHJJPFa+3gUeSKW3ahdlijKyctI7cFNU
vNthOF/w30293wHHSvh+yLBQzw7f6UKHQJhOkyBfkID7luBIvpVHWxdo1wlLF5Iz9dZSQzRJ6BRu
RcH/z1KN3dIQAowol0o4W5Wf8/g8Bkw0tsHBb6tjuY29E8IPkwfdoJkM9uoP1OLmnFhJ4ExHDCdT
6SlHJu2kLuzErglRNSdxS7/Ls+XFTvinWn+SgtKk4XFCRUdD44QxbXtM87HWtdOukC4OkPmCtIt4
Y2RrIETxfGKF6oFfF9w7LQ3pukP+/vzMXd9qhkEQrZQ5FuQhRV/4Otc5U03K1zIgoo+YDQyo+2pD
51W6uvOz9qSh9Y1TjCnkV2U4loYUXb2YCfoinLN17aPbjnE/ajFkfOaflEZJ+IrXXdljeQ07AtOf
CzO1MgtSOKChXWGVPvIb0pEKyk7JZV8pfwqw7Dg9TMgJQl061HVmTvDSwfrZguQPr5sD5uQt/hwe
FcbAIY4+RRtjm1Q8R46roSe4gX5JfhsXzmI+cb8gSgf15QXz609m7KoOB3+tFQi2s9ZsHdmNyY1X
PIaL5ISzaIg3yjzENNg29ikcN/wMXFlFuswYdR4UUZVlSz/FfKHZsQmiTeBsRJzE7HXH0adZkgMQ
I+ptmz6avj3JiRrAeK/zXsxUNZ407XlHp8DM0RymZ/o/7vNARmqg3uUltj51fve4ubE1GaNFS5Z9
Ltyr+OSoJGa6oCprDl12ipudwduKaURx/8rB7jX1tqx/N2043gja7IUhRJGqSXq9yXrsqHQ94tXV
Or/TpwSyTFWCen0aHxxUqUiYGQjHiqoFlr6juelFuio8WUKencOLi3ugXOXtRdYFQU0b/7SalQLq
m9QRxontr2zslyMjAr8n5+FuJVua9M7cl4Wk+GSrQfZkzeqyZvgg/6YpxJ2Xn18sqlJfLuGEHO5m
JN7BzS4hg69fB9meyWi+/UqiIRTV4jxPQhDmaaNkZTxZcabYxlw/9RuCx9MPCULQDguL75NYRO87
5N4uF8aZYeZj47iZzFKYEtrYWF8nf5qf+xEV4fV/DBzHhpyPGk6oEYdy3cixz0nH1MmsXOTYUq8L
yCLjKqff4B40iLS56LK9kFnzYczIeVfpmrQWESI/5rQoKA7GZRVsfuaAlMTtNnN96+Z90EPBmCE5
/JlA9xlGaa3EAHKgkDk8zbLxDCY4Ql4IQnIocnYXbFvUTaqBjvzkTFH1nQgL8l4N3mK+/VUuHv3F
P2ccYmNOkem71083U0NuynTJE0JCMCNGM4HZHxxnOpdocwrWsFaLoABMyOyGxxUhahAI5DAsjDEa
H74Hpgms9UPQW9Vvwnl9nnLP5EuvSgqE4ZcgZI9pwwEy2Ut06Ohp5EJLejBPIdPbkOTA9aUxz+OL
2Za3tVwuPW5+ok1amC+fozAcbOSLPJ31tdaVQoi3D43o6ozT9tXvF3O1Jsm5K6/H/ewPSoGs8T3D
utkaTbXmpR7uqzNIbptnv2wAMZcnmWHYcdtjSdLZ11EZL0lSG4lfudhuP5Sif42CIGSBKusDrJhW
VvzwswJVCBLfia6DwQocTD+MSlHFBybqXOX1hRnLHZ37I6g85EOzo0n6oEW0Li6FkCXtI6NEEpAN
QjGAOgRRUuL5fIj+jFPDcjw82CJ6+0/k7V/bZncdFofo5ta9HBAN2BIum3/PQT4QYD22y5b+FIP4
bva6owJ4FywLFOLIhXThgidzpOh9lAPvqJjxT+mpg5nOW6RvcxDQWpMCE2PsM8yD59eJnVFFJsiY
m/9X0Avx0Gja2KagKrVHSRdRbWrhR59B0bSKIvJJ0dEzhA0n54wBEdnC8/KavDGIVtm/FW4Xdif3
kJ5t7JvFXCqmbd0pYXmeYUpB5ApOnaJQ5XZCEAsGhzsNYtmdKHthTMtzsu3oZioUL2FMdB7L8MJO
PxX7uVZVxgLoZKd0pnnddj32hkJRLx0CH0aXuBk0jEJBDzm0sR+03sf+LWLfZ+oYki1S43MKtqaw
FfoZnifaDVd2Io/g3sYdG5PBX9z4d4fgiSP3j5ByQiCQ5rqK7Rv4kCa7GX4WlphwT5qxTMi91tfI
MaNMlZDuVwf2aTgDun98VavxdawqsGIQTKIX9vNgxRBHLncp0tAUUrKKulrwh8b5ZPs3NIGB9xKc
h5a78UUuoVQs4NvPa77dLhMS4ZnrgZBVJhsPPe7dnVWuralFE4qSFJ1OiPllY3ePis7sD3/hEJJa
MmWJs4pZwqkB5ZWAfAInJz9lNAxxp1/E46hpwZR3DQYay6IepRjImswX8CZot2+oxveKwYhrG5yh
+lujX1pdVXe495hglbUfm2ugipNnFBwNa4nM8faSbSSlGC82xUdHo8Bw6Gh8mTqTKjREiBOy8fyM
b7t77o+4Mej7jap0Thp5BOYfz0eJFrUvsS2FnPhXGnixKQulD2QreLUQlZ0tAuEzY9WHKHuu8FOd
OPI+hnY8tfxn6XG9/rbOs1f0hblUxiecZNjdna6vVB3/yahZor2fTTz0opbIopOhMV4HXwmLYUPN
EEF1Pf/odRY2HdURHBLiL4zLShw0SlgY6Qaor7wsBVEbghiMrSbUan1I3USDqkMKN+ZsbQCkK2mg
k8JFxgogPRkHc7HJBPMuMTh/eOavGE1+R6CGiiaat3nxYV2N2S9kDUWQKlTX2cIDhU8++GU7xULy
PHLn2c+XcQhGzmYI7MIVJ87kghDxsLRNfrSa+/vPb3ZzZLAv1+vHQrkS8C1Nz8lTZKk33tHPUZqe
BOoBQoUOU1Z8XLTZhsDWhoSZC9O3ae77Qch0zGhYRp0lLmfKW7518D/LbjlopF5M4/ssD1hT/POc
DeUQqXf0vKWPuMOSmxyTfPNL8G17FftjoDnJIgl2SGNmrft3iEzjO3aRWxRS/Ihg+NB6EXrbyQHY
HJUioxsA0DdqENpqoz5JOpk0FuAg0R9C7PcIZMrgkkg9EcRkai8N6cQF6j3I+P3qMdUJfRGgvF3T
EZ5FhaQK8lXMPbI83hmyno2y+BEoCdQ0wGew8fIWk21RbtZrd/Z0aqBLEqtXqn3I2zY+FvZloSv+
Jk39dGJC+6cWb+1nu83xWvA5lxqwU5i9qrsMTv2XH2984GEIwhye6NnyHVIJ+vGLXJ3Zv/0z/sKL
iW6r01UiEHgmnkh9WZBNdHFnumE34wUrJnuH0bSJiQ+FYe1XxPeSVYArf+m07f32eUSy5YSge4LQ
O6ln+dvX2ylTy2Lq0vBWwxIJdEunjn5C8jJo7wUgsm6djn2q9VrLtc5xkx1fatwZfb55ydWH++49
UOSVLRbhRP3V7zWxdnnYCgvnHRTpuYVSymcUrvVMI5EvSR5EFfVvz+TwaEIrDR95UV4f0+ElTzL/
MEi8pSq3FXHDj6AhrNVALNqbbBTk3g7VA1s7Wuf7L3WKkdJHBFfkBq+LE1++gvrlOUWSVp0jp2jM
INNcGCLx9HT+QbPoFKBx9e+b2oli7rYzNY0ZzrGTAk691LCJejhwyh9XaF7FdtNbzlnLJ+/ztQNE
oLtFeOr8SHVdM+jFKIXD74YNnYEl8ZkMAzgW7R+9HNqUNrpdV7MzpfG8aXySwOVspuPRrpRRCwiD
s8pw5elpnw33WXouisFhhfQ8RIN2F6oIjiWOlZGgkoVcZJ8AWf+7J9H8OqvzNZLlsXqApVZQbOqJ
y4Yd+yzdSSmqGjZCXpMMnDxBSzuoz6vDlDB0FDxr4TKQV7bJqunq4NUsWz/fPE+3fFp2scCXPDqC
WN6Mi5gtb9yNMO+Ts3JYguXwz1HQcYT8EApHPaWf+CZnzGP4geEtcIng5CXVY8jNgqLFjsYThGDU
xD/99/gaDCsVtP712Ol96nPw4KRIxf5V/5ONCoIbBJjAGcReLQQUXe+N3oNmhpaXwDAeXxDdwdSt
gt3gRfeWQZjYzjMysd4c+nyByJVz7gItAJXFOKJZwdHQHKwVGgPclpQwjP/wGjqtveiJgi4ltrxI
A7oy7X1tTAASzCYy7TbjO+fBPbP98CQbR01pqiQ/DKuIwRu3C9ppEJSj6WNz9JDTwYGniZSmyEa9
2IWy5YjmYMWhe4pEZ26+5oXEuYGE8q1oEoXBYqppCLwP6UBLpZ0vmHWGv4naE3z2ox/1E2kMfcSx
x7b7Xwj3+C0+7Wml/yVswqfSZij3QmeSOBwKX3XIkeQ2nAIp+v0o7ynUvshMGSdMDirADoBLCrOT
1PedqV6m51qsOOIFYSAugOhl5XrmVmBdmG+dBqkBL661k9QXZcRY4AXHMtq7MXG3qLGKsIgba/GJ
gOoNwMi6/TMrmnpnw+YMGMs2iIOLMKsOrzZIUSEAk7e42bmEgPYfcGZt/w8f4DAhAXw2zphXYDCl
HhfpXjEuZG5WU3Woli6yAfOCDm9px7WYDyygunRncAxiB7K75Gyq2NIxOVCEP35F4IGvIfaiXVcJ
eCYnKTKHkJaEwRKD1tzrfOyop5GMH/ryDXnX1qVySpgkFSsQ3SNr0fqnw4hXGHj4NAKPRPbGNy4J
e5W/UYHZ960TVOJt+GNFdcgVnylmNrvgIAxFleQ7LogHMTeMFjffu30dXWDiyW6W1KsWKYKO4a8R
NYlixGeLUwRKvYXIG/348heLOD0jqFUlhefjiyhz4OV1zb3JXx3/aAWqaeK1kkmc7v0Fs7+nQgYn
WgyNiiF3YxX7wOmpwlcXcsdmRIdAxNz4KGacpNDUUbE65fpgpdMu43uBDMZx9LCnWmFf4iJDSrFR
+ClJdhbdkgdMrGe1hftgEc29XQBdgFn37bdi/l3xQeQuLp/IfJE9JcTIK2wlBdp19rELWC73fzsE
Z+p59jUgHWHQWSnB01pgdZJ4Hxg0LIMEyDkUkKfhewdlA93gRgcnFmmDi40bF/X2ysJzq+w4qguE
9SZobGt+HzIpESlapNQwCyJ4FdyO+0/2tC9lix2YuW7xhTHGjS++3SVtQETHIyBrrRwIbIBhv5N5
O6BtkCayy5QFTgL3V3se8vdqtc0uzvfz6YkhW763yYbteB6bCgzzJk+gQ15qAFRn9miMGevTt1r5
fkWAr4+e4ykdOW0FbbrKBKj6cLf2hYGnmntIYYjTCDWV4GXB+Zc00kgRe1GIqJe8shOmH0RGPnNG
nv8h1B1g1Fih4gb1ELExzrE6Xwg4ee1fsrggEIF4OuzgRizBRrTVlyANttsNblx4Q7PwypvRMOwK
+yxahKMUE123ji/JzSG6OA2igavazMNa2FDz5QwRO40prvaehi3mjzo79otqyCBe/XgI29qKfrbG
nqSxCsoN9ArNL0QzRDspgmw1dee79FzG/ZMk460CPmWvhqkj5++1yWrFnMYBhbZqxnMYUD53X05H
S+iNPG42i9oPQWmufMv2N3NlBJKyuhpL5oxD+XcLt7bo0IfgegAFSO2yHHCzomMM8qICiwHCCHwq
gXQ2xrUiXwtrUggGNdPktX3x17fYJMnPoHG4jCNeJjEfZ03Pk1eMnrFmVMCLe6tY3xpJN+Zju1aT
9Yq+jxSiIlHjbaH/l2hVgVAwnE9E9QbcjL+UpdPofso1dnq7Tg3D8IAcmtPLfJsaGvXVBV4aXqxg
3SG2R3NDBMIhBppIiB4UPM6jlbBYg7x0t84U/ynRJ5B/uIyT4wp5Q9F1gazuK2IpwIWuGEAn6AFS
o3bF3Qg9uZJBYqGbFbadQTSO0R9T9wcsxBQshTj9/w23iKRBGZ2JzC3gYed92YffHKnThaLSz0k9
hZ2BYQaTDiHuuh6cgeKn1qezkHFGgbXeMo4rCHAq/5h9gQ+rOs5i1nkvt9tme+ym53cIJVyeO4WL
JXJ22MguH32RiW/oF3xGhtLVGi/JgGeAGIjiR6EW0ctVZpKO8znduP+aUggU7DzXqoiX4BwOOzPn
LGLf2UXLQsODpW/O8RvunQguCNgIEdU9a+oG7hQOOMihnKvewUVmbYEIAMr6CSFqKyuZqNBStiYE
yZhslGupehcMkGulFLLWx5gUZ1Ls6waLmMu44qvRBbJymFfadpkTn+PQThSgdQG1m/W2I/mIQK3M
v/MYJDTtRtWxBZqACp44wR3rIL3QcqP0Dy35hyr8R+2yYMqf9Tn8eLVbgChoMj6O1JkHqk1RB59y
/+og6e4SzwvSWGNYPnZtZ/UwA/XL5yGgn5RIlJXzcHvAvMhSQDg4+V8pMlV94+mwHIhZOUdYzqqM
0ceMSZaT2b6/Xs9D35yEj+vYUy5YrieWvumc4WTjqBinM9JZ6ZDDRmMqWu1kLDsDOyZFuFDzCZH3
eiuF3IqVjogMDlCnYOju4VKUKf/LK9Db3s7zNwjtyBBNnNDx/or/nyJt2QXXWG9U2gJsf7YmySeR
ptJGaNy4EwAz26p9SUQYY7oN1Bmr87joQQtSoEh0X1DqgoV21RvKS12n2+xCZOHhpacijBnCg20d
6aP/F5Ed5ukrt4EwpLsqoopJmOCeBQGQnRtvAhb6SAajpdIqAbPQ89GV4bY/lfA58x+foDOaBIB9
6P47uUn/u59gEjr7ldTCf8HINZecCYUuLuVV4TncR+6vaZeRpvaBdSqcTaZm7+G5bttHPgemkHJd
5uAJd/iwYXrdbwY2z6s2D9fME28PhQ4j7FbuCVApPf/5bTYh95gKmoD6spejso+zFtCoJu7Vk2am
DW7dbaY7ERY8H2Rsw6gNtt/Z0Qw3ljcs4JRThVtLc2Y1AP5uZTFSA9ucXInDiu1X1fSMFV+xIwJz
qby9aUFWsqQiKr8AlfvBjZpsVMXitYIct2O3fzROqJ7EoASn7Fs/JE8+viGl4Su+w2TcB8EELHy1
ANHU4x3PEywDCF2sfxwZuJU+PkcRne/N6AQr6WdpbnVoSMylTE2oCIFKbZRT9w5rUM/AsBPv7AFM
zfWH0RqAzVpNXsr0yW6hWJEe12IX6dEdu1VRUraHhsVCMAsDdXWWu9lsNscAGfkglntKk8TkDmIc
1QK55p0JLa5b++g3x43tztpIFqRKRHKBhIqWSmqgdoVlcLcMoHlWzZ/siZOZzZG36ElXhquod+ax
1/vGUkwcoS5QfV8T4v/poL++EzhlTljNOexMFP1CgeZ81sRdL3j4WuP0NOLMXALEcI1NUpkWo9jA
b49CUlUu2v5bT/K77v6YtlqnVD80naWFMWsTm6QEMZdgmK0osVoxSBRvic/cX11jisDm4twVrQIX
7ioXWc/gtSHBXZIzqONIwLyt6XyNg7KZXpzOCFvKdf868TUzvH+VfrNbX9omkJFNhvu15+BwaMWh
6JV9458LT1fzIvKuJZckj64HJu2dWxRF6ffUNDgkro3xlAGNJ0yqqKbvCVblkEz1GZUn+EnIqDp2
A3E5I9Igbuz2HybFU2smjhT7PaVIhSEjilEgu7xJrhAxzVm0lM9EGTRSTaCFH+ru1vulFKAi2dYK
xOukVuFuKDXb3ptQoRLujETv3KgHSW3I/OqTLSCzKVjJ42P/DVoZOfppAg/3zRzZu3F0iNIrIfW2
EPDoDGPAgRFDFrrCTUYYSrq9+ErsA0rshfp16GoFZWfvmphvJ2x8OxvFG9/ZGbtvh9A8w/x08oFN
Z3msed9fSqxqOQ18t5UqgY9vC8D01aILtnrAqgRaW815yKMudx9N4GVD9jTGxBUDhLaeDEUFpPX7
XRR7gMMRow1DZoraDF8bWbH7b90m2XEfqEF8sszAh7KiXfLKlXoHU/TZ/JFgsJbbIAK5v5FakdYK
kLQzGAOeuggIRc3+8M5J8+s2XDyF5IVQIk+Zbfu0b8OwGi6x7rYyah5ZdJhmGhqTTnFcxok5QFVR
2E2xwhoTrIsMJhuXSVk2OE8Lb11MPitDF9mQAIhZCEiF29Vj51plm2wSUAXo3eEedRGrzBqnN9YK
gBzm1Y+sU0vy9q72PdTKxQ9t1yt33jXCJ/zKjjTiY0MPoLZdl+0pqfQ0DOch2J/n3t5DfmNzjNNX
PuDbBuexaqqimC6XMkAcJiT0WSKlidw/4H+Kxyw/2VbrGZFECohuUWH5BbHccknOQYO42nQQJ50A
ugvakDgMMnxix9z2nZZBcciDwJENTHI5Dlj0xQxiMaKEgQKxyp1ruWcgJ7IkMPWv5SRhmwEuLgJg
K6uXIZO/fzWtG7fpj0Ko1L1UMQoOfh3V3vQ2LoNs2F8B9y4k5GgMmIj0X0k2jR1/W0beEccEoCqB
xklbNwDNFg7b5ZqPKZ50Wha6CpgQmNCBdsYd3Rra/qGdrXXdIR+gCv/9HG+BVd1AU37L3oOv/Oc9
2AXzCqE+tjH7Nz8armTb5+SnVazgJXeSoyUxXkEb5fvAcUQoEdL5teVJq0ZoPNf1kRWwbIvbNioY
JhGooakF4M0W1DnKffEZKmcSvxKEQt1tkS7bFHNpRFZB5rzDW4hQjnK3/i4oQVf4EyuDnsYAoKuP
LAXH3YLbAqhG9cxvF8BsH0nMvhxUP6ZlAMGCF7eb67ic8LNsXJ+3pcKQLYfH/Sfn8+1R7xFK+SUa
ZO7BaZzpMZMbkmzXC2evk45lEvBV+2dV9tcuzKBenETyflDA3yVkVmABD55sB9l4d7IO7fWQlvhX
Cv/aTQ0iD2OoXox8Mpuq6e6NpFMB9pVOIKP0YMDInpvvZuz4UkFzBYIza1sE0OWIV6Ijedt3Qw8x
S54hKBYaHLlpN/tXap8TUQMVNhTveFCiy3sf3/T8zWNIDQINdYCQnO9E0w3lu1cxO3/80TR2WbC2
Ult351B1IbwkxObqRhFzUgm+NG5z3cGFXzrwCb2J/abuzK1EikpSjuZQMwwRQMeLXRK5fcbezQsN
GFz/YmvcbepfbIavJfvtftrESu6MIeJ2TIdrO5Iq1nvIfVRcPi4qMT0xjMmsny2UkAU1MDd4XCuI
JMHlERZFia3xte4nzcqy2kA5hlg3bczo6FiusrurQBaV/cL4Cn/r0dj+Su3f5e9J99t8lh6I375q
d6hrp/J/zNJwxzHr3SInhfiRK7r83rOShqRhipQyHDIXu/JFQDHR7bPR2LOCStzc/+f0AOwGADZF
6YFv5DrjKpKFpYGjBrv9gyDjvVrykwZDkJ07Ls03x3mBrNe/BsBi1BUXYS035PsnJHzHyj9yA6Ui
gqMhW8dAZWOE/WPswcVFQJYRa7kCMAcge2TeaJAUHCTxAG7+KX26NnGq5dHAlRiLi6kmTnzj26/h
jf0iQMDcPuGxI0rVm9/F/Ar/TIc+kV85whRDDTb2vmcsef7UAoO63ejV4XEemcbgmGUU5RxFndPy
oDpJ6Fp9ZWa/drUJkubifBv9kyfibLCFOjPIFrmC+fyOs4/GKIHtj0y9mEVFXpNV018uflalycYq
AZBOAf2gQEbhh7ylcHcMvXM17bAb5vWm2K8DuQ1hhK0u2Ek3ZEXR9r5BLIVJiurvfU/2zo/ao1Le
CgSEy2CZN7Aw1OwrzXLJCICcZpZc5QopmUpTE9PKtAzB7oBfnan3PxPoD/Pyl7ud12zy+hfT/Seu
eRkiHtgj6KwwmJcXrNP+DEZNj9cYoVEZU7DHu4GZ+u64N01Dq98adAWZ+bj99EgkfQwc10eA+Sjr
Z5Kye7S3l8NkfbVJrhrnbjtzuIM6w7c6TzE9UhULmtWbvxIGzamEBBR4B8nrQ0bCpMaHHG+z6uSA
sgv8jKxnBIogdVwJJ9k8HzcHRLmi69EBtFJ1i6CjE43Utfp3jPTZuVrj/lmq01INdgoA+LEI3Wda
Rw9TqsUMdi3r5P9IR98I1MmbGF6kLOlkyKUZn55PXWlv4U7aN5Wzf+iH+7aM5HwabfsbXtxnCk1/
JeVlyLY1dWtdiMQZkDoa9AEN79h2dp/4WoBNCJVfWjGz346k5Bn6W7dRDSgK+UrXjEBa4QTCYBX2
x79q2fsmxfUdkf/+yrXL0wdkNrAq+Tkxk5ET7/v9VtTCTH+nKxrA8sSfdRpQre9xxyzk+8yhul69
A3glDcN4ZTgRJ6anTjEpwc1LW1hEkQH/18KkQ8+gWvMUi6d+XZzfDc7ONzZm+p1sy6CyQngmxe0X
P6XiJKT9ZFjKYNNb7kGPf7ctJ0JADV2yYSvS7FOoCmFYC2Oq4qWESjhw2mqvHiDzNIsHm0vr6D30
qI+o68y+z9uj9BlrOoBZa82qkbnAo2/mPsLQ/DHUoYC9FNVsM9vRcWpxqY0kfn7TGCDygy6TdUdq
rJnlkH8R+zntMsNHeDBUrUR2tsLK+h2qq/GUWiYahpNRYXh2EaSaskVva1hGYORlX67989hCXDas
uA0joTYxhxh0OUh71v0/JvVhmQDSPx0w+4bHydqw9U7n3UsyikNzvnpjPk2L0WzED36QrSfGx2PY
goi4F6gLpJIxI9qWX1xwSTSuoWsgJpA8arxh1zxGYC2lk2u6yl3pcgX84xKjabYTBLcL2qEKpgSB
+sM4P2KCOrPT/PJCIfi3FkovgMn3OqDacMmSJlOIcj1HAk88kufuTxIwcvid1O6zKa6fAeUisfVU
bnpRIgj24hdglrRIe0cNT7oellRwCdTnz1Tw5DfyTsxiNJohdSOGGzKJ2dWCPwjsXvVSUs3/09hs
SsgJtIXE9F36kMwGs1YQx6A+7goRGt95F5vf7/sOYSP1+7k7DTnWI6QrZCOfQoEdhlPbESeGmoeP
9IQFokfvOxKpqbbFXBa8Ca2qmP1xFaj9TLHw0fAFWrMOH/tJ/bHPvr6kz1MW+xd0l7zsAu083Z2s
PuqbOZN4CwpWx+naRhA0UdHom65g+ytBQvZgLeEfm3F6Uazv2W6pKS1yN9aiCNihkvbjuvoxvhbH
tpSlB08VzjyNW8wjJAhMyGW3gU9utny2gKtKNKReoYdiOawmZ+glpZK1mjYie4AikI5sndGkBAls
POm+4qTntptg5hCzjR41/UBgpXHC2oI9WimPocz8iQ49N1oxAEEshFvF87mvCo9uCOiw6UIsiwvC
ESdAaRaO8BZhxxJglII2Ex5U7q/d2s3FR4lJnzjHKvfTArQLk4hm/Dhd1mjplThBPk7cfKBW20b5
k835Yp/jtFej9r0PacVKLM+PDL3jcsvo8qPFuNAM2G89XGuFe54WnG7pX7KsapIKxrqZt1Rne7x8
4Aud1v6QhWvB/NU6Vw/HT6KQ5SM0JLdBrA+WiTZIxNgf/T7tNTROsNkL2fA7+GXP/mVcSI5oi3pd
T/Wa2CGbxlM5wQd7e32F9x1uXJJCPX37mSyV3SPWeJo7UrWrfsEppeY8aOhUYW0mCcD+t8R5xXNq
PHMaHuCfdmTXRQPGPriRNmtSHImIG2uT9Gz8toM9bP50NVWxNoZZeeMlTW8IwYtaINoHVyXAXjbY
ZRg5fDtcUKTLaouHcpEEQ1CiSZ2mnQQoFxVj20tD3+aOVhVgnut3dMJ5lSryrKtdBoAKlPRxOAUw
D4rXllbpN7peJJQTpS13lBMyFsUmOzXJvYb6K/LXknsyKPLWaRgs2kPyGb2e/b36nHC3t/NX/811
gDR+hS673RRE9rUUq3YZKTXJZx3J67sDq38jrU+Ru3Y9HwrsXGyZF2YhLruUz0z+7p9hh0kfpMOu
tIN+PsBeQwqkMQtYbPdWOXo5I+11yM4/3WnRggeZB94l7IbNaIK0NbMIzxsFz3NXwtjI5xhokTP9
wi+nlyq7tslYfD/w8r1Z3SmaDzQuUV535S66uunz/JLchjDBZqFO2Sr0smjhtCB/GvCcGRKhfFFQ
LyaUdfHOI+MNgz3lv0b37YfJlr69NzZep7pto5hG6DsAMG3Pljp46T64A5DFUoCnTHi4gh69HoJE
YVd0G5vaZ4i2bWG2ApQXreyy9FrKoH/9uheAPTcbd4/8Z5XFjIf0QvUu0CHyXq0IHbBRrbfMXrqg
80NbYzg0dWj52ex+8vE/VdTFr8RuZYHWsZwSx0fabHC9ob2gtDOTdcnVXlME5r7Piwhw7P+xhetH
AWaqwzx5EFQl+4KYtNdIBwUW2WtdquYKvJfJ2gvXhSO1jdoHO0eZhfx2PhNhFQ1jdlTpzEUikbqq
dmnw2qUTPzqDYvotXC0fc1EGuudDGlVacr1DaHiSJ0RD1QJf5+tgzJS1FpP76u2jV7tdxghd305P
snETwQwg88WV12lpf0967Lg+bABWDh+rDO8/5+I2loWrs26QyxawTwn7MVbbiaCx0HXpseDNt9hR
4W1AtqMWR8FxZSwngCv99WLMF+V12ymY5o154N3dcsh9XqdOftcthfJNva9o/WmGDwbzPboKztEB
f3pf385sZ2MHUYqPuZ0rnkB4/NN8yX7HrhQrtjUojYuxhKbXAGgXzMr2NcT6/0i9Oc9xpjtoBOMW
mKP16LYGluPvaDq2W80Oc0gzY+ne/z0JFcic8szKdsLjuwPjmXXtzTj6Z9KhWL0z+2uDxHFxrG8r
Ii22/NdW77bjQj6YeGN465+dCbb0b3KRquzqGChkSqzQzEAc6cpexGqI0chxAOR7oOVDtk+Ei1Gx
Sh4tm8RVH9ZrIDs2fUvxHa0feXa704v5lhpKZbGRTNXecHIyy8f9NAqJolLkjZMYWlfyTGsgK6J+
5ipn/luDGyRpb0I7B3C3CqgcDrLOnj4WoV6PLSpeZ3En+jwZY3KKDa+ymYzsDwzNPZnRV5fYYDOE
TH2MTbvUDzYPolKglPPr4zffC380iSi7mvsrpTKkkEHI+5x/phd8WPWaayS/MoyfbiEkiPKfDv2Q
ErOypjRbt4gTu+pbjWIcdag8a55nPfeJbtx0/hLsY94yuemaIbACeOzo2KQ7piEiXHnZAVQ7sBJz
KxOd12caTUlDqbSgajIzsfGmhJhz0jiOIxvyOMLL7zmUpP9mf8DNKJcExnKGS+osMOy4p/aWRyE7
m2L3mKb5T+mxQR1bSVqdnQiuQz/bChVKCX21fai+zkBWpIuiMsXsNHhNGHNpU4sq2EaHOlgs/1D6
IJIl02tAq/Rk/EW6LETeoEJNXM16MsweNMOa54IADh/KepkcfEQrBKSCSipPn7iRNX2oPRoHLVHb
N9JbUk3aW+IovQ7K7H9GB48R8vOPVfsgkEKY+OHv1Cn9snI/lFQU2ht0JzjggAODtSJiueIgbIRz
EZFvJ7ALVs9F3oD1sO05PRv5WaSeQUS/LfI4E6sIsHo16Czr5dVYPRNQ4g+yqMf23khcjx8Kgg68
HLhGg82NXKhhzDSFzzDRUqp6/byXmJc=

`pragma protect end_protected
////////////////////////////////////////////////////////////////////////////////////////////////////////////


`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-1", key_method="rsa"
`pragma protect key_block
WPJG34g1IbOSE0VpbA+jzDpWiUgr59F3WTebCeym0EepnLxRoPkdrRQ5HCslLKaof0aU2iKLVe9/
xiUVEZlG9xGxIeDpDI18kx8Jt+SEYV8EUM5F9pg19Mu6OMFU2CQw6fu9JOiMFazdStRxt56QnvSH
NITOYWziWD6SQjowtSE=

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Synopsys", key_keyname="SNPS-VCS-RSA-1", key_method="rsa"
`pragma protect key_block
U8yl3g6oC8k3YIr20MwIWdaBluANjax3DChH3fk6+gdAgA8Xhrnf1inJb4JovZtjpUouRBs9+Yeu
7xpXx17uk9vlM6vJxLinhZNeu3Idmd61tv0DRvA9y7HaIPxxWxLfLhABtmjLjxKHX5UsRO/lvsRS
ItawJpxuTH1bFirPDOI=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=2576)
`pragma protect data_block
Afn9oeHxDxdYDfO6rRoB9A1M3QoUzWVuoA7oi3o5+/j5SFJLata0MK3w4acZgppr9BJrXDx3I5Tu
gVsP9QnQQWATr5dUSOHznWPTyT8FeGddTEzpRu52qRckhxYKezi46ITCVXM/vDzVzmyr6Voh3IFS
OKdP+qOUkZuxm6XUs7/f3OzD34xBe+rAP/xa1KyWkcZw/ZNC9dxAJNFLjL6DXM2ja8M8ONAO88Pd
vwoMYIKYK6j7GINWmZHcbuf7lvHOnxjnnCZGlPQXGBp8L9UyM5o0l61UHR9XSWRUH2TRRO2nnk8A
Y8hGbQvLoOVjbCJWV7P9Os1pYX9poQuPRV97JTUh+YA2dAeJMWkOC6kVE3tZ+KyDwULNpaSv/lhu
QrbrY65bBIFFAt2KXGQBN5e6SqmPLh3NP3G4p5yF0wwbB70Co+mo/jldKpoJmBGGWVN6byuqySRX
YpAjuIz9TXgy3qWmNwPDIW0Sihh2Sexj9JaI/Gik495UBIVF9p3HGx2kQqbafGAeVYwyAOGHs/lC
2TlnEMuOtFwYgh4EyyDgy6RGj79nOJj6UWdSiydRqsBjtB1ebs+VWYg1zlkvaVs0UxDBYYo0qRQ3
3kbQpXK77Od5vNITauygS3Hp2Xk4/Bq+EFeAZJ/irtBu1IBUo/Ny/qqqofForn4p7NPDuDnSlKsJ
O8OOIta+1w+crF69STTWind+51QTQ3SOczDQ/+wIFBBglahdfwK963DKRKkI9fhESgGtrcga6mHJ
bU0rYX8Xi6gF19T8Z9I7TsSw5r4rbfA62DQvWrKKzg4O/00S4ir0s20tJRIJfEm+9FVwTkji4N1i
Mi25aUz64A19QuGyPlwAAoEshvFdVgCNiBjjexFys13zRxoLV4I5pC5QDdZBKqlKjfS3Zuo7ZXBe
5lIxX43Je1D1CQXYCSW26x3Jun/SRNXr7k2RXTXc3OWbBT6fSiRYHsEZ5NiUfmEY0NSD6yVTWQR7
gj7YIICrs1XPcRWx8TMYsZ5RN6Aa27jKERXwTyGgwxv7AWI0LMyxJ38N17EpJL2L9eO5OpTQiJbW
7COviE86fm31RHdpYgZu+70gIAyvv7BylIuwE5J/LIiElPNq7JmgGVAIJ/+ealF69lA1t6jTajTj
KCc3Ia5XlQXIYdrPE0ilaN3ia8FeA9IXU/dOp4potHCciBJG3PRRgMI9g/tCJASS5t5ulCu9a3Q1
3S4E0ougbnzd1KUiWJ2AKxSBYafETCASk2kLpM8qTbDu9Cb0HoC352MXfCvJIuM3YLWVfwgciuIt
L6zgTNhxc92MFq6yh3Q8LAqLfJY+og8K31YvEtcZRtwDgpTfkUqzUJ1n3fLTmiAZs0FbwotM37DE
/qNiKLLoE/Us+vk5IN0oKboZH9/oZ+mGvyabiHiZcCNjTHw464YA57dVO2aMSBx4ve9IPwImNI8F
+4/aRADEMYT1U/NUgrTeTkVAyJgKExN6WJoTqOXbom7LQbQ1tPtTXcOxYrWA+Xjm6Xn/O34AOjYu
RGNWY5kVzp+EgiDQbG0GUq3oHjqkKoCMg+ixOsLQskEIS+2cq6YmVzMw2DbsAS2cOzxnMauJHYMb
MKn2IS78el/B1OZif+c5Ykk14WPI501gLeUwieN+a7TsnBIG6sGminl95nz0ANlHcL7NDGJjvo4f
nrBmjYZLp12p6Ozbhq1wlpedd3dR+86SuyZJQnEvE66iakujCoB2qa7NaHYDZNkgrVW18Ha38B7M
m1dvQ/K8ocx9vejLxn5oelrEURlPm+QJ8Zae9DM6O9gtyVf1JeB3Vu7+brlenOAlkHbI1dyuFOlT
rJP7fyaWDcvx6D4X83LY1SvbwVfw7CoYv9ovw24fO89WTdPepVWuLhJUuIQG5nv50bBfUNupWNkw
hzrj9GcbOX1gX6DJOQyfjwG55JdPu1CbGmFUTMcOn4NkyjXJRMbn+LCOPAeEPWT02yJn7CW+6VrX
rqRr0PrHe6cVYTlWMzN1PXwQXv5WFg5cRSXASo9bc6GCXfcG0wtH+koZGDK6F10ppeG7WN92AisH
dPCVf8h0K3Lj51gdXj4rAMDtxjlQpJOdyYd8Vvjljv8mgceAuFjmLNt019CXEJgM5C+5lNwu48Zo
JDFOns4ZtM4VeJyr54ohgChF2alJrZVHDna1zuiTxVL+MYstQXoDo34hcsTtXT3RGBKKYaqnYOuW
Q7p0ssxLu6MzLrBh/6DGFPKJEK/qmcsfSrfkLBlXnyernmw3NZIV/iEJ3vGISE0tNlw5supWFBw2
8Qz6WTGYrSiU7SOo3ntwc22G9RMOmFi57+GFhy6hNjClX7UAWWbEpSGO13hOmmhKnt/meDu7zD6S
xrYQY8GYmOxegZtS1SQaUSTWLopoQh1YkqXtIH3F8E4Y9FNAt8RYVPsoldFDaBJZwjrsCHuvAicK
EmjX4M9SwaOAbmxBt8UDMXsK0S933BzUfVlEUMebUHNQY/0o+6V1J3LnPBThLJ/EgTTkAFNCaiY8
vUtjzYJe/gPCQFqEo2bd/NMlm2N7mZfxXxWlQkBucW09srQv2FeLEK8UAxmlqvngO38/UZ22CL7f
oDA4f00D/p80JAs5qBDw0PF0zHQ1Z3LQ9KtBaGzNUWYl/zMxkbDNy05BhxBsm7Xwwc5/M4QuQNtD
sjZouiEtVy4N1TTdrdam4l2gywLm5zioI/ijlNCac3igD5RmFVxzB0GTayuWXqC11Yyx3wxU2OMG
d/CrtfBg7dNWL5iRxqX/RX0VKuXfIGQWdStnAyGyqJ6lLiQNlG9CuBnV96V266c2/Io5k4iSwl9B
L1Qy4lFYpj4B727+V6BGAYAs5Tu9+qYo29NGobzA4roQ2umr7hi7C0OtxcLTqvHT3ufwjHVsGkZ1
2LXa7HuWSEz2tVPX64eSpLQnya9tqU13Nj8Q1lCmjzPtwZtxGEPfM89D6WX0lnQPjehLsuVg2KaE
LFlnm5Qe0vCxL1JAWmx3h54buXxPmNKJAsPHPUWmelgdBz96FXHUuBkiojgx915DCd2nVL0vnvOp
VShBOcZG+Ak1E798p0Veg3oBmgT7joo9cTqJJNhaxj1T1192GRCafGGDPMA1CBR5IKEqn3aC34qQ
j0Akf2iRpLjgxh2JXWzfQAJGBucGQvG2K0bL/rWeWcYhDALMIuNP+ugrP8glVVcHFVaVaYQe+ogS
zf1Bb3kMtWWZlv2g+a2PKo+HI/jd6xYfIcvToHcDE0DITEuHfFf6fdtFPdCVk53niK98mIBkaBBO
wB+kVlU/FEM+oGMdY1duh0LEJOkoFpcR4X7rmpzoSmdg24n/nWcIKuYqPd8DgOGmJfMqnlq4riX3
kRM8OZfcRlj4JqJQEdaSYvkgYYJIupvm5pxo/XpqEv0qXRygkBC2pRKaD1m6C+gbJ/eDK97MofQ/
C99/cHEcC5AnZew=

`pragma protect end_protected
////////////////////////////////////////////////////////////////////////////////////////////////////////////


`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-1", key_method="rsa"
`pragma protect key_block
SMb1p9ylkdc+u6WbH9CRPYeu4Ya363Ddv1SPZcP1uXmOuG+rR5DiLM0b/UK1SgeKeOM0l9kFvXTw
GGBMKjbqIo08tYiFsLv5CRaGGhZ4WZlk4v9wxpDFWY+ngDHlGNRMkSEfF1+CzVyubsQ5QSby96Eb
Ypma/UJXYdEBccHeHCg=

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Synopsys", key_keyname="SNPS-VCS-RSA-1", key_method="rsa"
`pragma protect key_block
zhEmnfZLR9cUZjOcxc+4Z/ohG76lN23cZe6+7fZeI8jGTR8XmuDmGqCozXT728ccJN4GTUqsomdo
EYrCY4viiERWdHx3irL5viNm8usm0emPQzIyjA2ECrZERb9A4ae8NlCpu8erEiehPk9AjzHAR3A0
gEBNVIBzYn6dmNX0D1w=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=13664)
`pragma protect data_block
M2KGn8k9D2oWQPr07pIp92qIb/IHY94FiWD0RQuMmSYuJG6oYT4nDgxbPLCE5ms1kL4pNcAjGZ3u
lj21XrbTD7TuY5tWJ38ZJRfpAG70buqhtaVm1xG/QUs6q9MgQF1xyARgCbhqnSveHcf/TDe1J5Ls
kyit3YDKcuGn00nszGSH7gqjycCRrTRaWMGZvIw4o8xXx8q5/p3fn+p+T5dsjKQ0OkWghoZBxAaB
EtuvXqR4c1/WNf3F30qEQbT2gC3hD8HU+jvAteKxVrPOXVAxn0qHuzycY2OZpWOnUZw6uSVyVzLh
1nw9v1wt1+6cwIdlUkb/D6LJiPVQWFUkjIvGnZzVFdnKBFsF/t11wRipx35R7gV7yLUQHevslG9J
ofI5kQLb6t1Iup78fPOGlxDOd4N0Trc5rMlr4oXbdqJeJ0c0wCNZfxCxZK+qFdVZIMLMJE92SmPc
+dptOwXs0OSDamjPaPzrWlevrvfU5eNnDb3hlkcpIY1ai39GCO5cIOeb9fJO5sNqEI05pO1kfsl2
QF2/YvgImjqDSVJoh0I3xK9rx7ksKtwAeoSe5Wdx3ZZeIymU3qPzWGLdHSw3sqEMNvafI9AiNq7r
rixcUqQGM3h+rZ1+rJmTkLUVOj5hy9qNeoFjBVrP2dbCP7EBjyG507XMoSJl7so6y1kQufBap3BD
k7aRzDIAP0F2VoSDaf+xpHZyIXXNQWSpg8sNvGrN4m33dHb6AFTYdxfF3MWrCmfZuK6vcsH2JQKN
pNidhxXHTDtpMgQcQM1/YxiZg0mYHAPICPETCVfV9EQmKSvT/cxeRFnNCuzjW9TycPM4ZidqtOA4
dB2MkZTZglcbN7QLbpyvNUURXZ4cpM2QRPyMD0ltbpu8NDWX2a7GYr0R3iatZljlHdOstLmpWTNn
1LYV/0qXECRbNRu4u8twdCR2QL/qjWoTmFq9PbqeYm569RvVetWFBWtr+I4HIn6vjf38AaTtIs/l
6qs498YFHm/I9YObuoHyYd9r6ANdVjUChjvPps6bubVXzdXn5OWc5SnKYLoqzDP32abtRh5asT+x
5EtlyDA7TZ/M3cB/bIdSCkxGufPpUZtXTIMQuBXXFtdBLm4iLqThsN9H64M6cbPVcOmbxidl0iWQ
yJmNi8Bzjl+5GtFoAMQFmFf34bNSbKFmUS/CtAWruS5lhR969I52Ok4jrM2RHLzzlZoHALkTTeJH
w8Kv7YT9kCnNgulQqprLhPgB8RNhK/46KLF564RDdvYQiuG1z6TCSXG5dMwnqZ56uyx+eMC9A0YE
rd2IiJlSSQkCS93rAKzj4cGBMZ/HLbKv/hoWDN/VwmpwF5VuWqyhPqvp5gFWu/o5uiL9uWY6Vh95
HNwCnQAhJ+a8BlK73ank11XgR0YkVtbGzWmgDgyoYSytHTfzJ7lzk6aRMe/oIufA29sWFQFbAak3
kyre61I8stD14WLwwaWALIJf73NcEUsDqe0fgc8sR3dL1yiyl1TEeJD123Tba04zqL4gusHN3Cfd
zygE7pL8vJsw9F5kQoSxnZ6+NkLVmnljaL6RD0T5tMagYIE7wkldDmz9Y5CZlJZMhgni1kiHKkec
JDBwvwEkGBJw/7/a3M5mpy4T9gPHN+Vtdo+28vBYwnW2s7ZqxpkaT90Kn8uuN58B5HujY0a8eu+R
dNgb9G8IhW7CANe8F8JeCfVBgFFvBrLKhVEBABwDRvwSIV6RJ+FhElGvqRaeT+1ofogbRvcuKtrI
Jx/Hcnt5htkzEjCkFX8bBjgtSsTgWkMujeVvl6T+mMbgMDyiETtjrX8j2Ra7crI9rqJyxQbmq3G6
InwAzt2PbQ1VguKIM5fp1Q70vEuyiSI9e9MuYw0EibLH+gJ8sv8r829m3ZWQpB56VH83q0njvuFr
/0IZArdyDC7AEqLDpJGKf1s1RylQk9QdbXClB6+PlR+eV/4hzinAh3Ibm/WF4TkbGJlOPmcXR2hh
HMykvf4RJeCCo/iGzqQxFccy/jFWoHsC/Y8Iguwy3IePde0jmge8lmorW/0eH9N5vE/UuiH8DtBE
yR16HweQWW4YxwsEtd/o5kp7qhD7zw3lhqfSJgzk5/eLsgJ0iPihGMMclCrbuuHnwhek9OqPQJq4
CrK2Jrc7l5HLxso+XPvPLFjqG2uI+ruKeoe60QMooAAT2nwcBoN6kYq1WIphHd3a9R9PRnxksrdP
8jX09KFMzNm9WyK3qEDFyS1FfkFvoHvA3sbf4WbqT8lKAWohHpVm115kEh51v48jFS4tqxp41Ern
L9SX43lS+ejM92a5BA8vmJUqDYBZ/EyIZJ3vnlzLQ2UXlcAUhNKC4yKhC7Klu3J/JPV/mrIiczLe
AxHWuxzXFee79PSnWOHpQSZUL4/jHO0N982teCnmYH2kG5WRwm8lewN1ZsGsjsnUvrUwwRqwekIp
73d+/wpk1FLfRqGzKYs5UYkBfQxt8kOA4f+MAhhMKn84SWGSzNx/LuP8wIxrWpTl+RY5OidW6Kvn
jzJ6qjGe7IK+zVYMQ4SDeoc1m+nRl/mthoxJDajSxWZxodxCURP3Mqh+NCM/JSSXEpZE4iFqY4TG
l9zJxVZ5DyCPqJNf1x+NGXpgLiOsYFRpDw3dX08/czaONmwZSbUNZEv4TOXj9IC8B6wbsKBpLtUv
E3MfDPtDh+wCd/GsQW7k8w02XFhxdo/n/9AiuCMo8+feeTnfOcE1S+e2LWkcEI9Zr+PFMcyV6/ES
9RRRyK4cFqHO0Rqo1HnPCMyJEpzB16I84RYwfA6V+yaZPkRsr9ZOisYyKHgYhbeJlqh5Q1BBCXIo
OulT36U1iWVFFIqpMwe3bJDSYlPgcKfwXYCV0OKDyfUGVBu2nasXEhi6zEbbxZEFogOpFunkxt+X
rOOfgvFyT/bcFbcBmS1lo0o9B9R3N/T4imCaO/cGlNRXgnMOLrSiZaienfpLwD2uKIUxrPTnbU89
pBThNb1+hJVki9m/TEntZf+Llez3sxMkyc3lmtKvbBgx4O90TKg9ap8DQRQiJArhWoDMzDEFovS0
lHfBs3ncMlDOKWYEOIfcYkouVIM7fwYhsQLGhoto6d2KJkh3pA5pTChc1yUX79JcPAby0gl1Yxw7
IKG9PDM/XX8gVY6xigeXwE5L18NqK/SFKs+P0sxBaKmAsBOCBoK7QaUq4k2Tk7SCG77756HOqX1/
aE9ogGNHsBE/gTRmJVaVRcvx+WVgCObklCD7QFbJ8AYi7DSSoDRKR84HRwOLAYrIKGSPYsisAMFc
JJu+eB0R/HdcNXD32hs4bbDK9/TFXcTyTMYzYuLKqg9hYMZ+wuyBof8w5CxcWviUi+bRv+KPAKSz
tUXQ0JloOlowpk5XbmGXPuUiLnYlogGWpfzC24/Mna4uL9OzLdkdN0bN+hjCY8u5fhLCuS8eBbhb
PVWmdtL+IHMfO7HZF8iDYZNQBss4h0lBHFAmQKhRZ5o7ZKNvPovCuL4XimQUx0pcEXoH8UJHrloK
0zgGoopPAQThLSunkc9EjG+MVY3Zgj/pOb6gRcXHd2aMZcSUzhjEsvq87rCfkr7tsxt6rw9i8d89
d7ZyIL6OktIearEKKm6ofImJAnzexOvZD5OHtsbOtaDFpbU79D40NquIXpKYcVH/UksrAUdoALgt
Wb12HewLfvX308G+H3QAHQaATksDg8TO3fjD3JFgLgFeRN8w16b6Srua0XhI0VRSAIEA4KKzhc/F
Ep6QZ0VSNjy+NyZaGKo/EannKnW4DoA9Dgqqilz0h9UlRnx7Jkr4PS0nCfTGyPvo8bqfa+gbCCn1
tuhU5KnIo+F0LHqLpSyYaj4yRQuqPSjoATNA20KYzr/xv6tAAdqg+IaHUSC9YsLnlVCD9jkweTDt
3YqqS2Ko9phX49U3gB3sLTRYzp0tAcbcnlE+5KO9hwG12BIvFQYxyWjHSX+vn8D05NFANzLCoQuN
XK5BlaBQDZ69xl7b3CoK2MH3o3H7D6qzHBWU+iVxSVayprsFQZt+DDz/wv6TnIk+2bTFHEhjzfg8
drBo0yhj/64cf0BoAm3apLZZtOmqKf8NnrzqsSslhLRmJn3XHQtJPBPEdtNC53sV4qV8THbJh21b
HnzxAjSDYQg4wScZ8wpaPhNRXpaq4Mmbm4JhGxDmeigjJl/WqB3XUb8hSRJJsVUomRoVmKqlL3dT
F5/eurPLAVhUYc8+oy6l2WjJEQKsefJM/RsXLa0UlhXDmnGJ0ApPjKXxd88TT3QZ3Y37uAHyUK6e
6s5mlNw3TexMlhSSGunMjVV1Gx1X3ZZmWYbbLWRP9FSAnMV9itC2EledxCMr88MApcfLi4U5gNu6
rWuyg4vwxOnLDMYIRDL4RYEYsgRaeVQiwodVWYtzNPw0ys4JYz7BnNrBehIScFmG3kaC+T4Dv2HA
q903MpPVdsUPSQHBp1gxJ/8SpISw6EYJ55woZaHmwQ/KhpXpbbzKZgXUUBkYcEbIEaOOGrko0dva
DH2eXklXU8vleIVxhHVwxNKGDyfj/hULpFQU61WzqY7WP0DL8nLw/faUXfY8/PE7OnZWecXOX5EL
Bpn/Toyl0xg1DbgZrdo3ztV0DCEjULXrSi9I/8tp1jJHq6VC8Kz5j77Opc/Fs/UVCS+Fmav4EbWA
43rsOKKiLuPPdvuPeR4d6335jvZ4Z+n5PRyezXoKrMveyWNV6McOGaEeQfdg4ox7HrozYvPcc6pA
9u9G9lXlIelVZebaIiTODma1sH1cQCY7PNNeQQ1BTCdQZzu+dItsxhQVUHaxmHkGhCSkVuBtyvF4
KEqSqdYS74mQ4rKdlTdHSiYmmpyVQelkg0gIXRd6Y1q6rzJsn0DkTuxaF9k/RVORtc6BBeHwL8CM
jn78OZAbSogmAXS9w+o6x0klsZi3mLekPIzTowU+oWPyMtyK1JMeHP3oh6LWFLj/nCBeVOuIC/eZ
dKjnfc1QdhxcFDNp3w1bj8gFQYbvItr1YFc2VDdZJrbomPlZ+OL+ivJ2PfgQ04rjCJ1vAYADxmu0
4l2ZOTm267Yi5Iz+6FXDNZ0RoHyCA0lAwgNzDE3E3YcAm1LBLASbixmUst00hOId1QF4BDP9NUCU
3UIjkMYZ4zZnkTpdjn2mHoI2rH5OyIAhmccUYJBIH7gXjPP8/vi86WXFk3c0LY5lYmYrI81pL5vt
vEY/pLoRseybG0F01RirY+SWU6Qa0jFZI6KOrXU7bHOHQ9rK1To9XS824Oopq8o0lqlPKCTsFuDE
L90aIlnLAylbH20FQa7l7WMn3D6cDFsCL+hYesuC0SBlY+8/hk6Oa9rGk0Bin96IFa+jhjqzVJ/A
3nkeUIsOXTcg5eohiwmwX+nOVvx/xoxVOn2QYgTMJEyuyDfMflzXI+PwNULjlc3mAWx/RdcANeL2
mGOvql1VcDcHOEUWI8vM9mFY1LHlY0IzGYFVV7qe2RR6HfAlRAljfHxv4DrlwSMPtzeVjW/6MSyR
4ou79KT5SIk8o7V9t7wfAtdcTFI+8AXlugOOeLmih1RhkNPyu20q0ktgENeyDliq4tQhIwmWSbPv
y2tjKJoo8Ucu3fzin2VrvELF9HfPhNbXPv4UsLV5Lx8aU94hN7zcBz5rWNCWbIR9azov/1kOfRFu
mOoh6QQEKZZtIcFDcX/P2Dm/yeq/GqTdX9Dfb++ouox7pWGfJBZavega+MzDwggLcXx3oIUrorLk
PwJpGB7HdiYH3fmjg7WVGtxLAfTdYTDgaIbb6d2781pNWN2cXWgDrzQrJHI5zXHG6yf1P26+EEsV
AeI+LHEuYWSy5dpbfiRi1yfZJJ9rIssm01zQQOnJfqNg8UVdwg4b8AEezkPBixSWtOoC3biaE6Q7
VNxAIiDHtKOJbD5J/v8K6BKNQfJW8yDFevQa8Ng4WyZGBusZezmr1u/giknajxe9wEW6GrrOOiyh
K49uAVxowT8Bq8w7ufUjxmsuEuTejWZUwXTvFXnjLx98b05Sswr6+X+wpY/PHRrX/DEYcF5o5nag
jWf+4kcN+oICyt+bJjaAB2by/WdGCFyw6DLXCvyDIDWgYd5AAUKFFc3M697doMInpf7PNbcgeBZT
m/4YnEWbCd0COwTDF6VkdP1sGhX8K1ahkUMIgp9EchgkBaITEFaaPCtvz88xFgBthWzHnpTtzCAy
NqwhAX9uJaZ9z5+bCtmyBVFq398OKx1Ry0ChOa2izi6XcRdDv5QSKVcNApcGVgYn2p1oR9VV2V22
TK8NjqtgQHAQucBn5S8TU5Q2ISPlB7WmZjOy9rJ1EeNQY/AQRXGDYFTS9V9/kiyx9O+01PsVbkT+
HbL7/VlBCl6z3Xtq8mDo3Zq/w925Ky5oPN2PoEZY1yN3IW4Z3ga4ExhjwR7uo3pqGu0lEvr7hd7U
KnOVd+7RTYhhMGxtt/K3U+jwb9s2QJ6VatduGxoE87awVeVfLUrIlYNvyCoED1n/UK7+cs+iUP2u
Rm/qbXv3f+zBCAYYx6CkpilF4FDXYIg5JwTEF/lxTir9z2ItFqDC9l+pbna7KkbivekfX/j8Y0oY
k7Ym+ge/CSHd+IQIKA9rGeRnyd4wMSphMPTcJMz3fur0A30pIanXEcV5KQMjzZBLHXDG+CBG2fGB
Jx5z7qXB4whXoMrJP0WiI3dMA6zHUsJlgIjxVu4f4X2lCjmFRpzy+iooPt29MAKhpsxO3FLMHbAp
+K8UV28q/KUZySkHop+SoW3QRSB8j1/36JdeFT6pmLIMUqHcmtToiRJbiTwcpGGHD10HkhgXMxQl
E4PIbrk8nSvxLcKtIwhzGuAlP3RO8lBCnwEDQSXRyG5ab/QN5szUM0zDSl4xWeKCXM4TYh0+q/Is
fHo2ltz6HIJUET0M303w/LtdCxocXwbKrvoZICSsqDi5YLOVZWqVKy6OIFynmX/NGJOJx9G9Ls9z
tdrN2h8k7LhJPXrd+DTvZs+BS2QXKBZsddqYZ3EciGXipDf23YsxjaecyxQvLwhPD0aJIG0936ek
x51ui3aBNlxZBlk0T5z29Ha4M1biYuEXfEgeVhMDPA779AbsgkBg63vIA4maSKChZn2xpEjkCXQl
9Apg8v0c+MKuGX5gceQPWy2XeYl0CPFdNN748DAKFSRQMzxtFnJ586LgHi7ipk2o5mlX6DD0ToNi
2UzaqkgHvCIYqYJkxNiEk8NNOnDImpxi7e1uP24Jh1cD+AFi8JshfQZ5ZSCi/R40f2adW7PP4MHR
hGPpc0067XptIEULeRi2j524tI94uPW4IjQaTT7IkAjBFP6RKWQ83wECVBEfck2y8PJxpvLTmYK9
2pQGNpNCQnU3EGwIsDW3s1jB+5Ibv0pp4YlbvbVD+JOxLVq9+5dx+C/Kb3sgUjpBn7GkzoTumlgZ
EgNAUFQ2E4SScR1FTv+RFq80Gf75QSDLsM+G9Z92v+RSuBdc6WSGBUwOmIZ1yQxRLUIfzZec2sPr
CREcJaAn4Epal/QEobMSRZCQcg+9QEko52od7l+JMY60dBDY3bMRtsshj6rd5UfYoffrbtUaRnfB
UfLcusnmBT+qODunJQmMVxqWTaph9XgkYWe004zbclB2SplJmK1edVLMTX/V+Z2b2o/EOlrGenpz
qBVrQ7cAnR5UqznFzfRsU+iJs2d3hzgUUlg6qIJxhKO3rsqlK/OLGovTBeU3Eu918oIHN0Mmry/4
5pxzMtbF1S6ce3XpWxUF49htSD9kaGiG3R9uOPAvhishL7+yWjNvaDqJ6H2a4e1aNnVZdElim6xR
iYHme43Qi3UapqssiRvSplayOSSBV5gzpXQ0/uS23VAsyIfOR+oQzg91iyPOCv6dp0eWreCmgR7B
gX3xNn3nw3AjX+Gwmid8BvfxvyQPhzQqR8sOU548GeL/SI88xTx3v5Jq+5vMiI+AJe+l4awn8S3K
4F1GkZewT5JtIogEggBRBY+MlMmyZNBHZvGiuShi83rM1sxQjk+ibLzx8AKLjjTPvWQQf6dpLY75
NJwtCwb9573o9etzdyzOF+8/Atq6vZsJVz2WZcS/0/xYjJTfTbirhKEp5qmW1YQV4DUtg5loKSYu
IbXGWb4ike8DYQbjmJ7TeLl330hEYeX/9BdfvDV+T47dBQeBgStkL+d2DOozVKVL+P2i7ESaZovR
+d1/affuk7QDTCTJdeh+Y3bSEUINLlxxI75gqZEAE2DO2HKgvZV0cBuuXoXQLlgOQmhzmSAL5kqT
YlcTywoZSR7MbMrzP4I3cuCusZEqvz0lz1Gq0EhAYlNvUCY6YiET+qkfOpOgwL+k0+1+LXiNXYnd
tgtXjevxz8CVzn4burmPrMIjGQd29dapwTrx2r4yu9Ck2HMdfRZi4blSZQCoofxDW9pMOpAb2LyN
xQT/rnDT7IwiY+F2LZXfeII6x0ERQUEKabU4O/rqDKsyHmmeHKt1o1mmUGi5Z7jL+Fj1k7QBtY3I
8XRaBHjUz6BezOg/30ICY8yRzagABvLPe7U0AxHRhfAyuQUrTH6MQ1VMicimStwOfL/2Avg3X+pe
3W7zJ0a0pFRj5h9pNrr5+gxbVNYvgrB7Y7Rwwl+X/Q8Dm+HI5PYP7Rm6kUh6ckdvwIVCrNpltLLs
ndkzdWI1g7tZpHu9UXcL+h13m+Za1vO9Gv/JZkKgP52El8P1PnYf+USa+aowglXr4gHjKNl5AJhn
wfvCNo1Hm9wYnKJi+OKuIUtCZB5sqHtXKF7PlxwGAc+UBEHqkQmZ/ylc2z1z1535VwIL4kgsLk9h
am8gcvj82/U3yG7v2WN9QwQu01eWruCDRawZgLz5DPuhNTzxQdjpCzPpjVU/CH9KqSfgO3CVA5pR
E9Iz82zydRmpKCutupwSbHfLAeeDX4aUaaeE8o3MmlxGCqLq7Zud+qyzqqwDdKgab1j55nzr1vUa
tX8c3bdzZULh+32AF4Oaxxuay7lYFFhiBhk83LfvvCXZ6SjkNpSJNcQB17M1Gt2gWSeBJvWs13WC
1A33li8HiSwXeONZRi3M8Z46q9dZDNy3lWvfrUHKSHoplb+GXKPdmkKmN73vUPWV+JG0z2iwm9r7
I3mBV+zSny2W2pz7HaaqdQiBGTkvj9BGp+ATi81d5fU5CoMGOqgufzFtkiANUumDVNZUo45z779E
NohK36NsC+oTB3zsFot7rv3+Foh1zoN4vViQK7DVJ5Pb9Gyg9mkcZVh+GWM7ygaea/XIUQeiLW0x
4dKsH1DHOgm9yPzrQO2YoHqzcDVvemjyeW3PBoSKqHQPO3YOzN896YgaAD20slw3RYuk9TmB/6L+
vMlElCJJsNpORHRz52N/VrYXLJExY77svKIFcpcBb7GsNzONP5CI2qekeu1Qtn3d2FwytWJPJcRS
CHWKpxVgvYvlMqUCu25F0RhtXn4J4Cqeb0KZOVn7ju6etnplJb4ZUjImf9yV5Jrxj17FSyHexITi
klx8qebBxVt6NlwGaHD9ryQsurzobMu6397MzbIbnmN5Oa/O2/sLpQYcBYzdk4St1qLaVuwPWIKn
LsfNsnqv2kAhfbyynFED5isv0qe+Sf9M5i4BV/AnbmsuMAW+kUGJ/Xd1wfjoqJNiiKygffmSMU5j
TOGO8xPfePlndkFkBjNSRmitsmFimFiwQwAUwWPZp27p/0T1hIzkjCtEyz8QsC2P3MEfrmFpJ1lR
CMcg9zLD6WSNc3KgYX+3ieCoKMBOkMh+AvHO8ymE3vgFo2C9/fxtfEkr7/c3nI9YGU5QyUKW8YUO
52RlZL8NuLt5njTf2Xkdy0hD5AVN21mdth/5EnLtY4P5kBZr1Uyx+7lMmjjH8sFE+QNH+UMlOT7G
Z3NzrSYBNh8uO+DN9KP4yM4WwAQZMQxCRJ0IUw7V0loQesyQ1lFV4MTKwRRPJAqlpiXQtZTdG3jJ
fBEFnBKLJ1KCZZJOPDYNYSP8ERdAj2FnabZVvaUhN8Q1WTBEeq2GbqZxm78qLq2zguYwBxruVnr9
5C32I0y7QnjpFihw4auL6YVw6DoAp8FHE99HrTic+T2lLA4or9j0esayxnQeU+sVGEfBof61PPoE
ZBhqCDavWnCRQfsuTOPN5FEvsCoU8RhD3WXQ1PC0SFxSpKAAgoOHAc8dwsPRJH/wUEb4ifCwQx7p
WLDenHr7re9U+VU0AeGn+4oKyFqVxqd8EOT3hGrqTl6MbFzTjQjC+q4IxEnoE2DfR+aEXfAVJWjv
msfO1g0S0sAATDb+fpZqFPSNY/s2nbBsfeC3th3fipR+JmwhcC3mCsBdDALwxLklfkKnOa+76msj
Z24IyWMeuaKzKCbYj2INSpU3fDZEGey4APcBr6vCsHvEf5PwfFW57kejzVKpz3G2EOPWf0Q3r5IJ
MPlZ0WaR6t945fyQUgTkYiCWWdbEe4HIxqN7L51C/z8s2qerqo2OuNmphP9IYW+9Zij6zU4hbyMP
VM6C04gh3pMr7J85qe+/8KimgRMi6grffJlVE98xLnNwBznml43py7A8jdWTxOOdYLqVXrUluUum
JJsVCQYEboT5h98YgD9xa6a2xK+PFsQ7B923U40Y7F2KnC/Z/O0qH/0/XCb9AZQPlOUoc9JfabFD
xlnZ/KdM1diFAkIO2fJDTQAg2kyXDgjL0FqZ2L3LP4FLxFsAjQlRsSGdlb58GvI3tPqVJEAKh70m
kIxnp2H26gyvdX+g4US/u+1hIMh2XUnDFwrZGPF1/8yEyjdqxoO07ojYXv3YhiV3gyBfkJUKSBs4
JM+4H+G5QpElNl4GMtnVs8JBiW3tr6fR1NPuDQnae6EsTMkMkwrQt+kIZLNbQm1ihTK2SAOg8HIf
LEQXS5i88sngtb8f6snxncK8h5IgqX+WzXlBlsmzgzbuWBoTM2AItr30AsMM7NxfEceE+4tPScKQ
zIpesLRaYwEjX93uP2LTGuKGQhQ1cboXfHlI8DFdgcRHocJyNRjHJp1BU2VH0zxWGoCX6hIaTih0
ZoL+JfYA+oKi7Jo8ypTulNc0ppSYCFH1dvKnTzZgRWELzkUG6Wv2yqMBWAAQwdW9yq+VIFWmNRJV
yx33oX/cznG13QbzdpcAuf/wogrhj3jAA7MJASnYfg3fGsSY6G/mpDV0UdHDZxmQFlpGsDeBCmjx
i+CHjbnS7J15NSHcRhNmoJBazeroKBZ/iPlSPZsXeA4I9Eac1ZmLIcTn6Kjr2gVvYhANUQLy7IYe
QNutEmDM9UbOKkHhD5QMzEFDcJgFr7DwZRRN6FSuCOyy6aJWrb6sgLwjPU92kHeisRU5HCLtZ4T+
8gn+RlS/DlcMpD1R0QkV5/HryBuIm99BqhX+8cMmkztRenVtx963mux33Dewfjfkr4fEz+UlsV0Q
GQDUH5ZKScT6AfJG9/NKZhZHP9nfrDx81mTL0pvOyyIS8/P1E4c7qJs8ybAuY83wtuF2P81P0skx
eRDB0/EsfDGzBYLP73qgByTsY/f4NA8wWQaepaq2izqojyx4yYMmj/JFHDszXpS73Mu41q0nsb5L
UvItjRf5MiOrmjEBJdzscOCEcEWK3+MPwSvVbKPkR6fh7lLZM3wuQMzROjG8XrEIEbaEXi2gEI4M
T1DrB5uocU9XxE95d6mcWvwtfDJyDulqOhWDUhc9yQ86OOB++cW0pd4hQoUiOOQtEcwOkA7134wh
yR3QaPrLEchLyeAO0DNnZpglc/Oi3yIGSg3e59NQVkhAhQFr65+bQwCGFkKJVHWtn7Qqu+XWay9j
AeD+w5IJlV/DVKBq1M55ITU3LX0BVPfk5Jjd8xdBCVOzWpiw+rjH9zgAZJ0sPIk6eXMrgOLXnEF9
fnqaJL/PEB0oVs7Kskxv++aPoA/FaQVnvWykjDPFuLLgx7JsO+6WfjF2XU5QKFLwLs8yMiEf+kPm
kRap5BB6ZvbRyLiFRZ608Zo1Sy9r4F0iFpF0u+AeGOe3On5pWkMjgLOD/9tVlNM+8vktH+LCoDR/
riv5ORPTxatqbnX9v+4n9727h+ojjTzbKiaiVzVNBede/z0vw7PgF/iX+zoTWsRSIA5R7c9PJ0Fh
XMPrgtrxGv5iExMsboFXixi3hi/4xxxXkUTFC2vOmqa9H9LfuBje4v4AMeY0VwIvu0DnlesBznex
zC25dQEwRZQINRi7+76sPsnYrqZ3QiWqijnhiyPGY8Mt0Vjhz+U8sgx0cFxLiuljdvUosrZEoa4R
8xDeFGrvS6UkEUEpx0Qr0GlwWAYUWPP4mhEvVWsLzGXAr/LbOJez0mGvBO8n9NgM1dRUh7eWFjI/
8u5hz2r4Gn4/3GXKYDHhZNrMV5fYQa9rpeZvuE9Gw5bCjtfHgNhTqnXdBiGuFl0XSfFKX6hDJ6eU
ooxiRcJI4RmOTTPgPaTAK298rfpqCGQsMDOMPVFyHJwBDH3XngNc2h969gFM6LbGRu4bd9y8OUWH
hsZErmJ6SpjOrUPCRr8oLD7qRwrOcEGh0F7qKAQrCH8+XwdJuX5pQaJETeetOz8w+Mm06HodLecZ
UUE3WGFomq0DICSiuaO0gSnujLbhMia3wtXQKEJHjALL1i7QHZ5hZpJV/t4GzCb0Ecr1j2gVSOQB
dJfYfwXEM2izfuW1GyMKnd9dBJq68932uxIJRboWdAZ1BrovXaUV99aV+DPQFcvN8Gtmx88pqo1e
LLFaAmRV0iPpqKIKJ7fZfh3/T7tkk9sa6yPDipqW1ZJIExoDbCqQmXXkWTrATn4KlUIkDgkPaRrt
YorY0IIjo0OD59NxFvJ9j9qwUBm+j5C1k2dXYuDf2BGznIgqPVNZ1UXczV5xWNv1RRwSxyCboBOX
DkBuXPVKIhVKss6pdVj5jMn+0r+RZdIMT7KHh96l6EXIYbnVqN9Dfbp1mlSA84pyrdDyD3MpSw9l
2uLnnwZncZgtEDjFPCJ+h8r8+fyR5TFlB8Ypv9TbOFBGNWlKZcW9uRsmrIvAiwRreLhHUQzZ/Fqy
dsKD2i2T+1RXn46mx+PLLAfcgdkImhAlVkZxl9bY1QryUDGqlALPcjwP3c5Bxe1FSHH+4QwN6yLZ
lnlgwnaiCNbo0TE9L9us/1sg96pAfLepvG3YmEKBwZ8wKOtZJygNGddRYaQ0bTQS+d4CKAmehy7e
Hf+BX0KSMBX4/R4GYLLSRrSxNV8+gDG1WsKom9re+yRhsm/o51b3vbOG939hQW/yARuOkAGTbUKH
UIPFBUKcRtIDV7oGcdUSzmtdCeUP2m/qq0ztVlMgmcPE/Ewi+Zy/nP1wzk+Owv4L5y0TVxVcGkH9
zP9CYmzEEBxSttRbxzi3CeB5GWMxfFkdByLQm/DFa+VYaZ0hDOIee0CsBMQVnFb5LH578Qp0dMle
2h/0jV9s8HXmHSbpOH0XhtH8KX1ldn/y9zNQrMRpceyjWfGvB0ahUcfOTumP538X7d3F+2/1sLtg
ckd94xwtR44xo/6+R04f0DBSRPuX6bDfP4ABhXuEeqYL5y0XqBeYMOmnx+RZnHyxDq9J/36niv5b
RZ7gyWZjRqpYTe+hh0aEvTc2uAhn+73Jqgqanm81FvlUL/X+qHl7V05ej1oYSaKrTKZFW5lk/y4z
M/WkKcjk18yAJc406wFk6aCYLHismrPg40yGm17onAe999v8wo0KBm8fvO/duzH49VI2Lx7aTDMg
4MoZ2FFo1dWWTRPCAGlTsJuH6MevxVX/bh7uGB6Eb0XUxmEGqrDG2RLqxSBwSGetQh3uLRN1wsnN
sUoQhL26guQ0EDHBn0xyR60NoD89+ot4f1oNJ6DcjXpzh7SpZ1DmhvSac6s6kxdghGV6JY/Xtidj
a3FM8bBu7/0nU3LhbILzP7kIUOzrYGCcafV/4+h58CS3OlhkzJRvcjItSc3Wtr3E2GoP/LlIWOK/
1GHwDNf0dheAEKsKc8ZoVgfFIXON6JUI6hQlWUg3tAZhyBwJ+id4WnuH0hancAAJ/F9QCiNt7Swt
2ehZt64YtzozZF2f3JNny/qgOKhe5vHqU4WRS2QJDdCxtlJzi+oYCPhkd03X+JarNYSsyLaRYCD8
0tLwdsIUVx/iCTM+bFmHVCVg3YNa8V+8Msvr+KyMOXNFif4UnVAjQBPl89RqajAjqVkpTyiKbcZf
G1916Q6E2qoCaZ2WROSCMpASAAILc+8vE34oPzN6daeUQjIx3AmMVcRjWk8g1TpmjGTE4eMQL7IP
odYKO68HlbiggzQt3Y4A1VL0jQhI0Mk3eRcam4YhEtqi4jBQveewE/KCfuun47bD/dqnM8Gf1awS
7Lk0+ih9vPnndP4wztiOZxBjnt1+i2zFo0wy3misaH/NUJhMiF2TuA3/8BT1TqUN7TDvuD4dSPeY
da3IGdU1YouFQce6a1nhaYRRGqiJgqt0vKmdtbT6hMf7IlNPToBnoP9xTtHWa3dq/voKFTitpPu2
0e4S5uZCXWVH8S6SEI3f7vq/Ln01KOALjjTVWF3WbkKgYIZ1A2rr+ZG3bo6b0TY8lmVeolU52Og7
z2aTim/Dm5Nxpp3Lfx94P3dmzTq0D7pVx52cz12nkIBSd+TLa38rFTiXItV5YUo2FK+XC/TCCmPj
oK2ITSrwJ1eXbo27vC3iz9zV3W6qTLXWLOPWjtOQoN4yctXVUejRBP4NI9WAhMif/1Gf0eQ3NweR
jbYdeqEz6NIEGpqoTKI4uMR5t2zcasMqi0JPfX43bFaQlt2mhPuEQYjxFrRLr1QNtG1LpewAfqEH
jaMOAKMbwrmW9paQk27HJ7wX3vb9FI/WtXjbCSp6CaRLDf5YfUZjBd4QPOcOg/E9JVYM0LO/zB8/
FbFJe32B1C7VGZk0ePOBZTcemQVeKkMR2PMT2v8q1C/RCJw3MVKWRKaTkWScTGl3xs8Oxss0Ed1+
ynmrstNGvdPugbQmzhAsFqRRwv6GpVKpHC9y9sAU3Pkd/m7btvLY5FgBGIxnvDJrOCCz9RwsQRG6
rn/0RDkAECLOr27UgrF0oBi3TeN8uTnF9YMUVYE7J6l5tqrpzZ2h3pxpNAcN6s6YfV3mm73Ixpla
Nxvgb16WJ6iEz9mnMydm7u4spAcFX8nrtcGdgyGfiAUj13OMev3ND8Ja7dzjdJrVQJR6lzQlUrZ+
dRoRCghGT5R2CmSvdDydcX0DcdlT1LLhSBo1sWcpSqwDfpOEK3Tub4onlouCii5wWX55Gd8f3wSx
X+6SZBF9Ftf5gAhwuUP6v9Fq84y8HovOTbOhFAdLg93N2lP8cF2xxwjo0R4kMt65+BpGAovN2oQC
57hIW738wh9FCTYNxFW8qLgASlH8qUwMSk1Wlc0IjifsCQPQk2qvAhFfpfSfz76iBhlJYgiTiPZD
GSx09UDSfyx2V6M88EDSuQ/NsKyyMjwYusW6voSHPW+NKaHXlINHrTxHW43BLHL5tenCJedPqWS7
X12DsQ2JchkAdA2tBUGImtcSg8lg6tPHL70tYKLnSOgrThCbrrMDonmon2g/AB7QsA8alPZiOjML
svk0AQdU2cDNZQN/4i8ts6k4GFeihuD6edE3peGIAYzXsUBV5zXBDSA+E26zwCP6Q1skaAZuXoHK
kugPm9eoHkraN+zPJR/jfK8n9f4JBBb7GIlqHZ3Bi+r6Se9aiObMuT+Bdz87GxhAA9HmTxZR0kzh
RL7jLqbCr40Q+Rr9C4mYHQW76SInhFmmt16T2vj61NxEkP1caSApDhTFgT9Z2xoieH8Vbk9lNfqQ
ZI+CZcq3JBVb3KKhHwzayRb10PxXqeNu1dj56gSDU2y8BZQznZ0O1vF/GmPue3b463Df0OeAivlz
03aRy6d2xEkMDwaxjuzie3lAHE/Cia9tQdsSaipxPSwyUQn5l6bAgZSl+Ute44x9Vn+p3+y7Zwr5
WupOZ6mS2YZxIVa/cd2dPfOwtjihCvO/H9g+YY8KvFtPtGp61/cSmPpsI99AHjibP6sgorILyBfL
Bc27j8lhgGBIWBcsaOQ6zhj0ZFPf2I69gDA46kj0OZOqCOqeHstEyecH7x/CbWOFNsEtsZ8xk25t
k/WSC/ocRo+llV0rG8zLhAr+Fqs7BhKS3oV27+QgLt4C6kaE6Gpa1WPhgCa9vo9VUU/RwB6UnMDr
AlQZIxPY/McXTdS3Wxgz6KUE+6tY4ayDyk//0x1JNf2yEFdeuyqJgpP3YKPvgzAkvnuItBrUycGL
5u5ZZt/wH7x1xtvFuAF+Pzg+dcIOWgUQwxZ4cuqhDBqd1bVt5/LI5DLT2lKWsZaYZmP12+W2xVFk
vJPigm+95knibAW8S6MyNG7jPQxfZAZSBU8WJCa1C+wZssfcJnjxsYOB7wnCDgxrsrpd2vG+/baa
akGCvC4B6GcOatcYMuLCAYbHxHXB/a6G+RSHw5dAnKOJioMgBCjCqFLno6bSXGDM3Vbo+amMIBWq
Ii+3wFUHyjP/hDF+PFZ1iBU579D2bEvs+mBN7GHKLphJQAaOPB2fkmOm7EfS2gZ9CMx7+Qo7vxm9
PsTa52SU2/KeQ+p03Is2866GJhmqhfjHcUc4HkZMK8WDKKD+fTPRPSnWPfW+C/wxqGWFn1rUgtJh
HjkF9h3Ng2XIjBXW1t6I8GeXJvN/42Nke2nkKTzE/Jhh3fpz4a6EKxNjI4cVehOiKjoH+cN4KWCK
IzOSKwi05D28g5ktwe1dwpZDbyJYavKUYf0FTPUB9rH46JfdDTQLZNXTH5NCSvWDLmf8F3oB294O
LX8Fh8nxA9jKa7KVl4Q899bk+hHfG9E8yB1v0sfnp8NAR9KtfabnUjg9ugfV5rooGIWT0tfJ4/bu
G/zqNKHOMKYYoV+wA98JrnyeHwoAFdmWPnYmBW3H+pD7XfdSVJwiojTCjibDmYL+3PQl9ye1HXo0
MnS4WXA71zZf11WRgYiqGVwlIF/X8gRwmLXemIrzwvHHjuu8Wp9Pjdkiw75/tdyvRqbHZS7Bdqr5
mOcam1+f5CFFT1cDgcf+ibAfAPfPhTcZqF4/jWkfSsozm2uVMtwhl6vE6DSLpO1Q99tmIono+i+2
YFcEFXsY4LHA9G5hg1mTSRLe3qk6cBG8gubGM/6h9SeBuVNra2N9wrxdWmPPheCEboPCElVbLceN
gF4lZcARDHqsVUoN77bwfwlSXIO3wZFCG0xwTNQ0v5g+tVW/e+hGvu2BQt0Eu4NgvuOl/jBNsmGY
qqIit+hFKzL3az8lj25Wksk6YDtVFmZivZ1Vm7hpOgOoWZYo8H8+VTkBcJrGwey+lG81kZmE3Zop
eO9S7bFULSLIYtca3T9RVdgM+t9ar5DGWx1gexdw0EfAT+4VbDDrs8eqRbLVWzureYjWxuhXm+qu
Sy+fPXqJobDG/kwtYwXBziOrAG84/f76c5pHRDFC18RGMnqaiCNscGN9pMOsQzPF6/m1yoO1RrS8
XKaE/WTj1LOZLkRb1PhTO4vVX4nTilMOIsgTEL2hRzLD97C6wrYeC5n64lDn7RMLzgUGh4m0Ejus
FcpdLhiCPbm/ryne7CGdIzShHySmKYXLK3J7aXl+Sa3dxKRmrZhJN6ZbXZ/iwSHe9PE1+HFGraMM
uVDg2kl3YjIuNtaqj1zY5EXwdc+AXQNQ+kniqIDfUorgGUwTiUU5iMxxKsVjoa43LRRAbDws98BE
PjcOGYTMhRmCjCC7XGBu3viI32wbwCB5yWqWyp3bPZADxBNFYGiLo4V8TE8Pxet8rEeSJwZoQb1S
wPHQLfktgkg0/QhUS0d0Saf9fKlj+BYgXI7/+6sSxrC2eVVPOjLJEVb+cqJ9dkyb0w359f6XxWc0
1ox0j2hvGZkgVahOc9JDYrRMn09xJCEU2Kms9gOwcFaald7ZEPh9ugxegoHqHVs+r1DYzJFWivtL
MnvT/P/1tjAjifowsL8zlWnuDi0TKBqf78K3UaFb0DaiKGjRyjK2Jwimw5xRfkGakYjMrpbH5sD1
6Wb3C/2kG9zayj0HmAERrfxP/uqw4BeyeVZM0ScDh0oQ2P01CRWU3m50f/T7yIh+wwHDXR95x63X
1eAL+WvS82xjUqk7HKFf/7tiGlC4Rbxu1YoVOj5hW2ON5xPlL5P0UKHCHd+yjAMnOtsG0kQ0Yy+Q
hg/UMqf0KdG4cX+5uTXp9qETUl2JVFrpPXB9J7tWkp59H4GkYxbgV0ZdogOAq2CORzzE1xY/VsuZ
MmBw+AtZsLdyX9pR/CiBa/wKDC91XICQlxacAWAr2awScmi6SMPLQYZ53g8LZxbHS2jlusbGSY3S
18rO/8JnGE7dNtGoyA3ppquxl7eLES68S7858TJTUlycS4qMRLZHh4k=

`pragma protect end_protected
////////////////////////////////////////////////////////////////////////////////////////////////////////////


`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-1", key_method="rsa"
`pragma protect key_block
pZhvvXE274Dh9fxV8MKnncyzx5m1BiU6jS9ZB5o465fCSeGNLwwrqNl1THm0QNSmRKth7uCrb1u9
gZIagEIJ1otjDIUaZ30Gvyt3JCc/+6C22hl5ZiHTKVzTRtIVSHl5WOUCdEWhN/RGvV13n1hI9DKO
R/81go3t2CmE/x73fGo=

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Synopsys", key_keyname="SNPS-VCS-RSA-1", key_method="rsa"
`pragma protect key_block
WHaTqwGItFKTOYORlChmgExL2caRMh1Ohj7wzQPWUyaKLU4EDo5jBziIsdukPeAYzTVqF3XbV84H
MvaASdlNXyX79txhbdnU8RH3Y2NRR6LZOxEYVZ6UnQL7LoZe3DLOscWREJg1431sHllAvoGLyHtJ
UFJTyFs+eXCxchwrQKw=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=7056)
`pragma protect data_block
a4F/5OH1VkZ5efm0rXi5N74qnEf7FJWP+FMfmyCT9n2MBhW32JKIeaYHIiYxkYvYlQXF+LygzWh7
6VbehWnMomCFTnpFGx/eJbW60KQmNlLWXEi9Iq8/Xv3gKZLhNaca6c8cf1LiNyFWNrhQT0oiBD/b
C1z7lH1sAN0h+chnFSyxeHBf/nIY+DsORRjE3ks0BPi+tJFwD4nX+cOamE7xUPP+vzXTE4Rfs8rm
UlqBkXvxnatOO2KDxdYudzxrIkEqn49FJn2YITGykIEva2GlzsHj1LgQt23IPu+7uO5URtUR16AQ
kGEXe4XPlyCUwdhASAWJEPK41G5uQ2gKWP7+e4AbtNdZHXQ+bf7U4k224wxZ9TJZ9sCiGpRckf6O
q1MGsBHsxV2Kx3fdh3FekmAEcVqnm6nAlES5soM1rxs5AkN1/SmU/zBKT4x+71pcsuvDmac5DeZE
U28vV2OECAXAhcdac4sd4oimY083apTAby5zt2cBcrWbpJZlOIJBOOSOkhtrj/LU6kZC3dpWyB9h
5A/ox8B2IamLmuirZt2rDHD3oOMPw+IQp0bXZ/pBJ5OLUHtU9patix2h4TgcR5GCczd/I4474haj
SyXj/pPocuDMCjjKnjgQA35A1S6iU8uafaRPWksicePlWBkMz+iezpg4Ciea3dDoaC6mpXtDVCPK
Cn5xOVOtQrvyAMeiKuQJIiki/e+uv/JWQFkfPGoCHUwkxQJctzpj+iIlXoX4YMtsxtRRzpcevhbn
Pc0ti9hU6hIETCBWTM0Vsb2Wb4k+VUyZDqjaOOpzVmxhxVob1kqGrEu7s6niEoTesDSS2XwwpTBj
q1n7xQDFYxvcEpsnhvMkAaQ4a8rNFRpHXahICNJBFTbkMLBmCsbKYGkhDVImrTv4EdZYbs6ThjgU
qwcDDBUg6p8FhAY7pwMj02Wdpezqf/GsIaxR+ykf6nJ7ivvxpQYAIyJUNqD6N1NEgykEpS3hJQuE
eF9zm6xjlP39BLoCD6FWTTdewuhk9tDD0IJB4H8+l9uwMjgzhB6xI82gCLT9tSQzk6Pe5o8YoXSn
mtoMNJUQpoWX4MgcX339GIik1rm9NTOts3Xakmbd2IVtJ7+mXxU1XXK/7I23d6/wsp0ocsIL37PX
NozOhpUdUUGGgjraqpcoGC8sx7VEJkKfgZc6uuc7x7GNfN1NlJdPpWXfCEY9H5a3talcT40avM4M
Um2ubmCXmvuP7li7qwvhvzGICqwJ8StCgR5khn2PhNp/efreOAPDGjV3CbM3YAXIxS6qo8YcWms7
RClt/fpEhOUBOJNoGatyCFPmQMrtmSWrWA8IuhX6R10guN4XtqCp2KHCs6tUPQqdCcEdXm3J0G31
aKzOMpgZlpD4BLaQQOBKX7WP0EQ8U9lzGI/0R/L1pHKXWVnZiQLkrTHLavIvuWmrSqpx0vBlddf4
Mox7WE/w2315pdgu7MuM9RLZezmyAVsDBzG0NJXu3wCvqNChgfD79rEf4CcxJoTy+kGzvpUOtX9x
9caT1XZl6OCx3DxWWyOURbPxHwFLlI6rYw8urTHwMNwaTsllQgUti7vX9knNZA91xqnDJD68aj40
mdSpp1UNZ9w1KjddR1lxBLq9hH4SM4SyCLMoLS0rheIaSX5rz/wZtHq3X+XicbtLT/4dzwFPC0Cn
emuxWMLw/6p9Icm881tlwjEXCuOIvr7uqiEsU14DkAQCfHUlk2rdpZR2rYv3B9zHclM96/Go2KrR
kVR9dqmu36c58o5cubaGi3vsE7uXNbCnqdXbG/kTU807aUcC+a0li63cD21lDSIEpzWHdu8FkZG5
D64xdZBD5HvdoSU8VpuI/jEzYUDlHF+SwTUINl5sj+buGW632X5d56Ho2Wvlz0KmIyzrLg1uVgRO
jZCPZ7aNRyr1VcdBKrCgnztBsYMTXlke51P/oYzdr+JxXYnyUdsimMLyk69cuMxy2XH4mxPpysPZ
dcrNFLkzH207/KXOY1smY6l7qiyMoqUuzW2BaZnN2Swh4g34L5P9osTzTG/xv2OGGg8HzzaIp7sh
3ekSbwyR3fcsvf1gCrp5jStMZDb5RSr2rwIC4Ho0z3wuhc2St17D8qlJcih8qAT3ZXRbUB96AAxX
i0ADoz1bSkvfdI1YAezMAnnKemq25OU3rUsJbGE/CRHKIcRpxGRI3i5k/61k6jjoXsMRHUPWW8To
9zCOUgXLWcJGxf2Ujq6vi+HJvCNLYwKSYywcbkhrrXKJCM36PvThSbCHgxjnpgRHMBqS4WsET4Wi
yuueWy4xpDaZ7CulQMRFVpfwX5zh+X+gSFuoiFJKPJQ2HQQrO9KKZ7mAEUjMwI8B0h/P3p/g0aY4
WxoR0hGUInGy439pvt7ZRrqbaK2Sn6x6fkjAlsn+b5WFlqbR3LreFYt9NWVZpMA2BHCfNqWG/yQ/
ivTopU8WIry9Aefn8UJneADlKblQxQIUWdM8MhkCcP2qpr8bGrSpICowMoe6U33U4izq/1qHsv4l
STeWR7BRnQzY5j0hLhzsv6byg0GdQZIJhoE5aCBDcdUklCWLuo+r/Efh+RR+rfFw0IXFPpi+dGxp
bYMtkbz/gsAFXbKMATzPPecsCanU9DZ/NcdcqZ6koiCUVZfqFTAJX1JHolDARNAlBL94Mev4BWOX
8PCpPuURMHeuhjK6+tIP345iyhCGdiiIKhxBhPvGuy/TcCmddcv3bzmuHaTvvx/QA4lb1NHTQlo4
V94sg/x65uIPMPQwsupoRoyQYKanSfEdcQHFIAsjZcFxtLJBDq7Pmed5UdE88n1lXNtps4fQdfjx
r9iOn0nTXvk050KYXiZXMgqWmneGRRiig4jdn4O0oegaMjgDIw/eYxgApk7fusm6tF5q0CHEiurP
XdKYpjuqDFT0ya+ggOkAUBt8adeCH1JwxCaOBFHSCFmJok4UBXyK0HlIBlQXU1BUGLpk2lfT5ONo
kUEtX6YW5hnb3cjtP8tyKeRaQYiLG+ZvbDTLmPPsWI3Ey+JE/+BrUtQ9e4mGvGoJKSwzdqPldsVb
odake12Yi1BkbVzXMZqg3wTtMNzHQFCItUNr1hjhnWtbOAuMiKpnxi+nz4vAW0dc7QQvWVVwwKSf
lmGPzesLJNc+qWeCmRNTAKEHP9mmSNlqvxtstlI94/9rh2jOa5iqN11TP1PZ0hAuybh/niCYcg0/
Ir2tiWtRAlIO4scvNzqhdjT1HuywMLwtbh0agtTry0K5DcsW4qATC2q15aezKm4mOzVIYAGOKYJ/
snIHMquFINVUKMY1U7Ee/ACVYu2+leuutQjwgeuqpx39I9daUj2D1jFpUjkxk9G0usQHuJoPu766
RGZ069ujEZqONE3GsrrSiNW1JdNLyYCRFlGhghUnuFiW4GlxJi6UDqZRneNxRupRxKyhHNBw4glW
PA+M3wduUCt72bM4FWFJKj8ppNjKnXwmsxK4pqKmV11Y+azhmUB/mqK2/tkdwfPXetmp0RlTilmB
1+ssJx6nCyKL0LtaQqNNbPnCewu9n5GH/kZwZ/6oFh7pF6rW3LPwyAh/f6KGosxPWcuqNttZqaMU
sK8evVECIxw99QjLb2etjSv2AVCb7yziIvWxsDgIHG94YKu/91lLPvnYHVEEk9I55iau4oGCXhvr
uIURw7w4ZmER2j4+RY+DC7JO1WwuKcMmb5wvs9RIgBT1dThIabggcnvXB5nnUfdI766SxlI9ZkHC
yvlvVmFB4CqIR2HWLk/Laqnf8r9I4ceozxd7GSfldEP19akytxsBOH2knKwe/RLkD4Lmo8IHL8p5
9RfEdkeNP6EiTnstIoabFNLIZPUCtnFIctXK+LmUh10it6l/V/KNoKw4/EPKoExxvyVOWBcGMd4s
J9kjDt+INr6NmC+5lm7IwQNp7HSQ0lJpLIy2fS/nIRkPgulIhA6nQTZ6yBe6EiKHvejseOwv+ZJA
h41wM2dLmP3pZOCvEemFmsdXjU4FIgPWH/vP0bEYLH6JTtO+fWcHBKlBbwaNhVnhefLnsTsAOE8T
vq1rFPOlygiNFSPi4JDO4phjh28kiLzIeH3JI0f9kRaQDBbP6n8qrSh4GX4kfZhNd8sjR5AW+UTK
SMxsy5ZHHqGgYv1R9J0CT+bsnw6ZXfHLMHtSe3LO28l007LFNmFqLEEmWCylOIiJgwH9U87HRuEn
laNFTe5pE78LY/b+f076xjRBzZqwvJvh8gacHQmRJ3yW4EpF6G97DaRIxwnmY+PE1lvtd/SQtY7V
YSvqwFbgFQC4KYaj1WgPV/OprezN7n34FVLKsp7ocfvhfokMkNJle2BQ0LyzOi1MtIoqJMfZ4SZL
loU0RoY0XHrYqYQVl5Lrq0N4zNS0vD7ICZFyF9TQbwijs9G3OItTCxHZNKWIMsenzYaeRS75GtZ3
qZSmYoUB2GMggtsvDY2ckNlzfue/oJtvFh5GzgBrl2eAbCTvCAC3TPsFhHZ+gt7vubMgQeRh4ozc
Ht1rgxH+ttsOBVWZr60dAVEmL6heB4wd9xU/Ovw8+wNT2xeOQy3Vg6/ccmNIUAkLp3pqyyeNricT
XEi1ikkCkoFf4qzZ1C/hnm0ZpPfBX0r5khu/NG5G6yteVITshYXc/4mAONhFagEXiydZFP4JEtWA
8Eyt6v8N3Bhy94mRpSnvdOMl5lVQOe4bm052O0gkBuSpzzeQLY0nAWBnwuo2P6yuvwOlQ+musHSx
xATwUHfUXuvbxrWLBBuTWQdKdA5SXdgppOJad0rbBz0qfFkMJcw1U3FSLu/s/jKvzAb0OOOMvzz7
ag7J2DgTE8T8PTiHqvstXxYHf9/PJkhSRmZtCiCiqQ1v1t1L0if4yrQIHtDnddmrH13T0Lq/AXfr
VdLmbKfbc+0krwO1/BsIroghLuC7TN1yStaB+Wm+Q2YEYSB4vBgrbj/ohaLh0fZqb0AVWTgD0Nw2
y56xX+HovU4UhkqPgYen2Mv1NlAcHgdFSwYL2ZhPVb7cOi9oAQyGHXpH1qbbyzdLR3q6Le1gxKwA
KOtv0ylOnjshfhAExGiYWn4lbbj8IpiWdXFDpVI+qWAX11zQMkvisGv/UAPnDD7VnkFksdMb5KAZ
vgHkkJ5LY0XnD4oPP4io5qc68u131zMSD8/avn4OPHpITcddiY8t3v6MY2/w52x44JdD26p358Ae
Zfe7CCuNAHtIfLlTKDOH85L1guDhadsBFKKUnA7XPZenD47Uye5HqBncACWv5mOEN+co5lcUNdAY
r3iRzYJMuuAhFr6HLYRJtxkjnlSZ4YaObCpfLXB61QR9PJYQBYHiDXZ342pz6RtL810abhymu3mY
zqG5P273x11ylifq+96uc4iQpjNgV5TwB9HtkqWPRt4FXrgB+RWwroH++hh8HjxSaT33dYxB4wGl
Yrxct1TVK8LPIZ/yG2/K/CMCK95e6oErZQ+qtuCYiFu0wK3GZZD1fx274Bw50UooG1owGvHuH89D
aJfK1wzoliiZXBREDRAbvU8aBnUZ0i9pujUAisJR7Kbegi7kApfVgtaFnDGsL7E44vuVF6qbNflL
w6mjhzw+X+YZ9NXXr/RlHGQq/TEFtllNfjSRI8Bgunds9df3hX1pwSGbNuHEQ5qheGqqw5MerL4w
ZyazaRa7mtYGDBvCKLNy3a5lVOD6+wb4jbWfzg+STDRhZP6hwDa57xsHeERZkotwdpHiJtqO3EKG
61rKSQNX6KDmP0kZTDUpKXdBm+2gmmNBcijF4hsVmm3M/NtIS03duXodFWbuG4+O/5rHcpMqkzny
VwZNdWvb6IDkSUbcTqztC3JHjE/JcJQonn+cnZccSTp931Kle7VqyYhpmKE6MtK85t2iDyosPyf9
6Jw14TP5KNIwCzkvRZKs6R95RLabLfJJSh0DAkkH1gYOkjQKWDE9ASnGo+Yv56xeFJePIgEN1FI1
nzu43J++v4p40IGev81En8pDj28m8Ii3RPFE+Npay1O1nytPb6VFJDqhTttT5WP32y0FQMnWMYoP
idunUdAMThIutl8lOyaYhvJD1xWLjAhxHO32pWXwBfA5SbQyk+YL8ihcIYQv1NlkSdOpCsm0nQDi
TaBYR0lSho4cA+zRYOiMgQEKecNWGDasSnlX9+hYOteMitnuKkYcSTM5+F1ycqvLKxIB57Szt/VS
LszH7ixSnYU/j4HkON1GNfClmIvOFFUb5kyhsUX0NRaQBkbf16YsKzwpOvGt7qAOZZW1ig5EymEF
BSZ3M010V9rc9t0l2Vmba5Nm0pLFx16feCxH4HOd5SIk4H6ExfakAWQXdXIIEBYxkWrV+Sk3yJi0
AdQQvYjoKf6KcPJ9VUmtZj9kG1jYCvaAAX7Ud9d3o2+HdBhp81t06oUCYTHv74yXmctduP1JpNSd
k7szdWYYNZFGxpnlbk0dn7344FgBOW/NQnwwLiP+RfTmjlU9JU07tUtzV4QASm2DvremBRM2Cj64
sqpVG1ssSK7IFj/43f4aKYHrYtVhPqF8aJlRBQtUepDDK0u3gAIvJFLs6cB0bmNSBmYYZnEHDH9o
SJ10S5lrB2kxUfKuBJSAI+UB3+vtMEYo+LqZ11kZkAILvHIM9gtq6DJ1nbbS1uynTw9yBatgQAC3
7NloAU5wNAGoygJuuG1oBEnx2WQ6ARpFlP4/ytSTwxGR6pLun1ES+tXMc8MffEVr4/CNhD7fkjd2
tkJvtSJTDv1NXjUFmYc9r7A6sMhQ69TO638A6Bk1pGnLvLGJn/PQnhyqOPOo92JZu7zHjcoqHN+E
lkAhzuSC99+e9wfdbtHmQCYcUrhFAvMUk7WmeBsAA8kKCUmjJ6vSxVN0dE3/KRN9YKi6yxSVwikD
TdpOp2AZcj7aTJUC8jncW8DfRPAp8uNBEoTcEYHm2qr0wbxllhunmTUoz+HmRdf37bCRLYu3XXvQ
nYyCR1YjNCpWo+tO/j8gyNS9WsdAf4K24Y6fQkGf6jzYFrYsmX45GnKgPMOgGWk+rQSfvAAemuhq
JreOA79bhZfPIze2Su9gMDjByDHn8EBbfeQ1QnNxv7vWdeQTUgdKFNigVUMlcAS2MZxVvq5S3tly
NGtvfpO+wFrqMpXhZxqgnT3g3aa6x1K4NoGhPd+dfd2kSptMRr2LPKZSk4IAXk9rmed2l71ug+8i
8+W69/u3CMOuk2fWzwLwMVQ9doeaAskqjz7t17K9M7WMz5P8CW0PMDhv02ENfNxdrE25mGyBMZ+z
AHfAV4YOZdch7AR7061FjXX8t64L1OnSTVGA5mmT6nNyzP/MH8AcheIVVecY+/UpvQvn0mghToKs
/nevOd+Jvccl633/KlqEc5FZ90+lrLLzAZ0/gcy+1+Pl4ZV6FwEqT4HZSe5yHqGbsD/ZoZw8MPSQ
xlVjskDvvBrPwT+MMg8vk+Yv2Eb0ZlQHdm3HggaGgotEXuC3XdiOFpctfnl/UMH2gzDNl6NUxNqL
NUBOYreGDKNGisAnvhivyFYUO6sspGDkeDHK0Hlm1OaXHf3tV8AEq2iOc8kMoK/GwJNcdo0BIAWC
Zxk4QGrgBA2um3WyaQfvmLBFzQZMmXTlTSsm68C9K8EyRNELB1atp3Bm73kLTlL36I6EGfrYgOPP
5FzzmA+a/8Rp3QjPHCDg0WwB3m+dkS6XxbI0zCZilD3spttMtFdjjlrTvtdTci+NN4hLPKSRiSnv
I3HeYtZI5ctWJ6Zci3s7CcZibJLA1TX3oppPOGGEk68kN8Eml+9tN44G63z/WMcXB+jnk0eYYyXZ
/POoR3/Oq+G3kJcHyEON0sFOXZP7yC47ac6kpsu7Veh4o89RkygGYDtq2MmmFvkw2VWoetgE5b6T
KFZpwFK9vjcIwweGQpciVr6nns5QzxJTEC/mWVH5J+Ywt5XCRbkUFEl2A5vllYAKDa9flHMfQo9c
1yRzFxj8ldWXteqI3zTfCvlPgeh3MdWmxZbUtQSujGbn6R/yTiW0UL1Gf3EbEyR9JMMPwVSWfyi/
Z8T9AgjabGKqrhwp0Gkk9jre85Rh/aXa4qI5aSgm9DlXbF6fZQNZx2zw3hieR7p9/0BEieaUjxGZ
d3kYS84gzHMK4iOqZ4x/hgbxtCZEuyUj2iapmpoXl+2HiuFz+tNddMOiYpEcje+9YgeMnIusSPcG
MXd5PwNBL46ee4NDfXEEWOS0fHozLRj6n5lVKcPOJnVx0d7OWDTHxx7UqNec00QvSRVh5692krcY
yDtnowOW9SinIPnr8GX8Ehw85BaT+EHDg2qhnQXgCJklPH49k+q8JcDt8nFNVlYHY+DVIFzXcD++
THmFfKVYeJIkrpUgslBB6Bfu3wWW6Jf8G4euKkxYmresDrK9zBQ0o1YFXednjzn9DK+xXS66/Aqt
QsmKAtniFMFgZbT0kTFpfq26e9y2MitE9BGwGHr4cADNnnrGx4gVv9Zi1BCxytjAZkLkvDEw7XHL
ED0hylXSscHPP/9GYHLSanIhlGNRiXOz1MPFXU8HOlOedFlNF1fKMDaJ/nJzTdzXXta90m+ZkIvq
d4OXWzrnrT2/zG+iJEUBHtsV/dypOBUpofgSkKIYGIqzpgq41PIH8JtB4FpLZj1qo0+TzX7Y+MbM
j4TFBxVe5jTW84satmEkq75x7BD3AXb/V0wrAXt1ZPHCzAjTTrSwl4hvGEZhZ0ClPTO742sHzxyv
5tapLPUFQStHjOAFKMjIrDJdtK47/oEmmdHtIsD4hoEbv2n5DVVC2cenvw+3lsmcsm05O4OpkwGL
tt6quOo6B0VzgZjX2iNy5ewvtiT3U+nGy22NclB2T9yfzOh2HtW4wnmi0naMgEKVkiaZeIoRSwHQ
UsF3y5gQewB0jjihgHPHDw+R/gH9/pLXBQGzzRPFnk2HreGgeVOfF8aIaYVNU+XNXdCifUfbuiaV
psHk/SHRGKhaqDG6gPZBx1gh5+Q/cKK+e3WWbDGcmEQ6dfvuMsbM6GG8o4rPZBtEQDfay0BD4uHA
62edaLqjrCUi2EdKf+/oe2whYVkjEOPwqRALw0ciINPC8bPgHK2oaIVdROJx1A/d/M4FSjDHGaZn
5+inNqrq8rNm1M7uDcmnvadKpAg5GTuaWHzeyZvFwuYt+7vAhXovqlk5ICbg403Bi6UD8u1k9PLx
W/PgU53RYh1JzQE3aBCmTDbEBXs6VA4MN7kXIaW7kMync1yTAIHZOTsNVercONzumtRpckEREDOd
RPb6I1pk+fPiX9RBGxB12JMuxtwxt8iLc0BEy4WxoxW7aftSLOeMX378SBl8XsR8LE5BmLCpcJwH
l203BSEEI/t478s8O5o3eNPZC4Ep3sNe2edZOHARTBdkYXyQCAsLbmwbgByUQyqBiQn1jAxoKuu2
+c0/iCJ4pMXTWUcV0K5oXm47FCpqFyWTGywL2gfr8hz4QpwKOrUTvJGnbHp1

`pragma protect end_protected
////////////////////////////////////////////////////////////////////////////////////////////////////////////


`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-1", key_method="rsa"
`pragma protect key_block
XF1x53/U06/1bd88EIerWO7hHedcd7Qh6/izaG0ralUp/wwhTUTDNmrpTtKak8RE/pjVdj1lY9lF
gSM8/Yu0LvLDbNrFBUWihO3qHmXpfxCIrAxcfyL+YChDPy3jUWgsTBx9Mum+QXr/fdgvc4/NvzET
uJoxxE4RAO7roLLIw1w=

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Synopsys", key_keyname="SNPS-VCS-RSA-1", key_method="rsa"
`pragma protect key_block
ceOcqDuViZ/DSDOdRcGKe9B/T47xyhT7wnsMit9Q2GAgesPPaUqDfduplGVzSnFI8nJQ6e9T+7uY
f5GG7PIIZDujHa3kAPkauWX1RsgtFmnoKWxLvQq6jhYaPqC/zYkDC4/E26t4XkXdLV/Ub2sIAi6z
tVxZz71PQCaMUQQgfEM=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=7664)
`pragma protect data_block
EYFDKCnB0FTqvbXjvQF3lL7FvQI/1A3J4eP+U177tzFcfOgg0uuta1Fj4yPeT11fBV7XUgaqqFm5
0qczHxjvpVnWprWstBOqgWR+R4njlkDOSt76c31my7j/vFgS+6+tsBK/DAilDdZ6YuuX7BfnOuoE
wMUd80O9SMrp2m5SiXZXlb/UmDXQTbRvIOfATSAbwAPrcor/LzipTc2LsDSUanG3K9RnHwhCIEgh
qjUXDAtNEyrGM4x5G2bM4pZZWYHxA0KemSRn2KnuOzrkmNEHGOSsr+IYxBS90YNx0Bsoi331h6JC
Kc4dqokgH0IOaYT7TyHouR/gZvogANZs/lbQgdXBVNLop9S0Tf4k2tFbaaNO/GJss+SeRqqmmsze
U1dzjyLkhvgOgUfTOAzDxSaRE9MEf2+yWHeyWYAt9BHLpAdGp2vDNotwPeLG7XfyxQ76kC14jli4
wjlLynCgbVxLwpw32+AXWpHvErDReQlZd50YwwfkSesrJP7e1RpfjuV8J6gchTef4r1tL43ZUEHo
aTL3WMB0T6NvnobMuanx41CkhA/jhrcIB9buUi0kFu5ZXTmipvMbIivIjh55uik95T6Nd6F6eh2M
CEdbX4GpVm+OEBy65/V9t/qUr8KC2dYfRL3eO94TuiFU6d4JQNMjAtLWXFmlv+0mNazThrj+k87C
b7bE0p5Lr29Lp2bnSwYvJmN42EmvnRTJH5zMDFsVtRG70doRwprZUZcH4wLSsy8+1qu6p1L7gGVB
Heg8pgejJHuN4SnVyQkCbOfT8deEY8t0fYjstA+z5God3ihfotrKHsqWPDB+4sMdCYqZrUM7Wab9
YdFNAXJV5WDPxXhZ/XgNsV5dsr8dsFekqOScea9ZEIFMv1D86mQ8XlOcBs7IcV2tT8mnt0BXrlS8
1Xvx7SPLgFhkymtJHhrCMplpiPr+gTUh/wOoyIsSijVMNhns8wa4NLMpiDIXBuyTGc2mQjYaN/h9
0qeroaQ9dXRQiOlFAy0uw+LEXHjI9ywaRAHhc8cUsR3hwKwVguWFNBXTdc+waKQzqRuZ6UoXSKqh
/yr6NK/9cBx/UAkhcOaUr+pWnLTaTSWS7Xo4u9gg7Tmwk4M6UpC3B+nmEAGvvZ1xbSfer3f74rCR
r2c4uw+VcXDF4Aj/FpCe7POOHSLTrmj4A/cIuORBHGfYEW10ZH/vqGpTpkw1eBlXqHn3eJ12oAf4
IuhSu/eHDBHOBh8pzbtianrFNYUVWbOpmXs2oQXTnGuMOECoTwkfE3pwrDh14IIppGxZ6utlXsiD
r8MiO/ykfokF1URbWZRseIWHXVJhObA5gamP3FP6lsBVevww/EejOjSlKdvdBNbGaUYuoBIc3330
kIRWFHcSGKbD4myobQX+CXWu2XlyzcAxQ46Yt+e//v5ewynpqNJUOS3bcLJdtt9/7ys1+0gDPEw2
QGwSyp0oIhkXMa4WRNHn/3ilfYYDJBpOIsCFWfEL7Vx9krp4oWHQGCvkokg2BKE+uTVsfkuoW2R6
2YEW8sCmO0tYFpdssCh+83eJWFhpbCpB3l/bkYmoR9Rt/fgR/LZvt2/lBfHIwNVWLQCnqAqaAgmd
3XhIPO9gt4bY4BjIccABnvXzFmJCy7UL4Cnq2X1KwLB4b7/e5udVMGGSrToiEWGwyx8hevh6lvA4
iv2kabbVDDLYlaMmqSVB1uRDUwLo2jTrY27PkKK+IFLNhhdmkkEhyTFaAfIqw/0Nfm3zxaM1xSeg
ulIN/LKZYwh2Bcy4IkHbA5z5Yrxok2Acc73NfkZEj3NwBIham3+xTUxU9ie6Z70ho8s/6frwejga
P9oObjBvcDU/F4jYlKnCOEW4UewSz84W5Yd9qgfD49fYb37QP4wpUVA5YwIye8zHJZa+BmXWGobR
fPbIN5FPK59cqsPGXvVm7eDKes4rabPR0mrK3nb2kKgklk4TqBolhy1pYY39k1fvStWUqRtPwCFT
ecVgLgnjcG8dY37byhsqDOHiKEV753sgqaJNYqXG8IrXbS9dlXLMd3NWGIF0Q0wh2UgVg5it4uvo
ZzuuWYvW0n7he+kINS/0wyb2HRH9ZoY7ERVBDKyG0fAwtrLStcSBQMm0WOHy8UiuzPSD9Rferwwy
1KdtwaIQUTNGT0xdBWszA/dHCqXAOY6lEjwkzFh590KwxNlOne+e4eIBUAMRxmIP4m/KDXcIEoGa
sAKSK/+6VW9gbEPeiKzqBJ6EOaAp4fyCvFamyyd3EmC0gMeJ2Ku304s/x91oTAmQK9EDyJUevyaS
grLj2O0AbW/sq2JkwFyJjtWeTwjlDHlICn6GN3PEz4TBo3372HmMQaY1jmK+W8Ps/Zibf1bpQYbn
rpZtuvKRnwd/6lhm8ePgjw/RXrFHN+K3NPXKDT1P/fi/Am3hB7eFCKDnzaPWwtP4HRV5P1zgVpcZ
myTSMC2o/OQGhyKJVsS40ic23oNAwnZNTwglt4XzfXVNfn8enokgS5CUnv5NA7B4Cw0i1fV5qwmm
4LLCjCCJeIHid1jFz6m1qO1e+DS5KvMzTS9JxDPKlLZwSYtrA7P9G9xFNr1y8sSRaDCxWgXplDyd
k/A7lGK0Unw0fTskz72e0eXk3GzbnDSOYUyzY7ZaKmzf5nwbJYTZUQc0E55EJgdQvS0kwZ3UBgLm
c785yiej/K8xVm0u7xY4c5pyDqvaO7Gxvrs79aRJOCyTYVLbIVKlFes2wwssdvLaPJFceNYT0frT
73weWlL73dhGY+hu9t3gnNxNw3iSAWPKg7G6bfMUp9E7PyipNH4wwq0Rk/YDYq9IUiXI56efogyP
RdJWiGZLOH0Yn73K9rE1nWVnVNDZBHaRn3s0GJdHkCamZJ1WTqMW3aTA8qZtRChS7AhphT7DbeTY
/MPh7oVc+A1a07TIKhN828PWa8VnwD4NVUL+84Qy262UkkG+Tuoq1uu3EMBu196ZnJfJt14xuaMA
Lh429AK/5pVfGrx0Psd7Eldg/M3gXaLRWCdiY7PLLmnOqncd4QaD/VmAAPODXOjUnOb4IcJ34kKM
SVS9b7nxJk75TMRtGzSim1e8F04SwL7uEI942JYVFOMM8TxxawLosodUAQESPaissGD87HNgeh1w
hBHX35v/aOKGdUNBlenbmfLgCHOy/GvqIRcFdLr+lh77A1nV4LY88Nay3Po2EEAqTh/nS3i7x2cw
7XV4OcrA9mMmqU+axQB8gTgAzuiF4ZusnH5UGYkdPFhH9z5KO4wRnvfJ3bsMKDbD+qE6xEntabnl
A3qCJDw39zL82Ze8KMHkMOuPWno4KmQ+kce+i1/FFcq9RteviN+qN3HMxs6tV8B3v/qztUgQE6/C
N6blBp5bPmcek48t44v01Ll6iNpqC56gyWplqT+rA7ij3GXEM+SJJBeSHQY0OL+ACJyYqDP18YAw
ZCpN2pTjjkEyq1rMGTFe6PVVUNV/aqWLCNflrbIDn6AK+pEzsXxCegL30uLWGz1QoKDENR228Zf0
SbGKcUsLzxdTGPvqxcFIzbgIO5GQfA8PbGQ4UfrLqvr6qRwWwQEAnFToyUnRAy6hZ7kv4M1Can4L
hCMG5PKib20WVAwSkq66NM/NNCh0wlkNwTPXAczt/U07c6pXv4VUIEuo7nyQ/o0iv9qALV02yffv
Ca1OR/zM+ncViW7ZW/d+orGGhzsdEQ3DnlVeyWvrKofU/fX1VVdIMd05fyCcJNvPAPK2QLP1I3mP
LohUjmwyIrNUWQj68fVlrCXl5o3kRpccx/jtFFN/UUga1I5JCfHaGK7A7nTAOmh0gIhumJPeFAfy
87Lg8+eoNJp2ednRbesOobe30wYj8px6XP5wjuYp2AwLkfggfPGFhXLsVCKEcWQDe5KOjrQt4WBx
wZ+QxgVL0dol49mYauRWGZY5Oor2m8R/E2kLsffQ4oO3lsOWVMZiuxc6eQ6T9FMUiN1PQRMr1p4/
cSwuyw+kmkBXUxKOr04z95akhhYmAbeLq6/MDScri9u/SD8BNC4H4KlVUqvD1/RDYNrAZoZLMtVT
FfzvwwwCqBbdl6s8lH0O8KHlyiYST5wO5W0JuvJVn3TmYoxdb8X33SoCRjxN9PVYQ+UE0aOZhi8D
WizQzIzQsearmR8Z/cOD6FFoM6t6TFJtAIzaytlO6zIlWpN6/YuUXEBAfbG6X1LfHl+YWMeOFoBC
XzOWktJqcqkHQ7OVxsVM4ZcxuGDH1gfDI1s2yrWzi8W2+C6p1VXDtkjW4VSgVwPnY/+fHkb6F/XJ
mV4l8KJzQxSld0nW3qu+isMhst29tZu614rdWFMWqHOfBYaEDMu8HlekmhsUTKSiOO0RPSiQrvdz
ceiR9I1uW6YYM0SKBLC1PJNa13dDKpSotarIiwkOHZmjatH++2EGPFKviBvucU4hxsCjHr9hvvF0
cDdnCSSFnMrPrGeZkiWkxpLP/y7ZQ69sH+G5feCBlw0LT+f8Xxif0riwWGk6hdaOxVEndy+BBota
wSFFYqAkweW5FqAw0dR8AU8ya3I1uvP+hdw3F781N83wlWL130tf7E/jYXPhVzldLOhkFbU2sjoe
RPmBxvqttGKdiaxvUmLD0A6gw2j+fSnPjoxA/JOI8Da7JqEMUGUrfoVidCKMcezyPIdsk+o8HYu8
XmgQwbSJE1GVQbBcYdM2Dr4cRlNsXjDfPRHf1EMGHEwnQIn/i0W9DdcdXYkLUa53rg+sS8ZHX5ri
JqpMJqm71vouLWCaueRCHhldR4GelKgTpGRzDURS1Rd/alfBbPaoMHC1Ep5Yk8TiBCwNjJjbeTKA
B+kZKMTAjRDpwyVEs1DeLc4/jUcHzoZiiLGIupreX0WH1/onIlbwNGTZGfHfAjUmXHh7i78MWNdt
JuPGhX4xhDK5d9IKtGwbfd6zQagYRtGjT8ADVLBMJG+zjBksPnzJO1XvTBn6+6B0h3Is58mEeQwZ
Le+atHfKKLR0ORhC58alPXu8DJY4qlbP5YKwsWAllDnMh207kDQ9TSLui3AzaBDeIftnNZDyAO48
h8/Ywb8QKWsWMdHSUk8MYAoWJ3zDiWMFWyu9gheHs0krzNxZbagrBuhZ2jMaehB387iM1oAegD8D
zA68Ft6fpKPJKNKcUPJWJArJ2qJkg9jcH6vJtQKbhdy7MpGBEwpuWpoTGfviDDr36/fedMKHEZYj
htdZUI4IhrxcdoeaJ79AkmGL+5tgPpBLvNIaIwP0G6pWIQX73DwB4C+XCbZElBy/RD5pSDsZqGWG
sv9vQzPZIQb6YDK2VHB1Z0LIi0XEv50je1/EYPf0833KL17zD/GN+hde3t9iJ/ZWLBTthVtvLixG
4HMaVtyVfeWK/LEwv5m2yP7BBaEVLYsmphsWUoaHtmugwPU8wusunS+zdrp93uJtDTeoo1MHlZHe
ijQTdYifqttR7OL3JBeqAlQ0D5kiGXF0EWl0O0PnXbB5uUSl0EY4MaD0rnzbcnc5dO8OvVNOEuOW
Vm6Zndw3BSQYD4IadsTWuG5sklRPAEp129hbEXXobW1yBHZx0GlZ9Egl1me67YmzZLRc1m7QUHE8
PIzhVg+2qMA3th3CBLC9w/sXsmWOdHt7vhl0m7KA2tWlDZ2LO9W8FTEa3NQCInxj93FwdMRptMM4
6gBZ9i/x9ausSgMIYSGg+Z3x+8V/qET5d3uOR1S836Dk/ofPU+LiK+NyPUJaa/N/9vfJ5fbocpfr
vQGsFoMC8aDTxcrTs93ElwL2eJ2ZztVPuaajwD4yperf7Ir3kdeQWCPvZBGOMTYGEI2deLl2WWUZ
Rzq6/ZxQTFICmMllQgeKkqwYBwBjMg99PI7XDRLGR0kwgEd1nrzkzamOm7WtaaLbaFYQHGdJdK9h
2PuGnYI52YFLkgPEDQbJXr/QS6S2VEJo0AJrcibmHYb5JakzdodTwtUask7wqtGFMp5lkGj+2F7W
2Y+nIpZeuYmxpbxwoGducHVN9gbbKiurglmXlbU/epTDJlIQ4uYLE2hobuc+tnapa/tKeRR69ty6
qOI3PuqrdYlNwd0ohrCyTuO0JlAb/iFhgr013NNWfItso00XTUBuhNd6/iyENpYg2RWDxB7eHh97
+iI11sj4xNIXqw26+Ib19WaWAmiAZxQvwkal0Qt0f2Hq/CmMk4dHKC/FVRYTlByuSBpE/aSck7t3
5A02eL+Z0XRYjOmDQQh4J9ASW3Bgb5tgxirHhPdPz3c0pjGAPD242giV8/sByvkwQfFh+cqAjCKB
Myp8CSHwwAdF1SdQniy0rkq+/HILcUQm67idpZQo0O4yJegdY52BbD3ybQnJwX7bsMYed93geZKY
M0X77kZ83q9Gm7gmaaIUQM98AAj4yX249oW83fOfAKvE3gU+btBLCqBMYpuQZF6kVEUgA/z4i1jz
1mrDH0M5ywlmXqN1Qq2gqa4t7KVilsJZnw4vwTD7O5VeKl1z0U+/d+5C0wXqoEaIdgXN1+NkwLhr
wjpOpIYhTkcsOAo9d7OK3495XsKKafy85/ITwLFolC33vwxraH0COpCIUMgJbJ0wkwKr173Llfj2
eCDDxXB9A/eJcsyc47ekSywNiuoPFKVcZZnEiiEk0UfITOvcY+V95iLevMP43SQwZBwS29N0jpLX
zis6uu+1rVHQxF6nA4FbO+CLh1uyfzbD7U/hW1o1s/qQCQCT0Piy0CJout376ZI1AZcqIIb4+EZw
Kj1XF5h0xOOpZ5COZ8kM6Jltg3Rno7C6pC+d/IxP5stsJaEfjlDlmlveiLK9o1P3gxy1A6OMXWjD
sOBLupdA3Wacc9mYN1XqIsQ/csw67msW99D9Ek9UoTPw416+LPq+hTC4xAntHecqcfgF6u4TmpSg
l5Nqjy+Z++zqbd28/2hX7Q+w1S0aDawr8MXMh/INbUWpjT//c4lIxy4BF7BKKu3cV0Iccl0hqX4o
0GANjpQt8KqfRvZeS4cI2YqNPEPYBPRZEYHgO9G1os2hojy2shH6jqqvQhT8I2S5H+b99UMIr+zC
V5FxEzFaGiFbeIFSr2pxroWhHBDtjjIVh8eyDcXvgcRVFyGECHFz2ZhhAOnF5jSkCOeeiKEeeOEp
WVEmch6M2nOVQevHc0lBULtxdDsMPcbMbFCzpciPFPXUrjgaABv9sq3a3YIoWMoXahFg+O+DpNaR
9oE4rgb4CjUg0PiB6D0yr0RdJh/vZE7MOy+0hWB5LOAX/QbcV04fdnSZ3+0XttlKuZmF7w1bDGYf
a73ve7s49n8ZOWp69KCMWWUmsK+NjiO6ntwkCCnFdMdu33x37Uspw4BCq0ZMUSMbedGHDn0KdOrs
3aLjgvoFnyJ4bhcqhV/gt7kB8BPzNkgHDIHkciCxbYSbiqu36kewe3AFYkdBcHoUjBvp6DLZgMVX
pEZLuk+KgcyXdlaIAxsfX6KnaVl3XrF4YmAN7JJZjaZOajVbNb0Snm3Stpk7haw0QPakmU6/7aF0
rNXbdlfPp9C6/uAQyEnDevrg8eReVzBbTBRX2UVlY0YaI9kBCCwnfZXE/iVhjjTESka4zZhMJbbr
DJ3EnVJWwbORf7Agpvlu8a/jjk0HvWbpmFbAqzHnOx/Gs/5liVrvpRbN0R2AovabU1ER/kyuFXkE
VqPSE/rze4Gv23mLBwxToWmudwJJig/g7V7Tfe2LjlGS5Db12L36xob7leT/EwaE1Grgwkz2OXEJ
wIWM1cDKF7Gu5FwAuVzzVhF2TCbYgMg/6IOgU08mmER4Ui1ZFn5tHHMxBqkLvGXBh/XtrRZt1rqx
XHFgoxk2kFXKY+wj7COFBlykKK2FPcDKCpBkgpH4SgM0pGFh/9JcG+FoOra6Wkrbr03vzyJLQ9xM
fbBz/BRnILTz2P3JJWa0/TkQ7ohZIA7P48UhV/BbmtE/EL4zgwTpgEEz9ewAJtmABqiIp7mnxKdB
ubks0wQ+VIvDRPjBNjVtyq6YvNHDN37qAt4AuafKQ+9PYtEZkhdGvi4dG51EPGsF4k/DfxDP1wI+
SmUCrYy+lYnMqYEnSQFZbnkj51F4tgqLpz2LVYFWBEJx5KskGRHl1IDrTcz8AS09WmYV1v/kuOZ+
5mfFlhLA4TvQvSFI6+Tf9RNypGG4SQrAQwSW9z3fIbH8EIgRx/ACWXWOaqDl6kWM7PpBb/QJma9Q
AEP9uhRdYl/xA357SiecUUiVgkTw97xaecAmTz9n8LhBM8gPVTRVb+tWt/1ooq+YF5wZBta57DNi
HDTYCv1be+mUmkhE/0dlfkfyFJm58QLrOJUnPBM7ucjG41RAkTxxq71JJwmhFX+c12B10KvJGKo7
R735C6PkAekX3u4pO7rPmUbmFk8dXNnz9nvxxtg9G8uPudONOyS8IgA5e4PEKelKPj9nXehKwGIJ
2T1Ag4wB/jlQ0d0GUxMmLY+K4Q7BMXhJpEc1N9YU2wFb3P24ShAx8n2J6g3QqbtHTKbP8qY6MDhC
DRbAKZ3ycC5+32RWczm+6TztQyDlfxiK+VPBMtRvk1BH9FvgP0TdOT2toUQBH6MG9II0R/pKOEeG
U8NAcaBKDOuPwPnueci1aVcsnKe9R4wLAjO96LTTxIi108J7V92u3+tbq0lbK/JukFDRk2A3nfAS
MefoTRCttcLQujSA2pcpy+BTdc+38MIMusHWpAJYaD9ZspteM+1AVJTQ+QlBMSWBVh+vQ16cyU9H
WYT2PFrs7/p+fpfbM4KbUZDWH7On4DKqZYC9KcUtRGAzTuwXvydkn4PaMsF7kOzWFQBYDRz2pjuF
p5SAHpCKnfYgmHt5eRQydW/auaOqkY+mX4dR1UHV7nWgTqAB/JzPTO+sXoOcnhfoswvGm/7ha5X6
5bQvCwep71Pz1MzXJwhbxKTAEYNVvqDNZx4shAWRAfQQzpOzr8mbv227XZu9Bfy6Scrd1N8VqoBw
vYOEjAoXn20vFAJfPd0yuLT5SKUTh5r1dbPAmexJycd2Hmyh66pvOVfPtaKEtiGwGNm5SqTGY5HS
cJtDxyfF4ZpJ7s9E3mXDPohtYMIA44ms+5mJ1p0uR3fsNomfnFOEsqDIMb0mX27FkfxT/lnj/gyv
/YL8dBZI/9WI0hfAsATIO/TkTVEZSGSlWexQUZrf4q9/z12w9aA/QQPnsPk/yeloiJh37VAbcrYA
12283URWmnl/c/ZBjUEh1Ogz1SdaOww+eGI0HlWfH/BAiCO1SvghTizuU4uBTdwf/EaRWgZls40l
b7auJWu/NMpaWgDc2COplRIGvRcCp9p0LwSNG0KENHvUnvfUAjHZyAPe/eTyz0wIBjqhcpnRMQUT
KlEfEY+kI2/iUT9wJXl3oTt/97IiDDaGbz63BzeL8gfZFuy2ivzDbup+5Za6rlD51iE/GkfDJ+lD
LC2UnTf6nMb1kstrG/6ejJV9LPYC/5tijkHK07mBO29s4eW9+TT0Iraf5ztbjiHCFz7ByoST8jrQ
YZgTRpyK7XOOA9h/eFaktqsA6EL/RDSHr7uCjvfIzeWV4WNilKo3+3pbDeyI9dNCVTrEjbbrUp4e
MoQYomr2D1vMACXuykeI8OTRuUcidmCpwI2eqBW9Ya/cPe5erenE64EPLK1Xl8Laa+NUOLxFVndD
a4UiH20ZE6gSZDY4wl17WOWPT17l2uVONNqtG2YRTy+J/NYeF4m+mitqTAfbxlQpeiduIeQVYZ7Z
qgLdoq4VRpxhhvotLYiRFttScbvQz2+2w7L0RJ3fdXxBrcIoFt5Al+Yvl86mgCYuSQ3DQxwVzbOo
a8tRvxyEowfL/Vn4w10GR2jXncucFqFBkqf67NQ8xG9PTZTJ29ObS78rO7J47UJVki6LK/1YN46j
iuav0GxOzsur8pGvLJxCN1p7HBkOoCAwrwnrPrEfbneWsh0SYiO6pxccczh7waJhurRTlhr9/ov0
XP0fQR0BEQjcncDfB2widcy2zVCfiveWYRgHhQK5993pqAOXtqsstLlSOt7Qc9f8c/Ihda3dWjWr
NnXWZmmOVzZ4leVSaF8/l63wis4eNj4V4M2bvrzdDLM/azwJjskJ8U0btxhwNeQBCGQR06S/tDf2
H/6BokNTiAd1guHk5Nu0oLJ8ZLD73LiA+JevyxX09b37ZTAxrEN3Jbw6D1HKB/vXkSGWIVcs1gZ/
MvoTAVn74HgpyDUTh2Jv8O0S4BxiDcVeTnrpv8U6fzSxKlnZvBgKFuM486Tezh25bNvEqyalcLlJ
6wz/Ys0b6mgsc0btLyWiDOlh//TTlmoSsv8=

`pragma protect end_protected
////////////////////////////////////////////////////////////////////////////////////////////////////////////


`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-1", key_method="rsa"
`pragma protect key_block
XKvMsEObhXCxaQCYged0pxsBPW5WOPVZ3UtuHa3cP+2VojMocgKllSWImURfGZJYE4I6wEz5TssP
QzmLpqMrfYDdgM7AfRYRwudB7P+xINB2wn2MNHAyJylVflXM4y2LEpuK0EJupVCabLK78599A2Ms
PTaoZlNJ9EyVEVdpt64=

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Synopsys", key_keyname="SNPS-VCS-RSA-1", key_method="rsa"
`pragma protect key_block
bmjn9NEtNwVJC5+uWEBZguLiQvlhuPetz3wNUvOGiNGc/UtvKvbbGv7vH0EyikYyqSFQNmBAw0Fc
8ktlXz54rIWmlbt12o4hlxcHKwS1ZLgIsdTb1zcz/ll6Xa+rt1lXd6nxbHi5Q5czjtr+p5q7MCvQ
bD+YmU6GASOn0rihqqs=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=2176)
`pragma protect data_block
PwtnI4y/xfhUaqvLckH3UOd6ogtB9UWFFi4yp8J0oWCqFCNmZvo+N0eSaEk746reJlec0GYPV/k6
M58HsnWfXwPt1ygfWQlojy/Xp07wrq5Ks1JCD7iNKGnBF7/3a+wyJbQlOKCzBUvdalt0YrwlnegN
0S4TibB9jYuIhD9iucPBuErmzf7ZEf6wbhMHOYBnYfmq6W5wKamn1ObWPhAiFgWHV+u5v+Gz0dq4
bboTCU6OsGRpXVkGVv7Q758IpEZDajPDjzrTAwC4yGQp1ksCSrCD/sgYJd/DDwcQ50TSu1S9gmZG
A6aD7BHqgkiGQ0nE+h3VK58UesgjJBToSinZYci5N35xS4GON1XWYCR4mvAW2BNtJEKzVEN6SXQy
VcgSgbaaOw4Nj/hA8n1VP8kWHTXC+7z4dWSHEw/HQX7aXqI7CHqrjHZVBiOEy/4fqN7qwXORpHB4
npxthqVrri7IRLe2q9fdMPyRjjhrzviRZQ1oF7OQoQ34YjRM5noYXkk5YYG8HQfLemw3mQA17MoJ
QTvN6toOgMMrGO6oqDVCKVsLdx6jjZcsVFFC33RVoKgRySgXpXBiQT3BMgVd0gPEMIXKbC4KxzWv
qzis9pclbrwbn0jcBRKYH3t1ZzIeFKsRmuohM70AWTKtLGfmoH00UNLzeGXSQYw0juh/sUmh+wCr
RkKaf3qqkOClL1ayLttFo3iu7iUyqu9iY8N02+AFpRgJU7131zp/S5G7yR0QHJpXXSHhU5tKl03O
GfG18SqwmqzgoWGtt9rXm2i/vWHzo/5gkKIarl6U/5qYEKBF5Z1MWJ7tCbQXr4N/gQ9UsG3K6ElL
2JpEfgQAbfSNGTE2XdYkLHLo72F3T2sYtDvKhry2SP0AOQD/1pPTjyYl0LmNWpvHqBvRpptqeUaY
KHQ3Xd+bcyRChOYRzqDhh0osmlY9znVMcWZAli+JiHnFDnMYjj1N0Qflg/J9xfYKmuNKjiG8yXB9
aZX9nqVAHbjzDBN4E7wb8b488VRHGIw82Jw+oluzp4/k3GHB6LOL5HnTPik6WrQjt+Aa36iPoggz
L2RuOxgHQTFyY+/78FKRxwWBxX6ibHfT2v5JJ4x2LClV4Dnug1PH8krCOqjRlEz8hBeRO4hn95yo
9ZIB4CDbbbNL8va5Fr3JNh7FtrAnWAM6EOba8RFLTF11GAbt5ksItXNoJig3wxx9r2mID73M2Hxw
uPL+qD9dThbmQy0kR4+YjQGC0vqPZYOpZ66ZC1p/++HChq7BkDNot2eXknsUw8ZBA9ShQt/8E3gy
KEC5apSjcGcFnNcf1CBWrwlHF1zOakvb4EX4i+w7wmjayUbFS19t9sp1etemaWI/un3dFIgPLTrI
fe7M6yXgP1fize+GQRRV9BHqIr8+LeRIdU9YfYMDko2gfSZPi2XchWECYENZN+a0kMJpmT9oYL6X
VNrhqMJ3FvbiMdNr0P/w5wVuNWp3SMZ7UjtyFtS10I2pVhdE76ZA8fcsEulAH1N1D8ZuWvqcv8SJ
RC9tjG9DFlSGB+zeaffkHhR9gJj+V6ds07j4YaUKVc6rk6CROTqIcejcR08y+IctfWR2JhHFXg9c
CUPVVReXUk+ATlGBMxrYcHFW/K3M+d+J8qxVasuP/MYRvr5BNRDiIeICvNlLZ1ToJT3nyewgxpk4
1JiInVYBGj3EW+DO/IJlXKgEhSj0hXDh0YgmefcPznceVunNDM2nzmYZ2tcGdaxbka9YsdGffPwW
wMpDhhJXLo8K9oxuBXjnDsWfargA01+x1BvNxYBMEOQf/wKVU91Q77xkbh1Tq/Uj0fu5KhmCn1v1
5RrTBd5D9YMwosyoEL8EHFz79+kIeuRQYv0do7h9ZKBFgs9KIGTuKmM69JBO2hLj/hC8UnfmpVRv
h3JQICksXYHxPiwmU1D9lox7XiOuz//GObYJAmrU5orT6bWD4M30I7gbC4/cOHZ8oTRjPQ01bpAP
5naqpw5U8GN5ggZQ2fMe9B1MzXSAf0Vo4eAbdOYErA3Bzzasp891lJexRApsDq3gXeIpmo34ppAz
za+9Cx6HSgt9klfcTyUO/wPSyF035u3zqVaFOur/ISKAvt0oLCnDm8ORGU4H8gzJjr3OSeY8E3dW
5CPU2O/jcee5HneerUtcpoADkzrAu3f8BY61fD3VA/T5DPUPkYucbABCH9LbKTHB+xmuAPtphYwX
pAw0qCFZnGAYTLY42TVUx+c7PMnEGU2sTLHaBeD8FfDWrm3R8+RIFvDd+n6J2FwRNttIHZ5CwG1j
SKy3AVTszS2Kh27lfw8tHpgCkoLm4QI8/xDxVUWpktMJMrw7L9IbbFRuj53w3EIoyqt+nxSuE3ga
/DEPzNuWd/J4fTH7bw5NZ23SnOWPFP1ruVLGDIWIku8WnozpeD1nZXx3Mjt+wRzu/izjx18qqnDB
vQ9oyFjXbh5Ak0m/m0Y5tfji9WU2EP2YMHLVQi2/Mgec7bmjP/IqGFBz4LgGTCN6QDqT6ov2V40F
tfcQzPYSNnLj9+FsIJ1S8ClZHpOWYLh3JxQqDQBWT1aCzsDsqnVUCbxdg28YE8AeZLUbrpn1clhC
WcwYKJ021FZCQ+jOstC3bNZhDVkddO1fAEtC52Ri21fZMaCfHloxqGEqA5p5tUvFqkw+Q5qvOeAc
B5Usb19sYKjvC6FJ+VEPdOEq9w+byATKzWRQy3PHaDVcjhkjbUYLqU8HRPhLaRFVZEldfC7axISP
lGp8yPJ8oS6x67tQJv+Yi2woESyTTk0KX2+DDOIwePOTC8sLlq4CUc1cGpDqrIuAoGN7LfhV4Pwq
Y60ZmWHS8cUtjAk3yxjfhD/D94qyLcWufLXVCZhCnB/RGof0D6+iFL/C/7aGw1XvebERpkFuaXLR
sCnBKTgESJdzhg==

`pragma protect end_protected
////////////////////////////////////////////////////////////////////////////////////////////////////////////


`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-1", key_method="rsa"
`pragma protect key_block
fHvAQs1ZxNRwNdljJiGiblmKTKefnn7aw+tKed9I05LdpPoK5dVdslcywSC9ADg1r1DbRlcbP6mQ
3Q7VipoAhajD5PLPp7+AjQQhoIPhOLgYUUK4FupPoa/myaB/6rRaGZ+7U2Tcio9nJ2cctulYEJoN
Le4P5Qer62itlNPiuuo=

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Synopsys", key_keyname="SNPS-VCS-RSA-1", key_method="rsa"
`pragma protect key_block
afr5D6x5CIFkpnVHvT1VNUfxk3XqWu7hzythw2l6cwYG013HrnfyMHJq25V3doIe5ANdHz67sizJ
Auqy3/Ad25ONpbBSHrNJ5heDTzEWhL1CHrXPBcMb3Ea4x/aE/0nxdJ7InlBWTYti8nWK4SszIuLV
cbD6xRxMQ2jgJglCaJg=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=6112)
`pragma protect data_block
xEE12fXHoQn6WTB4SguiK76XW7EMR0D6bbRjH/6FBnrfPNBBb4VLxhYO+VgfrHHjNhZkQ5/AKvrL
/fF75PYoO+yoy5bmNJgRY0WdrApjt8qKqjW7Nhfy3303BWABQB1eroCxjCmarzbpXlvt8RPpxZsR
iu72U30Kdxil+k5quXBwq+mfiaR5HTASeQVsdwQnivxYvgvdz1cx0OBz3UWqsf0NjDO9OU4VuAgB
0pupShw3BLxE3QiY1TNPWrSSqskWGEL4eY3b+LXDWwvEgxFC5JjLH27GTftfPaW4wLv2BrZkg7h2
DWw9dXmeshvMXsVG5oF7PXhY1Xnotdo9t4qPunaBVORCQtp+AaXqwOyibvOBvj63NAd/mF2oHNQT
9WGBUz0X8ZeQZH1ps/zPl8EiuF2nX9h+S4Tl6oO38gdSMZhGbEjH7h0REVLHP2V2j6mWqy5ssvKY
JQYTACyV/OV19k6gdJQisNqQ1dZixtwmFpCfL6au1cRq8T4IJzSMebDdU8xSYIPvY0jstlfWVxc1
2s12uqD5ExWPtIPGWBd7V5zdXzRf1lmYx6IbB/JR1qvDU85sXuImJadeo1NH+/v0rjM4qTBL51ah
YfQ6UvivT4qYwC7JyDNQDdjCg6ySSAqIySuPZ5SyuzHdMQvKReWo21syssCc7M+fmzwzBFRFF+BY
mlkM3wBJjeTmQYEtM7Q1GCAqAiFKcE31ySr9Hif6h+Y3Ff9JsSheJs6UTHU/XdUzOuIVIbCOx1xB
Vv//s0uOlTPZvKd2qTxJRakUqWjN0u55jpy4y2vTVUmaLmEUkqagJO1YYFJEl+dOMpJumlivO4hY
AM30b0ciwDY1781yM/gZpY8Wyga8ykVMuz1ydVk0mcacOA9NoNAhgSnrE4YaV9m357rVmpxG6ile
/swun/tCa22pResLHsH9SvFKLz++DzZKmesY96UIrTS5NLqcY+RoGJkHkOowxOJNl4CyiiF65Edb
3T3t+w/5oafd4HTK5mX52hUFP7AXFo2MBHO0w62wNnlEsgDGYr25lsieB1RtBlcxfWqpdlqZeE8c
F4er3g/J0EG6NTCAOB1vVc4Nn8w6znQ9J61vvmAD8/QHelN7Keg3tMcqRfHfKFyqfvS8gGP+c/wm
czcAZedMqWxTN7BXLuRzMuo4bwaZXGv488Dq62PvapC/FIayj0SxXzvEPFKA5C2AyqLXzjGhKpoD
qvIAz9iTV3Z3rPEIp5CkCJH4r4QEuW2cHeZXqf3WKWRQXxd8hnfdsuPNRiz4eWMHXNpLNM0n02Wp
+clUCkviAfxraorhdj2PubQwIy2VVj76VVIBysTIVCen6vAF6yZUZvbQYkkzX8N/+o0rVeI4TGxh
y4X0W0urUPE1Bby/H08ToSJ/ifG0JlZCk9PCNtlPqXV5P8aEr5uTTSOdNTf1H2iKhabTxQWypH8R
alXJKENmUYhfLrzta8kSpH1SGwWdzZ7pmNR0RaNyrKET7wqZVsO3ZrGvJRLSTbQrenp4jFHQ/pv9
dH+epWq3wdZqVJJXpG+SRphhcMceTXeYh9GKG8OcknneQCXcO0C1FYRipWmpg66gQVPH5NUI3wgE
wYV7F1Jc42ti+GdrxsR1tx+dpuM3FB0ANG5/LmBKP1D3zASiWWgsJYL/2NvoGS5rBiShrRXwTYb5
TtPaXI1l5MZ3ZOW8oCIEugQViwrwQsy+W9DeDb981rwLt8LwpjpCeIoW4Q88eEUFNjQ0Xom6NACp
2kPwe7TUWQ7Hdx/eSw/GJHx7bJqS/ex0t54TBMRwL5fIvgcCe7TlK8K/UdY9INFPQz44xGc4grxY
pl6Xa6mxK8EiPXhAZiclZEQIe5EFI3vA8jr4p09eg3Jlh1i8ZcCsffR97We/d/MUiCtdwmMODFqE
f/VyUgEOv6gzV6wjUQaQobNxCphnlOUOMd0iYGuBsvvSVTZQVt7vkvkI4GW7bPedAvQLkBPuF4Aq
Fsj3NdubJ9H0WPn9T3vBxZbjoVp8ulY+h4tTJ6ll7Mt1+VkEe1tohSlLiAnbMmuOVBcmetfQVs9o
d5EFI6w9igmHqRE6zGvaUmxndhxYeZ/r1ITsQlJepQY7kWuSt8XyjHM0FCJLWqWbj+/Ji6VEzmEr
1/2vXUVBpQxrXSYECDeO9OYgebmdgw9SrXRDZAMW9i3n6QmA9E+UH62X/1OfMLRE6kxtiaDmewB5
BI+XP9+2LIHZips6NIi747wJVXfBBV2q+uMDuN7QbgfYeJjqqC1YixVE7/sYMEifOM+nbtH6HrkL
yNVccVzW44iErNA02gKHgBZJFrcjjrN9WMzDnJ+BFIkjt1Wq6NTuLdWjcFdS6kt3byhUujmKcd9w
mm0iJVjMwvAaK/90IIw0aJa3Ph3r7yt540AaSopIfBlvp5Se4tFofUKBYhOGaOKEkUrTPEUEPrDr
19++uv11CUAC6wt1y2G1Ug8WiLuXoLYL44XWeIvHjT7VzRWk3mXeEPYpG/d21/4M9SOvZmmSMj9n
0UTyIKTOWVS/sYa7iJ514ehgqhVKUIXzRLZh6Wi7AiBxQDgzDqodYJPJ+EM0ZD3IhZzyBIgcj3N5
69FVe7ChZ86MkGhKjvJuh2Ff788Xx7Y80lJitvGVclttPpOB4snXPx4UkVELz+VYwOsYQGbYh7Db
fCZTPIQk1scxtjsGZBl3kKBsxkZj/m7FM9lts5M5I0HfE3yr8JN2PTPRi5iTSOWoB9c3kOiziLR9
sohS/TdxwvwD+T/DcbyCaIuhgEdcSQtrcnylLKRlNegaT7d1jABVhLgt/I9E1DN9OYs4b70wsAwV
8IrFvWycdRQWc4fFpycR8wQ7DcW31MWR0rywmpDM9TRNTzTG6jParj4+y1qc4tUBUhNVfOgGXkFR
Kt3a/77jkXmqLWQ/5NGTW0BBckpm+UfZACXNWscLx+uygcTwQDro+iNOmG4pvLgRoEJVXb+v73yw
ZNsNhpV4HxO7ID4noboMVrgbz4G67ipvQnLo51XGKVcnKmQMzBKgNXnK9uozYdpz212gdCUIlSLZ
eHf9Kd0SX3GcFjC1YkxTdo/ukBh1CHpRF127OnKwNwOaWieK1wZQb0ijaupfSvpPqOAe1q97hUhB
JNgU0HQ4zfbZFl43HErgmnIPK7gc70rsu/sqq8mN16HVP3AGtpM8STl5MQZztYkwK+XdKHoNPg+R
aq2wXPFA4CGmY1V5EXX2AbLlrt3Zd3MZ/rj+0I4id7YqPi1hpI8Ur/Nh+RNSl4Xa6iSI94nCrYBi
jYtqG9ZehwwKaxSJfPejkzj0ccEE1QD2w2nf4DndEhEmF1D3i8D1yn4DDNLDQ0C/nT3U4gbK29Zc
+j+5N8VoRSttEXpHRVA4XPGKtIIBNwJkB+wTDs8Q8wj6yXpWyuKL4t51ksqvaQWTZlNEtrTfHzeT
qrTAjFtc1Dvo1rTfcmSXNAkkbOvi8ULY5f7kscKd12CpL4ILbDr/i0HjERYR+CElxqiF9wqPpJkH
igj34dR+toVgGH0K6ko2soSAU7R5k0hc1B5aT/8P1PvkeYkMsIGS2LVGgy99eAJfjbz09XiVBXs7
kRTWXuAEfUB6W0dKQtZp12e4rDgFTwp1maQQ8AxebmDOHVT7WvCzIF+bcKWEnBeJ2e3Vh9527oGr
w94Mh7BqY87xp3t4EjAEqnpAnnMBIjG6SQf2yOkLY32Qr8xm/99vvul52aMtUxT+f/v7szY0K72r
kt5MnPPmePTydUh/nqEKtl7mL05BV88iB8BuHfetYkdzMs8QCn+35dFJyLQhlnx3/nIwH2D/3D/a
hjBksuix8R4CFM861b6wcF7tdaor41CGcCp5nXOzYUv1QNzHXgfBa6jEXh2oKeWcDQbNfPECHWeE
p8yuIV/1FPjBDo44IxOMvEbRXK5y1oTDnq2DdZ6lH/vtJGNYNyDkU+UmaOnqQeMtpEQPsQTqLkvs
JnD70neKxKRhtAB6+mdhd76QuN9eyRthIm9Gksxaw62Z+oq1nEVqfoKEe75nY6E8lHaqkRmCXGBj
ZhudPl88/9k7SBh0eq3o85srCcMnC3H/70pb0cqrYrRyX9TiC9fmq8lasg4dpX9fVyerMacrGaYO
J0WzoNpY2gKzhp0ZukZ9R4pvSWzR3iW5N3z0TYKHNPIjFadqabuQhLNWdQ1wLvhx1AHIGsMke6H+
SBu2Dhs9w5o5ozxqyRuICWn7azWpfAkUzFYmA4pagpOZRdhexfVUgpxKwJkeTYogGz1fi/J46yyB
5yXpgD+/ErvD682zFRdM7HyOTxIWHgbxrI5G0zMK4lDCKasoufmjN+Kn2kr8GPPdRk2ElA6y9N5T
YTY25BfbVBwRsL9A9j7JGnqUPabvefVRjD8A15iu0pUcPXR/gRcewNdnomRsPEXKSIgKFC9Gz7T/
LqylRUFT9BVi6zPf4KcrgkDqONv84ZrL+JE79gimT0yscd8jFy597Zv8E4DIzRQPL+ob4Ljt1zcW
2TLhiItQ9pIc73qNYQKiE1k2iOGKIWnxnN2FWO3GztjPN13TxXJY9wEeqJZFFQmsvPGvHHvbg+xQ
HBOicBSOtBmZ6Zlouwd0EaZNYwV2kzM1zF1gLB9liLpmrgSRviVBAmP+47BnGYhV4pUVhiERbdMV
hV2X7HHtBNi33rfCV/lCDUVSJfbFOtbefGTSya9cQkqoi6adO4+Xwi4s4Rt1CKLfO6xAsl0c0s8V
dJxmTZbPu/TAbPGRO7N34mxXoMecSVUZVNhReJO0H+WUdl4Rvikv7klCOah66RW6bukIKi5UOBUu
bIZ+ArQBxzRGGq+tAZpTS8y2SgMmadRJ1v41PgtOovk2ycm6bSrGNy6CHE9CerBJ0tFFycmTzCoZ
WcYLCA+9PRxra/1cyOsYT2adRPw+KVrxKhG4KWbnaCgKA1uOXFR4wvnpCQ+yTLOsLkqioI83HI5f
yFR4Haw33U//mUSa05CuXwmN/aiop/8Z3purtHmV37sXpjy/91dfAzRW1AqEWivpkrVfslGEvrVL
7dxFw3KfZD5Q0pZK845I6FkJggsjgOPKGUnAfmG0+kX7wuTPqS3/xfU2xrqZf9pNAbN0cnQkN/l6
HzouRPP8ZIO829m6aElzaM9e2i8iSCjjx2YiLANNZY406gS7QkEPy4qpeDitqEoHEiNT0kzJQDnJ
VSo+REIDCiJUEUPVFVSHivV6URH3bW6CpyBYz2ZXp2OMMhZZRdI5WbX2r8vsOpaYX+MRLJ6sR9eW
CDaAsi3whHhrEe8sqaeS8HJX6vKuoqiYT51aYh4fvUmkdbRLiQB6mSIP0dgUQfjnFGRW8wJEsHDZ
3i4RSIewhuzuhRSGZvMVHUMhs3rcJrkabKUJbaX7Bt+3TNtDMvCcyflcXEjpBVGr+EUY0qWlRwTQ
tpqmRFHkqzDMjq01FbaTY4vMUldLC1sEvm3oywarOo4eqeLjjCVcp09UUgLnXH5BMHtIwG9mXDFn
wSwavcfrqIc0fkkIx7A+O5Xsdpr//vWh61vNUPvwczJ4GIvqSwqX3F36W3tkOlplCYHmtxWN2BFn
iRv5jqEIoA77B0hyFhpgeG7/bNg4FRpv4qZD/OO96JWsTEznDZuZxwHj5g8i7Ra/qCrFLyaOY5rO
KJ0+6PvJS9KIqSKnCsiMiNglRH//Y+GH+fKUr8nvJjzYyR72EMdcgqdPFeaQDJhWsY7AuG4SZ6li
YrgXa/OMgAwY7vjyi9IdF3aGQ/9a051LsoUtbFAmxa27BzlQXcW5nsyw9Px0NInJzYxpQ4YIFk2v
zIs9RgJIC47qHXj4oTt3FqFwuG9NnU6DwzzOgHsOJHaDNOSjab7UHTXFl2fjkL+46FZsyFlqYaHx
uDVdljlCkynWkv75G8Zzkf+dUR2JfYiDIt32yGamnKpKhO9rrjq+w3uHvE5p8SmyYHHxg1uP7kJp
qhhuo7zbwv3MrZtEzqHChUj5XHsIvqD7mbweNgGsBEcDV3YPzBJtK13F5RVfFJv3sTOb1e5pjuDE
e4cFJuaXWJNGW5VmeBSV1XLZyvCDMe84iMLMn9bPucB324KA7oIodVQe8eVa5eRVsUkwRqdt+7XK
zeF/gfjLAHA87jFBdIU/yHiypL1E32mi9/pySsuQAao37LatqOW09+mrWUXikebVvifyENle3awS
8MS8aUhnLppJg1JP3IYDE3zTH89/rima/ltvBvutOiPRPakRY3t1fadiSHRSw4GPHfhSWuJVgkfa
bOQZr3gjN1BFlnRKPMFJPiosPM3E/F4r7JqqzpwEKMXf/NHpgieMDw/dlLif6vWrT2Bs+ykieZN7
/tWy8VrhagpyD+jNhT+4c30cr44WkmGnAw8samitI2PWKNml35t9TOwH50z3xZFKExKyedX+JbBa
Jk9rgJAxp9BtCD8gLSG9afWre4z8yCH3Bj70i8biVVUmGXyvhHC2zuHMUYD5Z+ROokWxtZ4BUF1N
yIF+SL3I8ajn4jlEvyt/OTPiKGCjJ3Kyg+VL5pUprn8l51Mxhygi0KqT3yCWvQRKrTByS85i5Cic
5SDjM3uPHO7o4EP+z/kWuykwYt9Pf9QDwMqWIuSGyA2+3pA4B6Wb5BYtHwLxBc4YCuHp7KMgbaZe
8wx4IOvjqVaASsF+zQakL4D/gA45qdhfa5EYHHZDnNog7fnkpaPJJYo/PB63Vhr1KNRTtwCQGmkH
TXkZvksoi7dhjPSbPJ5Nt60kcHpYhIYPgHSMTjQ0wXqdFRD4r/2wu6mkVocQJvJspo4Jqf6/ZHz0
bY9tf91YDGml1nlYpwp1OnHvj9L3eqssFK2Dk07STSV7BENqhlrbPa2QPtdEwxO7w2HVslnTBRu2
z7M+dN4hIUKLY95PmCzTZydbe0URRwQBj/V8JAMrG4nPqcFHV0vzDU5NwG1PNBpLjpmDzevxGGP2
+SV+74pcrE7bqLw/OT0zGXoU+sfUz0VW8l3qvfcTQKO8RfQORM7bl+EfvAyNKIgtD6JyOZdQpvQQ
bW5PenIEmBUhV6wcUgD9G7R3jnOuZS4D2pu65hcEH2X1uShQQ7VToTaqMgdyyaivZ0YWigber7XL
2HNZi5hP3knO6fZxM/NMinc1ZMpFJWO4og9aKyXCJQFM8YjKh4SZ6neD3nNfSueDJb0FXZk8QpII
eMOL7nLq+1sww1uwD46LYgLMnRLwUthgPBKxx1plfirSHbqe8i0rdW8hfo3aCmC20yrtPgxvGeL7
5suxEl6QHwpAJZn1wPMAofYA0kpjHeiI8wb+M4HbsV9sR/i0165vLL3ER72l9qr4Xfp15I7vBg4T
zbcwkpKk/AZVHiHkk92k2KxChxbZXAZ4gVThZTEFKBIbebhG+Mjr3wyc2h0yK00oTVZ7Gj7iw/F5
lYXVf8VLkHtZpSXVhMd1lJbAU02NkjPoULRQiGHwJEeZ3g5HdjIKsBnkxIOI93OkA5JPKnjuyyPH
fkVPIN94uAGxmdALAUGl4YiXa2kSUqZoozcU0VxKM52A/BGvqjo5ufApWOZI+3Nz8DvJnXHCu1kC
Q5hjRNctTGqJj3ek/SYC6w6SwSsaXyr70LtI+ugaywy2WkUG7r+/6bMherid0o/WwhwE6T4yh3XV
W7NcDjPUIlycEevoFp8Cpbdu3wKHuuyJD4ZMGa93uawiRrlV/im8jpixt7zCskYcaPTyn0A4bGus
sY2JjacGghgQ0/Lh7+ThrpGTMHM84o/2J5h63XCQIEBVuJFjQwj20oCVpq0sr9uTiQJQeMfB0O69
E7cAsmmjtTQY0SIyECwnMz4tT9qUdpp02p6MSp//hPyJkjnddTp3H8+xx2FP8G+C0zwqdhgQ9tnW
3icOrQKdZUaxnoQRtEytI4s+wtieHNhpxFyX0qq+0iH788op8CeFwc0io+6fF9AIgySPpWNF/6a7
ZkXapB24CPEzXlzawduR//IjyFimaQXbAHtocZ1ODa2WDcu/sQOreVO5NzR6rzlAR+c/eTvsSOA6
vjcpegmBTkkyvK1SU2pBGtEl8ZiF8R+LLtv52FfYcaQqS7ONKsZsTELoDg3D+0sDhcknpy5WrqXR
WTbKqgHVtuvKvfuqVyJz8srbreCLc56TmDpg70Tn+2/lO2vzM8VlSCq1CZOLG9GvM20ssf7njPeh
AaWUK7WZ1f7YYfh91Q==

`pragma protect end_protected
////////////////////////////////////////////////////////////////////////////////////////////////////////////


`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-1", key_method="rsa"
`pragma protect key_block
Ri4Vkk5EC0VoSLPDDt48B9w2ILPOnzT8hojbR3HUc3f0DdQXkNrUGOrMp55i7uR4KsIo6NF/NEpR
rjueU/SD12jLABU6yNTiqNalcIr2ldYhnG8K+WyFT9w7A5wfFp5sInRRNIuPUabkP+ancT5DZTEq
2Oj9o5VkICFCZA5M6tc=

`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_keyowner="Synopsys", key_keyname="SNPS-VCS-RSA-1", key_method="rsa"
`pragma protect key_block
3/txWaBoR7MVACedo8p2/hNqGDUkWVaklBDA1NY6Foauvphw5CJTm0CohEu80mRh7aLuxCZaoDuZ
yWXvT/3Yj6wrJcVVwre5RRR45W65fWxNJVzdd5Rti2zhpX+BN+5FMlp2Y3Ga3dkasmu8SfqwlGbF
0IlTamNJJNrMgoO+rlI=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=13344)
`pragma protect data_block
cHv6Z0ZFAOum+6IggIXHurnr/tinj0ZnyyHVwddLNpdelXyMHfpwOWGPmQFSGJEthblSfjFbzw+s
LsO1n+k1MoiylrHgRewjeWLH3PTK6UmkeReSozyDk6ddZ8th1ij7IJg2nscfdhUyl6NtBiIEhD3i
vVuG1eev0IxwckWtWn/H+/ZZYZZTLrnTLpPyZJfnZKJU8POCKlUx5+guSwCt2qCX/l1cnRwoiiMR
sPbk62lFbReUNiSNxZze534jud2u6dQ3YOgkhJjtQvl8g9xRVRmpjQ/+g6ALQt/s1W2MqhsZwidJ
dLx3EQ7D49D5scl/IiqNy2XLOL7cHeX3EPBDv1YURt7xvQkpXqjkP4UIIr/e/klkvT72b8jBZlMD
xZMZkd+5qolG5NiBUxStP5I+OiNowhg38b61LWD+pC2YfM2svF3O9kvdxWVrn8i8jhvkYg6FAOsi
LcE29WQ/C6v/PdfIZEQMuCiA5e6+KP5eH9O2XIF32jwr0dTGOLHC4dYUZm2udEUSqrBgW2fivtvV
H5X6zHXhiGchofCSjBGVNHFy3xEM89guORnyzOSjrESkb72V29HwHlFts9vUP0ngtlrZJZRHnlMG
9LE+iNF6kijYHP5lYAO+iNU9aAzxAWzcR9WHAVa/DDWdkfa5ncsw+LSdllLLQDz5EbN56GTkQfCv
q/M1u/jrkNS5cUoOo6boPzwVbEmf5IaqKcd92H3dKOmbuQgJDzq2z3OJGj59E/cCFUyJ0372ymCT
4WCBFsC8OelhutBF2eiTQSuwF55TjOJ/myXrXIg2FIHk2+nOmOzupf+cnrm7wJ/rYCHISPjnCyf+
xErgK8bUWObOPSs/IiF/kRkb0D8ZC5+21uu4O06FCwGc9mQvkZ7pj0ep31/5rfrySZVtsSbvdCy2
b21ikeXcIAt44gc/GLss1V6Hbg4RCH7hPRfVwIEw8nZXIc4RrVdP/sjkiyGKUbETplMsh9BhYA4d
T3tBChZW2vH9gJZafzng9SdzUjnW+xlhsFmK/7DXW+fQRi/AKoWXYxymRGdHmeQ04poH0zBxrPrQ
jAbALpDipS0FyNhvhlv4ukEs3i/GpnXz6qYUXAV5uKX4M/lzKE7lCt7Q395VHe8Cmp6gmXtX4cqX
x56JfQsKcfo42ug9IpZDezRL6orVV8Y7hqrA5ci7EweYkZiv5vbwbZDIgPyXCNnPbc1WLIPoD/Zr
/pED+PTx4x0BMFyrpz1YZR0/JLKUM9CyDXGOIIU/HMf6+9Neei/4D4yDE+UOWUj6Fom9/022Wxsf
8Hz/KBXKr9GCrVUz2wQvfrzYkPKF/sQNl7ikkF79Qlps103SToAuYhDRSp8vZ2AbrkcEtMuF5spW
23m1584cD9+8kMhi1TPeVtlcTemBsHrQVsmY17ZhCGYGhYGlmzthDB/vnlxWfu+jVSIo2LIw4o0q
QP5xS0eYIMXI3q3CCzm28hAiko/d8kcyRAgdxv1rS1iN6XFAWTUg/BfoIVPp8mzdTmic9cl4y9W3
fK/KZH42z7+QizJWuLSjbGXPVmaL1csLqtoDbEfBHesenDiNSEKYKOcMiR7+0AnVr4TqzwUB1FGV
KCkzjvJCeWO1u5AC7I+tB2YjlY61Wg4LmHnLing85RGO5+4/rHspro7OcMoeGRE0sWqBineaRFxx
aq7WWYNqrdagNlbxDJFbkmoAMNsi/XUZ1KYE0b9XW/MtrFTstUfYouS33G7qfjfeS5BU5k8yddAg
LlMKP1ooQCj0YNmnXK5LS0GGDB9lGuGpcueDVivGP5urYC8EULoL1XvioVKCwMi8u3gVNfMPCPgL
szNAQkXYEqhyH0Ss+cHvvhytkCvZzbNrqHBR41uVT3vXNw5+CdDz0Kgkxy/CB0iE1BUKroEVPtcv
6cSsBfToVDmP7YPbHx4EqN+ov7bYt05gkaZ1RABrwCxjlyBLl1Aawbs3Z6EqTIeI+jFviwrH5Wp2
nWPb+RzsvLYpIiiWRlTc9EIYaMyL/a6m02VO8DZ78jxW8WINEHdxP4o+Z/CWaaHojh8BIsjMqOYT
IeAwEQ53NFCHM87AAog/8Z2T7aQqxon7KWqE0xnvac5XMBv3+kFfKckRE8xDsqcym9v9rF1t9RbJ
bJixQilJu+GMdr0DbcreR4MacZBoD3NGiJrPFTRjTXKyVhAg7qbKC+18lJ/kM504L00dPFvLgPXL
dJ3ohW51dDOL2HDJsUPqr7mKmOT+34k2w8JRFsQFRaOR6GZtPRAn3v25oK2zwTxx+DDD2NkhOI/B
70LksdwIaI4U+l4LZGVwbOECUkbnOaSZbIMV7otZ4VGWreFWtdIYAtlIKE+aB8CXVPpHG33Sr6M5
mvLCy2JDgWXWTuLvPU+3ZAU9JyZYdQHf1UDECkeMzPV1UvZ+l0vMvep0tlMz4U/iYJsDBX4ircwi
Kry3UwL++5zwejlY0R2/9xd8mTa8Uxpf3tF0hakztaA9z+SNJR6pZd9dEV8Rrd+t0SBBIa98r5KY
WNHYXHd3yDSxcZ+6GX1tUD3K/FE1mZ5pFpS67YC01KLYFmJL0ZiiZyhK5LdG8v64FC2enZzt1Eae
5JhR0xL6fIuYueYoBOqKW9+ZBKr5uFBJOS3Ma3TxvUw5Kj7fuTEjNnciFFhoaRTLm/cXNQplnDoK
nvtUE1RnvpkUgqiag49m4bFcLZ3eIASuMNT8hc5HZ3yxuiexk1XFSz+65mbMuNs5WNyOjoEY+jQ9
c+wdnYhvmbeACDMoljp/0yYizezYktpEReev8fejdrRAQ68WJRFWYj1xj4kLH1uEuyuyj0EL2k6V
DSmFVdTZMJQPyAs+OfwCS1dlOfMvzIQh2UHo0F6s2wzpRbn64h2juXeMmCLegqYh+OAEGoL1+RTE
lqePORzMATgXGek5/fpECFB5jDytsyBbp8JwjrHkpUZ/AlqQlJN335awB3vpFSpr7v4zBoJrn45H
YM5jaf8m/2T3Woe0iVIcaAqp/v3DAejC3d1zvTTTR8maZqeF1oOqV4rnUWiE8GZBnSo6F0/xKgNR
BU4sUotFgPtRBFpPP34iOW20FH1G9OSX7zvMgxK1b0o5dnfnWVCfae4CsjEB4SDbIFlmShUZjIPt
Oi1smf8kLyMDA4D7EmOr+oirO01Z0wrAe0GjUeGzbGJDELfN2BIkYi0utHuOUJq0q+VvkOayBMUU
qJI1VBvt1Wehud/A8RS7N98K/TUv/pq3V8xUndOOPAceqtR+1/9lWhenfsBTQbm6eOZCNBTxI+i5
/4rsb0gQZaeoV3WU5iwXIEb7SLTxleLsw/wDk+JGBHy/s+Orwamu9oGMEy9UEXQUMyUeGANPpdDx
eDph3RfzKL5n4EQchwLUO/ZkjK+Tb0uSJgRhX1s8XR36eY0Bifggt2zBnb0BADM4E1xyFZH0tn6Y
N4oLqJ8hrJgNkN1UPqXYRoWdIK9lsQFqSBAgGtAkKQRN+RPojTtJYaPgn7tFAqkDJWi+wJpc/3QK
30GLcn8dfCWipriwwmiVf4txRua0bZRQUXM64/9AMw59BqfRhYT7swTKK5tOD6etL2IUcIAg5/QG
yeVKoNob/gSFsPIYgKH4v63X3x+GGs8IL8eHYx2MBV2EkH5MkInif5NIyQC91/nOPRckn72JYcMz
7PDBLvYnDO+U0xM/0hzKO6uJ1MqtSpRiGEMAxTzOHhDGn7BQuEE4U3z+Hihbw9aaL4aEaR08lqR8
y93j3CUXgGcdUSnfJSdqxKxgLe6Ki+o3O9D6s7ctIDXwLdnqcK2hGJ/WuahdjJsKHDLTLolh0HRe
5u1o7isDPB1zXQZVg/73Pz0+53pLSfjUG7iLBdpvA/DiCFovHXRoG9i8caXnp7yjDVgbQdPi+uXX
aEJACKy30oeDhfKP0+0FgvNSm3yL89Wh26lbVkbPD/dCKI8Dh67pp0AwZPGOOFYMjVMH0vz+y/D5
zAvSZ7RwmNeRbFsMlIChh9jiCnFA5VgmEBCLL/FRo9VZS5F/2FltwlmQKvszrhnp7KHtJZxEUWc0
w8MdznIqspYI9clT+/ZBmhfOnBQYsn4bYIBlfLyThYTcQztoo2o/xe5toZPkU3ywYOIa4qcvi1Nq
NGqjXxdcFsnwL/Wip9jHGaa4JjKPpVSIvE8VrDCLtbXkWWD8IKMYd+m0v10EvyEmP0u54T3nehfB
Bn10qRT6AetV0NKp9YgE5TXDi44KTTndXRmuA09LEB6AiYl0JEfCjk5p5mKVYCPKexnBkAvoUOPp
PSpz7fqAQNPvRkXoCcgb7PSeMTpyfsQDuvy/ePVwigJsuwR6yiY+GbIpc+6dGqZTRoaVZZ4VnXBz
DqfhMtl31tZMO/FXr9VK0gKNdRd/J4sEtHL1MqpOSp4/4NrdEAVFSkMjgjMSyB192qCjtgJpCHuM
KouXH/SIYV3URVEflu2zShLjpUAYsCuRil5IFa1sAmACLWDSJ84MVs0wGnv7kYUmW5M4guytrR58
aoJPGT6D+2D6yzeKFhhOfJElnOuiq/r78ad2BdUp9WAWTmmodrtU0Ma2f4NWSttUIPJ8pAEO5CYX
bja1dX++A8LKT8xfnlrFD6g2rqnxdthzOwzGQZ5MgEUpWtxY75BYTRyxk2JwOA6OYSqA/9riYSkC
COzXVFr+/yE3ePR7x0waUxkA6vpV2wmIvaPYeQ+5LLpI5ish5rh6NwrWQxjjOb23lKzwpVNaUKeX
BWx2PKO8fixn8/3W25zIXhW2CAg7sTDfZjSykW1oKwovIklOmtRHFNc/mAduUYAnbSSrqA5rIm2u
iaV01cjud0jIEodUMpPYzDxjp7CqgYbcs6JMlOtJ8nyYMRKo5x6u+zeyRUumQGtX58sA1LdHA/A1
Mma8YJLMbKZ41syooIPkgJhrDKOrnu4+0sOlvutuZC8rDy2VDoZT8dbIy7Cyq64tWme1oCLeyOX0
Z1VqlrDi8GDsBonrXVhcx+LnaLblnOJXgXWAwOLQw5tSuT4DjYEFiXHJuWVLQCJPURaHvF4wax+S
klk5dsWcO8BDFUBJ6ZyDukMmSYP2syWX25XO26dKdTLud+CI5J2ExP5eAz5mUrKJHN+xdZRwx0n0
QUZraRew/Jmj1/Ze/PxlFIYp5FFGOYSLjDDoVUsNBpvT3Es6xDMfOtjTEt3Ju70/LgD5pBdqjw7j
FlXR9tuRMEID0jHZJV3kThqQrwDpeOG3eyUZiDmQAdmcuHVexgCGRA8fBhUpy+ewakEUVpBzy6jO
WeTeP3gYPnLWOk8GRNuIaAUZXV5KJUmdkdzOB9ySjfu7fyrd1U7p755IRJa+Zksk3Q9PCuTR+2nT
y+y6WpvIdUi/GR5bvzVxw2ZW2Jz9SBhr2QMKu8dIXaVBztEauM8MV1Cq6+7Gb5gGN03phm+1pvid
dt6PSz2hNydCp+j4WMYemrScIhnaGHr1ImaBS4xIsBnCWZJpenKk4FSC0n1d0EmBRj2e2On+l23G
J7UOAoBetv4LZcvi/WKdEvEr+sGruHgZJ0h0dtvo9XNEF5qFDblh6HUxpfuzr/NfYCSWJSH8sER1
Vkx/TVeHKPpea02M4HJPs1kEqIfOqp70g0JnLaW1Jbx4qXc+HI0wKrsvOsPpFcyMmV3oF4Q9MEft
Ktm1EGBZdMVT8s89Res32J+lM427V2iPSkBg4tFwX+su4DNFd9JcLfd+I8VRWS9rZvJIfqCmdXU7
+H8BIB7E8DZ/06JUm5fenFlisv4evZJjBcccie2IV8w3JWs33Ua5+5lIhowUoDooWhAIKXXjio3o
88EZSCfAklw12ZuslNN1c5bXsCwDiZlPU0M++gOvSSZllvk/XskTvdrIwYjmGcq5qlPT+Z5tdjyj
K0xncgE4yw5x3brM57Ekky0sQksTYiCVWLbtYxvf41X9IjN+UO5u04ky1nL2NzFq7+G87+R6b4fL
jNXXJ1aqOdyqcWS+KmUyOy65wkBnQEFV7T8Wx1EGZ98MOZNknnNTFBCns72ITFAXs+QEuH6jHkRC
cBCONZrYk/fe5c7wYAQrIfPotYh4/J0q90L5wJG+rkCjoy/Fj9ey/kKJb2aI1q1mJYMAObdUhpEQ
Jc4TXCcOuY1BZVSPJ/bpp5nxJRyaDu7Vnv9pFWn0uRDb2BvMsj4zLJFSS6ytm3v/2TnjDKza1ib3
1Yrz4K2YaHFnUNa4Y5/cnHhIlfzQYXsqDjOS218QQ1PMb0YOViSLDuFrwCr1uNwzcRx1uMem9K8R
KnF0D2OH1FD6fMuwxm4vQ6j5iBzgZ0Vg4WCdxQl1rFIpx2RbccPrBBqqtdboRO/jWnGD+PbmKjvE
yzqyvpRVneCh2MOnBErGEBgkKOZM2AGIIDU9UyuTufB3bKke7Try6CZLbuHWd4zrRHlHVGh22uYf
crRaGPnl2DpfvbIApd3FSnCEcSVHCj4HfKuNL5tLttN5RlL2yjrb795NLl0CIRfW7W2MVB7+NTDx
vWuK/O3mzWvwExoiov3BzmLyXl19I9lfLwGCGUDfI9tKOJ4R/DJSSrAQC+0aUgfnt04+o33xWmn8
9qx0gGx8U2Zw0R/L7nQDDLHh3TDiap4Q4L4E3QUAynYiy2fcXxIijDRXSbY4uIu2PDs+u2IlVi6l
CxdJPX5pYM3dpCSIYfx9PIWLwEVB5cGB8xFHG6Rhcohv/zcE+V21Pw6zgGXN1MyxiIjZ3yd8jyQa
iS/RGFPACSIIioFiHE7GOMM7yFrT9u9/1EXdkEY+7QbuzwmUJX2RzlrBevb9YG7xZzlEPgDU7EFO
Ns4AOHeN0Yw2viYRqr8Vohsg0aActMwx4U+KjWCbf1IqcBF/xYLtDfizhIHgWclstoEEUBBTFDkD
jM+bfptKsh2q7nEFhgxJfkgX8mronLosE6W9p/17M46890K/B1hKg1stCa5cagqTVUnGx1P1gfrX
GxXmz3Q2BAOLdXjrthsFd0hNt6nCHlAqI0Iy/VS4nB55ojSUDlKYTzg2khNNc6aPdel8y6jnhhpr
A5FGzf7ImvJExYNA3mApjR7bQfGcH2ciRYKsq3BArRbk+DlkNj0GJf45j4xTcN8u2ehiIOput3mr
XW/P8xvAKdkev4NE/cNmuCt/h72JvwVX2OMNaLs7RQ2S0IgnxIodzJQ8xPDYAZY1nDyubl3low80
KDeQkpQgfArt2a21SnqMaMJ2xuU2h3AfgDWDZhjpMYWXTl3KNHj/EyvzAsCKn183u/QsfQbL7P//
hGHhg4vdOP3z3bVieKT1TKIVI6ulXsrsj7F9ZKrcKqG5+/pi8fe31pqyx4kAe6MzBa4//Y0yPulU
8nhMG0RqQfmADxz53BehoboROr2JnOEtnfuij+hviU43bdqtfvz9qim74QHb9pK1mvEk510fbKSX
hm/yvaoUTj3z9q7hfBC5W/BFLmGqjnURn//++e12iBlZAFZyslY+jvGHPBsjdGrswgIDYqthEIt6
SLt34mpD/52ID4ZbHAG/QiSiLRIiMsUOK0vyxPmccKsYnychxPXqWoxripylaGw6saJXBlfgwtaR
vEG1UhdOsbyOBAxrMEj12oqoALA/G3IRBM4tBJUt4fqK5OEzW8SPi7ipjYFN3KSoxLI1K8zlTzWf
KYayBYKSkwseeCxOz4dhfJAgoO/sRZKwBN0f2zlz10qIof0FGLjiq/uneqL5l42ijwoc9YjGO+TX
DKpoxfcHX6qC6rUNiaYAQfECUw2somDdXMa1hOS5H0eV/eOhdN4RGyAHqYf5c87ep77whn7OyK0X
8qFy2DlurXoeEDBDbPYN7DHWqLt0ci6ItqzFBSC3u5y6P0WOC44B+zASawNL2Wi+bJRrEjebET7B
EL6imRQjVDp0gj5jSrhSVBdMkBBTtPwTXv1LXAyye35hCIckAH3sRD7ZbfkLHAbsjbgEcVDXLdNm
AD94fANdYYxe8SJnS0whUeqcrjXWEbMJxYnz26SLDk5k/6hqkfjnKVd65Su1nJZYkiASqO6pYAKm
biZf8gh2XTudXtM1JslOeKA5cjbCdGoiJoDw2tVCLrAbNNyZPURWV8eoAkLWeKAQ5Vaa3QznJjKs
wFslwr2fvRhzJL/DMrgxxFcPR6ehGoBrztXAVCioijGUJPnren1yTHgD9ZqeC8k/PDp/2Qf+ZWK+
yZh7vih4p7Tz5d3Or8eltjt2bGZunYcbSCrv5sbEhv2QKz3JLBWNOJxzozDYecVixYviiNilaMqr
Jh9NjB1IZZI9o/IznY0stjyZbK2MZiNQjG0yc7+XaMkQMMvS3s/HLtKtJ52U0ocV6ubCM4OzsSTw
Ll1d0BJ2vSCrYVa4PaTVXaTBUp0AVJxB2sR9DVizM2oloBTZoBbaw63f3Jw62g8pCE8WaPqsBjj2
xlolX40pBPXbF861beBzGP5W4NJa44ZOXr2tlLkRvueaGncBgUXhDl2D7llAc3+VDpBrUO6xn1QL
VuvEr0QLv5Xc++QkdIAX6Y3Ef8FuuEGqJ70Qx1k9v5E2RYDPkDbpVRlE3NEqIxG0U3/4PjkFZcsp
cOAij+dHYnHaB5ddLY1SQ0CmP5M5GrXPN5YSknq1AP0640Z3GWYsbmY47JZtACK8ZK7G+q+4GYQS
Xi+M81rBSAhDpeAxT/lklhucteLLay4nZgjFret1SFUTDRhb2aF23LPieJz888imG69+mnvKB/NS
sPqhDLP7PHiGeqK57llVik9Q/FiqolVNoIr/EzOPQhfExtoiXGS5joV/LVFOfGfVkorZI2QCfcqj
xkeL27NbzQ+3sOvRZoiLgMpQ8a3c0OBWs1gXBrsrlIjlfLMHEptI5yE0qllDNnVrfTf/ZDDDFlxc
bhftzj8OGW6wrWnoPbIIVBBqGbjSTY7HCpCeViurz8vG1hT5Fe7qNy3jRtQBpTfc4+XlxG/a1zBy
ePjvUWgRWMroa07ZysdOj9orO3He90Bmaxj9H+D86OEcjT8bpBDaL/IztzBx7Na8umIL29jev/Oj
BTT1ADulDs6tnRlmjVXV4t6s9rbV3CmZbOavrKlwimnQWQmCC2egs142FjXh96yVepfqIwqVKsM7
+FI5PHTuwEI9yGNAw2azzzKfWcDd4WQEhBE15+7vQo8MyDRllnsv/PFVb91lfzEto/MHeVOVLrCY
z52Zx4i4NbNCAWGJ+AwP77dQRMTaKI1tswq6+mnCq4ZPqQSSVFh818O5XfEHztT1G1oJs8UfwEfE
A504xIF4AEb4AwAWQ1nJVeHGg/6xtFxI3aaHKZB5sAuWu8h5aSWm10Ig33O98kXugMvRk54od1Q7
V8joMaFBwSLirVRDDv0iHMgFcpymG7L+vsf9iCVObA6RSjJu0T8FlpyXlA1RSm3YtKi34kghU/yJ
p/WPI/v+5JSbBEOOVt5EdScVcITd/TsRCLhlkUOOnich91DcCsS3MUH/79Acs/XitQ7XyJN23Hmx
4Hbbdyz7qXZwfSh2S53uG611VXkPE3HQxZm9HTWD5577E2HAFdiYCeToalo4AgDdYz2fgF3Y9dmu
hYaARSBWqHe7VLdFsbuRFZIUBA0Nux+Jb2PUNENRz/Ff/jGJ+ZZmjb8XCFNhwDORw1fZ4m9DUben
bhVMg/ugL6pSaXlVVscXwGQMPiV+xbpccgyYVywb+NIBTn0lJgaLBX0Oh3dV/Sig2U8lcKy3oJ+N
KCI48lTNDD7Bwtw05PnW7Xfn3ME2yciv6X+MPRF8yMaQepKrMk30i9bF9INzRVbYARvaScofQotD
3LaFahkguz6qFVVRg7BBGq93H4gwTXVE0EdHXnf1tHlCPa4CNgkis6FyfMVyvx88GUHjaMK65AVt
F6zFz582jrB0n/Olic6I5SuBePeAIdBtxmHg10siQZ4i+y/q0mqsjqlO3EtHr2pGJ/maZ8xnSfdt
tQzmLtkK6O1vyUtpYsmVhY+FPbeSpC0VNaZkQSni2SVIbgjzvKVb6y9hDN7ZqhfAQc+rXQwsqXM/
KyHNXueLEjfwZPQn8ia6+fKjWJ2XePkfUMBEguhwphSB9X8StrMrgoBK128kosKCPdMlBD1PBS22
w7sNOjbjTbo/SPIwBwrKGzS7lSTEYUHGJILjJCe26KjA1z3n52kjO7cKb0sGmlutwHFWPLJgQ7Gc
9Ls1wLgtmX7YNfhnNFp2WMdDdOohWV0z9c/hi+ObW8DBOVhb/Bk6i/BQA69fZgPBHDP1/QK5wUih
I73+yi0mtObooU3YWVOGGXoiniqGTAXfbW1QA8naGcPaoo3aKMDls79W0GIFx+mvYEr+Z4m/bfNW
X/uLSIXcjfZtABJnTQgMcIgeCthI0BReGgZu7H9s2zb10L6SPghEGJtEmSxvE25AKRseeWSDilbJ
3qHmYqBDB6NfbOnUW5Yvq2PwQdVzjYPfxERqQAvbRdQwjpCX0o18r0ZgWT3d8KsnoaQ971WRYp2H
lYW0nPHDSFydFSTrTZWbXkNiMPcdzqwtuVr3e/rCY5aec/ZTOurlCsqNuCc3OKRnXE3RZuW22qYs
R8GyGyVdeFQ616FUeQqyxxR5rGZhoAaukf4Q/YeXQYKvTZopBth8tx6RvbZ5ZPaIvZ7fCuO3X86k
i2p6LXV4zdTy4bc8rjkYdZR3PwYTU9Sh+IFLHaF20yyDdBrLM7EUhmz8qWgEgr7Jue9W5E71XHpt
QCCIQdHtUwDVnAmVZcXLo4DwMw0zr52PhK6NWpTwcnRV6aB7tLNNi6gP6eks6PFH45FB7WYIRNch
Fq5BaggG5jPd0kbBWX9Em/uiYBOBTKkY2pNIoNYPPLtA1wwbv9AEhXEhmiNjdL1dAXkQLOiBkQpf
0Nstz6QVQNenz6bKwmRGRiZZAtkXJRX9UfAoP+jJ4neCbOqVd2on3YiLLXSYiHWT1rJ1n/WGusIJ
NA4adpmWarOmJ5TpfO8o4iH+QzU/zTfHkJvP38ZEL+GgLJQYQ6Wb7i3M1sYaDoCfoqzwsprOWiY8
7FpYJ0Q0v74UpXtIxp99gKskLfAOD9Tz8eFQmtqA44HISi9js15hqyjsgkbV+r+ODxp2g6LfXH0i
D/z+O1xA4R44bUtJxgfWJYVxGN3pj7ygFuY6c1/3UMSFE8mXSPfH2Rzi+p5P0cak5COVkVIO5hkd
Yy0g2jW1MOE/2OY3buXfONAp6/XfelyYgdFUPe3aYfbtXNtXyqbjWUGVyFNhvW0k7IUA7w6maJcA
UK9l2MrpPYqGmNGc+e1tEC9bnz+zund4OpF40y3+OPCV3FahR4Gi1ycgFyhlZznjyXBlQckvnqaL
/tILd9wZgTN63hPN/qStyEIO4JXoDCsWWET01M/dXvkfbXOhdKSWhKpCM/5XxxccSVK5OfJeP5Di
Yuk2p6lS/eO4VbTTVUL3awtPZPqgkMdfqKyBEVcmSGGmd9LHE5ewm4FllOSOXsDSX6tIQA40lX6b
NHpRy89RVkri5WOw6LhHE+6nOFqh12Iv2gQLczm5KLKIopG1FEx+F/kQo0KX2UKR5xMsE1hIo0e7
LGyR1x2dX6HfEk5oPPdR15nZF0WNX+tu5TEti+CKYOC++uMHrSlYj26m5rkbvWabnCP0su9xjVat
B9T1t8MHIyJUZaLDa6u76c5Uy/zhzoOPUIopeuv6R+pCK4icRHdgYso+jTwBbFyjRiFYTZehu3XH
Sn8Hhe2LiR+COzPFkbbGsuMoNXt7bzDssrXlgrD7HFtSU18vRBLPPNxgobi9n7VTmNXZmaH8txLM
qnRN4C/2vjgpKvw/ei/bEqhnzy6doagHfxTgys3vI/F9jNZu3eYGEST86fKno0+n4ubrfQvZB1YO
0lQitW5R7KQ5ZujrJPB+e2YBbBtvpPuwrzSnTImmxhmikII7cv9GbIcvRQW6bD8BGmmAGWEP0wuB
Wglhwehux7IoUFkHt48YuYV98pXcvTXjE/TissXiGLcpALC88Dk+cpsMMHSQJ/ZUQcx853JN3lqZ
fzt3jIdZkeo9xFcnG0rvTAs9JaX2mlejflX19yHqkZtsx5NbZ3RbJuAiBJSsdqGrgxEoY7EUbVnD
1pwUcCMmLCJXRPSys19God3f2ciXijp2BPBamEqqWXPOwA5iSUePm0PkuA7oSoscnByyHuweOsRC
HtHtTC/glio/c14qQS50wA3cogCSL4XqA1+w/l++n3FL+TEe9X9vlOP5pfX/3kB0zyGhdgJn+4p+
cKbSXBoXM62mVf3n/JIdHD0Td8Yk0vqlVCNlMCE04yoionGNbRkaoxTj/DTRs0py/0UGmAjfNSIF
QsGcfoE2+hBVUHShMF6WVGv1deel42A8q0ZJNmc96OBW8JAn7SjqPalYP7kaO3IcravXZVzCzVHw
jInx+UlQ00kBFJmNlwdreTK1/5lKC4IOZRsYkXUqneYV9Tiv9CEvSKWob6qWOe0CV7cGnbbVKBAB
CWGjqLkk0oh+NX7Lq10cq+qHcy2GWTUAu+RhttxLM0wXp6jjDtKcIQYh6KVgCxzoucmxgkYjG3qM
bVXWmHN4iEOXT+sGbzHzelMmDdJ2pOHnGPBoFaBG6cVu8zHkqjCGHDiK/dqsJGemy+/HzrpyTOiM
bRZprrG9ZDPRh/ZqpWu+SeN1mTmU1Jc+PXa3q/fxjBOHkqSrca498gNkQZgAlIIIr3EL36uXf/f7
DB/kg+pBuEIsgaekxpGCJapzAYtZAxQME58XYNqqG1ff9LCZcF0iS60X91vphzJY7qOVUeG7wSwV
GiVQkJwm1nzfzMwlslGQCyF0I+zI3szk00h6D5z3iWfIBxJqi5K4QPLX9kiMxVEKI4nas3AWnT7C
WOU6jMS9pqzU4f7+k8UlisO7kizLPahDXMbTSW/m4DQGPF8anVpEssMMFYqgfujIEIQTGWC0orBP
BksqwPJIneTbZToi43Z0FsF8Wx+kA9krr4TamKl8HAPIQM5QYt3+TaWPzv4yzzT4xU1WeCnu3kKX
9fpy9jTkX1oVbynG/EbCXuRy8wm70EzpbTw0xwV8pIzYq/TmSn+EWM3TO8yqoe0ca6CpAfUyUKk2
4spT4ZVPVC8yOCOJqoR5xPWmo0JtB+ZlC0f+qc/6Jw/5wgUHab79avEf3Q+7rd85OvdvXLq4s9Ap
h30MCeh/0ZkCuevFspX3ZRjQ7Lz5s8rL8jQPxOvYvznoL9RjjaGu+ex2klV1jNti37ASoRjLThij
G0q8gT1lpTvxi0EufYrfl1K7G1Y3jhLHqCUtn4cFSvo9DdnHzzfj2wAmrzCtXcl3I0BD4kE4nVaR
mlLP68WEzGvvJ84p/qtiuPNcBq8U28CH/cRTZU8mpQw65UMq3bqNWgIiRI5d2DOnDIJWgQaXKKLv
JKAVdhrwNWO6+mSUKxfOWqNLXI28jVb7sSoEWSxdFmg6OgdBPEPl5UNGfvp6ilv/udiXrZrvwSBS
W7WABInEW+mUO2NmKO4n+0tTGPjWGPJnQh8atfZ8EXHCtQSDyXCSFKVgxt3Uhy2aOex9afEOCZfV
FPrCM1ec31LL17E6ty+Ty/zD8GAH6+7Qy9Z/WGhLBcQG3wWiHxpajo4mwuSCqdIIojOsnUxmVadu
56jBSCs7Q4T/X3n/pRRkwjjY3zryeGKR9imHk6IfVg60t6cPOd5RWi9t+Rd+JmlXRt5d900f7G0p
bNWS49ak8NEqTbyJ0TsrfPkXXMDQkqUv/DZwWLhJZZTXjpOMZmzVKxvbxrwCCtWcoVgrMBtgrrq+
JNEbwNg58xcdJkZ4S5jbo2FrYB8xh4bYBC9RPh1y+NuQNg4v8hx1GzeyUg5FP81STw0vDLeZyTfn
wmZD1RFPkvGPm7/8de85AjUT8OpqCa6eTmQi+PMjM0X57QHoQHiB7Bd1+zCrwswv5b5V/prKXby8
KBRk0jX63/YFqSYEdFlIHekHEgkb+Lyx+CerSNzS6eHqMmm5li0SWgYQLWmU9EXokQ7V0jWqP16o
HhIdPLxQnniBL3vI1KCZ07d6KpfqyQVYkaY94ZnKtnzBh2RbaFtr+tuLaN+W0vDADvR6lPvXTkUM
0KKHKPz8Pu8N4s3woJnZ853nLLYeQJ7g7trXuEAX+S5FRfyruN6yoWx2Tq69/c3GOjCm58VAG3C9
LDCUapCHNXDaAY/i1Mbpxw/zN1BlbpOFIkaHEygF4AqLoAhmKFZZVsZxMUfRVBvEzFOwzXmNVZl4
/zH0wfB+Oo9QEW1T3bUndi4pJMeNveY9l/pKogVevFQWJdeIE6XamZHRnR65Lttppfvm4JEDh52i
63NRLrL4w4CbhflNdXi36J4Rq8Kqhz0VOdndrNAojXmkyhhC8cauLNF4TWJ2Q6pafo0UCLD3i4/m
Qet+8hGu7Ruje8bYmq4LgI+cAWWNajLSU8GFyBkrHV+ZdlLf5mfPdrFTQAplRysSOr5ZKPkk7yS8
5iBthWzpipnzcIoDEt4Gjj0olN/Qkv5dPwD6DxKiUbuFuPYRBHM7pDwJh7PrVAvX6xyYHQ9b4EC9
QL9LOfPOlGgbds8bSjTIMQmIvP7Pp4SvOOyxSRl+rlYV7hDV69/z/IrNhBvgiaa+MHJfBeHfaEza
IY1bfpE5XrMWyjyYxnd72HvTm0mMLCNcxbG9a1iUnuk7/XAPNMSvZaP8g8qI1cG31eTZTc9FI/lY
DyJJRrvlO02tVVL4x3lICuBmQftGPQoLXqW3CMypjqHeowaSyAFH8XMGUgifb5YkbpPPz1JKFoZx
WpDGUZ+uzjEKuAZOL6mfgkT5i4KHQtV7Cl6bMtHE1omes8rIDjS3KbCDWd9R1L3cMDhSd8esIKg/
5PRfozUMJiC9dW7b82hhcFaFLHzwprMY3hw0v+TiT7Y9YErKW4EixmACV93vnrNWxEX1JD4mbGvj
kqUiwRteOiZVkpotRIKzB3mLjcMrW4yMMsBicYpBaMg0V1RfIU8lU5ukOh+6S2eo5MhsdknvQ+yl
Kp/iB2EWXm8t+tMieXHKc0Yrx6Byaun6BmAFWq9/loREIBZY8V4QEBMB2NG3w+QOcI2fqYkldFI/
P+CD0Gwh6xINGlunAI5M2PKYCkf7nOIlJ0iYRAOlItg8HwbY4c+mvr6u+xq1SqbIuEAKDUTEzZJv
1yUVi+ny5oBOuI2m2gBJNAxJ1t9fm4gTh/MZPJxjqCeNYzFP/VNaqu5R/jXkskAMe7PHjllMuduq
LFGMxD/ux4/Hd3tFx5eeQmD1HxG44QgqW+50VOt3I/Gg/aL3jkwMOnEEs6uczuT++TljW3xmjll4
OU0ZKwx6d4sEUECepo8+A2KA6vAhHQB0AdOsFpKFKCQdzDKUqetl4my9BLZVxNgxHi/qEnR6kcg/
kOHNk6KwUr7Ec/UP6HQDWf/9mitCag0BAFxexor4wTwGBef1RuVl7UnUg7573mk784tpKjE146qw
P/8fQS+2NoKYqO1IGRqbDHyIyueHuTFBcBi1iy96U+jQ+xccLyjJnr98XFpuu5zQtjQKyS9NH8f3
HLclGdsD7cUy+Vef0NogJBbl+zj3M0t71ga/Ev5LtIFf7YuY+mNP4Nh9XA5qt6LBYZMfPKjc3xTm
TpBgBXn0/G2Nhs2HRoLYHepGgdQAlhIZ+zvUPMwy1c0uePTlFtZ4YE4rFft+qeMdT+wQ9QlF9V8R
ibDLmuNUenfLTzO46RvDS3u1QEUNYQk0lIP2KL/erHVvJNY23dJ4j6HmL8lx5Bj+TaUlxagCcvVq
BtKMvK5HJGjaKxOocfnuPZnrz0m1Dd1KynCilNiizjz1x3SB7Lcw7E5jvqeD64qVrMvdxmbeGq6m
Yq2VRG7eeJibqVPKebGsIzqmXh4SJU3eG09y0SIPKHh7FEQ/M07Ql9FJOQs0Vo5goePsqBi68zW9
NH0OwRwFcFblEDNWe6QhZT5dII+UFUW2co1d0Oi3l3rIi3id77Ee4mChscmc2ifGAFOegZzU/XXW
x5hk+sjJ9jbsiY+REZsuZwEzwP+m/lRutdQdolrijV+j/zMIx4lHzX7XaAuEXIp2hJN4UlviZ8tP
zRynvHd00CV2welMyoa4RnexbKMsVn7N6pPWmLyDo4jU9Qa6ec0RkUSntK0He84l/zTrTZwsSuzL
GYYAV71eqr+bL02zzTZghuUj+pg6uX74xF1UVzxJb71MQcUqlygRY1jD+3mdS91vjqJBp/7zWQbt
8GTsbP19AuaKDNhA7oNFyWh1bTLUu//gdISmfoEsr7Ee5a40AVugUwDlZU+RsHzWShH9fqdvgzHN
DTxKVaoFTYMLaYedjx+AiBGnjmD1xJ/XqJRd+03ptxaSt7iOf/KwTEbHP+gNLpNXVarfHL0g/II3
VEl01vJR6ghs7cuoo3IeW2CFyA0TryUla+z+aKKU+vcZjh7lLFixgpf0JyRJd2FkOoSwOjsl3lYD
EQiKe95RXgXL1fGUmvXCsY7FMcyrpJqynR4IUdPSfQrqRzuEyM5nqzKWvX/if/pObI0COnzilSYS
PhMuCbCb/QgH3gpHmKON0iXYo6I4LmBj/M7Jclw+JZWscTbENeLFjBZ/oPX8ZKuV9tK+hHRSvK5i
6753vIHYKC6y3GQ3Bmne5bNWnvRWcZiDme8QcWFiwKa7L2lkErFJM8uNpVsfTTMVcPocs41vSREQ
b2p7CdbdVL+C3kuUsziMog5cRrvhosgbOb+WTiYM/jZ5TyWsld+hRjtdQG6w1qko8ANWwO83znSk
Tq7DzGqplHpFUYn3NylYybVLegLCENj6wLmiRoiZciiECgQIEnF+lcI/t8pftcV0LE8mmhrd6dCA
Zlo5D1pKeHTP9wYVXattbQXLZgpNoyRWFzrfrvw81NYt0nc+hfsIcjKy7Y3R4uHvPvA276ktPOC6
DOb2jZOy+z60Kl/ZWS+m869GNkp4+/estSW4z5ZzL7FUFzSntz/4z3rL+Upe3t2WTJFSSpCkXEA9
z1iKYVhEdFcpJn2dcpxd3JkrOEbU/qGC3hmGGnQMXYL2zn/iZy5LjFoNFYZXey2PxsXiesOOv6el
33vB49+KE7K6NVqQC6TDM3ekTch2H2nn44b+f9AdaTnRnhYp/AKF8noM9WmO/P4YajDlzuId56xz
a3OMkQarKWLVnTAnkz0xl0cREd5bcLMwV99TzwxnO1wt0RJUsecNX81hAqmypdp724VLUbN2x1v+
hqTWlFDjQizor3szhS7U82JnGF2gI86n9wZL9+nATyEHx1OyGexwYU1mM4mMfnYsgp4tl9oVsoOK
Gxunj9SdQ5WOSVAx2aFZ2GH/ZbQk63Dfwl6xLNz9Bn1HobW3n8AAabjyM7YCI5cq5ptSaVrYafQh
DdEjaylo8jp6JgYgiLAx6eRfnjOC6VWRsWSIksyRmWn8gMVu3XbGlvD8Rf5WzEvJs2W9RGvHceZO
lRqhCy9+zy4CawXYcg4BzA4Fd0PqRziLfNC8rILR/e8MLtObYvY6D1Roe1kh/nA2Ee/rTq+JeEJQ
XCaBMRmq4pl/pH/PQFhDOiI3Zr+wg031OgAYi2TkDtR93iGDUWBjZs9HPa3RpDzQRsPLMckRFe4A
DiBrXasAYdZgUkwEXa4C1kCEm02yI5Eun9wWnJV/FFrh8ckUAtWdyN0vQzNt3b4qaPy/BasKsJPt
+10GPSSYm0DFLYhSwdi3kw3sGIhjzA7dvpFv4TViykrayVEv/ev/QMZ0BHTNsIRdMsPC7obOcjH5
DfE8yGSGeND6UAMx4WZQ57mOam/p6Y22ZzzPX9Q2z3+TVqCIyfZmXSBVx2Wwse8p0P57qH/9UZim
4JbdA2tCHPIC/g9jfiHEuBMpWAUtUta1QHL6TJg7q/xWwyRZ5+2RInCTGw7a7cpJFwtISZQ1UU1u
tthHWUDb

`pragma protect end_protected
////////////////////////////////////////////////////////////////////////////////////////////////////////////


