







//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library:
// Filename: GTP_IOCLKDELAY.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_IOCLKDELAY
#(
    parameter DELAY_STEP_VALUE  = 8'd0,
    parameter DELAY_STEP_SEL = "PARAMETER" //"PARAMETER"/ "PORT"    ,pgh "PARAMETER"-->1'b1-->delay_step_value    pgl  "PARAMETER"-->1'b0-->delay_step_value
) (
    output CLKOUT,
    output DELAY_OB,
    input  CLKIN,
    input  [7:0] DELAY_STEP,
    input  DIRECTION,
    input  LOAD,
    input  MOVE
);

//synthesis translate_off
reg [7:0] CLK_DLY_UNIT;

initial begin
   CLK_DLY_UNIT = 0;
end

initial 
begin
    if ((DELAY_STEP_SEL == "PARAMETER") || (DELAY_STEP_SEL == "PORT")) begin
    end
    else
    $display ("GTP_IOCLKDELAY error : illegal setting for DELAY_STEP_SEL");
end




wire [7:0] DELAY_STEP_CHOSEN = (DELAY_STEP_SEL == "PORT") ? DELAY_STEP : DELAY_STEP_VALUE;

    always @( LOAD or DELAY_STEP_CHOSEN ) begin
        if (LOAD)
            CLK_DLY_UNIT <= DELAY_STEP_CHOSEN;
    end

    always @(negedge MOVE )
    begin
        if (LOAD)
            CLK_DLY_UNIT <= DELAY_STEP_CHOSEN;
        else if (DIRECTION && (CLK_DLY_UNIT != 8'd0))
            CLK_DLY_UNIT <= CLK_DLY_UNIT - 1;
        else if ((~DIRECTION) && (CLK_DLY_UNIT != 8'd255))
            CLK_DLY_UNIT <= CLK_DLY_UNIT + 1;
    end

assign DELAY_OB = (DIRECTION && (CLK_DLY_UNIT == 8'd0)) || ((~DIRECTION) && (CLK_DLY_UNIT == 8'd255));

wire [255:0] clkdelay_chain;
assign clkdelay_chain[0] = CLKIN;
genvar gen_i;
generate
   for(gen_i=1;gen_i<256;gen_i=gen_i+1) begin
      assign #0.025 clkdelay_chain[gen_i] =  clkdelay_chain[gen_i-1];
   end
endgenerate

assign CLKOUT = clkdelay_chain[CLK_DLY_UNIT];

//synthesis translate_on

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

primitive INT_LUTMUX4_UDP (dout, s1, s0, di3, di2, di1, di0);
    output dout;
    input s1, s0, di3, di2, di1, di0;

    table
    //  s1  s0  di3 di2 di1 di0 : dout
        0   0   ?   ?   ?   0   : 0 ;
        0   0   ?   ?   ?   1   : 1 ;
        0   1   ?   ?   0   ?   : 0 ;
        0   1   ?   ?   1   ?   : 1 ;
        0   x   ?   ?   0   0   : 0 ;
        0   x   ?   ?   1   1   : 1 ;
        1   0   ?   0   ?   ?   : 0 ;
        1   0   ?   1   ?   ?   : 1 ;
        1   1   0   ?   ?   ?   : 0 ;
        1   1   1   ?   ?   ?   : 1 ;
        1   x   0   0   ?   ?   : 0 ;
        1   x   1   1   ?   ?   : 1 ;
        x   0   ?   0   ?   0   : 0 ;
        x   0   ?   1   ?   1   : 1 ;
        x   1   0   ?   0   ?   : 0 ;
        x   1   1   ?   1   ?   : 1 ;
        x   x   0   0   0   0   : 0 ;
        x   x   1   1   1   1   : 1 ;
    endtable

endprimitive





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_PREADD_MULTACC18.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

//P = MAC + (A*(B+C))
`timescale 1 ns / 1 ps

module GTP_PREADD_MULTACC18 #(
    parameter GRS_EN                = "TRUE", //"TRUE"; "FALSE"
    parameter SYNC_RST              = "FALSE", //"TRUE"; "FALSE"
    parameter INREG_EN              = "FALSE",  //"TRUE"; "FALSE"
    parameter PREREG_EN             = "FALSE",  //"TRUE"; "FALSE"
    parameter PIPEREG_EN            = "FALSE",   //"TRUE"; "FALSE"
    parameter ACC_ADDSUB_OP         = 0,
    parameter DYN_ACC_ADDSUB_OP     = 1,     //Select parameter ADDSUB or input ADDSUB
    parameter OVERFLOW_MASK         = 64'h0, //PSIZE = 64 OVERflow setting= 'h10000_0000_0000_0000, bit width = PSIZE
    parameter PATTERN               = 64'h0, //compare pattern
    parameter MASKPAT               = 64'h0, //pattern mask
    parameter ACC_INIT_VALUE        = 64'h0  //ACC_INIT_VALUE value
) (
    output  [63:0] P,
    output  OVER,
    output  UNDER,
    output  EQZ,
    output  EQZM,
    output  EQOM,
    output  EQPAT,
    output  EQPATN,

    input   CE,
    input   RST,
    input   CLK,
    input   [17:0] A,
    input   [17:0] B,
    input   A_SIGNED,
    input   B_SIGNED,
    input   C_SIGNED,
    input   [17:0] C,
    input   PREADDSUB,
    input   ACC_ADDSUB,
    input   RELOAD
);

    wire [63:0] R;

    INT_PREADD_MULTACC #(
        . GRS_EN(GRS_EN),      
        . SYNC_RST(SYNC_RST),    
        . INREG_EN(INREG_EN),    
        . PREREG_EN(PREREG_EN),    
        . PIPEREG_EN(PIPEREG_EN),  
        . ACCUMADDSUB_OP(ACC_ADDSUB_OP), 
        . DYN_OP_SEL(DYN_ACC_ADDSUB_OP),    
        . ASIZE(18), 
        . BSIZE(18), 
        . PSIZE(64), 
        . MASK(OVERFLOW_MASK),
        . DYN_ACC_INIT(0),
        . ACC_INIT_VALUE(ACC_INIT_VALUE)
    ) U_MACC (
        . CE(CE),
        . RST(RST),
        . CLK(CLK),
        . A(A),
        . B(B),
        . A_SIGNED(A_SIGNED),
        . B_SIGNED(B_SIGNED),
        . C_SIGNED(C_SIGNED),
        . C(C),
        . PREADDSUB(PREADDSUB),
        . ACCUM_INIT(64'b0),
        . ACCUMADDSUB(ACC_ADDSUB),
        . RELOAD(RELOAD),
        . P(P),
        . OVER(OVER),
        . UNDER(UNDER),
        . R(R)
    );

    INT_FLAG #(
        . GRS_EN(GRS_EN),
        . SYNC_RST(SYNC_RST),
        . PSIZE(64),
        . PATSIZE(64),
        . MASKPATSIZE(64),
        . OUTREG_EN("TRUE")
    ) U_FLAG (
        . CE(CE),
        . RST(RST),
        . CLK(CLK),
        . P(P),
        . PATTERN(PATTERN),
        . MASKPAT(MASKPAT),
        . OVERFLOW_MASK(OVERFLOW_MASK),
        . R(R),
        . eqz(EQZ),
        . eqzm(EQZM),
        . eqom(EQOM),
        . eqpat(EQPAT),
        . eqpatn(EQPATN)
    );

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

primitive INT_LUTMUX2_UDP (dout, sel, di1, di0);
    output dout;
    input sel, di1, di0;

    table
    //  sel di1 di0 : dout
        0   ?   0   : 0 ;
        0   ?   1   : 1 ;
        1   0   ?   : 0 ;
        1   1   ?   : 1 ;
        x   0   0   : 0 ;
        x   1   1   : 1 ;
    endtable

endprimitive





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2015 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_FIFO18K_E1.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_FIFO18K_E1
#(
    parameter GRS_EN = "TRUE",
    parameter integer DATA_WIDTH = 18,//1,2,4,8,9,16,18
    parameter integer DO_REG = 0,
    parameter [13:0]  ALMOST_FULL_OFFSET  = 14'h0000,
    parameter [13:0]  ALMOST_EMPTY_OFFSET = 14'h0000,
    parameter [35:0]  RST_VAL = 36'b0,
    parameter integer USE_EMPTY = 0,
    parameter integer USE_FULL = 0,
    parameter SYNC_FIFO = "FALSE"

) (
    output        ALMOST_EMPTY,
    output        ALMOST_FULL,
    output        EMPTY,
    output        FULL,
    output [35:0] DO,
    input  [35:0] DI,
    input         WCLK,
    input         RCLK,
    input         WCE,
    input         RCE,
    input         ORCE,
    input         RST
);
// synthesis translate_off
    reg  [14:0]   rd_binary;
    reg  [14:0]   wr_binary;
    reg  [13:0]   wcnt;
    reg  [13:0]   rcnt;
    reg  [14:0]   wr_binary_next;
    reg  [14:0]   rd_binary_next;
    reg           empty_reg;
    reg           full_reg;
    reg           full_val;
    reg           almost_full_val;
    reg           almost_full_reg;
    reg           almost_empty_reg;
    reg           flagempty_en;
    reg           flagfull_en;
    reg           dout_reg_en;
    reg           sync_fifo;
    reg           grs_en;
    reg  [35:0]   dout;
    reg  [35:0]   dout_reg;

    wire [14:0]   wptr_next;
    wire [14:0]   rptr_next;
    reg  [14:0]   wptr_rclk;
    reg  [14:0]   rptr_wclk;
    wire [14:0]   wptr_next_gray;
    reg  [14:0]   wdata_buf;
    reg  [14:0]   wdata_buf_d1;
    reg  [14:0]   wdata_buf_d2;
    wire [14:0]   rptr_next_gray;
    reg  [14:0]   rdata_buf;
    reg  [14:0]   rdata_buf_d1;
    reg  [14:0]   rdata_buf_d2;
    wire          wclk,rclk;
    wire          wr_en,rd_en;
    wire          rstw,rstr;
    wire          full,empty;
    wire [35:0]   din;
    wire [35:0]   dout_int;
    wire          almost_empty,almost_full;
    wire          global_rstn;

    reg  [(DATA_WIDTH-1):0] mem [16383 : 0];//16383
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
    initial   
    begin
        case(SYNC_FIFO)
            "FALSE" : sync_fifo = 0;
            "TRUE"  : sync_fifo = 1;
            default : begin
                $display ("ERROR: GTP_FIFO18K_E1 instance %m parameter SYNC_FIFO:%s, The legal values are FALSE or TRUE.",SYNC_FIFO);
                $finish;
            end
        endcase
        
        case(USE_EMPTY)
            1'b0 : flagempty_en = 0;
            1'b1 : flagempty_en = 1;
            default : begin
                $display ("ERROR: GTP_FIFO18K_E1 instance %m parameter USE_EMPTY:%d, The legal values are 0 or 1.",USE_EMPTY);
                $finish;
            end
        endcase
        
        case(USE_FULL)
            1'b0 : flagfull_en = 0;
            1'b1 : flagfull_en = 1;
            default : begin
                $display ("ERROR: GTP_FIFO18K_E1 instance %m parameter USE_FULL:%d, The legal values are 0 or 1.",USE_FULL);
                $finish;
            end
        endcase
        
        case(DO_REG)
            1'b0 : dout_reg_en = 0;
            1'b1 : dout_reg_en = 1;
            default : begin
                $display ("ERROR: GTP_FIFO18K_E1 instance %m parameter DO_REG:%d, The legal values are 0 or 1.",DO_REG);
                $finish;
            end
        endcase

        case(GRS_EN)
            "FALSE" : grs_en = 0;
            "TRUE"  : grs_en = 1;
            default : begin
                $display ("ERROR: GTP_FIFO36K instance %m parameter GRS_EN:%s, The legal values are FALSE or TRUE.",GRS_EN);
                $finish;
            end
        endcase

        dout_reg =36'b0;
    end
//////////////////////////////////////////////////////////////////////////////////////
    assign orce_in = ORCE;
    assign din = DI;
    assign wclk = WCLK;
    assign rclk = RCLK;
    assign wr_en = WCE;
    assign rd_en = RCE;
    assign rstw = ~RST & global_rstn;
    assign rstr = ~RST & global_rstn;
    assign EMPTY = empty;
    assign FULL  = full;
    assign ALMOST_EMPTY = almost_empty;
    assign ALMOST_FULL = almost_full;
    assign WCNT = wcnt;
    assign RCNT = rcnt;
    
    always @(posedge rclk or negedge rstr )
    begin
        if(rstr == 1'b0)
            dout_reg <= RST_VAL;
        else if(orce_in)
            dout_reg <= dout_int;
    end    
    
    assign DO = dout_reg_en ? dout_reg : dout_int;
    
    assign global_rstn = grs_en ? GRS_INST.GRSNET : 1'b1;
//////////////////////////////////////////////////////////////////////////////////////
    always @ (posedge wclk or negedge rstw )  //////wr binary addr
    begin
        if (rstw == 1'b0)
             wr_binary <= 0;
        else
             wr_binary <= wr_binary_next;
    end
    
    always @ (*)
    begin
        if (full == 1'b0)
             wr_binary_next = wr_binary + wr_en;
        else
             wr_binary_next = wr_binary;
    end
    
    assign wptr_next = wr_binary_next;
//////////////////////////////////////////////////////////////////////////////////////

    always @ (*) begin
        case(DATA_WIDTH)
        1: begin
             full_val = (wr_binary_next[14:0] == {~rptr_wclk[14],rptr_wclk[13:0]});
             almost_full_val = ~rptr_wclk[14]&((({~rptr_wclk[14],rptr_wclk[13:0]} - wr_binary_next[14:0]) <= ALMOST_FULL_OFFSET) | (({~wr_binary_next[14],wr_binary_next[13:0]}) - rptr_wclk[14:0]) <= ALMOST_FULL_OFFSET) | rptr_wclk[14]&(((wr_binary_next[14:0] - {~rptr_wclk[14],rptr_wclk[13:0]}) <= ALMOST_FULL_OFFSET) | ((rptr_wclk[14:0] - {~wr_binary_next[14],wr_binary_next[13:0]}) <= ALMOST_FULL_OFFSET));
        end
        2: begin
             full_val = (wr_binary_next[13:0] == {~rptr_wclk[13],rptr_wclk[12:0]});
             almost_full_val = ~rptr_wclk[13]&((({~rptr_wclk[13],rptr_wclk[12:0]} - wr_binary_next[13:0]) <= ALMOST_FULL_OFFSET) | (({~wr_binary_next[13],wr_binary_next[12:0]}) - rptr_wclk[13:0]) <= ALMOST_FULL_OFFSET) | rptr_wclk[13]&(((wr_binary_next[13:0] - {~rptr_wclk[13],rptr_wclk[12:0]}) <= ALMOST_FULL_OFFSET) | ((rptr_wclk[13:0] - {~wr_binary_next[13],wr_binary_next[12:0]}) <= ALMOST_FULL_OFFSET));
        end
        4: begin
             full_val = (wr_binary_next[12:0] == {~rptr_wclk[12],rptr_wclk[11:0]});
             almost_full_val = ~rptr_wclk[12]&((({~rptr_wclk[12],rptr_wclk[11:0]} - wr_binary_next[12:0]) <= ALMOST_FULL_OFFSET) | (({~wr_binary_next[12],wr_binary_next[11:0]}) - rptr_wclk[12:0]) <= ALMOST_FULL_OFFSET) | rptr_wclk[12]&(((wr_binary_next[12:0] - {~rptr_wclk[12],rptr_wclk[11:0]}) <= ALMOST_FULL_OFFSET) | ((rptr_wclk[12:0] - {~wr_binary_next[12],wr_binary_next[11:0]}) <= ALMOST_FULL_OFFSET));
        end
        8, 9: begin
             full_val = (wr_binary_next[11:0] == {~rptr_wclk[11],rptr_wclk[10:0]});
             almost_full_val = ~rptr_wclk[11]&((({~rptr_wclk[11],rptr_wclk[10:0]} - wr_binary_next[11:0]) <= ALMOST_FULL_OFFSET) | (({~wr_binary_next[11],wr_binary_next[10:0]}) - rptr_wclk[11:0]) <= ALMOST_FULL_OFFSET) | rptr_wclk[11]&(((wr_binary_next[11:0] - {~rptr_wclk[11],rptr_wclk[10:0]}) <= ALMOST_FULL_OFFSET) | ((rptr_wclk[11:0] - {~wr_binary_next[11],wr_binary_next[10:0]}) <= ALMOST_FULL_OFFSET));
        end
        16, 18: begin
             full_val = (wr_binary_next[10:0] == {~rptr_wclk[10],rptr_wclk[9:0]});
             almost_full_val = ~rptr_wclk[10]&((({~rptr_wclk[10],rptr_wclk[9:0]} - wr_binary_next[10:0]) <= ALMOST_FULL_OFFSET) | (({~wr_binary_next[10],wr_binary_next[9:0]}) - rptr_wclk[10:0]) <= ALMOST_FULL_OFFSET) | rptr_wclk[10]&(((wr_binary_next[10:0] - {~rptr_wclk[10],rptr_wclk[9:0]}) <= ALMOST_FULL_OFFSET) | ((rptr_wclk[10:0] - {~wr_binary_next[10],wr_binary_next[9:0]}) <= ALMOST_FULL_OFFSET));
        end
        32, 36: begin
             full_val = (wr_binary_next[9:0] == {~rptr_wclk[9],rptr_wclk[8:0]});
             almost_full_val = ~rptr_wclk[9]&((({~rptr_wclk[9],rptr_wclk[8:0]} - wr_binary_next[9:0]) <= ALMOST_FULL_OFFSET) | (({~wr_binary_next[9],wr_binary_next[8:0]}) - rptr_wclk[9:0]) <= ALMOST_FULL_OFFSET) | rptr_wclk[9]&(((wr_binary_next[9:0] - {~rptr_wclk[9],rptr_wclk[8:0]}) <= ALMOST_FULL_OFFSET) | ((rptr_wclk[9:0] - {~wr_binary_next[9],wr_binary_next[8:0]}) <= ALMOST_FULL_OFFSET));
             //almost_full_val = (({~rptr_wclk[9],rptr_wclk[8:0]} - wr_binary_next[9:0]) <= ALMOST_FULL_OFFSET) | ((wr_binary_next[9:0] - {~rptr_wclk[9],rptr_wclk[8:0]}) <= ALMOST_FULL_OFFSET);
        end
        default: begin  //default x18
             full_val = (wr_binary_next[10:0] == {~rptr_wclk[10],rptr_wclk[9:0]});
             almost_full_val = ~rptr_wclk[10]&((({~rptr_wclk[10],rptr_wclk[9:0]} - wr_binary_next[10:0]) <= ALMOST_FULL_OFFSET) | (({~wr_binary_next[10],wr_binary_next[9:0]}) - rptr_wclk[10:0]) <= ALMOST_FULL_OFFSET) | rptr_wclk[10]&(((wr_binary_next[10:0] - {~rptr_wclk[10],rptr_wclk[9:0]}) <= ALMOST_FULL_OFFSET) | ((rptr_wclk[10:0] - {~wr_binary_next[10],wr_binary_next[9:0]}) <= ALMOST_FULL_OFFSET));
        end
        endcase
    end
    
    always @ (posedge wclk or negedge rstw) begin //////write full flag
        if (rstw == 1'b0)
             full_reg <= 1'b0;
        else
             full_reg <= full_val;
    end
    
    assign full = flagfull_en & full_reg;

    wire [14:0] write_water_level;
    assign write_water_level = wr_binary_next - rptr_wclk;
    always @ (posedge wclk or negedge rstw) begin //////write almost_full flag
        if (rstw == 1'b0)
             almost_full_reg <= 1'b0;
        else
             almost_full_reg <= (write_water_level >= ALMOST_FULL_OFFSET);
    end
    
    assign almost_full = flagfull_en & almost_full_reg;
//////////////////////////////////////////////////////////////////////////////////////
    always @ (posedge rclk or negedge rstr) begin
        if(rstr == 1'b0)
             rd_binary <= 0;
        else
             rd_binary <= rd_binary_next;
    end

    
    wire empty_int;
    assign empty_int = wptr_rclk==rd_binary_next;
    always @ (*) begin
          if ((~empty_reg) & rd_en)
             rd_binary_next = rd_binary + 1;
          else
             rd_binary_next = rd_binary;
    end
    
    assign rptr_next = rd_binary_next;
    
    always @ (posedge rclk or negedge rstr) begin
          if (rstr == 1'b0) begin
              empty_reg <= 1'b1;
          end
          else begin
              empty_reg <= wptr_rclk == rd_binary_next;
          end
    end
    
    assign empty = ~flagempty_en |empty_reg;
    
    always @ (posedge rclk or negedge rstr) begin
          if (rstr == 1'b0) begin
              almost_empty_reg <= 1'b1;
          end
          else begin
              almost_empty_reg <= (wptr_rclk - rd_binary_next) <= ALMOST_EMPTY_OFFSET;
          end
    end
    
    assign almost_empty = ~flagempty_en |almost_empty_reg;
//////////////////////////////////////////////////////////////////////////////////////
    always @ (wr_binary) begin
        case(DATA_WIDTH)
             1:     wcnt <=  wr_binary[13:0];
             2:     wcnt <= {wr_binary[12:0],1'b1};
             4:     wcnt <= {wr_binary[11:0],2'b11};
             8:     wcnt <= {wr_binary[10:0],3'b111};
             9:     wcnt <= {wr_binary[10:0],3'b111};
             16:    wcnt <= {wr_binary[9:0],4'b1111};
             18:    wcnt <= {wr_binary[9:0],4'b1111};
             32:    wcnt <= {wr_binary[8:0],5'b1111};
             36:    wcnt <= {wr_binary[8:0],5'b1111};
             default:
                    wcnt <= 14'b0;
        endcase
    end
    
    always @ (rd_binary) begin
        case(DATA_WIDTH)
             1:     rcnt <=  rd_binary[13:0];
             2:     rcnt <= {rd_binary[12:0],1'b1};
             4:     rcnt <= {rd_binary[11:0],2'b11};
             8:     rcnt <= {rd_binary[10:0],3'b111};
             9:     rcnt <= {rd_binary[10:0],3'b111};
             16:    rcnt <= {rd_binary[9:0],4'b1111};
             18:    rcnt <= {rd_binary[9:0],4'b1111};
             32:    rcnt <= {rd_binary[8:0],5'b1111};
             36:    rcnt <= {rd_binary[8:0],5'b1111};
             default:
                    rcnt <= 14'b0;
        endcase
    end
//////////////////////////////////////////////////////////////////////////////////////
    assign wptr_next_gray = (wptr_next>>1)^wptr_next;
    assign rptr_next_gray = (rptr_next>>1)^rptr_next;
    
    always @(posedge wclk or negedge rstw)
    begin
        if(rstw == 1'b0)
        begin 
            wdata_buf <= 0;
            rdata_buf_d1 <= 0;
            rdata_buf_d2 <= 0;
        end else begin
            wdata_buf <= wptr_next_gray;
            rdata_buf_d1 <= rdata_buf;
            if(sync_fifo)
                rdata_buf_d2 <= rptr_next_gray;
            else
                rdata_buf_d2 <= rdata_buf_d1;
        end
    end
    
    always @(posedge rclk or negedge rstr)
    begin
        if(rstr == 1'b0)
        begin
            wdata_buf_d1 <= 0;
            wdata_buf_d2 <= 0;
            rdata_buf <= 0;
        end else begin
            wdata_buf_d1 <= wdata_buf;
            rdata_buf <= rptr_next_gray;
            if(sync_fifo)
                wdata_buf_d2 <= wptr_next_gray;
            else
                wdata_buf_d2 <= wdata_buf_d1;
        end
    end
    
    integer i,j,k;
    
    always @(wdata_buf_d2) begin
       for (i=0; i< 15;i=i+1)
           wptr_rclk[i] = ^(wdata_buf_d2>>i);
    end
    
    always @(rdata_buf_d2) begin
       for (j=0; j< 15;j=j+1)
           rptr_wclk[j] = ^(rdata_buf_d2>>j);
    end
//////////////////////////////////////////////////////////////////////////////////////
    initial
    begin
        for(k=0;k<(1<<14);k=k+1)
            mem[k] <= {DATA_WIDTH{1'b0}};
    end
    
    always @(posedge rclk or negedge rstr)
    begin
        if(rstr == 1'b0)
            dout <= RST_VAL;
        else if(rd_en)
            dout <= mem[rcnt];
    end

    assign dout_int = dout;

    always @(posedge wclk)
    begin
        if(wr_en && !full_reg)
            mem[wcnt] <= din;
    end


// synthesis translate_on
endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_OGSER7.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_OGSER7 #(
parameter GRS_EN = "TRUE", //"TRUE"; "FALSE"  
parameter LRS_EN = "TRUE"   //"TRUE"; "FALSE"  
)(
output PADO,
input [6:0] D,
input SERCLK,
input RCLK,
input RST
);

//synthesis translate_off
reg [6:0] d_rclk;
reg [2:0] cnt;
reg shift_en;
reg [7:0] capture_d_reg;
reg [7:0] shift_d_reg;
reg PADO_POS;
reg PADO_NEG;


initial begin
d_rclk          = 0;
cnt             = 0;
shift_en        = 0;
capture_d_reg   = 0;
shift_d_reg     = 0;
PADO_POS        = 0;
PADO_NEG        = 0;  
end
assign global_rstn = (GRS_EN == "TRUE") ? GRS_INST.GRSNET : 1'b1;
assign lsr_rstn = LRS_EN == "TRUE" ? (~RST) : 1'b1;

always @(posedge RCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      d_rclk <= 0;
   else if (!lsr_rstn)
      d_rclk <= 0;
   else
      d_rclk <= D;
      
always @(posedge SERCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      cnt <= 0;
   else if (!lsr_rstn)
      cnt <= 0;
   else if (cnt == 6)
      cnt <= 0;
   else
      cnt <= cnt + 1;   
      
assign capture_en_0 = cnt == 3;
assign capture_en_1 = cnt == 6;

always @(posedge SERCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      shift_en <= 0;
   else if (!lsr_rstn)
      shift_en <= 0;
   else 
      shift_en <= capture_en_0 | capture_en_1;
      
always @(posedge SERCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      capture_d_reg <= 0;
   else if (!lsr_rstn)
      capture_d_reg <= 0;
   else if (capture_en_0)
      capture_d_reg <= {1'b0, d_rclk[6:0]};
   else if (capture_en_1)
      capture_d_reg <= {d_rclk[6:0], capture_d_reg[6]};
      
always @(posedge SERCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      shift_d_reg <= 0;
   else if (!lsr_rstn)
      shift_d_reg <= 0;
   else if (shift_en)
      shift_d_reg <= capture_d_reg;
   else
      shift_d_reg <= {2'd0, shift_d_reg[7:2]};
      
always @(posedge SERCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      PADO_POS <= 0;
   else if (!lsr_rstn)
      PADO_POS <= 0;
   else
      PADO_POS <= shift_d_reg[1];
   
always @(negedge SERCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      PADO_NEG <= 0;
   else if (!lsr_rstn)
      PADO_NEG <= 0;
   else
      PADO_NEG <= shift_d_reg[0];
   
assign PADO =  SERCLK ? PADO_NEG : PADO_POS;
//synthesis translate_on

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_OGDDR.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_OGDDR #(
parameter GRS_EN = "TRUE", //"TRUE"; "FALSE"
parameter LRS_EN = "TRUE"   //"TRUE"; "FALSE"
)(
output  PADO,
output  PADT,
input [1:0] D,
input T,
input RCLK,
input RST
);

//synthesis translate_off
reg [1:0] d_rclk;
reg t_rclk;
reg [1:0] shift_d_reg;
reg shift_t_reg;
reg PADO_POS;
reg PADT_reg;
reg PADO_NEG;

initial begin
d_rclk      = 0;
t_rclk      = 0;
shift_d_reg = 0;
shift_t_reg = 0;
PADO_POS    = 0;
PADT_reg    = 0;
PADO_NEG    = 0;
end
assign global_rstn = (GRS_EN == "TRUE") ? GRS_INST.GRSNET : 1'b1;
assign lsr_rstn = LRS_EN == "TRUE" ? (~RST) : 1'b1;

always @(posedge RCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn) begin
      d_rclk <= 0;
      t_rclk <= 0;
   end   
   else if (!lsr_rstn) begin
      d_rclk <= 0;
      t_rclk <= 0;
   end   
   else begin
      d_rclk <= D;
      t_rclk <= T;
   end   

always @(posedge RCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn) begin
      shift_d_reg <= 0;
      shift_t_reg <= 0;
   end   
   else if (!lsr_rstn) begin
      shift_d_reg <= 0;
      shift_t_reg <= 0;
   end   
   else begin
      shift_d_reg <= d_rclk;
      shift_t_reg <= t_rclk;
   end   
   
always @(posedge RCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn) begin
      PADO_POS <= 0;
      PADT_reg <= 0;
   end
   else if (!lsr_rstn) begin
      PADO_POS <= 0;
      PADT_reg <= 0;
   end
   else begin
      PADO_POS <= shift_d_reg[1];
      PADT_reg <= shift_t_reg;    
   end           
   
always @(negedge RCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn) begin
      PADO_NEG <= 0;
   end
   else if (!lsr_rstn) begin
      PADO_NEG <= 0;
   end
   else begin
      PADO_NEG <= shift_d_reg[0];
   end           


assign PADO =  RCLK ? PADO_NEG : PADO_POS;
assign PADT = PADT_reg;
//synthesis translate_on

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_MULTADD18.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

//P = A0*B0 +/- A1*B1
module GTP_MULTADD18 #(
    parameter GRS_EN      = "TRUE", //"TRUE"; "FALSE"
    parameter SYNC_RST    = "FALSE", //"TRUE"; "FALSE"
    parameter INREG_EN    = "FALSE", //"TRUE"; "FALSE"
    parameter PIPEREG_EN  = "FALSE", //"TRUE"; "FALSE"
    parameter OUTREG_EN   = "FALSE", //"TRUE"; "FALSE"
    parameter ADDSUB_OP     = 0 ,
    parameter DYN_ADDSUB_OP = 1
)(
    output  [37-1:0] P,          //product
    input   CE,
    input   RST,
    input   CLK,
    input   A_SIGNED,
    input   [18-1:0] A0,
    input   [18-1:0] A1,
    input   B_SIGNED,
    input   [18-1:0] B0,
    input   [18-1:0] B1,
    input   ADDSUB
);

    INT_PREADD_MULTADD #(
        . GRS_EN(GRS_EN),
        . SYNC_RST(SYNC_RST),   
        . INREG_EN(INREG_EN),   
        . PIPEREG_EN(PIPEREG_EN), 
        . OUTREG_EN(OUTREG_EN),  
        . ADDSUB_OP(ADDSUB_OP),  
        . DYN_OP_ADDSUB(DYN_ADDSUB_OP), 
        . ASIZE(18), 
        . BSIZE(18),
        . PREADD_EN(0)
    ) U_MULTADD18 (
        . CE(CE),
        . RST(RST),
        . CLK(CLK),
        . A_SIGNED(A_SIGNED),
        . A0(A0),
        . A1(A1),
        . B_SIGNED(B_SIGNED),
        . B0(B0),
        . B1(B1),
        . C_SIGNED(B_SIGNED),
        . C0(18'b0),
        . C1(18'b0),
        . PREADDSUB(2'b0),
        . ADDSUB(ADDSUB),
        . P(P)
    );

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_PREADD_MULT27.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

//P = A*(B+C)
`timescale 1 ns / 1 ps

module GTP_PREADD_MULT27 #(
    parameter GRS_EN      = "TRUE", //"TRUE"; "FALSE"
    parameter SYNC_RST    = "FALSE", //"TRUE"; "FALSE"
    parameter INREG_EN    = "FALSE", //"TRUE"; "FALSE"
    parameter PREREG_EN   = "FALSE", //"TRUE"; "FALSE"
    parameter OUTREG_EN   = "FALSE"  //"TRUE"; "FALSE"
)(
    output  [54-1:0] P,
    input   CE,
    input   RST,
    input   CLK,
    input   A_SIGNED,
    input   [27-1:0] A,
    input   B_SIGNED,
    input   [26-1:0] B,
    input   C_SIGNED,
    input   [26-1:0] C,
    input   PREADDSUB
);

    INT_PREADD_MULT  #(.GRS_EN(GRS_EN),
        .SYNC_RST(SYNC_RST),    
        .INREG_EN(INREG_EN),    
        .PREREG_EN(PREREG_EN),    
        .OUTREG_EN(OUTREG_EN),   
        .ASIZE(27),  
        .BSIZE(26)
    ) U_INT_PREADD_MULT (
        .CE(CE),
        .RST(RST),
        .CLK(CLK),
        .A_SIGNED(A_SIGNED),
        .A(A),
        .B_SIGNED(B_SIGNED),
        .B(B),
        .C_SIGNED(C_SIGNED),
        .C(C),
        .PREADDSUB(PREADDSUB),
        .P(P)
    );

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_DDC.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_DDC #(
parameter GRS_EN = "TRUE",             //"TRUE"; "FALSE"
parameter DDC_MODE = "FULL_RATE", //"FULL_RATE"; "HALF_RATE"; "QUAD_RATE"
parameter IFIFO_GENERIC  ="FALSE",       //"TRUE"; "FALSE"
parameter WCLK_DELAY_OFFSET = 9'd0,          //0~255 for posedge adjust; 256~511 for negedge adjust; bit[8] used as signed flag
parameter DQSI_DELAY_OFFSET = 9'd0,          //0~255 for posedge adjust; 256~511 for negedge adjust; bit[8] used as signed flag
parameter CLKA_GATE_EN = "FALSE",
parameter R_DELAY_STEP_EN = "TRUE", //"TRUE"; "FALSE"
parameter R_MOVE_EN = "FALSE", //"TRUE"; "FALSE"
parameter W_MOVE_EN = "FALSE", //"TRUE"; "FALSE"
parameter R_EXTEND = "FALSE", //"TRUE"; "FALSE"
parameter RADDR_INIT = 3'd0
)(
    //output
    output WDELAY_OB,
    output WCLK,
    output WCLK_DELAY,
    output RDELAY_OB,
    output DQSI_DELAY,
    output DGTS,
    output READ_VALID,
    output [2:0] IFIFO_WADDR,
    output [2:0] IFIFO_RADDR,
    //input
    input RST,
    input CLKB,
    input CLKA,
    input CLKA_GATE,
    input [7:0] DELAY_STEP1,
    input [7:0] DELAY_STEP0,
    input       W_DIRECTION,
    input       W_MOVE,
    input       W_LOAD_N,
    input [3:0] DQS_GATE_CTRL,
    input [2:0] READ_CLK_CTRL,
    input DQSI,
    input      R_DIRECTION,
    input      R_MOVE,
    input      R_LOAD_N
)/* synthesis syn_black_box */;

//synthesis translate_off
    //reg statement
    reg [1:0] DQS_GATE_CTRL_gate_d;
    reg [1:0] DQS_GATE_CTRL_gate_dd;
    reg [3:0] DQS_GATE_CTRL_d1;
    reg [3:0] DQS_GATE_CTRL_d2;
    reg [3:0] DQS_GATE_CTRL_d3;
    reg gate_st;
    reg [3:0] DQS_GATE_CTRL_d4;
    reg DQS_GATE_CTRL_d5;
    reg DQS_GATE_CTRL_d6;
    reg sel_gate_clk;
    reg DQS_GATE_CTRL_gate;
    reg DQS_GATE_CTRL_comb_d1;
    reg DQS_GATE_CTRL_comb_d2;
    reg [1:0] DQS_GATE_CTRL_comb_and_d;
    reg start_wr;
    reg [2:0] WADDR_reg;
    reg [2:0] IFIFO_WADDR_reg;
    reg start_rd;
    reg [2:0] RADDR_reg;
    reg RDVALID_reg;
    reg DQSIN_gated_reg;
    reg [7:0] adj_dly_wclk_del;
    reg [7:0] adj_dly_dqsi;
    reg read_enable_tmp;
    reg new_st;
    reg new_transfer_d;
    reg read_enable_d1;
    reg read_enable_d2;
    reg [1:0] cnt;
    reg [1:0] gate_cnt;
    reg [1:0] new_cnt;
    reg [7:0] gate_d;
    reg [2:0] WADDR_reg_d1;
    reg [2:0] WADDR_reg_d2;
    reg [2:0] RADDR_reg_plus1;
    reg new_rd_en_reg;
    //wire statement
    wire DQSIN_gated;
    wire new_transfer;

initial 
begin
    if ((GRS_EN == "TRUE")  || (GRS_EN == "FALSE")) 
    begin
    end
    else
    begin
        $display (" GTP_DDC error: illegal setting for GRS_EN"); 
    end
    if ((DDC_MODE == "FULL_RATE") || (DDC_MODE == "HALF_RATE")  || (DDC_MODE == "QUAD_RATE")) 
    begin
    end
    else 
    begin
        $display (" GTP_DDC error: illegal setting for DDC_MODE");
    end
    if ((IFIFO_GENERIC == "TRUE") || (IFIFO_GENERIC == "FALSE")) 
    begin
    end
    else
    begin
       $display (" GTP_DDC error: illegal setting for IFIFO_GENERIC");
    end
    if ((CLKA_GATE_EN == "TRUE")   || (CLKA_GATE_EN == "FALSE")) 
    begin
    end
    else
    begin
        $display (" GTP_DDC error: illegal setting for CLKA_GATE_EN");
    end
    if ((R_DELAY_STEP_EN == "TRUE")   || (R_DELAY_STEP_EN == "FALSE")) 
    begin
    end
    else
    begin
        $display (" GTP_DDC error: illegal setting for R_DELAY_STEP_EN");
    end
    if ((R_MOVE_EN == "TRUE")   || (R_MOVE_EN == "FALSE")) 
    begin
    end
    else
    begin
        $display (" GTP_DDC error: illegal setting for R_MOVE_EN");
    end
    if ((W_MOVE_EN == "TRUE")   || (W_MOVE_EN == "FALSE")) 
    begin
    end
    else
    begin
        $display (" GTP_DDC error: illegal setting for W_MOVE_EN");
    end
    if ((R_EXTEND == "TRUE")   || (R_EXTEND == "FALSE")) 
    begin
    end
    else
    begin
        $display (" GTP_DDC error: illegal setting for R_EXTEND");
    end

    DQSIN_gated_reg = 1'b0;  
    DQS_GATE_CTRL_gate_d = 0;
    DQS_GATE_CTRL_gate_dd = 0;
    DQS_GATE_CTRL_d1 = 0;
    DQS_GATE_CTRL_d2 = 0;
    DQS_GATE_CTRL_d3 = 0;
    gate_st          = 0;
    DQS_GATE_CTRL_d4 = 0;
    DQS_GATE_CTRL_d5 = 0;
    DQS_GATE_CTRL_d6 = 0;
    sel_gate_clk = 0;
    DQS_GATE_CTRL_gate = 0;
    DQS_GATE_CTRL_comb_d1 = 0;
    DQS_GATE_CTRL_comb_d2 = 0;
    DQS_GATE_CTRL_comb_and_d = 0;
    start_wr  = 0;
    WADDR_reg = 0;
    IFIFO_WADDR_reg = 0;
    start_rd  = 0;
    RADDR_reg = RADDR_INIT;
    RDVALID_reg = 0;
    DQSIN_gated_reg = 0;
    adj_dly_wclk_del = 0;
    adj_dly_dqsi = 0;
    read_enable_tmp = 0;
    new_st = 0;
    new_transfer_d = 0;
    read_enable_d1 = 0;
    read_enable_d2 = 0;
    cnt = 0;
    gate_cnt = 0;
    new_cnt = 0;  
    gate_d = 0;
    WADDR_reg_d1 = 0;
    WADDR_reg_d2 = 0;
    RADDR_reg_plus1 = 0;
    new_rd_en_reg = 0;
end

assign global_rstn = GRS_EN == "TRUE" ? GRS_INST.GRSNET : 1'b1;
assign lsr_rstn = ~RST;

wire global_rstn_cgn;
wire lsr_rstn_cgn;
wire gatein;


assign gatein = CLKA_GATE_EN == "TRUE" ? (~CLKA_GATE) : 1'b1;

assign rstn_fifo = (lsr_rstn & global_rstn) & gatein;

assign rst_start_rd = start_rd & rstn_fifo;

always @(negedge CLKA or posedge RST)
begin
    if (RST) 
    begin
        gate_d <= 8'd0;
    end
    else if (CLKA_GATE_EN == "TRUE")
        gate_d <= {gate_d[6:0], CLKA_GATE};
    else
        gate_d <= 8'd0;
end

assign ioclk_gated = CLKA & (~gate_d[2]);

wire [255:0] wclk_delay_chain;
assign #0.3 wclk_delay_chain[0] = (DDC_MODE == "FULL_RATE") ? CLKB : ioclk_gated;
genvar gen_i;
generate  
    for(gen_i=1;gen_i<256;gen_i=gen_i+1) 
    begin
        assign #0.025 wclk_delay_chain[gen_i] =  wclk_delay_chain[gen_i-1];
    end
endgenerate

assign WCLK_comb = wclk_delay_chain[DELAY_STEP0];

assign WCLK = WCLK_comb;

assign WL_CTRL_b0_tmp = W_MOVE_EN == "TRUE" ? W_LOAD_N : 1'b0;
wire [8:0]  WCLK_DEL_OFFSET_tmp = WCLK_DELAY_OFFSET;

//wire [7:0] DLL_STEP_PLUS_WCLK_DEL_OFFSET = WCLK_DEL_OFFSET_tmp[8] ? (DLL_STEP - WCLK_DEL_OFFSET_tmp[7:0]) : (DLL_STEP + WCLK_DEL_OFFSET_tmp[7:0]);
wire [7:0] DLL_STEP_PLUS_WCLK_DEL_OFFSET = DELAY_STEP1 + WCLK_DEL_OFFSET_tmp[7:0];

wire DLL_STEP_PLUS_WCLK_DEL_OFFSET_co_0 = DELAY_STEP1[0] && WCLK_DEL_OFFSET_tmp[0];
wire DLL_STEP_PLUS_WCLK_DEL_OFFSET_co_1 = (DELAY_STEP1[1] && WCLK_DEL_OFFSET_tmp[1]) || ((DELAY_STEP1[1] || WCLK_DEL_OFFSET_tmp[1]) && DLL_STEP_PLUS_WCLK_DEL_OFFSET_co_0);
wire DLL_STEP_PLUS_WCLK_DEL_OFFSET_co_2 = (DELAY_STEP1[2] && WCLK_DEL_OFFSET_tmp[2]) || ((DELAY_STEP1[2] || WCLK_DEL_OFFSET_tmp[2]) && DLL_STEP_PLUS_WCLK_DEL_OFFSET_co_1);
wire DLL_STEP_PLUS_WCLK_DEL_OFFSET_co_3 = (DELAY_STEP1[3] && WCLK_DEL_OFFSET_tmp[3]) || ((DELAY_STEP1[3] || WCLK_DEL_OFFSET_tmp[3]) && DLL_STEP_PLUS_WCLK_DEL_OFFSET_co_2);
wire DLL_STEP_PLUS_WCLK_DEL_OFFSET_co_4 = (DELAY_STEP1[4] && WCLK_DEL_OFFSET_tmp[4]) || ((DELAY_STEP1[4] || WCLK_DEL_OFFSET_tmp[4]) && DLL_STEP_PLUS_WCLK_DEL_OFFSET_co_3);
wire DLL_STEP_PLUS_WCLK_DEL_OFFSET_co_5 = (DELAY_STEP1[5] && WCLK_DEL_OFFSET_tmp[5]) || ((DELAY_STEP1[5] || WCLK_DEL_OFFSET_tmp[5]) && DLL_STEP_PLUS_WCLK_DEL_OFFSET_co_4);
wire DLL_STEP_PLUS_WCLK_DEL_OFFSET_co_6 = (DELAY_STEP1[6] && WCLK_DEL_OFFSET_tmp[6]) || ((DELAY_STEP1[6] || WCLK_DEL_OFFSET_tmp[6]) && DLL_STEP_PLUS_WCLK_DEL_OFFSET_co_5);
wire DLL_STEP_PLUS_WCLK_DEL_OFFSET_co_7 = (DELAY_STEP1[7] && WCLK_DEL_OFFSET_tmp[7]) || ((DELAY_STEP1[7] || WCLK_DEL_OFFSET_tmp[7]) && DLL_STEP_PLUS_WCLK_DEL_OFFSET_co_6);


assign DLL_STEP_PLUS_WCLK_DEL_OFFSET_sel= ~(WCLK_DEL_OFFSET_tmp[8] ^ DLL_STEP_PLUS_WCLK_DEL_OFFSET_co_7);


wire [7:0] DLL_STEP_WCLK_DEL = WCLK_DEL_OFFSET_tmp[8] ? (DLL_STEP_PLUS_WCLK_DEL_OFFSET_sel ? DLL_STEP_PLUS_WCLK_DEL_OFFSET[7:0] : 8'd0) :
                              (DLL_STEP_PLUS_WCLK_DEL_OFFSET_sel ? DLL_STEP_PLUS_WCLK_DEL_OFFSET[7:0] : 8'd255);

wire [7:0] WL_STEP_24 = (DDC_MODE == "FULL_RATE") ? 8'd0 : DELAY_STEP0; 

wire [7:0] adj_dly_wclk_del_9b = DLL_STEP_WCLK_DEL + WL_STEP_24;

wire DLL_STEP_PLUS_WCLK_DEL_OFFSET2_co_0 = DLL_STEP_WCLK_DEL[0] && WL_STEP_24[0];
wire DLL_STEP_PLUS_WCLK_DEL_OFFSET2_co_1 = (DLL_STEP_WCLK_DEL[1] && WL_STEP_24[1]) || ((DLL_STEP_WCLK_DEL[1] || WL_STEP_24[1]) && DLL_STEP_PLUS_WCLK_DEL_OFFSET2_co_0);
wire DLL_STEP_PLUS_WCLK_DEL_OFFSET2_co_2 = (DLL_STEP_WCLK_DEL[2] && WL_STEP_24[2]) || ((DLL_STEP_WCLK_DEL[2] || WL_STEP_24[2]) && DLL_STEP_PLUS_WCLK_DEL_OFFSET2_co_1);
wire DLL_STEP_PLUS_WCLK_DEL_OFFSET2_co_3 = (DLL_STEP_WCLK_DEL[3] && WL_STEP_24[3]) || ((DLL_STEP_WCLK_DEL[3] || WL_STEP_24[3]) && DLL_STEP_PLUS_WCLK_DEL_OFFSET2_co_2);
wire DLL_STEP_PLUS_WCLK_DEL_OFFSET2_co_4 = (DLL_STEP_WCLK_DEL[4] && WL_STEP_24[4]) || ((DLL_STEP_WCLK_DEL[4] || WL_STEP_24[4]) && DLL_STEP_PLUS_WCLK_DEL_OFFSET2_co_3);
wire DLL_STEP_PLUS_WCLK_DEL_OFFSET2_co_5 = (DLL_STEP_WCLK_DEL[5] && WL_STEP_24[5]) || ((DLL_STEP_WCLK_DEL[5] || WL_STEP_24[5]) && DLL_STEP_PLUS_WCLK_DEL_OFFSET2_co_4);
wire DLL_STEP_PLUS_WCLK_DEL_OFFSET2_co_6 = (DLL_STEP_WCLK_DEL[6] && WL_STEP_24[6]) || ((DLL_STEP_WCLK_DEL[6] || WL_STEP_24[6]) && DLL_STEP_PLUS_WCLK_DEL_OFFSET2_co_5);
wire DLL_STEP_PLUS_WCLK_DEL_OFFSET2_co_7 = (DLL_STEP_WCLK_DEL[7] && WL_STEP_24[7]) || ((DLL_STEP_WCLK_DEL[7] || WL_STEP_24[7]) && DLL_STEP_PLUS_WCLK_DEL_OFFSET2_co_6);

assign DLL_STEP_PLUS_WCLK_DEL_OFFSET_sel2= ~(1'b0 ^ DLL_STEP_PLUS_WCLK_DEL_OFFSET2_co_7);

wire [7:0] adj_dly_wclk_del_init = DLL_STEP_PLUS_WCLK_DEL_OFFSET_sel2 ? adj_dly_wclk_del_9b[7:0] : 8'd255;



always @(WL_CTRL_b0_tmp or adj_dly_wclk_del_init) 
begin
    if (!WL_CTRL_b0_tmp) 
        adj_dly_wclk_del <= adj_dly_wclk_del_init;    
end
      
always @(negedge W_MOVE) 
begin
    if (!WL_CTRL_b0_tmp)
        adj_dly_wclk_del <= adj_dly_wclk_del_init;
    else if (W_DIRECTION && (adj_dly_wclk_del != 8'd0))
        adj_dly_wclk_del <= adj_dly_wclk_del - 1;
    else if ((~W_DIRECTION) && (adj_dly_wclk_del != 8'd255))
        adj_dly_wclk_del <= adj_dly_wclk_del + 1;
end


assign WDELAY_OB = (W_DIRECTION && (adj_dly_wclk_del == 8'd0)) || ((~W_DIRECTION) && (adj_dly_wclk_del == 8'd255));

wire [255:0] wclk_del_delay_chain;
assign #0.3 wclk_del_delay_chain[0] = (DDC_MODE == "FULL_RATE") ? CLKB : ioclk_gated;
genvar gen_j;
generate  
    for(gen_j=1;gen_j<256;gen_j=gen_j+1) 
    begin
        assign #0.025 wclk_del_delay_chain[gen_j] =  wclk_del_delay_chain[gen_j-1];
    end
endgenerate

assign WCLK_DEL_TMP = ~wclk_del_delay_chain[adj_dly_wclk_del];
assign WCLK_DELAY = wclk_del_delay_chain[adj_dly_wclk_del];

always @(posedge CLKB or negedge global_rstn or negedge lsr_rstn)
begin
    if (!global_rstn) 
    begin
        DQS_GATE_CTRL_d1 <= 0;
        DQS_GATE_CTRL_d2 <= 0;
    end
    else if (!lsr_rstn) 
    begin
        DQS_GATE_CTRL_d1 <= 0;
        DQS_GATE_CTRL_d2 <= 0;
    end
    else 
    begin
        if (DDC_MODE == "QUAD_RATE")
            DQS_GATE_CTRL_d2 <= DQS_GATE_CTRL;
        else 
        begin
            DQS_GATE_CTRL_d1 <= DQS_GATE_CTRL;
            DQS_GATE_CTRL_d2 <= #1 DQS_GATE_CTRL_d1;   
        end
    end
end

always @(posedge CLKA or negedge global_rstn or negedge lsr_rstn)
begin
    if (!global_rstn) 
    begin
        cnt <= 0;
    end
    else if (!lsr_rstn) 
    begin
        cnt <= 0;
    end
    else 
    begin
      cnt <= cnt + 1;
    end
end

assign capture = (DDC_MODE == "HALF_RATE") ? (~cnt[0]) : cnt == 3;

always @(posedge CLKA or negedge global_rstn or negedge lsr_rstn)
begin
    if (!global_rstn)
        DQS_GATE_CTRL_d3 <= 0;
    else if (!lsr_rstn)
        DQS_GATE_CTRL_d3 <= 0;
    else if (capture)
        DQS_GATE_CTRL_d3 <= #0.2 DQS_GATE_CTRL_d2;
end

assign WCLK_sel = WCLK;

always @(posedge WCLK_sel or negedge global_rstn or negedge lsr_rstn)
begin
    if (!global_rstn) 
    begin
        gate_st       <= 0;
        gate_cnt      <= 0;
    end
    else if (!lsr_rstn) 
    begin
        gate_st       <= 0;
        gate_cnt      <= 0;
    end
    else 
    begin
        gate_st       <= 1;
        if (gate_st)
            gate_cnt   <= gate_cnt + 1;
    end
end

assign shift = R_EXTEND == "TRUE" ? ((DDC_MODE == "HALF_RATE") ? gate_cnt[0] : (gate_cnt == 2)) :
                 ((DDC_MODE == "HALF_RATE") ? ~gate_cnt[0] : (gate_cnt == 1));

always @(posedge WCLK_sel or negedge global_rstn or negedge lsr_rstn)
begin
    if (!global_rstn)
        DQS_GATE_CTRL_d4 <= 0;
    else if (!lsr_rstn)
        DQS_GATE_CTRL_d4 <= 0;
    else if (shift)
        DQS_GATE_CTRL_d4 <= #0.2 DQS_GATE_CTRL_d3;     
    else
        DQS_GATE_CTRL_d4 <= {1'b0, DQS_GATE_CTRL_d4[3:1]};
end

always @(posedge WCLK_sel or negedge global_rstn or negedge lsr_rstn)
begin
    if (!global_rstn) 
    begin
        DQS_GATE_CTRL_d5 <= 0;
        DQS_GATE_CTRL_d6 <= 0;
    end
    else if (!lsr_rstn) 
    begin
        DQS_GATE_CTRL_d5 <= 0;
        DQS_GATE_CTRL_d6 <= 0;
    end   
    else 
    begin     
        DQS_GATE_CTRL_d5 <= DQS_GATE_CTRL_d4[0];
        if (DDC_MODE == "FULL_RATE")
            DQS_GATE_CTRL_d6 <= #0.1 DQS_GATE_CTRL_d2[0];
        else
            DQS_GATE_CTRL_d6 <= #0.1 DQS_GATE_CTRL_d5;
    end
end

always @(READ_CLK_CTRL or WCLK_sel or WCLK_DEL_TMP) 
begin
    case (READ_CLK_CTRL[1:0])
        2'd0: sel_gate_clk = ~ WCLK_DEL_TMP;
        2'd1: sel_gate_clk = ~ WCLK_sel;
        2'd2: sel_gate_clk = WCLK_DEL_TMP;
        2'd3: sel_gate_clk = WCLK_sel;
    endcase
end

always @(posedge sel_gate_clk or negedge global_rstn or negedge lsr_rstn)
begin
    if (!global_rstn)
        DQS_GATE_CTRL_comb_d1 <= 0;
    else if (!lsr_rstn)
        DQS_GATE_CTRL_comb_d1 <= 0;
    else 
    begin
        if (READ_CLK_CTRL[2])
            DQS_GATE_CTRL_comb_d1 <= DQS_GATE_CTRL_d6;
        else if (DDC_MODE == "FULL_RATE")
            DQS_GATE_CTRL_comb_d1 <= DQS_GATE_CTRL_d2[0];
        else   
            DQS_GATE_CTRL_comb_d1 <= DQS_GATE_CTRL_d5;
    end
end

always @(negedge sel_gate_clk or negedge global_rstn or negedge lsr_rstn)
begin
    if (!global_rstn)
        DQS_GATE_CTRL_comb_d2 <= 0;
    else if (!lsr_rstn)
        DQS_GATE_CTRL_comb_d2 <= 0;
    else
        DQS_GATE_CTRL_comb_d2 <= DQS_GATE_CTRL_comb_d1;
end

assign dqs_gate_ctrl_comb = DQS_GATE_CTRL_comb_d1 & DQS_GATE_CTRL_comb_d2;

always @(negedge DQSIN_gated or negedge global_rstn or negedge lsr_rstn or posedge dqs_gate_ctrl_comb)
begin
    if (!global_rstn)
        DQS_GATE_CTRL_gate <= 1'b0;
    else if (!lsr_rstn)
        DQS_GATE_CTRL_gate <= 1'b0;
    else if (dqs_gate_ctrl_comb)
        DQS_GATE_CTRL_gate <= 1'b1;
    else
        DQS_GATE_CTRL_gate <= 1'b0;
end

assign DQSIN_gated = DQS_GATE_CTRL_gate & DQSI;
//
wire [7:0] DLL_STEP_tmp = R_DELAY_STEP_EN == "TRUE" ? DELAY_STEP1 :8'd0;
wire RDEL_CTRL_b0_tmp = R_MOVE_EN == "TRUE" ? R_LOAD_N : 1'b0;

wire [8:0] DQSI_DEL_OFFSET_tmp = DQSI_DELAY_OFFSET;

//wire [7:0] tmp_dqsi_del = DQSI_DEL_OFFSET_tmp[8] ? (DLL_STEP_tmp - DQSI_DEL_OFFSET_tmp[7:0]) : (DLL_STEP_tmp + DQSI_DEL_OFFSET_tmp[7:0]);
wire [7:0] tmp_dqsi_del = (DLL_STEP_tmp + DQSI_DEL_OFFSET_tmp[7:0]);

wire tmp_dqsi_del_co_0 = DLL_STEP_tmp[0] && DQSI_DEL_OFFSET_tmp[0];
wire tmp_dqsi_del_co_1 = (DLL_STEP_tmp[1] && DQSI_DEL_OFFSET_tmp[1]) || ((DLL_STEP_tmp[1] || DQSI_DEL_OFFSET_tmp[1]) && tmp_dqsi_del_co_0);
wire tmp_dqsi_del_co_2 = (DLL_STEP_tmp[2] && DQSI_DEL_OFFSET_tmp[2]) || ((DLL_STEP_tmp[2] || DQSI_DEL_OFFSET_tmp[2]) && tmp_dqsi_del_co_1);
wire tmp_dqsi_del_co_3 = (DLL_STEP_tmp[3] && DQSI_DEL_OFFSET_tmp[3]) || ((DLL_STEP_tmp[3] || DQSI_DEL_OFFSET_tmp[3]) && tmp_dqsi_del_co_2);
wire tmp_dqsi_del_co_4 = (DLL_STEP_tmp[4] && DQSI_DEL_OFFSET_tmp[4]) || ((DLL_STEP_tmp[4] || DQSI_DEL_OFFSET_tmp[4]) && tmp_dqsi_del_co_3); 
wire tmp_dqsi_del_co_5 = (DLL_STEP_tmp[5] && DQSI_DEL_OFFSET_tmp[5]) || ((DLL_STEP_tmp[5] || DQSI_DEL_OFFSET_tmp[5]) && tmp_dqsi_del_co_4);
wire tmp_dqsi_del_co_6 = (DLL_STEP_tmp[6] && DQSI_DEL_OFFSET_tmp[6]) || ((DLL_STEP_tmp[6] || DQSI_DEL_OFFSET_tmp[6]) && tmp_dqsi_del_co_5);
wire tmp_dqsi_del_co_7 = (DLL_STEP_tmp[7] && DQSI_DEL_OFFSET_tmp[7]) || ((DLL_STEP_tmp[7] || DQSI_DEL_OFFSET_tmp[7]) && tmp_dqsi_del_co_6);


assign tmp_dqsi_del_sel= ~(DQSI_DEL_OFFSET_tmp[8] ^ tmp_dqsi_del_co_7);
wire [7:0] adj_dly_dqsi_tmp = DQSI_DEL_OFFSET_tmp[8] ? (tmp_dqsi_del_sel ?  tmp_dqsi_del[7:0] : 8'd0) :
                              (tmp_dqsi_del_sel ? tmp_dqsi_del[7:0] : 8'd255);

always @(*) 
begin
    if (!RDEL_CTRL_b0_tmp)
        adj_dly_dqsi <= adj_dly_dqsi_tmp;
end

always @(negedge R_MOVE)
begin
    if (!RDEL_CTRL_b0_tmp)
        adj_dly_dqsi <= adj_dly_dqsi_tmp;
    else if (R_DIRECTION && (adj_dly_dqsi != 8'd0))
        adj_dly_dqsi <= adj_dly_dqsi - 1;
    else if ((~R_DIRECTION) && (adj_dly_dqsi != 8'd255))
        adj_dly_dqsi <= adj_dly_dqsi + 1;
end

assign RDELAY_OB = (R_DIRECTION && (adj_dly_dqsi == 8'd0)) || ((~R_DIRECTION) && (adj_dly_dqsi == 8'd255));

wire [255:0] dqsi_delay_chain;
assign #0.3 dqsi_delay_chain[0] = DQSIN_gated;
genvar gen_k;
generate  
    for(gen_k=1;gen_k<256;gen_k=gen_k+1) 
    begin
        assign #0.025 dqsi_delay_chain[gen_k] =  dqsi_delay_chain[gen_k-1];
    end
endgenerate

assign DQSI_DELAY = dqsi_delay_chain[adj_dly_dqsi];


assign #0.2 DQS_GATE_CTRL_gate_dly = DQS_GATE_CTRL_gate;
assign DQS_GATE_CTRL_gate_rising = DQS_GATE_CTRL_gate & (~DQS_GATE_CTRL_gate_dly);

always @(posedge DQSIN_gated or posedge DQS_GATE_CTRL_gate_rising or negedge global_rstn or negedge lsr_rstn)
begin
    if (!global_rstn)
        DQS_GATE_CTRL_gate_d <= 1'b0;
    else if (!lsr_rstn)
        DQS_GATE_CTRL_gate_d <= 1'b0;
    else if (DQS_GATE_CTRL_gate_rising)
        DQS_GATE_CTRL_gate_d <= 1'b0;
    else if (DQS_GATE_CTRL_gate) 
    begin
        DQS_GATE_CTRL_gate_d[0] <= ~ DQS_GATE_CTRL_gate_d[0];
        DQS_GATE_CTRL_gate_d[1] <= DQS_GATE_CTRL_gate_d[0];
    end
end

always @(negedge DQSIN_gated or posedge DQS_GATE_CTRL_gate_rising or negedge global_rstn or negedge lsr_rstn)
begin
    if (!global_rstn)
        DQS_GATE_CTRL_gate_dd <= 1'b0;
    else if (!lsr_rstn)
        DQS_GATE_CTRL_gate_dd <= 1'b0;
    else if (DQS_GATE_CTRL_gate_rising)
        DQS_GATE_CTRL_gate_dd <= 1'b0;
    else if (DQS_GATE_CTRL_gate) 
    begin
        DQS_GATE_CTRL_gate_dd[0] <= ~ DQS_GATE_CTRL_gate_dd[0];
        DQS_GATE_CTRL_gate_dd[1] <= DQS_GATE_CTRL_gate_dd[0];
    end
end

always @(negedge DQSI_DELAY or posedge DQS_GATE_CTRL_gate_rising or negedge global_rstn or negedge lsr_rstn)
begin
    if (!global_rstn)
        DQS_GATE_CTRL_comb_and_d <= 1'b0;
    else if (!lsr_rstn)
        DQS_GATE_CTRL_comb_and_d <= 1'b0;
    else if (DQS_GATE_CTRL_gate_rising)
        DQS_GATE_CTRL_comb_and_d <= 1'b0;
    else if (dqs_gate_ctrl_comb) 
    begin
        DQS_GATE_CTRL_comb_and_d[0] <= ~ DQS_GATE_CTRL_comb_and_d[0];
        DQS_GATE_CTRL_comb_and_d[1] <= DQS_GATE_CTRL_comb_and_d[0];
    end
end

assign DGTS_a = (~DQS_GATE_CTRL_gate) && (DQS_GATE_CTRL_gate_d == 2'b10);
assign DGTS_b = (DQS_GATE_CTRL_gate_dd == 2'b10) &&  (DQS_GATE_CTRL_comb_and_d == 2'b01);

assign DGTS = DGTS_a & DGTS_b;


always @(posedge DQSI_DELAY or negedge rstn_fifo)
begin
    if (!rstn_fifo)
        start_wr <= 0;
    else
        start_wr <= rstn_fifo;
end

assign start_wr_comb = (IFIFO_GENERIC == "TRUE") ?  start_wr : rstn_fifo;

always @(posedge DQSI_DELAY or negedge start_wr_comb)
begin
    if (!start_wr_comb)
        WADDR_reg <= 0;
    else 
    begin
        case (WADDR_reg)
            3'b000: WADDR_reg <= 3'b001;
            3'b001: WADDR_reg <= 3'b011;
            3'b011: WADDR_reg <= 3'b010;
            3'b010: WADDR_reg <= 3'b110;
            3'b110: WADDR_reg <= 3'b111;
            3'b111: WADDR_reg <= 3'b101;
            3'b101: WADDR_reg <= 3'b100;
            3'b100: WADDR_reg <= 3'b000;
        endcase
    end
end

always @(negedge DQSI_DELAY or negedge start_wr_comb)
begin
    if (!start_wr_comb)
        IFIFO_WADDR_reg <= 0;
    else
        IFIFO_WADDR_reg <= WADDR_reg;
end

assign IFIFO_WADDR = IFIFO_WADDR_reg;

assign rd_clk = (DDC_MODE == "FULL_RATE") ? CLKB : CLKA;

always @(posedge rd_clk or negedge rstn_fifo)
begin
    if (!rstn_fifo)
        start_rd <= 0;
    else
        start_rd <= rstn_fifo;
end

always @(posedge rd_clk or negedge rst_start_rd)
begin
    if (!rst_start_rd)
        WADDR_reg_d1 <= 3'd0;
    else
        WADDR_reg_d1 <= WADDR_reg;
end

always @(posedge rd_clk or negedge rst_start_rd)
begin
    if (!rst_start_rd)
        WADDR_reg_d2 <= 3'd0;
    else
        WADDR_reg_d2 <= WADDR_reg_d1;
end

assign buffer_empty = WADDR_reg_d2 == RADDR_reg;
assign buffer_almost_empty = WADDR_reg_d2 == RADDR_reg_plus1;


always @(posedge rd_clk or negedge rstn_fifo)
begin
    if (!rstn_fifo) 
    begin
        new_st         <= 0;
        new_cnt        <= 0;
        new_transfer_d <= 0;
    end
    else 
    begin
        new_st       <= 1;
        if (new_st)
            new_cnt      <= new_cnt + 1;
            new_transfer_d <= new_transfer;
    end
end

assign  new_transfer =  (DDC_MODE == "HALF_RATE") ? new_cnt[0] : (new_cnt == 2);

always @(posedge rd_clk or negedge rst_start_rd)
begin
    if (!rst_start_rd) 
    begin
        new_rd_en_reg <= 0;
    end
    else if ((DDC_MODE == "FULL_RATE") || new_transfer) 
    begin //sel port
        if (new_rd_en_reg) 
        begin
            if (buffer_almost_empty)
                new_rd_en_reg <= 1'b0;
        end
        else 
        begin
            if (~buffer_empty)
                new_rd_en_reg <= 1'b1;
        end
    end
end

wire read_enable = (new_rd_en_reg && (~buffer_empty)) || (IFIFO_GENERIC == "TRUE");

wire start_generic_read = (IFIFO_GENERIC == "TRUE") ? new_st : (~buffer_empty);


always @(posedge rd_clk or negedge rst_start_rd)
begin
    if (!rst_start_rd)
        RADDR_reg <= RADDR_INIT;
    else if (read_enable && start_generic_read) 
    begin
        case (RADDR_reg)
            3'b000: RADDR_reg <= 3'b001;
            3'b001: RADDR_reg <= 3'b011;
            3'b011: RADDR_reg <= 3'b010;
            3'b010: RADDR_reg <= 3'b110;
            3'b110: RADDR_reg <= 3'b111;
            3'b111: RADDR_reg <= 3'b101;
            3'b101: RADDR_reg <= 3'b100;
            3'b100: RADDR_reg <= 3'b000;
        endcase
    end
end

always @(*) 
begin
    case (RADDR_reg)
        3'b000: RADDR_reg_plus1 <= 3'b001;
        3'b001: RADDR_reg_plus1 <= 3'b011;
        3'b011: RADDR_reg_plus1 <= 3'b010;
        3'b010: RADDR_reg_plus1 <= 3'b110;
        3'b110: RADDR_reg_plus1 <= 3'b111;
        3'b111: RADDR_reg_plus1 <= 3'b101;
        3'b101: RADDR_reg_plus1 <= 3'b100;
        3'b100: RADDR_reg_plus1 <= 3'b000;
    endcase
end

assign IFIFO_RADDR = RADDR_reg;

always @(posedge rd_clk or negedge rst_start_rd)
begin
    if (!rst_start_rd) 
    begin
        read_enable_d1 <= 0;
        read_enable_d2 <= 0;
    end
    else 
    begin
        read_enable_d1 <= (new_rd_en_reg && (~buffer_empty));
        if (new_transfer_d)
            read_enable_d2 <= read_enable_d1;
    end
end

always @(posedge CLKB or negedge rst_start_rd)
begin
    if (!rst_start_rd)
        RDVALID_reg <= 0;
    else if (DDC_MODE == "FULL_RATE") 
    begin
        if (IFIFO_GENERIC == "TRUE")
            RDVALID_reg <= 1'b1;
        else
            RDVALID_reg <=  (new_rd_en_reg && (~buffer_empty));
    end
    else 
        RDVALID_reg <= read_enable_d2;
end

assign READ_VALID = RDVALID_reg;
//synthesis translate_on

endmodule





































//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_PREADD_MULT9.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

//P = A*(B+C)
`timescale 1 ns / 1 ps

module GTP_PREADD_MULT9 #(
    parameter GRS_EN      = "TRUE", //"TRUE"; "FALSE"
    parameter SYNC_RST    = "FALSE", //"TRUE"; "FALSE"
    parameter INREG_EN    = "FALSE",  //"TRUE"; "FALSE"
    parameter PREREG_EN   = "FALSE",  //"TRUE"; "FALSE"
    parameter OUTREG_EN   = "FALSE"    //"TRUE"; "FALSE"
)(
    output  [18-1:0] P,
    input   CE,
    input   RST,
    input   CLK,
    input   A_SIGNED,
    input   [9-1:0] A,
    input   B_SIGNED,
    input   [8-1:0] B,
    input   C_SIGNED,
    input   [8-1:0] C,
    input   PREADDSUB
);

    INT_PREADD_MULT  #(.GRS_EN(GRS_EN),
        .SYNC_RST(SYNC_RST),    
        .INREG_EN(INREG_EN),    
        .PREREG_EN(PREREG_EN),    
        .OUTREG_EN(OUTREG_EN),   
        .ASIZE(9),  
        .BSIZE(8)
    )  U_INT_PREADD_MULT (
        .CE(CE),
        .RST(RST),
        .CLK(CLK),
        .A_SIGNED(A_SIGNED),
        .A(A),
        .B_SIGNED(B_SIGNED),
        .B(B),
        .C_SIGNED(C_SIGNED),
        .C(C),
        .PREADDSUB(PREADDSUB),
        .P(P)
    );

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_DFF_S.v
//
// Functional description: D-type flip-flop with sync set
//
// Parameter description:
//      INIT: init value
//
// Port description:
//      S: synchronous set
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_DFF_S
#(
    parameter GRS_EN = "TRUE",
    parameter INIT = 1'b1
) (
    output reg Q,
    input wire D,
    input wire CLK, S
);

    wire grs_n;
    wire RS;

    tri1 grsnet = GRS_INST.GRSNET;
    assign grs_n=(GRS_EN=="TRUE")?grsnet:1'b1;

    not (RS, grs_n);

    initial Q = 1'bx;

    always @(posedge CLK or posedge RS) begin
        if (RS)
            Q <= 1'b1;
        else if (S)
            Q <= 1'b1;
        else
            Q <= D;
    end

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_DLATCH_P.v
//
// Functional description: D-type latch with set
//
// Parameter description:
//      INIT: init value
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_DLATCH_P
#(
    parameter GRS_EN = "TRUE",
    parameter INIT = 1'b1
) (
    output reg Q,
    input wire D,
    input wire G, P
);

    wire grs_n;
    wire grs, RS;

    tri1 grsnet = GRS_INST.GRSNET;
    assign grs_n=(GRS_EN=="TRUE")?grsnet:1'b1;

    not (grs, grs_n);
    or (RS, grs, P);

    initial Q = 1'bx;

    always @(D or G or RS) begin
        if (RS)
            Q <= 1'b1;
        else if (G)
            Q <= D;
    end

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_OUTBUFTDS.v
//
// Functional description: Differential Signaling Tristate Output Buffer
//
// Parameter description:
//      
//
// Port description:
//
// Revision:
//    06/18/14 - Initial version.
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_OUTBUFTDS #(
    parameter IOSTANDARD = "DEFAULT"
)(
    output O,
    output OB,
    input I,
    input T
) /* synthesis syn_black_box */ ;
  
  initial begin
    case (IOSTANDARD)
    "LVDS", "MINI-LVDS", "SUB-LVDS","TMDS", "DEFAULT" :;
    default : begin
           $display("Attribute Syntax Error : The attribute IOSTANDARD on GTP_OUTBUFTDS instance %m is set to %s.", IOSTANDARD);
           $finish;
              end
    endcase
    end
    bufif0 (O, I, T);
    notif0 (OB, I, T);

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_DLATCH_PE.v
//
// Functional description: D-type latch with set and enable
//
// Parameter description:
//      INIT: init value
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_DLATCH_PE
#(
    parameter GRS_EN = "TRUE",
    parameter INIT = 1'b1
) (
    output reg Q,
    input wire D,
    input wire G, P, GE
);

    wire grs_n;
    wire grs, RS;

    tri1 grsnet = GRS_INST.GRSNET;
    assign grs_n=(GRS_EN=="TRUE")?grsnet:1'b1;

    not (grs, grs_n);
    or (RS, grs, P);

    initial Q = 1'bx;

    always @(D or G or RS or GE) begin
        if (RS)
            Q <= 1'b1;
        else if (G && GE)
            Q <= D;
    end

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_PREADD_MULTADD9.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

//P = A0*(B0+-C0) +/- A1*(B1+-C1)
`timescale 1 ns / 1 ps

module GTP_PREADD_MULTADD9 #(
    parameter GRS_EN           = "TRUE", //"TRUE"; "FALSE"
    parameter SYNC_RST         = "FALSE", //"TRUE"; "FALSE"  
    parameter INREG_EN         = "FALSE", //"TRUE"; "FALSE"
    parameter PREREG_EN        = "FALSE", //"TRUE"; "FALSE"
    parameter PIPEREG_EN       = "FALSE", //"TRUE"; "FALSE"
    parameter OUTREG_EN        = "FALSE", //"TRUE"; "FALSE"
    parameter ADDSUB_OP        = 0 ,
    parameter DYN_ADDSUB_OP    = 1
)(
    output  [19-1:0] P,
    input   CE,
    input   RST,
    input   CLK,
    input   [9-1:0] A0,
    input   [9-1:0] A1,
    input   [8-1:0] B0,
    input   [8-1:0] B1,
    input   [8-1:0] C0,
    input   [8-1:0] C1,
    input   A_SIGNED,
    input   B_SIGNED,
    input   C_SIGNED,
    input   [1:0] PREADDSUB,
    input   ADDSUB
);


    INT_PREADD_MULTADD #(
        . GRS_EN(GRS_EN),    
        . SYNC_RST(SYNC_RST),  
        . INREG_EN(INREG_EN), 
        . PREREG_EN(PREREG_EN), 
        . PIPEREG_EN(PIPEREG_EN),
        . OUTREG_EN(OUTREG_EN), 
        . ADDSUB_OP(ADDSUB_OP),   
        . DYN_OP_ADDSUB(DYN_ADDSUB_OP),
        . ASIZE(9), 
        . BSIZE(8)
    ) U_INT_PREADD_MULTADD(
        . CE(CE),
        . RST(RST),
        . CLK(CLK),
        . A0(A0),
        . A1(A1),
        . B0(B0),
        . B1(B1),
        . C0(C0),
        . C1(C1),
        . A_SIGNED(A_SIGNED),
        . B_SIGNED(B_SIGNED),
        . C_SIGNED(C_SIGNED),
        . PREADDSUB(PREADDSUB),
        . ADDSUB(ADDSUB),
        . P(P)
    );   

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_MULTADD9.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

//P = A0*B0 +/- A1*B1
module GTP_MULTADD9 #(
    parameter GRS_EN        = "TRUE", //"TRUE"; "FALSE"
    parameter SYNC_RST      = "FALSE", //"TRUE"; "FALSE"
    parameter INREG_EN      = "FALSE",  //"TRUE"; "FALSE"
    parameter PIPEREG_EN    = "FALSE",  //"TRUE"; "FALSE"
    parameter OUTREG_EN     = "FALSE",  //"TRUE"; "FALSE"
    parameter ADDSUB_OP     = 0 ,
    parameter DYN_ADDSUB_OP = 1
)(
    output  [19-1:0] P,          //product
    input   CE,
    input   RST,
    input   CLK,
    input   A_SIGNED,
    input   [9-1:0] A0,
    input   [9-1:0] A1,
    input   B_SIGNED,
    input   [9-1:0] B0,
    input   [9-1:0] B1,
    input   ADDSUB
);

    INT_PREADD_MULTADD #(
        . GRS_EN(GRS_EN),
        . SYNC_RST(SYNC_RST),   
        . INREG_EN(INREG_EN),   
        . PIPEREG_EN(PIPEREG_EN), 
        . OUTREG_EN(OUTREG_EN),  
        . ADDSUB_OP(ADDSUB_OP),  
        . DYN_OP_ADDSUB(DYN_ADDSUB_OP), 
        . ASIZE(9), 
        . BSIZE(9),
        . PREADD_EN(0)
    ) U_MULTADD9 (
        . CE(CE),
        . RST(RST),
        . CLK(CLK),
        . A_SIGNED(A_SIGNED),
        . A0(A0),
        . A1(A1),
        . B_SIGNED(B_SIGNED),
        . B0(B0),
        . B1(B1),
        . C_SIGNED(B_SIGNED),
        . C0(9'b0),
        . C1(9'b0),
        . PREADDSUB(2'b0),
        . ADDSUB(ADDSUB),
        . P(P)
    );

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_TIMER.v
//
// Functional description: Timer Circuit
//
// Parameter description:
//      
//
// Port description:
//      
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////


`timescale 1 ns / 1 ps
module GTP_TIMER
(
input         RST_N,
input         CLK,
input         STAMP,
output        PWM,
output        IRQ
);

assign  GTP_GRS.timer_rstn  = RST_N;
assign  GTP_GRS.timer_clk   = CLK;
assign  GTP_GRS.timer_stamp = STAMP;
assign  PWM = GTP_GRS.timer_pwm;
assign  IRQ = GTP_GRS.irq_timer;

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2016 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_RAM128X1DP.v
//
// Functional description: simple-dual-port 128x1 distributed ram
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_RAM128X1DP
#(
    parameter [127:0] INIT = 128'h0000_0000_0000_0000_0000_0000_0000_0000
) (
    output  DO,
    input   DI,
    input [6:0] RADDR,
    input [6:0] WADDR,
    input WCLK,
    input WE
);
//synthesis translate_off
    reg [127:0] mem ;

    initial begin
        mem = INIT;
    end

    always @(posedge WCLK) begin
        if (WE == 1'b1) begin
            mem[WADDR] <= DI;
        end
    end

    assign DO = mem[RADDR];
//synthesis translate_on
endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2019 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_PPLL.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1ns/10fs
module GTP_PPLL #(
    parameter real CLKIN_FREQ = 50.0,    //19MHz~800MHz
    parameter LOCK_MODE       = 1'b0,    //1'b0~1'b1
    parameter integer STATIC_RATIOI   = 1, //1~128
    parameter integer STATIC_RATIOM   = 1, //1~128
    parameter integer STATIC_RATIO0   = 1, //1~128
    parameter integer STATIC_RATIO1   = 1, //1~128
    parameter integer STATIC_RATIO2   = 1, //1~128
    parameter integer STATIC_RATIO3   = 1, //1~128
    parameter integer STATIC_RATIO4   = 1, //1~128
    parameter integer STATIC_RATIOPHY = 1, //1~128
    parameter integer STATIC_RATIOF   = 1, //1~128
    parameter integer STATIC_DUTY0   = 2, //2<=STATIC_DUTY0<=2*STATIC_RATIO0-1
    parameter integer STATIC_DUTY1   = 2, //2<=STATIC_DUTY1<=2*STATIC_RATIO1-1
    parameter integer STATIC_DUTY2   = 2, //2<=STATIC_DUTY2<=2*STATIC_RATIO2-1
    parameter integer STATIC_DUTY3   = 2, //2<=STATIC_DUTY3<=2*STATIC_RATIO3-1
    parameter integer STATIC_DUTY4   = 2, //2<=STATIC_DUTY4<=2*STATIC_RATIO4-1
    parameter integer STATIC_DUTYPHY = 2, //2<=STATIC_DUTY5<=2*STATIC_RATIO5-1
    parameter integer STATIC_DUTYF   = 2, //2<=STATIC_DUTYF<=2*STATIC_RATIOF-1
    parameter integer STATIC_PHASE0   = 0, //0~7
    parameter integer STATIC_PHASE1   = 0, //0~7
    parameter integer STATIC_PHASE2   = 0, //0~7
    parameter integer STATIC_PHASE3   = 0, //0~7
    parameter integer STATIC_PHASE4   = 0, //0~7
    parameter integer STATIC_PHASEPHY = 0, //0~7
    parameter integer STATIC_PHASEF    = 0, //0~7
    parameter integer STATIC_CPHASE0   = 0, //0~127
    parameter integer STATIC_CPHASE1   = 0, //0~127
    parameter integer STATIC_CPHASE2   = 0, //0~127
    parameter integer STATIC_CPHASE3   = 0, //0~127
    parameter integer STATIC_CPHASE4   = 0, //0~127
    parameter integer STATIC_CPHASEPHY = 0, //0~127
    parameter integer STATIC_CPHASEF   = 0, //0~127
    parameter CLKOUT0_SYN_EN   = "FALSE", //"TRUE"; "FALSE"
    parameter CLKOUT1_SYN_EN   = "FALSE", //"TRUE"; "FALSE"
    parameter CLKOUT2_SYN_EN   = "FALSE", //"TRUE"; "FALSE"
    parameter CLKOUT3_SYN_EN   = "FALSE", //"TRUE"; "FALSE"
    parameter CLKOUT4_SYN_EN   = "FALSE", //"TRUE"; "FALSE"
    parameter CLKOUTPHY_SYN_EN = "FALSE", //"TRUE"; "FALSE"
    parameter CLKOUTF_SYN_EN   = "FALSE", //"TRUE"; "FALSE"
    parameter INTERNAL_FB = "CLKOUTF",  //"CLKOUT0"; "CLKOUT1"; "CLKOUT2"; "CLKOUT3"; "CLKOUT4"; "CLKOUTF"; "DISABLE";
    parameter EXTERNAL_FB = "DISABLE",  //"CLKOUT0"; "CLKOUT1"; "CLKOUT2"; "CLKOUT3"; "CLKOUT4"; "CLKOUTF"; "DISABLE";
    parameter BANDWIDTH   = "OPTIMIZED" //"LOW"; "OPTIMIZED"; "HIGH"
    )(
    output CLKOUT0,
    output CLKOUT0N,
    output CLKOUT1,
    output CLKOUT1N,
    output CLKOUT2,
    output CLKOUT2N,
    output CLKOUT3,
    output CLKOUT3N,
    output CLKOUT4,
    output CLKOUTPHY,
    output CLKOUTPHYN,
    output CLKOUTF,
    output CLKOUTFN,
    output LOCK,
    output [15:0] APB_RDATA,
    output APB_READY,
    input CLKIN1,
    input CLKIN2,
    input CLKFB,
    input CLKIN_SEL,
    input CLKOUT0_SYN,
    input CLKOUT1_SYN,
    input CLKOUT2_SYN,
    input CLKOUT3_SYN,
    input CLKOUT4_SYN,
    input CLKOUTPHY_SYN,
    input CLKOUTF_SYN,
    input PLL_PWD,
    input RST,
    input APB_CLK,
    input APB_RST_N,
    input [4:0] APB_ADDR,
    input APB_SEL,
    input APB_EN,
    input APB_WRITE,
    input [15:0] APB_WDATA
    );

    initial
    begin
        if((CLKOUT0_SYN_EN == "TRUE") || (CLKOUT0_SYN_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PPLL error: illegal setting for CLKOUT0_SYN_EN");

        if((CLKOUT1_SYN_EN == "TRUE") || (CLKOUT1_SYN_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PPLL error: illegal setting for CLKOUT1_SYN_EN");

        if((CLKOUT2_SYN_EN == "TRUE") || (CLKOUT2_SYN_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PPLL error: illegal setting for CLKOUT2_SYN_EN");

        if((CLKOUT3_SYN_EN == "TRUE") || (CLKOUT3_SYN_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PPLL error: illegal setting for CLKOUT3_SYN_EN");

        if((CLKOUT4_SYN_EN == "TRUE") || (CLKOUT4_SYN_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PPLL error: illegal setting for CLKOUT4_SYN_EN");

        if((CLKOUTPHY_SYN_EN == "TRUE") || (CLKOUTPHY_SYN_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PPLL error: illegal setting for CLKOUTPHY_SYN_EN");

        if((CLKOUTF_SYN_EN == "TRUE") || (CLKOUTF_SYN_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PPLL error: illegal setting for CLKOUTF_SYN_EN");

        if((INTERNAL_FB == "CLKOUT0") || (INTERNAL_FB == "CLKOUT1") || (INTERNAL_FB == "CLKOUT2") || (INTERNAL_FB == "CLKOUT3") || (INTERNAL_FB == "CLKOUT4") || (INTERNAL_FB == "CLKOUTF") || (INTERNAL_FB == "DISABLE"))
        begin
        end
        else
            $display ("GTP_PPLL error: illegal setting for INTERNAL_FB");

        if((EXTERNAL_FB == "CLKOUT0") || (EXTERNAL_FB == "CLKOUT1") || (EXTERNAL_FB == "CLKOUT2") || (EXTERNAL_FB == "CLKOUT3") || (EXTERNAL_FB == "CLKOUT4") || (EXTERNAL_FB == "CLKOUTF") || (EXTERNAL_FB == "DISABLE"))
        begin
        end
        else
            $display ("GTP_PPLL error: illegal setting for EXTERNAL_FB");

        if((BANDWIDTH == "LOW") || (BANDWIDTH == "OPTIMIZED") || (BANDWIDTH == "HIGH"))
        begin
        end
        else
            $display ("GTP_PPLL error: illegal setting for BANDWIDTH");
    end
///////////////////////////////////////////////////////
////INITIAL////////////////////////////////////////////
    reg [7:0] ratioi_i, ratiom_i, ratiof_i, ratio0_i, ratio1_i, ratio2_i, ratio3_i, ratio4_i, ratiophy_i;
    reg [7:0] dutyf_i, duty0_i, duty1_i, duty2_i, duty3_i, duty4_i, dutyphy_i;
    reg [6:0] odiv0_cphase_i, odiv1_cphase_i, odiv2_cphase_i, odiv3_cphase_i, odiv4_cphase_i, odivphy_cphase_i, fdiv_cphase_i;
    reg [2:0] odiv0_fphase_i, odiv1_fphase_i, odiv2_fphase_i, odiv3_fphase_i, odiv4_fphase_i, odivphy_fphase_i, fdiv_fphase_i;

    reg muxsel0_en_i, muxsel1_en_i, muxsel2_en_i, muxsel3_en_i, muxsel4_en_i, muxselphy_en_i, muxself_en_i;

    reg [15:0] mem0, mem1, mem2, mem3, mem4, mem5, mem6, mem7, mem8, mem9, mem10, mem11, mem12, mem13, mem14, mem15, mem16, mem17;
    reg [1:0] vctrl_i;
    reg [1:0] cp_selbias_i, cp_base_i;
    reg [3:0] cp_cur_i;
    reg [2:0] lpf_r_i;
    reg lpf_c_i;
    reg [5:0] lock_set_i;
    reg lockfilter_pd_i;

    wire [7:0] ratioi, ratiom, ratiof, ratio0, ratio1, ratio2, ratio3, ratio4, ratiophy;
    wire [7:0] dutyf, duty0, duty1, duty2, duty3, duty4, dutyphy;
    wire [6:0] odiv0_cphase, odiv1_cphase, odiv2_cphase, odiv3_cphase, odiv4_cphase, odivphy_cphase, fdiv_cphase;
    wire [2:0] odiv0_fphase, odiv1_fphase, odiv2_fphase, odiv3_fphase, odiv4_fphase, odivphy_fphase, fdiv_fphase;

    initial
    begin
        ratioi_i   = STATIC_RATIOI;
        ratiom_i   = STATIC_RATIOM;
        ratiof_i   = STATIC_RATIOF;
        ratio0_i   = STATIC_RATIO0;
        ratio1_i   = STATIC_RATIO1;
        ratio2_i   = STATIC_RATIO2;
        ratio3_i   = STATIC_RATIO3;
        ratio4_i   = STATIC_RATIO4;
        ratiophy_i = STATIC_RATIOPHY;
        dutyf_i    = STATIC_DUTYF;
        duty0_i    = STATIC_DUTY0;
        duty1_i    = STATIC_DUTY1;
        duty2_i    = STATIC_DUTY2;
        duty3_i    = STATIC_DUTY3;
        duty4_i    = STATIC_DUTY4;
        dutyphy_i  = STATIC_DUTYPHY;
        odiv0_cphase_i   = STATIC_CPHASE0;
        odiv1_cphase_i   = STATIC_CPHASE1;
        odiv2_cphase_i   = STATIC_CPHASE2;
        odiv3_cphase_i   = STATIC_CPHASE3;
        odiv4_cphase_i   = STATIC_CPHASE4;
        odivphy_cphase_i = STATIC_CPHASEPHY;
        fdiv_cphase_i    = STATIC_CPHASEF;
        odiv0_fphase_i   = STATIC_PHASE0;
        odiv1_fphase_i   = STATIC_PHASE1;
        odiv2_fphase_i   = STATIC_PHASE2;
        odiv3_fphase_i   = STATIC_PHASE3;
        odiv4_fphase_i   = STATIC_PHASE4;
        odivphy_fphase_i = STATIC_PHASEPHY;
        fdiv_fphase_i    = STATIC_PHASEF;
        muxsel0_en_i   = 1'b1;
        muxsel1_en_i   = 1'b1;
        muxsel2_en_i   = 1'b1;
        muxsel3_en_i   = 1'b1;
        muxsel4_en_i   = 1'b1;
        muxselphy_en_i = 1'b1;
        muxself_en_i   = 1'b1;
        vctrl_i        = 2'b00;
        cp_selbias_i   = 2'b01;
        cp_base_i      = 2'b10;
        cp_cur_i       = 4'b0001;
        lpf_r_i        = 3'b001;
        lpf_c_i        = 1'b0;
        lock_set_i      = 5'h0;
        lockfilter_pd_i = 1'b1;

        mem0  = {ratio0_i, duty0_i};
        mem1  = {5'h0, muxsel0_en_i, odiv0_fphase_i, odiv0_cphase_i};
        mem2  = {ratio1_i, duty1_i};
        mem3  = {5'h0, muxsel1_en_i, odiv1_fphase_i, odiv1_cphase_i};
        mem4  = {ratio2_i, duty2_i};
        mem5  = {5'h0, muxsel2_en_i, odiv2_fphase_i, odiv2_cphase_i};
        mem6  = {ratio3_i, duty3_i};
        mem7  = {5'h0, muxsel3_en_i, odiv3_fphase_i, odiv3_cphase_i};
        mem8  = {ratio4_i, duty4_i};
        mem9  = {5'h0, muxsel4_en_i, odiv4_fphase_i, odiv4_cphase_i};
        mem10 = {ratiophy_i, dutyphy_i};
        mem11 = {5'h0, muxselphy_en_i, odivphy_fphase_i, odivphy_cphase_i};
        mem12 = {ratiof_i, dutyf_i};
        mem13 = {5'h0, muxself_en_i, fdiv_fphase_i, fdiv_cphase_i};
        mem14 = {8'h0, ratioi_i};
        mem15 = {8'h0, ratiom_i};
        mem16 = {2'b00, vctrl_i, cp_selbias_i, cp_base_i, cp_cur_i, lpf_r_i, lpf_c_i};
        mem17 = {10'h0, lockfilter_pd_i, lock_set_i};
    end

    assign ratioi   = mem14[7:0];
    assign ratiom   = mem15[7:0];
    assign ratiof   = mem12[15:8];
    assign ratio0   = mem0[15:8];
    assign ratio1   = mem2[15:8];
    assign ratio2   = mem4[15:8];
    assign ratio3   = mem6[15:8];
    assign ratio4   = mem8[15:8];
    assign ratiophy = mem10[15:8];
    assign dutyf    = mem12[7:0];
    assign duty0    = mem0[7:0];
    assign duty1    = mem2[7:0];
    assign duty2    = mem4[7:0];
    assign duty3    = mem6[7:0];
    assign duty4    = mem8[7:0];
    assign dutyphy  = mem10[7:0];
    assign odiv0_cphase   = mem1[6:0];
    assign odiv1_cphase   = mem3[6:0];
    assign odiv2_cphase   = mem5[6:0];
    assign odiv3_cphase   = mem7[6:0];
    assign odiv4_cphase   = mem9[6:0];
    assign odivphy_cphase = mem11[6:0];
    assign fdiv_cphase    = mem13[6:0];
    assign odiv0_fphase   = mem1[9:7];
    assign odiv1_fphase   = mem3[9:7];
    assign odiv2_fphase   = mem5[9:7];
    assign odiv3_fphase   = mem7[9:7];
    assign odiv4_fphase   = mem9[9:7];
    assign odivphy_fphase = mem11[9:7];
    assign fdiv_fphase    = mem13[9:7];
    assign muxsel0_en   = mem1[10];
    assign muxsel1_en   = mem3[10];
    assign muxsel2_en   = mem5[10];
    assign muxsel3_en   = mem7[10];
    assign muxsel4_en   = mem9[10];
    assign muxselphy_en = mem11[10];
    assign muxself_en   = mem13[10];
///////////////////////////////////////////////////////
    wire rst_n;
    reg inner_rstn;
///////////////////////////////////////////////////////
    wire clk_in;
///////////////////////////////////////////////////////
    reg clk_in_first_time, clk_fb_first_time;
    realtime clk_in_first_edge, clk_fb_first_edge;
    reg adjust;
    realtime fb_route_delay, virtual_delay1;
    integer tmp_ratio;
    realtime tmp_delay, real_delay;
///////////////////////////////////////////////////////
    reg clk_test;
    reg clkref_wo, clkfb_wo;
    realtime clkref_test_time1 , clkref_test_time2, clkref_test_time3;
    realtime clkfb_rtime_last, clkfb_rtime_next;
    realtime clkfb_test_time1 , clkfb_test_time2, clkfb_test_time3;
    wire clkwo;
///////////////////////////////////////////////////////
    wire [7:0] idivider, mdivider, fdivider, divider0, divider1, divider2, divider3, divider4, dividerphy;
    real fsdiv_set_int, fbdiv_set_int;

    wire rstanalog_n;
    realtime clkin_rtime_last, clkin_rtime_next;
    realtime clkin_time, clkin_time1, clkin_time2, clkin_time3;
    reg clkout_lock;
    realtime vcoclk_period, vcoclk_period_half;
    realtime clkout0_time, clkout1_time, clkout2_time, clkout3_time, clkout4_time, clkoutphy_time, clkoutf_time;
    integer  vcoclk_period_amp;
    realtime vcoclk_period_real, vcoclk_period_dev;

    reg done;
    integer idiv_set;
    integer fdiv_set;
    integer swap_set;
    integer midd_set;
    integer fdiv_int;
    realtime offset;

    real cnt_fdiv;
    reg clk_gate, inner_clk;
    reg vcoclk;
///////////////////////////////////////////////////////
    wire clk_lock;
    reg [2:0] cnt_clkfb;
    reg start_clk;
    reg [10:0] cnt_lock;
    reg lock_wait;
    reg lock_reg;
///////////////////////////////////////////////////////
    wire odiv0_clkin, odiv1_clkin, odiv2_clkin, odiv3_clkin, odiv4_clkin, odivphy_clkin, fdiv_clkin;
    reg [7:0] odiv0_counter, odiv1_counter, odiv2_counter, odiv3_counter, odiv4_counter, odivphy_counter, fdiv_counter;
    reg odiv0_out_reg, odiv1_out_reg, odiv2_out_reg, odiv3_out_reg, odiv4_out_reg, odivphy_out_reg, fdiv_out_reg;
    wire odiv0_out, odiv1_out, odiv2_out, odiv3_out, odiv4_out, odivphy_out, fdiv_out;
///////////////////////////////////////////////////////
    realtime vco_fphase_delay0, vco_fphase_delay1, vco_fphase_delay2, vco_fphase_delay3, vco_fphase_delay4, vco_fphase_delayphy, vco_fphase_delayf;
    integer cphase0, cphase1, cphase2, cphase3, cphase4, cphasephy, cphasef;
    realtime cphase_delay0, cphase_delay1, cphase_delay2, cphase_delay3, cphase_delay4, cphase_delayphy, cphase_delayf;
    reg odiv0_out_delay1, odiv1_out_delay1, odiv2_out_delay1, odiv3_out_delay1, odiv4_out_delay1, odivphy_out_delay1, fdiv_out_delay1;
    reg odiv0_out_delay, odiv1_out_delay, odiv2_out_delay, odiv3_out_delay, odiv4_out_delay, odivphy_out_delay, fdiv_out_delay;
///////////////////////////////////////////////////////
    reg [2:0] clk_out0_gate, clk_out1_gate, clk_out2_gate, clk_out3_gate, clk_out4_gate, clk_outphy_gate, clk_outf_gate;
    wire clkout0_gate, clkout1_gate, clkout2_gate, clkout3_gate, clkout4_gate, clkoutphy_gate, clkoutf_gate;
///////////////////////////////////////////////////////
    reg [1:0] apb_rstn_sync;
    reg ready;
    reg [15:0] rdata;
///////////////////////////////////////////////////////
    initial
    begin
        inner_rstn = 1'b0;
        clk_in_first_time = 1'b0;
        clk_fb_first_time = 1'b0;
        clk_in_first_edge = 0.0;
        clk_fb_first_edge = 0.0;
        fb_route_delay = 0.0;
        tmp_ratio      = 0;
        tmp_delay      = 0.0;
        real_delay     = 0.0;
        clk_test = 1'b0;
        fsdiv_set_int = 0;
        fbdiv_set_int = 0;
        done = 1'b0;
        idiv_set = 0;
        fdiv_set = 0;
        swap_set = 0;
        midd_set = 0;
        fdiv_int = 0;
        offset = 0;
        cnt_fdiv  = 0;
        clk_gate  = 1'b1;
        inner_clk = 1'b0;
        vcoclk    = 1'b0;
        vco_fphase_delay0   = 0.0;
        vco_fphase_delay1   = 0.0;
        vco_fphase_delay2   = 0.0;
        vco_fphase_delay3   = 0.0;
        vco_fphase_delay4   = 0.0;
        vco_fphase_delayphy = 0.0;
        vco_fphase_delayf   = 0.0;
        cphase_delay0   = 0.0;
        cphase_delay1   = 0.0;
        cphase_delay2   = 0.0;
        cphase_delay3   = 0.0;
        cphase_delay4   = 0.0;
        cphase_delayphy = 0.0;
        cphase_delayf   = 0.0;
        odiv0_out_delay1   = 1'b0;
        odiv1_out_delay1   = 1'b0;
        odiv2_out_delay1   = 1'b0;
        odiv3_out_delay1   = 1'b0;
        odiv4_out_delay1   = 1'b0;
        odivphy_out_delay1 = 1'b0;
        fdiv_out_delay1    = 1'b0;
        odiv0_out_delay    = 1'b0;
        odiv1_out_delay    = 1'b0;
        odiv2_out_delay    = 1'b0;
        odiv3_out_delay    = 1'b0;
        odiv4_out_delay    = 1'b0;
        odivphy_out_delay  = 1'b0;
        fdiv_out_delay     = 1'b0;
        clk_out0_gate   = 3'b000;
        clk_out1_gate   = 3'b000;
        clk_out2_gate   = 3'b000;
        clk_out3_gate   = 3'b000;
        clk_out4_gate   = 3'b000;
        clk_outphy_gate = 3'b000;
        clk_outf_gate   = 3'b000;
        #1;
        inner_rstn = 1'b1;
        clk_in_first_time = 1'b1;
        clk_fb_first_time = 1'b1;
    end
///////////////////////////////////////////////////////
////RESET//////////////////////////////////////////////
    assign rst_n = ~(PLL_PWD | RST) & inner_rstn;
///////////////////////////////////////////////////////
////INPUT_CLK_SEL//////////////////////////////////////
    assign clk_in = (CLKIN_SEL == 1'b0) ? CLKIN1 : CLKIN2;
///////////////////////////////////////////////////////
////FBCK_DELAY/////////////////////////////////////////
    always @(posedge clk_in or negedge rst_n)
    begin
        if(!rst_n)
        begin
            clk_in_first_time = 1'b1;
            clk_in_first_edge = 0.0;
        end
        else
        begin
            if(clk_in_first_time == 1'b1)
                clk_in_first_edge = $realtime;
            clk_in_first_time = 1'b0;
        end
    end

    always @(posedge CLKFB or negedge rst_n)
    begin
        if(!rst_n)
        begin
            clk_fb_first_time = 1'b1;
            clk_fb_first_edge = 0.0;
        end
        else
        begin
            if(clk_fb_first_time == 1'b1)
                clk_fb_first_edge = $realtime;
            clk_fb_first_time = 1'b0;
        end
    end
///////////////////////////////////////////////////////
////CLK_TEST///////////////////////////////////////////
    always #200 clk_test = ~clk_test;

    always @(posedge clk_test or negedge rst_n)
    begin
        if(!rst_n)
        begin
            clkref_wo <= 1'b0;
            clkref_test_time1 = 0;
            clkref_test_time2 = 0;
            clkref_test_time3 = 0;
        end
        else
        begin
            clkref_test_time3 = clkref_test_time2;
            clkref_test_time2 = clkref_test_time1;
            clkref_test_time1 = clkin_rtime_next;
            if(clkref_test_time3 == clkref_test_time1)
                clkref_wo <= 1'b1;
            else
                clkref_wo <= 1'b0;
        end
    end

    always @(posedge CLKFB or negedge rst_n)
    begin
        if(!rst_n)
        begin
            clkfb_rtime_last = 0.0;
            clkfb_rtime_next = 0.0;
        end
        else
        begin
            clkfb_rtime_last = clkin_rtime_next;
            clkfb_rtime_next = $realtime;
        end
    end

    always @(posedge clk_test or negedge rst_n)
    begin
        if(!rst_n)
        begin
            clkfb_wo <= 1'b0;
            clkfb_test_time3 = 0;
            clkfb_test_time2 = 0;
            clkfb_test_time1 = 0;
        end
        else
        begin
            if(clk_fb_first_time == 1'b0)
            begin
                clkfb_test_time3 = clkfb_test_time2;
                clkfb_test_time2 = clkfb_test_time1;
                clkfb_test_time1 = clkfb_rtime_next;
                if(clkfb_test_time3 == clkfb_test_time1)
                    clkfb_wo <= 1'b1;
                else
                    clkfb_wo <= 1'b0;
            end
        end
    end

    assign clkwo = clkref_wo | clkfb_wo;
///////////////////////////////////////////////////////
////PLL_ANALOG/////////////////////////////////////////
////FEEDBACK_DIVIDER_CAL///////////////////////////////
    assign idivider   = ratioi;
    assign mdivider   = ratiom;
    assign fdivider   = ratiof;
    assign divider0   = ratio0;
    assign divider1   = ratio1;
    assign divider2   = ratio2;
    assign divider3   = ratio3;
    assign divider4   = ratio4;
    assign dividerphy = ratiophy;

    always @(*)
    begin
    	if(INTERNAL_FB == "CLKOUTF" || EXTERNAL_FB == "CLKOUTF")
            fsdiv_set_int = fdivider;
        else if(INTERNAL_FB == "CLKOUT0" || EXTERNAL_FB == "CLKOUT0")
            fsdiv_set_int = divider0;
        else if(INTERNAL_FB == "CLKOUT1" || EXTERNAL_FB == "CLKOUT1")
            fsdiv_set_int = divider1;
        else if(INTERNAL_FB == "CLKOUT2" || EXTERNAL_FB == "CLKOUT2")
            fsdiv_set_int = divider2;
        else if(INTERNAL_FB == "CLKOUT3" || EXTERNAL_FB == "CLKOUT3")
            fsdiv_set_int = divider3;
        else if(INTERNAL_FB == "CLKOUT4" || EXTERNAL_FB == "CLKOUT4")
            fsdiv_set_int = divider4;
    end

    always @(*)
    begin
        fbdiv_set_int = mdivider * fsdiv_set_int;
    end
////PLL_VCO_CAL////////////////////////////////////////
    assign rstanalog_n = rst_n;

    always @(posedge clk_in or negedge rstanalog_n)
    begin
        if(!rstanalog_n)
        begin
            clkin_rtime_last = 0.0;
            clkin_rtime_next = 0.0;
            clkin_time  <= 0.0;
            clkin_time1 <= 0.0;
            clkin_time2 <= 0.0;
            clkin_time3 <= 0.0;
            clkout_lock <= 0.0;
            vcoclk_period <= 1'b0;
            vcoclk_period_half <= 0.0;
            clkout0_time       <= 0.0;
            clkout1_time       <= 0.0;
            clkout2_time       <= 0.0;
            clkout3_time       <= 0.0;
            clkout4_time       <= 0.0;
            vcoclk_period_amp  <= 0.0;
            vcoclk_period_real <= 0.0;
            vcoclk_period_dev  <= 0.0;
        end
        else
        begin
            clkin_rtime_last = clkin_rtime_next;
            clkin_rtime_next = $realtime;
            if(clkin_rtime_last > 0)
            begin
                clkin_time  <= clkin_rtime_next-clkin_rtime_last;
                clkin_time1 <= clkin_time;
                clkin_time2 <= clkin_time1;
                clkin_time3 <= clkin_time2;
            end
            if(clkin_time > 0)
            begin
                clkout_lock <= (clkin_time  > 0) &&
                               (clkin_time1 > 0) &&
                               (clkin_time2 > 0) &&
                               (clkin_time3 > 0) &&
                               ((clkin_time - clkin_time1)  < 0.0001) &&
                               ((clkin_time1 - clkin_time)  < 0.0001) &&
                               ((clkin_time1 - clkin_time2) < 0.0001) &&
                               ((clkin_time2 - clkin_time1) < 0.0001) &&
                               ((clkin_time2 - clkin_time3) < 0.0001) &&
                               ((clkin_time3 - clkin_time2) < 0.0001);
            end
            if(clkin_time > 0)
            begin
                vcoclk_period      = (clkin_time * idivider) / fbdiv_set_int;
                vcoclk_period_half = vcoclk_period / 2;
                clkout0_time       = vcoclk_period * divider0;
                clkout1_time       = vcoclk_period * divider1;
                clkout2_time       = vcoclk_period * divider2;
                clkout3_time       = vcoclk_period * divider3;
                clkout4_time       = vcoclk_period * divider4;
                clkoutphy_time     = vcoclk_period * dividerphy;
                clkoutf_time       = vcoclk_period * fdivider;
                vcoclk_period_amp  = vcoclk_period_half * 100000;
                vcoclk_period_real = vcoclk_period_amp / 100000.0;
                vcoclk_period_dev  = (clkin_time - (vcoclk_period_real * 2 * fbdiv_set_int) / idivider) / 2;
            end
        end
    end

    always @(*)
    begin
        if(!rst_n)
        begin
            done = 1'b0;
            idiv_set = 0;
            fdiv_set = 0;
            swap_set = 0;
            midd_set = 0;
            offset = 0;
        end
        else
        begin
            idiv_set = idivider;
            fdiv_set = $rtoi(fbdiv_set_int);
            while(!done)
            begin
                if(idiv_set < fdiv_set)
                begin
                    swap_set = idiv_set;
                    idiv_set = fdiv_set;
                    fdiv_set = swap_set;
                end
                else
                    if(fdiv_set != 0)
                        idiv_set = idiv_set - fdiv_set;
                    else
                    begin
                        done = 1;
                        midd_set = idiv_set;
                    end
            end
        end
    end

    always @(*)
    begin
        if(!rst_n)
        begin
            fdiv_int = 0;
            offset = 0;
        end
        else
            begin
                fdiv_int = midd_set;
                offset = vcoclk_period_dev * idivider/midd_set;
            end
    end

    always @(clkout_lock or inner_clk or clkwo)
    begin
        if(clkout_lock == 1'b0 || clkwo == 1'b1)
        begin
            inner_clk <= 1'b0;
            clk_gate  <= 1'b1;
            cnt_fdiv   = 0;
        end
        else
            if(clk_gate == 1)
            begin
                inner_clk <= 1'b1;
                clk_gate  <= 1'b0;
                cnt_fdiv   = 0;
            end
            else
            begin
                cnt_fdiv = cnt_fdiv + 1;
                if(cnt_fdiv  == fbdiv_set_int/fdiv_int)
                begin
                    inner_clk <= #(vcoclk_period_half + offset) ~inner_clk;
                    cnt_fdiv = 0;
                end
                else
                    inner_clk <= #vcoclk_period_half ~inner_clk;
            end
    end

    always @(clk_in or CLKFB or negedge rst_n)
    begin
        if(!rst_n)
        begin
            adjust <= 1'b1;
            fb_route_delay = 0.0;
            tmp_ratio  = 0;
            tmp_delay  = 0.0;
            real_delay = 0.0;
        end
        else
            if(adjust == 1'b1)
            begin
                fb_route_delay = clk_fb_first_edge - clk_in_first_edge;
                if((clkin_time > 0) && (fb_route_delay > 0))
                begin
                    tmp_ratio  = fb_route_delay / clkin_time;
                    tmp_delay  = fb_route_delay - (clkin_time * tmp_ratio);
                    real_delay = clkin_time - tmp_delay;
                    adjust <= 1'b0;
                end
            end
    end

    always @(inner_clk)
    begin
        if(EXTERNAL_FB == "CLKOUTF" || EXTERNAL_FB == "CLKOUT0" || EXTERNAL_FB == "CLKOUT1" || EXTERNAL_FB == "CLKOUT2" || EXTERNAL_FB == "CLKOUT3" || EXTERNAL_FB == "CLKOUT4")
            vcoclk <= #real_delay inner_clk;
        else
            vcoclk <= inner_clk;
    end
///////////////////////////////////////////////////////
////PLL_LOCK///////////////////////////////////////////
    assign clk_lock = (INTERNAL_FB == "DISABLE") ? CLKFB : clk_in;
    
    always @(posedge clk_lock or negedge rstanalog_n or clk_gate)
    begin
        if(!rstanalog_n)
        begin
            start_clk <= 1'b0;
            cnt_clkfb <= 2'b00;
        end
        else
            if(!clk_gate)
                if(cnt_clkfb == 2'b11)
                    start_clk = 1'b1;
                else
                    cnt_clkfb = cnt_clkfb + 1'b1;
            else
            begin
                start_clk <= 1'b0;
                cnt_clkfb <= 2'b00;
            end 
    end

    always @(posedge clk_in or negedge rstanalog_n or clk_gate)
    begin
        if(!rstanalog_n)
        begin
            cnt_lock  <= 8'h1;
            lock_wait <= 1'b0;
        end
        else
            if(!clk_gate && start_clk)
                if(cnt_lock == idivider * 3)
                    lock_wait <= 1'b1;
                else
                    cnt_lock <= cnt_lock + 1'b1;
            else
            begin
                cnt_lock <= 8'h1;
                lock_wait <= 1'b0;
            end
    end

    always @(posedge clk_in or negedge rst_n or clk_gate)
    begin
        if(!rst_n)
            lock_reg <= 1'b0;
        else
            if(LOCK_MODE == 1'b0)
                if(!clk_gate)
                    lock_reg <= lock_wait;
                else
                    lock_reg <= 1'b0;
            else
                lock_reg <= lock_reg | lock_wait;
    end

    assign LOCK = lock_reg;
///////////////////////////////////////////////////////
////PLL_ODIV///////////////////////////////////////////
////ODIV0//////////////////////////////////////////////
    assign odiv0_clkin = (muxsel0_en) ? vcoclk : 1'b0;

    always @(posedge odiv0_clkin or negedge odiv0_clkin or negedge rst_n)
    begin
        if(!rst_n)
        begin
            odiv0_counter <= 8'h0;
            odiv0_out_reg <= 1'b0;
        end
        else
        begin
            if(divider0 == 8'h1)
            begin
                odiv0_counter <= 8'h0;
                odiv0_out_reg <= 1'b0;
            end
            else
            begin
                if(odiv0_counter < ({divider0, 1'b0} - 1'b1))
                    odiv0_counter <= odiv0_counter + 1'b1;
                else
                    odiv0_counter <= 8'h0;

                if(odiv0_counter < duty0)
                    odiv0_out_reg <= 1'b1;
                else
                    odiv0_out_reg <= 1'b0;
            end
        end
    end

    assign odiv0_out = (divider0 == 8'h1) ? odiv0_clkin : odiv0_out_reg;
////ODIV1//////////////////////////////////////////////
    assign odiv1_clkin = (muxsel1_en) ? vcoclk : 1'b0;

    always @(posedge odiv1_clkin or negedge odiv1_clkin or negedge rst_n)
    begin
        if(!rst_n)
        begin
            odiv1_counter <= 8'h0;
            odiv1_out_reg <= 1'b0;
        end
        else
        begin
            if(divider1 == 8'h1)
            begin
                odiv1_counter <= 8'h0;
                odiv1_out_reg <= 1'b0;
            end
            else
            begin
                if(odiv1_counter < ({divider1, 1'b0} - 1'b1))
                    odiv1_counter <= odiv1_counter + 1'b1;
                else
                    odiv1_counter <= 8'h0;

                if(odiv1_counter < duty1)
                    odiv1_out_reg <= 1'b1;
                else
                    odiv1_out_reg <= 1'b0;
            end
        end
    end

    assign odiv1_out = (divider1 == 8'h1) ? odiv1_clkin : odiv1_out_reg;
////ODIV2//////////////////////////////////////////////
    assign odiv2_clkin = (muxsel2_en) ? vcoclk : 1'b0;

    always @(posedge odiv2_clkin or negedge odiv2_clkin or negedge rst_n)
    begin
        if(!rst_n)
        begin
            odiv2_counter <= 8'h0;
            odiv2_out_reg <= 1'b0;
        end
        else
        begin
            if(divider2 == 8'h1)
            begin
                odiv2_counter <= 8'h0;
                odiv2_out_reg <= 1'b0;
            end
            else
            begin
                if(odiv2_counter < ({divider2, 1'b0} - 1'b1))
                    odiv2_counter <= odiv2_counter + 1'b1;
                else
                    odiv2_counter <= 8'h0;

                if(odiv2_counter < duty2)
                    odiv2_out_reg <= 1'b1;
                else
                    odiv2_out_reg <= 1'b0;
            end
        end
    end

    assign odiv2_out = (divider2 == 8'h1) ? odiv2_clkin : odiv2_out_reg;
////ODIV3//////////////////////////////////////////////
    assign odiv3_clkin = (muxsel3_en) ? vcoclk : 1'b0;

    always @(posedge odiv3_clkin or negedge odiv3_clkin or negedge rst_n)
    begin
        if(!rst_n)
        begin
            odiv3_counter <= 8'h0;
            odiv3_out_reg <= 1'b0;
        end
        else
        begin
            if(divider3 == 8'h1)
            begin
                odiv3_counter <= 8'h0;
                odiv3_out_reg <= 1'b0;
            end
            else
            begin
                if(odiv3_counter < ({divider3, 1'b0} - 1'b1))
                    odiv3_counter <= odiv3_counter + 1'b1;
                else
                    odiv3_counter <= 8'h0;

                if(odiv3_counter < duty3)
                    odiv3_out_reg <= 1'b1;
                else
                    odiv3_out_reg <= 1'b0;
            end
        end
    end

    assign odiv3_out = (divider3 == 8'h1) ? odiv3_clkin : odiv3_out_reg;
////ODIV4//////////////////////////////////////////////
    assign odiv4_clkin = (muxsel4_en) ? vcoclk : 1'b0;

    always @(posedge odiv4_clkin or negedge odiv4_clkin or negedge rst_n)
    begin
        if(!rst_n)
        begin
            odiv4_counter <= 8'h0;
            odiv4_out_reg <= 1'b0;
        end
        else
        begin
            if(divider4 == 8'h1)
            begin
                odiv4_counter <= 8'h0;
                odiv4_out_reg <= 1'b0;
            end
            else
            begin
                if(odiv4_counter < ({divider4, 1'b0} - 1'b1))
                    odiv4_counter <= odiv4_counter + 1'b1;
                else
                    odiv4_counter <= 8'h0;

                if(odiv4_counter < duty4)
                    odiv4_out_reg <= 1'b1;
                else
                    odiv4_out_reg <= 1'b0;
            end
        end
    end

    assign odiv4_out = (divider4 == 8'h1) ? odiv4_clkin : odiv4_out_reg;
////ODIVPHY////////////////////////////////////////////
    assign odivphy_clkin = (muxselphy_en) ? vcoclk : 1'b0;

    always @(posedge odivphy_clkin or negedge odivphy_clkin or negedge rst_n)
    begin
        if(!rst_n)
        begin
            odivphy_counter <= 8'h0;
            odivphy_out_reg <= 1'b0;
        end
        else
        begin
            if(dividerphy == 8'h1)
            begin
                odivphy_counter <= 8'h0;
                odivphy_out_reg <= 1'b0;
            end
            else
            begin
                if(odivphy_counter < ({dividerphy, 1'b0} - 1'b1))
                    odivphy_counter <= odivphy_counter + 1'b1;
                else
                    odivphy_counter <= 8'h0;

                if(odivphy_counter < dutyphy)
                    odivphy_out_reg <= 1'b1;
                else
                    odivphy_out_reg <= 1'b0;
            end
        end
    end

    assign odivphy_out = (dividerphy == 8'h1) ? odivphy_clkin : odivphy_out_reg;
////FDIV///////////////////////////////////////////////
    assign fdiv_clkin = (muxself_en) ? vcoclk : 1'b0;

    always @(posedge fdiv_clkin or negedge fdiv_clkin or negedge rst_n)
    begin
        if(!rst_n)
        begin
            fdiv_counter <= 8'h0;
            fdiv_out_reg <= 1'b0;
        end
        else
        begin
            if(fdivider == 8'h1)
            begin
                fdiv_counter <= 8'h0;
                fdiv_out_reg <= 1'b0;
            end
            else
            begin
                if(fdiv_counter < ({fdivider, 1'b0} - 1'b1))
                    fdiv_counter <= fdiv_counter + 1'b1;
                else
                    fdiv_counter <= 8'h0;

                if(fdiv_counter < dutyf)
                    fdiv_out_reg <= 1'b1;
                else
                    fdiv_out_reg <= 1'b0;
            end
        end
    end

    assign fdiv_out = (fdivider == 8'h1) ? fdiv_clkin : fdiv_out_reg;
///////////////////////////////////////////////////////
////PHASE_SHIFT////////////////////////////////////////
    always @(*)
    begin
        if(clkout0_time > 0)
            vco_fphase_delay0 <= (odiv0_fphase * clkout0_time) / (8 * divider0);

        if(clkout1_time > 0)
            vco_fphase_delay1 <= (odiv1_fphase * clkout1_time) / (8 * divider1);

        if(clkout2_time > 0)
            vco_fphase_delay2 <= (odiv2_fphase * clkout2_time) / (8 * divider2);

        if(clkout3_time > 0)
            vco_fphase_delay3 <= (odiv3_fphase * clkout3_time) / (8 * divider3);

        if(clkout4_time > 0)
            vco_fphase_delay4 <= (odiv4_fphase * clkout4_time) / (8 * divider4);

        if(clkoutphy_time > 0)
            vco_fphase_delayphy <= (odivphy_fphase * clkoutphy_time) / (8 * dividerphy);

        if(clkoutf_time > 0)
            vco_fphase_delayf <= (fdiv_fphase * clkoutf_time) / (8 * fdivider);
    end

    always @(*)
    begin
        if(divider0 > odiv0_cphase)
            cphase0 = odiv0_cphase;
        else
            cphase0 = odiv0_cphase - (odiv0_cphase / divider0) * divider0;

        if(divider1 > odiv1_cphase)
            cphase1 = odiv1_cphase;
        else
            cphase1 = odiv1_cphase - (odiv1_cphase / divider1) * divider1;

        if(divider2 > odiv2_cphase)
            cphase2 = odiv2_cphase;
        else
            cphase2 = odiv2_cphase - (odiv2_cphase / divider2) * divider2;

        if(divider3 > odiv3_cphase)
            cphase3 = odiv3_cphase;
        else
            cphase3 = odiv3_cphase - (odiv3_cphase / divider3) * divider3;

        if(divider4 > odiv4_cphase)
            cphase4 = odiv4_cphase;
        else
            cphase4 = odiv4_cphase - (odiv4_cphase / divider4) * divider4;

        if(dividerphy > odivphy_cphase)
            cphasephy = odivphy_cphase;
        else
            cphasephy = odivphy_cphase - (odivphy_cphase / dividerphy) * dividerphy;

        if(fdivider > fdiv_cphase)
            cphasef = fdiv_cphase;
        else
            cphasef = fdiv_cphase - (fdiv_cphase / fdivider) * fdivider;
    end

    always @(*)
    begin
        if(clkout0_time > 0)
            cphase_delay0 <= clkout0_time - (((divider0 - cphase0) * clkout0_time) / divider0);
        else
            cphase_delay0 <= 0.0;

        if(clkout1_time > 0)
            cphase_delay1 <= clkout1_time - (((divider1 - cphase1) * clkout1_time) / divider1);
        else
            cphase_delay1 <= 0.0;

        if(clkout2_time > 0)
            cphase_delay2 <= clkout2_time - (((divider2 - cphase2) * clkout2_time) / divider2);
        else
            cphase_delay2 <= 0.0;

        if(clkout3_time > 0)
            cphase_delay3 <= clkout3_time - (((divider3 - cphase3) * clkout3_time) / divider3);
        else
            cphase_delay3 <= 0.0;

        if(clkout4_time > 0)
            cphase_delay4 <= clkout4_time - (((divider4 - cphase4) * clkout4_time) / divider4);
        else
            cphase_delay4 <= 0.0;

        if(clkoutphy_time > 0)
            cphase_delayphy <= clkoutphy_time - (((dividerphy - cphasephy) * clkoutphy_time) / dividerphy);
        else
            cphase_delayphy <= 0.0;

        if(clkoutf_time > 0)
            cphase_delayf <= clkoutf_time - (((fdivider - cphasef) * clkoutf_time) / fdivider);
        else
            cphase_delayf <= 0.0;
    end
////PHASE_SHIFT_DLY////////////////////////////////////
    always @(odiv0_out or negedge rst_n)
    begin
        if(!rst_n)
            odiv0_out_delay1 <= 1'b0;
        else
            odiv0_out_delay1 <= #vco_fphase_delay0 odiv0_out;
    end

    always @(odiv0_out_delay1 or negedge rst_n)
    begin
        if(!rst_n)
            odiv0_out_delay <= 1'b0;
        else
            odiv0_out_delay <= #cphase_delay0 odiv0_out_delay1;
    end

    always @(odiv1_out or negedge rst_n)
    begin
        if(!rst_n)
            odiv1_out_delay1 <= 1'b0;
        else
            odiv1_out_delay1 <= #vco_fphase_delay1 odiv1_out;
    end

    always @(odiv1_out_delay1 or negedge rst_n)
    begin
        if(!rst_n)
            odiv1_out_delay <= 1'b0;
        else
            odiv1_out_delay <= #cphase_delay1 odiv1_out_delay1;
    end

    always @(odiv2_out or negedge rst_n)
    begin
        if(!rst_n)
            odiv2_out_delay1 <= 1'b0;
        else
            odiv2_out_delay1 <= #vco_fphase_delay2 odiv2_out;
    end

    always @(odiv2_out_delay1 or negedge rst_n)
    begin
        if(!rst_n)
            odiv2_out_delay <= 1'b0;
        else
            odiv2_out_delay <= #cphase_delay2 odiv2_out_delay1;
    end

    always @(odiv3_out or negedge rst_n)
    begin
        if(!rst_n)
            odiv3_out_delay1 <= 1'b0;
        else
            odiv3_out_delay1 <= #vco_fphase_delay3 odiv3_out;
    end

    always @(odiv3_out_delay1 or negedge rst_n)
    begin
        if(!rst_n)
            odiv3_out_delay <= 1'b0;
        else
            odiv3_out_delay <= #cphase_delay3 odiv3_out_delay1;
    end

    always @(odiv4_out or negedge rst_n)
    begin
        if(!rst_n)
            odiv4_out_delay1 <= 1'b0;
        else
            odiv4_out_delay1 <= #vco_fphase_delay4 odiv4_out;
    end

    always @(odiv4_out_delay1 or negedge rst_n)
    begin
        if(!rst_n)
            odiv4_out_delay <= 1'b0;
        else
            odiv4_out_delay <= #cphase_delay4 odiv4_out_delay1;
    end

    always @(odivphy_out or negedge rst_n)
    begin
        if(!rst_n)
            odivphy_out_delay1 <= 1'b0;
        else
            odivphy_out_delay1 <= #vco_fphase_delayphy odivphy_out;
    end

    always @(odivphy_out_delay1 or negedge rst_n)
    begin
        if(!rst_n)
            odivphy_out_delay <= 1'b0;
        else
            odivphy_out_delay <= #cphase_delayphy odivphy_out_delay1;
    end

    always @(fdiv_out or negedge rst_n)
    begin
        if(!rst_n)
            fdiv_out_delay1 <= 1'b0;
        else
            fdiv_out_delay1 <= #vco_fphase_delayf fdiv_out;
    end

    always @(fdiv_out_delay1 or negedge rst_n)
    begin
        if(!rst_n)
            fdiv_out_delay <= 1'b0;
        else
            fdiv_out_delay <= #cphase_delayf fdiv_out_delay1;
    end
///////////////////////////////////////////////////////
////PLL_GATE///////////////////////////////////////////
    assign clkout0_gate = (CLKOUT0_SYN_EN == "TRUE") ? CLKOUT0_SYN : 1'b0;

    always @(negedge odiv0_out_delay or negedge rst_n)
    begin
        if(!rst_n)
            clk_out0_gate <= 3'b000;
        else
            clk_out0_gate <= {clk_out0_gate[1:0], ~clkout0_gate};
    end

    assign CLKOUT0  = odiv0_out_delay & clk_out0_gate[2];
    assign CLKOUT0N = ~CLKOUT0;

    assign clkout1_gate = (CLKOUT1_SYN_EN == "TRUE") ? CLKOUT1_SYN : 1'b0;

    always @(negedge odiv1_out_delay or negedge rst_n)
    begin
        if(!rst_n)
            clk_out1_gate <= 3'b000;
        else
            clk_out1_gate <= {clk_out1_gate[1:0], ~clkout1_gate};
    end

    assign CLKOUT1  = odiv1_out_delay & clk_out1_gate[2];
    assign CLKOUT1N = ~CLKOUT1;    

    assign clkout2_gate = (CLKOUT2_SYN_EN == "TRUE") ? CLKOUT2_SYN : 1'b0;

    always @(negedge odiv2_out_delay or negedge rst_n)
    begin
        if(!rst_n)
            clk_out2_gate <= 3'b000;
        else
            clk_out2_gate <= {clk_out2_gate[1:0], ~clkout2_gate};
    end

    assign CLKOUT2  = odiv2_out_delay & clk_out2_gate[2];
    assign CLKOUT2N = ~CLKOUT2;

    assign clkout3_gate = (CLKOUT3_SYN_EN == "TRUE") ? CLKOUT3_SYN : 1'b0;

    always @(negedge odiv3_out_delay or negedge rst_n)
    begin
        if(!rst_n)
            clk_out3_gate <= 3'b000;
        else
            clk_out3_gate <= {clk_out3_gate[1:0], ~clkout3_gate};
    end

    assign CLKOUT3  = odiv3_out_delay & clk_out3_gate[2];
    assign CLKOUT3N = ~CLKOUT3;

    assign clkout4_gate = (CLKOUT4_SYN_EN == "TRUE") ? CLKOUT4_SYN : 1'b0;

    always @(negedge odiv4_out_delay or negedge rst_n)
    begin
        if(!rst_n)
            clk_out4_gate <= 3'b000;
        else
            clk_out4_gate <= {clk_out4_gate[1:0], ~clkout4_gate};
    end

    assign CLKOUT4  = odiv4_out_delay & clk_out4_gate[2];

    assign clkoutphy_gate = (CLKOUTPHY_SYN_EN == "TRUE") ? CLKOUTPHY_SYN : 1'b0;

    always @(negedge odivphy_out_delay or negedge rst_n)
    begin
        if(!rst_n)
            clk_outphy_gate <= 3'b000;
        else
            clk_outphy_gate <= {clk_outphy_gate[1:0], ~clkoutphy_gate};
    end

    assign CLKOUTPHY  = odivphy_out_delay & clk_outphy_gate[2];
    assign CLKOUTPHYN = ~CLKOUTPHY;

    assign clkoutf_gate = (CLKOUTF_SYN_EN == "TRUE") ? CLKOUTF_SYN: 1'b0;

    always @(negedge fdiv_out_delay or negedge rst_n)
    begin
        if(!rst_n)
            clk_outf_gate <= 3'b000;
        else
            clk_outf_gate <= {clk_outf_gate[1:0], ~clkoutf_gate};
    end

    assign CLKOUTF  = fdiv_out_delay & clk_outf_gate[2];
    assign CLKOUTFN = ~CLKOUTF;
///////////////////////////////////////////////////////
////APB////////////////////////////////////////////////
    always @(posedge APB_CLK or negedge APB_RST_N)
    begin
       if(!APB_RST_N)
           apb_rstn_sync <= 2'b00;
       else
           apb_rstn_sync <= {apb_rstn_sync[0], 1'b1};
    end

    always @(posedge APB_CLK or negedge apb_rstn_sync[1])
    begin
        if(!apb_rstn_sync[1])
            ready <= 1'b0;
        else
            if(APB_SEL && !APB_EN)
                ready <= 1'b1;
            else
                ready <= 1'b0;
    end

    always @(posedge APB_CLK)
    begin
        if(APB_WRITE && APB_SEL && APB_EN)
            case(APB_ADDR)
                5'h0 : mem0  <= APB_WDATA;
                5'h1 : mem1  <= APB_WDATA[10:0];
                5'h2 : mem2  <= APB_WDATA;
                5'h3 : mem3  <= APB_WDATA[10:0];
                5'h4 : mem4  <= APB_WDATA;
                5'h5 : mem5  <= APB_WDATA[10:0];
                5'h6 : mem6  <= APB_WDATA;
                5'h7 : mem7  <= APB_WDATA[10:0];
                5'h8 : mem8  <= APB_WDATA;
                5'h9 : mem9  <= APB_WDATA[10:0];
                5'hA : mem10 <= APB_WDATA;
                5'hB : mem11 <= APB_WDATA[10:0];
                5'hC : mem12 <= APB_WDATA;
                5'hD : mem13 <= APB_WDATA[10:0];
                5'hE : mem14 <= APB_WDATA[7:0];
                5'hF : mem15 <= APB_WDATA[7:0];
                5'h10: mem16 <= APB_WDATA[13:0];
                5'h11: mem17 <= APB_WDATA[5:0];
            endcase
    end

    always @(posedge APB_CLK or negedge apb_rstn_sync[1])
    begin
        if(!apb_rstn_sync[1])
            rdata <= 16'h0;
        else
            if(!APB_WRITE && APB_SEL && !APB_EN)
                case(APB_ADDR)
                    5'h0 : rdata <= mem0;
                    5'h1 : rdata <= mem1;
                    5'h2 : rdata <= mem2;
                    5'h3 : rdata <= mem3;
                    5'h4 : rdata <= mem4;
                    5'h5 : rdata <= mem5;
                    5'h6 : rdata <= mem6;
                    5'h7 : rdata <= mem7;
                    5'h8 : rdata <= mem8;
                    5'h9 : rdata <= mem9;
                    5'hA : rdata <= mem10;
                    5'hB : rdata <= mem11;
                    5'hC : rdata <= mem12;
                    5'hD : rdata <= mem13;
                    5'hE : rdata <= mem14;
                    5'hF : rdata <= mem15;
                    5'h10: rdata <= mem16;
                    5'h11: rdata <= mem17;
                endcase
            else
                rdata <= 16'h0;
    end

    assign APB_READY = ready;
    assign APB_RDATA = rdata;
endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_ROM32X1.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_ROM32X1
#(
    parameter [31:0] INIT = 32'h0000_0000
) (
    output Z,
    input I0, I1, I2, I3, I4
);

   reg [31:0] mem;
   wire [4:0] addr;

   initial mem = INIT;

   assign addr = {I4, I3, I2, I1, I0};
   //assign Z = mem[addr];
   assign Z = INIT[addr];

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_RAM32X2DP.v
//
// Functional description: simple-dual-port 32x2 distributed ram
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_RAM32X2DP
#(
    parameter [31:0] INIT_0 = 32'h00000000 ,
    parameter [31:0] INIT_1 = 32'h00000000
) (
    output [1:0] DO,
    input  [1:0] DI,
    input [4:0] RADDR, WADDR,
    input WCLK, WE
);

    reg [31:0] mem [1:0];

    initial begin
        mem[0] = INIT_0;
        mem[1] = INIT_1;
    end

    always @(posedge WCLK) begin
        if (WE == 1'b1) begin
            mem[0][WADDR] <= DI[0];
            mem[1][WADDR] <= DI[1];
        end
    end

    assign DO[0] = mem[0][RADDR];
    assign DO[1] = mem[1][RADDR];

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2019 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_GPLL.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1ns/1fs
module GTP_GPLL #(
    parameter real CLKIN_FREQ = 50.0,    //10MHz~800MHz
    parameter LOCK_MODE       = 1'b0,    //1'b0~1'b1
    parameter integer STATIC_RATIOI = 1,   //1~128
    parameter integer STATIC_RATIOM = 1,   //1~128
    parameter real    STATIC_RATIO0 = 1.0, //1~128 or 2.000~128.000
    parameter integer STATIC_RATIO1 = 1,   //1~128
    parameter integer STATIC_RATIO2 = 1,   //1~128
    parameter integer STATIC_RATIO3 = 1,   //1~128
    parameter integer STATIC_RATIO4 = 1,   //1~128
    parameter integer STATIC_RATIO5 = 1,   //1~128
    parameter integer STATIC_RATIO6 = 1,   //1~128
    parameter real    STATIC_RATIOF = 1.0, //1~128 or 2.000~128.000
    parameter integer STATIC_DUTY0 = 2, //2<=STATIC_DUTY0<=2*STATIC_RATIO0-1
    parameter integer STATIC_DUTY1 = 2, //2<=STATIC_DUTY1<=2*STATIC_RATIO1-1
    parameter integer STATIC_DUTY2 = 2, //2<=STATIC_DUTY2<=2*STATIC_RATIO2-1
    parameter integer STATIC_DUTY3 = 2, //2<=STATIC_DUTY3<=2*STATIC_RATIO3-1
    parameter integer STATIC_DUTY4 = 2, //2<=STATIC_DUTY4<=2*STATIC_RATIO4-1
    parameter integer STATIC_DUTY5 = 2, //2<=STATIC_DUTY5<=2*STATIC_RATIO5-1
    parameter integer STATIC_DUTY6 = 2, //2<=STATIC_DUTY6<=2*STATIC_RATIO6-1
    parameter integer STATIC_DUTYF = 2, //2<=STATIC_DUTYF<=2*STATIC_RATIOF-1
    parameter integer STATIC_PHASE   = 0, //0~63
    parameter integer STATIC_PHASE0  = 0, //0~7
    parameter integer STATIC_PHASE1  = 0, //0~7
    parameter integer STATIC_PHASE2  = 0, //0~7
    parameter integer STATIC_PHASE3  = 0, //0~7
    parameter integer STATIC_PHASE4  = 0, //0~7
    parameter integer STATIC_PHASE5  = 0, //0~7
    parameter integer STATIC_PHASE6  = 0, //0~7
    parameter integer STATIC_PHASEF  = 0, //0~7
    parameter integer STATIC_CPHASE0 = 0, //0~127
    parameter integer STATIC_CPHASE1 = 0, //0~127
    parameter integer STATIC_CPHASE2 = 0, //0~127
    parameter integer STATIC_CPHASE3 = 0, //0~127
    parameter integer STATIC_CPHASE4 = 0, //0~127
    parameter integer STATIC_CPHASE5 = 0, //0~127
    parameter integer STATIC_CPHASE6 = 0, //0~127
    parameter integer STATIC_CPHASEF = 0, //0~127
    parameter CLK_DPS0_EN = "FALSE", //"TRUE"; "FALSE"
    parameter CLK_DPS1_EN = "FALSE", //"TRUE"; "FALSE"
    parameter CLK_DPS2_EN = "FALSE", //"TRUE"; "FALSE"
    parameter CLK_DPS3_EN = "FALSE", //"TRUE"; "FALSE"
    parameter CLK_DPS4_EN = "FALSE", //"TRUE"; "FALSE"
    parameter CLK_DPS5_EN = "FALSE", //"TRUE"; "FALSE"
    parameter CLK_DPS6_EN = "FALSE", //"TRUE"; "FALSE"
    parameter CLK_DPSF_EN = "FALSE", //"TRUE"; "FALSE"
    parameter CLK_CAS5_EN  = "FALSE", //"TRUE"; "FALSE"
    parameter CLKOUT0_SYN_EN = "FALSE", //"TRUE"; "FALSE"
    parameter CLKOUT1_SYN_EN = "FALSE", //"TRUE"; "FALSE"
    parameter CLKOUT2_SYN_EN = "FALSE", //"TRUE"; "FALSE"
    parameter CLKOUT3_SYN_EN = "FALSE", //"TRUE"; "FALSE"
    parameter CLKOUT4_SYN_EN = "FALSE", //"TRUE"; "FALSE"
    parameter CLKOUT5_SYN_EN = "FALSE", //"TRUE"; "FALSE"
    parameter CLKOUT6_SYN_EN = "FALSE", //"TRUE"; "FALSE"
    parameter CLKOUTF_SYN_EN = "FALSE", //"TRUE"; "FALSE"
    parameter SSC_MODE      = "DISABLE",//"DOWN_LOW"; "DOWN_HIGH"; "CENTER_LOW"; "CENTER_HIGH"; "DISABLE";
    parameter real SSC_FREQ = 50.0,     //25KHz~250KHz;
    parameter INTERNAL_FB = "CLKOUTF",  //"CLKOUT0"; "CLKOUT1"; "CLKOUT2"; "CLKOUT3"; "CLKOUT4"; "CLKOUT5"; "CLKOUT6"; "CLKOUTF"; "DISABLE";
    parameter EXTERNAL_FB = "DISABLE",  //"CLKOUT0"; "CLKOUT1"; "CLKOUT2"; "CLKOUT3"; "CLKOUT4"; "CLKOUT5"; "CLKOUT6"; "CLKOUTF"; "DISABLE";
    parameter BANDWIDTH   = "OPTIMIZED" //"LOW"; "OPTIMIZED"; "HIGH"
    )(
    output CLKOUT0,
    output CLKOUT0N,
    output CLKOUT1,
    output CLKOUT1N,
    output CLKOUT2,
    output CLKOUT2N,
    output CLKOUT3,
    output CLKOUT3N,
    output CLKOUT4,
    output CLKOUT5,
    output CLKOUT6,
    output CLKOUTF,
    output CLKOUTFN,
    output LOCK,
    output DPS_DONE,
    output [15:0] APB_RDATA,
    output APB_READY,
    input CLKIN1,
    input CLKIN2,
    input CLKFB,
    input CLKIN_SEL,
    input DPS_CLK,
    input DPS_EN,
    input DPS_DIR,
    input CLKOUT0_SYN,
    input CLKOUT1_SYN,
    input CLKOUT2_SYN,
    input CLKOUT3_SYN,
    input CLKOUT4_SYN,
    input CLKOUT5_SYN,
    input CLKOUT6_SYN,
    input CLKOUTF_SYN,
    input PLL_PWD,
    input RST,
    input APB_CLK,
    input APB_RST_N,
    input [4:0] APB_ADDR,
    input APB_SEL,
    input APB_EN,
    input APB_WRITE,
    input [15:0] APB_WDATA
    );

    initial
    begin
        if((CLK_DPS0_EN == "TRUE") || (CLK_DPS0_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_GPLL error: illegal setting for CLKOUT0_DPS_EN");

        if((CLK_DPS1_EN == "TRUE") || (CLK_DPS1_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_GPLL error: illegal setting for CLKOUT1_DPS_EN");

        if((CLK_DPS2_EN == "TRUE") || (CLK_DPS2_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_GPLL error: illegal setting for CLKOUT2_DPS_EN");

        if((CLK_DPS3_EN == "TRUE") || (CLK_DPS3_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_GPLL error: illegal setting for CLKOUT3_DPS_EN");

        if((CLK_DPS4_EN == "TRUE") || (CLK_DPS4_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_GPLL error: illegal setting for CLKOUT4_DPS_EN");

        if((CLK_DPS5_EN == "TRUE") || (CLK_DPS5_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_GPLL error: illegal setting for CLKOUT5_DPS_EN");

        if((CLK_DPS6_EN == "TRUE") || (CLK_DPS6_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_GPLL error: illegal setting for CLKOUT6_DPS_EN");

        if((CLK_DPSF_EN == "TRUE") || (CLK_DPSF_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_GPLL error: illegal setting for CLK_DPSF_EN");

        if((CLK_CAS5_EN  == "TRUE") || (CLK_CAS5_EN  == "FALSE"))
        begin
        end
        else
            $display ("GTP_GPLL error: illegal setting for CLK_CAS5_EN ");

        if((CLKOUT0_SYN_EN == "TRUE") || (CLKOUT0_SYN_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_GPLL error: illegal setting for CLKOUT0_SYN_EN");

        if((CLKOUT1_SYN_EN == "TRUE") || (CLKOUT1_SYN_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_GPLL error: illegal setting for CLKOUT1_SYN_EN");

        if((CLKOUT2_SYN_EN == "TRUE") || (CLKOUT2_SYN_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_GPLL error: illegal setting for CLKOUT2_SYN_EN");

        if((CLKOUT3_SYN_EN == "TRUE") || (CLKOUT3_SYN_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_GPLL error: illegal setting for CLKOUT3_SYN_EN");

        if((CLKOUT4_SYN_EN == "TRUE") || (CLKOUT4_SYN_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_GPLL error: illegal setting for CLKOUT4_SYN_EN");

        if((CLKOUT5_SYN_EN == "TRUE") || (CLKOUT5_SYN_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_GPLL error: illegal setting for CLKOUT5_SYN_EN");

        if((CLKOUT6_SYN_EN == "TRUE") || (CLKOUT6_SYN_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_GPLL error: illegal setting for CLKOUT6_SYN_EN");

        if((CLKOUTF_SYN_EN == "TRUE") || (CLKOUTF_SYN_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_GPLL error: illegal setting for CLKOUTF_SYN_EN");

        if((INTERNAL_FB == "CLKOUT0") || (INTERNAL_FB == "CLKOUT1") || (INTERNAL_FB == "CLKOUT2") || (INTERNAL_FB == "CLKOUT3") || (INTERNAL_FB == "CLKOUT4") || (INTERNAL_FB == "CLKOUT5") || (INTERNAL_FB == "CLKOUT6") || (INTERNAL_FB == "CLKOUTF") || (INTERNAL_FB == "DISABLE"))
        begin
        end
        else
            $display ("GTP_GPLL error: illegal setting for INTERNAL_FB");

        if((EXTERNAL_FB == "CLKOUT0") || (EXTERNAL_FB == "CLKOUT1") || (EXTERNAL_FB == "CLKOUT2") || (EXTERNAL_FB == "CLKOUT3") || (EXTERNAL_FB == "CLKOUT4") || (EXTERNAL_FB == "CLKOUT5") || (INTERNAL_FB == "CLKOUT6") || (EXTERNAL_FB == "CLKOUTF") || (EXTERNAL_FB == "DISABLE"))
        begin
        end
        else
            $display ("GTP_GPLL error: illegal setting for EXTERNAL_FB");

        if((BANDWIDTH == "LOW") || (BANDWIDTH == "OPTIMIZED") || (BANDWIDTH == "HIGH"))
        begin
        end
        else
            $display ("GTP_GPLL error: illegal setting for BANDWIDTH");
    end
///////////////////////////////////////////////////////
////INITIAL////////////////////////////////////////////
    reg [7:0] ratioi_i, ratiom_i, ratiof_i, ratio0_i, ratio1_i, ratio2_i, ratio3_i, ratio4_i, ratio5_i, ratio6_i;
    reg [7:0] dutyf_i, duty0_i, duty1_i, duty2_i, duty3_i, duty4_i, duty5_i, duty6_i;
    reg [6:0] odiv0_cphase_i, odiv1_cphase_i, odiv2_cphase_i, odiv3_cphase_i, odiv4_cphase_i, odiv5_cphase_i, odiv6_cphase_i, fdiv_cphase_i;
    reg [2:0] odiv0_fphase_i, odiv1_fphase_i, odiv2_fphase_i, odiv3_fphase_i, odiv4_fphase_i, odiv5_fphase_i, odiv6_fphase_i, fdiv_fphase_i;

    reg [2:0] ratio0_frac_i, ratiof_frac_i;
    reg [2:0] psoffset0_i, psoffsetf_i;

    reg muxsel0_en_i, muxsel1_en_i, muxsel2_en_i, muxsel3_en_i, muxsel4_en_i, muxsel5_en_i, muxsel6_en_i, muxself_en_i;
    reg [1:0] muxsel0_i, muxsel1_i, muxsel2_i, muxsel3_i, muxsel4_i, muxsel5_i, muxsel6_i, muxself_i;

    reg odiv0_frac_en_i, fdiv_frac_en_i;
    reg [1:0] odiv0_frac_adjust_i, fdiv_frac_adjust_i;

    reg [15:0] mem0, mem1, mem2, mem3, mem4, mem5, mem6, mem7, mem8, mem9, mem10, mem11, mem12, mem13, mem14, mem15, mem16, mem17, mem18, mem19, mem20, mem21;
    reg [1:0] vctrl_i;
    reg [1:0] cp_selbias_i, cp_base_i;
    reg [3:0] cp_cur_i;
    reg [2:0] lpf_r_i;
    reg lpf_c_i;
    reg [5:0] lock_set_i;
    reg lockfilter_pd_i;

    integer dps_init;
    reg odiv0_dps_en, odiv1_dps_en, odiv2_dps_en, odiv3_dps_en, odiv4_dps_en, odiv5_dps_en, odiv6_dps_en, fdiv_dps_en;
    reg div_dps_en;

    integer ratio0_int, ratiof_int;
    real ratio0_fra, ratiof_fra;

    wire [7:0] ratioi, ratiom, ratiof, ratio0, ratio1, ratio2, ratio3, ratio4, ratio5, ratio6;
    wire [7:0] dutyf, duty0, duty1, duty2, duty3, duty4, duty5, duty6;
    wire [6:0] odiv0_cphase, odiv1_cphase, odiv2_cphase, odiv3_cphase, odiv4_cphase, odiv5_cphase, odiv6_cphase, fdiv_cphase;
    wire [2:0] odiv0_fphase, odiv1_fphase, odiv2_fphase, odiv3_fphase, odiv4_fphase, odiv5_fphase, odiv6_fphase, fdiv_fphase;
    
    wire [2:0] ratio0_frac, ratiof_frac;
    wire [2:0] psoffset0, psoffsetf;

    wire muxsel0_en, muxsel1_en, muxsel2_en, muxsel3_en, muxsel4_en, muxsel5_en, muxsel6_en, muxself_en;
    wire [1:0] muxsel0, muxsel1, muxsel2, muxsel3, muxsel4, muxsel5, muxsel6, muxself;

    wire odiv0_frac_en, fdiv_frac_en;
    wire [1:0] odiv0_frac_adjust, fdiv_frac_adjust;

    initial
    begin
        ratioi_i = STATIC_RATIOI;
        ratiom_i = STATIC_RATIOM;
        ratiof_i = $rtoi(STATIC_RATIOF);
        ratio0_i = $rtoi(STATIC_RATIO0);
        ratio1_i = STATIC_RATIO1;
        ratio2_i = STATIC_RATIO2;
        ratio3_i = STATIC_RATIO3;
        ratio4_i = STATIC_RATIO4;
        ratio5_i = STATIC_RATIO5;
        ratio6_i = STATIC_RATIO6;
        dutyf_i = STATIC_DUTYF;
        duty0_i = STATIC_DUTY0;
        duty1_i = STATIC_DUTY1;
        duty2_i = STATIC_DUTY2;
        duty3_i = STATIC_DUTY3;
        duty4_i = STATIC_DUTY4;
        duty5_i = STATIC_DUTY5;
        duty6_i = STATIC_DUTY6;
        odiv0_cphase_i = STATIC_CPHASE0;
        odiv1_cphase_i = STATIC_CPHASE1;
        odiv2_cphase_i = STATIC_CPHASE2;
        odiv3_cphase_i = STATIC_CPHASE3;
        odiv4_cphase_i = STATIC_CPHASE4;
        odiv5_cphase_i = STATIC_CPHASE5;
        odiv6_cphase_i = STATIC_CPHASE6;
        fdiv_cphase_i  = STATIC_CPHASEF;
        odiv0_fphase_i = STATIC_PHASE0;
        odiv1_fphase_i = STATIC_PHASE1;
        odiv2_fphase_i = STATIC_PHASE2;
        odiv3_fphase_i = STATIC_PHASE3;
        odiv4_fphase_i = STATIC_PHASE4;
        odiv5_fphase_i = STATIC_PHASE5;
        odiv6_fphase_i = STATIC_PHASE6;
        fdiv_fphase_i  = STATIC_PHASEF;
        muxsel0_en_i = 1'b1;
        muxsel1_en_i = 1'b1;
        muxsel2_en_i = 1'b1;
        muxsel3_en_i = 1'b1;
        muxsel4_en_i = 1'b1;
        muxsel5_en_i = 1'b1;
        muxsel6_en_i = 1'b1;
        muxself_en_i = 1'b1;
        vctrl_i        = 2'b00;
        cp_selbias_i   = 2'b01;
        cp_base_i      = 2'b10;
        cp_cur_i       = 4'b0001;
        lpf_r_i        = 3'b001;
        lpf_c_i        = 1'b0;
        lock_set_i      = 5'h0;
        lockfilter_pd_i = 1'b1;

        dps_init = STATIC_PHASE;

        if(CLK_DPS0_EN == "TRUE")
        begin
            muxsel0_i    = 2'b01;
            odiv0_dps_en = 1'b1;
        end
        else
        begin
            muxsel0_i    = 2'b00;
            odiv0_dps_en = 1'b0;
        end

        if(CLK_DPS1_EN == "TRUE")
        begin
            muxsel1_i    = 2'b01;
            odiv1_dps_en = 1'b1;
        end
        else
        begin
            muxsel1_i    = 2'b00;
            odiv1_dps_en = 1'b0;
        end

        if(CLK_DPS2_EN == "TRUE")
        begin
            muxsel2_i    = 2'b01;
            odiv2_dps_en = 1'b1;
        end
        else
        begin
            muxsel2_i    = 2'b00;
            odiv2_dps_en = 1'b0;
        end

        if(CLK_DPS3_EN == "TRUE")
        begin
            muxsel3_i    = 2'b01;
            odiv3_dps_en = 1'b1;
        end
        else
        begin
            muxsel3_i    = 2'b00;
            odiv3_dps_en = 1'b0;
        end

        if(CLK_DPS4_EN == "TRUE")
        begin
            muxsel4_i    = 2'b01;
            odiv4_dps_en = 1'b1;
        end
        else
        begin
            muxsel4_i    = 2'b00;
            odiv4_dps_en = 1'b0;
        end

        if(CLK_DPS5_EN == "TRUE")
        begin
            muxsel5_i    = 2'b01;
            odiv5_dps_en = 1'b1;
        end
        else if(CLK_CAS5_EN == "TRUE")
        begin
            muxsel5_i    = 2'b10;
            odiv5_dps_en = 1'b0;
        end
        else
        begin
            muxsel5_i    = 2'b00;
            odiv5_dps_en = 1'b0;
        end

        if(CLK_DPS6_EN == "TRUE")
        begin
            muxsel6_i    = 2'b01;
            odiv6_dps_en = 1'b1;
        end
        else
        begin
            muxsel6_i    = 2'b00;
            odiv6_dps_en = 1'b0;
        end

        if(CLK_DPSF_EN == "TRUE")
        begin
            muxself_i   = 2'b01;
            fdiv_dps_en = 1'b1;
        end
        else
        begin
            muxself_i   = 2'b00;
            fdiv_dps_en = 1'b0;
        end

        div_dps_en = odiv0_dps_en || odiv1_dps_en || odiv2_dps_en || odiv3_dps_en || odiv4_dps_en || odiv5_dps_en || odiv6_dps_en || fdiv_dps_en;

        ratio0_int    = $rtoi(STATIC_RATIO0);
        ratio0_fra    = STATIC_RATIO0 - ratio0_int;
        ratio0_frac_i = ratio0_fra * 8;
        
        if(ratio0_fra > 0.000)
        begin
            odiv0_frac_en_i = 1'b1;
            if(!ratio0_i[0])
            begin
                psoffset0_i = (ratio0_frac_i + 1'b1) / 2 + odiv0_fphase_i;
                if(ratio0_fra > 0.000 && ratio0_fra < 0.875)
                    odiv0_frac_adjust_i = 2'b11;
                else
                    odiv0_frac_adjust_i = 2'b10;
            end
            else
            begin
                psoffset0_i = ({1'b0, ratio0_frac_i} + 4'd9) / 2 + odiv0_fphase_i;
                if(ratio0_fra > 0.000 && ratio0_fra < 0.875)
                    odiv0_frac_adjust_i = 2'b00;
                else
                    odiv0_frac_adjust_i = 2'b01;
            end
        end
        else
        begin
            odiv0_frac_en_i     = 1'b0;
            psoffset0_i         = 3'b000;
            odiv0_frac_adjust_i = 2'b00;
        end

        ratiof_int    = $rtoi(STATIC_RATIOF);
        ratiof_fra    = STATIC_RATIOF - ratiof_int;
        ratiof_frac_i = ratiof_fra * 8;
        
        if(ratiof_fra > 0.000)
        begin
            fdiv_frac_en_i = 1'b1;
            if(!ratiof_i[0])
            begin
                psoffsetf_i = (ratiof_frac_i + 1'b1) / 2 + fdiv_fphase_i;
                if(ratiof_fra > 0.000 && ratiof_fra < 0.875)
                    fdiv_frac_adjust_i = 2'b11;
                else
                    fdiv_frac_adjust_i = 2'b10;
            end
            else
            begin
                psoffsetf_i = ({1'b0, ratiof_frac_i} + 4'd9) / 2 + fdiv_fphase_i;
                if(ratiof_fra > 0.000 && ratiof_fra < 0.875)
                    fdiv_frac_adjust_i = 2'b00;
                else
                    fdiv_frac_adjust_i = 2'b01;
            end
        end
        else
        begin
            fdiv_frac_en_i     = 1'b0;
            psoffsetf_i        = 3'b000;
            fdiv_frac_adjust_i = 2'b00;
        end

        mem0  = {ratio0_i, duty0_i};
        mem1  = {ratio0_frac_i, psoffset0_i, odiv0_fphase_i, odiv0_cphase_i};
        mem2  = {10'h0, odiv0_frac_adjust_i, odiv0_frac_en_i, muxsel0_i, muxsel0_en_i};
        mem3  = {ratio1_i, duty1_i};
        mem4  = {3'h0, muxsel1_i, muxsel1_en_i, odiv1_fphase_i, odiv1_cphase_i};
        mem5  = {ratio2_i, duty2_i};
        mem6  = {3'h0, muxsel2_i, muxsel2_en_i, odiv2_fphase_i, odiv2_cphase_i};
        mem7  = {ratio3_i, duty3_i};
        mem8  = {3'h0, muxsel3_i, muxsel3_en_i, odiv3_fphase_i, odiv3_cphase_i};
        mem9  = {ratio4_i, duty4_i};
        mem10 = {3'h0, muxsel4_i, muxsel4_en_i, odiv4_fphase_i, odiv4_cphase_i};
        mem11 = {ratio5_i, duty5_i};
        mem12 = {3'h0, muxsel5_i, muxsel5_en_i, odiv5_fphase_i, odiv5_cphase_i};
        mem13 = {ratio6_i, duty6_i};
        mem14 = {3'h0, muxsel6_i, muxsel6_en_i, odiv6_fphase_i, odiv6_cphase_i};
        mem15 = {ratiof_i, dutyf_i};
        mem16 = {ratiof_frac_i, psoffsetf_i, fdiv_fphase_i, fdiv_cphase_i};
        mem17 = {10'h0, fdiv_frac_adjust_i, fdiv_frac_en_i, muxself_i, muxself_en_i};
        mem18 = {8'h0, ratioi_i};
        mem19 = {8'h0, ratiom_i};
        mem20 = {2'b00, vctrl_i, cp_selbias_i, cp_selbias_i, cp_base_i, cp_cur_i, lpf_r_i, lpf_c_i};
        mem21 = {10'h0, lockfilter_pd_i, lock_set_i};
    end

    assign ratioi = mem18[7:0];
    assign ratiom = mem19[7:0];
    assign ratiof = mem15[15:8];
    assign ratio0 = mem0[15:8];
    assign ratio1 = mem3[15:8];
    assign ratio2 = mem5[15:8];
    assign ratio3 = mem7[15:8];
    assign ratio4 = mem9[15:8];
    assign ratio5 = mem11[15:8];
    assign ratio6 = mem13[15:8];
    assign dutyf  = mem15[7:0];
    assign duty0  = mem0[7:0];
    assign duty1  = mem3[7:0];
    assign duty2  = mem5[7:0];
    assign duty3  = mem7[7:0];
    assign duty4  = mem9[7:0];
    assign duty5  = mem11[7:0];
    assign duty6  = mem13[7:0];
    assign odiv0_cphase = mem1[6:0];
    assign odiv1_cphase = mem4[6:0];
    assign odiv2_cphase = mem6[6:0];
    assign odiv3_cphase = mem8[6:0];
    assign odiv4_cphase = mem10[6:0];
    assign odiv5_cphase = mem12[6:0];
    assign odiv6_cphase = mem14[6:0];
    assign fdiv_cphase  = mem16[6:0];
    assign odiv0_fphase = mem1[9:7];
    assign odiv1_fphase = mem4[9:7];
    assign odiv2_fphase = mem6[9:7];
    assign odiv3_fphase = mem8[9:7];
    assign odiv4_fphase = mem10[9:7];
    assign odiv5_fphase = mem12[9:7];
    assign odiv6_fphase = mem14[9:7];
    assign fdiv_fphase  = mem16[9:7];
    assign ratio0_frac  = mem1[15:13];
    assign ratiof_frac  = mem16[15:13];
    assign psoffset0    = mem1[12:10];
    assign psoffsetf    = mem16[12:10];
    assign muxsel0_en = mem2[0];
    assign muxsel1_en = mem4[10];
    assign muxsel2_en = mem6[10];
    assign muxsel3_en = mem8[10];
    assign muxsel4_en = mem10[10];
    assign muxsel5_en = mem12[10];
    assign muxsel6_en = mem14[10];
    assign muxself_en = mem17[0];
    assign muxsel0    = mem2[2:1];
    assign muxsel1    = mem4[12:11];
    assign muxsel2    = mem6[12:11];
    assign muxsel3    = mem8[12:11];
    assign muxsel4    = mem10[12:11];
    assign muxsel5    = mem12[12:11];
    assign muxsel6    = mem14[12:11];
    assign muxself    = mem17[2:1];
    assign odiv0_frac_en     = mem2[3];
    assign fdiv_frac_en      = mem17[3];
    assign odiv0_frac_adjust = mem2[5:4];
    assign fdiv_frac_adjust  = mem17[5:4];
///////////////////////////////////////////////////////
    wire rst_n;
    reg inner_rstn;
///////////////////////////////////////////////////////
    wire clk_in;
///////////////////////////////////////////////////////
    reg clk_in_first_time, clk_fb_first_time;
    realtime clk_in_first_edge, clk_fb_first_edge;
    reg adjust;
    realtime fb_route_delay, virtual_delay1;
    integer tmp_ratio;
    realtime tmp_delay, real_delay;
///////////////////////////////////////////////////////
    reg clk_test;
    reg clkref_wo, clkfb_wo;
    realtime clkref_test_time1 , clkref_test_time2, clkref_test_time3;
    realtime clkfb_rtime_last, clkfb_rtime_next;
    realtime clkfb_test_time1 , clkfb_test_time2, clkfb_test_time3;
    wire clkwo;
///////////////////////////////////////////////////////
    wire [7:0] idivider, mdivider, fdivider, divider0, divider1, divider2, divider3, divider4, divider5, divider6;
    real fsdiv_set_int, fbdiv_set_int;

    wire rstanalog_n;
    realtime clkin_rtime_last, clkin_rtime_next;
    realtime clkin_time, clkin_time1, clkin_time2, clkin_time3;
    reg clkout_lock;
    realtime vcoclk_period, vcoclk_period_half;
    realtime clkout0_time, clkout1_time, clkout2_time, clkout3_time, clkout4_time, clkout5_time, clkout6_time, clkoutf_time;
    integer  vcoclk_period_amp;
    realtime vcoclk_period_real, vcoclk_period_dev;

    reg done;
    integer idiv_set;
    integer fdiv_set;
    integer swap_set;
    integer midd_set;
    integer fdiv_int;
    realtime offset;

    real cnt_fdiv;
    reg clk_gate, inner_clk;
    reg vcoclk;

    real new_delay;
    wire adjust_dly, frac_restart;
///////////////////////////////////////////////////////
    wire clk_lock;
    reg [2:0] cnt_clkfb;
    reg start_clk;
    reg [10:0] cnt_lock;
    reg lock_wait;
    reg lock_reg;
///////////////////////////////////////////////////////
    reg [5:0] dps_cnt;
    reg dps_cnt_finish;
    reg dps_done_reg;
    integer dps_done_cnt;
    wire [63:0] vcoclk_dps_dly;
    reg vcoclk_dps_adjust;
    integer dps_cnt_dly0, dps_cnt_dly1;
    wire vcoclk_dps;
///////////////////////////////////////////////////////
    reg odiv0_clkin, odiv1_clkin, odiv2_clkin, odiv3_clkin, odiv4_clkin, odiv5_clkin, odiv6_clkin, fdiv_clkin;
    reg [7:0] odiv0_counter, odiv1_counter, odiv2_counter, odiv3_counter, odiv4_counter, odiv5_counter, odiv6_counter, fdiv_counter;
    reg odiv0_out_reg, odiv1_out_reg, odiv2_out_reg, odiv3_out_reg, odiv4_out_reg, odiv5_out_reg, odiv6_out_reg, fdiv_out_reg;
    wire odiv0_out, odiv1_out, odiv2_out, odiv3_out, odiv4_out, odiv5_out, odiv6_out, fdiv_out;

    wire odiv0_int_out, fdiv_int_out;
    wire [2:0] divider0_frac, fdivider_frac;
    integer odiv0_p_int, odiv0_hp_frac, odiv0_lp_frac, fdiv_p_int, fdiv_hp_frac, fdiv_lp_frac;
    real odiv0_frac_hp, odiv0_frac_lp, fdiv_frac_hp, fdiv_frac_lp;
    integer i,j;
    reg odiv0_frac_out, fdiv_frac_out;
///////////////////////////////////////////////////////
    realtime vco_fphase_delay0, vco_fphase_delay1, vco_fphase_delay2, vco_fphase_delay3, vco_fphase_delay4, vco_fphase_delay5, vco_fphase_delay6, vco_fphase_delayf;
    integer cphase0, cphase1, cphase2, cphase3, cphase4, cphase5, cphase6, cphasef;
    realtime cphase_delay0, cphase_delay1, cphase_delay2, cphase_delay3, cphase_delay4, cphase_delay5, cphase_delay6, cphase_delayf;
    reg odiv0_out_delay1, odiv1_out_delay1, odiv2_out_delay1, odiv3_out_delay1, odiv4_out_delay1, odiv5_out_delay1, odiv6_out_delay1, fdiv_out_delay1;
    reg odiv0_out_delay, odiv1_out_delay, odiv2_out_delay, odiv3_out_delay, odiv4_out_delay, odiv5_out_delay, odiv6_out_delay, fdiv_out_delay;
///////////////////////////////////////////////////////
    reg [2:0] clk_out0_gate, clk_out1_gate, clk_out2_gate, clk_out3_gate, clk_out4_gate, clk_out5_gate, clk_out6_gate, clk_outf_gate;
    wire clkout0_gate, clkout1_gate, clkout2_gate, clkout3_gate, clkout4_gate, clkout5_gate, clkout6_gate, clkoutf_gate;
///////////////////////////////////////////////////////
    reg [1:0] apb_rstn_sync;
    reg ready;
    reg [15:0] rdata;
///////////////////////////////////////////////////////
    initial
    begin
        inner_rstn = 1'b0;
        clk_in_first_time = 1'b0;
        clk_fb_first_time = 1'b0;
        clk_in_first_edge = 0.0;
        clk_fb_first_edge = 0.0;
        fb_route_delay = 0.0;
        tmp_ratio      = 0;
        tmp_delay      = 0.0;
        real_delay     = 0.0;
        clk_test = 1'b0;
        fsdiv_set_int = 0;
        fbdiv_set_int = 0;
        done = 1'b0;
        idiv_set = 0;
        fdiv_set = 0;
        swap_set = 0;
        midd_set = 0;
        fdiv_int = 0;
        offset = 0;
        cnt_fdiv  = 0;
        clk_gate  = 1'b1;
        inner_clk = 1'b0;
        vcoclk    = 1'b0;
        i = 1;
        j = 1;
        vco_fphase_delay0 = 0.0;
        vco_fphase_delay1 = 0.0;
        vco_fphase_delay2 = 0.0;
        vco_fphase_delay3 = 0.0;
        vco_fphase_delay4 = 0.0;
        vco_fphase_delay5 = 0.0;
        vco_fphase_delay6 = 0.0;
        vco_fphase_delayf = 0.0;
        cphase_delay0 = 0.0;
        cphase_delay1 = 0.0;
        cphase_delay2 = 0.0;
        cphase_delay3 = 0.0;
        cphase_delay4 = 0.0;
        cphase_delay5 = 0.0;
        cphase_delay6 = 0.0;
        cphase_delayf = 0.0;
        odiv0_out_delay1 = 1'b0;
        odiv1_out_delay1 = 1'b0;
        odiv2_out_delay1 = 1'b0;
        odiv3_out_delay1 = 1'b0;
        odiv4_out_delay1 = 1'b0;
        odiv5_out_delay1 = 1'b0;
        odiv6_out_delay1 = 1'b0;
        fdiv_out_delay1  = 1'b0;
        odiv0_out_delay  = 1'b0;
        odiv1_out_delay  = 1'b0;
        odiv2_out_delay  = 1'b0;
        odiv3_out_delay  = 1'b0;
        odiv4_out_delay  = 1'b0;
        odiv5_out_delay  = 1'b0;
        odiv6_out_delay  = 1'b0;
        fdiv_out_delay   = 1'b0;
        clk_out0_gate = 3'b000;
        clk_out1_gate = 3'b000;
        clk_out2_gate = 3'b000;
        clk_out3_gate = 3'b000;
        clk_out4_gate = 3'b000;
        clk_out5_gate = 3'b000;
        clk_out6_gate = 3'b000;
        clk_outf_gate = 3'b000;
        #1;
        inner_rstn = 1'b1;
        clk_in_first_time = 1'b1;
        clk_fb_first_time = 1'b1;
    end
///////////////////////////////////////////////////////
////RESET//////////////////////////////////////////////
    assign rst_n = ~(PLL_PWD | RST) & inner_rstn;
///////////////////////////////////////////////////////
////INPUT_CLK_SEL//////////////////////////////////////
    assign clk_in = (CLKIN_SEL == 1'b0) ? CLKIN1 : CLKIN2;
///////////////////////////////////////////////////////
////FBCK_DELAY/////////////////////////////////////////
    always @(posedge clk_in or negedge rst_n)
    begin
        if(!rst_n)
        begin
            clk_in_first_time = 1'b1;
            clk_in_first_edge = 0.0;
        end
        else
        begin
            if(clk_in_first_time == 1'b1)
                clk_in_first_edge = $realtime;
            clk_in_first_time = 1'b0;
        end
    end

    always @(posedge CLKFB or negedge rst_n)
    begin
        if(!rst_n)
        begin
            clk_fb_first_time = 1'b1;
            clk_fb_first_edge = 0.0;
        end
        else
        begin
            if(clk_fb_first_time == 1'b1)
                clk_fb_first_edge = $realtime;
            clk_fb_first_time = 1'b0;
        end
    end
///////////////////////////////////////////////////////
////CLK_TEST///////////////////////////////////////////
    always #200 clk_test = ~clk_test;

    always @(posedge clk_test or negedge rst_n)
    begin
        if(!rst_n)
        begin
            clkref_wo <= 1'b0;
            clkref_test_time1 = 0;
            clkref_test_time2 = 0;
            clkref_test_time3 = 0;
        end
        else
        begin
            clkref_test_time3 = clkref_test_time2;
            clkref_test_time2 = clkref_test_time1;
            clkref_test_time1 = clkin_rtime_next;
            if(clkref_test_time3 == clkref_test_time1)
                clkref_wo <= 1'b1;
            else
                clkref_wo <= 1'b0;
        end
    end

    always @(posedge CLKFB or negedge rst_n)
    begin
        if(!rst_n)
        begin
            clkfb_rtime_last = 0.0;
            clkfb_rtime_next = 0.0;
        end
        else
        begin
            clkfb_rtime_last = clkin_rtime_next;
            clkfb_rtime_next = $realtime;
        end
    end

    always @(posedge clk_test or negedge rst_n)
    begin
        if(!rst_n)
        begin
            clkfb_wo <= 1'b0;
            clkfb_test_time3 = 0;
            clkfb_test_time2 = 0;
            clkfb_test_time1 = 0;
        end
        else
        begin
            if(clk_fb_first_time == 1'b0)
            begin
                clkfb_test_time3 = clkfb_test_time2;
                clkfb_test_time2 = clkfb_test_time1;
                clkfb_test_time1 = clkfb_rtime_next;
                if(clkfb_test_time3 == clkfb_test_time1)
                    clkfb_wo <= 1'b1;
                else
                    clkfb_wo <= 1'b0;
            end
        end
    end

    assign clkwo = clkref_wo | clkfb_wo;
///////////////////////////////////////////////////////
////PLL_ANALOG/////////////////////////////////////////
////FEEDBACK_DIVIDER_CAL///////////////////////////////
    assign idivider = ratioi;
    assign mdivider = ratiom;
    assign fdivider = ratiof;
    assign divider0 = ratio0;
    assign divider1 = ratio1;
    assign divider2 = ratio2;
    assign divider3 = ratio3;
    assign divider4 = ratio4;
    assign divider5 = ratio5;
    assign divider6 = ratio6;

    always @(*)
    begin
    	if((INTERNAL_FB == "CLKOUTF" || EXTERNAL_FB == "CLKOUTF") && fdiv_frac_en == 1'b0)
            fsdiv_set_int = fdivider;
    	else if((INTERNAL_FB == "CLKOUTF" || EXTERNAL_FB == "CLKOUTF") && fdiv_frac_en == 1'b1)
            fsdiv_set_int = fdivider + ratiof_frac * 0.125;
        else if((INTERNAL_FB == "CLKOUT0" || EXTERNAL_FB == "CLKOUT0") && odiv0_frac_en == 1'b0)
            fsdiv_set_int = divider0;
        else if((INTERNAL_FB == "CLKOUT0" || EXTERNAL_FB == "CLKOUT0") && odiv0_frac_en == 1'b1)
            fsdiv_set_int = divider0 + ratio0_frac * 0.125;
        else if(INTERNAL_FB == "CLKOUT1" || EXTERNAL_FB == "CLKOUT1")
            fsdiv_set_int = divider1;
        else if(INTERNAL_FB == "CLKOUT2" || EXTERNAL_FB == "CLKOUT2")
            fsdiv_set_int = divider2;
        else if(INTERNAL_FB == "CLKOUT3" || EXTERNAL_FB == "CLKOUT3")
            fsdiv_set_int = divider3;
        else if(INTERNAL_FB == "CLKOUT4" || EXTERNAL_FB == "CLKOUT4")
            fsdiv_set_int = divider4;
        else if(INTERNAL_FB == "CLKOUT5" || EXTERNAL_FB == "CLKOUT5")
            fsdiv_set_int = divider5;
        else if(INTERNAL_FB == "CLKOUT6" || EXTERNAL_FB == "CLKOUT6")
            fsdiv_set_int = divider6;
    end

    always @(*)
    begin
        fbdiv_set_int = mdivider * fsdiv_set_int;
    end
////PLL_VCO_CAL////////////////////////////////////////
    assign rstanalog_n = rst_n;

    always @(posedge clk_in or negedge rstanalog_n)
    begin
        if(!rstanalog_n)
        begin
            clkin_rtime_last = 0.0;
            clkin_rtime_next = 0.0;
            clkin_time  <= 0.0;
            clkin_time1 <= 0.0;
            clkin_time2 <= 0.0;
            clkin_time3 <= 0.0;
            clkout_lock <= 0.0;
            vcoclk_period <= 1'b0;
            vcoclk_period_half <= 0.0;
            clkout0_time       <= 0.0;
            clkout1_time       <= 0.0;
            clkout2_time       <= 0.0;
            clkout3_time       <= 0.0;
            clkout4_time       <= 0.0;
            vcoclk_period_amp  <= 0.0;
            vcoclk_period_real <= 0.0;
            vcoclk_period_dev  <= 0.0;
        end
        else
        begin
            clkin_rtime_last = clkin_rtime_next;
            clkin_rtime_next = $realtime;
            if(clkin_rtime_last > 0)
            begin
                clkin_time  <= clkin_rtime_next-clkin_rtime_last;
                clkin_time1 <= clkin_time;
                clkin_time2 <= clkin_time1;
                clkin_time3 <= clkin_time2;
            end
            if(clkin_time > 0)
            begin
                clkout_lock <= (clkin_time  > 0) &&
                               (clkin_time1 > 0) &&
                               (clkin_time2 > 0) &&
                               (clkin_time3 > 0) &&
                               ((clkin_time - clkin_time1)  < 0.0001) &&
                               ((clkin_time1 - clkin_time)  < 0.0001) &&
                               ((clkin_time1 - clkin_time2) < 0.0001) &&
                               ((clkin_time2 - clkin_time1) < 0.0001) &&
                               ((clkin_time2 - clkin_time3) < 0.0001) &&
                               ((clkin_time3 - clkin_time2) < 0.0001);
            end
            if(clkin_time > 0)
            begin
                vcoclk_period      = (clkin_time * idivider) / fbdiv_set_int;
                vcoclk_period_half = vcoclk_period / 2;
                clkout0_time       = vcoclk_period * divider0;
                clkout1_time       = vcoclk_period * divider1;
                clkout2_time       = vcoclk_period * divider2;
                clkout3_time       = vcoclk_period * divider3;
                clkout4_time       = vcoclk_period * divider4;
                clkout5_time       = vcoclk_period * divider5;
                clkout6_time       = vcoclk_period * divider6;
                clkoutf_time       = vcoclk_period * fdivider;
                vcoclk_period_amp  = vcoclk_period_half * 1000000;
                vcoclk_period_real = vcoclk_period_amp / 1000000.0;
                vcoclk_period_dev  = (clkin_time - (vcoclk_period_real * 2 * fbdiv_set_int) / idivider) / 2;
            end
        end
    end

    always @(*)
    begin
        if(!rst_n)
        begin
            done = 1'b0;
            idiv_set = 0;
            fdiv_set = 0;
            swap_set = 0;
            midd_set = 0;
            offset = 0;
        end
        else
        begin
            idiv_set = idivider;
            fdiv_set = $rtoi(fbdiv_set_int);
            while(!done)
            begin
                if(idiv_set < fdiv_set)
                begin
                    swap_set = idiv_set;
                    idiv_set = fdiv_set;
                    fdiv_set = swap_set;
                end
                else
                    if(fdiv_set != 0)
                        idiv_set = idiv_set - fdiv_set;
                    else
                    begin
                        done = 1;
                        midd_set = idiv_set;
                    end
            end
        end
    end

    always @(*)
    begin
        if(!rst_n)
        begin
            fdiv_int = 0;
            offset = 0;
        end
        else
            begin
                fdiv_int = midd_set;
                offset = vcoclk_period_dev * idivider/midd_set;
            end
    end

    always @(clkout_lock or inner_clk or clkwo)
    begin
        if(clkout_lock == 1'b0 || clkwo == 1'b1)
        begin
            inner_clk <= 1'b0;
            clk_gate  <= 1'b1;
            cnt_fdiv   = 0;
        end
        else
            if(clk_gate == 1)
            begin
                inner_clk <= 1'b1;
                clk_gate  <= 1'b0;
                cnt_fdiv   = 0;
            end
            else
            begin
                cnt_fdiv = cnt_fdiv + 1;
                if(cnt_fdiv == $rtoi(fbdiv_set_int)/fdiv_int)
                begin
                    inner_clk <= #(vcoclk_period_half + offset) ~inner_clk;
                    cnt_fdiv = 0;
                end
                else
                    inner_clk <= #vcoclk_period_half ~inner_clk;
            end
    end

    always @(posedge clk_in or CLKFB or negedge rst_n)
    begin
        if(!rst_n)
        begin
            adjust <= 1'b1;
            fb_route_delay = 0.0;
            tmp_ratio  = 0;
            tmp_delay  = 0.0;
            real_delay = 0.0;
        end
        else
            if(adjust == 1'b1)
            begin
                fb_route_delay = clk_fb_first_edge - clk_in_first_edge;
                if((clkin_time > 0) && (fb_route_delay > 0))
                begin
                    tmp_ratio  = fb_route_delay / clkin_time;
                    tmp_delay  = fb_route_delay - (clkin_time * tmp_ratio);
                    real_delay = clkin_time - tmp_delay;
                    adjust <= 1'b0;
                end
            end
    end

    always @(inner_clk)
    begin
        if(EXTERNAL_FB == "CLKOUTF" || EXTERNAL_FB == "CLKOUT0" || EXTERNAL_FB == "CLKOUT1" || EXTERNAL_FB == "CLKOUT2" || EXTERNAL_FB == "CLKOUT3" || EXTERNAL_FB == "CLKOUT4" || EXTERNAL_FB == "CLKOUT5" || EXTERNAL_FB == "CLKOUT6")
            vcoclk <= #real_delay inner_clk;
        else
            vcoclk <= inner_clk;
    end

    always @(*)
    begin
        if(!rst_n)
            new_delay = 0;
        else
            new_delay = (clkin_time * idivider) / mdivider;
    end

    assign #(real_delay + new_delay) adjust_dly = adjust; 
    assign frac_restart = ~adjust & adjust_dly;
///////////////////////////////////////////////////////
////PLL_LOCK///////////////////////////////////////////
    assign clk_lock = (INTERNAL_FB == "DISABLE") ? CLKFB : clk_in;

    always @(posedge clk_lock or negedge rstanalog_n or clk_gate)
    begin
        if(!rstanalog_n)
        begin
            start_clk <= 1'b0;
            cnt_clkfb <= 2'b00;
        end
        else
            if(!clk_gate)
                if(cnt_clkfb == 2'b11)
                    start_clk = 1'b1;
                else
                    cnt_clkfb = cnt_clkfb + 1'b1;
            else
            begin
                start_clk <= 1'b0;
                cnt_clkfb <= 2'b00;
            end
    end

    always @(posedge clk_in or negedge rstanalog_n or clk_gate)
    begin
        if(!rstanalog_n)
        begin
            cnt_lock  <= 8'h1;
            lock_wait <= 1'b0;
        end
        else
            if(!clk_gate && start_clk)
                if(cnt_lock == idivider * 3)
                    lock_wait <= 1'b1;
                else
                    cnt_lock <= cnt_lock + 1'b1;
            else
            begin
                cnt_lock <= 8'h1;
                lock_wait <= 1'b0;
            end
    end

    always @(posedge clk_in or negedge rst_n or clk_gate)
    begin
        if(!rst_n)
            lock_reg <= 1'b0;
        else
            if(LOCK_MODE == 1'b0)
                if(!clk_gate)
                    lock_reg <= lock_wait;
                else
                    lock_reg <= 1'b0;
            else
                lock_reg <= lock_reg | lock_wait;
    end

    assign LOCK = lock_reg;
///////////////////////////////////////////////////////
////DPS////////////////////////////////////////////////
    always @(posedge DPS_CLK or negedge rst_n)
    begin
        if(!rst_n)
        begin
            dps_cnt <= dps_init;
            dps_cnt_finish <= 1'b0;
        end
        else
        begin
            if(div_dps_en == 1'b1 && DPS_EN == 1'b1)
                if(DPS_DIR == 1'b0)
                begin
                    if(dps_cnt < 6'd63)
                        dps_cnt <= dps_cnt + 1'b1;
                    else
                        dps_cnt <= 0;

                    dps_cnt_finish <= 1'b1;
                end
                else
                    if(DPS_DIR == 1'b1)
                    begin
                        if(dps_cnt > 0)
                            dps_cnt <= dps_cnt - 1'b1;
                        else
                            dps_cnt <= 6'd63;

                        dps_cnt_finish <= 1'b1;
                    end

             if(dps_done_reg == 1'b1)
                  dps_cnt_finish <= 1'b0;
        end
    end

    always @(posedge DPS_CLK or negedge rst_n)
    begin
        if(!rst_n)
        begin
            dps_done_cnt <= 1;
            dps_done_reg <= 1'b0;
        end
        else
            if(dps_cnt_finish)
                if(dps_done_cnt < 13)
                begin
                    dps_done_cnt <= dps_done_cnt + 1;
                    dps_done_reg <= 1'b0;
                end
                else
                begin
                    dps_done_cnt <= 0;
                    dps_done_reg <= 1'b1;
                end
    end

    assign DPS_DONE = dps_done_reg;

    assign vcoclk_dps_dly[0] = vcoclk;

    genvar gen_j;

    generate
        for(gen_j=1; gen_j<64; gen_j=gen_j+1'b1)
        begin
            assign #(vcoclk_period/64) vcoclk_dps_dly[gen_j] = vcoclk_dps_dly[gen_j-1];
        end
    endgenerate

    always @(*)
    begin
        if(DPS_DIR == 1'b1)
            vcoclk_dps_adjust = vcoclk_dps_dly[dps_cnt];
        else
            if(dps_cnt == 6'd63)
                vcoclk_dps_adjust = vcoclk_dps_dly[0];
            else
                vcoclk_dps_adjust = vcoclk_dps_dly[dps_cnt + 1];
    end

    always @(negedge vcoclk_dps_adjust or negedge rst_n)
    begin
        if(!rst_n)
        begin
            dps_cnt_dly0 = dps_cnt;
            dps_cnt_dly1 = dps_cnt;
        end
        else
        begin
            dps_cnt_dly0 <= dps_cnt;
            dps_cnt_dly1 <= dps_cnt_dly0;
        end
    end

    assign vcoclk_dps = vcoclk_dps_dly[dps_cnt_dly1];
///////////////////////////////////////////////////////
////PLL_ODIV///////////////////////////////////////////
////ODIV0//////////////////////////////////////////////
    always @(*)
    begin
        if(muxsel0_en)
            case(muxsel0)
                2'b00: odiv0_clkin = vcoclk;
                2'b01: odiv0_clkin = vcoclk_dps;
                default: odiv0_clkin = 1'b0;
            endcase
        else
            odiv0_clkin = 1'b0;
    end

    always @(posedge odiv0_clkin or negedge odiv0_clkin or negedge rst_n)
    begin
        if(!rst_n)
        begin
            odiv0_counter <= 8'h0;
            odiv0_out_reg <= 1'b0;
        end
        else
        begin
            if(divider0 == 8'h1)
            begin
                odiv0_counter <= 8'h0;
                odiv0_out_reg <= 1'b0;
            end
            else
            begin
                if(odiv0_counter < ({divider0, 1'b0} - 1'b1))
                    odiv0_counter <= odiv0_counter + 1'b1;
                else
                    odiv0_counter <= 8'h0;

                if(odiv0_counter < duty0)
                    odiv0_out_reg <= 1'b1;
                else
                    odiv0_out_reg <= 1'b0;
            end
        end
    end

    assign odiv0_int_out = (divider0 == 8'h1) ? odiv0_clkin : odiv0_out_reg;

    assign divider0_frac = ratio0_frac;

    always @(*)
    begin
        if(odiv0_frac_en == 1'b1)
        begin
            odiv0_p_int = divider0 / 2;

            if(!divider0[0])
                if(!divider0_frac[0])
                begin
                    odiv0_hp_frac = divider0_frac / 2;
                    odiv0_lp_frac = divider0_frac / 2;
                end
                else
                begin
                    odiv0_hp_frac = (divider0_frac + 1'b1) / 2;
                    odiv0_lp_frac = divider0_frac / 2;
                end
            else
                if(!divider0_frac[0])
                begin
                    odiv0_hp_frac = divider0_frac / 2 + 3'b100;
                    odiv0_lp_frac = divider0_frac / 2 + 3'b100;
                end
                else
                begin
                    odiv0_hp_frac = divider0_frac / 2 + 3'b101;
                    odiv0_lp_frac = divider0_frac / 2 + 3'b100;
                end
        end
        else
        begin
             odiv0_p_int   = 0;
             odiv0_hp_frac = 0;
             odiv0_lp_frac = 0;
        end
    end

    always @(*)
    begin
        odiv0_frac_hp = vcoclk_period * odiv0_p_int + (vcoclk_period * odiv0_hp_frac) / 8;
        odiv0_frac_lp = vcoclk_period * odiv0_p_int + (vcoclk_period * odiv0_lp_frac) / 8;
    end

    always @(clk_gate or odiv0_frac_out or negedge rst_n)
    begin
        if(!rst_n)
            odiv0_frac_out <= 1'b0;
        else
            if(!clk_gate && odiv0_frac_en && odiv0_dps_en == 1'b0)
            begin
                odiv0_frac_out <= 1'b1;
                for(i = 1; i < 8; i = i+1)
                begin: loop1
                    if(frac_restart)
                    begin
                        #(real_delay);
                        #(odiv0_frac_hp) odiv0_frac_out <= 1'b0;
                        #(odiv0_frac_lp) odiv0_frac_out <= 1'b1;
                    end
                    else
                    begin
                        #(odiv0_frac_hp) odiv0_frac_out <= 1'b0;
                        #(odiv0_frac_lp) odiv0_frac_out <= 1'b1;
                    end
                end
                #(odiv0_frac_hp) odiv0_frac_out <= 1'b0;
                #(odiv0_frac_lp);
                i = 1;
                odiv0_frac_out <= 1'b1;
            end
            else
                odiv0_frac_out <= 1'b0;
    end

    assign odiv0_out = (odiv0_frac_en) ? odiv0_frac_out : odiv0_int_out;
////ODIV1//////////////////////////////////////////////
    always @(*)
    begin
        if(muxsel1_en)
            case(muxsel1)
                2'b00: odiv1_clkin = vcoclk;
                2'b01: odiv1_clkin = vcoclk_dps;
                default: odiv1_clkin = 1'b0;
            endcase
        else
            odiv1_clkin = 1'b0;
    end

    always @(posedge odiv1_clkin or negedge odiv1_clkin or negedge rst_n)
    begin
        if(!rst_n)
        begin
            odiv1_counter <= 8'h0;
            odiv1_out_reg <= 1'b0;
        end
        else
        begin
            if(divider1 == 8'h1)
            begin
                odiv1_counter <= 8'h0;
                odiv1_out_reg <= 1'b0;
            end
            else
            begin
                if(odiv1_counter < ({divider1, 1'b0} - 1'b1))
                    odiv1_counter <= odiv1_counter + 1'b1;
                else
                    odiv1_counter <= 8'h0;

                if(odiv1_counter < duty1)
                    odiv1_out_reg <= 1'b1;
                else
                    odiv1_out_reg <= 1'b0;
            end
        end
    end

    assign odiv1_out = (divider1 == 8'h1) ? odiv1_clkin : odiv1_out_reg;
////ODIV2//////////////////////////////////////////////
    always @(*)
    begin
        if(muxsel2_en)
            case(muxsel2)
                2'b00: odiv2_clkin = vcoclk;
                2'b01: odiv2_clkin = vcoclk_dps;
                default: odiv2_clkin = 1'b0;
            endcase
        else
            odiv2_clkin = 1'b0;
    end

    always @(posedge odiv2_clkin or negedge odiv2_clkin or negedge rst_n)
    begin
        if(!rst_n)
        begin
            odiv2_counter <= 8'h0;
            odiv2_out_reg <= 1'b0;
        end
        else
        begin
            if(divider2 == 8'h1)
            begin
                odiv2_counter <= 8'h0;
                odiv2_out_reg <= 1'b0;
            end
            else
            begin
                if(odiv2_counter < ({divider2, 1'b0} - 1'b1))
                    odiv2_counter <= odiv2_counter + 1'b1;
                else
                    odiv2_counter <= 8'h0;

                if(odiv2_counter < duty2)
                    odiv2_out_reg <= 1'b1;
                else
                    odiv2_out_reg <= 1'b0;
            end
        end
    end

    assign odiv2_out = (divider2 == 8'h1) ? odiv2_clkin : odiv2_out_reg;
////ODIV3//////////////////////////////////////////////
    always @(*)
    begin
        if(muxsel3_en)
            case(muxsel3)
                2'b00: odiv3_clkin = vcoclk;
                2'b01: odiv3_clkin = vcoclk_dps;
                default: odiv3_clkin = 1'b0;
            endcase
        else
            odiv3_clkin = 1'b0;
    end

    always @(posedge odiv3_clkin or negedge odiv3_clkin or negedge rst_n)
    begin
        if(!rst_n)
        begin
            odiv3_counter <= 8'h0;
            odiv3_out_reg <= 1'b0;
        end
        else
        begin
            if(divider3 == 8'h1)
            begin
                odiv3_counter <= 8'h0;
                odiv3_out_reg <= 1'b0;
            end
            else
            begin
                if(odiv3_counter < ({divider3, 1'b0} - 1'b1))
                    odiv3_counter <= odiv3_counter + 1'b1;
                else
                    odiv3_counter <= 8'h0;

                if(odiv3_counter < duty3)
                    odiv3_out_reg <= 1'b1;
                else
                    odiv3_out_reg <= 1'b0;
            end
        end
    end

    assign odiv3_out = (divider3 == 8'h1) ? odiv3_clkin : odiv3_out_reg;
////ODIV4//////////////////////////////////////////////
    always @(*)
    begin
        if(muxsel4_en)
            case(muxsel4)
                2'b00: odiv4_clkin = vcoclk;
                2'b01: odiv4_clkin = vcoclk_dps;
                default: odiv4_clkin = 1'b0;
            endcase
        else
            odiv4_clkin = 1'b0;
    end


    always @(posedge odiv4_clkin or negedge odiv4_clkin or negedge rst_n)
    begin
        if(!rst_n)
        begin
            odiv4_counter <= 8'h0;
            odiv4_out_reg <= 1'b0;
        end
        else
        begin
            if(divider4 == 8'h1)
            begin
                odiv4_counter <= 8'h0;
                odiv4_out_reg <= 1'b0;
            end
            else
            begin
                if(odiv4_counter < ({divider4, 1'b0} - 1'b1))
                    odiv4_counter <= odiv4_counter + 1'b1;
                else
                    odiv4_counter <= 8'h0;

                if(odiv4_counter < duty4)
                    odiv4_out_reg <= 1'b1;
                else
                    odiv4_out_reg <= 1'b0;
            end
        end
    end

    assign odiv4_out = (divider4 == 8'h1) ? odiv4_clkin : odiv4_out_reg;
////odiv5////////////////////////////////////////////
    always @(*)
    begin
        if(muxsel5_en)
            case(muxsel5)
                2'b00: odiv5_clkin = vcoclk;
                2'b01: odiv5_clkin = vcoclk_dps;
                2'b10: odiv5_clkin = odiv6_out;
                default: odiv5_clkin = 1'b0;
            endcase
        else
            odiv5_clkin = 1'b0;
    end

    always @(posedge odiv5_clkin or negedge odiv5_clkin or negedge rst_n)
    begin
        if(!rst_n)
        begin
            odiv5_counter <= 8'h0;
            odiv5_out_reg <= 1'b0;
        end
        else
        begin
            if(divider5 == 8'h1)
            begin
                odiv5_counter <= 8'h0;
                odiv5_out_reg <= 1'b0;
            end
            else
            begin
                if(odiv5_counter < ({divider5, 1'b0} - 1'b1))
                    odiv5_counter <= odiv5_counter + 1'b1;
                else
                    odiv5_counter <= 8'h0;

                if(odiv5_counter < duty5)
                    odiv5_out_reg <= 1'b1;
                else
                    odiv5_out_reg <= 1'b0;
            end
        end
    end

    assign odiv5_out = (divider5 == 8'h1) ? odiv5_clkin : odiv5_out_reg;
////odiv6////////////////////////////////////////////
    always @(*)
    begin
        if(muxsel6_en)
            case(muxsel6)
                2'b00: odiv6_clkin = vcoclk;
                2'b01: odiv6_clkin = vcoclk_dps;
                default: odiv6_clkin = 1'b0;
            endcase
        else
            odiv6_clkin = 1'b0;
    end

    always @(posedge odiv6_clkin or negedge odiv6_clkin or negedge rst_n)
    begin
        if(!rst_n)
        begin
            odiv6_counter <= 8'h0;
            odiv6_out_reg <= 1'b0;
        end
        else
        begin
            if(divider6 == 8'h1)
            begin
                odiv6_counter <= 8'h0;
                odiv6_out_reg <= 1'b0;
            end
            else
            begin
                if(odiv6_counter < ({divider6, 1'b0} - 1'b1))
                    odiv6_counter <= odiv6_counter + 1'b1;
                else
                    odiv6_counter <= 8'h0;

                if(odiv6_counter < duty6)
                    odiv6_out_reg <= 1'b1;
                else
                    odiv6_out_reg <= 1'b0;
            end
        end
    end

    assign odiv6_out = (divider6 == 8'h1) ? odiv6_clkin : odiv6_out_reg;
////FDIV///////////////////////////////////////////////
    always @(*)
    begin
        if(muxself_en)
            case(muxself)
                2'b00: fdiv_clkin = vcoclk;
                2'b01: fdiv_clkin = vcoclk_dps;
                default: fdiv_clkin = 1'b0;
            endcase
        else
            fdiv_clkin = 1'b0;
    end

    always @(posedge fdiv_clkin or negedge fdiv_clkin or negedge rst_n)
    begin
        if(!rst_n)
        begin
            fdiv_counter <= 8'h0;
            fdiv_out_reg <= 1'b0;
        end
        else
        begin
            if(fdivider == 8'h1)
            begin
                fdiv_counter <= 8'h0;
                fdiv_out_reg <= 1'b0;
            end
            else
            begin
                if(fdiv_counter < ({fdivider, 1'b0} - 1'b1))
                    fdiv_counter <= fdiv_counter + 1'b1;
                else
                    fdiv_counter <= 8'h0;

                if(fdiv_counter < dutyf)
                    fdiv_out_reg <= 1'b1;
                else
                    fdiv_out_reg <= 1'b0;
            end
        end
    end

    assign fdiv_int_out = (fdivider == 8'h1) ? fdiv_clkin : fdiv_out_reg;

    assign fdivider_frac = ratiof_frac;

    always @(*)
    begin
        if(fdiv_frac_en == 1'b1)
        begin
            fdiv_p_int = fdivider / 2;

            if(!fdivider[0])
                if(!fdivider_frac[0])
                begin
                    fdiv_hp_frac = fdivider_frac / 2;
                    fdiv_lp_frac = fdivider_frac / 2;
                end
                else
                begin
                    fdiv_hp_frac = fdivider_frac / 2 + 3'b001;
                    fdiv_lp_frac = fdivider_frac / 2;
                end
            else
                if(!fdivider_frac[0])
                begin
                    fdiv_hp_frac = fdivider_frac / 2 + 3'b100;
                    fdiv_lp_frac = fdivider_frac / 2 + 3'b100;
                end
                else
                begin
                    fdiv_hp_frac = fdivider_frac / 2 + 3'b101;
                    fdiv_lp_frac = fdivider_frac / 2 + 3'b100;
                end
        end
        else
        begin
             fdiv_p_int   = 0;
             fdiv_hp_frac = 0;
             fdiv_lp_frac = 0;
        end
    end

    always @(*)
    begin
        fdiv_frac_hp = vcoclk_period * fdiv_p_int + (vcoclk_period * fdiv_hp_frac) / 8;
        fdiv_frac_lp = vcoclk_period * fdiv_p_int + (vcoclk_period * fdiv_lp_frac) / 8;
    end

    always @(clk_gate or fdiv_frac_out or negedge rst_n)
    begin
        if(!rst_n)
            fdiv_frac_out <= 1'b0;
        else
            if(!clk_gate && fdiv_frac_en && fdiv_dps_en == 1'b0)
            begin
                fdiv_frac_out <= 1'b1;
                for(j = 1; j < 8; j = j+1)
                begin: loop2
                    if(frac_restart)
                    begin
                        #(real_delay);
                        #(fdiv_frac_hp) fdiv_frac_out <= 1'b0;
                        #(fdiv_frac_lp) fdiv_frac_out <= 1'b1;
                    end
                    else
                    begin
                        #(fdiv_frac_hp) fdiv_frac_out <= 1'b0;
                        #(fdiv_frac_lp) fdiv_frac_out <= 1'b1;
                    end
                end
                #(fdiv_frac_hp) fdiv_frac_out <= 1'b0;
                #(fdiv_frac_lp);
                j = 1;
                fdiv_frac_out <= 1'b1;
            end
            else
                fdiv_frac_out <= 1'b0;
    end

    assign fdiv_out = (fdiv_frac_en) ? fdiv_frac_out : fdiv_int_out;
///////////////////////////////////////////////////////
////PHASE_SHIFT////////////////////////////////////////
    always @(*)
    begin
        if(clkout0_time > 0 && odiv0_dps_en == 1'b0)
            vco_fphase_delay0 <= (odiv0_fphase * clkout0_time) / (8 * divider0);
        else
            vco_fphase_delay0 <= 0.0;

        if(clkout1_time > 0 && odiv1_dps_en == 1'b0)
            vco_fphase_delay1 <= (odiv1_fphase * clkout1_time) / (8 * divider1);
        else
            vco_fphase_delay1 <= 0.0;

        if(clkout2_time > 0 && odiv2_dps_en == 1'b0)
            vco_fphase_delay2 <= (odiv2_fphase * clkout2_time) / (8 * divider2);
        else
            vco_fphase_delay2 <= 0.0;

        if(clkout3_time > 0 && odiv3_dps_en == 1'b0)
            vco_fphase_delay3 <= (odiv3_fphase * clkout3_time) / (8 * divider3);
        else
            vco_fphase_delay3 <= 0.0;

        if(clkout4_time > 0 && odiv4_dps_en == 1'b0)
            vco_fphase_delay4 <= (odiv4_fphase * clkout4_time) / (8 * divider4);
        else
            vco_fphase_delay4 <= 0.0;

        if(clkout5_time > 0 && odiv5_dps_en == 1'b0)
            vco_fphase_delay5 <= (odiv5_fphase * clkout5_time) / (8 * divider5);
        else
            vco_fphase_delay5 <= 0.0;

        if(clkout6_time > 0 && odiv6_dps_en == 1'b0)
            vco_fphase_delay6 <= (odiv6_fphase * clkout6_time) / (8 * divider6);
        else
            vco_fphase_delay6 <= 0.0;

        if(clkoutf_time > 0 && fdiv_dps_en == 1'b0)
            vco_fphase_delayf <= (fdiv_fphase * clkoutf_time) / (8 * fdivider);
        else
            vco_fphase_delayf <= 0.0;
    end

    always @(*)
    begin
        if(divider0 > odiv0_cphase)
            cphase0 = odiv0_cphase;
        else
            cphase0 = odiv0_cphase - (odiv0_cphase / divider0) * divider0;

        if(divider1 > odiv1_cphase)
            cphase1 = odiv1_cphase;
        else
            cphase1 = odiv1_cphase - (odiv1_cphase / divider1) * divider1;

        if(divider2 > odiv2_cphase)
            cphase2 = odiv2_cphase;
        else
            cphase2 = odiv2_cphase - (odiv2_cphase / divider2) * divider2;

        if(divider3 > odiv3_cphase)
            cphase3 = odiv3_cphase;
        else
            cphase3 = odiv3_cphase - (odiv3_cphase / divider3) * divider3;

        if(divider4 > odiv4_cphase)
            cphase4 = odiv4_cphase;
        else
            cphase4 = odiv4_cphase - (odiv4_cphase / divider4) * divider4;

        if(divider5 > odiv5_cphase)
            cphase5 = odiv5_cphase;
        else
            cphase5 = odiv5_cphase - (odiv5_cphase / divider5) * divider5;

        if(divider6 > odiv6_cphase)
            cphase6 = odiv6_cphase;
        else
            cphase5 = odiv6_cphase - (odiv6_cphase / divider6) * divider6;

        if(fdivider > fdiv_cphase)
            cphasef = fdiv_cphase;
        else
            cphasef = fdiv_cphase - (fdiv_cphase / fdivider) * fdivider;
    end

    always @(*)
    begin
        if(clkout0_time > 0)
            cphase_delay0 <= clkout0_time - (((divider0 - cphase0) * clkout0_time) / divider0);
        else
            cphase_delay0 <= 0.0;

        if(clkout1_time > 0)
            cphase_delay1 <= clkout1_time - (((divider1 - cphase1) * clkout1_time) / divider1);
        else
            cphase_delay1 <= 0.0;

        if(clkout2_time > 0)
            cphase_delay2 <= clkout2_time - (((divider2 - cphase2) * clkout2_time) / divider2);
        else
            cphase_delay2 <= 0.0;

        if(clkout3_time > 0)
            cphase_delay3 <= clkout3_time - (((divider3 - cphase3) * clkout3_time) / divider3);
        else
            cphase_delay3 <= 0.0;

        if(clkout4_time > 0)
            cphase_delay4 <= clkout4_time - (((divider4 - cphase4) * clkout4_time) / divider4);
        else
            cphase_delay4 <= 0.0;

        if(clkout5_time > 0)
            cphase_delay5 <= clkout5_time - (((divider5 - cphase5) * clkout5_time) / divider5);
        else
            cphase_delay5 <= 0.0;

        if(clkout6_time > 0)
            cphase_delay6 <= clkout6_time - (((divider6 - cphase6) * clkout6_time) / divider6);
        else
            cphase_delay6 <= 0.0;

        if(clkoutf_time > 0)
            cphase_delayf <= clkoutf_time - (((fdivider - cphasef) * clkoutf_time) / fdivider);
        else
            cphase_delayf <= 0.0;
    end
////PHASE_SHIFT_DLY////////////////////////////////////
    always @(odiv0_out or negedge rst_n)
    begin
        if(!rst_n)
            odiv0_out_delay1 <= 1'b0;
        else
            odiv0_out_delay1 <= #vco_fphase_delay0 odiv0_out;
    end

    always @(odiv0_out_delay1 or negedge rst_n)
    begin
        if(!rst_n)
            odiv0_out_delay <= 1'b0;
        else
            odiv0_out_delay <= #cphase_delay0 odiv0_out_delay1;
    end

    always @(odiv1_out or negedge rst_n)
    begin
        if(!rst_n)
            odiv1_out_delay1 <= 1'b0;
        else
            odiv1_out_delay1 <= #vco_fphase_delay1 odiv1_out;
    end

    always @(odiv1_out_delay1 or negedge rst_n)
    begin
        if(!rst_n)
            odiv1_out_delay <= 1'b0;
        else
            odiv1_out_delay <= #cphase_delay1 odiv1_out_delay1;
    end

    always @(odiv2_out or negedge rst_n)
    begin
        if(!rst_n)
            odiv2_out_delay1 <= 1'b0;
        else
            odiv2_out_delay1 <= #vco_fphase_delay2 odiv2_out;
    end

    always @(odiv2_out_delay1 or negedge rst_n)
    begin
        if(!rst_n)
            odiv2_out_delay <= 1'b0;
        else
            odiv2_out_delay <= #cphase_delay2 odiv2_out_delay1;
    end

    always @(odiv3_out or negedge rst_n)
    begin
        if(!rst_n)
            odiv3_out_delay1 <= 1'b0;
        else
            odiv3_out_delay1 <= #vco_fphase_delay3 odiv3_out;
    end

    always @(odiv3_out_delay1 or negedge rst_n)
    begin
        if(!rst_n)
            odiv3_out_delay <= 1'b0;
        else
            odiv3_out_delay <= #cphase_delay3 odiv3_out_delay1;
    end

    always @(odiv4_out or negedge rst_n)
    begin
        if(!rst_n)
            odiv4_out_delay1 <= 1'b0;
        else
            odiv4_out_delay1 <= #vco_fphase_delay4 odiv4_out;
    end

    always @(odiv4_out_delay1 or negedge rst_n)
    begin
        if(!rst_n)
            odiv4_out_delay <= 1'b0;
        else
            odiv4_out_delay <= #cphase_delay4 odiv4_out_delay1;
    end

    always @(odiv5_out or negedge rst_n)
    begin
        if(!rst_n)
            odiv5_out_delay1 <= 1'b0;
        else
            odiv5_out_delay1 <= #vco_fphase_delay5 odiv5_out;
    end

    always @(odiv5_out_delay1 or negedge rst_n)
    begin
        if(!rst_n)
            odiv5_out_delay <= 1'b0;
        else
            odiv5_out_delay <= #cphase_delay5 odiv5_out_delay1;
    end

    always @(odiv6_out or negedge rst_n)
    begin
        if(!rst_n)
            odiv6_out_delay1 <= 1'b0;
        else
            odiv6_out_delay1 <= #vco_fphase_delay6 odiv6_out;
    end

    always @(odiv6_out_delay1 or negedge rst_n)
    begin
        if(!rst_n)
            odiv6_out_delay <= 1'b0;
        else
            odiv6_out_delay <= #cphase_delay6 odiv6_out_delay1;
    end

    always @(fdiv_out or negedge rst_n)
    begin
        if(!rst_n)
            fdiv_out_delay1 <= 1'b0;
        else
            fdiv_out_delay1 <= #vco_fphase_delayf fdiv_out;
    end

    always @(fdiv_out_delay1 or negedge rst_n)
    begin
        if(!rst_n)
            fdiv_out_delay <= 1'b0;
        else
            fdiv_out_delay <= #cphase_delayf fdiv_out_delay1;
    end
///////////////////////////////////////////////////////
////PLL_GATE///////////////////////////////////////////
    assign clkout0_gate = (CLKOUT0_SYN_EN == "TRUE") ? CLKOUT0_SYN : 1'b0;

    always @(negedge odiv0_out_delay or negedge rst_n)
    begin
        if(!rst_n)
            clk_out0_gate <= 3'b000;
        else
            clk_out0_gate <= {clk_out0_gate[1:0], ~clkout0_gate};
    end

    assign CLKOUT0  = odiv0_out_delay & clk_out0_gate[2];
    assign CLKOUT0N = ~CLKOUT0;

    assign clkout1_gate = (CLKOUT1_SYN_EN == "TRUE") ? CLKOUT1_SYN : 1'b0;

    always @(negedge odiv1_out_delay or negedge rst_n)
    begin
        if(!rst_n)
            clk_out1_gate <= 3'b000;
        else
            clk_out1_gate <= {clk_out1_gate[1:0], ~clkout1_gate};
    end

    assign CLKOUT1  = odiv1_out_delay & clk_out1_gate[2];
    assign CLKOUT1N = ~CLKOUT1;

    assign clkout2_gate = (CLKOUT2_SYN_EN == "TRUE") ? CLKOUT2_SYN : 1'b0;

    always @(negedge odiv2_out_delay or negedge rst_n)
    begin
        if(!rst_n)
            clk_out2_gate <= 3'b000;
        else
            clk_out2_gate <= {clk_out2_gate[1:0], ~clkout2_gate};
    end

    assign CLKOUT2  = odiv2_out_delay & clk_out2_gate[2];
    assign CLKOUT2N = ~CLKOUT2;

    assign clkout3_gate = (CLKOUT3_SYN_EN == "TRUE") ? CLKOUT3_SYN : 1'b0;

    always @(negedge odiv3_out_delay or negedge rst_n)
    begin
        if(!rst_n)
            clk_out3_gate <= 3'b000;
        else
            clk_out3_gate <= {clk_out3_gate[1:0], ~clkout3_gate};
    end

    assign CLKOUT3  = odiv3_out_delay & clk_out3_gate[2];
    assign CLKOUT3N = ~CLKOUT3;

    assign clkout4_gate = (CLKOUT4_SYN_EN == "TRUE") ? CLKOUT4_SYN : 1'b0;

    always @(negedge odiv4_out_delay or negedge rst_n)
    begin
        if(!rst_n)
            clk_out4_gate <= 3'b000;
        else
            clk_out4_gate <= {clk_out4_gate[1:0], ~clkout4_gate};
    end

    assign CLKOUT4 = odiv4_out_delay & clk_out4_gate[2];

    assign clkout5_gate = (CLKOUT5_SYN_EN == "TRUE") ? CLKOUT5_SYN : 1'b0;

    always @(negedge odiv5_out_delay or negedge rst_n)
    begin
        if(!rst_n)
            clk_out5_gate <= 3'b000;
        else
            clk_out5_gate <= {clk_out5_gate[1:0], ~clkout5_gate};
    end

    assign CLKOUT5 = odiv5_out_delay & clk_out5_gate[2];

    assign clkout6_gate = (CLKOUT6_SYN_EN == "TRUE") ? CLKOUT6_SYN : 1'b0;

    always @(negedge odiv6_out_delay or negedge rst_n)
    begin
        if(!rst_n)
            clk_out6_gate <= 3'b000;
        else
            clk_out6_gate <= {clk_out6_gate[1:0], ~clkout6_gate};
    end

    assign CLKOUT6 = odiv6_out_delay & clk_out6_gate[2];

    assign clkoutf_gate = (CLKOUTF_SYN_EN == "TRUE") ? CLKOUTF_SYN: 1'b0;

    always @(negedge fdiv_out_delay or negedge rst_n)
    begin
        if(!rst_n)
            clk_outf_gate <= 3'b000;
        else
            clk_outf_gate <= {clk_outf_gate[1:0], ~clkoutf_gate};
    end

    assign CLKOUTF  = fdiv_out_delay & clk_outf_gate[2];
    assign CLKOUTFN = ~CLKOUTF;
///////////////////////////////////////////////////////
////APB////////////////////////////////////////////////
    always @(posedge APB_CLK or negedge APB_RST_N)
    begin
       if(!APB_RST_N)
           apb_rstn_sync <= 2'b00;
       else
           apb_rstn_sync <= {apb_rstn_sync[0], 1'b1};
    end

    always @(posedge APB_CLK or negedge apb_rstn_sync[1])
    begin
        if(!apb_rstn_sync[1])
            ready <= 1'b0;
        else
            if(APB_SEL && !APB_EN)
                ready <= 1'b1;
            else
                ready <= 1'b0;
    end

    always @(posedge APB_CLK)
    begin
        if(APB_WRITE && APB_SEL && APB_EN)
            case(APB_ADDR)
                5'h0 : mem0  <= APB_WDATA;
                5'h1 : mem1  <= APB_WDATA;
                5'h2 : mem2  <= APB_WDATA[5:0];
                5'h3 : mem3  <= APB_WDATA;
                5'h4 : mem4  <= APB_WDATA[12:0];
                5'h5 : mem5  <= APB_WDATA;
                5'h6 : mem6  <= APB_WDATA[12:0];
                5'h7 : mem7  <= APB_WDATA;
                5'h8 : mem8  <= APB_WDATA[12:0];
                5'h9 : mem9  <= APB_WDATA;
                5'hA : mem10 <= APB_WDATA[12:0];
                5'hB : mem11 <= APB_WDATA;
                5'hC : mem12 <= APB_WDATA[12:0];
                5'hD : mem13 <= APB_WDATA;
                5'hE : mem14 <= APB_WDATA[12:0];
                5'hF : mem15 <= APB_WDATA;
                5'h10: mem16 <= APB_WDATA;
                5'h11: mem17 <= APB_WDATA[5:0];
                5'h12: mem18 <= APB_WDATA[7:0];
                5'h13: mem19 <= APB_WDATA[7:0];
                5'h14: mem20 <= APB_WDATA[13:0];
                5'h15: mem21 <= APB_WDATA[5:0];
            endcase
    end

    always @(posedge APB_CLK or negedge apb_rstn_sync[1])
    begin
        if(!apb_rstn_sync[1])
            rdata <= 16'h0;
        else
            if(!APB_WRITE && APB_SEL && !APB_EN)
                case(APB_ADDR)
                    5'h0 : rdata <= mem0;
                    5'h1 : rdata <= mem1;
                    5'h2 : rdata <= mem2;
                    5'h3 : rdata <= mem3;
                    5'h4 : rdata <= mem4;
                    5'h5 : rdata <= mem5;
                    5'h6 : rdata <= mem6;
                    5'h7 : rdata <= mem7;
                    5'h8 : rdata <= mem8;
                    5'h9 : rdata <= mem9;
                    5'hA : rdata <= mem10;
                    5'hB : rdata <= mem11;
                    5'hC : rdata <= mem12;
                    5'hD : rdata <= mem13;
                    5'hE : rdata <= mem14;
                    5'hF : rdata <= mem15;
                    5'h10: rdata <= mem16;
                    5'h11: rdata <= mem17;
                    5'h12: rdata <= mem18;
                    5'h13: rdata <= mem19;
                    5'h14: rdata <= mem20;
                    5'h15: rdata <= mem21;
                endcase
            else
                rdata <= 16'h0;
    end

    assign APB_READY = ready;
    assign APB_RDATA = rdata;
endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_ZERO.v
//
// Functional description: constant zero
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_ZERO
(
    output wire Z
);

    supply0 VSS;
    buf (Z, VSS);

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_PREADD_MULTADD18.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

//P = A0*(B0+-C0) +/- A1*(B1+-C1)
`timescale 1 ns / 1 ps

module GTP_PREADD_MULTADD18 #(
    parameter GRS_EN            = "TRUE", //"TRUE"; "FALSE"
    parameter SYNC_RST          = "FALSE", //"TRUE"; "FALSE"  
    parameter INREG_EN          = "FALSE", //"TRUE"; "FALSE"
    parameter PREREG_EN         = "FALSE", //"TRUE"; "FALSE"
    parameter PIPEREG_EN        = "FALSE", //"TRUE"; "FALSE"
    parameter OUTREG_EN         = "FALSE", //"TRUE"; "FALSE"
    parameter ADDSUB_OP         = 0,
    parameter DYN_ADDSUB_OP     = 1
)(
    output  [38-1:0] P,
    input   CE,
    input   RST,
    input   CLK,
    input   [18-1:0] A0,
    input   [18-1:0] A1,
    input   [18-1:0] B0,
    input   [18-1:0] B1,
    input   [18-1:0] C0,
    input   [18-1:0] C1,
    input   A_SIGNED,
    input   B_SIGNED,
    input   C_SIGNED,
    input   [1:0] PREADDSUB,
    input   ADDSUB
);


    INT_PREADD_MULTADD #(
        . GRS_EN(GRS_EN),    
        . SYNC_RST(SYNC_RST),  
        . INREG_EN(INREG_EN), 
        . PREREG_EN(PREREG_EN), 
        . PIPEREG_EN(PIPEREG_EN),
        . OUTREG_EN(OUTREG_EN), 
        . ADDSUB_OP(ADDSUB_OP),   
        . DYN_OP_ADDSUB(DYN_ADDSUB_OP),
        . ASIZE(18), 
        . BSIZE(18)
    ) U_INT_PREADD_MULTADD(
        . CE(CE),
        . RST(RST),
        . CLK(CLK),
        . A0(A0),
        . A1(A1),
        . B0(B0),
        . B1(B1),
        . C0(C0),
        . C1(C1),
        . A_SIGNED(A_SIGNED),
        . B_SIGNED(B_SIGNED),
        . C_SIGNED(C_SIGNED),
        . PREADDSUB(PREADDSUB),
        . ADDSUB(ADDSUB),
        . P(P)
    );   


endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
//  REVISION:
//  10/10/15   - Initial version
//  10/13/15   - Change sram bits of "other" blocks parameter type from integer to string
//             - Remove ports "P_DATA/N", "P_VSSM/P_VCCM", "P_ADDR_T/B"                     
//  10/22/15   - Based on 10-14 Schematic
//             - Parameter newly refreshed
//             - New PMA model of 10-14
//  10/29/15   - Based on 10-14 Schematic
//             - Parameter newly refreshed
//             - Removed Power related IOs
//             - Removed Bscan related IOs
//             - Removed DFT related IOs
//  11/04/15   - Correct "db" to upper case "DB"
//             - Corresponding wrap file updated of rule process
//  12/04/15   - Add one missing parameter for 4 channels 
//             - PCS_CH0_PCIE_SLAVE
//             - PCS_CH1_PCIE_SLAVE
//             - PCS_CH2_PCIE_SLAVE
//             - PCS_CH3_PCIE_SLAVE
//  12/10/15   - Removed "TAB" space 
//  01/14/16   - BASE-ED ON PMA VENDOR V1.4 register table 
//             - add one parameter "PMA_QUAD_LF_TEST_EN" on txpll[3] 
//             - add one parameter "PMA_QUAD_LF_TESTBY2" on txpll[10] 
//             - correct name on txpll[0] 
//             - correct name on txpll[1] 
//             - correct name on refclk[1] 
//             - correct name on refclk[17:18] 
//  03/18/16   - Optimize the parameter's value adjustment
//             - As, PMA_CH[0-3]_CDR_TEST_OUT_SELECT:  value "FB_CK"2"FBCK" 
//             - As, PMA_CH1_EQ1_CURRENT_SETTING: value "1111"2"15"  
//             - As, PMA_QUAD_FREQ_LKO/I: value "100PCT"2"10PCT" 

 

`timescale 1ns/100fs

module GTP_HSST 

#(
// PARAMETER  PART BEGINS ////////////////////////////////////////////////////////////////////
// PARAMETER  PART BEGINS ////////////////////////////////////////////////////////////////////
// PARAMETER  PART BEGINS ////////////////////////////////////////////////////////////////////



parameter        PCS_CH0_BYPASS_WORD_ALIGN    = "FALSE",        // FALSE,TRUE
parameter           PCS_CH0_BYPASS_DENC    = "FALSE",        // FALSE,TRUE
parameter           PCS_CH0_BYPASS_BONDING    = "FALSE",        // FALSE,TRUE
parameter           PCS_CH0_BYPASS_CTC    = "FALSE",        // FALSE,TRUE
parameter           PCS_CH0_BYPASS_GEAR    = "FALSE",        // FALSE,TRUE
parameter           PCS_CH0_BYPASS_BRIDGE    = "FALSE",        // FALSE,TRUE
parameter           PCS_CH0_DATA_MODE    = "X8",        // 8bit,10bit,16bit,20bit
parameter           PCS_CH0_RX_POLARITY_INV    = "DELAY",        // 00: delay 01: bit polarity inversion 10: bit reversal 11: polarity inversion and bit reversal
parameter           PCS_CH0_ALIGN_MODE    = "1GB",        // 1GB,10GB,RAPIDIO,OUTSIDE
parameter           PCS_CH0_SAMP_16B = "X16",        // 16bit,20bit
parameter   integer PCS_CH0_COMMA_REG0 = 0,        // 
parameter   integer PCS_CH0_COMMA_MASK = 0,        // 
parameter        PCS_CH0_CEB_MODE = "10GB",        // 10GB,RAPIDIO,OUTSIDE
parameter           PCS_CH0_CTC_MODE = "1SKIP",        // 00: add or del 1 skip,01: add or del 2 skips,10: reserved ,11:4 skips
parameter   integer PCS_CH0_A_REG = 0,        // 
parameter        PCS_CH0_GE_AUTO_EN = "FALSE",        // CTC,FALSE,TRUE
parameter   integer PCS_CH0_SKIP_REG0 = 0,        // 
parameter   integer PCS_CH0_SKIP_REG1 = 0,        // 
parameter   integer PCS_CH0_SKIP_REG2 = 0,        // 
parameter   integer PCS_CH0_SKIP_REG3 = 0,        // 
parameter        PCS_CH0_DEC_DUAL = "FALSE",        // signal for 8b10b decoder module
parameter           PCS_CH0_SPLIT = "FALSE",        // signal for RX GEAR split, 1:split  0:no split, 
parameter           PCS_CH0_FIFOFLAG_CTC = "FALSE",        // FALSE,TRUE
parameter           PCS_CH0_COMMA_DET_MODE = "COMMA_PATTERN",        // 0: comma pattern mode  1: RX_CLK_SLIP mode 
parameter           PCS_CH0_ERRDETECT_SILENCE = "FALSE",        // 0: comma pattern mode  1: RX_CLK_SLIP mode 
parameter           PCS_CH0_PMA_RCLK_POLINV = "PMA_RCLK",        // 1'b0:pma_rclk 1'b1:reverse of pma_rclk
parameter           PCS_CH0_PCS_RCLK_SEL = "PMA_RCLK",        // 1'b0:pma_rclk,1'b1:pma_tclk,
parameter           PCS_CH0_MCB_RCLK_POLINV = "MCB_RCLK",        // 1'b0:mcb_rclk 1'b1:reverse of mcb_rclk
parameter        PCS_CH0_CB_RCLK_SEL = "PMA_RCLK",        // 2'b00:pma_rclk,2'b01:pma_tclk,2'b10:mcb_rclk,2'b11:reserved
parameter           PCS_CH0_AFTER_CTC_RCLK_SEL = "PMA_RCLK",        // 2'b00:pma_rclk,2'b01:pma_tclk,2'b10:mcb_rclk,2'b11:reserved
parameter           PCS_CH0_RCLK_POLINV = "RCLK",        // 1'b0:rclk 1'b1:reverse of rclk
parameter           PCS_CH0_BRIDGE_RCLK_SEL = "PMA_RCLK",        // 2'b00:pma_rclk,2'b01:pma_tclk,2'b10:mcb_rclk,2'b11:rclk
parameter           PCS_CH0_PCS_RCLK_EN = "FALSE",        // FALSE,TRUE
parameter           PCS_CH0_CB_RCLK_EN = "FALSE",        // FALSE,TRUE
parameter           PCS_CH0_AFTER_CTC_RCLK_EN = "FALSE",        // FALSE,TRUE
parameter           PCS_CH0_AFTER_CTC_RCLK_EN_GB = "FALSE",        // FALSE,TRUE
parameter           PCS_CH0_BRIDGE_RCLK_EN = "FALSE",        // FALSE,TRUE
parameter           PCS_CH0_PCS_RX_RSTN = "FALSE",        // 1:pcs_rx_rstn is valued,is 0,0:pcs_rx_rstn is released
parameter           PCS_CH0_SLAVE = "MASTER",        // 1:slave channel 0:master channel
parameter           PCS_CH0_PCIE_SLAVE = "MASTER",        // 1:slave channel 0:master channel
parameter           PCS_CH0_PCS_CB_RSTN = "FALSE",        // 1: pcs_cb_rstn is valued,is 0,0: pcs_cb_rstn is released
parameter           PCS_CH0_TX_BYPASS_BRIDGE_UINT    = "FALSE",        // FALSE,TRUE
parameter           PCS_CH0_TX_BYPASS_GEAR    = "FALSE",        // FALSE,TRUE
parameter           PCS_CH0_TX_BYPASS_ENC    = "FALSE",        // FALSE,TRUE
parameter           PCS_CH0_TX_BYPASS_BIT_SLIP    = "FALSE",        // FALSE,TRUE
parameter           PCS_CH0_TX_GEAR_SPLIT    = "FALSE",        // 1:spilt 44bits data to 22bits data,0: no spilt
parameter        PCS_CH0_TX_DRIVE_REG_MODE    = "NO_CHANGE",        // 00:no change, 01:enable polarity reverse,10:enable bit reverse, 11:enable both
parameter   integer PCS_CH0_TX_BIT_SLIP_CYCLES = 0,        // 
parameter        PCS_CH0_INT_TX_MASK_0 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by tx_bridge_unit async fifo overflow
parameter              PCS_CH0_INT_TX_MASK_1 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by tx bridge unit underflow,
parameter              PCS_CH0_INT_TX_MASK_2 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by tx_invalid_k 
parameter              PCS_CH0_INT_TX_CLR_0 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by tx bridge unit overflow,
parameter              PCS_CH0_INT_TX_CLR_1 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by tx_bridge_unit async fifo underflow
parameter              PCS_CH0_INT_TX_CLR_2 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by tx_invalid_k
parameter        PCS_CH0_TX_PMA_TCLK_POLINV = "PMA_TCLK",        // 1'b0:pma_tclk 1'b1:reverse of pma_tclk
parameter        PCS_CH0_TX_PCS_CLK_EN_SEL = "FALSE",        // FALSE,TRUE
parameter        PCS_CH0_TX_BRIDGE_TCLK_SEL = "PCS_TCLK",        // 1'b0: pcs_tclk 1'b1:tclk
parameter        PCS_CH0_TX_TCLK_POLINV = "TCLK",        // 1'b0:tclk 1'b1:reverse of tclk
parameter        PCS_CH0_TX_PCS_TX_RSTN = "FALSE",        // 1:pcs_tx_rstn is valued,is 0,0:pcs_tx_rstn is released
parameter        PCS_CH0_TX_SLAVE = "SLAVE",        // 1:slave channel,0:master channel
parameter        PCS_CH0_TX_BRIDGE_CLK_EN_SEL = "FALSE",        // FALSE,TRUE
parameter        PCS_CH0_DATA_WIDTH_MODE    = "X20",        // 20bit,16bit,10bit,8bit
parameter        PCS_CH0_TX_TCLK2FABRIC_SEL = "FALSE",        // FALSE,TRUE
parameter        PCS_CH0_TX_OUTZZ = "FALSE",        // 1:16bit/32bit only,0:20bit/40bit only
parameter        PCS_CH0_ENC_DUAL = "FALSE",        // FALSE,TRUE
parameter        PCS_CH0_TX_BITSLIP_DATA_MODE = "X10",        // 1: 20bit,0: 10bit
parameter   integer PCS_CH0_COMMA_REG1 = 0,        // 
parameter   integer PCS_CH0_RAPID_IMAX = 0,        // 
parameter   integer PCS_CH0_RAPID_VMIN_1 = 0,        // 
parameter   integer PCS_CH0_RAPID_VMIN_2 = 0,        // 
parameter        PCS_CH0_RX_PRBS_MODE = "DISABLE",        // Mode select:4'd0: reserved,4'd1: PRBS-7,4'd2: PRBS-15,4'd3: PRBS-23,4'd4: PRBS-31,4'd5: long "1",4'd6: long "0",4'd7: 20UI square wave,4'd8: D10_2,4'd9: PCIe complianece pattern,Others: reserved
parameter        PCS_CH0_RX_ERRCNT_CLR = "FALSE",        // FALSE,TRUE
parameter        PCS_CH0_TX_PRBS_MODE = "DISABLE",        // Mode select:4'd0: reserved,4'd1: PRBS-7,4'd2: PRBS-15,4'd3: PRBS-23,4'd4: PRBS-31,4'd5: long "1",4'd6: long "0",4'd7: 20UI square wave,4'd8: D10_2,4'd9: PCIe complianece pattern,Others: reserved
parameter        PCS_CH0_TX_INSERT_ER = "FALSE",        // FALSE,TRUE
parameter        PCS_CH0_ENABLE_PRBS_GEN = "FALSE",        // FALSE,TRUE
parameter   integer PCS_CH0_ERR_CNT = 0,        // 
parameter   integer PCS_CH0_DEFAULT_RADDR = 0,        // 
parameter   integer PCS_CH0_MASTER_CHECK_OFFSET = 0,        // 
parameter   integer PCS_CH0_DELAY_SET = 0,        // 
parameter        PCS_CH0_SEACH_OFFSET = "20BIT",        // 20bit,30bit,40bit,50bit,60bit,70bit
parameter   integer PCS_CH0_CEB_RAPIDLS_MMAX = 0,        // 
parameter   integer PCS_CH0_CTC_AFULL = 0,        // 
parameter   integer PCS_CH0_CTC_AEMPTY = 0,        // 
parameter        PCS_CH0_FAR_LOOP = "FALSE",        // FALSE,TRUE
parameter              PCS_CH0_NEAR_LOOP = "FALSE",        // FALSE,TRUE
parameter              PCS_CH0_INT_RX_MASK_0 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by pcs_lsm_synced
parameter              PCS_CH0_INT_RX_MASK_1 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by pcs_rx_mcb_status
parameter              PCS_CH0_INT_RX_MASK_2 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by channel bonding async fifo overflow
parameter              PCS_CH0_INT_RX_MASK_3 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by channel bonding async fifo underflow
parameter              PCS_CH0_INT_RX_MASK_4 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by ctc unit async fifo overflow
parameter              PCS_CH0_INT_RX_MASK_5 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by ctc unit async fifo underflow
parameter              PCS_CH0_INT_RX_MASK_6 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by rx_bridge_unit async fifo overflow
parameter              PCS_CH0_INT_RX_MASK_7 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by rx_bridge_unit async fifo underflow
parameter              PCS_CH0_INT_RX_CLR_0 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by pcs_lsm_synced
parameter              PCS_CH0_INT_RX_CLR_1 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by pcs_rx_mcb_status
parameter              PCS_CH0_INT_RX_CLR_2 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by channel bonding async fifo overflow
parameter              PCS_CH0_INT_RX_CLR_3 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by channel bonding async fifo underflow
parameter              PCS_CH0_INT_RX_CLR_4 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by ctc unit async fifo overflow
parameter              PCS_CH0_INT_RX_CLR_5 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by ctc unit async fifo underflow
parameter              PCS_CH0_INT_RX_CLR_6 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by rx_bridge_unit async fifo overflow
parameter              PCS_CH0_INT_RX_CLR_7 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by rx_bridge_unit async fifo underflow



parameter        PCS_CH1_BYPASS_WORD_ALIGN    = "FALSE",        // FALSE,TRUE
parameter           PCS_CH1_BYPASS_DENC    = "FALSE",        // FALSE,TRUE
parameter           PCS_CH1_BYPASS_BONDING    = "FALSE",        // FALSE,TRUE
parameter           PCS_CH1_BYPASS_CTC    = "FALSE",        // FALSE,TRUE
parameter           PCS_CH1_BYPASS_GEAR    = "FALSE",        // FALSE,TRUE
parameter           PCS_CH1_BYPASS_BRIDGE    = "FALSE",        // FALSE,TRUE
parameter           PCS_CH1_DATA_MODE    = "X8",        // 8bit,10bit,16bit,20bit
parameter           PCS_CH1_RX_POLARITY_INV    = "DELAY",        // 00: delay 01: bit polarity inversion 10: bit reversal 11: polarity inversion and bit reversal
parameter           PCS_CH1_ALIGN_MODE    = "1GB",        // 1GB,10GB,RAPIDIO,OUTSIDE
parameter           PCS_CH1_SAMP_16B = "X16",        // 16bit,20bit
parameter   integer PCS_CH1_COMMA_REG0 = 0,        // 
parameter   integer PCS_CH1_COMMA_MASK = 0,        // 
parameter        PCS_CH1_CEB_MODE = "10GB",        // 10GB,RAPIDIO,OUTSIDE
parameter           PCS_CH1_CTC_MODE = "1SKIP",        // 00: add or del 1 skip,01: add or del 2 skips,10: reserved ,11:4 skips
parameter   integer PCS_CH1_A_REG = 0,        // 
parameter        PCS_CH1_GE_AUTO_EN = "FALSE",        // CTC,FALSE,TRUE
parameter   integer PCS_CH1_SKIP_REG0 = 0,        // 
parameter   integer PCS_CH1_SKIP_REG1 = 0,        // 
parameter   integer PCS_CH1_SKIP_REG2 = 0,        // 
parameter   integer PCS_CH1_SKIP_REG3 = 0,        // 
parameter        PCS_CH1_DEC_DUAL = "FALSE",        // signal for 8b10b decoder module
parameter           PCS_CH1_SPLIT = "FALSE",        // signal for RX GEAR split, 1:split  0:no split, 
parameter           PCS_CH1_FIFOFLAG_CTC = "FALSE",        // FALSE,TRUE
parameter           PCS_CH1_COMMA_DET_MODE = "COMMA_PATTERN",        // 0: comma pattern mode  1: RX_CLK_SLIP mode 
parameter           PCS_CH1_ERRDETECT_SILENCE = "FALSE",        // 0: comma pattern mode  1: RX_CLK_SLIP mode 
parameter           PCS_CH1_PMA_RCLK_POLINV = "PMA_RCLK",        // 1'b0:pma_rclk 1'b1:reverse of pma_rclk
parameter           PCS_CH1_PCS_RCLK_SEL = "PMA_RCLK",        // 1'b0:pma_rclk,1'b1:pma_tclk,
parameter           PCS_CH1_MCB_RCLK_POLINV = "MCB_RCLK",        // 1'b0:mcb_rclk 1'b1:reverse of mcb_rclk
parameter        PCS_CH1_CB_RCLK_SEL = "PMA_RCLK",        // 2'b00:pma_rclk,2'b01:pma_tclk,2'b10:mcb_rclk,2'b11:reserved
parameter           PCS_CH1_AFTER_CTC_RCLK_SEL = "PMA_RCLK",        // 2'b00:pma_rclk,2'b01:pma_tclk,2'b10:mcb_rclk,2'b11:reserved
parameter           PCS_CH1_RCLK_POLINV = "RCLK",        // 1'b0:rclk 1'b1:reverse of rclk
parameter           PCS_CH1_BRIDGE_RCLK_SEL = "PMA_RCLK",        // 2'b00:pma_rclk,2'b01:pma_tclk,2'b10:mcb_rclk,2'b11:rclk
parameter           PCS_CH1_PCS_RCLK_EN = "FALSE",        // FALSE,TRUE
parameter           PCS_CH1_CB_RCLK_EN = "FALSE",        // FALSE,TRUE
parameter           PCS_CH1_AFTER_CTC_RCLK_EN = "FALSE",        // FALSE,TRUE
parameter           PCS_CH1_AFTER_CTC_RCLK_EN_GB = "FALSE",        // FALSE,TRUE
parameter           PCS_CH1_BRIDGE_RCLK_EN = "FALSE",        // FALSE,TRUE
parameter           PCS_CH1_PCS_RX_RSTN = "FALSE",        // 1:pcs_rx_rstn is valued,is 0,0:pcs_rx_rstn is released
parameter           PCS_CH1_SLAVE = "MASTER",        // 1:slave channel 0:master channel
parameter           PCS_CH1_PCIE_SLAVE = "MASTER",        // 1:slave channel 0:master channel
parameter           PCS_CH1_PCS_CB_RSTN = "FALSE",        // 1: pcs_cb_rstn is valued,is 0,0: pcs_cb_rstn is released
parameter           PCS_CH1_TX_BYPASS_BRIDGE_UINT    = "FALSE",        // FALSE,TRUE
parameter           PCS_CH1_TX_BYPASS_GEAR    = "FALSE",        // FALSE,TRUE
parameter           PCS_CH1_TX_BYPASS_ENC    = "FALSE",        // FALSE,TRUE
parameter           PCS_CH1_TX_BYPASS_BIT_SLIP    = "FALSE",        // FALSE,TRUE
parameter           PCS_CH1_TX_GEAR_SPLIT    = "FALSE",        // 1:spilt 44bits data to 22bits data,0: no spilt
parameter        PCS_CH1_TX_DRIVE_REG_MODE    = "NO_CHANGE",        // 00:no change, 01:enable polarity reverse,10:enable bit reverse, 11:enable both
parameter   integer PCS_CH1_TX_BIT_SLIP_CYCLES = 0,        // 
parameter        PCS_CH1_INT_TX_MASK_0 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by tx_bridge_unit async fifo overflow
parameter              PCS_CH1_INT_TX_MASK_1 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by tx bridge unit underflow,
parameter              PCS_CH1_INT_TX_MASK_2 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by tx_invalid_k 
parameter              PCS_CH1_INT_TX_CLR_0 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by tx bridge unit overflow,
parameter              PCS_CH1_INT_TX_CLR_1 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by tx_bridge_unit async fifo underflow
parameter              PCS_CH1_INT_TX_CLR_2 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by tx_invalid_k
parameter        PCS_CH1_TX_PMA_TCLK_POLINV = "PMA_TCLK",        // 1'b0:pma_tclk 1'b1:reverse of pma_tclk
parameter        PCS_CH1_TX_PCS_CLK_EN_SEL = "FALSE",        // FALSE,TRUE
parameter        PCS_CH1_TX_BRIDGE_TCLK_SEL = "PCS_TCLK",        // 1'b0: pcs_tclk 1'b1:tclk
parameter        PCS_CH1_TX_TCLK_POLINV = "TCLK",        // 1'b0:tclk 1'b1:reverse of tclk
parameter        PCS_CH1_TX_PCS_TX_RSTN = "FALSE",        // 1:pcs_tx_rstn is valued,is 0,0:pcs_tx_rstn is released
parameter        PCS_CH1_TX_SLAVE = "SLAVE",        // 1:slave channel,0:master channel
parameter        PCS_CH1_TX_BRIDGE_CLK_EN_SEL = "FALSE",        // FALSE,TRUE
parameter        PCS_CH1_DATA_WIDTH_MODE    = "X20",        // 20bit,16bit,10bit,8bit
parameter        PCS_CH1_TX_TCLK2FABRIC_SEL = "FALSE",        // FALSE,TRUE
parameter        PCS_CH1_TX_OUTZZ = "FALSE",        // 1:16bit/32bit only,0:20bit/40bit only
parameter        PCS_CH1_ENC_DUAL = "FALSE",        // FALSE,TRUE
parameter        PCS_CH1_TX_BITSLIP_DATA_MODE = "X10",        // 1: 20bit,0: 10bit
parameter   integer PCS_CH1_COMMA_REG1 = 0,        // 
parameter   integer PCS_CH1_RAPID_IMAX = 0,        // 
parameter   integer PCS_CH1_RAPID_VMIN_1 = 0,        // 
parameter   integer PCS_CH1_RAPID_VMIN_2 = 0,        // 
parameter        PCS_CH1_RX_PRBS_MODE = "DISABLE",        // Mode select:4'd0: reserved,4'd1: PRBS-7,4'd2: PRBS-15,4'd3: PRBS-23,4'd4: PRBS-31,4'd5: long "1",4'd6: long "0",4'd7: 20UI square wave,4'd8: D10_2,4'd9: PCIe complianece pattern,Others: reserved
parameter        PCS_CH1_RX_ERRCNT_CLR = "FALSE",        // FALSE,TRUE
parameter        PCS_CH1_TX_PRBS_MODE = "DISABLE",        // Mode select:4'd0: reserved,4'd1: PRBS-7,4'd2: PRBS-15,4'd3: PRBS-23,4'd4: PRBS-31,4'd5: long "1",4'd6: long "0",4'd7: 20UI square wave,4'd8: D10_2,4'd9: PCIe complianece pattern,Others: reserved
parameter        PCS_CH1_TX_INSERT_ER = "FALSE",        // FALSE,TRUE
parameter        PCS_CH1_ENABLE_PRBS_GEN = "FALSE",        // FALSE,TRUE
parameter   integer PCS_CH1_ERR_CNT = 0,        // 
parameter   integer PCS_CH1_DEFAULT_RADDR = 0,        // 
parameter   integer PCS_CH1_MASTER_CHECK_OFFSET = 0,        // 
parameter   integer PCS_CH1_DELAY_SET = 0,        // 
parameter        PCS_CH1_SEACH_OFFSET = "20BIT",        // 20bit,30bit,40bit,50bit,60bit,70bit
parameter   integer PCS_CH1_CEB_RAPIDLS_MMAX = 0,        // 
parameter   integer PCS_CH1_CTC_AFULL = 0,        // 
parameter   integer PCS_CH1_CTC_AEMPTY = 0,        // 
parameter        PCS_CH1_FAR_LOOP = "FALSE",        // FALSE,TRUE
parameter              PCS_CH1_NEAR_LOOP = "FALSE",        // FALSE,TRUE
parameter              PCS_CH1_INT_RX_MASK_0 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by pcs_lsm_synced
parameter              PCS_CH1_INT_RX_MASK_1 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by pcs_rx_mcb_status
parameter              PCS_CH1_INT_RX_MASK_2 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by channel bonding async fifo overflow
parameter              PCS_CH1_INT_RX_MASK_3 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by channel bonding async fifo underflow
parameter              PCS_CH1_INT_RX_MASK_4 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by ctc unit async fifo overflow
parameter              PCS_CH1_INT_RX_MASK_5 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by ctc unit async fifo underflow
parameter              PCS_CH1_INT_RX_MASK_6 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by rx_bridge_unit async fifo overflow
parameter              PCS_CH1_INT_RX_MASK_7 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by rx_bridge_unit async fifo underflow
parameter              PCS_CH1_INT_RX_CLR_0 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by pcs_lsm_synced
parameter              PCS_CH1_INT_RX_CLR_1 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by pcs_rx_mcb_status
parameter              PCS_CH1_INT_RX_CLR_2 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by channel bonding async fifo overflow
parameter              PCS_CH1_INT_RX_CLR_3 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by channel bonding async fifo underflow
parameter              PCS_CH1_INT_RX_CLR_4 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by ctc unit async fifo overflow
parameter              PCS_CH1_INT_RX_CLR_5 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by ctc unit async fifo underflow
parameter              PCS_CH1_INT_RX_CLR_6 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by rx_bridge_unit async fifo overflow
parameter              PCS_CH1_INT_RX_CLR_7 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by rx_bridge_unit async fifo underflow



parameter        PCS_CH2_BYPASS_WORD_ALIGN    = "FALSE",        // FALSE,TRUE
parameter           PCS_CH2_BYPASS_DENC    = "FALSE",        // FALSE,TRUE
parameter           PCS_CH2_BYPASS_BONDING    = "FALSE",        // FALSE,TRUE
parameter           PCS_CH2_BYPASS_CTC    = "FALSE",        // FALSE,TRUE
parameter           PCS_CH2_BYPASS_GEAR    = "FALSE",        // FALSE,TRUE
parameter           PCS_CH2_BYPASS_BRIDGE    = "FALSE",        // FALSE,TRUE
parameter           PCS_CH2_DATA_MODE    = "X8",        // 8bit,10bit,16bit,20bit
parameter           PCS_CH2_RX_POLARITY_INV    = "DELAY",        // 00: delay 01: bit polarity inversion 10: bit reversal 11: polarity inversion and bit reversal
parameter           PCS_CH2_ALIGN_MODE    = "1GB",        // 1GB,10GB,RAPIDIO,OUTSIDE
parameter           PCS_CH2_SAMP_16B = "X16",        // 16bit,20bit
parameter   integer PCS_CH2_COMMA_REG0 = 0,        // 
parameter   integer PCS_CH2_COMMA_MASK = 0,        // 
parameter        PCS_CH2_CEB_MODE = "10GB",        // 10GB,RAPIDIO,OUTSIDE
parameter           PCS_CH2_CTC_MODE = "1SKIP",        // 00: add or del 1 skip,01: add or del 2 skips,10: reserved ,11:4 skips
parameter   integer PCS_CH2_A_REG = 0,        // 
parameter        PCS_CH2_GE_AUTO_EN = "FALSE",        // CTC,FALSE,TRUE
parameter   integer PCS_CH2_SKIP_REG0 = 0,        // 
parameter   integer PCS_CH2_SKIP_REG1 = 0,        // 
parameter   integer PCS_CH2_SKIP_REG2 = 0,        // 
parameter   integer PCS_CH2_SKIP_REG3 = 0,        // 
parameter        PCS_CH2_DEC_DUAL = "FALSE",        // signal for 8b10b decoder module
parameter           PCS_CH2_SPLIT = "FALSE",        // signal for RX GEAR split, 1:split  0:no split, 
parameter           PCS_CH2_FIFOFLAG_CTC = "FALSE",        // FALSE,TRUE
parameter           PCS_CH2_COMMA_DET_MODE = "COMMA_PATTERN",        // 0: comma pattern mode  1: RX_CLK_SLIP mode 
parameter           PCS_CH2_ERRDETECT_SILENCE = "FALSE",        // 0: comma pattern mode  1: RX_CLK_SLIP mode 
parameter           PCS_CH2_PMA_RCLK_POLINV = "PMA_RCLK",        // 1'b0:pma_rclk 1'b1:reverse of pma_rclk
parameter           PCS_CH2_PCS_RCLK_SEL = "PMA_RCLK",        // 1'b0:pma_rclk,1'b1:pma_tclk,
parameter           PCS_CH2_MCB_RCLK_POLINV = "MCB_RCLK",        // 1'b0:mcb_rclk 1'b1:reverse of mcb_rclk
parameter        PCS_CH2_CB_RCLK_SEL = "PMA_RCLK",        // 2'b00:pma_rclk,2'b01:pma_tclk,2'b10:mcb_rclk,2'b11:reserved
parameter           PCS_CH2_AFTER_CTC_RCLK_SEL = "PMA_RCLK",        // 2'b00:pma_rclk,2'b01:pma_tclk,2'b10:mcb_rclk,2'b11:reserved
parameter           PCS_CH2_RCLK_POLINV = "RCLK",        // 1'b0:rclk 1'b1:reverse of rclk
parameter           PCS_CH2_BRIDGE_RCLK_SEL = "PMA_RCLK",        // 2'b00:pma_rclk,2'b01:pma_tclk,2'b10:mcb_rclk,2'b11:rclk
parameter           PCS_CH2_PCS_RCLK_EN = "FALSE",        // FALSE,TRUE
parameter           PCS_CH2_CB_RCLK_EN = "FALSE",        // FALSE,TRUE
parameter           PCS_CH2_AFTER_CTC_RCLK_EN = "FALSE",        // FALSE,TRUE
parameter           PCS_CH2_AFTER_CTC_RCLK_EN_GB = "FALSE",        // FALSE,TRUE
parameter           PCS_CH2_BRIDGE_RCLK_EN = "FALSE",        // FALSE,TRUE
parameter           PCS_CH2_PCS_RX_RSTN = "FALSE",        // 1:pcs_rx_rstn is valued,is 0,0:pcs_rx_rstn is released
parameter           PCS_CH2_SLAVE = "MASTER",        // 1:slave channel 0:master channel
parameter           PCS_CH2_PCIE_SLAVE = "MASTER",        // 1:slave channel 0:master channel
parameter           PCS_CH2_PCS_CB_RSTN = "FALSE",        // 1: pcs_cb_rstn is valued,is 0,0: pcs_cb_rstn is released
parameter           PCS_CH2_TX_BYPASS_BRIDGE_UINT    = "FALSE",        // FALSE,TRUE
parameter           PCS_CH2_TX_BYPASS_GEAR    = "FALSE",        // FALSE,TRUE
parameter           PCS_CH2_TX_BYPASS_ENC    = "FALSE",        // FALSE,TRUE
parameter           PCS_CH2_TX_BYPASS_BIT_SLIP    = "FALSE",        // FALSE,TRUE
parameter           PCS_CH2_TX_GEAR_SPLIT    = "FALSE",        // 1:spilt 44bits data to 22bits data,0: no spilt
parameter        PCS_CH2_TX_DRIVE_REG_MODE    = "NO_CHANGE",        // 00:no change, 01:enable polarity reverse,10:enable bit reverse, 11:enable both
parameter   integer PCS_CH2_TX_BIT_SLIP_CYCLES = 0,        // 
parameter        PCS_CH2_INT_TX_MASK_0 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by tx_bridge_unit async fifo overflow
parameter              PCS_CH2_INT_TX_MASK_1 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by tx bridge unit underflow,
parameter              PCS_CH2_INT_TX_MASK_2 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by tx_invalid_k 
parameter              PCS_CH2_INT_TX_CLR_0 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by tx bridge unit overflow,
parameter              PCS_CH2_INT_TX_CLR_1 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by tx_bridge_unit async fifo underflow
parameter              PCS_CH2_INT_TX_CLR_2 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by tx_invalid_k
parameter        PCS_CH2_TX_PMA_TCLK_POLINV = "PMA_TCLK",        // 1'b0:pma_tclk 1'b1:reverse of pma_tclk
parameter        PCS_CH2_TX_PCS_CLK_EN_SEL = "FALSE",        // FALSE,TRUE
parameter        PCS_CH2_TX_BRIDGE_TCLK_SEL = "PCS_TCLK",        // 1'b0: pcs_tclk 1'b1:tclk
parameter        PCS_CH2_TX_TCLK_POLINV = "TCLK",        // 1'b0:tclk 1'b1:reverse of tclk
parameter        PCS_CH2_TX_PCS_TX_RSTN = "FALSE",        // 1:pcs_tx_rstn is valued,is 0,0:pcs_tx_rstn is released
parameter        PCS_CH2_TX_SLAVE = "SLAVE",        // 1:slave channel,0:master channel
parameter        PCS_CH2_TX_BRIDGE_CLK_EN_SEL = "FALSE",        // FALSE,TRUE
parameter        PCS_CH2_DATA_WIDTH_MODE    = "X20",        // 20bit,16bit,10bit,8bit
parameter        PCS_CH2_TX_TCLK2FABRIC_SEL = "FALSE",        // FALSE,TRUE
parameter        PCS_CH2_TX_OUTZZ = "FALSE",        // 1:16bit/32bit only,0:20bit/40bit only
parameter        PCS_CH2_ENC_DUAL = "FALSE",        // FALSE,TRUE
parameter        PCS_CH2_TX_BITSLIP_DATA_MODE = "X10",        // 1: 20bit,0: 10bit
parameter   integer PCS_CH2_COMMA_REG1 = 0,        // 
parameter   integer PCS_CH2_RAPID_IMAX = 0,        // 
parameter   integer PCS_CH2_RAPID_VMIN_1 = 0,        // 
parameter   integer PCS_CH2_RAPID_VMIN_2 = 0,        // 
parameter        PCS_CH2_RX_PRBS_MODE = "DISABLE",        // Mode select:4'd0: reserved,4'd1: PRBS-7,4'd2: PRBS-15,4'd3: PRBS-23,4'd4: PRBS-31,4'd5: long "1",4'd6: long "0",4'd7: 20UI square wave,4'd8: D10_2,4'd9: PCIe complianece pattern,Others: reserved
parameter        PCS_CH2_RX_ERRCNT_CLR = "FALSE",        // FALSE,TRUE
parameter        PCS_CH2_TX_PRBS_MODE = "DISABLE",        // Mode select:4'd0: reserved,4'd1: PRBS-7,4'd2: PRBS-15,4'd3: PRBS-23,4'd4: PRBS-31,4'd5: long "1",4'd6: long "0",4'd7: 20UI square wave,4'd8: D10_2,4'd9: PCIe complianece pattern,Others: reserved
parameter        PCS_CH2_TX_INSERT_ER = "FALSE",        // FALSE,TRUE
parameter        PCS_CH2_ENABLE_PRBS_GEN = "FALSE",        // FALSE,TRUE
parameter   integer PCS_CH2_ERR_CNT = 0,        // 
parameter   integer PCS_CH2_DEFAULT_RADDR = 0,        // 
parameter   integer PCS_CH2_MASTER_CHECK_OFFSET = 0,        // 
parameter   integer PCS_CH2_DELAY_SET = 0,        // 
parameter        PCS_CH2_SEACH_OFFSET = "20BIT",        // 20bit,30bit,40bit,50bit,60bit,70bit
parameter   integer PCS_CH2_CEB_RAPIDLS_MMAX = 0,        // 
parameter   integer PCS_CH2_CTC_AFULL = 0,        // 
parameter   integer PCS_CH2_CTC_AEMPTY = 0,        // 
parameter        PCS_CH2_FAR_LOOP = "FALSE",        // FALSE,TRUE
parameter              PCS_CH2_NEAR_LOOP = "FALSE",        // FALSE,TRUE
parameter              PCS_CH2_INT_RX_MASK_0 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by pcs_lsm_synced
parameter              PCS_CH2_INT_RX_MASK_1 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by pcs_rx_mcb_status
parameter              PCS_CH2_INT_RX_MASK_2 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by channel bonding async fifo overflow
parameter              PCS_CH2_INT_RX_MASK_3 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by channel bonding async fifo underflow
parameter              PCS_CH2_INT_RX_MASK_4 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by ctc unit async fifo overflow
parameter              PCS_CH2_INT_RX_MASK_5 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by ctc unit async fifo underflow
parameter              PCS_CH2_INT_RX_MASK_6 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by rx_bridge_unit async fifo overflow
parameter              PCS_CH2_INT_RX_MASK_7 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by rx_bridge_unit async fifo underflow
parameter              PCS_CH2_INT_RX_CLR_0 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by pcs_lsm_synced
parameter              PCS_CH2_INT_RX_CLR_1 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by pcs_rx_mcb_status
parameter              PCS_CH2_INT_RX_CLR_2 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by channel bonding async fifo overflow
parameter              PCS_CH2_INT_RX_CLR_3 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by channel bonding async fifo underflow
parameter              PCS_CH2_INT_RX_CLR_4 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by ctc unit async fifo overflow
parameter              PCS_CH2_INT_RX_CLR_5 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by ctc unit async fifo underflow
parameter              PCS_CH2_INT_RX_CLR_6 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by rx_bridge_unit async fifo overflow
parameter              PCS_CH2_INT_RX_CLR_7 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by rx_bridge_unit async fifo underflow



parameter        PCS_CH3_BYPASS_WORD_ALIGN    = "FALSE",        // FALSE,TRUE
parameter           PCS_CH3_BYPASS_DENC    = "FALSE",        // FALSE,TRUE
parameter           PCS_CH3_BYPASS_BONDING    = "FALSE",        // FALSE,TRUE
parameter           PCS_CH3_BYPASS_CTC    = "FALSE",        // FALSE,TRUE
parameter           PCS_CH3_BYPASS_GEAR    = "FALSE",        // FALSE,TRUE
parameter           PCS_CH3_BYPASS_BRIDGE    = "FALSE",        // FALSE,TRUE
parameter           PCS_CH3_DATA_MODE    = "X8",        // 8bit,10bit,16bit,20bit
parameter           PCS_CH3_RX_POLARITY_INV    = "DELAY",        // 00: delay 01: bit polarity inversion 10: bit reversal 11: polarity inversion and bit reversal
parameter           PCS_CH3_ALIGN_MODE    = "1GB",        // 1GB,10GB,RAPIDIO,OUTSIDE
parameter           PCS_CH3_SAMP_16B = "X16",        // 16bit,20bit
parameter   integer PCS_CH3_COMMA_REG0 = 0,        // 
parameter   integer PCS_CH3_COMMA_MASK = 0,        // 
parameter        PCS_CH3_CEB_MODE = "10GB",        // 10GB,RAPIDIO,OUTSIDE
parameter           PCS_CH3_CTC_MODE = "1SKIP",        // 00: add or del 1 skip,01: add or del 2 skips,10: reserved ,11:4 skips
parameter   integer PCS_CH3_A_REG = 0,        // 
parameter        PCS_CH3_GE_AUTO_EN = "FALSE",        // CTC,FALSE,TRUE
parameter   integer PCS_CH3_SKIP_REG0 = 0,        // 
parameter   integer PCS_CH3_SKIP_REG1 = 0,        // 
parameter   integer PCS_CH3_SKIP_REG2 = 0,        // 
parameter   integer PCS_CH3_SKIP_REG3 = 0,        // 
parameter        PCS_CH3_DEC_DUAL = "FALSE",        // signal for 8b10b decoder module
parameter           PCS_CH3_SPLIT = "FALSE",        // signal for RX GEAR split, 1:split  0:no split, 
parameter           PCS_CH3_FIFOFLAG_CTC = "FALSE",        // FALSE,TRUE
parameter           PCS_CH3_COMMA_DET_MODE = "COMMA_PATTERN",        // 0: comma pattern mode  1: RX_CLK_SLIP mode 
parameter           PCS_CH3_ERRDETECT_SILENCE = "FALSE",        // 0: comma pattern mode  1: RX_CLK_SLIP mode 
parameter           PCS_CH3_PMA_RCLK_POLINV = "PMA_RCLK",        // 1'b0:pma_rclk 1'b1:reverse of pma_rclk
parameter           PCS_CH3_PCS_RCLK_SEL = "PMA_RCLK",        // 1'b0:pma_rclk,1'b1:pma_tclk,
parameter           PCS_CH3_MCB_RCLK_POLINV = "MCB_RCLK",        // 1'b0:mcb_rclk 1'b1:reverse of mcb_rclk
parameter        PCS_CH3_CB_RCLK_SEL = "PMA_RCLK",        // 2'b00:pma_rclk,2'b01:pma_tclk,2'b10:mcb_rclk,2'b11:reserved
parameter           PCS_CH3_AFTER_CTC_RCLK_SEL = "PMA_RCLK",        // 2'b00:pma_rclk,2'b01:pma_tclk,2'b10:mcb_rclk,2'b11:reserved
parameter           PCS_CH3_RCLK_POLINV = "RCLK",        // 1'b0:rclk 1'b1:reverse of rclk
parameter           PCS_CH3_BRIDGE_RCLK_SEL = "PMA_RCLK",        // 2'b00:pma_rclk,2'b01:pma_tclk,2'b10:mcb_rclk,2'b11:rclk
parameter           PCS_CH3_PCS_RCLK_EN = "FALSE",        // FALSE,TRUE
parameter           PCS_CH3_CB_RCLK_EN = "FALSE",        // FALSE,TRUE
parameter           PCS_CH3_AFTER_CTC_RCLK_EN = "FALSE",        // FALSE,TRUE
parameter           PCS_CH3_AFTER_CTC_RCLK_EN_GB = "FALSE",        // FALSE,TRUE
parameter           PCS_CH3_BRIDGE_RCLK_EN = "FALSE",        // FALSE,TRUE
parameter           PCS_CH3_PCS_RX_RSTN = "FALSE",        // 1:pcs_rx_rstn is valued,is 0,0:pcs_rx_rstn is released
parameter           PCS_CH3_SLAVE = "MASTER",        // 1:slave channel 0:master channel
parameter           PCS_CH3_PCIE_SLAVE = "MASTER",        // 1:slave channel 0:master channel
parameter           PCS_CH3_PCS_CB_RSTN = "FALSE",        // 1: pcs_cb_rstn is valued,is 0,0: pcs_cb_rstn is released
parameter           PCS_CH3_TX_BYPASS_BRIDGE_UINT    = "FALSE",        // FALSE,TRUE
parameter           PCS_CH3_TX_BYPASS_GEAR    = "FALSE",        // FALSE,TRUE
parameter           PCS_CH3_TX_BYPASS_ENC    = "FALSE",        // FALSE,TRUE
parameter           PCS_CH3_TX_BYPASS_BIT_SLIP    = "FALSE",        // FALSE,TRUE
parameter           PCS_CH3_TX_GEAR_SPLIT    = "FALSE",        // 1:spilt 44bits data to 22bits data,0: no spilt
parameter        PCS_CH3_TX_DRIVE_REG_MODE    = "NO_CHANGE",        // 00:no change, 01:enable polarity reverse,10:enable bit reverse, 11:enable both
parameter   integer PCS_CH3_TX_BIT_SLIP_CYCLES = 0,        // 
parameter        PCS_CH3_INT_TX_MASK_0 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by tx_bridge_unit async fifo overflow
parameter              PCS_CH3_INT_TX_MASK_1 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by tx bridge unit underflow,
parameter              PCS_CH3_INT_TX_MASK_2 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by tx_invalid_k 
parameter              PCS_CH3_INT_TX_CLR_0 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by tx bridge unit overflow,
parameter              PCS_CH3_INT_TX_CLR_1 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by tx_bridge_unit async fifo underflow
parameter              PCS_CH3_INT_TX_CLR_2 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by tx_invalid_k
parameter        PCS_CH3_TX_PMA_TCLK_POLINV = "PMA_TCLK",        // 1'b0:pma_tclk 1'b1:reverse of pma_tclk
parameter        PCS_CH3_TX_PCS_CLK_EN_SEL = "FALSE",        // FALSE,TRUE
parameter        PCS_CH3_TX_BRIDGE_TCLK_SEL = "PCS_TCLK",        // 1'b0: pcs_tclk 1'b1:tclk
parameter        PCS_CH3_TX_TCLK_POLINV = "TCLK",        // 1'b0:tclk 1'b1:reverse of tclk
parameter        PCS_CH3_TX_PCS_TX_RSTN = "FALSE",        // 1:pcs_tx_rstn is valued,is 0,0:pcs_tx_rstn is released
parameter        PCS_CH3_TX_SLAVE = "SLAVE",        // 1:slave channel,0:master channel
parameter        PCS_CH3_TX_BRIDGE_CLK_EN_SEL = "FALSE",        // FALSE,TRUE
parameter        PCS_CH3_DATA_WIDTH_MODE    = "X20",        // 20bit,16bit,10bit,8bit
parameter        PCS_CH3_TX_TCLK2FABRIC_SEL = "FALSE",        // FALSE,TRUE
parameter        PCS_CH3_TX_OUTZZ = "FALSE",        // 1:16bit/32bit only,0:20bit/40bit only
parameter        PCS_CH3_ENC_DUAL = "FALSE",        // FALSE,TRUE
parameter        PCS_CH3_TX_BITSLIP_DATA_MODE = "X10",        // 1: 20bit,0: 10bit
parameter   integer PCS_CH3_COMMA_REG1 = 0,        // 
parameter   integer PCS_CH3_RAPID_IMAX = 0,        // 
parameter   integer PCS_CH3_RAPID_VMIN_1 = 0,        // 
parameter   integer PCS_CH3_RAPID_VMIN_2 = 0,        // 
parameter        PCS_CH3_RX_PRBS_MODE = "DISABLE",        // Mode select:4'd0: reserved,4'd1: PRBS-7,4'd2: PRBS-15,4'd3: PRBS-23,4'd4: PRBS-31,4'd5: long "1",4'd6: long "0",4'd7: 20UI square wave,4'd8: D10_2,4'd9: PCIe complianece pattern,Others: reserved
parameter        PCS_CH3_RX_ERRCNT_CLR = "FALSE",        // FALSE,TRUE
parameter        PCS_CH3_TX_PRBS_MODE = "DISABLE",        // Mode select:4'd0: reserved,4'd1: PRBS-7,4'd2: PRBS-15,4'd3: PRBS-23,4'd4: PRBS-31,4'd5: long "1",4'd6: long "0",4'd7: 20UI square wave,4'd8: D10_2,4'd9: PCIe complianece pattern,Others: reserved
parameter        PCS_CH3_TX_INSERT_ER = "FALSE",        // FALSE,TRUE
parameter        PCS_CH3_ENABLE_PRBS_GEN = "FALSE",        // FALSE,TRUE
parameter   integer PCS_CH3_ERR_CNT = 0,        // 
parameter   integer PCS_CH3_DEFAULT_RADDR = 0,        // 
parameter   integer PCS_CH3_MASTER_CHECK_OFFSET = 0,        // 
parameter   integer PCS_CH3_DELAY_SET = 0,        // 
parameter        PCS_CH3_SEACH_OFFSET = "20BIT",        // 20bit,30bit,40bit,50bit,60bit,70bit
parameter   integer PCS_CH3_CEB_RAPIDLS_MMAX = 0,        // 
parameter   integer PCS_CH3_CTC_AFULL = 0,        // 
parameter   integer PCS_CH3_CTC_AEMPTY = 0,        // 
parameter        PCS_CH3_FAR_LOOP = "FALSE",        // FALSE,TRUE
parameter              PCS_CH3_NEAR_LOOP = "FALSE",        // FALSE,TRUE
parameter              PCS_CH3_INT_RX_MASK_0 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by pcs_lsm_synced
parameter              PCS_CH3_INT_RX_MASK_1 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by pcs_rx_mcb_status
parameter              PCS_CH3_INT_RX_MASK_2 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by channel bonding async fifo overflow
parameter              PCS_CH3_INT_RX_MASK_3 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by channel bonding async fifo underflow
parameter              PCS_CH3_INT_RX_MASK_4 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by ctc unit async fifo overflow
parameter              PCS_CH3_INT_RX_MASK_5 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by ctc unit async fifo underflow
parameter              PCS_CH3_INT_RX_MASK_6 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by rx_bridge_unit async fifo overflow
parameter              PCS_CH3_INT_RX_MASK_7 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by rx_bridge_unit async fifo underflow
parameter              PCS_CH3_INT_RX_CLR_0 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by pcs_lsm_synced
parameter              PCS_CH3_INT_RX_CLR_1 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by pcs_rx_mcb_status
parameter              PCS_CH3_INT_RX_CLR_2 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by channel bonding async fifo overflow
parameter              PCS_CH3_INT_RX_CLR_3 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by channel bonding async fifo underflow
parameter              PCS_CH3_INT_RX_CLR_4 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by ctc unit async fifo overflow
parameter              PCS_CH3_INT_RX_CLR_5 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by ctc unit async fifo underflow
parameter              PCS_CH3_INT_RX_CLR_6 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by rx_bridge_unit async fifo overflow
parameter              PCS_CH3_INT_RX_CLR_7 = "FALSE",        // FALSE,TRUE  active high to clr int triggered by rx_bridge_unit async fifo underflow



parameter   PMA_CH0_TXDATA_WIDTH    = "8_BIT",        // 8_BIT:2'b00, 10_BIT:2'b01, 16_BIT:2'b10, 20_BIT:2'b11
parameter   integer PMA_CH0_TX_TESTPATTERN    = 0,        // 0 to 3
parameter   PMA_CH0_TESTPATTERN_O_ENABLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH0_DISABLE_BSMODE_DRVAMP    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH0_FORCE_BIST_ENABLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH0_FORCE_ELECTRICAL_IDLE    = "FALSE",    // TRUE , FALSE 
parameter   PMA_CH0_FORCE_RXDCT_ENABLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH0_FORCE_EXTLB_ENABLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH0_DISABLE_LANE_SYNC    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH0_DISABLE_ELECTRICAL_IDLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH0_DISABLE_RXDCT_ENABLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH0_DISABLE_EXTLB_ENABLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH0_DISABLE_LOW_SPEED_PATH_ENABLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH0_FORCE_LANE_ENABLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH0_FORCE_LANE_RESETB_DISABLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH0_RXDCT_LGBW_ENABLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH0_RXDCT_VTH    = "MINUS_300MV",    // MINUS_300MV:1'b00 ,MINUS_375MV:1'b01 ,MINUS_150MV:1'b10 ,MINUS_225MV:1'b11 
parameter   PMA_CH0_DE_EMPHASIS_ADDITIONAL_CONTROL    = "0DB",        // 0db:1'b00 ,0_7db:1'b01 ,1_4db:1'b11 
parameter   PMA_CH0_DRV_RTERM_CONTROL    = "100PCT",        //  100PCT , 95PCT , 91PCT , 87PCT , 105PCT , 111PCT , 117PCT ,highZ
parameter   PMA_CH0_FDRV_AMP_CONTROL    = "100PCT",    // 100PCT , 92PCT , 109PCT , 120PCT
parameter   PMA_CH0_PREPC_AMP_CONTROL    = "100PCT",    // 100PCT , 83PCT , 133PCT , 117PCT
parameter   PMA_CH0_PREMC_AMP_CONTROL    = "100PCT",    // 100PCT , 83PCT , 133PCT , 117PCT
parameter   PMA_CH0_SER_AMP_CONTROL    = "100PCT",    // 100PCT , 83PCT , 133PCT , 117PCT
parameter   integer PMA_CH0_PFD_LOOP_RESISTOR_SETTING    = 0,        // 0 to 15
parameter   integer PMA_CH0_PD_LOOP_RESISTOR_SETTING    = 0,        // 0 to 15
parameter   PMA_CH0_CDR_TEST_OUT_SELECT    = "FBCK",    // FBCK , PD
parameter   PMA_CH0_PI_DIV1_BP    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH0_PI_TEST_FOR_CKI    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH0_PI_CURRENT_SETTING    = "100PCT",        // 100PCT,80PCT,140PCT,120PCT,160PCT,120PCTr,200PCT,180PCT
parameter   integer PMA_CH0_PI_FREQUENCY_SETTING    = 0,        // 0 to 3
parameter   PMA_CH0_TEST_OUT_SELECT_FOR_RCK    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH0_TEST_OUT_SELECT_SOURCE    = "SLPI1UI",    // SLPI1UI , PD1
parameter   PMA_CH0_TEST_DATA_OUT_SELECT_SOURCE    = "DO",    // DO , DE
parameter   PMA_CH0_TEST_CK_OUT_SELECT_SOURCE    = "DATA",    // DATA , CLOCK
parameter   PMA_CH0_ENABLE_SLIP1UI_MODULE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH0_PN_SWAP_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH0_SIPO_BIT_SETTING    = "10_BIT",        // 10_BIT:2'b00, 8_BIT:2'b01, 20_BIT:2'b10, 16_BIT:2'b11
parameter   PMA_CH0_OOB_EN    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH0_ALOS_EN    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH0_LFMODE    = "HIGH",    // HIGH , LOW
parameter   PMA_CH0_TSO_HS_SEL    = "CDR",    // CDR , EQ
parameter   PMA_CH0_LX_SELLC    = "RING",            // RING , LC
parameter   integer PMA_CH0_LX_RXPLL_DIVSEL45_FB    = 4,            // 4 , 5
parameter   integer PMA_CH0_LX_RXPLL_DIVSEL_FB    = 2,        // 2,4,5,8,10
parameter   integer PMA_CH0_LX_RXPLL_DIVSEL_REF    = 1,        // 1:2'b00 ,2:1'b01 ,4:2'b10 ,4:2'b11 
parameter   integer PMA_CH0_PICODE    = 0,        // 0 to 255 
parameter   integer PMA_CH0_RX_REFCK_SEL    = 0,        // 0 to 3
parameter   PMA_CH0_PFDLPEN_REGISTER_CONTROL_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH0_PFDLPEN_REGISTER_SETTING    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH0_PDLPEN_REGISTER_CONTROL_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH0_PDLPEN_REGISTER_SETTING    = "FALSE",    // TRUE , FALSE
parameter   integer PMA_CH0_DIV_CHANGE_ENABLE_DELAY_TIMER    = 0,        // 0 to 3
parameter   PMA_CH0_DIV_CHANGE_ENABLE_SIGNAL_GATING    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH0_CDR_ALIGN_REGISTER_SETTING_VALUE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH0_FORCE_CDR_ALIGN_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH0_SELLC_REGISTER_SETTING_VALUE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH0_SELLC_CONTROL_BY_REGISTER    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH0_REG_PLLI_LDO_VREF_SETTING    = "0_9V",        //  000:0_9V , 001:0_95V , 010:1_00V , 011:1_05V , 100: 1_1V(DF) , 101:1_15V , 110:1_20V , 111:1_25V
parameter   integer PMA_CH0_REG_PLLI_LDO_BYPASS_CURRENT    = 0,        //  0 to 7
parameter   PMA_CH0_REG_PLL_HSTEST_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH0_REG_PLL_ISNK_CURRENT_CONTROL    = "5U",        // 5U:1'B00 ,15U:1'B01 ,25U:1'B10 ,35U:1'B11 
parameter   integer PMA_CH0_REG_PLL_PFD_LOOP_CP0_CURRENT_SETTING    = 0,        // 0 to 31 
parameter   PMA_CH0_REG_PLL_PD_LOOP_PLLGM_SETTING    = "100PCT",        //  100PCT , 89PCT , 122PCT , 111PCT , 144PCT , 133PCT , 167PCT ,156PCT
parameter   integer PMA_CH0_REG_PLL_PFD_LOOP_CP1_CURRENT_SETTING    = 0,        // 0 to 31 
parameter   PMA_CH0_REG_PLL_CP0_BIAS_CONTROL    = "100PCT",        //  100PCT , 111PCT , 125PCT , 143PCT , 71PCT , 77PCT , 83PCT ,91PCT
parameter   integer PMA_CH0_REG_PLL_PD_LOOP_CP0_CURRENT_SETTING    = 0,        // 0 to 31 
parameter   PMA_CH0_REG_PLL_CP1_BIAS_CONTROL    = "100PCT",        //  100PCT , 111PCT , 125PCT , 143PCT , 71PCT , 77PCT , 83PCT ,91PCT
parameter   integer PMA_CH0_REG_PLL_PD_LOOP_CP1_CURRENT_SETTING    = 0,        // 0 to 31 
parameter   PMA_CH0_REG_PLL_CP0_CURRENT_SETTING    = "100PCT",        //  100PCT , 20PCT , 140PCT , 60PCT , 160PCT , 80PCT , 200PCT ,120PCT
parameter   PMA_CH0_REG_PLL_CP1_CURRENT_SETTING    = "100PCT",        //  100PCT , 20PCT , 140PCT , 60PCT , 160PCT , 80PCT , 200PCT ,120PCT
parameter   PMA_CH0_REG_PLL_GM1_CURRENT_SETTING    = "100PCT",        //  100PCT , 67PCT , 167PCT , 133PCT , 300PCT , 267PCT , 367PCT ,333PCT
parameter   PMA_CH0_REG_PLL_LC_BF2_CURRENT_SETTING    = "100PCT",        //  100PCT , 20PCT , 140PCT , 60PCT , 160PCT , 80PCT , 200PCT ,120PCT
parameter   PMA_CH0_REG_PLL_LC_BF2_CURRENT_SETTING_LOW    = "100PCT",        //  100PCT , 20PCT , 140PCT , 60PCT , 160PCT , 80PCT , 200PCT ,120PCT
parameter   PMA_CH0_REG_PLL_REG_CUR    = "100PCT",        //  100PCT , 80PCT , 140PCT , 120PCT , 180PCT , 160PCT , 220PCT ,200PCT
parameter   PMA_CH0_REG_PLL_LCCUR    = "DEFAULT",        //  DEFAULT , MINUS_1MA , 2MA , 1MA , 4MA , 3MA , 6MA ,5MA
parameter   PMA_CH0_REG_PLL_LCOBAS    = "100PCT",        // 100PCT , 75PCT , 150PCT , 125PCT 
parameter   PMA_CH0_REG_PLL_FB_CK_TEST_OUT_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   integer PMA_CH0_CDR_ALIGN_TIMER    = 0,        // 0 to 3
parameter   integer PMA_CH0_CALIB_WAIT    = 1024,        // 1024 , 2048 , 4096 , 512 
parameter   integer PMA_CH0_CALIB_TIMER    = 512,        // 512 , 1024 , 2048 , 4096 
parameter   integer PMA_CH0_TOT_RANGE    = 0,        // 0 to 3
parameter   integer PMA_CH0_SUB_RANGE    = 0,        // 0 to 3
parameter   integer PMA_CH0_OVLP    = 0,        // 0 to 3
parameter   integer PMA_CH0_BIST_WAIT    = 1024,        // 1024 , 2048 , 4096 , 512 
parameter   integer PMA_CH0_BIST_TIMER    = 512,        // 512 , 1024 , 2048 , 4096 
parameter   integer PMA_CH0_BAND_LB    = 0,        // 0 to 7 
parameter   integer PMA_CH0_BAND_HB    = 0,        // 0 to 31 
parameter   integer PMA_CH0_FREQ_LOCK_ACCURACY    = 0,        // 0 to 7
parameter   integer PMA_CH0_REG_SET_LC_BAND    = 0,        // 0 to 31 
parameter   integer PMA_CH0_REG_SET_VCODIV    = 0,        // 0 to 3
parameter   PMA_CH0_REGISTER_SET_VCODIV_BAND_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH0_REG_SET_PLL_LOCK    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH0_REGISTER_SET_PLL_LOCK_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH0_REG_SET_VCO_HI    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH0_REG_SET_VCO_LO    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH0_REGISTER_SET_VCO_HI_VCO_LO_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH0_FORCE_LC_PLL_LOOP_EN_H    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH0_FORCE_LC_PLL_LOOP_EN_L    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH0_VCO_DIV_CALI_BYPASS    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH0_BIST_EN    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH0_PLL_LOOP_EN_SETTING_FROM_REGISTER_ENABLE     = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH0_FREQ_DETECT_ENABLE_SOURCE     = "DISABLE",    // DISABLE , ENABLE
parameter   integer PMA_CH0_REG_SET_DIVSEL_REF    = 0,        // 0 to 3
parameter   PMA_CH0_REG_SET_DIVSEL45_FB    = "FALSE",    // TRUE , FALSE
parameter   integer PMA_CH0_REG_SET_DIVSEL_FB    = 0,        // 0 to 7  
parameter   PMA_CH0_PLL_LOOP_EN_SETTING     = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH0_REGISTER_SET_TXPLL_DIV_ENABLE     = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH0_FORCE_RXPLL_RESET    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH0_FORCE_RXPLL_ON    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH0_DPCK_DIV2    = "FALSE",    // TRUE , FALSE
parameter   integer PMA_CH0_LFO_SETTING    = 0,        // 0 to 7
parameter   PMA_CH0_ALOS_COUNTER_CLOCK_SELECTION    = "LOCAL",    // LOCAL , GLOBAL25M
parameter   PMA_CH0_RX_BIAS_CURRENT_ADJUSTMENT    = "100PCT",        //  100PCT , 111PCT , 125PCT , 143PCT , 71PCT , 77PCT , 83PCT ,91PCT
parameter   integer PMA_CH0_OOB_ENTER_DELAY_SETTING    = 0,        // 0 to 3
parameter   integer PMA_CH0_ALOS_LOW_TO_HIGH_COUNTER_SETTING    = 0,        // 0 to 3
parameter   PMA_CH0_ENABLE_ALOS_RESULT_AUTOMATICALLY_ENABLE_CHANNEL     = "DISABLE",    // DISABLE , ENABLE
parameter   integer PMA_CH0_ALOS_EXIT_COUNTER_CLOCK_DIVIDER    = 0,        // 0 to 3
parameter   integer PMA_CH0_OOB_OSCILATER_FREQUENCY_SETTING    = 0,        // 0 to 3
parameter   PMA_CH0_FORCE_OOB    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH0_OOB_VTH_SET    = "27MV",        // 27MV, 30MV, 35MV, 42_5MV, 52MV, 68MV 
parameter   PMA_CH0_FORCE_DET_FORCE_ALOS_LOW    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH0_ALOS_THRESHOLD_VOLTAGE    = "27MV",        // 27MV, 30MV, 35MV, 42_5MV, 52MV, 68MV 
parameter   integer PMA_CH0_WAKEUP_VCM_RX_COMMON_MODE_VOLTAGE    = 0,        // 0 to 3
parameter   PMA_CH0_REGR_NEGATIVE_HYSTERESIS_SETTING    = "100MV",        // 100MV, 75MV, 50MV, 25MV, 25MV, 0MV 
parameter   PMA_CH0_REGL_POSITIVE_HYSTERESIS_SETTING    = "100MV",        // 100MV, 75MV, 50MV, 25MV, 25MV, 0MV 
parameter   PMA_CH0_REG_EN    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH0_REGREF_SEL    = "VREF",    // VREF , SELF_DC
parameter   PMA_CH0_DC496    = "39_6MHZ",        // 5MHZ, 8MHZ, 11_5MHZ, 20_6MHZ, 39_6MHZ 
parameter   integer PMA_CH0_EQ2_AC_VAR_SETTING    = 0,        // 255,254,252,248,240,224,192,128,0
parameter   integer PMA_CH0_EQ2_AC_RES_SETTING    = 0,        // 0 to 31 
parameter   integer PMA_CH0_EQ2_DC_RESTOP_SETTING    = 0,        // 0 to 3
parameter   integer PMA_CH0_EQ1_DC_RESTOP_SETTING    = 50,        //  50, 60, 71, 78, 107 
parameter   integer PMA_CH0_EQ1_AC_VAR_SETTING    = 0,        // 255,254,252,248,240,224,192,128,0
parameter   integer PMA_CH0_EQ2_CURRENT_SETTING    = 0,        // 0,1,3,7
parameter   integer PMA_CH0_EQ1_AC_RES_SETTING    = 0,        // 0 to 31 
parameter   integer PMA_CH0_EQ1_CURRENT_SETTING    = 0,        // 15,7,3,9,1,0 
parameter   integer PMA_CH0_RPLUS    = 0,        // 0,1,3,7,15
parameter   integer PMA_CH0_RMINUS    = 0,        // 0,1,3,7,15
parameter   integer PMA_CH0_RVALSET    = 0,        // 0 to 3
parameter   integer PMA_CH0_RTERM    = 0,        // 0 to 3
parameter   PMA_CH0_DCFB_EN    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH0_DCCOUP    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH0_3G    = "FALSE",    // TRUE , FALSE

parameter   PMA_CH1_TXDATA_WIDTH    = "8_BIT",        // 8_BIT:2'b00, 10_BIT:2'b01, 16_BIT:2'b10, 20_BIT:2'b11
parameter   integer PMA_CH1_TX_TESTPATTERN    = 0,        // 0 to 3
parameter   PMA_CH1_TESTPATTERN_O_ENABLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH1_DISABLE_BSMODE_DRVAMP    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH1_FORCE_BIST_ENABLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH1_FORCE_ELECTRICAL_IDLE    = "FALSE",    // TRUE , FALSE 
parameter   PMA_CH1_FORCE_RXDCT_ENABLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH1_FORCE_EXTLB_ENABLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH1_DISABLE_LANE_SYNC    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH1_DISABLE_ELECTRICAL_IDLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH1_DISABLE_RXDCT_ENABLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH1_DISABLE_EXTLB_ENABLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH1_DISABLE_LOW_SPEED_PATH_ENABLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH1_FORCE_LANE_ENABLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH1_FORCE_LANE_RESETB_DISABLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH1_RXDCT_LGBW_ENABLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH1_RXDCT_VTH    = "MINUS_300MV",    // MINUS_300MV:1'b00 ,MINUS_375MV:1'b01 ,MINUS_150MV:1'b10 ,MINUS_225MV:1'b11 
parameter   PMA_CH1_DE_EMPHASIS_ADDITIONAL_CONTROL    = "0DB",        // 0db:1'b00 ,0_7db:1'b01 ,1_4db:1'b11 
parameter   PMA_CH1_DRV_RTERM_CONTROL    = "100PCT",        //  100PCT , 95PCT , 91PCT , 87PCT , 105PCT , 111PCT , 117PCT ,highZ
parameter   PMA_CH1_FDRV_AMP_CONTROL    = "100PCT",    // 100PCT , 92PCT , 109PCT , 120PCT
parameter   PMA_CH1_PREPC_AMP_CONTROL    = "100PCT",    // 100PCT , 83PCT , 133PCT , 117PCT
parameter   PMA_CH1_PREMC_AMP_CONTROL    = "100PCT",    // 100PCT , 83PCT , 133PCT , 117PCT
parameter   PMA_CH1_SER_AMP_CONTROL    = "100PCT",    // 100PCT , 83PCT , 133PCT , 117PCT
parameter   integer PMA_CH1_PFD_LOOP_RESISTOR_SETTING    = 0,        // 0 to 15
parameter   integer PMA_CH1_PD_LOOP_RESISTOR_SETTING    = 0,        // 0 to 15
parameter   PMA_CH1_CDR_TEST_OUT_SELECT    = "FBCK",    // FBCK , PD
parameter   PMA_CH1_PI_DIV1_BP    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH1_PI_TEST_FOR_CKI    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH1_PI_CURRENT_SETTING    = "100PCT",        // 100PCT,80PCT,140PCT,120PCT,160PCT,120PCTr,200PCT,180PCT
parameter   integer PMA_CH1_PI_FREQUENCY_SETTING    = 0,        // 0 to 3
parameter   PMA_CH1_TEST_OUT_SELECT_FOR_RCK    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH1_TEST_OUT_SELECT_SOURCE    = "SLPI1UI",    // SLPI1UI , PD1
parameter   PMA_CH1_TEST_DATA_OUT_SELECT_SOURCE    = "DO",    // DO , DE
parameter   PMA_CH1_TEST_CK_OUT_SELECT_SOURCE    = "DATA",    // DATA , CLOCK
parameter   PMA_CH1_ENABLE_SLIP1UI_MODULE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH1_PN_SWAP_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH1_SIPO_BIT_SETTING    = "10_BIT",        // 10_BIT:2'b00, 8_BIT:2'b01, 20_BIT:2'b10, 16_BIT:2'b11
parameter   PMA_CH1_OOB_EN    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH1_ALOS_EN    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH1_LFMODE    = "HIGH",    // HIGH , LOW
parameter   PMA_CH1_TSO_HS_SEL    = "CDR",    // CDR , EQ
parameter   PMA_CH1_LX_SELLC    = "RING",            // RING , LC
parameter   integer PMA_CH1_LX_RXPLL_DIVSEL45_FB    = 4,            // 4 , 5
parameter   integer PMA_CH1_LX_RXPLL_DIVSEL_FB    = 2,        // 2,4,5,8,10
parameter   integer PMA_CH1_LX_RXPLL_DIVSEL_REF    = 1,        // 1:2'b00 ,2:1'b01 ,4:2'b10 ,4:2'b11 
parameter   integer PMA_CH1_PICODE    = 0,        // 0 to 255 
parameter   integer PMA_CH1_RX_REFCK_SEL    = 0,        // 0 to 3
parameter   PMA_CH1_PFDLPEN_REGISTER_CONTROL_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH1_PFDLPEN_REGISTER_SETTING    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH1_PDLPEN_REGISTER_CONTROL_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH1_PDLPEN_REGISTER_SETTING    = "FALSE",    // TRUE , FALSE
parameter   integer PMA_CH1_DIV_CHANGE_ENABLE_DELAY_TIMER    = 0,        // 0 to 3
parameter   PMA_CH1_DIV_CHANGE_ENABLE_SIGNAL_GATING    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH1_CDR_ALIGN_REGISTER_SETTING_VALUE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH1_FORCE_CDR_ALIGN_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH1_SELLC_REGISTER_SETTING_VALUE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH1_SELLC_CONTROL_BY_REGISTER    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH1_REG_PLLI_LDO_VREF_SETTING    = "0_9V",        //  000:0_9V , 001:0_95V , 010:1_00V , 011:1_05V , 100: 1_1V(DF) , 101:1_15V , 110:1_20V , 111:1_25V
parameter   integer PMA_CH1_REG_PLLI_LDO_BYPASS_CURRENT    = 0,        //  0 to 7
parameter   PMA_CH1_REG_PLL_HSTEST_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH1_REG_PLL_ISNK_CURRENT_CONTROL    = "5U",        // 5U:1'B00 ,15U:1'B01 ,25U:1'B10 ,35U:1'B11 
parameter   integer PMA_CH1_REG_PLL_PFD_LOOP_CP0_CURRENT_SETTING    = 0,        // 0 to 31 
parameter   PMA_CH1_REG_PLL_PD_LOOP_PLLGM_SETTING    = "100PCT",        //  100PCT , 89PCT , 122PCT , 111PCT , 144PCT , 133PCT , 167PCT ,156PCT
parameter   integer PMA_CH1_REG_PLL_PFD_LOOP_CP1_CURRENT_SETTING    = 0,        // 0 to 31 
parameter   PMA_CH1_REG_PLL_CP0_BIAS_CONTROL    = "100PCT",        //  100PCT , 111PCT , 125PCT , 143PCT , 71PCT , 77PCT , 83PCT ,91PCT
parameter   integer PMA_CH1_REG_PLL_PD_LOOP_CP0_CURRENT_SETTING    = 0,        // 0 to 31 
parameter   PMA_CH1_REG_PLL_CP1_BIAS_CONTROL    = "100PCT",        //  100PCT , 111PCT , 125PCT , 143PCT , 71PCT , 77PCT , 83PCT ,91PCT
parameter   integer PMA_CH1_REG_PLL_PD_LOOP_CP1_CURRENT_SETTING    = 0,        // 0 to 31 
parameter   PMA_CH1_REG_PLL_CP0_CURRENT_SETTING    = "100PCT",        //  100PCT , 20PCT , 140PCT , 60PCT , 160PCT , 80PCT , 200PCT ,120PCT
parameter   PMA_CH1_REG_PLL_CP1_CURRENT_SETTING    = "100PCT",        //  100PCT , 20PCT , 140PCT , 60PCT , 160PCT , 80PCT , 200PCT ,120PCT
parameter   PMA_CH1_REG_PLL_GM1_CURRENT_SETTING    = "100PCT",        //  100PCT , 67PCT , 167PCT , 133PCT , 300PCT , 267PCT , 367PCT ,333PCT
parameter   PMA_CH1_REG_PLL_LC_BF2_CURRENT_SETTING    = "100PCT",        //  100PCT , 20PCT , 140PCT , 60PCT , 160PCT , 80PCT , 200PCT ,120PCT
parameter   PMA_CH1_REG_PLL_LC_BF2_CURRENT_SETTING_LOW    = "100PCT",        //  100PCT , 20PCT , 140PCT , 60PCT , 160PCT , 80PCT , 200PCT ,120PCT
parameter   PMA_CH1_REG_PLL_REG_CUR    = "100PCT",        //  100PCT , 80PCT , 140PCT , 120PCT , 180PCT , 160PCT , 220PCT ,200PCT
parameter   PMA_CH1_REG_PLL_LCCUR    = "DEFAULT",        //  DEFAULT , MINUS_1MA , 2MA , 1MA , 4MA , 3MA , 6MA ,5MA
parameter   PMA_CH1_REG_PLL_LCOBAS    = "100PCT",        // 100PCT , 75PCT , 150PCT , 125PCT 
parameter   PMA_CH1_REG_PLL_FB_CK_TEST_OUT_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   integer PMA_CH1_CDR_ALIGN_TIMER    = 0,        // 0 to 3
parameter   integer PMA_CH1_CALIB_WAIT    = 1024,        // 1024 , 2048 , 4096 , 512 
parameter   integer PMA_CH1_CALIB_TIMER    = 512,        // 512 , 1024 , 2048 , 4096 
parameter   integer PMA_CH1_TOT_RANGE    = 0,        // 0 to 3
parameter   integer PMA_CH1_SUB_RANGE    = 0,        // 0 to 3
parameter   integer PMA_CH1_OVLP    = 0,        // 0 to 3
parameter   integer PMA_CH1_BIST_WAIT    = 1024,        // 1024 , 2048 , 4096 , 512 
parameter   integer PMA_CH1_BIST_TIMER    = 512,        // 512 , 1024 , 2048 , 4096 
parameter   integer PMA_CH1_BAND_LB    = 0,        // 0 to 7 
parameter   integer PMA_CH1_BAND_HB    = 0,        // 0 to 31 
parameter   integer PMA_CH1_FREQ_LOCK_ACCURACY    = 0,        // 0 to 7
parameter   integer PMA_CH1_REG_SET_LC_BAND    = 0,        // 0 to 31 
parameter   integer PMA_CH1_REG_SET_VCODIV    = 0,        // 0 to 3
parameter   PMA_CH1_REGISTER_SET_VCODIV_BAND_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH1_REG_SET_PLL_LOCK    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH1_REGISTER_SET_PLL_LOCK_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH1_REG_SET_VCO_HI    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH1_REG_SET_VCO_LO    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH1_REGISTER_SET_VCO_HI_VCO_LO_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH1_FORCE_LC_PLL_LOOP_EN_H    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH1_FORCE_LC_PLL_LOOP_EN_L    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH1_VCO_DIV_CALI_BYPASS    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH1_BIST_EN    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH1_PLL_LOOP_EN_SETTING_FROM_REGISTER_ENABLE     = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH1_FREQ_DETECT_ENABLE_SOURCE     = "DISABLE",    // DISABLE , ENABLE
parameter   integer PMA_CH1_REG_SET_DIVSEL_REF    = 0,        // 0 to 3
parameter   PMA_CH1_REG_SET_DIVSEL45_FB    = "FALSE",    // TRUE , FALSE
parameter   integer PMA_CH1_REG_SET_DIVSEL_FB    = 0,        // 0 to 7  
parameter   PMA_CH1_PLL_LOOP_EN_SETTING     = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH1_REGISTER_SET_TXPLL_DIV_ENABLE     = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH1_FORCE_RXPLL_RESET    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH1_FORCE_RXPLL_ON    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH1_DPCK_DIV2    = "FALSE",    // TRUE , FALSE
parameter   integer PMA_CH1_LFO_SETTING    = 0,        // 0 to 7
parameter   PMA_CH1_ALOS_COUNTER_CLOCK_SELECTION    = "LOCAL",    // LOCAL , GLOBAL25M
parameter   PMA_CH1_RX_BIAS_CURRENT_ADJUSTMENT    = "100PCT",        //  100PCT , 111PCT , 125PCT , 143PCT , 71PCT , 77PCT , 83PCT ,91PCT
parameter   integer PMA_CH1_OOB_ENTER_DELAY_SETTING    = 0,        // 0 to 3
parameter   integer PMA_CH1_ALOS_LOW_TO_HIGH_COUNTER_SETTING    = 0,        // 0 to 3
parameter   PMA_CH1_ENABLE_ALOS_RESULT_AUTOMATICALLY_ENABLE_CHANNEL     = "DISABLE",    // DISABLE , ENABLE
parameter   integer PMA_CH1_ALOS_EXIT_COUNTER_CLOCK_DIVIDER    = 0,        // 0 to 3
parameter   integer PMA_CH1_OOB_OSCILATER_FREQUENCY_SETTING    = 0,        // 0 to 3
parameter   PMA_CH1_FORCE_OOB    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH1_OOB_VTH_SET    = "27MV",        // 27MV, 30MV, 35MV, 42_5MV, 52MV, 68MV 
parameter   PMA_CH1_FORCE_DET_FORCE_ALOS_LOW    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH1_ALOS_THRESHOLD_VOLTAGE    = "27MV",        // 27MV, 30MV, 35MV, 42_5MV, 52MV, 68MV 
parameter   integer PMA_CH1_WAKEUP_VCM_RX_COMMON_MODE_VOLTAGE    = 0,        // 0 to 3
parameter   PMA_CH1_REGR_NEGATIVE_HYSTERESIS_SETTING    = "100MV",        // 100MV, 75MV, 50MV, 25MV, 25MV, 0MV 
parameter   PMA_CH1_REGL_POSITIVE_HYSTERESIS_SETTING    = "100MV",        // 100MV, 75MV, 50MV, 25MV, 25MV, 0MV 
parameter   PMA_CH1_REG_EN    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH1_REGREF_SEL    = "VREF",    // VREF , SELF_DC
parameter   PMA_CH1_DC496    = "39_6MHZ",        // 5MHZ, 8MHZ, 11_5MHZ, 20_6MHZ, 39_6MHZ 
parameter   integer PMA_CH1_EQ2_AC_VAR_SETTING    = 0,        // 255,254,252,248,240,224,192,128,0
parameter   integer PMA_CH1_EQ2_AC_RES_SETTING    = 0,        // 0 to 31 
parameter   integer PMA_CH1_EQ2_DC_RESTOP_SETTING    = 0,        // 0 to 3
parameter   integer PMA_CH1_EQ1_DC_RESTOP_SETTING    = 50,        //  50, 60, 71, 78, 107 
parameter   integer PMA_CH1_EQ1_AC_VAR_SETTING    = 0,        // 255,254,252,248,240,224,192,128,0
parameter   integer PMA_CH1_EQ2_CURRENT_SETTING    = 0,        // 0,1,3,7
parameter   integer PMA_CH1_EQ1_AC_RES_SETTING    = 0,        // 0 to 31 
parameter   integer PMA_CH1_EQ1_CURRENT_SETTING    = 0,        // 15,7,3,9,1,0 
parameter   integer PMA_CH1_RPLUS    = 0,        // 0,1,3,7,15
parameter   integer PMA_CH1_RMINUS    = 0,        // 0,1,3,7,15
parameter   integer PMA_CH1_RVALSET    = 0,        // 0 to 3
parameter   integer PMA_CH1_RTERM    = 0,        // 0 to 3
parameter   PMA_CH1_DCFB_EN    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH1_DCCOUP    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH1_3G    = "FALSE",    // TRUE , FALSE

parameter   PMA_CH2_TXDATA_WIDTH    = "8_BIT",        // 8_BIT:2'b00, 10_BIT:2'b01, 16_BIT:2'b10, 20_BIT:2'b11
parameter   integer PMA_CH2_TX_TESTPATTERN    = 0,        // 0 to 3
parameter   PMA_CH2_TESTPATTERN_O_ENABLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH2_DISABLE_BSMODE_DRVAMP    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH2_FORCE_BIST_ENABLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH2_FORCE_ELECTRICAL_IDLE    = "FALSE",    // TRUE , FALSE 
parameter   PMA_CH2_FORCE_RXDCT_ENABLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH2_FORCE_EXTLB_ENABLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH2_DISABLE_LANE_SYNC    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH2_DISABLE_ELECTRICAL_IDLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH2_DISABLE_RXDCT_ENABLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH2_DISABLE_EXTLB_ENABLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH2_DISABLE_LOW_SPEED_PATH_ENABLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH2_FORCE_LANE_ENABLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH2_FORCE_LANE_RESETB_DISABLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH2_RXDCT_LGBW_ENABLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH2_RXDCT_VTH    = "MINUS_300MV",    // MINUS_300MV:1'b00 ,MINUS_375MV:1'b01 ,MINUS_150MV:1'b10 ,MINUS_225MV:1'b11 
parameter   PMA_CH2_DE_EMPHASIS_ADDITIONAL_CONTROL    = "0DB",        // 0db:1'b00 ,0_7db:1'b01 ,1_4db:1'b11 
parameter   PMA_CH2_DRV_RTERM_CONTROL    = "100PCT",        //  100PCT , 95PCT , 91PCT , 87PCT , 105PCT , 111PCT , 117PCT ,highZ
parameter   PMA_CH2_FDRV_AMP_CONTROL    = "100PCT",    // 100PCT , 92PCT , 109PCT , 120PCT
parameter   PMA_CH2_PREPC_AMP_CONTROL    = "100PCT",    // 100PCT , 83PCT , 133PCT , 117PCT
parameter   PMA_CH2_PREMC_AMP_CONTROL    = "100PCT",    // 100PCT , 83PCT , 133PCT , 117PCT
parameter   PMA_CH2_SER_AMP_CONTROL    = "100PCT",    // 100PCT , 83PCT , 133PCT , 117PCT
parameter   integer PMA_CH2_PFD_LOOP_RESISTOR_SETTING    = 0,        // 0 to 15
parameter   integer PMA_CH2_PD_LOOP_RESISTOR_SETTING    = 0,        // 0 to 15
parameter   PMA_CH2_CDR_TEST_OUT_SELECT    = "FBCK",    // FBCK , PD
parameter   PMA_CH2_PI_DIV1_BP    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH2_PI_TEST_FOR_CKI    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH2_PI_CURRENT_SETTING    = "100PCT",        // 100PCT,80PCT,140PCT,120PCT,160PCT,120PCTr,200PCT,180PCT
parameter   integer PMA_CH2_PI_FREQUENCY_SETTING    = 0,        // 0 to 3
parameter   PMA_CH2_TEST_OUT_SELECT_FOR_RCK    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH2_TEST_OUT_SELECT_SOURCE    = "SLPI1UI",    // SLPI1UI , PD1
parameter   PMA_CH2_TEST_DATA_OUT_SELECT_SOURCE    = "DO",    // DO , DE
parameter   PMA_CH2_TEST_CK_OUT_SELECT_SOURCE    = "DATA",    // DATA , CLOCK
parameter   PMA_CH2_ENABLE_SLIP1UI_MODULE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH2_PN_SWAP_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH2_SIPO_BIT_SETTING    = "10_BIT",        // 10_BIT:2'b00, 8_BIT:2'b01, 20_BIT:2'b10, 16_BIT:2'b11
parameter   PMA_CH2_OOB_EN    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH2_ALOS_EN    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH2_LFMODE    = "HIGH",    // HIGH , LOW
parameter   PMA_CH2_TSO_HS_SEL    = "CDR",    // CDR , EQ
parameter   PMA_CH2_LX_SELLC    = "RING",            // RING , LC
parameter   integer PMA_CH2_LX_RXPLL_DIVSEL45_FB    = 4,            // 4 , 5
parameter   integer PMA_CH2_LX_RXPLL_DIVSEL_FB    = 2,        // 2,4,5,8,10
parameter   integer PMA_CH2_LX_RXPLL_DIVSEL_REF    = 1,        // 1:2'b00 ,2:1'b01 ,4:2'b10 ,4:2'b11 
parameter   integer PMA_CH2_PICODE    = 0,        // 0 to 255 
parameter   integer PMA_CH2_RX_REFCK_SEL    = 0,        // 0 to 3
parameter   PMA_CH2_PFDLPEN_REGISTER_CONTROL_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH2_PFDLPEN_REGISTER_SETTING    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH2_PDLPEN_REGISTER_CONTROL_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH2_PDLPEN_REGISTER_SETTING    = "FALSE",    // TRUE , FALSE
parameter   integer PMA_CH2_DIV_CHANGE_ENABLE_DELAY_TIMER    = 0,        // 0 to 3
parameter   PMA_CH2_DIV_CHANGE_ENABLE_SIGNAL_GATING    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH2_CDR_ALIGN_REGISTER_SETTING_VALUE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH2_FORCE_CDR_ALIGN_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH2_SELLC_REGISTER_SETTING_VALUE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH2_SELLC_CONTROL_BY_REGISTER    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH2_REG_PLLI_LDO_VREF_SETTING    = "0_9V",        //  000:0_9V , 001:0_95V , 010:1_00V , 011:1_05V , 100: 1_1V(DF) , 101:1_15V , 110:1_20V , 111:1_25V
parameter   integer PMA_CH2_REG_PLLI_LDO_BYPASS_CURRENT    = 0,        //  0 to 7
parameter   PMA_CH2_REG_PLL_HSTEST_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH2_REG_PLL_ISNK_CURRENT_CONTROL    = "5U",        // 5U:1'B00 ,15U:1'B01 ,25U:1'B10 ,35U:1'B11 
parameter   integer PMA_CH2_REG_PLL_PFD_LOOP_CP0_CURRENT_SETTING    = 0,        // 0 to 31 
parameter   PMA_CH2_REG_PLL_PD_LOOP_PLLGM_SETTING    = "100PCT",        //  100PCT , 89PCT , 122PCT , 111PCT , 144PCT , 133PCT , 167PCT ,156PCT
parameter   integer PMA_CH2_REG_PLL_PFD_LOOP_CP1_CURRENT_SETTING    = 0,        // 0 to 31 
parameter   PMA_CH2_REG_PLL_CP0_BIAS_CONTROL    = "100PCT",        //  100PCT , 111PCT , 125PCT , 143PCT , 71PCT , 77PCT , 83PCT ,91PCT
parameter   integer PMA_CH2_REG_PLL_PD_LOOP_CP0_CURRENT_SETTING    = 0,        // 0 to 31 
parameter   PMA_CH2_REG_PLL_CP1_BIAS_CONTROL    = "100PCT",        //  100PCT , 111PCT , 125PCT , 143PCT , 71PCT , 77PCT , 83PCT ,91PCT
parameter   integer PMA_CH2_REG_PLL_PD_LOOP_CP1_CURRENT_SETTING    = 0,        // 0 to 31 
parameter   PMA_CH2_REG_PLL_CP0_CURRENT_SETTING    = "100PCT",        //  100PCT , 20PCT , 140PCT , 60PCT , 160PCT , 80PCT , 200PCT ,120PCT
parameter   PMA_CH2_REG_PLL_CP1_CURRENT_SETTING    = "100PCT",        //  100PCT , 20PCT , 140PCT , 60PCT , 160PCT , 80PCT , 200PCT ,120PCT
parameter   PMA_CH2_REG_PLL_GM1_CURRENT_SETTING    = "100PCT",        //  100PCT , 67PCT , 167PCT , 133PCT , 300PCT , 267PCT , 367PCT ,333PCT
parameter   PMA_CH2_REG_PLL_LC_BF2_CURRENT_SETTING    = "100PCT",        //  100PCT , 20PCT , 140PCT , 60PCT , 160PCT , 80PCT , 200PCT ,120PCT
parameter   PMA_CH2_REG_PLL_LC_BF2_CURRENT_SETTING_LOW    = "100PCT",        //  100PCT , 20PCT , 140PCT , 60PCT , 160PCT , 80PCT , 200PCT ,120PCT
parameter   PMA_CH2_REG_PLL_REG_CUR    = "100PCT",        //  100PCT , 80PCT , 140PCT , 120PCT , 180PCT , 160PCT , 220PCT ,200PCT
parameter   PMA_CH2_REG_PLL_LCCUR    = "DEFAULT",        //  DEFAULT , MINUS_1MA , 2MA , 1MA , 4MA , 3MA , 6MA ,5MA
parameter   PMA_CH2_REG_PLL_LCOBAS    = "100PCT",        // 100PCT , 75PCT , 150PCT , 125PCT 
parameter   PMA_CH2_REG_PLL_FB_CK_TEST_OUT_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   integer PMA_CH2_CDR_ALIGN_TIMER    = 0,        // 0 to 3
parameter   integer PMA_CH2_CALIB_WAIT    = 1024,        // 1024 , 2048 , 4096 , 512 
parameter   integer PMA_CH2_CALIB_TIMER    = 512,        // 512 , 1024 , 2048 , 4096 
parameter   integer PMA_CH2_TOT_RANGE    = 0,        // 0 to 3
parameter   integer PMA_CH2_SUB_RANGE    = 0,        // 0 to 3
parameter   integer PMA_CH2_OVLP    = 0,        // 0 to 3
parameter   integer PMA_CH2_BIST_WAIT    = 1024,        // 1024 , 2048 , 4096 , 512 
parameter   integer PMA_CH2_BIST_TIMER    = 512,        // 512 , 1024 , 2048 , 4096 
parameter   integer PMA_CH2_BAND_LB    = 0,        // 0 to 7 
parameter   integer PMA_CH2_BAND_HB    = 0,        // 0 to 31 
parameter   integer PMA_CH2_FREQ_LOCK_ACCURACY    = 0,        // 0 to 7
parameter   integer PMA_CH2_REG_SET_LC_BAND    = 0,        // 0 to 31 
parameter   integer PMA_CH2_REG_SET_VCODIV    = 0,        // 0 to 3
parameter   PMA_CH2_REGISTER_SET_VCODIV_BAND_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH2_REG_SET_PLL_LOCK    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH2_REGISTER_SET_PLL_LOCK_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH2_REG_SET_VCO_HI    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH2_REG_SET_VCO_LO    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH2_REGISTER_SET_VCO_HI_VCO_LO_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH2_FORCE_LC_PLL_LOOP_EN_H    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH2_FORCE_LC_PLL_LOOP_EN_L    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH2_VCO_DIV_CALI_BYPASS    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH2_BIST_EN    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH2_PLL_LOOP_EN_SETTING_FROM_REGISTER_ENABLE     = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH2_FREQ_DETECT_ENABLE_SOURCE     = "DISABLE",    // DISABLE , ENABLE
parameter   integer PMA_CH2_REG_SET_DIVSEL_REF    = 0,        // 0 to 3
parameter   PMA_CH2_REG_SET_DIVSEL45_FB    = "FALSE",    // TRUE , FALSE
parameter   integer PMA_CH2_REG_SET_DIVSEL_FB    = 0,        // 0 to 7  
parameter   PMA_CH2_PLL_LOOP_EN_SETTING     = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH2_REGISTER_SET_TXPLL_DIV_ENABLE     = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH2_FORCE_RXPLL_RESET    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH2_FORCE_RXPLL_ON    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH2_DPCK_DIV2    = "FALSE",    // TRUE , FALSE
parameter   integer PMA_CH2_LFO_SETTING    = 0,        // 0 to 7
parameter   PMA_CH2_ALOS_COUNTER_CLOCK_SELECTION    = "LOCAL",    // LOCAL , GLOBAL25M
parameter   PMA_CH2_RX_BIAS_CURRENT_ADJUSTMENT    = "100PCT",        //  100PCT , 111PCT , 125PCT , 143PCT , 71PCT , 77PCT , 83PCT ,91PCT
parameter   integer PMA_CH2_OOB_ENTER_DELAY_SETTING    = 0,        // 0 to 3
parameter   integer PMA_CH2_ALOS_LOW_TO_HIGH_COUNTER_SETTING    = 0,        // 0 to 3
parameter   PMA_CH2_ENABLE_ALOS_RESULT_AUTOMATICALLY_ENABLE_CHANNEL     = "DISABLE",    // DISABLE , ENABLE
parameter   integer PMA_CH2_ALOS_EXIT_COUNTER_CLOCK_DIVIDER    = 0,        // 0 to 3
parameter   integer PMA_CH2_OOB_OSCILATER_FREQUENCY_SETTING    = 0,        // 0 to 3
parameter   PMA_CH2_FORCE_OOB    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH2_OOB_VTH_SET    = "27MV",        // 27MV, 30MV, 35MV, 42_5MV, 52MV, 68MV 
parameter   PMA_CH2_FORCE_DET_FORCE_ALOS_LOW    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH2_ALOS_THRESHOLD_VOLTAGE    = "27MV",        // 27MV, 30MV, 35MV, 42_5MV, 52MV, 68MV 
parameter   integer PMA_CH2_WAKEUP_VCM_RX_COMMON_MODE_VOLTAGE    = 0,        // 0 to 3
parameter   PMA_CH2_REGR_NEGATIVE_HYSTERESIS_SETTING    = "100MV",        // 100MV, 75MV, 50MV, 25MV, 25MV, 0MV 
parameter   PMA_CH2_REGL_POSITIVE_HYSTERESIS_SETTING    = "100MV",        // 100MV, 75MV, 50MV, 25MV, 25MV, 0MV 
parameter   PMA_CH2_REG_EN    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH2_REGREF_SEL    = "VREF",    // VREF , SELF_DC
parameter   PMA_CH2_DC496    = "39_6MHZ",        // 5MHZ, 8MHZ, 11_5MHZ, 20_6MHZ, 39_6MHZ 
parameter   integer PMA_CH2_EQ2_AC_VAR_SETTING    = 0,        // 255,254,252,248,240,224,192,128,0
parameter   integer PMA_CH2_EQ2_AC_RES_SETTING    = 0,        // 0 to 31 
parameter   integer PMA_CH2_EQ2_DC_RESTOP_SETTING    = 0,        // 0 to 3
parameter   integer PMA_CH2_EQ1_DC_RESTOP_SETTING    = 50,        //  50, 60, 71, 78, 107 
parameter   integer PMA_CH2_EQ1_AC_VAR_SETTING    = 0,        // 255,254,252,248,240,224,192,128,0
parameter   integer PMA_CH2_EQ2_CURRENT_SETTING    = 0,        // 0,1,3,7
parameter   integer PMA_CH2_EQ1_AC_RES_SETTING    = 0,        // 0 to 31 
parameter   integer PMA_CH2_EQ1_CURRENT_SETTING    = 0,        // 15,7,3,9,1,0 
parameter   integer PMA_CH2_RPLUS    = 0,        // 0,1,3,7,15
parameter   integer PMA_CH2_RMINUS    = 0,        // 0,1,3,7,15
parameter   integer PMA_CH2_RVALSET    = 0,        // 0 to 3
parameter   integer PMA_CH2_RTERM    = 0,        // 0 to 3
parameter   PMA_CH2_DCFB_EN    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH2_DCCOUP    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH2_3G    = "FALSE",    // TRUE , FALSE

parameter   PMA_CH3_TXDATA_WIDTH    = "8_BIT",        // 8_BIT:2'b00, 10_BIT:2'b01, 16_BIT:2'b10, 20_BIT:2'b11
parameter   integer PMA_CH3_TX_TESTPATTERN    = 0,        // 0 to 3
parameter   PMA_CH3_TESTPATTERN_O_ENABLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH3_DISABLE_BSMODE_DRVAMP    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH3_FORCE_BIST_ENABLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH3_FORCE_ELECTRICAL_IDLE    = "FALSE",    // TRUE , FALSE 
parameter   PMA_CH3_FORCE_RXDCT_ENABLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH3_FORCE_EXTLB_ENABLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH3_DISABLE_LANE_SYNC    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH3_DISABLE_ELECTRICAL_IDLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH3_DISABLE_RXDCT_ENABLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH3_DISABLE_EXTLB_ENABLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH3_DISABLE_LOW_SPEED_PATH_ENABLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH3_FORCE_LANE_ENABLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH3_FORCE_LANE_RESETB_DISABLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH3_RXDCT_LGBW_ENABLE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH3_RXDCT_VTH    = "MINUS_300MV",    // MINUS_300MV:1'b00 ,MINUS_375MV:1'b01 ,MINUS_150MV:1'b10 ,MINUS_225MV:1'b11 
parameter   PMA_CH3_DE_EMPHASIS_ADDITIONAL_CONTROL    = "0DB",        // 0db:1'b00 ,0_7db:1'b01 ,1_4db:1'b11 
parameter   PMA_CH3_DRV_RTERM_CONTROL    = "100PCT",        //  100PCT , 95PCT , 91PCT , 87PCT , 105PCT , 111PCT , 117PCT ,highZ
parameter   PMA_CH3_FDRV_AMP_CONTROL    = "100PCT",    // 100PCT , 92PCT , 109PCT , 120PCT
parameter   PMA_CH3_PREPC_AMP_CONTROL    = "100PCT",    // 100PCT , 83PCT , 133PCT , 117PCT
parameter   PMA_CH3_PREMC_AMP_CONTROL    = "100PCT",    // 100PCT , 83PCT , 133PCT , 117PCT
parameter   PMA_CH3_SER_AMP_CONTROL    = "100PCT",    // 100PCT , 83PCT , 133PCT , 117PCT
parameter   integer PMA_CH3_PFD_LOOP_RESISTOR_SETTING    = 0,        // 0 to 15
parameter   integer PMA_CH3_PD_LOOP_RESISTOR_SETTING    = 0,        // 0 to 15
parameter   PMA_CH3_CDR_TEST_OUT_SELECT    = "FBCK",    // FBCK , PD
parameter   PMA_CH3_PI_DIV1_BP    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH3_PI_TEST_FOR_CKI    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH3_PI_CURRENT_SETTING    = "100PCT",        // 100PCT,80PCT,140PCT,120PCT,160PCT,120PCTr,200PCT,180PCT
parameter   integer PMA_CH3_PI_FREQUENCY_SETTING    = 0,        // 0 to 3
parameter   PMA_CH3_TEST_OUT_SELECT_FOR_RCK    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH3_TEST_OUT_SELECT_SOURCE    = "SLPI1UI",    // SLPI1UI , PD1
parameter   PMA_CH3_TEST_DATA_OUT_SELECT_SOURCE    = "DO",    // DO , DE
parameter   PMA_CH3_TEST_CK_OUT_SELECT_SOURCE    = "DATA",    // DATA , CLOCK
parameter   PMA_CH3_ENABLE_SLIP1UI_MODULE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH3_PN_SWAP_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH3_SIPO_BIT_SETTING    = "10_BIT",        // 10_BIT:2'b00, 8_BIT:2'b01, 20_BIT:2'b10, 16_BIT:2'b11
parameter   PMA_CH3_OOB_EN    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH3_ALOS_EN    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH3_LFMODE    = "HIGH",    // HIGH , LOW
parameter   PMA_CH3_TSO_HS_SEL    = "CDR",    // CDR , EQ
parameter   PMA_CH3_LX_SELLC    = "RING",            // RING , LC
parameter   integer PMA_CH3_LX_RXPLL_DIVSEL45_FB    = 4,            // 4 , 5
parameter   integer PMA_CH3_LX_RXPLL_DIVSEL_FB    = 2,        // 2,4,5,8,10
parameter   integer PMA_CH3_LX_RXPLL_DIVSEL_REF    = 1,        // 1:2'b00 ,2:1'b01 ,4:2'b10 ,4:2'b11 
parameter   integer PMA_CH3_PICODE    = 0,        // 0 to 255 
parameter   integer PMA_CH3_RX_REFCK_SEL    = 0,        // 0 to 3
parameter   PMA_CH3_PFDLPEN_REGISTER_CONTROL_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH3_PFDLPEN_REGISTER_SETTING    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH3_PDLPEN_REGISTER_CONTROL_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH3_PDLPEN_REGISTER_SETTING    = "FALSE",    // TRUE , FALSE
parameter   integer PMA_CH3_DIV_CHANGE_ENABLE_DELAY_TIMER    = 0,        // 0 to 3
parameter   PMA_CH3_DIV_CHANGE_ENABLE_SIGNAL_GATING    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH3_CDR_ALIGN_REGISTER_SETTING_VALUE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH3_FORCE_CDR_ALIGN_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH3_SELLC_REGISTER_SETTING_VALUE    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH3_SELLC_CONTROL_BY_REGISTER    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH3_REG_PLLI_LDO_VREF_SETTING    = "0_9V",        //  000:0_9V , 001:0_95V , 010:1_00V , 011:1_05V , 100: 1_1V(DF) , 101:1_15V , 110:1_20V , 111:1_25V
parameter   integer PMA_CH3_REG_PLLI_LDO_BYPASS_CURRENT    = 0,        //  0 to 7
parameter   PMA_CH3_REG_PLL_HSTEST_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH3_REG_PLL_ISNK_CURRENT_CONTROL    = "5U",        // 5U:1'B00 ,15U:1'B01 ,25U:1'B10 ,35U:1'B11 
parameter   integer PMA_CH3_REG_PLL_PFD_LOOP_CP0_CURRENT_SETTING    = 0,        // 0 to 31 
parameter   PMA_CH3_REG_PLL_PD_LOOP_PLLGM_SETTING    = "100PCT",        //  100PCT , 89PCT , 122PCT , 111PCT , 144PCT , 133PCT , 167PCT ,156PCT
parameter   integer PMA_CH3_REG_PLL_PFD_LOOP_CP1_CURRENT_SETTING    = 0,        // 0 to 31 
parameter   PMA_CH3_REG_PLL_CP0_BIAS_CONTROL    = "100PCT",        //  100PCT , 111PCT , 125PCT , 143PCT , 71PCT , 77PCT , 83PCT ,91PCT
parameter   integer PMA_CH3_REG_PLL_PD_LOOP_CP0_CURRENT_SETTING    = 0,        // 0 to 31 
parameter   PMA_CH3_REG_PLL_CP1_BIAS_CONTROL    = "100PCT",        //  100PCT , 111PCT , 125PCT , 143PCT , 71PCT , 77PCT , 83PCT ,91PCT
parameter   integer PMA_CH3_REG_PLL_PD_LOOP_CP1_CURRENT_SETTING    = 0,        // 0 to 31 
parameter   PMA_CH3_REG_PLL_CP0_CURRENT_SETTING    = "100PCT",        //  100PCT , 20PCT , 140PCT , 60PCT , 160PCT , 80PCT , 200PCT ,120PCT
parameter   PMA_CH3_REG_PLL_CP1_CURRENT_SETTING    = "100PCT",        //  100PCT , 20PCT , 140PCT , 60PCT , 160PCT , 80PCT , 200PCT ,120PCT
parameter   PMA_CH3_REG_PLL_GM1_CURRENT_SETTING    = "100PCT",        //  100PCT , 67PCT , 167PCT , 133PCT , 300PCT , 267PCT , 367PCT ,333PCT
parameter   PMA_CH3_REG_PLL_LC_BF2_CURRENT_SETTING    = "100PCT",        //  100PCT , 20PCT , 140PCT , 60PCT , 160PCT , 80PCT , 200PCT ,120PCT
parameter   PMA_CH3_REG_PLL_LC_BF2_CURRENT_SETTING_LOW    = "100PCT",        //  100PCT , 20PCT , 140PCT , 60PCT , 160PCT , 80PCT , 200PCT ,120PCT
parameter   PMA_CH3_REG_PLL_REG_CUR    = "100PCT",        //  100PCT , 80PCT , 140PCT , 120PCT , 180PCT , 160PCT , 220PCT ,200PCT
parameter   PMA_CH3_REG_PLL_LCCUR    = "DEFAULT",        //  DEFAULT , MINUS_1MA , 2MA , 1MA , 4MA , 3MA , 6MA ,5MA
parameter   PMA_CH3_REG_PLL_LCOBAS    = "100PCT",        // 100PCT , 75PCT , 150PCT , 125PCT 
parameter   PMA_CH3_REG_PLL_FB_CK_TEST_OUT_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   integer PMA_CH3_CDR_ALIGN_TIMER    = 0,        // 0 to 3
parameter   integer PMA_CH3_CALIB_WAIT    = 1024,        // 1024 , 2048 , 4096 , 512 
parameter   integer PMA_CH3_CALIB_TIMER    = 512,        // 512 , 1024 , 2048 , 4096 
parameter   integer PMA_CH3_TOT_RANGE    = 0,        // 0 to 3
parameter   integer PMA_CH3_SUB_RANGE    = 0,        // 0 to 3
parameter   integer PMA_CH3_OVLP    = 0,        // 0 to 3
parameter   integer PMA_CH3_BIST_WAIT    = 1024,        // 1024 , 2048 , 4096 , 512 
parameter   integer PMA_CH3_BIST_TIMER    = 512,        // 512 , 1024 , 2048 , 4096 
parameter   integer PMA_CH3_BAND_LB    = 0,        // 0 to 7 
parameter   integer PMA_CH3_BAND_HB    = 0,        // 0 to 31 
parameter   integer PMA_CH3_FREQ_LOCK_ACCURACY    = 0,        // 0 to 7
parameter   integer PMA_CH3_REG_SET_LC_BAND    = 0,        // 0 to 31 
parameter   integer PMA_CH3_REG_SET_VCODIV    = 0,        // 0 to 3
parameter   PMA_CH3_REGISTER_SET_VCODIV_BAND_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH3_REG_SET_PLL_LOCK    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH3_REGISTER_SET_PLL_LOCK_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH3_REG_SET_VCO_HI    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH3_REG_SET_VCO_LO    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH3_REGISTER_SET_VCO_HI_VCO_LO_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH3_FORCE_LC_PLL_LOOP_EN_H    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH3_FORCE_LC_PLL_LOOP_EN_L    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH3_VCO_DIV_CALI_BYPASS    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH3_BIST_EN    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH3_PLL_LOOP_EN_SETTING_FROM_REGISTER_ENABLE     = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH3_FREQ_DETECT_ENABLE_SOURCE     = "DISABLE",    // DISABLE , ENABLE
parameter   integer PMA_CH3_REG_SET_DIVSEL_REF    = 0,        // 0 to 3
parameter   PMA_CH3_REG_SET_DIVSEL45_FB    = "FALSE",    // TRUE , FALSE
parameter   integer PMA_CH3_REG_SET_DIVSEL_FB    = 0,        // 0 to 7  
parameter   PMA_CH3_PLL_LOOP_EN_SETTING     = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH3_REGISTER_SET_TXPLL_DIV_ENABLE     = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH3_FORCE_RXPLL_RESET    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH3_FORCE_RXPLL_ON    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH3_DPCK_DIV2    = "FALSE",    // TRUE , FALSE
parameter   integer PMA_CH3_LFO_SETTING    = 0,        // 0 to 7
parameter   PMA_CH3_ALOS_COUNTER_CLOCK_SELECTION    = "LOCAL",    // LOCAL , GLOBAL25M
parameter   PMA_CH3_RX_BIAS_CURRENT_ADJUSTMENT    = "100PCT",        //  100PCT , 111PCT , 125PCT , 143PCT , 71PCT , 77PCT , 83PCT ,91PCT
parameter   integer PMA_CH3_OOB_ENTER_DELAY_SETTING    = 0,        // 0 to 3
parameter   integer PMA_CH3_ALOS_LOW_TO_HIGH_COUNTER_SETTING    = 0,        // 0 to 3
parameter   PMA_CH3_ENABLE_ALOS_RESULT_AUTOMATICALLY_ENABLE_CHANNEL     = "DISABLE",    // DISABLE , ENABLE
parameter   integer PMA_CH3_ALOS_EXIT_COUNTER_CLOCK_DIVIDER    = 0,        // 0 to 3
parameter   integer PMA_CH3_OOB_OSCILATER_FREQUENCY_SETTING    = 0,        // 0 to 3
parameter   PMA_CH3_FORCE_OOB    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH3_OOB_VTH_SET    = "27MV",        // 27MV, 30MV, 35MV, 42_5MV, 52MV, 68MV 
parameter   PMA_CH3_FORCE_DET_FORCE_ALOS_LOW    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH3_ALOS_THRESHOLD_VOLTAGE    = "27MV",        // 27MV, 30MV, 35MV, 42_5MV, 52MV, 68MV 
parameter   integer PMA_CH3_WAKEUP_VCM_RX_COMMON_MODE_VOLTAGE    = 0,        // 0 to 3
parameter   PMA_CH3_REGR_NEGATIVE_HYSTERESIS_SETTING    = "100MV",        // 100MV, 75MV, 50MV, 25MV, 25MV, 0MV 
parameter   PMA_CH3_REGL_POSITIVE_HYSTERESIS_SETTING    = "100MV",        // 100MV, 75MV, 50MV, 25MV, 25MV, 0MV 
parameter   PMA_CH3_REG_EN    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH3_REGREF_SEL    = "VREF",    // VREF , SELF_DC
parameter   PMA_CH3_DC496    = "39_6MHZ",        // 5MHZ, 8MHZ, 11_5MHZ, 20_6MHZ, 39_6MHZ 
parameter   integer PMA_CH3_EQ2_AC_VAR_SETTING    = 0,        // 255,254,252,248,240,224,192,128,0
parameter   integer PMA_CH3_EQ2_AC_RES_SETTING    = 0,        // 0 to 31 
parameter   integer PMA_CH3_EQ2_DC_RESTOP_SETTING    = 0,        // 0 to 3
parameter   integer PMA_CH3_EQ1_DC_RESTOP_SETTING    = 50,        //  50, 60, 71, 78, 107 
parameter   integer PMA_CH3_EQ1_AC_VAR_SETTING    = 0,        // 255,254,252,248,240,224,192,128,0
parameter   integer PMA_CH3_EQ2_CURRENT_SETTING    = 0,        // 0,1,3,7
parameter   integer PMA_CH3_EQ1_AC_RES_SETTING    = 0,        // 0 to 31 
parameter   integer PMA_CH3_EQ1_CURRENT_SETTING    = 0,        // 15,7,3,9,1,0 
parameter   integer PMA_CH3_RPLUS    = 0,        // 0,1,3,7,15
parameter   integer PMA_CH3_RMINUS    = 0,        // 0,1,3,7,15
parameter   integer PMA_CH3_RVALSET    = 0,        // 0 to 3
parameter   integer PMA_CH3_RTERM    = 0,        // 0 to 3
parameter   PMA_CH3_DCFB_EN    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_CH3_DCCOUP    = "FALSE",    // TRUE , FALSE
parameter   PMA_CH3_3G    = "FALSE",    // TRUE , FALSE

parameter   PMA_QUAD_TURN_ON_BANDGAP_AT_AOS_ON    = "FALSE",    // TRUE , FALSE
parameter   PMA_QUAD_TURN_ON_BANDGAP_AT_RX_DETECTION_ON    = "FALSE",    // TRUE , FALSE
parameter   PMA_QUAD_TURN_ON_BANDGAP_AT_BOUNDARY_SCAN_ON    = "FALSE",    // TRUE , FALSE
parameter   PMA_QUAD_CFG_HSST_RSTN    = "FALSE",    // TRUE , FALSE
parameter   PMA_QUAD_SELECT_LANE_TCK_FOR_QUAD_SYNC    = "LANE0",        // LANE0,LANE1,LANE2,LANE3 
parameter   PMA_QUAD_CK_REN    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_QUAD_C1_EN    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_QUAD_C2_EN    = "DISABLE",    // DISABLE , ENABLE
parameter   integer PMA_QUAD_CLK_DIVIDER_SETTING_FROM_25M_TO_200K    = 0,        // 0 to 3 
parameter   PMA_QUAD_ACMODE_SCANMODE_EN    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_QUAD_REGISTER_ACMODE    = "FALSE",    // TRUE , FALSE
parameter   PMA_QUAD_REGISTER_SCANMODE    = "FALSE",    // TRUE , FALSE
parameter   PMA_QUAD_REFCK2CORE_EN    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_QUAD_REG_EN    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_QUAD_REGR    = "100MV",        // 100MV, 75MV, 50MV, 25MV, 0MV
parameter   PMA_QUAD_REGL    = "100MV",        // 100MV, 75MV, 50MV, 25MV, 0MV
parameter   integer PMA_QUAD_DPCK_SEL    = 0,        // 0 to 3
parameter   PMA_QUAD_TX_REFCK_SEL    = "FALSE",    // TRUE , FALSE
parameter   PMA_QUAD_REFCK_SRC_SEL    = "FALSE",    // TRUE , FALSE
parameter   PMA_QUAD_RREFCK_PWRUP    = "FALSE",    // TRUE , FALSE
parameter   PMA_QUAD_REFCK_SK_SEL       = "BOTH",    // BOTH, UP, DOWN, NONE
parameter   PMA_QUAD_REFCK_DIV2_SEL    = "FALSE",    // TRUE , FALSE
parameter   PMA_QUAD_REFCK_TO_NQ_EN    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_QUAD_AUXI_ADJ    = "100PCT",        //  100PCT , 111PCT , 125PCT , 143PCT , 71PCT , 77PCT , 83PCT ,91PCT
parameter   PMA_QUAD_DC496    = "39_6MHZ",        // 5MHZ, 8MHZ, 11_5MHZ, 20_6MHZ, 39_6MHZ 
parameter   integer PMA_QUAD_REG_FDET_TIMER    = 512,        // 256, 512 , 1024 , 2048 
parameter   PMA_QUAD_FREQ_LKO    = "10PCT",    // 1PCT , 2PCT , 5PCT , 10PCT
parameter   PMA_QUAD_FREQ_LKI    = "10PCT",    // 1PCT , 2PCT , 5PCT , 10PCT
parameter   PMA_QUAD_CLOCK_SRC_SEL    = "LOCAL",    // LOCAL, NEIGHBOR 
parameter   PMA_QUAD_FRE_DET_EN    = "DISABLE",    // DISABLE , ENABLE
parameter   integer PMA_QUAD_TSO_LS_SEL    = 0,        // 0 to 127 
parameter   PMA_QUAD_TXPLL_START    = "FALSE",    // TRUE , FALSE
parameter   integer PMA_QUAD_VCODIV    = 0,        // 0 to 3
parameter   integer PMA_QUAD_LC_BAND    = 0,        // 0 to 31 
parameter   PMA_QUAD_SET_VCO_HI    = "FALSE",    // TRUE , FALSE
parameter   PMA_QUAD_SET_VCO_LO    = "FALSE",    // TRUE , FALSE
parameter   PMA_QUAD_CALIB_FAIL    = "FALSE",    // TRUE , FALSE
parameter   PMA_QUAD_CALIB_DONE    = "FALSE",    // TRUE , FALSE
parameter   PMA_QUAD_BIST_DONE    = "FALSE",    // TRUE , FALSE
parameter   PMA_QUAD_TOTRANGE_FAIL    = "FALSE",    // TRUE , FALSE
parameter   PMA_QUAD_SUBRANGE_FAIL    = "FALSE",    // TRUE , FALSE
parameter   PMA_QUAD_OVLP_FAIL    = "FALSE",    // TRUE , FALSE
parameter   PMA_QUAD_TXPLL_LOCK    = "FALSE",    // TRUE , FALSE
parameter   PMA_QUAD_TXPLL_LOOP_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   integer PMA_QUAD_TXPLL_DIVSEL_REF_STA    = 0,        // 0 to 3
parameter   PMA_QUAD_TXPLL_DIVSEL45_FB_STA    = "FALSE",    // TRUE , FALSE
parameter   integer PMA_QUAD_TXPLL_DIVSEL_FB_STA    = 0,        // 0 to 7 
parameter   PMA_QUAD_TXPLL_DIVSEL45_FB    = "FALSE",    // TRUE , FALSE
parameter   integer PMA_QUAD_TXPLL_DIVSEL_FB    = 0,        // 0 to 7 
parameter   integer PMA_QUAD_TXPLL_DIVSEL_REF    = 0,        // 0 to 3
parameter   PMA_QUAD_REG_DISABLE_HOLDCLK    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_QUAD_REG_DISABLE_SYNC    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_QUAD_FORCE_OUTPUT_PLL_LOCK    = "FALSE",    // TRUE , FALSE
parameter   PMA_QUAD_REGISTER_SET_SYNCTCK_SEL_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_QUAD_REG_SET_SYNCTCK_SEL    = "LANE0",        // LANE0,LANE1,LANE2,LANE3 
parameter   PMA_QUAD_CK4TEST_OUTPUT_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_QUAD_RSTGENBAS    = "100PCT",    // 100PCT , 83PCT , 133PCT , 117PCT
parameter   PMA_QUAD_LCBUFBAS    = "100PCT",    // 100PCT , 83PCT , 133PCT , 117PCT
parameter   PMA_QUAD_REGISTER_SET_CPCUR_ENABEL    = "DISABLE",    // DISABLE , ENABLE
parameter   integer PMA_QUAD_REG_SET_CPCUR    = 0,        // 0 to 31 
parameter   PMA_QUAD_CPBAS    = "100PCT",        //  100PCT , 111PCT , 125PCT , 143PCT , 71PCT , 77PCT , 83PCT ,91PCT
parameter   PMA_QUAD_LCOBAS    = "100PCT",    // 100PCT , 75PCT , 150PCT , 125PCT
parameter   PMA_QUAD_LCCUR    = "DEFAULT",        //  DEFAULT , _1MA , 2MA , 1MA , 4MA , 3MA , 6MA ,5MA
parameter   PMA_QUAD_ENABLE_REGISTER_SETTING_BAND    = "DISABLE",    // DISABLE , ENABLE
parameter   integer PMA_QUAD_CALIB_WAIT    = 1024,        // 1024 , 2048 , 4096 , 512 
parameter   integer PMA_QUAD_CALIB_TIMER    = 512,        // 512 , 1024 , 2048 , 4096 
parameter   integer PMA_QUAD_TOT_RANGE    = 0,        // 0 to 3
parameter   integer PMA_QUAD_SUB_RANGE    = 0,        // 0 to 3
parameter   integer PMA_QUAD_OVLP    = 0,        // 0 to 3
parameter   integer PMA_QUAD_BIST_WAIT    = 1024,        // 1024 , 2048 , 4096 , 512 
parameter   integer PMA_QUAD_BIST_TIMER    = 512,        // 512 , 1024 , 2048 , 4096 
parameter   integer PMA_QUAD_BAND_LB    = 0,        // 0 to 7 
parameter   integer PMA_QUAD_BAND_HB    = 0,        // 0 to 31 
parameter   integer PMA_QUAD_FREQ_LOCK_ACCURACY    = 0,        //  0 to 7
parameter   integer PMA_QUAD_REG_SET_LC_BAND    = 0,        // 0 to 31 
parameter   integer PMA_QUAD_REG_SET_VCODIV    = 0,        // 0 to 3
parameter   PMA_QUAD_REGISTER_SET_VCODIV_BAND_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_QUAD_REG_SET_PLL_LOCK    = "FALSE",    // TRUE , FALSE
parameter   PMA_QUAD_REGISTER_SET_PLL_LOCK_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_QUAD_REG_SET_VCO_HI    = "FALSE",    // TRUE , FALSE
parameter   PMA_QUAD_REG_SET_VCO_LO    = "FALSE",    // TRUE , FALSE
parameter   PMA_QUAD_REGISTER_SET_VCO_HI_VCO_LO_ENABLE    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_QUAD_FORCE_LC_PLL_LOOP_EN_H    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_QUAD_FORCE_LC_PLL_LOOP_EN_L    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_QUAD_VCO_DIV_CALI_BYPASS    = "FALSE",    // TRUE , FALSE
parameter   PMA_QUAD_BIST_EN    = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_QUAD_ENABLE_TXPLL_BIST_BLOCK_CLOCKS     = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_QUAD_LF_TESTBY2     = "DISABLE",    // DISABLE , ENABLE
parameter   integer PMA_QUAD_REG_SET_DIVSEL_REF    = 0,        // 0 to 3
parameter   PMA_QUAD_REG_SET_DIVSEL45_FB    = "FALSE",    // TRUE , FALSE
parameter   integer PMA_QUAD_REG_SET_DIVSEL_FB    = 0,        // 0 to 7  
parameter   PMA_QUAD_LF_TEST_EN     = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_QUAD_REGISTER_SET_TXPLL_DIV_ENABLE     = "DISABLE",    // DISABLE , ENABLE
parameter   PMA_QUAD_FORCE_TXPLL_RESET    = "FALSE",    // TRUE , FALSE
parameter   PMA_QUAD_FORCE_TXPLL_ON    = "FALSE",    // TRUE , FALSE



parameter integer  CLK_ALIGNER_RX0    = 0,        // 
parameter integer  CLK_ALIGNER_RX1    = 0,        // 
parameter integer  CLK_ALIGNER_RX2    = 0,        // 
parameter integer  CLK_ALIGNER_RX3    = 0,        // 
parameter integer  CLK_ALIGNER_TX0    = 0,        // 
parameter integer  CLK_ALIGNER_TX1    = 0,        // 
parameter integer  CLK_ALIGNER_TX2    = 0,        // 
parameter integer  CLK_ALIGNER_TX3    = 0,        // 
parameter          DYN_DLY_EN_RX0    = "FALSE",        // 
parameter          DYN_DLY_EN_RX1    = "FALSE",        // 
parameter          DYN_DLY_EN_RX2    = "FALSE",        // 
parameter          DYN_DLY_EN_RX3    = "FALSE",        // 
parameter          DYN_DLY_EN_TX0    = "FALSE",        // 
parameter          DYN_DLY_EN_TX1    = "FALSE",        // 
parameter          DYN_DLY_EN_TX2    = "FALSE",        // 
parameter          DYN_DLY_EN_TX3    = "FALSE",        // 
parameter          DYN_DLY_SEL_RX0    = "FALSE",        // 
parameter          DYN_DLY_SEL_RX1    = "FALSE",        // 
parameter          DYN_DLY_SEL_RX2    = "FALSE",        // 
parameter          DYN_DLY_SEL_RX3    = "FALSE",        // 
parameter          DYN_DLY_SEL_TX0    = "FALSE",        // 
parameter          DYN_DLY_SEL_TX1    = "FALSE",        // 
parameter          DYN_DLY_SEL_TX2    = "FALSE",        // 
parameter          DYN_DLY_SEL_TX3    = "FALSE",        // 
parameter integer  CLK_ALIGNER_RSTN_RX    = 0,        // 
parameter integer  CLK_ALIGNER_RSTN_TX    = 0,        // 
parameter integer  LX_BISTLB_EN    = 0,        // 
parameter integer  LX_ELECIDLE_EN_MSB    = 0,        // 
parameter integer  LX_EXTLB_EN    = 0,        // 
parameter integer  LX_RXDCT_EN    = 0,        // 
parameter integer  LX_TX_LFMODE    = 0,        // 
parameter integer  RX_LANE_POWERUP    = 0,        // 
parameter integer  TX_LANE_POWERUP    = 0,        // 
parameter          PLL_RSTN    = "FALSE",        // 
parameter          PLLPOWERDOWN    = "FALSE",        // 
parameter          QUAD_PWRUP    = "FALSE",        // 
parameter          GRSN_DIS    = "FALSE",        // 
parameter          HSST_RSTN    = "FALSE",        // 
parameter          CFG_RSTN    = "FALSE"        // 





 )


(


 output         P_AFTER_CTC_RCLK_EN_COUT    ,
 output         P_AFTER_CTC_RCLK_EN_GB_COUT    ,
 output         P_APATTERN_MATCH_LSB_COUT    ,
 output         P_APATTERN_MATCH_MSB_COUT    ,
 output         P_APATTERN_SEACHING_PROC_COUT    ,
 output         P_APATTERN_STATUS_COUT    ,
 output         P_BRIDGE_RCLK_EN_COUT    ,
 output         P_BRIDGE_TCLK_EN_COUT    ,
 output         P_CB_RCLK_EN_COUT    ,
 output         P_CFG_INT    ,
 output         P_CFG_READY    ,
 output         P_CTC_RD_FIFO_COUT    ,
 output         P_L0TXN    ,
 output         P_L0TXP    ,
 output         P_L1TXN    ,
 output         P_L1TXP    ,
 output         P_L2TXN    ,
 output         P_L2TXP    ,
 output         P_L3TXN    ,
 output         P_L3TXP    ,
 output         P_LX_ALOS_STA_0    ,
 output         P_LX_ALOS_STA_1    ,
 output         P_LX_ALOS_STA_2    ,
 output         P_LX_ALOS_STA_3    ,
 output         P_LX_CDR_ALIGN_0    ,
 output         P_LX_CDR_ALIGN_1    ,
 output         P_LX_CDR_ALIGN_2    ,
 output         P_LX_CDR_ALIGN_3    ,
 output         P_LX_LFO_0    ,
 output         P_LX_LFO_1    ,
 output         P_LX_LFO_2    ,
 output         P_LX_LFO_3    ,
 output         P_LX_OOB_STA_0    ,
 output         P_LX_OOB_STA_1    ,
 output         P_LX_OOB_STA_2    ,
 output         P_LX_OOB_STA_3    ,
 output         P_LX_RXDCT_DONE_0    ,
 output         P_LX_RXDCT_DONE_1    ,
 output         P_LX_RXDCT_DONE_2    ,
 output         P_LX_RXDCT_DONE_3    ,
 output         P_LX_RXDCT_OUT_0    ,
 output         P_LX_RXDCT_OUT_1    ,
 output         P_LX_RXDCT_OUT_2    ,
 output         P_LX_RXDCT_OUT_3    ,
 output         P_PCS_TCLK_EN_COUT    ,
 output         P_PLL_LOCK    ,
 output         P_REFCK2CORE    ,
 output         P_REFCK_2NMQ    ,
 output         P_REFCK_2NPQ    ,
 output         P_REXT    ,
 output         P_RFIFO_EN_AFTER_CTC_COUT    ,
 output         P_RFIFO_EN_AFTER_CTC_GB_COUT    ,
 output         P_RFIFO_EN_BRIDGE_COUT    ,
 output         P_RFIFO_EN_CB_COUT    ,
 output         P_SKIP_ADD_LSB_MCB_COUT    ,
 output         P_SKIP_ADD_MCB_COUT    ,
 output         P_SKIP_DEL_LSB_MCB_COUT    ,
 output         P_SKIP_DEL_MCB_COUT    ,
 output         P_TFIFO_EN_BRIDGE_COUT    ,
 output         P_TFIFO_EN_PCS_TX_COUT    ,
 output         P_TSO_LS_OUT    ,





 input         P_AFTER_CTC_RCLK_EN_CIN    ,
 input         P_AFTER_CTC_RCLK_EN_GB_CIN    ,
 input         P_APATTERN_MATCH_LSB_CIN    ,
 input         P_APATTERN_MATCH_MSB_CIN    ,
 input         P_APATTERN_SEACHING_PROC_CIN    ,
 input         P_APATTERN_STATUS_CIN    ,
 input         P_BRIDGE_RCLK_EN_CIN    ,
 input         P_BRIDGE_TCLK_EN_CIN    ,
 input         P_CB_RCLK_EN_CIN    ,
 input         P_CFG_CLK    ,
 input         P_CFG_ENABLE    ,
 input         P_CFG_RSTN    ,
 input         P_CFG_WRITE    ,
 input         P_COMPRESSION_MODE    ,
 input         P_CTC_RD_FIFO_CIN    ,
 input         P_HSST_RSTN    ,
 input         P_L0RXN    ,
 input         P_L0RXP    ,
 input         P_L1RXN    ,
 input         P_L1RXP    ,
 input         P_L2RXN    ,
 input         P_L2RXP    ,
 input         P_L3RXN    ,
 input         P_L3RXP    ,
 input         P_LANE_SYNC_EN_0    ,
 input         P_LANE_SYNC_EN_1    ,
 input         P_LANE_SYNC_EN_2    ,
 input         P_LANE_SYNC_EN_3    ,
 input         P_LX_LFD_FRCORE_0    ,
 input         P_LX_LFD_FRCORE_1    ,
 input         P_LX_LFD_FRCORE_2    ,
 input         P_LX_LFD_FRCORE_3    ,
 input         P_LX_RX_CKDIV_DYNSEL_0    ,
 input         P_LX_RX_CKDIV_DYNSEL_1    ,
 input         P_LX_RX_CKDIV_DYNSEL_2    ,
 input         P_LX_RX_CKDIV_DYNSEL_3    ,
 input         P_MCB_CLK_FRNQ    ,
 input         P_PCS_RX_RSTN_0    ,
 input         P_PCS_RX_RSTN_1    ,
 input         P_PCS_RX_RSTN_2    ,
 input         P_PCS_RX_RSTN_3    ,
 input         P_PCS_TCLK_EN_CIN    ,
 input         P_PCS_TX_RSTN_0    ,
 input         P_PCS_TX_RSTN_1    ,
 input         P_PCS_TX_RSTN_2    ,
 input         P_PCS_TX_RSTN_3    ,
 input         P_PLL_BYPASS    ,
 input         P_PLL_REF_CLK    ,
 input         P_PLL_RESET    ,
 input         P_PLL_RSTN    ,
 input         P_PLLPOWERDOWN    ,
 input         P_QUAD_PWRUP    ,
 input         P_REFCK_FRNMQ    ,
 input         P_REFCK_FRNPQ    ,
 input         P_REFCKN    ,
 input         P_REFCKP    ,
 input         P_RFIFO_EN_AFTER_CTC_CIN    ,
 input         P_RFIFO_EN_AFTER_CTC_GB_CIN    ,
 input         P_RFIFO_EN_BRIDGE_CIN    ,
 input         P_RFIFO_EN_CB_CIN    ,
 input         P_RX0_CLK_FR_CORE    ,
 input         P_RX1_CLK_FR_CORE    ,
 input         P_RX2_CLK_FR_CORE    ,
 input         P_RX3_CLK_FR_CORE    ,
 input         P_RX_PLL_RSTN_0    ,
 input         P_RX_PLL_RSTN_1    ,
 input         P_RX_PLL_RSTN_2    ,
 input         P_RX_PLL_RSTN_3    ,
 input         P_RX_PMA_RSTN_0    ,
 input         P_RX_PMA_RSTN_1    ,
 input         P_RX_PMA_RSTN_2    ,
 input         P_RX_PMA_RSTN_3    ,
 input         P_RX_REF_CLK_0    ,
 input         P_RX_REF_CLK_1    ,
 input         P_RX_REF_CLK_2    ,
 input         P_RX_REF_CLK_3    ,
 input         P_SEL_SYNC_NXQ    ,
 input         P_SKIP_ADD_LSB_MCB_CIN    ,
 input         P_SKIP_ADD_MCB_CIN    ,
 input         P_SKIP_DEL_LSB_MCB_CIN    ,
 input         P_SKIP_DEL_MCB_CIN    ,
 input         P_SYNC_TOGGLE    ,
 input         P_TFIFO_EN_BRIDGE_CIN    ,
 input         P_TFIFO_EN_PCS_TX_CIN    ,
 input         P_TWOQUAD_SYNC_EN    ,
 input         P_TX0_CLK_FR_CORE    ,
 input         P_TX1_CLK_FR_CORE    ,
 input         P_TX2_CLK_FR_CORE    ,
 input         P_TX3_CLK_FR_CORE    ,
 input         P_TX_PMA_RSTN_0    ,
 input         P_TX_PMA_RSTN_1    ,
 input         P_TX_PMA_RSTN_2    ,
 input         P_TX_PMA_RSTN_3    ,
 input         P_TXCKDIV_DYNSEL    ,



output [46:0]  P_RDATA_0,
output [46:0]  P_RDATA_1,
output [3:0]  P_PCS_LSM_SYNCED,
output [46:0]  P_RDATA_2,
output [3:0]  P_ALIGN_TX,
output [3:0]  P_ALIGN_RX,
output [46:0]  P_RDATA_3,
output [3:0]  P_CLK2CORE_TX,
output [3:0]  P_CLK2CORE_RX,
output [7:0]  P_CFG_RDATA,
output [3:0]  P_PCS_RX_MCB_STATUS,
input [7:0]  P_CIM_CLK_ALIGNER_TX3,
input [1:0]  P_TX_CKDIV_1,
input [2:0]  P_LX_DEEMP_CTL_1,
input [3:0]  P_LX_TX_LFMODE,
input [3:0]  P_LX_AMP_CTL_0,
input [3:0]  P_LX_RXDCT_EN,
input [1:0]  P_TX_CKDIV_0,
input [1:0]  P_LX_RX_CKDIV_3,
input [3:0]  P_PCS_MCB_EXT_EN,
input [7:0]  P_CIM_CLK_ALIGNER_TX0,
input [2:0]  P_LX_DEEMP_CTL_0,
input [43:0]  P_TDATA_2,
input [3:0]  P_LX_AMP_CTL_3,
input [7:0]  P_CIM_CLK_ALIGNER_TX1,
input [1:0]  P_LX_RX_CKDIV_2,
input [3:0]  P_CEB_ADETECT_EN,
input [1:0]  P_TX_CKDIV_3,
input [7:0]  P_CIM_CLK_ALIGNER_RX1,
input [7:0]  P_CFG_WDATA,
input [3:0]  P_TX_LANE_POWERUP,
input [43:0]  P_TDATA_1,
input [3:0]  P_LX_EXTLB_EN,
input [15:0]  P_CFG_ADDR,
input [7:0]  P_CIM_CLK_ALIGNER_RX0,
input [3:0]  P_LX_ELECIDLE_EN_MSB,
input [3:0]  P_PCS_NEAREND_LOOP,
input [1:0]  P_LX_ELECIDLE_EN_0,
input [1:0]  P_LX_ELECIDLE_EN_3,
input [3:0]  P_CIM_CLK_DYN_DLY_SEL_RX,
input [2:0]  P_LX_DEEMP_CTL_3,
input [1:0]  P_LX_ELECIDLE_EN_1,
input [3:0]  P_CIM_CLK_START_ALIGN_TX,
input [3:0]  P_LX_BISTLB_EN,
input [43:0]  P_TDATA_0,
input [7:0]  P_CIM_CLK_ALIGNER_RX3,
input [3:0]  P_CIM_CLK_DYN_DLY_SEL_TX,
input [7:0]  P_CIM_CLK_ALIGNER_TX2,
input [1:0]  P_LX_ELECIDLE_EN_2,
input [3:0]  P_RX_LANE_POWERUP,
input [1:0]  P_TX_CKDIV_2,
input [3:0]  P_PCS_WORD_ALIGN_EN,
input [3:0]  P_LX_AMP_CTL_1,
input [7:0]  P_CIM_CLK_ALIGNER_RX2,
input [3:0]  P_RX_POLARITY_INVERT,
input [2:0]  P_LX_DEEMP_CTL_2,
input [3:0]  P_LX_AMP_CTL_2,
input [1:0]  P_LX_RX_CKDIV_1,
input [43:0]  P_TDATA_3,
input [3:0]  P_PCS_FAREND_LOOP,
input [3:0]  P_CIM_CLK_START_ALIGN_RX,
input [1:0]  P_LX_RX_CKDIV_0


);

supply0 REP0;
supply1 REP1;
reg P_CK25M;
initial begin 
        P_CK25M=0; 
        forever #20 P_CK25M = ~P_CK25M;
        end

hsst_gtp_wrap 
#(

 .PCS_CH0_BYPASS_WORD_ALIGN(PCS_CH0_BYPASS_WORD_ALIGN), 
 .PCS_CH0_BYPASS_DENC(PCS_CH0_BYPASS_DENC), 
 .PCS_CH0_BYPASS_BONDING(PCS_CH0_BYPASS_BONDING), 
 .PCS_CH0_BYPASS_CTC(PCS_CH0_BYPASS_CTC), 
 .PCS_CH0_BYPASS_GEAR(PCS_CH0_BYPASS_GEAR), 
 .PCS_CH0_BYPASS_BRIDGE(PCS_CH0_BYPASS_BRIDGE), 
 .PCS_CH0_DATA_MODE(PCS_CH0_DATA_MODE), 
 .PCS_CH0_RX_POLARITY_INV(PCS_CH0_RX_POLARITY_INV), 
 .PCS_CH0_ALIGN_MODE(PCS_CH0_ALIGN_MODE), 
 .PCS_CH0_SAMP_16B(PCS_CH0_SAMP_16B), 
 .PCS_CH0_COMMA_REG0(PCS_CH0_COMMA_REG0), 
 .PCS_CH0_COMMA_MASK(PCS_CH0_COMMA_MASK), 
 .PCS_CH0_CEB_MODE(PCS_CH0_CEB_MODE), 
 .PCS_CH0_CTC_MODE(PCS_CH0_CTC_MODE), 
 .PCS_CH0_A_REG(PCS_CH0_A_REG), 
 .PCS_CH0_GE_AUTO_EN(PCS_CH0_GE_AUTO_EN), 
 .PCS_CH0_SKIP_REG0(PCS_CH0_SKIP_REG0), 
 .PCS_CH0_SKIP_REG1(PCS_CH0_SKIP_REG1), 
 .PCS_CH0_SKIP_REG2(PCS_CH0_SKIP_REG2), 
 .PCS_CH0_SKIP_REG3(PCS_CH0_SKIP_REG3), 
 .PCS_CH0_DEC_DUAL(PCS_CH0_DEC_DUAL), 
 .PCS_CH0_SPLIT(PCS_CH0_SPLIT), 
 .PCS_CH0_FIFOFLAG_CTC(PCS_CH0_FIFOFLAG_CTC), 
 .PCS_CH0_COMMA_DET_MODE(PCS_CH0_COMMA_DET_MODE), 
 .PCS_CH0_ERRDETECT_SILENCE(PCS_CH0_ERRDETECT_SILENCE), 
 .PCS_CH0_PMA_RCLK_POLINV(PCS_CH0_PMA_RCLK_POLINV), 
 .PCS_CH0_PCS_RCLK_SEL(PCS_CH0_PCS_RCLK_SEL), 
 .PCS_CH0_MCB_RCLK_POLINV(PCS_CH0_MCB_RCLK_POLINV), 
 .PCS_CH0_CB_RCLK_SEL(PCS_CH0_CB_RCLK_SEL), 
 .PCS_CH0_AFTER_CTC_RCLK_SEL(PCS_CH0_AFTER_CTC_RCLK_SEL), 
 .PCS_CH0_RCLK_POLINV(PCS_CH0_RCLK_POLINV), 
 .PCS_CH0_BRIDGE_RCLK_SEL(PCS_CH0_BRIDGE_RCLK_SEL), 
 .PCS_CH0_PCS_RCLK_EN(PCS_CH0_PCS_RCLK_EN), 
 .PCS_CH0_CB_RCLK_EN(PCS_CH0_CB_RCLK_EN), 
 .PCS_CH0_AFTER_CTC_RCLK_EN(PCS_CH0_AFTER_CTC_RCLK_EN), 
 .PCS_CH0_AFTER_CTC_RCLK_EN_GB(PCS_CH0_AFTER_CTC_RCLK_EN_GB), 
 .PCS_CH0_BRIDGE_RCLK_EN(PCS_CH0_BRIDGE_RCLK_EN), 
 .PCS_CH0_PCS_RX_RSTN(PCS_CH0_PCS_RX_RSTN), 
 .PCS_CH0_SLAVE(PCS_CH0_SLAVE), 
 .PCS_CH0_PCIE_SLAVE(PCS_CH0_PCIE_SLAVE), 
 .PCS_CH0_PCS_CB_RSTN(PCS_CH0_PCS_CB_RSTN), 
 .PCS_CH0_TX_BYPASS_BRIDGE_UINT(PCS_CH0_TX_BYPASS_BRIDGE_UINT), 
 .PCS_CH0_TX_BYPASS_GEAR(PCS_CH0_TX_BYPASS_GEAR), 
 .PCS_CH0_TX_BYPASS_ENC(PCS_CH0_TX_BYPASS_ENC), 
 .PCS_CH0_TX_BYPASS_BIT_SLIP(PCS_CH0_TX_BYPASS_BIT_SLIP), 
 .PCS_CH0_TX_GEAR_SPLIT(PCS_CH0_TX_GEAR_SPLIT), 
 .PCS_CH0_TX_DRIVE_REG_MODE(PCS_CH0_TX_DRIVE_REG_MODE), 
 .PCS_CH0_TX_BIT_SLIP_CYCLES(PCS_CH0_TX_BIT_SLIP_CYCLES), 
 .PCS_CH0_INT_TX_MASK_0(PCS_CH0_INT_TX_MASK_0), 
 .PCS_CH0_INT_TX_MASK_1(PCS_CH0_INT_TX_MASK_1), 
 .PCS_CH0_INT_TX_MASK_2(PCS_CH0_INT_TX_MASK_2), 
 .PCS_CH0_INT_TX_CLR_0(PCS_CH0_INT_TX_CLR_0), 
 .PCS_CH0_INT_TX_CLR_1(PCS_CH0_INT_TX_CLR_1), 
 .PCS_CH0_INT_TX_CLR_2(PCS_CH0_INT_TX_CLR_2), 
 .PCS_CH0_TX_PMA_TCLK_POLINV(PCS_CH0_TX_PMA_TCLK_POLINV), 
 .PCS_CH0_TX_PCS_CLK_EN_SEL(PCS_CH0_TX_PCS_CLK_EN_SEL), 
 .PCS_CH0_TX_BRIDGE_TCLK_SEL(PCS_CH0_TX_BRIDGE_TCLK_SEL), 
 .PCS_CH0_TX_TCLK_POLINV(PCS_CH0_TX_TCLK_POLINV), 
 .PCS_CH0_TX_PCS_TX_RSTN(PCS_CH0_TX_PCS_TX_RSTN), 
 .PCS_CH0_TX_SLAVE(PCS_CH0_TX_SLAVE), 
 .PCS_CH0_TX_BRIDGE_CLK_EN_SEL(PCS_CH0_TX_BRIDGE_CLK_EN_SEL), 
 .PCS_CH0_DATA_WIDTH_MODE(PCS_CH0_DATA_WIDTH_MODE), 
 .PCS_CH0_TX_TCLK2FABRIC_SEL(PCS_CH0_TX_TCLK2FABRIC_SEL), 
 .PCS_CH0_TX_OUTZZ(PCS_CH0_TX_OUTZZ), 
 .PCS_CH0_ENC_DUAL(PCS_CH0_ENC_DUAL), 
 .PCS_CH0_TX_BITSLIP_DATA_MODE(PCS_CH0_TX_BITSLIP_DATA_MODE), 
 .PCS_CH0_COMMA_REG1(PCS_CH0_COMMA_REG1), 
 .PCS_CH0_RAPID_IMAX(PCS_CH0_RAPID_IMAX), 
 .PCS_CH0_RAPID_VMIN_1(PCS_CH0_RAPID_VMIN_1), 
 .PCS_CH0_RAPID_VMIN_2(PCS_CH0_RAPID_VMIN_2), 
 .PCS_CH0_RX_PRBS_MODE(PCS_CH0_RX_PRBS_MODE), 
 .PCS_CH0_RX_ERRCNT_CLR(PCS_CH0_RX_ERRCNT_CLR), 
 .PCS_CH0_TX_PRBS_MODE(PCS_CH0_TX_PRBS_MODE), 
 .PCS_CH0_TX_INSERT_ER(PCS_CH0_TX_INSERT_ER), 
 .PCS_CH0_ENABLE_PRBS_GEN(PCS_CH0_ENABLE_PRBS_GEN), 
 .PCS_CH0_ERR_CNT(PCS_CH0_ERR_CNT), 
 .PCS_CH0_DEFAULT_RADDR(PCS_CH0_DEFAULT_RADDR), 
 .PCS_CH0_MASTER_CHECK_OFFSET(PCS_CH0_MASTER_CHECK_OFFSET), 
 .PCS_CH0_DELAY_SET(PCS_CH0_DELAY_SET), 
 .PCS_CH0_SEACH_OFFSET(PCS_CH0_SEACH_OFFSET), 
 .PCS_CH0_CEB_RAPIDLS_MMAX(PCS_CH0_CEB_RAPIDLS_MMAX), 
 .PCS_CH0_CTC_AFULL(PCS_CH0_CTC_AFULL), 
 .PCS_CH0_CTC_AEMPTY(PCS_CH0_CTC_AEMPTY), 
 .PCS_CH0_FAR_LOOP(PCS_CH0_FAR_LOOP), 
 .PCS_CH0_NEAR_LOOP(PCS_CH0_NEAR_LOOP), 
 .PCS_CH0_INT_RX_MASK_0(PCS_CH0_INT_RX_MASK_0), 
 .PCS_CH0_INT_RX_MASK_1(PCS_CH0_INT_RX_MASK_1), 
 .PCS_CH0_INT_RX_MASK_2(PCS_CH0_INT_RX_MASK_2), 
 .PCS_CH0_INT_RX_MASK_3(PCS_CH0_INT_RX_MASK_3), 
 .PCS_CH0_INT_RX_MASK_4(PCS_CH0_INT_RX_MASK_4), 
 .PCS_CH0_INT_RX_MASK_5(PCS_CH0_INT_RX_MASK_5), 
 .PCS_CH0_INT_RX_MASK_6(PCS_CH0_INT_RX_MASK_6), 
 .PCS_CH0_INT_RX_MASK_7(PCS_CH0_INT_RX_MASK_7), 
 .PCS_CH0_INT_RX_CLR_0(PCS_CH0_INT_RX_CLR_0), 
 .PCS_CH0_INT_RX_CLR_1(PCS_CH0_INT_RX_CLR_1), 
 .PCS_CH0_INT_RX_CLR_2(PCS_CH0_INT_RX_CLR_2), 
 .PCS_CH0_INT_RX_CLR_3(PCS_CH0_INT_RX_CLR_3), 
 .PCS_CH0_INT_RX_CLR_4(PCS_CH0_INT_RX_CLR_4), 
 .PCS_CH0_INT_RX_CLR_5(PCS_CH0_INT_RX_CLR_5), 
 .PCS_CH0_INT_RX_CLR_6(PCS_CH0_INT_RX_CLR_6), 
 .PCS_CH0_INT_RX_CLR_7(PCS_CH0_INT_RX_CLR_7), 
 .PCS_CH1_BYPASS_WORD_ALIGN(PCS_CH1_BYPASS_WORD_ALIGN), 
 .PCS_CH1_BYPASS_DENC(PCS_CH1_BYPASS_DENC), 
 .PCS_CH1_BYPASS_BONDING(PCS_CH1_BYPASS_BONDING), 
 .PCS_CH1_BYPASS_CTC(PCS_CH1_BYPASS_CTC), 
 .PCS_CH1_BYPASS_GEAR(PCS_CH1_BYPASS_GEAR), 
 .PCS_CH1_BYPASS_BRIDGE(PCS_CH1_BYPASS_BRIDGE), 
 .PCS_CH1_DATA_MODE(PCS_CH1_DATA_MODE), 
 .PCS_CH1_RX_POLARITY_INV(PCS_CH1_RX_POLARITY_INV), 
 .PCS_CH1_ALIGN_MODE(PCS_CH1_ALIGN_MODE), 
 .PCS_CH1_SAMP_16B(PCS_CH1_SAMP_16B), 
 .PCS_CH1_COMMA_REG0(PCS_CH1_COMMA_REG0), 
 .PCS_CH1_COMMA_MASK(PCS_CH1_COMMA_MASK), 
 .PCS_CH1_CEB_MODE(PCS_CH1_CEB_MODE), 
 .PCS_CH1_CTC_MODE(PCS_CH1_CTC_MODE), 
 .PCS_CH1_A_REG(PCS_CH1_A_REG), 
 .PCS_CH1_GE_AUTO_EN(PCS_CH1_GE_AUTO_EN), 
 .PCS_CH1_SKIP_REG0(PCS_CH1_SKIP_REG0), 
 .PCS_CH1_SKIP_REG1(PCS_CH1_SKIP_REG1), 
 .PCS_CH1_SKIP_REG2(PCS_CH1_SKIP_REG2), 
 .PCS_CH1_SKIP_REG3(PCS_CH1_SKIP_REG3), 
 .PCS_CH1_DEC_DUAL(PCS_CH1_DEC_DUAL), 
 .PCS_CH1_SPLIT(PCS_CH1_SPLIT), 
 .PCS_CH1_FIFOFLAG_CTC(PCS_CH1_FIFOFLAG_CTC), 
 .PCS_CH1_COMMA_DET_MODE(PCS_CH1_COMMA_DET_MODE), 
 .PCS_CH1_ERRDETECT_SILENCE(PCS_CH1_ERRDETECT_SILENCE), 
 .PCS_CH1_PMA_RCLK_POLINV(PCS_CH1_PMA_RCLK_POLINV), 
 .PCS_CH1_PCS_RCLK_SEL(PCS_CH1_PCS_RCLK_SEL), 
 .PCS_CH1_MCB_RCLK_POLINV(PCS_CH1_MCB_RCLK_POLINV), 
 .PCS_CH1_CB_RCLK_SEL(PCS_CH1_CB_RCLK_SEL), 
 .PCS_CH1_AFTER_CTC_RCLK_SEL(PCS_CH1_AFTER_CTC_RCLK_SEL), 
 .PCS_CH1_RCLK_POLINV(PCS_CH1_RCLK_POLINV), 
 .PCS_CH1_BRIDGE_RCLK_SEL(PCS_CH1_BRIDGE_RCLK_SEL), 
 .PCS_CH1_PCS_RCLK_EN(PCS_CH1_PCS_RCLK_EN), 
 .PCS_CH1_CB_RCLK_EN(PCS_CH1_CB_RCLK_EN), 
 .PCS_CH1_AFTER_CTC_RCLK_EN(PCS_CH1_AFTER_CTC_RCLK_EN), 
 .PCS_CH1_AFTER_CTC_RCLK_EN_GB(PCS_CH1_AFTER_CTC_RCLK_EN_GB), 
 .PCS_CH1_BRIDGE_RCLK_EN(PCS_CH1_BRIDGE_RCLK_EN), 
 .PCS_CH1_PCS_RX_RSTN(PCS_CH1_PCS_RX_RSTN), 
 .PCS_CH1_SLAVE(PCS_CH1_SLAVE), 
 .PCS_CH1_PCIE_SLAVE(PCS_CH1_PCIE_SLAVE), 
 .PCS_CH1_PCS_CB_RSTN(PCS_CH1_PCS_CB_RSTN), 
 .PCS_CH1_TX_BYPASS_BRIDGE_UINT(PCS_CH1_TX_BYPASS_BRIDGE_UINT), 
 .PCS_CH1_TX_BYPASS_GEAR(PCS_CH1_TX_BYPASS_GEAR), 
 .PCS_CH1_TX_BYPASS_ENC(PCS_CH1_TX_BYPASS_ENC), 
 .PCS_CH1_TX_BYPASS_BIT_SLIP(PCS_CH1_TX_BYPASS_BIT_SLIP), 
 .PCS_CH1_TX_GEAR_SPLIT(PCS_CH1_TX_GEAR_SPLIT), 
 .PCS_CH1_TX_DRIVE_REG_MODE(PCS_CH1_TX_DRIVE_REG_MODE), 
 .PCS_CH1_TX_BIT_SLIP_CYCLES(PCS_CH1_TX_BIT_SLIP_CYCLES), 
 .PCS_CH1_INT_TX_MASK_0(PCS_CH1_INT_TX_MASK_0), 
 .PCS_CH1_INT_TX_MASK_1(PCS_CH1_INT_TX_MASK_1), 
 .PCS_CH1_INT_TX_MASK_2(PCS_CH1_INT_TX_MASK_2), 
 .PCS_CH1_INT_TX_CLR_0(PCS_CH1_INT_TX_CLR_0), 
 .PCS_CH1_INT_TX_CLR_1(PCS_CH1_INT_TX_CLR_1), 
 .PCS_CH1_INT_TX_CLR_2(PCS_CH1_INT_TX_CLR_2), 
 .PCS_CH1_TX_PMA_TCLK_POLINV(PCS_CH1_TX_PMA_TCLK_POLINV), 
 .PCS_CH1_TX_PCS_CLK_EN_SEL(PCS_CH1_TX_PCS_CLK_EN_SEL), 
 .PCS_CH1_TX_BRIDGE_TCLK_SEL(PCS_CH1_TX_BRIDGE_TCLK_SEL), 
 .PCS_CH1_TX_TCLK_POLINV(PCS_CH1_TX_TCLK_POLINV), 
 .PCS_CH1_TX_PCS_TX_RSTN(PCS_CH1_TX_PCS_TX_RSTN), 
 .PCS_CH1_TX_SLAVE(PCS_CH1_TX_SLAVE), 
 .PCS_CH1_TX_BRIDGE_CLK_EN_SEL(PCS_CH1_TX_BRIDGE_CLK_EN_SEL), 
 .PCS_CH1_DATA_WIDTH_MODE(PCS_CH1_DATA_WIDTH_MODE), 
 .PCS_CH1_TX_TCLK2FABRIC_SEL(PCS_CH1_TX_TCLK2FABRIC_SEL), 
 .PCS_CH1_TX_OUTZZ(PCS_CH1_TX_OUTZZ), 
 .PCS_CH1_ENC_DUAL(PCS_CH1_ENC_DUAL), 
 .PCS_CH1_TX_BITSLIP_DATA_MODE(PCS_CH1_TX_BITSLIP_DATA_MODE), 
 .PCS_CH1_COMMA_REG1(PCS_CH1_COMMA_REG1), 
 .PCS_CH1_RAPID_IMAX(PCS_CH1_RAPID_IMAX), 
 .PCS_CH1_RAPID_VMIN_1(PCS_CH1_RAPID_VMIN_1), 
 .PCS_CH1_RAPID_VMIN_2(PCS_CH1_RAPID_VMIN_2), 
 .PCS_CH1_RX_PRBS_MODE(PCS_CH1_RX_PRBS_MODE), 
 .PCS_CH1_RX_ERRCNT_CLR(PCS_CH1_RX_ERRCNT_CLR), 
 .PCS_CH1_TX_PRBS_MODE(PCS_CH1_TX_PRBS_MODE), 
 .PCS_CH1_TX_INSERT_ER(PCS_CH1_TX_INSERT_ER), 
 .PCS_CH1_ENABLE_PRBS_GEN(PCS_CH1_ENABLE_PRBS_GEN), 
 .PCS_CH1_ERR_CNT(PCS_CH1_ERR_CNT), 
 .PCS_CH1_DEFAULT_RADDR(PCS_CH1_DEFAULT_RADDR), 
 .PCS_CH1_MASTER_CHECK_OFFSET(PCS_CH1_MASTER_CHECK_OFFSET), 
 .PCS_CH1_DELAY_SET(PCS_CH1_DELAY_SET), 
 .PCS_CH1_SEACH_OFFSET(PCS_CH1_SEACH_OFFSET), 
 .PCS_CH1_CEB_RAPIDLS_MMAX(PCS_CH1_CEB_RAPIDLS_MMAX), 
 .PCS_CH1_CTC_AFULL(PCS_CH1_CTC_AFULL), 
 .PCS_CH1_CTC_AEMPTY(PCS_CH1_CTC_AEMPTY), 
 .PCS_CH1_FAR_LOOP(PCS_CH1_FAR_LOOP), 
 .PCS_CH1_NEAR_LOOP(PCS_CH1_NEAR_LOOP), 
 .PCS_CH1_INT_RX_MASK_0(PCS_CH1_INT_RX_MASK_0), 
 .PCS_CH1_INT_RX_MASK_1(PCS_CH1_INT_RX_MASK_1), 
 .PCS_CH1_INT_RX_MASK_2(PCS_CH1_INT_RX_MASK_2), 
 .PCS_CH1_INT_RX_MASK_3(PCS_CH1_INT_RX_MASK_3), 
 .PCS_CH1_INT_RX_MASK_4(PCS_CH1_INT_RX_MASK_4), 
 .PCS_CH1_INT_RX_MASK_5(PCS_CH1_INT_RX_MASK_5), 
 .PCS_CH1_INT_RX_MASK_6(PCS_CH1_INT_RX_MASK_6), 
 .PCS_CH1_INT_RX_MASK_7(PCS_CH1_INT_RX_MASK_7), 
 .PCS_CH1_INT_RX_CLR_0(PCS_CH1_INT_RX_CLR_0), 
 .PCS_CH1_INT_RX_CLR_1(PCS_CH1_INT_RX_CLR_1), 
 .PCS_CH1_INT_RX_CLR_2(PCS_CH1_INT_RX_CLR_2), 
 .PCS_CH1_INT_RX_CLR_3(PCS_CH1_INT_RX_CLR_3), 
 .PCS_CH1_INT_RX_CLR_4(PCS_CH1_INT_RX_CLR_4), 
 .PCS_CH1_INT_RX_CLR_5(PCS_CH1_INT_RX_CLR_5), 
 .PCS_CH1_INT_RX_CLR_6(PCS_CH1_INT_RX_CLR_6), 
 .PCS_CH1_INT_RX_CLR_7(PCS_CH1_INT_RX_CLR_7), 
 .PCS_CH2_BYPASS_WORD_ALIGN(PCS_CH2_BYPASS_WORD_ALIGN), 
 .PCS_CH2_BYPASS_DENC(PCS_CH2_BYPASS_DENC), 
 .PCS_CH2_BYPASS_BONDING(PCS_CH2_BYPASS_BONDING), 
 .PCS_CH2_BYPASS_CTC(PCS_CH2_BYPASS_CTC), 
 .PCS_CH2_BYPASS_GEAR(PCS_CH2_BYPASS_GEAR), 
 .PCS_CH2_BYPASS_BRIDGE(PCS_CH2_BYPASS_BRIDGE), 
 .PCS_CH2_DATA_MODE(PCS_CH2_DATA_MODE), 
 .PCS_CH2_RX_POLARITY_INV(PCS_CH2_RX_POLARITY_INV), 
 .PCS_CH2_ALIGN_MODE(PCS_CH2_ALIGN_MODE), 
 .PCS_CH2_SAMP_16B(PCS_CH2_SAMP_16B), 
 .PCS_CH2_COMMA_REG0(PCS_CH2_COMMA_REG0), 
 .PCS_CH2_COMMA_MASK(PCS_CH2_COMMA_MASK), 
 .PCS_CH2_CEB_MODE(PCS_CH2_CEB_MODE), 
 .PCS_CH2_CTC_MODE(PCS_CH2_CTC_MODE), 
 .PCS_CH2_A_REG(PCS_CH2_A_REG), 
 .PCS_CH2_GE_AUTO_EN(PCS_CH2_GE_AUTO_EN), 
 .PCS_CH2_SKIP_REG0(PCS_CH2_SKIP_REG0), 
 .PCS_CH2_SKIP_REG1(PCS_CH2_SKIP_REG1), 
 .PCS_CH2_SKIP_REG2(PCS_CH2_SKIP_REG2), 
 .PCS_CH2_SKIP_REG3(PCS_CH2_SKIP_REG3), 
 .PCS_CH2_DEC_DUAL(PCS_CH2_DEC_DUAL), 
 .PCS_CH2_SPLIT(PCS_CH2_SPLIT), 
 .PCS_CH2_FIFOFLAG_CTC(PCS_CH2_FIFOFLAG_CTC), 
 .PCS_CH2_COMMA_DET_MODE(PCS_CH2_COMMA_DET_MODE), 
 .PCS_CH2_ERRDETECT_SILENCE(PCS_CH2_ERRDETECT_SILENCE), 
 .PCS_CH2_PMA_RCLK_POLINV(PCS_CH2_PMA_RCLK_POLINV), 
 .PCS_CH2_PCS_RCLK_SEL(PCS_CH2_PCS_RCLK_SEL), 
 .PCS_CH2_MCB_RCLK_POLINV(PCS_CH2_MCB_RCLK_POLINV), 
 .PCS_CH2_CB_RCLK_SEL(PCS_CH2_CB_RCLK_SEL), 
 .PCS_CH2_AFTER_CTC_RCLK_SEL(PCS_CH2_AFTER_CTC_RCLK_SEL), 
 .PCS_CH2_RCLK_POLINV(PCS_CH2_RCLK_POLINV), 
 .PCS_CH2_BRIDGE_RCLK_SEL(PCS_CH2_BRIDGE_RCLK_SEL), 
 .PCS_CH2_PCS_RCLK_EN(PCS_CH2_PCS_RCLK_EN), 
 .PCS_CH2_CB_RCLK_EN(PCS_CH2_CB_RCLK_EN), 
 .PCS_CH2_AFTER_CTC_RCLK_EN(PCS_CH2_AFTER_CTC_RCLK_EN), 
 .PCS_CH2_AFTER_CTC_RCLK_EN_GB(PCS_CH2_AFTER_CTC_RCLK_EN_GB), 
 .PCS_CH2_BRIDGE_RCLK_EN(PCS_CH2_BRIDGE_RCLK_EN), 
 .PCS_CH2_PCS_RX_RSTN(PCS_CH2_PCS_RX_RSTN), 
 .PCS_CH2_SLAVE(PCS_CH2_SLAVE), 
 .PCS_CH2_PCIE_SLAVE(PCS_CH2_PCIE_SLAVE), 
 .PCS_CH2_PCS_CB_RSTN(PCS_CH2_PCS_CB_RSTN), 
 .PCS_CH2_TX_BYPASS_BRIDGE_UINT(PCS_CH2_TX_BYPASS_BRIDGE_UINT), 
 .PCS_CH2_TX_BYPASS_GEAR(PCS_CH2_TX_BYPASS_GEAR), 
 .PCS_CH2_TX_BYPASS_ENC(PCS_CH2_TX_BYPASS_ENC), 
 .PCS_CH2_TX_BYPASS_BIT_SLIP(PCS_CH2_TX_BYPASS_BIT_SLIP), 
 .PCS_CH2_TX_GEAR_SPLIT(PCS_CH2_TX_GEAR_SPLIT), 
 .PCS_CH2_TX_DRIVE_REG_MODE(PCS_CH2_TX_DRIVE_REG_MODE), 
 .PCS_CH2_TX_BIT_SLIP_CYCLES(PCS_CH2_TX_BIT_SLIP_CYCLES), 
 .PCS_CH2_INT_TX_MASK_0(PCS_CH2_INT_TX_MASK_0), 
 .PCS_CH2_INT_TX_MASK_1(PCS_CH2_INT_TX_MASK_1), 
 .PCS_CH2_INT_TX_MASK_2(PCS_CH2_INT_TX_MASK_2), 
 .PCS_CH2_INT_TX_CLR_0(PCS_CH2_INT_TX_CLR_0), 
 .PCS_CH2_INT_TX_CLR_1(PCS_CH2_INT_TX_CLR_1), 
 .PCS_CH2_INT_TX_CLR_2(PCS_CH2_INT_TX_CLR_2), 
 .PCS_CH2_TX_PMA_TCLK_POLINV(PCS_CH2_TX_PMA_TCLK_POLINV), 
 .PCS_CH2_TX_PCS_CLK_EN_SEL(PCS_CH2_TX_PCS_CLK_EN_SEL), 
 .PCS_CH2_TX_BRIDGE_TCLK_SEL(PCS_CH2_TX_BRIDGE_TCLK_SEL), 
 .PCS_CH2_TX_TCLK_POLINV(PCS_CH2_TX_TCLK_POLINV), 
 .PCS_CH2_TX_PCS_TX_RSTN(PCS_CH2_TX_PCS_TX_RSTN), 
 .PCS_CH2_TX_SLAVE(PCS_CH2_TX_SLAVE), 
 .PCS_CH2_TX_BRIDGE_CLK_EN_SEL(PCS_CH2_TX_BRIDGE_CLK_EN_SEL), 
 .PCS_CH2_DATA_WIDTH_MODE(PCS_CH2_DATA_WIDTH_MODE), 
 .PCS_CH2_TX_TCLK2FABRIC_SEL(PCS_CH2_TX_TCLK2FABRIC_SEL), 
 .PCS_CH2_TX_OUTZZ(PCS_CH2_TX_OUTZZ), 
 .PCS_CH2_ENC_DUAL(PCS_CH2_ENC_DUAL), 
 .PCS_CH2_TX_BITSLIP_DATA_MODE(PCS_CH2_TX_BITSLIP_DATA_MODE), 
 .PCS_CH2_COMMA_REG1(PCS_CH2_COMMA_REG1), 
 .PCS_CH2_RAPID_IMAX(PCS_CH2_RAPID_IMAX), 
 .PCS_CH2_RAPID_VMIN_1(PCS_CH2_RAPID_VMIN_1), 
 .PCS_CH2_RAPID_VMIN_2(PCS_CH2_RAPID_VMIN_2), 
 .PCS_CH2_RX_PRBS_MODE(PCS_CH2_RX_PRBS_MODE), 
 .PCS_CH2_RX_ERRCNT_CLR(PCS_CH2_RX_ERRCNT_CLR), 
 .PCS_CH2_TX_PRBS_MODE(PCS_CH2_TX_PRBS_MODE), 
 .PCS_CH2_TX_INSERT_ER(PCS_CH2_TX_INSERT_ER), 
 .PCS_CH2_ENABLE_PRBS_GEN(PCS_CH2_ENABLE_PRBS_GEN), 
 .PCS_CH2_ERR_CNT(PCS_CH2_ERR_CNT), 
 .PCS_CH2_DEFAULT_RADDR(PCS_CH2_DEFAULT_RADDR), 
 .PCS_CH2_MASTER_CHECK_OFFSET(PCS_CH2_MASTER_CHECK_OFFSET), 
 .PCS_CH2_DELAY_SET(PCS_CH2_DELAY_SET), 
 .PCS_CH2_SEACH_OFFSET(PCS_CH2_SEACH_OFFSET), 
 .PCS_CH2_CEB_RAPIDLS_MMAX(PCS_CH2_CEB_RAPIDLS_MMAX), 
 .PCS_CH2_CTC_AFULL(PCS_CH2_CTC_AFULL), 
 .PCS_CH2_CTC_AEMPTY(PCS_CH2_CTC_AEMPTY), 
 .PCS_CH2_FAR_LOOP(PCS_CH2_FAR_LOOP), 
 .PCS_CH2_NEAR_LOOP(PCS_CH2_NEAR_LOOP), 
 .PCS_CH2_INT_RX_MASK_0(PCS_CH2_INT_RX_MASK_0), 
 .PCS_CH2_INT_RX_MASK_1(PCS_CH2_INT_RX_MASK_1), 
 .PCS_CH2_INT_RX_MASK_2(PCS_CH2_INT_RX_MASK_2), 
 .PCS_CH2_INT_RX_MASK_3(PCS_CH2_INT_RX_MASK_3), 
 .PCS_CH2_INT_RX_MASK_4(PCS_CH2_INT_RX_MASK_4), 
 .PCS_CH2_INT_RX_MASK_5(PCS_CH2_INT_RX_MASK_5), 
 .PCS_CH2_INT_RX_MASK_6(PCS_CH2_INT_RX_MASK_6), 
 .PCS_CH2_INT_RX_MASK_7(PCS_CH2_INT_RX_MASK_7), 
 .PCS_CH2_INT_RX_CLR_0(PCS_CH2_INT_RX_CLR_0), 
 .PCS_CH2_INT_RX_CLR_1(PCS_CH2_INT_RX_CLR_1), 
 .PCS_CH2_INT_RX_CLR_2(PCS_CH2_INT_RX_CLR_2), 
 .PCS_CH2_INT_RX_CLR_3(PCS_CH2_INT_RX_CLR_3), 
 .PCS_CH2_INT_RX_CLR_4(PCS_CH2_INT_RX_CLR_4), 
 .PCS_CH2_INT_RX_CLR_5(PCS_CH2_INT_RX_CLR_5), 
 .PCS_CH2_INT_RX_CLR_6(PCS_CH2_INT_RX_CLR_6), 
 .PCS_CH2_INT_RX_CLR_7(PCS_CH2_INT_RX_CLR_7), 
 .PCS_CH3_BYPASS_WORD_ALIGN(PCS_CH3_BYPASS_WORD_ALIGN), 
 .PCS_CH3_BYPASS_DENC(PCS_CH3_BYPASS_DENC), 
 .PCS_CH3_BYPASS_BONDING(PCS_CH3_BYPASS_BONDING), 
 .PCS_CH3_BYPASS_CTC(PCS_CH3_BYPASS_CTC), 
 .PCS_CH3_BYPASS_GEAR(PCS_CH3_BYPASS_GEAR), 
 .PCS_CH3_BYPASS_BRIDGE(PCS_CH3_BYPASS_BRIDGE), 
 .PCS_CH3_DATA_MODE(PCS_CH3_DATA_MODE), 
 .PCS_CH3_RX_POLARITY_INV(PCS_CH3_RX_POLARITY_INV), 
 .PCS_CH3_ALIGN_MODE(PCS_CH3_ALIGN_MODE), 
 .PCS_CH3_SAMP_16B(PCS_CH3_SAMP_16B), 
 .PCS_CH3_COMMA_REG0(PCS_CH3_COMMA_REG0), 
 .PCS_CH3_COMMA_MASK(PCS_CH3_COMMA_MASK), 
 .PCS_CH3_CEB_MODE(PCS_CH3_CEB_MODE), 
 .PCS_CH3_CTC_MODE(PCS_CH3_CTC_MODE), 
 .PCS_CH3_A_REG(PCS_CH3_A_REG), 
 .PCS_CH3_GE_AUTO_EN(PCS_CH3_GE_AUTO_EN), 
 .PCS_CH3_SKIP_REG0(PCS_CH3_SKIP_REG0), 
 .PCS_CH3_SKIP_REG1(PCS_CH3_SKIP_REG1), 
 .PCS_CH3_SKIP_REG2(PCS_CH3_SKIP_REG2), 
 .PCS_CH3_SKIP_REG3(PCS_CH3_SKIP_REG3), 
 .PCS_CH3_DEC_DUAL(PCS_CH3_DEC_DUAL), 
 .PCS_CH3_SPLIT(PCS_CH3_SPLIT), 
 .PCS_CH3_FIFOFLAG_CTC(PCS_CH3_FIFOFLAG_CTC), 
 .PCS_CH3_COMMA_DET_MODE(PCS_CH3_COMMA_DET_MODE), 
 .PCS_CH3_ERRDETECT_SILENCE(PCS_CH3_ERRDETECT_SILENCE), 
 .PCS_CH3_PMA_RCLK_POLINV(PCS_CH3_PMA_RCLK_POLINV), 
 .PCS_CH3_PCS_RCLK_SEL(PCS_CH3_PCS_RCLK_SEL), 
 .PCS_CH3_MCB_RCLK_POLINV(PCS_CH3_MCB_RCLK_POLINV), 
 .PCS_CH3_CB_RCLK_SEL(PCS_CH3_CB_RCLK_SEL), 
 .PCS_CH3_AFTER_CTC_RCLK_SEL(PCS_CH3_AFTER_CTC_RCLK_SEL), 
 .PCS_CH3_RCLK_POLINV(PCS_CH3_RCLK_POLINV), 
 .PCS_CH3_BRIDGE_RCLK_SEL(PCS_CH3_BRIDGE_RCLK_SEL), 
 .PCS_CH3_PCS_RCLK_EN(PCS_CH3_PCS_RCLK_EN), 
 .PCS_CH3_CB_RCLK_EN(PCS_CH3_CB_RCLK_EN), 
 .PCS_CH3_AFTER_CTC_RCLK_EN(PCS_CH3_AFTER_CTC_RCLK_EN), 
 .PCS_CH3_AFTER_CTC_RCLK_EN_GB(PCS_CH3_AFTER_CTC_RCLK_EN_GB), 
 .PCS_CH3_BRIDGE_RCLK_EN(PCS_CH3_BRIDGE_RCLK_EN), 
 .PCS_CH3_PCS_RX_RSTN(PCS_CH3_PCS_RX_RSTN), 
 .PCS_CH3_SLAVE(PCS_CH3_SLAVE), 
 .PCS_CH3_PCIE_SLAVE(PCS_CH3_PCIE_SLAVE), 
 .PCS_CH3_PCS_CB_RSTN(PCS_CH3_PCS_CB_RSTN), 
 .PCS_CH3_TX_BYPASS_BRIDGE_UINT(PCS_CH3_TX_BYPASS_BRIDGE_UINT), 
 .PCS_CH3_TX_BYPASS_GEAR(PCS_CH3_TX_BYPASS_GEAR), 
 .PCS_CH3_TX_BYPASS_ENC(PCS_CH3_TX_BYPASS_ENC), 
 .PCS_CH3_TX_BYPASS_BIT_SLIP(PCS_CH3_TX_BYPASS_BIT_SLIP), 
 .PCS_CH3_TX_GEAR_SPLIT(PCS_CH3_TX_GEAR_SPLIT), 
 .PCS_CH3_TX_DRIVE_REG_MODE(PCS_CH3_TX_DRIVE_REG_MODE), 
 .PCS_CH3_TX_BIT_SLIP_CYCLES(PCS_CH3_TX_BIT_SLIP_CYCLES), 
 .PCS_CH3_INT_TX_MASK_0(PCS_CH3_INT_TX_MASK_0), 
 .PCS_CH3_INT_TX_MASK_1(PCS_CH3_INT_TX_MASK_1), 
 .PCS_CH3_INT_TX_MASK_2(PCS_CH3_INT_TX_MASK_2), 
 .PCS_CH3_INT_TX_CLR_0(PCS_CH3_INT_TX_CLR_0), 
 .PCS_CH3_INT_TX_CLR_1(PCS_CH3_INT_TX_CLR_1), 
 .PCS_CH3_INT_TX_CLR_2(PCS_CH3_INT_TX_CLR_2), 
 .PCS_CH3_TX_PMA_TCLK_POLINV(PCS_CH3_TX_PMA_TCLK_POLINV), 
 .PCS_CH3_TX_PCS_CLK_EN_SEL(PCS_CH3_TX_PCS_CLK_EN_SEL), 
 .PCS_CH3_TX_BRIDGE_TCLK_SEL(PCS_CH3_TX_BRIDGE_TCLK_SEL), 
 .PCS_CH3_TX_TCLK_POLINV(PCS_CH3_TX_TCLK_POLINV), 
 .PCS_CH3_TX_PCS_TX_RSTN(PCS_CH3_TX_PCS_TX_RSTN), 
 .PCS_CH3_TX_SLAVE(PCS_CH3_TX_SLAVE), 
 .PCS_CH3_TX_BRIDGE_CLK_EN_SEL(PCS_CH3_TX_BRIDGE_CLK_EN_SEL), 
 .PCS_CH3_DATA_WIDTH_MODE(PCS_CH3_DATA_WIDTH_MODE), 
 .PCS_CH3_TX_TCLK2FABRIC_SEL(PCS_CH3_TX_TCLK2FABRIC_SEL), 
 .PCS_CH3_TX_OUTZZ(PCS_CH3_TX_OUTZZ), 
 .PCS_CH3_ENC_DUAL(PCS_CH3_ENC_DUAL), 
 .PCS_CH3_TX_BITSLIP_DATA_MODE(PCS_CH3_TX_BITSLIP_DATA_MODE), 
 .PCS_CH3_COMMA_REG1(PCS_CH3_COMMA_REG1), 
 .PCS_CH3_RAPID_IMAX(PCS_CH3_RAPID_IMAX), 
 .PCS_CH3_RAPID_VMIN_1(PCS_CH3_RAPID_VMIN_1), 
 .PCS_CH3_RAPID_VMIN_2(PCS_CH3_RAPID_VMIN_2), 
 .PCS_CH3_RX_PRBS_MODE(PCS_CH3_RX_PRBS_MODE), 
 .PCS_CH3_RX_ERRCNT_CLR(PCS_CH3_RX_ERRCNT_CLR), 
 .PCS_CH3_TX_PRBS_MODE(PCS_CH3_TX_PRBS_MODE), 
 .PCS_CH3_TX_INSERT_ER(PCS_CH3_TX_INSERT_ER), 
 .PCS_CH3_ENABLE_PRBS_GEN(PCS_CH3_ENABLE_PRBS_GEN), 
 .PCS_CH3_ERR_CNT(PCS_CH3_ERR_CNT), 
 .PCS_CH3_DEFAULT_RADDR(PCS_CH3_DEFAULT_RADDR), 
 .PCS_CH3_MASTER_CHECK_OFFSET(PCS_CH3_MASTER_CHECK_OFFSET), 
 .PCS_CH3_DELAY_SET(PCS_CH3_DELAY_SET), 
 .PCS_CH3_SEACH_OFFSET(PCS_CH3_SEACH_OFFSET), 
 .PCS_CH3_CEB_RAPIDLS_MMAX(PCS_CH3_CEB_RAPIDLS_MMAX), 
 .PCS_CH3_CTC_AFULL(PCS_CH3_CTC_AFULL), 
 .PCS_CH3_CTC_AEMPTY(PCS_CH3_CTC_AEMPTY), 
 .PCS_CH3_FAR_LOOP(PCS_CH3_FAR_LOOP), 
 .PCS_CH3_NEAR_LOOP(PCS_CH3_NEAR_LOOP), 
 .PCS_CH3_INT_RX_MASK_0(PCS_CH3_INT_RX_MASK_0), 
 .PCS_CH3_INT_RX_MASK_1(PCS_CH3_INT_RX_MASK_1), 
 .PCS_CH3_INT_RX_MASK_2(PCS_CH3_INT_RX_MASK_2), 
 .PCS_CH3_INT_RX_MASK_3(PCS_CH3_INT_RX_MASK_3), 
 .PCS_CH3_INT_RX_MASK_4(PCS_CH3_INT_RX_MASK_4), 
 .PCS_CH3_INT_RX_MASK_5(PCS_CH3_INT_RX_MASK_5), 
 .PCS_CH3_INT_RX_MASK_6(PCS_CH3_INT_RX_MASK_6), 
 .PCS_CH3_INT_RX_MASK_7(PCS_CH3_INT_RX_MASK_7), 
 .PCS_CH3_INT_RX_CLR_0(PCS_CH3_INT_RX_CLR_0), 
 .PCS_CH3_INT_RX_CLR_1(PCS_CH3_INT_RX_CLR_1), 
 .PCS_CH3_INT_RX_CLR_2(PCS_CH3_INT_RX_CLR_2), 
 .PCS_CH3_INT_RX_CLR_3(PCS_CH3_INT_RX_CLR_3), 
 .PCS_CH3_INT_RX_CLR_4(PCS_CH3_INT_RX_CLR_4), 
 .PCS_CH3_INT_RX_CLR_5(PCS_CH3_INT_RX_CLR_5), 
 .PCS_CH3_INT_RX_CLR_6(PCS_CH3_INT_RX_CLR_6), 
 .PCS_CH3_INT_RX_CLR_7(PCS_CH3_INT_RX_CLR_7), 
 .PMA_CH0_TXDATA_WIDTH(PMA_CH0_TXDATA_WIDTH), 
 .PMA_CH0_TX_TESTPATTERN(PMA_CH0_TX_TESTPATTERN), 
 .PMA_CH0_TESTPATTERN_O_ENABLE(PMA_CH0_TESTPATTERN_O_ENABLE), 
 .PMA_CH0_DISABLE_BSMODE_DRVAMP(PMA_CH0_DISABLE_BSMODE_DRVAMP), 
 .PMA_CH0_FORCE_BIST_ENABLE(PMA_CH0_FORCE_BIST_ENABLE), 
 .PMA_CH0_FORCE_ELECTRICAL_IDLE(PMA_CH0_FORCE_ELECTRICAL_IDLE), 
 .PMA_CH0_FORCE_RXDCT_ENABLE(PMA_CH0_FORCE_RXDCT_ENABLE), 
 .PMA_CH0_FORCE_EXTLB_ENABLE(PMA_CH0_FORCE_EXTLB_ENABLE), 
 .PMA_CH0_DISABLE_LANE_SYNC(PMA_CH0_DISABLE_LANE_SYNC), 
 .PMA_CH0_DISABLE_ELECTRICAL_IDLE(PMA_CH0_DISABLE_ELECTRICAL_IDLE), 
 .PMA_CH0_DISABLE_RXDCT_ENABLE(PMA_CH0_DISABLE_RXDCT_ENABLE), 
 .PMA_CH0_DISABLE_EXTLB_ENABLE(PMA_CH0_DISABLE_EXTLB_ENABLE), 
 .PMA_CH0_DISABLE_LOW_SPEED_PATH_ENABLE(PMA_CH0_DISABLE_LOW_SPEED_PATH_ENABLE), 
 .PMA_CH0_FORCE_LANE_ENABLE(PMA_CH0_FORCE_LANE_ENABLE), 
 .PMA_CH0_FORCE_LANE_RESETB_DISABLE(PMA_CH0_FORCE_LANE_RESETB_DISABLE), 
 .PMA_CH0_RXDCT_LGBW_ENABLE(PMA_CH0_RXDCT_LGBW_ENABLE), 
 .PMA_CH0_RXDCT_VTH(PMA_CH0_RXDCT_VTH), 
 .PMA_CH0_DE_EMPHASIS_ADDITIONAL_CONTROL(PMA_CH0_DE_EMPHASIS_ADDITIONAL_CONTROL), 
 .PMA_CH0_DRV_RTERM_CONTROL(PMA_CH0_DRV_RTERM_CONTROL), 
 .PMA_CH0_FDRV_AMP_CONTROL(PMA_CH0_FDRV_AMP_CONTROL), 
 .PMA_CH0_PREPC_AMP_CONTROL(PMA_CH0_PREPC_AMP_CONTROL), 
 .PMA_CH0_PREMC_AMP_CONTROL(PMA_CH0_PREMC_AMP_CONTROL), 
 .PMA_CH0_SER_AMP_CONTROL(PMA_CH0_SER_AMP_CONTROL), 
 .PMA_CH0_PFD_LOOP_RESISTOR_SETTING(PMA_CH0_PFD_LOOP_RESISTOR_SETTING), 
 .PMA_CH0_PD_LOOP_RESISTOR_SETTING(PMA_CH0_PD_LOOP_RESISTOR_SETTING), 
 .PMA_CH0_CDR_TEST_OUT_SELECT(PMA_CH0_CDR_TEST_OUT_SELECT), 
 .PMA_CH0_PI_DIV1_BP(PMA_CH0_PI_DIV1_BP), 
 .PMA_CH0_PI_TEST_FOR_CKI(PMA_CH0_PI_TEST_FOR_CKI), 
 .PMA_CH0_PI_CURRENT_SETTING(PMA_CH0_PI_CURRENT_SETTING), 
 .PMA_CH0_PI_FREQUENCY_SETTING(PMA_CH0_PI_FREQUENCY_SETTING), 
 .PMA_CH0_TEST_OUT_SELECT_FOR_RCK(PMA_CH0_TEST_OUT_SELECT_FOR_RCK), 
 .PMA_CH0_TEST_OUT_SELECT_SOURCE(PMA_CH0_TEST_OUT_SELECT_SOURCE), 
 .PMA_CH0_TEST_DATA_OUT_SELECT_SOURCE(PMA_CH0_TEST_DATA_OUT_SELECT_SOURCE), 
 .PMA_CH0_TEST_CK_OUT_SELECT_SOURCE(PMA_CH0_TEST_CK_OUT_SELECT_SOURCE), 
 .PMA_CH0_ENABLE_SLIP1UI_MODULE(PMA_CH0_ENABLE_SLIP1UI_MODULE), 
 .PMA_CH0_PN_SWAP_ENABLE(PMA_CH0_PN_SWAP_ENABLE), 
 .PMA_CH0_SIPO_BIT_SETTING(PMA_CH0_SIPO_BIT_SETTING), 
 .PMA_CH0_OOB_EN(PMA_CH0_OOB_EN), 
 .PMA_CH0_ALOS_EN(PMA_CH0_ALOS_EN), 
 .PMA_CH0_LFMODE(PMA_CH0_LFMODE), 
 .PMA_CH0_TSO_HS_SEL(PMA_CH0_TSO_HS_SEL), 
 .PMA_CH0_LX_SELLC(PMA_CH0_LX_SELLC), 
 .PMA_CH0_LX_RXPLL_DIVSEL45_FB(PMA_CH0_LX_RXPLL_DIVSEL45_FB), 
 .PMA_CH0_LX_RXPLL_DIVSEL_FB(PMA_CH0_LX_RXPLL_DIVSEL_FB), 
 .PMA_CH0_LX_RXPLL_DIVSEL_REF(PMA_CH0_LX_RXPLL_DIVSEL_REF), 
 .PMA_CH0_PICODE(PMA_CH0_PICODE), 
 .PMA_CH0_RX_REFCK_SEL(PMA_CH0_RX_REFCK_SEL), 
 .PMA_CH0_PFDLPEN_REGISTER_CONTROL_ENABLE(PMA_CH0_PFDLPEN_REGISTER_CONTROL_ENABLE), 
 .PMA_CH0_PFDLPEN_REGISTER_SETTING(PMA_CH0_PFDLPEN_REGISTER_SETTING), 
 .PMA_CH0_PDLPEN_REGISTER_CONTROL_ENABLE(PMA_CH0_PDLPEN_REGISTER_CONTROL_ENABLE), 
 .PMA_CH0_PDLPEN_REGISTER_SETTING(PMA_CH0_PDLPEN_REGISTER_SETTING), 
 .PMA_CH0_DIV_CHANGE_ENABLE_DELAY_TIMER(PMA_CH0_DIV_CHANGE_ENABLE_DELAY_TIMER), 
 .PMA_CH0_DIV_CHANGE_ENABLE_SIGNAL_GATING(PMA_CH0_DIV_CHANGE_ENABLE_SIGNAL_GATING), 
 .PMA_CH0_CDR_ALIGN_REGISTER_SETTING_VALUE(PMA_CH0_CDR_ALIGN_REGISTER_SETTING_VALUE), 
 .PMA_CH0_FORCE_CDR_ALIGN_ENABLE(PMA_CH0_FORCE_CDR_ALIGN_ENABLE), 
 .PMA_CH0_SELLC_REGISTER_SETTING_VALUE(PMA_CH0_SELLC_REGISTER_SETTING_VALUE), 
 .PMA_CH0_SELLC_CONTROL_BY_REGISTER(PMA_CH0_SELLC_CONTROL_BY_REGISTER), 
 .PMA_CH0_REG_PLLI_LDO_VREF_SETTING(PMA_CH0_REG_PLLI_LDO_VREF_SETTING), 
 .PMA_CH0_REG_PLLI_LDO_BYPASS_CURRENT(PMA_CH0_REG_PLLI_LDO_BYPASS_CURRENT), 
 .PMA_CH0_REG_PLL_HSTEST_ENABLE(PMA_CH0_REG_PLL_HSTEST_ENABLE), 
 .PMA_CH0_REG_PLL_ISNK_CURRENT_CONTROL(PMA_CH0_REG_PLL_ISNK_CURRENT_CONTROL), 
 .PMA_CH0_REG_PLL_PFD_LOOP_CP0_CURRENT_SETTING(PMA_CH0_REG_PLL_PFD_LOOP_CP0_CURRENT_SETTING), 
 .PMA_CH0_REG_PLL_PD_LOOP_PLLGM_SETTING(PMA_CH0_REG_PLL_PD_LOOP_PLLGM_SETTING), 
 .PMA_CH0_REG_PLL_PFD_LOOP_CP1_CURRENT_SETTING(PMA_CH0_REG_PLL_PFD_LOOP_CP1_CURRENT_SETTING), 
 .PMA_CH0_REG_PLL_CP0_BIAS_CONTROL(PMA_CH0_REG_PLL_CP0_BIAS_CONTROL), 
 .PMA_CH0_REG_PLL_PD_LOOP_CP0_CURRENT_SETTING(PMA_CH0_REG_PLL_PD_LOOP_CP0_CURRENT_SETTING), 
 .PMA_CH0_REG_PLL_CP1_BIAS_CONTROL(PMA_CH0_REG_PLL_CP1_BIAS_CONTROL), 
 .PMA_CH0_REG_PLL_PD_LOOP_CP1_CURRENT_SETTING(PMA_CH0_REG_PLL_PD_LOOP_CP1_CURRENT_SETTING), 
 .PMA_CH0_REG_PLL_CP0_CURRENT_SETTING(PMA_CH0_REG_PLL_CP0_CURRENT_SETTING), 
 .PMA_CH0_REG_PLL_CP1_CURRENT_SETTING(PMA_CH0_REG_PLL_CP1_CURRENT_SETTING), 
 .PMA_CH0_REG_PLL_GM1_CURRENT_SETTING(PMA_CH0_REG_PLL_GM1_CURRENT_SETTING), 
 .PMA_CH0_REG_PLL_LC_BF2_CURRENT_SETTING(PMA_CH0_REG_PLL_LC_BF2_CURRENT_SETTING), 
 .PMA_CH0_REG_PLL_LC_BF2_CURRENT_SETTING_LOW(PMA_CH0_REG_PLL_LC_BF2_CURRENT_SETTING_LOW), 
 .PMA_CH0_REG_PLL_REG_CUR(PMA_CH0_REG_PLL_REG_CUR), 
 .PMA_CH0_REG_PLL_LCCUR(PMA_CH0_REG_PLL_LCCUR), 
 .PMA_CH0_REG_PLL_LCOBAS(PMA_CH0_REG_PLL_LCOBAS), 
 .PMA_CH0_REG_PLL_FB_CK_TEST_OUT_ENABLE(PMA_CH0_REG_PLL_FB_CK_TEST_OUT_ENABLE), 
 .PMA_CH0_CDR_ALIGN_TIMER(PMA_CH0_CDR_ALIGN_TIMER), 
 .PMA_CH0_CALIB_WAIT(PMA_CH0_CALIB_WAIT), 
 .PMA_CH0_CALIB_TIMER(PMA_CH0_CALIB_TIMER), 
 .PMA_CH0_TOT_RANGE(PMA_CH0_TOT_RANGE), 
 .PMA_CH0_SUB_RANGE(PMA_CH0_SUB_RANGE), 
 .PMA_CH0_OVLP(PMA_CH0_OVLP), 
 .PMA_CH0_BIST_WAIT(PMA_CH0_BIST_WAIT), 
 .PMA_CH0_BIST_TIMER(PMA_CH0_BIST_TIMER), 
 .PMA_CH0_BAND_LB(PMA_CH0_BAND_LB), 
 .PMA_CH0_BAND_HB(PMA_CH0_BAND_HB), 
 .PMA_CH0_FREQ_LOCK_ACCURACY(PMA_CH0_FREQ_LOCK_ACCURACY), 
 .PMA_CH0_REG_SET_LC_BAND(PMA_CH0_REG_SET_LC_BAND), 
 .PMA_CH0_REG_SET_VCODIV(PMA_CH0_REG_SET_VCODIV), 
 .PMA_CH0_REGISTER_SET_VCODIV_BAND_ENABLE(PMA_CH0_REGISTER_SET_VCODIV_BAND_ENABLE), 
 .PMA_CH0_REG_SET_PLL_LOCK(PMA_CH0_REG_SET_PLL_LOCK), 
 .PMA_CH0_REGISTER_SET_PLL_LOCK_ENABLE(PMA_CH0_REGISTER_SET_PLL_LOCK_ENABLE), 
 .PMA_CH0_REG_SET_VCO_HI(PMA_CH0_REG_SET_VCO_HI), 
 .PMA_CH0_REG_SET_VCO_LO(PMA_CH0_REG_SET_VCO_LO), 
 .PMA_CH0_REGISTER_SET_VCO_HI_VCO_LO_ENABLE(PMA_CH0_REGISTER_SET_VCO_HI_VCO_LO_ENABLE), 
 .PMA_CH0_FORCE_LC_PLL_LOOP_EN_H(PMA_CH0_FORCE_LC_PLL_LOOP_EN_H), 
 .PMA_CH0_FORCE_LC_PLL_LOOP_EN_L(PMA_CH0_FORCE_LC_PLL_LOOP_EN_L), 
 .PMA_CH0_VCO_DIV_CALI_BYPASS(PMA_CH0_VCO_DIV_CALI_BYPASS), 
 .PMA_CH0_BIST_EN(PMA_CH0_BIST_EN), 
 .PMA_CH0_PLL_LOOP_EN_SETTING_FROM_REGISTER_ENABLE(PMA_CH0_PLL_LOOP_EN_SETTING_FROM_REGISTER_ENABLE), 
 .PMA_CH0_FREQ_DETECT_ENABLE_SOURCE(PMA_CH0_FREQ_DETECT_ENABLE_SOURCE), 
 .PMA_CH0_REG_SET_DIVSEL_REF(PMA_CH0_REG_SET_DIVSEL_REF), 
 .PMA_CH0_REG_SET_DIVSEL45_FB(PMA_CH0_REG_SET_DIVSEL45_FB), 
 .PMA_CH0_REG_SET_DIVSEL_FB(PMA_CH0_REG_SET_DIVSEL_FB), 
 .PMA_CH0_PLL_LOOP_EN_SETTING(PMA_CH0_PLL_LOOP_EN_SETTING), 
 .PMA_CH0_REGISTER_SET_TXPLL_DIV_ENABLE(PMA_CH0_REGISTER_SET_TXPLL_DIV_ENABLE), 
 .PMA_CH0_FORCE_RXPLL_RESET(PMA_CH0_FORCE_RXPLL_RESET), 
 .PMA_CH0_FORCE_RXPLL_ON(PMA_CH0_FORCE_RXPLL_ON), 
 .PMA_CH0_DPCK_DIV2(PMA_CH0_DPCK_DIV2), 
 .PMA_CH0_LFO_SETTING(PMA_CH0_LFO_SETTING), 
 .PMA_CH0_ALOS_COUNTER_CLOCK_SELECTION(PMA_CH0_ALOS_COUNTER_CLOCK_SELECTION), 
 .PMA_CH0_RX_BIAS_CURRENT_ADJUSTMENT(PMA_CH0_RX_BIAS_CURRENT_ADJUSTMENT), 
 .PMA_CH0_OOB_ENTER_DELAY_SETTING(PMA_CH0_OOB_ENTER_DELAY_SETTING), 
 .PMA_CH0_ALOS_LOW_TO_HIGH_COUNTER_SETTING(PMA_CH0_ALOS_LOW_TO_HIGH_COUNTER_SETTING), 
 .PMA_CH0_ENABLE_ALOS_RESULT_AUTOMATICALLY_ENABLE_CHANNEL(PMA_CH0_ENABLE_ALOS_RESULT_AUTOMATICALLY_ENABLE_CHANNEL), 
 .PMA_CH0_ALOS_EXIT_COUNTER_CLOCK_DIVIDER(PMA_CH0_ALOS_EXIT_COUNTER_CLOCK_DIVIDER), 
 .PMA_CH0_OOB_OSCILATER_FREQUENCY_SETTING(PMA_CH0_OOB_OSCILATER_FREQUENCY_SETTING), 
 .PMA_CH0_FORCE_OOB(PMA_CH0_FORCE_OOB), 
 .PMA_CH0_OOB_VTH_SET(PMA_CH0_OOB_VTH_SET), 
 .PMA_CH0_FORCE_DET_FORCE_ALOS_LOW(PMA_CH0_FORCE_DET_FORCE_ALOS_LOW), 
 .PMA_CH0_ALOS_THRESHOLD_VOLTAGE(PMA_CH0_ALOS_THRESHOLD_VOLTAGE), 
 .PMA_CH0_WAKEUP_VCM_RX_COMMON_MODE_VOLTAGE(PMA_CH0_WAKEUP_VCM_RX_COMMON_MODE_VOLTAGE), 
 .PMA_CH0_REGR_NEGATIVE_HYSTERESIS_SETTING(PMA_CH0_REGR_NEGATIVE_HYSTERESIS_SETTING), 
 .PMA_CH0_REGL_POSITIVE_HYSTERESIS_SETTING(PMA_CH0_REGL_POSITIVE_HYSTERESIS_SETTING), 
 .PMA_CH0_REG_EN(PMA_CH0_REG_EN), 
 .PMA_CH0_REGREF_SEL(PMA_CH0_REGREF_SEL), 
 .PMA_CH0_DC496(PMA_CH0_DC496), 
 .PMA_CH0_EQ2_AC_VAR_SETTING(PMA_CH0_EQ2_AC_VAR_SETTING), 
 .PMA_CH0_EQ2_AC_RES_SETTING(PMA_CH0_EQ2_AC_RES_SETTING), 
 .PMA_CH0_EQ2_DC_RESTOP_SETTING(PMA_CH0_EQ2_DC_RESTOP_SETTING), 
 .PMA_CH0_EQ1_DC_RESTOP_SETTING(PMA_CH0_EQ1_DC_RESTOP_SETTING), 
 .PMA_CH0_EQ1_AC_VAR_SETTING(PMA_CH0_EQ1_AC_VAR_SETTING), 
 .PMA_CH0_EQ2_CURRENT_SETTING(PMA_CH0_EQ2_CURRENT_SETTING), 
 .PMA_CH0_EQ1_AC_RES_SETTING(PMA_CH0_EQ1_AC_RES_SETTING), 
 .PMA_CH0_EQ1_CURRENT_SETTING(PMA_CH0_EQ1_CURRENT_SETTING), 
 .PMA_CH0_RPLUS(PMA_CH0_RPLUS), 
 .PMA_CH0_RMINUS(PMA_CH0_RMINUS), 
 .PMA_CH0_RVALSET(PMA_CH0_RVALSET), 
 .PMA_CH0_RTERM(PMA_CH0_RTERM), 
 .PMA_CH0_DCFB_EN(PMA_CH0_DCFB_EN), 
 .PMA_CH0_DCCOUP(PMA_CH0_DCCOUP), 
 .PMA_CH0_3G(PMA_CH0_3G), 
 .PMA_CH1_TXDATA_WIDTH(PMA_CH1_TXDATA_WIDTH), 
 .PMA_CH1_TX_TESTPATTERN(PMA_CH1_TX_TESTPATTERN), 
 .PMA_CH1_TESTPATTERN_O_ENABLE(PMA_CH1_TESTPATTERN_O_ENABLE), 
 .PMA_CH1_DISABLE_BSMODE_DRVAMP(PMA_CH1_DISABLE_BSMODE_DRVAMP), 
 .PMA_CH1_FORCE_BIST_ENABLE(PMA_CH1_FORCE_BIST_ENABLE), 
 .PMA_CH1_FORCE_ELECTRICAL_IDLE(PMA_CH1_FORCE_ELECTRICAL_IDLE), 
 .PMA_CH1_FORCE_RXDCT_ENABLE(PMA_CH1_FORCE_RXDCT_ENABLE), 
 .PMA_CH1_FORCE_EXTLB_ENABLE(PMA_CH1_FORCE_EXTLB_ENABLE), 
 .PMA_CH1_DISABLE_LANE_SYNC(PMA_CH1_DISABLE_LANE_SYNC), 
 .PMA_CH1_DISABLE_ELECTRICAL_IDLE(PMA_CH1_DISABLE_ELECTRICAL_IDLE), 
 .PMA_CH1_DISABLE_RXDCT_ENABLE(PMA_CH1_DISABLE_RXDCT_ENABLE), 
 .PMA_CH1_DISABLE_EXTLB_ENABLE(PMA_CH1_DISABLE_EXTLB_ENABLE), 
 .PMA_CH1_DISABLE_LOW_SPEED_PATH_ENABLE(PMA_CH1_DISABLE_LOW_SPEED_PATH_ENABLE), 
 .PMA_CH1_FORCE_LANE_ENABLE(PMA_CH1_FORCE_LANE_ENABLE), 
 .PMA_CH1_FORCE_LANE_RESETB_DISABLE(PMA_CH1_FORCE_LANE_RESETB_DISABLE), 
 .PMA_CH1_RXDCT_LGBW_ENABLE(PMA_CH1_RXDCT_LGBW_ENABLE), 
 .PMA_CH1_RXDCT_VTH(PMA_CH1_RXDCT_VTH), 
 .PMA_CH1_DE_EMPHASIS_ADDITIONAL_CONTROL(PMA_CH1_DE_EMPHASIS_ADDITIONAL_CONTROL), 
 .PMA_CH1_DRV_RTERM_CONTROL(PMA_CH1_DRV_RTERM_CONTROL), 
 .PMA_CH1_FDRV_AMP_CONTROL(PMA_CH1_FDRV_AMP_CONTROL), 
 .PMA_CH1_PREPC_AMP_CONTROL(PMA_CH1_PREPC_AMP_CONTROL), 
 .PMA_CH1_PREMC_AMP_CONTROL(PMA_CH1_PREMC_AMP_CONTROL), 
 .PMA_CH1_SER_AMP_CONTROL(PMA_CH1_SER_AMP_CONTROL), 
 .PMA_CH1_PFD_LOOP_RESISTOR_SETTING(PMA_CH1_PFD_LOOP_RESISTOR_SETTING), 
 .PMA_CH1_PD_LOOP_RESISTOR_SETTING(PMA_CH1_PD_LOOP_RESISTOR_SETTING), 
 .PMA_CH1_CDR_TEST_OUT_SELECT(PMA_CH1_CDR_TEST_OUT_SELECT), 
 .PMA_CH1_PI_DIV1_BP(PMA_CH1_PI_DIV1_BP), 
 .PMA_CH1_PI_TEST_FOR_CKI(PMA_CH1_PI_TEST_FOR_CKI), 
 .PMA_CH1_PI_CURRENT_SETTING(PMA_CH1_PI_CURRENT_SETTING), 
 .PMA_CH1_PI_FREQUENCY_SETTING(PMA_CH1_PI_FREQUENCY_SETTING), 
 .PMA_CH1_TEST_OUT_SELECT_FOR_RCK(PMA_CH1_TEST_OUT_SELECT_FOR_RCK), 
 .PMA_CH1_TEST_OUT_SELECT_SOURCE(PMA_CH1_TEST_OUT_SELECT_SOURCE), 
 .PMA_CH1_TEST_DATA_OUT_SELECT_SOURCE(PMA_CH1_TEST_DATA_OUT_SELECT_SOURCE), 
 .PMA_CH1_TEST_CK_OUT_SELECT_SOURCE(PMA_CH1_TEST_CK_OUT_SELECT_SOURCE), 
 .PMA_CH1_ENABLE_SLIP1UI_MODULE(PMA_CH1_ENABLE_SLIP1UI_MODULE), 
 .PMA_CH1_PN_SWAP_ENABLE(PMA_CH1_PN_SWAP_ENABLE), 
 .PMA_CH1_SIPO_BIT_SETTING(PMA_CH1_SIPO_BIT_SETTING), 
 .PMA_CH1_OOB_EN(PMA_CH1_OOB_EN), 
 .PMA_CH1_ALOS_EN(PMA_CH1_ALOS_EN), 
 .PMA_CH1_LFMODE(PMA_CH1_LFMODE), 
 .PMA_CH1_TSO_HS_SEL(PMA_CH1_TSO_HS_SEL), 
 .PMA_CH1_LX_SELLC(PMA_CH1_LX_SELLC), 
 .PMA_CH1_LX_RXPLL_DIVSEL45_FB(PMA_CH1_LX_RXPLL_DIVSEL45_FB), 
 .PMA_CH1_LX_RXPLL_DIVSEL_FB(PMA_CH1_LX_RXPLL_DIVSEL_FB), 
 .PMA_CH1_LX_RXPLL_DIVSEL_REF(PMA_CH1_LX_RXPLL_DIVSEL_REF), 
 .PMA_CH1_PICODE(PMA_CH1_PICODE), 
 .PMA_CH1_RX_REFCK_SEL(PMA_CH1_RX_REFCK_SEL), 
 .PMA_CH1_PFDLPEN_REGISTER_CONTROL_ENABLE(PMA_CH1_PFDLPEN_REGISTER_CONTROL_ENABLE), 
 .PMA_CH1_PFDLPEN_REGISTER_SETTING(PMA_CH1_PFDLPEN_REGISTER_SETTING), 
 .PMA_CH1_PDLPEN_REGISTER_CONTROL_ENABLE(PMA_CH1_PDLPEN_REGISTER_CONTROL_ENABLE), 
 .PMA_CH1_PDLPEN_REGISTER_SETTING(PMA_CH1_PDLPEN_REGISTER_SETTING), 
 .PMA_CH1_DIV_CHANGE_ENABLE_DELAY_TIMER(PMA_CH1_DIV_CHANGE_ENABLE_DELAY_TIMER), 
 .PMA_CH1_DIV_CHANGE_ENABLE_SIGNAL_GATING(PMA_CH1_DIV_CHANGE_ENABLE_SIGNAL_GATING), 
 .PMA_CH1_CDR_ALIGN_REGISTER_SETTING_VALUE(PMA_CH1_CDR_ALIGN_REGISTER_SETTING_VALUE), 
 .PMA_CH1_FORCE_CDR_ALIGN_ENABLE(PMA_CH1_FORCE_CDR_ALIGN_ENABLE), 
 .PMA_CH1_SELLC_REGISTER_SETTING_VALUE(PMA_CH1_SELLC_REGISTER_SETTING_VALUE), 
 .PMA_CH1_SELLC_CONTROL_BY_REGISTER(PMA_CH1_SELLC_CONTROL_BY_REGISTER), 
 .PMA_CH1_REG_PLLI_LDO_VREF_SETTING(PMA_CH1_REG_PLLI_LDO_VREF_SETTING), 
 .PMA_CH1_REG_PLLI_LDO_BYPASS_CURRENT(PMA_CH1_REG_PLLI_LDO_BYPASS_CURRENT), 
 .PMA_CH1_REG_PLL_HSTEST_ENABLE(PMA_CH1_REG_PLL_HSTEST_ENABLE), 
 .PMA_CH1_REG_PLL_ISNK_CURRENT_CONTROL(PMA_CH1_REG_PLL_ISNK_CURRENT_CONTROL), 
 .PMA_CH1_REG_PLL_PFD_LOOP_CP0_CURRENT_SETTING(PMA_CH1_REG_PLL_PFD_LOOP_CP0_CURRENT_SETTING), 
 .PMA_CH1_REG_PLL_PD_LOOP_PLLGM_SETTING(PMA_CH1_REG_PLL_PD_LOOP_PLLGM_SETTING), 
 .PMA_CH1_REG_PLL_PFD_LOOP_CP1_CURRENT_SETTING(PMA_CH1_REG_PLL_PFD_LOOP_CP1_CURRENT_SETTING), 
 .PMA_CH1_REG_PLL_CP0_BIAS_CONTROL(PMA_CH1_REG_PLL_CP0_BIAS_CONTROL), 
 .PMA_CH1_REG_PLL_PD_LOOP_CP0_CURRENT_SETTING(PMA_CH1_REG_PLL_PD_LOOP_CP0_CURRENT_SETTING), 
 .PMA_CH1_REG_PLL_CP1_BIAS_CONTROL(PMA_CH1_REG_PLL_CP1_BIAS_CONTROL), 
 .PMA_CH1_REG_PLL_PD_LOOP_CP1_CURRENT_SETTING(PMA_CH1_REG_PLL_PD_LOOP_CP1_CURRENT_SETTING), 
 .PMA_CH1_REG_PLL_CP0_CURRENT_SETTING(PMA_CH1_REG_PLL_CP0_CURRENT_SETTING), 
 .PMA_CH1_REG_PLL_CP1_CURRENT_SETTING(PMA_CH1_REG_PLL_CP1_CURRENT_SETTING), 
 .PMA_CH1_REG_PLL_GM1_CURRENT_SETTING(PMA_CH1_REG_PLL_GM1_CURRENT_SETTING), 
 .PMA_CH1_REG_PLL_LC_BF2_CURRENT_SETTING(PMA_CH1_REG_PLL_LC_BF2_CURRENT_SETTING), 
 .PMA_CH1_REG_PLL_LC_BF2_CURRENT_SETTING_LOW(PMA_CH1_REG_PLL_LC_BF2_CURRENT_SETTING_LOW), 
 .PMA_CH1_REG_PLL_REG_CUR(PMA_CH1_REG_PLL_REG_CUR), 
 .PMA_CH1_REG_PLL_LCCUR(PMA_CH1_REG_PLL_LCCUR), 
 .PMA_CH1_REG_PLL_LCOBAS(PMA_CH1_REG_PLL_LCOBAS), 
 .PMA_CH1_REG_PLL_FB_CK_TEST_OUT_ENABLE(PMA_CH1_REG_PLL_FB_CK_TEST_OUT_ENABLE), 
 .PMA_CH1_CDR_ALIGN_TIMER(PMA_CH1_CDR_ALIGN_TIMER), 
 .PMA_CH1_CALIB_WAIT(PMA_CH1_CALIB_WAIT), 
 .PMA_CH1_CALIB_TIMER(PMA_CH1_CALIB_TIMER), 
 .PMA_CH1_TOT_RANGE(PMA_CH1_TOT_RANGE), 
 .PMA_CH1_SUB_RANGE(PMA_CH1_SUB_RANGE), 
 .PMA_CH1_OVLP(PMA_CH1_OVLP), 
 .PMA_CH1_BIST_WAIT(PMA_CH1_BIST_WAIT), 
 .PMA_CH1_BIST_TIMER(PMA_CH1_BIST_TIMER), 
 .PMA_CH1_BAND_LB(PMA_CH1_BAND_LB), 
 .PMA_CH1_BAND_HB(PMA_CH1_BAND_HB), 
 .PMA_CH1_FREQ_LOCK_ACCURACY(PMA_CH1_FREQ_LOCK_ACCURACY), 
 .PMA_CH1_REG_SET_LC_BAND(PMA_CH1_REG_SET_LC_BAND), 
 .PMA_CH1_REG_SET_VCODIV(PMA_CH1_REG_SET_VCODIV), 
 .PMA_CH1_REGISTER_SET_VCODIV_BAND_ENABLE(PMA_CH1_REGISTER_SET_VCODIV_BAND_ENABLE), 
 .PMA_CH1_REG_SET_PLL_LOCK(PMA_CH1_REG_SET_PLL_LOCK), 
 .PMA_CH1_REGISTER_SET_PLL_LOCK_ENABLE(PMA_CH1_REGISTER_SET_PLL_LOCK_ENABLE), 
 .PMA_CH1_REG_SET_VCO_HI(PMA_CH1_REG_SET_VCO_HI), 
 .PMA_CH1_REG_SET_VCO_LO(PMA_CH1_REG_SET_VCO_LO), 
 .PMA_CH1_REGISTER_SET_VCO_HI_VCO_LO_ENABLE(PMA_CH1_REGISTER_SET_VCO_HI_VCO_LO_ENABLE), 
 .PMA_CH1_FORCE_LC_PLL_LOOP_EN_H(PMA_CH1_FORCE_LC_PLL_LOOP_EN_H), 
 .PMA_CH1_FORCE_LC_PLL_LOOP_EN_L(PMA_CH1_FORCE_LC_PLL_LOOP_EN_L), 
 .PMA_CH1_VCO_DIV_CALI_BYPASS(PMA_CH1_VCO_DIV_CALI_BYPASS), 
 .PMA_CH1_BIST_EN(PMA_CH1_BIST_EN), 
 .PMA_CH1_PLL_LOOP_EN_SETTING_FROM_REGISTER_ENABLE(PMA_CH1_PLL_LOOP_EN_SETTING_FROM_REGISTER_ENABLE), 
 .PMA_CH1_FREQ_DETECT_ENABLE_SOURCE(PMA_CH1_FREQ_DETECT_ENABLE_SOURCE), 
 .PMA_CH1_REG_SET_DIVSEL_REF(PMA_CH1_REG_SET_DIVSEL_REF), 
 .PMA_CH1_REG_SET_DIVSEL45_FB(PMA_CH1_REG_SET_DIVSEL45_FB), 
 .PMA_CH1_REG_SET_DIVSEL_FB(PMA_CH1_REG_SET_DIVSEL_FB), 
 .PMA_CH1_PLL_LOOP_EN_SETTING(PMA_CH1_PLL_LOOP_EN_SETTING), 
 .PMA_CH1_REGISTER_SET_TXPLL_DIV_ENABLE(PMA_CH1_REGISTER_SET_TXPLL_DIV_ENABLE), 
 .PMA_CH1_FORCE_RXPLL_RESET(PMA_CH1_FORCE_RXPLL_RESET), 
 .PMA_CH1_FORCE_RXPLL_ON(PMA_CH1_FORCE_RXPLL_ON), 
 .PMA_CH1_DPCK_DIV2(PMA_CH1_DPCK_DIV2), 
 .PMA_CH1_LFO_SETTING(PMA_CH1_LFO_SETTING), 
 .PMA_CH1_ALOS_COUNTER_CLOCK_SELECTION(PMA_CH1_ALOS_COUNTER_CLOCK_SELECTION), 
 .PMA_CH1_RX_BIAS_CURRENT_ADJUSTMENT(PMA_CH1_RX_BIAS_CURRENT_ADJUSTMENT), 
 .PMA_CH1_OOB_ENTER_DELAY_SETTING(PMA_CH1_OOB_ENTER_DELAY_SETTING), 
 .PMA_CH1_ALOS_LOW_TO_HIGH_COUNTER_SETTING(PMA_CH1_ALOS_LOW_TO_HIGH_COUNTER_SETTING), 
 .PMA_CH1_ENABLE_ALOS_RESULT_AUTOMATICALLY_ENABLE_CHANNEL(PMA_CH1_ENABLE_ALOS_RESULT_AUTOMATICALLY_ENABLE_CHANNEL), 
 .PMA_CH1_ALOS_EXIT_COUNTER_CLOCK_DIVIDER(PMA_CH1_ALOS_EXIT_COUNTER_CLOCK_DIVIDER), 
 .PMA_CH1_OOB_OSCILATER_FREQUENCY_SETTING(PMA_CH1_OOB_OSCILATER_FREQUENCY_SETTING), 
 .PMA_CH1_FORCE_OOB(PMA_CH1_FORCE_OOB), 
 .PMA_CH1_OOB_VTH_SET(PMA_CH1_OOB_VTH_SET), 
 .PMA_CH1_FORCE_DET_FORCE_ALOS_LOW(PMA_CH1_FORCE_DET_FORCE_ALOS_LOW), 
 .PMA_CH1_ALOS_THRESHOLD_VOLTAGE(PMA_CH1_ALOS_THRESHOLD_VOLTAGE), 
 .PMA_CH1_WAKEUP_VCM_RX_COMMON_MODE_VOLTAGE(PMA_CH1_WAKEUP_VCM_RX_COMMON_MODE_VOLTAGE), 
 .PMA_CH1_REGR_NEGATIVE_HYSTERESIS_SETTING(PMA_CH1_REGR_NEGATIVE_HYSTERESIS_SETTING), 
 .PMA_CH1_REGL_POSITIVE_HYSTERESIS_SETTING(PMA_CH1_REGL_POSITIVE_HYSTERESIS_SETTING), 
 .PMA_CH1_REG_EN(PMA_CH1_REG_EN), 
 .PMA_CH1_REGREF_SEL(PMA_CH1_REGREF_SEL), 
 .PMA_CH1_DC496(PMA_CH1_DC496), 
 .PMA_CH1_EQ2_AC_VAR_SETTING(PMA_CH1_EQ2_AC_VAR_SETTING), 
 .PMA_CH1_EQ2_AC_RES_SETTING(PMA_CH1_EQ2_AC_RES_SETTING), 
 .PMA_CH1_EQ2_DC_RESTOP_SETTING(PMA_CH1_EQ2_DC_RESTOP_SETTING), 
 .PMA_CH1_EQ1_DC_RESTOP_SETTING(PMA_CH1_EQ1_DC_RESTOP_SETTING), 
 .PMA_CH1_EQ1_AC_VAR_SETTING(PMA_CH1_EQ1_AC_VAR_SETTING), 
 .PMA_CH1_EQ2_CURRENT_SETTING(PMA_CH1_EQ2_CURRENT_SETTING), 
 .PMA_CH1_EQ1_AC_RES_SETTING(PMA_CH1_EQ1_AC_RES_SETTING), 
 .PMA_CH1_EQ1_CURRENT_SETTING(PMA_CH1_EQ1_CURRENT_SETTING), 
 .PMA_CH1_RPLUS(PMA_CH1_RPLUS), 
 .PMA_CH1_RMINUS(PMA_CH1_RMINUS), 
 .PMA_CH1_RVALSET(PMA_CH1_RVALSET), 
 .PMA_CH1_RTERM(PMA_CH1_RTERM), 
 .PMA_CH1_DCFB_EN(PMA_CH1_DCFB_EN), 
 .PMA_CH1_DCCOUP(PMA_CH1_DCCOUP), 
 .PMA_CH1_3G(PMA_CH1_3G), 
 .PMA_CH2_TXDATA_WIDTH(PMA_CH2_TXDATA_WIDTH), 
 .PMA_CH2_TX_TESTPATTERN(PMA_CH2_TX_TESTPATTERN), 
 .PMA_CH2_TESTPATTERN_O_ENABLE(PMA_CH2_TESTPATTERN_O_ENABLE), 
 .PMA_CH2_DISABLE_BSMODE_DRVAMP(PMA_CH2_DISABLE_BSMODE_DRVAMP), 
 .PMA_CH2_FORCE_BIST_ENABLE(PMA_CH2_FORCE_BIST_ENABLE), 
 .PMA_CH2_FORCE_ELECTRICAL_IDLE(PMA_CH2_FORCE_ELECTRICAL_IDLE), 
 .PMA_CH2_FORCE_RXDCT_ENABLE(PMA_CH2_FORCE_RXDCT_ENABLE), 
 .PMA_CH2_FORCE_EXTLB_ENABLE(PMA_CH2_FORCE_EXTLB_ENABLE), 
 .PMA_CH2_DISABLE_LANE_SYNC(PMA_CH2_DISABLE_LANE_SYNC), 
 .PMA_CH2_DISABLE_ELECTRICAL_IDLE(PMA_CH2_DISABLE_ELECTRICAL_IDLE), 
 .PMA_CH2_DISABLE_RXDCT_ENABLE(PMA_CH2_DISABLE_RXDCT_ENABLE), 
 .PMA_CH2_DISABLE_EXTLB_ENABLE(PMA_CH2_DISABLE_EXTLB_ENABLE), 
 .PMA_CH2_DISABLE_LOW_SPEED_PATH_ENABLE(PMA_CH2_DISABLE_LOW_SPEED_PATH_ENABLE), 
 .PMA_CH2_FORCE_LANE_ENABLE(PMA_CH2_FORCE_LANE_ENABLE), 
 .PMA_CH2_FORCE_LANE_RESETB_DISABLE(PMA_CH2_FORCE_LANE_RESETB_DISABLE), 
 .PMA_CH2_RXDCT_LGBW_ENABLE(PMA_CH2_RXDCT_LGBW_ENABLE), 
 .PMA_CH2_RXDCT_VTH(PMA_CH2_RXDCT_VTH), 
 .PMA_CH2_DE_EMPHASIS_ADDITIONAL_CONTROL(PMA_CH2_DE_EMPHASIS_ADDITIONAL_CONTROL), 
 .PMA_CH2_DRV_RTERM_CONTROL(PMA_CH2_DRV_RTERM_CONTROL), 
 .PMA_CH2_FDRV_AMP_CONTROL(PMA_CH2_FDRV_AMP_CONTROL), 
 .PMA_CH2_PREPC_AMP_CONTROL(PMA_CH2_PREPC_AMP_CONTROL), 
 .PMA_CH2_PREMC_AMP_CONTROL(PMA_CH2_PREMC_AMP_CONTROL), 
 .PMA_CH2_SER_AMP_CONTROL(PMA_CH2_SER_AMP_CONTROL), 
 .PMA_CH2_PFD_LOOP_RESISTOR_SETTING(PMA_CH2_PFD_LOOP_RESISTOR_SETTING), 
 .PMA_CH2_PD_LOOP_RESISTOR_SETTING(PMA_CH2_PD_LOOP_RESISTOR_SETTING), 
 .PMA_CH2_CDR_TEST_OUT_SELECT(PMA_CH2_CDR_TEST_OUT_SELECT), 
 .PMA_CH2_PI_DIV1_BP(PMA_CH2_PI_DIV1_BP), 
 .PMA_CH2_PI_TEST_FOR_CKI(PMA_CH2_PI_TEST_FOR_CKI), 
 .PMA_CH2_PI_CURRENT_SETTING(PMA_CH2_PI_CURRENT_SETTING), 
 .PMA_CH2_PI_FREQUENCY_SETTING(PMA_CH2_PI_FREQUENCY_SETTING), 
 .PMA_CH2_TEST_OUT_SELECT_FOR_RCK(PMA_CH2_TEST_OUT_SELECT_FOR_RCK), 
 .PMA_CH2_TEST_OUT_SELECT_SOURCE(PMA_CH2_TEST_OUT_SELECT_SOURCE), 
 .PMA_CH2_TEST_DATA_OUT_SELECT_SOURCE(PMA_CH2_TEST_DATA_OUT_SELECT_SOURCE), 
 .PMA_CH2_TEST_CK_OUT_SELECT_SOURCE(PMA_CH2_TEST_CK_OUT_SELECT_SOURCE), 
 .PMA_CH2_ENABLE_SLIP1UI_MODULE(PMA_CH2_ENABLE_SLIP1UI_MODULE), 
 .PMA_CH2_PN_SWAP_ENABLE(PMA_CH2_PN_SWAP_ENABLE), 
 .PMA_CH2_SIPO_BIT_SETTING(PMA_CH2_SIPO_BIT_SETTING), 
 .PMA_CH2_OOB_EN(PMA_CH2_OOB_EN), 
 .PMA_CH2_ALOS_EN(PMA_CH2_ALOS_EN), 
 .PMA_CH2_LFMODE(PMA_CH2_LFMODE), 
 .PMA_CH2_TSO_HS_SEL(PMA_CH2_TSO_HS_SEL), 
 .PMA_CH2_LX_SELLC(PMA_CH2_LX_SELLC), 
 .PMA_CH2_LX_RXPLL_DIVSEL45_FB(PMA_CH2_LX_RXPLL_DIVSEL45_FB), 
 .PMA_CH2_LX_RXPLL_DIVSEL_FB(PMA_CH2_LX_RXPLL_DIVSEL_FB), 
 .PMA_CH2_LX_RXPLL_DIVSEL_REF(PMA_CH2_LX_RXPLL_DIVSEL_REF), 
 .PMA_CH2_PICODE(PMA_CH2_PICODE), 
 .PMA_CH2_RX_REFCK_SEL(PMA_CH2_RX_REFCK_SEL), 
 .PMA_CH2_PFDLPEN_REGISTER_CONTROL_ENABLE(PMA_CH2_PFDLPEN_REGISTER_CONTROL_ENABLE), 
 .PMA_CH2_PFDLPEN_REGISTER_SETTING(PMA_CH2_PFDLPEN_REGISTER_SETTING), 
 .PMA_CH2_PDLPEN_REGISTER_CONTROL_ENABLE(PMA_CH2_PDLPEN_REGISTER_CONTROL_ENABLE), 
 .PMA_CH2_PDLPEN_REGISTER_SETTING(PMA_CH2_PDLPEN_REGISTER_SETTING), 
 .PMA_CH2_DIV_CHANGE_ENABLE_DELAY_TIMER(PMA_CH2_DIV_CHANGE_ENABLE_DELAY_TIMER), 
 .PMA_CH2_DIV_CHANGE_ENABLE_SIGNAL_GATING(PMA_CH2_DIV_CHANGE_ENABLE_SIGNAL_GATING), 
 .PMA_CH2_CDR_ALIGN_REGISTER_SETTING_VALUE(PMA_CH2_CDR_ALIGN_REGISTER_SETTING_VALUE), 
 .PMA_CH2_FORCE_CDR_ALIGN_ENABLE(PMA_CH2_FORCE_CDR_ALIGN_ENABLE), 
 .PMA_CH2_SELLC_REGISTER_SETTING_VALUE(PMA_CH2_SELLC_REGISTER_SETTING_VALUE), 
 .PMA_CH2_SELLC_CONTROL_BY_REGISTER(PMA_CH2_SELLC_CONTROL_BY_REGISTER), 
 .PMA_CH2_REG_PLLI_LDO_VREF_SETTING(PMA_CH2_REG_PLLI_LDO_VREF_SETTING), 
 .PMA_CH2_REG_PLLI_LDO_BYPASS_CURRENT(PMA_CH2_REG_PLLI_LDO_BYPASS_CURRENT), 
 .PMA_CH2_REG_PLL_HSTEST_ENABLE(PMA_CH2_REG_PLL_HSTEST_ENABLE), 
 .PMA_CH2_REG_PLL_ISNK_CURRENT_CONTROL(PMA_CH2_REG_PLL_ISNK_CURRENT_CONTROL), 
 .PMA_CH2_REG_PLL_PFD_LOOP_CP0_CURRENT_SETTING(PMA_CH2_REG_PLL_PFD_LOOP_CP0_CURRENT_SETTING), 
 .PMA_CH2_REG_PLL_PD_LOOP_PLLGM_SETTING(PMA_CH2_REG_PLL_PD_LOOP_PLLGM_SETTING), 
 .PMA_CH2_REG_PLL_PFD_LOOP_CP1_CURRENT_SETTING(PMA_CH2_REG_PLL_PFD_LOOP_CP1_CURRENT_SETTING), 
 .PMA_CH2_REG_PLL_CP0_BIAS_CONTROL(PMA_CH2_REG_PLL_CP0_BIAS_CONTROL), 
 .PMA_CH2_REG_PLL_PD_LOOP_CP0_CURRENT_SETTING(PMA_CH2_REG_PLL_PD_LOOP_CP0_CURRENT_SETTING), 
 .PMA_CH2_REG_PLL_CP1_BIAS_CONTROL(PMA_CH2_REG_PLL_CP1_BIAS_CONTROL), 
 .PMA_CH2_REG_PLL_PD_LOOP_CP1_CURRENT_SETTING(PMA_CH2_REG_PLL_PD_LOOP_CP1_CURRENT_SETTING), 
 .PMA_CH2_REG_PLL_CP0_CURRENT_SETTING(PMA_CH2_REG_PLL_CP0_CURRENT_SETTING), 
 .PMA_CH2_REG_PLL_CP1_CURRENT_SETTING(PMA_CH2_REG_PLL_CP1_CURRENT_SETTING), 
 .PMA_CH2_REG_PLL_GM1_CURRENT_SETTING(PMA_CH2_REG_PLL_GM1_CURRENT_SETTING), 
 .PMA_CH2_REG_PLL_LC_BF2_CURRENT_SETTING(PMA_CH2_REG_PLL_LC_BF2_CURRENT_SETTING), 
 .PMA_CH2_REG_PLL_LC_BF2_CURRENT_SETTING_LOW(PMA_CH2_REG_PLL_LC_BF2_CURRENT_SETTING_LOW), 
 .PMA_CH2_REG_PLL_REG_CUR(PMA_CH2_REG_PLL_REG_CUR), 
 .PMA_CH2_REG_PLL_LCCUR(PMA_CH2_REG_PLL_LCCUR), 
 .PMA_CH2_REG_PLL_LCOBAS(PMA_CH2_REG_PLL_LCOBAS), 
 .PMA_CH2_REG_PLL_FB_CK_TEST_OUT_ENABLE(PMA_CH2_REG_PLL_FB_CK_TEST_OUT_ENABLE), 
 .PMA_CH2_CDR_ALIGN_TIMER(PMA_CH2_CDR_ALIGN_TIMER), 
 .PMA_CH2_CALIB_WAIT(PMA_CH2_CALIB_WAIT), 
 .PMA_CH2_CALIB_TIMER(PMA_CH2_CALIB_TIMER), 
 .PMA_CH2_TOT_RANGE(PMA_CH2_TOT_RANGE), 
 .PMA_CH2_SUB_RANGE(PMA_CH2_SUB_RANGE), 
 .PMA_CH2_OVLP(PMA_CH2_OVLP), 
 .PMA_CH2_BIST_WAIT(PMA_CH2_BIST_WAIT), 
 .PMA_CH2_BIST_TIMER(PMA_CH2_BIST_TIMER), 
 .PMA_CH2_BAND_LB(PMA_CH2_BAND_LB), 
 .PMA_CH2_BAND_HB(PMA_CH2_BAND_HB), 
 .PMA_CH2_FREQ_LOCK_ACCURACY(PMA_CH2_FREQ_LOCK_ACCURACY), 
 .PMA_CH2_REG_SET_LC_BAND(PMA_CH2_REG_SET_LC_BAND), 
 .PMA_CH2_REG_SET_VCODIV(PMA_CH2_REG_SET_VCODIV), 
 .PMA_CH2_REGISTER_SET_VCODIV_BAND_ENABLE(PMA_CH2_REGISTER_SET_VCODIV_BAND_ENABLE), 
 .PMA_CH2_REG_SET_PLL_LOCK(PMA_CH2_REG_SET_PLL_LOCK), 
 .PMA_CH2_REGISTER_SET_PLL_LOCK_ENABLE(PMA_CH2_REGISTER_SET_PLL_LOCK_ENABLE), 
 .PMA_CH2_REG_SET_VCO_HI(PMA_CH2_REG_SET_VCO_HI), 
 .PMA_CH2_REG_SET_VCO_LO(PMA_CH2_REG_SET_VCO_LO), 
 .PMA_CH2_REGISTER_SET_VCO_HI_VCO_LO_ENABLE(PMA_CH2_REGISTER_SET_VCO_HI_VCO_LO_ENABLE), 
 .PMA_CH2_FORCE_LC_PLL_LOOP_EN_H(PMA_CH2_FORCE_LC_PLL_LOOP_EN_H), 
 .PMA_CH2_FORCE_LC_PLL_LOOP_EN_L(PMA_CH2_FORCE_LC_PLL_LOOP_EN_L), 
 .PMA_CH2_VCO_DIV_CALI_BYPASS(PMA_CH2_VCO_DIV_CALI_BYPASS), 
 .PMA_CH2_BIST_EN(PMA_CH2_BIST_EN), 
 .PMA_CH2_PLL_LOOP_EN_SETTING_FROM_REGISTER_ENABLE(PMA_CH2_PLL_LOOP_EN_SETTING_FROM_REGISTER_ENABLE), 
 .PMA_CH2_FREQ_DETECT_ENABLE_SOURCE(PMA_CH2_FREQ_DETECT_ENABLE_SOURCE), 
 .PMA_CH2_REG_SET_DIVSEL_REF(PMA_CH2_REG_SET_DIVSEL_REF), 
 .PMA_CH2_REG_SET_DIVSEL45_FB(PMA_CH2_REG_SET_DIVSEL45_FB), 
 .PMA_CH2_REG_SET_DIVSEL_FB(PMA_CH2_REG_SET_DIVSEL_FB), 
 .PMA_CH2_PLL_LOOP_EN_SETTING(PMA_CH2_PLL_LOOP_EN_SETTING), 
 .PMA_CH2_REGISTER_SET_TXPLL_DIV_ENABLE(PMA_CH2_REGISTER_SET_TXPLL_DIV_ENABLE), 
 .PMA_CH2_FORCE_RXPLL_RESET(PMA_CH2_FORCE_RXPLL_RESET), 
 .PMA_CH2_FORCE_RXPLL_ON(PMA_CH2_FORCE_RXPLL_ON), 
 .PMA_CH2_DPCK_DIV2(PMA_CH2_DPCK_DIV2), 
 .PMA_CH2_LFO_SETTING(PMA_CH2_LFO_SETTING), 
 .PMA_CH2_ALOS_COUNTER_CLOCK_SELECTION(PMA_CH2_ALOS_COUNTER_CLOCK_SELECTION), 
 .PMA_CH2_RX_BIAS_CURRENT_ADJUSTMENT(PMA_CH2_RX_BIAS_CURRENT_ADJUSTMENT), 
 .PMA_CH2_OOB_ENTER_DELAY_SETTING(PMA_CH2_OOB_ENTER_DELAY_SETTING), 
 .PMA_CH2_ALOS_LOW_TO_HIGH_COUNTER_SETTING(PMA_CH2_ALOS_LOW_TO_HIGH_COUNTER_SETTING), 
 .PMA_CH2_ENABLE_ALOS_RESULT_AUTOMATICALLY_ENABLE_CHANNEL(PMA_CH2_ENABLE_ALOS_RESULT_AUTOMATICALLY_ENABLE_CHANNEL), 
 .PMA_CH2_ALOS_EXIT_COUNTER_CLOCK_DIVIDER(PMA_CH2_ALOS_EXIT_COUNTER_CLOCK_DIVIDER), 
 .PMA_CH2_OOB_OSCILATER_FREQUENCY_SETTING(PMA_CH2_OOB_OSCILATER_FREQUENCY_SETTING), 
 .PMA_CH2_FORCE_OOB(PMA_CH2_FORCE_OOB), 
 .PMA_CH2_OOB_VTH_SET(PMA_CH2_OOB_VTH_SET), 
 .PMA_CH2_FORCE_DET_FORCE_ALOS_LOW(PMA_CH2_FORCE_DET_FORCE_ALOS_LOW), 
 .PMA_CH2_ALOS_THRESHOLD_VOLTAGE(PMA_CH2_ALOS_THRESHOLD_VOLTAGE), 
 .PMA_CH2_WAKEUP_VCM_RX_COMMON_MODE_VOLTAGE(PMA_CH2_WAKEUP_VCM_RX_COMMON_MODE_VOLTAGE), 
 .PMA_CH2_REGR_NEGATIVE_HYSTERESIS_SETTING(PMA_CH2_REGR_NEGATIVE_HYSTERESIS_SETTING), 
 .PMA_CH2_REGL_POSITIVE_HYSTERESIS_SETTING(PMA_CH2_REGL_POSITIVE_HYSTERESIS_SETTING), 
 .PMA_CH2_REG_EN(PMA_CH2_REG_EN), 
 .PMA_CH2_REGREF_SEL(PMA_CH2_REGREF_SEL), 
 .PMA_CH2_DC496(PMA_CH2_DC496), 
 .PMA_CH2_EQ2_AC_VAR_SETTING(PMA_CH2_EQ2_AC_VAR_SETTING), 
 .PMA_CH2_EQ2_AC_RES_SETTING(PMA_CH2_EQ2_AC_RES_SETTING), 
 .PMA_CH2_EQ2_DC_RESTOP_SETTING(PMA_CH2_EQ2_DC_RESTOP_SETTING), 
 .PMA_CH2_EQ1_DC_RESTOP_SETTING(PMA_CH2_EQ1_DC_RESTOP_SETTING), 
 .PMA_CH2_EQ1_AC_VAR_SETTING(PMA_CH2_EQ1_AC_VAR_SETTING), 
 .PMA_CH2_EQ2_CURRENT_SETTING(PMA_CH2_EQ2_CURRENT_SETTING), 
 .PMA_CH2_EQ1_AC_RES_SETTING(PMA_CH2_EQ1_AC_RES_SETTING), 
 .PMA_CH2_EQ1_CURRENT_SETTING(PMA_CH2_EQ1_CURRENT_SETTING), 
 .PMA_CH2_RPLUS(PMA_CH2_RPLUS), 
 .PMA_CH2_RMINUS(PMA_CH2_RMINUS), 
 .PMA_CH2_RVALSET(PMA_CH2_RVALSET), 
 .PMA_CH2_RTERM(PMA_CH2_RTERM), 
 .PMA_CH2_DCFB_EN(PMA_CH2_DCFB_EN), 
 .PMA_CH2_DCCOUP(PMA_CH2_DCCOUP), 
 .PMA_CH2_3G(PMA_CH2_3G), 
 .PMA_CH3_TXDATA_WIDTH(PMA_CH3_TXDATA_WIDTH), 
 .PMA_CH3_TX_TESTPATTERN(PMA_CH3_TX_TESTPATTERN), 
 .PMA_CH3_TESTPATTERN_O_ENABLE(PMA_CH3_TESTPATTERN_O_ENABLE), 
 .PMA_CH3_DISABLE_BSMODE_DRVAMP(PMA_CH3_DISABLE_BSMODE_DRVAMP), 
 .PMA_CH3_FORCE_BIST_ENABLE(PMA_CH3_FORCE_BIST_ENABLE), 
 .PMA_CH3_FORCE_ELECTRICAL_IDLE(PMA_CH3_FORCE_ELECTRICAL_IDLE), 
 .PMA_CH3_FORCE_RXDCT_ENABLE(PMA_CH3_FORCE_RXDCT_ENABLE), 
 .PMA_CH3_FORCE_EXTLB_ENABLE(PMA_CH3_FORCE_EXTLB_ENABLE), 
 .PMA_CH3_DISABLE_LANE_SYNC(PMA_CH3_DISABLE_LANE_SYNC), 
 .PMA_CH3_DISABLE_ELECTRICAL_IDLE(PMA_CH3_DISABLE_ELECTRICAL_IDLE), 
 .PMA_CH3_DISABLE_RXDCT_ENABLE(PMA_CH3_DISABLE_RXDCT_ENABLE), 
 .PMA_CH3_DISABLE_EXTLB_ENABLE(PMA_CH3_DISABLE_EXTLB_ENABLE), 
 .PMA_CH3_DISABLE_LOW_SPEED_PATH_ENABLE(PMA_CH3_DISABLE_LOW_SPEED_PATH_ENABLE), 
 .PMA_CH3_FORCE_LANE_ENABLE(PMA_CH3_FORCE_LANE_ENABLE), 
 .PMA_CH3_FORCE_LANE_RESETB_DISABLE(PMA_CH3_FORCE_LANE_RESETB_DISABLE), 
 .PMA_CH3_RXDCT_LGBW_ENABLE(PMA_CH3_RXDCT_LGBW_ENABLE), 
 .PMA_CH3_RXDCT_VTH(PMA_CH3_RXDCT_VTH), 
 .PMA_CH3_DE_EMPHASIS_ADDITIONAL_CONTROL(PMA_CH3_DE_EMPHASIS_ADDITIONAL_CONTROL), 
 .PMA_CH3_DRV_RTERM_CONTROL(PMA_CH3_DRV_RTERM_CONTROL), 
 .PMA_CH3_FDRV_AMP_CONTROL(PMA_CH3_FDRV_AMP_CONTROL), 
 .PMA_CH3_PREPC_AMP_CONTROL(PMA_CH3_PREPC_AMP_CONTROL), 
 .PMA_CH3_PREMC_AMP_CONTROL(PMA_CH3_PREMC_AMP_CONTROL), 
 .PMA_CH3_SER_AMP_CONTROL(PMA_CH3_SER_AMP_CONTROL), 
 .PMA_CH3_PFD_LOOP_RESISTOR_SETTING(PMA_CH3_PFD_LOOP_RESISTOR_SETTING), 
 .PMA_CH3_PD_LOOP_RESISTOR_SETTING(PMA_CH3_PD_LOOP_RESISTOR_SETTING), 
 .PMA_CH3_CDR_TEST_OUT_SELECT(PMA_CH3_CDR_TEST_OUT_SELECT), 
 .PMA_CH3_PI_DIV1_BP(PMA_CH3_PI_DIV1_BP), 
 .PMA_CH3_PI_TEST_FOR_CKI(PMA_CH3_PI_TEST_FOR_CKI), 
 .PMA_CH3_PI_CURRENT_SETTING(PMA_CH3_PI_CURRENT_SETTING), 
 .PMA_CH3_PI_FREQUENCY_SETTING(PMA_CH3_PI_FREQUENCY_SETTING), 
 .PMA_CH3_TEST_OUT_SELECT_FOR_RCK(PMA_CH3_TEST_OUT_SELECT_FOR_RCK), 
 .PMA_CH3_TEST_OUT_SELECT_SOURCE(PMA_CH3_TEST_OUT_SELECT_SOURCE), 
 .PMA_CH3_TEST_DATA_OUT_SELECT_SOURCE(PMA_CH3_TEST_DATA_OUT_SELECT_SOURCE), 
 .PMA_CH3_TEST_CK_OUT_SELECT_SOURCE(PMA_CH3_TEST_CK_OUT_SELECT_SOURCE), 
 .PMA_CH3_ENABLE_SLIP1UI_MODULE(PMA_CH3_ENABLE_SLIP1UI_MODULE), 
 .PMA_CH3_PN_SWAP_ENABLE(PMA_CH3_PN_SWAP_ENABLE), 
 .PMA_CH3_SIPO_BIT_SETTING(PMA_CH3_SIPO_BIT_SETTING), 
 .PMA_CH3_OOB_EN(PMA_CH3_OOB_EN), 
 .PMA_CH3_ALOS_EN(PMA_CH3_ALOS_EN), 
 .PMA_CH3_LFMODE(PMA_CH3_LFMODE), 
 .PMA_CH3_TSO_HS_SEL(PMA_CH3_TSO_HS_SEL), 
 .PMA_CH3_LX_SELLC(PMA_CH3_LX_SELLC), 
 .PMA_CH3_LX_RXPLL_DIVSEL45_FB(PMA_CH3_LX_RXPLL_DIVSEL45_FB), 
 .PMA_CH3_LX_RXPLL_DIVSEL_FB(PMA_CH3_LX_RXPLL_DIVSEL_FB), 
 .PMA_CH3_LX_RXPLL_DIVSEL_REF(PMA_CH3_LX_RXPLL_DIVSEL_REF), 
 .PMA_CH3_PICODE(PMA_CH3_PICODE), 
 .PMA_CH3_RX_REFCK_SEL(PMA_CH3_RX_REFCK_SEL), 
 .PMA_CH3_PFDLPEN_REGISTER_CONTROL_ENABLE(PMA_CH3_PFDLPEN_REGISTER_CONTROL_ENABLE), 
 .PMA_CH3_PFDLPEN_REGISTER_SETTING(PMA_CH3_PFDLPEN_REGISTER_SETTING), 
 .PMA_CH3_PDLPEN_REGISTER_CONTROL_ENABLE(PMA_CH3_PDLPEN_REGISTER_CONTROL_ENABLE), 
 .PMA_CH3_PDLPEN_REGISTER_SETTING(PMA_CH3_PDLPEN_REGISTER_SETTING), 
 .PMA_CH3_DIV_CHANGE_ENABLE_DELAY_TIMER(PMA_CH3_DIV_CHANGE_ENABLE_DELAY_TIMER), 
 .PMA_CH3_DIV_CHANGE_ENABLE_SIGNAL_GATING(PMA_CH3_DIV_CHANGE_ENABLE_SIGNAL_GATING), 
 .PMA_CH3_CDR_ALIGN_REGISTER_SETTING_VALUE(PMA_CH3_CDR_ALIGN_REGISTER_SETTING_VALUE), 
 .PMA_CH3_FORCE_CDR_ALIGN_ENABLE(PMA_CH3_FORCE_CDR_ALIGN_ENABLE), 
 .PMA_CH3_SELLC_REGISTER_SETTING_VALUE(PMA_CH3_SELLC_REGISTER_SETTING_VALUE), 
 .PMA_CH3_SELLC_CONTROL_BY_REGISTER(PMA_CH3_SELLC_CONTROL_BY_REGISTER), 
 .PMA_CH3_REG_PLLI_LDO_VREF_SETTING(PMA_CH3_REG_PLLI_LDO_VREF_SETTING), 
 .PMA_CH3_REG_PLLI_LDO_BYPASS_CURRENT(PMA_CH3_REG_PLLI_LDO_BYPASS_CURRENT), 
 .PMA_CH3_REG_PLL_HSTEST_ENABLE(PMA_CH3_REG_PLL_HSTEST_ENABLE), 
 .PMA_CH3_REG_PLL_ISNK_CURRENT_CONTROL(PMA_CH3_REG_PLL_ISNK_CURRENT_CONTROL), 
 .PMA_CH3_REG_PLL_PFD_LOOP_CP0_CURRENT_SETTING(PMA_CH3_REG_PLL_PFD_LOOP_CP0_CURRENT_SETTING), 
 .PMA_CH3_REG_PLL_PD_LOOP_PLLGM_SETTING(PMA_CH3_REG_PLL_PD_LOOP_PLLGM_SETTING), 
 .PMA_CH3_REG_PLL_PFD_LOOP_CP1_CURRENT_SETTING(PMA_CH3_REG_PLL_PFD_LOOP_CP1_CURRENT_SETTING), 
 .PMA_CH3_REG_PLL_CP0_BIAS_CONTROL(PMA_CH3_REG_PLL_CP0_BIAS_CONTROL), 
 .PMA_CH3_REG_PLL_PD_LOOP_CP0_CURRENT_SETTING(PMA_CH3_REG_PLL_PD_LOOP_CP0_CURRENT_SETTING), 
 .PMA_CH3_REG_PLL_CP1_BIAS_CONTROL(PMA_CH3_REG_PLL_CP1_BIAS_CONTROL), 
 .PMA_CH3_REG_PLL_PD_LOOP_CP1_CURRENT_SETTING(PMA_CH3_REG_PLL_PD_LOOP_CP1_CURRENT_SETTING), 
 .PMA_CH3_REG_PLL_CP0_CURRENT_SETTING(PMA_CH3_REG_PLL_CP0_CURRENT_SETTING), 
 .PMA_CH3_REG_PLL_CP1_CURRENT_SETTING(PMA_CH3_REG_PLL_CP1_CURRENT_SETTING), 
 .PMA_CH3_REG_PLL_GM1_CURRENT_SETTING(PMA_CH3_REG_PLL_GM1_CURRENT_SETTING), 
 .PMA_CH3_REG_PLL_LC_BF2_CURRENT_SETTING(PMA_CH3_REG_PLL_LC_BF2_CURRENT_SETTING), 
 .PMA_CH3_REG_PLL_LC_BF2_CURRENT_SETTING_LOW(PMA_CH3_REG_PLL_LC_BF2_CURRENT_SETTING_LOW), 
 .PMA_CH3_REG_PLL_REG_CUR(PMA_CH3_REG_PLL_REG_CUR), 
 .PMA_CH3_REG_PLL_LCCUR(PMA_CH3_REG_PLL_LCCUR), 
 .PMA_CH3_REG_PLL_LCOBAS(PMA_CH3_REG_PLL_LCOBAS), 
 .PMA_CH3_REG_PLL_FB_CK_TEST_OUT_ENABLE(PMA_CH3_REG_PLL_FB_CK_TEST_OUT_ENABLE), 
 .PMA_CH3_CDR_ALIGN_TIMER(PMA_CH3_CDR_ALIGN_TIMER), 
 .PMA_CH3_CALIB_WAIT(PMA_CH3_CALIB_WAIT), 
 .PMA_CH3_CALIB_TIMER(PMA_CH3_CALIB_TIMER), 
 .PMA_CH3_TOT_RANGE(PMA_CH3_TOT_RANGE), 
 .PMA_CH3_SUB_RANGE(PMA_CH3_SUB_RANGE), 
 .PMA_CH3_OVLP(PMA_CH3_OVLP), 
 .PMA_CH3_BIST_WAIT(PMA_CH3_BIST_WAIT), 
 .PMA_CH3_BIST_TIMER(PMA_CH3_BIST_TIMER), 
 .PMA_CH3_BAND_LB(PMA_CH3_BAND_LB), 
 .PMA_CH3_BAND_HB(PMA_CH3_BAND_HB), 
 .PMA_CH3_FREQ_LOCK_ACCURACY(PMA_CH3_FREQ_LOCK_ACCURACY), 
 .PMA_CH3_REG_SET_LC_BAND(PMA_CH3_REG_SET_LC_BAND), 
 .PMA_CH3_REG_SET_VCODIV(PMA_CH3_REG_SET_VCODIV), 
 .PMA_CH3_REGISTER_SET_VCODIV_BAND_ENABLE(PMA_CH3_REGISTER_SET_VCODIV_BAND_ENABLE), 
 .PMA_CH3_REG_SET_PLL_LOCK(PMA_CH3_REG_SET_PLL_LOCK), 
 .PMA_CH3_REGISTER_SET_PLL_LOCK_ENABLE(PMA_CH3_REGISTER_SET_PLL_LOCK_ENABLE), 
 .PMA_CH3_REG_SET_VCO_HI(PMA_CH3_REG_SET_VCO_HI), 
 .PMA_CH3_REG_SET_VCO_LO(PMA_CH3_REG_SET_VCO_LO), 
 .PMA_CH3_REGISTER_SET_VCO_HI_VCO_LO_ENABLE(PMA_CH3_REGISTER_SET_VCO_HI_VCO_LO_ENABLE), 
 .PMA_CH3_FORCE_LC_PLL_LOOP_EN_H(PMA_CH3_FORCE_LC_PLL_LOOP_EN_H), 
 .PMA_CH3_FORCE_LC_PLL_LOOP_EN_L(PMA_CH3_FORCE_LC_PLL_LOOP_EN_L), 
 .PMA_CH3_VCO_DIV_CALI_BYPASS(PMA_CH3_VCO_DIV_CALI_BYPASS), 
 .PMA_CH3_BIST_EN(PMA_CH3_BIST_EN), 
 .PMA_CH3_PLL_LOOP_EN_SETTING_FROM_REGISTER_ENABLE(PMA_CH3_PLL_LOOP_EN_SETTING_FROM_REGISTER_ENABLE), 
 .PMA_CH3_FREQ_DETECT_ENABLE_SOURCE(PMA_CH3_FREQ_DETECT_ENABLE_SOURCE), 
 .PMA_CH3_REG_SET_DIVSEL_REF(PMA_CH3_REG_SET_DIVSEL_REF), 
 .PMA_CH3_REG_SET_DIVSEL45_FB(PMA_CH3_REG_SET_DIVSEL45_FB), 
 .PMA_CH3_REG_SET_DIVSEL_FB(PMA_CH3_REG_SET_DIVSEL_FB), 
 .PMA_CH3_PLL_LOOP_EN_SETTING(PMA_CH3_PLL_LOOP_EN_SETTING), 
 .PMA_CH3_REGISTER_SET_TXPLL_DIV_ENABLE(PMA_CH3_REGISTER_SET_TXPLL_DIV_ENABLE), 
 .PMA_CH3_FORCE_RXPLL_RESET(PMA_CH3_FORCE_RXPLL_RESET), 
 .PMA_CH3_FORCE_RXPLL_ON(PMA_CH3_FORCE_RXPLL_ON), 
 .PMA_CH3_DPCK_DIV2(PMA_CH3_DPCK_DIV2), 
 .PMA_CH3_LFO_SETTING(PMA_CH3_LFO_SETTING), 
 .PMA_CH3_ALOS_COUNTER_CLOCK_SELECTION(PMA_CH3_ALOS_COUNTER_CLOCK_SELECTION), 
 .PMA_CH3_RX_BIAS_CURRENT_ADJUSTMENT(PMA_CH3_RX_BIAS_CURRENT_ADJUSTMENT), 
 .PMA_CH3_OOB_ENTER_DELAY_SETTING(PMA_CH3_OOB_ENTER_DELAY_SETTING), 
 .PMA_CH3_ALOS_LOW_TO_HIGH_COUNTER_SETTING(PMA_CH3_ALOS_LOW_TO_HIGH_COUNTER_SETTING), 
 .PMA_CH3_ENABLE_ALOS_RESULT_AUTOMATICALLY_ENABLE_CHANNEL(PMA_CH3_ENABLE_ALOS_RESULT_AUTOMATICALLY_ENABLE_CHANNEL), 
 .PMA_CH3_ALOS_EXIT_COUNTER_CLOCK_DIVIDER(PMA_CH3_ALOS_EXIT_COUNTER_CLOCK_DIVIDER), 
 .PMA_CH3_OOB_OSCILATER_FREQUENCY_SETTING(PMA_CH3_OOB_OSCILATER_FREQUENCY_SETTING), 
 .PMA_CH3_FORCE_OOB(PMA_CH3_FORCE_OOB), 
 .PMA_CH3_OOB_VTH_SET(PMA_CH3_OOB_VTH_SET), 
 .PMA_CH3_FORCE_DET_FORCE_ALOS_LOW(PMA_CH3_FORCE_DET_FORCE_ALOS_LOW), 
 .PMA_CH3_ALOS_THRESHOLD_VOLTAGE(PMA_CH3_ALOS_THRESHOLD_VOLTAGE), 
 .PMA_CH3_WAKEUP_VCM_RX_COMMON_MODE_VOLTAGE(PMA_CH3_WAKEUP_VCM_RX_COMMON_MODE_VOLTAGE), 
 .PMA_CH3_REGR_NEGATIVE_HYSTERESIS_SETTING(PMA_CH3_REGR_NEGATIVE_HYSTERESIS_SETTING), 
 .PMA_CH3_REGL_POSITIVE_HYSTERESIS_SETTING(PMA_CH3_REGL_POSITIVE_HYSTERESIS_SETTING), 
 .PMA_CH3_REG_EN(PMA_CH3_REG_EN), 
 .PMA_CH3_REGREF_SEL(PMA_CH3_REGREF_SEL), 
 .PMA_CH3_DC496(PMA_CH3_DC496), 
 .PMA_CH3_EQ2_AC_VAR_SETTING(PMA_CH3_EQ2_AC_VAR_SETTING), 
 .PMA_CH3_EQ2_AC_RES_SETTING(PMA_CH3_EQ2_AC_RES_SETTING), 
 .PMA_CH3_EQ2_DC_RESTOP_SETTING(PMA_CH3_EQ2_DC_RESTOP_SETTING), 
 .PMA_CH3_EQ1_DC_RESTOP_SETTING(PMA_CH3_EQ1_DC_RESTOP_SETTING), 
 .PMA_CH3_EQ1_AC_VAR_SETTING(PMA_CH3_EQ1_AC_VAR_SETTING), 
 .PMA_CH3_EQ2_CURRENT_SETTING(PMA_CH3_EQ2_CURRENT_SETTING), 
 .PMA_CH3_EQ1_AC_RES_SETTING(PMA_CH3_EQ1_AC_RES_SETTING), 
 .PMA_CH3_EQ1_CURRENT_SETTING(PMA_CH3_EQ1_CURRENT_SETTING), 
 .PMA_CH3_RPLUS(PMA_CH3_RPLUS), 
 .PMA_CH3_RMINUS(PMA_CH3_RMINUS), 
 .PMA_CH3_RVALSET(PMA_CH3_RVALSET), 
 .PMA_CH3_RTERM(PMA_CH3_RTERM), 
 .PMA_CH3_DCFB_EN(PMA_CH3_DCFB_EN), 
 .PMA_CH3_DCCOUP(PMA_CH3_DCCOUP), 
 .PMA_CH3_3G(PMA_CH3_3G), 
 .PMA_QUAD_TURN_ON_BANDGAP_AT_AOS_ON(PMA_QUAD_TURN_ON_BANDGAP_AT_AOS_ON), 
 .PMA_QUAD_TURN_ON_BANDGAP_AT_RX_DETECTION_ON(PMA_QUAD_TURN_ON_BANDGAP_AT_RX_DETECTION_ON), 
 .PMA_QUAD_TURN_ON_BANDGAP_AT_BOUNDARY_SCAN_ON(PMA_QUAD_TURN_ON_BANDGAP_AT_BOUNDARY_SCAN_ON), 
 .PMA_QUAD_CFG_HSST_RSTN(PMA_QUAD_CFG_HSST_RSTN), 
 .PMA_QUAD_SELECT_LANE_TCK_FOR_QUAD_SYNC(PMA_QUAD_SELECT_LANE_TCK_FOR_QUAD_SYNC), 
 .PMA_QUAD_CK_REN(PMA_QUAD_CK_REN), 
 .PMA_QUAD_C1_EN(PMA_QUAD_C1_EN), 
 .PMA_QUAD_C2_EN(PMA_QUAD_C2_EN), 
 .PMA_QUAD_CLK_DIVIDER_SETTING_FROM_25M_TO_200K(PMA_QUAD_CLK_DIVIDER_SETTING_FROM_25M_TO_200K), 
 .PMA_QUAD_ACMODE_SCANMODE_EN(PMA_QUAD_ACMODE_SCANMODE_EN), 
 .PMA_QUAD_REGISTER_ACMODE(PMA_QUAD_REGISTER_ACMODE), 
 .PMA_QUAD_REGISTER_SCANMODE(PMA_QUAD_REGISTER_SCANMODE), 
 .PMA_QUAD_REFCK2CORE_EN(PMA_QUAD_REFCK2CORE_EN), 
 .PMA_QUAD_REG_EN(PMA_QUAD_REG_EN), 
 .PMA_QUAD_REGR(PMA_QUAD_REGR), 
 .PMA_QUAD_REGL(PMA_QUAD_REGL), 
 .PMA_QUAD_DPCK_SEL(PMA_QUAD_DPCK_SEL), 
 .PMA_QUAD_TX_REFCK_SEL(PMA_QUAD_TX_REFCK_SEL), 
 .PMA_QUAD_REFCK_SRC_SEL(PMA_QUAD_REFCK_SRC_SEL), 
 .PMA_QUAD_RREFCK_PWRUP(PMA_QUAD_RREFCK_PWRUP), 
 .PMA_QUAD_REFCK_SK_SEL(PMA_QUAD_REFCK_SK_SEL),
 .PMA_QUAD_REFCK_DIV2_SEL(PMA_QUAD_REFCK_DIV2_SEL), 
 .PMA_QUAD_REFCK_TO_NQ_EN(PMA_QUAD_REFCK_TO_NQ_EN), 
 .PMA_QUAD_AUXI_ADJ(PMA_QUAD_AUXI_ADJ), 
 .PMA_QUAD_DC496(PMA_QUAD_DC496), 
 .PMA_QUAD_REG_FDET_TIMER(PMA_QUAD_REG_FDET_TIMER), 
 .PMA_QUAD_FREQ_LKO(PMA_QUAD_FREQ_LKO), 
 .PMA_QUAD_FREQ_LKI(PMA_QUAD_FREQ_LKI), 
 .PMA_QUAD_CLOCK_SRC_SEL(PMA_QUAD_CLOCK_SRC_SEL), 
 .PMA_QUAD_FRE_DET_EN(PMA_QUAD_FRE_DET_EN), 
 .PMA_QUAD_TSO_LS_SEL(PMA_QUAD_TSO_LS_SEL), 
 .PMA_QUAD_TXPLL_START(PMA_QUAD_TXPLL_START), 
 .PMA_QUAD_VCODIV(PMA_QUAD_VCODIV), 
 .PMA_QUAD_LC_BAND(PMA_QUAD_LC_BAND), 
 .PMA_QUAD_SET_VCO_HI(PMA_QUAD_SET_VCO_HI), 
 .PMA_QUAD_SET_VCO_LO(PMA_QUAD_SET_VCO_LO), 
 .PMA_QUAD_CALIB_FAIL(PMA_QUAD_CALIB_FAIL), 
 .PMA_QUAD_CALIB_DONE(PMA_QUAD_CALIB_DONE), 
 .PMA_QUAD_BIST_DONE(PMA_QUAD_BIST_DONE), 
 .PMA_QUAD_TOTRANGE_FAIL(PMA_QUAD_TOTRANGE_FAIL), 
 .PMA_QUAD_SUBRANGE_FAIL(PMA_QUAD_SUBRANGE_FAIL), 
 .PMA_QUAD_OVLP_FAIL(PMA_QUAD_OVLP_FAIL), 
 .PMA_QUAD_TXPLL_LOCK(PMA_QUAD_TXPLL_LOCK), 
 .PMA_QUAD_TXPLL_LOOP_ENABLE(PMA_QUAD_TXPLL_LOOP_ENABLE), 
 .PMA_QUAD_TXPLL_DIVSEL_REF_STA(PMA_QUAD_TXPLL_DIVSEL_REF_STA), 
 .PMA_QUAD_TXPLL_DIVSEL45_FB_STA(PMA_QUAD_TXPLL_DIVSEL45_FB_STA), 
 .PMA_QUAD_TXPLL_DIVSEL_FB_STA(PMA_QUAD_TXPLL_DIVSEL_FB_STA), 
 .PMA_QUAD_TXPLL_DIVSEL45_FB(PMA_QUAD_TXPLL_DIVSEL45_FB), 
 .PMA_QUAD_TXPLL_DIVSEL_FB(PMA_QUAD_TXPLL_DIVSEL_FB), 
 .PMA_QUAD_TXPLL_DIVSEL_REF(PMA_QUAD_TXPLL_DIVSEL_REF), 
 .PMA_QUAD_REG_DISABLE_HOLDCLK(PMA_QUAD_REG_DISABLE_HOLDCLK), 
 .PMA_QUAD_REG_DISABLE_SYNC(PMA_QUAD_REG_DISABLE_SYNC), 
 .PMA_QUAD_FORCE_OUTPUT_PLL_LOCK(PMA_QUAD_FORCE_OUTPUT_PLL_LOCK), 
 .PMA_QUAD_REGISTER_SET_SYNCTCK_SEL_ENABLE(PMA_QUAD_REGISTER_SET_SYNCTCK_SEL_ENABLE), 
 .PMA_QUAD_REG_SET_SYNCTCK_SEL(PMA_QUAD_REG_SET_SYNCTCK_SEL), 
 .PMA_QUAD_CK4TEST_OUTPUT_ENABLE(PMA_QUAD_CK4TEST_OUTPUT_ENABLE), 
 .PMA_QUAD_RSTGENBAS(PMA_QUAD_RSTGENBAS), 
 .PMA_QUAD_LCBUFBAS(PMA_QUAD_LCBUFBAS), 
 .PMA_QUAD_REGISTER_SET_CPCUR_ENABEL(PMA_QUAD_REGISTER_SET_CPCUR_ENABEL), 
 .PMA_QUAD_REG_SET_CPCUR(PMA_QUAD_REG_SET_CPCUR), 
 .PMA_QUAD_CPBAS(PMA_QUAD_CPBAS), 
 .PMA_QUAD_LCOBAS(PMA_QUAD_LCOBAS), 
 .PMA_QUAD_LCCUR(PMA_QUAD_LCCUR), 
 .PMA_QUAD_ENABLE_REGISTER_SETTING_BAND(PMA_QUAD_ENABLE_REGISTER_SETTING_BAND), 
 .PMA_QUAD_CALIB_WAIT(PMA_QUAD_CALIB_WAIT), 
 .PMA_QUAD_CALIB_TIMER(PMA_QUAD_CALIB_TIMER), 
 .PMA_QUAD_TOT_RANGE(PMA_QUAD_TOT_RANGE), 
 .PMA_QUAD_SUB_RANGE(PMA_QUAD_SUB_RANGE), 
 .PMA_QUAD_OVLP(PMA_QUAD_OVLP), 
 .PMA_QUAD_BIST_WAIT(PMA_QUAD_BIST_WAIT), 
 .PMA_QUAD_BIST_TIMER(PMA_QUAD_BIST_TIMER), 
 .PMA_QUAD_BAND_LB(PMA_QUAD_BAND_LB), 
 .PMA_QUAD_BAND_HB(PMA_QUAD_BAND_HB), 
 .PMA_QUAD_FREQ_LOCK_ACCURACY(PMA_QUAD_FREQ_LOCK_ACCURACY), 
 .PMA_QUAD_REG_SET_LC_BAND(PMA_QUAD_REG_SET_LC_BAND), 
 .PMA_QUAD_REG_SET_VCODIV(PMA_QUAD_REG_SET_VCODIV), 
 .PMA_QUAD_REGISTER_SET_VCODIV_BAND_ENABLE(PMA_QUAD_REGISTER_SET_VCODIV_BAND_ENABLE), 
 .PMA_QUAD_REG_SET_PLL_LOCK(PMA_QUAD_REG_SET_PLL_LOCK), 
 .PMA_QUAD_REGISTER_SET_PLL_LOCK_ENABLE(PMA_QUAD_REGISTER_SET_PLL_LOCK_ENABLE), 
 .PMA_QUAD_REG_SET_VCO_HI(PMA_QUAD_REG_SET_VCO_HI), 
 .PMA_QUAD_REG_SET_VCO_LO(PMA_QUAD_REG_SET_VCO_LO), 
 .PMA_QUAD_REGISTER_SET_VCO_HI_VCO_LO_ENABLE(PMA_QUAD_REGISTER_SET_VCO_HI_VCO_LO_ENABLE), 
 .PMA_QUAD_FORCE_LC_PLL_LOOP_EN_H(PMA_QUAD_FORCE_LC_PLL_LOOP_EN_H), 
 .PMA_QUAD_FORCE_LC_PLL_LOOP_EN_L(PMA_QUAD_FORCE_LC_PLL_LOOP_EN_L), 
 .PMA_QUAD_VCO_DIV_CALI_BYPASS(PMA_QUAD_VCO_DIV_CALI_BYPASS), 
 .PMA_QUAD_BIST_EN(PMA_QUAD_BIST_EN), 
 .PMA_QUAD_ENABLE_TXPLL_BIST_BLOCK_CLOCKS(PMA_QUAD_ENABLE_TXPLL_BIST_BLOCK_CLOCKS), 
 .PMA_QUAD_LF_TESTBY2(PMA_QUAD_LF_TESTBY2), 
 .PMA_QUAD_REG_SET_DIVSEL_REF(PMA_QUAD_REG_SET_DIVSEL_REF), 
 .PMA_QUAD_REG_SET_DIVSEL45_FB(PMA_QUAD_REG_SET_DIVSEL45_FB), 
 .PMA_QUAD_REG_SET_DIVSEL_FB(PMA_QUAD_REG_SET_DIVSEL_FB), 
 .PMA_QUAD_LF_TEST_EN(PMA_QUAD_LF_TEST_EN), 
 .PMA_QUAD_REGISTER_SET_TXPLL_DIV_ENABLE(PMA_QUAD_REGISTER_SET_TXPLL_DIV_ENABLE), 
 .PMA_QUAD_FORCE_TXPLL_RESET(PMA_QUAD_FORCE_TXPLL_RESET), 
 .PMA_QUAD_FORCE_TXPLL_ON(PMA_QUAD_FORCE_TXPLL_ON), 
 .CLK_ALIGNER_RX0(CLK_ALIGNER_RX0), 
 .CLK_ALIGNER_RX1(CLK_ALIGNER_RX1), 
 .CLK_ALIGNER_RX2(CLK_ALIGNER_RX2), 
 .CLK_ALIGNER_RX3(CLK_ALIGNER_RX3), 
 .CLK_ALIGNER_TX0(CLK_ALIGNER_TX0), 
 .CLK_ALIGNER_TX1(CLK_ALIGNER_TX1), 
 .CLK_ALIGNER_TX2(CLK_ALIGNER_TX2), 
 .CLK_ALIGNER_TX3(CLK_ALIGNER_TX3), 
 .DYN_DLY_EN_RX0(DYN_DLY_EN_RX0), 
 .DYN_DLY_EN_RX1(DYN_DLY_EN_RX1), 
 .DYN_DLY_EN_RX2(DYN_DLY_EN_RX2), 
 .DYN_DLY_EN_RX3(DYN_DLY_EN_RX3), 
 .DYN_DLY_EN_TX0(DYN_DLY_EN_TX0), 
 .DYN_DLY_EN_TX1(DYN_DLY_EN_TX1), 
 .DYN_DLY_EN_TX2(DYN_DLY_EN_TX2), 
 .DYN_DLY_EN_TX3(DYN_DLY_EN_TX3), 
 .DYN_DLY_SEL_RX0(DYN_DLY_SEL_RX0), 
 .DYN_DLY_SEL_RX1(DYN_DLY_SEL_RX1), 
 .DYN_DLY_SEL_RX2(DYN_DLY_SEL_RX2), 
 .DYN_DLY_SEL_RX3(DYN_DLY_SEL_RX3), 
 .DYN_DLY_SEL_TX0(DYN_DLY_SEL_TX0), 
 .DYN_DLY_SEL_TX1(DYN_DLY_SEL_TX1), 
 .DYN_DLY_SEL_TX2(DYN_DLY_SEL_TX2), 
 .DYN_DLY_SEL_TX3(DYN_DLY_SEL_TX3), 
 .CLK_ALIGNER_RSTN_RX(CLK_ALIGNER_RSTN_RX), 
 .CLK_ALIGNER_RSTN_TX(CLK_ALIGNER_RSTN_TX), 
 .LX_BISTLB_EN(LX_BISTLB_EN), 
 .LX_ELECIDLE_EN_MSB(LX_ELECIDLE_EN_MSB), 
 .LX_EXTLB_EN(LX_EXTLB_EN), 
 .LX_RXDCT_EN(LX_RXDCT_EN), 
 .LX_TX_LFMODE(LX_TX_LFMODE), 
 .RX_LANE_POWERUP(RX_LANE_POWERUP), 
 .TX_LANE_POWERUP(TX_LANE_POWERUP), 
 .PLL_RSTN(PLL_RSTN), 
 .PLLPOWERDOWN(PLLPOWERDOWN), 
 .QUAD_PWRUP(QUAD_PWRUP), 
 .GRSN_DIS(GRSN_DIS), 
 .HSST_RSTN(HSST_RSTN), 
 .CFG_RSTN(CFG_RSTN) 
)
 

GTP_HSST(

 .after_ctc_rclk_en_cout        (P_AFTER_CTC_RCLK_EN_COUT),
 .after_ctc_rclk_en_gb_cout        (P_AFTER_CTC_RCLK_EN_GB_COUT),
 .align_rx        (P_ALIGN_RX),
 .align_tx        (P_ALIGN_TX),
 .apattern_match_lsb_cout        (P_APATTERN_MATCH_LSB_COUT),
 .apattern_match_msb_cout        (P_APATTERN_MATCH_MSB_COUT),
 .apattern_seaching_proc_cout        (P_APATTERN_SEACHING_PROC_COUT),
 .apattern_status_cout        (P_APATTERN_STATUS_COUT),
 .bridge_rclk_en_cout        (P_BRIDGE_RCLK_EN_COUT),
 .bridge_tclk_en_cout        (P_BRIDGE_TCLK_EN_COUT),
 .bs_ac_ts_o        (P_BS_AC_TS_O),
 .bs_acmode_o        (P_BS_ACMODE_O),
 .bs_shift_o        (P_BS_SHIFT_O),
 .bs_tck_o        (P_BS_TCK_O),
 .bs_tdo        (P_BS_TDO),
 .bs_update_o        (P_BS_UPDATE_O),
 .bsmode_o        (P_BSMODE_O),
 .bsmode_rx_o        (P_BSMODE_RX_O),
 .cb_rclk_en_cout        (P_CB_RCLK_EN_COUT),
 .cfg_int        (P_CFG_INT),
 .cfg_rdata        (P_CFG_RDATA),
 .cfg_ready        (P_CFG_READY),
 .clk2core_rx        (P_CLK2CORE_RX),
 .clk2core_tx        (P_CLK2CORE_TX),
 .ctc_rd_fifo_cout        (P_CTC_RD_FIFO_COUT),
 .l0txn        (P_L0TXN),
 .l0txp        (P_L0TXP),
 .l1txn        (P_L1TXN),
 .l1txp        (P_L1TXP),
 .l2txn        (P_L2TXN),
 .l2txp        (P_L2TXP),
 .l3txn        (P_L3TXN),
 .l3txp        (P_L3TXP),
 .lx_alos_sta_0        (P_LX_ALOS_STA_0),
 .lx_alos_sta_1        (P_LX_ALOS_STA_1),
 .lx_alos_sta_2        (P_LX_ALOS_STA_2),
 .lx_alos_sta_3        (P_LX_ALOS_STA_3),
 .lx_cdr_align_0        (P_LX_CDR_ALIGN_0),
 .lx_cdr_align_1        (P_LX_CDR_ALIGN_1),
 .lx_cdr_align_2        (P_LX_CDR_ALIGN_2),
 .lx_cdr_align_3        (P_LX_CDR_ALIGN_3),
 .lx_lfo_0        (P_LX_LFO_0),
 .lx_lfo_1        (P_LX_LFO_1),
 .lx_lfo_2        (P_LX_LFO_2),
 .lx_lfo_3        (P_LX_LFO_3),
 .lx_oob_sta_0        (P_LX_OOB_STA_0),
 .lx_oob_sta_1        (P_LX_OOB_STA_1),
 .lx_oob_sta_2        (P_LX_OOB_STA_2),
 .lx_oob_sta_3        (P_LX_OOB_STA_3),
 .lx_rxdct_done_0        (P_LX_RXDCT_DONE_0),
 .lx_rxdct_done_1        (P_LX_RXDCT_DONE_1),
 .lx_rxdct_done_2        (P_LX_RXDCT_DONE_2),
 .lx_rxdct_done_3        (P_LX_RXDCT_DONE_3),
 .lx_rxdct_out_0        (P_LX_RXDCT_OUT_0),
 .lx_rxdct_out_1        (P_LX_RXDCT_OUT_1),
 .lx_rxdct_out_2        (P_LX_RXDCT_OUT_2),
 .lx_rxdct_out_3        (P_LX_RXDCT_OUT_3),
 .pcs_lsm_synced        (P_PCS_LSM_SYNCED),
 .pcs_rx_mcb_status        (P_PCS_RX_MCB_STATUS),
 .pcs_tclk_en_cout        (P_PCS_TCLK_EN_COUT),
 .pll_lock        (P_PLL_LOCK),
 .rdata_0        (P_RDATA_0),
 .rdata_1        (P_RDATA_1),
 .rdata_2        (P_RDATA_2),
 .rdata_3        (P_RDATA_3),
 .refck2core        (P_REFCK2CORE),
 .refck_2nmq        (P_REFCK_2NMQ),
 .refck_2npq        (P_REFCK_2NPQ),
 .rext        (P_REXT),
 .rfifo_en_after_ctc_cout        (P_RFIFO_EN_AFTER_CTC_COUT),
 .rfifo_en_after_ctc_gb_cout        (P_RFIFO_EN_AFTER_CTC_GB_COUT),
 .rfifo_en_bridge_cout        (P_RFIFO_EN_BRIDGE_COUT),
 .rfifo_en_cb_cout        (P_RFIFO_EN_CB_COUT),
 .serdes_bscan_memint_o        (P_SERDES_BSCAN_MEMINT_O),
 .skip_add_lsb_mcb_cout        (P_SKIP_ADD_LSB_MCB_COUT),
 .skip_add_mcb_cout        (P_SKIP_ADD_MCB_COUT),
 .skip_del_lsb_mcb_cout        (P_SKIP_DEL_LSB_MCB_COUT),
 .skip_del_mcb_cout        (P_SKIP_DEL_MCB_COUT),
 .test_so0        (),
 .test_so1        (),
 .test_so2        (),
 .test_so3        (),
 .test_so4        (),
 .test_so5        (),
 .test_so6        (),
 .test_so7        (),
 .tfifo_en_bridge_cout        (P_TFIFO_EN_BRIDGE_COUT),
 .tfifo_en_pcs_tx_cout        (P_TFIFO_EN_PCS_TX_COUT),
 .tso_ls_out        (P_TSO_LS_OUT),
 .apown_r        ({REP0,REP0,REP0,REP0}),
 .apown_t        (REP0),
 .apowp11_r        ({REP1,REP1,REP1,REP1}),
 .apowp11_t        (REP1),
 .pown        (REP0),
 .pown_bg        (REP0),
 .pown_nmq        (REP0),
 .pown_npq        (REP0),
 .powp11_r        ({REP1,REP1,REP1,REP1}),
 .powp11_refck        (REP1),
 .powp11_refck_nmq        (REP1),
 .powp11_refck_npq        (REP1),
 .powp11_t        (REP1),
 .powp12_r        ({REP1,REP1,REP1,REP1}),
 .powp12_t        ({REP1,REP1,REP1,REP1}),
 .vccm        (),
 .vdd33a        (REP1),
 .vssm        (),
 .ac_ts        (1'b0),
 .addr_b        (),
 .addr_t        (),
 .after_ctc_rclk_en_cin        (P_AFTER_CTC_RCLK_EN_CIN),
 .after_ctc_rclk_en_gb_cin        (P_AFTER_CTC_RCLK_EN_GB_CIN),
 .apattern_match_lsb_cin        (P_APATTERN_MATCH_LSB_CIN),
 .apattern_match_msb_cin        (P_APATTERN_MATCH_MSB_CIN),
 .apattern_seaching_proc_cin        (P_APATTERN_SEACHING_PROC_CIN),
 .apattern_status_cin        (P_APATTERN_STATUS_CIN),
 .bridge_rclk_en_cin        (P_BRIDGE_RCLK_EN_CIN),
 .bridge_tclk_en_cin        (P_BRIDGE_TCLK_EN_CIN),
 .bs_acmode        (1'b0),
 .bs_shift        (1'b1),
 .bs_tck_i        (1'b0),
 .bs_tdi        (1'b0),
 .bs_update        (1'b0),
 .bsmode        (1'b0),
 .bsmode_rx        (1'b0),
 .cb_rclk_en_cin        (P_CB_RCLK_EN_CIN),
 .ceb_adetect_en        (P_CEB_ADETECT_EN),
 .cfg_addr        (P_CFG_ADDR),
 .cfg_clk        (P_CFG_CLK),
 .cfg_enable        (P_CFG_ENABLE),
 .cfg_rstn        (P_CFG_RSTN),
 .cfg_wdata        (P_CFG_WDATA),
 .cfg_write        (P_CFG_WRITE),
 .cim_clk_aligner_rx0        (P_CIM_CLK_ALIGNER_RX0),
 .cim_clk_aligner_rx1        (P_CIM_CLK_ALIGNER_RX1),
 .cim_clk_aligner_rx2        (P_CIM_CLK_ALIGNER_RX2),
 .cim_clk_aligner_rx3        (P_CIM_CLK_ALIGNER_RX3),
 .cim_clk_aligner_tx0        (P_CIM_CLK_ALIGNER_TX0),
 .cim_clk_aligner_tx1        (P_CIM_CLK_ALIGNER_TX1),
 .cim_clk_aligner_tx2        (P_CIM_CLK_ALIGNER_TX2),
 .cim_clk_aligner_tx3        (P_CIM_CLK_ALIGNER_TX3),
 .cim_clk_dyn_dly_sel_rx        (P_CIM_CLK_DYN_DLY_SEL_RX),
 .cim_clk_dyn_dly_sel_tx        (P_CIM_CLK_DYN_DLY_SEL_TX),
 .cim_clk_start_align_rx        (P_CIM_CLK_START_ALIGN_RX),
 .cim_clk_start_align_tx        (P_CIM_CLK_START_ALIGN_TX),
 .ck25m        (P_CK25M),
 .compression_mode        (P_COMPRESSION_MODE),
 .ctc_rd_fifo_cin        (P_CTC_RD_FIFO_CIN),
 .data        (),
 .datan        (),
 .glogen        (1'b1),
 .grsn        (1'b1),
 .hsst_rstn        (P_HSST_RSTN),
 .l0rxn        (P_L0RXN),
 .l0rxp        (P_L0RXP),
 .l1rxn        (P_L1RXN),
 .l1rxp        (P_L1RXP),
 .l2rxn        (P_L2RXN),
 .l2rxp        (P_L2RXP),
 .l3rxn        (P_L3RXN),
 .l3rxp        (P_L3RXP),
 .lane_sync_en_0        (P_LANE_SYNC_EN_0),
 .lane_sync_en_1        (P_LANE_SYNC_EN_1),
 .lane_sync_en_2        (P_LANE_SYNC_EN_2),
 .lane_sync_en_3        (P_LANE_SYNC_EN_3),
 .lx_amp_ctl_0        (P_LX_AMP_CTL_0),
 .lx_amp_ctl_1        (P_LX_AMP_CTL_1),
 .lx_amp_ctl_2        (P_LX_AMP_CTL_2),
 .lx_amp_ctl_3        (P_LX_AMP_CTL_3),
 .lx_bistlb_en        (P_LX_BISTLB_EN),
 .lx_deemp_ctl_0        (P_LX_DEEMP_CTL_0),
 .lx_deemp_ctl_1        (P_LX_DEEMP_CTL_1),
 .lx_deemp_ctl_2        (P_LX_DEEMP_CTL_2),
 .lx_deemp_ctl_3        (P_LX_DEEMP_CTL_3),
 .lx_elecidle_en_0        (P_LX_ELECIDLE_EN_0),
 .lx_elecidle_en_1        (P_LX_ELECIDLE_EN_1),
 .lx_elecidle_en_2        (P_LX_ELECIDLE_EN_2),
 .lx_elecidle_en_3        (P_LX_ELECIDLE_EN_3),
 .lx_elecidle_en_msb        (P_LX_ELECIDLE_EN_MSB),
 .lx_extlb_en        (P_LX_EXTLB_EN),
 .lx_lfd_frcore_0        (P_LX_LFD_FRCORE_0),
 .lx_lfd_frcore_1        (P_LX_LFD_FRCORE_1),
 .lx_lfd_frcore_2        (P_LX_LFD_FRCORE_2),
 .lx_lfd_frcore_3        (P_LX_LFD_FRCORE_3),
 .lx_rx_ckdiv_0        (P_LX_RX_CKDIV_0),
 .lx_rx_ckdiv_1        (P_LX_RX_CKDIV_1),
 .lx_rx_ckdiv_2        (P_LX_RX_CKDIV_2),
 .lx_rx_ckdiv_3        (P_LX_RX_CKDIV_3),
 .lx_rx_ckdiv_dynsel_0        (P_LX_RX_CKDIV_DYNSEL_0),
 .lx_rx_ckdiv_dynsel_1        (P_LX_RX_CKDIV_DYNSEL_1),
 .lx_rx_ckdiv_dynsel_2        (P_LX_RX_CKDIV_DYNSEL_2),
 .lx_rx_ckdiv_dynsel_3        (P_LX_RX_CKDIV_DYNSEL_3),
 .lx_rxdct_en        (P_LX_RXDCT_EN),
 .lx_tx_lfmode        (P_LX_TX_LFMODE),
 .mcb_clk_frnq        (P_MCB_CLK_FRNQ),
 .pcs_farend_loop        (P_PCS_FAREND_LOOP),
 .pcs_mcb_ext_en        (P_PCS_MCB_EXT_EN),
 .pcs_nearend_loop        (P_PCS_NEAREND_LOOP),
 .pcs_rx_rstn_0        (P_PCS_RX_RSTN_0),
 .pcs_rx_rstn_1        (P_PCS_RX_RSTN_1),
 .pcs_rx_rstn_2        (P_PCS_RX_RSTN_2),
 .pcs_rx_rstn_3        (P_PCS_RX_RSTN_3),
 .pcs_tclk_en_cin        (P_PCS_TCLK_EN_CIN),
 .pcs_tx_rstn_0        (P_PCS_TX_RSTN_0),
 .pcs_tx_rstn_1        (P_PCS_TX_RSTN_1),
 .pcs_tx_rstn_2        (P_PCS_TX_RSTN_2),
 .pcs_tx_rstn_3        (P_PCS_TX_RSTN_3),
 .pcs_word_align_en        (P_PCS_WORD_ALIGN_EN),
 .pll_bypass        (P_PLL_BYPASS),
 .pll_ref_clk        (P_PLL_REF_CLK),
 .pll_reset        (P_PLL_RESET),
 .pll_rstn        (P_PLL_RSTN),
 .pllpowerdown        (P_PLLPOWERDOWN),
 .quad_pwrup        (P_QUAD_PWRUP),
 .refck_frnmq        (P_REFCK_FRNMQ),
 .refck_frnpq        (P_REFCK_FRNPQ),
 .refckn        (P_REFCKN),
 .refckp        (P_REFCKP),
 .rfifo_en_after_ctc_cin        (P_RFIFO_EN_AFTER_CTC_CIN),
 .rfifo_en_after_ctc_gb_cin        (P_RFIFO_EN_AFTER_CTC_GB_CIN),
 .rfifo_en_bridge_cin        (P_RFIFO_EN_BRIDGE_CIN),
 .rfifo_en_cb_cin        (P_RFIFO_EN_CB_CIN),
 .rx0_clk_fr_core        (P_RX0_CLK_FR_CORE),
 .rx1_clk_fr_core        (P_RX1_CLK_FR_CORE),
 .rx2_clk_fr_core        (P_RX2_CLK_FR_CORE),
 .rx3_clk_fr_core        (P_RX3_CLK_FR_CORE),
 .rx_lane_powerup        (P_RX_LANE_POWERUP),
 .rx_pll_rstn_0        (P_RX_PLL_RSTN_0),
 .rx_pll_rstn_1        (P_RX_PLL_RSTN_1),
 .rx_pll_rstn_2        (P_RX_PLL_RSTN_2),
 .rx_pll_rstn_3        (P_RX_PLL_RSTN_3),
 .rx_pma_rstn_0        (P_RX_PMA_RSTN_0),
 .rx_pma_rstn_1        (P_RX_PMA_RSTN_1),
 .rx_pma_rstn_2        (P_RX_PMA_RSTN_2),
 .rx_pma_rstn_3        (P_RX_PMA_RSTN_3),
 .rx_polarity_invert        (P_RX_POLARITY_INVERT),
 .rx_ref_clk_0        (P_RX_REF_CLK_0),
 .rx_ref_clk_1        (P_RX_REF_CLK_1),
 .rx_ref_clk_2        (P_RX_REF_CLK_2),
 .rx_ref_clk_3        (P_RX_REF_CLK_3),
 .sel_sync_nxq        (P_SEL_SYNC_NXQ),
 .serdes_bs_meminit        (1'b0),
 .skip_add_lsb_mcb_cin        (P_SKIP_ADD_LSB_MCB_CIN),
 .skip_add_mcb_cin        (P_SKIP_ADD_MCB_CIN),
 .skip_del_lsb_mcb_cin        (P_SKIP_DEL_LSB_MCB_CIN),
 .skip_del_mcb_cin        (P_SKIP_DEL_MCB_CIN),
 .sync_toggle        (P_SYNC_TOGGLE),
 .tdata_0        (P_TDATA_0),
 .tdata_1        (P_TDATA_1),
 .tdata_2        (P_TDATA_2),
 .tdata_3        (P_TDATA_3),
 .test_clk        (),
 .test_mode        (1'b0),
 .test_rstn        (1'b1),
 .test_se        (),
 .test_si0        (),
 .test_si1        (),
 .test_si2        (),
 .test_si3        (),
 .test_si4        (),
 .test_si5        (),
 .test_si6        (),
 .test_si7        (),
 .tfifo_en_bridge_cin        (P_TFIFO_EN_BRIDGE_CIN),
 .tfifo_en_pcs_tx_cin        (P_TFIFO_EN_PCS_TX_CIN),
 .twoquad_sync_en        (P_TWOQUAD_SYNC_EN),
 .tx0_clk_fr_core        (P_TX0_CLK_FR_CORE),
 .tx1_clk_fr_core        (P_TX1_CLK_FR_CORE),
 .tx2_clk_fr_core        (P_TX2_CLK_FR_CORE),
 .tx3_clk_fr_core        (P_TX3_CLK_FR_CORE),
 .tx_ckdiv_0        (P_TX_CKDIV_0),
 .tx_ckdiv_1        (P_TX_CKDIV_1),
 .tx_ckdiv_2        (P_TX_CKDIV_2),
 .tx_ckdiv_3        (P_TX_CKDIV_3),
 .tx_lane_powerup        (P_TX_LANE_POWERUP),
 .tx_pma_rstn_0        (P_TX_PMA_RSTN_0),
 .tx_pma_rstn_1        (P_TX_PMA_RSTN_1),
 .tx_pma_rstn_2        (P_TX_PMA_RSTN_2),
 .tx_pma_rstn_3        (P_TX_PMA_RSTN_3),
 .txckdiv_dynsel        (P_TXCKDIV_DYNSEL)

);


endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_PREADD_FIR_B.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_PREADD_FIR_B
#(
    parameter GRS_EN    = "TRUE", //"TRUE"; "FALSE"
    parameter SYNC_RST  = "FALSE", //"TRUE"; "FALSE"
    parameter INREG_EN  = "TRUE",
    parameter INREG_Z0_EN  = "TRUE",
    parameter OUTREG_EN = "TRUE",
    parameter INPUT_OP    = 4'b1111,
    parameter DYN_OP_SEL  = 4'b1111,
    parameter OPCD_DYN_SEL = 1'b0,
    parameter OPCD_CPI_SEL = 1'b0
) (
    output  [25:0] CYO,
    output         CYO_SIGNED,
    output [25:0]  CZO,
    output         CZO_SIGNED,
    output  [63:0] CPO,                  //p
    output         CPO_SIGNED,
    output  [63:0] P,

    input   CE,
    input   RST,
    input   CLK,
    input [25:0] CYI,
    input        CYI_SIGNED,
    input [25:0] CZI,
    input        CZI_SIGNED,
    input [25:0] Y0,                  //y0 ,DYIB,DYIA
    input        Y0_SIGNED,
    input [25:0] Z0,                  //z0 ,DZIB,DZIA
    input        Z0_SIGNED,            
    input [26:0] H0,                  //h0 ,DXIB,DXIA
    input        H0_SIGNED,
    input [63:0] CPI,
    input        CPI_SIGNED,
    input        S0,
    input        S1,
    input [1:0]  DYN_OP,
    input        OPCD_CPI_DYN
);

//PSE parameters
localparam [24:0] SC_PSE_Y0 = 25'b0;  //SC_PSE = 0, disable PSE, parameter bit width=25
localparam [24:0] SC_PSE_Z0 = 25'b0;  //SC_PSE = 0, disable PSE, parameter bit width=25
localparam [25:0] SC_PSE_H0 = 26'b0;  //SC_PSE = 0, disable PSE, parameter bit width=26

initial begin
    if ((GRS_EN != "TRUE") && (GRS_EN != "FALSE")) begin
        $display("GRS_EN error");
        $finish;
    end
    if ((SYNC_RST != "TRUE") && (SYNC_RST != "FALSE")) begin
        $display("SYNC_RST error");
        $finish;
    end

    if (DYN_OP_SEL[3] != 1'b1 || DYN_OP_SEL[1] != 1'b1) begin
        $display("DRC ERROR");
        $finish;
    end
end

wire [3:0] dyn_op;
reg [26:0] h0_d;
reg        h0_signed_d;
reg [25:0] y0_d;
reg [25:0] y1_d;
reg        y0_signed_d;
reg        y1_signed_d;

wire [25:0] y0_sel;
wire        y0_signed_sel;

wire [25:0] czi_sel;
wire        czi_signed_sel;

reg [25:0] z0_d;
reg        z0_signed_d;

wire [25:0] z0_sel;
wire        z0_signed_sel;

wire [26:0] preadd_1;
wire        preadd_1_signed;

wire [53:0] mult1_in1;
wire [53:0] mult1_in2;

wire [53:0] mult1;
wire        mult1_signed;

wire [63:0] sum;
wire        sum_signed;

wire [3:0]  INPUT_OP_CODE;

reg  [63:0] CPO_d;                  //p
reg         CPO_SIGNED_d;

wire [26:0]  h0_d_sel;
wire  h0_signed_d_sel;
wire [25:0]  y0_d_sel;
wire  y0_signed_d_sel;
wire [25:0]  z0_d_sel;
wire  z0_signed_d_sel;

wire global_rstn ;
wire RST_sync ;
wire RST_async;
wire rst_asyncomb ;

wire [63:0] CPI_SEL;
wire        OPCD_SEL;


assign global_rstn = GRS_EN == "TRUE" ? GRS_INST.GRSNET : 1'b1;
assign RST_sync = (SYNC_RST == "TRUE") ? RST : 1'b0;
assign RST_async = (SYNC_RST == "FALSE") ? RST : 1'b0;
assign rst_asyncomb = RST_async | (~global_rstn);

wire [25:0] Y0_PSE;
wire [25:0] Z0_PSE;
wire [26:0] H0_PSE;

INT_PSE #(.ASIZE(27),.SC_PSE(SC_PSE_H0)) U1_PSE(.A(H0),    .SIGN(H0_SIGNED),    .A_PSE(H0_PSE));
INT_PSE #(.ASIZE(26),.SC_PSE(SC_PSE_Y0)) U2_PSE(.A(y0_sel),.SIGN(y0_signed_sel),.A_PSE(Y0_PSE));
INT_PSE #(.ASIZE(26),.SC_PSE(SC_PSE_Z0)) U3_PSE(.A(z0_sel),.SIGN(z0_signed_sel),.A_PSE(Z0_PSE));

INT_REG #(.SIZE(4)) USEL (.Q(dyn_op),
    .BYPASS(INREG_EN == "TRUE" ? 1'b0 : 1'b1),
    .D({DYN_OP, S1, S0}),
    .CLK(CLK), .CE(CE), .ARST(rst_asyncomb), .SRST(RST_sync)
);
assign INPUT_OP_CODE[0] = (DYN_OP_SEL[0] ==1'b1) ? dyn_op[0] : INPUT_OP[0]; // ir_op[0,3]
assign INPUT_OP_CODE[1] = (DYN_OP_SEL[1] ==1'b1) ? dyn_op[1] : INPUT_OP[1]; // ir_op[5]
assign INPUT_OP_CODE[2] = (DYN_OP_SEL[2] ==1'b1) ? dyn_op[2] : INPUT_OP[2]; // ir_op[1,7]
assign INPUT_OP_CODE[3] = (DYN_OP_SEL[3] ==1'b1) ? dyn_op[3] : INPUT_OP[3]; // ir_op[6]

assign OPCD_SEL = (OPCD_DYN_SEL == 1'b1)?OPCD_CPI_DYN :OPCD_CPI_SEL;
assign CPI_SEL  = (OPCD_SEL == 1'b1)? 64'b0 : CPI;

initial begin
    {h0_signed_d, h0_d} = 'b0;
    {y0_signed_d, y0_d} = 'b0;
    {y1_signed_d, y1_d} = 'b0;
    {z0_signed_d, z0_d} = 'b0;
    {CPO_SIGNED_d, CPO_d} = 65'b0;
end

always @(posedge CLK or posedge rst_asyncomb)
    if (rst_asyncomb || RST_sync) begin
        {h0_signed_d, h0_d} <= 'b0;
        {y0_signed_d, y0_d} <= 'b0;
        {y1_signed_d, y1_d} <= 'b0;
        {z0_signed_d, z0_d} <= 'b0;
    end
    else if (CE) begin
        {h0_signed_d, h0_d} <= {H0_SIGNED, H0_PSE};
        {y0_signed_d, y0_d} <= {y0_signed_sel, Y0_PSE};
        {y1_signed_d, y1_d} <= {y0_signed_d_sel, y0_d_sel};
        {z0_signed_d, z0_d} <= {z0_signed_sel, Z0_PSE};
    end

assign  {h0_signed_d_sel, h0_d_sel} = (INREG_EN=="TRUE")? {h0_signed_d, h0_d} : {H0_SIGNED, H0_PSE};
assign  {y0_signed_d_sel, y0_d_sel} = (INREG_EN=="TRUE")? {y0_signed_d, y0_d} : {y0_signed_sel, Y0_PSE};
assign  {z0_signed_d_sel, z0_d_sel} = (INREG_Z0_EN=="TRUE")? {z0_signed_d, z0_d} : {z0_signed_sel, Z0_PSE};

assign {y0_signed_sel, y0_sel} = (INPUT_OP_CODE[0] == 1'b1)? {CYI_SIGNED, CYI} : {Y0_SIGNED, Y0};  // default S0 = 1 
assign {z0_signed_sel, z0_sel} = (INPUT_OP_CODE[2] == 1'b1)? {czi_signed_sel, czi_sel} : {Z0_SIGNED, Z0};

assign {czi_signed_sel, czi_sel} = (INPUT_OP_CODE[3] == 1'b0)? {CZI_SIGNED, CZI} : {CYO_SIGNED, CYO};


assign preadd_1 = {y0_d_sel[25]&y0_signed_d_sel,y0_d_sel} + {z0_d_sel[25]&z0_signed_d_sel, z0_d_sel}; 
assign preadd_1_signed = y0_signed_d_sel | z0_signed_d_sel;

reg preadd_over_flag;
always @(*)begin
    if((y0_signed_d_sel==1'b1 && y0_d_sel[25]==1'b0 && z0_signed_d_sel==1'b0 && preadd_1[26]==1'b1) || (y0_signed_d_sel==1'b0 && z0_signed_d_sel==1'b1 && z0_d_sel[25]==1'b0 && preadd_1[26]==1'b1))begin
      preadd_over_flag = 1'b1;
    end
    else begin
      preadd_over_flag = 1'b0;
    end
  end

always @(preadd_over_flag) begin
    if (preadd_over_flag==1)
    $display("Error: PREADD result is overflow!");
end

assign mult1_in1 = {{27{preadd_1_signed & preadd_1[26]}},preadd_1};
assign mult1_in2 = {{27{h0_signed_d_sel & h0_d_sel[26]}},h0_d_sel};

assign mult1 = mult1_in1 * mult1_in2;
assign mult1_signed = preadd_1_signed | h0_signed_d_sel;

assign sum = {{10{mult1_signed & mult1[53]}},mult1} + CPI_SEL;
assign sum_signed = mult1_signed | CPI_SIGNED;


always @(posedge CLK or posedge rst_asyncomb)
    if (rst_asyncomb || RST_sync) begin
        {CPO_SIGNED_d, CPO_d} <= 65'b0;
    end
    else if (CE) begin
        {CPO_SIGNED_d, CPO_d} <= {sum_signed, sum};
    end

assign {CYO_SIGNED, CYO} = (INPUT_OP_CODE[1] == 1'b1)? {y0_signed_d_sel, y0_d_sel} : {y1_signed_d, y1_d}; //default s1 = 1
assign {CZO_SIGNED, CZO} = {z0_signed_d_sel, z0_d_sel};
assign {CPO_SIGNED, CPO} = (OUTREG_EN == "TRUE") ? {CPO_SIGNED_d, CPO_d} : {sum_signed, sum};
assign P = CPO;

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2017 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_PLL_E2.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1ns/10fs
module GTP_PLL_E2 #(
    parameter real CLKIN_FREQ = 50.0,
    parameter PFDEN_EN        = "FALSE", //"TRUE"; "FALSE"
    parameter PFDEN_APB_EN    = "FALSE", //"TRUE"; "FALSE"
    parameter LOCK_MODE       = 1'b0,    //1'b0~1'b1
    parameter integer STATIC_RATIOI = 1, //1~128, step=1
    parameter integer STATIC_RATIO0 = 1, //1~128, step=1
    parameter integer STATIC_RATIO1 = 1, //1~128, step=1
    parameter integer STATIC_RATIO2 = 1, //1~128, step=1
    parameter integer STATIC_RATIO3 = 1, //1~128, step=1
    parameter integer STATIC_RATIOF = 1, //1~128, step=1
    parameter FRACN_EN          = "FALSE", //"TRUE"; "FALSE"
    parameter integer FRACN_DIV = 0,       //0~65535
    parameter PHASE_APB_EN      = "FALSE", //"TRUE"; "FALSE"
    parameter integer STATIC_PHASE0  = 0, //0~7
    parameter integer STATIC_PHASE1  = 0, //0~7
    parameter integer STATIC_PHASE2  = 0, //0~7
    parameter integer STATIC_PHASE3  = 0, //0~7
    parameter integer STATIC_CPHASE0 = 0, //0~127
    parameter integer STATIC_CPHASE1 = 0, //0~127
    parameter integer STATIC_CPHASE2 = 0, //0~127
    parameter integer STATIC_CPHASE3 = 0, //0~127
    parameter VCOCLK_BYPASS0 = "FALSE", //"TRUE"; "FALSE"
    parameter VCOCLK_BYPASS1 = "FALSE", //"TRUE"; "FALSE"
    parameter VCOCLK_BYPASS2 = "FALSE", //"TRUE"; "FALSE"
    parameter VCOCLK_BYPASS3 = "FALSE", //"TRUE"; "FALSE"
    parameter integer ODIV0_CLKIN_SEL = 0, //0~3
    parameter integer ODIV1_CLKIN_SEL = 0, //0~3
    parameter integer ODIV2_CLKIN_SEL = 0, //0~3
    parameter integer ODIV3_CLKIN_SEL = 0, //0~3
    parameter CLKOUT0_SEL = 0, //0~4
    parameter CLKOUT1_SEL = 0, //0~4
    parameter CLKOUT2_SEL = 0, //0~4
    parameter CLKOUT3_SEL = 0, //0~4
    parameter CLKOUT0_SYN_EN = "TRUE", //"TRUE"; "FALSE"
    parameter CLKOUT1_SYN_EN = "TRUE", //"TRUE"; "FALSE"
    parameter CLKOUT2_SYN_EN = "TRUE", //"TRUE"; "FALSE"
    parameter CLKOUT3_SYN_EN = "TRUE", //"TRUE"; "FALSE"
    parameter INTERNAL_FB = "CLKOUT0", //"CLKOUT0"; "CLKOUT1"; "CLKOUT2"; "CLKOUT3"; "DISABLE";
    parameter EXTERNAL_FB = "DISABLE", //"CLKOUT0"; "CLKOUT1"; "CLKOUT2"; "CLKOUT3"; "DISABLE";
    parameter BANDWIDTH   = "OPTIMIZED", //"LOW"; "OPTIMIZED"; "HIGH"
    parameter STDBY_EN     = "FALSE", //"TRUE"; "FALSE"
    parameter RST_INNER_EN = "TRUE",  //"TRUE"; "FALSE"
    parameter RSTODIV_EN   = "TRUE",  //"TRUE"; "FALSE"
    parameter RSTODIV2_EN  = "FALSE", //"TRUE"; "FALSE"
    parameter RSTODIV3_EN  = "FALSE"  //"TRUE"; "FALSE"
    )(
    output CLKOUT,
    output CLKOUT0,
    output CLKOUT1,
    output CLKOUT2,
    output CLKOUT3,
    output PHASE_SOURCE,
    output LOCK,
    input CLKIN1,
    input CLKIN2,
    input CLKFB,
    input CLKIN_SEL,
    input PFDEN,
    input [1:0] PHASE_SEL,
    input PHASE_DIR,
    input PHASE_STEP_N,
    input LOAD_PHASE,
    input CPHASE_STEP_N,
    input CLKOUT0_SYN,
    input CLKOUT1_SYN,
    input CLKOUT2_SYN,
    input CLKOUT3_SYN,
    input STDBY,
    input PLL_PWD,
    input RST,
    input RSTODIV,
    input RSTODIV2,
    input RSTODIV3,
    input APB_CLK,
    input APB_RST_N,
    input [4:0] APB_ADDR,
    input APB_SEL,
    input APB_EN,
    input APB_WRITE,
    input [7:0] APB_WDATA
    );

    initial
    begin
        if((PFDEN_EN == "TRUE") || (PFDEN_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E2 error: illegal setting for PFDEN_EN");

        if((PFDEN_APB_EN == "TRUE") || (PFDEN_APB_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E2 error: illegal setting for PFDEN_APB_EN");

        if((FRACN_EN == "TRUE") || (FRACN_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E2 error: illegal setting for FRACN_EN");

        if((PHASE_APB_EN == "TRUE") || (PHASE_APB_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E2 error: illegal setting for PHASE_APB_EN");

        if((VCOCLK_BYPASS0 == "TRUE") || (VCOCLK_BYPASS0 == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E2 error: illegal setting for VCOCLK_BYPASS0");

        if((VCOCLK_BYPASS1 == "TRUE") || (VCOCLK_BYPASS1 == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E2 error: illegal setting for VCOCLK_BYPASS1");

        if((VCOCLK_BYPASS2 == "TRUE") || (VCOCLK_BYPASS2 == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E2 error: illegal setting for VCOCLK_BYPASS2");

        if((VCOCLK_BYPASS3 == "TRUE") || (VCOCLK_BYPASS3 == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E2 error: illegal setting for VCOCLK_BYPASS3");

        if((CLKOUT0_SYN_EN == "TRUE") || (CLKOUT0_SYN_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E2 error: illegal setting for CLKOUT0_SYN_EN");

        if((CLKOUT1_SYN_EN == "TRUE") || (CLKOUT1_SYN_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E2 error: illegal setting for CLKOUT1_SYN_EN");

        if((CLKOUT2_SYN_EN == "TRUE") || (CLKOUT2_SYN_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E2 error: illegal setting for CLKOUT2_SYN_EN");

        if((CLKOUT3_SYN_EN == "TRUE") || (CLKOUT3_SYN_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E2 error: illegal setting for CLKOUT3_SYN_EN");

        if((INTERNAL_FB == "CLKOUT0") || (INTERNAL_FB == "CLKOUT1") || (INTERNAL_FB == "CLKOUT2") || (INTERNAL_FB == "CLKOUT3") || (INTERNAL_FB == "DISABLE"))
        begin
        end
        else
            $display ("GTP_PLL_E2 error: illegal setting for INTERNAL_FB");

        if((EXTERNAL_FB == "CLKOUT0") || (EXTERNAL_FB == "CLKOUT1") || (EXTERNAL_FB == "CLKOUT2") || (EXTERNAL_FB == "CLKOUT3") || (EXTERNAL_FB == "DISABLE"))
        begin
        end
        else
            $display ("GTP_PLL_E2 error: illegal setting for EXTERNAL_FB");

        if((STDBY_EN == "TRUE") || (STDBY_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E2 error: illegal setting for STDBY_EN");

        if((RST_INNER_EN == "TRUE") || (RST_INNER_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E2 error: illegal setting for RST_INNER_EN");

        if((RSTODIV_EN == "TRUE") || (RSTODIV_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E2 error: illegal setting for RSTODIV_EN");

        if((RSTODIV2_EN == "TRUE") || (RSTODIV2_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E2 error: illegal setting for RSTODIV2_EN");

        if((RSTODIV3_EN == "TRUE") || (RSTODIV3_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E2 error: illegal setting for RSTODIV3_EN");
    end
///////////////////////////////////////////////////////
////INITIAL////////////////////////////////////////////
    reg [15:0] fracn_div;
    reg [7:0]  idivider, fdivider, ratio0, ratio1, ratio2, ratio3;
    reg [7:0]  odiv0_cphase, odiv1_cphase, odiv2_cphase, odiv3_cphase;
    reg [2:0]  odiv0_fphase, odiv1_fphase, odiv2_fphase, odiv3_fphase;
    reg        clkout0_gate_en, clkout1_gate_en, clkout2_gate_en, clkout3_gate_en;
    reg [1:0]  odiv0_clkin_sel, odiv1_clkin_sel, odiv2_clkin_sel, odiv3_clkin_sel;
    reg        vcoclk_bypass0, vcoclk_bypass1, vcoclk_bypass2, vcoclk_bypass3;
    reg [2:0]  clkout0_sel, clkout1_sel, clkout2_sel, clkout3_sel;
    reg        stdby_en, pwd_en, rstodiv_en, rst_en, rstodiv2_en, rstodiv3_en;
    reg        rstodiv_apb, pwd_apb;
    reg [1:0]  phasesel_apb;
    reg        fphasedir_apb, fphasestep_n_apb, load_fphase_apb, cphasestep_n_apb;
    reg        phase_apb_en, pfden_apb_en, pfden_en, pfden_apb;
    reg        lock_mode;
    reg [2:0]  lock_accuracy;
    reg        fracn_en;
    reg        icp_base_trim;

    initial
    begin
        fracn_div    = FRACN_DIV    ;
        idivider     = STATIC_RATIOI;
        fdivider     = STATIC_RATIOF;
        ratio0       = STATIC_RATIO0;
        ratio1       = STATIC_RATIO1;
        ratio2       = STATIC_RATIO2;
        ratio3       = STATIC_RATIO3;
        odiv0_cphase = STATIC_CPHASE0;
        odiv1_cphase = STATIC_CPHASE1;
        odiv2_cphase = STATIC_CPHASE2;
        odiv3_cphase = STATIC_CPHASE3;
        odiv0_fphase = STATIC_PHASE0;
        odiv1_fphase = STATIC_PHASE1;
        odiv2_fphase = STATIC_PHASE2;
        odiv3_fphase = STATIC_PHASE3;

        if(CLKOUT0_SYN_EN == "TRUE")
            clkout0_gate_en = 1'b1;
        else
            clkout0_gate_en = 1'b0;

        if(CLKOUT1_SYN_EN == "TRUE")
            clkout1_gate_en = 1'b1;
        else
            clkout1_gate_en = 1'b0;

        if(CLKOUT2_SYN_EN == "TRUE")
            clkout2_gate_en = 1'b1;
        else
            clkout2_gate_en = 1'b0;

        if(CLKOUT3_SYN_EN == "TRUE")
            clkout3_gate_en = 1'b1;
        else
            clkout3_gate_en = 1'b0;

        odiv0_clkin_sel = ODIV0_CLKIN_SEL;
        odiv1_clkin_sel = ODIV1_CLKIN_SEL;
        odiv2_clkin_sel = ODIV2_CLKIN_SEL;
        odiv3_clkin_sel = ODIV3_CLKIN_SEL;

        if(VCOCLK_BYPASS0 == "TRUE")
            vcoclk_bypass0 = 1'b1;
        else
            vcoclk_bypass0 = 1'b0;

        if(VCOCLK_BYPASS1 == "TRUE")
            vcoclk_bypass1 = 1'b1;
        else
            vcoclk_bypass1 = 1'b0;

        if(VCOCLK_BYPASS2 == "TRUE")
            vcoclk_bypass2 = 1'b1;
        else
            vcoclk_bypass2 = 1'b0;

        if(VCOCLK_BYPASS3 == "TRUE")
            vcoclk_bypass3 = 1'b1;
        else
            vcoclk_bypass3 = 1'b0;

        clkout0_sel = CLKOUT0_SEL;
        clkout1_sel = CLKOUT1_SEL;
        clkout2_sel = CLKOUT2_SEL;
        clkout3_sel = CLKOUT3_SEL;

        if(STDBY_EN == "TRUE")
            stdby_en = 1'b1;
        else
            stdby_en = 1'b0;

        pwd_en = 1'b1;

        if(RSTODIV_EN== "TRUE")
            rstodiv_en = 1'b1;
        else
            rstodiv_en = 1'b0;

        if(RST_INNER_EN == "TRUE")
            rst_en = 1'b1;
        else
            rst_en = 1'b0;

        if(RSTODIV2_EN == "TRUE")
            rstodiv2_en = 1'b1;
        else
            rstodiv2_en = 1'b0;

        if(RSTODIV3_EN == "TRUE")
            rstodiv3_en = 1'b1;
        else
            rstodiv3_en = 1'b0;

        rstodiv_apb      = 1'b0;
        pwd_apb          = 1'b0;
        phasesel_apb     = 2'b11;
        fphasedir_apb    = 1'b1;
        fphasestep_n_apb = 1'b1;
        load_fphase_apb  = 1'b1;
        cphasestep_n_apb = 1'b1;

        if(PHASE_APB_EN == "TRUE")
            phase_apb_en = 1'b1;
        else
            phase_apb_en = 1'b0;

        if(PFDEN_APB_EN == "TRUE")
            pfden_apb_en = 1'b1;
        else     
            pfden_apb_en = 1'b0;

        if(PFDEN_EN == "TRUE")
            pfden_en = 1'b1;
        else
            pfden_en = 1'b0;

        pfden_apb     = 1'b1;
        lock_mode     = LOCK_MODE;
        lock_accuracy = 3'b000;

        if(FRACN_EN == "TRUE")
            fracn_en = 1'b1;
        else     
            fracn_en = 1'b0;

        icp_base_trim = 1'b0;
    end
///////////////////////////////////////////////////////
    wire pll_stdby, pll_pwd;
    wire pll_rst, pll_rstodiv, pll_rstodiv2, pll_rstodiv3;
    wire rst_n, rstodiv2_n, rstodiv3_n;
///////////////////////////////////////////////////////
    wire clk_in;
///////////////////////////////////////////////////////
    reg clk_in_first_time, clk_fb_first_time;
    realtime clk_in_first_edge, clk_fb_first_edge;
    reg adjust;
    realtime fb_route_delay, virtual_delay1;
    integer tmp_ratio;
    realtime tmp_delay, real_delay;
///////////////////////////////////////////////////////
    wire pfden, pfden1;
    reg clk_pfd, vcolow;
    integer cnt;

    reg clk_test, clkwo;
    realtime clk_test_time1 , clk_test_time2, clk_test_time3;
///////////////////////////////////////////////////////
    wire [7:0] divider0, divider1, divider2, divider3;
    real dividerf, frac_div, fsdiv_set_int, fbdiv_set_int;

    wire rstanalog_n;
    realtime clkin_rtime_last, clkin_rtime_next;
    realtime clkin_time, clkin_time1, clkin_time2, clkin_time3;
    reg clkout_lock;
    realtime vcoclk_period, vcoclk_period_half, clkout0_time, clkout1_time, clkout2_time, clkout3_time;
    integer  vcoclk_period_amp;
    realtime vcoclk_period_real, vcoclk_period_dev;

    real cnt_fdiv;
    reg clk_gate, inner_clk;
    reg vcoclk;
    wire pha, phb, phc, phd;
///////////////////////////////////////////////////////
    wire clk_lock;
    reg [2:0] cnt_clkfb;
    reg start_clk;
    reg [9:0] cnt_lock;
    reg lock_wait, lock_reg;
///////////////////////////////////////////////////////
    reg muxa0_out, muxa1_out, muxa2_out, muxa3_out;
    reg muxb0_out, muxb1_out, muxb2_out, muxb3_out;
///////////////////////////////////////////////////////
    reg [2:0] enclk_b0, enclk_b1, enclk_b2, enclk_b3;
    wire b0out, b1out, b2out, b3out;
    reg [7:0] odiv0_cnt, odiv1_cnt, odiv2_cnt, odiv3_cnt;
    reg clkdivr_odiv0, clkdivr_odiv1, clkdivr_odiv2, clkdivr_odiv3;
    reg clkdivf_odiv0, clkdivf_odiv1, clkdivf_odiv2, clkdivf_odiv3;
    wire odiv0_out, odiv1_out, odiv2_out, odiv3_out;
///////////////////////////////////////////////////////
    reg [1:0] phase_sel;
    reg fphase_dir, fphase_step, load_fphase, cphase_step;

    reg last_fphase_step, fphase_overband;
    integer step_odiv0, step_odiv1, step_odiv2, step_odiv3;
    integer step_odiv0_1, step_odiv1_1, step_odiv2_1, step_odiv3_1;
    integer step_odiv0_2, step_odiv1_2, step_odiv2_2, step_odiv3_2;
    integer step_odiv0_3, step_odiv1_3, step_odiv2_3, step_odiv3_3;
    integer step_odiv0_4, step_odiv1_4, step_odiv2_4, step_odiv3_4;
    integer step_odiv0_5, step_odiv1_5, step_odiv2_5, step_odiv3_5;

    reg cphase_step_odiv0, cphase_step_odiv0_1, cphase_step_odiv0_2;
    reg cphase_step_odiv1, cphase_step_odiv1_1, cphase_step_odiv1_2;
    reg cphase_step_odiv2, cphase_step_odiv2_1, cphase_step_odiv2_2;
    reg cphase_step_odiv3, cphase_step_odiv3_1, cphase_step_odiv3_2;

    integer cnt_odiv0, cnt_odiv1, cnt_odiv2, cnt_odiv3;
    integer cnt_odiv0_1, cnt_odiv1_1, cnt_odiv2_1, cnt_odiv3_1;
    integer cnt_odiv0_2, cnt_odiv1_2, cnt_odiv2_2, cnt_odiv3_2;

    realtime vco_fphase_delay0, vco_fphase_delay1, vco_fphase_delay2, vco_fphase_delay3;
    realtime cphase_delay0, cphase_delay1, cphase_delay2, cphase_delay3;
    realtime cphase_delay0_1, cphase_delay1_1, cphase_delay2_1, cphase_delay3_1;
    reg odiv0_out_delay1, odiv1_out_delay1, odiv2_out_delay1, odiv3_out_delay1;
    reg odiv0_out_delay, odiv1_out_delay, odiv2_out_delay, odiv3_out_delay;
///////////////////////////////////////////////////////
    reg clkout0_reg, clkout1_reg, clkout2_reg, clkout3_reg;
///////////////////////////////////////////////////////
    wire clkout0_gate, clkout1_gate, clkout2_gate, clkout3_gate;
    reg [2:0] clkout0_gate_d, clkout1_gate_d, clkout2_gate_d, clkout3_gate_d;
    reg inner_rstn;
///////////////////////////////////////////////////////
    reg rstn_apb, rstn_apb_syn;
///////////////////////////////////////////////////////
    initial
    begin
        clk_in_first_time = 1'b0;
        clk_fb_first_time = 1'b0;
        clk_in_first_edge = 0.0;
        clk_fb_first_edge = 0.0;
        fb_route_delay = 0.0;
        tmp_ratio  = 0;
        tmp_delay  = 0.0;
        real_delay = 0.0;
        clk_pfd  = 1'b0;
        clk_test = 1'b0;
        vcolow   = 1'b0;
        cnt      = 0;
        fsdiv_set_int = 0.0;
        fbdiv_set_int = 0.0;
        clkin_rtime_last = 0.0;
        clkin_rtime_next = 0.0;
        clkin_time  = 0.0;
        clkin_time1 = 0.0;
        clkin_time2 = 0.0;
        clkin_time3 = 0.0;
        clkout_lock = 1'b0;
        vcoclk_period = 0.0;
        vcoclk_period_half = 0.0;
        clkout0_time = 0.0;
        clkout1_time = 0.0;
        clkout2_time = 0.0;
        clkout3_time = 0.0;
        vcoclk_period_amp  = 0;
        vcoclk_period_real = 0.0;
        vcoclk_period_dev  = 0.0;
        cnt_fdiv = 0;
        clk_gate = 1'b0;
        inner_clk = 1'b0;
        vcoclk    = 1'b0;
        cnt_clkfb = 3'b000;
        start_clk = 1'b0;
        cnt_lock  = 10'b00_0000_0000;
        lock_wait = 1'b0;
        lock_reg  = 1'b0;
        muxa0_out = 1'b0;
        muxa1_out = 1'b0;
        muxa2_out = 1'b0;
        muxa3_out = 1'b0;
        muxb0_out = 1'b0;
        muxb1_out = 1'b0;
        muxb2_out = 1'b0;
        muxb3_out = 1'b0;
        enclk_b0  = 3'b000;
        enclk_b1  = 3'b000;
        enclk_b2  = 3'b000;
        enclk_b3  = 3'b000;
        odiv0_cnt = 8'b0000_0000;
        odiv1_cnt = 8'b0000_0000;
        odiv2_cnt = 8'b0000_0000;
        odiv3_cnt = 8'b0000_0000;
        clkdivr_odiv0 = 1'b0;
        clkdivr_odiv1 = 1'b0;
        clkdivr_odiv2 = 1'b0;
        clkdivr_odiv3 = 1'b0;
        clkdivf_odiv0 = 1'b0;
        clkdivf_odiv1 = 1'b0;
        clkdivf_odiv2 = 1'b0;
        clkdivf_odiv3 = 1'b0;
        phase_sel   = 2'b00;
        fphase_dir  = 1'b0;
        fphase_step = 1'b0;
        load_fphase = 1'b0;
        cphase_step = 1'b0;
        last_fphase_step = 1'b0;
        fphase_overband  = 1'b0;
        step_odiv0 = 0;
        step_odiv1 = 0;
        step_odiv2 = 0;
        step_odiv3 = 0;
        step_odiv0_1 = odiv0_fphase;
        step_odiv1_1 = odiv1_fphase;
        step_odiv2_1 = odiv2_fphase;
        step_odiv3_1 = odiv3_fphase;
        step_odiv0_2 = odiv0_fphase;
        step_odiv1_2 = odiv1_fphase;
        step_odiv2_2 = odiv2_fphase;
        step_odiv3_2 = odiv3_fphase;
        step_odiv0_3 = odiv0_fphase;
        step_odiv1_3 = odiv1_fphase;
        step_odiv2_3 = odiv2_fphase;
        step_odiv3_3 = odiv3_fphase;
        step_odiv0_4 = odiv0_fphase;
        step_odiv1_4 = odiv1_fphase;
        step_odiv2_4 = odiv2_fphase;
        step_odiv3_4 = odiv3_fphase;
        cphase_step_odiv0   = 1'b1;
        cphase_step_odiv0_1 = 1'b1;
        cphase_step_odiv0_2 = 1'b1;
        cphase_step_odiv1   = 1'b1;
        cphase_step_odiv1_1 = 1'b1;
        cphase_step_odiv1_2 = 1'b1;
        cphase_step_odiv2   = 1'b1;
        cphase_step_odiv2_1 = 1'b1;
        cphase_step_odiv2_2 = 1'b1;
        cphase_step_odiv3   = 1'b1;
        cphase_step_odiv3_1 = 1'b1;
        cphase_step_odiv3_2 = 1'b1;
        cnt_odiv0 = 1;
        cnt_odiv1 = 1;
        cnt_odiv2 = 1;
        cnt_odiv3 = 1;
        cnt_odiv0_1 = 1;
        cnt_odiv1_1 = 1;
        cnt_odiv2_1 = 1;
        cnt_odiv3_1 = 1;
        cnt_odiv0_2 = 1;
        cnt_odiv1_2 = 1;
        cnt_odiv2_2 = 1;
        cnt_odiv3_2 = 1;
        vco_fphase_delay0 = 0.0;
        vco_fphase_delay1 = 0.0;
        vco_fphase_delay2 = 0.0;
        vco_fphase_delay3 = 0.0;
        cphase_delay0 = 0.0;
        cphase_delay1 = 0.0;
        cphase_delay2 = 0.0;
        cphase_delay3 = 0.0;
        cphase_delay0_1 = 0.0;
        cphase_delay1_1 = 0.0;
        cphase_delay2_1 = 0.0;
        cphase_delay3_1 = 0.0;
        odiv0_out_delay1 = 1'b0;
        odiv1_out_delay1 = 1'b0;
        odiv2_out_delay1 = 1'b0;
        odiv3_out_delay = 1'b0;
        odiv0_out_delay = 1'b0;
        odiv1_out_delay = 1'b0;
        odiv2_out_delay = 1'b0;
        odiv3_out_delay = 1'b0;
        clkout0_reg = 1'b0;
        clkout1_reg = 1'b0;
        clkout2_reg = 1'b0;
        clkout3_reg = 1'b0;
        clkout0_gate_d = 1'b0;
        clkout1_gate_d = 1'b0;
        clkout2_gate_d = 1'b0;
        clkout3_gate_d = 1'b0;
        rstn_apb     = 1'b0;
        rstn_apb_syn = 1'b0;
        inner_rstn = 1'b0;
        #1;
        inner_rstn = 1'b1;
        clk_in_first_time = 1'b1;
        clk_fb_first_time = 1'b1;
    end
///////////////////////////////////////////////////////
////RESET//////////////////////////////////////////////
    assign pll_stdby = (stdby_en == 1'b1) ? STDBY   : 1'b0;
    assign pll_pwd   = (pwd_en   == 1'b1) ? PLL_PWD : 1'b0;

    assign pll_rst      = (rst_en      == 1'b1) ? RST      : 1'b0;
    assign pll_rstodiv  = (rstodiv_en  == 1'b1) ? RSTODIV  : 1'b0;
    assign pll_rstodiv2 = (rstodiv2_en == 1'b1) ? RSTODIV2 : 1'b0;
    assign pll_rstodiv3 = (rstodiv3_en == 1'b1) ? RSTODIV3 : 1'b0;

    assign rst_n = ~pll_stdby & (~pll_pwd & ~pwd_apb) & ~pll_rst & (~pll_rstodiv & ~rstodiv_apb) & inner_rstn;
    assign rstodiv2_n = rst_n & ~pll_rstodiv2;
    assign rstodiv3_n = rst_n & ~pll_rstodiv3;
///////////////////////////////////////////////////////
////INPUT_CLK_SEL//////////////////////////////////////
    assign clk_in = (CLKIN_SEL == 1'b0) ? CLKIN1 : CLKIN2;
///////////////////////////////////////////////////////
////FBCK_DELAY/////////////////////////////////////////
    always @(posedge clk_in or negedge rst_n)
    begin
        if(!rst_n)
        begin
            clk_in_first_time = 1'b1;
            clk_in_first_edge = 0.0;
        end
        else
        begin
            if(clk_in_first_time == 1'b1)
                clk_in_first_edge = $realtime;
            clk_in_first_time = 1'b0;
        end
    end

    always @(posedge CLKFB or negedge rst_n)
    begin
        if(!rst_n)
        begin
            clk_fb_first_time = 1'b1;
            clk_fb_first_edge = 0.0;
        end
        else
        begin
           if(clk_fb_first_time == 1'b1)
                clk_fb_first_edge = $realtime;
            clk_fb_first_time = 1'b0;
        end
    end
////////////////////////////////////////////////////////////////////////////////////
////PFD_ENABLE//////////////////////////////////////////////////////////////////////
    assign pfden  = (pfden_en     == 1'b1) ? PFDEN     : 1'b1 ;
    assign pfden1 = (pfden_apb_en == 1'b1) ? pfden_apb : pfden;

    always #0.5 clk_pfd = ~clk_pfd;

    always @(posedge clk_pfd or negedge rst_n)
    begin
        if(!rst_n)
        begin
            vcolow <= 0;
            cnt = 0;
        end
        else
            if(pfden1)
            begin
                vcolow <= 0;
                cnt = 0;
            end
            else
            begin
                cnt = cnt + 1;
                if(cnt == 500000)
                vcolow <= 1;
            end
    end

    always #200 clk_test = ~clk_test;

    always @(posedge clk_test or negedge rst_n)
    begin
        if(!rst_n)
        begin
            clkwo <= 1'b0;
            clk_test_time1 = 0;
            clk_test_time2 = 0;
            clk_test_time3 = 0;

        end
        else
        begin
            clk_test_time3 = clk_test_time2;
            clk_test_time2 = clk_test_time1;
            clk_test_time1 = clkin_rtime_next;
            if(clk_test_time3 == clk_test_time1)
                clkwo <= 1'b1;
            else
                clkwo <= 1'b0;
        end
    end
///////////////////////////////////////////////////////
////PLL_ANALOG/////////////////////////////////////////
////FEEDBACK_DIVIDER_CAL///////////////////////////////
    assign divider0 = ratio0;
    assign divider1 = ratio1;
    assign divider2 = ratio2;
    assign divider3 = ratio3;

    always @(*)
    begin
        dividerf = fdivider;
        frac_div = fracn_div;

        if(INTERNAL_FB == "CLKOUT0" || EXTERNAL_FB == "CLKOUT0")
            fsdiv_set_int = divider0;
        else if(INTERNAL_FB == "CLKOUT1" || EXTERNAL_FB == "CLKOUT1")
            fsdiv_set_int = divider1;
        else if(INTERNAL_FB == "CLKOUT2" || EXTERNAL_FB == "CLKOUT2")
            fsdiv_set_int = divider2;
        else if(INTERNAL_FB == "CLKOUT3" || EXTERNAL_FB == "CLKOUT3")
            fsdiv_set_int = divider3;
    end

    always @(*)
    begin
        if(fracn_en == 1'b1)
            fbdiv_set_int = fsdiv_set_int * (dividerf + (frac_div / 65536));
        else
            fbdiv_set_int = dividerf * fsdiv_set_int;
    end
////PLL_VCO_CAL////////////////////////////////////////
    assign rstanalog_n = rst_n & ~vcolow;

    always @(posedge clk_in or negedge rstanalog_n)
    begin
        if(!rstanalog_n)
        begin
            clkin_rtime_last = 0.0;
            clkin_rtime_next = 0.0;
            clkin_time  <= 0.0;
            clkin_time1 <= 0.0;
            clkin_time2 <= 0.0;
            clkin_time3 <= 0.0;
            clkout_lock <= 0.0;
            vcoclk_period <= 1'b0;
            vcoclk_period_half <= 0.0;
            vcoclk_period_amp  <= 0.0;
            vcoclk_period_real <= 0.0;
            vcoclk_period_dev  <= 0.0;
        end
        else
        begin
            clkin_rtime_last = clkin_rtime_next;
            clkin_rtime_next = $realtime;
            if(clkin_rtime_last > 0)
            begin
                clkin_time  <= clkin_rtime_next-clkin_rtime_last;
                clkin_time1 <= clkin_time;
                clkin_time2 <= clkin_time1;
                clkin_time3 <= clkin_time2;
            end
            if(clkin_time > 0)
            begin
                clkout_lock <= (clkin_time  > 0) &&
                               (clkin_time1 > 0) &&
                               (clkin_time2 > 0) &&
                               (clkin_time3 > 0) &&
                               ((clkin_time - clkin_time1)  < 0.0001) &&
                               ((clkin_time1 - clkin_time)  < 0.0001) &&
                               ((clkin_time1 - clkin_time2) < 0.0001) &&
                               ((clkin_time2 - clkin_time1) < 0.0001) &&
                               ((clkin_time2 - clkin_time3) < 0.0001) &&
                               ((clkin_time3 - clkin_time2) < 0.0001);
            end
            if(clkin_time > 0)
            begin
                vcoclk_period      = (clkin_time * idivider) / fbdiv_set_int;
                vcoclk_period_half = vcoclk_period / 2;
                clkout0_time       = vcoclk_period * divider0;
                clkout1_time       = vcoclk_period * divider1;
                clkout2_time       = vcoclk_period * divider2;
                clkout3_time       = vcoclk_period * divider3;
                vcoclk_period_amp  = vcoclk_period_half * 100000;
                vcoclk_period_real = vcoclk_period_amp / 100000.0;
                vcoclk_period_dev  = (clkin_time - (vcoclk_period_real * 2 * fbdiv_set_int) / idivider) / 2;
            end
        end
    end

    always @(clkout_lock or inner_clk or clkwo)
    begin
        if(clkout_lock == 1'b0 || clkwo == 1'b1)
        begin
            inner_clk <= 1'b0;
            clk_gate  <= 1'b1;
            cnt_fdiv   = 0;
        end
        else
            if(clk_gate == 1)
            begin
                inner_clk <= 1'b1;
                clk_gate  <= 1'b0;
                cnt_fdiv   = 0;
            end
            else
            begin
                cnt_fdiv = cnt_fdiv + 1;
                if(cnt_fdiv  == fbdiv_set_int)
                begin
                    inner_clk <= #(vcoclk_period_half + vcoclk_period_dev) ~inner_clk;
                    cnt_fdiv = 0;
                end
                else
                    inner_clk <= #vcoclk_period_half ~inner_clk;
            end
    end

    always @(clk_in or CLKFB or negedge rst_n)
    begin
        if(!rst_n)
        begin
            adjust <= 1'b1;
            fb_route_delay = 0.0;
            tmp_ratio  = 0;
            tmp_delay  = 0.0;
            real_delay = 0.0;
        end
        else
            if(adjust == 1'b1)
            begin
                fb_route_delay = clk_fb_first_edge - clk_in_first_edge;
                if((clkin_time > 0) && (fb_route_delay > 0))
                begin
                    tmp_ratio  = fb_route_delay / clkin_time;
                    tmp_delay  = fb_route_delay - (clkin_time * tmp_ratio);
                    real_delay = clkin_time - tmp_delay;
                    adjust <= 1'b0;
                end
            end
    end

    always @(inner_clk)
    begin
        if(INTERNAL_FB == "DISABLE")
            vcoclk <= #real_delay inner_clk;
        else
            vcoclk <= inner_clk;
    end

    assign pha = vcoclk;
    assign phb = vcoclk;
    assign phc = vcoclk;
    assign phd = vcoclk;
///////////////////////////////////////////////////////
////PLL_LOCK///////////////////////////////////////////
    assign clk_lock = (INTERNAL_FB == "DISABLE") ? CLKFB : clk_in;

    always @(posedge clk_lock or negedge rstanalog_n)
    begin
        if(!rstanalog_n)
        begin
            start_clk <= 1'b0;
            cnt_clkfb <= 2'b00;
        end
        else
            if(cnt_clkfb == 3)
                start_clk = 1'b1;
            else
                cnt_clkfb = cnt_clkfb + 1;
    end

    always @(posedge clk_in or negedge rstanalog_n or clk_gate)
    begin
        if(!rstanalog_n)
        begin
            cnt_lock  <= 8'h1;
            lock_wait <= 1'b0;
        end
        else
            if(!clk_gate && start_clk)
                if(cnt_lock == idivider * 3)
                    lock_wait <= 1'b1;
                else
                    cnt_lock <= cnt_lock + 1'b1;
            else
            begin
                cnt_lock <= 8'h1;
                lock_wait <= 1'b0;
            end
    end

    always @(posedge clk_in or negedge rstanalog_n or clk_gate)
    begin
        if(!rst_n)
            lock_reg <= 1'b0;
        else
            if(LOCK_MODE == 1'b0)
                if(!clk_gate)
                    lock_reg <= lock_wait;
                else
                    lock_reg <= 1'b0;
            else
                lock_reg <= lock_reg | lock_wait;
    end

    assign LOCK = lock_reg;
///////////////////////////////////////////////////////
////ODIV_CAS///////////////////////////////////////////
    always @(*)
    begin
        if(vcoclk_bypass0 == 1'b0)
            muxa0_out <= pha;
        else if(vcoclk_bypass0 == 1'b1)
            muxa0_out <= clk_in;
    end

    always @(*)
    begin
        if(vcoclk_bypass1 == 1'b0)
            muxa1_out <= phb;
        else if(vcoclk_bypass1 == 1'b1)
            muxa1_out <= clk_in;
    end

    always @(*)
    begin
        if(vcoclk_bypass2 == 1'b0)
            muxa2_out <= phc;
        else if(vcoclk_bypass2 == 1'b1)
            muxa2_out <= clk_in;
    end

    always @(*)
    begin
        if(vcoclk_bypass3 == 1'b0)
            muxa3_out <= phd;
        else if(vcoclk_bypass3 == 1'b1)
            muxa3_out <= clk_in;
    end

    always @(*)
    begin
        if(odiv0_clkin_sel == 2'b00)
            muxb0_out <= muxa0_out;
        else if(odiv0_clkin_sel == 2'b01)
            muxb0_out <= odiv3_out_delay;
        else if(odiv0_clkin_sel == 2'b10)
            muxb0_out <= odiv1_out_delay;
        else if(odiv0_clkin_sel == 2'b11)
            muxb0_out <= odiv2_out_delay;
    end

    always @(*)
    begin
        if(odiv1_clkin_sel == 2'b00)
            muxb1_out <= muxa1_out;
        else if(odiv1_clkin_sel == 2'b01)
            muxb1_out <= odiv0_out_delay;
        else if(odiv1_clkin_sel == 2'b10)
            muxb1_out <= odiv3_out_delay;
        else if(odiv1_clkin_sel == 2'b11)
            muxb1_out <= odiv2_out_delay;
    end

    always @(*)
    begin
        if(odiv2_clkin_sel == 2'b00)
            muxb2_out <= muxa2_out;
        else if(odiv2_clkin_sel == 2'b01)
            muxb2_out <= odiv0_out_delay;
        else if(odiv2_clkin_sel == 2'b10)
            muxb2_out <= odiv1_out_delay;
        else if(odiv2_clkin_sel == 2'b11)
            muxb2_out <= odiv3_out_delay;
    end

    always @(*)
    begin
        if(odiv3_clkin_sel == 2'b00)
            muxb3_out <= muxa3_out;
        else if(odiv3_clkin_sel == 2'b01)
            muxb3_out <= odiv0_out_delay;
        else if(odiv3_clkin_sel == 2'b10)
            muxb3_out <= odiv1_out_delay;
        else if(odiv3_clkin_sel == 2'b11)
            muxb3_out <= odiv2_out_delay;
    end
///////////////////////////////////////////////////////
////PLL_ODIV///////////////////////////////////////////
////ODIV0//////////////////////////////////////////////
    always @(negedge muxb0_out or negedge rst_n)
    begin
        if(!rst_n)
            enclk_b0 <= 3'b000;
        else
            enclk_b0 <= {enclk_b0[1:0],1'b1};
    end

    assign b0out = muxb0_out & enclk_b0[2];

    always @(posedge b0out or negedge rst_n)
    begin
        if(!rst_n)
            odiv0_cnt <= 8'b0000_0000;
        else
            if(odiv0_cnt == divider0 - 1'b1)
                odiv0_cnt <= 10'b00_0000_0000;
            else
                odiv0_cnt <= odiv0_cnt + 1'b1;
    end

    always @(posedge b0out or negedge rst_n)
    begin
        if(!rst_n)
            clkdivr_odiv0 <= 1'b0;
        else
            if(odiv0_cnt < {1'b0,divider0[7:1]})
                clkdivr_odiv0 <= 1'b1;
            else
                clkdivr_odiv0 <= 1'b0;
    end

    always @(negedge b0out or negedge rst_n)
    begin
        if(!rst_n)
            clkdivf_odiv0 <= 1'b0;
        else
            if(divider0[0] == 1'b0)
                clkdivf_odiv0 <= 1'b0;
            else
                clkdivf_odiv0 <= clkdivr_odiv0;
    end

    assign odiv0_out = (divider0 == 7'd1) ? b0out : (clkdivr_odiv0 | clkdivf_odiv0);
////ODIV1//////////////////////////////////////////////
    always @(negedge muxb1_out or negedge rst_n)
    begin
        if(!rst_n)
            enclk_b1 <= 3'b000;
        else
            enclk_b1 <= {enclk_b1[1:0],1'b1};
    end

    assign b1out = muxb1_out & enclk_b1[2];

    always @(posedge b1out or negedge rst_n)
    begin
        if(!rst_n)
            odiv1_cnt <= 8'b0000_0000;
        else
            if(odiv1_cnt == divider1 - 1'b1)
                odiv1_cnt <= 10'b00_0000_0000;
            else
                odiv1_cnt <= odiv1_cnt + 1'b1;
    end

    always @(posedge b1out or negedge rst_n)
    begin
        if(!rst_n)
            clkdivr_odiv1 <= 1'b0;
        else
            if(odiv1_cnt < {1'b0,divider1[7:1]})
                clkdivr_odiv1 <= 1'b1;
            else
                clkdivr_odiv1 <= 1'b0;
    end

    always @(negedge b1out or negedge rst_n)
    begin
        if(!rst_n)
            clkdivf_odiv1 <= 1'b0;
        else
            if(divider1[0] == 1'b0)
                clkdivf_odiv1 <= 1'b0;
            else
                clkdivf_odiv1 <= clkdivr_odiv1;
    end

    assign odiv1_out = (divider1 == 7'd1) ? b1out : (clkdivr_odiv1 | clkdivf_odiv1);
////ODIV2//////////////////////////////////////////////
    always @(negedge muxb2_out or negedge rstodiv2_n)
    begin
        if(!rstodiv2_n)
            enclk_b2 <= 3'b000;
        else
            enclk_b2 <= {enclk_b2[1:0],1'b1};
    end

    assign b2out = muxb2_out & enclk_b2[2];

    always @(posedge b2out or negedge rstodiv2_n)
    begin
        if(!rstodiv2_n)
            odiv2_cnt <= 8'b0000_0000;
        else
            if(odiv2_cnt == divider2 - 1'b1)
                odiv2_cnt <= 10'b00_0000_0000;
            else
                odiv2_cnt <= odiv2_cnt + 1'b1;
    end

    always @(posedge b2out or negedge rstodiv2_n)
    begin
        if(!rstodiv2_n)
            clkdivr_odiv2 <= 1'b0;
        else
            if(odiv2_cnt < {1'b0,divider2[7:1]})
                clkdivr_odiv2 <= 1'b1;
            else
                clkdivr_odiv2 <= 1'b0;
    end

    always @(negedge b2out or negedge rst_n)
    begin
        if(!rstodiv2_n)
            clkdivf_odiv2 <= 1'b0;
        else
            if(divider2[0] == 1'b0)
                clkdivf_odiv2 <= 1'b0;
            else
                clkdivf_odiv2 <= clkdivr_odiv2;
    end

    assign odiv2_out = (divider2 == 7'd1) ? b2out : (clkdivr_odiv2 | clkdivf_odiv2);
////ODIV3//////////////////////////////////////////////
    always @(negedge muxb3_out or negedge rstodiv3_n)
    begin
        if(!rstodiv3_n)
            enclk_b3 <= 3'b000;
        else
            enclk_b3 <= {enclk_b3[1:0],1'b1};
    end

    assign b3out = muxb3_out & enclk_b3[2];

    always @(posedge b3out or negedge rstodiv3_n)
    begin
        if(!rstodiv3_n)
            odiv3_cnt <= 8'b0000_0000;
        else
            if(odiv3_cnt == divider3 - 1'b1)
                odiv3_cnt <= 10'b00_0000_0000;
            else
                odiv3_cnt <= odiv3_cnt + 1'b1;
    end

    always @(posedge b3out or negedge rstodiv3_n)
    begin
        if(!rstodiv3_n)
            clkdivr_odiv3 <= 1'b0;
        else
            if(odiv3_cnt < {1'b0,divider3[7:1]})
                clkdivr_odiv3 <= 1'b1;
            else
                clkdivr_odiv3 <= 1'b0;
    end

    always @(negedge b3out or negedge rst_n)
    begin
        if(!rstodiv3_n)
            clkdivf_odiv3 <= 1'b0;
        else
            if(divider3[0] == 1'b0)
                clkdivf_odiv3 <= 1'b0;
            else
                clkdivf_odiv3 <= clkdivr_odiv3;
    end

    assign odiv3_out = (divider3 == 7'd1) ? b3out : (clkdivr_odiv3 | clkdivf_odiv3);
///////////////////////////////////////////////////////
////PHASE_SHIFT////////////////////////////////////////
    assign PHASE_SOURCE = phase_apb_en;

    always @(*)
    begin
        if(phase_apb_en == 1'b0)
        begin
            phase_sel   = PHASE_SEL;
            fphase_dir  = PHASE_DIR;
            fphase_step = PHASE_STEP_N;
            load_fphase = LOAD_PHASE;
            cphase_step = CPHASE_STEP_N;
        end
        else
        begin
            phase_sel   = phasesel_apb;
            fphase_dir  = fphasedir_apb;
            fphase_step = fphasestep_n_apb;
            load_fphase = load_fphase_apb;
            cphase_step = cphasestep_n_apb;
        end
    end

    always @(fphase_step)
    begin
        last_fphase_step <= fphase_step;
    end

    always @(*)
    begin
        if(load_fphase == 1'b1)
        begin
            step_odiv0  = step_odiv0_1;
            step_odiv1  = step_odiv1_1;
            step_odiv2 = step_odiv2_1;
            step_odiv3 = step_odiv3_1;
        end
        else
            if(phase_sel == 2'b00)
            begin
                if(fphase_step === 1'b0 && last_fphase_step === 1'b1)
                    if(fphase_dir == 1'b0)
                        step_odiv0 <= step_odiv0 + 1;
                    else
                        step_odiv0 <= step_odiv0 - 1;
            end
            else if(phase_sel == 2'b11)
            begin
                if(fphase_step === 1'b0 && last_fphase_step === 1'b1)
                    if(fphase_dir == 1'b0)
                        step_odiv1 <= step_odiv1 + 1;
                    else
                        step_odiv1 <= step_odiv1 - 1;
            end
            else if(phase_sel == 2'b10)
            begin
                if(fphase_step === 1'b0 && last_fphase_step === 1'b1)
                    if(fphase_dir == 1'b0)
                        step_odiv2 <= step_odiv2 + 1;
                    else
                        step_odiv2 <= step_odiv2 - 1;
            end
            else if(phase_sel == 2'b01)
            begin
                if(fphase_step === 1'b0 && last_fphase_step === 1'b1)
                    if(fphase_dir == 1'b0)
                        step_odiv3 <= step_odiv3 + 1;
                    else
                        step_odiv3 <= step_odiv3 - 1;
            end
    end

    always @(*)
    begin
        if(phase_sel == 2'b00)
        begin
            if((fphase_dir == 1'b0 && step_odiv0 == 7) || (fphase_dir == 1'b1 && step_odiv0 == 0))
                fphase_overband = 1'b1;
            else
                fphase_overband = 1'b0;
        end
        else if(phase_sel == 2'b11)
        begin
            if((fphase_dir == 1'b0 && step_odiv1 == 7) || (fphase_dir == 1'b1 && step_odiv1 == 0))
                fphase_overband = 1'b1;
            else
                fphase_overband = 1'b0;
        end
        else if(phase_sel == 2'b10)
        begin
            if((fphase_dir == 1'b0 && step_odiv2 == 7) || (fphase_dir == 1'b1 && step_odiv2 == 0))
                fphase_overband = 1'b1;
            else
                fphase_overband = 1'b0;
        end
        else if(phase_sel == 2'b01)
        begin
            if((fphase_dir == 1'b0 && step_odiv3 == 7) || (fphase_dir == 1'b1 && step_odiv3 == 0))
                fphase_overband = 1'b1;
            else
                fphase_overband = 1'b0;
        end
    end

    always @(posedge last_fphase_step or negedge rst_n)
    begin
        if(!rst_n)
        begin
            step_odiv0_1 <= odiv0_fphase;
            step_odiv1_1 <= odiv1_fphase;
            step_odiv2_1 <= odiv2_fphase;
            step_odiv3_1 <= odiv3_fphase;
        end
        else
        begin
            step_odiv0_1 <= step_odiv0;
            step_odiv1_1 <= step_odiv1;
            step_odiv2_1 <= step_odiv2;
            step_odiv3_1 <= step_odiv3;
        end
    end

    always @(posedge inner_clk)
    begin
        step_odiv0_2 <= step_odiv0_1;
        step_odiv0_3 <= step_odiv0_2;
        step_odiv1_2 <= step_odiv1_1;
        step_odiv1_3 <= step_odiv1_2;
        step_odiv2_2 <= step_odiv2_1;
        step_odiv2_3 <= step_odiv2_2;
        step_odiv3_2 <= step_odiv3_1;
        step_odiv3_3 <= step_odiv3_2;
    end

    always @(negedge inner_clk)
    begin
        step_odiv0_4 <= step_odiv0_3;
        step_odiv1_4 <= step_odiv1_3;
        step_odiv2_4 <= step_odiv2_3;
        step_odiv3_4 <= step_odiv3_3;
    end

    always @(posedge odiv0_out)
    begin
        cphase_step_odiv0   <= cphase_step;
        cphase_step_odiv0_1 <= cphase_step_odiv0;
    end

    always @(negedge odiv0_out_delay1)
    begin
        cphase_step_odiv0_2 <= cphase_step_odiv0_1;
    end

    always @(posedge odiv1_out)
    begin
        cphase_step_odiv1   <= cphase_step;
        cphase_step_odiv1_1 <= cphase_step_odiv1;
    end

    always @(negedge odiv1_out_delay1)
    begin
        cphase_step_odiv1_2 <= cphase_step_odiv1_1;
    end

    always @(posedge odiv2_out)
    begin

        cphase_step_odiv2   <= cphase_step;
        cphase_step_odiv2_1 <= cphase_step_odiv2;
    end

    always @(negedge odiv2_out_delay1)
    begin
        cphase_step_odiv2_2 <= cphase_step_odiv2_1;
    end

    always @(posedge odiv3_out)
    begin

        cphase_step_odiv3   <= cphase_step;
        cphase_step_odiv3_1 <= cphase_step_odiv3;
    end

    always @(negedge odiv3_out_delay1)
    begin
        cphase_step_odiv3_2 <= cphase_step_odiv3_1;
    end

    always @(negedge cphase_step_odiv0_2)
    begin
        if(phase_sel == 2'b00)
            cnt_odiv0 <= cnt_odiv0 + 1;
    end

    always @(negedge cphase_step_odiv1_2)
    begin
        if(phase_sel == 2'b11)
            cnt_odiv1 <= cnt_odiv1 + 1;
    end

    always @(negedge cphase_step_odiv2_2)
    begin
        if(phase_sel == 2'b10)
            cnt_odiv2 <= cnt_odiv2 + 1;
    end

    always @(negedge cphase_step_odiv3_2)
    begin
        if(phase_sel == 2'b01)
            cnt_odiv3 <= cnt_odiv3 + 1;
    end

    always @(posedge cphase_step_odiv0_2 or negedge rst_n)
    begin
        if(!rst_n)
            cnt_odiv0_1 <= 1;
        else
            cnt_odiv0_1 <= cnt_odiv0;
    end

    always @(posedge cphase_step_odiv1_2 or negedge rst_n)
    begin
        if(!rst_n)
            cnt_odiv1_1 <= 1;
        else
            cnt_odiv1_1 <= cnt_odiv1;
    end

    always @(posedge cphase_step_odiv2_2 or negedge rst_n)
    begin
        if(!rst_n)
            cnt_odiv2_1 <= 1;
        else
            cnt_odiv2_1 <= cnt_odiv2;
    end

    always @(posedge cphase_step_odiv3_2 or negedge rst_n)
    begin
        if(!rst_n)
            cnt_odiv3_1 <= 1;
        else
            cnt_odiv3_1 <= cnt_odiv3;
    end

////PHASE_SHIFT_CAL////////////////////////////////////
    always @(*)
    begin
        if(step_odiv0_4 >= 0)
            step_odiv0_5 <= step_odiv0_4;
        else
            step_odiv0_5 <= step_odiv0_4 + (~step_odiv0_4/(8*divider0))*8*divider0;

        if(step_odiv1_4 >= 0)
            step_odiv1_5 <= step_odiv1_4;
        else
            step_odiv1_5 <= step_odiv1_4 + (~step_odiv1_4/(8*divider1))*8*divider1;

        if(step_odiv2_4 >= 0)
            step_odiv2_5 <= step_odiv2_4;
        else
            step_odiv2_5 <= step_odiv2_4 + (~step_odiv2_4/(8*divider2))*8*divider2;

        if(step_odiv3_4 >= 0)
            step_odiv3_5 <= step_odiv3_4;
        else
            step_odiv3_5 <= step_odiv3_4 + (~step_odiv3_4/(8*divider3))*8*divider3;
    end

    always @(*)
    begin      
        if(clkout0_time > 0)
            if(step_odiv0_5 >= 0)
                vco_fphase_delay0 <= (step_odiv0_5 * clkout0_time) / (8 * divider0);
            else
                vco_fphase_delay0 <= clkout0_time + (step_odiv0_5 * clkout0_time) / (8 * divider0);

        if(clkout1_time > 0)
            if(step_odiv1_5 >= 0)
                vco_fphase_delay1 <= (step_odiv1_5 * clkout1_time) / (8 * divider1);
            else
                vco_fphase_delay1 <= clkout1_time + (step_odiv1_5 * clkout1_time) / (8 * divider1);

        if(clkout2_time > 0)
            if(step_odiv2_5 >= 0)
                vco_fphase_delay2 <= (step_odiv2_5 * clkout2_time) / (8 * divider2);
            else
                vco_fphase_delay2 <= clkout2_time + (step_odiv2_5 * clkout2_time) / (8 * divider2);

        if(clkout3_time > 0)
            if(step_odiv3_5 >= 0)
                vco_fphase_delay3 <= (step_odiv3_5 * clkout3_time) / (8 * divider3);
            else
                vco_fphase_delay3 <= clkout3_time + (step_odiv3_5 * clkout3_time) / (8 * divider3);
    end

    always @(*)
    begin
        if(clkout0_time > 0)
            if(divider0 >= odiv0_cphase)
                cphase_delay0 <= clkout0_time - (((divider0 - odiv0_cphase) * clkout0_time) / divider0);
            else
                cphase_delay0 <= ((odiv0_cphase - divider0) * clkout0_time) / divider0;
        else
            cphase_delay0 <= 0.0;

        if(clkout1_time > 0)
            if(divider1 >= odiv1_cphase)
                cphase_delay1 <= clkout1_time - (((divider1 - odiv1_cphase) * clkout1_time) / divider1);
            else
                cphase_delay1 <= ((odiv1_cphase - divider1) * clkout1_time)/ divider1;
        else
            cphase_delay1 <= 0.0;

        if(clkout2_time > 0)
            if(divider2 >= odiv2_cphase)
                cphase_delay2 <= clkout2_time - (((divider2 - odiv2_cphase) * clkout2_time) / divider2);
            else
                cphase_delay2 <= ((odiv2_cphase - divider2) * clkout2_time) / divider2;
        else
            cphase_delay2 <= 0.0;

        if(clkout3_time > 0)
            if(divider3 >= odiv3_cphase)
                cphase_delay3 <= clkout3_time - (((divider3 - odiv3_cphase) * clkout3_time) / divider3);
            else
                cphase_delay3 <= ((odiv3_cphase - divider3) * clkout3_time) / divider3;
        else
                cphase_delay3 <= 0.0;
    end
////PHASE_SHIFT_DLY////////////////////////////////////
    always @(odiv0_out)
    begin
        odiv0_out_delay1 <= #(vco_fphase_delay0) odiv0_out;
    end

    always @(*)
    begin
        if(divider0 >= cnt_odiv0_1)
            cnt_odiv0_2 <= cnt_odiv0_1;
        else
            cnt_odiv0_2 <= cnt_odiv0_1 - (cnt_odiv0_1/divider0)*divider0;
    end

    always @(*)
    begin
        cphase_delay0_1 <= cnt_odiv0_2 * cphase_delay0;
    end

    always @(odiv0_out_delay1)
    begin
        odiv0_out_delay <= #(cphase_delay0_1) odiv0_out_delay1;
    end

    always @(odiv1_out)
    begin
        odiv1_out_delay1 <= #(vco_fphase_delay1) odiv1_out;
    end

    always @(*)
    begin
        if(divider1 >= cnt_odiv1_1)
            cnt_odiv1_2 <= cnt_odiv1_1;
        else
            cnt_odiv1_2 <= cnt_odiv1_1 - (cnt_odiv1_1/divider1)*divider1;
    end

    always @(*)
    begin
        cphase_delay1_1 <= cnt_odiv1_2 * cphase_delay1;
    end

    always @(odiv1_out_delay1)
    begin
        odiv1_out_delay <= #(cphase_delay1_1) odiv1_out_delay1;
    end

    always @(odiv2_out)
    begin
        odiv2_out_delay1 <= #(vco_fphase_delay2) odiv2_out;
    end

    always @(*)
    begin
        if(divider2 >= cnt_odiv2_1)
            cnt_odiv2_2 <= cnt_odiv2_1;
        else
            cnt_odiv2_2 <= cnt_odiv2_1 - (cnt_odiv2_1/divider2)*divider2;
    end

    always @(*)
    begin
        cphase_delay2_1 <= cnt_odiv2_2 * cphase_delay2;
    end

    always @(odiv2_out_delay1)
    begin
        odiv2_out_delay <= #(cphase_delay2_1) odiv2_out_delay1;
    end

    always @(odiv3_out)
    begin
        odiv3_out_delay1 <= #(vco_fphase_delay3) odiv3_out;
    end

    always @(*)
    begin
        if(divider3 >= cnt_odiv3_1)
            cnt_odiv3_2 <= cnt_odiv3_1;
        else
            cnt_odiv3_2 <= cnt_odiv3_1 - (cnt_odiv3_1/divider3)*divider3;
    end

    always @(*)
    begin
        cphase_delay3_1 <= cnt_odiv3_2 * cphase_delay3;
    end

    always @(odiv3_out_delay1)
    begin
        odiv3_out_delay <= #(cphase_delay3_1) odiv3_out_delay1;
    end
///////////////////////////////////////////////////////
////CLKOUT_SEL/////////////////////////////////////////
    always @(*)
    begin
        case(clkout0_sel)
            3'b000: clkout0_reg = odiv0_out_delay;
            3'b001: clkout0_reg = odiv1_out_delay;
            3'b010: clkout0_reg = odiv2_out_delay;
            3'b011: clkout0_reg = odiv3_out_delay;
            3'b100: clkout0_reg = clk_in;
        endcase
    end

    always @(*)
    begin
        case(clkout1_sel)
            3'b000: clkout1_reg = odiv1_out_delay;
            3'b001: clkout1_reg = odiv2_out_delay;
            3'b010: clkout1_reg = odiv3_out_delay;
            3'b011: clkout1_reg = odiv0_out_delay;
            3'b100: clkout1_reg = clk_in;
        endcase
    end

    always @(*)
    begin
        case(clkout2_sel)
            3'b000: clkout2_reg = odiv2_out_delay;
            3'b001: clkout2_reg = odiv3_out_delay;
            3'b010: clkout2_reg = odiv0_out_delay;
            3'b011: clkout2_reg = odiv1_out_delay;
            3'b100: clkout2_reg = clk_in;
        endcase
    end

    always @(*)
    begin
        case(clkout3_sel)
            3'b000: clkout3_reg = odiv3_out_delay;
            3'b001: clkout3_reg = odiv0_out_delay;
            3'b010: clkout3_reg = odiv1_out_delay;
            3'b011: clkout3_reg = odiv2_out_delay;
            3'b100: clkout3_reg = clk_in;
        endcase
    end
////////////////////////////////////////////////////////////////////////////////////
////CLK_ENABLE//////////////////////////////////////////////////////////////////////
    assign clkout0_gate = clkout0_gate_en & CLKOUT0_SYN ;
    assign clkout1_gate = clkout1_gate_en & CLKOUT1_SYN ;
    assign clkout2_gate = clkout2_gate_en & CLKOUT2_SYN;
    assign clkout3_gate = clkout3_gate_en & CLKOUT3_SYN;
    
    always @(negedge clkout0_reg or negedge rst_n)
    begin
        if(!rst_n)
            clkout0_gate_d <= 3'b000;
        else
            clkout0_gate_d <= {clkout0_gate_d[1:0],~clkout0_gate};
    end

    always @(negedge clkout1_reg or negedge rst_n)
    begin
        if(!rst_n)
            clkout1_gate_d <= 3'b000;
        else
            clkout1_gate_d <= {clkout1_gate_d[1:0],~clkout1_gate};
    end

    always @(negedge clkout2_reg or negedge rst_n)
    begin
        if(!rst_n)
            clkout2_gate_d <= 3'b000;
        else
            clkout2_gate_d <= {clkout2_gate_d[1:0],~clkout2_gate};
    end
    always @(negedge clkout3_reg or negedge rst_n)
    begin
        if(!rst_n)
            clkout3_gate_d <= 3'b000;
        else
            clkout3_gate_d <= {clkout3_gate_d[1:0],~clkout3_gate};
    end

    assign CLKOUT = clk_in;
    assign CLKOUT0 = clkout0_reg & clkout0_gate_d[2];
    assign CLKOUT1 = clkout1_reg & clkout1_gate_d[2];
    assign CLKOUT2 = clkout2_reg & clkout2_gate_d[2];
    assign CLKOUT3 = clkout3_reg & clkout3_gate_d[2];
///////////////////////////////////////////////////////
////APB////////////////////////////////////////////////
    always @(posedge APB_CLK or negedge APB_RST_N)
    begin
        if(!APB_RST_N)
        begin
            rstn_apb     <= 1'b0;
            rstn_apb_syn <= 1'b0;
        end
        else
        begin
            rstn_apb     <= 1'b1;
            rstn_apb_syn <= rstn_apb;
        end
    end

    always @(posedge APB_CLK)
    begin
        if(APB_WRITE && APB_SEL)
        begin
            case(APB_ADDR)
                5'h0  : fracn_div[7:0]    <= APB_WDATA;
                5'h1  : fracn_div[15:8]   <= APB_WDATA;
                5'h2  : idivider[7:0]     <= APB_WDATA;
                5'h3  : fdivider[7:0]     <= APB_WDATA;
                5'h4  : ratio0[7:0]       <= APB_WDATA;
                5'h5  : ratio1[7:0]       <= APB_WDATA;
                5'h6  : ratio2[7:0]       <= APB_WDATA;
                5'h7  : ratio3[7:0]       <= APB_WDATA;
                5'h8  : odiv0_cphase[7:0] <= APB_WDATA;
                5'h9  : odiv1_cphase[7:0] <= APB_WDATA;
                5'ha  : odiv2_cphase[7:0] <= APB_WDATA;
                5'hb  : odiv3_cphase[7:0] <= APB_WDATA;
                5'hc  : {clkout1_gate_en, clkout0_gate_en, odiv1_fphase[2:0], odiv0_fphase[2:0]} <= APB_WDATA;
                5'hd  : {clkout3_gate_en, clkout2_gate_en, odiv3_fphase[2:0], odiv2_fphase[2:0]} <= APB_WDATA;
                5'he  : {odiv3_clkin_sel[1:0], odiv2_clkin_sel[1:0], odiv1_clkin_sel[1:0], odiv0_clkin_sel[1:0]} <= APB_WDATA;
                5'hf  : {vcoclk_bypass1, vcoclk_bypass0, clkout1_sel[2:0], clkout0_sel[2:0]} <= APB_WDATA;
                5'h10 : {vcoclk_bypass3, vcoclk_bypass2, clkout3_sel[2:0], clkout2_sel[2:0]} <= APB_WDATA;
                5'h11 : {pwd_apb, rstodiv_apb, rstodiv3_en, rstodiv2_en, rst_en, rstodiv_en, pwd_en, stdby_en} <= APB_WDATA;
                5'h12 : {pfden_apb_en, phase_apb_en, cphasestep_n_apb, load_fphase_apb, fphasestep_n_apb, fphasedir_apb, phasesel_apb[1:0]} <= APB_WDATA;
                5'h13 : {pfden_en, pfden_apb, lock_mode, lock_accuracy[2:0], fracn_en, icp_base_trim} <= APB_WDATA;
            endcase
        end
    end
endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_OMSER8.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_OMSER8 #(
parameter WL_EXTEND = "FALSE",     //"TRUE"; "FALSE"
parameter GRS_EN = "TRUE", //"TRUE"; "FALSE" 
parameter LRS_EN = "TRUE"   //"TRUE"; "FALSE" 
)(
output  PADO,
output  PADT,
input [7:0] D,
input [3:0] T,
input RCLK,
input SERCLK,
input OCLK,
input RST
);

//synthesis translate_off
reg [7:0] d_rclk;
reg [3:0] t_rclk;
reg [7:0] capture_d_reg;
reg [3:0] capture_t_reg;
reg [7:0] shift_d_reg;
reg [3:0] shift_t_reg;
reg PADO_POS;
reg PADT_reg;
reg PADO_NEG;
wire shift_en_oclk;
reg [1:0] cnt;
reg [1:0] cnt_oclk;
reg shift_en_oclk_d;

initial begin
d_rclk           = 0;
t_rclk           = 0;
capture_d_reg    = 0;
capture_t_reg    = 0;
shift_d_reg      = 0;
shift_t_reg      = 0;
PADO_POS         = 0;
PADT_reg         = 0;
PADO_NEG         = 0;
cnt              = 0;
cnt_oclk         = 0;
shift_en_oclk_d  = 0;
end


assign global_rstn = (GRS_EN == "TRUE") ? GRS_INST.GRSNET : 1'b1; 
assign lsr_rstn = LRS_EN == "TRUE" ? (~RST) : 1'b1;

always @(posedge RCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn) begin
      d_rclk <= 0;
      t_rclk <= 0;
   end   
   else if (!lsr_rstn) begin
      d_rclk <= 0;
      t_rclk <= 0;
   end   
   else begin
      d_rclk <= D;
      t_rclk <= T;
   end   

always @(posedge SERCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn) begin
      cnt       <= 0;
   end
   else if (!lsr_rstn) begin
      cnt       <= 0;
   end   
   else begin
      cnt       <= cnt + 1;
   end
   
assign  capture_en  = cnt == 3;

always @(posedge SERCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn) begin
      capture_d_reg <= 0;
      capture_t_reg <= 0;
   end
   else if (!lsr_rstn) begin
      capture_d_reg <= 0;
      capture_t_reg <= 0;
   end   
   else begin
      if (capture_en) begin
         capture_d_reg <= d_rclk;
         capture_t_reg <= t_rclk;     
      end
   end 

always @(posedge OCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn) begin
      cnt_oclk        <= 0;
      shift_en_oclk_d <= 0;
   end
   else if (!lsr_rstn) begin
      cnt_oclk        <= 0;
      shift_en_oclk_d <= 0;
   end   
   else begin
      cnt_oclk        <= cnt_oclk + 1;
      shift_en_oclk_d <= shift_en_oclk;
   end

assign shift_en_oclk = cnt_oclk == 2;
assign shift_en = (WL_EXTEND == "FALSE") ? shift_en_oclk : shift_en_oclk_d;
   
always @(posedge OCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn) begin
      shift_d_reg <= 0;
      shift_t_reg <= 0;
   end   
   else if (!lsr_rstn) begin
      shift_d_reg <= 0;
      shift_t_reg <= 0;
   end   
   else if (shift_en) begin
      shift_d_reg <= capture_d_reg;
      shift_t_reg <= capture_t_reg;
   end
   else begin
      shift_d_reg <= {2'd0, shift_d_reg[7:2]};
      shift_t_reg <= {1'b0, shift_t_reg[3:1]};        
   end
   
always @(posedge OCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn) begin
      PADO_POS <= 0;
      PADT_reg <= 0;
   end
   else if (!lsr_rstn) begin
      PADO_POS <= 0;
      PADT_reg <= 0;
   end
   else begin
      PADO_POS <= shift_d_reg[1];
      PADT_reg <= shift_t_reg[0];     
   end           
   
always @(negedge OCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn) begin
      PADO_NEG <= 0;
   end
   else if (!lsr_rstn) begin
      PADO_NEG <= 0;
   end
   else begin
      PADO_NEG <= shift_d_reg[0];
   end           
   
assign PADO =  OCLK ? PADO_NEG : PADO_POS;
assign PADT = PADT_reg;

//synthesis translate_on

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_RES_CAL.v
//
// Functional description: IO buffer driver and termination impedance calibration in each bank.
//
// Parameter description:
//
// Port description:
//    CAL_DONE: it refers to whether calibration is done or not. 1:done, 0: in progress.
//    CLK: on die clock used to do calibration, it runs at 50MHz.
//    CAL_REQ: request signal, this is set by usr and need to be a pulse.
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_RES_CAL #(
    parameter BANK_LOC = "L0", // IO Bank location: L0/L1/L2/R0/R1/R2
    parameter [19:0] CAL_CODE = 20'b11111_11111_10000_10000,  // static code to set resistor at "STATIC_MODE"
    parameter CAL_MODE = "STATIC_MODE", //"STATIC_MODE","DYNAMIC_MODE","AUTO_MODE","AUTO_MODE2"
    parameter DDR_RES = "50" // "75","60","50","40"
)(
    output reg CAL_DONE,  // see "Port description" above 
    input CAL_REQ
) /* synthesis syn_black_box */ ;
  
    reg cal_en;
    reg cal_start;
    reg [10:0] counter;
    reg CLK;

  initial begin
    CLK = 1'b0;
    CAL_DONE = 1'b1;
    cal_start = 1'b0;
    counter = 11'b000_000_000_00;  
    cal_en = 1'b1;

    end

 always #10 CLK = ~CLK;

 always @( negedge CAL_REQ)
   begin
    if (cal_en == 1'b1) 
      begin
       CAL_DONE <= 1'b0;
      end
    else if(cal_en == 1'b0)
      begin
       CAL_DONE <= 1'b1;
      end
    else begin 
         end
   end

 always @( posedge CAL_REQ)
   begin
    if (cal_en == 1'b1) 
    cal_start <= 1'b1;
    else
    cal_start <= 1'b0;
   end

 always @(posedge CLK )
  begin
    if (!cal_start)
        counter <= 0;
    else 
        counter <= counter + 1;      
 end

 always @(*)
  begin
   if (counter == 11'b10000011010)  // 1050 cycle
   CAL_DONE = 1'b1;
  end

 always @(posedge CAL_DONE )
  begin
  cal_start <= 1'b0;
  end

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_DFF_E.v
//
// Functional description: D-type flip-flop with enable
//
// Parameter description:
//      INIT: init value
//
// Port description:
//      CE  : enable
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_DFF_E
#(
    parameter GRS_EN = "TRUE",
    parameter INIT = 1'b0
) (
    output reg Q,
    input wire D,
    input wire CLK, CE
);

    wire grs_n;
    wire RS;

    tri1 grsnet = GRS_INST.GRSNET;
    assign grs_n=(GRS_EN=="TRUE")?grsnet:1'b1;

    not (RS, grs_n);

    initial Q = 1'bx;

    always @(posedge CLK or posedge RS) begin
        if (RS)
            Q <= 1'b0;
        else if (CE)
            Q <= D;
    end

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_IODELAY.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_IODELAY #(
parameter [6:0] DELAY_STEP = 7'h00,
parameter integer DELAY_DEPTH = 7 
)(
output DO,
output DELAY_OB,
input  DI,
input  LOAD_N,
input  MOVE,
input  DIRECTION
) /* synthesis syn_black_box */ ;

//synthesis translate_off
reg [DELAY_DEPTH-1:0] DELAY_UNIT;

localparam integer DELAY_UB = 2**DELAY_DEPTH-1;

initial begin
   if(DELAY_DEPTH != 7 && DELAY_DEPTH != 4)
   begin
     $display("GTP_IODELAY Error: Illegal setting of DELAY_DEPTH %s, ONLY 7 or 4 supported",DELAY_DEPTH);
     $finish;
   end
   if(DELAY_STEP > DELAY_UB || DELAY_STEP < 0)
   begin
     $display("GTP_IODELAY Error: Illegal range of DELAY_STEP %s", DELAY_STEP);
     $finish;
   end
   DELAY_UNIT = 0;
end

always @(DELAY_STEP or LOAD_N) 
begin
   if (!LOAD_N)
      DELAY_UNIT <= DELAY_STEP;
end

always @(negedge MOVE)
begin
   if (!LOAD_N)
      DELAY_UNIT <= DELAY_STEP;
   else if (DIRECTION && (DELAY_UNIT != 0))
      DELAY_UNIT <= DELAY_UNIT - 1;
   else if ((~DIRECTION) && (DELAY_UNIT != DELAY_UB))
      DELAY_UNIT <= DELAY_UNIT + 1;
end

assign DELAY_OB = (DIRECTION && (DELAY_UNIT == 0)) || ((~DIRECTION) && (DELAY_UNIT == DELAY_UB));

wire [DELAY_UB:0] delay_chain;
assign delay_chain[0] = DI;
genvar gen_i;
generate  
   for(gen_i=1;gen_i< DELAY_UB + 1;gen_i=gen_i+1) 
   begin
      assign #0.025 delay_chain[gen_i] =  delay_chain[gen_i-1];
   end
endgenerate

assign DO = delay_chain[DELAY_UNIT];

//synthesis translate_on

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: Internal simulation model
// Filename: GTP_IOBUF.v
//
// Functional description: Input/Output Buffer
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_IOBUF #(
    parameter IOSTANDARD = "DEFAULT",
    parameter SLEW_RATE = "SLOW",
    parameter DRIVE_STRENGTH = "8",
    parameter TERM_DDR = "ON"
)(
    output O,
    inout IO,
    input I,
    input T
) /* synthesis syn_black_box */ ;

  initial begin
    case (IOSTANDARD)
    "LVTTL33", "PCI33", "LVCMOS33", "LVCMOS25", "LVCMOS18", "LVCMOS15", "LVCMOS12", "SSTL25_I", "SSTL25_II", "SSTL18_I", "SSTL18_II", "SSTL15_I", "SSTL15_II", "HSTL18_I", "HSTL18_II", "HSTL15_I", "SSTL15_I_CAL", "SSTL15_II_CAL", "HSTL15_I_CAL", "DEFAULT" :;
    default : begin
           $display("Attribute Syntax Error : The attribute IOSTANDARD on GTP_IOBUF instance %m is set to %s.", IOSTANDARD);
           $finish;
              end
    endcase

    case (SLEW_RATE)
    "FAST", "SLOW":;
    default : begin
           $display("Attribute Syntax Error : The attribute SLEW_RATE on GTP_IOBUF instance %m is set to %s.", SLEW_RATE);
           $finish;
              end
    endcase

    case (DRIVE_STRENGTH)
    "2", "4", "6", "8", "12", "16", "24":;
    default : begin
           $display("Attribute Syntax Error : The attribute DRIVE_STRENGTH on GTP_IOBUF instance %m is set to %s.", DRIVE_STRENGTH);
           $finish;
              end
    endcase

    case (TERM_DDR)
    "ON", "OFF" :;
    default : begin
           $display("Attribute Syntax Error : The attribute TERM_DDR on GTP_IOBUF instance %m is set to %s.", TERM_DDR);
           $finish;
              end
    endcase
    end

    buf (O, IO);

    bufif0 (IO, I, T);

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2016 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_OSERDES_E2.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//////////////////////////////////////////////////////////////////////////////
`timescale 1ps / 1ps

module GTP_OSERDES_E2 #(
	parameter         GRS_EN          =  "TRUE",        // "TRUE","FALSE"   
	parameter         OSERDES_MODE    =  "SDR4TO1",     // "SDR2TO1","SDR3TO1","SDR4TO1","SDR5TO1","SDR6TO1","SDR7TO1","SDR8TO1",
                                                        // "DDR2TO1_SAME_EDGE","DDR2TO1_OPPOSITE_EDGE",
                                                        // "DDR4TO1","DDR8TO1","DDR10TO1","DDR14TO1",
                                                        // "HMSDR4TO1","HMSDR8TO1","OLATCH","ODFF",
                                                        
	parameter         TSERDES_EN      =  "FALSE",     // "FALSE","TRUE"
	parameter         UPD0_SHIFT_EN   =  "FALSE",     // "FALSE","TRUE"
	parameter         UPD1_SHIFT_EN   =  "FALSE",     // "FALSE","TRUE"
	parameter [1:0]   INIT_SET        =  2'b00,         // 2'b00,2'b01,2'b10,2'b11
	parameter         GRS_TYPE_DQ     =  "RESET",       // "RESET" "SET"
	parameter         LRS_TYPE_DQ0    =  "ASYNC_RESET", // ASYNC_SET  ASYNC_RESET  SYNC_SET SYNC_RESET  
	parameter         LRS_TYPE_DQ1    =  "ASYNC_RESET", // ASYNC_SET  ASYNC_RESET  SYNC_SET SYNC_RESET
	parameter         LRS_TYPE_DQ2    =  "ASYNC_RESET", // ASYNC_SET  ASYNC_RESET  SYNC_SET SYNC_RESET
	parameter         LRS_TYPE_DQ3    =  "ASYNC_RESET", // ASYNC_SET  ASYNC_RESET  SYNC_SET SYNC_RESET
	parameter         GRS_TYPE_TQ     =  "RESET",       // "RESET" "SET"
	parameter         LRS_TYPE_TQ0    =  "ASYNC_RESET", // ASYNC_SET  ASYNC_RESET  SYNC_SET SYNC_RESET    
	parameter         LRS_TYPE_TQ1    =  "ASYNC_RESET", // ASYNC_SET  ASYNC_RESET  SYNC_SET SYNC_RESET
	parameter         LRS_TYPE_TQ2    =  "ASYNC_RESET", // ASYNC_SET  ASYNC_RESET  SYNC_SET SYNC_RESET
	parameter         LRS_TYPE_TQ3    =  "ASYNC_RESET", // ASYNC_SET  ASYNC_RESET  SYNC_SET SYNC_RESET
	parameter         TRI_EN          =  "FALSE",     // "FALSE","TRUE"
	parameter         TBYTE_EN        =  "FALSE",     // "FALSE","TRUE"
	parameter         MIPI_EN         =  "FALSE",     // "FALSE","TRUE"
	parameter         OCASCADE_EN     =  "FALSE"      // "FALSE","TRUE"

)(
    //input         GRS_N,
    input         RST,
    input         OCE,
    input         TCE,
    input         OCLKDIV,
    //input         OCLKDIVB,
    input         SERCLK,
    //input         SERCLKB,
    input         OCLK,
    //input         OCLKB,
    input         MIPI_CTRL,
    input         UPD0_SHIFT,
    input         UPD1_SHIFT,
    input         OSHIFTIN0,
    input         OSHIFTIN1,
    input [7:0]   DI,
    input [1:0]   TI,
    input         TBYTE_IN,
    output        OSHIFTOUT0,
    output        OSHIFTOUT1,
    output        TQ,
    output        DO

);

wire         osr_iolhr;
wire         gwen;
wire         glogen;
wire         grs_n;
wire         oce;
wire         tce;
wire         oclkdiv;
wire         oclkdivb;
wire         serclk;
wire         serclkb;
wire         oclk;
wire         oclkb;
wire         mipi_sw_dyn_i;
wire         inbuf_dyn_dis_n_i;
wire         upd0_shift;
wire         upd1_shift;
wire         do_cas_in;
wire         oshiftin0;
wire         oshiftin1;
wire [7:0]   tx_data;
wire [1:0]   ts_ctrl;
wire         tbyte_in;
wire         termbyte_in;      
wire         to_cas_in;
wire         term_cas_in;
wire         dly_odly_in;
wire         oshiftout0;
wire         oshiftout1;
wire         do_p;
wire         to;
///////////////////////////////////////////// sc --> cp /////////////
reg  [3:0]   sc_oserdes_mode;
wire         sc_osr_pol;
wire         sc_sro_en;
wire         sc_srt_en;
//wire         sc_t_sync;
wire         sc_grs_dis;
wire         sc_clk_pol4;
wire         sc_clk_pol5;
wire         sc_clk_pol6;
wire         sc_upd0_shiften;
wire         sc_upd1_shiften;
wire [1:0]   sc_init_set;
wire         sc_tbyte_en;
wire         sc_mipi_en;
wire         sc_pdiff;
wire         sc_do_sel;       //used in mipi application
wire         sc_ocascade_en;
wire         sc_tri_en;
wire         sc_odly_en;
wire [1:0]   sc_dqmode;

reg  [1:0]   sc_dqmode_reg;
reg  [1:0]   sc_tqmode;
reg          sc_o_sync;
reg          sc_t_sync;
reg          sc_init_dq;
reg          sc_init_tq;
reg  [3:0]   sc_srval_dq;
reg  [3:0]   sc_srval_tq;
reg          sc_oserdes_en;
reg          sc_ser_ddren;
reg          sc_ser_sdren;
reg          sc_ohsmem_en;
reg          sc_opposite_en;
reg          sc_olthen;
reg          sc_odffen;


// parameter
assign  sc_osr_pol       =  1'b0;
assign  sc_sro_en		 =  1'b1;
assign  sc_srt_en		 =  1'b1;
//assign  sc_t_sync		 =  1'b0;
assign  sc_grs_dis		 = (GRS_EN=="TRUE")    ? 1'b0 : 1'b1;
assign  sc_clk_pol4		 =  1'b0;
assign  sc_clk_pol5		 =  1'b0;
assign  sc_clk_pol6		 =  1'b0;
assign  sc_upd0_shiften	 = (UPD0_SHIFT_EN=="FALSE") ? 1'b0 : 1'b1;
assign  sc_upd1_shiften	 = (UPD1_SHIFT_EN=="FALSE") ? 1'b0 : 1'b1;
assign  sc_init_set		 =  INIT_SET;
assign  sc_tbyte_en		 = (TBYTE_EN    =="FALSE") ? 1'b0 : 1'b1;
assign  sc_mipi_en		 = (MIPI_EN     =="FALSE") ? 1'b0 : 1'b1;
assign  sc_pdiff		 =  1'b0;
assign  sc_do_sel		 =  1'b0;       //used in mipi application
assign  sc_ocascade_en	 = (OCASCADE_EN =="FALSE") ? 1'b0 : 1'b1;
assign  sc_tri_en   	 = (TRI_EN =="FALSE") ? 1'b0 : 1'b1;
assign  sc_odly_en		 = 1'b0;
assign  sc_dqmode	     = sc_mipi_en ? 2'b00 : sc_dqmode_reg;



// input
assign  gwen             = 1'b1;
assign  glogen           = 1'b1;
assign  grs_n            = (GRS_EN == "TRUE") ? GRS_INST.GRSNET : 1'b1;
//assign  grs_n            =  1'b1;
//assign  grs_n            =  GRS_N;

assign  osr_iolhr	      = RST;
assign  oce		          = OCE;
assign  tce		          = TCE;
assign  oclkdiv		      = OCLKDIV;
assign  oclkdivb	      = ~OCLKDIV;
assign  serclk		      = SERCLK;
assign  serclkb		      = ~SERCLK;
assign  oclk		      = OCLK;
assign  oclkb		      = ~OCLK;
assign  mipi_sw_dyn_i     = MIPI_CTRL;
assign  inbuf_dyn_dis_n_i = 1'b0;
assign  upd0_shift		  = UPD0_SHIFT;
assign  upd1_shift		  = UPD1_SHIFT;
assign  do_cas_in		  = 1'b0;
assign  oshiftin0		  = OSHIFTIN0;
assign  oshiftin1		  = OSHIFTIN1;
assign  tx_data		      = DI;
assign  ts_ctrl		      = TI;
assign  tbyte_in		  = TBYTE_IN;
assign  termbyte_in		  = 1'b0;      
assign  to_cas_in		  = 1'b0;
assign  term_cas_in		  = 1'b0;
assign  dly_odly_in		  = 1'b0;

// output
assign  OSHIFTOUT0		  = oshiftout0;
assign  OSHIFTOUT1		  = oshiftout1;
assign  DO		          = do_p;
assign  TQ		          = to;

initial begin
    if(GRS_EN != "TRUE" && GRS_EN != "FALSE")
    begin $display("Error: Illegal setting GRS_EN of %s",GRS_EN);$finish;end

    if(UPD0_SHIFT_EN != "TRUE" && UPD0_SHIFT_EN != "FALSE")
    begin $display("Error: Illegal setting UPD0_SHIFT_EN of %s",UPD0_SHIFT_EN);$finish;end

    if(UPD1_SHIFT_EN != "TRUE" && UPD1_SHIFT_EN != "FALSE")
    begin $display("Error: Illegal setting UPD1_SHIFT_EN of %s",UPD1_SHIFT_EN);$finish;end

    if(INIT_SET != 2'b00 && INIT_SET != 2'b01 && INIT_SET != 2'b10 && INIT_SET != 2'b11)
    begin $display("Error: Illegal setting INIT_SET of %b",INIT_SET);$finish;end

    if(GRS_TYPE_DQ != "RESET" && GRS_TYPE_DQ != "SET")
    begin $display("Error: Illegal setting GRS_TYPE_DQ of %s",GRS_TYPE_DQ);$finish;end



    if(LRS_TYPE_DQ0 != "ASYNC_RESET" && LRS_TYPE_DQ0 != "ASYNC_SET" && LRS_TYPE_DQ0 != "SYNC_RESET" && LRS_TYPE_DQ0 != "SYNC_SET")
    begin $display("Error: Illegal setting LRS_TYPE_DQ0 of %s",LRS_TYPE_DQ0);$finish;end

    if(LRS_TYPE_DQ1 != "ASYNC_RESET" && LRS_TYPE_DQ1 != "ASYNC_SET" && LRS_TYPE_DQ1 != "SYNC_RESET" && LRS_TYPE_DQ1 != "SYNC_SET")
    begin $display("Error: Illegal setting LRS_TYPE_DQ1 of %s",LRS_TYPE_DQ1);$finish;end

    if(LRS_TYPE_DQ2 != "ASYNC_RESET" && LRS_TYPE_DQ2 != "ASYNC_SET" && LRS_TYPE_DQ2 != "SYNC_RESET" && LRS_TYPE_DQ2 != "SYNC_SET")
    begin $display("Error: Illegal setting LRS_TYPE_DQ2 of %s",LRS_TYPE_DQ2);$finish;end

    if(LRS_TYPE_DQ3 != "ASYNC_RESET" && LRS_TYPE_DQ3 != "ASYNC_SET" && LRS_TYPE_DQ3 != "SYNC_RESET" && LRS_TYPE_DQ3 != "SYNC_SET")
    begin $display("Error: Illegal setting LRS_TYPE_DQ3 of %s",LRS_TYPE_DQ3);$finish;end



    if(GRS_TYPE_TQ != "RESET" && GRS_TYPE_TQ != "SET")
    begin $display("Error: Illegal setting GRS_TYPE_TQ of %s",GRS_TYPE_TQ);$finish;end



    if(LRS_TYPE_TQ0 != "ASYNC_RESET" && LRS_TYPE_TQ0 != "ASYNC_SET" && LRS_TYPE_TQ0 != "SYNC_RESET" && LRS_TYPE_TQ0 != "SYNC_SET")
    begin $display("Error: Illegal setting LRS_TYPE_TQ0 of %s",LRS_TYPE_TQ0);$finish;end

    if(LRS_TYPE_TQ1 != "ASYNC_RESET" && LRS_TYPE_TQ1 != "ASYNC_SET" && LRS_TYPE_TQ1 != "SYNC_RESET" && LRS_TYPE_TQ1 != "SYNC_SET")
    begin $display("Error: Illegal setting LRS_TYPE_TQ1 of %s",LRS_TYPE_TQ1);$finish;end

    if(LRS_TYPE_TQ2 != "ASYNC_RESET" && LRS_TYPE_TQ2 != "ASYNC_SET" && LRS_TYPE_TQ2 != "SYNC_RESET" && LRS_TYPE_TQ2 != "SYNC_SET")
    begin $display("Error: Illegal setting LRS_TYPE_TQ2 of %s",LRS_TYPE_TQ2);$finish;end

    if(LRS_TYPE_TQ3 != "ASYNC_RESET" && LRS_TYPE_TQ3 != "ASYNC_SET" && LRS_TYPE_TQ3 != "SYNC_RESET" && LRS_TYPE_TQ3 != "SYNC_SET")
    begin $display("Error: Illegal setting LRS_TYPE_TQ3 of %s",LRS_TYPE_TQ3);$finish;end



    if((LRS_TYPE_DQ0 == "ASYNC_RESET" || LRS_TYPE_DQ0 == "ASYNC_SET" || LRS_TYPE_DQ1 == "ASYNC_RESET" || LRS_TYPE_DQ1 == "ASYNC_SET" 
        || LRS_TYPE_DQ2 == "ASYNC_RESET" || LRS_TYPE_DQ2 == "ASYNC_SET" || LRS_TYPE_DQ3 == "ASYNC_RESET" || LRS_TYPE_DQ3 == "ASYNC_SET") 
        && (LRS_TYPE_DQ0 == "SYNC_RESET" || LRS_TYPE_DQ0 == "SYNC_SET" || LRS_TYPE_DQ1 == "SYNC_RESET" || LRS_TYPE_DQ1 == "SYNC_SET" 
        ||  LRS_TYPE_DQ2 == "SYNC_RESET" || LRS_TYPE_DQ2 == "SYNC_SET" || LRS_TYPE_DQ3 == "SYNC_RESET" || LRS_TYPE_DQ3 == "SYNC_SET"))
    begin $display("Error: LRS_TYPE_DQx must be all of ASYNC_ or SYNC_.");$finish;end


    if((LRS_TYPE_TQ0 == "ASYNC_RESET" || LRS_TYPE_TQ0 == "ASYNC_SET" || LRS_TYPE_TQ1 == "ASYNC_RESET" || LRS_TYPE_TQ1 == "ASYNC_SET" 
        || LRS_TYPE_TQ2 == "ASYNC_RESET" || LRS_TYPE_TQ2 == "ASYNC_SET" || LRS_TYPE_TQ3 == "ASYNC_RESET" || LRS_TYPE_TQ3 == "ASYNC_SET") 
        && (LRS_TYPE_TQ0 == "SYNC_RESET" || LRS_TYPE_TQ0 == "SYNC_SET" || LRS_TYPE_TQ1 == "SYNC_RESET" || LRS_TYPE_TQ1 == "SYNC_SET" 
        ||  LRS_TYPE_TQ2 == "SYNC_RESET" || LRS_TYPE_TQ2 == "SYNC_SET" || LRS_TYPE_TQ3 == "SYNC_RESET" || LRS_TYPE_TQ3 == "SYNC_SET"))
    begin $display("Error: LRS_TYPE_TQx must be all of ASYNC_ or SYNC_.");$finish;end



    if(TBYTE_EN != "TRUE" && TBYTE_EN != "FALSE")
    begin $display("Error: Illegal setting TBYTE_EN of %s",TBYTE_EN);$finish;end

    if(MIPI_EN != "TRUE" && MIPI_EN != "FALSE")
    begin $display("Error: Illegal setting MIPI_EN of %s",MIPI_EN);$finish;end

    if(OCASCADE_EN != "TRUE" && OCASCADE_EN != "FALSE")
    begin $display("Error: Illegal setting OCASCADE_EN of %s",OCASCADE_EN);$finish;end

    if(TRI_EN != "TRUE" && TRI_EN != "FALSE")
    begin $display("Error: Illegal setting TRI_EN of %s",TRI_EN);$finish;end

    if((TSERDES_EN == "TRUE")) begin
        if(OSERDES_MODE == "SDR2TO1" || OSERDES_MODE == "SDR4TO1" || OSERDES_MODE == "SDR8TO1" 
            || OSERDES_MODE == "DDR4TO1" || OSERDES_MODE == "DDR8TO1" 
            || OSERDES_MODE == "HMSDR4TO1" || OSERDES_MODE == "HMSDR8TO1")
            ;
        else begin $display("Error: Illegal setting OSERDES_MODE of %s when TSERDES_EN == TRUE",OSERDES_MODE);$finish;end
    end
end


// sc_oserdes_mode
initial begin
// default value
    sc_oserdes_mode = 4'b0000;
    sc_dqmode_reg	= 2'b00;
    sc_tqmode       = 2'b00;
    sc_oserdes_en   = 1'b0;
    sc_ser_sdren    = 1'b0;
    sc_ser_ddren    = 1'b0;
    sc_ohsmem_en    = 1'b0;
    sc_opposite_en  = 1'b0;
    sc_olthen       = 1'b0;
    sc_odffen       = 1'b0;
//
    case (OSERDES_MODE)
// SDR
        "SDR2TO1" :begin
                    sc_oserdes_mode = 4'b0101;
                    sc_dqmode_reg	= 2'b01;
                    sc_tqmode       = 2'b01;
                    sc_oserdes_en   = 1'b1;
                    sc_ser_sdren    = 1'b1;
                   end 
        "SDR3TO1" :begin
                    sc_oserdes_mode = 4'b0110;
                    sc_dqmode_reg	= 2'b01;
                    sc_tqmode       = 2'b01;
                    sc_oserdes_en   = 1'b1;
                    sc_ser_sdren    = 1'b1;
                   end 
        "SDR4TO1" :begin
                    sc_oserdes_mode = 4'b0000;
                    sc_dqmode_reg	= 2'b01;
                    sc_tqmode       = 2'b01;
                    sc_oserdes_en   = 1'b1;
                    sc_ser_sdren    = 1'b1;
                   end 
        "SDR5TO1" :begin
                    sc_oserdes_mode = 4'b0011;
                    sc_dqmode_reg	= 2'b01;
                    sc_tqmode       = 2'b01;
                    sc_oserdes_en   = 1'b1;
                    sc_ser_sdren    = 1'b1;
                   end 
        "SDR6TO1" :begin
                    sc_oserdes_mode = 4'b1000;
                    sc_dqmode_reg	= 2'b01;
                    sc_tqmode       = 2'b01;
                    sc_oserdes_en   = 1'b1;
                    sc_ser_sdren    = 1'b1;
                   end 
        "SDR7TO1" :begin
                    sc_oserdes_mode = 4'b0010;
                    sc_dqmode_reg	= 2'b01;
                    sc_tqmode       = 2'b01;
                    sc_oserdes_en   = 1'b1;
                    sc_ser_sdren    = 1'b1;
                   end 
        "SDR8TO1" :begin
                    sc_oserdes_mode = 4'b0001;
                    sc_dqmode_reg	= 2'b01;
                    sc_tqmode       = 2'b01;
                    sc_oserdes_en   = 1'b1;
                    sc_ser_sdren    = 1'b1;
                   end 
// DDR  
        "OLATCH" :begin
                    sc_dqmode_reg	= 2'b01;
                    sc_tqmode       = 2'b01;
                    sc_oserdes_en   = 1'b0;
                    sc_olthen       = 1'b1;
                   end 
        "ODFF" :begin
                    sc_dqmode_reg	= 2'b01;
                    sc_tqmode       = 2'b01;
                    sc_oserdes_en   = 1'b0;
                    sc_odffen       = 1'b1;
                   end 
        "DDR2TO1_SAME_EDGE" :begin
                    sc_oserdes_en   = 1'b0;
                    sc_dqmode_reg	= 2'b10;
                    sc_tqmode       = 2'b10;
                    sc_ser_ddren    = 1'b1;
                    sc_opposite_en  = 1'b0;
                   end 
        "DDR2TO1_OPPOSITE_EDGE" :begin
                    sc_oserdes_en   = 1'b0;
                    sc_dqmode_reg	= 2'b10;
                    sc_tqmode       = 2'b10;
                    sc_ser_ddren    = 1'b1;
                    sc_opposite_en  = 1'b1;
                   end 
        "DDR4TO1" :begin
                    sc_oserdes_mode = 4'b0000;
                    sc_dqmode_reg	= 2'b10;
                    sc_tqmode       = 2'b10;
                    sc_oserdes_en   = 1'b1;
                    sc_ser_ddren    = 1'b1;
                   end 
        "DDR6TO1" :begin
                    sc_oserdes_mode = 4'b1000;
                    sc_dqmode_reg	= 2'b10;
                    sc_tqmode       = 2'b10;
                    sc_oserdes_en   = 1'b1;
                    sc_ser_ddren    = 1'b1;
                   end 
        "DDR8TO1" :begin
                    sc_oserdes_mode = 4'b0001;
                    sc_dqmode_reg	= 2'b10;
                    sc_tqmode       = 2'b10;
                    sc_oserdes_en   = 1'b1;
                    sc_ser_ddren    = 1'b1;
                   end 
        "DDR10TO1" :begin
                    sc_oserdes_mode = 4'b0100;
                    sc_dqmode_reg	= 2'b10;
                    sc_tqmode       = 2'b10;
                    sc_oserdes_en   = 1'b1;
                    sc_ser_ddren    = 1'b1;
                   end 
        "DDR14TO1" :begin
                    sc_oserdes_mode = 4'b0111;
                    sc_dqmode_reg	= 2'b10;
                    sc_tqmode       = 2'b10;
                    sc_oserdes_en   = 1'b1;
                    sc_ser_ddren    = 1'b1;
                   end 
// High Speed Memory 
//         "HMSDR2TO1" :begin
//                     sc_ser_sdren    = 1'b1;
//                     sc_ohsmem_en    = 1'b1;
//                    end 
        "HMSDR4TO1" :begin
                    sc_oserdes_mode = 4'b0000;
                    sc_dqmode_reg	= 2'b01;
                    sc_tqmode       = 2'b01;
                    sc_oserdes_en   = 1'b1;
                    sc_ser_sdren    = 1'b1;
                    sc_ohsmem_en    = 1'b1;
                   end
        "HMSDR8TO1" :begin
                    sc_oserdes_mode = 4'b0001;
                    sc_dqmode_reg	= 2'b01;
                    sc_tqmode       = 2'b01;
                    sc_oserdes_en   = 1'b1;
                    sc_ser_sdren    = 1'b1;
                    sc_ohsmem_en    = 1'b1;
                   end
        default:    begin 
                    sc_oserdes_mode = 4'b0000; 
                    $display("Error: Illegal setting OSERDES_MODE of %s",OSERDES_MODE);
                    $finish; 
                    end
        endcase
end

initial begin
    case (GRS_TYPE_DQ)
        "SET"  :begin sc_init_dq=1'b1; end
        "RESET":begin sc_init_dq=1'b0; end
    endcase
end

initial begin
    case (LRS_TYPE_DQ0)
        "ASYNC_SET"  :begin sc_o_sync=1'b0; sc_srval_dq[0]=1'b1; end
        "ASYNC_RESET":begin sc_o_sync=1'b0; sc_srval_dq[0]=1'b0; end
        "SYNC_SET"   :begin sc_o_sync=1'b1; sc_srval_dq[0]=1'b1; end
        "SYNC_RESET" :begin sc_o_sync=1'b1; sc_srval_dq[0]=1'b0; end
    endcase
end

initial begin
    case (LRS_TYPE_DQ1)
        "ASYNC_SET"  :begin sc_o_sync=1'b0; sc_srval_dq[1]=1'b1; end
        "ASYNC_RESET":begin sc_o_sync=1'b0; sc_srval_dq[1]=1'b0; end
        "SYNC_SET"   :begin sc_o_sync=1'b1; sc_srval_dq[1]=1'b1; end
        "SYNC_RESET" :begin sc_o_sync=1'b1; sc_srval_dq[1]=1'b0; end
    endcase
end

initial begin
    case (LRS_TYPE_DQ2)
        "ASYNC_SET"  :begin sc_o_sync=1'b0; sc_srval_dq[2]=1'b1; end
        "ASYNC_RESET":begin sc_o_sync=1'b0; sc_srval_dq[2]=1'b0; end
        "SYNC_SET"   :begin sc_o_sync=1'b1; sc_srval_dq[2]=1'b1; end
        "SYNC_RESET" :begin sc_o_sync=1'b1; sc_srval_dq[2]=1'b0; end
    endcase
end

initial begin
    case (LRS_TYPE_DQ3)
        "ASYNC_SET"  :begin sc_o_sync=1'b0; sc_srval_dq[3]=1'b1; end
        "ASYNC_RESET":begin sc_o_sync=1'b0; sc_srval_dq[3]=1'b0; end
        "SYNC_SET"   :begin sc_o_sync=1'b1; sc_srval_dq[3]=1'b1; end
        "SYNC_RESET" :begin sc_o_sync=1'b1; sc_srval_dq[3]=1'b0; end
    endcase
end

initial begin
    case (GRS_TYPE_TQ)
        "SET"  :begin sc_init_tq=1'b1; end
        "RESET":begin sc_init_tq=1'b0; end
    endcase
end

initial begin
    case (LRS_TYPE_TQ0)
        "ASYNC_SET"  :begin sc_t_sync=1'b0; sc_srval_tq[0]=1'b1; end
        "ASYNC_RESET":begin sc_t_sync=1'b0; sc_srval_tq[0]=1'b0; end
        "SYNC_SET"   :begin sc_t_sync=1'b1; sc_srval_tq[0]=1'b1; end
        "SYNC_RESET" :begin sc_t_sync=1'b1; sc_srval_tq[0]=1'b0; end
    endcase
end

initial begin
    case (LRS_TYPE_TQ1)
        "ASYNC_SET"  :begin sc_t_sync=1'b0; sc_srval_tq[1]=1'b1; end
        "ASYNC_RESET":begin sc_t_sync=1'b0; sc_srval_tq[1]=1'b0; end
        "SYNC_SET"   :begin sc_t_sync=1'b1; sc_srval_tq[1]=1'b1; end
        "SYNC_RESET" :begin sc_t_sync=1'b1; sc_srval_tq[1]=1'b0; end
    endcase
end

initial begin
    case (LRS_TYPE_TQ2)
        "ASYNC_SET"  :begin sc_t_sync=1'b0; sc_srval_tq[2]=1'b1; end
        "ASYNC_RESET":begin sc_t_sync=1'b0; sc_srval_tq[2]=1'b0; end
        "SYNC_SET"   :begin sc_t_sync=1'b1; sc_srval_tq[2]=1'b1; end
        "SYNC_RESET" :begin sc_t_sync=1'b1; sc_srval_tq[2]=1'b0; end
    endcase
end

initial begin
    case (LRS_TYPE_TQ3)
        "ASYNC_SET"  :begin sc_t_sync=1'b0; sc_srval_tq[3]=1'b1; end
        "ASYNC_RESET":begin sc_t_sync=1'b0; sc_srval_tq[3]=1'b0; end
        "SYNC_SET"   :begin sc_t_sync=1'b1; sc_srval_tq[3]=1'b1; end
        "SYNC_RESET" :begin sc_t_sync=1'b1; sc_srval_tq[3]=1'b0; end
    endcase
end

oserdes_e2_iolhr_ol xoserdes_e2_iolhr_ol(
               .sc_osr_pol(sc_osr_pol),
               .sc_sro_en(sc_sro_en),
               .sc_o_sync(sc_o_sync),
               .sc_srt_en(sc_srt_en),
               .sc_t_sync(sc_t_sync),
               .sc_grs_dis(sc_grs_dis),
               .sc_clk_pol4(sc_clk_pol4),
               .sc_clk_pol5(sc_clk_pol5),
               .sc_clk_pol6(sc_clk_pol6),
               .sc_opposite_en(sc_opposite_en),
               .sc_ohsmem_en(sc_ohsmem_en),
               .sc_oserdes_en(sc_oserdes_en),
               .sc_ser_ddren(sc_ser_ddren),
               .sc_ser_sdren(sc_ser_sdren),
               .sc_olthen(sc_olthen),
               .sc_odffen(sc_odffen),
               .sc_oserdes_mode(sc_oserdes_mode),
               .sc_upd0_shiften(sc_upd0_shiften),
               .sc_upd1_shiften(sc_upd1_shiften),
               .sc_init_set(sc_init_set),
               .sc_init_dq(sc_init_dq),
               .sc_srval_dq(sc_srval_dq),
               .sc_mipi_en(sc_mipi_en),
               .sc_pdiff(sc_pdiff),
               .sc_do_sel(sc_do_sel),       //used in mipi application
               .sc_ocascade_en(sc_ocascade_en),
               .sc_dqmode(sc_dqmode),
               .sc_tri_en(sc_tri_en),
               .sc_odly_en(sc_odly_en),
               .osr_iolhr(osr_iolhr),
                .gwen(gwen),
               .glogen(glogen),
               .grs_n(grs_n),
               //.por_n(por_n),
               .oce(oce),
               .tce(tce),
               .oclkdiv(oclkdiv),
               .oclkdivb(oclkdivb),
               .serclk(serclk),
               .serclkb(serclkb),
               .oclk(oclk),
               .oclkb(oclkb),
               .upd0_shift(upd0_shift),
               .upd1_shift(upd1_shift),
               .do_cas_in(do_cas_in),
               .oshiftin0(oshiftin0),
               .oshiftin1(oshiftin1),
               .tx_data(tx_data),
               .mipi_sw_dyn_i(mipi_sw_dyn_i),
               .inbuf_dyn_dis_n_i(inbuf_dyn_dis_n_i),
               .sc_srval_tq(sc_srval_tq),
               .sc_init_tq(sc_init_tq),
               .sc_tqmode(sc_tqmode),
               .sc_tbyte_en(sc_tbyte_en),
               .ts_ctrl(ts_ctrl),
               .tbyte_in(tbyte_in),
               .termbyte_in(termbyte_in),      
               .to_cas_in(to_cas_in),
               .term_cas_in(term_cas_in),
               .dly_odly_in(dly_odly_in),
               .term(),
               .tfb(),
               .term_fb(),
               .to_cas_out(),
               .term_cas_out(),
               .oshiftout0(oshiftout0),
               .oshiftout1(oshiftout1),
               .do_p(do_p),
               .do_n(),
               .to(to),
               .do_cas_out(),
               .ofb(),
               .mipi_sw_dyn_o(),
               .inbuf_dyn_dis_n_o()
              );

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_ROM256X1.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_ROM256X1
#(
    parameter [255:0] INIT = 256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000
) (
    output Z,
    input I0, I1, I2, I3, I4, I5, I6, I7
);

   reg [255:0] mem;
   wire [8:0] addr;

   initial mem = INIT;

   assign addr = {I7, I6, I5, I4, I3, I2, I1, I0};
   //assign Z = mem[addr];
   assign Z = INIT[addr];

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_LUT5M.v
//
// Functional description: 5-input Look-Up-Table for 4-to-1 Mux
//
// Parameter description:
//      INIT: init value
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_LUT5M
#(
    parameter [31:0] INIT = 32'h0000_0000
) (
    output wire Z,
    input wire I0, ID, I1, I2, I3, I4
);

    wire x7, x6, x5, x4, y1;
    wire x3, x2, x1, x0, y0;

    INT_LUTMUX4_UDP (x7, I1, I0, INIT[31], INIT[30], INIT[29], INIT[28]);
    INT_LUTMUX4_UDP (x6, I1, I0, INIT[27], INIT[26], INIT[25], INIT[24]);
    INT_LUTMUX4_UDP (x5, I1, I0, INIT[23], INIT[22], INIT[21], INIT[20]);
    INT_LUTMUX4_UDP (x4, I1, I0, INIT[19], INIT[18], INIT[17], INIT[16]);
    INT_LUTMUX4_UDP (y1, I3, I2, x7, x6, x5, x4);

    INT_LUTMUX4_UDP (x3, I1, ID, INIT[15], INIT[14], INIT[13], INIT[12]);
    INT_LUTMUX4_UDP (x2, I1, ID, INIT[11], INIT[10], INIT[9], INIT[8]);
    INT_LUTMUX4_UDP (x1, I1, ID, INIT[7], INIT[6], INIT[5], INIT[4]);
    INT_LUTMUX4_UDP (x0, I1, ID, INIT[3], INIT[2], INIT[1], INIT[0]);
    INT_LUTMUX4_UDP (y0, I3, I2, x3, x2, x1, x0);

    INT_LUTMUX2_UDP (Z, I4, y1, y0);

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_MULTADDACC18.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

//P = MAC + (A0*B0 + A1*B1)
module GTP_MULTADDACC18 #(
    parameter  GRS_EN            = "TRUE", //"TRUE"; "FALSE"
    parameter  SYNC_RST          = "FALSE", //"TRUE"; "FALSE"
    parameter  INREG_EN          = "FALSE",  //"TRUE"; "FALSE"
    parameter  PIPEREG_EN        = "FALSE",//"TRUE"; "FALSE"
    parameter  ADDSUB_OP         = 0 ,
    parameter  ACC_ADDSUB_OP     = 0,
    parameter  DYN_ADDSUB_OP     = 1,
    parameter  DYN_ACC_ADDSUB_OP = 1,
    parameter  OVERFLOW_MASK     = 64'h0, //PSZIE = 64 OVERflow setting = 'h20_0000_0000_0000, bit width = PSIZE
    parameter  PATTERN           = 64'h0,  //compare pattern
    parameter  MASKPAT           = 64'h0,  //pattern mask
    parameter  DYN_ACC_INIT      = 0,  //acc init value dynamic input
    parameter  ACC_INIT_VALUE    = 64'h0   //acc init value parameter
) (
    output  [63:0] P,
    output  OVER,
    output  UNDER,
    output  EQZ,
    output  EQZM,
    output  EQOM,
    output  EQPAT,
    output  EQPATN,

    input   CE,
    input   RST,
    input   CLK,
    input   A_SIGNED,
    input   [17:0] A0,
    input   [17:0] A1,
    input   B_SIGNED,
    input   [17:0] B0,
    input   [17:0] B1,
    input   [63:0] ACC_INIT,
    input   ADDSUB,
    input   ACC_ADDSUB,
    input   RELOAD
);

    wire [63:0] R;

    INT_PREADD_MULTADDACC #(
        . GRS_EN(GRS_EN),     
        . SYNC_RST(SYNC_RST),   
        . INREG_EN(INREG_EN),   
        . PIPEREG_EN(PIPEREG_EN), 
        . ADDSUB_OP(ADDSUB_OP),    
        . ACCUMADDSUB_OP(ACC_ADDSUB_OP),
        . DYN_OP_ADDSUB(DYN_ADDSUB_OP),   
        . DYN_OP_ACC(DYN_ACC_ADDSUB_OP),  
        . ASIZE(18), 
        . BSIZE(18), 
        . PSIZE(64), 
        . PREADD_EN(0),
        . MASK(OVERFLOW_MASK), 
        . DYN_ACC_INIT(DYN_ACC_INIT),
        . ACC_INIT_VALUE(ACC_INIT_VALUE)
    ) U_MACC (
        . CE(CE),
        . RST(RST),
        . CLK(CLK),
        . A_SIGNED(A_SIGNED),
        . A0(A0),
        . A1(A1),
        . B_SIGNED(B_SIGNED),
        . B0(B0),
        . B1(B1),
        . C_SIGNED(B_SIGNED),
        . C0(18'b0),
        . C1(18'b0),
        . PREADDSUB(2'b0),
        . ACCUM_INIT(ACC_INIT),
        . ADDSUB(ADDSUB),
        . ACCUMADDSUB(ACC_ADDSUB),
        . RELOAD(RELOAD),
        . P(P),
        . OVER(OVER),
        . UNDER(UNDER),
        . R(R) 
    );

    INT_FLAG #(
        . GRS_EN(GRS_EN),
        . SYNC_RST(SYNC_RST),
        . PSIZE(64),
        . PATSIZE(64),
        . MASKPATSIZE(64),
        . OUTREG_EN("TRUE")
    ) U_FLAG (
        . CE(CE),
        . RST(RST),
        . CLK(CLK),
        . P(P),
        . PATTERN(PATTERN),
        . MASKPAT(MASKPAT),
        . OVERFLOW_MASK(OVERFLOW_MASK),
        . R(R),
        . eqz(EQZ),
        . eqzm(EQZM),
        . eqom(EQOM),
        . eqpat(EQPAT),
        . eqpatn(EQPATN)
    );

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_LUT8.v
//
// Functional description: 8-input Look-Up-Table
//
// Parameter description:
//      INIT: init value
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_LUT8
#(
    parameter [255:0] INIT = 256'h0000000000000000_0000000000000000_0000000000000000_0000000000000000
) (
    output wire Z,
    input wire I0, I1, I2, I3, I4, I5, I6, I7
);

    wire z6a, z6b, z6c, z6d;
    wire z7ab, z7cd;

    GTP_LUT6 #(.INIT(INIT[63:0]))
        l6a (.I0(I0), .I1(I1), .I2(I2), .I3(I3), .I4(I4), .I5(I5), .Z(z6a));

    GTP_LUT6 #(.INIT(INIT[127:64]))
        l6b (.I0(I0), .I1(I1), .I2(I2), .I3(I3), .I4(I4), .I5(I5), .Z(z6b));

    GTP_MUX2LUT7 mxl7ab (.I0(z6a), .I1(z6b), .S(I6), .Z(z7ab));

    GTP_LUT6 #(.INIT(INIT[191:128]))
        l6c (.I0(I0), .I1(I1), .I2(I2), .I3(I3), .I4(I4), .I5(I5), .Z(z6c));

    GTP_LUT6 #(.INIT(INIT[255:192]))
        l6d (.I0(I0), .I1(I1), .I2(I2), .I3(I3), .I4(I4), .I5(I5), .Z(z6d));

    GTP_MUX2LUT7 mxl7cd (.I0(z6c), .I1(z6d), .S(I6), .Z(z7cd));

    GTP_MUX2LUT8 mxl8 (.I0(z7ab), .I1(z7cd), .S(I7), .Z(Z));

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_MUX2LUT8.v
//
// Functional description: 2-to-1 MUX to generate LUT8 func
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_MUX2LUT8
(
    output wire Z,
    input wire I0, I1, S
);

    INT_LUTMUX2_UDP (Z, S, I1, I0);

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////

//P = A0*(B0+-C0) +/- A1*(B1+-C1)
`timescale 1 ns / 1 ps

module INT_PREADD_MULTADD
#(
    parameter GRS_EN        = "FALSE", //"TRUE"; "FALSE"
    parameter SYNC_RST      = "FALSE", //"TRUE"; "FALSE"  
    parameter SIC0_EN       = "FALSE", //"TRUE"; "FALSE"  
    parameter SIB1_EN       = "FALSE", //"TRUE"; "FALSE"  
    parameter SIC1_EN       = "FALSE", //"TRUE"; "FALSE"  
    parameter INREG_EN      = "FALSE",  //"TRUE"; "FALSE"
    parameter PREREG_EN     = "FALSE",  //"TRUE"; "FALSE"
    parameter PIPEREG_EN    = "FALSE",  //"TRUE"; "FALSE"
    parameter OUTREG_EN     = "FALSE",   //"TRUE"; "FALSE"
    parameter ADDSUB_OP     = 0 ,
    parameter DYN_OP_ADDSUB = 1,
    parameter ASIZE         = 9,              // LEGAL ASIZE = 9,18,27,36
    parameter BSIZE         = 8,              // LEGAL BSIZE = 8,18,26,18
    //PSE parameters
    parameter [ASIZE-2:0] SC_PSE_A0 = 0, //SC_PSE = 0, disable PSE,  bit width = ASIZE-1
    parameter [ASIZE-2:0] SC_PSE_A1 = 0, //SC_PSE = 0, disable PSE,  bit width = ASIZE-1
    parameter [BSIZE-2:0] SC_PSE_B0 = 0, //SC_PSE = 0, disable PSE,  bit width = BSIZE-1
    parameter [BSIZE-2:0] SC_PSE_B1 = 0, //SC_PSE = 0, disable PSE,  bit width = BSIZE-1
    parameter [BSIZE-2:0] SC_PSE_C0 = 0, //SC_PSE = 0, disable PSE,  bit width = BSIZE-1
    parameter [BSIZE-2:0] SC_PSE_C1 = 0, //SC_PSE = 0, disable PSE,  bit width = BSIZE-1
    parameter integer PREADD_EN = 1,
    parameter integer PSIZE = ASIZE + BSIZE + 1 + PREADD_EN
) (
    input   CE,
    input   RST,
    input   CLK,
    input   [ASIZE-1:0] A0,
    input   [ASIZE-1:0] A1,
    input   [BSIZE-1:0] B0,
    input   [BSIZE-1:0] B1,
    input   [BSIZE-1:0] C0,
    input   [BSIZE-1:0] C1,
    input   A_SIGNED,
    input   B_SIGNED,
    input   C_SIGNED,
    input   [1:0] PREADDSUB,
    input   ADDSUB,
    output  [PSIZE-1:0] P
);

initial begin
    if ((PREADD_EN != 0) && (PREADD_EN != 1))
    begin
        $finish;
    end
    case (ASIZE)
        9:  if ((BSIZE + PREADD_EN) != 9)
            begin
                $finish;
            end
        18, 36: if (BSIZE != 18)
            begin
                $finish;
            end
        27: if ((BSIZE + PREADD_EN) != 27)
            begin
                $finish;
            end
        default :
            $finish;
    endcase
    //  $display (" INT_PREADD_MULTADD error :illegal setting of ASIZE or BSIZE");

    if ((GRS_EN != "TRUE") && (GRS_EN != "FALSE")) begin
        $display("GRS_EN error");
        $finish;
    end
    if ((SYNC_RST != "TRUE") && (SYNC_RST != "FALSE")) begin
        $display("SYNC_RST error");
        $finish;
    end

    if ((INREG_EN != "TRUE") && (INREG_EN != "FALSE")) begin
        $display("INREG_EN error");
        $finish;
    end
    if ((PREREG_EN != "TRUE") && (PREREG_EN != "FALSE")) begin
        $display("PREREG_EN error");
        $finish;
    end
    if ((PIPEREG_EN != "TRUE") && (PIPEREG_EN != "FALSE")) begin
        $display("PIPEREG_EN error");
        $finish;
    end
    if ((OUTREG_EN != "TRUE") && (OUTREG_EN != "FALSE")) begin
        $display("OUTREG_EN error");
        $finish;
    end

    if (SIB1_EN != "FALSE" || SIC0_EN != "FALSE" || SIC1_EN != "FALSE") begin
        $display("DRC error");
        $finish;
    end
end

wire [ASIZE-1:0] A0_PSE;
wire [ASIZE-1:0] A1_PSE;
wire [BSIZE-1:0] B0_PSE;
wire [BSIZE-1:0] B1_PSE;
wire [BSIZE-1:0] C0_PSE;
wire [BSIZE-1:0] C1_PSE;

wire [PSIZE-1:0] P_OUT;
wire [PSIZE-1:0] P_ROUND;

reg  [ASIZE-1:0] a0_ireg, a1_ireg;
reg  [BSIZE-1:0] b0_ireg, b1_ireg;
reg  [BSIZE-1:0] c0_ireg, c1_ireg;
reg  asign_ireg, bsign_ireg, csign_ireg;
reg  addsub_ireg;
reg  [1:0] preaddsub_ireg;

wire [ASIZE-1:0] a0_in, a1_in;
wire [BSIZE-1:0] b0_in, b1_in;
wire [BSIZE-1:0] c0_in, c1_in;
wire asign_in, bsign_in, csign_in;
wire addsub_in;
wire [1:0] preaddsub_in;

wire [BSIZE:0] prad_b0, prad_c0, prad_sum0;
wire [BSIZE:0] prad_b1, prad_c1, prad_sum1;
wire prad_sign;
wire [BSIZE:0] b0_inmux;
wire [BSIZE:0] b1_inmux;
wire bsign_inmux;

reg  [ASIZE-1:0] a1_pareg, a0_pareg;
reg  [BSIZE:0]   b1_pareg, b0_pareg;
reg  asign_pareg, bsign_pareg;
wire [ASIZE-1:0] mult_a1, mult_a0;
wire [BSIZE:0]   mult_b1, mult_b0;
wire mult_asign, mult_bsign;

wire [PSIZE-1:0] mult_a1ext, mult_a0ext;
wire [PSIZE-1:0] mult_b1ext, mult_b0ext;
wire [PSIZE-1:0] PRODUCT_0;
wire [PSIZE-1:0] PRODUCT_1;
reg  [PSIZE-1:0] P2_reg_PRODUCT_0;
reg  [PSIZE-1:0] P2_reg_PRODUCT_1;
reg  P2_reg_ADDSUB;
wire P2_reg_ADDSUB_comb;

wire [PSIZE-1:0] P2_reg_PRODUCT_0_comb;
wire [PSIZE-1:0] P2_reg_PRODUCT_1_comb;
wire [PSIZE-1:0] sum;
reg  [PSIZE-1:0] P_reg;
wire [BSIZE-1:0]  b1_mux;
wire [BSIZE-1:0]  c0_mux;
wire [BSIZE-1:0]  c1_mux;
wire        csign_mux;
wire global_rstn, RST_sync, RST_async, rst_asyncomb;

assign global_rstn = GRS_EN == "TRUE" ? GRS_INST.GRSNET : 1'b1;
assign RST_sync = (SYNC_RST == "TRUE") ? RST : 1'b0;
assign RST_async = (SYNC_RST == "FALSE") ? RST : 1'b0;
assign rst_asyncomb = RST_async | (~global_rstn);

assign b1_mux = (SIB1_EN == "TRUE") ?  b0_in :  B1_PSE;
assign c0_mux = (SIC0_EN == "TRUE") ?  b0_in :  C0_PSE;
assign c1_mux = (SIC1_EN == "TRUE") ?  c0_in :  C1_PSE; // FIXME
assign csign_mux = (SIC0_EN == "TRUE") ?  bsign_in : C_SIGNED ;

INT_PSE #(.ASIZE(ASIZE),.SC_PSE(SC_PSE_A0)) U1_PSE( .A(A0), .SIGN(A_SIGNED), .A_PSE(A0_PSE) );
INT_PSE #(.ASIZE(ASIZE),.SC_PSE(SC_PSE_A1)) U2_PSE( .A(A1), .SIGN(A_SIGNED), .A_PSE(A1_PSE) );
INT_PSE #(.ASIZE(BSIZE),.SC_PSE(SC_PSE_B0)) U3_PSE( .A(B0), .SIGN(B_SIGNED), .A_PSE(B0_PSE) );
INT_PSE #(.ASIZE(BSIZE),.SC_PSE(SC_PSE_B1)) U4_PSE( .A(B1), .SIGN(B_SIGNED), .A_PSE(B1_PSE) );
INT_PSE #(.ASIZE(BSIZE),.SC_PSE(SC_PSE_C0)) U5_PSE( .A(C0), .SIGN(C_SIGNED), .A_PSE(C0_PSE) );
INT_PSE #(.ASIZE(BSIZE),.SC_PSE(SC_PSE_C1)) U6_PSE( .A(C1), .SIGN(C_SIGNED), .A_PSE(C1_PSE) );

initial begin
    {asign_ireg, a1_ireg, a0_ireg} = 'b0;
    {bsign_ireg, b1_ireg, b0_ireg} = 'b0;
    {csign_ireg, c1_ireg, c0_ireg} = 'b0;
     addsub_ireg = 0;
     preaddsub_ireg = 0;
     P2_reg_PRODUCT_0 = 0;
     P2_reg_PRODUCT_1 = 0;
     P2_reg_ADDSUB   = 0;
     P_reg    = 0;
end

always @(posedge CLK or posedge rst_asyncomb)
    if (rst_asyncomb || RST_sync) begin
        {asign_ireg, a1_ireg, a0_ireg} <= 'b0;
        {bsign_ireg, b1_ireg, b0_ireg} <= 'b0;
        {csign_ireg, c1_ireg, c0_ireg} <= 'b0;
         addsub_ireg    <= 0;
         preaddsub_ireg <= 0;
    end
    else if (CE) begin
        {asign_ireg, a1_ireg, a0_ireg} <= {A_SIGNED, A1_PSE, A0_PSE};
        {bsign_ireg, b1_ireg, b0_ireg} <= {B_SIGNED, b1_mux, B0_PSE};
        {csign_ireg, c1_ireg, c0_ireg} <= {csign_mux, c1_mux, c0_mux};
         addsub_ireg    <= (DYN_OP_ADDSUB == 1'b1)? ADDSUB : ADDSUB_OP;
         preaddsub_ireg <=  PREADDSUB;
    end

assign {asign_in, a1_in, a0_in} = (INREG_EN == "TRUE") ? {asign_ireg, a1_ireg, a0_ireg} : {A_SIGNED, A1_PSE, A0_PSE};
assign {bsign_in, b1_in, b0_in} = (INREG_EN == "TRUE") ? {bsign_ireg, b1_ireg, b0_ireg} : {B_SIGNED, b1_mux, B0_PSE};
assign {csign_in, c1_in, c0_in} = (INREG_EN == "TRUE") ? {csign_ireg, c1_ireg, c0_ireg} : {csign_mux, c1_mux, c0_mux};
assign preaddsub_in = (INREG_EN == "TRUE") ? preaddsub_ireg : PREADDSUB;
assign addsub_in    = (INREG_EN == "TRUE") ? addsub_ireg : (DYN_OP_ADDSUB == 1'b1)? ADDSUB : ADDSUB_OP;

always @(*) begin
    if (PREADD_EN && (BSIZE == 26) && (prad_sign == 1'b0))
        if ((preaddsub_in[0] == 1'b1 && prad_sum0[BSIZE] == 1'b1) ||
            (preaddsub_in[1] == 1'b1 && prad_sum1[BSIZE] == 1'b1) ) begin
            $display("PG30-ERROR: Unexpected function mismatch.");
        end
end

assign prad_b0 = {(bsign_in & b0_in[BSIZE-1]), b0_in};
assign prad_c0 = {(csign_in & c0_in[BSIZE-1]), c0_in};
assign prad_b1 = {(bsign_in & b1_in[BSIZE-1]), b1_in};
assign prad_c1 = {(csign_in & c1_in[BSIZE-1]), c1_in};
assign prad_sum0 = preaddsub_in[0] ? (prad_b0 - prad_c0) : (prad_b0 + prad_c0);
assign prad_sum1 = preaddsub_in[1] ? (prad_b1 - prad_c1) : (prad_b1 + prad_c1);
assign prad_sign = bsign_in | csign_in;

reg preadd_over_flag0;
always @(*)begin
  if(preaddsub_in[0]==1'b0 &&  PREADD_EN==1)begin
    if((bsign_in==1'b1 && b0_in[BSIZE-1]==1'b0 && csign_in==1'b0 && prad_sum0[BSIZE]==1'b1) || (bsign_in==1'b0 && csign_in==1'b1 && c0_in[BSIZE-1]==1'b0 && prad_sum0[BSIZE]==1'b1))begin
      preadd_over_flag0 = 1'b1;
    end
    else begin
      preadd_over_flag0 = 1'b0;
    end
  end
  else if(preaddsub_in[0]==1'b1 && PREADD_EN==1)begin
    if((bsign_in==1'b1 && b0_in[BSIZE-1]==1'b1 && csign_in==1'b0 && prad_sum0[BSIZE]==1'b0) || (bsign_in==1'b0 && csign_in==1'b1 && c0_in[BSIZE-1]==1'b1 && prad_sum0[BSIZE]==1'b1) ||
      (bsign_in ==1'b0 && csign_in==1'b0 && (b0_in<c0_in)))begin
      preadd_over_flag0 = 1'b1;
    end
    else begin
      preadd_over_flag0 = 1'b0;
    end
  end
end

reg preadd_over_flag1;
always @(*)begin
  if(preaddsub_in[1]==1'b0 && PREADD_EN==1)begin
    if((bsign_in==1'b1 && b1_in[BSIZE-1]==1'b0 && csign_in==1'b0 && prad_sum1[BSIZE]==1'b1) || (bsign_in==1'b0 && csign_in==1'b1 && c1_in[BSIZE-1]==1'b0 && prad_sum1[BSIZE]==1'b1))begin
      preadd_over_flag1 = 1'b1;
    end
    else begin
      preadd_over_flag1 = 1'b0;
    end
  end
  else if(preaddsub_in[1]==1'b1 && PREADD_EN==1)begin
    if((bsign_in==1'b1 && b1_in[BSIZE-1]==1'b1 && csign_in==1'b0 && prad_sum1[BSIZE]==1'b0) || (bsign_in==1'b0 && csign_in==1'b1 && c1_in[BSIZE-1]==1'b1 && prad_sum1[BSIZE]==1'b1) ||
      (bsign_in ==1'b0 && csign_in==1'b0 && (b1_in<c1_in)))begin
      preadd_over_flag1 = 1'b1;
    end
    else begin
      preadd_over_flag1 = 1'b0;
    end
  end
end

always @(preadd_over_flag0 or preadd_over_flag1) begin
    if ((preadd_over_flag0==1 || preadd_over_flag1==1) && PREADD_EN==1)
    $display("Error: PREADD result is overflow!");
end

assign b0_inmux    = PREADD_EN ? prad_sum0 : {1'b0, b0_in};
assign b1_inmux    = PREADD_EN ? prad_sum1 : {1'b0, b1_in};
assign bsign_inmux = PREADD_EN ? prad_sign : bsign_in;
always @(posedge CLK or posedge rst_asyncomb)
    if (rst_asyncomb || RST_sync) begin
        {asign_pareg, a1_pareg, a0_pareg} <= 'b0;
        {bsign_pareg, b1_pareg, b0_pareg} <= 'b0;
    end
    else if (CE) begin
        {asign_pareg, a1_pareg, a0_pareg} <= {asign_in, a1_in, a0_in};
        {bsign_pareg, b1_pareg, b0_pareg} <= {bsign_inmux, b1_inmux, b0_inmux};
    end

assign {mult_asign, mult_a1, mult_a0} = (PREREG_EN == "TRUE") ? {asign_pareg, a1_pareg, a0_pareg} : {asign_in, a1_in, a0_in};
assign {mult_bsign, mult_b1, mult_b0} = (PREREG_EN == "TRUE") ? {bsign_pareg, b1_pareg, b0_pareg} : {bsign_inmux, b1_inmux, b0_inmux};

assign mult_a0ext = {{(PSIZE-ASIZE){mult_asign & mult_a0[ASIZE-1]}}, mult_a0};
assign mult_a1ext = {{(PSIZE-ASIZE){mult_asign & mult_a1[ASIZE-1]}}, mult_a1};
assign mult_b0ext = {{(PSIZE-BSIZE-PREADD_EN){mult_bsign & mult_b0[BSIZE+PREADD_EN-1]}}, mult_b0[BSIZE+PREADD_EN-1:0]};
assign mult_b1ext = {{(PSIZE-BSIZE-PREADD_EN){mult_bsign & mult_b1[BSIZE+PREADD_EN-1]}}, mult_b1[BSIZE+PREADD_EN-1:0]};

assign PRODUCT_0 = mult_a0ext * mult_b0ext;
assign PRODUCT_1 = mult_a1ext * mult_b1ext;

always @(posedge CLK or posedge rst_asyncomb)
    if (rst_asyncomb || RST_sync) begin
        P2_reg_PRODUCT_0 <= 0;
        P2_reg_PRODUCT_1 <= 0;
        P2_reg_ADDSUB    <= 0;
    end
    else if (CE) begin
        P2_reg_PRODUCT_0 <= PRODUCT_0;
        P2_reg_PRODUCT_1 <= PRODUCT_1;
        P2_reg_ADDSUB    <= addsub_in;
    end
assign P2_reg_PRODUCT_0_comb = (PIPEREG_EN == "TRUE") ? P2_reg_PRODUCT_0 : PRODUCT_0;
assign P2_reg_PRODUCT_1_comb = (PIPEREG_EN == "TRUE") ? P2_reg_PRODUCT_1 : PRODUCT_1;
assign P2_reg_ADDSUB_comb    = (PIPEREG_EN == "TRUE") ? P2_reg_ADDSUB : addsub_in;

assign sum = (P2_reg_ADDSUB_comb == 0) ? (P2_reg_PRODUCT_0_comb + P2_reg_PRODUCT_1_comb) : 
                                   (P2_reg_PRODUCT_0_comb - P2_reg_PRODUCT_1_comb);

always @(posedge CLK or posedge rst_asyncomb)
    if (rst_asyncomb || RST_sync) begin
        P_reg <= 0;
    end
    else if (CE) begin
        P_reg <= sum;             
    end
assign P_OUT = (OUTREG_EN == "TRUE") ? P_reg : sum;

assign P = P_OUT;

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_DFF.v
//
// Functional description: D-type flip-flop
//
// Parameter description:
//      INIT: init value
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_DFF
#(
    parameter GRS_EN = "TRUE",
    parameter INIT = 1'b0
) (
    output reg Q,
    input wire D,
    input wire CLK
);

    wire grs_n;
    wire RS;

    tri1 grsnet = GRS_INST.GRSNET;

    assign grs_n=(GRS_EN=="TRUE")?grsnet:1'b1;

    not (RS, grs_n);

    initial Q = 1'bx;

    always @(posedge CLK or posedge RS) begin
        if (RS)
            Q <= 1'b0;
        else
            Q <= D;
    end

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_CLKBUFGMUX.v
//
// Functional description: Global Clock Mux Buffer
//
// Parameter description:
//      xxxx
//
// Port description:
//
// Revision:
//    06/18/14 - Initial version.
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_CLKBUFGMUX
#(
    parameter TRIGGER_MODE = "NORMAL",  // "NORMAL", "NEGEDGE", "POSEDGE"
    parameter SIM_DEVICE = "TITAN" //
)(
    output reg CLKOUT,
    input CLKIN0,
    input CLKIN1,
    input SEL
);

    reg  NEG_O, POS_O, NORMAL_O;    
    reg SEL_NEG1, SEL_NEG2, SEL_POS1, SEL_POS2;
    reg SEL_NEG1_D, SEL_NEG2_D, SEL_POS1_D, SEL_POS2_D;
    reg init;
    reg SWITCH;

    initial 
    begin
       CLKOUT = 1'b0;
       SEL_NEG1 = SEL;//1'b0;
       SEL_NEG2 = SEL;//1'b0;
       SEL_POS1 = SEL;//1'b0;     
       SEL_POS2 = SEL;//1'b0;
       SEL_NEG1_D = SEL;//1'b0;
       SEL_NEG2_D = SEL;//1'b0;
       SEL_POS1_D = SEL;//1'b0;     
       SEL_POS2_D = SEL;//1'b0;
       init = 1;
        #0.1;
       SEL_NEG1 = SEL;//1'b0;
       SEL_NEG2 = SEL;//1'b0;
       SEL_POS1 = SEL;//1'b0;     
       SEL_POS2 = SEL;//1'b0;
       SEL_NEG1_D = SEL;//1'b0;
       SEL_NEG2_D = SEL;//1'b0;
       SEL_POS1_D = SEL;//1'b0;     
       SEL_POS2_D = SEL;//1'b0;
       init = 0;

    end
    
    initial begin
       if ((TRIGGER_MODE == "NORMAL") || (TRIGGER_MODE == "NEGEDGE") || (TRIGGER_MODE == "POSEDGE")) begin
       end
       else
          $display ("GTP_CLKBUFGMUX error : illegal setting for TRIGGER_MODE");

       case (SIM_DEVICE)
            "TITAN": SWITCH = 0;
            "LOGOS","COMPACT","LOGOS2": SWITCH = 1;         
            default: begin
                $display("ERROR: GTP_CLKBUFGMUX instance %m parameter SIM_DEVICE value: %s is illegal. The legal values are TITAN or LOGOS or COMPACT or LOGOS2.", SIM_DEVICE);
                $finish;
            end
       endcase


    end



  
    always@ (negedge CLKIN0)
    begin
        if (SEL == 1'b1) begin
            SEL_NEG1 <= SEL;
            if(SWITCH)
                SEL_NEG1_D <= SEL_NEG1;
        end
    end
    
    always@ (negedge CLKIN1)
    begin
        if (SEL_NEG1 == 1'b1) begin
            if(!SWITCH)
                SEL_NEG2 <= SEL_NEG1;    
            else begin
                SEL_NEG2 <= SEL_NEG1_D;
                SEL_NEG2_D <= SEL_NEG2;
            end
        end
    end
  
    always@ (negedge CLKIN1)
    begin
        if (SEL == 1'b0) begin
            SEL_NEG1 <= SEL;
            if(SWITCH)
                SEL_NEG1_D <= SEL_NEG1;
        end
    end
  
    always@ (negedge CLKIN0)
    begin
        if (SEL_NEG1 == 1'b0) begin
            if(!SWITCH)
                SEL_NEG2 <= SEL_NEG1;
            else begin
                SEL_NEG2 <= SEL_NEG1_D;
                SEL_NEG2_D <= SEL_NEG2;
            end
        end
    end
    
    always@(*) begin
        if(SWITCH) begin
            if({SEL_NEG1_D, SEL_NEG2_D} == 2'b00)
                NEG_O = CLKIN0;
            else if({SEL_NEG1_D, SEL_NEG2_D} == 2'b11)
                NEG_O = CLKIN1;
            else
                NEG_O = 1'b0; 
        end
        else begin
            if ({SEL_NEG1, SEL_NEG2} == 2'b00)
                NEG_O = CLKIN0;
            else if({SEL_NEG1, SEL_NEG2} == 2'b11)
                NEG_O = CLKIN1;
            else 
                NEG_O = 1'b0;
        end
    end
  
    always@ (posedge CLKIN0)
    begin
        if (SEL == 1'b1) begin
            SEL_POS1 <= SEL;
            if(SWITCH)
                SEL_POS1_D <= SEL_POS1;
        end
    end
    
    always@ (posedge CLKIN1)
    begin
        if (SEL == 1'b1) begin
            if(!SWITCH)
                SEL_POS2 <= SEL_POS1;
            else begin
                SEL_POS2 <= SEL_POS1_D;
                SEL_POS2_D <= SEL_POS2;
            end
        end
    end
  
    always@ (posedge CLKIN1)
    begin
        if (SEL == 1'b0) begin
            SEL_POS1 <= SEL;
            if(SWITCH)
                SEL_POS1_D <= SEL_POS1;
        end
    end
  
    always@ (posedge CLKIN0)
    begin
        if (SEL == 1'b0) begin
            if(!SWITCH)
                SEL_POS2 <= SEL_POS1;
            else begin
                SEL_POS2 <= SEL_POS1_D;
                SEL_POS2_D <= SEL_POS2;
            end
        end
    end
    
    always@(*) begin
        if(SWITCH) begin
            if({SEL_POS1_D, SEL_POS2_D} == 2'b00)
                POS_O = CLKIN0;
            else if({SEL_POS1_D, SEL_POS2_D} == 2'b11)
                POS_O = CLKIN1;
            else 
                POS_O = 1'b1;
        end
        else begin
            if ({SEL_POS1, SEL_POS2} == 2'b00)
                POS_O = CLKIN0;
            else if({SEL_POS1, SEL_POS2} == 2'b11)
                POS_O = CLKIN1;
            else 
                POS_O = 1'b1;
        end
    end

    always@(*)
    begin
        if (SEL == 1'b0)
            NORMAL_O = CLKIN0;
        else
            NORMAL_O = CLKIN1;
    end
  
    always @ (*)
    begin
        if(!init) begin
            if (TRIGGER_MODE == "NORMAL")
                CLKOUT = NORMAL_O;
            else if (TRIGGER_MODE == "NEGEDGE")
                CLKOUT = NEG_O;
            else if (TRIGGER_MODE == "POSEDGE")
                CLKOUT = POS_O;
        end
    end   

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library:
// Filename: GTP_IOCLKDIV_E1.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_IOCLKDIV_E1 #(
parameter DIV_FACTOR = "DIV_DIS", //"DIV_DIS";"2"; "3.5"; "4"; 
parameter GRS_EN = "TRUE" //"TRUE"; "FALSE"
)(
output CLKDIVOUT,
output CLKOUT,
input CLKIN,
input RST_N,
input ALIGNWD
);                        // synthesis syn_black_box

//synthesis translate_off
assign global_rstn = ((GRS_EN == "TRUE" )? GRS_INST.GRSNET : 1'b1);

initial 
begin
if ((DIV_FACTOR == "2") || (DIV_FACTOR == "3.5") ||  (DIV_FACTOR == "4") || (DIV_FACTOR == "DIV_DIS")) begin
end
else
   $display (" GTP_IOCLKDIV_E1 error: illegal setting for DIV_FACTOR");
end




reg [1:0] ctl_div;



initial
begin
    casex(DIV_FACTOR)
    "DIV_DIS":ctl_div=2'b00;
    "2"      :ctl_div=2'b01;
    "3.5"    :ctl_div=2'b10;
    "4"      :ctl_div=2'b11;
     default:ctl_div=2'b00;
    endcase
end

wire rst_div;

assign rst_div = !((!RST_N)|(!global_rstn));


  reg [2:0] counter_h;
  reg [2:0] counter_l;
  reg temp1;
  reg temp2;
  reg rst_n;
  wire temp3;
  wire divmode_cut ;
  assign divmode_cut = ((DIV_FACTOR =="2")? 1'b1:1'b0)|((DIV_FACTOR =="3.5")? 1'b1:1'b0)|((DIV_FACTOR =="4")? 1'b1:1'b0);
  assign CLKDIVOUT = (divmode_cut==1'b1) ? (temp1|temp2):temp3;

assign temp3 = (rst_n == 1'b0) ? 1'b0 : 1'b1;




wire temp7;
  assign temp7 = (ctl_div==2'b00)?1'b1:CLKIN;

assign CLKOUT = (rst_n & temp7);



  
//  assign CLKDIVOUT = temp1|temp2;
 
  always @( negedge CLKIN or negedge rst_div )  
           begin
              if (rst_div == 1'b1)   //rst_loc_n =1,work;rst_loc_n=0,rst
                rst_n <= 1'b1;
              else
                rst_n <= 1'b0;
           end


reg out_reg0_0;

  always @( posedge CLKIN or negedge rst_n )
           begin
              if (rst_n == 1'b0)
                out_reg0_0 <= 1'b0;
              else begin
                     if(ALIGNWD==1'b1)
                         out_reg0_0 <=1'b1;
                      else out_reg0_0 <=1'b0;
                    end
           end


reg out_reg0_0_bak;

  always @( posedge CLKIN or negedge rst_n )
           begin
              if (rst_n == 1'b0)
                out_reg0_0_bak <= 1'b0;
              else begin
                     if(out_reg0_0==1'b1)
                         out_reg0_0_bak <=1'b1;
                      else out_reg0_0_bak <=1'b0;
                    end
           end




reg out_reg0;

  always @( posedge CLKIN or negedge rst_n )  
           begin
              if (rst_n == 1'b0) 
                out_reg0 <= 1'b0;
              else begin
                     if(out_reg0_0_bak==1'b1)
                         out_reg0 <=1'b1;
                      else out_reg0 <=1'b0;
                    end
           end



reg out_reg1;

  always @( posedge CLKIN or negedge rst_n )  
           begin
              if (rst_n == 1'b0) 
                out_reg1 <= 1'b0;
              else begin
                     if(out_reg0==1'b1)
                         out_reg1 <=1'b1;
                      else out_reg1 <=1'b0;
                    end
           end


reg out_reg2;


  always @( negedge CLKIN or negedge rst_n )  
           begin
              if (rst_n == 1'b0) 
                out_reg2 <= 1'b0;
              else begin
                     if(out_reg1==1'b1)
                         out_reg2 <=1'b1;
                      else out_reg2<=1'b0;
                    end
           end



reg out_reg3;

  always @( negedge CLKIN or negedge rst_n )  
           begin
              if (rst_n == 1'b0) 
                out_reg3 <= 1'b0;
              else begin
                     if(out_reg0==1'b1)
                         out_reg3 <=1'b1;
                      else out_reg3<=1'b0;
                    end
           end

wire ALIGNWD_TMP;

assign out_reg2_n = ~out_reg2;

assign ALIGNWD_TMP=~(out_reg2_n&out_reg3);



reg ALIGN0;
wire ALIGN0_N;
wire ALIGNWD_TMP_N ;
assign ALIGNWD_TMP_N=~ALIGNWD_TMP;
assign ALIGN0_N=~ALIGN0;

  always @( posedge ALIGNWD_TMP_N or negedge rst_n )  
           begin
              if (rst_n == 1'b0) 
                ALIGN0 <= 1'b0;
              else begin
                     if(ALIGN0_N==1'b1)
                         ALIGN0 <=1'b1;
                      else ALIGN0<=1'b0;
                    end
           end


reg out_reg4;
assign out_reg4_n=~out_reg4;
  always @( posedge ALIGNWD_TMP or negedge rst_n )  
           begin
              if (rst_n == 1'b0) 
                out_reg4 <= 1'b0;
              else begin
                     if(out_reg4_n==1'b1)
                         out_reg4 <=1'b1;
                      else out_reg4<=1'b0;
                    end
           end


wire BLOCK1;
assign BLOCK1= ~(ALIGN0_N&out_reg4);










wire ali_ctl_b;
wire clk_in_b;


assign ali_ctl_b = ((ctl_div==2'b01)? 1'b1:1'b0)| ((ctl_div==2'b11)? 1'b1:1'b0) ;

assign clk_in_b = ((ali_ctl_b==1'b1)? BLOCK1:ALIGNWD_TMP)&CLKIN&rst_n;

  always @(posedge clk_in_b or negedge rst_n)                //counter created
    if(~rst_n) begin
      counter_h <= 3'b000;
      temp1 <= 0;
    end else 
      case(DIV_FACTOR)
        "2":                                            //create DIV2 counter
          temp1 <= ~temp1;
        "3.5":                                           //create DIV35 counter
          if(counter_h == 3'b110)
            counter_h <= 3'b000;
          else begin
            temp1 <= ~(counter_h[2]|counter_h[1]);
            counter_h <= counter_h+1;
          end 
        "4":                                           //create DIV4 counter
          if(counter_h == 3'b011)
            counter_h <= 3'b000;
          else begin
            temp1 <= ~counter_h[1];
            counter_h <= counter_h+1;  
          end                               
      endcase
      
  always @(negedge clk_in_b or negedge rst_n)
    if(~rst_n) begin
      counter_l <= 3'b000;
      temp2 <= 0;
    end else 
      case(DIV_FACTOR)
        "3.5":                                        //create DIV35 clock
              temp2 <= counter_h[2]&(~counter_h[1]);
      endcase         







//synthesis translate_on


endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_RBCRC.v
//
// Functional description: RBCRC Circuit
//
// Parameter description:
//      
//
// Port description:
//      
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 10 fs
module GTP_RBCRC
(
input         RST,
input         START,
input         SEC_START,
output        ERR,
output        VALID,
output        SEC_OVER
);

wire            init_complete;
wire            done;

wire    [1:0]   cmem_type;
wire            erase_en;
wire            wl_on;
wire            wlsrce;

wire            prog_on;
wire            prog_cap;
wire    [4:0]   region_sel;
wire            region_rw_en;
wire   [31:0]   blsrin;

wire            prechge;
wire            read;
wire            rdbk_cap;
wire            clk_cram;
wire            clk_drm;
wire    [7:0]   frame_addr;
wire            ndrm_column_inc;
wire    [7:0]   column;
wire            ndrm_region_inc;
wire            ndrm_region_end;
wire            mce;
wire            mwr;
wire   [31:0]   databack;

reg  clk;
wire rbcrc_clk;
reg  rstn;

reg  clk_532_reg;
reg  [6:0] cnt_sed_reg;
reg  clk_sed_reg;
wire [6:0] clk_sed_div;
wire [31:0] optionr0;

always #24.438 clk = ~clk;
always #0.94 clk_532_reg = ~clk_532_reg;

initial 
    begin
        clk = 1'b0;
        rstn = 1'b0;
        clk_532_reg = 1'b0;
        #10;
        rstn = 1'b1;
    end



INT_RBCRC_CCS  INT_RBCRC_CCS (

.idcode               (32'h0),

.por_n                (rstn),
.rst_n                (rstn),

.init_n               (init_complete),
.init_complete        (init_complete),

.done_i               (done),
.done                 (done),

.fpclk                (1'b1),
.dout                 (32'd0),

.clk_cram             (clk_cram),
.clk_drm              (clk_drm),
.cmem_type            (cmem_type),
.erase_en             (erase_en     ),
.wl_on                (wl_on        ),

.frame_addr           (frame_addr),
.ndrm_column_inc      (ndrm_column_inc),
.column               (column),

.prog_on              (prog_on      ),
.prog_cap             (prog_cap     ),
.ndrm_region_end      (ndrm_region_end),

.region_rw_en         (region_rw_en ),
.blsrin               (blsrin       ),
                                    
.databack             (databack),
.prechge              (prechge      ),
.read                 (read         ),
.rdbk_cap             (rdbk_cap     ),
.mce                  (mce),
.mwr                  (mwr),

.glogen_fb            (glogen),
.glogen               (glogen),

.clk                  (clk),

.pctlr_clk            (1'b1),

.pclk                 (1'b1),
.presetn              (1'b1),
.paddr                (5'h1F),
.psel_ccs             (1'b1),
.psel_spi             (1'b1),
.psel_i2c0            (1'b1),
.psel_i2c1            (1'b1),
.psel_timer           (1'b1),
.psel_pll0            (1'b1),
.psel_pll1            (1'b1),
.penable              (1'b1),
.pwrite               (1'b1),
.pwdata               (8'hFF),
.prdata               (),
.pready               (),

.pll0_prdata          (8'hFF),
.pll0_pready          (1'b1),

.pll1_prdata          (8'h0),
.pll1_pready          (1'b0),

.rbcrc_clk            (rbcrc_clk),
.rbcrc_rst            (RST),
.rbcrc_start          (START),
.rbcrc_err            (ERR),
.rbcrc_valid          (VALID),

.spi_ss_i_n           (1'b1),
.spi_ss_o_n           (),
.spi_sck_oe_n         (),
.spi_sck_i            (1'b1),
.spi_sck_o            (),
.spi_mosi_oe_n        (),
.spi_mosi_i           (1'b1),
.spi_mosi_o           (),
.spi_miso_oe_n        (),
.spi_miso_i           (1'b1),
.spi_miso_o           (),
.irq_spi              (),

.i2c0_scl_i           (1'b1),
.i2c0_scl_o           (),
.i2c0_sda_i           (1'b1),
.i2c0_sda_o           (),
.irq_i2c0             (),

.i2c1_scl_i           (1'b1),
.i2c1_scl_o           (),
.i2c1_sda_i           (1'b1),
.i2c1_sda_o           (),
.irq_i2c1             (),

.timer_rstn           (1'b1),
.timer_clk            (1'b1),
.timer_stamp          (1'b1),
.timer_pwm            (),
.irq_timer            ()

);

assign clk_sed_div = optionr0[30:24];

INT_RBCRC_CRAM  INT_RBCRC_CRAM (
.cmem_type          (cmem_type[0]),
.wl_on              (wl_on),
.clk_cram           (clk_cram),
.clk_drm            (clk_drm),
.read               (read),
.rdbk_cap           (rdbk_cap),
.erase_en           (erase_en),
.prog_cap           (prog_cap),
.prog_on            (prog_on),
.blsrin             (blsrin),
.frame_addr         (frame_addr),
.prechg             (prechge),
.ndrm_column_inc    (ndrm_column_inc),
.column             (column),
.ndrm_region_end    (ndrm_region_end),
.region_rw_en       (region_rw_en),
.por_n              (rstn),
.mce                (mce),
.mwr                (mwr),
.databack           (databack),
.optionr0           (optionr0)

);

always @(posedge clk_532_reg or negedge rstn)
begin
    if (!rstn)
    begin
        cnt_sed_reg <= 7'b000_0000;
        clk_sed_reg <= 1'b0;
    end
    else 
        if(cnt_sed_reg == clk_sed_div - 7'b1)
        begin
            cnt_sed_reg <= 7'b000000;
            clk_sed_reg <= ~clk_sed_reg;
        end
        else
        begin
            cnt_sed_reg <= cnt_sed_reg + 1'b1;
            clk_sed_reg <= clk_sed_reg;
    end
end

assign rbcrc_clk = clk_sed_reg;


endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_MULTACC36.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

//P = MAC + A*B
module GTP_MULTACC36 #(
    parameter GRS_EN              = "TRUE", //"TRUE"; "FALSE"
    parameter SYNC_RST            = "FALSE", //"TRUE"; "FALSE"
    parameter INREG_EN            = "FALSE",  //"TRUE"; "FALSE"
    parameter PIPEREG_EN          = "FALSE",   //"TRUE"; "FALSE"
    parameter ACC_ADDSUB_OP       = 0,
    parameter DYN_ACC_ADDSUB_OP   = 1,     //Select parameter ADDSUB or input ADDSUB
    parameter OVERFLOW_MASK       = 64'h0, //PSIZE = 64 OVERflow setting =  'h8000_0000_0000_00XX , bit width = PSIZE
    parameter PATTERN             = 64'h0, //compare pattern
    parameter MASKPAT             = 64'h0, //pattern mask
    parameter DYN_ACC_INIT        = 0,  //acc init value dynamic input
    parameter ACC_INIT_VALUE      = 64'h0  //acc init value parameter
) (
    output  [63:0] P,
    output  OVER,
    output  UNDER,
    output  EQZ,
    output  EQZM,
    output  EQOM,
    output  EQPAT,
    output  EQPATN,

    input   CE,
    input   RST,
    input   CLK,
    input   [35:0] A,
    input   [17:0] B,
    input   A_SIGNED,
    input   B_SIGNED,
    input   [63:0] ACC_INIT,
    input   ACC_ADDSUB,
    input   RELOAD
);

    wire [63:0] R;

    INT_PREADD_MULTACC #(
        . GRS_EN(GRS_EN),     
        . SYNC_RST(SYNC_RST),   
        . INREG_EN(INREG_EN),   
        . PIPEREG_EN(PIPEREG_EN), 
        . ACCUMADDSUB_OP(ACC_ADDSUB_OP), 
        . DYN_OP_SEL(DYN_ACC_ADDSUB_OP),     
        . ASIZE(36),    
        . BSIZE(18),    
        . PSIZE(64),    
        . PREADD_EN(0),
        . MASK(OVERFLOW_MASK),      
        . DYN_ACC_INIT(DYN_ACC_INIT),
        . ACC_INIT_VALUE(ACC_INIT_VALUE)
    ) U_MACC (
        .CE(CE),
        .RST(RST),
        .CLK(CLK),
        .A(A),
        .B(B),
        .A_SIGNED(A_SIGNED),
        .B_SIGNED(B_SIGNED),
        .C_SIGNED(B_SIGNED),
        .C(18'b0),
        .PREADDSUB(1'b0),
        .ACCUM_INIT(ACC_INIT),
        .ACCUMADDSUB(ACC_ADDSUB),
        .RELOAD(RELOAD),
        .P(P),
        .OVER(OVER),
        .UNDER(UNDER),     
        .R(R)
    );

    INT_FLAG #(
        . GRS_EN(GRS_EN),
        . SYNC_RST(SYNC_RST),
        . PSIZE(64),
        . PATSIZE(64),
        . MASKPATSIZE(64),
        . OUTREG_EN("TRUE")
    ) U_FLAG (
        . CE(CE),
        . RST(RST),
        . CLK(CLK),
        . P(P),
        . PATTERN(PATTERN),
        . MASKPAT(MASKPAT),
        . OVERFLOW_MASK(OVERFLOW_MASK),
        . R(R),
        . eqz(EQZ),
        . eqzm(EQZM),
        . eqom(EQOM),
        . eqpat(EQPAT),
        . eqpatn(EQPATN)
    );

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_MULTADD36.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

//P = A0*B0 +/- A1*B1
module GTP_MULTADD36 #(
    parameter GRS_EN        = "TRUE", //"TRUE"; "FALSE"
    parameter SYNC_RST      = "FALSE", //"TRUE"; "FALSE"
    parameter INREG_EN      = "FALSE", //"TRUE"; "FALSE"
    parameter PIPEREG_EN    = "FALSE", //"TRUE"; "FALSE"
    parameter OUTREG_EN     = "FALSE", //"TRUE"; "FALSE"
    parameter ADDSUB_OP     = 0 ,
    parameter DYN_ADDSUB_OP = 1
)(
    output  [55-1:0] P,           //product
    input   CE,
    input   RST,
    input   CLK,
    input   A_SIGNED,
    input   [36-1:0] A0,
    input   [36-1:0] A1,
    input   B_SIGNED,
    input   [18-1:0] B0,
    input   [18-1:0] B1,
    input   ADDSUB
);

    INT_PREADD_MULTADD #(
        . GRS_EN(GRS_EN),
        . SYNC_RST(SYNC_RST),   
        . INREG_EN(INREG_EN),   
        . PIPEREG_EN(PIPEREG_EN), 
        . OUTREG_EN(OUTREG_EN),  
        . ADDSUB_OP(ADDSUB_OP),  
        . DYN_OP_ADDSUB(DYN_ADDSUB_OP), 
        . ASIZE(36), 
        . BSIZE(18),
        . PREADD_EN(0)
    ) U_MULTADD36 (
        . CE(CE),
        . RST(RST),
        . CLK(CLK),
        . A_SIGNED(A_SIGNED),
        . A0(A0),
        . A1(A1),
        . B_SIGNED(B_SIGNED),
        . B0(B0),
        . B1(B1),
        . C_SIGNED(B_SIGNED),
        . C0(18'b0),
        . C1(18'b0),
        . PREADDSUB(2'b0),
        . ADDSUB(ADDSUB),
        . P(P)
    );

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2016 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_CLKBUFMCE.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_CLKBUFMCE
#(
    parameter TRIGGER_MODE = "POSEDGE",
    parameter CE_TYPE = "SYNC",
    parameter CE_INV = "FALSE"

) (
    output CLKOUT,
    input CLKIN,
    input CE
);

//synthesis translate_off

    initial begin
        if(CE_TYPE != "SYNC" && CE_TYPE != "ASYNC") begin
            $display("ERROR: The attribute CE_TYPE on instance %m is %s. Legal value are SYNC or ASYNC.", CE_TYPE);
            $finish;
        end
        if(TRIGGER_MODE != "POSEDGE" && TRIGGER_MODE != "NEGEDGE") begin
            $display("ERROR: The attribute TRIGGER_MODE on instance %m is %s. Legal value are POSEDGE or NEGEDGE.", TRIGGER_MODE);
            $finish;
        end
        if(CE_INV != "TRUE" && CE_INV != "FALSE") begin
            $display("ERROR: The attribute CE_INV on instance %m is %s. Legal value are TRUE or FALSE.", CE_INV);
            $finish;
        end        
    end

    wire ce;
    wire outs;
    wire outps;
    wire outns;
    wire outa;
    wire outpa;
    wire outna;
    
    reg flag1;
    reg flag2;
    reg mid1;
    reg mid2;

    initial 
    begin
        flag1 = 0;
        flag2 = 0;
        mid1 = 0;
        mid2 = 0;
        #0.1 ;
        flag1 = 0;
        flag2 = 0;
        mid1 = 0;
        mid2 = 0;
    end

    assign ce = (CE_INV == "FALSE")? CE : !CE;
    assign CLKOUT = (CE_TYPE == "SYNC")? outs : outa;
    assign outs = (TRIGGER_MODE == "POSEDGE")? outps : outns;
    assign outps = flag1? CLKIN : 1'b1;
    assign outns = flag2? CLKIN : 1'b0;
    assign outa = (TRIGGER_MODE == "POSEDGE")? outpa : outna;
    assign outpa = ce? CLKIN : 1'b1;
    assign outna = ce? CLKIN : 1'b0;

    always@(posedge CLKIN) begin
        if(ce) begin
            flag1 <= mid1;
            mid1 <= 1;
        end        
        else begin
            flag1 <= mid1;
            mid1 <= 0;
        end
    end

    always@(negedge CLKIN) begin
        if(ce) begin
            flag2 <= mid2;
            mid2 <= 1;
    
        end
        else begin
            flag2 <= mid2;
            mid2 <= 0;
        end        
    end


//synthesis translate_on

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2017 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_ADC_E1.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1ns/1ps

module GTP_ADC_E1 #(
     parameter AVERAGE      = "1",   ///  1/16/64/256
     parameter CALIB        = "NONE",///  NONE/OFFSET/OFFSET_GAIN
     parameter REFERENCE       = "INTERNAL", ///  INTERNAL/EXTERNAL
     parameter CALIB_REFERENCE = "INTERNAL", ///  INTERNAL/EXTERNAL
     parameter FULL_SWING   = "0.5V",///  0.5/0.6/0.7/0.8/0.9/1.0/1.1/1.2
     parameter VCM          = "0.8V",///  0.8/0.9/1.0/1.1/1.2/1.3/1.4/1.5
     parameter DIVIDER      = "2",   ///  2/3/4/5/6/7/8/9/10/11/12/13/14/15/16

     parameter ADC_MODE       = "DEFAULT",///  DEFAULT/SINGLE_PASS/CONTINUE_SEQ/SINGLE_CHANNEL
     parameter EVENT_DRIVE    = "FALSE",///  FALSE/TRUE
     parameter ADC_MODE_1MSPS = "FALSE",///  FALSE/TRUE
     parameter CLKSWITCH      = "FALSE",///  FALSE/TRUE
     parameter INTERNAL_VOL_SEL = "VDD33",  ///  VDD33/VDD11/VDDM
     parameter SINGLE_CH_SEL    = "0", ///  0/1/2/3/4/5/6/7/8/9/10/11/12/13/14/15/
     parameter SINGLE_CH_IN     = "SINGLE_END",///  SINGLE_END/UNIPOLAR/BIPOLAR

     parameter SEQ_CH11_10_SEL  = "NONE",///  NONE/CH10/CH11/ALL
     parameter SEQ_CH9_8_SEL    = "NONE",///  NONE/CH8/CH9/ALL
     parameter SEQ_CH7_6_SEL    = "NONE",///  NONE/CH6/CH7/ALL
     parameter SEQ_CH5_4_SEL    = "NONE",///  NONE/CH4/CH5/ALL
     parameter SEQ_CH3_2_SEL    = "NONE",///  NONE/CH2/CH3/ALL
     parameter SEQ_CH1_0_SEL    = "NONE",///  NONE/CH0/CH1/ALL

     parameter SEQ_CH11_10_IN   = "SINGLE_END",///  SINGLE_END/UNIPOLAR/BIPOLAR
     parameter SEQ_CH9_8_IN     = "SINGLE_END",///  SINGLE_END/UNIPOLAR/BIPOLAR
     parameter SEQ_CH7_6_IN     = "SINGLE_END",///  SINGLE_END/UNIPOLAR/BIPOLAR
     parameter SEQ_CH5_4_IN     = "SINGLE_END",///  SINGLE_END/UNIPOLAR/BIPOLAR
     parameter SEQ_CH3_2_IN     = "SINGLE_END",///  SINGLE_END/UNIPOLAR/BIPOLAR
     parameter SEQ_CH1_0_IN     = "SINGLE_END",///  SINGLE_END/UNIPOLAR/BIPOLAR
    
     parameter integer TEMP_SENSOR_HIGH = 0,//0~255
     parameter integer TEMP_SENSOR_LOW  = 0,//0~255

     parameter ADC_EN_ENABLE = "FALSE" // FALSE/TRUE

     ) (
     input  [9:0]  VAUX,
     input  [1:0]  VA,
     input         RST_N,
     input         LOADSC_N,
     input         DCLK,
     input         DEN,
     input  [15:0] DI,
     input         DWE,
     input  [7:0]  DADDR,
     input         CONVST,

     input         ADC_EN,

     output        DBUSY,
     output [15:0] DO,
     output        DRDY,
     output        DMODIFIED,
     output        LOGIC_DONE,
     output        OVER_TEMP
     );

    // pragma translate_off
    /////signal begin/////
    wire           ad_done;
    wire  [11:0]   ad_dat;

    ////out
    wire           ad_clk;
    wire           ad_rstn;
    wire           ad_do_offset;
    wire           ad_do_gain;
    wire   [1:0]   ad_offset;
    wire           ad_mode_diff_en;
    wire   [1:0]   ad_mux;
    wire   [3:0]   ad_sela;
    wire   [3:0]   ad_selb;
    wire           ad_bias_pd;
    wire           ad_clk_en;
    wire   [2:0]   ad_fs_g;
    wire   [2:0]   ad_vcm_g;
    wire           ad_ref_sel;
    wire           ad_cref_sel;
    wire           over_temp_ccs;

    reg   [15:0]  sc_reg0   ;
    reg   [15:0]  sc_reg1   ;
    reg   [15:0]  sc_reg2   ;
    reg   [15:0]  sc_reg3   ;
    reg   [15:0]  sc_reg4   ;

    reg sc_ad_en_enable;
    /////signal end/////

    ///////////////////////////////////
    reg                TCK       ;
    reg                FLG_JDRP  ;
    reg                CLOCKDR   ;
    reg                CAPTUREDR ;
    reg                SHIFTDR   ;
    reg                UPDATEDR  ;
    reg                TDI       ;
    reg                GLOGEN    ;
    reg                CLK_OSC   ;
    reg                POR_N     ;
    reg                VDD33A    ;
    reg                VDD33     ;
    reg                VDD11     ;
    reg                VDDM      ;
    reg                VTEMP_P   ;
    reg                VTEMP_N   ;
    reg                VREF_EXT  ;
    reg                IBREF10U  ;
    reg                IB10U_IN  ;
    reg                VSSA      ;
    reg                VSS       ;

    wire               TDO;
    wire               ad_vref_test;
    ///////////////////////////////////

    initial
    begin
                sc_reg0      <= 16'b0000_0000_0000_0000;
                sc_reg1      <= 16'b0000_0000_0000_0000;
                sc_reg2      <= 16'b0000_0000_0000_0000;
                sc_reg3      <= 16'b0000_0000_0000_0000;
                sc_reg4      <= 16'b0000_0000_0000_0000;

                sc_ad_en_enable <= 1'b0;
              
                TCK          <= 0;
                FLG_JDRP     <= 0;
                CLOCKDR      <= 0;
                CAPTUREDR    <= 0;
                SHIFTDR      <= 0;
                UPDATEDR     <= 0;
                TDI          <= 0;
                GLOGEN       <= 0;
                CLK_OSC      <= 0;
                POR_N        <= 0;
                VDD33A       <= 1;
                VDD33        <= 1;
                VDD11        <= 1;
                VDDM         <= 1;
                VTEMP_P      <= 1;
                VTEMP_N      <= 1;
                VREF_EXT     <= 1;
                IBREF10U     <= 1;
                IB10U_IN     <= 1;
                VSSA         <= 0;
                VSS          <= 0;
                #500;
                POR_N        <= 1;
                #200000;
                GLOGEN       <= 1;
    end

    always #10 CLK_OSC = ~CLK_OSC & GLOGEN;

    //////parameter to sc signal//////
    always @(GLOGEN)
    begin
        if(GLOGEN)
            case(AVERAGE)
                "1"  : sc_reg0[15:14] = 2'b00;
                "16" : sc_reg0[15:14] = 2'b01;
                "64" : sc_reg0[15:14] = 2'b10;
                "256": sc_reg0[15:14] = 2'b11;
                default:
                begin
                    $display ("GTP_ADC_E1 error: illegal setting for AVERAGE");
                    $stop;
                end
            endcase
        else
            sc_reg0[15:14] = 2'b00;
    end

    always @(GLOGEN)
    begin
        if(GLOGEN)
            case(CALIB)
                "NONE"        : sc_reg0[13:12] = 2'b00;
                "OFFSET"      : sc_reg0[13:12] = 2'b01;
                "OFFSET_GAIN" : sc_reg0[13:12] = 2'b11;
                default:
                begin
                    $display ("GTP_ADC_E1 error: illegal setting for CALIB");
                    $stop;
                end
            endcase
        else
            sc_reg0[13:12] = 2'b00;
    end

    always @(GLOGEN)
    begin
        if(GLOGEN)
            case(REFERENCE)
                "INTERNAL" : sc_reg0[11] = 1'b0;
                "EXTERNAL" : sc_reg0[11] = 1'b1;
                default:
                begin
                    $display ("GTP_ADC_E1 error: illegal setting for REFERENCE");
                    $stop;
                end
            endcase
        else
            sc_reg0[11] = 1'b0;
    end

    always @(GLOGEN)
    begin
        if(GLOGEN)
            case(CALIB_REFERENCE)
                "INTERNAL" : sc_reg0[10] = 1'b0;
                "EXTERNAL" : sc_reg0[10] = 1'b1;
                default:
                begin
                    $display ("GTP_ADC_E1 error: illegal setting for CALIB_REFERENCE");
                    $stop;
                end
            endcase
        else
            sc_reg0[10] = 1'b0;
    end

    always @(GLOGEN)
    begin
        if(GLOGEN)
            case(FULL_SWING)
                "0.5V" : sc_reg0[9:7] = 3'b000;
                "0.6V" : sc_reg0[9:7] = 3'b001;
                "0.7V" : sc_reg0[9:7] = 3'b010;
                "0.8V" : sc_reg0[9:7] = 3'b011;
                "0.9V" : sc_reg0[9:7] = 3'b100;
                "1.0V" : sc_reg0[9:7] = 3'b101;
                "1.1V" : sc_reg0[9:7] = 3'b110;
                "1.2V" : sc_reg0[9:7] = 3'b111;
                default:
                begin
                    $display ("GTP_ADC_E1 error: illegal setting for FULL_SWING");
                    $stop;
                end
            endcase
        else
            sc_reg0[9:7] = 3'b000;
    end

    always @(GLOGEN)
    begin
        if(GLOGEN)
            case(VCM)
                "0.8V" : sc_reg0[6:4] = 3'b000;
                "0.9V" : sc_reg0[6:4] = 3'b001;
                "1.0V" : sc_reg0[6:4] = 3'b010;
                "1.1V" : sc_reg0[6:4] = 3'b011;
                "1.2V" : sc_reg0[6:4] = 3'b100;
                "1.3V" : sc_reg0[6:4] = 3'b101;
                "1.4V" : sc_reg0[6:4] = 3'b110;
                "1.5V" : sc_reg0[6:4] = 3'b111;
                default:
                begin
                    $display ("GTP_ADC_E1 error: illegal setting for VCM");
                    $stop;
                end
            endcase
        else
            sc_reg0[6:4] = 3'b000;
    end

    always @(GLOGEN)
    begin
        if(GLOGEN)
            case(DIVIDER)
                "2" : sc_reg0[3:0] = 4'b0001;
                "3" : sc_reg0[3:0] = 4'b0010;
                "4" : sc_reg0[3:0] = 4'b0011;
                "5" : sc_reg0[3:0] = 4'b0100;
                "6" : sc_reg0[3:0] = 4'b0101;
                "7" : sc_reg0[3:0] = 4'b0110;
                "8" : sc_reg0[3:0] = 4'b0111;
                "9" : sc_reg0[3:0] = 4'b1000;
                "10": sc_reg0[3:0] = 4'b1001;
                "11": sc_reg0[3:0] = 4'b1010;
                "12": sc_reg0[3:0] = 4'b1011;
                "13": sc_reg0[3:0] = 4'b1100;
                "14": sc_reg0[3:0] = 4'b1101;
                "15": sc_reg0[3:0] = 4'b1110;
                "16": sc_reg0[3:0] = 4'b1111;
                default:
                begin
                    $display ("GTP_ADC_E1 error: illegal setting for DIVIDER");
                    $stop;
                end
            endcase
        else
            sc_reg0[3:0] = 4'b0000;
    end

    always @(GLOGEN)
    begin
        if(GLOGEN)
            case(ADC_MODE)
                "DEFAULT"       : sc_reg1[15:14] = 2'b00;
                "SINGLE_PASS"   : sc_reg1[15:14] = 2'b01;
                "CONTINUE_SEQ"  : sc_reg1[15:14] = 2'b10;
                "SINGLE_CHANNEL": sc_reg1[15:14] = 2'b11;
                default:
                begin
                    $display ("GTP_ADC_E1 error: illegal setting for ADC_MODE");
                    $stop;
                end
            endcase
        else
            sc_reg1[15:14] = 2'b00;
    end

    always @(GLOGEN)
    begin
        if(GLOGEN)
            case(EVENT_DRIVE)
                "FALSE" : sc_reg1[13] = 1'b0;
                "TRUE"  : sc_reg1[13] = 1'b1;
                default:
                begin
                    $display ("GTP_ADC_E1 error: illegal setting for EVENT_DRIVE");
                    $stop;
                end
            endcase
        else
            sc_reg1[13] = 1'b0;
    end

    always @(GLOGEN)
    begin
        if(GLOGEN)
            case(ADC_MODE_1MSPS)
                "FALSE" : sc_reg1[12] = 1'b0;
                "TRUE"  : sc_reg1[12] = 1'b1;
                default:
                begin
                    $display ("GTP_ADC_E1 error: illegal setting for ADC_MODE_1MSPS");
                    $stop;
                end
            endcase
        else
            sc_reg1[12] = 1'b0;
    end

    always @(GLOGEN)
    begin
        if(GLOGEN)
            case(CLKSWITCH)
                "FALSE" : sc_reg1[11] = 1'b0;
                "TRUE"  : sc_reg1[11] = 1'b1;
                default:
                begin
                    $display ("GTP_ADC_E1 error: illegal setting for CLKSWITCH");
                    $stop;
                end
            endcase
        else
            sc_reg1[11] = 1'b0;
    end

    always @(GLOGEN)
    begin
        if(GLOGEN)
            case(INTERNAL_VOL_SEL)
                "VDD33" : sc_reg1[7:6] = 2'b01;
                "VDD11" : sc_reg1[7:6] = 2'b10;
                "VDDM"  : sc_reg1[7:6] = 2'b11;
                default:
                begin
                    $display ("GTP_ADC_E1 error: illegal setting for INTERNAL_VOL_SEL");
                    $stop;
                end
            endcase
        else
            sc_reg1[7:6] = 2'b00;
    end

    always @(GLOGEN)
    begin
        if(GLOGEN)
            case(SINGLE_CH_SEL)
                "0" : sc_reg1[5:2] = 4'b0000;
                "1" : sc_reg1[5:2] = 4'b0001;
                "2" : sc_reg1[5:2] = 4'b0010;
                "3" : sc_reg1[5:2] = 4'b0011;
                "4" : sc_reg1[5:2] = 4'b0100;
                "5" : sc_reg1[5:2] = 4'b0101;
                "6" : sc_reg1[5:2] = 4'b0110;
                "7" : sc_reg1[5:2] = 4'b0111;
                "8" : sc_reg1[5:2] = 4'b1000;
                "9" : sc_reg1[5:2] = 4'b1001;
                "10": sc_reg1[5:2] = 4'b1010;
                "11": sc_reg1[5:2] = 4'b1011;
                "12": sc_reg1[5:2] = 4'b1100;
                "13": sc_reg1[5:2] = 4'b1101;
                "14": sc_reg1[5:2] = 4'b1110;
                "15": sc_reg1[5:2] = 4'b1111;
                default:
                begin
                    $display ("GTP_ADC_E1 error: illegal setting for SINGLE_CH_SEL");
                    $stop;
                end
            endcase
        else
            sc_reg1[5:2] = 4'b0000;
    end

    always @(GLOGEN)
    begin
        if(GLOGEN)
            case(SINGLE_CH_IN)
                "SINGLE_END" : sc_reg1[1:0] = 2'b00;
                "UNIPOLAR"   : sc_reg1[1:0] = 2'b01;
                "BIPOLAR"    : sc_reg1[1:0] = 2'b11;
                default:
                begin
                    $display ("GTP_ADC_E1 error: illegal setting for SINGLE_CH_IN");
                    $stop;
                end
            endcase
        else
            sc_reg1[1:0] = 2'b00;
    end

    always @(GLOGEN)
    begin
        if(GLOGEN)
            case(SEQ_CH11_10_SEL)
                "NONE" : sc_reg2[11:10] = 2'b00;
                "CH10" : sc_reg2[11:10] = 2'b01;
                "CH11" : sc_reg2[11:10] = 2'b10;
                "ALL"  : sc_reg2[11:10] = 2'b11;
                default:
                begin
                    $display ("GTP_ADC_E1 error: illegal setting for SEQ_CH11_10_SEL");
                    $stop;
                end
            endcase
        else
            sc_reg2[11:10] = 2'b00;
    end

    always @(GLOGEN)
    begin
        if(GLOGEN)
            case(SEQ_CH9_8_SEL)
                "NONE" : sc_reg2[9:8] = 2'b00;
                "CH8"  : sc_reg2[9:8] = 2'b01;
                "CH9"  : sc_reg2[9:8] = 2'b10;
                "ALL"  : sc_reg2[9:8] = 2'b11;
                default:
                begin
                    $display ("GTP_ADC_E1 error: illegal setting for SEQ_CH9_8_SEL");
                    $stop;
                end
            endcase
        else
            sc_reg2[9:8] = 2'b00;
    end

    always @(GLOGEN)
    begin
        if(GLOGEN)
            case(SEQ_CH7_6_SEL)
                "NONE" : sc_reg2[7:6] = 2'b00;
                "CH6"  : sc_reg2[7:6] = 2'b01;
                "CH7"  : sc_reg2[7:6] = 2'b10;
                "ALL"  : sc_reg2[7:6] = 2'b11;
                default:
                begin
                    $display ("GTP_ADC_E1 error: illegal setting for SEQ_CH7_6_SEL");
                    $stop;
                end
            endcase
        else
            sc_reg2[7:6] = 2'b00;
    end

    always @(GLOGEN)
    begin
        if(GLOGEN)
            case(SEQ_CH5_4_SEL)
                "NONE" : sc_reg2[5:4] = 2'b00;
                "CH4"  : sc_reg2[5:4] = 2'b01;
                "CH5"  : sc_reg2[5:4] = 2'b10;
                "ALL"  : sc_reg2[5:4] = 2'b11;
                default:
                begin
                    $display ("GTP_ADC_E1 error: illegal setting for SEQ_CH5_4_SEL");
                    $stop;
                end
            endcase
        else
            sc_reg2[5:4] = 2'b00;
    end

    always @(GLOGEN)
    begin
        if(GLOGEN)
            case(SEQ_CH3_2_SEL)
                "NONE" : sc_reg2[3:2] = 2'b00;
                "CH2"  : sc_reg2[3:2] = 2'b01;
                "CH3"  : sc_reg2[3:2] = 2'b10;
                "ALL"  : sc_reg2[3:2] = 2'b11;
                default:
                begin
                    $display ("GTP_ADC_E1 error: illegal setting for SEQ_CH3_2_SEL");
                    $stop;
                end
            endcase
        else
            sc_reg2[3:2] = 2'b00;
    end

    always @(GLOGEN)
    begin
        if(GLOGEN)
            case(SEQ_CH1_0_SEL)
                "NONE" : sc_reg2[1:0] = 2'b00;
                "CH0"  : sc_reg2[1:0] = 2'b01;
                "CH1"  : sc_reg2[1:0] = 2'b10;
                "ALL"  : sc_reg2[1:0] = 2'b11;
                default:
                begin
                    $display ("GTP_ADC_E1 error: illegal setting for SEQ_CH1_0_SEL");
                    $stop;
                end
            endcase
        else
            sc_reg2[1:0] = 2'b00;
    end

    always @(GLOGEN)
    begin
        if(GLOGEN)
            case(SEQ_CH11_10_IN)
                "SINGLE_END" : sc_reg3[11:10] = 2'b00;
                "UNIPOLAR"   : sc_reg3[11:10] = 2'b01;
                "BIPOLAR"    : sc_reg3[11:10] = 2'b11;
                default:
                begin
                    $display ("GTP_ADC_E1 error: illegal setting for SEQ_CH11_10_IN");
                    $stop;
                end
            endcase
        else
            sc_reg3[11:10] = 2'b00;
    end

    always @(GLOGEN)
    begin
        if(GLOGEN)
            case(SEQ_CH9_8_IN)
                "SINGLE_END" : sc_reg3[9:8] = 2'b00;
                "UNIPOLAR"   : sc_reg3[9:8] = 2'b01;
                "BIPOLAR"    : sc_reg3[9:8] = 2'b11;
                default:
                begin
                    $display ("GTP_ADC_E1 error: illegal setting for SEQ_CH9_8_IN");
                    $stop;
                end
            endcase
        else
            sc_reg3[9:8] = 2'b00;
    end

    always @(GLOGEN)
    begin
        if(GLOGEN)
            case(SEQ_CH7_6_IN)
                "SINGLE_END" : sc_reg3[7:6] = 2'b00;
                "UNIPOLAR"   : sc_reg3[7:6] = 2'b01;
                "BIPOLAR"    : sc_reg3[7:6] = 2'b11;
                default:
                begin
                    $display ("GTP_ADC_E1 error: illegal setting for SEQ_CH7_6_IN");
                    $stop;
                end
            endcase
        else
            sc_reg3[7:6] = 2'b00;
    end

    always @(GLOGEN)
    begin
        if(GLOGEN)
            case(SEQ_CH5_4_IN)
                "SINGLE_END" : sc_reg3[5:4] = 2'b00;
                "UNIPOLAR"   : sc_reg3[5:4] = 2'b01;
                "BIPOLAR"    : sc_reg3[5:4] = 2'b11;
                default:
                begin
                    $display ("GTP_ADC_E1 error: illegal setting for SEQ_CH5_4_IN");
                    $stop;
                end
            endcase
        else
            sc_reg3[5:4] = 2'b00;
    end

    always @(GLOGEN)
    begin
        if(GLOGEN)
            case(SEQ_CH3_2_IN)
                "SINGLE_END" : sc_reg3[3:2] = 2'b00;
                "UNIPOLAR"   : sc_reg3[3:2] = 2'b01;
                "BIPOLAR"    : sc_reg3[3:2] = 2'b11;
                default:
                begin
                    $display ("GTP_ADC_E1 error: illegal setting for SEQ_CH3_2_IN");
                    $stop;
                end
            endcase
        else
            sc_reg3[3:2] = 2'b00;
    end

    always @(GLOGEN)
    begin
        if(GLOGEN)
            case(SEQ_CH1_0_IN)
                "SINGLE_END" : sc_reg3[1:0] = 2'b00;
                "UNIPOLAR"   : sc_reg3[1:0] = 2'b01;
                "BIPOLAR"    : sc_reg3[1:0] = 2'b11;
                default:
                begin
                    $display ("GTP_ADC_E1 error: illegal setting for SEQ_CH1_0_IN");
                    $stop;
                end
            endcase
        else
            sc_reg3[1:0] = 2'b00;
    end

    always @(GLOGEN)
    begin
        if(GLOGEN)
        begin
            sc_reg4[15:8] = TEMP_SENSOR_HIGH;
            sc_reg4[7:0]  = TEMP_SENSOR_LOW;
        end
        else
            sc_reg4[15:0] = 16'h0000;
    end

    always @(GLOGEN)
    begin
        if(GLOGEN)
            if(ADC_EN_ENABLE == "TRUE")
                sc_ad_en_enable = 1'b1;
            else if(ADC_EN_ENABLE == "FALSE")
                sc_ad_en_enable = 1'b0;
            else
                begin
                    $display ("GTP_ADC_E1 error: illegal setting for ADC_EN_ENABLE");
                    $stop;
                end
        else
            sc_ad_en_enable = 1'b0;
    end

    /////rtl code begin/////
    adc_logic_top   adc_logic_top(
        .sc_reg0         (sc_reg0    ),
        .sc_reg1         (sc_reg1    ),
        .sc_reg2         (sc_reg2    ),
        .sc_reg3         (sc_reg3    ),
        .sc_reg4         (sc_reg4    ),

        .sc_ad_en_enable (sc_ad_en_enable),

        .ad_en           (ADC_EN     ),
        .rst_n           (RST_N      ),
        .loadn_sc        (LOADSC_N   ),
        .dclk            (DCLK       ),
        .den             (DEN        ),
        .di              (DI         ),
        .dwe             (DWE        ),
        .daddr           (DADDR      ),
        .tck             (TCK        ),
        .flg_jdrp        (FLG_JDRP   ),
        .clockdr         (CLOCKDR    ),
        .capturedr       (CAPTUREDR  ),
        .shiftdr         (SHIFTDR    ),
        .updatedr        (UPDATEDR   ),
        .tdi             (TDI        ),
        .glogen          (GLOGEN     ),
        .convst          (CONVST     ),
        .clk_osc         (CLK_OSC    ),
        .por_n           (POR_N      ),

    ///////////////to adc_core_top///////////////
        .ad_done         (ad_done    ),
        .ad_dat          (ad_dat     ),

    ////out
        .ad_clk          (ad_clk     ),
        .ad_rstn         (ad_rstn    ),
        .ad_do_offset    (ad_do_offset),
        .ad_do_gain      (ad_do_gain  ),
        .ad_offset       (ad_offset   ),
        .ad_mode_diff_en (ad_mode_diff_en),
        .ad_mux          (ad_mux      ),
        .ad_sela         (ad_sela     ),
        .ad_selb         (ad_selb     ),
        .ad_bias_pd      (ad_bias_pd  ),
        .ad_clk_en       (ad_clk_en   ),
        .ad_fs_g         (ad_fs_g     ),
        .ad_vcm_g        (ad_vcm_g    ),
        .ad_ref_sel      (ad_ref_sel  ),
        .ad_cref_sel     (ad_cref_sel ),

    /////////////////////////////////////////

        .over_temp       (OVER_TEMP   ),
        .over_temp_ccs   (over_temp_ccs),

        .logic_done      (LOGIC_DONE  ),
        .dbusy           (DBUSY       ),
        .dataout         (DO          ),
        .drdy            (DRDY        ),
        .dmodified       (DMODIFIED   ),
        .tdo             (TDO         )
        );

    /////instance/////
    ADC_CORE_TOP ADC_CORE_TOP(
        .VAUX                (VAUX           ),
        .VA                  (VA             ),
        .VREF_EXT            (VREF_EXT       ),
        .VDD33               (VDD33          ),
        .VDD11               (VDD11          ),
        .VDDM                (VDDM           ),
        .VDD33A              (VDD33A         ),
        .VSSA                (VSSA           ),
        .VSS                 (VSS            ),
        .VTEMP_N             (VTEMP_N        ),
        .VTEMP_P             (VTEMP_P        ),
        .IBREF10U            (IBREF10U       ),
        .IB10U_IN            (IB10U_IN       ),
        .AD_CLK              (ad_clk         ),
        .AD_RSTN             (ad_rstn        ),
        .AD_MUX              (ad_mux         ),
        .AD_SELA             (ad_sela        ),
        .AD_SELB             (ad_selb        ),
        .AD_MODE_DIFF_EN     (ad_mode_diff_en),
        .AD_BIAS_PD          (ad_bias_pd     ),
        .AD_CLK_EN           (ad_clk_en      ),
        .AD_OFFSET           (ad_offset      ),
        .AD_FS_G             (ad_fs_g        ),
        .AD_VCM_G            (ad_vcm_g       ),
        .AD_GAIN_SEL         ({VSSA,VSSA}    ),
        .AD_REF_SEL          (ad_ref_sel     ),
        .AD_CREF_SEL         (ad_cref_sel    ),
        .AD_DO_OFFSET        (ad_do_offset   ),
        .AD_DO_GAIN          (ad_do_gain     ),
        .AD_DAT              (ad_dat         ),
        .AD_DONE             (ad_done        ),
        .VREF_BUF            (ad_vref_test   )
        );

    // pragma translate_on
endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: Internal simulation model
// Filename: GTP_IOBUFE.v
//
// Functional description: Input/Output Buffer
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_IOBUFE #(
    parameter IOSTANDARD = "DEFAULT",
    parameter SLEW_RATE = "SLOW",
    parameter DRIVE_STRENGTH = "8",
    parameter TERM_DDR = "ON"
)(
    output reg O,
    inout IO,
    input I,
    input EN,                    // 1: enable inbuf, normal mode; 0: disable inbuf, standby mode.
    input T
) /* synthesis syn_black_box */ ;

  initial begin
    case (IOSTANDARD)
    "LVTTL33", "PCI33", "LVCMOS33", "LVCMOS25", "LVCMOS18", "LVCMOS15", "LVCMOS12", "SSTL25_I", "SSTL25_II", "SSTL18_I", "SSTL18_II", "SSTL15_I", "SSTL15_II", "HSTL18_I", "HSTL18_II", "HSTL15_I", "SSTL15_I_CAL", "SSTL15_II_CAL", "HSTL15_I_CAL", "DEFAULT" :;
    default : begin
           $display("Attribute Syntax Error : The attribute IOSTANDARD on GTP_IOBUFE instance %m is set to %s.", IOSTANDARD);
           $finish;
              end
    endcase

    case (SLEW_RATE)
    "FAST", "SLOW":;
    default : begin
           $display("Attribute Syntax Error : The attribute SLEW_RATE on GTP_IOBUFE instance %m is set to %s.", SLEW_RATE);
           $finish;
              end
    endcase

    case (DRIVE_STRENGTH)
    "2", "4", "6", "8", "12", "16", "24":;
    default : begin
           $display("Attribute Syntax Error : The attribute DRIVE_STRENGTH on GTP_IOBUFE instance %m is set to %s.", DRIVE_STRENGTH);
           $finish;
              end
    endcase

    case (TERM_DDR)
    "ON", "OFF" :;
    default : begin
           $display("Attribute Syntax Error : The attribute TERM_DDR on GTP_IOBUFE instance %m is set to %s.", TERM_DDR);
           $finish;
              end
    endcase
    end

//    buf (O, IO);

    bufif0 (IO, I, T);

    always @(*)
    begin
        if (EN == 1'b1)
            O = IO;
        else
            O = 1'b1;
    end

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_IPAL.v
//
// Functional description: the simulation model of configuration and readback
//
// Parameter description:
//      
//
// Port description:
//      
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_IPAL
#(
    parameter DATA_WIDTH = "X8",
    parameter [31:0] IDCODE = 32'haaaa5555,
    parameter MEM_DEPTH = 1616
)
(
    input             RST_N  ,
    
    input             CLK   ,
    input      [7:0]  DI   ,
    input             CS_N  ,
    input             RW_SEL,
    output     [7:0]  DO  ,
    output            BUSY
);

ipal_gtp_wrap
#(
.DATA_WIDTH       (DATA_WIDTH),
.IDCODE           (IDCODE    ),
.MEM_DEPTH        (MEM_DEPTH )
)
GTP_IPAL_WRAP
(
.RST_N            (RST_N     ),
.CLK              (CLK       ),
.DI               (DI        ),
.CS_N             (CS_N      ),
.RW_SEL           (RW_SEL    ),
.DO               (DO        ),
.BUSY             (BUSY      )
);

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_IGDES4.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_IGDES4 #(
parameter GRS_EN = "TRUE", //"TRUE"; "FALSE"
parameter LRS_EN = "TRUE",  //"TRUE"; "FALSE"
parameter DPI_EN = "FALSE"  //"TRUE"; "FALSE"
)(
output [3:0] Q,
output [1:0] DPI_STS,
input [1:0] DPI_CTRL,
input DPI_STS_CLR_N,
input PADI,
input DESCLK,
input RCLK,
input RST
);

//synthesis translate_off
wire [7:0] PADI_D;
reg DPI_P;
reg [1:0] DPI_STS_R;
wire COMP_BEFORE;
wire COMP_AFTER;
wire COMP_BEFORE_D;
wire COMP_AFTER_D;
wire PD_BEFORE;
wire PD_AFTER;
wire DPI_BEFORE_POS_REG_T;
wire DPI_AFTER_POS_REG_T;
wire DPI_BEFORE_NEG_REG_T;
wire DPI_AFTER_NEG_REG_T;
wire AFTER_POS;
wire BEFORE_POS;
wire AFTER_NEG;
wire BEFORE_NEG;
reg DPI_N_reg;
reg DPI_BEFORE;
reg DPI_AFTER;
reg DPI_BEFORE_POS_REG;
reg DPI_BEFORE_NEG_REG;
reg DPI_AFTER_POS_REG;
reg DPI_AFTER_NEG_REG;
reg [3:0] shift_reg;
reg [3:0] capture_reg;
reg capture_en_b;
reg capture_en;
reg [3:0] Q_reg;

initial begin
DPI_P                = 0;
DPI_STS_R            = 0;
DPI_N_reg            = 0;
DPI_BEFORE           = 0;
DPI_AFTER            = 0;
DPI_BEFORE_POS_REG   = 0;
DPI_BEFORE_NEG_REG   = 0;
DPI_AFTER_POS_REG    = 0;
DPI_AFTER_NEG_REG    = 0;
shift_reg            = 0;
capture_reg          = 0;
capture_en_b         = 0;
capture_en           = 0;
Q_reg                = 0; 
end


assign global_rstn = (GRS_EN == "TRUE") ? GRS_INST.GRSNET : 1'b1;
assign lsr_rstn = LRS_EN == "TRUE" ? (~RST) : 1'b1;


assign  #0.05 PADI_D[0] =  PADI;
assign  #0.05 PADI_D[1] =  PADI_D[0];
assign  #0.05 PADI_D[2] =  PADI_D[1];
assign  #0.05 PADI_D[3] =  PADI_D[2];
assign  #0.05 PADI_D[4] =  PADI_D[3];
assign  #0.05 PADI_D[5] =  PADI_D[4];
assign  #0.05 PADI_D[6] =  PADI_D[5];
assign  #0.05 PADI_D[7] =  PADI_D[6];

assign PADI_SAMPLE = (DPI_EN == "TRUE") ? PADI_D[3] : PADI;

always @(posedge DESCLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_P <= 0;
   else if (!lsr_rstn)
      DPI_P <= 0;
   else
      DPI_P <= PADI_SAMPLE;
end

always @(negedge DESCLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_N_reg <= 0;
   else if (!lsr_rstn)
      DPI_N_reg <= 0;
   else 
      DPI_N_reg <= PADI_SAMPLE;
end

always @(*) begin
   case (DPI_CTRL[1:0])
      2'd0:    begin DPI_BEFORE = PADI_D[2];  DPI_AFTER = PADI_D[4]; end
      2'd1:    begin DPI_BEFORE = PADI_D[1];  DPI_AFTER = PADI_D[5]; end
      2'd2:    begin DPI_BEFORE = PADI_D[0];  DPI_AFTER = PADI_D[6]; end
      default: begin DPI_BEFORE = PADI;       DPI_AFTER = PADI_D[7]; end
   endcase
end

always @(posedge DESCLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_BEFORE_POS_REG <= 0;
   else if (!lsr_rstn)
      DPI_BEFORE_POS_REG <= 0;
   else   
      DPI_BEFORE_POS_REG <= DPI_BEFORE;
end

always @(negedge DESCLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_BEFORE_NEG_REG <= 0;
   else if (!lsr_rstn)
      DPI_BEFORE_NEG_REG <= 0;
   else     
      DPI_BEFORE_NEG_REG <= DPI_BEFORE;
end


always @(posedge DESCLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_AFTER_POS_REG <= 0;
   else if (!lsr_rstn)
      DPI_AFTER_POS_REG <= 0;
   else   
      DPI_AFTER_POS_REG <= DPI_AFTER;
end


always @(negedge DESCLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_AFTER_NEG_REG <= 0;
   else if (!lsr_rstn)
      DPI_AFTER_NEG_REG <= 0;
   else     
      DPI_AFTER_NEG_REG <= DPI_AFTER;
end


assign BEFORE_POS = DPI_BEFORE_POS_REG_T ^ DPI_P;
assign DPI_BEFORE_POS_REG_T = (DPI_EN == "TRUE") ? DPI_BEFORE_POS_REG : 0;

assign AFTER_POS = DPI_AFTER_POS_REG_T ^ DPI_P;
assign DPI_AFTER_POS_REG_T = (DPI_EN == "TRUE") ? DPI_AFTER_POS_REG : 0;

assign BEFORE_NEG = DPI_BEFORE_NEG_REG_T ^ DPI_N_reg;
assign DPI_BEFORE_NEG_REG_T = (DPI_EN == "TRUE") ? DPI_BEFORE_NEG_REG : 0;

assign AFTER_NEG = DPI_AFTER_NEG_REG_T ^ DPI_N_reg;
assign DPI_AFTER_NEG_REG_T = (DPI_EN == "TRUE") ? DPI_AFTER_NEG_REG : 0;


assign COMP_BEFORE = BEFORE_POS || BEFORE_NEG;
assign COMP_AFTER = AFTER_POS || AFTER_NEG;

assign #0.1 COMP_BEFORE_D = COMP_BEFORE;
assign #0.1 COMP_AFTER_D = COMP_AFTER;

assign PD_BEFORE = COMP_BEFORE && COMP_BEFORE_D;
assign PD_AFTER = COMP_AFTER && COMP_AFTER_D;

always @(posedge DPI_STS_CLR_N or negedge global_rstn or negedge lsr_rstn or posedge PD_BEFORE) begin
   if (!global_rstn)
      DPI_STS_R[0] <= 0;
   else if (!lsr_rstn)
      DPI_STS_R[0] <= 0;
   else if (PD_BEFORE)
      DPI_STS_R[0] <= 1;
   else
      DPI_STS_R[0] <= 1'b0;
end

always @(posedge DPI_STS_CLR_N or negedge global_rstn or negedge lsr_rstn or posedge PD_AFTER) begin
   if (!global_rstn)
      DPI_STS_R[1] <= 0;
   else if (!lsr_rstn)
      DPI_STS_R[1] <= 0;
   else if (PD_AFTER)
      DPI_STS_R[1] <= 1;
   else
      DPI_STS_R[1] <= 1'b0;
end


assign DPI_STS[0] = DPI_STS_R[0];
assign DPI_STS[1] = DPI_STS_R[1];

//assign DPI_STS[0] = (DPI_EN == "TRUE") ? DPI_STS_T[0] : 1;
//assign DPI_STS[1] = (DPI_EN == "TRUE") ? DPI_STS_T[1] : 1;

always @(posedge DESCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      shift_reg <= 0;
   else if (!lsr_rstn)
      shift_reg <= 0;
   else
      shift_reg <= {DPI_N_reg, DPI_P, shift_reg[3:2]};

always @(posedge DESCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn) begin
      capture_en_b <= 0;
      capture_en   <= 0;
   end   
   else if (!lsr_rstn) begin
      capture_en_b <= 0;
      capture_en   <= 0;      
   end
   else begin
      capture_en_b <= ~ capture_en_b;
      capture_en   <= capture_en_b;            
   end   

always @(posedge DESCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      capture_reg <= 0;
   else if (!lsr_rstn)
      capture_reg <= 0;
   else if (capture_en)
      capture_reg <= shift_reg;
      
always @(posedge RCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      Q_reg <= 0;
   else if (!lsr_rstn)
      Q_reg <= 0;
   else
      Q_reg <= capture_reg;      

assign Q = Q_reg;      
//synthesis translate_on

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_CLKBUFGCE.v
//
// Functional description: Global Clock Buffer
//
// Parameter description:
//      DEFAULT_VALUE
//
// Port description:
//
// Revision:
//    06/18/14 - Initial version.
//    05/11/14 - 
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_CLKBUFGCE
#(
    parameter DEFAULT_VALUE = 1'b0,  //1'b0, 1'b1
    parameter SIM_DEVICE = "TITAN"   //"TITAN", "LOGOS", "COMPACT", "LOGOS2"
) (
    output wire CLKOUT ,
    input CLKIN,
    input CE
);
    wire clkout0;
    wire clkout1;
    wire clkout1_pos;
    wire clkout1_neg;

    reg  SWITCH;
    reg  ce_d_pos;
    reg  ce_2d_pos;
    reg  ce_d_neg;
    reg  ce_2d_neg;
    reg  init_set;

    initial begin
       case (SIM_DEVICE)
            "TITAN": SWITCH = 0;
            "LOGOS","COMPACT","LOGOS2": SWITCH = 1;         
            default: begin
                $display("ERROR: GTP_CLKBUFGMUX instance %m parameter SIM_DEVICE value: %s is illegal. The legal values are TITAN or LOGOS or COMPACT or LOGOS2.", SIM_DEVICE);
                $finish;
            end
       endcase
    end

    initial begin
        ce_d_pos <= CE;
        ce_2d_pos <= CE;
        ce_d_neg <= CE;
        ce_2d_neg <= CE;
        init_set <= 1;
        #0.1 init_set <= 0;
    end

    assign CLKOUT = SIM_DEVICE == "TITAN" ? clkout0 : clkout1;
    assign clkout0 = CE ? CLKIN:DEFAULT_VALUE;
    assign clkout1 = DEFAULT_VALUE ? clkout1_pos : clkout1_neg;
    assign clkout1_pos = ce_2d_pos ? CLKIN : 1'b1;
    assign clkout1_neg = ce_2d_neg ? CLKIN : 1'b0;
    
    always@(posedge CLKIN) begin
        if(DEFAULT_VALUE && !init_set) begin
            ce_d_pos <= CE;
            ce_2d_pos <= ce_d_pos;
        end
        else begin
            ce_d_pos <= CE;
            ce_2d_pos <= CE;
        end
    end

    always@(negedge CLKIN) begin
        if(!DEFAULT_VALUE && !init_set) begin
            ce_d_neg <= CE;
            ce_2d_neg <= ce_d_neg;
        end
        else begin
            ce_d_neg <= CE;
            ce_2d_neg <= CE;
        end
    end
endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: Internal simulation model
// Filename: GTP_BANKCTL.v
//
// Functional description: Bank controller 
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_BANKCTL #(
    parameter DIFFO_DYN_EN = "FALSE",
    parameter DIFFI_DYN_EN = "FLASE",
    parameter BANK_LOC = "BK0" // IO Bank location: "BK0", "BK1", "BK2", "BK3", "BK4", "BK5"
)(
    input OE_N,
    input IE_N
) /* synthesis syn_black_box */ ;
  
  initial begin
    case (DIFFO_DYN_EN)
    "TRUE", "FALSE"  :;
    default : begin
           $display("Attribute Syntax Error : The attribute DIFFO_DYN_EN on GTP_BANKCTL instance %m is set to %s.", DIFFO_DYN_EN);
           $finish;
              end
    endcase

    case (DIFFI_DYN_EN)
    "TRUE", "FALSE" :;
    default : begin
           $display("Attribute Syntax Error : The attribute DIFFI_DYN_EN on GTP_BANKCTL instance %m is set to %s.", DIFFI_DYN_EN);
           $finish;
              end
    endcase
    end


endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_IOCLKMUX.v
//
// Functional description: io Clock iockbrgmux
//
// Parameter description:
//      xxxx
//
// Port description:
//
// Revision:
//    10/10/18 - Initial version.
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_IOCLKMUX
    (
    output  CLKOUT,
    input CLKIN0,
    input CLKIN1,
    input SEL
);



reg sel_d_a;
reg sel_d_b;
reg [1:0] glitch_free_sel;
reg clk_sel;

wire [1:0] selector;
wire iockbrgsel_ctrl;
wire sel_a2b;
wire sel_b2a;
wire clk_a_buf;
wire clk_b_buf;
wire iockbrgsel_buf;
wire iockbrgsel_ctrl_b;
reg [2:0] iockbrg_mode;
wire reg1_out;
wire reg0_out;


initial
begin
 iockbrg_mode = 3'b000;
end

assign  selector = glitch_free_sel;
assign iockbrgsel_ctrl = ( iockbrg_mode[1] &  iockbrg_mode[2] )? 1'b1:1'b0;
assign iockbrgsel_ctrl_b = ~iockbrgsel_ctrl;
assign sel_a2b = (iockbrgsel_ctrl & iockbrg_mode[0])? 1'b1:1'b0;
assign sel_b2a = (iockbrgsel_ctrl_b | iockbrg_mode[0])? 1'b1:1'b0;

assign  clk_a_buf = sel_a2b?CLKIN1:CLKIN0;
assign  clk_b_buf = sel_b2a?CLKIN1:CLKIN0;
assign  iockbrgsel_buf = SEL;



wire clk_sel_reg;
assign clk_sel_reg = iockbrgsel_buf? clk_a_buf:clk_b_buf;

wire iockbrgsel_delay;
assign #0.2 iockbrgsel_delay = iockbrgsel_buf; 


reg sel_reg0;


initial begin
  sel_reg0 = 1'b0;
  sel_d_a = 1'b0;
  sel_d_b = 1'b0;
end


  always@ (negedge clk_sel_reg )        
  begin                                       
     if (iockbrgsel_delay == 1'b1)
        sel_reg0 <= 1'b1;
     else
        sel_reg0 <= 1'b0;
  end    


  always@ (negedge clk_sel_reg )         
  begin
     if (sel_reg0 == 1'b0)
        sel_d_a <= 1'b0;
      else
        sel_d_a <= 1'b1;
  end


wire clk_reg2;
reg  sel_reg2;
wire sel_in_buf;

initial begin
   sel_reg2 =1'b0;
end


assign sel_in_buf = iockbrgsel_buf;
assign clk_reg2 = sel_in_buf? clk_b_buf: clk_a_buf;

  always@ (negedge clk_reg2  )        
    begin
          if (sel_d_a == 1'b0)
          sel_reg2 <= 1'b0;
          else
          sel_reg2 <= 1'b1;
    end





wire clk_reg3;

assign clk_reg3 = sel_in_buf? clk_b_buf: clk_a_buf;

  always@ (negedge clk_reg3 )          
    begin
          if (sel_reg2 == 1'b0)
          sel_d_b <= 1'b0;
          else
          sel_d_b <= 1'b1;
    end







always@ (*) 
begin
   casex ({sel_d_b, sel_d_a})
      2'b00: glitch_free_sel = 2'b00; 
      2'b01: glitch_free_sel = 2'b11;
      2'b10: glitch_free_sel = 2'b11;
      2'b11: glitch_free_sel = 2'b01;
      default: glitch_free_sel = 2'b00;
   endcase
end



always @(*) begin
   case (selector)
      2'b00: clk_sel = CLKIN0;
      2'b01: clk_sel = CLKIN1;
      2'b10: clk_sel = 1'b0;
      2'b11: clk_sel = 1'b0;
      default: clk_sel = CLKIN0;
   endcase   
end


assign reg1_out= reg0_out?1'b0:1'b1;
assign reg0_out = (sel_d_b | iockbrgsel_ctrl_b )? 1'b0:1'b1;


assign  CLKOUT = reg1_out? clk_sel : 1'b0;




endmodule







//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_OGSER10.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_OGSER10 #(
parameter GRS_EN = "TRUE", //"TRUE"; "FALSE"  
parameter LRS_EN = "TRUE"   //"TRUE"; "FALSE"  
)(
output  PADO,
input [9:0] D,
input RCLK,
input SERCLK,
input RST
);

//synthesis translate_off
reg [9:0] d_rclk;
reg [2:0] cnt;                                     
reg [9:0] capture_r_reg;
reg [9:0] shift_r_reg;
wire capture_en;
reg PADO_POS;
reg PADO_NEG;

initial begin
d_rclk        = 0;
cnt           = 0;                                     
capture_r_reg = 0;
shift_r_reg   = 0;
PADO_POS      = 0;
PADO_NEG      = 0;
end

assign global_rstn = (GRS_EN == "TRUE") ? GRS_INST.GRSNET : 1'b1; 
assign lsr_rstn = LRS_EN == "TRUE" ? (~RST) : 1'b1;                

always @(posedge RCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      d_rclk <= 0;
   else if (!lsr_rstn)
      d_rclk <= 0;
   else
      d_rclk <= D;
   
always @(posedge SERCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      cnt <= 0;
   else if (!lsr_rstn)
      cnt <= 0;
   else if (cnt == 4)
      cnt <= 0;
   else
      cnt <= cnt + 1;

assign capture_en = cnt == 4;      
assign shift_en = cnt == 4;
 
always @(posedge SERCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      capture_r_reg <= 0;
   else if (!lsr_rstn)
      capture_r_reg <= 0;
   else if (capture_en)
      capture_r_reg <= d_rclk;
   
always @(posedge SERCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      shift_r_reg <= 0;
   else if (!lsr_rstn)
      shift_r_reg <= 0;
   else if (capture_en)
      shift_r_reg <= capture_r_reg;
   else
      shift_r_reg <= {2'd0, shift_r_reg[9:2]};
   
always @(posedge SERCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      PADO_POS <= 0;
   else if (!lsr_rstn)
      PADO_POS <= 0;
   else
      PADO_POS <= shift_r_reg[1];
   
always @(negedge SERCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      PADO_NEG <= 0;
   else if (!lsr_rstn)
      PADO_NEG <= 0;
   else
      PADO_NEG <= shift_r_reg[0];
   
assign PADO =  SERCLK ? PADO_NEG : PADO_POS;

//synthesis translate_on

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_LUT7.v
//
// Functional description: 7-input Look-Up-Table
//
// Parameter description:
//      INIT: init value
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_LUT7
#(
    parameter [127:0] INIT = 128'h00000000_00000000_00000000_00000000
) (
    output wire Z,
    input wire I0, I1, I2, I3, I4, I5, I6
);

    wire z6a, z6b;

    GTP_LUT6 #(.INIT(INIT[63:0]))
        l6a (.I0(I0), .I1(I1), .I2(I2), .I3(I3), .I4(I4), .I5(I5), .Z(z6a));

    GTP_LUT6 #(.INIT(INIT[127:64]))
        l6b (.I0(I0), .I1(I1), .I2(I2), .I3(I3), .I4(I4), .I5(I5), .Z(z6b));

    GTP_MUX2LUT7 mxl7 (.I0(z6a), .I1(z6b), .S(I6), .Z(Z));

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_DLATCH_C.v
//
// Functional description: D-type latch with clear
//
// Parameter description:
//      INIT: init value
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_DLATCH_C
#(
    parameter GRS_EN = "TRUE",
    parameter INIT = 1'b0
) (
    output reg Q,
    input wire D,
    input wire G, C
);

    wire grs_n;
    wire grs, RS;

    tri1 grsnet = GRS_INST.GRSNET;
    assign grs_n=(GRS_EN=="TRUE")?grsnet:1'b1;

    not (grs, grs_n);
    or (RS, grs, C);

    initial Q = 1'bx;

    always @(D or G or RS) begin
        if (RS)
            Q <= 1'b0;
        else if (G)
            Q <= D;
    end

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_DFF_SE.v
//
// Functional description: D-type flip-flop with sync set and enable
//
// Parameter description:
//      INIT: init value
//
// Port description:
//      S: synchronous set
//      CE  : enable
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_DFF_SE
#(
    parameter GRS_EN = "TRUE",
    parameter INIT = 1'b1
) (
    output reg Q,
    input wire D,
    input wire CLK, S, CE
);

    wire grs_n;
    wire RS;

    tri1 grsnet = GRS_INST.GRSNET;
    assign grs_n=(GRS_EN=="TRUE")?grsnet:1'b1;

    not (RS, grs_n);

    initial Q = 1'bx;

    always @(posedge CLK or posedge RS) begin
        if (RS)
            Q <= 1'b1;
        else if (S)
            Q <= 1'b1;
        else if (CE)
            Q <= D;
    end

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_OSERDES.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//   2016/10/18: Remove OSERDES_MODE parameter value "NONE"
//   2018/03/14: ADD DYNAMIC MIPI SELECT
//   2018/03/29: delete MIPI_sel and MIPI_sel ctrl for DO
//   2018/08/17: change OGSER4/7/8 to OSER4/7/8
//               change OGDDR to ODDR 
//               by xxma
////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_OSERDES #(
parameter OSERDES_MODE = "ODDR",  //"ODDR","OMDDR","OSER4","OMSER4","OSER7","OSER8",OMSER8"
parameter WL_EXTEND = "FALSE",     //"TRUE"; "FALSE"
parameter GRS_EN = "TRUE",         //"TRUE"; "FALSE"
parameter LRS_EN = "TRUE",          //"TRUE"; "FALSE"
parameter TSDDR_INIT = 1'b0         //1'b0;1'b1
)(
output      DO,
output      TQ,
input [7:0] DI,
input [3:0] TI,
input       RCLK,
input       SERCLK,
input       OCLK,
input       RST
);  // synthesis syn_black_box

//synthesis translate_off
///////////////////////////////////////////////////////////////////////////
reg  [7:0] d_rclk;
reg  [3:0] t_rclk;
reg  [7:0] capture_d_reg;
reg  [3:0] capture_t_reg;
reg  [7:0] shift_d_reg;
reg  [3:0] shift_t_reg;
reg        DO_POS;
reg        TO_reg;
reg        DO_NEG;
wire       shift_en_oclk;
reg  [2:0] cnt;
reg  [1:0] cnt_oclk;
wire       cnt_rst;
wire       capture_en0;
wire       capture_en1;
reg        shift_en_oclk_d;

reg        rstn_dly;
reg        rstn_dly_oclk;
reg  [7:0] in_en;
wire [3:0] int_en;
reg        omem_mode;
reg  [3:0] odata_width;
wire       RCLK_buf;
wire       SERCLK_buf;
wire       OCLK_buf;
wire       DO_buf;
wire       TO_buf;
wire [7:0] DI_buf;
wire [3:0] TI_buf;
///////////////////////////////////////////////////////////////////////////
initial begin
    if(GRS_EN != "TRUE" && GRS_EN != "FALSE")
    begin
      $display("GTP_OSERDES Error: Illegal setting of GRS_EN %s",GRS_EN);
      $finish;
    end
    if(LRS_EN != "TRUE" && LRS_EN != "FALSE")
    begin
      $display("GTP_OSERDES Error: Illegal setting of LRS_EN %s",LRS_EN);
      $finish;
    end
    case(OSERDES_MODE)
        "ODDR":   begin
                     omem_mode = 0;
                     odata_width = 2;
                     in_en = 8'b0000_0011;
                   end
        "OMDDR":   begin
                     omem_mode = 1;
                     odata_width = 2;
                     in_en = 8'b0000_0011;
                   end
        "OSER4":  begin
                     omem_mode = 0;
                     odata_width = 4;
                     in_en = 8'b0000_1111;
                   end
        "OMSER4":  begin
                     omem_mode = 1;
                     odata_width = 4;
                     in_en = 8'b0000_1111;
                   end
        "OSER7":  begin
                     omem_mode = 0;
                     odata_width = 7;
                     in_en = 8'b0111_1111;
                   end
        "OSER8":  begin
                     omem_mode = 0;
                     odata_width = 8;
                     in_en = 8'b1111_1111;
                   end
        "OMSER8":  begin
                     omem_mode = 1;
                     odata_width = 8;
                     in_en = 8'b1111_1111;
                   end
        default:   begin
                     $display("GTP_OSERDES Error: Illegal setting of OSERDES_MODE %s",OSERDES_MODE);
                     $finish;
                   end
    endcase
end

initial begin
d_rclk           = 0;
t_rclk           = 0;
capture_d_reg    = 0;
capture_t_reg    = 0;
shift_d_reg      = 0;
shift_t_reg      = 0;
DO_POS         = 0;
TO_reg         = 0;
DO_NEG         = 0;
cnt              = 0;
cnt_oclk         = 0;
shift_en_oclk_d  = 0;
end

///////////////////////////////////////////////////////////////////////////
assign DI_buf = in_en & DI;
assign TI_buf = {in_en[6],in_en[4],in_en[2],in_en[0]} & TI;
assign RCLK_buf = RCLK;
assign SERCLK_buf = (odata_width == 2) ? ((omem_mode) ? OCLK : RCLK) : SERCLK;
assign OCLK_buf =  (omem_mode) ? OCLK : ((odata_width == 2) ? RCLK : SERCLK);
assign DO = DO_buf;
assign TQ = TO_buf;

assign init = (TSDDR_INIT == 1'b0) ? 1'b0 : 1'b1;
///////////////////////////////////////////////////////////////////////////
assign global_rstn = (GRS_EN == "TRUE") ? GRS_INST.GRSNET : 1'b1;
assign lrs_rstn = (LRS_EN == "TRUE") ? (~RST) : 1'b1;
///////////////////////////////////////////////////////////////////////////
always @(posedge RCLK_buf or negedge global_rstn or negedge lrs_rstn) begin
   if (!global_rstn) begin
      d_rclk <= 0;
      t_rclk <= {4{init}};
   end
   else if (!lrs_rstn) begin
      d_rclk <= 0;
      t_rclk <= {4{init}};
   end
   else begin
      d_rclk <= DI_buf;
      t_rclk <= TI_buf;
   end
end
///////////////////////////////////////////////////////////////////////////
always @(posedge SERCLK_buf or negedge global_rstn or negedge lrs_rstn)
begin
   if (!global_rstn)
      rstn_dly <= 0;
   else if (!lrs_rstn)
      rstn_dly <= 0;
   else
      rstn_dly <= 1'b1;
end
always @(posedge SERCLK_buf or negedge global_rstn or negedge lrs_rstn)
begin
   if (!global_rstn)
      cnt <= 0;
   else if (!lrs_rstn || cnt_rst)
      cnt <= 0;
   else if (rstn_dly)
      cnt <= cnt + 1;
end

assign cnt_rst = (odata_width == 4) ? (cnt == 1) :
                ((odata_width == 8) ? (cnt == 3) :
                ((odata_width == 7) ? (cnt == 6) : 1'b1));
assign capture_en0 = (odata_width == 4) ? (cnt == 1) :
                    ((odata_width == 8) ? (cnt == 2) :
                    ((odata_width == 7) ? (cnt == 2) : 1'b1));
assign capture_en1 = cnt == 5;

always @(posedge SERCLK_buf or negedge global_rstn or negedge lrs_rstn)
begin
   if (!global_rstn)
   begin
      capture_d_reg <= 0;
      capture_t_reg <= {4{init}};
   end else if (!lrs_rstn)
   begin
      capture_d_reg <= 0;
      capture_t_reg <= {4{init}};
   end else
   begin
      if (capture_en0)
      begin
         capture_d_reg <= d_rclk;
         capture_t_reg <= t_rclk;
      end else if (capture_en1 && (odata_width == 7))
         capture_d_reg <= {d_rclk[6:0], capture_d_reg[6]};
   end
end
///////////////////////////////////////////////////////////////////////////
wire cnt_rst_oclk;
wire shift_en;
reg  shift_en_v;

always @(posedge OCLK_buf or negedge global_rstn or negedge lrs_rstn)
begin
   if (!global_rstn)
      rstn_dly_oclk <= 0;
   else if (!lrs_rstn)
      rstn_dly_oclk <= 0;
   else
      rstn_dly_oclk <= 1'b1;
end

always @(posedge OCLK_buf or negedge global_rstn or negedge lrs_rstn)
begin
   if (!global_rstn)
      cnt_oclk <= 0;
   else if (!lrs_rstn)
      cnt_oclk <= 0;
   else if (rstn_dly_oclk)
      cnt_oclk <= cnt_oclk + 1;
end

assign shift_en_oclk = (odata_width == 4) ? (cnt_oclk == 2 | cnt_oclk == 0 & rstn_dly_oclk) :
                      ((odata_width == 8) ? (cnt_oclk == 1) :
                      ((odata_width == 7) ? shift_en_v : 1'b0));

always @(posedge OCLK_buf or negedge global_rstn or negedge lrs_rstn)
begin
   if (!global_rstn)
   begin
      shift_en_v <= 0;
      shift_en_oclk_d <= 0;
   end else if (!lrs_rstn)
   begin
      shift_en_v <= 0;
      shift_en_oclk_d <= 0;
   end else begin
      shift_en_v <= capture_en0 | capture_en1;
      shift_en_oclk_d <= shift_en_oclk;
   end
end

assign shift_en = (WL_EXTEND == "FALSE") ? shift_en_oclk : shift_en_oclk_d;

always @(posedge OCLK_buf or negedge global_rstn or negedge lrs_rstn)
   if (!global_rstn) begin
      shift_d_reg <= 0;
      shift_t_reg <= {4{init}};
   end
   else if (!lrs_rstn) begin
      shift_d_reg <= 0;
      shift_t_reg <= {4{init}};
   end
   else if (shift_en) begin
      shift_d_reg <= capture_d_reg;
      shift_t_reg <= capture_t_reg;
   end
   else begin
      shift_d_reg <= {2'd0, shift_d_reg[7:2]};
      shift_t_reg <= {init, shift_t_reg[3:1]};
   end
///////////////////////////////////////////////////////////////////////////
always @(posedge OCLK_buf or negedge global_rstn or negedge lrs_rstn)
begin
   if (!global_rstn) begin
      DO_POS <= 0;
      TO_reg <= init;
   end else if (!lrs_rstn) begin
      DO_POS <= 0;
      TO_reg <= init;
   end else if(odata_width == 2)
   begin
      DO_POS <= capture_d_reg[1];
      TO_reg <= capture_t_reg[0];
   end else
   begin
      DO_POS <= shift_d_reg[1];
      TO_reg <= shift_t_reg[0];
   end
end

always @(negedge OCLK_buf or negedge global_rstn or negedge lrs_rstn)
begin
   if (!global_rstn) begin
      DO_NEG <= 0;
   end else if (!lrs_rstn) begin
      DO_NEG <= 0;
   end else if(odata_width == 2)
      DO_NEG <= capture_d_reg[0];
   else
      DO_NEG <= shift_d_reg[0];
end

assign DO_buf = OCLK_buf ? DO_NEG : DO_POS;
assign TO_buf = TO_reg;

//synthesis translate_on

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_MULTACC27.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

//P = MAC + A*B
module GTP_MULTACC27 #(
    parameter GRS_EN            = "TRUE", //"TRUE"; "FALSE"
    parameter SYNC_RST          = "FALSE", //"TRUE"; "FALSE"
    parameter INREG_EN          = "FALSE",  //"TRUE"; "FALSE"
    parameter PIPEREG_EN        = "FALSE",   //"TRUE"; "FALSE"
    parameter ACC_ADDSUB_OP     = 0,
    parameter DYN_ACC_ADDSUB_OP = 1,     //Select parameter ADDSUB or input ADDSUB
    parameter OVERFLOW_MASK     = 64'h0, //PSIZE = 64 OVERflow setting =  'h8000_0000_0000_00XX , bit width = PSIZE
    parameter PATTERN           = 64'h0, //compare pattern
    parameter MASKPAT           = 64'h0, //pattern mask
    parameter DYN_ACC_INIT      = 0,   //acc init value dynamic input
    parameter ACC_INIT_VALUE    = 64'h0  //acc init value parameter
) (
    output  [63:0] P,
    output  OVER,
    output  UNDER,
    output  EQZ,
    output  EQZM,
    output  EQOM,
    output  EQPAT,
    output  EQPATN,

    input   CE,
    input   RST,
    input   CLK,
    input   [26:0] A,
    input   [26:0] B,
    input   A_SIGNED,
    input   B_SIGNED,
    input   [63:0] ACC_INIT,
    input   ACC_ADDSUB,
    input   RELOAD
);

    wire [63:0] R;

    INT_PREADD_MULTACC #(
        . GRS_EN(GRS_EN),     
        . SYNC_RST(SYNC_RST),   
        . INREG_EN(INREG_EN),   
        . PIPEREG_EN(PIPEREG_EN), 
        . ACCUMADDSUB_OP(ACC_ADDSUB_OP), 
        . DYN_OP_SEL(DYN_ACC_ADDSUB_OP),     
        . ASIZE(27),    
        . BSIZE(27),    
        . PSIZE(64),    
        . PREADD_EN(0),
        . MASK(OVERFLOW_MASK),      
        . DYN_ACC_INIT(DYN_ACC_INIT),
        . ACC_INIT_VALUE(ACC_INIT_VALUE)               
    ) U_MACC (
        .CE(CE),
        .RST(RST),
        .CLK(CLK),
        .A(A),
        .B(B),
        .A_SIGNED(A_SIGNED),
        .B_SIGNED(B_SIGNED),
        .C_SIGNED(B_SIGNED),
        .C(27'b0),
        .PREADDSUB(1'b0),
        .ACCUM_INIT(ACC_INIT),
        .ACCUMADDSUB(ACC_ADDSUB),
        .RELOAD(RELOAD),
        .P(P),
        .OVER(OVER),
        .UNDER(UNDER),
        .R(R)     
    );

    INT_FLAG #(
        . GRS_EN(GRS_EN),
        . SYNC_RST(SYNC_RST),
        . PSIZE(64),
        . PATSIZE(64),
        . MASKPATSIZE(64),
        . OUTREG_EN("TRUE")
    ) U_FLAG (
        . CE(CE),
        . RST(RST),
        . CLK(CLK),
        . P(P),
        . PATTERN(PATTERN),
        . MASKPAT(MASKPAT),
        . OVERFLOW_MASK(OVERFLOW_MASK),
        . R(R),
        . eqz(EQZ),
        . eqzm(EQZM),
        . eqom(EQOM),
        . eqpat(EQPAT),
        . eqpatn(EQPATN)
    );

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_OSERDES_E1.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//2017/12/20 : initial version
//2018/01/02 : delete RST_EN & RSTC_EN
//             update ODDR_MODE
//2018/03/20 : fix bug2861
//2018/03/27 : change ODDR_MODE to OSERDES_MODE
//2018/03/30 : fix bug 2961
//2018/10/16 : fix bug 7114
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_OSERDES_E1 #(
parameter OSERDES_MODE = "OSER4", //"OSER4","OSER7","OSER8"
parameter GRS_EN = "TRUE"         //"TRUE"; "FALSE"
)(
output      DO,
input [7:0] DI,
input       RCLK,
input       OCLK,
input       RST
);  // synthesis syn_black_box

//synthesis translate_off
///////////////////////////////////////////////////////////////////////////
wire global_rstn;
wire local_rstn;
wire upd_stage0;
wire upd_stage1;
wire sel;
wire update0;
wire update1;

reg [7:0] t_r;
reg [7:0] m;
reg [7:0] up_r0;
reg [7:0] up_r1;
reg       f_reg;
reg       rstn_sync;
reg [1:0] cnt;
reg       select_reg;
reg       update0_reg;
reg       update1_reg;

initial begin
    if(GRS_EN != "TRUE" && GRS_EN != "FALSE")
    begin
      $display("GTP_OSERDES Error: Illegal setting of GRS_EN %s",GRS_EN);
      $finish;
    end
    if(OSERDES_MODE != "OSER4" && OSERDES_MODE != "OSER7" && OSERDES_MODE != "OSER8")
    begin
    $display("GTP_OSERDES Error: Illegal setting of OSERDES_MODE %s",OSERDES_MODE);
    $finish;
    end

end

initial
begin
   t_r           = 8'b0;
   m             = 8'b0;
   up_r0         = 8'b0;
   up_r1         = 8'b0;
   f_reg       = 1'b0;
   rstn_sync   = 1'b0;
   cnt         = 2'b0;
   select_reg    = 1'b0;
   update0_reg = 1'b0;
   update1_reg = 1'b0;
end
///////////////////////////////////////////////////////////////////////////
assign global_rstn = (GRS_EN == "TRUE") ? GRS_INST.GRSNET : 1'b1;
assign local_rstn = ~RST;
///////////////////////////////////////////////////////////////////////////

assign upd_stage0 = update0;
assign upd_stage1 = (OSERDES_MODE == "OSER7") ? update1 : update0;
///////////////////////////stage 1/////////////////////////////////////////
always @(posedge RCLK or negedge global_rstn or negedge local_rstn)
begin
   if (!global_rstn)
       t_r <= 8'b0;
   else if (!local_rstn) 
       t_r <= 8'b0;
   else 
       t_r <= DI;
end

////////////////////////////stage 2///////////////////////////////////////
always @(*)
begin
    case(sel)
        1'b0 : m[3:0] = t_r[3:0];
        1'b1 : m[3:0] = {t_r[2:0],up_r0[6]};
        default : m[3:0] = 4'bx;
    endcase
end

always @(*)
begin
    case(sel)
        1'b0 : m[7:4] = (OSERDES_MODE == "OSER7") ? {1'b0,t_r[6:4]} : t_r[7:4];
        1'b1 : m[7:4] = t_r[6:3];
        default : m[7:4] = 4'bx;
    endcase
end

always @(posedge OCLK or negedge global_rstn or negedge local_rstn)
begin
   if (!global_rstn)
       up_r0 <= 8'b0;
   else if (!local_rstn)
       up_r0 <= 8'b0;
   else if(upd_stage0)
       up_r0 <= m;
end

//////////////////////////stage 3/////////////////////////////////////
always @(posedge OCLK or negedge global_rstn or negedge local_rstn)
begin
   if (!global_rstn)
       up_r1 <= 8'b0;
   else if (!local_rstn)
       up_r1 <= 8'b0;
   else
   begin
        if(upd_stage1)
            up_r1 <= up_r0;
        else
        begin
            up_r1[7:6] <= 2'b0;
            up_r1[5:4] <= up_r1[7:6];
            up_r1[3:2] <= (OSERDES_MODE == "OSER4") ? 2'b0 : up_r1[5:4];
            up_r1[1:0] <= up_r1[3:2];
        end
    end
end

////////////////////parallel to serial//////////////////////////////
always @(negedge OCLK or negedge global_rstn or negedge local_rstn)
begin
   if (!global_rstn)
       f_reg <= 'b0;
   else if (!local_rstn)
       f_reg <= 'b0;
   else
       f_reg <= up_r1[1];
end

assign DO = OCLK ? up_r1[0] : f_reg;
/////////////////////////update & sel function //////////////////
always @(posedge OCLK or negedge global_rstn or negedge local_rstn)
begin
   if (!global_rstn)
        rstn_sync <= 1'b0;
   else if (!local_rstn)
        rstn_sync <= 1'b0;
    else
        rstn_sync <= 1'b1;
end

always @(posedge OCLK or negedge rstn_sync)
begin
    if (!rstn_sync)
        cnt <= 2'b0;
    else if(OSERDES_MODE == "OSER4")
        cnt[0] <= cnt[0] + 1;
    else begin
        if((OSERDES_MODE == "OSER7") && select_reg && (cnt == 2'b10))
            cnt <= 2'b0;
        else
            cnt <= cnt + 1;
    end
end

always @(posedge OCLK or negedge rstn_sync)
begin
    if (!rstn_sync)
        select_reg <= 0;
    else if(OSERDES_MODE == "OSER7")
    begin
        if((cnt == 2'b10) && select_reg)
            select_reg <= ~select_reg;
        else if((cnt == 2'b11) && (~select_reg))
            select_reg <= ~select_reg;
    end
end

always @(posedge OCLK or negedge rstn_sync)
begin
    if (!rstn_sync)
    begin
        update0_reg <= 1'b0;
        update1_reg <= 1'b0;
    end
    else
    begin
        if(OSERDES_MODE == "OSER7")
        begin
            if(select_reg) begin
                update0_reg <= (~cnt[1])&(~cnt[0]);
                update1_reg <= (~cnt[1])& cnt[0];
            end
            else begin
                update0_reg <= (~cnt[1])&cnt[0];
                update1_reg <= cnt[1]&(~cnt[0]);
            end
        end
        else if(OSERDES_MODE == "OSER4")
        begin
            update0_reg <= ~cnt[0];
        end
        else if(OSERDES_MODE == "OSER8")
        begin
            update0_reg <= (~cnt[1])&&cnt[0];
        end
    end
end

assign update0 = update0_reg;
assign update1 = update1_reg;
assign sel       = select_reg;

//synthesis translate_on

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_IGDES8.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_IGDES8 #(
parameter GRS_EN = "TRUE", //"TRUE"; "FALSE"
parameter LRS_EN = "TRUE",  //"TRUE"; "FALSE"
parameter DPI_EN = "FALSE"  //"TRUE"; "FALSE"
)(
output [7:0] Q,
output [1:0] DPI_STS,
input [1:0] DPI_CTRL,
input DPI_STS_CLR_N,
input PADI,
input DESCLK,
input RCLK,
input RST
);

//synthesis translate_off
reg PADI_POS;
reg PADI_NEG;
reg [7:0] shift_reg;
reg [7:0] capture_reg;
reg [1:0] cnt;
wire capture_en;
reg [7:0] Q_reg;
wire [7:0] PADI_D;
reg DPI_P;
reg [1:0] DPI_STS_R;
wire COMP_BEFORE;
wire COMP_AFTER;
wire COMP_BEFORE_D;
wire COMP_AFTER_D;
wire PD_BEFORE;
wire PD_AFTER;
wire DPI_BEFORE_POS_REG_T;
wire DPI_AFTER_POS_REG_T;
wire DPI_BEFORE_NEG_REG_T;
wire DPI_AFTER_NEG_REG_T;
wire AFTER_POS;
wire BEFORE_POS;
wire AFTER_NEG;
wire BEFORE_NEG;
reg DPI_N_reg;
reg DPI_BEFORE;
reg DPI_AFTER;
reg DPI_BEFORE_POS_REG;
reg DPI_BEFORE_NEG_REG;
reg DPI_AFTER_POS_REG;
reg DPI_AFTER_NEG_REG;

initial begin
PADI_POS            = 0;
PADI_NEG            = 0;
shift_reg           = 0;
capture_reg         = 0;
cnt                 = 0;
Q_reg               = 0;
DPI_P               = 0;
DPI_STS_R           = 0;
DPI_N_reg           = 0;
DPI_BEFORE          = 0;
DPI_AFTER           = 0;
DPI_BEFORE_POS_REG  = 0;
DPI_BEFORE_NEG_REG  = 0;
DPI_AFTER_POS_REG   = 0;
DPI_AFTER_NEG_REG   = 0;  
end
assign global_rstn = (GRS_EN == "TRUE") ? GRS_INST.GRSNET : 1'b1;
assign lsr_rstn = LRS_EN == "TRUE" ? (~RST) : 1'b1;


assign  #0.05 PADI_D[0] =  PADI;
assign  #0.05 PADI_D[1] =  PADI_D[0];
assign  #0.05 PADI_D[2] =  PADI_D[1];
assign  #0.05 PADI_D[3] =  PADI_D[2];
assign  #0.05 PADI_D[4] =  PADI_D[3];
assign  #0.05 PADI_D[5] =  PADI_D[4];
assign  #0.05 PADI_D[6] =  PADI_D[5];
assign  #0.05 PADI_D[7] =  PADI_D[6];

assign PADI_SAMPLE = (DPI_EN == "TRUE") ? PADI_D[3] : PADI;

always @(posedge DESCLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_P <= 0;
   else if (!lsr_rstn)
      DPI_P <= 0;
   else
      DPI_P <= PADI_SAMPLE;
end

always @(negedge DESCLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_N_reg <= 0;
   else if (!lsr_rstn)
      DPI_N_reg <= 0;
   else 
      DPI_N_reg <= PADI_SAMPLE;
end

always @(*) begin
   case (DPI_CTRL[1:0])
      2'd0:    begin DPI_BEFORE = PADI_D[2];  DPI_AFTER = PADI_D[4]; end
      2'd1:    begin DPI_BEFORE = PADI_D[1];  DPI_AFTER = PADI_D[5]; end
      2'd2:    begin DPI_BEFORE = PADI_D[0];  DPI_AFTER = PADI_D[6]; end
      default: begin DPI_BEFORE = PADI;       DPI_AFTER = PADI_D[7]; end
   endcase
end

always @(posedge DESCLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_BEFORE_POS_REG <= 0;
   else if (!lsr_rstn)
      DPI_BEFORE_POS_REG <= 0;
   else   
      DPI_BEFORE_POS_REG <= DPI_BEFORE;
end

always @(negedge DESCLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_BEFORE_NEG_REG <= 0;
   else if (!lsr_rstn)
      DPI_BEFORE_NEG_REG <= 0;
   else     
      DPI_BEFORE_NEG_REG <= DPI_BEFORE;
end


always @(posedge DESCLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_AFTER_POS_REG <= 0;
   else if (!lsr_rstn)
      DPI_AFTER_POS_REG <= 0;
   else   
      DPI_AFTER_POS_REG <= DPI_AFTER;
end


always @(negedge DESCLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_AFTER_NEG_REG <= 0;
   else if (!lsr_rstn)
      DPI_AFTER_NEG_REG <= 0;
   else     
      DPI_AFTER_NEG_REG <= DPI_AFTER;
end

assign BEFORE_POS = DPI_BEFORE_POS_REG_T ^ DPI_P;
assign DPI_BEFORE_POS_REG_T = (DPI_EN == "TRUE") ? DPI_BEFORE_POS_REG : 0;

assign AFTER_POS = DPI_AFTER_POS_REG_T ^ DPI_P;
assign DPI_AFTER_POS_REG_T = (DPI_EN == "TRUE") ? DPI_AFTER_POS_REG : 0;

assign BEFORE_NEG = DPI_BEFORE_NEG_REG_T ^ DPI_N_reg;
assign DPI_BEFORE_NEG_REG_T = (DPI_EN == "TRUE") ? DPI_BEFORE_NEG_REG : 0;

assign AFTER_NEG = DPI_AFTER_NEG_REG_T ^ DPI_N_reg;
assign DPI_AFTER_NEG_REG_T = (DPI_EN == "TRUE") ? DPI_AFTER_NEG_REG : 0;

assign COMP_BEFORE = BEFORE_POS || BEFORE_NEG;
assign COMP_AFTER = AFTER_POS || AFTER_NEG;

assign #0.1 COMP_BEFORE_D = COMP_BEFORE;
assign #0.1 COMP_AFTER_D = COMP_AFTER;

assign PD_BEFORE = COMP_BEFORE && COMP_BEFORE_D;
assign PD_AFTER = COMP_AFTER && COMP_AFTER_D;


always @(posedge DPI_STS_CLR_N or negedge global_rstn or negedge lsr_rstn or posedge PD_BEFORE) begin
   if (!global_rstn)
      DPI_STS_R[0] <= 0;
   else if (!lsr_rstn)
      DPI_STS_R[0] <= 0;
   else if (PD_BEFORE)     
      DPI_STS_R[0] <= 1'b1;
   else
      DPI_STS_R[0] <= 1'b0;
end

always @(posedge DPI_STS_CLR_N or negedge global_rstn or negedge lsr_rstn or posedge PD_AFTER) begin
   if (!global_rstn)
      DPI_STS_R[1] <= 0;
   else if (!lsr_rstn)
      DPI_STS_R[1] <= 0;
   else if (PD_AFTER)     
      DPI_STS_R[1] <= 1'b1;
   else
      DPI_STS_R[1] <= 1'b0;
end


assign DPI_STS[0] = DPI_STS_R[0];
assign DPI_STS[1] = DPI_STS_R[1];

always @(posedge DESCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      shift_reg <= 0;
   else if (!lsr_rstn)
      shift_reg <= 0;
   else
      shift_reg <= {DPI_N_reg, DPI_P, shift_reg[7:2]};

always @(posedge DESCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      cnt <= 0;
   else if (!lsr_rstn)
      cnt <= 0;
   else
      cnt <= cnt + 1;

assign capture_en = cnt == 3;

always @(posedge DESCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      capture_reg <= 0;
   else if (!lsr_rstn)
      capture_reg <= 0;
   else if (capture_en)
      capture_reg <= shift_reg;
      
always @(posedge RCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      Q_reg <= 0;
   else if (!lsr_rstn)
      Q_reg <= 0;
   else
      Q_reg <= capture_reg;      

assign Q = Q_reg;
//synthesis translate_on

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////

//P = (A0*(B0+/-C0) +/- A1*(B1 +/-C1)) +- (A2*(B2+/-C2) +/- A3*(B3+/-C3))
`timescale 1 ns / 1 ps

module INT_PREADD_MULTADDSUM #(
parameter GRS_EN      = "FALSE", //"TRUE"; "FALSE"
parameter SYNC_RST    = "FALSE", //"TRUE"; "FALSE"
parameter SIB1_EN     = "FALSE", //"TRUE"; "FALSE"
parameter SIB2_EN     = "FALSE", //"TRUE"; "FALSE"
parameter SIB3_EN     = "FALSE", //"TRUE"; "FALSE"
parameter SIC0_EN     = "FALSE", //"TRUE"; "FALSE"
parameter SIC1_EN     = "FALSE", //"TRUE"; "FALSE"
parameter SIC2_EN     = "FALSE", //"TRUE"; "FALSE"
parameter SIC3_EN     = "FALSE", //"TRUE"; "FALSE"
parameter INREG_EN    = "FALSE",  //"TRUE"; "FALSE"
parameter PREREG_EN = "FALSE",  //"TRUE"; "FALSE"
parameter PIPEREG_EN  = "FALSE",  //"TRUE"; "FALSE"
parameter OUTREG_EN   = "FALSE",   //"TRUE"; "FALSE"
parameter ADDSUB_OP01     = 0 ,
parameter ADDSUB_OP23     = 0 ,
parameter ADDSUBSUM_OP     = 0 ,
parameter DYN_OP_SEL0  = 1,
parameter DYN_OP_SEL1  = 1,
parameter DYN_OP_SEL2  = 1,
parameter ASIZE = 9,               // LEGAL ASIZE = 9, 18
parameter BSIZE = 8,               // LEGAL BSIZE = 8, 18
parameter CSIZE = BSIZE,
parameter PSIZE = ASIZE + BSIZE +2,
parameter SC_PSE_A0 = 0, //SC_PSE = 0, disable PSE,  bit width = ASIZE-1
parameter SC_PSE_A1 = 0, //SC_PSE = 0, disable PSE,  bit width = ASIZE-1
parameter SC_PSE_A2 = 0, //SC_PSE = 0, disable PSE,  bit width = ASIZE-1
parameter SC_PSE_A3 = 0, //SC_PSE = 0, disable PSE,  bit width = ASIZE-1
parameter SC_PSE_B0 = 0, //SC_PSE = 0, disable PSE,  bit width = BSIZE-1 
parameter SC_PSE_B1 = 0, //SC_PSE = 0, disable PSE,  bit width = BSIZE-1
parameter SC_PSE_B2 = 0, //SC_PSE = 0, disable PSE,  bit width = BSIZE-1
parameter SC_PSE_B3 = 0, //SC_PSE = 0, disable PSE,  bit width = BSIZE-1
parameter SC_PSE_C0 = 0, //SC_PSE = 0, disable PSE,  bit width = CSIZE-1
parameter SC_PSE_C1 = 0, //SC_PSE = 0, disable PSE,  bit width = CSIZE-1
parameter SC_PSE_C2 = 0, //SC_PSE = 0, disable PSE,  bit width = CSIZE-1
parameter SC_PSE_C3 = 0  //SC_PSE = 0, disable PSE,  bit width = CSIZE-1 
)(
input   CE,
input   RST,
input   CLK,
input   A_SIGNED01,
input   A_SIGNED23,
input   [ASIZE-1:0] A0,
input   [ASIZE-1:0] A1,
input   [ASIZE-1:0] A2,
input   [ASIZE-1:0] A3,
input   B_SIGNED01,
input   B_SIGNED23,
input   C_SIGNED01,
input   C_SIGNED23,
input   [BSIZE-1:0] B0,
input   [BSIZE-1:0] B1,
input   [BSIZE-1:0] B2,
input   [BSIZE-1:0] B3,
input   [CSIZE-1:0] C0,
input   [CSIZE-1:0] C1,
input   [CSIZE-1:0] C2,
input   [CSIZE-1:0] C3,
input   [1:0] PREADDSUB01,
input   [1:0] PREADDSUB23,
input   ADDSUB01,
input   ADDSUB23,
input   ADDSUBSUM,
output  [PSIZE:0] P
);

initial begin
    if ((ASIZE == 9 && BSIZE == 8) || (ASIZE == 18 && BSIZE == 18))
    begin 
    end
    else
        $display (" GTP_PREADD_MULTADDSUM error: illegal setting of ASZIE or BSIZE");

    if (SIB1_EN != "FALSE" || SIB2_EN != "FALSE" || SIB3_EN != "FALSE") begin
        $display("DRC error");
        $finish;
    end
    if (SIC0_EN != "FALSE" || SIC1_EN != "FALSE" || SIC2_EN != "FALSE" || SIC3_EN != "FALSE") begin
        $display("DRC error");
        $finish;
    end
end

parameter PRODUCT_SIZE = (ASIZE + BSIZE +1 )*2; 
parameter P_EXT1 = BSIZE +3;
parameter P_EXT2 = ASIZE +2;

wire [ASIZE-1:0] A0_PSE;
wire [ASIZE-1:0] A1_PSE;
wire [ASIZE-1:0] A2_PSE;
wire [ASIZE-1:0] A3_PSE;
wire [BSIZE-1:0] B0_PSE;
wire [BSIZE-1:0] B1_PSE;
wire [BSIZE-1:0] B2_PSE;
wire [BSIZE-1:0] B3_PSE;
wire [CSIZE-1:0] C0_PSE;
wire [CSIZE-1:0] C1_PSE;
wire [CSIZE-1:0] C2_PSE;
wire [CSIZE-1:0] C3_PSE;

reg  [ASIZE-1:0] P1_reg_A0;
reg  [ASIZE-1:0] P1_reg_A1;
reg  [ASIZE-1:0] P1_reg_A2;
reg  [ASIZE-1:0] P1_reg_A3;
reg  P1_reg_A_SIGNED01;
reg  P1_reg_A_SIGNED23;
reg  [BSIZE-1:0] P1_reg_B0;
reg  [BSIZE-1:0] P1_reg_B1;
reg  [BSIZE-1:0] P1_reg_B2;
reg  [BSIZE-1:0] P1_reg_B3;
reg  [CSIZE-1:0] P1_reg_C0;
reg  [CSIZE-1:0] P1_reg_C1;
reg  [CSIZE-1:0] P1_reg_C2;
reg  [CSIZE-1:0] P1_reg_C3;
reg  P1_reg_B_SIGNED01;
reg  P1_reg_B_SIGNED23;
reg  P1_reg_C_SIGNED01;
reg  P1_reg_C_SIGNED23;
reg  P1_reg_ADDSUB01;
reg  P1_reg_ADDSUB23;
reg  P1_reg_ADDSUBSUM;
reg  [1:0] P1_reg_PREADDSUB01;
reg  [1:0] P1_reg_PREADDSUB23;
wire P1_reg_ADDSUB01_comb;
wire P1_reg_ADDSUB23_comb;
wire P1_reg_ADDSUBSUM_comb;
wire [1:0] P1_reg_PREADDSUB01_comb;
wire [1:0] P1_reg_PREADDSUB23_comb;

wire [ASIZE-1:0] P1_reg_A0_comb;
wire [ASIZE-1:0] P1_reg_A1_comb;
wire [ASIZE-1:0] P1_reg_A2_comb;
wire [ASIZE-1:0] P1_reg_A3_comb;
wire P1_reg_A_SIGNED01_comb;
wire P1_reg_A_SIGNED23_comb;
wire [BSIZE-1:0] P1_reg_B0_comb;
wire [BSIZE-1:0] P1_reg_B1_comb;
wire [BSIZE-1:0] P1_reg_B2_comb;
wire [BSIZE-1:0] P1_reg_B3_comb;
wire [CSIZE-1:0] P1_reg_C0_comb;
wire [CSIZE-1:0] P1_reg_C1_comb;
wire [CSIZE-1:0] P1_reg_C2_comb;
wire [CSIZE-1:0] P1_reg_C3_comb;
wire P1_reg_B_SIGNED01_comb;
wire P1_reg_B_SIGNED23_comb;
wire P1_reg_C_SIGNED01_comb;
wire P1_reg_C_SIGNED23_comb;
reg  [PSIZE:0] P1_reg_A0_comb_ext;
reg  [PSIZE:0] P1_reg_A1_comb_ext;
reg  [PSIZE:0] P1_reg_A2_comb_ext;
reg  [PSIZE:0] P1_reg_A3_comb_ext;
reg  [PSIZE:0] P1_reg_B0_comb_ext;
reg  [PSIZE:0] P1_reg_B1_comb_ext;
reg  [PSIZE:0] P1_reg_B2_comb_ext;
reg  [PSIZE:0] P1_reg_B3_comb_ext;
reg  [PSIZE:0] P1_reg_A0_comb_ext_d;
reg  [PSIZE:0] P1_reg_A1_comb_ext_d;
reg  [PSIZE:0] P1_reg_A2_comb_ext_d;
reg  [PSIZE:0] P1_reg_A3_comb_ext_d;
reg  [PSIZE:0] P1_reg_B0_comb_ext_d;
reg  [PSIZE:0] P1_reg_B1_comb_ext_d;
reg  [PSIZE:0] P1_reg_B2_comb_ext_d;
reg  [PSIZE:0] P1_reg_B3_comb_ext_d;
wire  [PSIZE:0] P1_reg_A0_comb_ext_d_sel;
wire  [PSIZE:0] P1_reg_A1_comb_ext_d_sel;
wire  [PSIZE:0] P1_reg_A2_comb_ext_d_sel;
wire  [PSIZE:0] P1_reg_A3_comb_ext_d_sel;
wire  [PSIZE:0] P1_reg_B0_comb_ext_d_sel;
wire  [PSIZE:0] P1_reg_B1_comb_ext_d_sel;
wire  [PSIZE:0] P1_reg_B2_comb_ext_d_sel;
wire  [PSIZE:0] P1_reg_B3_comb_ext_d_sel;
wire [PRODUCT_SIZE-1:0] PRODUCT_0;
wire [PRODUCT_SIZE-1:0] PRODUCT_1;
wire [PRODUCT_SIZE-1:0] PRODUCT_2;
wire [PRODUCT_SIZE-1:0] PRODUCT_3;
wire  PRODUCT0_signed;
wire  PRODUCT1_signed;
wire  PRODUCT2_signed;
wire  PRODUCT3_signed;

reg  [PSIZE:0] P2_reg_PRODUCT_0;
reg  [PSIZE:0] P2_reg_PRODUCT_1;
reg  [PSIZE:0] P2_reg_PRODUCT_2;
reg  [PSIZE:0] P2_reg_PRODUCT_3;
reg  P2_reg_ADDSUB01;
wire P2_reg_ADDSUB01_comb;
reg  P2_reg_ADDSUB23;
wire P2_reg_ADDSUB23_comb;
reg  P2_reg_ADDSUBSUM;
wire P2_reg_ADDSUBSUM_comb;
wire [PSIZE:0] P2_reg_PRODUCT_0_comb;
wire [PSIZE:0] P2_reg_PRODUCT_1_comb;
wire [PSIZE:0] P2_reg_PRODUCT_2_comb;
wire [PSIZE:0] P2_reg_PRODUCT_3_comb;
wire [PSIZE:0] sum01;
wire [PSIZE:0] sum23;
wire [PSIZE:0] sum;
reg  [PSIZE:0] P_reg;
wire [ASIZE-1:0]  A1_comb;
wire [ASIZE-1:0]  A2_comb;
wire [ASIZE-1:0]  A3_comb;
wire [BSIZE-1:0]  B1_comb;
wire [BSIZE-1:0]  B2_comb;
wire [BSIZE-1:0]  B3_comb;
wire [CSIZE-1:0]  C0_comb;
wire [CSIZE-1:0]  C1_comb;
wire [CSIZE-1:0]  C2_comb;
wire [CSIZE-1:0]  C3_comb;
wire        C_SIGNED_comb01;
wire        C_SIGNED_comb23;


wire [BSIZE:0] P1_preadd_BC0;
wire       P1_preadd_BC0_SIGNED;
wire [BSIZE:0] P1_preadd_BC1;
wire       P1_preadd_BC1_SIGNED;
wire [BSIZE:0] P1_preadd_BC2;
wire       P1_preadd_BC2_SIGNED;
wire [BSIZE:0] P1_preadd_BC3;
wire       P1_preadd_BC3_SIGNED;

INT_PSE #(.ASIZE(ASIZE),.SC_PSE(SC_PSE_A0)) U1_PSE (.A(A0), .SIGN(A_SIGNED01), .A_PSE(A0_PSE));
INT_PSE #(.ASIZE(ASIZE),.SC_PSE(SC_PSE_A1)) U2_PSE (.A(A1), .SIGN(A_SIGNED01), .A_PSE(A1_PSE));
INT_PSE #(.ASIZE(ASIZE),.SC_PSE(SC_PSE_A2)) U3_PSE (.A(A2), .SIGN(A_SIGNED23), .A_PSE(A2_PSE));
INT_PSE #(.ASIZE(ASIZE),.SC_PSE(SC_PSE_A3)) U4_PSE (.A(A3), .SIGN(A_SIGNED23), .A_PSE(A3_PSE));

INT_PSE #(.ASIZE(BSIZE),.SC_PSE(SC_PSE_B0)) U5_PSE (.A(B0), .SIGN(B_SIGNED01), .A_PSE(B0_PSE));
INT_PSE #(.ASIZE(BSIZE),.SC_PSE(SC_PSE_B1)) U6_PSE (.A(B1), .SIGN(B_SIGNED01), .A_PSE(B1_PSE));
INT_PSE #(.ASIZE(BSIZE),.SC_PSE(SC_PSE_B2)) U7_PSE (.A(B2), .SIGN(B_SIGNED23), .A_PSE(B2_PSE));
INT_PSE #(.ASIZE(BSIZE),.SC_PSE(SC_PSE_B3)) U8_PSE (.A(B3), .SIGN(B_SIGNED23), .A_PSE(B3_PSE));

INT_PSE #(.ASIZE(CSIZE),.SC_PSE(SC_PSE_C0)) U9_PSE (.A(C0), .SIGN(C_SIGNED01), .A_PSE(C0_PSE));
INT_PSE #(.ASIZE(CSIZE),.SC_PSE(SC_PSE_C1)) U10_PSE(.A(C1), .SIGN(C_SIGNED01), .A_PSE(C1_PSE));
INT_PSE #(.ASIZE(CSIZE),.SC_PSE(SC_PSE_C2)) U11_PSE(.A(C2), .SIGN(C_SIGNED23), .A_PSE(C2_PSE));
INT_PSE #(.ASIZE(CSIZE),.SC_PSE(SC_PSE_C3)) U12_PSE(.A(C3), .SIGN(C_SIGNED23), .A_PSE(C3_PSE));

wire global_rstn, RST_sync, RST_async, rst_asyncomb;

assign global_rstn = GRS_EN == "TRUE" ? GRS_INST.GRSNET : 1'b1;
assign RST_sync = (SYNC_RST == "TRUE") ? RST : 1'b0;
assign RST_async = (SYNC_RST == "FALSE") ? RST : 1'b0;
assign rst_asyncomb = RST_async | (~global_rstn);

assign A1_comb = A1_PSE;
assign B1_comb = (SIB1_EN == "TRUE") ?  P1_reg_B0_comb :  B1_PSE;
assign C0_comb = (SIC0_EN == "TRUE") ?  P1_reg_B0_comb :  C0_PSE;
assign C1_comb = (SIC1_EN == "TRUE") ?  P1_reg_B1_comb :  C1_PSE;
assign A2_comb = A2_PSE;
assign B2_comb = (SIB2_EN == "TRUE") ?  P1_reg_B1_comb :  B2_PSE;
assign C2_comb = (SIC2_EN == "TRUE") ?  P1_reg_B1_comb :  C2_PSE;
assign A3_comb = A3_PSE;
assign B3_comb = (SIB3_EN == "TRUE") ?  P1_reg_B2_comb :  B3_PSE;
assign C3_comb = (SIC3_EN == "TRUE") ?  P1_reg_B2_comb :  C3_PSE;
assign C_SIGNED_comb01 = (SIC0_EN == "TRUE") ?  P1_reg_B_SIGNED01_comb :  C_SIGNED01 ;
assign C_SIGNED_comb23 = (SIC2_EN == "TRUE") ?  P1_reg_B_SIGNED23_comb :  C_SIGNED23 ;

initial begin
      P1_reg_A0        = 0;
      P1_reg_A1        = 0;
      P1_reg_A2        = 0;
      P1_reg_A3        = 0;      
      P1_reg_A_SIGNED01 = 0;
      P1_reg_A_SIGNED23 = 0;
      P1_reg_B0        = 0;
      P1_reg_B1        = 0;
      P1_reg_B2        = 0;
      P1_reg_B3        = 0;      
      P1_reg_C0        = 0;
      P1_reg_C1        = 0;
      P1_reg_C2        = 0;
      P1_reg_C3        = 0;      
      P1_reg_B_SIGNED01 = 0;
      P1_reg_B_SIGNED23 = 0;
      P1_reg_C_SIGNED01 = 0;
      P1_reg_C_SIGNED23 = 0;
      P1_reg_ADDSUB01 = 0;
      P1_reg_ADDSUB23 = 0;
      P1_reg_ADDSUBSUM = 0;      
      P1_reg_PREADDSUB01 = 0;
      P1_reg_PREADDSUB23 = 0;
         P2_reg_PRODUCT_0 = 0;
         P2_reg_PRODUCT_1 = 0;
         P2_reg_PRODUCT_2 = 0;
         P2_reg_PRODUCT_3 = 0;         
         P2_reg_ADDSUB01 = 0;
         P2_reg_ADDSUB23 = 0;
          P2_reg_ADDSUBSUM =0 ;
      P_reg    = 0;             
end
always @(posedge CLK or posedge rst_asyncomb)
   if (rst_asyncomb || RST_sync) begin
      P1_reg_A0        <= 0;
      P1_reg_A1        <= 0;
      P1_reg_A2        <= 0;
      P1_reg_A3        <= 0;      
      P1_reg_A_SIGNED01 <= 0;
      P1_reg_A_SIGNED23 <= 0;
      P1_reg_B0        <= 0;
      P1_reg_B1        <= 0;
      P1_reg_B2        <= 0;
      P1_reg_B3        <= 0;      
      P1_reg_C0        <= 0;
      P1_reg_C1        <= 0;
      P1_reg_C2        <= 0;
      P1_reg_C3        <= 0;      
      P1_reg_B_SIGNED01 <= 0;
      P1_reg_B_SIGNED23 <= 0;
      P1_reg_C_SIGNED01 <= 0;
      P1_reg_C_SIGNED23 <= 0;
      P1_reg_ADDSUB01 <= 0;
      P1_reg_ADDSUB23 <= 0;
      P1_reg_ADDSUBSUM <= 0;      
      P1_reg_PREADDSUB01 <= 0;
      P1_reg_PREADDSUB23 <= 0;
   end
      else if (CE) begin
         P1_reg_A0        <= A0;
         P1_reg_A1        <= A1_comb;
         P1_reg_A2        <= A2_comb;
         P1_reg_A3        <= A3_comb;
         P1_reg_A_SIGNED01 <= A_SIGNED01;
         P1_reg_A_SIGNED23 <= A_SIGNED23;
         P1_reg_B0        <= B0;
         P1_reg_B1        <= B1_comb;
         P1_reg_B2        <= B2_comb;         
         P1_reg_B3        <= B3_comb;         
         P1_reg_C0        <= C0_comb;
         P1_reg_C1        <= C1_comb;
         P1_reg_C2        <= C2_comb;
         P1_reg_C3        <= C3_comb;      
         P1_reg_B_SIGNED01 <= B_SIGNED01;
         P1_reg_B_SIGNED23 <= B_SIGNED23;
         P1_reg_C_SIGNED01 <= C_SIGNED_comb01;
         P1_reg_C_SIGNED23 <= C_SIGNED_comb23;
         P1_reg_ADDSUB01 <= (DYN_OP_SEL0 == 1'b1)? ADDSUB01 : ADDSUB_OP01;
         P1_reg_ADDSUB23 <= (DYN_OP_SEL1 == 1'b1)? ADDSUB23 : ADDSUB_OP23;
     P1_reg_ADDSUBSUM <=(DYN_OP_SEL2 == 1'b1)? ADDSUBSUM:ADDSUBSUM_OP;
         P1_reg_PREADDSUB01 <= PREADDSUB01;
         P1_reg_PREADDSUB23 <= PREADDSUB23;
   end
   
assign P1_reg_A0_comb        = (INREG_EN == "TRUE") ? P1_reg_A0        : A0_PSE;
assign P1_reg_A1_comb        = (INREG_EN == "TRUE") ? P1_reg_A1        : A1_comb;
assign P1_reg_A2_comb        = (INREG_EN == "TRUE") ? P1_reg_A2        : A2_comb;
assign P1_reg_A3_comb        = (INREG_EN == "TRUE") ? P1_reg_A3        : A3_comb;
assign P1_reg_A_SIGNED01_comb = (INREG_EN == "TRUE") ? P1_reg_A_SIGNED01 : A_SIGNED01;
assign P1_reg_A_SIGNED23_comb = (INREG_EN == "TRUE") ? P1_reg_A_SIGNED23 : A_SIGNED23;
assign P1_reg_B0_comb        = (INREG_EN == "TRUE") ? P1_reg_B0        : B0_PSE;
assign P1_reg_B1_comb        = (INREG_EN == "TRUE") ? P1_reg_B1        : B1_comb;
assign P1_reg_B2_comb        = (INREG_EN == "TRUE") ? P1_reg_B2        : B2_comb;
assign P1_reg_B3_comb        = (INREG_EN == "TRUE") ? P1_reg_B3        : B3_comb;
assign P1_reg_C0_comb        = (INREG_EN == "TRUE") ? P1_reg_C0        : C0_comb;
assign P1_reg_C1_comb        = (INREG_EN == "TRUE") ? P1_reg_C1        : C1_comb;
assign P1_reg_C2_comb        = (INREG_EN == "TRUE") ? P1_reg_C2        : C2_comb;
assign P1_reg_C3_comb        = (INREG_EN == "TRUE") ? P1_reg_C3        : C3_comb;
assign P1_reg_B_SIGNED01_comb = (INREG_EN == "TRUE") ? P1_reg_B_SIGNED01 : B_SIGNED01;
assign P1_reg_B_SIGNED23_comb = (INREG_EN == "TRUE") ? P1_reg_B_SIGNED23 : B_SIGNED23;
assign P1_reg_C_SIGNED01_comb = (INREG_EN == "TRUE") ? P1_reg_C_SIGNED01 : C_SIGNED01;
assign P1_reg_C_SIGNED23_comb = (INREG_EN == "TRUE") ? P1_reg_C_SIGNED23 : C_SIGNED23;
assign P1_reg_ADDSUB01_comb = (INREG_EN == "TRUE") ? P1_reg_ADDSUB01 :(DYN_OP_SEL0 == 1'b1)? ADDSUB01 : ADDSUB_OP01;
assign P1_reg_ADDSUB23_comb = (INREG_EN == "TRUE") ? P1_reg_ADDSUB23 :(DYN_OP_SEL1 == 1'b1)? ADDSUB23 : ADDSUB_OP23;
assign P1_reg_ADDSUBSUM_comb = (INREG_EN == "TRUE") ? P1_reg_ADDSUBSUM : (DYN_OP_SEL2 == 1'b1)? ADDSUBSUM:ADDSUBSUM_OP;
assign P1_reg_PREADDSUB01_comb = (INREG_EN == "TRUE") ? P1_reg_PREADDSUB01 : PREADDSUB01;
assign P1_reg_PREADDSUB23_comb = (INREG_EN == "TRUE") ? P1_reg_PREADDSUB23 : PREADDSUB23;

assign P1_preadd_BC0 = (P1_reg_PREADDSUB01_comb[0] == 1'b0)? {P1_reg_B_SIGNED01_comb&P1_reg_B0_comb[BSIZE-1],P1_reg_B0_comb} + {P1_reg_C_SIGNED01_comb&P1_reg_C0_comb[CSIZE-1],P1_reg_C0_comb} : {P1_reg_B_SIGNED01_comb&P1_reg_B0_comb[BSIZE-1],P1_reg_B0_comb} - {P1_reg_C_SIGNED01_comb&P1_reg_C0_comb[CSIZE-1],P1_reg_C0_comb} ;
assign P1_preadd_BC0_SIGNED = P1_reg_B_SIGNED01_comb | P1_reg_C_SIGNED01_comb;
assign P1_preadd_BC1 = (P1_reg_PREADDSUB01_comb[1] == 1'b0)?{P1_reg_B_SIGNED01_comb&P1_reg_B1_comb[BSIZE-1],P1_reg_B1_comb}+ {P1_reg_C_SIGNED01_comb&P1_reg_C1_comb[CSIZE-1],P1_reg_C1_comb}:{P1_reg_B_SIGNED01_comb&P1_reg_B1_comb[BSIZE-1],P1_reg_B1_comb} - {P1_reg_C_SIGNED01_comb&P1_reg_C1_comb[CSIZE-1],P1_reg_C1_comb} ;
assign P1_preadd_BC1_SIGNED = P1_reg_B_SIGNED01_comb | P1_reg_C_SIGNED01_comb;


assign P1_preadd_BC2 = (P1_reg_PREADDSUB23_comb[0] == 1'b0)? {P1_reg_B_SIGNED23_comb&P1_reg_B2_comb[BSIZE-1],P1_reg_B2_comb} + {P1_reg_C_SIGNED23_comb&P1_reg_C2_comb[CSIZE-1],P1_reg_C2_comb} : {P1_reg_B_SIGNED23_comb&P1_reg_B2_comb[BSIZE-1],P1_reg_B2_comb} - {P1_reg_C_SIGNED23_comb&P1_reg_C2_comb[CSIZE-1],P1_reg_C2_comb} ;
assign P1_preadd_BC2_SIGNED = P1_reg_B_SIGNED23_comb | P1_reg_C_SIGNED23_comb;
assign P1_preadd_BC3 = (P1_reg_PREADDSUB23_comb[1] == 1'b0)?{P1_reg_B_SIGNED23_comb&P1_reg_B3_comb[BSIZE-1],P1_reg_B3_comb}+ {P1_reg_C_SIGNED23_comb&P1_reg_C3_comb[CSIZE-1],P1_reg_C3_comb}:{P1_reg_B_SIGNED23_comb&P1_reg_B3_comb[BSIZE-1],P1_reg_B3_comb} - {P1_reg_C_SIGNED23_comb&P1_reg_C3_comb[CSIZE-1],P1_reg_C3_comb} ;
assign P1_preadd_BC3_SIGNED = P1_reg_B_SIGNED23_comb | P1_reg_C_SIGNED23_comb;

reg preadd_over_flag0;
always @(*)begin
  if(P1_reg_PREADDSUB01_comb[0]==1'b0)begin
    if((P1_reg_B_SIGNED01_comb==1'b1 && P1_reg_B0_comb[BSIZE-1]==1'b0 && P1_reg_C_SIGNED01_comb==1'b0 && P1_preadd_BC0[BSIZE]==1'b1) || (P1_reg_B_SIGNED01_comb==1'b0 && P1_reg_C_SIGNED01_comb==1'b1 && P1_reg_C0_comb[CSIZE-1]==1'b0 && P1_preadd_BC0[BSIZE]==1'b1))begin
      preadd_over_flag0 = 1'b1;
    end
    else begin
      preadd_over_flag0 = 1'b0;
    end
  end
  else if(P1_reg_PREADDSUB01_comb[0]==1'b1)begin
    if((P1_reg_B_SIGNED01_comb==1'b1 && P1_reg_B0_comb[BSIZE-1]==1'b1 && P1_reg_C_SIGNED01_comb==1'b0 && P1_preadd_BC0[BSIZE]==1'b0) || (P1_reg_B_SIGNED01_comb==1'b0 && P1_reg_C_SIGNED01_comb==1'b1 && P1_reg_C0_comb[CSIZE-1]==1'b1 && P1_preadd_BC0[BSIZE]==1'b1) || (P1_reg_B_SIGNED01_comb ==1'b0 && P1_reg_C_SIGNED01_comb==1'b0 && (P1_reg_B0_comb<P1_reg_C0_comb)))begin
      preadd_over_flag0 = 1'b1;
    end
    else begin
      preadd_over_flag0 = 1'b0;
    end
  end
end

reg preadd_over_flag1;
always @(*)begin
  if(P1_reg_PREADDSUB01_comb[1]==1'b0)begin
    if((P1_reg_B_SIGNED01_comb==1'b1 && P1_reg_B1_comb[BSIZE-1]==1'b0 && P1_reg_C_SIGNED01_comb==1'b0 && P1_preadd_BC1[BSIZE]==1'b1) || (P1_reg_B_SIGNED01_comb==1'b0 && P1_reg_C_SIGNED01_comb==1'b1 && P1_reg_C1_comb[CSIZE-1]==1'b0 && P1_preadd_BC1[BSIZE]==1'b1))begin
      preadd_over_flag1 = 1'b1;
    end
    else begin
      preadd_over_flag1 = 1'b0;
    end
  end
  else if(P1_reg_PREADDSUB01_comb[1]==1'b1)begin
    if((P1_reg_B_SIGNED01_comb==1'b1 && P1_reg_B1_comb[BSIZE-1]==1'b1 && P1_reg_C_SIGNED01_comb==1'b0 && P1_preadd_BC1[BSIZE]==1'b0) || (P1_reg_B_SIGNED01_comb==1'b0 && P1_reg_C_SIGNED01_comb==1'b1 && P1_reg_C1_comb[CSIZE-1]==1'b1 && P1_preadd_BC1[BSIZE]==1'b1) || (P1_reg_B_SIGNED01_comb ==1'b0 && P1_reg_C_SIGNED01_comb==1'b0 && (P1_reg_B1_comb<P1_reg_C1_comb)))begin
      preadd_over_flag1 = 1'b1;
    end
    else begin
      preadd_over_flag1 = 1'b0;
    end
  end
end

reg preadd_over_flag2;
always @(*)begin
  if(P1_reg_PREADDSUB23_comb[0]==1'b0)begin
    if((P1_reg_B_SIGNED23_comb==1'b1 && P1_reg_B2_comb[BSIZE-1]==1'b0 && P1_reg_C_SIGNED23_comb==1'b0 && P1_preadd_BC2[BSIZE]==1'b1) || (P1_reg_B_SIGNED23_comb==1'b0 && P1_reg_C_SIGNED23_comb==1'b1 && P1_reg_C2_comb[CSIZE-1]==1'b0 && P1_preadd_BC2[BSIZE]==1'b1))begin
      preadd_over_flag2 = 1'b1;
    end
    else begin
      preadd_over_flag2 = 1'b0;
    end
  end
  else if(P1_reg_PREADDSUB23_comb[0]==1'b1)begin
    if((P1_reg_B_SIGNED23_comb==1'b1 && P1_reg_B2_comb[BSIZE-1]==1'b1 && P1_reg_C_SIGNED23_comb==1'b0 && P1_preadd_BC2[BSIZE]==1'b0) || (P1_reg_B_SIGNED23_comb==1'b0 && P1_reg_C_SIGNED23_comb==1'b1 && P1_reg_C2_comb[CSIZE-1]==1'b1 && P1_preadd_BC2[BSIZE]==1'b1) || (P1_reg_B_SIGNED23_comb ==1'b0 && P1_reg_C_SIGNED23_comb==1'b0 && (P1_reg_B2_comb<P1_reg_C2_comb)))begin
      preadd_over_flag2 = 1'b1;
    end
    else begin
      preadd_over_flag2 = 1'b0;
    end
  end
end

reg preadd_over_flag3;
always @(*)begin
  if(P1_reg_PREADDSUB23_comb[1]==1'b0)begin
    if((P1_reg_B_SIGNED23_comb==1'b1 && P1_reg_B3_comb[BSIZE-1]==1'b0 && P1_reg_C_SIGNED23_comb==1'b0 && P1_preadd_BC3[BSIZE]==1'b1) || (P1_reg_B_SIGNED23_comb==1'b0 && P1_reg_C_SIGNED23_comb==1'b1 && P1_reg_C3_comb[CSIZE-1]==1'b0 && P1_preadd_BC3[BSIZE]==1'b1))begin
      preadd_over_flag3 = 1'b1;
    end
    else begin
      preadd_over_flag3 = 1'b0;
    end
  end
  else if(P1_reg_PREADDSUB23_comb[1]==1'b1)begin
    if((P1_reg_B_SIGNED23_comb==1'b1 && P1_reg_B3_comb[BSIZE-1]==1'b1 && P1_reg_C_SIGNED23_comb==1'b0 && P1_preadd_BC3[BSIZE]==1'b0) || (P1_reg_B_SIGNED23_comb==1'b0 && P1_reg_C_SIGNED23_comb==1'b1 && P1_reg_C3_comb[CSIZE-1]==1'b1 && P1_preadd_BC3[BSIZE]==1'b1) || (P1_reg_B_SIGNED23_comb ==1'b0 && P1_reg_C_SIGNED23_comb==1'b0 && (P1_reg_B3_comb<P1_reg_C3_comb)))begin
      preadd_over_flag3 = 1'b1;
    end
    else begin
      preadd_over_flag3 = 1'b0;
    end
  end
end

always @(preadd_over_flag0 or preadd_over_flag1 or preadd_over_flag2 or preadd_over_flag3) begin
    if (preadd_over_flag0==1 || preadd_over_flag1==1 || preadd_over_flag2==1 || preadd_over_flag3==1)
    $display("Error: PREADD result is overflow!");
end

always @(*) begin
   if (P1_reg_A_SIGNED01_comb) begin
      P1_reg_A0_comb_ext = {{P_EXT1{P1_reg_A0_comb[ASIZE-1]}}, P1_reg_A0_comb};
      P1_reg_A1_comb_ext = {{P_EXT1{P1_reg_A1_comb[ASIZE-1]}}, P1_reg_A1_comb};
   end
   else begin
      P1_reg_A0_comb_ext = {{P_EXT1{1'd0}}, P1_reg_A0_comb};
      P1_reg_A1_comb_ext = {{P_EXT1{1'd0}}, P1_reg_A1_comb};
   end
end

always @(*) begin
   if (P1_reg_A_SIGNED23_comb) begin
      P1_reg_A2_comb_ext = {{P_EXT1{P1_reg_A2_comb[ASIZE-1]}}, P1_reg_A2_comb};
      P1_reg_A3_comb_ext = {{P_EXT1{P1_reg_A3_comb[ASIZE-1]}}, P1_reg_A3_comb};
   end
   else begin
      P1_reg_A2_comb_ext = {{P_EXT1{1'd0}}, P1_reg_A2_comb};
      P1_reg_A3_comb_ext = {{P_EXT1{1'd0}}, P1_reg_A3_comb};
   end
end

always @(*) begin
   if (P1_preadd_BC0_SIGNED) begin
      P1_reg_B0_comb_ext = {{P_EXT2{P1_preadd_BC0[BSIZE]}}, P1_preadd_BC0};
      P1_reg_B1_comb_ext = {{P_EXT2{P1_preadd_BC1[BSIZE]}}, P1_preadd_BC1};
   end
   else begin
      P1_reg_B0_comb_ext = {{P_EXT2{1'd0}}, P1_preadd_BC0};
      P1_reg_B1_comb_ext = {{P_EXT2{1'd0}}, P1_preadd_BC1};
   end
end
always @(*) begin
   if (P1_preadd_BC2_SIGNED) begin
      P1_reg_B2_comb_ext = {{P_EXT2{P1_preadd_BC2[BSIZE]}}, P1_preadd_BC2};
      P1_reg_B3_comb_ext = {{P_EXT2{P1_preadd_BC3[BSIZE]}}, P1_preadd_BC3};
   end
   else begin
      P1_reg_B2_comb_ext = {{P_EXT2{1'd0}}, P1_preadd_BC2};
      P1_reg_B3_comb_ext = {{P_EXT2{1'd0}}, P1_preadd_BC3};
   end
end

always @(posedge CLK or posedge rst_asyncomb)
   if (rst_asyncomb || RST_sync) begin
          P1_reg_A0_comb_ext_d <= 0;
          P1_reg_A1_comb_ext_d <= 0;
          P1_reg_A2_comb_ext_d <= 0;
          P1_reg_A3_comb_ext_d <= 0;
          P1_reg_B0_comb_ext_d <= 0;
          P1_reg_B1_comb_ext_d <= 0;
          P1_reg_B2_comb_ext_d <= 0;
          P1_reg_B3_comb_ext_d <= 0;
   end
         else if (CE) begin
          P1_reg_A0_comb_ext_d <=P1_reg_A0_comb_ext;
          P1_reg_A1_comb_ext_d <=P1_reg_A1_comb_ext;
          P1_reg_A2_comb_ext_d <=P1_reg_A2_comb_ext;
          P1_reg_A3_comb_ext_d <=P1_reg_A3_comb_ext;
          P1_reg_B0_comb_ext_d <=P1_reg_B0_comb_ext;
          P1_reg_B1_comb_ext_d <=P1_reg_B1_comb_ext;
          P1_reg_B2_comb_ext_d <=P1_reg_B2_comb_ext;
          P1_reg_B3_comb_ext_d <=P1_reg_B3_comb_ext;
   end
         
   
assign P1_reg_A0_comb_ext_d_sel =  (PREREG_EN == "TRUE")? P1_reg_A0_comb_ext_d:P1_reg_A0_comb_ext; 
assign P1_reg_A1_comb_ext_d_sel =  (PREREG_EN == "TRUE")? P1_reg_A1_comb_ext_d:P1_reg_A1_comb_ext;
assign P1_reg_A2_comb_ext_d_sel =  (PREREG_EN == "TRUE")? P1_reg_A2_comb_ext_d:P1_reg_A2_comb_ext;
assign P1_reg_A3_comb_ext_d_sel =  (PREREG_EN == "TRUE")? P1_reg_A3_comb_ext_d:P1_reg_A3_comb_ext;
assign P1_reg_B0_comb_ext_d_sel =  (PREREG_EN == "TRUE")? P1_reg_B0_comb_ext_d:P1_reg_B0_comb_ext;
assign P1_reg_B1_comb_ext_d_sel =  (PREREG_EN == "TRUE")? P1_reg_B1_comb_ext_d:P1_reg_B1_comb_ext;
assign P1_reg_B2_comb_ext_d_sel =  (PREREG_EN == "TRUE")? P1_reg_B2_comb_ext_d:P1_reg_B2_comb_ext;
assign P1_reg_B3_comb_ext_d_sel =  (PREREG_EN == "TRUE")? P1_reg_B3_comb_ext_d:P1_reg_B3_comb_ext;

assign PRODUCT_0 = P1_reg_A0_comb_ext_d_sel * P1_reg_B0_comb_ext_d_sel;
assign PRODUCT_1 = P1_reg_A1_comb_ext_d_sel * P1_reg_B1_comb_ext_d_sel;
assign PRODUCT_2 = P1_reg_A2_comb_ext_d_sel * P1_reg_B2_comb_ext_d_sel;
assign PRODUCT_3 = P1_reg_A3_comb_ext_d_sel * P1_reg_B3_comb_ext_d_sel;
assign PRODUCT0_signed = P1_reg_A_SIGNED01_comb | P1_preadd_BC0_SIGNED;
assign PRODUCT1_signed = P1_reg_A_SIGNED01_comb | P1_preadd_BC0_SIGNED;
assign PRODUCT2_signed = P1_reg_A_SIGNED23_comb | P1_preadd_BC2_SIGNED;
assign PRODUCT3_signed = P1_reg_A_SIGNED23_comb | P1_preadd_BC2_SIGNED;


always @(posedge CLK or posedge rst_asyncomb)
   if (rst_asyncomb || RST_sync) begin
         P2_reg_PRODUCT_0 <= 0;
         P2_reg_PRODUCT_1 <= 0;
         P2_reg_PRODUCT_2 <= 0;
         P2_reg_PRODUCT_3 <= 0;         
         P2_reg_ADDSUB01 <= 0;
         P2_reg_ADDSUB23 <= 0;
          P2_reg_ADDSUBSUM <=0 ;
   end
         else if (CE) begin
            P2_reg_PRODUCT_0 <= PRODUCT_0;
            P2_reg_PRODUCT_1 <= PRODUCT_1;
            P2_reg_PRODUCT_2 <= PRODUCT_2;
            P2_reg_PRODUCT_3 <= PRODUCT_3;          
            P2_reg_ADDSUB01 <= P1_reg_ADDSUB01_comb;
            P2_reg_ADDSUB23 <= P1_reg_ADDSUB23_comb;
            P2_reg_ADDSUBSUM <=P1_reg_ADDSUBSUM_comb ;
   end


assign P2_reg_PRODUCT_0_comb = (PIPEREG_EN == "TRUE") ? P2_reg_PRODUCT_0 : PRODUCT_0;
assign P2_reg_PRODUCT_1_comb = (PIPEREG_EN == "TRUE") ? P2_reg_PRODUCT_1 : PRODUCT_1;
assign P2_reg_PRODUCT_2_comb = (PIPEREG_EN == "TRUE") ? P2_reg_PRODUCT_2 : PRODUCT_2;
assign P2_reg_PRODUCT_3_comb = (PIPEREG_EN == "TRUE") ? P2_reg_PRODUCT_3 : PRODUCT_3;   
assign P2_reg_ADDSUB01_comb = (PIPEREG_EN == "TRUE") ? P2_reg_ADDSUB01 : P1_reg_ADDSUB01_comb;
assign P2_reg_ADDSUB23_comb = (PIPEREG_EN == "TRUE") ? P2_reg_ADDSUB23 : P1_reg_ADDSUB23_comb;
assign P2_reg_ADDSUBSUM_comb = (PIPEREG_EN == "TRUE") ? P2_reg_ADDSUBSUM : P1_reg_ADDSUBSUM_comb;

assign sum01 = (P2_reg_ADDSUB01_comb == 0) ? (P2_reg_PRODUCT_0_comb + P2_reg_PRODUCT_1_comb) : 
                                       (P2_reg_PRODUCT_0_comb - P2_reg_PRODUCT_1_comb);
assign sum23 = (P2_reg_ADDSUB23_comb == 0) ? (P2_reg_PRODUCT_2_comb + P2_reg_PRODUCT_3_comb) : 
                                       (P2_reg_PRODUCT_2_comb - P2_reg_PRODUCT_3_comb);                                       
assign sum =   (P2_reg_ADDSUBSUM_comb == 0)? (sum01 + sum23) : (sum01 - sum23);

always @(posedge CLK or posedge rst_asyncomb)
   if (rst_asyncomb || RST_sync) begin
         P_reg    <= 0;
   end
         else if (CE) begin
         P_reg    <= sum;             
   end
   
assign P = (OUTREG_EN == "TRUE") ? P_reg : sum;

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module INT_FLAG #(
    parameter GRS_EN    = "FALSE",  //"TRUE"; "FALSE"
    parameter SYNC_RST  = "FALSE",  //"TRUE"; "FALSE"
    parameter PSIZE     = 64,       //APM calculate product size
    parameter PATSIZE   = 64,       //compare pattern size
    parameter MASKPATSIZE = 64,     //pattern mask size
    parameter OUTREG_EN = "TRUE"
) (
    input   CE,
    input   RST,
    input   CLK,
    input [PSIZE-1:0] P,            //APM calculate product
    input [PATSIZE-1:0] PATTERN,    //compare pattern
    input [MASKPATSIZE-1:0] MASKPAT, //pattern mask
    input [PSIZE-1:0] OVERFLOW_MASK, //pattern mask
    input [PSIZE-1:0] R,

    output  eqz,
    output  eqzm,
    output  eqom,
    output  eqpat,
    output  eqpatn
);

initial begin
    if ((GRS_EN != "TRUE") && (GRS_EN != "FALSE")) begin
        $display("GRS_EN error");
        $finish;
    end
    if ((SYNC_RST != "TRUE") && (SYNC_RST != "FALSE")) begin
        $display("SYNC_RST error");
        $finish;
    end
    if ((OUTREG_EN != "TRUE") && (OUTREG_EN != "FALSE")) begin
        $display("OUTREG_EN error");
        $finish;
    end
end

wire eqzero;
wire eqzero_mask;
wire eqone_mask;
wire eqpattern;
wire eqpattern_n;

wire global_rstn, RST_sync, RST_async, rst_asyncomb;
assign global_rstn = GRS_EN == "TRUE" ? GRS_INST.GRSNET : 1'b1;
assign RST_sync = (SYNC_RST == "TRUE") ? RST : 1'b0;
assign RST_async = (SYNC_RST == "FALSE") ? RST : 1'b0;
assign rst_asyncomb = RST_async | (~global_rstn);

assign eqzero = (R == 0);
assign eqone_mask  = &( R | OVERFLOW_MASK);
assign eqzero_mask = &(~R | OVERFLOW_MASK);
assign eqpattern   = &((R[PATSIZE-1:0] ~^ PATTERN) | MASKPAT);
assign eqpattern_n = &((R[PATSIZE-1:0] ^ PATTERN)  | MASKPAT);

INT_REG #(.SIZE(5)) UFLAG (
    .Q({eqpatn, eqpat, eqom, eqzm, eqz}),
    .BYPASS((OUTREG_EN == "TRUE") ? 1'b0 : 1'b1),
    .D({eqpattern_n, eqpattern, eqone_mask, eqzero_mask, eqzero}),
    .CLK(CLK), .CE(CE), .ARST(rst_asyncomb), .SRST(RST_sync));

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2019 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_ROM32X2.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_ROM32X2
#(
    parameter [31:0] INIT_0 = 32'h00000000,
    parameter [31:0] INIT_1 = 32'h00000000
) (
    output [1:0] Z,
    input        I0,
    input        I1,
    input        I2,
    input        I3,
    input        I4
);
//synthesis translate_off
   reg [31:0] mem [1:0];
   wire [4:0] addr;

   initial begin
       mem[0] = INIT_0;
       mem[1] = INIT_1;
   end

   assign addr = {I4, I3, I2, I1, I0};
   //assign Z = mem[addr];
   assign Z[0] = INIT_0[addr];
   assign Z[1] = INIT_1[addr];
//synthesis translate_on
endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2019 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_DDC_E2.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//////////////////////////////////////////////////////////////////////////////
//
`timescale 1 ns / 1 ps

module GTP_DDC_E2 #(
parameter CLKA_GATE_EN = "FALSE",         //"TRUE":GATEI available; "FALSE":GATEI disable;
parameter WCLK_DELAY_SEL = "FALSE",         //"TRUE":Phase shift = 90; "FALSE":Phase shift = -90;
parameter DDC_MODE = "QUAD_RATE",         //"HALF_RATE"; "QUAD_RATE";
parameter R_EXTEND = "FALSE",         //"TRUE":gate delay; "FALSE": gate no delay;
parameter DELAY_SEL = 1'b0,         //1'b0: 1x delay range (~0.9ns); 1'b1: 2x delay range (~1.8-2.5ns);
parameter GRS_EN ="TRUE",         //"TRUE":GRS_N is available;"FALSE":GRS_N is disable;
parameter IFIFO_GENERIC = "FALSE",          //"TRUE":GENERIC mode;"FALSE":DDR MEM mode
parameter [2:0] RADDR_INIT = 3'b000,           //The initial value of read address in GENERIC mode
parameter [1:0] DATA_RATE = 2'b00              //2'b00, IO data rate: 533-2133Mbps;2'b01, IO data rate: 400Mbps;
)(
    //output
    output WCLK,
    output WCLK_DELAY,
    output DQSI_DELAY,
    output DQSIB_DELAY,
    output DGTS,
    output [2:0] IFIFO_WADDR,
    output [2:0] IFIFO_RADDR,
    output READ_VALID,
    output [1:0] DQS_DRIFT,
    output DRIFT_DETECT_ERR,
    output DQS_DRIFT_STATUS,
    output DQS_SAMPLE,
    //input
    input RST,
    input RST_TRAINING_N,
    input CLKA,
    input CLKB,
    input DQSI,
    input DQSIB,
    input [7:0] DELAY_STEP0,
    input [7:0] DELAY_STEP1,
    input [7:0] DELAY_STEP2,
    input [7:0] DELAY_STEP3,
    input [7:0] DELAY_STEP4,
    input [3:0] DQS_GATE_CTRL,
    input GATE_SEL,
    input [1:0] CLK_GATE_CTRL,
    input CLKA_GATE
)/* synthesis syn_black_box */;

//synthesis translate_off
    //reg statement
    reg [2:0]sc_dqs_mode;
   //wire statement
    wire [7:0] dqs_even_code;
    wire [7:0] dqs_odd_code;
    wire [7:0] wl_step;
    wire [7:0] wl_p_dllcode;
    wire [3:0] dqs_gate_ctrl;
    wire sc_gate_en;
    wire sc_wclkdel_sel;
//    wire sc_clkr_sel;
    wire sc_wl_extend;
    wire sc_dly_2x;
    wire [1:0] sc_rst_ctrl;
    wire [4:0] sc_en_ctrl;
    wire sc_fifomode_sel;
    wire sc_ififo_generic;
    wire [2:0]sc_rd_addr_init;
    wire ldo_ctrl;
    wire grs_n;
    wire [2:0] read_clk_ctrl;
    wire SC_DQS_GATE_SEL;
    wire GLOGEN;
    wire VCC_IO;
    wire VSS;
// DQSL.v
    wire [3:0] q;
    wire dqs_gate_ctrl_gate_dly;
    wire dqs_clean;
    reg new_transfer;
    wire set_en;
    wire rst_en;
    wire s0;
    wire s1;
    wire s2;
    wire wclk_sel_div2;
    wire clk_io_div2;
    reg wclk_source_dly;
    reg wclk_del_source_dly;
    reg dqsin_gated_dly;
    reg [1:0] dqs_gate_ctrl_gate_d;
    reg [1:0] dqs_gate_ctrl_gate_dd;
    reg [3:0] dqs_gate_ctrl_d1;
    reg [3:0] dqs_gate_ctrl_d2;
    reg [3:0] dqs_gate_ctrl_d3;
    reg gate_st;
    reg [3:0] dqs_gate_ctrl_d4;
    reg dqs_gate_ctrl_d5;
    reg dqs_gate_ctrl_d6;
    reg sel_gate_clk;
    reg dqs_ena;
    reg dqs_gate_ctrl_comb_d1;
    reg dqs_gate_ctrl_comb_d2;
    reg dqs_gate_ctrl_comb_d3;
    reg [1:0] dqs_gate_ctrl_comb_and_d;
    reg start_wr;
    reg [2:0] waddr_reg;
    reg [2:0] ififo_waddr_reg;
    reg start_rd;
    reg [2:0] raddr_reg;
    reg rdvalid_reg;
    reg [7:0] adj_dly_wclk_del; //kylau: dll_code+wl_code
    reg [7:0] adj_dly_dqsi;
    reg read_enable_tmp;
    reg new_st;
    reg new_transfer_d;
    reg read_enable_d1;
    reg read_enable_d2;
    reg [1:0] cnt;
    reg [1:0] gate_cnt;
    reg [1:0] new_cnt;
    reg [2:0] gate_d;
    reg [2:0] waddr_reg_d1;
    reg [2:0] waddr_reg_d2;
    reg [2:0] raddr_reg_plus1;
    reg new_rd_en_reg;
    reg [1:0] cnt_gate;
    reg [2:0] fifo_state_check_reg;
    reg init_rd_en_reg;
    reg init_rd_en;
    reg new_cnt_reg;
    //reg [3:0] q;
    reg [1:0] dqs_drift_reg;
    reg drift_status_reg; 
    reg drift_detect_err_reg;
    reg w_move_enable;
    reg r_move_enable;
    reg init_rd_en_x1;

initial
begin
    if ((CLKA_GATE_EN == "TRUE")  || (CLKA_GATE_EN == "FALSE")) begin
    end
    else
        $display (" GTP_DDC_E2 error: illegal setting for CLKA_GATE_EN");

    if ((GRS_EN == "TRUE")  || (GRS_EN == "FALSE")) begin
    end
    else
        $display (" GTP_DDC_E2 error: illegal setting for GRS_EN");

    if ((WCLK_DELAY_SEL == "TRUE")  || (WCLK_DELAY_SEL == "FALSE")) begin
    end
    else
        $display (" GTP_DDC_E2 error: illegal setting for WCLK_DELAY_SEL");

    if ((DDC_MODE == "HALF_RATE") || (DDC_MODE == "QUAD_RATE")) begin
    end
    else
        $display (" GTP_DDC_E2 error: illegal setting for DDC_MODE");

    if ((R_EXTEND == "TRUE")  || (R_EXTEND == "FALSE")) begin
    end
    else
        $display (" GTP_DDC_E2 error: illegal setting for R_EXTEND");

    if ((DELAY_SEL == 1'b1)  || (DELAY_SEL == 1'b0)) begin
    end
    else
        $display (" GTP_DDC_E2 error: illegal setting for DELAY_SEL");

    if ((DATA_RATE == 2'b00)  || (DATA_RATE == 2'b01)) begin
    end
    else
        $display (" GTP_DDC_E2 error: illegal setting for DATA_RATE");

    if ((IFIFO_GENERIC == "TRUE")  || (IFIFO_GENERIC == "FALSE")) begin
    end
    else
        $display (" GTP_DDC_E2 error: illegal setting for IFIFO_GENERIC");

    if ((RADDR_INIT == 3'b000)  || (RADDR_INIT == 3'b001) || (RADDR_INIT == 3'b010) || (RADDR_INIT == 3'b011) || (RADDR_INIT == 3'b100) || (RADDR_INIT == 3'b101) || (RADDR_INIT == 3'b110) || (RADDR_INIT == 3'b111)) begin
    end
    else
        $display (" GTP_DDC_E2 error: illegal setting for RADDR_INIT");
end

    initial 
    begin  
       dqs_gate_ctrl_gate_d = 2'b00;
       dqs_gate_ctrl_gate_dd = 2'b00;
       dqs_gate_ctrl_d1 = 4'b0000;
       dqs_gate_ctrl_d2 = 4'b0000;
       dqs_gate_ctrl_d3 = 4'b0000;
       gate_st          = 1'b0;
       dqs_gate_ctrl_d4 = 4'b0000;
       dqs_gate_ctrl_d5 = 1'b0;
       dqs_gate_ctrl_d6 = 1'b0;
       sel_gate_clk = 1'b0;
       dqs_ena = 1'b0;
       dqs_gate_ctrl_comb_d1 = 1'b0;
       dqs_gate_ctrl_comb_d2 = 1'b0;
       dqs_gate_ctrl_comb_d3 = 1'b0;
       dqs_gate_ctrl_comb_and_d = 2'b00;
       start_wr  = 1'b0;
       waddr_reg = 3'b000;
       ififo_waddr_reg = 3'b000;
       start_rd  = 1'b0;
       raddr_reg = sc_rd_addr_init;
       rdvalid_reg = 1'b0;
       adj_dly_wclk_del = 8'b00000000;
       adj_dly_dqsi = 8'b00000000;
       read_enable_tmp = 1'b0;
       new_st = 1'b0;
       new_transfer_d = 1'b0;
       read_enable_d1 = 1'b0;
       read_enable_d2 = 1'b0;
       cnt = 2'b00;
       gate_cnt = 2'b00;
       new_cnt = 2'b00;  
       gate_d = 3'b000;
       waddr_reg_d1 = 3'b000;
       waddr_reg_d2 = 3'b000;
       raddr_reg_plus1 = 3'b000;
       new_rd_en_reg = 1'b0;
       cnt_gate = 2'b00;
       fifo_state_check_reg = 3'b000;
       init_rd_en_reg = 1'b0;
       init_rd_en = 1'b0;
       new_cnt_reg = 1'b0;
       //q = 4'b0000;
       dqs_drift_reg = 2'b00;
       drift_detect_err_reg = 1'b0;
       dqsin_gated_dly = 1'b0;
       wclk_source_dly = 1'b0;
       wclk_del_source_dly = 1'b0;
       w_move_enable = 1'b0;
       r_move_enable = 1'b0;
    end

    wire nextrd_eq_wr;
    wire rd_eq_wr;
    wire fifo_state_check;
    wire r_qq_en;
    wire r_en;
    wire lsr_rst_n;
    wire gatein;
    wire rst_fifo_n;
    wire rst_global;
    wire rst_local;
    wire rst;
    wire [1:0] cnt_gate_next;
    wire dqs_gate_ctrl_d2_d;
    wire rst_transfer_n;
    wire dqsw;
    wire dqsw90;

    assign rst_global = (sc_rst_ctrl[1] && GLOGEN) ? 1'b0 : (~grs_n);
    assign rst_local = sc_rst_ctrl[0] ? RST : ~RST;
    assign rst = rst_local||rst_global;
    assign lsr_rst_n = ~rst;     
    assign gatein = sc_gate_en ? (~CLKA_GATE) : 1'b1;
    assign rst_fifo_n = sc_en_ctrl[1] ? lsr_rst_n & gatein & RST_TRAINING_N : 1'b0;
    assign rst_transfer_n = sc_en_ctrl[1] ? lsr_rst_n : 1'b0;
    assign rst_start_rd = start_rd & rst_fifo_n;
//    assign TIE_HI = 1'b1;
//    assign TIE_LO = 1'b0;
    assign WCLK = dqsw && GLOGEN;
    assign WCLK_DELAY = GLOGEN? (sc_wclkdel_sel? ~dqsw90 : dqsw90) : 1'b0;



assign sc_gate_en          =(CLKA_GATE_EN    == "TRUE"   ) ? 1'b1 : 1'b0;
assign sc_wclkdel_sel      =(WCLK_DELAY_SEL == "TRUE"   ) ? 1'b1 : 1'b0;
assign sc_wl_extend        =(R_EXTEND     == "TRUE"   ) ? 1'b1 : 1'b0;
assign sc_dly_2x           =DELAY_SEL;
assign sc_fifomode_sel     =1'b1;
assign sc_ififo_generic    =(IFIFO_GENERIC == "TRUE"   ) ? 1'b1 : 1'b0;
assign sc_rd_addr_init	   = RADDR_INIT;
assign ldo_ctrl            = DATA_RATE;
assign grs_n               =(GRS_EN       == "TRUE" ) ? GRS_INST.GRSNET : 1'b1;
//assign grs_n               =1'b1;
assign sc_rst_ctrl[0]      =1'b1;
assign sc_rst_ctrl[1]      =(GRS_EN       == "TRUE"   ) ? 1'b0 : 1'b1;
assign read_clk_ctrl[2]    =GATE_SEL;
assign read_clk_ctrl[1]    =CLK_GATE_CTRL[1];
assign read_clk_ctrl[0]    =CLK_GATE_CTRL[0];
assign sc_en_ctrl          =5'b01110;
assign SC_DQS_GATE_SEL     =1'b1;
assign GLOGEN              =1'b1;
assign VCC_IO              =1'b1;
assign VSS                 =1'b0;

initial
begin
     case (DDC_MODE)
//        "FULL_RATE": sc_dqs_mode = 3'b000;
        "HALF_RATE": sc_dqs_mode = 3'b010;
        "QUAD_RATE": sc_dqs_mode = 3'b111;
        default:
             begin sc_dqs_mode = 3'b111;
             $display (" DDC_MODE error: illegal setting for DDC_MODE");
             $finish;
             end
     endcase
end
    ///////////////clock gate////////////////////////
    always @(negedge CLKA or posedge rst)
    begin
       if(rst) 
       begin
          gate_d <= 3'd0;
       end
       else
       begin
          gate_d <= {gate_d[1:0], ~gatein};
       end
    end
    always @(negedge CLKA or posedge rst)
    begin
       if(rst) 
       begin
          cnt_gate <= 2'b0;
       end
       else if((gate_d[2]==1'b1)||(cnt_gate!=2'b00))
       begin
          cnt_gate <= cnt_gate_next;
       end
    end

    assign cnt_gate_next[0] = ~cnt_gate[0];
    assign cnt_gate_next[1] = cnt_gate[0] ? ~cnt_gate[1] : cnt_gate[1];
    assign ioclk_gated = (gate_d[2]==1'b1)||(cnt_gate!=2'b0) ? 0 : CLKA;

////////////////////////////////write clock part//////////////////////////
    wire wclk_source;
    wire  [63:0] wl_code_therm;
    wire  [63:0] dll_45code_therm;
    wire  [63:0] wl_p_dllcode_therm;

    assign wclk_source = (sc_dqs_mode == 3'b000) ? CLKB : ioclk_gated;

    ddc_e2_ddrphy_gray2therm gray2therm0(.gray_code(DELAY_STEP0),       .therm_code(wl_code_therm), .vcc(VCC_IO), .vss(VSS));
    ddc_e2_ddrphy_gray2therm gray2therm1(.gray_code(DELAY_STEP3),   .therm_code(dll_45code_therm), .vcc(VCC_IO), .vss(VSS));
    ddc_e2_ddrphy_gray2therm gray2therm2(.gray_code(DELAY_STEP4), .therm_code(wl_p_dllcode_therm), .vcc(VCC_IO), .vss(VSS));

    ddc_e2_dly_chain  dly_chain0(.dly_en(sc_en_ctrl[3]), .dly_sel(sc_dly_2x), .therm_code(wl_code_therm),       .din(wclk_source), .ldo_ctrl(ldo_ctrl), .d_dly(dqsw));
    ddc_e2_dly_chain  dly_chain1(.dly_en(sc_en_ctrl[3]), .dly_sel(1'b0),      .therm_code({64{1'b0}}),          .din(wclk_source), .ldo_ctrl(ldo_ctrl), .d_dly(clk_r0));
    ddc_e2_dly_chain  dly_chain2(.dly_en(sc_en_ctrl[3]), .dly_sel(sc_dly_2x), .therm_code(wl_p_dllcode_therm),  .din(wclk_source), .ldo_ctrl(ldo_ctrl), .d_dly(dqsw90));
    //ddc_e2_dly_chain  dly_chain3(.dly_en(sc_en_ctrl[3]), .dly_sel(sc_dly_2x), .therm_code(dll_45code_therm),    .din(wclk_source), .d_dly(clk_r90));
    ddc_e2_dly_chain  dly_chain3(.dly_en(sc_en_ctrl[3]), .dly_sel(1'b0), .therm_code(dll_45code_therm),    .din(wclk_source), .ldo_ctrl(ldo_ctrl), .d_dly(clk_r90));

/////////////////////////read clock part//////////////////////////////////
    wire [3:0] dqs_gate_ctrl_tmp;
    wire sel_x1;
    wire sel_x2;
    wire sel_x4;
    wire sel_x2x4;
    wire gate_reg_x1;
    reg  gate_reg;

    assign sel_x1 = (sc_dqs_mode==0)? 1'b1:1'b0;
    assign sel_x2 = (sc_dqs_mode==2)? 1'b1:1'b0;
    assign sel_x4 = (sc_dqs_mode==7)? 1'b1:1'b0;
    assign sel_x2x4 = (sc_dqs_mode[1:0]== 2'b00)? 1'b0 : 1'b1; 

    assign dqs_gate_ctrl_tmp = sc_en_ctrl[0] ? 4'b1111 : DQS_GATE_CTRL;
    
    assign gate_reg_x1 = dqs_gate_ctrl_d2_d;

    always @(posedge CLKB or negedge lsr_rst_n)
    begin
       if(!lsr_rst_n) 
       begin
          dqs_gate_ctrl_d1 <= 4'b0000;
          dqs_gate_ctrl_d2 <= 4'b0000;
       end
       else 
       begin
          if(sel_x4)
          begin
             dqs_gate_ctrl_d2 <= dqs_gate_ctrl_tmp;
          end
          else 
          begin
             dqs_gate_ctrl_d1 <= {2'b00,dqs_gate_ctrl_tmp[1:0]};
             dqs_gate_ctrl_d2 <= dqs_gate_ctrl_d1;   
          end
       end
    end

   wire  dqsw_tree;
   wire  dqsw_ls;
   wire  dqsw270_tree;
   wire  dqsw270_ls;

   assign dqsw_tree = clk_r0;
   assign dqsw270_tree = ~clk_r90;
   assign dqsw_ls = GLOGEN? dqsw_tree : 1'b0;
   assign dqsw270_ls = GLOGEN? dqsw270_tree : 1'b0;
   assign wclk_sel = sel_x1? CLKB : dqsw_ls;

   reg wclk_cnt;
   wire wclk_clk;
   always @(posedge wclk_sel or negedge lsr_rst_n)
   begin
      if(!lsr_rst_n)
          wclk_cnt <= 1'b0;
      else
          wclk_cnt <= wclk_cnt + 1'b1;
   end
   assign wclk_sel_div2 = wclk_cnt;

   assign wclk_clk = sel_x1 ? wclk_sel : wclk_sel_div2;

   /////uqdate_0///
   wire uqdate_rstn;
   wire uqdate_0_sel;
   wire cnt_0;
   wire cnt_1;
   wire cnt_1_in;
   wire cnt_1_rstn;
   reg  uqdate_0;

   assign cnt_1_in   = cnt_0 ^ cnt_1;
   assign cnt_1_rstn = uqdate_rstn & (~sel_x2);
   assign uqdate_0_sel = (~cnt_0 & sel_x2) | (cnt_0 & ~cnt_1 & sel_x4);

    reg dout;
always @(posedge wclk_clk or negedge lsr_rst_n)
begin
   if (!lsr_rst_n)
      dout <= 1'b0;
   else
      dout <= 1'b1;
   end
   assign uqdate_rstn = dout;

    reg dout_1;
always @(posedge wclk_clk or negedge uqdate_rstn)
begin
   if (!uqdate_rstn)
      dout_1 <= 1'b0;
   else
      dout_1 <= ~cnt_0;
   end
   assign cnt_0 = dout_1;

    reg dout_2;
always @(posedge wclk_clk or negedge cnt_1_rstn)
begin
   if (!cnt_1_rstn)
      dout_2 <= 1'b0;
   else
      dout_2 <= cnt_1_in;
   end
   assign cnt_1 = dout_2;



   always @(posedge wclk_clk or negedge uqdate_rstn)
   begin
      if(!uqdate_rstn) 
      begin
         uqdate_0 <= 0;
      end 
      else if(uqdate_0_sel)
      begin
         uqdate_0 <=  1;
      end
      else
      begin
         uqdate_0 <=  0;
      end
   end
   /////uqdate_1///
   wire uqdate_1_sel;
   wire uqdate_1_sel_a;
   wire uqdate_1_sel_b;
   wire uqdate_1;
   reg  uqdate_1_reg;

   assign uqdate_1_sel_a = (cnt_0 & sel_x2) | (~cnt_0 & ~cnt_1 & sel_x4);
   assign uqdate_1_sel_b = (~cnt_0 & sel_x2) | (cnt_0 & ~cnt_1 & sel_x4);
   assign uqdate_1_sel   = (sc_wl_extend==0) ? uqdate_1_sel_a:uqdate_1_sel_b;
   assign uqdate_1 = uqdate_1_reg | sel_x1;

   always @(posedge wclk_clk or negedge uqdate_rstn)
   begin
      if(!uqdate_rstn) 
      begin
         uqdate_1_reg <= 0;
      end 
      else
      begin
        uqdate_1_reg <= uqdate_1_sel;
      end
      //else if(uqdate_1_sel)
      //begin
      //   uqdate_1_reg <=  1;
      //end
      //else 
      //begin
      //   uqdate_1_reg <=  0;
      //end
   end

   always @(posedge wclk_clk or negedge lsr_rst_n)
   begin   
      if(!lsr_rst_n)
      begin
         dqs_gate_ctrl_d3 <= 4'b0;
      end
      else if (uqdate_0)
      begin
         dqs_gate_ctrl_d3 <= dqs_gate_ctrl_d2;
      end
   end

   //assign #0.2 dqs_gate_ctrl_d3_d = dqs_gate_ctrl_d3;
   //assign #0.2 dqs_gate_ctrl_d2_d = dqs_gate_ctrl_d2[0];
   wire [3:0] dqs_gate_ctrl_d3_d;
   assign dqs_gate_ctrl_d3_d = dqs_gate_ctrl_d3;
   assign dqs_gate_ctrl_d2_d = dqs_gate_ctrl_d2[0];

   always @(posedge wclk_clk or negedge lsr_rst_n) //KY
   begin
      if(!lsr_rst_n)
      begin
         dqs_gate_ctrl_d4 <= 4'b0000;
      end
      else if (uqdate_1)
      begin
        dqs_gate_ctrl_d4 <= dqs_gate_ctrl_d3_d;     
      end
      else
      begin
         if(sel_x4)
         begin
            dqs_gate_ctrl_d4 <= {1'b0, dqs_gate_ctrl_d4[3:1]};
         end
         else
         begin
            dqs_gate_ctrl_d4 <= {1'b0, dqs_gate_ctrl_d4[3],1'b0,dqs_gate_ctrl_d4[1]};
         end
      end
   end

   always @(posedge wclk_sel or negedge lsr_rst_n)
   begin   
      if(!lsr_rst_n)
      begin
         gate_reg <= 1'b0;
      end
      else
      begin
      gate_reg<=dqs_gate_ctrl_d4[0];
      end
   end

   
   always @(posedge wclk_sel or negedge lsr_rst_n)
   begin   
      if (!lsr_rst_n) 
      begin
         dqs_gate_ctrl_d5 <= 1'b0;
      end   
      else 
      begin      
         if (sel_x2x4)
         begin
            dqs_gate_ctrl_d5 <= gate_reg;
         end
         else
         begin
            dqs_gate_ctrl_d5 <= gate_reg_x1;
         end
      end
   end

   always @( * )  
   begin
      case (read_clk_ctrl[1:0])
         2'b00: sel_gate_clk = ~dqsw270_ls;
         2'b01: sel_gate_clk = ~wclk_sel;
         2'b10: sel_gate_clk = dqsw270_ls;
         2'b11: sel_gate_clk = wclk_sel;
      endcase
   end

   always @( * )
   begin
      case ({read_clk_ctrl[2], sel_x2x4})
         2'b00: dqs_gate_ctrl_d6 = gate_reg_x1;
         2'b01: dqs_gate_ctrl_d6 = gate_reg;
         2'b10: dqs_gate_ctrl_d6 = dqs_gate_ctrl_d5;
         2'b11: dqs_gate_ctrl_d6 = dqs_gate_ctrl_d5;
      endcase    
   end

   always @(posedge sel_gate_clk or negedge lsr_rst_n)
   begin
      if (!lsr_rst_n)
      begin
         dqs_gate_ctrl_comb_d1 <= 1'b0;
       //  dqs_gate_ctrl_comb_d2 <= 1'b0;
      end
      else 
      begin
         dqs_gate_ctrl_comb_d1 <= dqs_gate_ctrl_d6;
      //   dqs_gate_ctrl_comb_d2 <= dqs_gate_ctrl_comb_d1;
      end
   end

   always @(negedge sel_gate_clk or negedge lsr_rst_n)
   begin
      if (!lsr_rst_n)
      begin
         //dqs_gate_ctrl_comb_d1 <= 1'b0;
         dqs_gate_ctrl_comb_d2 <= 1'b0;
      end
      else 
      begin
         //dqs_gate_ctrl_comb_d1 <= dqs_gate_ctrl_d6;
         dqs_gate_ctrl_comb_d2 <= dqs_gate_ctrl_comb_d1;
      end
   end
   
   always @(posedge sel_gate_clk or negedge lsr_rst_n)
   begin
      if (!lsr_rst_n)
      begin
         //dqs_gate_ctrl_comb_d1 <= 1'b0;
         dqs_gate_ctrl_comb_d3 <= 1'b0;
      end
      else 
      begin
         //dqs_gate_ctrl_comb_d1 <= dqs_gate_ctrl_d6;
         dqs_gate_ctrl_comb_d3 <= dqs_gate_ctrl_comb_d2;
      end
   end

   wire read_ena;
   //assign read_ena =  dqs_gate_ctrl_comb_d1 && dqs_gate_ctrl_comb_d2 ;
   assign read_ena =  dqs_gate_ctrl_comb_d1 && dqs_gate_ctrl_comb_d3;
   assign set_en = read_ena && rst_en;
   assign rst_en = lsr_rst_n && RST_TRAINING_N ;
   always @(negedge dqs_clean or negedge rst_en or posedge set_en)
   begin   
      if (!rst_en)
      begin
         dqs_ena <= 1'b0;
      end
      else if (set_en)
      begin
        dqs_ena <= 1'b1;
      end
      else
      begin
         if(SC_DQS_GATE_SEL)
         begin
            dqs_ena <= read_ena;
         end
         else
         begin
            dqs_ena <= 1'b0;
         end
      end
   end

   wire          dqs_cleanb;
   wire   [7:0]  dqs_even_code_g;
   wire   [7:0]  dqs_odd_code_g;
   wire   [63:0] dqs_even_code_t;
   wire   [63:0] dqs_odd_code_t;
   wire          dqsi_del;
   wire          dqsib_del;
   
   assign DQSI_DELAY  = GLOGEN? dqsi_del  : 1'b0;
   assign DQSIB_DELAY = GLOGEN? dqsib_del : 1'b0;
   assign dqs_clean = dqs_ena && DQSI;
   //assign dqs_cleanb = dqs_ena & DQSIB;
   assign dqs_cleanb = ~dqs_ena || DQSIB;
   assign dqs_even_code_g = sc_en_ctrl[4]? 8'b00000000 : DELAY_STEP1;
   assign dqs_odd_code_g = sc_en_ctrl[4]? 8'b00000000 : DELAY_STEP2;

   ddc_e2_ddrphy_gray2therm gray2therm3(.gray_code(dqs_even_code_g),  .therm_code(dqs_even_code_t), .vcc(VCC_IO), .vss(VSS));
   ddc_e2_ddrphy_gray2therm gray2therm4(.gray_code(dqs_odd_code_g),   .therm_code(dqs_odd_code_t),  .vcc(VCC_IO), .vss(VSS));
   
   //ddc_e2_dly_chain  dly_chain4(.dly_en(sc_en_ctrl[2]), .dly_sel(sc_dly_2x), .therm_code(dqs_even_code_t), .din(dqs_clean), .d_dly(DQSI_DELAY));
   //ddc_e2_dly_chain  dly_chain5(.dly_en(sc_en_ctrl[2]), .dly_sel(sc_dly_2x), .therm_code(dqs_odd_code_t),  .din(dqs_cleanb), .d_dly(DQSIB_DELAY));

   ddc_e2_dly_chain  dly_chain4(.dly_en(sc_en_ctrl[2]), .dly_sel(sc_dly_2x), .therm_code(dqs_even_code_t), .din(dqs_clean), .ldo_ctrl(ldo_ctrl), .d_dly(dqsi_del));
   ddc_e2_dly_chain  dly_chain5(.dly_en(sc_en_ctrl[2]), .dly_sel(sc_dly_2x), .therm_code(dqs_odd_code_t),  .din(dqs_cleanb), .ldo_ctrl(ldo_ctrl), .d_dly(dqsib_del));

   //KYLAU: sample DQSI for DQS_gate training
   wire s0_dly;


   
    reg dout_3;
always @(posedge read_ena or negedge rst_en)
begin
   if (!rst_en)
      dout_3 <= 1'b0;
   else
      dout_3 <= DQSI;
   end
   assign s0 = dout_3;


   assign #0.00001  s0_dly = s0;



    reg dout_4;
always @(posedge dqsw_ls or negedge rst_en)
begin
   if (!rst_en)
      dout_4 <= 1'b0;
   else
      dout_4 <= s0_dly;
   end
   assign s1 = dout_4;




    reg dout_5;
always @(posedge dqsw_ls or negedge rst_en)
begin
   if (!rst_en)
      dout_5 <= 1'b0;
   else
      dout_5 <= s1;
   end
   assign s2 = dout_5;



    reg dout_6;
always @(posedge dqsw_ls or negedge rst_en)
begin
   if (!rst_en)
      dout_6 <= 1'b0;
   else
      dout_6 <= s2;
   end
   assign DQS_SAMPLE = dout_6;


   ////////////////////Drift detection/////////////////////////////  
   
   reg [3:0] q_reg;
   always@(posedge read_ena or negedge lsr_rst_n) 
   begin
      if(!lsr_rst_n)
      begin
         drift_status_reg <= 1'b0;
      end
      else
      begin
         drift_status_reg <=DQSI;
      end
   end

   always @(posedge dqs_clean or negedge lsr_rst_n)
   begin
      if(!lsr_rst_n)
      begin
         q_reg <= 4'b0000;
      end
      else
      begin
         q_reg <= {~dqsw270_ls, ~wclk_sel, dqsw270_ls, wclk_sel};
      end
   end
   
   assign q = q_reg;

   always @(posedge dqs_clean or negedge lsr_rst_n)
   begin
      if(!lsr_rst_n)
      begin
         dqs_drift_reg <= 2'b00;
         drift_detect_err_reg <= 1'b0;
      end
      else
      begin
         case(q)
            4'b0000:begin
               drift_detect_err_reg <= 1'b0;
            end
            4'b0001:begin
               dqs_drift_reg <= 2'b00;
               drift_detect_err_reg <= 1'b0;
            end
            4'b1001:begin
               dqs_drift_reg <= 2'b00;
               drift_detect_err_reg <= 1'b0;
            end
            4'b1101:begin
               dqs_drift_reg <= 2'b00;
               drift_detect_err_reg <= 1'b0;
            end
            4'b1000:begin
               dqs_drift_reg <= 2'b01;
               drift_detect_err_reg <= 1'b0;
            end
            4'b1100:begin
               dqs_drift_reg <= 2'b01;
               drift_detect_err_reg <= 1'b0;
            end
            4'b1110:begin
               dqs_drift_reg <= 2'b01;
               drift_detect_err_reg <= 1'b0;
            end
            4'b0100:begin
               dqs_drift_reg <= 2'b11;
               drift_detect_err_reg <= 1'b0;
            end
            4'b0110:begin
               dqs_drift_reg <= 2'b11;
               drift_detect_err_reg <= 1'b0;
            end
            4'b0111:begin
               dqs_drift_reg <= 2'b11;
               drift_detect_err_reg <= 1'b0;
            end
            4'b1011:begin
               dqs_drift_reg <= 2'b10;
               drift_detect_err_reg <= 1'b0;
            end
            4'b0010:begin
               dqs_drift_reg <= 2'b10;
               drift_detect_err_reg <= 1'b0;
            end
            4'b0011:begin
               dqs_drift_reg <= 2'b10;
               drift_detect_err_reg <= 1'b0;
            end
            4'b0101:begin
               drift_detect_err_reg <= 1'b1;
            end
            4'b1010:begin
               drift_detect_err_reg <= 1'b1;
            end
            4'b1111:begin
               drift_detect_err_reg <= 1'b1;
            end
            default:begin
               dqs_drift_reg <= 2'b00;
               drift_detect_err_reg <= 1'b0;
            end 
         endcase   
      end
   end

   assign DQS_DRIFT = GLOGEN ? dqs_drift_reg : 2'b11;
   assign DRIFT_DETECT_ERR = GLOGEN ? drift_detect_err_reg : 1'b1;
   assign DQS_DRIFT_STATUS = GLOGEN ? drift_status_reg : 1'b1;
//////////////////////////////busrt_det/////////////////////////////////
   
   wire  dqs_gate_ctrl_comb_d1_dly;
   assign #0.2 dqs_gate_ctrl_comb_d1_dly = dqs_gate_ctrl_comb_d1;
   assign dqs_gate_ctrl_comb_d1_rising = dqs_gate_ctrl_comb_d1 & (~dqs_gate_ctrl_comb_d1_dly);
   assign dqs_gate_ctrl_gate_dly = dqs_ena;
   //assign #0.1 dqs_gate_ctrl_gate_dly = dqs_ena;
   
   //assign dqs_gate_ctrl_comb_d1_dly = dqs_gate_ctrl_comb_d1;
   //assign dqs_gate_ctrl_comb_d1_rising = dqs_gate_ctrl_comb_d1 & (~dqs_gate_ctrl_comb_d1_dly);
   //assign dqs_gate_ctrl_gate_dly = dqs_ena;
   //counter0
   always @(posedge dqs_clean or posedge dqs_gate_ctrl_comb_d1_rising or negedge lsr_rst_n or negedge RST_TRAINING_N)
   begin
      if (!lsr_rst_n)
      begin
         dqs_gate_ctrl_gate_d <= 2'b00;
      end
      else if (!RST_TRAINING_N)
      begin
         dqs_gate_ctrl_gate_d <= 2'b00;
      end
      else if (dqs_gate_ctrl_comb_d1_rising)
      begin
         dqs_gate_ctrl_gate_d <= 2'b00;
      end
      else if (dqs_gate_ctrl_gate_dly) 
      begin
        dqs_gate_ctrl_gate_d <= dqs_gate_ctrl_gate_d + 1;  
      end
   end

   //counter1
   always @(negedge dqs_clean or posedge dqs_gate_ctrl_comb_d1_rising or negedge lsr_rst_n or negedge RST_TRAINING_N)
   begin   
      if (!lsr_rst_n)
      begin
         dqs_gate_ctrl_gate_dd <= 2'b00;
      end
      else if (!RST_TRAINING_N)
      begin
         dqs_gate_ctrl_gate_dd <= 2'b00;
      end
      else if (dqs_gate_ctrl_comb_d1_rising)
      begin
          dqs_gate_ctrl_gate_dd <= 2'b00;
      end
      else
      begin
         dqs_gate_ctrl_gate_dd <= dqs_gate_ctrl_gate_dd + 1;
      end
   end

   //counter2
   always @(negedge dqs_clean or posedge dqs_gate_ctrl_comb_d1_rising or negedge lsr_rst_n or negedge RST_TRAINING_N)
   begin
      if (!lsr_rst_n)
      begin
         dqs_gate_ctrl_comb_and_d <= 2'b00;
      end
      else if (!RST_TRAINING_N)
      begin
         dqs_gate_ctrl_comb_and_d <= 2'b00;
      end
      else if (dqs_gate_ctrl_comb_d1_rising)
      begin
         dqs_gate_ctrl_comb_and_d <= 2'b00;
      end
      else if (read_ena) 
      begin
         dqs_gate_ctrl_comb_and_d <= dqs_gate_ctrl_comb_and_d + 1;
      end
   end
 
   assign dgts_a = (~dqs_gate_ctrl_gate_dly) && (dqs_gate_ctrl_gate_d == 2'b00);
   assign dgts_b = (dqs_gate_ctrl_gate_dd == 2'b00) &&  (dqs_gate_ctrl_comb_and_d == 2'b11);
   assign DGTS = GLOGEN ? dgts_a & dgts_b : 1'b1;

/////////////////////////////ififo management////////////////////////
   ///ififo_w
   always @(posedge DQSI_DELAY or negedge rst_fifo_n)
   begin   
      if (!rst_fifo_n)
      begin
         start_wr <= 1'b0;
      end
      else
      begin
         start_wr <= rst_fifo_n;
      end
   end

   assign start_wr_comb = (sc_ififo_generic == 1'b1) ?  start_wr : rst_fifo_n;

   always @(posedge DQSI_DELAY or negedge start_wr_comb)
   begin
      if (!start_wr_comb)
      begin
         waddr_reg <= 3'b000;
      end
      else 
      begin
         case (waddr_reg)
            3'b000: waddr_reg <= 3'b001;
            3'b001: waddr_reg <= 3'b011;
            3'b011: waddr_reg <= 3'b010;
            3'b010: waddr_reg <= 3'b110;
            3'b110: waddr_reg <= 3'b111;
            3'b111: waddr_reg <= 3'b101;
            3'b101: waddr_reg <= 3'b100;
            3'b100: waddr_reg <= 3'b000;
         endcase
      end
   end

   always @(negedge DQSI_DELAY or negedge start_wr_comb)
   begin
      if (!start_wr_comb)
      begin
         ififo_waddr_reg <= 3'b000;
      end
      else
      begin
        ififo_waddr_reg <= waddr_reg;
      end
   end

   assign IFIFO_WADDR = ififo_waddr_reg;

   //clk_io_div2 generation 
    reg dout_7;
always @(posedge CLKA or negedge lsr_rst_n)
begin
   if (!lsr_rst_n)
      dout_7 <= 1'b0;
   else
      dout_7 <= ~clk_io_div2;
   end
   assign clk_io_div2 = dout_7;


   //mode1
   assign rd_clk = sel_x1? CLKB : clk_io_div2;

   always @(posedge rd_clk or negedge rst_fifo_n)
   begin
      if (!rst_fifo_n)
      begin
        start_rd <= 1'b0;
      end
      else
      begin
         start_rd <= rst_fifo_n;
      end
   end
   
   always @(posedge rd_clk or negedge rst_start_rd)
   begin
      if (!rst_start_rd)
      begin
        waddr_reg_d1 <= 3'b000;
      end
      else
      begin
         waddr_reg_d1 <= waddr_reg;
      end
   end

   always @(posedge rd_clk or negedge rst_start_rd)
   begin
      if (!rst_start_rd)
      begin
         waddr_reg_d2 <= 3'b000;
      end
      else
      begin
         waddr_reg_d2 <= waddr_reg_d1;
      end
   end

   assign buffer_empty = (waddr_reg_d2 == raddr_reg) ? 1'b1 : 1'b0;
   assign buffer_almost_empty = (waddr_reg_d2 == raddr_reg_plus1) ? 1'b1 : 1'b0;

   //ififo_mgt_update
   always @(posedge rd_clk or negedge rst_transfer_n)
   begin
      if (!rst_transfer_n) 
      begin
         new_st         <= 1'b0;
         new_cnt        <= 2'b00;
         new_transfer_d <= 1'b0;
      end
      else 
      begin
         new_st       <= 1'b1;
         new_transfer_d <= new_transfer;
         if (new_st)
         begin
            new_cnt[0]      <= new_cnt[0] + 1;
            if(~sel_x2)
            begin
               new_cnt[1] <= new_cnt[1] ^ new_cnt[0];
            end
            else
            begin
               new_cnt[1] <= 1'b0;
            end
         end
      end
   end
   
   wire   transfer_sel;
   always @(posedge rd_clk or negedge new_st)
   begin
     if (!new_st)
      begin
         new_transfer <= 1'b0;
      end
      else
      begin
         if(transfer_sel)
         begin
            new_transfer  <= 1'b1;
         end
         else
         begin
            new_transfer  <= 1'b0;            
         end
      end
   end

   assign  transfer_sel  =  (sel_x2 && new_cnt[0]) || (new_cnt[0] && ~new_cnt[1] && sel_x4);

   
   always @(posedge rd_clk or negedge rst_start_rd)
   begin
      if (!rst_start_rd) 
      begin
         new_rd_en_reg <= 1'b0;
      end
      else if (sel_x1 || new_transfer)  //sel port
      begin  
         if (new_rd_en_reg) 
         begin
            if (buffer_almost_empty)
            begin
               new_rd_en_reg <= 1'b0;
            end
         end
         else 
         begin
            if (~buffer_empty)
            begin
               new_rd_en_reg <= 1'b1;
            end
         end
      end
   end

   //mode0
   assign rd_eq_wr =  (waddr_reg == raddr_reg) ? 1'b0 : 1'b1;
   assign nextrd_eq_wr = (waddr_reg  == raddr_reg_plus1) ? 1'b0 : 1'b1;

   assign fifo_state_check = (~sc_ififo_generic) && ((~init_rd_en_x1 && rd_eq_wr) || (init_rd_en_x1 && nextrd_eq_wr));

   always @(*)
   begin
      if(!rst_start_rd)
      begin
        fifo_state_check_reg[0] <= 1'b0;
      end
      else if(!rd_clk)
      begin
         fifo_state_check_reg[0] <= fifo_state_check;
      end
   end

   always @(negedge rd_clk or negedge rst_start_rd)
   begin
      if(!rst_start_rd)
      begin
        fifo_state_check_reg[1] <= 1'b0;
      end
      else
      begin
         fifo_state_check_reg[1] <= (~init_rd_en_x1)&&fifo_state_check_reg[0];
      end
   end

   always @(*)
   begin
      if(!rst_start_rd)
      begin
         fifo_state_check_reg[2] <= 1'b0;
      end
      else if(rd_clk)
      begin
         fifo_state_check_reg[2] <= fifo_state_check;    
      end
   end
   
   assign fifo_state_check_out = fifo_state_check_reg[2] && (sel_x1 || fifo_state_check_reg[1] || init_rd_en_x1);
   always @(posedge rd_clk or negedge rst_start_rd)
   begin
      if(!rst_start_rd)
      begin
        init_rd_en_x1 <= 1'b0;
      end
      else
      begin
        init_rd_en_x1 <= fifo_state_check_out;
      end
   end

   always @(posedge rd_clk or negedge rst_start_rd)
   begin
    if(!rst_start_rd)
    begin
       init_rd_en <= 1'b0;
    end
    else if(new_transfer)
    begin
       init_rd_en <= fifo_state_check_out;
    end
   end

    //ififo_r
   assign r_en = (sc_ififo_generic== 1'b1) ? 1'b1 : (sc_fifomode_sel ? new_rd_en_reg && (~buffer_empty) : init_rd_en_x1);
   assign r_qq_en = (sc_ififo_generic== 1'b1) ? 1'b1 : (sc_fifomode_sel ? new_rd_en_reg && (~buffer_empty) : init_rd_en);

   assign read_enable = sel_x1? r_en : r_qq_en;

   always @(posedge rd_clk or negedge rst_start_rd)
   begin
      if (!rst_start_rd)
      begin
         raddr_reg <= sc_rd_addr_init;
      end
      else if (read_enable) 
      begin
         case (raddr_reg)
            3'b000: raddr_reg <= 3'b001;
            3'b001: raddr_reg <= 3'b011;
            3'b011: raddr_reg <= 3'b010;
            3'b010: raddr_reg <= 3'b110;
            3'b110: raddr_reg <= 3'b111;
            3'b111: raddr_reg <= 3'b101;
            3'b101: raddr_reg <= 3'b100;
            3'b100: raddr_reg <= 3'b000;
         endcase
      end
      else
      begin
         raddr_reg <= raddr_reg;
      end
   end

   always @(*) 
   begin
      case (raddr_reg)
         3'b000: raddr_reg_plus1 = 3'b001;
         3'b001: raddr_reg_plus1 = 3'b011;
         3'b011: raddr_reg_plus1 = 3'b010;
         3'b010: raddr_reg_plus1 = 3'b110;
         3'b110: raddr_reg_plus1 = 3'b111;
         3'b111: raddr_reg_plus1 = 3'b101;
         3'b101: raddr_reg_plus1 = 3'b100;
         3'b100: raddr_reg_plus1 = 3'b000;
      endcase
   end

   assign IFIFO_RADDR = raddr_reg;
    
   //Read_valid
   always @(posedge rd_clk or negedge rst_start_rd)
   begin   
      if (!rst_start_rd) 
      begin
         read_enable_d1 <= 1'b0;
         read_enable_d2 <= 1'b0;
      end
      else 
      begin 
        if(sc_fifomode_sel)
        begin
           read_enable_d1 <= new_rd_en_reg && (~buffer_empty);
           if(new_transfer_d)
           begin
              read_enable_d2 <= read_enable_d1;
           end
        end
        else
        begin
           read_enable_d1 <= init_rd_en;
           if(new_transfer_d)
           begin
              read_enable_d2 <= read_enable_d1;
           end
        end
      end
   end


   always @(posedge CLKB or negedge rst_start_rd)
   begin
      if (!rst_start_rd)
      begin
         rdvalid_reg <= 1'b0;
      end
      else if (sel_x1) 
      begin
         rdvalid_reg <= r_en;
      end
      else
      begin
         rdvalid_reg <= read_enable_d2;
      end
   end

   assign READ_VALID = GLOGEN ? rdvalid_reg : 1'b1;
   //pragma translate_on
endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2016 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_KEYRAM.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_KEYRAM
#(

) (
    input   ERASE_KEY_N
);
//synthesis translate_off

    reg     [7:0]      net_addr;
    reg     [31:0]     net_data;
    wire    [31:0]     mem [7:0];
    wire            ERASE_KEY_N_A;
    wire            ERASE_KEY_N_D;

    assign ERASE_KEY_N_A = ERASE_KEY_N;
    assign #2 ERASE_KEY_N_D = ERASE_KEY_N_A;

    always@(*)begin
        if(!ERASE_KEY_N_A)
            net_addr = 8'b1111_1111;
        else
            net_addr = 8'b0000_0000;

        if(!ERASE_KEY_N_D)
            net_data = 32'b0;
    end

    assign mem[7] = net_addr[7] ? net_data : mem[7];
    assign mem[6] = net_addr[6] ? net_data : mem[6];
    assign mem[5] = net_addr[5] ? net_data : mem[5];
    assign mem[4] = net_addr[4] ? net_data : mem[4];
    assign mem[3] = net_addr[3] ? net_data : mem[3];
    assign mem[2] = net_addr[2] ? net_data : mem[2];
    assign mem[1] = net_addr[1] ? net_data : mem[1];
    assign mem[0] = net_addr[0] ? net_data : mem[0];


//synthesis translate_on
endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2016 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_OSC_E4
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_OSC_E4
(
    output     CLKOUT,
    input      EN_N
);
//synthesis translate_off

    //////////////////////////// OSC ///////////////////////////////////////////////////
    wire osc_en_cfg ;
    wire clk_cfg ;
    reg  POR_N;
    initial
    begin
    POR_N=1'b0;
    #0.1;
    POR_N=1'b1;
    end
    
    assign osc_en_cfg  = !EN_N;
    ////////////adc_syn////////////////////
    wire cfg_en_syn;
    wire cfgs_disable;
    reg [1:0] cfg_en_dly_cfgs;
    
    assign cfgs_disable = osc_en_cfg | cfg_en_dly_cfgs[1];
    assign cfg_en_syn   = cfgs_disable ;

    always @(negedge CLKOUT or negedge POR_N)
    begin
        if(!POR_N)
            cfg_en_dly_cfgs <= 0;
        else 
            cfg_en_dly_cfgs <= {cfg_en_dly_cfgs[0],osc_en_cfg};
    end 
    //OSC_CORE osc_cfg  (.OSCEN(cfg_en_syn ), .POR_N(POR_N), .OSC_ADC(1'b0), .OSC_FREQ_CTRL(4'h0 ), .CLKOUT(clk_cfg ));
    //OSC_DIV osc_div_cfg (.POR_N(POR_N), .OSCEN(cfgs_disable), .OSC_DIV_EN(1'b1), .CLKIN(clk_cfg ), .CLKOUT(CLKOUT));



//////////////////////////////////////////OSC_CORE///////////////////////////////////////////

    wire        OSCEN_CORE;
    wire        OSC_ADC;
    wire  [3:0] OSC_FREQ_CTRL;
    wire        CLKOUT_CORE;

    assign OSCEN_CORE = cfg_en_syn;
    assign OSC_ADC = 1'b0;
    assign OSC_FREQ_CTRL = 4'h0;
    assign clk_cfg = CLKOUT_CORE;

    wire        osc_rstn;
    reg         clk_reg;
    reg [3:0]   freq_ctrl;
    realtime clkout_time_half;
    assign CLKOUT_CORE =  clk_reg;
    assign osc_rstn = POR_N & OSCEN_CORE;
    
    
    initial begin
        clk_reg = 1'b0;
    end
    always@(*)
    begin
        if(OSC_ADC==0)
            freq_ctrl = OSC_FREQ_CTRL + 5;
        else 
            freq_ctrl = OSC_FREQ_CTRL;
    end
    always@(*)
    begin
        case(freq_ctrl) 
            4'h0:clkout_time_half = 2.40 ;
            4'h1:clkout_time_half = 2.42 ;
            4'h2:clkout_time_half = 2.44 ;
            4'h3:clkout_time_half = 2.46 ;
            4'h4:clkout_time_half = 2.48 ;
            4'h5:clkout_time_half = 2.50 ;
            4'h6:clkout_time_half = 2.52 ;
            4'h7:clkout_time_half = 2.54 ;
            4'h8:clkout_time_half = 2.56 ;
            4'h9:clkout_time_half = 2.58 ;
            4'ha:clkout_time_half = 2.60 ;
            4'hb:clkout_time_half = 2.62 ;
            4'hc:clkout_time_half = 2.64 ;
            4'hd:clkout_time_half = 2.68 ;
            4'he:clkout_time_half = 2.70 ;
            4'hf:clkout_time_half = 2.72 ;
            default: clkout_time_half = 2.5 ;
        endcase
    end

    always begin
        wait (osc_rstn == 1'b1) begin
            clk_reg = 1'b0;
            #clkout_time_half;
            clk_reg = 1'b1;
            #clkout_time_half;
        end
    end

    always begin
        wait (osc_rstn != 1'b1) begin
            force clk_reg = 1'b0;
            #2 release clk_reg;
        end
    end


///////////////////////////////////////////OSC_DIV///////////////////////////////////////////
    wire    OSCEN_DIV;
    wire    OSC_DIV_EN;
    wire    CLKIN;
    wire    CLKOUT_DIV;
    
    assign OSCEN_DIV = cfgs_disable;
    assign OSC_DIV_EN = 1'b1;
    assign CLKIN = clk_cfg;
    assign CLKOUT = CLKOUT_DIV;
   
    wire cfgs_rstn;
    wire div_en_syn;
    wire clk_out;
    reg  div_start;
    reg [1:0] div_en_dly;
    reg [1:0] div ;
    
    assign cfgs_rstn = POR_N & OSCEN_DIV;
    assign div_en_syn = OSC_DIV_EN | div_en_dly[1];
    assign clk_out = div[1];
    assign CLKOUT_DIV = clk_out & div_en_syn;


    always @(posedge CLKIN or negedge POR_N)
    begin
        if(!POR_N)
            div_start <= 1;
        else 
            div_start <= div_en_syn;
    end

    always @(posedge CLKIN or negedge cfgs_rstn)
    begin
        if(!cfgs_rstn)
            div<=0;
        else
        begin
            if(div_start)
                div<=div + 1'b1;
            else
                div<=0;
        end
    end

    always @(negedge clk_out or negedge cfgs_rstn)
    begin
        if(!cfgs_rstn)
            div_en_dly <= 0;
        else 
            div_en_dly <= {div_en_dly[0],OSC_DIV_EN};
    end
//synthesis translate_on
endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2016 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_IPAL_E2
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_IPAL_E2
#(
    parameter            SIM_DEVICE = "PG2L100H",// for cmem
    parameter     [31:0] IDCODE = 32'haaaa5555,
    parameter            DATA_WIDTH = "X8" //X8, X16, X32, Ipal data width select
) (
    output        [31:0] DO,//Ipal data out
    output               RBCRC_ERR,//readback CRC error flag
    output               RBCRC_VALID,//readback CRC result valid
    output               ECC_VALID,//SEU result valid
    output        [11:0] ECC_INDEX,//address of single error bit
    output               SERROR,//single-bit error flag
    output               DERROR,//double-bit error flag
    output   reg  [7:0]  SEU_FRAME_ADDR,//current frame address of SEU
    output   reg  [7:0]  SEU_COLUMN_ADDR,//current column address of SEU
    output   reg  [4:0]  SEU_REGION_ADDR,//current region address of SEU
    output   reg  [7:0]  SEU_FRAME_NADDR,//next frame address of SEU
    output   reg  [7:0]  SEU_COLUMN_NADDR,//next column address of SEU
    output   reg  [4:0]  SEU_REGION_NADDR,//next region address of SEU
    output               PRCFG_OVER,// Partial reconfiguration over pulse
    output               PRCFG_ERR,// Partial reconfiguration error flag
    output               DRCFG_OVER,
    output               DRCFG_ERR,
    
    input                RST_N,
    input                CLK,// 50M system clock
    input                CS_N,// chip select to enable the pal data bus, active low
    input                RW_SEL,//Ipal rdw, 0: write, 1: read
    input        [31:0]  DI//Ipal data in
 
);



//synthesis translate_off
    localparam          HEADER       =  1'b0;
    localparam          DAT          =  1'b1;

    wire    [31:0]  data; //aligned 32-bit input data
    wire            data_valid;
    wire            flg_rcmem;
    wire            flg_read_tmp;
    wire            flg_write_tmp;
    wire            flg_type1;
    wire            flg_type2;
    wire    [26:0]  word_count_tmp;
    wire            flg_desync;
    wire            flg_prcfgen;
    wire            flg_prcfgdis;
    wire            flg_drcfgen;
    wire            flg_drcfgdis;
    wire            flg_rbcrc;
    wire            flg_rrbcrc;
    wire            rbcrc_en;
    wire            seu_en;
    wire            re_rb;
    wire            we;
    wire            flg_rb_reg;
    wire    [1:0]   cmemtype;
    wire    [4:0]   addr_region;
    wire    [7:0]   addr_column;
    wire    [7:0]   addr_frame;
    wire            region0;
    wire            region1;
    wire            region2;
    wire            region3;
    wire            serror;
    wire            derror;
    wire    [11:0]  index; 
    wire            cmemclk;
    wire            crc_err;
    wire            flg_rstcrc;
    wire            prcfg_err;
    wire            drcfg_err;
    


    reg     [31:0]  data_rb;
    reg     [1:0]   ipal_m;
    reg     [4:0]   regaddr;
    reg             flg_write;
    reg             flg_rb_cmem;
    reg             flg_rb_cmem_d;
    reg             s;
    reg             ns;
    reg     [26:0]  word_count;
    reg     [26:0]  word_count_rb;
    reg             prcfg_en;
    reg             prcfg_en_d;
    reg             prcfg_over;
    reg             drcfg_en; 
    reg             drcfg_en_d;   
    reg             drcfg_over;
    
    reg     [4:0]   reg_cmd;
    reg     [31:0]  data_rb_reg;  
    reg             serror_d;
    reg             derror_d;
    reg     [3231:0]cmem [0:7999];
    reg             [13:0] addr_row;
    reg             [13:0] naddr_row;
    reg             [6:0] addr_word;
    reg             flg_region_end;
    reg             flg_column_end;
    reg             flg_frame_end;


    reg     [31:0]  reg_crcr;
    reg     [31:0]  reg_idr;
    reg     [31:0]  reg_cmdr;
    reg     [31:0]  reg_ctrl0r;
    reg     [31:0]  reg_ctrl1r;
    reg     [31:0]  reg_cmemir;
    reg     [31:0]  reg_mfwriter;
    reg     [95:0]  reg_ivr;
    reg     [31:0]  reg_chainr;
    reg     [31:0]  reg_adrr;
    reg     [31:0]  reg_sbpir;
    reg     [31:0]  reg_seur;
    reg     [31:0]  reg_irstctrlr;
    reg     [31:0]  reg_irstadrr;
    reg     [31:0]  reg_watchdogr;
    reg     [31:0]  reg_cmaskr;
    reg     [255:0]  reg_keyr;
    reg     [31:0]  reg_option0r;
    reg     [31:0]  reg_option1r;
    reg     [31:0]  reg_rcrr;
    reg     [8383:0]  reg_autr;
    reg     [31:0]  reg_seuaddr;
    reg     [31:0]  reg_seunaddr;

    reg     [31:0]  reg_cmemor;
    reg     [31:0]  reg_statusr;
    reg     [31:0]  reg_seustatusr;
    reg     [31:0]  reg_hstatusr;
    reg     [31:0]  reg_adrr_seu;

    integer         i;




///////////////////////////////////////////////////ISPAL/////////////////////////////////////////////////////////////
    integer count_csn;
    always@(posedge CLK or negedge CS_N) begin
        if(!CS_N) begin
            count_csn <= 0;
        end
        else begin
            count_csn <= count_csn + 1;
        end
    end

    always@(negedge CS_N) begin
        if(RW_SEL && flg_rcmem && count_csn < 40) begin
            $display("[Warning] : In GTP_IPAL_E2, CS_N = 1 must last for at least 40 CLK cycle when reading back configuration memory. at time%t",$realtime);                  
        end
        else if(RW_SEL && flg_rb_reg && count_csn < 20) begin
            $display("[Warning] : In GTP_IPAL_E2, CS_N = 1 must last for at least 20 CLK cycle when reading back configuration register. at time%t",$realtime);                
        end
    end

    initial begin
        case(DATA_WIDTH)
            "X8"  :  ipal_m = 2'd0;
            "X16" :  ipal_m = 2'd1;
            "X32" :  ipal_m = 2'd2;
          default :  begin
                     ipal_m = 2'd0;
                     $display("Setting Error : The DATA_WIDTH is set to %s. Legal values is X8,X16,X32",DATA_WIDTH);
                     $finish;                  
          end
        endcase
        count_csn <= 0; 
    end



    always@(*) begin
        if(RW_SEL&&!CS_N) begin
            if(flg_rb_reg && !flg_rb_cmem)
                data_rb = data_rb_reg;
            else if(flg_rb_cmem && !flg_rb_reg)
                data_rb = reg_cmemor;
            else 
                data_rb = 32'hFFFF_FFFF;
        end
        else begin
            data_rb = 32'hFFFF_FFFF;
        end
    end


    ipal_e2_ispal CCS_IF_ISPAL (

        .rstn               (RST_N),
        .clk                (CLK), 
        .en                 (1'b1), 
        .m                  (ipal_m), 
        .din                (DI), 
        .cs_n               (CS_N), 
        .rdwr_n             (RW_SEL), 
        .flg_desync         (flg_desync),
        .data_rb            (data_rb), 

        .dout               (DO),  
        .data               (data), 
        .data_valid         (data_valid), 
        .re_rb              (re_rb));


///////////////////////////////packet processor////////////////////////////////////////

//    assign flg_read_tmp   = (data[28:27] == 2'b10);
//    assign flg_write_tmp  = (data[28:27] == 2'b01);
//    assign flg_type1      = (data[31:29] == 3'b101);
//    assign flg_type2      = (data[31:29] == 3'b010);
//    assign word_count_tmp = flg_type1 ? {5'd0, data[21:0]} : data[26:0];
//    assign flg_rb_reg = ~CS_N & RW_SEL & (~flg_rb_cmem);

    assign flg_read_tmp   = (data_valid==1)?(data[28:27] == 2'b10):flg_read_tmp;
    assign flg_write_tmp  = (data_valid==1)?(data[28:27] == 2'b01):flg_write_tmp;
    assign flg_type1      = (data_valid==1)?(data[31:29] == 3'b101):flg_type1;
    assign flg_type2      = (data_valid==1)?(data[31:29] == 3'b010):flg_type2;
    assign word_count_tmp = (flg_type1==1&&data_valid==1)?{5'd0, data[21:0]} : data[26:0]; 
    assign flg_rb_reg = ~CS_N & RW_SEL & (~flg_rb_cmem);


//State machine to indicate HEADER or DATA for current data
    always @(posedge CLK or negedge RST_N)begin
        if(RST_N == 1'b0)
            s <= HEADER;
        else if(data_valid||re_rb)
            s <= ns;
    end

    always @(*) begin
        case(s)
            HEADER: begin
                if(((flg_type1 || flg_type2) && (flg_read_tmp || flg_write_tmp)) && (word_count_tmp != 27'd0))
                    ns = DAT;
                else
                    ns = HEADER;
            end

            DAT:  begin
                if((data_valid && (word_count == 27'd0)) || (re_rb && (word_count_rb == 27'd0)))
                    ns = HEADER;
                else
                    ns = DAT;
            end
        endcase
    end

//get address
    always @(posedge CLK or negedge RST_N) begin
        if(RST_N == 1'b0)
            regaddr <= 5'd0;
        else if((data_valid || re_rb) && (s == HEADER) && flg_type1 && (flg_read_tmp || flg_write_tmp))
            regaddr <= data[26:22];
    end

//write flag
    always @(posedge CLK or negedge RST_N) begin
        if(RST_N == 1'b0)
            flg_write <= 1'b0;
        else if(data_valid) begin
            if((s == HEADER) && (flg_type1 || flg_type2) && flg_write_tmp && (word_count_tmp != 27'd0))
                flg_write <= 1'b1;
            else if(word_count == 27'd0)
                flg_write <= 1'b0;
        end
    end

//write operation count
    always @(posedge CLK or negedge RST_N) begin
        if(RST_N == 1'b0)
            word_count <= 27'd0;
        else if(data_valid) begin
            if((s == HEADER) && (flg_type1 || flg_type2) && flg_write_tmp && (word_count_tmp != 27'd0))
                word_count <= word_count_tmp - 1'b1;
            else if((s == DAT) && (word_count != 27'd0))
                word_count <= word_count - 1'b1;
            else
                word_count <= 27'd0;
        end
    end

//cmem readback count
    always @(posedge CLK or negedge RST_N) begin   
        if(RST_N == 1'b0)
            word_count_rb <= 27'd0;
        else if(/*re_rb && */(s == HEADER) && (flg_type1 || flg_type2) && flg_read_tmp && (word_count_tmp != 27'd0) && flg_rcmem&&data_valid==1)
            word_count_rb <= word_count_tmp - 1;
        else if((re_rb || flg_rb_reg) && (word_count_rb != 27'd0))
            word_count_rb <= word_count_rb - 1'b1;
    end

//cmem readback flag

    assign flg_rcmem   = (reg_cmd == 5'b00110);//read cmem, 
    always @(posedge CLK or negedge RST_N) begin
        if(RST_N == 1'b0)
            flg_rb_cmem <= 1'b0;
        else if(RW_SEL) begin
            if((flg_type1 || flg_type2) && flg_read_tmp && (word_count_rb != 27'd0) && flg_rcmem && (regaddr == 5'b0_0111))
                flg_rb_cmem <= 1'b1;
            //else if(word_count_rb == 27'd0)
                //flg_rb_cmem <= 1'b0;
            else if((re_rb || flg_rb_reg) && (word_count_rb == 27'd0))
                flg_rb_cmem <= 1'b0;
        end
        else begin
            flg_rb_cmem <= 1'b0;
        end
    end

    always @(posedge CLK or negedge RST_N) begin
        if(RST_N == 1'b0)
            flg_rb_cmem_d <= 1'b0;
        else 
            flg_rb_cmem_d <= flg_rb_cmem;
    end

    wire flg_rb_cmem_seu;
    assign flg_rb_cmem_seu = !flg_rb_cmem_d&flg_rb_cmem;

//command
    always@(*) begin
        if(!RST_N)
            reg_cmd = 0;
        else if(data_valid && flg_write && regaddr == 5'b00010)
            reg_cmd <= data[4:0];
    end

    assign flg_desync  = (reg_cmd == 5'b01011);//DESYNC


//////////////////////////////////////////////////reg array////////////////////////////////////////////////////////////////////

    always@(*) begin
        if(!RST_N) begin
            reg_crcr <= 0;
            reg_idr <= 0;
            reg_cmdr <= 0;
            reg_ctrl0r <= 0;
            reg_ctrl1r <= 0;
            reg_cmemir <= 0;
            reg_mfwriter <= 0;
            reg_ivr <= 0;
            reg_chainr <= 0;
            reg_adrr <= 0;
            reg_sbpir <= 0;
            reg_seur <= 0;
            reg_irstctrlr <= 0;
            reg_irstadrr <= 0;
            reg_watchdogr <= 0;
            reg_cmaskr <= 0;
            reg_keyr <= 0;
            reg_option0r <= 0;
            reg_option1r <= 0;
            reg_rcrr <= 0;
            reg_autr <= 0;
            reg_cmemor <= 32'hFFFF_FFFF;
            reg_seustatusr <= 0;
            reg_seuaddr <= 0;
            reg_seunaddr <= 0;
        end
        else begin
            if(data_valid && flg_write) begin
                case(regaddr)
                5'b00000 : reg_crcr <= data;
                5'b00001 : reg_idr <= IDCODE;
                5'b00010 : reg_cmdr <= data;
                5'b00011 : reg_ctrl0r <= data;
                5'b00100 : reg_ctrl1r <= data;
                5'b00101 : reg_cmemir <= data;
                5'b00110 : reg_mfwriter <= data;
                5'b01000 : reg_ivr <= data;
                5'b01010 : reg_chainr <= data;
                5'b01011 : begin 
                                reg_adrr <= data;
                                reg_adrr_seu <= data;
                           end
                5'b01100 : reg_sbpir <= data;
                5'b01101 : reg_seur <= data;
                5'b01111 : reg_irstctrlr <= data;
                5'b10000 : reg_irstadrr <= data;
                5'b10001 : reg_watchdogr <= data;
                5'b10111 : reg_cmaskr <= data;
                5'b11000 : reg_keyr <= data;
                5'b11001 : reg_option0r <= data;
                5'b11010 : reg_option1r <= data;
                5'b11011 : reg_rcrr <= data;
                5'b11110 : reg_autr <= data;
                endcase
            end
            else if(!CS_N && flg_rb_reg) begin
                case(regaddr)
                5'b00000 : data_rb_reg <= reg_crcr;
                5'b00001 : data_rb_reg <= IDCODE;
                5'b00010 : data_rb_reg <= reg_cmdr;
                5'b00011 : data_rb_reg <= 32'h0000_0010;//reg_ctrl0r;
                5'b00100 : data_rb_reg <= reg_ctrl1r;
                5'b00111 : data_rb_reg <= reg_cmemor;
                5'b01001 : data_rb_reg <= reg_statusr;
                5'b01011 : data_rb_reg <= reg_adrr;
                5'b01100 : data_rb_reg <= reg_sbpir;
                5'b01101 : data_rb_reg <= reg_seur;
                5'b01110 : data_rb_reg <= reg_seustatusr;
                5'b01111 : data_rb_reg <= reg_irstctrlr;
                5'b10000 : data_rb_reg <= reg_irstadrr;
                5'b10001 : data_rb_reg <= 32'h3FFF_FFFF;//reg_watchdogr;
                5'b10010 : data_rb_reg <= reg_hstatusr;
                5'b10111 : data_rb_reg <= reg_cmaskr;
                5'b11001 : data_rb_reg <= reg_option0r;
                5'b11010 : data_rb_reg <= reg_option1r;
                5'b11011 : data_rb_reg <= 32'h0360_0000;//reg_rcrr;
                5'b11110 : data_rb_reg <= reg_autr;
                5'b11101 : data_rb_reg <= reg_seuaddr;
                5'b11111 : data_rb_reg <= reg_seunaddr;
                default  : data_rb_reg <= 32'hFFFF_FFFF;
                endcase                
            end
        end                    
    end

////////////////////////////////////////////////cmem_e2////////////////////////////////////////////////


    assign cmemclk = CLK && (data_valid || re_rb);
    assign we = (flg_write == 1 && regaddr == 5'b00101 && reg_cmd == 5'b00100) ? 1'b1 : 1'b0;
    assign cmemtype = reg_adrr[26:25];
    assign addr_region = reg_adrr[24:20];
    assign addr_column = reg_adrr[17:10];
    assign addr_frame = reg_adrr[7:0];
    assign region0 = (addr_region == 5'd0) ? 1 : 0;
    assign region1 = (addr_region == 5'd1) ? 1 : 0;
    assign region2 = (addr_region == 5'd2) ? 1 : 0;
    assign region3 = (addr_region == 5'd3) ? 1 : 0;

    initial begin
        for(i = 0; i < 7328; i = i + 1)
            cmem[i] <= 0;
    end

    always@(posedge CLK or negedge RST_N) begin
        if(!RST_N) begin
            addr_word <= 0; 
            flg_frame_end <= 0;
            flg_column_end <= 0;
            flg_region_end <= 0;
            for(i = 0; i < 8000; i = i + 1)
                cmem[i] <= 0;
        end
        else if((we && data_valid) || (flg_rb_cmem && re_rb)) begin
            addr_word <= addr_word + 1;
            if(addr_word == 100) begin
                addr_word <= 0;   
                flg_frame_end <= 1;
                reg_adrr[7:0] <= reg_adrr[7:0] + 1;//addr_frame + 1
            end
            else
                flg_frame_end <= 0;
        end
    end

    always@(posedge flg_rcmem) begin
        if(seu_en)
            flg_frame_end = 1;
    end


    always@(negedge CLK) begin//CLK
            if(we && data_valid) begin
                    cmem[addr_row][(100 - addr_word)*32] <= reg_cmemir[0];
                    cmem[addr_row][(100 - addr_word)*32 + 1] <= reg_cmemir[1];
                    cmem[addr_row][(100 - addr_word)*32 + 2] <= reg_cmemir[2];
                    cmem[addr_row][(100 - addr_word)*32 + 3] <= reg_cmemir[3];
                    cmem[addr_row][(100 - addr_word)*32 + 4] <= reg_cmemir[4];
                    cmem[addr_row][(100 - addr_word)*32 + 5] <= reg_cmemir[5];
                    cmem[addr_row][(100 - addr_word)*32 + 6] <= reg_cmemir[6];
                    cmem[addr_row][(100 - addr_word)*32 + 7] <= reg_cmemir[7];
                    cmem[addr_row][(100 - addr_word)*32 + 8] <= reg_cmemir[8];
                    cmem[addr_row][(100 - addr_word)*32 + 9] <= reg_cmemir[9];
                    cmem[addr_row][(100 - addr_word)*32 + 10] <= reg_cmemir[10];
                    cmem[addr_row][(100 - addr_word)*32 + 11] <= reg_cmemir[11];
                    cmem[addr_row][(100 - addr_word)*32 + 12] <= reg_cmemir[12];
                    cmem[addr_row][(100 - addr_word)*32 + 13] <= reg_cmemir[13];
                    cmem[addr_row][(100 - addr_word)*32 + 14] <= reg_cmemir[14];
                    cmem[addr_row][(100 - addr_word)*32 + 15] <= reg_cmemir[15];
                    cmem[addr_row][(100 - addr_word)*32 + 16] <= reg_cmemir[16];
                    cmem[addr_row][(100 - addr_word)*32 + 17] <= reg_cmemir[17];
                    cmem[addr_row][(100 - addr_word)*32 + 18] <= reg_cmemir[18];
                    cmem[addr_row][(100 - addr_word)*32 + 19] <= reg_cmemir[19];
                    cmem[addr_row][(100 - addr_word)*32 + 20] <= reg_cmemir[20];
                    cmem[addr_row][(100 - addr_word)*32 + 21] <= reg_cmemir[21];
                    cmem[addr_row][(100 - addr_word)*32 + 22] <= reg_cmemir[22];
                    cmem[addr_row][(100 - addr_word)*32 + 23] <= reg_cmemir[23];
                    cmem[addr_row][(100 - addr_word)*32 + 24] <= reg_cmemir[24];
                    cmem[addr_row][(100 - addr_word)*32 + 25] <= reg_cmemir[25];
                    cmem[addr_row][(100 - addr_word)*32 + 26] <= reg_cmemir[26];
                    cmem[addr_row][(100 - addr_word)*32 + 27] <= reg_cmemir[27];
                    cmem[addr_row][(100 - addr_word)*32 + 28] <= reg_cmemir[28];
                    cmem[addr_row][(100 - addr_word)*32 + 29] <= reg_cmemir[29];
                    cmem[addr_row][(100 - addr_word)*32 + 30] <= reg_cmemir[30];
                    cmem[addr_row][(100 - addr_word)*32 + 31] <= reg_cmemir[31];
                end
        end
        always@(*) begin
                if(flg_rb_cmem && !CS_N) begin
                    reg_cmemor[0] <= cmem[addr_row][(100 - addr_word)*32];
                    reg_cmemor[1] <= cmem[addr_row][(100 - addr_word)*32 + 1];
                    reg_cmemor[2] <= cmem[addr_row][(100 - addr_word)*32 + 2];
                    reg_cmemor[3] <= cmem[addr_row][(100 - addr_word)*32 + 3];
                    reg_cmemor[4] <= cmem[addr_row][(100 - addr_word)*32 + 4];
                    reg_cmemor[5] <= cmem[addr_row][(100 - addr_word)*32 + 5];
                    reg_cmemor[6] <= cmem[addr_row][(100 - addr_word)*32 + 6];
                    reg_cmemor[7] <= cmem[addr_row][(100 - addr_word)*32 + 7];
                    reg_cmemor[8] <= cmem[addr_row][(100 - addr_word)*32 + 8];
                    reg_cmemor[9] <= cmem[addr_row][(100 - addr_word)*32 + 9];
                    reg_cmemor[10] <= cmem[addr_row][(100 - addr_word)*32 + 10];
                    reg_cmemor[11] <= cmem[addr_row][(100 - addr_word)*32 + 11];
                    reg_cmemor[12] <= cmem[addr_row][(100 - addr_word)*32 + 12];
                    reg_cmemor[13] <= cmem[addr_row][(100 - addr_word)*32 + 13];
                    reg_cmemor[14] <= cmem[addr_row][(100 - addr_word)*32 + 14];
                    reg_cmemor[15] <= cmem[addr_row][(100 - addr_word)*32 + 15];
                    reg_cmemor[16] <= cmem[addr_row][(100 - addr_word)*32 + 16];
                    reg_cmemor[17] <= cmem[addr_row][(100 - addr_word)*32 + 17];
                    reg_cmemor[18] <= cmem[addr_row][(100 - addr_word)*32 + 18];
                    reg_cmemor[19] <= cmem[addr_row][(100 - addr_word)*32 + 19];
                    reg_cmemor[20] <= cmem[addr_row][(100 - addr_word)*32 + 20];
                    reg_cmemor[21] <= cmem[addr_row][(100 - addr_word)*32 + 21];
                    reg_cmemor[22] <= cmem[addr_row][(100 - addr_word)*32 + 22];
                    reg_cmemor[23] <= cmem[addr_row][(100 - addr_word)*32 + 23];
                    reg_cmemor[24] <= cmem[addr_row][(100 - addr_word)*32 + 24];
                    reg_cmemor[25] <= cmem[addr_row][(100 - addr_word)*32 + 25];
                    reg_cmemor[26] <= cmem[addr_row][(100 - addr_word)*32 + 26];
                    reg_cmemor[27] <= cmem[addr_row][(100 - addr_word)*32 + 27];
                    reg_cmemor[28] <= cmem[addr_row][(100 - addr_word)*32 + 28];
                    reg_cmemor[29] <= cmem[addr_row][(100 - addr_word)*32 + 29];
                    reg_cmemor[30] <= cmem[addr_row][(100 - addr_word)*32 + 30];
                    reg_cmemor[31] <= cmem[addr_row][(100 - addr_word)*32 + 31];
                end
    end


    always@(negedge we) begin
        #0.1;
        $writememb("cmem.txt", cmem);
        addr_word <= 0;
    end

    always@(posedge flg_rb_cmem) begin
        $readmemb("cmem.txt", cmem);  
    end

    always@(negedge flg_rb_cmem) begin
        addr_word <= 0;
        reg_cmemor <= 32'hFFFF_FFFF;
    end


    always@(*)begin
        case(addr_region)
            0:  case (addr_column)
                    2, 3, 4, 6, 7, 8, 9, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 24, 25, 26, 27, 28, 29, 30, 31, 32, 34, 35, 36, 38, 39, 41, 42, 43, 45, 46, 48, 49, 50, 52, 53, 54, 55, 56, 57: begin //CLM
                        if(addr_frame < 36) begin
                            addr_row = 0 + 36* addr_column + addr_frame;
                            if(addr_frame == 35) begin
                                flg_column_end = 1;
                                flg_region_end = 0;                                
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0;
                            end
                        end
                        else if(addr_frame == 36) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end
                    5, 40, 47, 51: begin // DRM
                        if(addr_frame < 28) begin
                            addr_row = 0 + 36*addr_column + addr_frame;
                            if(addr_frame == 27) begin
                                flg_column_end = 1;
                                flg_region_end = 0;
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0;
                            end
                        end
                        else if(addr_frame == 28) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end    
                    10, 37, 44: begin //APM
                        if(addr_frame < 28) begin
                            addr_row = 0 + 36*addr_column + addr_frame;
                            if(addr_frame == 27) begin
                                flg_column_end = 1;
                                flg_region_end = 0;                
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0;
                            end
                        end
                        else if(addr_frame == 28) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;                        
                        end
                    end  
                    1: begin //IOL
                        if(addr_frame < 34) begin
                            addr_row = 0 + 36*addr_column + addr_frame;
                            if(addr_frame == 33) begin
                                flg_column_end = 1;
                                flg_region_end = 0;  
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0;
                            end
                        end
                        else if(addr_frame == 34) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end 
                    0: begin //IOB
                        if(addr_frame < 2) begin
                            addr_row = 0 + 36*addr_column + addr_frame;
                            if(addr_frame == 1) begin
                                flg_column_end = 1;
                                flg_region_end = 0;  
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0;
                            end
                        end
                        else if(addr_frame == 2) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;

                        end
                    end 

                    23, 33: begin //CLK or ADC
                        if(addr_frame < 28) begin
                            addr_row = 0 + 36*addr_column + addr_frame;
                            if(addr_frame == 27) begin
                                flg_column_end = 1;
                                flg_region_end = 0;  
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0;
                            end
                        end
                        else if(addr_frame == 28) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end 
                    58: begin // HSST
                        if(addr_frame < 28) begin
                            addr_row = 0 + 36*addr_column + addr_frame;
                            if(addr_frame == 27) begin
                                flg_column_end = 1;
                                flg_region_end = 1;  
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0;
                            end
                        end
                        else if(addr_frame == 28) begin
                                reg_adrr[7:0] = 0;
                                reg_adrr[17:10] = 0;
                                reg_adrr[24:20] = 1;
                        end
                    end 
                endcase
            1:  case(addr_column)
                    2, 3, 4, 6, 7, 8, 9, 11, 12, 14, 15, 16, 17, 18, 19, 20, 21, 22, 24, 25, 26, 28, 29, 31, 32, 33, 35, 36, 38, 39, 40, 42, 43, 44, 45, 46, 47:begin //CLM
                        if(addr_frame < 36) begin
                            addr_row = 36*59 + 36*addr_column + addr_frame;
                            if(addr_frame == 35) begin
                                flg_region_end = 0;
                                flg_column_end = 1;
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0;
                            end
                        end
                        else if(addr_frame == 36)begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end
                    5, 30, 37, 41: begin //DRM
                        if(addr_frame < 28) begin
                            addr_row = 36*59 + 36*addr_column + addr_frame;
                            if(addr_frame == 27) begin
                                flg_region_end = 0;
                                flg_column_end = 1;   
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0;     
                            end                       
                        end
                        else if(addr_frame == 28) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;                         
                        end
                    end
                    10, 27, 34: begin //APM
                        if(addr_frame < 28) begin
                            addr_row = 36*59 + 36*addr_column + addr_frame;
                            if(addr_frame == 27) begin
                                flg_region_end = 0;
                                flg_column_end = 1;    
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0;  
                            end

                        end
                        else if(addr_frame == 28) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;                      
                        end
                    end
                    1, 48: begin //IOL
                        if(addr_frame < 34) begin
                            addr_row = 36*59 + 36*addr_column + addr_frame;
                            if(addr_frame == 33) begin
                                flg_region_end = 0;
                                flg_column_end = 1;  
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0;  
                            end
                        end
                        else if(addr_frame == 34)begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1; 
                        end
                    end
                    0, 49: begin //IOB
                        if(addr_frame < 2) begin
                            addr_row = 36*59 + 36*addr_column + addr_frame;
                            if(addr_frame == 1) begin
                                if(addr_column == 49) begin
                                    flg_region_end = 1;
                                    flg_column_end = 1;  
                                end
                                else begin
                                    flg_region_end = 0;
                                    flg_column_end = 1;  
                                end
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0;  
                            end
                        end
                        else if(addr_frame == 2) begin
                            if(addr_column == 49) begin
                                reg_adrr[7:0] = 0;
                                reg_adrr[17:10] = 0;
                                reg_adrr[24:20] = 2;
                            end
                            else begin
                                reg_adrr[7:0] = 0;
                                reg_adrr[17:10] = reg_adrr[17:10] + 1;
                            end
                        end
                    end
                    13, 23: begin //CLK and ADC
                        if(addr_frame < 28) begin
                            addr_row = 36*59 + 36*addr_column + addr_frame;
                            if(addr_frame == 27) begin
                                flg_region_end = 0;
                                flg_column_end = 1;
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0;  
                            end
                        end
                        else if(addr_frame == 28) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end   
                    end             
                endcase
            2:  case(addr_column)
                    2, 3, 4, 6, 7, 8, 9, 11, 12, 14, 15, 16, 17, 18, 19, 20, 21, 22, 24, 25, 26, 28, 29, 31, 32, 33, 35, 36, 38, 39, 40, 42, 43, 44, 45, 46, 47:begin //CLM
                        if(addr_frame < 36) begin
                            addr_row = 36*(59 + 50) + 36*addr_column + addr_frame;
                            if(addr_frame == 35) begin
                                flg_region_end = 0;
                                flg_column_end = 1;
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0;
                            end
                        end
                        else if(addr_frame == 36)begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end
                    5, 30, 37, 41: begin //DRM
                        if(addr_frame < 28) begin
                            addr_row = 36*(59 + 50) + 36*addr_column + addr_frame;
                            if(addr_frame == 27) begin
                                flg_region_end = 0;
                                flg_column_end = 1; 
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0;    
                            end                        
                        end
                        else if(addr_frame == 28) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;                           
                        end
                    end
                    10, 27, 34: begin //APM
                        if(addr_frame < 28) begin
                            addr_row = 36*(59 + 50) + 36*addr_column + addr_frame;
                            if(addr_frame == 27) begin
                                flg_region_end = 0;
                                flg_column_end = 1;  
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0; 
                            end
                        end
                        else if(addr_frame == 28) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;                        
                        end
                    end
                    1, 48: begin //IOL
                        if(addr_frame < 34) begin
                            addr_row = 36*(59 + 50) + 36*addr_column + addr_frame;
                            if(addr_frame == 33) begin
                                flg_region_end = 0;
                                flg_column_end = 1;   
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0;  
                            end
                        end
                        else if(addr_frame == 34)begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end
                    0, 49: begin //IOB
                        if(addr_frame < 2) begin
                            addr_row = 36*(59 + 50) + 36*addr_column + addr_frame;
                            if(addr_frame == 1) begin
                                if(addr_column == 49) begin
                                    flg_region_end = 1;
                                    flg_column_end = 1;  
                                end
                                else begin
                                    flg_region_end = 0;
                                    flg_column_end = 1;  
                                end
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0;  
                            end
                        end
                        else if(addr_frame == 2) begin
                            if(addr_column == 49) begin
                                reg_adrr[7:0] = 0;
                                reg_adrr[17:10] = 0;
                                reg_adrr[24:20] = 3;
                            end
                            else begin
                                reg_adrr[7:0] = 0;
                                reg_adrr[17:10] = reg_adrr[17:10] + 1;
                            end
                        end
                    end
                    13, 23: begin //CLK and ADC
                        if(addr_frame < 28) begin
                            addr_row = 36*(59 + 50) + 36*addr_column + addr_frame;
                            if(addr_frame == 27) begin
                                flg_region_end = 0;
                                flg_column_end = 1;
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0;  
                            end
                        end
                        else if(addr_frame == 28) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end   
                    end             
                endcase

            3:  case (addr_column)
                    2, 3, 4, 6, 7, 8, 9, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 24, 25, 26, 27, 28, 29, 30, 31, 32, 34, 35, 36, 38, 39, 41, 42, 43, 45, 46, 48, 49, 50, 52, 53, 54, 55, 56, 57: begin //CLM
                        if(addr_frame < 36) begin
                            addr_row = 36*(59 + 50 + 50) + 36* addr_column + addr_frame;
                            if(addr_frame == 35) begin
                                flg_column_end = 1;
                                flg_region_end = 0;
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0;
                            end
                        end
                        else if(addr_frame == 36) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end
                    5, 40, 47, 51: begin // DRM
                        if(addr_frame < 28) begin
                            addr_row = 36*(59 + 50 + 50) + 36*addr_column + addr_frame;
                            if(addr_frame == 27) begin
                                flg_column_end = 1;
                                flg_region_end = 0;
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0;
                            end
                        end
                        else if(addr_frame == 28) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end    
                    10, 37, 44: begin //APM
                        if(addr_frame < 28) begin
                            addr_row = 36*(59 + 50 + 50) + 36*addr_column + addr_frame;
                            if(addr_frame == 27) begin
                                flg_column_end = 1;
                                flg_region_end = 0;  
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0;
                            end
                        end
                        else if(addr_frame == 28) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;                          
                        end
                    end  
                    1: begin //IOL
                        if(addr_frame < 34) begin
                            addr_row = 36*(59 + 50 + 50) + 36*addr_column + addr_frame;
                            if(addr_frame == 33) begin
                                flg_column_end = 1;
                                flg_region_end = 0;  
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0;
                            end
                        end
                        else if(addr_frame == 34) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end 
                    0: begin //IOB
                        if(addr_frame < 2) begin
                            addr_row = 36*(59 + 50 + 50) + 36*addr_column + addr_frame;
                            if(addr_frame == 1) begin
                                flg_column_end = 1;
                                flg_region_end = 0;  
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0;
                            end
                        end
                        else if(addr_frame == 2) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end 

                    23, 33: begin //CLK or ADC
                        if(addr_frame < 28) begin
                            addr_row = 36*(59 + 50 + 50) + 36*addr_column + addr_frame;
                            if(addr_frame == 27) begin
                                flg_column_end = 1;
                                flg_region_end = 0;  
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0;
                            end
                        end
                        else if(addr_frame == 28) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end 
                    58: begin // HSST
                        if(addr_frame < 28) begin
                            addr_row = 36*(59 + 50 + 50) + 36*addr_column + addr_frame;
                            if(addr_frame == 27) begin
                                flg_column_end = 1;
                                flg_region_end = 1;  
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0;
                            end
                        end
                        else if(addr_frame == 28) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = 0;
                            reg_adrr[24:20] = 0;
                        end
                    end 
                endcase
        endcase
    end    

///////////////////////////////////////////rb_crc///////////////////////////////////////////////////
    assign rbcrc_en = reg_seur[0];
    assign seu_en = (cmemtype == 2'b00) ? reg_seur[1] : 0;
    assign flg_rrbcrc = (rbcrc_en && (reg_cmd == 5'b01101)) ? 1 : 0;//reset readback CRC
    assign flg_rbcrc = (rbcrc_en && (reg_cmd == 5'b01110)) ? 1 : 0;//readback CRC

    ipal_e2_rbcrc CCS_RBCRC(

        .rstn               (RST_N),
        .clk                (CLK & (re_rb | data_valid)),
        .rbcrc_en           (rbcrc_en),
        .data               (reg_cmemor),
        .data_valid         (flg_rb_cmem),//
        .flg_rrbcrc         (flg_rrbcrc),
        .flg_rbcrc          (flg_rbcrc),
        .irstn              (RST_N),
        .iclk               (CLK & (re_rb | data_valid)),

        .rbcrc_err          (RBCRC_ERR),
        .rbcrc_valid        (RBCRC_VALID)
    );

///////////////////////////////////////seu///////////////////////////////////////////////////////////


    wire seu_we;
    wire ecc_valid_tmp;
    wire seu_clk;
    wire [31:0] seu_din;
    wire [6:0] seu_addr;
    reg  seu_we_d;
    reg  seu_we_d2;
    //reg  [6:0] addr_word_d;
    reg re_rb_d;
    reg re_rb_d2;
    reg re_rb_d3;
    reg re_rb_d4;
    wire clk_div;
    always@(posedge CLK or negedge RST_N) begin
        if(!RST_N) begin
            re_rb_d <= 0;
            re_rb_d2 <= 0;
            re_rb_d3 <= 0;
            re_rb_d4 <= 0;
        end
        else begin
            re_rb_d <= re_rb;
            re_rb_d2 <= re_rb_d;
            re_rb_d3 <= re_rb_d2;
            re_rb_d4 <= re_rb_d3;
        end
    end
    assign clk_div = (DATA_WIDTH == "X16") ? (re_rb | re_rb_d2) : (re_rb | re_rb_d4);
    assign seu_we = (DATA_WIDTH == "X32") ? flg_rb_cmem : re_rb;    
    assign seu_clk = (DATA_WIDTH == "X32") ? CLK : flg_rb_cmem ? clk_div : CLK;
    always@(negedge RST_N or posedge ECC_VALID or negedge CS_N) begin
        if(!RST_N) begin
            seu_we_d <= 0;
        end
        else if(ECC_VALID)
            seu_we_d <= 0;
        else begin
            if(!CS_N && RW_SEL && addr_word == 0 && seu_en)
                #0.1 seu_we_d <= 1;//seu_we;
            //else
                //seu_we_d <= 0;

            //addr_word_d <= addr_word;
        end
    end


    assign #0.1 seu_addr = addr_word;
    assign #0.1 seu_din = reg_cmemor;

    ipal_e2_secded CCS_SECDED (
        .rstn               (RST_N),
        .clk                (seu_clk),//seu_clk
        .en                 (seu_en),
        .addr               (seu_addr),//addr_word_d
        .we                 (seu_we_d),
        .din                (seu_din),//reg_cmemor

        .flg_ecc_over       (ecc_valid_tmp),
        .flg_sec            (serror),
        .flg_ded            (derror),
        .index              (ECC_INDEX)
    );
    reg ecc_valid_tmp_d;
    wire ecc_valid_tmp_p;
    always@(posedge CLK or negedge RST_N) begin
        if(!RST_N)
            ecc_valid_tmp_d <= 0;
        else
            ecc_valid_tmp_d <= ecc_valid_tmp;
    end
    assign ecc_valid_tmp_p = !ecc_valid_tmp_d&ecc_valid_tmp;
    assign ECC_VALID = ecc_valid_tmp_p&flg_rcmem; 

    always@(posedge CLK or negedge RST_N) begin
        if(!RST_N) begin
            serror_d <= 0;
            derror_d <= 0;
        end
        else begin
            serror_d <= serror;
            derror_d <= derror;
        end
    end

    assign SERROR = serror; //(!serror_d && serror) ? 1 : 0;
    assign DERROR = derror; //(!derror_d && derror) ? 1 : 0;



    
    reg serror_reg;
    reg derror_reg;
    reg [11:0]ecc_index_reg;
    reg ecc_valid_reg;

    always@(posedge ECC_VALID or negedge RST_N) begin
        if(!RST_N) begin
            serror_reg <= 0;
            derror_reg <= 0;
            ecc_index_reg <= 0;
            ecc_valid_reg <= 0;
        end
        else begin
            serror_reg <= SERROR;
            derror_reg <= DERROR;
            ecc_index_reg <= ECC_INDEX;
            ecc_valid_reg <= 1'b1;
        end
    end

    reg drcfg_over_reg;
    reg drcfg_err_reg;

    always@(posedge DRCFG_OVER or negedge RST_N) begin
        if(!RST_N) begin
            drcfg_over_reg <= 0;
            drcfg_err_reg <= 0;
        end
        else begin
            drcfg_over_reg <= DRCFG_OVER;
            drcfg_err_reg <= DRCFG_ERR;
        end
    end


    always@(*) begin
        if(RST_N) begin
            reg_seustatusr[31:17] = 0;
            reg_seustatusr[16] = drcfg_over_reg;
            reg_seustatusr[15] = drcfg_err_reg;
            reg_seustatusr[14:3] = ecc_index_reg;
            reg_seustatusr[2] = derror_reg;
            reg_seustatusr[1] = serror_reg;
            reg_seustatusr[0] = ecc_valid_reg;
        end
    end

/////////////////////////////////////////prcfg and drcfg/////////////////////////////////////////


    assign flg_prcfgen    = (reg_cmd == 5'b10100);
    assign flg_prcfgdis   = (reg_cmd == 5'b10101);
    assign flg_drcfgen    = (reg_cmd == 5'b10110);
    assign flg_drcfgdis   = (reg_cmd == 5'b10111);
    assign flg_rstcrc     = (reg_cmd == 5'b00001);
 
    assign PRCFG_OVER     = prcfg_over;
    assign PRCFG_ERR      = PRCFG_OVER ? prcfg_err : 0;
    assign DRCFG_OVER     = drcfg_over;
    assign DRCFG_ERR      = DRCFG_OVER ? drcfg_err : 0;

    always @(posedge CLK or negedge RST_N) begin
        if(RST_N == 1'b0)
            prcfg_en <= 1'b0;
        else if(flg_prcfgen)
            prcfg_en <= 1'b1;
        else if(flg_prcfgdis)
            prcfg_en <= 1'b0;
    end

    always@(posedge CLK or negedge RST_N) begin
        if(!RST_N)
            drcfg_en <= 0;
        else if(flg_drcfgen)
            drcfg_en <= 1;
        else if(flg_drcfgdis)
            drcfg_en <= 0;
    end

    always @(posedge CLK or negedge RST_N) begin
        if(RST_N == 1'b0)
            prcfg_en_d <= 1'b0;
        else
            prcfg_en_d <= prcfg_en;
    end

    always@(posedge CLK or negedge RST_N) begin
        if(!RST_N)
            drcfg_en_d <= 0;
        else
            drcfg_en_d <= drcfg_en;
    end

    always @(posedge CLK or negedge RST_N) begin
        if(RST_N == 1'b0)
            prcfg_over <= 1'b0;
        else if(!prcfg_en && prcfg_en_d)
            prcfg_over <= 1'b1;
        else
            prcfg_over <= 1'b0;
    end

    always@(posedge CLK or negedge RST_N) begin
        if(!RST_N)
            drcfg_over <= 0;
        else if(!drcfg_en && drcfg_en_d)
            drcfg_over <= 1;
        else 
            drcfg_over <= 0;
    end



    ipal_e2_crc  crc (

        .rstn                   (RST_N),
        .clk                    (CLK),
        
        .regaddr                (regaddr),
        .id_err                 (1'b0),
        .crc_disable            (reg_option1r[0]),//
        .data                   (data),
        .data_valid             (data_valid),
        .flg_write              (flg_write),
        .flg_rstcrc             (flg_rstcrc),//
        .reg_crc                (reg_crcr),
        .prcfg_en               (prcfg_en),
        .prcfg_err              (prcfg_err),
        .drcfg_en               (drcfg_en),
        .drcfg_err              (drcfg_err),
        .crc_err                (crc_err)//floating

);
/////////////////////////////////////////FRAME\COLUMN\REGION/////////////////////////////////////////
    reg [7:0] addr_frame_seu;
    reg [7:0] addr_column_seu;
    reg [4:0] addr_region_seu;
    initial begin
        addr_frame_seu <= 0;
        addr_column_seu <= 0;
        addr_region_seu <= 0;
        reg_adrr_seu <= 0;
    end
    always@(reg_adrr) begin
        if(seu_en) begin
            addr_frame_seu <= reg_adrr_seu[7:0];
            addr_column_seu <= reg_adrr_seu[17:10];
            addr_region_seu <= reg_adrr_seu[24:20];
        end
    end

    //assign SEU_FRAME_ADDR = seu_en ? reg_adrr_seu[7:0] : 0;
    //assign SEU_COLUMN_ADDR = seu_en ? reg_adrr_seu[17:10] : 0;
    //assign SEU_REGION_ADDR = seu_en ? reg_adrr_seu[24:20] : 0;


    //assign SEU_FRAME_NADDR = seu_en ? (flg_column_end ? 0: SEU_FRAME_ADDR + flg_frame_end) : 0;
    //assign SEU_COLUMN_NADDR = seu_en ? (flg_region_end ? 0: SEU_COLUMN_ADDR + flg_column_end) : 0;
    //assign SEU_REGION_NADDR = seu_en ? (SEU_REGION_ADDR != 3 ? SEU_REGION_ADDR + flg_region_end : 0) : 0;


    initial begin
        SEU_REGION_ADDR = 0;
        SEU_COLUMN_ADDR = 0;
        SEU_FRAME_ADDR = 0;
        SEU_REGION_NADDR = 0;
        SEU_COLUMN_NADDR = 0;
        SEU_FRAME_NADDR = 0;   
    end

    always@(posedge CLK or negedge RST_N) begin
        if(!RST_N) begin
            SEU_REGION_ADDR = 0;
            SEU_COLUMN_ADDR = 0;
            SEU_FRAME_ADDR = 0;

            SEU_REGION_NADDR = 0;
            SEU_COLUMN_NADDR = 0;
            SEU_FRAME_NADDR = 0;
        end
        else if(flg_rb_cmem_seu && addr_word == 0)begin
            SEU_FRAME_ADDR = seu_en ? reg_adrr[7:0] : 0;
            SEU_COLUMN_ADDR = seu_en ? reg_adrr[17:10] : 0;
            SEU_REGION_ADDR = seu_en ? reg_adrr[24:20] : 0;

            SEU_FRAME_NADDR = seu_en ? (flg_column_end ? 0: SEU_FRAME_ADDR + flg_frame_end) : 0;
            SEU_COLUMN_NADDR = seu_en ? (flg_region_end ? 0: SEU_COLUMN_ADDR + flg_column_end) : 0;
            SEU_REGION_NADDR[1:0] = seu_en ? SEU_REGION_ADDR + flg_region_end : 0;  
        end
    end

    always@(*) begin
        reg_seuaddr <= {10'b0, SEU_REGION_ADDR, SEU_COLUMN_ADDR, SEU_FRAME_ADDR};
        reg_seunaddr <= {10'b0, SEU_REGION_NADDR, SEU_COLUMN_NADDR, SEU_FRAME_NADDR};
    end
//synthesis translate_on
endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_DLATCH_E.v
//
// Functional description: D-type latch with enable
//
// Parameter description:
//      INIT: init value
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_DLATCH_E
#(
    parameter GRS_EN = "TRUE",
    parameter INIT = 1'b0
) (
    output reg Q,
    input wire D,
    input wire G, GE
);

    wire grs_n;
    wire RS;

    tri1 grsnet = GRS_INST.GRSNET;
    assign grs_n=(GRS_EN=="TRUE")?grsnet:1'b1;

    not (RS, grs_n);

    initial Q = 1'bx;

    always @(D or G or GE or RS) begin
        if (RS)
            Q <= 1'b0;
        else if (G && GE)
            Q <= D;
    end

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_DRM9K_E1.v
//
// Functional description:
//
// Parameter  description:
//
// Port description:
//
// Revision history:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_DRM9K_E1
#(
    parameter GRS_EN = "TRUE",
    parameter [2:0] CSA_MASK = 3'b000,
    parameter [2:0] CSB_MASK = 3'b000,
    parameter integer DATA_WIDTH_A = 9,
    parameter integer DATA_WIDTH_B = 9,
    parameter WRITE_MODE_A = "NORMAL_WRITE",
    parameter WRITE_MODE_B = "NORMAL_WRITE",
    parameter integer DOA_REG = 0,
    parameter integer DOB_REG = 0,
    parameter integer DOA_REG_CLKINV = 0,
    parameter integer DOB_REG_CLKINV = 0,
    parameter [8:0] RSTA_VAL = 9'b000000000,
    parameter [8:0] RSTB_VAL = 9'b000000000,
    parameter RST_TYPE = "SYNC",
    parameter RAM_MODE = "TRUE_DUAL_PORT",
    parameter RAM_CASCADE = "NONE",
    parameter [287:0] INIT_00 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_01 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_02 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_03 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_04 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_05 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_06 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_07 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_08 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_09 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_10 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_11 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_12 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_13 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_14 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_15 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_16 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_17 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_18 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_19 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_FILE = "NONE",
    parameter integer BLOCK_X = 0,
    parameter integer BLOCK_Y = 0,
    parameter integer RAM_DATA_WIDTH = 9,
    parameter integer RAM_ADDR_WIDTH = 10,
    parameter INIT_FORMAT = "BIN"
) (
    output [8:0] DOA,
    output [8:0] DOB,
    input [8:0] DIA,
    input [8:0] DIB,
    input [13:0] ADDRA,
    input ADDRA_HOLD,
    input [13:0] ADDRB,
    input ADDRB_HOLD,
    input [2:0] CSA,
    input [2:0] CSB,
    input [1:0] BWEA,
    input CLKA,
    input CLKB,
    input CEA,
    input CEB,
    input WEA,
    input WEB,
    input ORCEA,
    input ORCEB,
    input RSTA,
    input RSTB,
    input CINA,
    input CINB,
    output COUTA,
    output COUTB
);

    localparam  BLOCK_DEPTH = 2**(DATA_WIDTH_A == 1 ? 13 :
                                  DATA_WIDTH_A == 2 ? 12 :
                                  DATA_WIDTH_A == 4 ? 11 :
                                  DATA_WIDTH_A <= 9 ? 10 : 9);

    localparam  BLOCK_WIDTH =   DATA_WIDTH_A;             //block memory data width

    localparam MEM_SIZE = 9216;
    localparam width_a = (DATA_WIDTH_A == 18) ? 9 : (DATA_WIDTH_A == 16) ? 8 : DATA_WIDTH_A;
    localparam width_b = (DATA_WIDTH_B == 18) ? 9 : (DATA_WIDTH_B == 16) ? 8 : DATA_WIDTH_B;

    integer  cnt;
    reg [9-1:0] mem [MEM_SIZE/9-1:0];

    reg csa_reg = 1'b0, csb_reg = 1'b0;
    reg [13:0] ada_reg = 13'b0, adb_reg = 13'b0;
    reg [8:0] da_reg = 9'b0, db_reg = 9'b0;
    reg wea_reg = 1'b0, web_reg = 1'b0;
    reg [1:0] bea_reg;
    wire write_en_a, write_en_b, read_en_a, read_en_b;

    reg [8:0] a_out;
    reg [8:0] a_out_reg;
    reg [8:0] b_out;
    reg [8:0] b_out_reg;

    wire grs, rsta_grs, rstb_grs;
    wire rsta_grs_sync;
    wire rstb_grs_sync;
    wire rsta_grs_async;
    wire rstb_grs_async;
    
    reg [8:0] doa;
    reg [8:0] dob;

    reg [1:0] cas_en;
    wire cas_inta,cas_intb;
    reg  cas_sela,cas_selb;
    wire [8:0] a_out_mux;
    wire [8:0] b_out_mux;
    wire CLKA_for_or,CLKB_for_or;
    wire rsta_int,rstb_int;

    initial begin
        doa = RSTA_VAL;
        dob = RSTB_VAL;
        a_out = RSTA_VAL[width_a-1:0];
        a_out_reg = RSTA_VAL;
        b_out = RSTB_VAL[width_b-1:0];
        b_out_reg = RSTB_VAL;
    end

// synthesis translate_off

   reg [RAM_DATA_WIDTH-1:0] ini_mem [2**RAM_ADDR_WIDTH-1:0];
   integer p;
   initial
   begin
      if(INIT_FILE != "NONE")
      begin
          if(INIT_FORMAT == "BIN")
              $readmemb(INIT_FILE,ini_mem);
          else
              $readmemh(INIT_FILE,ini_mem);
          for(p=0;p<20;p=p+1)
              $display("ini_mem[%d] = %b",p,ini_mem[p]);
      end
   end
///////////////////
// parameter check
///////////////////
    initial begin
        case (DATA_WIDTH_A)
            1, 2, 4, 8, 16: begin
                case (DATA_WIDTH_B)
                    1, 2, 4, 8, 16:  ; //null
                    default: begin
                        $display("ERROR: GTP_DRM9K_E1 instance %m parameter DATA_WIDTH_B:%d is illegal. The legal values are 1,2,4,8 or 16.",DATA_WIDTH_B);
                        $finish;
                    end
                endcase
            end
            9, 18: begin
                case (DATA_WIDTH_B)
                    9, 18:    ; //null
                    default: begin
                        $display("ERROR: GTP_DRM9K_E1 instance %m parameter DATA_WIDTH_B:%d is illegal. The legal values are 9 or 18.",DATA_WIDTH_B);
                        $finish;
                    end
                endcase
            end
            default: begin
                $display("ERROR: GTP_DRM9K_E1 instance %m parameter DATA_WIDTH_A:%d is illegal. The legal values are 1,2,4,8,9,16 or 18.",DATA_WIDTH_A);
                $finish;
            end
        endcase

        case (WRITE_MODE_A)
            "NORMAL_WRITE",
            "TRANSPARENT_WRITE",
            "READ_BEFORE_WRITE":    ; //null 
            default: begin
                $display("ERROR: GTP_DRM9K_E1 instance %m parameter WRITE_MODE_A: %s is illegal. The legal values are NORMAL_WRITE,TRANSPARENT_WRITE or READ_BEFORE_WRITE.", WRITE_MODE_A);
                $finish;
            end
        endcase

        case (WRITE_MODE_B)
            "NORMAL_WRITE",
            "TRANSPARENT_WRITE",
            "READ_BEFORE_WRITE":    ; //null  
            default: begin
                $display("ERROR: GTP_DRM9K_E1 instance %m parameter WRITE_MODE_B: %s is illegal. The legal values are NORMAL_WRITE,TRANSPARENT_WRITE or READ_BEFORE_WRITE.", WRITE_MODE_B);
                $finish;
            end
        endcase

        case (DOA_REG)
            0,1:     ;//null
            default: begin
                $display("ERROR: GTP_DRM9K_E1 instance %m parameter DOA_REG: %s is illegal. The legal values are 0 or 1.", DOA_REG);
                $finish;
            end
        endcase

        case (DOB_REG)
            0,1:     ;//null
            default: begin
                $display("ERROR: GTP_DRM9K_E1 instance %m parameter DOB_REG: %s is illegal. The legal values are 0 or 1.", DOB_REG);
                $finish;
            end
        endcase

        case (DOA_REG_CLKINV)
            0,1:     ;//null
            default: begin
                $display("ERROR: GTP_DRM9K_E1 instance %m parameter DOA_REG_CLKINV: %s is illegal. The legal values are 0 or 1.", DOA_REG_CLKINV);
                $finish;
            end
        endcase

        case (DOB_REG_CLKINV)
            0,1:     ;//null
            default: begin
                $display("ERROR: GTP_DRM9K_E1 instance %m parameter DOB_REG_CLKINV: %s is illegal. The legal values are 0 or 1.", DOB_REG_CLKINV);
                $finish;
            end
        endcase

        case (RST_TYPE)
            "ASYNC",
            "SYNC":     ;//null
            default: begin
                $display("ERROR: GTP_DRM9K_E1 instance %m parameter RST_TYPE: %s is illegal. The legal values are ASYNC or SYNC.", RST_TYPE);
                $finish;
            end
        endcase

        case (RAM_MODE)
            "ROM",
            "SINGLE_PORT":      ;//null
            "SIMPLE_DUAL_PORT": begin
                if (DATA_WIDTH_A < 16 && WRITE_MODE_A != "NORMAL_WRITE") begin
                    $display("Warrning: GTP_DRM9K_E1 instance %m suggest to use TRUE_DUAL_PORT RAM_MODE if DATA_WIDTH_A and WRITE_MODE_A: %d,%s.",DATA_WIDTH_A,WRITE_MODE_A);
                end
            end
            "TRUE_DUAL_PORT": begin
                if (DATA_WIDTH_A > 18 || DATA_WIDTH_B > 18) begin
                    $display("ERROR: GTP_DRM9K_E1 instance %m parameter DATA_WIDTH_A and DATA_WIDTH_B in TRUE_DUAL_PORT MODE:%d,%d is illegal. The legal values are 1,2,4,8,9,16 or 18.",DATA_WIDTH_A,DATA_WIDTH_B);
                    $finish;
                end
            end
            default: begin
                $display("ERROR: GTP_DRM9K_E1 instance %m parameter RAM_MODE value: %s is illegal. The legal values are ROM or SINGLE_PORT, SIMPLE_DUAL_PORT or TRUE_DUAL_PORT.", RAM_MODE);
                $finish;
            end
        endcase
        
        case (RAM_CASCADE)
            "NONE": begin
                cas_en = 2'b00;
            end
            "LOWER": begin
                if (DATA_WIDTH_A != 1 || DATA_WIDTH_B != 1) begin
                    $display("ERROR: GTP_DRM9K_E1 instance %m parameter DATA_WIDTH_A and DATA_WIDTH_B:%s,%s in CASCADING MODE:%s are illegal, then DATA_WIDTH_A and DATA_WIDTH_B have to be set to 1.",DATA_WIDTH_A,DATA_WIDTH_B,RAM_CASCADE);
                    $finish;
                end
                cas_en = 2'b01;
            end
            "UPPER": begin
                if (DATA_WIDTH_A != 1 || DATA_WIDTH_B != 1) begin
                    $display("ERROR: GTP_DRM9K_E1 instance %m parameter DATA_WIDTH_A and DATA_WIDTH_B:%s,%s in CASCADING MODE:%s are illegal, then DATA_WIDTH_A and DATA_WIDTH_B have to be set to 1.",DATA_WIDTH_A,DATA_WIDTH_B,RAM_CASCADE);
                    $finish;
                end
                cas_en = 2'b11;
            end
            default: begin
                $display("ERROR: GTP_DRM9K_E1 instance %m parameter RAM_CASCADE: %s is illegal, the legal values are NONE,LOWER or UPPER", RAM_CASCADE);
                $finish;
            end
        endcase
    end

/////////////////
// initialization
/////////////////

    initial begin
        if (INIT_FILE == "NONE") begin
            for (cnt = 0; cnt < 32; cnt = cnt + 1) begin
                mem[32*0 + cnt] = INIT_00[cnt*9 +: 9];
                mem[32*1 + cnt] = INIT_01[cnt*9 +: 9];
                mem[32*2 + cnt] = INIT_02[cnt*9 +: 9];
                mem[32*3 + cnt] = INIT_03[cnt*9 +: 9];
                mem[32*4 + cnt] = INIT_04[cnt*9 +: 9];
                mem[32*5 + cnt] = INIT_05[cnt*9 +: 9];
                mem[32*6 + cnt] = INIT_06[cnt*9 +: 9];
                mem[32*7 + cnt] = INIT_07[cnt*9 +: 9];
                mem[32*8 + cnt] = INIT_08[cnt*9 +: 9];
                mem[32*9 + cnt] = INIT_09[cnt*9 +: 9];
                mem[32*10 + cnt] = INIT_0A[cnt*9 +: 9];
                mem[32*11 + cnt] = INIT_0B[cnt*9 +: 9];
                mem[32*12 + cnt] = INIT_0C[cnt*9 +: 9];
                mem[32*13 + cnt] = INIT_0D[cnt*9 +: 9];
                mem[32*14 + cnt] = INIT_0E[cnt*9 +: 9];
                mem[32*15 + cnt] = INIT_0F[cnt*9 +: 9];
                mem[32*16 + cnt] = INIT_10[cnt*9 +: 9];
                mem[32*17 + cnt] = INIT_11[cnt*9 +: 9];
                mem[32*18 + cnt] = INIT_12[cnt*9 +: 9];
                mem[32*19 + cnt] = INIT_13[cnt*9 +: 9];
                mem[32*20 + cnt] = INIT_14[cnt*9 +: 9];
                mem[32*21 + cnt] = INIT_15[cnt*9 +: 9];
                mem[32*22 + cnt] = INIT_16[cnt*9 +: 9];
                mem[32*23 + cnt] = INIT_17[cnt*9 +: 9];
                mem[32*24 + cnt] = INIT_18[cnt*9 +: 9];
                mem[32*25 + cnt] = INIT_19[cnt*9 +: 9];
                mem[32*26 + cnt] = INIT_1A[cnt*9 +: 9];
                mem[32*27 + cnt] = INIT_1B[cnt*9 +: 9];
                mem[32*28 + cnt] = INIT_1C[cnt*9 +: 9];
                mem[32*29 + cnt] = INIT_1D[cnt*9 +: 9];
                mem[32*30 + cnt] = INIT_1E[cnt*9 +: 9];
                mem[32*31 + cnt] = INIT_1F[cnt*9 +: 9];
            end
        end
        else  begin      // INIT_FILE 
            case(DATA_WIDTH_A)
                1: begin  //DRM TYPE 8K*1
                   for(cnt=0; cnt<1024;cnt = cnt+1)
                       mem[cnt][7:0] = {ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*8+7][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*8+6][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*8+5][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*8+4][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*8+3][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*8+2][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*8+1][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*8][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH]};
                end
                2: begin //DRM TYPE 4K*2
                   for(cnt=0; cnt<1024;cnt = cnt+1)
                       mem[cnt][7:0] = {ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*4+3][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*4+2][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*4+1][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*4][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH]};
                end
                4: begin //DRM TYPE 2K*4
                   for(cnt=0; cnt<1024;cnt = cnt+1)
                       {mem[cnt][7:0]} = {ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*2+1][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                          ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*2][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH]};
                end
                8: begin //DRM TYPE 1K*8
                   for(cnt=0; cnt<1024;cnt = cnt+1)
                       mem[cnt][7:0] = ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH];
                end
                9: begin //DRM TYPE 1K*9
                   for(cnt=0; cnt<1024;cnt = cnt+1)
                       mem[cnt] = ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH];
                end
                16:begin //DRM TYPE 512*16
                   for(cnt=0; cnt<512;cnt = cnt+1)
                       {mem[cnt*2+1][7:0], mem[cnt*2][7:0]} = ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH];
                end
                18:begin //DRM TYPE 512*18
                   for(cnt=0; cnt<512;cnt = cnt+1)
                       {mem[cnt*2+1], mem[cnt*2]} = ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH];
                end
            endcase
        end
    end

    always @(posedge CLKA) begin
        if (CEA) begin
            // high to hold the address
            if (ADDRA_HOLD == 1'b0) begin
                ada_reg <= ADDRA;
                csa_reg <= CSA == CSA_MASK;
                bea_reg <= BWEA;
            end
            da_reg[8:0] <= DIA[8:0];
            wea_reg <= WEA;
        end
    end

    always @(posedge CLKB) begin
        if (CEB) begin
            // high to hold the address
            if (ADDRB_HOLD == 1'b0) begin
                adb_reg <= ADDRB;
                csb_reg <= CSB == CSB_MASK;
            end
                web_reg <= WEB;
        end
    end
    ///////////////////
    // task & function
    ///////////////////
    function [DATA_WIDTH_A-1:0] mem_read_a;
        input [12:0]  addr;
    begin
        case (DATA_WIDTH_A)
            1: mem_read_a = mem[addr[12:3]][addr[2:0]];
            2: mem_read_a = mem[addr[12:3]][addr[2:1]*2 +: 2];
            4: mem_read_a = mem[addr[12:3]][addr[2]*4 +: 4];
            8: mem_read_a = mem[addr[12:3]][7:0];
            9: mem_read_a = mem[addr[12:3]];
            default:      ;//null 
        endcase
    end
    endfunction

    function [DATA_WIDTH_B-1:0] mem_read_b;
        input [12:0] addr;
    begin
        case (DATA_WIDTH_B)
            1: mem_read_b = mem[addr[12:3]][addr[2:0]];
            2: mem_read_b = mem[addr[12:3]][addr[2:1]*2 +: 2];
            4: mem_read_b = mem[addr[12:3]][addr[2]*4 +: 4];
            8: mem_read_b = mem[addr[12:3]][7:0];
            9: mem_read_b = mem[addr[12:3]];
            16: mem_read_b = {mem[addr[12:4]*2+1][7:0], mem[addr[12:4]*2][7:0]};
            18: mem_read_b = {mem[addr[12:4]*2+1],      mem[addr[12:4]*2]};
            default:      ;//null
        endcase
    end
    endfunction

    task mem_write_a;
        input [12:0] addr;
        input [17:0] data;
        input [1:0]  byte_en;
    begin
        case (DATA_WIDTH_A)
            1: mem[addr[12:3]][addr[2:0]] = data[0];
            2: mem[addr[12:3]][addr[2:1]*2 +: 2] = data[1:0];
            4: mem[addr[12:3]][addr[2]*4 +: 4] = data[3:0];
            8: mem[addr[12:3]][7:0] = data[7:0];
            9: mem[addr[12:3]] = data[8:0];
            16: begin
                if (byte_en[1])
                    mem[addr[12:4]*2+1][7:0] = data[16:9];
                if (byte_en[0])
                    mem[addr[12:4]*2][7:0]   = data[7:0];
            end
            18: begin
                if (byte_en[1])
                    mem[addr[12:4]*2+1] = data[17:9];
                if (byte_en[0])
                    mem[addr[12:4]*2]   = data[8:0];
            end
            default:     ;//null
        endcase
    end
    endtask

    task mem_write_b;
        input [12:0] addr;
        input [8:0] data;
    begin
        case (DATA_WIDTH_B)
            1: mem[addr[12:3]][addr[2:0]] = data[0];
            2: mem[addr[12:3]][addr[2:1]*2 +: 2] = data[1:0];
            4: mem[addr[12:3]][addr[2]*4 +: 4] = data[3:0];
            8: mem[addr[12:3]][7:0] = data[7:0];
            9: mem[addr[12:3]] = data[8:0];
            default:     ;//null
        endcase
    end
    endtask

    ///////////////
    // memory core
    ///////////////
reg CLKA_active;
reg CLKB_active;
initial begin
  CLKA_active = 1'b0;
  CLKB_active = 1'b0;
end
always @(posedge CLKA) begin
   if (CEA) begin
      CLKA_active <= 1'b1;
      #0.2 CLKA_active = 1'b0;
   end
   else
      CLKA_active <= 1'b0;
end
always @(posedge CLKB) begin
   if (CEB) begin
      CLKB_active <= 1'b1;
      #0.2 CLKB_active = 1'b0;
   end
   else
      CLKB_active <= 1'b0;
end

////////////////////////////////////////////////////////////////////////////////////////////
//
////////////////////////////////////////////////////////////////////////////////////////////
//assign cas_inta = cas_en[0] ? (cas_en[1] ? ~ada_reg[13] : ada_reg[13]) : 1'b1;
//assign cas_intb = cas_en[0] ? (cas_en[1] ? ~adb_reg[13] : adb_reg[13]) : 1'b1;
assign cas_inta = cas_en[1] ? ~ada_reg[13] : ada_reg[13];
assign cas_intb = cas_en[1] ? ~adb_reg[13] : adb_reg[13];

always @(*) begin
    if(WRITE_MODE_A == "NORMAL_WRITE" && wea_reg == 1'b1) begin
        cas_sela = cas_sela;
    end else begin
        cas_sela = cas_inta;
    end
end
always @(*) begin
    if(WRITE_MODE_B == "NORMAL_WRITE" && web_reg == 1'b1) begin
        cas_selb = cas_selb;
    end else begin
        cas_selb = cas_intb;
    end
end

assign a_out_mux[0] = ((cas_sela == 1'b0) && cas_en == 2'b11) ? CINA : a_out[0];
assign a_out_mux[8:1] = a_out[8:1];
assign b_out_mux[0] = ((cas_selb == 1'b0) && cas_en == 2'b11) ? CINB : b_out[0];
assign b_out_mux[8:1] = b_out[8:1];

assign COUTA = a_out_mux[0];
assign COUTB = b_out_mux[0];

generate
////////////////////////////////////////////////////////////////////////////////////////////
// ROM or SINGLE_PORT 
////////////////////////////////////////////////////////////////////////////////////////////
if(RAM_MODE == "ROM" || RAM_MODE == "SINGLE_PORT") begin:ROMorSP_MODE

    always @(posedge CLKA) begin
        if (CEA)
            db_reg[8:0] <= DIB[8:0];
    end
    if (DATA_WIDTH_A >= 16 || DATA_WIDTH_B >= 16) begin

        assign write_en_a = csa_reg && cas_inta && (wea_reg == 1'b1);
        assign read_en_b  = csb_reg && cas_intb && (web_reg == 1'b0);
        // Port A operations
        always @(negedge CLKA_active)
        begin
            if (write_en_a) begin  // write
                mem_write_a(ada_reg[12:0], {db_reg[8:0], da_reg[8:0]}, bea_reg[1:0]);
            end
        end
        // Port B operations
        always @(negedge CLKB_active or posedge rstb_int)
        begin
            if (rstb_int)
               {b_out[width_b-1:0], a_out[width_b-1:0]} = {RSTB_VAL[width_b-1:0],RSTA_VAL[width_b-1:0]};
            else if(read_en_b)
               {b_out[width_b-1:0], a_out[width_b-1:0]} = mem_read_b(adb_reg[12:0]);
        end

    end
    else  begin   //x1 x2 x4 x8 x9

        assign write_en_a = csa_reg && cas_inta && (wea_reg == 1'b1);
        assign read_en_a  = csa_reg && cas_inta && (wea_reg == 1'b0);
        // Port A operations
        always @(negedge CLKA_active)
        begin
            if (write_en_a)  begin  // write
               // read during write
               if (WRITE_MODE_A == "TRANSPARENT_WRITE") begin
                   a_out[width_a-1:0] = da_reg[width_a-1:0];
               end
               else if (WRITE_MODE_A == "READ_BEFORE_WRITE")
                   a_out[width_a-1:0] = mem_read_a(ada_reg[12:0]);

               mem_write_a(ada_reg[12:0], da_reg[8:0], 2'b0);
            end
        end

        always @(negedge CLKA_active or posedge rsta_int)
        begin
            if (rsta_int)
               a_out[width_a-1:0] = RSTA_VAL[width_a-1 : 0];
            else if (read_en_a)          // read 
               a_out[width_a-1:0] = mem_read_a(ada_reg[12:0]);
        end
    end
end
////////////////////////////////////////////////////////////////////////////////////////////
//SIMPLE_DUAL_PORT
////////////////////////////////////////////////////////////////////////////////////////////
else if(RAM_MODE == "SIMPLE_DUAL_PORT")begin:SDP_MODE
    //port_A operation: only write in SDP MODE
    if (DATA_WIDTH_A >= 16) begin:PORTA

        assign write_en_a = csa_reg && cas_inta && (wea_reg == 1'b1);

        always @(posedge CLKA) begin
           if (CEA)
              db_reg[8:0]  <= DIB[8:0];
        end
        always @(negedge CLKA_active) begin
           if (write_en_a)    // write 
              mem_write_a(ada_reg[12:0], {db_reg[8:0], da_reg[8:0]},bea_reg[1:0]);
        end
    end
    else  begin:PORTA    //  x1 x2 x4 x8 x9

        assign write_en_a = csa_reg && cas_inta && (wea_reg == 1'b1);
        assign read_en_a  = csa_reg && cas_inta && (wea_reg == 1'b0) ;

        always @(negedge CLKA_active) begin
           if (write_en_a)     // write
           begin
              if (WRITE_MODE_A == "TRANSPARENT_WRITE")
              begin
                 a_out[width_a-1:0] = da_reg[width_a-1:0];
              end
              else if (WRITE_MODE_A == "READ_BEFORE_WRITE")
                 a_out[width_a-1 : 0] = mem_read_a(ada_reg[12:0]);

              mem_write_a(ada_reg[12:0], da_reg[8:0], 2'b0);
           end
        end
        if(DATA_WIDTH_B <16) begin
           always @(negedge CLKA_active or posedge rsta_int)
           begin
               if (rsta_int)
                  a_out[width_a-1 : 0] = RSTA_VAL[width_a-1:0];
               else if (read_en_a)
                  a_out[width_a-1 : 0] = mem_read_a(ada_reg[12:0]);
           end
        end
    end
    //port_B operation:only read in SDP MODE
    if (DATA_WIDTH_B >= 16) begin:PORTB
    // SIMPLE_DUAL_PORT 
        assign read_en_b  = csb_reg && cas_intb && (web_reg == 1'b0);

        always @(negedge CLKB_active or posedge rstb_int)
        begin
           if (rstb_int)
              {b_out[width_b-1 : 0], a_out[width_b-1 : 0]} = {RSTB_VAL[width_b-1:0],RSTA_VAL[width_b-1:0]};
           else if (read_en_b)       // read 
              {b_out[width_b-1 : 0], a_out[width_b-1 : 0]} = mem_read_b(adb_reg[12:0]);
        end
    end
    else  begin:PORTB  //  x1 x2 x4 x8 x9

        assign read_en_b  = csb_reg && cas_intb && (web_reg == 1'b0);

        always @(negedge CLKB_active or posedge rstb_int)
        begin
           if (rstb_int)
              b_out[width_b-1 : 0] = RSTB_VAL[width_b-1:0];
           else if (read_en_b)   //  read 
              b_out[width_b-1 : 0] = mem_read_b(adb_reg[12:0]);
        end
    end
end
////////////////////////////////////////////////////////////////////////////////////////////
//DP_MODE
////////////////////////////////////////////////////////////////////////////////////////////
else   begin:DP_MODE   //  --x1 x2 x4 x8 x9 
    assign write_en_a = csa_reg && cas_inta && (wea_reg == 1'b1) ;
    assign read_en_a  = csa_reg && cas_inta && (wea_reg == 1'b0) ;
    assign write_en_b = csb_reg && cas_intb && (web_reg == 1'b1) ;
    assign read_en_b  = csb_reg && cas_intb && (web_reg == 1'b0) ;
    // Port A operations
    always @(negedge CLKA_active)
    begin
        if (write_en_a)  begin  // write
            // read during write
            if (WRITE_MODE_A == "TRANSPARENT_WRITE")
            begin
               a_out[width_a-1:0] = da_reg[width_a-1:0];
            end
            else if (WRITE_MODE_A == "READ_BEFORE_WRITE")
               a_out[width_a-1 : 0] = mem_read_a(ada_reg[12:0]);

            mem_write_a(ada_reg[12:0], da_reg[8:0], 2'b0);
        end
    end

    always @(negedge CLKA_active or posedge rsta_int)
    begin
        if (rsta_int)
           a_out[width_a-1 : 0] = RSTA_VAL[width_a-1:0];
        else if (read_en_a)
           a_out[width_a-1 : 0] = mem_read_a(ada_reg[12:0]);
    end
    // Port B operations
    always @(posedge CLKB) begin
         if (CEB)
            db_reg[8:0] <= DIB[8:0];
    end

    always @(negedge CLKB_active)
    begin
        if (write_en_b)  begin  // write
            // read during write
            if (WRITE_MODE_B == "TRANSPARENT_WRITE")
            begin
                b_out[width_b-1:0] = db_reg[width_b-1:0];
            end
            else if (WRITE_MODE_B == "READ_BEFORE_WRITE")
                b_out[width_b-1 : 0] = mem_read_b(adb_reg[12:0]);

            mem_write_b(adb_reg[12:0], db_reg[8:0]);
        end
    end

    always @(negedge CLKB_active or posedge rstb_int)
    begin
        if (rstb_int)
           b_out[width_b-1 : 0] = RSTB_VAL[width_b-1:0];
        else if (read_en_b)
           b_out[width_b-1 : 0] = mem_read_b(adb_reg[12:0]);
    end
end

endgenerate

//////////////
// core latch
//////////////
assign grsn =  (GRS_EN == "TRUE") ? GRS_INST.GRSNET : 1'b1;
assign grs =  ~grsn;
or (rsta_grs, grs, RSTA);
or (rstb_grs, grs, RSTB);

reg rsta_grsn_d;

    always @(posedge CLKA_for_or) begin
        if (RSTA) begin
            rsta_grsn_d   <= 1'b1;
        end
        else begin
            rsta_grsn_d   <= 1'b0;
        end
    end

reg rstb_grsn_d;
    
    always @(posedge CLKB_for_or) begin
        if (RSTB) begin
            rstb_grsn_d   <= 1'b1;
        end
        else begin
            rstb_grsn_d   <= 1'b0;
        end
    end

initial begin
    rsta_grsn_d = 1'b1;
    rstb_grsn_d = 1'b1;
end

assign rsta_grs_sync  = (RST_TYPE == "SYNC") ? rsta_grsn_d : 1'b0;
assign rstb_grs_sync  = (RST_TYPE == "SYNC") ? rstb_grsn_d : 1'b0;
assign rsta_grs_async = (RST_TYPE == "ASYNC") ? rsta_grs : grs;
assign rstb_grs_async = (RST_TYPE == "ASYNC") ? rstb_grs : grs;

assign rsta_int = rsta_grs_sync | rsta_grs_async;
assign rstb_int = rstb_grs_sync | rstb_grs_async;
/////////////////////////////////////////////////////////////////////
//port out
assign CLKA_for_or = (DOA_REG_CLKINV == 1) ? ~CLKA : CLKA;
assign CLKB_for_or = (DOB_REG_CLKINV == 1) ? ~CLKB : CLKB;

generate
if (DATA_WIDTH_B >= 16)
begin:FAKE_DP_OUT
    //port_A output
    always @(posedge CLKB_for_or or posedge rstb_int)
    begin
        if (rstb_int)
            a_out_reg <= RSTA_VAL;
        else if (ORCEB)
            a_out_reg <= a_out;
    end

    //doa combination logic
    always @(*)
    begin
        if (DOB_REG == 0)
        begin
            case(DATA_WIDTH_B)
                16: doa[8:0] = a_out_mux[8:0];
                18: doa[width_b-1:0] = a_out_mux[width_b-1:0];
            endcase
        end
        else
        begin
            case(DATA_WIDTH_B)
                16: doa[8:0] = a_out_reg[8:0];
                18: doa[width_b-1:0] = a_out_reg[width_b-1 : 0];
            endcase
        end
    end

    always @(posedge CLKB_for_or or posedge rstb_int)
    begin
        if (rstb_int)
            b_out_reg <= RSTB_VAL;
        else if (ORCEB)
            b_out_reg <= b_out;
    end

    //dob combination logic
    always @(*)
    begin
        if (DOB_REG == 0)
        begin
            case(DATA_WIDTH_B)
                16: dob[8:0] = b_out_mux[8:0];
                18: dob[width_b-1:0] = b_out_mux[width_b-1 : 0];
            endcase
        end
        else
        begin
            case(DATA_WIDTH_B)
                16: dob[8:0] = b_out_reg[8:0];
                18: dob[width_b-1:0] = b_out_reg[width_b-1 : 0];
            endcase
        end
    end
end
else
begin:TRUE_DP_OUT
    //port_A output

    always @(posedge CLKA_for_or or posedge rsta_int)
    begin
        if (rsta_int)
            a_out_reg <= RSTA_VAL;
        else if (ORCEA)
            a_out_reg <= a_out_mux;
    end

    //doa combination logic
    always @(*)
    begin
        if (DOA_REG == 0)
        begin
            case(DATA_WIDTH_A)   
               1: doa[8:0] = {{8{1'b0}},a_out_mux[width_a-1:0]};
               2: doa[8:0] = {{7{1'b0}},a_out_mux[width_a-1:0]};
               4: doa[8:0] = {{5{1'b0}},a_out_mux[width_a-1:0]};
               8: doa[8:0] = a_out_mux[8:0];
               9: doa[8:0] = a_out_mux[8:0];
            endcase
        end
        else
        begin
            doa = a_out_reg;
        end
    end
    ////port_B output

    always @(posedge CLKB_for_or or posedge rstb_int)
    begin
        if (rstb_int)
            b_out_reg <= RSTB_VAL;
        else if (ORCEB)
            b_out_reg <= b_out_mux;
    end

    //dob combination logic
    always @(*)
    begin
        if (DOB_REG == 0)
        begin
            case(DATA_WIDTH_B)  
               1: dob[8:0] = {{8{1'b0}},b_out_mux[width_b-1:0]};
               2: dob[8:0] = {{7{1'b0}},b_out_mux[width_b-1:0]};
               4: dob[8:0] = {{5{1'b0}},b_out_mux[width_b-1:0]};
               8: dob[8:0] = b_out_mux[8:0];
               9: dob[8:0] = b_out_mux[8:0];
            endcase
        end
        else
            dob = b_out_reg;
    end
end
endgenerate

assign DOA = doa;
assign DOB = dob;

// synthesis translate_on
endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_OUTBUFDS.v
//
// Functional description: Differential Signaling Output Buffer
//
// Parameter description:
//      
//
// Port description:
//
// Revision:
//    06/18/14 - Initial version.
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_OUTBUFDS #(
    parameter IOSTANDARD = "DEFAULT"
)(
    output O,
    output OB,
    input I
) /* synthesis syn_black_box */ ;
  
  initial begin
    case (IOSTANDARD)
    "LVDS", "MINI-LVDS", "SUB-LVDS","TMDS", "DEFAULT" :;
    default : begin
           $display("Attribute Syntax Error : The attribute IOSTANDARD on GTP_OUTBUFDS instance %m is set to %s.", IOSTANDARD);
           $finish;
              end
    endcase
    end

    buf (O, I);
    not (OB, I);

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2015 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_FIFO18K.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//      2018/01/09: Update display informations.
//      2018/06/28: timescale defined
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps
 
module  GTP_FIFO18K
#(
    parameter GRS_EN = "TRUE",
    parameter integer DATA_WIDTH = 18,
    parameter integer DO_REG = 0,
    parameter [13:0] ALMOST_FULL_OFFSET = 14'h0000,
    parameter [13:0] ALMOST_EMPTY_OFFSET = 14'h0000,
    parameter integer USE_EMPTY = 0,
    parameter integer USE_FULL = 0,
    parameter REWRITE_EN = "FALSE",
    parameter RESEND_EN = "FALSE",
    parameter SYNC_FIFO = "FALSE"
) (
    output ALMOST_EMPTY,
    output ALMOST_FULL,
    output EMPTY,
    output FULL,
    output [35:0] DO,
    input [35:0] DI,
    input WCLK,
    input RCLK,
    input WCE,
    input RCE,
    input WERR,
    input WEOP,
    input RNAK,
    input ORCE,
    input RST
);

        reg  [14:0]             wptr_next;
        reg  [14:0]             rptr_next;
        reg  [14:0]             rd_binary;
        reg  [14:0]             wr_binary;
        reg  [13:0]             wcnt;
        reg  [13:0]             rcnt;
        reg  [14:0]             wr_binary_next;
        reg  [14:0]             rd_binary_next;
        reg                     empty_reg;
        reg                     full_reg;
        reg                     full_val;
        reg                     almost_full_reg;
        reg                     almost_empty_reg;
        reg  [14:0]             wr_addr_sop;
        reg  [14:0]             rd_addr_sop;
        reg                     resend_en;
        reg                     rewrite_en;
        reg                     flagempty_en;
        reg                     flagfull_en;
        reg                     dout_reg_en;
        reg                     sync_fifo;
        reg                     grs_en;
        reg                     rd_eop;  
        reg [35:0]              dout_reg;

      

        wire                    resend;
        wire                    rewrite;
        wire [14:0]             wptr_rclk;
        wire [14:0]             rptr_wclk;
        wire                    wclk,rclk;
        wire                    wr_en,rd_en;
        wire                    rstw,rstr;
        wire                    wr_err,wr_eop;
        wire                    rd_nak;
        wire                    full,empty;
        wire                    almost_empty,almost_full;
        wire  [13:0]            waddr,raddr;         
        wire  [35:0]            dout;
        wire                    dout_reg_in;
        wire  [35:0]            din;
        wire                    global_rstn;




initial   
  begin

        case(SYNC_FIFO)
                    "FALSE" : sync_fifo = 0;
                    "TRUE"  : sync_fifo = 1;
                    default : begin
                        $display ("ERROR: GTP_FIFO18K instance %m parameter SYNC_FIFO:%s, The legal values are FALSE or TRUE.",SYNC_FIFO);
                        $finish;
                    end
        endcase

        case(REWRITE_EN)
                    "FALSE" : rewrite_en = 0;
                    "TRUE"  : rewrite_en = 1;
                    default : begin
                        $display ("ERROR: GTP_FIFO18K instance %m parameter REWRITE_EN:%s, The legal values are FALSE or TRUE.",REWRITE_EN);
                        $finish;
                    end
        endcase

        case(RESEND_EN)
                    "FALSE" : resend_en = 0;
                    "TRUE"  : resend_en = 1;
                    default : begin
                        $display ("ERROR: GTP_FIFO18K instance %m parameter RESEND_EN:%s, The legal values are FALSE or TRUE.",RESEND_EN);
                        $finish;
                    end
        endcase

        case(USE_EMPTY)
                    1'b0 : flagempty_en = 0;
                    1'b1 : flagempty_en = 1;
                    default : begin
                        $display ("ERROR: GTP_FIFO18K instance %m parameter USE_EMPTY:%d, The legal values are 0 or 1.",USE_EMPTY);
                        $finish;
                    end
        endcase

        case(USE_FULL)
                    1'b0 : flagfull_en = 0;
                    1'b1 : flagfull_en = 1;
                    default : begin
                        $display ("ERROR: GTP_FIFO18K instance %m parameter USE_FULL:%d, The legal values are 0 or 1.",USE_FULL);
                        $finish;
                    end
        endcase

        case(DO_REG)
                    1'b0 : dout_reg_en = 0;
                    1'b1 : dout_reg_en = 1;
                    default : begin
                        $display ("ERROR: GTP_FIFO18K instance %m parameter DO_REG:%d, The legal values are 0 or 1.",DO_REG);
                        $finish;
                    end
        endcase


        case(GRS_EN)
                    "FALSE" : grs_en = 0;
                    "TRUE"  : grs_en = 1;
                    default : begin
                        $display ("ERROR: GTP_FIFO18K instance %m parameter GRS_EN:%s, The legal values are FALSE or TRUE.",GRS_EN);
                        $finish;
                    end
        endcase

        case(DATA_WIDTH)
                    1,2,4,8,9,16,18,32,36: ;
                    default : begin
                        $display ("ERROR: GTP_FIFO18K instance %m parameter DATA_WIDTH:%d, The legal values are 1,2,4,8,9,16,18,32 or 36.",DATA_WIDTH);
                        $finish;
                    end
        endcase

      dout_reg ='b0;
  end

assign dout_reg_in = ORCE;
assign din = DI;
assign wclk = WCLK;
assign rclk = RCLK;
assign wr_en = WCE;
assign rd_en = RCE;
assign rstw = !RST & global_rstn;
assign rstr = !RST & global_rstn;
assign wr_err = WERR;
assign wr_eop = WEOP;
assign rd_nak = RNAK;
assign EMPTY = empty;
assign FULL  = full;
assign ALMOST_EMPTY = almost_empty;
assign ALMOST_FULL = almost_full;


always @(posedge rclk or negedge rstr )
  begin
    if(!rstr)
      dout_reg <= 'b0;
      
    else if(dout_reg_in)
      dout_reg <= dout;
    else
     dout_reg <= dout_reg;
end    

assign DO = dout_reg_en ? dout_reg : dout;

always @(DATA_WIDTH or DO)
   begin 
     case(DATA_WIDTH)
    'd9  :   rd_eop = DO[8];
    'd18 :   rd_eop = DO[8];
    'd36 :   rd_eop = DO[26];
   default:
    rd_eop = 0;
endcase
end


assign global_rstn = grs_en ? GRS_INST.GRSNET : 1'b1;


//*************************************************************************************
//main code
//************************************************************************************* 
always @ (posedge wclk or negedge rstw )      //wr binary addr
  begin 
    if (rstw == 1'b0)
         wr_binary <= 15'd0;
    else
         wr_binary <= wr_binary_next;
  end

always @ (*) 
  begin
    if (rewrite == 1'b1)
         wr_binary_next = wr_addr_sop;
    else if (full == 1'b0)
         wr_binary_next = wr_binary + wr_en;
    else
         wr_binary_next = wr_binary;
  end

always @ (*)
  begin
    if (rewrite_en == 1'b1)
        wptr_next = wr_addr_sop;
    else
        wptr_next = wr_binary_next;
  end
//**************************************************************
reg wr_eop_d;
always @(posedge wclk or negedge rstw)
  begin
   if (rstw == 1'b0)
      wr_eop_d <= 1'b0;
   else
      wr_eop_d <= wr_eop;  //it's user's reponsibility to have wr_en == 1'b1 when wr_eop  == 1'b1
  end

reg wr_err_d;

assign wr_eop_in = rewrite_en && wr_eop_d && (~ wr_err_d);

always @ (posedge wclk or negedge rstw) 
  begin
    if (rstw == 1'b0)
        wr_err_d <= 1'b0;
    else
        wr_err_d <= wr_err; //it's user's reponsibility to have wr_en == 1'b1 when wr_en  == 1'b1
  end

assign rewrite = rewrite_en & wr_err_d;

always @ (posedge wclk or negedge rstw)
  begin
    if (rstw == 1'b0)
        wr_addr_sop <= 'd0;
    else if (wr_eop_in)  //it's user's responsibility to have wr_en == 1'b1 && wr_err == 1'b0 when wr_eop_in == 1'b1  
        wr_addr_sop <= wr_binary;
  end

localparam ASIZE = ((DATA_WIDTH == 32) || (DATA_WIDTH == 36)) ? 'd8 :
                   ((DATA_WIDTH == 16) || (DATA_WIDTH == 18)) ? 'd9 :
                   ((DATA_WIDTH == 8) || (DATA_WIDTH == 9)) ? 'd10 :
                   (DATA_WIDTH == 4) ? 'd11 :
                   (DATA_WIDTH == 2) ? 'd12 : 
                   (DATA_WIDTH == 1) ? 'd13 : 'bx;


//initial  
//  begin
//    case (ASIZE)
//     'd8 : 
//     if(DATA_WIDTH != 32 && DATA_WIDTH != 36)  begin
//         $display ("The ASIZE is mismatched with DATA_WIDTH,The legal input is  32 or 36");
//  end
//     'd9 :
//      if(DATA_WIDTH != 18 && DATA_WIDTH != 16 )  begin
//         $display ("The ASIZE is mismatched with DATA_WIDTH,The legal input is  18 or 16");
//  end
//     'd10 :
//      if(DATA_WIDTH != 9 && DATA_WIDTH != 8) begin
//         $display ("The ASIZE is mismatched with DATA_WIDTH,The legal input is 8 or 9");
//  end
//     'd11 : 
//      if(DATA_WIDTH != 4)   begin 
//         $display ("The ASIZE is mismatched with DATA_WIDTH,The legal input is 4");
//  end
//
//     'd12 :
//      if(DATA_WIDTH != 2)   begin
//         $display ("The ASIZE is mismatched with DATA_WIDTH,The legal input is 2");
//  end
// 
//     'd13 : 
//      if(DATA_WIDTH != 1)  begin
//         $display ("The ASIZE is mismatched with DATA_WIDTH,The legal input is 1");
//  end
//
//    default :
//         $display("the input DATA_WIDTH illegal.");
//      endcase
//  end


     
//***********************************************************************************************
always @ (*) begin
    case(ASIZE)
    'd13: begin
        full_val = (wr_binary_next[14:0] == {~rptr_wclk[14],rptr_wclk[13:0]});
    end
    'd12: begin
        full_val = (wr_binary_next[13:0] == {~rptr_wclk[13],rptr_wclk[12:0]});
    end
    'd11: begin
        full_val = (wr_binary_next[12:0] == {~rptr_wclk[12],rptr_wclk[11:0]});
    end
    'd10: begin
        full_val = (wr_binary_next[11:0] == {~rptr_wclk[11],rptr_wclk[10:0]});
    end
    'd9: begin
        full_val = (wr_binary_next[10:0] == {~rptr_wclk[10],rptr_wclk[9:0]});
    end
    default: begin
        full_val = (wr_binary_next[9:0] == {~rptr_wclk[9],rptr_wclk[8:0]});
    end
    endcase
end

always @ (posedge wclk or negedge rstw) begin     //write full flag
    if (rstw == 1'b0)
         full_reg <= 1'b0;
    else
         full_reg <= full_val; 
end

assign full=~flagfull_en |full_reg;
wire [14:0]  write_water_level = wr_binary_next- rptr_wclk;
wire [14:0]  write_water_level_gud = wr_binary- rptr_wclk;
always @ (posedge wclk or negedge rstw) begin     //write almost_full flag
    if (rstw == 1'b0)
         almost_full_reg <= 1'b0;
    else
         almost_full_reg <= write_water_level >= ALMOST_FULL_OFFSET;
  end

assign almost_full=~flagfull_en |almost_full_reg;
//****************************************************************************************************************************************
INT_FIFO18K_SYNCLOGIC #(
.c_DW (15)
) w2r_sync_logic (
//configuration
.sync_fifo       (sync_fifo),
.gray_en         (~rewrite_en),

.src_clk         (wclk),
.rstn_src        (rstw),
.src_data        (wptr_next), //binary
.des_clk         (rclk),
.rstn_des        (rstr),
.des_data        (wptr_rclk)//binary
);
//****************************************************************************************************************************************
INT_FIFO18K_SYNCLOGIC #(
.c_DW (15)
)r2w_sync_logic(
//configuration
.sync_fifo       (sync_fifo),
.gray_en         (~resend_en),
//
.src_clk         (rclk),
.rstn_src        (rstr),
.src_data        (rptr_next), //binary
.des_clk         (wclk),
.rstn_des        (rstw),
.des_data        (rptr_wclk)//binary
);
//****************************************************************************************************************************************
    INT_FIFO18K_MEM #(
        DATA_WIDTH , ASIZE
    ) fifomem1 (
        .dout(dout), .din(din),
        .waddr(waddr), .raddr(raddr),
        .wr_en(wr_en), .wclk(wclk), 
        .full(full),   .rstr(rstr),
        .rd_en(rd_en),  .rclk(rclk));

//*************************************************************************************************************************
wire [14:0] read_water_level; 
wire [14:0] read_water_level_gud; 

always @ (posedge rclk or negedge rstr) begin
    if(rstr == 1'b0)
    
         rd_binary <= 15'd0;
        
     
    else 
         rd_binary <= rd_binary_next;
end

wire [14:0] rd_binary_inc = rd_binary + 1;

always @ (*) begin
      if (resend)
         rd_binary_next = rd_addr_sop;
      else if ((~empty) & rd_en)
         rd_binary_next = rd_binary_inc;
      else
         rd_binary_next = rd_binary;
end
       

always @ (*) begin
    if (resend_en == 1'b1) 
        rptr_next = rd_addr_sop;
    else
        rptr_next = rd_binary_next;
end 
       
always @ (posedge rclk or negedge rstr) begin
      if (rstr == 1'b0) begin
          empty_reg <= 1'b1;
      end
      else begin
          empty_reg <= wptr_rclk == rd_binary_next;
      end
end

assign empty=~flagempty_en |empty_reg;
assign read_water_level = wptr_rclk - rd_binary_next; 
assign read_water_level_gud = wptr_rclk - rd_binary;
 
always @ (posedge rclk or negedge rstr) begin
      if (rstr == 1'b0) begin
          almost_empty_reg <= 1'b1;
      end
      else begin
          almost_empty_reg <= read_water_level <= ALMOST_EMPTY_OFFSET;
      end
end

assign almost_empty=~flagempty_en |almost_empty_reg;
//*****************************************************************************                   
always @ (*) begin
case(ASIZE) 
     'd13: wcnt <= wr_binary[13:0];
     'd12: wcnt <= {wr_binary[12:0],1'b1};
     'd11: wcnt <= {wr_binary[11:0],2'b11};
     'd10: wcnt <= {wr_binary[10:0],3'b111};
     'd9:  wcnt <= {wr_binary[9:0],4'b1111}; 
     'd8:  wcnt <= {wr_binary[8:0],5'b11111};
     default: 
      $display("ERROR: GTP_FIFO18K instance %m local parameter ASIZE:%d is illegal. The legal value is 8,9,19,11,12 or 13",ASIZE);

endcase
end

                   
always @ (*) begin
case(ASIZE) 
     4'd13: rcnt <=  rd_binary[13:0];
     4'd12: rcnt <= {rd_binary[12:0],1'b1};
     4'd11: rcnt <= {rd_binary[11:0],2'b11};
     4'd10: rcnt <= {rd_binary[10:0],3'b111};
     4'd9:  rcnt <= {rd_binary[9:0],4'b1111};
     4'd8:  rcnt <= {rd_binary[8:0],5'b11111};
     default:
      $display("ERROR: GTP_FIFO18K instance %m local parameter ASIZE:%d is illegal. The legal value is 8,9,19,11,12 or 13",ASIZE);

endcase
end

assign #0 waddr = wcnt;
assign #0 raddr = rcnt;
//****************************************************************

reg rd_nak_d; 
always @ (posedge rclk or negedge rstr) begin
    if (rstr == 1'b0) 
         rd_nak_d <= 1'b0;
    else
         rd_nak_d <= rd_nak; //it is user's responsibility to have rd_en == 1'b1 when rd_nak == 1'b1
end

assign resend = resend_en & rd_nak_d;

reg [1:0] rd_en_d;
always @ (posedge rclk or negedge rstr) begin
   if (!rstr) begin
      rd_en_d <= 2'd0;
   end
   else begin
      if (resend)
         rd_en_d <= 2'd0;
      else if (rd_en)
         rd_en_d <= {rd_en_d[0], (~empty)};
   end
end

assign rd_valid = dout_reg_en ? rd_en_d[1] : rd_en_d[0];


always @ (posedge rclk or negedge rstr) begin
    if (rstr == 1'b0) 
        rd_addr_sop <= 'd0;
    else if (rd_eop & rd_valid & (~resend)) begin
        if (dout_reg_en) begin
           if (~rd_en_d[0])
              rd_addr_sop <= rd_binary;
           else
              rd_addr_sop <= rd_binary - 1;
        end  
        else
           rd_addr_sop <= rd_binary; 
    end
    else 
        rd_addr_sop <= rd_addr_sop;
end 
        
         
endmodule

module INT_FIFO18K_SYNCLOGIC #(
    parameter ASIZE = 12,// 8 9 10 11 12 13 
    parameter c_DW =  15 
)(
//configuration
    input sync_fifo,
    input gray_en,

    input src_clk,
    input rstn_src,
    input [c_DW-1:0] src_data, //binary
    input des_clk,
    input rstn_des,
    output reg [c_DW-1:0] des_data //binary
);

        wire [c_DW-1:0] src_data_gray;
        reg [1:0] update_ack_dly;
        reg [c_DW-1:0] data_buf;
        reg update_ack;
        reg update_strobe;

assign src_data_gray = (src_data>>1)^src_data;
//source clk domain
always @(posedge src_clk or negedge rstn_src)
   if (!rstn_src) begin
      update_ack_dly <= 0;
      update_strobe  <= 0;
      data_buf       <= 0;
   end
   else begin
      update_ack_dly <= {update_ack_dly[0], update_ack};

      //latch new data
      if (update_strobe == update_ack_dly[1]) begin
         data_buf <= src_data_gray;  //need to convert into gray code
         if (gray_en)
            update_strobe <= 1'b0;
         else
            update_strobe <= ~ update_strobe;
      end
   end

//**********************************************************************
        reg [c_DW-1:0] data_buf_d1;
        reg [c_DW-1:0] data_buf_d2;
        reg  [1:0] update_strobe_dly;

always @(posedge des_clk or negedge rstn_des)
   if (!rstn_des) begin
      data_buf_d1 <= 0;
      data_buf_d2 <= 0;
      update_strobe_dly <= 0;
      update_ack <= 1'b0;
   end
   else begin
      update_strobe_dly <= {update_strobe_dly[0], update_strobe};
      data_buf_d1 <= data_buf;
      if (sync_fifo)
         data_buf_d2 <= src_data_gray;
      else if (gray_en)
         data_buf_d2 <= data_buf_d1;
      else if (update_strobe_dly[1] !=  update_ack) begin
         data_buf_d2 <= data_buf_d1;
         update_ack <= ~ update_ack;
      end
   end

integer i;

always @(*) begin
   for (i=0; i< c_DW;i=i+1)
       des_data[i] = ^(data_buf_d2>>i);
end

endmodule


//*********************************THE MEM MODULE*****************************
module INT_FIFO18K_MEM (dout, din, waddr, raddr, wr_en, wclk,full,rstr,rd_en,rclk);

        parameter DATA_WIDTH = 2; // Memory data word width
        parameter ASIZE = 12; // Number of memory address bits

        output [35:0] dout;
        input rstr;
        input rd_en;
        input [35:0] din;
        input [13:0] waddr, raddr;
        input wr_en, wclk,rclk;
        input full;

        reg [(DATA_WIDTH-1):0] MEM [0:(1<<14)-1];  
        integer k;      
        reg [35:0] dout;  
initial
   begin                   
      for(k=0;k<(1<<14);k=k+1)   
         MEM[k]<={DATA_WIDTH{1'b0}};
     dout <='b0;
     end
    

//assign dout = rd_en ? MEM[raddr]:dout;
always @(posedge rclk or negedge rstr)
    begin
      if(!rstr)
       dout <= 'b0;
      else if(rd_en )
    dout <= MEM[raddr];
  else
    dout <= dout;
end
always @(posedge wclk )
    begin 
    if (wr_en && !full) MEM[waddr] <= din;
end
endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_RAM32X1SP.v
//
// Functional description: single-port 32x1 distributed ram
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_RAM32X1SP
#(
    parameter [31:0] INIT = 32'h00000000
) (
    output  DO,
    input   DI,
    input [4:0] ADDR,
    input WCLK, WE
);

    reg [31:0] mem ;

    initial begin
        mem = INIT;
    end

    always @(posedge WCLK) begin
        if (WE == 1'b1) begin
            mem[ADDR] <= DI;
        end
    end

    assign DO = mem[ADDR];

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_DFF_RE.v
//
// Functional description: D-type flip-flop with sync clear and enable
//
// Parameter description:
//      INIT: init value
//
// Port description:
//      R: synchronous clear
//      CE  : enable
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_DFF_RE
#(
    parameter GRS_EN = "TRUE",
    parameter INIT = 1'b0
) (
    output reg Q,
    input wire D,
    input wire CLK, R, CE
);

    wire grs_n;
    wire RS;

    tri1 grsnet = GRS_INST.GRSNET;
    assign grs_n=(GRS_EN=="TRUE")?grsnet:1'b1;

    not (RS, grs_n);

    initial Q = 1'bx;

    always @(posedge CLK or posedge RS) begin
        if (RS)
            Q <= 1'b0;
        else if (R)
            Q <= 1'b0;
        else if (CE)
            Q <= D;
    end

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_EFUSECODE.v
//
// Functional description: efuse for user
//
// Parameter description:
//      
//
// Port description:
//      
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps 

module GTP_EFUSECODE
#(
    parameter [31:0] SIM_EFUSE_VALUE = 32'h12345678
)
(
    output [31:0] EFUSE_CODE// EFUSECODE signals
);

assign EFUSE_CODE = SIM_EFUSE_VALUE;

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_ISERDES.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//   2016/10/18: Remove ISERDES_MODE parameter value "NONE"
//   2018/08/17: change IGDES4/7/8 to IDES4/7/8
//               change IGDDR to IDDR
//               by xxma
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_ISERDES #(
parameter ISERDES_MODE = "IDDR",   //"IDDR","IMDDR","IDES4","IMDES4","IDES7","IDES8","IMDES8"
parameter GRS_EN = "TRUE",          //"TRUE"; "FALSE"
parameter LRS_EN = "TRUE"           //"TRUE"; "FALSE"
)(
input        DI,
input        ICLK,
input        DESCLK,
input        RCLK,
input  [2:0] WADDR,
input  [2:0] RADDR,
input        RST,
output [7:0] DO
)/* synthesis syn_black_box */;

//synthesis translate_off

reg        DI_P_reg;
reg        DI_N_reg;
reg  [7:0] DI_P_mem;
reg  [7:0] DI_N_mem;
reg  [7:0] DO_reg;
reg  [7:0] shift_reg;
reg  [7:0] capture_reg;
wire       capture_en0;
wire       capture_en1;
wire       cnt_rst;
reg  [2:0] cnt;
reg        rstn_dly;
reg  [7:0] out_en;
reg        imem_mode;
reg  [3:0] idata_width;

wire [7:0] DO_int;
wire       RCLK_buf;
wire       ICLK_buf;
wire       DESCLK_buf;
wire       DI_buf;
wire [2:0] WADDR_buf;
wire [2:0] RADDR_buf;

initial begin
    if(GRS_EN != "TRUE" && GRS_EN != "FALSE")
    begin
      $display("GTP_ISERDES Error: Illegal setting of GRS_EN %s",GRS_EN);
      $finish;
    end
    if(LRS_EN != "TRUE" && LRS_EN != "FALSE")
    begin
      $display("GTP_ISERDES Error: Illegal setting of LRS_EN %s",LRS_EN);
      $finish;
    end
    case(ISERDES_MODE)
        "IDDR":   begin
                     imem_mode = 0;
                     idata_width = 2;
                     out_en = 8'b1100_0000;
                   end
        "IMDDR":   begin
                     imem_mode = 1;
                     idata_width = 2;
                     out_en = 8'b1100_0000;
                   end
        "IDES4":  begin
                     imem_mode = 0;
                     idata_width = 4;
                     out_en = 8'b1111_0000;
                   end
        "IMDES4":  begin
                     imem_mode = 1;
                     idata_width = 4;
                     out_en = 8'b1111_0000;
                   end
        "IDES7":  begin
                     imem_mode = 0;
                     idata_width = 7;
                     out_en = 8'b1111_1110;
                   end
        "IDES8":  begin
                     imem_mode = 0;
                     idata_width = 8;
                     out_en = 8'b1111_1111;
                   end
        "IMDES8":  begin
                     imem_mode = 1;
                     idata_width = 8;
                     out_en = 8'b1111_1111;
                   end
        default:   begin
                     $display("GTP_ISERDES Error: Illegal setting of ISERDES_MODE %s",ISERDES_MODE);
                     $finish;
                   end
    endcase
end
///////////////////////////////////////////////////////////////////////////
assign DI_buf = DI;
assign WADDR_buf = WADDR;
assign RADDR_buf = RADDR;
assign ICLK_buf =  (imem_mode) ? ICLK : ((idata_width == 2) ? RCLK : DESCLK);
assign DESCLK_buf = (idata_width == 2) ? RCLK : DESCLK;
assign RCLK_buf = RCLK;
assign DO = DO_int;
///////////////////////////////////////////////////////////////////////////
assign global_rstn = (GRS_EN == "TRUE") ? GRS_INST.GRSNET : 1'b1;
assign lrs_rstn = (LRS_EN == "TRUE") ? (~RST) : 1'b1;
///////////////////////////////////////////////////////////////////////////
//for input dule data rate
always @(posedge ICLK_buf or negedge global_rstn or negedge lrs_rstn) 
begin
   if (!global_rstn)
      DI_P_reg <= 0;
   else if (!lrs_rstn)
      DI_P_reg <= 0;
   else
      DI_P_reg <= DI_buf;
end
always @(negedge ICLK_buf or negedge global_rstn or negedge lrs_rstn) 
begin
   if (!global_rstn)
      DI_N_reg <= 0;
   else if (!lrs_rstn)
      DI_N_reg <= 0;
   else
      DI_N_reg <= DI_buf;
end
///////////////////////////////////////////////////////////////////////////
//for input dule data rate in mem mode
always @(negedge ICLK_buf or negedge global_rstn or negedge lrs_rstn)
begin
   if (!global_rstn)
      DI_P_mem <= 0;
   else if (!lrs_rstn)
      DI_P_mem <= 0;
   else
      DI_P_mem[WADDR_buf] <= DI_P_reg;
end
always @(negedge ICLK_buf or negedge global_rstn or negedge lrs_rstn)
begin
   if (!global_rstn)
      DI_N_mem <= 0;
   else if (!lrs_rstn)
      DI_N_mem <= 0;
   else
      DI_N_mem[WADDR_buf] <= DI_buf; 
end
///////////////////////////////////////////////////////////////////////////
wire q_pos,q_neg;
assign q_pos=DI_P_mem[RADDR_buf];
assign q_neg=DI_N_mem[RADDR_buf];

always @(posedge DESCLK_buf or negedge global_rstn or negedge lrs_rstn)
begin
   if (!global_rstn)
      shift_reg <= 0;
   else if (!lrs_rstn)
      shift_reg <= 0;
   else
   begin
      if(imem_mode)
          shift_reg <= {DI_N_mem[RADDR_buf], DI_P_mem[RADDR_buf], shift_reg[7:2]};
      else
          shift_reg <= {DI_N_reg, DI_P_reg, shift_reg[7:2]};
   end
end
///////////////////////////////////////////////////////////////////////////
always @(posedge DESCLK_buf or negedge global_rstn or negedge lrs_rstn)
begin
   if (!global_rstn)
      rstn_dly <= 0;
   else if (!lrs_rstn)
      rstn_dly <= 0;
   else
      rstn_dly <= 1'b1;
end
///////////////////////////////////////////////////////////////////////////
always @(posedge DESCLK_buf or negedge global_rstn or negedge lrs_rstn)
begin
   if (!global_rstn)
      cnt <= 0;
   else if (!lrs_rstn || cnt_rst)
      cnt <= 0;
   else if (rstn_dly)
      cnt <= cnt + 1;
end

assign cnt_rst = (idata_width == 4) ? (cnt == 1) :
                 ((idata_width == 8) ? (cnt == 3) :
                 ((idata_width == 7) ? (cnt == 6) : 1'b0));
assign capture_en0 = (idata_width == 4) ? (cnt == 1) :
                    ((idata_width == 8) ? (cnt == 3) :
                    ((idata_width == 7) ? (cnt == 2) : 1'b0));
assign capture_en1 = cnt == 5;
///////////////////////////////////////////////////////////////////////////
always @(posedge DESCLK_buf or negedge global_rstn or negedge lrs_rstn)
begin
   if (!global_rstn)
      capture_reg <= 0;
   else if (!lrs_rstn)
      capture_reg <= 0;
   else if (capture_en0)
      capture_reg <= shift_reg;
   else if (capture_en1 && (idata_width == 7))
      capture_reg <= {DI_P_reg, shift_reg[7:1]};
end
///////////////////////////////////////////////////////////////////////////
always @(posedge RCLK_buf or negedge global_rstn or negedge lrs_rstn)
begin
   if (!global_rstn)
      DO_reg <= 0;
   else if (!lrs_rstn)
      DO_reg <= 0;
   else
      DO_reg <= capture_reg;      
end
assign DO_int = out_en & ((idata_width == 2) ? shift_reg : DO_reg);

//synthesis translate_on

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_DLL_E1.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//2018/01/03: initial version
//2018/03/12: fix error
//2018/04/02: change DELAY_STEP0 to DELAY_STEP for compatibility 
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps
module GTP_DLL_E1 #(
parameter GRS_EN = "TRUE", //TRUE, FALSE;
parameter FAST_LOCK = "TRUE", //FALSE, TRUE
parameter DELAY_STEP_OFFSET = 0  //-4, -3,-2, -1, 0, 1, 2, 3, 4
)(
output [7:0] DELAY_STEP,
output [7:0] DELAY_STEP1,
output LOCK,
input CLKIN,
input UPDATE_N,
input RST,
input PWD
)/* synthesis syn_black_box */;

//synthesis translate_off
reg        clk_osc;
reg [1:0]  pwd_clkosc;
reg [1:0]  pwd_clkin;
reg [10:0] cnt_div;
reg [1:0]  clkin_div_d;
reg [11:0] cnt;
reg [1:0]  state;
reg [1:0]  next_state;
reg [2:0]  stop;
reg [11:0] lth_code;
reg [1:0]  lock_update;
reg [7:0]  code_scaled_d;
reg [1:0]  updncnt_reg;
reg [7:0]  ctrl_code_reg;

reg clkin_update;
reg lth_en;
reg carry_en;
reg rstn_counter;
reg carry_q;
reg div_osc_lock;
reg lock_reg;

wire global_rstn;
wire lsr_rstn;
wire clk_osc_tmp;
wire clkin_tmp;
wire clkin_div;
wire counter_en;
wire carry_d;
wire [11:0] scaled_code_0;
wire [8:0]  scaled_code_1;
wire [7:0]  code_scaled;

initial
begin
    if ((GRS_EN == "TRUE")  || (GRS_EN == "FALSE")) begin
    end
    else
        $display (" GTP_DLL error: illegal setting for GRS_EN");

    if ((FAST_LOCK == "TRUE")  || (FAST_LOCK == "FALSE")) begin
    end
    else
        $display (" GTP_DLL error: illegal setting for FAST_LOCK");

    if ((DELAY_STEP_OFFSET == -4)  || (DELAY_STEP_OFFSET == -3) || (DELAY_STEP_OFFSET == -2)  || (DELAY_STEP_OFFSET == -1) ||(DELAY_STEP_OFFSET == 0)  || (DELAY_STEP_OFFSET == 1) ||(DELAY_STEP_OFFSET == 2)  || (DELAY_STEP_OFFSET == 3) ||(DELAY_STEP_OFFSET == 4)) begin
    end
    else
        $display (" GTP_DLL error: illegal setting for DELAY_STEP_OFFSET");
end

initial
begin
    clk_osc       = 1'b0;
    pwd_clkosc    = 2'b0;
    pwd_clkin     = 2'b0;
    cnt_div       = 11'b0;
    clkin_div_d   = 2'b0;
    cnt           = 12'b0;
    state         = 2'b0;
    next_state    = 2'b0;
    stop          = 3'b0;
    lth_code      = 12'b0;
    lock_update   = 2'b0;
    code_scaled_d = 8'b0;
    updncnt_reg   = 2'b0;
    ctrl_code_reg = 8'b0;
    clkin_update  = 1'b0;
    lth_en        = 1'b0;
    carry_en      = 1'b0;
    rstn_counter  = 1'b0;
    carry_q       = 1'b0;
    div_osc_lock  = 1'b0;
    lock_reg      = 1'b0;
end


assign global_rstn = (GRS_EN == "TRUE") ? GRS_INST.GRSNET : 1'b1;
assign lsr_rstn    = ~RST;

always #6.4 clk_osc = ~ clk_osc;

always @(negedge clk_osc or negedge global_rstn or negedge lsr_rstn)
begin
    if(!global_rstn)
        pwd_clkosc <= 2'b0;
    else if(!lsr_rstn)
        pwd_clkosc <= 2'b0;
    else
        pwd_clkosc <={pwd_clkosc[0],PWD};
end 
    
always @(negedge CLKIN or negedge global_rstn or negedge lsr_rstn)
begin
    if(!global_rstn)
        pwd_clkin <= 2'b0;
    else if(!lsr_rstn)
        pwd_clkin <= 2'b0;
    else
        pwd_clkin <= {pwd_clkin[0],PWD};
end

assign clk_osc_tmp = (~pwd_clkosc[1])&clk_osc;
    
assign clkin_tmp = (~pwd_clkin[1])&CLKIN;

always @(posedge clkin_tmp or negedge global_rstn or negedge lsr_rstn)
begin
    if (!global_rstn)
        cnt_div <= 0;
    else if (!lsr_rstn)
        cnt_div <= 0;
    else
        cnt_div <= cnt_div + 1;
end

assign clkin_div = cnt_div[10];

always @(posedge clk_osc_tmp or negedge global_rstn or negedge lsr_rstn)
begin
    if (!global_rstn)
        clkin_div_d <= 0;
    else if (!lsr_rstn)
        clkin_div_d <= 0;
    else
        clkin_div_d <= {clkin_div_d[0], clkin_div};
end

assign counter_en = clkin_div_d[1];

always @(posedge clk_osc_tmp or negedge global_rstn or negedge lsr_rstn)
begin
    if (!global_rstn)
        cnt <= 0;
    else if (!lsr_rstn)
        cnt <= 0;
    else if (!rstn_counter)
        cnt <= 0;
    else if (counter_en)
        cnt <= cnt + 1;
end

always @(posedge clk_osc_tmp or negedge global_rstn or negedge lsr_rstn)
begin
    if(!global_rstn)
        state <= 2'b00;
    else if(!lsr_rstn)
        state <= 2'b00;
    else
        state <= next_state;
end

always @(state or counter_en or stop)
begin
    case(state)
        2'b00: if(counter_en)
                next_state = 2'b01;
            else
                next_state = 2'b00;
        2'b01: if(counter_en == 1'b0)
                next_state = 2'b10;
            else
                next_state = 2'b01;
        2'b10: if(counter_en == 1'b0 && stop == 3'h7)
                next_state = 2'b11;
            else
                next_state = 2'b10;
        2'b11: begin
                next_state = 2'b00;
            end
    endcase
end

always @(posedge clk_osc_tmp or negedge global_rstn or negedge lsr_rstn)
begin
    if(!global_rstn)
        stop <= 3'b0;
    else if(!lsr_rstn)
        stop <= 3'b0;
    else if(state == 2'b10)
        stop <= stop + 1;
    else
        stop <= 3'b0;
end

always @(state or stop or div_osc_lock)
begin
    clkin_update   = 1'b0;
    lth_en         = 1'b0;
    carry_en       = 1'b0;
    rstn_counter   = 1'b1;
    case(state)
    2'b00: begin
           if(div_osc_lock)
               clkin_update = 1'b1;
           else
               clkin_update = 1'b0;
           end
    2'b01: ;
    2'b10: begin
               if(stop == 3'b000) begin
                   lth_en = 1'b1;
               end
               else if(stop == 3'b100) begin
                   carry_en = 1'b1;
                end
           end

    2'b11: rstn_counter = 1'b0;
    endcase
end

always @(posedge clk_osc_tmp or negedge global_rstn or negedge lsr_rstn)
begin
    if(!global_rstn)
        lth_code <= 12'b0;
    else if(!lsr_rstn)
        lth_code <= 12'b0;
    else if(lth_en)
        lth_code <= cnt;
end

assign scaled_code_0 = lth_code[10:0]*(8+DELAY_STEP_OFFSET)/8;

always @(posedge clk_osc_tmp or negedge global_rstn or negedge lsr_rstn)
begin
    if(!global_rstn)
        carry_q <= 1'b0;
    else if(!lsr_rstn)
        carry_q <= 1'b0;
    else if(carry_en)
        carry_q <= carry_d;
end

assign carry_d = carry_q ? scaled_code_0[2]|scaled_code_0[1] : scaled_code_0[2]&scaled_code_0[1];

assign scaled_code_1 = scaled_code_0[10:3] + carry_q;

assign over_flow = lth_code[11]|scaled_code_0[11]|scaled_code_1[8];

assign code_scaled = over_flow ? 8'hFF : scaled_code_1[7:0];

always @(posedge clk_osc_tmp or negedge global_rstn or negedge lsr_rstn)
begin
    if(!global_rstn)
        div_osc_lock <= 1'b0;
    else if(!lsr_rstn)
        div_osc_lock <= 1'b0;
    else if(state == 2'b11)
        div_osc_lock <= 1'b1;
end

always @(posedge CLKIN or negedge global_rstn or negedge lsr_rstn)
begin
    if (!global_rstn)
        lock_update <= 2'b0;
    else if(!lsr_rstn)
        lock_update <= 2'b0;
    else
        lock_update <= {lock_update[0],clkin_update};
end

always @(posedge CLKIN or negedge global_rstn or negedge lsr_rstn)
begin
    if (!global_rstn)
        code_scaled_d <= 8'd0;
    else if(!lsr_rstn)
        code_scaled_d <= 8'd0;
    else if (lock_update[1])
        code_scaled_d <= code_scaled;
end

always @(posedge CLKIN or negedge global_rstn or negedge lsr_rstn)
begin
    if (!global_rstn)
        lock_reg <= 1'b0;
    else if(!lsr_rstn)
        lock_reg <= 1'b0;
    else if(lock_update[1])
        lock_reg <= div_osc_lock;
end

always @(posedge CLKIN or negedge global_rstn or negedge lsr_rstn)
begin
    if(!global_rstn)
        updncnt_reg <= 2'b0;
    else if(!lsr_rstn)
        updncnt_reg <= 2'b0;
    else
       updncnt_reg <= {updncnt_reg[0], ~UPDATE_N};
end 

always@(posedge CLKIN or negedge global_rstn or negedge lsr_rstn)
begin
    if(!global_rstn)
        ctrl_code_reg <= 8'b0;
    else if(!lsr_rstn)
        ctrl_code_reg <= 8'b0;
    else if(updncnt_reg[1])
        ctrl_code_reg <= code_scaled_d;
end

assign DELAY_STEP = ctrl_code_reg;

assign DELAY_STEP1 = code_scaled_d;

assign LOCK = lock_reg;

//pragma translate_on 
endmodule







//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_LUT5.v
//
// Functional description: 5-input Look-Up-Table
//
// Parameter description:
//      INIT: init value
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_LUT5
#(
    parameter [31:0] INIT = 32'h0000_0000
) (
    output wire Z,
    input wire I0, I1, I2, I3, I4
);

    wire x7, x6, x5, x4, y1;
    wire x3, x2, x1, x0, y0;

    INT_LUTMUX4_UDP (x7, I1, I0, INIT[31], INIT[30], INIT[29], INIT[28]);
    INT_LUTMUX4_UDP (x6, I1, I0, INIT[27], INIT[26], INIT[25], INIT[24]);
    INT_LUTMUX4_UDP (x5, I1, I0, INIT[23], INIT[22], INIT[21], INIT[20]);
    INT_LUTMUX4_UDP (x4, I1, I0, INIT[19], INIT[18], INIT[17], INIT[16]);
    INT_LUTMUX4_UDP (y1, I3, I2, x7, x6, x5, x4);

    INT_LUTMUX4_UDP (x3, I1, I0, INIT[15], INIT[14], INIT[13], INIT[12]);
    INT_LUTMUX4_UDP (x2, I1, I0, INIT[11], INIT[10], INIT[9], INIT[8]);
    INT_LUTMUX4_UDP (x1, I1, I0, INIT[7], INIT[6], INIT[5], INIT[4]);
    INT_LUTMUX4_UDP (x0, I1, I0, INIT[3], INIT[2], INIT[1], INIT[0]);
    INT_LUTMUX4_UDP (y0, I3, I2, x3, x2, x1, x0);

    INT_LUTMUX2_UDP (Z, I4, y1, y0);

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: Internal simulation model
// Filename: GTP_OUTBUF.v
//
// Functional description: output buffer
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_OUTBUF #(
    parameter IOSTANDARD = "DEFAULT",
    parameter SLEW_RATE = "SLOW",
    parameter DRIVE_STRENGTH = "8"
)(
    output O,
    input I
) /* synthesis syn_black_box */ ;

  initial begin
    case (IOSTANDARD)
    "LVTTL33", "PCI33", "LVCMOS33", "LVCMOS25", "LVCMOS18", "LVCMOS15", "LVCMOS12", "SSTL25_I", "SSTL25_II", "SSTL18_I", "SSTL18_II", "SSTL15_I", "SSTL15_II", "HSTL18_I", "HSTL18_II", "HSTL15_I", "SSTL15_I_CAL", "SSTL15_II_CAL", "HSTL15_I_CAL", "DEFAULT" :;
    default : begin
           $display("Attribute Syntax Error : The attribute IOSTANDARD on GTP_OUTBUF instance %m is set to %s.", IOSTANDARD);
           $finish;
              end
    endcase

    case (SLEW_RATE)
    "SLOW", "FAST":;
    default : begin
           $display("Attribute Syntax Error : The attribute SLEW_RATE on GTP_OUTBUF instance %m is set to %s.", SLEW_RATE);
           $finish;
              end
    endcase

    case (DRIVE_STRENGTH)
    "2", "4", "6", "8", "12", "16", "24":;
    default : begin
           $display("Attribute Syntax Error : The attribute DRIVE_STRENGTH on GTP_OUTBUF instance %m is set to %s.", DRIVE_STRENGTH);
           $finish;
              end
    endcase
    end

    buf (O, I);

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_SCANCHAIN_E1.v
//
// Functional description: JTAG TAP Controller simulation model
//
// Parameter description:
//      
//
// Port description:
//      
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale  1 ns / 1 ps

module GTP_SCANCHAIN_E1
#(
    parameter [31:0] IDCODE = 32'haaaa5555, //dr idcode
    parameter   CHAIN_NUM = 1 //1 2 3 4 available
)
(
    input      TCK      ,//JTAG signals
    input      TDI      ,
    input      TMS      ,
    output reg TDO      ,
    
    output reg CAPDR    ,//scanchain signals
    output     JCLK     ,
    output reg RST      ,
    output reg FLG_USER ,
    output reg SHFTDR   ,
    output     TDI_USER ,
    output     TCK_USER ,
    output     TMS_USER ,
    output reg JRTI     ,
    output reg UPDR     ,
    input      TDO_USER 
);

wire           flg_capture_ir  ;
wire           flg_shift_ir    ;
wire           flg_update_ir   ;
wire           flg_capture_dr  ;
wire           flg_shift_dr    ;
wire           flg_update_dr   ;
wire           flg_idcode      ;
wire           flg_bypass      ;
wire           flg_bypass_highz;

wire           irq             ;
wire           drq_bypass      ;
wire           drq_idcode      ;
wire	       flg_user        ;

reg    [3:0]   s               ;
reg    [3:0]   ns              ;

//reg            flg_jclk        ;
reg    [9:0]   USER	       ;
reg    [9:0]   shift_ir        ;
reg    [9:0]   update          ;

wire           flg_highz       ;


//////////JTAG signals///////////
reg            JTAG_USER = 1'bz;

localparam TEST_LOGIC_RESET  =  4'd0 ,
           RUN_TEST_IDLE     =  4'd1 ,
           SELECT_IR_SCAN    =  4'd2 ,
           CAPTURE_IR        =  4'd3 ,
           SHIFT_IR          =  4'd4 ,
           EXIT1_IR          =  4'd5 ,
           PAUSE_IR          =  4'd6 ,
           EXIT2_IR          =  4'd7 ,
           UPDATE_IR         =  4'd8 ,
           SELECT_DR_SCAN    =  4'd9 ,
           CAPTURE_DR        =  4'd10,
           SHIFT_DR          =  4'd11,
           EXIT1_DR          =  4'd12,
           PAUSE_DR          =  4'd13,
           EXIT2_DR          =  4'd14,
           UPDATE_DR         =  4'd15;

localparam USER1                =  10'b10_1000_0110, // Access user-defined register 1
           USER2                =  10'b10_1000_0111, // Access user-defined register 2
           USER3                =  10'b10_1000_1000, // Access user-defined register 3
           USER4                =  10'b10_1000_1001, // Access user-defined register 4
           ID_CODE               =  10'b10_1000_0011, // Enables shifting out of ID code
           HIGHZ                =  10'b10_1000_0101, // 3-state output pins while enabling
           BYPASS               =  10'b11_1111_1111; // Enables BYPASS


                    
initial 
     begin
       case (CHAIN_NUM)
           1: USER <= USER1;
           2: USER <= USER2;
           3: USER <= USER3;
           4: USER <= USER4;
     default: 
            $display("Error: CHAIN_NUM is not available");
endcase
end
           


/*always @(posedge TCK)
       begin
          scanchain <= SCANCHAIN;
end
*/
always @(posedge TCK)
    begin
        s <= ns;
    end

always @(*)
    begin
        case(s)
            TEST_LOGIC_RESET:
                begin
                    if(TMS)
                        ns = TEST_LOGIC_RESET;
                    else
                        ns = RUN_TEST_IDLE;
                end

            RUN_TEST_IDLE:
                begin
                    if(TMS)
                        ns = SELECT_DR_SCAN;
                    else
                        ns = RUN_TEST_IDLE;
                end

            SELECT_IR_SCAN:
                begin
                    if(TMS)
                        ns = TEST_LOGIC_RESET;
                    else
                        ns = CAPTURE_IR;
                end

            CAPTURE_IR, SHIFT_IR:
                begin
                    if(TMS)
                        ns = EXIT1_IR;
                    else
                        ns = SHIFT_IR;
                end
            
            EXIT1_IR:
                begin
                    if(TMS)
                        ns = UPDATE_IR;
                    else
                        ns = PAUSE_IR;
                end

            PAUSE_IR:
                begin
                    if(TMS)
                        ns = EXIT2_IR;
                    else
                        ns = PAUSE_IR;
                end

            EXIT2_IR:
                begin
                    if(TMS)
                        ns = UPDATE_IR;
                    else
                        ns = SHIFT_IR;
                end

            UPDATE_IR, UPDATE_DR:
                begin
                    if(TMS)
                        ns = SELECT_DR_SCAN;
                    else
                        ns = RUN_TEST_IDLE;
                end

            SELECT_DR_SCAN:
                begin
                    if(TMS)
                        ns = SELECT_IR_SCAN;
                    else
                        ns = CAPTURE_DR;
                end

            CAPTURE_DR, SHIFT_DR:
                begin
                    if(TMS)
                        ns = EXIT1_DR;
                    else
                        ns = SHIFT_DR;
                end

            EXIT1_DR:
                begin
                    if(TMS)
                        ns = UPDATE_DR;
                    else
                        ns = PAUSE_DR;
                end

            PAUSE_DR:
                begin
                    if(TMS)
                        ns = EXIT2_DR;
                    else
                        ns = PAUSE_DR;
                end

            EXIT2_DR:
                begin
                    if(TMS)
                        ns = UPDATE_DR;
                    else
                        ns = SHIFT_DR;
                end
        default: 
               ns = TEST_LOGIC_RESET;
        endcase
    end

always @(negedge TCK)
    begin
        if(s == TEST_LOGIC_RESET)
            RST <= 1'b1;
        else
            RST <= 1'b0;
    end
always @(negedge TCK)
    begin
        if(s == RUN_TEST_IDLE)
            JRTI <= 1'b1;
        else
            JRTI <= 1'b0;
    end       
assign flg_capture_ir = (s == CAPTURE_IR);
assign flg_shift_ir   = (s == SHIFT_IR  );
assign flg_update_ir  = (s == UPDATE_IR );
assign flg_capture_dr = (s == CAPTURE_DR);
assign flg_shift_dr   = (s == SHIFT_DR  );
assign flg_update_dr  = (s == UPDATE_DR );


always @(posedge TCK)
    begin
        if(RST)
            shift_ir <= 10'd0;
        else if(flg_capture_ir)
            shift_ir <= 10'd0;
        else if(flg_shift_ir)
            shift_ir <= {TDI, shift_ir[9:1]};
    end

assign irq = shift_ir[0];

always @(negedge TCK)
    begin
        if(RST)
            update <= ID_CODE;//ir idcode
        else if(flg_update_ir)
            update <= shift_ir;
    end

assign flg_user                 =  (update == USER );
assign flg_idcode               =  (update == ID_CODE);
assign flg_bypass               =  (update == BYPASS);
assign flg_highz                =  (update == HIGHZ );
assign flg_bypass_highz         =  flg_bypass | flg_highz;

reg    shift_bypass;
assign drq_bypass = shift_bypass;

always @(posedge TCK)
    begin
        if(RST)
            shift_bypass <= 1'b0;
        else if(flg_bypass_highz)
            begin
                if(flg_capture_dr)
                    shift_bypass <= 1'b0;
                else if(flg_shift_dr)
                    shift_bypass <= TDI;
            end
    end


reg    [31:0]    shift_id;
assign drq_idcode = shift_id[0];

always @(posedge TCK)
    begin
        if(RST)
            shift_id <= 32'd0;
        else if(flg_idcode)
            begin
                if(flg_capture_dr)
                    shift_id <= IDCODE;//dr idcode
                else if(flg_shift_dr)
                    shift_id <= {TDI, shift_id[31:1]};
                else
                    shift_id <= 32'd0;
            end
        else
            shift_id <= 32'd0;
    end


always @(negedge TCK)
    begin
        if(RST)
            begin
                CAPDR  <= 1'b0;
                SHFTDR <= 1'b0;
                UPDR   <= 1'b0;
            end
        else
            begin
                CAPDR  <= flg_capture_dr;
                SHFTDR <= flg_shift_dr  ;
                UPDR   <= flg_update_dr ;
            end
    end

//always @(negedge TCK)
//    begin
//        if(RST)
//            flg_jclk <= 1'b0;
//        else if(CAPDR)
//            flg_jclk <= 1'b1;
//        else if(UPDR)
//            flg_jclk <= 1'b0;
//    end

//assign JCLK = flg_user & (CAPDR | flg_jclk) & TCK;
assign JCLK = flg_user & (CAPDR | SHFTDR) & TCK;

always @(negedge TCK)
    begin
        if(RST)
            TDO <= 1'b0;
        else if(flg_shift_ir)
            TDO <= irq;
        else if(flg_shift_dr)
            case({flg_bypass_highz, flg_idcode, flg_user})
                3'b10_0: TDO <= drq_bypass;
                3'b01_0: TDO <= drq_idcode;
                3'b00_1: TDO <= TDO_USER;
                default: TDO <= 1'b0;
            endcase
    end
always@(*)

	begin 
		FLG_USER <= flg_user;
	end
////////////////////user tdo//////////
always@(*)
	begin
		JTAG_USER <= TDO_USER;
end
assign TDI_USER = TDI;
assign TCK_USER = TCK;
assign TMS_USER = TMS;

endmodule









//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS REVERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//Description:
//$Author: xqlin
//$Reversion:
//  2019/09/10: Initial Version.
//////////////////////////////////////////////////////////////////////////////
`timescale 1ns / 1ps
module GTP_DLL_E2 #(
    parameter           GRS_EN              = "TRUE",   //TRUE, FALSE;
    parameter   [7:0]   CAL_INIT            = 8'b00011111,
    parameter           DELAY_STEP_OFFSET   = 0,        // CP_CODE_OFFSET: -4 -3 -2 -1 0 1 2 3 4
    parameter           DELAY_SEL           = 1'b0,
    parameter           FAST_LOCK           = "FALSE",
    parameter   [1:0]   FDIV                = 2'b10, 
    parameter           INT_CLK             = 1'b0,
    parameter   [1:0]   UPD_DLY             = 2'b01
)(
    input           CLKIN,   // IOCLK_2X
    input           SYS_CLK,   // SYSCLK
    input           PWD,    // DLL_FREEZE
    input           RST,
    input           UPDATE_N,
    output          LOCK,
    output  [7:0]   DELAY_STEP,          // DLL_90CODE_GRAY
    output  [7:0]   DELAY_STEP1          // DLL_45CODE_GRAY
    )/* synthesis syn_black_box */;

   //synthesis translate_off


    wire   [7:0]    SC_CAL_INIT;
    reg    [3:0]    SC_CODE_OFFSET;
    wire            SC_DELAY_SEL;
    reg             SC_FAST_LOCK;
    wire   [1:0]    SC_FDIV;
    wire            SC_INT_CLK;
    wire   [1:0]    SC_UPD_DLY;
    wire   [1:0]    SC_LDO_CTRL;

    wire            grs_n;
    wire            dll_rstn;
    wire            ioclk_0p5x;
    wire            ioclk_0p5x_dly0;
    wire            ioclk_0p5x_dly1;
    wire            ioclk_0p5x_dly2;
    wire            ioclk_0p5x_dly;
    wire            ioclk_0p5x_mindly;
    wire    [63:0]  dly_cal_therm;
    wire            up_dnb;
    wire            rst_n;

    initial
        begin
            if ((GRS_EN == "TRUE")  || (GRS_EN == "FALSE")) begin
            end
            else
                $display ("error: illegal setting for GRS_EN");
        
            if ((FAST_LOCK == "TRUE")  || (FAST_LOCK == "FALSE")) begin
            end
            else
                $display ("error: illegal setting for FAST_LOCK");
        
            if ((DELAY_STEP_OFFSET == -4)  || (DELAY_STEP_OFFSET == -3) || (DELAY_STEP_OFFSET == -2)  || (DELAY_STEP_OFFSET == -1) ||(DELAY_STEP_OFFSET == 0)  || (DELAY_STEP_OFFSET == 1) ||(DELAY_STEP_OFFSET == 2)  || (DELAY_STEP_OFFSET == 3) ||(DELAY_STEP_OFFSET == 4)) begin
            end
            else
                $display ("error: illegal setting for DELAY_STEP_OFFSET");
        end


    assign grs_n    = (GRS_EN == "TRUE") ? GRS_INST.GRSNET : 1'b1;
    //assign grs_n    = 1'b1;
    assign dll_rstn = ~(~grs_n || RST);
    assign rst_n    = ~(PWD || ~dll_rstn);

    dll_e2_ddrphy_dll_fdiv fdiv(
	.ioclk_2x(CLKIN),
	.rst_n(rst_n),
	.sc_fdiv(SC_FDIV),
	.ioclk_div_out(ioclk_0p5x)
    );

    dll_e2_dly_chain #(.dly_en(1'b1), .dly_sel(DELAY_SEL))    U0_DLY(.therm_code(dly_cal_therm), .din(ioclk_0p5x),       .d_dly(ioclk_0p5x_dly0));
    dll_e2_dly_chain #(.dly_en(1'b1), .dly_sel(DELAY_SEL))    U1_DLY(.therm_code(dly_cal_therm), .din(ioclk_0p5x_dly0),  .d_dly(ioclk_0p5x_dly1));
    dll_e2_dly_chain #(.dly_en(1'b1), .dly_sel(DELAY_SEL))    U2_DLY(.therm_code(dly_cal_therm), .din(ioclk_0p5x_dly1),  .d_dly(ioclk_0p5x_dly2));
    dll_e2_dly_chain #(.dly_en(1'b1), .dly_sel(DELAY_SEL))    U3_DLY(.therm_code(dly_cal_therm), .din(ioclk_0p5x_dly2),  .d_dly(ioclk_0p5x_dly));
    dll_e2_dly_chain #(.dly_en(1'b1), .dly_sel(DELAY_SEL))    U4_DLY(.therm_code({64{1'b0}}),    .din(ioclk_0p5x),       .d_dly(ioclk_0p5x_mindly));
    dll_e2_DLL_DFF   U0_DFF(.CLK(ioclk_0p5x_dly),   .DIN(ioclk_0p5x_mindly),   .RSTN(!RST), .Q(up_dnb));
    
    dll_e2_ddrphy_dll_fsm  fsm(
    .sc_dll_force(1'b0),
    .sc_code_offset(SC_CODE_OFFSET),
    .sc_fast_lock(SC_FAST_LOCK),
    .sc_int_clk(SC_INT_CLK),
    .sc_cal_init(SC_CAL_INIT),
    .sc_upd_dly(SC_UPD_DLY),
    .sys_clk(SYS_CLK),
    .ioclk_2x(CLKIN),
    .rst_n(!RST),
    .glogen(1'b1),
    .up_dnb(up_dnb),
    .update_n(UPDATE_N),
    .dll_freeze(PWD),
    .dll_90code_gray(DELAY_STEP),
    .dll_45code_gray(DELAY_STEP1),
    .lock(LOCK),
    .therm_code(dly_cal_therm)
    );

    ////////////CP2SC/////////////////////////   
//    always @( * )                           //                        
//    begin                                   // 
//       if(DLL_FORCE == "FALSE")          // 
//       begin                                //
//           SC_DLL_FORCE = 1'b0;             //
//       end                                  //
//       else if(DLL_FORCE == "TRUE")      //
//       begin                                //
//           SC_DLL_FORCE = 1'b1;             //
//       end                                  //
//       else                                 //
//       begin                                //
//           SC_DLL_FORCE = 1'bx;             //
//       end                                  //
//    end                                     //
                                            //
initial begin                                   //
       if(FAST_LOCK == "FALSE")              //
       begin                                //
           SC_FAST_LOCK = 1'b0;             //
       end                                  //
       else if(FAST_LOCK == "TRUE")         //
       begin                                //
           SC_FAST_LOCK = 1'b1;             //
       end                                  //
       else                                 //
       begin                                //
           SC_FAST_LOCK = 1'bx;             //
       end                                  //
    end                                     //
                                            //
    assign  SC_FDIV[0]    = FDIV[0];     //
                                            //
    assign  SC_FDIV[1]    = FDIV[1];     //
                                            //
    assign  SC_INT_CLK    = INT_CLK;     //
                                            //
    assign  SC_UPD_DLY[0] = UPD_DLY[0];  //
                                            //
    assign  SC_UPD_DLY[1] = UPD_DLY[1];  //
                                            //
    assign  SC_DELAY_SEL      = DELAY_SEL;     //
                                            //
    assign  SC_CAL_INIT[0] = CAL_INIT[0];//
                                            //
    assign  SC_CAL_INIT[1] = CAL_INIT[1];//
                                            //
    assign  SC_CAL_INIT[2] = CAL_INIT[2];//
                                            //
    assign  SC_CAL_INIT[3] = CAL_INIT[3];//
                                            //
    assign  SC_CAL_INIT[4] = CAL_INIT[4];//
                                            //
    assign  SC_CAL_INIT[5] = CAL_INIT[5];//
                                            //
    assign  SC_CAL_INIT[6] = CAL_INIT[6];//
                                            //
    assign  SC_CAL_INIT[7] = CAL_INIT[7];//
                                            //////// 

    initial begin
        case (DELAY_STEP_OFFSET)
            -4 : SC_CODE_OFFSET = 4'b1111;
            -3 : SC_CODE_OFFSET = 4'b1110;
            -2 : SC_CODE_OFFSET = 4'b1101;
            -1 : SC_CODE_OFFSET = 4'b1100;
             0 : SC_CODE_OFFSET = 4'b0000;
             1 : SC_CODE_OFFSET = 4'b1000;
             2 : SC_CODE_OFFSET = 4'b1001;
             3 : SC_CODE_OFFSET = 4'b1010;
             4 : SC_CODE_OFFSET = 4'b1011;
            default :SC_CODE_OFFSET = 4'b0000;
        endcase
    end

//    assign  SC_CODE_OFFSET[0] = DELAY_STEP_OFFSET[0];//
//                                                  //
//    assign  SC_CODE_OFFSET[1] = DELAY_STEP_OFFSET[1];//
//                                                  //
//    assign  SC_CODE_OFFSET[2] = DELAY_STEP_OFFSET[2];//
//                                                  //
//    assign  SC_CODE_OFFSET[3] = DELAY_STEP_OFFSET[3];//
    ////////////////////////////////////////////////
    //synthesis translate_on
endmodule




    




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_IOBUFCO.v
//
// Functional description: Differential Signaling Input/Output Buffer
//
// Parameter description:
//
// Port description:
//
// Revision:
//    06/18/14 - Initial version.
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_IOBUFCO #(
    parameter IOSTANDARD = "DEFAULT",
    parameter TERM_DDR = "ON"
)(
    output reg O,
    inout IO,
    inout IOB,
    input I,
    input T
) /* synthesis syn_black_box */ ;
  
  initial begin
    case (IOSTANDARD)
    "SSTL18D_I", "SSTL18D_II", "SSTL15D_I", "SSTL15D_II", "HSTL15D_I", "SSTL25D_I", "SSTL25D_II", "SSTL15D_I_CAL", "SSTL15D_II_CAL", "HSTL15D_I_CAL", "LVPECL", "RSDS", "PPDS", "BLVDS", "LVCMOS25D", "LVCMOS33D","LVDS25E", "DEFAULT":;
    default : begin
           $display("Attribute Syntax Error : The attribute IOSTANDARD on GTP_IOBUFCO instance %m is set to %s.", IOSTANDARD);
           $finish;
              end
    endcase

    case (TERM_DDR)
    "ON", "OFF" :;
    default : begin
           $display("Attribute Syntax Error : The attribute TERM_DDR on GTP_IOBUFCO instance %m is set to %s.", TERM_DDR);
           $finish;
              end
    endcase
    end 
    bufif0 (IO, I, T);
    notif0 (IOB, I, T);

    always @(*)
    begin
        if (IO == 1'b1 && IOB == 1'b0)
            O = IO;
        else if (IO == 1'b0 && IOB == 1'b1)
            O = IO;
        else
            O = 1'bx;
    end

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2016 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_ISERDES_E2.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//////////////////////////////////////////////////////////////////////////////
`timescale 1ps / 1ps

module GTP_ISERDES_E2 #(
    parameter         ISERDES_MODE     =   "SDR1TO4",       // "SDR1TO2","SDR1TO3","SDR1TO4","SDR1TO5","SDR1TO6","SDR1TO7","SDR1TO8",
                                                            // "DDR1TO2_SAME_PIPELINED", "DDR1TO2_SAME_EDGE", "DDR1TO2_OPPOSITE_EDGE",
                                                            // "DDR1TO4","DDR1TO6","DDR1TO8","DDR1TO10","DDR1TO14",
                                                            // "HMDDR1TO4","HMDDR1TO8",
                                                            // "LMDDR1TO4","LMDDR1TO8",
                                                            // "OVERSAMPLE","ILATCH","IDFF",

    parameter         CASCADE_MODE     =   "MASTER",        // "MASTER" ,"SLAVE"
    parameter         BITSLIP_EN       =   "FALSE",       // "FALSE","TRUE"
    parameter         GRS_EN           =   "TRUE",          // "TRUE", "FALSE"
    parameter         NUM_ICE          =   1'b0,            // 1'b1 , 1'b0
    parameter         GRS_TYPE_Q0      =   "RESET",         // SET  RESET 
    parameter         GRS_TYPE_Q1      =   "RESET",         // SET  RESET 
    parameter         GRS_TYPE_Q2      =   "RESET",         // SET  RESET 
    parameter         GRS_TYPE_Q3      =   "RESET",         // SET  RESET 
    parameter         LRS_TYPE_Q0      =   "ASYNC_RESET",   // ASYNC_SET  ASYNC_RESET  SYNC_SET SYNC_RESET
    parameter         LRS_TYPE_Q1      =   "ASYNC_RESET",   // ASYNC_SET  ASYNC_RESET  SYNC_SET SYNC_RESET
    parameter         LRS_TYPE_Q2      =   "ASYNC_RESET",   // ASYNC_SET  ASYNC_RESET  SYNC_SET SYNC_RESET
    parameter         LRS_TYPE_Q3      =   "ASYNC_RESET"    // ASYNC_SET  ASYNC_RESET  SYNC_SET SYNC_RESET  

)(
    //input        GRS_N,
    input        RST,
    input        ICE0,
    input        ICE1,
    input        DESCLK,
    input        ICLK,
    //input        ICLKB,
    input        OCLK,
    //input        OCLKB,
    input        ICLKDIV,
    input        DI,
    input        BITSLIP,
    input        ISHIFTIN0,
    input        ISHIFTIN1,
    input  [2:0] IFIFO_WADDR,
    input  [2:0] IFIFO_RADDR,
    output [7:0] DO,
    output       ISHIFTOUT0,
    output       ISHIFTOUT1
);

wire        gwen;
wire        glogen;
wire        grs_n;
wire        isr_iolhr;
wire        ice0;
wire        ice1;
wire        desclk;
wire        iclk;
wire        iclkb;
wire        oclk;
wire        oclkb;
wire        iclkdiv;
wire        dyn_clkpol;
wire        dyn_clkdivpol;
wire        di;
wire        di_n;
wire        di_mipi;
wire        di_from_srb;
wire        ofb;
wire        tfb;
wire        bitslip;
wire        ishiftin0;
wire        ishiftin1;
wire  [2:0] ififo_waddr;
wire  [2:0] ififo_raddr;
wire        dly_idly_in;
wire        dly_zhold_in;
reg         desclk_reg;
reg         sc_div_en;

assign  gwen         =  1'b1;
assign  glogen       =  1'b1;
assign  grs_n        =  (GRS_EN == "TRUE") ? GRS_INST.GRSNET : 1'b1;
//assign  grs_n        =  1'b1;
//assign  grs_n        =  GRS_N;
assign  isr_iolhr    =  RST;
assign  ice0         =  ICE0;
assign  ice1         =  ICE1;
assign  desclk       =  sc_div_en ? desclk_reg : DESCLK;
assign  iclk         =  ICLK;
assign  iclkb        =  ~ICLK;
assign  oclk         =  OCLK;
assign  oclkb        =  ~OCLK;
assign  iclkdiv      =  ICLKDIV;
assign  dyn_clkpol   =  1'b1;
assign  dyn_clkdivpol=  1'b1;
assign  di           =  DI;
assign  di_n         =  ~DI;
assign  di_mipi      =  1'b0;
assign  di_from_srb  =  1'b0;
assign  ofb          =  1'b0;
assign  tfb          =  1'b0;
assign  bitslip      =  BITSLIP;
assign  ishiftin0    =  ISHIFTIN0;
assign  ishiftin1    =  ISHIFTIN1;
assign  ififo_waddr  =  IFIFO_WADDR;
assign  ififo_raddr  =  IFIFO_RADDR;

wire       rstn_out;
wire [7:0] rx_data;
wire       ishiftout0;
wire       ishiftout1;

assign  DO	         = rx_data;
assign  ISHIFTOUT0	 = ishiftout0;
assign  ISHIFTOUT1	 = ishiftout1;

wire      gsr;
//wire      rstn;
wire      lsr_sync;
wire      lsr_async;
wire      ce_hsmem;
wire      ce_out_0;
wire      ce_out_1;
wire      clk_stg0;
wire      clkb_stg0;
wire      hsmem_clk;
wire      hsmem_clkb;
wire      clk_stg1_0;
wire      clk_stg1_1;
wire      clk_stg1_2;
wire      clk_stg2_0;
wire      clk_stg2_1;
wire      clk_stg3;
wire      clk_for_bs;
wire       bsclk;
wire [4:0] sel0;
wire       sel1;
wire [2:0] sel2;
wire [1:0] sel3;
wire [2:0] sel4;
wire [3:0] sel5;
wire [1:0] sel6;
wire       sdr1to2;
wire       sdr1to3;
wire       sdr1to4;
wire       sdr1to5;
wire       sdr1to6;
wire       sdr1to7;
wire       sdr1to8;
wire       ddr1to4;
wire       ddr1to6;
wire       ddr1to8;
wire       ddr1to10;
wire       ddr1to14;


wire       di_to_gear;

wire        sc_dyn_clkpol;
wire        sc_dyn_clkdivpol;
wire        sc_clk_pol0;
wire        sc_clk_pol1;
wire        sc_clk_pol2;
wire        sc_clk_pol3;
wire        sc_oclkpol;
wire        sc_oclkbpol;
wire        sc_d_pol0;
wire        sc_d_pol1;
wire        sc_d_sel0;
wire        sc_d_sel1;
wire        sc_d_sel2;
wire        sc_d_sel3;
wire  [1:0] sc_d_sel4;
wire  [1:0] sc_d_sel5;
wire  [1:0] sc_d_sel6;
wire        sc_test_en0;
wire        sc_test_en1;
wire        sc_mipi_en;
wire        sc_master;
wire        sc_bitslip_en;
wire        sc_isr_pol;
wire        sc_isr_en;
wire        sc_grs_dis;
wire        sc_num_ice;

reg         sc_isr_sync;
reg   [3:0] sc_init_q;
reg   [3:0] sc_srval_q;

reg   [3:0] sc_iserdes_mode;
reg         sc_ddri_en;
reg         sc_des_sdren;
reg         sc_des_ddren;
reg         sc_networking_en;
reg         sc_ihsmem_en;
reg         sc_ififo_en;
reg         sc_lsmem_en;
reg         sc_oversample_en;
reg         sc_samepipeline_en;
reg         sc_isame_en;
reg         sc_iopposite_en;
reg         sc_ilthen;
reg         sc_idffen;

assign  sc_dyn_clkpol		 = 1'b0;
assign  sc_dyn_clkdivpol	 = 1'b0;
assign  sc_clk_pol0		     = 1'b0;
assign  sc_clk_pol1		     = 1'b0;
assign  sc_clk_pol2		     = 1'b0;
assign  sc_clk_pol3		     = 1'b0;
assign  sc_oclkpol		     = 1'b0;
assign  sc_oclkbpol		     = 1'b0;
assign  sc_d_pol0		     = 1'b0;
assign  sc_d_pol1		     = 1'b0;
assign  sc_d_sel0		     = 1'b0;    // di
assign  sc_d_sel1		     = 1'b0;
assign  sc_d_sel2		     = 1'b0;
assign  sc_d_sel3		     = 1'b0;
assign  sc_d_sel4		     = 2'b01;   // 00:zhold_delay; 01:IOB; 10:idelay; 11:set 0 
assign  sc_d_sel5		     = 2'b01;   // 00:zhold_delay; 01:IOB; 10:idelay; 11:set 0 
assign  sc_d_sel6		     = 2'b00;   // 00:IOB;         01:SRB; 10:ofb;    11:idelay
assign  sc_test_en0		     = 1'b0;
assign  sc_test_en1		     = 1'b0;
assign  sc_mipi_en		     = 1'b0;
assign  sc_master		     = (CASCADE_MODE    == "MASTER" ) ? 1'b0 : 1'b1;
assign  sc_bitslip_en		 = (BITSLIP_EN      == "FALSE") ? 1'b0 : 1'b1;
assign  sc_isr_pol           = 1'b0;
assign  sc_isr_en		     = 1'b1;
assign  sc_grs_dis		     = (GRS_EN          == "TRUE"  ) ? 1'b0 : 1'b1; // GRS_DIS --> GRS_EN
assign  sc_num_ice		     = NUM_ICE;

initial begin

//    if(MIPI_EN != "TRUE" && MIPI_EN != "FALSE")
//    begin $display("Error: Illegal setting MIPI_EN of %s",MIPI_EN);$finish;end

    if(CASCADE_MODE != "MASTER" && CASCADE_MODE != "SLAVE")
    begin $display("Error: Illegal setting CASCADE_MODE of %s",CASCADE_MODE);$finish;end

    if(BITSLIP_EN != "TRUE" && BITSLIP_EN != "FALSE")
    begin $display("Error: Illegal setting BITSLIP_EN of %s",BITSLIP_EN);$finish;end

    if(GRS_EN != "TRUE" && GRS_EN != "FALSE")
    begin $display("Error: Illegal setting GRS_EN of %s",GRS_EN);$finish;end

    if(NUM_ICE != 1'b0 && NUM_ICE != 1'b1)
    begin $display("Error: Illegal setting NUM_ICE of %b",NUM_ICE);$finish;end

    if(GRS_TYPE_Q0 != "SET" && GRS_TYPE_Q0 != "RESET")
    begin $display("Error: Illegal setting GRS_TYPE_Q0 of %s",GRS_TYPE_Q0);$finish;end

    if(GRS_TYPE_Q1 != "SET" && GRS_TYPE_Q1 != "RESET")
    begin $display("Error: Illegal setting GRS_TYPE_Q1 of %s",GRS_TYPE_Q1);$finish;end

    if(GRS_TYPE_Q2 != "SET" && GRS_TYPE_Q2 != "RESET")
    begin $display("Error: Illegal setting GRS_TYPE_Q2 of %s",GRS_TYPE_Q2);$finish;end

    if(GRS_TYPE_Q3 != "SET" && GRS_TYPE_Q3 != "RESET")
    begin $display("Error: Illegal setting GRS_TYPE_Q3 of %s",GRS_TYPE_Q3);$finish;end

    if(LRS_TYPE_Q0 != "ASYNC_SET" && LRS_TYPE_Q0 != "ASYNC_RESET" && LRS_TYPE_Q0 != "SYNC_SET" && LRS_TYPE_Q0 != "SYNC_RESET")
    begin $display("Error: Illegal setting LRS_TYPE_Q0 of %s",LRS_TYPE_Q0);$finish;end

    if(LRS_TYPE_Q1 != "ASYNC_SET" && LRS_TYPE_Q1 != "ASYNC_RESET" && LRS_TYPE_Q1 != "SYNC_SET" && LRS_TYPE_Q1 != "SYNC_RESET")
    begin $display("Error: Illegal setting LRS_TYPE_Q1 of %s",LRS_TYPE_Q1);$finish;end

    if(LRS_TYPE_Q2 != "ASYNC_SET" && LRS_TYPE_Q2 != "ASYNC_RESET" && LRS_TYPE_Q2 != "SYNC_SET" && LRS_TYPE_Q2 != "SYNC_RESET")
    begin $display("Error: Illegal setting LRS_TYPE_Q2 of %s",LRS_TYPE_Q2);$finish;end

    if(LRS_TYPE_Q3 != "ASYNC_SET" && LRS_TYPE_Q3 != "ASYNC_RESET" && LRS_TYPE_Q3 != "SYNC_SET" && LRS_TYPE_Q3 != "SYNC_RESET")
    begin $display("Error: Illegal setting LRS_TYPE_Q3 of %s",LRS_TYPE_Q3);$finish;end


    if((LRS_TYPE_Q0 == "ASYNC_RESET" || LRS_TYPE_Q0 == "ASYNC_SET" || LRS_TYPE_Q1 == "ASYNC_RESET" || LRS_TYPE_Q1 == "ASYNC_SET" 
        || LRS_TYPE_Q2 == "ASYNC_RESET" || LRS_TYPE_Q2 == "ASYNC_SET" || LRS_TYPE_Q3 == "ASYNC_RESET" || LRS_TYPE_Q3 == "ASYNC_SET") 
        && (LRS_TYPE_Q0 == "SYNC_RESET" || LRS_TYPE_Q0 == "SYNC_SET" || LRS_TYPE_Q1 == "SYNC_RESET" || LRS_TYPE_Q1 == "SYNC_SET" 
        ||  LRS_TYPE_Q2 == "SYNC_RESET" || LRS_TYPE_Q2 == "SYNC_SET" || LRS_TYPE_Q3 == "SYNC_RESET" || LRS_TYPE_Q3 == "SYNC_SET"))
    begin $display("Error: LRS_TYPE_Qx must be all of ASYNC_ or SYNC_.");$finish;end

end

// sc_iserdes_mode
initial begin
// default value
    sc_iserdes_mode  = 4'b0000; 
    sc_ddri_en       = 1'b0;
    sc_des_sdren     = 1'b0;
    sc_des_ddren     = 1'b0;
    sc_networking_en = 1'b0;
    sc_ihsmem_en     = 1'b0;
    sc_ififo_en      = 1'b0;
    sc_lsmem_en      = 1'b0;
    sc_oversample_en = 1'b0;
    sc_samepipeline_en = 1'b0;
    sc_isame_en		 = 1'b0;
    sc_iopposite_en	 = 1'b0;
    sc_ilthen		 = 1'b0;
    sc_idffen	     = 1'b0;
    sc_div_en	     = 1'b0;
    desclk_reg	     = 1'b0;

    case (ISERDES_MODE)
// Networking Mode
        "SDR1TO2" :begin 
                    sc_iserdes_mode  = 4'b0101;
                    sc_ddri_en       = 1'b1;
                    sc_des_sdren     = 1'b1;
                    sc_networking_en = 1'b1;
                    sc_div_en        = 1'b0;
                   end
        "SDR1TO3" :begin
                    sc_iserdes_mode  = 4'b0110;
                    sc_ddri_en       = 1'b1;
                    sc_des_sdren     = 1'b1;
                    sc_networking_en = 1'b1;
                    sc_div_en        = 1'b0;
                   end
        "SDR1TO4" :begin
                    sc_iserdes_mode  = 4'b0000;
                    sc_ddri_en       = 1'b1;
                    sc_des_sdren     = 1'b1;
                    sc_networking_en = 1'b1;
                    sc_div_en        = 1'b0;
                   end
        "SDR1TO5" :begin
                    sc_iserdes_mode  = 4'b0011;
                    sc_ddri_en       = 1'b1;
                    sc_des_sdren     = 1'b1;
                    sc_networking_en = 1'b1;
                    sc_div_en        = 1'b0;
                   end
        "SDR1TO6" :begin
                    sc_iserdes_mode  = 4'b1000;
                    sc_ddri_en       = 1'b1;
                    sc_des_sdren     = 1'b1;
                    sc_networking_en = 1'b1;
                    sc_div_en        = 1'b0;
                   end
        "SDR1TO7" :begin
                    sc_iserdes_mode  = 4'b0010;
                    sc_ddri_en       = 1'b1;
                    sc_des_sdren     = 1'b1;
                    sc_networking_en = 1'b1;
                    sc_div_en        = 1'b0;
                   end
        "SDR1TO8" :begin
                    sc_iserdes_mode  = 4'b0001;
                    sc_ddri_en       = 1'b1;
                    sc_des_sdren     = 1'b1;
                    sc_networking_en = 1'b1;
                    sc_div_en        = 1'b0;
                   end
// DDR 
        "ILATCH": begin
                    sc_ddri_en      = 1'b0;
                    sc_ilthen       = 1'b1;
                    sc_div_en       = 1'b0;
                   end
        "IDFF": begin
                    sc_ddri_en      = 1'b0;
                    sc_idffen       = 1'b1;
                    sc_div_en       = 1'b0;
                   end
        "DDR1TO2_SAME_PIPELINED": begin
                    sc_ddri_en          = 1'b0;
                    sc_des_ddren        = 1'b1;
                    sc_samepipeline_en  = 1'b1;
                    sc_div_en           = 1'b0;
                   end
        "DDR1TO2_SAME_EDGE": begin
                    sc_ddri_en       = 1'b0;
                    sc_des_ddren     = 1'b1;
                    sc_isame_en		 = 1'b1;
                    sc_div_en        = 1'b0;
                   end
        "DDR1TO2_OPPOSITE_EDGE": begin
                    sc_ddri_en       = 1'b0;
                    sc_des_ddren     = 1'b1;
                    sc_iopposite_en	 = 1'b1;
                    sc_div_en        = 1'b0;
                   end
        "DDR1TO4": begin
                    sc_iserdes_mode  = 4'b0000;
                    sc_ddri_en       = 1'b1;
                    sc_des_ddren     = 1'b1;
                    sc_networking_en = 1'b1;
                    sc_div_en        = 1'b0;
                   end
        "DDR1TO6": begin
                    sc_iserdes_mode  = 4'b1000;
                    sc_ddri_en       = 1'b1;
                    sc_des_ddren     = 1'b1;
                    sc_networking_en = 1'b1;
                    sc_div_en        = 1'b0;
                   end
        "DDR1TO8": begin
                    sc_iserdes_mode  = 4'b0001;
                    sc_ddri_en       = 1'b1;
                    sc_des_ddren     = 1'b1;
                    sc_networking_en = 1'b1;
                    sc_div_en        = 1'b0;
                   end
        "DDR1TO10":begin
                    sc_iserdes_mode  = 4'b0100;
                    sc_ddri_en       = 1'b1;
                    sc_des_ddren     = 1'b1;
                    sc_networking_en = 1'b1;
                    sc_div_en        = 1'b0;
                   end
        "DDR1TO14":begin
                    sc_iserdes_mode  = 4'b0111;
                    sc_ddri_en       = 1'b1;
                    sc_des_ddren     = 1'b1;
                    sc_networking_en = 1'b1;
                    sc_div_en        = 1'b0;
                   end
// High-Speed Memory DDR
        "HMDDR1TO4": begin
                    sc_iserdes_mode  = 4'b0000;
                    sc_ddri_en       = 1'b1;
                    sc_des_ddren     = 1'b1;
                    sc_ihsmem_en     = 1'b1;
                    sc_ififo_en      = 1'b1;
                    sc_div_en        = 1'b1;
                   end
        "HMDDR1TO8": begin
                    sc_iserdes_mode  = 4'b0001;
                    sc_ddri_en       = 1'b1;
                    sc_des_ddren     = 1'b1;
                    sc_ihsmem_en     = 1'b1;
                    sc_ififo_en      = 1'b1;
                    sc_div_en        = 1'b1;
                   end
// Low-Speed Memory DDR
        "LMDDR1TO4": begin
                    sc_iserdes_mode  = 4'b0000;
                    sc_ddri_en       = 1'b1;
                    sc_des_ddren     = 1'b1;
                    sc_lsmem_en      = 1'b1;
                    sc_div_en        = 1'b0;
                   end
        "LMDDR1TO8": begin
                    sc_iserdes_mode  = 4'b0001;
                    sc_ddri_en       = 1'b1;
                    sc_des_ddren     = 1'b1;
                    sc_lsmem_en      = 1'b1;
                    sc_div_en        = 1'b0;
                   end
// OVERSAMPLE
        "OVERSAMPLE": begin
                    sc_ddri_en       = 1'b1;
                    sc_oversample_en = 1'b1;
                    sc_div_en        = 1'b0;
                   end
        default:   begin 
                    sc_iserdes_mode  = 4'b0000; 
                    sc_ddri_en       = 1'b0;
                    sc_des_sdren     = 1'b0;
                    sc_des_ddren     = 1'b0;
                    sc_networking_en = 1'b0;
                    sc_ihsmem_en     = 1'b0;
                    sc_ififo_en      = 1'b0;
                    sc_lsmem_en      = 1'b0;
                    sc_oversample_en = 1'b0;
                    sc_samepipeline_en = 1'b0;
                    sc_isame_en		 = 1'b0;
                    sc_iopposite_en	 = 1'b0;
                    sc_div_en        = 1'b0;
                    $display("Error: Illegal setting ISERDES_MODE of %s",ISERDES_MODE);
                    $finish; 
                   end
        endcase
end

initial begin
    case (GRS_TYPE_Q0)
        "SET"  :begin sc_init_q[0]=1'b1; end
        "RESET":begin sc_init_q[0]=1'b0; end
    endcase
end

initial begin
    case (GRS_TYPE_Q1)
        "SET"  :begin sc_init_q[1]=1'b1; end
        "RESET":begin sc_init_q[1]=1'b0; end
    endcase
end

initial begin
    case (GRS_TYPE_Q2)
        "SET"  :begin sc_init_q[2]=1'b1; end
        "RESET":begin sc_init_q[2]=1'b0; end
    endcase
end

initial begin
    case (GRS_TYPE_Q3)
        "SET"  :begin sc_init_q[3]=1'b1; end
        "RESET":begin sc_init_q[3]=1'b0; end
    endcase
end

initial begin
    case (LRS_TYPE_Q0)
        "ASYNC_SET"  :begin sc_isr_sync=1'b0; sc_srval_q[0]=1'b1; end
        "ASYNC_RESET":begin sc_isr_sync=1'b0; sc_srval_q[0]=1'b0; end
        "SYNC_SET"   :begin sc_isr_sync=1'b1; sc_srval_q[0]=1'b1; end
        "SYNC_RESET" :begin sc_isr_sync=1'b1; sc_srval_q[0]=1'b0; end
    endcase
end

initial begin
    case (LRS_TYPE_Q1)
        "ASYNC_SET"  :begin sc_isr_sync=1'b0; sc_srval_q[1]=1'b1; end
        "ASYNC_RESET":begin sc_isr_sync=1'b0; sc_srval_q[1]=1'b0; end
        "SYNC_SET"   :begin sc_isr_sync=1'b1; sc_srval_q[1]=1'b1; end
        "SYNC_RESET" :begin sc_isr_sync=1'b1; sc_srval_q[1]=1'b0; end
    endcase
end

initial begin
    case (LRS_TYPE_Q2)
        "ASYNC_SET"  :begin sc_isr_sync=1'b0; sc_srval_q[2]=1'b1; end
        "ASYNC_RESET":begin sc_isr_sync=1'b0; sc_srval_q[2]=1'b0; end
        "SYNC_SET"   :begin sc_isr_sync=1'b1; sc_srval_q[2]=1'b1; end
        "SYNC_RESET" :begin sc_isr_sync=1'b1; sc_srval_q[2]=1'b0; end
    endcase
end

initial begin
    case (LRS_TYPE_Q3)
        "ASYNC_SET"  :begin sc_isr_sync=1'b0; sc_srval_q[3]=1'b1; end
        "ASYNC_RESET":begin sc_isr_sync=1'b0; sc_srval_q[3]=1'b0; end
        "SYNC_SET"   :begin sc_isr_sync=1'b1; sc_srval_q[3]=1'b1; end
        "SYNC_RESET" :begin sc_isr_sync=1'b1; sc_srval_q[3]=1'b0; end
    endcase
end

always @ (posedge DESCLK or posedge RST) begin
    if(RST)
        desclk_reg <= 0;
    else
        desclk_reg <= ~desclk_reg;
end

iserdes_e2_iolhr_il_clkgen xiserdes_e2_iolhr_il_clkgen(
                             .desclk(desclk),
                             .iclk(iclk),
                             .iclkb(iclkb),
                             .oclk(oclk),
                             .oclkb(oclkb),
                             .iclkdiv(iclkdiv),
                             .bsclk(bsclk),
                             .dyn_clkpol(dyn_clkpol),
                             .dyn_clkdivpol(dyn_clkdivpol),
                             .sc_dyn_clkpol(sc_dyn_clkpol),
                             .sc_dyn_clkdivpol(sc_dyn_clkdivpol),
                             .sc_clk_pol0(sc_clk_pol0),
                             .sc_clk_pol1(sc_clk_pol1),
                             .sc_clk_pol2(sc_clk_pol2),
                             .sc_clk_pol3(sc_clk_pol3),
                             .sc_oclkpol(sc_oclkpol),
                             .sc_oclkbpol(sc_oclkbpol),
                             .sc_lsmem_en(sc_lsmem_en),
                             .sc_ihsmem_en(sc_ihsmem_en),
                             .sc_oversample_en(sc_oversample_en),
                             .clk_stg0(clk_stg0),
                             .clkb_stg0(clkb_stg0),
                             .hsmem_clk(hsmem_clk),
                             .hsmem_clkb(hsmem_clkb),
                             .clk_stg1_0(clk_stg1_0),
                             .clk_stg1_1(clk_stg1_1),
                             .clk_stg1_2(clk_stg1_2),
                             .clk_stg2_0(clk_stg2_0),
                             .clk_stg2_1(clk_stg2_1),
                             .clk_stg3(clk_stg3),
                             .clk_for_bs(clk_for_bs)                             
                            );

iserdes_e2_iolhr_il_srce xiserdes_e2_iolhr_il_srce(
                        .sc_isr_pol(sc_isr_pol),
                        .sc_isr_sync(sc_isr_sync),
                        .sc_isr_en(sc_isr_en),
                        .sc_grs_dis(sc_grs_dis),
                        .sc_ihsmem_en(sc_ihsmem_en),
                        .sc_ddri_en(sc_ddri_en),
                        .sc_num_ice(sc_num_ice),
                        .gwen(gwen),
                        .glogen(glogen),
                        .grs_n(grs_n),
                        .isr_iolhr(isr_iolhr),
                        .ice0(ice0),
                        .ice1(ice1),
                        .clk_stg3(clk_stg3),
                        .gsr(gsr),
                        .rstn(rstn_out),
                        .lsr_sync(lsr_sync),
                        .lsr_async(lsr_async),
                        .ce_hsmem(ce_hsmem),
                        .ce_out_0(ce_out_0),
                        .ce_out_1(ce_out_1)
                        );

iserdes_e2_iolhr_il_data xiserdes_e2_iolhr_il_data(
                         .sc_d_pol0(sc_d_pol0),
                         .sc_d_pol1(sc_d_pol1),
                         .sc_d_sel0(sc_d_sel0),
                         .sc_d_sel1(sc_d_sel1),
                         .sc_d_sel2(sc_d_sel2),
                         .sc_d_sel3(sc_d_sel3),
                         .sc_d_sel4(sc_d_sel4),
                         .sc_d_sel5(sc_d_sel5),
                         .sc_d_sel6(sc_d_sel6),
                         .sc_test_en0(sc_test_en0),
                         .sc_test_en1(sc_test_en1),
                         .sc_mipi_en(sc_mipi_en),
                         .glogen(glogen),
                         .di(di),
                         .di_n(di_n),
                         .di_mipi(di_mipi),
                         .di_from_srb(di_from_srb),
                         .ofb(ofb),
                         .tfb(tfb),
                         .zhold_dly(dly_zhold_in),
                         .d_dly(dly_idly_in),
                         .di_to_clk(),
                         .di_to_clkb(),
                         .di_to_fabric(),
                         .di_to_gear(di_to_gear),
                         .di_to_zhold(),
                         .di_to_idly()
                        );


iserdes_e2_iolhr_il_gearctrl iserdes_e2_iolhr_il_gearctrl(
                                 .clk_for_bs(clk_for_bs),
                                 .clkdiv_for_bs(clk_stg3),
                                 .gwen(gwen),
                                 .rstn(rstn_out),
                                 .sc_ddri_en(sc_ddri_en),
                                 .sc_des_ddren(sc_des_ddren),
                                 .sc_des_sdren(sc_des_sdren),
                                 .sc_iserdes_mode(sc_iserdes_mode),
                                 .sc_ihsmem_en(sc_ihsmem_en),
                                 .sc_lsmem_en(sc_lsmem_en),
                                 .sc_samepipeline_en(sc_samepipeline_en),
                                 .sc_isame_en(sc_isame_en),
                                 .sc_iopposite_en(sc_iopposite_en),
                                 .sc_ilthen(sc_ilthen),
                                 .sc_idffen(sc_idffen),
                                 .sc_oversample_en(sc_oversample_en),
                                 .sc_master(sc_master),
                                 .sc_networking_en(sc_networking_en),
                                 .sc_bitslip_en(sc_bitslip_en),
                                 .bitslip(bitslip),
                                 .bsclk(bsclk),
                                 .sel0(sel0),
                                 .sel1(sel1),
                                 .sel2(sel2),
                                 .sel3(sel3),
                                 .sel4(sel4),
                                 .sel5(sel5),
                                 .sel6(sel6),
                                 .sdr1to2(sdr1to2),
                                 .sdr1to3(sdr1to3),
                                 .sdr1to4(sdr1to4),
                                 .sdr1to5(sdr1to5),
                                 .sdr1to6(sdr1to6),
                                 .sdr1to7(sdr1to7),
                                 .sdr1to8(sdr1to8),
                                 .ddr1to4(ddr1to4),
                                 .ddr1to6(ddr1to6),
                                 .ddr1to8(ddr1to8),
                                 .ddr1to10(ddr1to10),
                                 .ddr1to14(ddr1to14)
                                );


iserdes_e2_iolhr_il_gear xiserdes_e2_iolhr_il_gear(
                         .di(di_to_gear),
                         .clk_stg0(clk_stg0),
                         .clkb_stg0(clkb_stg0),
                         .hsmem_clk(hsmem_clk),
                         .hsmem_clkb(hsmem_clkb),
                         .ce_out_0(ce_out_0),
                         .ce_out_1(ce_out_1),
                         .ce_hsmem(ce_hsmem),
                         .clk_stg1_0(clk_stg1_0),
                         .clk_stg1_1(clk_stg1_1),
                         .clk_stg1_2(clk_stg1_2),
                         .clk_stg2_0(clk_stg2_0),
                         .clk_stg2_1(clk_stg2_1),
                         .clk_stg3(clk_stg3),
                         .ishiftin0(ishiftin0),
                         .ishiftin1(ishiftin1),
                         .sc_master(sc_master),
                         .sc_ddri_en(sc_ddri_en),
                         .sc_ihsmem_en(sc_ihsmem_en),
                         .sc_oversample_en(sc_oversample_en),
                         .sc_des_sdren(sc_des_sdren),
                         .sc_ififo_en(sc_ififo_en),
                         .sc_ilthen(sc_ilthen),
                         .sc_grs_dis(sc_grs_dis),
                         .sc_init_q(sc_init_q),
                         .sc_srval_q(sc_srval_q),
                         .lsr_async(lsr_async),
                         .lsr_sync(lsr_sync),
                         .gwen(gwen),
                         .gsr(gsr),
                         .rstn(rstn_out),
                         .sdr1to2(sdr1to2),
                         .sdr1to3(sdr1to3),
                         .sdr1to4(sdr1to4),
                         .sdr1to5(sdr1to5),
                         .sdr1to6(sdr1to6),
                         .sdr1to7(sdr1to7),
                         .sdr1to8(sdr1to8),
                         .ddr1to4(ddr1to4),
                         .ddr1to6(ddr1to6),
                         .ddr1to8(ddr1to8),
                         .ddr1to10(ddr1to10),
                         .ddr1to14(ddr1to14),
                         .sel0(sel0),
                         .sel1(sel1),
                         .sel2(sel2),
                         .sel3(sel3),
                         .sel4(sel4),
                         .sel5(sel5),
                         .sel6(sel6),
                         .ififo_waddr(ififo_waddr),
                         .ififo_raddr(ififo_raddr),
                         .rx_data(rx_data),
                         .ishiftout0(ishiftout0),
                         .ishiftout1(ishiftout1)
                        );


endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
//  REVISION:
//  06/03/2019  mm/dd/yy - Initial version,                                                   
///////////////////////////////////////////////////////////////////////////////
`timescale 1ns/100fs 

module GTP_HSST_E1 
#(   
// PARAMETER  PART BEGINS ////////////////////////////////////////////////////////////////////
// PARAMETER  PART BEGINS ////////////////////////////////////////////////////////////////////
// PARAMETER  PART BEGINS ////////////////////////////////////////////////////////////////////


parameter           PCS_CH0_BYPASS_WORD_ALIGN   = "FALSE",      // FALSE,TRUE
parameter           PCS_CH0_BYPASS_DENC = "FALSE",     // FALSE,TRUE
parameter           PCS_CH0_BYPASS_BONDING  = "FALSE",      // FALSE,TRUE
parameter           PCS_CH0_BYPASS_CTC  = "FALSE",      // FALSE,TRUE
parameter           PCS_CH0_BYPASS_GEAR = "FALSE",      // FALSE,TRUE
parameter           PCS_CH0_BYPASS_BRIDGE   = "FALSE",      // FALSE,TRUE
parameter           PCS_CH0_DATA_MODE   = "X8",     // 8bit,10bit,16bit,20bit
parameter           PCS_CH0_RX_POLARITY_INV = "DELAY",      // 00: delay 01: bit polarity inversion 10: bit reversal 11: polarity inversion and bit reversal
parameter           PCS_CH0_ALIGN_MODE  = "1GB",        // 1GB,10GB,RAPIDIO,OUTSIDE
parameter           PCS_CH0_SAMP_16B = "X16",       // 16bit,20bit
parameter   integer PCS_CH0_COMMA_REG0 = 0,     // 
parameter   integer PCS_CH0_COMMA_MASK = 0,     // 
parameter           PCS_CH0_CEB_MODE = "10GB",     // 10GB,RAPIDIO,OUTSIDE
parameter           PCS_CH0_CTC_MODE = "1SKIP",     // 00: add or del 1 skip;01: add or del 2 skips;10: reserved ;11:4 skips
parameter   integer PCS_CH0_A_REG = 0,      // 
parameter           PCS_CH0_GE_AUTO_EN = "FALSE",        // CTC,FALSE,TRUE
parameter   integer PCS_CH0_SKIP_REG0 = 0,      // 
parameter   integer PCS_CH0_SKIP_REG1 = 0,      // 
parameter   integer PCS_CH0_SKIP_REG2 = 0,      // 
parameter   integer PCS_CH0_SKIP_REG3 = 0,      // 
parameter           PCS_CH0_DEC_DUAL = "FALSE",      // signal for 8b10b decoder module
parameter           PCS_CH0_SPLIT = "FALSE",        // signal for RX GEAR split, 1:split  0:no split; 
parameter           PCS_CH0_FIFOFLAG_CTC = "FALSE",     // FALSE,TRUE
parameter           PCS_CH0_COMMA_DET_MODE = "COMMA_PATTERN",       // 0: comma pattern mode  1: RX_CLK_SLIP mode 
parameter           PCS_CH0_ERRDETECT_SILENCE = "FALSE",        // 0: comma pattern mode  1: RX_CLK_SLIP mode 
parameter           PCS_CH0_PMA_RCLK_POLINV = "PMA_RCLK",       // 1'b0:pma_rclk 1'b1:reverse of pma_rclk
parameter           PCS_CH0_PCS_RCLK_SEL = "PMA_RCLK",      // 1'b0:pma_rclk;1'b1:pma_tclk;
parameter           PCS_CH0_MCB_RCLK_POLINV = "MCB_RCLK",       // 1'b0:mcb_rclk 1'b1:reverse of mcb_rclk
parameter           PCS_CH0_CB_RCLK_SEL = "PMA_RCLK",       // 2'b00:pma_rclk;2'b01:pma_tclk;2'b10:mcb_rclk;2'b11:reserved
parameter           PCS_CH0_AFTER_CTC_RCLK_SEL = "PMA_RCLK",        // 2'b00:pma_rclk;2'b01:pma_tclk;2'b10:mcb_rclk;2'b11:reserved
parameter           PCS_CH0_RCLK_POLINV = "RCLK",       // 1'b0:rclk 1'b1:reverse of rclk
parameter           PCS_CH0_BRIDGE_RCLK_SEL = "PMA_RCLK",       // 2'b00:pma_rclk;2'b01:pma_tclk;2'b10:mcb_rclk;2'b11:rclk
parameter           PCS_CH0_PCS_RCLK_EN = "FALSE",      // FALSE,TRUE
parameter           PCS_CH0_CB_RCLK_EN = "FALSE",       // FALSE,TRUE
parameter           PCS_CH0_AFTER_CTC_RCLK_EN = "FALSE",        // FALSE,TRUE
parameter           PCS_CH0_AFTER_CTC_RCLK_EN_GB = "FALSE",     // FALSE,TRUE
parameter           PCS_CH0_BRIDGE_RCLK_EN = "FALSE",       // FALSE,TRUE
parameter           PCS_CH0_PCS_RX_RSTN = "FALSE",      // 1:pcs_rx_rstn is valued,is 0;0:pcs_rx_rstn is released
parameter           PCS_CH0_SLAVE = "MASTER",       // 1:slave channel 0:master channel
parameter           PCS_CH0_PCIE_SLAVE = "MASTER",  // 1:slave channel 0:master channel
parameter           PCS_CH0_PCS_CB_RSTN = "FALSE",      // 1: pcs_cb_rstn is valued,is 0;0: pcs_cb_rstn is released
parameter           PCS_CH0_TX_BYPASS_BRIDGE_UINT   = "FALSE",      // FALSE,TRUE
parameter           PCS_CH0_TX_BYPASS_GEAR  = "FALSE",      // FALSE,TRUE
parameter           PCS_CH0_TX_BYPASS_ENC   = "FALSE",      // FALSE,TRUE
parameter           PCS_CH0_TX_BYPASS_BIT_SLIP  = "FALSE",      // FALSE,TRUE
parameter           PCS_CH0_TX_GEAR_SPLIT   = "FALSE",      // 1:spilt 44bits data to 22bits data,0: no spilt
parameter           PCS_CH0_TX_DRIVE_REG_MODE    = "NO_CHANGE",      // 00:no change, 01:enable polarity reverse,10:enable bit reverse, 11:enable both
parameter   integer PCS_CH0_TX_BIT_SLIP_CYCLES = 0,     // 
parameter           PCS_CH0_INT_TX_MASK_0 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by tx_bridge_unit async fifo overflow
parameter           PCS_CH0_INT_TX_MASK_1 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by tx bridge unit underflow;
parameter           PCS_CH0_INT_TX_MASK_2 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by tx_invalid_k 
parameter           PCS_CH0_INT_TX_CLR_0 = "FALSE",     // FALSE,TRUE  active high to clr int triggered by tx bridge unit overflow;
parameter           PCS_CH0_INT_TX_CLR_1 = "FALSE",     // FALSE,TRUE  active high to clr int triggered by tx_bridge_unit async fifo underflow
parameter           PCS_CH0_INT_TX_CLR_2 = "FALSE",     // FALSE,TRUE  active high to clr int triggered by tx_invalid_k
parameter           PCS_CH0_TX_PMA_TCLK_POLINV = "PMA_TCLK",        // 1'b0:pma_tclk 1'b1:reverse of pma_tclk
parameter           PCS_CH0_TX_PCS_CLK_EN_SEL = "FALSE",        // FALSE,TRUE
parameter           PCS_CH0_TX_BRIDGE_TCLK_SEL = "PCS_TCLK",        // 1'b0: pcs_tclk 1'b1:tclk
parameter           PCS_CH0_TX_TCLK_POLINV = "TCLK",        // 1'b0:tclk 1'b1:reverse of tclk
parameter           PCS_CH0_TX_PCS_TX_RSTN = "FALSE",      // 1:pcs_tx_rstn is valued,is 0;0:pcs_tx_rstn is released
parameter           PCS_CH0_TX_SLAVE = "SLAVE",     // 1:slave channel,0:master channel
parameter           PCS_CH0_TX_BRIDGE_CLK_EN_SEL = "FALSE",     // FALSE,TRUE
parameter           PCS_CH0_DATA_WIDTH_MODE = "X20",        // 20bit,16bit,10bit,8bit
parameter           PCS_CH0_TX_TCLK2FABRIC_SEL = "FALSE",       // FALSE,TRUE
parameter           PCS_CH0_TX_OUTZZ = "FALSE",    // 1:16bit/32bit only;0:other data width mode
parameter           PCS_CH0_ENC_DUAL = "FALSE",    // FALSE,TRUE
parameter           PCS_CH0_TX_BITSLIP_DATA_MODE = "X10",       // 1: 20bit,0: 10bit
parameter   integer PCS_CH0_COMMA_REG1 = 0,     // 
parameter   integer PCS_CH0_RAPID_IMAX = 0,     // 
parameter   integer PCS_CH0_RAPID_VMIN_1 = 0,       // 
parameter   integer PCS_CH0_RAPID_VMIN_2 = 0,       // 
parameter           PCS_CH0_RX_PRBS_MODE = "DISABLE",       // Mode select:4'd0: reserved,4'd1: PRBS-7,4'd2: PRBS-15,4'd3: PRBS-23,4'd4: PRBS-31,4'd5: long "1",4'd6: long "0",4'd7: 20UI square wave,4'd8: D10_2,4'd9: PCIe complianece pattern,Others: reserved
parameter           PCS_CH0_RX_ERRCNT_CLR = "FALSE",        // FALSE,TRUE
parameter           PCS_CH0_TX_PRBS_MODE = "DISABLE",       // Mode select:4'd0: reserved,4'd1: PRBS-7,4'd2: PRBS-15,4'd3: PRBS-23,4'd4: PRBS-31,4'd5: long "1",4'd6: long "0",4'd7: 20UI square wave,4'd8: D10_2,4'd9: PCIe complianece pattern,Others: reserved
parameter           PCS_CH0_TX_INSERT_ER = "FALSE",     // FALSE,TRUE
parameter           PCS_CH0_ENABLE_PRBS_GEN = "FALSE",      // FALSE,TRUE
parameter   integer PCS_CH0_ERR_CNT = 0,        // 
parameter   integer PCS_CH0_DEFAULT_RADDR = 0,      // 
parameter   integer PCS_CH0_MASTER_CHECK_OFFSET = 0,        // 
parameter   integer PCS_CH0_DELAY_SET = 0,      // 
parameter           PCS_CH0_SEACH_OFFSET = "20BIT",     // 20bit,30bit,40bit,50bit,60bit,70bit
parameter   integer PCS_CH0_CEB_RAPIDLS_MMAX = 0,       // 
parameter   integer PCS_CH0_CTC_AFULL = 0,      // 
parameter   integer PCS_CH0_CTC_AEMPTY = 0,     // 
parameter   integer PCS_CH0_CTC_CONTI_SKP_SET  = 0,     //2018/7/18  
parameter           PCS_CH0_FAR_LOOP = "FALSE",     // FALSE,TRUE
parameter           PCS_CH0_NEAR_LOOP = "FALSE",        // FALSE,TRUE
parameter           PCS_CH0_INT_RX_MASK_0 = "FALSE",       // FALSE,TRUE  active high to mask int triggered by pcs_lsm_synced
parameter           PCS_CH0_INT_RX_MASK_1 = "FALSE",       // FALSE,TRUE  active high to mask int triggered by pcs_rx_mcb_status
parameter           PCS_CH0_INT_RX_MASK_2 = "FALSE",       // FALSE,TRUE  active high to mask int triggered by channel bonding async fifo overflow
parameter           PCS_CH0_INT_RX_MASK_3 = "FALSE",       // FALSE,TRUE  active high to mask int triggered by channel bonding async fifo underflow
parameter           PCS_CH0_INT_RX_MASK_4 = "FALSE",       // FALSE,TRUE  active high to mask int triggered by ctc unit async fifo overflow
parameter           PCS_CH0_INT_RX_MASK_5 = "FALSE",       // FALSE,TRUE  active high to mask int triggered by ctc unit async fifo underflow
parameter           PCS_CH0_INT_RX_MASK_6 = "FALSE",       // FALSE,TRUE  active high to mask int triggered by rx_bridge_unit async fifo overflow
parameter           PCS_CH0_INT_RX_MASK_7 = "FALSE",       // FALSE,TRUE  active high to mask int triggered by rx_bridge_unit async fifo underflow
parameter           PCS_CH0_INT_RX_CLR_0 = "FALSE",    // FALSE,TRUE  active high to clr int triggered by pcs_lsm_synced
parameter           PCS_CH0_INT_RX_CLR_1 = "FALSE",    // FALSE,TRUE  active high to clr int triggered by pcs_rx_mcb_status
parameter           PCS_CH0_INT_RX_CLR_2 = "FALSE",    // FALSE,TRUE  active high to clr int triggered by channel bonding async fifo overflow
parameter           PCS_CH0_INT_RX_CLR_3 = "FALSE",    // FALSE,TRUE  active high to clr int triggered by channel bonding async fifo underflow
parameter           PCS_CH0_INT_RX_CLR_4 = "FALSE",    // FALSE,TRUE  active high to clr int triggered by ctc unit async fifo overflow
parameter           PCS_CH0_INT_RX_CLR_5 = "FALSE",    // FALSE,TRUE  active high to clr int triggered by ctc unit async fifo underflow
parameter           PCS_CH0_INT_RX_CLR_6 = "FALSE",    // FALSE,TRUE  active high to clr int triggered by rx_bridge_unit async fifo overflow
parameter           PCS_CH0_INT_RX_CLR_7 = "FALSE",    // FALSE,TRUE  active high to clr int triggered by rx_bridge_unit async fifo underflow
//add for clk aligner@2018/1/23
parameter integer   PCS_CH0_CA_RX  = 0,        // 
parameter integer   PCS_CH1_CA_RX  = 0,        // 
parameter integer   PCS_CH2_CA_RX  = 0,        // 
parameter integer   PCS_CH3_CA_RX  = 0,        // 
parameter integer   PCS_CH0_CA_TX  = 0,        // 
parameter integer   PCS_CH1_CA_TX  = 0,        // 
parameter integer   PCS_CH2_CA_TX  = 0,        // 
parameter integer   PCS_CH3_CA_TX  = 0,        // 
parameter           PCS_CH0_CA_DYN_DLY_EN_RX   = "FALSE",      // 
parameter           PCS_CH1_CA_DYN_DLY_EN_RX   = "FALSE",      // 
parameter           PCS_CH2_CA_DYN_DLY_EN_RX   = "FALSE",      // 
parameter           PCS_CH3_CA_DYN_DLY_EN_RX   = "FALSE",      // 
parameter           PCS_CH0_CA_DYN_DLY_EN_TX   = "FALSE",      // 
parameter           PCS_CH1_CA_DYN_DLY_EN_TX   = "FALSE",      // 
parameter           PCS_CH2_CA_DYN_DLY_EN_TX   = "FALSE",      // 
parameter           PCS_CH3_CA_DYN_DLY_EN_TX   = "FALSE",      // 
parameter           PCS_CH0_CA_DYN_DLY_SEL_RX  = "FALSE",      // 
parameter           PCS_CH1_CA_DYN_DLY_SEL_RX  = "FALSE",      // 
parameter           PCS_CH2_CA_DYN_DLY_SEL_RX  = "FALSE",      // 
parameter           PCS_CH3_CA_DYN_DLY_SEL_RX  = "FALSE",      // 
parameter           PCS_CH0_CA_DYN_DLY_SEL_TX  = "FALSE",      // 
parameter           PCS_CH1_CA_DYN_DLY_SEL_TX  = "FALSE",      // 
parameter           PCS_CH2_CA_DYN_DLY_SEL_TX  = "FALSE",      // 
parameter           PCS_CH3_CA_DYN_DLY_SEL_TX  = "FALSE",      // 
parameter           PCS_CH0_CA_RSTN_RX         = "FALSE",      // 
parameter           PCS_CH1_CA_RSTN_RX         = "FALSE",      // 
parameter           PCS_CH2_CA_RSTN_RX         = "FALSE",      // 
parameter           PCS_CH3_CA_RSTN_RX         = "FALSE",      // 
parameter           PCS_CH0_CA_RSTN_TX         = "FALSE",      // 
parameter           PCS_CH1_CA_RSTN_TX         = "FALSE",      // 
parameter           PCS_CH2_CA_RSTN_TX         = "FALSE",      // 
parameter           PCS_CH3_CA_RSTN_TX         = "FALSE",      // 
                    
parameter           PCS_CH1_BYPASS_WORD_ALIGN   = "FALSE",      // FALSE,TRUE
parameter           PCS_CH1_BYPASS_DENC = "FALSE",      // FALSE,TRUE
parameter           PCS_CH1_BYPASS_BONDING  = "FALSE",      // FALSE,TRUE
parameter           PCS_CH1_BYPASS_CTC  = "FALSE",     // FALSE,TRUE
parameter           PCS_CH1_BYPASS_GEAR = "FALSE",     // FALSE,TRUE
parameter           PCS_CH1_BYPASS_BRIDGE   = "FALSE",      // FALSE,TRUE
parameter           PCS_CH1_DATA_MODE   = "X8",     // 8bit,10bit,16bit,20bit
parameter           PCS_CH1_RX_POLARITY_INV = "DELAY",      // 00: delay 01: bit polarity inversion 10: bit reversal 11: polarity inversion and bit reversal
parameter           PCS_CH1_ALIGN_MODE  = "1GB",        // 1GB,10GB,RAPIDIO,OUTSIDE
parameter           PCS_CH1_SAMP_16B = "X16",       // 16bit,20bit
parameter   integer PCS_CH1_COMMA_REG0 = 0,     // 
parameter   integer PCS_CH1_COMMA_MASK = 0,     // 
parameter           PCS_CH1_CEB_MODE = "10GB",      // 10GB,RAPIDIO,OUTSIDE
parameter           PCS_CH1_CTC_MODE = "1SKIP",     // 00: add or del 1 skip;01: add or del 2 skips;10: reserved ;11:4 skips
parameter   integer PCS_CH1_A_REG = 0,      // 
parameter           PCS_CH1_GE_AUTO_EN = "FALSE",       // CTC,FALSE,TRUE
parameter   integer PCS_CH1_SKIP_REG0 = 0,      // 
parameter   integer PCS_CH1_SKIP_REG1 = 0,      // 
parameter   integer PCS_CH1_SKIP_REG2 = 0,      // 
parameter   integer PCS_CH1_SKIP_REG3 = 0,      // 
parameter           PCS_CH1_DEC_DUAL = "FALSE",     // signal for 8b10b decoder module
parameter           PCS_CH1_SPLIT = "FALSE",       // signal for RX GEAR split, 1:split  0:no split; 
parameter           PCS_CH1_FIFOFLAG_CTC = "FALSE",     // FALSE,TRUE
parameter           PCS_CH1_COMMA_DET_MODE = "COMMA_PATTERN",       // 0: comma pattern mode  1: RX_CLK_SLIP mode 
parameter           PCS_CH1_ERRDETECT_SILENCE = "FALSE",        // 0: comma pattern mode  1: RX_CLK_SLIP mode 
parameter           PCS_CH1_PMA_RCLK_POLINV = "PMA_RCLK",      // 1'b0:pma_rclk 1'b1:reverse of pma_rclk
parameter           PCS_CH1_PCS_RCLK_SEL = "PMA_RCLK",      // 1'b0:pma_rclk;1'b1:pma_tclk;
parameter           PCS_CH1_MCB_RCLK_POLINV = "MCB_RCLK",       // 1'b0:mcb_rclk 1'b1:reverse of mcb_rclk
parameter           PCS_CH1_CB_RCLK_SEL = "PMA_RCLK",       // 2'b00:pma_rclk;2'b01:pma_tclk;2'b10:mcb_rclk;2'b11:reserved
parameter           PCS_CH1_AFTER_CTC_RCLK_SEL = "PMA_RCLK",        // 2'b00:pma_rclk;2'b01:pma_tclk;2'b10:mcb_rclk;2'b11:reserved
parameter           PCS_CH1_RCLK_POLINV = "RCLK",       // 1'b0:rclk 1'b1:reverse of rclk
parameter           PCS_CH1_BRIDGE_RCLK_SEL = "PMA_RCLK",       // 2'b00:pma_rclk;2'b01:pma_tclk;2'b10:mcb_rclk;2'b11:rclk
parameter           PCS_CH1_PCS_RCLK_EN = "FALSE",      // FALSE,TRUE
parameter           PCS_CH1_CB_RCLK_EN = "FALSE",       // FALSE,TRUE
parameter           PCS_CH1_AFTER_CTC_RCLK_EN = "FALSE",        // FALSE,TRUE
parameter           PCS_CH1_AFTER_CTC_RCLK_EN_GB = "FALSE",     // FALSE,TRUE
parameter           PCS_CH1_BRIDGE_RCLK_EN = "FALSE",       // FALSE,TRUE
parameter           PCS_CH1_PCS_RX_RSTN = "FALSE",      // 1:pcs_rx_rstn is valued,is 0;0:pcs_rx_rstn is released
parameter           PCS_CH1_SLAVE = "MASTER",       // 1:slave channel 0:master channel
parameter           PCS_CH1_PCIE_SLAVE = "MASTER",  // 1:slave channel 0:master channel
parameter           PCS_CH1_PCS_CB_RSTN = "FALSE",      // 1: pcs_cb_rstn is valued,is 0;0: pcs_cb_rstn is released
parameter           PCS_CH1_TX_BYPASS_BRIDGE_UINT   = "FALSE",      // FALSE,TRUE
parameter           PCS_CH1_TX_BYPASS_GEAR  = "FALSE",      // FALSE,TRUE
parameter           PCS_CH1_TX_BYPASS_ENC   = "FALSE",      // FALSE,TRUE
parameter           PCS_CH1_TX_BYPASS_BIT_SLIP  = "FALSE",      // FALSE,TRUE
parameter           PCS_CH1_TX_GEAR_SPLIT   = "FALSE",      // 1:spilt 44bits data to 22bits data,0: no spilt
parameter           PCS_CH1_TX_DRIVE_REG_MODE   = "NO_CHANGE",      // 00:no change, 01:enable polarity reverse,10:enable bit reverse, 11:enable both
parameter   integer PCS_CH1_TX_BIT_SLIP_CYCLES = 0,     // 
parameter           PCS_CH1_INT_TX_MASK_0 = "FALSE",       // FALSE,TRUE  active high to mask int triggered by tx_bridge_unit async fifo overflow
parameter           PCS_CH1_INT_TX_MASK_1 = "FALSE",       // FALSE,TRUE  active high to mask int triggered by tx bridge unit underflow;
parameter           PCS_CH1_INT_TX_MASK_2 = "FALSE",       // FALSE,TRUE  active high to mask int triggered by tx_invalid_k 
parameter           PCS_CH1_INT_TX_CLR_0 = "FALSE",     // FALSE,TRUE  active high to clr int triggered by tx bridge unit overflow;
parameter           PCS_CH1_INT_TX_CLR_1 = "FALSE",     // FALSE,TRUE  active high to clr int triggered by tx_bridge_unit async fifo underflow
parameter           PCS_CH1_INT_TX_CLR_2 = "FALSE",     // FALSE,TRUE  active high to clr int triggered by tx_invalid_k
parameter           PCS_CH1_TX_PMA_TCLK_POLINV = "PMA_TCLK",        // 1'b0:pma_tclk 1'b1:reverse of pma_tclk
parameter           PCS_CH1_TX_PCS_CLK_EN_SEL = "FALSE",        // FALSE,TRUE
parameter           PCS_CH1_TX_BRIDGE_TCLK_SEL = "PCS_TCLK",        // 1'b0: pcs_tclk 1'b1:tclk
parameter           PCS_CH1_TX_TCLK_POLINV = "TCLK",        // 1'b0:tclk 1'b1:reverse of tclk
parameter           PCS_CH1_TX_PCS_TX_RSTN = "FALSE",       // 1:pcs_tx_rstn is valued,is 0;0:pcs_tx_rstn is released
parameter           PCS_CH1_TX_SLAVE = "SLAVE",     // 1:slave channel,0:master channel
parameter           PCS_CH1_TX_BRIDGE_CLK_EN_SEL = "FALSE",     // FALSE,TRUE
parameter           PCS_CH1_DATA_WIDTH_MODE = "X20",        // 20bit,16bit,10bit,8bit
parameter           PCS_CH1_TX_TCLK2FABRIC_SEL = "FALSE",       // FALSE,TRUE
parameter           PCS_CH1_TX_OUTZZ = "FALSE",     // 1:16bit/32bit only;0:other data width mode
parameter           PCS_CH1_ENC_DUAL = "FALSE",     // FALSE,TRUE
parameter           PCS_CH1_TX_BITSLIP_DATA_MODE = "X10",       // 1: 20bit,0: 10bit
parameter   integer PCS_CH1_COMMA_REG1 = 0,     // 
parameter   integer PCS_CH1_RAPID_IMAX = 0,     // 
parameter   integer PCS_CH1_RAPID_VMIN_1 = 0,       // 
parameter   integer PCS_CH1_RAPID_VMIN_2 = 0,       // 
parameter           PCS_CH1_RX_PRBS_MODE = "DISABLE",       // Mode select:4'd0: reserved,4'd1: PRBS-7,4'd2: PRBS-15,4'd3: PRBS-23,4'd4: PRBS-31,4'd5: long "1",4'd6: long "0",4'd7: 20UI square wave,4'd8: D10_2,4'd9: PCIe complianece pattern,Others: reserved
parameter           PCS_CH1_RX_ERRCNT_CLR = "FALSE",        // FALSE,TRUE
parameter           PCS_CH1_TX_PRBS_MODE = "DISABLE",       // Mode select:4'd0: reserved,4'd1: PRBS-7,4'd2: PRBS-15,4'd3: PRBS-23,4'd4: PRBS-31,4'd5: long "1",4'd6: long "0",4'd7: 20UI square wave,4'd8: D10_2,4'd9: PCIe complianece pattern,Others: reserved
parameter           PCS_CH1_TX_INSERT_ER = "FALSE",     // FALSE,TRUE
parameter           PCS_CH1_ENABLE_PRBS_GEN = "FALSE",      // FALSE,TRUE
parameter   integer PCS_CH1_ERR_CNT = 0,        // 
parameter   integer PCS_CH1_DEFAULT_RADDR = 0,      // 
parameter   integer PCS_CH1_MASTER_CHECK_OFFSET = 0,        // 
parameter   integer PCS_CH1_DELAY_SET = 0,      // 
parameter           PCS_CH1_SEACH_OFFSET = "20BIT",     // 20bit,30bit,40bit,50bit,60bit,70bit
parameter   integer PCS_CH1_CEB_RAPIDLS_MMAX = 0,       // 
parameter   integer PCS_CH1_CTC_AFULL = 0,      // 
parameter   integer PCS_CH1_CTC_AEMPTY = 0,     // 
parameter   integer PCS_CH1_CTC_CONTI_SKP_SET  = 0,     //2018/7/18  
parameter           PCS_CH1_FAR_LOOP = "FALSE",     // FALSE,TRUE
parameter           PCS_CH1_NEAR_LOOP = "FALSE",        // FALSE,TRUE
parameter           PCS_CH1_INT_RX_MASK_0 = "FALSE",       // FALSE,TRUE  active high to mask int triggered by pcs_lsm_synced
parameter           PCS_CH1_INT_RX_MASK_1 = "FALSE",       // FALSE,TRUE  active high to mask int triggered by pcs_rx_mcb_status
parameter           PCS_CH1_INT_RX_MASK_2 = "FALSE",       // FALSE,TRUE  active high to mask int triggered by channel bonding async fifo overflow
parameter           PCS_CH1_INT_RX_MASK_3 = "FALSE",       // FALSE,TRUE  active high to mask int triggered by channel bonding async fifo underflow
parameter           PCS_CH1_INT_RX_MASK_4 = "FALSE",       // FALSE,TRUE  active high to mask int triggered by ctc unit async fifo overflow
parameter           PCS_CH1_INT_RX_MASK_5 = "FALSE",       // FALSE,TRUE  active high to mask int triggered by ctc unit async fifo underflow
parameter           PCS_CH1_INT_RX_MASK_6 = "FALSE",       // FALSE,TRUE  active high to mask int triggered by rx_bridge_unit async fifo overflow
parameter           PCS_CH1_INT_RX_MASK_7 = "FALSE",       // FALSE,TRUE  active high to mask int triggered by rx_bridge_unit async fifo underflow
parameter           PCS_CH1_INT_RX_CLR_0 = "FALSE",     // FALSE,TRUE  active high to clr int triggered by pcs_lsm_synced
parameter           PCS_CH1_INT_RX_CLR_1 = "FALSE",     // FALSE,TRUE  active high to clr int triggered by pcs_rx_mcb_status
parameter           PCS_CH1_INT_RX_CLR_2 = "FALSE",     // FALSE,TRUE  active high to clr int triggered by channel bonding async fifo overflow
parameter           PCS_CH1_INT_RX_CLR_3 = "FALSE",     // FALSE,TRUE  active high to clr int triggered by channel bonding async fifo underflow
parameter           PCS_CH1_INT_RX_CLR_4 = "FALSE",     // FALSE,TRUE  active high to clr int triggered by ctc unit async fifo overflow
parameter           PCS_CH1_INT_RX_CLR_5 = "FALSE",     // FALSE,TRUE  active high to clr int triggered by ctc unit async fifo underflow
parameter           PCS_CH1_INT_RX_CLR_6 = "FALSE",     // FALSE,TRUE  active high to clr int triggered by rx_bridge_unit async fifo overflow
parameter           PCS_CH1_INT_RX_CLR_7 = "FALSE",     // FALSE,TRUE  active high to clr int triggered by rx_bridge_unit async fifo underflow
                    
                    
                    
parameter           PCS_CH2_BYPASS_WORD_ALIGN   = "FALSE",      // FALSE,TRUE
parameter           PCS_CH2_BYPASS_DENC = "FALSE",      // FALSE,TRUE
parameter           PCS_CH2_BYPASS_BONDING  = "FALSE",      // FALSE,TRUE
parameter           PCS_CH2_BYPASS_CTC  = "FALSE",      // FALSE,TRUE
parameter           PCS_CH2_BYPASS_GEAR = "FALSE",      // FALSE,TRUE
parameter           PCS_CH2_BYPASS_BRIDGE   = "FALSE",      // FALSE,TRUE
parameter           PCS_CH2_DATA_MODE   = "X8",     // 8bit,10bit,16bit,20bit
parameter           PCS_CH2_RX_POLARITY_INV = "DELAY",      // 00: delay 01: bit polarity inversion 10: bit reversal 11: polarity inversion and bit reversal
parameter           PCS_CH2_ALIGN_MODE  = "1GB",        // 1GB,10GB,RAPIDIO,OUTSIDE
parameter           PCS_CH2_SAMP_16B = "X16",       // 16bit,20bit
parameter   integer PCS_CH2_COMMA_REG0 = 0,     // 
parameter   integer PCS_CH2_COMMA_MASK = 0,     // 
parameter           PCS_CH2_CEB_MODE = "10GB",      // 10GB,RAPIDIO,OUTSIDE
parameter           PCS_CH2_CTC_MODE = "1SKIP",     // 00: add or del 1 skip;01: add or del 2 skips;10: reserved ;11:4 skips
parameter   integer PCS_CH2_A_REG = 0,      // 
parameter           PCS_CH2_GE_AUTO_EN = "FALSE",       // CTC,FALSE,TRUE
parameter   integer PCS_CH2_SKIP_REG0 = 0,      // 
parameter   integer PCS_CH2_SKIP_REG1 = 0,      // 
parameter   integer PCS_CH2_SKIP_REG2 = 0,      // 
parameter   integer PCS_CH2_SKIP_REG3 = 0,      // 
parameter           PCS_CH2_DEC_DUAL = "FALSE",     // signal for 8b10b decoder module
parameter           PCS_CH2_SPLIT = "FALSE",        // signal for RX GEAR split, 1:split  0:no split; 
parameter           PCS_CH2_FIFOFLAG_CTC = "FALSE",     // FALSE,TRUE
parameter           PCS_CH2_COMMA_DET_MODE = "COMMA_PATTERN",       // 0: comma pattern mode  1: RX_CLK_SLIP mode 
parameter           PCS_CH2_ERRDETECT_SILENCE = "FALSE",        // 0: comma pattern mode  1: RX_CLK_SLIP mode 
parameter           PCS_CH2_PMA_RCLK_POLINV = "PMA_RCLK",       // 1'b0:pma_rclk 1'b1:reverse of pma_rclk
parameter           PCS_CH2_PCS_RCLK_SEL = "PMA_RCLK",      // 1'b0:pma_rclk;1'b1:pma_tclk;
parameter           PCS_CH2_MCB_RCLK_POLINV = "MCB_RCLK",       // 1'b0:mcb_rclk 1'b1:reverse of mcb_rclk
parameter           PCS_CH2_CB_RCLK_SEL = "PMA_RCLK",       // 2'b00:pma_rclk;2'b01:pma_tclk;2'b10:mcb_rclk;2'b11:reserved
parameter           PCS_CH2_AFTER_CTC_RCLK_SEL = "PMA_RCLK",        // 2'b00:pma_rclk;2'b01:pma_tclk;2'b10:mcb_rclk;2'b11:reserved
parameter           PCS_CH2_RCLK_POLINV = "RCLK",       // 1'b0:rclk 1'b1:reverse of rclk
parameter           PCS_CH2_BRIDGE_RCLK_SEL = "PMA_RCLK",       // 2'b00:pma_rclk;2'b01:pma_tclk;2'b10:mcb_rclk;2'b11:rclk
parameter           PCS_CH2_PCS_RCLK_EN = "FALSE",      // FALSE,TRUE
parameter           PCS_CH2_CB_RCLK_EN = "FALSE",      // FALSE,TRUE
parameter           PCS_CH2_AFTER_CTC_RCLK_EN = "FALSE",        // FALSE,TRUE
parameter           PCS_CH2_AFTER_CTC_RCLK_EN_GB = "FALSE",     // FALSE,TRUE
parameter           PCS_CH2_BRIDGE_RCLK_EN = "FALSE",       // FALSE,TRUE
parameter           PCS_CH2_PCS_RX_RSTN = "FALSE",      // 1:pcs_rx_rstn is valued,is 0;0:pcs_rx_rstn is released
parameter           PCS_CH2_SLAVE = "MASTER",       // 1:slave channel 0:master channel
parameter           PCS_CH2_PCIE_SLAVE = "MASTER", // 1:slave channel 0:master channel
parameter           PCS_CH2_PCS_CB_RSTN = "FALSE",     // 1: pcs_cb_rstn is valued,is 0;0: pcs_cb_rstn is released
parameter           PCS_CH2_TX_BYPASS_BRIDGE_UINT   = "FALSE",      // FALSE,TRUE
parameter           PCS_CH2_TX_BYPASS_GEAR  = "FALSE",      // FALSE,TRUE
parameter           PCS_CH2_TX_BYPASS_ENC   = "FALSE",      // FALSE,TRUE
parameter           PCS_CH2_TX_BYPASS_BIT_SLIP  = "FALSE",      // FALSE,TRUE
parameter           PCS_CH2_TX_GEAR_SPLIT   = "FALSE",      // 1:spilt 44bits data to 22bits data,0: no spilt
parameter           PCS_CH2_TX_DRIVE_REG_MODE   = "NO_CHANGE",      // 00:no change, 01:enable polarity reverse,10:enable bit reverse, 11:enable both
parameter   integer PCS_CH2_TX_BIT_SLIP_CYCLES = 0,     // 
parameter           PCS_CH2_INT_TX_MASK_0 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by tx_bridge_unit async fifo overflow
parameter           PCS_CH2_INT_TX_MASK_1 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by tx bridge unit underflow;
parameter           PCS_CH2_INT_TX_MASK_2 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by tx_invalid_k 
parameter           PCS_CH2_INT_TX_CLR_0 = "FALSE",     // FALSE,TRUE  active high to clr int triggered by tx bridge unit overflow;
parameter           PCS_CH2_INT_TX_CLR_1 = "FALSE",     // FALSE,TRUE  active high to clr int triggered by tx_bridge_unit async fifo underflow
parameter           PCS_CH2_INT_TX_CLR_2 = "FALSE",     // FALSE,TRUE  active high to clr int triggered by tx_invalid_k
parameter           PCS_CH2_TX_PMA_TCLK_POLINV = "PMA_TCLK",        // 1'b0:pma_tclk 1'b1:reverse of pma_tclk
parameter           PCS_CH2_TX_PCS_CLK_EN_SEL = "FALSE",        // FALSE,TRUE
parameter           PCS_CH2_TX_BRIDGE_TCLK_SEL = "PCS_TCLK",        // 1'b0: pcs_tclk 1'b1:tclk
parameter           PCS_CH2_TX_TCLK_POLINV = "TCLK",        // 1'b0:tclk 1'b1:reverse of tclk
parameter           PCS_CH2_TX_PCS_TX_RSTN = "FALSE",       // 1:pcs_tx_rstn is valued,is 0;0:pcs_tx_rstn is released
parameter           PCS_CH2_TX_SLAVE = "SLAVE",     // 1:slave channel,0:master channel
parameter           PCS_CH2_TX_BRIDGE_CLK_EN_SEL = "FALSE",     // FALSE,TRUE
parameter           PCS_CH2_DATA_WIDTH_MODE = "X20",        // 20bit,16bit,10bit,8bit
parameter           PCS_CH2_TX_TCLK2FABRIC_SEL = "FALSE",       // FALSE,TRUE
parameter           PCS_CH2_TX_OUTZZ = "FALSE",     // 1:16bit/32bit only;0:other data width mode
parameter           PCS_CH2_ENC_DUAL = "FALSE",     // FALSE,TRUE
parameter           PCS_CH2_TX_BITSLIP_DATA_MODE = "X10",       // 1: 20bit,0: 10bit
parameter   integer PCS_CH2_COMMA_REG1 = 0,     // 
parameter   integer PCS_CH2_RAPID_IMAX = 0,     // 
parameter   integer PCS_CH2_RAPID_VMIN_1 = 0,       // 
parameter   integer PCS_CH2_RAPID_VMIN_2 = 0,       // 
parameter           PCS_CH2_RX_PRBS_MODE = "DISABLE",       // Mode select:4'd0: reserved,4'd1: PRBS-7,4'd2: PRBS-15,4'd3: PRBS-23,4'd4: PRBS-31,4'd5: long "1",4'd6: long "0",4'd7: 20UI square wave,4'd8: D10_2,4'd9: PCIe complianece pattern,Others: reserved
parameter           PCS_CH2_RX_ERRCNT_CLR = "FALSE",        // FALSE,TRUE
parameter           PCS_CH2_TX_PRBS_MODE = "DISABLE",       // Mode select:4'd0: reserved,4'd1: PRBS-7,4'd2: PRBS-15,4'd3: PRBS-23,4'd4: PRBS-31,4'd5: long "1",4'd6: long "0",4'd7: 20UI square wave,4'd8: D10_2,4'd9: PCIe complianece pattern,Others: reserved
parameter           PCS_CH2_TX_INSERT_ER = "FALSE",     // FALSE,TRUE
parameter           PCS_CH2_ENABLE_PRBS_GEN = "FALSE",      // FALSE,TRUE
parameter   integer PCS_CH2_ERR_CNT = 0,        // 
parameter   integer PCS_CH2_DEFAULT_RADDR = 0,      // 
parameter   integer PCS_CH2_MASTER_CHECK_OFFSET = 0,        // 
parameter   integer PCS_CH2_DELAY_SET = 0,      // 
parameter           PCS_CH2_SEACH_OFFSET = "20BIT",     // 20bit,30bit,40bit,50bit,60bit,70bit
parameter   integer PCS_CH2_CEB_RAPIDLS_MMAX = 0,       // 
parameter   integer PCS_CH2_CTC_AFULL = 0,      // 
parameter   integer PCS_CH2_CTC_AEMPTY = 0,     // 
parameter   integer PCS_CH2_CTC_CONTI_SKP_SET  = 0,     //2018/7/18  
parameter           PCS_CH2_FAR_LOOP = "FALSE",     // FALSE,TRUE
parameter           PCS_CH2_NEAR_LOOP = "FALSE",        // FALSE,TRUE
parameter           PCS_CH2_INT_RX_MASK_0 = "FALSE",       // FALSE,TRUE  active high to mask int triggered by pcs_lsm_synced
parameter           PCS_CH2_INT_RX_MASK_1 = "FALSE",       // FALSE,TRUE  active high to mask int triggered by pcs_rx_mcb_status
parameter           PCS_CH2_INT_RX_MASK_2 = "FALSE",       // FALSE,TRUE  active high to mask int triggered by channel bonding async fifo overflow
parameter           PCS_CH2_INT_RX_MASK_3 = "FALSE",       // FALSE,TRUE  active high to mask int triggered by channel bonding async fifo underflow
parameter           PCS_CH2_INT_RX_MASK_4 = "FALSE",       // FALSE,TRUE  active high to mask int triggered by ctc unit async fifo overflow
parameter           PCS_CH2_INT_RX_MASK_5 = "FALSE",       // FALSE,TRUE  active high to mask int triggered by ctc unit async fifo underflow
parameter           PCS_CH2_INT_RX_MASK_6 = "FALSE",       // FALSE,TRUE  active high to mask int triggered by rx_bridge_unit async fifo overflow
parameter           PCS_CH2_INT_RX_MASK_7 = "FALSE",       // FALSE,TRUE  active high to mask int triggered by rx_bridge_unit async fifo underflow
parameter           PCS_CH2_INT_RX_CLR_0 = "FALSE",     // FALSE,TRUE  active high to clr int triggered by pcs_lsm_synced
parameter           PCS_CH2_INT_RX_CLR_1 = "FALSE",     // FALSE,TRUE  active high to clr int triggered by pcs_rx_mcb_status
parameter           PCS_CH2_INT_RX_CLR_2 = "FALSE",     // FALSE,TRUE  active high to clr int triggered by channel bonding async fifo overflow
parameter           PCS_CH2_INT_RX_CLR_3 = "FALSE",     // FALSE,TRUE  active high to clr int triggered by channel bonding async fifo underflow
parameter           PCS_CH2_INT_RX_CLR_4 = "FALSE",     // FALSE,TRUE  active high to clr int triggered by ctc unit async fifo overflow
parameter           PCS_CH2_INT_RX_CLR_5 = "FALSE",     // FALSE,TRUE  active high to clr int triggered by ctc unit async fifo underflow
parameter           PCS_CH2_INT_RX_CLR_6 = "FALSE",     // FALSE,TRUE  active high to clr int triggered by rx_bridge_unit async fifo overflow
parameter           PCS_CH2_INT_RX_CLR_7 = "FALSE",     // FALSE,TRUE  active high to clr int triggered by rx_bridge_unit async fifo underflow
                    
                    
                    
parameter           PCS_CH3_BYPASS_WORD_ALIGN   = "FALSE",      // FALSE,TRUE
parameter           PCS_CH3_BYPASS_DENC = "FALSE",      // FALSE,TRUE
parameter           PCS_CH3_BYPASS_BONDING  = "FALSE",      // FALSE,TRUE
parameter           PCS_CH3_BYPASS_CTC  = "FALSE",      // FALSE,TRUE
parameter           PCS_CH3_BYPASS_GEAR = "FALSE",      // FALSE,TRUE
parameter           PCS_CH3_BYPASS_BRIDGE   = "FALSE",      // FALSE,TRUE
parameter           PCS_CH3_DATA_MODE   = "X8",     // 8bit,10bit,16bit,20bit
parameter           PCS_CH3_RX_POLARITY_INV = "DELAY",      // 00: delay 01: bit polarity inversion 10: bit reversal 11: polarity inversion and bit reversal
parameter           PCS_CH3_ALIGN_MODE  = "1GB",        // 1GB,10GB,RAPIDIO,OUTSIDE
parameter           PCS_CH3_SAMP_16B = "X16",       // 16bit,20bit
parameter   integer PCS_CH3_COMMA_REG0 = 0,     // 
parameter   integer PCS_CH3_COMMA_MASK = 0,     // 
parameter           PCS_CH3_CEB_MODE = "10GB",      // 10GB,RAPIDIO,OUTSIDE
parameter           PCS_CH3_CTC_MODE = "1SKIP",     // 00: add or del 1 skip;01: add or del 2 skips;10: reserved ;11:4 skips
parameter   integer PCS_CH3_A_REG = 0,      // 
parameter           PCS_CH3_GE_AUTO_EN = "FALSE",       // CTC,FALSE,TRUE
parameter   integer PCS_CH3_SKIP_REG0 = 0,      // 
parameter   integer PCS_CH3_SKIP_REG1 = 0,      // 
parameter   integer PCS_CH3_SKIP_REG2 = 0,      // 
parameter   integer PCS_CH3_SKIP_REG3 = 0,      // 
parameter           PCS_CH3_DEC_DUAL = "FALSE",     // signal for 8b10b decoder module
parameter           PCS_CH3_SPLIT = "FALSE",        // signal for RX GEAR split, 1:split  0:no split; 
parameter           PCS_CH3_FIFOFLAG_CTC = "FALSE",     // FALSE,TRUE
parameter           PCS_CH3_COMMA_DET_MODE = "COMMA_PATTERN",       // 0: comma pattern mode  1: RX_CLK_SLIP mode 
parameter           PCS_CH3_ERRDETECT_SILENCE = "FALSE",        // 0: comma pattern mode  1: RX_CLK_SLIP mode 
parameter           PCS_CH3_PMA_RCLK_POLINV = "PMA_RCLK",       // 1'b0:pma_rclk 1'b1:reverse of pma_rclk
parameter           PCS_CH3_PCS_RCLK_SEL = "PMA_RCLK",      // 1'b0:pma_rclk;1'b1:pma_tclk;
parameter           PCS_CH3_MCB_RCLK_POLINV = "MCB_RCLK",       // 1'b0:mcb_rclk 1'b1:reverse of mcb_rclk
parameter           PCS_CH3_CB_RCLK_SEL = "PMA_RCLK",       // 2'b00:pma_rclk;2'b01:pma_tclk;2'b10:mcb_rclk;2'b11:reserved
parameter           PCS_CH3_AFTER_CTC_RCLK_SEL = "PMA_RCLK",        // 2'b00:pma_rclk;2'b01:pma_tclk;2'b10:mcb_rclk;2'b11:reserved
parameter           PCS_CH3_RCLK_POLINV = "RCLK",       // 1'b0:rclk 1'b1:reverse of rclk
parameter           PCS_CH3_BRIDGE_RCLK_SEL = "PMA_RCLK",       // 2'b00:pma_rclk;2'b01:pma_tclk;2'b10:mcb_rclk;2'b11:rclk
parameter           PCS_CH3_PCS_RCLK_EN = "FALSE",      // FALSE,TRUE
parameter           PCS_CH3_CB_RCLK_EN = "FALSE",       // FALSE,TRUE
parameter           PCS_CH3_AFTER_CTC_RCLK_EN = "FALSE",        // FALSE,TRUE
parameter           PCS_CH3_AFTER_CTC_RCLK_EN_GB = "FALSE",     // FALSE,TRUE
parameter           PCS_CH3_BRIDGE_RCLK_EN = "FALSE",       // FALSE,TRUE
parameter           PCS_CH3_PCS_RX_RSTN = "FALSE",      // 1:pcs_rx_rstn is valued,is 0;0:pcs_rx_rstn is released
parameter           PCS_CH3_SLAVE = "MASTER",       // 1:slave channel 0:master channel
parameter           PCS_CH3_PCIE_SLAVE = "MASTER",  // 1:slave channel 0:master channel
parameter           PCS_CH3_PCS_CB_RSTN = "FALSE",      // 1: pcs_cb_rstn is valued,is 0;0: pcs_cb_rstn is released
parameter           PCS_CH3_TX_BYPASS_BRIDGE_UINT   = "FALSE",      // FALSE,TRUE
parameter           PCS_CH3_TX_BYPASS_GEAR  = "FALSE",      // FALSE,TRUE
parameter           PCS_CH3_TX_BYPASS_ENC   = "FALSE",      // FALSE,TRUE
parameter           PCS_CH3_TX_BYPASS_BIT_SLIP  = "FALSE",      // FALSE,TRUE
parameter           PCS_CH3_TX_GEAR_SPLIT   = "FALSE",      // 1:spilt 44bits data to 22bits data,0: no spilt
parameter           PCS_CH3_TX_DRIVE_REG_MODE   = "NO_CHANGE",      // 00:no change, 01:enable polarity reverse,10:enable bit reverse, 11:enable both
parameter   integer PCS_CH3_TX_BIT_SLIP_CYCLES = 0,     // 
parameter           PCS_CH3_INT_TX_MASK_0 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by tx_bridge_unit async fifo overflow
parameter           PCS_CH3_INT_TX_MASK_1 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by tx bridge unit underflow;
parameter           PCS_CH3_INT_TX_MASK_2 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by tx_invalid_k 
parameter           PCS_CH3_INT_TX_CLR_0 = "FALSE",     // FALSE,TRUE  active high to clr int triggered by tx bridge unit overflow;
parameter           PCS_CH3_INT_TX_CLR_1 = "FALSE",     // FALSE,TRUE  active high to clr int triggered by tx_bridge_unit async fifo underflow
parameter           PCS_CH3_INT_TX_CLR_2 = "FALSE",     // FALSE,TRUE  active high to clr int triggered by tx_invalid_k
parameter           PCS_CH3_TX_PMA_TCLK_POLINV = "PMA_TCLK",        // 1'b0:pma_tclk 1'b1:reverse of pma_tclk
parameter           PCS_CH3_TX_PCS_CLK_EN_SEL = "FALSE",        // FALSE,TRUE
parameter           PCS_CH3_TX_BRIDGE_TCLK_SEL = "PCS_TCLK",        // 1'b0: pcs_tclk 1'b1:tclk
parameter           PCS_CH3_TX_TCLK_POLINV = "TCLK",        // 1'b0:tclk 1'b1:reverse of tclk
parameter           PCS_CH3_TX_PCS_TX_RSTN = "FALSE",       // 1:pcs_tx_rstn is valued,is 0;0:pcs_tx_rstn is released
parameter           PCS_CH3_TX_SLAVE = "SLAVE",     // 1:slave channel,0:master channel
parameter           PCS_CH3_TX_BRIDGE_CLK_EN_SEL = "FALSE",     // FALSE,TRUE
parameter           PCS_CH3_DATA_WIDTH_MODE = "X20",        // 20bit,16bit,10bit,8bit
parameter           PCS_CH3_TX_TCLK2FABRIC_SEL = "FALSE",       // FALSE,TRUE
parameter           PCS_CH3_TX_OUTZZ = "FALSE",     // 1:16bit/32bit only;0:other data width mode
parameter           PCS_CH3_ENC_DUAL = "FALSE",     // FALSE,TRUE
parameter           PCS_CH3_TX_BITSLIP_DATA_MODE = "X10",       // 1: 20bit,0: 10bit
parameter   integer PCS_CH3_COMMA_REG1 = 0,     // 
parameter   integer PCS_CH3_RAPID_IMAX = 0,     // 
parameter   integer PCS_CH3_RAPID_VMIN_1 = 0,       // 
parameter   integer PCS_CH3_RAPID_VMIN_2 = 0,       // 
parameter           PCS_CH3_RX_PRBS_MODE = "DISABLE",       // Mode select:4'd0: reserved,4'd1: PRBS-7,4'd2: PRBS-15,4'd3: PRBS-23,4'd4: PRBS-31,4'd5: long "1",4'd6: long "0",4'd7: 20UI square wave,4'd8: D10_2,4'd9: PCIe complianece pattern,Others: reserved
parameter           PCS_CH3_RX_ERRCNT_CLR = "FALSE",        // FALSE,TRUE
parameter           PCS_CH3_TX_PRBS_MODE = "DISABLE",       // Mode select:4'd0: reserved,4'd1: PRBS-7,4'd2: PRBS-15,4'd3: PRBS-23,4'd4: PRBS-31,4'd5: long "1",4'd6: long "0",4'd7: 20UI square wave,4'd8: D10_2,4'd9: PCIe complianece pattern,Others: reserved
parameter           PCS_CH3_TX_INSERT_ER = "FALSE",     // FALSE,TRUE
parameter           PCS_CH3_ENABLE_PRBS_GEN = "FALSE",      // FALSE,TRUE
parameter   integer PCS_CH3_ERR_CNT = 0,        // 
parameter   integer PCS_CH3_DEFAULT_RADDR = 0,      // 
parameter   integer PCS_CH3_MASTER_CHECK_OFFSET = 0,        // 
parameter   integer PCS_CH3_DELAY_SET = 0,      // 
parameter           PCS_CH3_SEACH_OFFSET = "20BIT",     // 20bit,30bit,40bit,50bit,60bit,70bit
parameter   integer PCS_CH3_CEB_RAPIDLS_MMAX = 0,       // 
parameter   integer PCS_CH3_CTC_AFULL = 0,      // 
parameter   integer PCS_CH3_CTC_AEMPTY = 0,     // 
parameter   integer PCS_CH3_CTC_CONTI_SKP_SET  = 0,     //2018/7/18  
parameter           PCS_CH3_FAR_LOOP = "FALSE",     // FALSE,TRUE
parameter           PCS_CH3_NEAR_LOOP = "FALSE",       // FALSE,TRUE
parameter           PCS_CH3_INT_RX_MASK_0 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by pcs_lsm_synced
parameter           PCS_CH3_INT_RX_MASK_1 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by pcs_rx_mcb_status
parameter           PCS_CH3_INT_RX_MASK_2 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by channel bonding async fifo overflow
parameter           PCS_CH3_INT_RX_MASK_3 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by channel bonding async fifo underflow
parameter           PCS_CH3_INT_RX_MASK_4 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by ctc unit async fifo overflow
parameter           PCS_CH3_INT_RX_MASK_5 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by ctc unit async fifo underflow
parameter           PCS_CH3_INT_RX_MASK_6 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by rx_bridge_unit async fifo overflow
parameter           PCS_CH3_INT_RX_MASK_7 = "FALSE",        // FALSE,TRUE  active high to mask int triggered by rx_bridge_unit async fifo underflow
parameter           PCS_CH3_INT_RX_CLR_0 = "FALSE",     // FALSE,TRUE  active high to clr int triggered by pcs_lsm_synced
parameter           PCS_CH3_INT_RX_CLR_1 = "FALSE",     // FALSE,TRUE  active high to clr int triggered by pcs_rx_mcb_status
parameter           PCS_CH3_INT_RX_CLR_2 = "FALSE",     // FALSE,TRUE  active high to clr int triggered by channel bonding async fifo overflow
parameter           PCS_CH3_INT_RX_CLR_3 = "FALSE",     // FALSE,TRUE  active high to clr int triggered by channel bonding async fifo underflow
parameter           PCS_CH3_INT_RX_CLR_4 = "FALSE",     // FALSE,TRUE  active high to clr int triggered by ctc unit async fifo overflow
parameter           PCS_CH3_INT_RX_CLR_5 = "FALSE",     // FALSE,TRUE  active high to clr int triggered by ctc unit async fifo underflow
parameter           PCS_CH3_INT_RX_CLR_6 = "FALSE",     // FALSE,TRUE  active high to clr int triggered by rx_bridge_unit async fifo overflow
parameter           PCS_CH3_INT_RX_CLR_7 = "FALSE",     // FALSE,TRUE  active high to clr int triggered by rx_bridge_unit async fifo underflow
///PCS LANE end     
                   
//PMA LANE0 begin   
//PMA LANE Rx begin 
parameter           PMA_CH0_REG_RX_PD                   = "ON",          //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_CH0_REG_RX_PD_EN                = "FALSE",       //FALSE,TRUE   
parameter           PMA_CH0_REG_RX_CLKPATH_PD           = "ON",          //ON,OFF   ON=poweron,OFF= powerdown,reserved
parameter           PMA_CH0_REG_RX_CLKPATH_PD_EN        = "FALSE",       //FALSE,TRUE  ,reserved
parameter           PMA_CH0_REG_RX_DATAPATH_PD          = "ON",          //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_CH0_REG_RX_DATAPATH_PD_EN       = "FALSE",       //FALSE,TRUE
parameter           PMA_CH0_REG_RX_SIGDET_PD            = "ON",          //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_CH0_REG_RX_SIGDET_PD_EN         = "FALSE",       //FALSE,TRUE 
parameter           PMA_CH0_REG_RX_DCC_RST_N            = "TRUE",        //FALSE,TRUE  FALSE=low, TRUE=high
parameter           PMA_CH0_REG_RX_DCC_RST_N_EN         = "FALSE",       //FALSE,TRUE
parameter           PMA_CH0_REG_RX_CDR_RST_N            = "TRUE",        //FALSE,TRUE  FALSE=low, TRUE=high
parameter           PMA_CH0_REG_RX_CDR_RST_N_EN         = "FALSE",       //FALSE,TRUE
parameter           PMA_CH0_REG_RX_SIGDET_RST_N         = "TRUE",        //FALSE,TRUE  FALSE=low, TRUE=high
parameter           PMA_CH0_REG_RX_SIGDET_RST_N_EN      = "FALSE",       //FALSE,TRUE
parameter           PMA_CH0_REG_RXPCLK_SLIP             = "FALSE",       //FALSE,TRUE
parameter           PMA_CH0_REG_RXPCLK_SLIP_OW          = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH0_REG_RX_PCLKSWITCH_RST_N     = "TRUE",        //FALSE,TRUE  FALSE=low, TRUE=high
parameter           PMA_CH0_REG_RX_PCLKSWITCH_RST_N_EN  = "FALSE",       //FALSE,TRUE
parameter           PMA_CH0_REG_RX_PCLKSWITCH           = "FALSE",       //FALSE,TRUE
parameter           PMA_CH0_REG_RX_PCLKSWITCH_EN        = "FALSE",       //FALSE,TRUE
parameter           PMA_CH0_REG_RX_HIGHZ                = "FALSE",       //FALSE,TRUE
parameter           PMA_CH0_REG_RX_HIGHZ_EN             = "FALSE",       //FALSE,TRUE
parameter   integer PMA_CH0_REG_RX_EQ_C_SET             = 8,             // 
parameter   integer PMA_CH0_REG_RX_EQ_R_SET             = 8,             // 
parameter           PMA_CH0_REG_RX_BUSWIDTH             = "20BIT" ,      //"8BIT","10BIT","16BIT","20BIT" 
parameter           PMA_CH0_REG_RX_BUSWIDTH_EN          = "FALSE",       //FALSE,TRUE
parameter           PMA_CH0_REG_RX_RATE                 = "DIV1",        //"DIV8","DIV4","DIV2","DIV1"           
parameter           PMA_CH0_REG_RX_RATE_EN              = "FALSE",       //FALSE,TRUE
parameter   integer PMA_CH0_REG_RX_RES_TRIM             = 51,            //
parameter           PMA_CH0_REG_RX_RES_TRIM_EN          = "FALSE",       //FALSE,TRUE
parameter           PMA_CH0_REG_RX_EQ_OFF               = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high
parameter   integer PMA_CH0_REG_RX_PREAMP_IC            = 1367,          //
parameter           PMA_CH0_REG_RX_PCLK_EDGE_SEL        = "POS_EDGE",    //"POS_EDGE","NEG_EDGE"
parameter   integer PMA_CH0_REG_RX_PIBUF_IC             = 2,             //
parameter   integer PMA_CH0_REG_RX_DCC_IC_RX            = 3,             //
parameter   integer PMA_CH0_REG_RX_DCC_IC_TX            = 3,             //
parameter           PMA_CH0_REG_RX_ICTRL_TRX            = "100PCT",      //"87_5PCT","100PCT","112_5PCT","125PCT" 
////parameter       PMA_CH0_REG_RX_ICTRL_SIGDET         = "100PCT",     //"87_5PCT","100PCT","112_5PCT","125PCT"  
parameter   integer PMA_CH0_REG_RX_ICTRL_SIGDET         = 5,
parameter           PMA_CH0_REG_RX_ICTRL_PREAMP         = "100PCT",      //"87_5PCT","100PCT","112_5PCT","125PCT"  
parameter           PMA_CH0_REG_RX_ICTRL_SLICER         = "100PCT",      //"87_5PCT","100PCT","112_5PCT","125PCT"  
parameter           PMA_CH0_REG_RX_ICTRL_PIBUF          = "100PCT",      //"87_5PCT","100PCT","112_5PCT","125PCT" 
parameter           PMA_CH0_REG_RX_ICTRL_PI             = "100PCT",      //"87_5PCT","100PCT","112_5PCT","125PCT" 
parameter           PMA_CH0_REG_RX_ICTRL_DCC            = "100PCT",      //"87_5PCT","100PCT","112_5PCT","125PCT"
parameter           PMA_CH0_REG_RX_ICTRL_PREDRV         = "100PCT",      //"87_5PCT","100PCT","112_5PCT","125PCT"
parameter           PMA_CH0_REG_TX_RATE                 = "DIV1",        //"DIV8","DIV4","DIV2","DIV1"  
parameter           PMA_CH0_REG_TX_RATE_EN              = "FALSE",       //FALSE,TRUE
parameter           PMA_CH0_REG_RX_TX2RX_PLPBK_RST_N    = "TRUE",        //FALSE,TRUE  FALSE=low, TRUE=high
parameter           PMA_CH0_REG_RX_TX2RX_PLPBK_RST_N_EN = "FALSE",       //FALSE,TRUE
parameter           PMA_CH0_REG_RX_TX2RX_PLPBK_EN       = "FALSE",       //FALSE,TRUE
parameter           PMA_CH0_REG_TXCLK_SEL               = "PLL",         //"PLL","RXCLK"
parameter           PMA_CH0_REG_RX_DATA_POLARITY        = "NORMAL",      //"NORMAL","REVERSE"
parameter           PMA_CH0_REG_RX_ERR_INSERT           = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high
parameter           PMA_CH0_REG_UDP_CHK_EN              = "FALSE",       //FALSE,TRUE
parameter           PMA_CH0_REG_PRBS_SEL                = "PRBS7",       //"PRBS7","PRBS15","PRBS23","PRBS31"
parameter           PMA_CH0_REG_PRBS_CHK_EN             = "FALSE",       //FALSE,TRUE
parameter           PMA_CH0_REG_PRBS_CHK_WIDTH_SEL      = "20BIT",       //"8BIT","10BIT","16BIT","20BIT"
parameter           PMA_CH0_REG_BIST_CHK_PAT_SEL        = "PRBS",        //"PRBS","CONSTANT"
parameter           PMA_CH0_REG_LOAD_ERR_CNT            = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH0_REG_CHK_COUNTER_EN          = "FALSE",       //FALSE,TRUE
parameter   integer PMA_CH0_REG_CDR_PROP_GAIN           = 2,             //
parameter   integer PMA_CH0_REG_CDR_PROP_TURBO_GAIN     = 6,             //
parameter   integer PMA_CH0_REG_CDR_INT_GAIN            = 2,             //
parameter   integer PMA_CH0_REG_CDR_INT_TURBO_GAIN      = 6,             //      
parameter   integer PMA_CH0_REG_CDR_INT_SAT_MAX         = 992,          //
parameter   integer PMA_CH0_REG_CDR_INT_SAT_MIN         = 32,            //
parameter           PMA_CH0_REG_CDR_INT_RST             = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high
parameter           PMA_CH0_REG_CDR_INT_RST_OW          = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH0_REG_CDR_PROP_RST            = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high 
parameter           PMA_CH0_REG_CDR_PROP_RST_OW         = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH0_REG_CDR_LOCK_RST            = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high 
parameter           PMA_CH0_REG_CDR_LOCK_RST_OW         = "DISABLE",     //DISABLE,ENABLE
parameter   integer PMA_CH0_REG_CDR_RX_PI_FORCE_SEL     = 0,             //
parameter   integer PMA_CH0_REG_CDR_RX_PI_FORCE_D       = 0,             //
parameter           PMA_CH0_REG_CDR_LOCK_TIMER          = "1_2U",        //"0_8U","1_2U","1_6U","2_4U","3_2U","4_8U","12_8U","25_6U"
parameter   integer PMA_CH0_REG_CDR_TURBO_MODE_TIMER    = 1,             //  
parameter           PMA_CH0_REG_CDR_LOCK_VAL            = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high 
parameter           PMA_CH0_REG_CDR_LOCK_OW             = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH0_REG_CDR_INT_SAT_DET_EN      = "TRUE",       //FALSE,TRUE
parameter           PMA_CH0_REG_CDR_SAT_DET_STATUS_EN   = "FALSE",       //FALSE,TRUE
parameter           PMA_CH0_REG_CDR_SAT_DET_STATUS_RESET_EN = "FALSE",       //FALSE,TRUE
parameter           PMA_CH0_REG_CDR_PI_CTRL_RST         = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high 
parameter           PMA_CH0_REG_CDR_PI_CTRL_RST_OW      = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH0_REG_CDR_SAT_DET_RST         = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high 
parameter           PMA_CH0_REG_CDR_SAT_DET_RST_OW      = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH0_REG_CDR_SAT_DET_STICKY_RST  = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high
parameter           PMA_CH0_REG_CDR_SAT_DET_STICKY_RST_OW = "DISABLE",   //DISABLE,ENABLE
parameter           PMA_CH0_REG_CDR_SIGDET_STATUS_DIS   = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high
parameter   integer PMA_CH0_REG_CDR_SAT_DET_TIMER       = 2,            //
parameter           PMA_CH0_REG_CDR_SAT_DET_STATUS_VAL  = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high
parameter           PMA_CH0_REG_CDR_SAT_DET_STATUS_OW   = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH0_REG_CDR_TURBO_MODE_EN       = "TRUE",       //FALSE,TRUE  
parameter   integer PMA_CH0_REG_CDR_STATUS_RADDR_INIT   = 0,             //
parameter           PMA_CH0_REG_CDR_STATUS_FIFO_EN      = "TRUE",       //FALSE,TRUE
parameter   integer PMA_CH0_REG_PMA_TEST_SEL            = 0,             //
parameter   integer PMA_CH0_REG_OOB_COMWAKE_GAP_MIN     = 3,             //
parameter   integer PMA_CH0_REG_OOB_COMWAKE_GAP_MAX     = 11,            //
parameter   integer PMA_CH0_REG_OOB_COMINIT_GAP_MIN     = 15,            //
parameter   integer PMA_CH0_REG_OOB_COMINIT_GAP_MAX     = 35,            //
parameter   integer PMA_CH0_REG_RX_PIBUF_IC_TX          = 1,            //
parameter   integer PMA_CH0_REG_COMWAKE_STATUS_CLEAR    = 0,            //
parameter   integer PMA_CH0_REG_COMINIT_STATUS_CLEAR    = 0,            //
parameter           PMA_CH0_REG_RX_SYNC_RST_N_EN        = "FALSE",       //FALSE,TRUE
parameter           PMA_CH0_REG_RX_SYNC_RST_N           = "TRUE",        //FALSE,TRUE  FALSE=low, TRUE=high           
parameter           PMA_CH0_REG_RX_SATA_COMINIT_OW      = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH0_REG_RX_SATA_COMINIT         = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high    
parameter           PMA_CH0_REG_RX_SATA_COMWAKE_OW      = "DISABLE",     //DISABLE,ENABLE      
parameter           PMA_CH0_REG_RX_SATA_COMWAKE         = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high          
parameter           PMA_CH0_REG_RX_DCC_DISABLE          = "ENABLE",      //DISABLE,ENABLE   
parameter           PMA_CH0_REG_TX_DCC_DISABLE          = "ENABLE",      //DISABLE,ENABLE  
parameter           PMA_CH0_REG_RX_SLIP_SEL_EN          = "FALSE",       //FALSE,TRUE
parameter   integer PMA_CH0_REG_RX_SLIP_SEL             = 0,            //
parameter           PMA_CH0_REG_RX_SLIP_EN              = "FALSE",       //FALSE,TRUE
parameter   integer PMA_CH0_REG_RX_SIGDET_STATUS_SEL    = 5,            //
parameter           PMA_CH0_REG_RX_SIGDET_FSM_RST_N     = "TRUE",        //FALSE,TRUE  FALSE=low, TRUE=high     
parameter           PMA_CH0_REG_RX_SIGDET_STATUS_OW     = "DISABLE",     //DISABLE,ENABLE    
parameter           PMA_CH0_REG_RX_SIGDET_STATUS        = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high         
parameter           PMA_CH0_REG_RX_SIGDET_VTH           = "50MV",        //"12_5MV","25MV","37_5MV","50MV","62_5MV","75MV","87_5MV","100MV"
parameter   integer PMA_CH0_REG_RX_SIGDET_GRM           = 0,             // 
parameter           PMA_CH0_REG_RX_SIGDET_PULSE_EXT     = "DISABLE",     //DISABLE,ENABLE  
parameter   integer PMA_CH0_REG_RX_SIGDET_CH2_SEL       = 0,             // 
parameter   integer PMA_CH0_REG_RX_SIGDET_CH2_CHK_WINDOW =3,             //
parameter           PMA_CH0_REG_RX_SIGDET_CHK_WINDOW_EN = "TRUE",       //FALSE,TRUE
parameter   integer PMA_CH0_REG_RX_SIGDET_NOSIG_COUNT_SETTING = 4,       //
parameter   integer PMA_CH0_REG_RX_SIGDET_OOB_DET_COUNT_VAL= 0,             //
parameter           PMA_CH0_REG_SLIP_FIFO_INV_EN        = "FALSE",       //FALSE,TRUE
parameter           PMA_CH0_REG_SLIP_FIFO_INV           = "POS_EDGE",    //POS_EDGE,NEG_EDGE
parameter   integer PMA_CH0_REG_RX_SIGDET_4OOB_DET_SEL  =7,              //
////parameter   integer PMA_CH0_REG_RX_SIGDET_CHK_WINDOW    = 5,             //
////parameter   integer PMA_CH0_REG_RX_SIGDET_CHK_WINDOW_COUNT =3,             //
////parameter           PMA_CH0_REG_RX_SIGDET_LONG_CHK_WINDOW_EN = "DISABLE",  //DISABLE,ENABLE  
////parameter   integer PMA_CH0_REG_RX_SIGDET_LONG_CHK_WINDOW = 25,          //
parameter   integer PMA_CH0_REG_RX_SIGDET_IC_I          = 10,            //
parameter           PMA_CH0_REG_RX_OOB_DETECTOR_RESET_N_OW = "DISABLE",  //DISABLE,ENABLE
parameter           PMA_CH0_REG_RX_OOB_DETECTOR_RESET_N = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high  
parameter           PMA_CH0_REG_RX_OOB_DETECTOR_PD_OW   = "DISABLE",     //DISABLE,ENABLE  
parameter           PMA_CH0_REG_RX_OOB_DETECTOR_PD      = "ON",          //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_CH0_REG_RX_TERM_CM_CTRL         = "5DIV7",       //"5DIV7","2DIV3","5DIV6","4DIV5"
//PMA LANE Rx end
//PMA LANE Tx begin  
parameter           PMA_CH0_REG_TX_PD                   = "ON",          //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_CH0_REG_TX_PD_OW                = "DISABLE",     //DISABLE,ENABLE       
parameter           PMA_CH0_REG_TX_CLKPATH_PD           = "ON",          //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_CH0_REG_TX_CLKPATH_PD_OW        = "DISABLE",     //DISABLE,ENABLE
parameter   integer PMA_CH0_REG_TX_BEACON_TIMER_SEL     = 0,            // 
parameter           PMA_CH0_REG_TX_RXDET_REQ_OW         = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH0_REG_TX_RXDET_REQ            = "FALSE",      //FALSE,TRUE FALSE=low, TRUE=high
parameter           PMA_CH0_REG_TX_BEACON_EN_OW         = "DISABLE",     //DISABLE,ENABLE         
parameter           PMA_CH0_REG_TX_BEACON_EN            = "FALSE",      //FALSE,TRUE
parameter           PMA_CH0_REG_TX_EI_EN_OW             = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH0_REG_TX_EI_EN                = "FALSE",      //FALSE,TRUE
parameter           PMA_CH0_REG_TX_RES_CAL_EN           = "FALSE",      //FALSE,TRUE
parameter   integer PMA_CH0_REG_TX_RES_CAL              = 51,           // 
parameter           PMA_CH0_REG_TX_BIAS_CAL_EN          = "FALSE",      //FALSE,TRUE
parameter   integer PMA_CH0_REG_TX_BIAS_CTRL            = 48,           //
parameter           PMA_CH0_REG_TX_RXDET_TIMER_SEL      = "12CYCLE",     //"3CYCLE","12CYCLE","24CYCLE","36CYCLE"
parameter           PMA_CH0_REG_TX_SYNC_OW              = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH0_REG_TX_SYNC                 = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH0_REG_TX_PD_POST              = "OFF",        //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_CH0_REG_TX_PD_POST_OW           = "DISABLE",      //DISABLE,ENABLE
parameter           PMA_CH0_REG_TX_RESET_N_OW           = "DISABLE",     //DISABLE,ENABLE     
parameter           PMA_CH0_REG_TX_RESET_N              = "TRUE",       //FALSE,TRUE FALSE=low, TRUE=high 
parameter           PMA_CH0_REG_TX_DCC_RESET_N_OW       = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH0_REG_TX_DCC_RESET_N          = "TRUE",        //FALSE,TRUE FALSE=low, TRUE=high
parameter           PMA_CH0_REG_TX_BUSWIDTH_OW          = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH0_REG_TX_BUSWIDTH             = "20BIT",       //"8BIT","10BIT","16BIT","20BIT"
parameter           PMA_CH0_REG_PLL_READY_OW            = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH0_REG_PLL_READY               = "TRUE",        //FALSE,TRUE FALSE=low, TRUE=high 
parameter           PMA_CH0_REG_TX_PCLK_SW_OW           = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH0_REG_TX_PCLK_SW              = "TRUE",        //FALSE,TRUE FALSE=low, TRUE=high 
parameter   integer PMA_CH0_REG_EI_PCLK_DELAY_SEL       = 0,             //
parameter   integer PMA_CH0_REG_TX_DRV01_DAC0           = 0,             //
parameter   integer PMA_CH0_REG_TX_DRV01_DAC1           = 10,            //
parameter   integer PMA_CH0_REG_TX_DRV01_DAC2           = 16,            //
parameter   integer PMA_CH0_REG_TX_DRV00_DAC0           = 63,            //
parameter   integer PMA_CH0_REG_TX_DRV00_DAC1           = 53,            //
parameter   integer PMA_CH0_REG_TX_DRV00_DAC2           = 48,            //
parameter   integer PMA_CH0_REG_TX_AMP0                 = 8,             //
parameter   integer PMA_CH0_REG_TX_AMP1                 = 16,            //
parameter   integer PMA_CH0_REG_TX_AMP2                 = 32,            //
parameter   integer PMA_CH0_REG_TX_AMP3                 = 48,            //
parameter   integer PMA_CH0_REG_TX_AMP4                 = 56,            //
parameter   integer PMA_CH0_REG_TX_MARGIN               = 0,             // 
parameter           PMA_CH0_REG_TX_MARGIN_OW            = "DISABLE",     //DISABLE,ENABLE
parameter   integer PMA_CH0_REG_TX_DEEMP                = 0,            // 
parameter           PMA_CH0_REG_TX_DEEMP_OW             = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH0_REG_TX_SWING                = "FALSE",      //FALSE,TRUE FALSE=low, TRUE=high
parameter           PMA_CH0_REG_TX_SWING_OW             = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH0_REG_TX_RXDET_THRESHOLD      = "100MV",       //"50MV","75MV","100MV","125MV"
parameter   integer PMA_CH0_REG_TX_BEACON_OSC_CTRL      = 4,            //
parameter   integer PMA_CH0_REG_TX_PREDRV_DAC           = 1,            //
parameter   integer PMA_CH0_REG_TX_PREDRV_CM_CTRL       = 1,            //
parameter           PMA_CH0_REG_TX_TX2RX_SLPBACK_EN     = "FALSE",      //FALSE,TRUE
parameter           PMA_CH0_REG_TX_PCLK_EDGE_SEL        = "POS_EDGE",    //"NEG_EDGE","POS_EDGE"
parameter           PMA_CH0_REG_TX_RXDET_STATUS_OW      = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH0_REG_TX_RXDET_STATUS         = "TRUE",        //FALSE,TRUE FALSE=low, TRUE=high 
parameter           PMA_CH0_REG_TX_PRBS_GEN_EN          = "FALSE",      //FALSE,TRUE     
parameter           PMA_CH0_REG_TX_PRBS_GEN_WIDTH_SEL   = "20BIT",       //"8BIT","10BIT","16BIT","20BIT"
parameter           PMA_CH0_REG_TX_PRBS_SEL             = "PRBS7",       //"PRBS7","PRBS15","PRBS23","PRBS31"
parameter   integer PMA_CH0_REG_TX_UDP_DATA             = 256773,        //
parameter           PMA_CH0_REG_TX_FIFO_RST_N           = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high 
parameter   integer PMA_CH0_REG_TX_FIFO_WP_CTRL         = 2,             //
parameter           PMA_CH0_REG_TX_FIFO_EN              = "FALSE",       //FALSE,TRUE         
parameter   integer PMA_CH0_REG_TX_DATA_MUX_SEL         = 2,             //
parameter           PMA_CH0_REG_TX_ERR_INSERT           = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high 
parameter           PMA_CH0_REG_TX_SATA_EN              = "FALSE",       //FALSE,TRUE                   
parameter           PMA_CH0_REG_RATE_CHANGE_TXPCLK_ON_OW = "DISABLE",    //DISABLE,ENABLE 
parameter           PMA_CH0_REG_RATE_CHANGE_TXPCLK_ON   = "ENABLE",      //DISABLE,ENABLE 
parameter   integer PMA_CH0_REG_TX_PULLUP_DAC0          = 8,             //
parameter   integer PMA_CH0_REG_TX_PULLUP_DAC1          = 8,             //
parameter   integer PMA_CH0_REG_TX_PULLUP_DAC2          = 8,             //
parameter   integer PMA_CH0_REG_TX_PULLUP_DAC3          = 8,             //
parameter   integer PMA_CH0_REG_TX_OOB_DELAY_SEL        = 0,             //
parameter           PMA_CH0_REG_TX_POLARITY             = "NORMAL",      //"NORMAL","REVERSE"
parameter   integer PMA_CH0_REG_TX_SLPBK_AMP            = 1,             //
parameter           PMA_CH0_REG_TX_LS_MODE_EN           = "FALSE",       //FALSE,TRUE   
parameter           PMA_CH0_REG_TX_JTAG_MODE_EN_OW      = "DISABLE",    //DISABLE,ENABLE 
parameter           PMA_CH0_REG_TX_JTAG_MODE_EN         = "FALSE",       //FALSE,TRUE
parameter           PMA_CH0_REG_RX_JTAG_MODE_EN_OW      = "DISABLE",    //DISABLE,ENABLE
parameter           PMA_CH0_REG_RX_JTAG_MODE_EN         = "FALSE",       //FALSE,TRUE
parameter           PMA_CH0_REG_RX_JTAG_OE              = "DISABLE",    //DISABLE,ENABLE 
parameter   integer PMA_CH0_REG_RX_ACJTAG_VHYSTSE       = 0,             //
parameter           PMA_CH0_REG_TX_FBCLK_FAR_EN         = "FALSE",       //FALSE,TRUE
parameter   integer PMA_CH0_REG_RX_TERM_MODE_CTRL       = 6,             //
parameter           PMA_CH0_REG_PLPBK_TXPCLK_EN         = "TRUE",        //FALSE,TRUE
//PMA LANE Tx end   
//PMA LANE CFG begin
parameter           PMA_CH0_CFG_LANE_POWERUP            = "OFF",         //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_CH0_CFG_PMA_POR_N               = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high    
parameter           PMA_CH0_CFG_RX_LANE_POWERUP         = "OFF",         //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_CH0_CFG_RX_PMA_RSTN             = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high   
parameter           PMA_CH0_CFG_TX_LANE_POWERUP         = "OFF",         //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_CH0_CFG_TX_PMA_RSTN             = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high
//PMA LANE CFG end  
////reserved reg    
parameter   integer PMA_CH0_REG_RESERVED_48_45          = 0,             //  
parameter   integer PMA_CH0_REG_RESERVED_69             = 0,             //
parameter   integer PMA_CH0_REG_RESERVED_77_76          = 0,             //
parameter   integer PMA_CH0_REG_RESERVED_171_164        = 0,             //
parameter   integer PMA_CH0_REG_RESERVED_175_172        = 0,             //
parameter   integer PMA_CH0_REG_RESERVED_190            = 0,             //
parameter   integer PMA_CH0_REG_RESERVED_233_232        = 0,             //
parameter   integer PMA_CH0_REG_RESERVED_235_234        = 0,             //
parameter   integer PMA_CH0_REG_RESERVED_241_240        = 0,             //
parameter   integer PMA_CH0_REG_RESERVED_285_283        = 0,             //
parameter   integer PMA_CH0_REG_RESERVED_286            = 0,             //
parameter   integer PMA_CH0_REG_RESERVED_295            = 0,             //
parameter   integer PMA_CH0_REG_RESERVED_298            = 0,             //
parameter   integer PMA_CH0_REG_RESERVED_332_325        = 0,             //
parameter   integer PMA_CH0_REG_RESERVED_340_333        = 0,             //
parameter   integer PMA_CH0_REG_RESERVED_348_341        = 0,             //
parameter   integer PMA_CH0_REG_RESERVED_354_349        = 0,             //
parameter   integer PMA_CH0_REG_RESERVED_373            = 0,             //
parameter   integer PMA_CH0_REG_RESERVED_376            = 0,             //
parameter   integer PMA_CH0_REG_RESERVED_452            = 0,             //
parameter   integer PMA_CH0_REG_RESERVED_502_499        = 0,             //
//parameter   integer PMA_CH0_REG_RESERVED_503            = 0,             // 
parameter   integer PMA_CH0_REG_RESERVED_506_505        = 0,            //
parameter   integer PMA_CH0_REG_RESERVED_550_549        = 0,            //
parameter   integer PMA_CH0_REG_RESERVED_556_552        = 0,            //
////reserved end    
//PMA LANE0 end   
                    
//PMA LANE1 begin   
//PMA LANE Rx begin 
parameter           PMA_CH1_REG_RX_PD                   = "ON",          //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_CH1_REG_RX_PD_EN                = "FALSE",       //FALSE,TRUE   
parameter           PMA_CH1_REG_RX_CLKPATH_PD           = "ON",         //ON,OFF   ON=poweron,OFF= powerdown,reserved
parameter           PMA_CH1_REG_RX_CLKPATH_PD_EN        = "FALSE",       //FALSE,TRUE  ,reserved
parameter           PMA_CH1_REG_RX_DATAPATH_PD          = "ON",         //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_CH1_REG_RX_DATAPATH_PD_EN       = "FALSE",       //FALSE,TRUE
parameter           PMA_CH1_REG_RX_SIGDET_PD            = "ON",         //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_CH1_REG_RX_SIGDET_PD_EN         = "FALSE",       //FALSE,TRUE
parameter           PMA_CH1_REG_RX_DCC_RST_N            = "TRUE",       //FALSE,TRUE  FALSE=low, TRUE=high
parameter           PMA_CH1_REG_RX_DCC_RST_N_EN         = "FALSE",       //FALSE,TRUE
parameter           PMA_CH1_REG_RX_CDR_RST_N            = "TRUE",       //FALSE,TRUE  FALSE=low, TRUE=high
parameter           PMA_CH1_REG_RX_CDR_RST_N_EN         = "FALSE",       //FALSE,TRUE
parameter           PMA_CH1_REG_RX_SIGDET_RST_N         = "TRUE",       //FALSE,TRUE  FALSE=low, TRUE=high
parameter           PMA_CH1_REG_RX_SIGDET_RST_N_EN      = "FALSE",       //FALSE,TRUE
parameter           PMA_CH1_REG_RXPCLK_SLIP             = "FALSE",      //FALSE,TRUE
parameter           PMA_CH1_REG_RXPCLK_SLIP_OW          = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH1_REG_RX_PCLKSWITCH_RST_N     = "TRUE",       //FALSE,TRUE  FALSE=low, TRUE=high
parameter           PMA_CH1_REG_RX_PCLKSWITCH_RST_N_EN  = "FALSE",       //FALSE,TRUE
parameter           PMA_CH1_REG_RX_PCLKSWITCH           = "FALSE",      //FALSE,TRUE
parameter           PMA_CH1_REG_RX_PCLKSWITCH_EN        = "FALSE",       //FALSE,TRUE
parameter           PMA_CH1_REG_RX_HIGHZ                = "FALSE",      //FALSE,TRUE
parameter           PMA_CH1_REG_RX_HIGHZ_EN             = "FALSE",       //FALSE,TRUE
parameter   integer PMA_CH1_REG_RX_EQ_C_SET             = 8,             // 
parameter   integer PMA_CH1_REG_RX_EQ_R_SET             = 8,             // 
parameter           PMA_CH1_REG_RX_BUSWIDTH             = "20BIT",       //"8BIT","10BIT","16BIT","20BIT" 
parameter           PMA_CH1_REG_RX_BUSWIDTH_EN          = "FALSE",       //FALSE,TRUE
parameter           PMA_CH1_REG_RX_RATE                 = "DIV1",       //"DIV8","DIV4","DIV2","DIV1"           
parameter           PMA_CH1_REG_RX_RATE_EN              = "FALSE",       //FALSE,TRUE
parameter   integer PMA_CH1_REG_RX_RES_TRIM             = 51,           //
parameter           PMA_CH1_REG_RX_RES_TRIM_EN          = "FALSE",       //FALSE,TRUE
parameter           PMA_CH1_REG_RX_EQ_OFF               = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high
parameter   integer PMA_CH1_REG_RX_PREAMP_IC            = 1367,          //
parameter           PMA_CH1_REG_RX_PCLK_EDGE_SEL        = "POS_EDGE",    //"POS_EDGE","NEG_EDGE"
parameter   integer PMA_CH1_REG_RX_PIBUF_IC             = 2,             //
parameter   integer PMA_CH1_REG_RX_DCC_IC_RX            = 3,             //
parameter   integer PMA_CH1_REG_RX_DCC_IC_TX            = 3,             //
parameter           PMA_CH1_REG_RX_ICTRL_TRX            = "100PCT",      //"87_5PCT","100PCT","112_5PCT","125PCT" 
////parameter           PMA_CH1_REG_RX_ICTRL_SIGDET         = "100PCT",      //"87_5PCT","100PCT","112_5PCT","125PCT"  
parameter   integer PMA_CH1_REG_RX_ICTRL_SIGDET         = 5,
parameter           PMA_CH1_REG_RX_ICTRL_PREAMP         = "100PCT",      //"87_5PCT","100PCT","112_5PCT","125PCT"  
parameter           PMA_CH1_REG_RX_ICTRL_SLICER         = "100PCT",      //"87_5PCT","100PCT","112_5PCT","125PCT"  
parameter           PMA_CH1_REG_RX_ICTRL_PIBUF          = "100PCT",      //"87_5PCT","100PCT","112_5PCT","125PCT" 
parameter           PMA_CH1_REG_RX_ICTRL_PI             = "100PCT",      //"87_5PCT","100PCT","112_5PCT","125PCT" 
parameter           PMA_CH1_REG_RX_ICTRL_DCC            = "100PCT",      //"87_5PCT","100PCT","112_5PCT","125PCT"
parameter           PMA_CH1_REG_RX_ICTRL_PREDRV         = "100PCT",      //"87_5PCT","100PCT","112_5PCT","125PCT"
parameter           PMA_CH1_REG_TX_RATE                 = "DIV1",        //"DIV8","DIV4","DIV2","DIV1"  
parameter           PMA_CH1_REG_TX_RATE_EN              = "FALSE",       //FALSE,TRUE
parameter           PMA_CH1_REG_RX_TX2RX_PLPBK_RST_N    = "TRUE",       //FALSE,TRUE  FALSE=low, TRUE=high
parameter           PMA_CH1_REG_RX_TX2RX_PLPBK_RST_N_EN = "FALSE",       //FALSE,TRUE
parameter           PMA_CH1_REG_RX_TX2RX_PLPBK_EN       = "FALSE",       //FALSE,TRUE
parameter           PMA_CH1_REG_TXCLK_SEL               = "PLL",         //"PLL","RXCLK"
parameter           PMA_CH1_REG_RX_DATA_POLARITY        = "NORMAL",      //"NORMAL","REVERSE"
parameter           PMA_CH1_REG_RX_ERR_INSERT           = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high
parameter           PMA_CH1_REG_UDP_CHK_EN              = "FALSE",       //FALSE,TRUE
parameter           PMA_CH1_REG_PRBS_SEL                = "PRBS7",       //"PRBS7","PRBS15","PRBS23","PRBS31"
parameter           PMA_CH1_REG_PRBS_CHK_EN             = "FALSE",       //FALSE,TRUE
parameter           PMA_CH1_REG_PRBS_CHK_WIDTH_SEL      = "20BIT",       //"8BIT","10BIT","16BIT","20BIT"
parameter           PMA_CH1_REG_BIST_CHK_PAT_SEL        = "PRBS",        //"PRBS","CONSTANT"
parameter           PMA_CH1_REG_LOAD_ERR_CNT            = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH1_REG_CHK_COUNTER_EN          = "FALSE",       //FALSE,TRUE 
parameter   integer PMA_CH1_REG_CDR_PROP_GAIN           = 2,             //
parameter   integer PMA_CH1_REG_CDR_PROP_TURBO_GAIN     = 6,             //
parameter   integer PMA_CH1_REG_CDR_INT_GAIN            = 2,             //
parameter   integer PMA_CH1_REG_CDR_INT_TURBO_GAIN      = 6,             //      
parameter   integer PMA_CH1_REG_CDR_INT_SAT_MAX         = 992,          //
parameter   integer PMA_CH1_REG_CDR_INT_SAT_MIN         = 32,            //
parameter           PMA_CH1_REG_CDR_INT_RST             = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high
parameter           PMA_CH1_REG_CDR_INT_RST_OW          = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH1_REG_CDR_PROP_RST            = "FALSE",      //FALSE,TRUE FALSE=low, TRUE=high 
parameter           PMA_CH1_REG_CDR_PROP_RST_OW         = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH1_REG_CDR_LOCK_RST            = "FALSE",      //FALSE,TRUE FALSE=low, TRUE=high 
parameter           PMA_CH1_REG_CDR_LOCK_RST_OW         = "DISABLE",     //DISABLE,ENABLE
parameter   integer PMA_CH1_REG_CDR_RX_PI_FORCE_SEL     = 0,             //
parameter   integer PMA_CH1_REG_CDR_RX_PI_FORCE_D       = 0,             //
parameter           PMA_CH1_REG_CDR_LOCK_TIMER          = "1_2U",        //"0_8U","1_2U","1_6U","2_4U","3_2U","4_8U","12_8U","25_6U"
parameter   integer PMA_CH1_REG_CDR_TURBO_MODE_TIMER    = 1,             //  
parameter           PMA_CH1_REG_CDR_LOCK_VAL            = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high 
parameter           PMA_CH1_REG_CDR_LOCK_OW             = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH1_REG_CDR_INT_SAT_DET_EN      = "TRUE",       //FALSE,TRUE
parameter           PMA_CH1_REG_CDR_SAT_DET_STATUS_EN   = "FALSE",       //FALSE,TRUE
parameter           PMA_CH1_REG_CDR_SAT_DET_STATUS_RESET_EN = "FALSE",       //FALSE,TRUE
parameter           PMA_CH1_REG_CDR_PI_CTRL_RST         = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high 
parameter           PMA_CH1_REG_CDR_PI_CTRL_RST_OW      = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH1_REG_CDR_SAT_DET_RST         = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high 
parameter           PMA_CH1_REG_CDR_SAT_DET_RST_OW      = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH1_REG_CDR_SAT_DET_STICKY_RST  = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high
parameter           PMA_CH1_REG_CDR_SAT_DET_STICKY_RST_OW = "DISABLE",   //DISABLE,ENABLE
parameter           PMA_CH1_REG_CDR_SIGDET_STATUS_DIS   = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high
parameter   integer PMA_CH1_REG_CDR_SAT_DET_TIMER       = 2,             //
parameter           PMA_CH1_REG_CDR_SAT_DET_STATUS_VAL  = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high
parameter           PMA_CH1_REG_CDR_SAT_DET_STATUS_OW   = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH1_REG_CDR_TURBO_MODE_EN       = "TRUE",       //FALSE,TRUE  
parameter   integer PMA_CH1_REG_CDR_STATUS_RADDR_INIT   = 0,             //
parameter           PMA_CH1_REG_CDR_STATUS_FIFO_EN      = "TRUE",       //FALSE,TRUE
parameter   integer PMA_CH1_REG_PMA_TEST_SEL            = 0,             //
parameter   integer PMA_CH1_REG_OOB_COMWAKE_GAP_MIN     = 3,             //
parameter   integer PMA_CH1_REG_OOB_COMWAKE_GAP_MAX     = 11,            //
parameter   integer PMA_CH1_REG_OOB_COMINIT_GAP_MIN     = 15,            //
parameter   integer PMA_CH1_REG_OOB_COMINIT_GAP_MAX     = 35,            //
parameter   integer PMA_CH1_REG_RX_PIBUF_IC_TX          = 1,             //
parameter   integer PMA_CH1_REG_COMWAKE_STATUS_CLEAR    = 0,             //
parameter   integer PMA_CH1_REG_COMINIT_STATUS_CLEAR    = 0,           //
parameter           PMA_CH1_REG_RX_SYNC_RST_N_EN        = "FALSE",       //FALSE,TRUE
parameter           PMA_CH1_REG_RX_SYNC_RST_N           = "TRUE",      //FALSE,TRUE  FALSE=low, TRUE=high           
parameter           PMA_CH1_REG_RX_SATA_COMINIT_OW      = "DISABLE",    //DISABLE,ENABLE
parameter           PMA_CH1_REG_RX_SATA_COMINIT         = "FALSE",     //FALSE,TRUE FALSE=low, TRUE=high    
parameter           PMA_CH1_REG_RX_SATA_COMWAKE_OW      = "DISABLE",    //DISABLE,ENABLE      
parameter           PMA_CH1_REG_RX_SATA_COMWAKE         = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high          
parameter           PMA_CH1_REG_RX_DCC_DISABLE          = "ENABLE",      //DISABLE,ENABLE   
parameter           PMA_CH1_REG_TX_DCC_DISABLE          = "ENABLE",      //DISABLE,ENABLE  
parameter           PMA_CH1_REG_RX_SLIP_SEL_EN          = "FALSE",       //FALSE,TRUE 
parameter   integer PMA_CH1_REG_RX_SLIP_SEL             = 0,             //
parameter           PMA_CH1_REG_RX_SLIP_EN              = "FALSE",       //FALSE,TRUE
parameter   integer PMA_CH1_REG_RX_SIGDET_STATUS_SEL    = 5,             //
parameter           PMA_CH1_REG_RX_SIGDET_FSM_RST_N     = "TRUE",        //FALSE,TRUE  FALSE=low, TRUE=high     
parameter           PMA_CH1_REG_RX_SIGDET_STATUS_OW     = "DISABLE",     //DISABLE,ENABLE    
parameter           PMA_CH1_REG_RX_SIGDET_STATUS        = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high         
parameter           PMA_CH1_REG_RX_SIGDET_VTH           = "50MV",        //"12_5MV","25MV","37_5MV","50MV","62_5MV","75MV","87_5MV","100MV"
parameter   integer PMA_CH1_REG_RX_SIGDET_GRM           = 0,             // 
parameter           PMA_CH1_REG_RX_SIGDET_PULSE_EXT     = "DISABLE",     //DISABLE,ENABLE  
parameter   integer PMA_CH1_REG_RX_SIGDET_CH2_SEL       = 0,             // 
parameter   integer PMA_CH1_REG_RX_SIGDET_CH2_CHK_WINDOW =3,             //
parameter           PMA_CH1_REG_RX_SIGDET_CHK_WINDOW_EN = "TRUE",       //FALSE,TRUE
parameter   integer PMA_CH1_REG_RX_SIGDET_NOSIG_COUNT_SETTING = 4,       //
parameter   integer PMA_CH1_REG_RX_SIGDET_OOB_DET_COUNT_VAL= 0,             //
parameter           PMA_CH1_REG_SLIP_FIFO_INV_EN        = "FALSE",       //FALSE,TRUE
parameter           PMA_CH1_REG_SLIP_FIFO_INV           = "POS_EDGE",    //POS_EDGE,NEG_EDGE
parameter   integer PMA_CH1_REG_RX_SIGDET_4OOB_DET_SEL   =7,             //
////parameter   integer PMA_CH1_REG_RX_SIGDET_CHK_WINDOW    = 5,             //
////parameter   integer PMA_CH1_REG_RX_SIGDET_CHK_WINDOW_COUNT =3,             //
////parameter           PMA_CH1_REG_RX_SIGDET_LONG_CHK_WINDOW_EN = "DISABLE",  //DISABLE,ENABLE  
////parameter   integer PMA_CH1_REG_RX_SIGDET_LONG_CHK_WINDOW = 25,          //
parameter   integer PMA_CH1_REG_RX_SIGDET_IC_I          = 10,            //
parameter           PMA_CH1_REG_RX_OOB_DETECTOR_RESET_N_OW = "DISABLE",  //DISABLE,ENABLE
parameter           PMA_CH1_REG_RX_OOB_DETECTOR_RESET_N = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high  
parameter           PMA_CH1_REG_RX_OOB_DETECTOR_PD_OW   = "DISABLE",     //DISABLE,ENABLE  
parameter           PMA_CH1_REG_RX_OOB_DETECTOR_PD      = "ON",          //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_CH1_REG_RX_TERM_CM_CTRL         = "5DIV7",       //"5DIV7","2DIV3","5DIV6","4DIV5"
//PMA LANE Rx end
//PMA LANE Tx begin  
parameter           PMA_CH1_REG_TX_PD                   = "ON",          //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_CH1_REG_TX_PD_OW                = "DISABLE",     //DISABLE,ENABLE       
parameter           PMA_CH1_REG_TX_CLKPATH_PD           = "ON",         //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_CH1_REG_TX_CLKPATH_PD_OW        = "DISABLE",     //DISABLE,ENABLE
parameter   integer PMA_CH1_REG_TX_BEACON_TIMER_SEL     = 0,            // 
parameter           PMA_CH1_REG_TX_RXDET_REQ_OW         = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH1_REG_TX_RXDET_REQ            = "FALSE",      //FALSE,TRUE FALSE=low, TRUE=high
parameter           PMA_CH1_REG_TX_BEACON_EN_OW         = "DISABLE",     //DISABLE,ENABLE         
parameter           PMA_CH1_REG_TX_BEACON_EN            = "FALSE",      //FALSE,TRUE
parameter           PMA_CH1_REG_TX_EI_EN_OW             = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH1_REG_TX_EI_EN                = "FALSE",      //FALSE,TRUE
parameter           PMA_CH1_REG_TX_RES_CAL_EN           = "FALSE",      //FALSE,TRUE
parameter   integer PMA_CH1_REG_TX_RES_CAL              = 51,           // 
parameter           PMA_CH1_REG_TX_BIAS_CAL_EN          = "FALSE",      //FALSE,TRUE
parameter   integer PMA_CH1_REG_TX_BIAS_CTRL            = 48,           //
parameter           PMA_CH1_REG_TX_RXDET_TIMER_SEL      = "12CYCLE",    //"3CYCLE","12CYCLE","24CYCLE","36CYCLE"
parameter           PMA_CH1_REG_TX_SYNC_OW              = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH1_REG_TX_SYNC                 = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH1_REG_TX_PD_POST              = "OFF",        //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_CH1_REG_TX_PD_POST_OW           = "DISABLE",      //DISABLE,ENABLE
parameter           PMA_CH1_REG_TX_RESET_N_OW           = "DISABLE",     //DISABLE,ENABLE     
parameter           PMA_CH1_REG_TX_RESET_N              = "TRUE",       //FALSE,TRUE FALSE=low, TRUE=high 
parameter           PMA_CH1_REG_TX_DCC_RESET_N_OW       = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH1_REG_TX_DCC_RESET_N          = "TRUE",       //FALSE,TRUE FALSE=low, TRUE=high
parameter           PMA_CH1_REG_TX_BUSWIDTH_OW          = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH1_REG_TX_BUSWIDTH             = "20BIT",      //"8BIT","10BIT","16BIT","20BIT"
parameter           PMA_CH1_REG_PLL_READY_OW            = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH1_REG_PLL_READY               = "TRUE",       //FALSE,TRUE FALSE=low, TRUE=high 
parameter           PMA_CH1_REG_TX_PCLK_SW_OW           = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH1_REG_TX_PCLK_SW              = "TRUE",        //FALSE,TRUE FALSE=low, TRUE=high 
parameter   integer PMA_CH1_REG_EI_PCLK_DELAY_SEL       = 0,             //
parameter   integer PMA_CH1_REG_TX_DRV01_DAC0           = 0,             //
parameter   integer PMA_CH1_REG_TX_DRV01_DAC1           = 10,            //
parameter   integer PMA_CH1_REG_TX_DRV01_DAC2           = 16,            //
parameter   integer PMA_CH1_REG_TX_DRV00_DAC0           = 63,            //
parameter   integer PMA_CH1_REG_TX_DRV00_DAC1           = 53,            //
parameter   integer PMA_CH1_REG_TX_DRV00_DAC2           = 48,            //
parameter   integer PMA_CH1_REG_TX_AMP0                 = 8,             //
parameter   integer PMA_CH1_REG_TX_AMP1                 = 16,            //
parameter   integer PMA_CH1_REG_TX_AMP2                 = 32,            //
parameter   integer PMA_CH1_REG_TX_AMP3                 = 48,            //
parameter   integer PMA_CH1_REG_TX_AMP4                 = 56,            //
parameter   integer PMA_CH1_REG_TX_MARGIN               = 0,             // 
parameter           PMA_CH1_REG_TX_MARGIN_OW            = "DISABLE",    //DISABLE,ENABLE
parameter   integer PMA_CH1_REG_TX_DEEMP                = 0,           // 
parameter           PMA_CH1_REG_TX_DEEMP_OW             = "DISABLE",    //DISABLE,ENABLE
parameter           PMA_CH1_REG_TX_SWING                = "FALSE",     //FALSE,TRUE FALSE=low, TRUE=high
parameter           PMA_CH1_REG_TX_SWING_OW             = "DISABLE",    //DISABLE,ENABLE
parameter           PMA_CH1_REG_TX_RXDET_THRESHOLD      = "100MV",       //"50MV","75MV","100MV","125MV"
parameter   integer PMA_CH1_REG_TX_BEACON_OSC_CTRL      = 4,             //
parameter   integer PMA_CH1_REG_TX_PREDRV_DAC           = 1,             //
parameter   integer PMA_CH1_REG_TX_PREDRV_CM_CTRL       = 1,             //
parameter           PMA_CH1_REG_TX_TX2RX_SLPBACK_EN     = "FALSE",      //FALSE,TRUE
parameter           PMA_CH1_REG_TX_PCLK_EDGE_SEL        = "POS_EDGE",    //"NEG_EDGE","POS_EDGE"
parameter           PMA_CH1_REG_TX_RXDET_STATUS_OW      = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH1_REG_TX_RXDET_STATUS         = "TRUE",        //FALSE,TRUE FALSE=low, TRUE=high 
parameter           PMA_CH1_REG_TX_PRBS_GEN_EN          = "FALSE",      //FALSE,TRUE     
parameter           PMA_CH1_REG_TX_PRBS_GEN_WIDTH_SEL   = "20BIT",       //"8BIT","10BIT","16BIT","20BIT"
parameter           PMA_CH1_REG_TX_PRBS_SEL             = "PRBS7",       //"PRBS7","PRBS15","PRBS23","PRBS31"
parameter   integer PMA_CH1_REG_TX_UDP_DATA             = 256773,        //
parameter           PMA_CH1_REG_TX_FIFO_RST_N           = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high 
parameter   integer PMA_CH1_REG_TX_FIFO_WP_CTRL         = 2,             //
parameter           PMA_CH1_REG_TX_FIFO_EN              = "FALSE",      //FALSE,TRUE         
parameter   integer PMA_CH1_REG_TX_DATA_MUX_SEL         = 2,             //
parameter           PMA_CH1_REG_TX_ERR_INSERT           = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high 
parameter           PMA_CH1_REG_TX_SATA_EN              = "FALSE",       //FALSE,TRUE                   
parameter           PMA_CH1_REG_RATE_CHANGE_TXPCLK_ON_OW = "DISABLE",    //DISABLE,ENABLE 
parameter           PMA_CH1_REG_RATE_CHANGE_TXPCLK_ON   = "ENABLE",      //DISABLE,ENABLE 
parameter   integer PMA_CH1_REG_TX_PULLUP_DAC0          = 8,             //
parameter   integer PMA_CH1_REG_TX_PULLUP_DAC1          = 8,             //
parameter   integer PMA_CH1_REG_TX_PULLUP_DAC2          = 8,             //
parameter   integer PMA_CH1_REG_TX_PULLUP_DAC3          = 8,             //
parameter   integer PMA_CH1_REG_TX_OOB_DELAY_SEL        = 0,             //
parameter           PMA_CH1_REG_TX_POLARITY             = "NORMAL",      //"NORMAL","REVERSE"
parameter   integer PMA_CH1_REG_TX_SLPBK_AMP            = 1,             //
parameter           PMA_CH1_REG_TX_LS_MODE_EN           = "FALSE",       //FALSE,TRUE   
parameter           PMA_CH1_REG_TX_JTAG_MODE_EN_OW      = "DISABLE",     //DISABLE,ENABLE 
parameter           PMA_CH1_REG_TX_JTAG_MODE_EN         = "FALSE",       //FALSE,TRUE
parameter           PMA_CH1_REG_RX_JTAG_MODE_EN_OW      = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH1_REG_RX_JTAG_MODE_EN         = "FALSE",       //FALSE,TRUE
parameter           PMA_CH1_REG_RX_JTAG_OE              = "DISABLE",     //DISABLE,ENABLE 
parameter   integer PMA_CH1_REG_RX_ACJTAG_VHYSTSE       = 0,             //
parameter           PMA_CH1_REG_TX_FBCLK_FAR_EN         = "FALSE",       //FALSE,TRUE
parameter   integer PMA_CH1_REG_RX_TERM_MODE_CTRL       = 6,             //
parameter           PMA_CH1_REG_PLPBK_TXPCLK_EN         = "TRUE",        //FALSE,TRUE
//PMA LANE Tx end
//PMA LANE CFG begin
parameter           PMA_CH1_CFG_LANE_POWERUP            = "OFF",         //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_CH1_CFG_PMA_POR_N               = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high    
parameter           PMA_CH1_CFG_RX_LANE_POWERUP         = "OFF",        //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_CH1_CFG_RX_PMA_RSTN             = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high   
parameter           PMA_CH1_CFG_TX_LANE_POWERUP         = "OFF",        //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_CH1_CFG_TX_PMA_RSTN             = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high
//PMA LANE CFG end
////reserved reg
parameter   integer PMA_CH1_REG_RESERVED_48_45          = 0,             //  
parameter   integer PMA_CH1_REG_RESERVED_69             = 0,             //
parameter   integer PMA_CH1_REG_RESERVED_77_76          = 0,             //
parameter   integer PMA_CH1_REG_RESERVED_171_164        = 0,             //
parameter   integer PMA_CH1_REG_RESERVED_175_172        = 0,             //
parameter   integer PMA_CH1_REG_RESERVED_190            = 0,             //
parameter   integer PMA_CH1_REG_RESERVED_233_232        = 0,             //
parameter   integer PMA_CH1_REG_RESERVED_235_234        = 0,             //
parameter   integer PMA_CH1_REG_RESERVED_241_240        = 0,             //
parameter   integer PMA_CH1_REG_RESERVED_285_283        = 0,             //
parameter   integer PMA_CH1_REG_RESERVED_286            = 0,             //
parameter   integer PMA_CH1_REG_RESERVED_295            = 0,             //
parameter   integer PMA_CH1_REG_RESERVED_298            = 0,             //
parameter   integer PMA_CH1_REG_RESERVED_332_325        = 0,             //
parameter   integer PMA_CH1_REG_RESERVED_340_333        = 0,             //
parameter   integer PMA_CH1_REG_RESERVED_348_341        = 0,             //
parameter   integer PMA_CH1_REG_RESERVED_354_349        = 0,             //
parameter   integer PMA_CH1_REG_RESERVED_373            = 0,             //
parameter   integer PMA_CH1_REG_RESERVED_376            = 0,             //
parameter   integer PMA_CH1_REG_RESERVED_452            = 0,             //
parameter   integer PMA_CH1_REG_RESERVED_502_499        = 0,             //
//parameter   integer PMA_CH1_REG_RESERVED_503            = 0,             // 
parameter   integer PMA_CH1_REG_RESERVED_506_505        = 0,             //
parameter   integer PMA_CH1_REG_RESERVED_550_549        = 0,             //
parameter   integer PMA_CH1_REG_RESERVED_556_552        = 0,             //
////reserved end
//PMA LANE1 end

//PMA LANE2 begin
//PMA LANE Rx begin 
parameter           PMA_CH2_REG_RX_PD                   = "ON",          //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_CH2_REG_RX_PD_EN                = "FALSE",       //FALSE,TRUE   
parameter           PMA_CH2_REG_RX_CLKPATH_PD           = "ON",         //ON,OFF   ON=poweron,OFF= powerdown,reserved
parameter           PMA_CH2_REG_RX_CLKPATH_PD_EN        = "FALSE",       //FALSE,TRUE  ,reserved 
parameter           PMA_CH2_REG_RX_DATAPATH_PD          = "ON",         //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_CH2_REG_RX_DATAPATH_PD_EN       = "FALSE",       //FALSE,TRUE
parameter           PMA_CH2_REG_RX_SIGDET_PD            = "ON",         //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_CH2_REG_RX_SIGDET_PD_EN         = "FALSE",       //FALSE,TRUE
parameter           PMA_CH2_REG_RX_DCC_RST_N            = "TRUE",       //FALSE,TRUE  FALSE=low, TRUE=high
parameter           PMA_CH2_REG_RX_DCC_RST_N_EN         = "FALSE",       //FALSE,TRUE
parameter           PMA_CH2_REG_RX_CDR_RST_N            = "TRUE",       //FALSE,TRUE  FALSE=low, TRUE=high
parameter           PMA_CH2_REG_RX_CDR_RST_N_EN         = "FALSE",       //FALSE,TRUE
parameter           PMA_CH2_REG_RX_SIGDET_RST_N         = "TRUE",       //FALSE,TRUE  FALSE=low, TRUE=high
parameter           PMA_CH2_REG_RX_SIGDET_RST_N_EN      = "FALSE",       //FALSE,TRUE
parameter           PMA_CH2_REG_RXPCLK_SLIP             = "FALSE",      //FALSE,TRUE
parameter           PMA_CH2_REG_RXPCLK_SLIP_OW          = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH2_REG_RX_PCLKSWITCH_RST_N     = "TRUE",       //FALSE,TRUE  FALSE=low, TRUE=high
parameter           PMA_CH2_REG_RX_PCLKSWITCH_RST_N_EN  = "FALSE",       //FALSE,TRUE
parameter           PMA_CH2_REG_RX_PCLKSWITCH           = "FALSE",      //FALSE,TRUE
parameter           PMA_CH2_REG_RX_PCLKSWITCH_EN        = "FALSE",       //FALSE,TRUE
parameter           PMA_CH2_REG_RX_HIGHZ                = "FALSE",      //FALSE,TRUE
parameter           PMA_CH2_REG_RX_HIGHZ_EN             = "FALSE",       //FALSE,TRUE
parameter   integer PMA_CH2_REG_RX_EQ_C_SET             = 8,            // 
parameter   integer PMA_CH2_REG_RX_EQ_R_SET             = 8,            // 
parameter           PMA_CH2_REG_RX_BUSWIDTH             = "20BIT",      //"8BIT","10BIT","16BIT","20BIT" 
parameter           PMA_CH2_REG_RX_BUSWIDTH_EN          = "FALSE",       //FALSE,TRUE
parameter           PMA_CH2_REG_RX_RATE                 = "DIV1",       //"DIV8","DIV4","DIV2","DIV1"           
parameter           PMA_CH2_REG_RX_RATE_EN              = "FALSE",       //FALSE,TRUE
parameter   integer PMA_CH2_REG_RX_RES_TRIM             = 51,           //
parameter           PMA_CH2_REG_RX_RES_TRIM_EN          = "FALSE",       //FALSE,TRUE
parameter           PMA_CH2_REG_RX_EQ_OFF               = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high
parameter   integer PMA_CH2_REG_RX_PREAMP_IC            = 1367,          //
parameter           PMA_CH2_REG_RX_PCLK_EDGE_SEL        = "POS_EDGE",    //"POS_EDGE","NEG_EDGE"
parameter   integer PMA_CH2_REG_RX_PIBUF_IC             = 2,             //
parameter   integer PMA_CH2_REG_RX_DCC_IC_RX            = 3,             //
parameter   integer PMA_CH2_REG_RX_DCC_IC_TX            = 3,             //
parameter           PMA_CH2_REG_RX_ICTRL_TRX            = "100PCT",      //"87_5PCT","100PCT","112_5PCT","125PCT" 
////parameter          PMA_CH2_REG_RX_ICTRL_SIGDET         = "100PCT",      //"87_5PCT","100PCT","112_5PCT","125PCT"  
parameter   integer PMA_CH2_REG_RX_ICTRL_SIGDET         = 5,      
parameter           PMA_CH2_REG_RX_ICTRL_PREAMP         = "100PCT",      //"87_5PCT","100PCT","112_5PCT","125PCT"  
parameter           PMA_CH2_REG_RX_ICTRL_SLICER         = "100PCT",      //"87_5PCT","100PCT","112_5PCT","125PCT"  
parameter           PMA_CH2_REG_RX_ICTRL_PIBUF          = "100PCT",      //"87_5PCT","100PCT","112_5PCT","125PCT" 
parameter           PMA_CH2_REG_RX_ICTRL_PI             = "100PCT",      //"87_5PCT","100PCT","112_5PCT","125PCT" 
parameter           PMA_CH2_REG_RX_ICTRL_DCC            = "100PCT",      //"87_5PCT","100PCT","112_5PCT","125PCT"
parameter           PMA_CH2_REG_RX_ICTRL_PREDRV         = "100PCT",      //"87_5PCT","100PCT","112_5PCT","125PCT"
parameter           PMA_CH2_REG_TX_RATE                 = "DIV1",        //"DIV8","DIV4","DIV2","DIV1"  
parameter           PMA_CH2_REG_TX_RATE_EN              = "FALSE",       //FALSE,TRUE
parameter           PMA_CH2_REG_RX_TX2RX_PLPBK_RST_N    = "TRUE",       //FALSE,TRUE  FALSE=low, TRUE=high
parameter           PMA_CH2_REG_RX_TX2RX_PLPBK_RST_N_EN = "FALSE",       //FALSE,TRUE
parameter           PMA_CH2_REG_RX_TX2RX_PLPBK_EN       = "FALSE",       //FALSE,TRUE
parameter           PMA_CH2_REG_TXCLK_SEL               = "PLL",         //"PLL","RXCLK"
parameter           PMA_CH2_REG_RX_DATA_POLARITY        = "NORMAL",      //"NORMAL","REVERSE"
parameter           PMA_CH2_REG_RX_ERR_INSERT           = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high
parameter           PMA_CH2_REG_UDP_CHK_EN              = "FALSE",       //FALSE,TRUE
parameter           PMA_CH2_REG_PRBS_SEL                = "PRBS7",       //"PRBS7","PRBS15","PRBS23","PRBS31"
parameter           PMA_CH2_REG_PRBS_CHK_EN             = "FALSE",       //FALSE,TRUE
parameter           PMA_CH2_REG_PRBS_CHK_WIDTH_SEL      = "20BIT",       //"8BIT","10BIT","16BIT","20BIT"
parameter           PMA_CH2_REG_BIST_CHK_PAT_SEL        = "PRBS",        //"PRBS","CONSTANT"
parameter           PMA_CH2_REG_LOAD_ERR_CNT            = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH2_REG_CHK_COUNTER_EN          = "FALSE",       //FALSE,TRUE 
parameter   integer PMA_CH2_REG_CDR_PROP_GAIN           = 2,            //
parameter   integer PMA_CH2_REG_CDR_PROP_TURBO_GAIN     = 6,            //
parameter   integer PMA_CH2_REG_CDR_INT_GAIN            = 2,            //
parameter   integer PMA_CH2_REG_CDR_INT_TURBO_GAIN      = 6,            //      
parameter   integer PMA_CH2_REG_CDR_INT_SAT_MAX         = 992,          //
parameter   integer PMA_CH2_REG_CDR_INT_SAT_MIN         = 32,           //
parameter           PMA_CH2_REG_CDR_INT_RST             = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high
parameter           PMA_CH2_REG_CDR_INT_RST_OW          = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH2_REG_CDR_PROP_RST            = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high 
parameter           PMA_CH2_REG_CDR_PROP_RST_OW         = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH2_REG_CDR_LOCK_RST            = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high 
parameter           PMA_CH2_REG_CDR_LOCK_RST_OW         = "DISABLE",     //DISABLE,ENABLE
parameter   integer PMA_CH2_REG_CDR_RX_PI_FORCE_SEL     = 0,             //
parameter   integer PMA_CH2_REG_CDR_RX_PI_FORCE_D       = 0,             //
parameter           PMA_CH2_REG_CDR_LOCK_TIMER          = "1_2U",        //"0_8U","1_2U","1_6U","2_4U","3_2U","4_8U","12_8U","25_6U"
parameter   integer PMA_CH2_REG_CDR_TURBO_MODE_TIMER    = 1,             //  
parameter           PMA_CH2_REG_CDR_LOCK_VAL            = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high 
parameter           PMA_CH2_REG_CDR_LOCK_OW             = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH2_REG_CDR_INT_SAT_DET_EN      = "TRUE",       //FALSE,TRUE
parameter           PMA_CH2_REG_CDR_SAT_DET_STATUS_EN   = "FALSE",       //FALSE,TRUE
parameter           PMA_CH2_REG_CDR_SAT_DET_STATUS_RESET_EN = "FALSE",       //FALSE,TRUE
parameter           PMA_CH2_REG_CDR_PI_CTRL_RST         = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high 
parameter           PMA_CH2_REG_CDR_PI_CTRL_RST_OW      = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH2_REG_CDR_SAT_DET_RST         = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high 
parameter           PMA_CH2_REG_CDR_SAT_DET_RST_OW      = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH2_REG_CDR_SAT_DET_STICKY_RST  = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high
parameter           PMA_CH2_REG_CDR_SAT_DET_STICKY_RST_OW = "DISABLE",   //DISABLE,ENABLE
parameter           PMA_CH2_REG_CDR_SIGDET_STATUS_DIS   = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high
parameter   integer PMA_CH2_REG_CDR_SAT_DET_TIMER       = 2,             //
parameter           PMA_CH2_REG_CDR_SAT_DET_STATUS_VAL  = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high
parameter           PMA_CH2_REG_CDR_SAT_DET_STATUS_OW   = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH2_REG_CDR_TURBO_MODE_EN       = "TRUE",       //FALSE,TRUE   
parameter   integer PMA_CH2_REG_CDR_STATUS_RADDR_INIT   = 0,             //
parameter           PMA_CH2_REG_CDR_STATUS_FIFO_EN      = "TRUE",       //FALSE,TRUE
parameter   integer PMA_CH2_REG_PMA_TEST_SEL            = 0,             //
parameter   integer PMA_CH2_REG_OOB_COMWAKE_GAP_MIN     = 3,             //
parameter   integer PMA_CH2_REG_OOB_COMWAKE_GAP_MAX     = 11,            //
parameter   integer PMA_CH2_REG_OOB_COMINIT_GAP_MIN     = 15,            //
parameter   integer PMA_CH2_REG_OOB_COMINIT_GAP_MAX     = 35,            //
parameter   integer PMA_CH2_REG_RX_PIBUF_IC_TX          = 1,             //
parameter   integer PMA_CH2_REG_COMWAKE_STATUS_CLEAR    = 0,             //
parameter   integer PMA_CH2_REG_COMINIT_STATUS_CLEAR    = 0,             //
parameter           PMA_CH2_REG_RX_SYNC_RST_N_EN        = "FALSE",       //FALSE,TRUE
parameter           PMA_CH2_REG_RX_SYNC_RST_N           = "TRUE",       //FALSE,TRUE  FALSE=low, TRUE=high           
parameter           PMA_CH2_REG_RX_SATA_COMINIT_OW      = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH2_REG_RX_SATA_COMINIT         = "FALSE",      //FALSE,TRUE FALSE=low, TRUE=high    
parameter           PMA_CH2_REG_RX_SATA_COMWAKE_OW      = "DISABLE",     //DISABLE,ENABLE      
parameter           PMA_CH2_REG_RX_SATA_COMWAKE         = "FALSE",      //FALSE,TRUE FALSE=low, TRUE=high          
parameter           PMA_CH2_REG_RX_DCC_DISABLE          = "ENABLE",     //DISABLE,ENABLE   
parameter           PMA_CH2_REG_TX_DCC_DISABLE          = "ENABLE",     //DISABLE,ENABLE  
parameter           PMA_CH2_REG_RX_SLIP_SEL_EN          = "FALSE",       //FALSE,TRUE 
parameter   integer PMA_CH2_REG_RX_SLIP_SEL             = 0,             //
parameter           PMA_CH2_REG_RX_SLIP_EN              = "FALSE",       //FALSE,TRUE
parameter   integer PMA_CH2_REG_RX_SIGDET_STATUS_SEL    = 5,             //
parameter           PMA_CH2_REG_RX_SIGDET_FSM_RST_N     = "TRUE",        //FALSE,TRUE  FALSE=low, TRUE=high     
parameter           PMA_CH2_REG_RX_SIGDET_STATUS_OW     = "DISABLE",     //DISABLE,ENABLE    
parameter           PMA_CH2_REG_RX_SIGDET_STATUS        = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high         
parameter           PMA_CH2_REG_RX_SIGDET_VTH           = "50MV",        //"12_5MV","25MV","37_5MV","50MV","62_5MV","75MV","87_5MV","100MV"
parameter   integer PMA_CH2_REG_RX_SIGDET_GRM           = 0,             // 
parameter           PMA_CH2_REG_RX_SIGDET_PULSE_EXT     = "DISABLE",     //DISABLE,ENABLE  
parameter   integer PMA_CH2_REG_RX_SIGDET_CH2_SEL       = 0,             // 
parameter   integer PMA_CH2_REG_RX_SIGDET_CH2_CHK_WINDOW =3,             //
parameter           PMA_CH2_REG_RX_SIGDET_CHK_WINDOW_EN = "TRUE",       //FALSE,TRUE
parameter   integer PMA_CH2_REG_RX_SIGDET_NOSIG_COUNT_SETTING = 4,       //
parameter   integer PMA_CH2_REG_RX_SIGDET_OOB_DET_COUNT_VAL= 0,             //
parameter           PMA_CH2_REG_SLIP_FIFO_INV_EN        = "FALSE",       //FALSE,TRUE
parameter           PMA_CH2_REG_SLIP_FIFO_INV           = "POS_EDGE",    //POS_EDGE,NEG_EDGE
parameter   integer PMA_CH2_REG_RX_SIGDET_4OOB_DET_SEL   =7,             //
////parameter   integer PMA_CH2_REG_RX_SIGDET_CHK_WINDOW    = 5,             //
////parameter   integer PMA_CH2_REG_RX_SIGDET_CHK_WINDOW_COUNT =3,             //
////parameter           PMA_CH2_REG_RX_SIGDET_LONG_CHK_WINDOW_EN = "DISABLE",  //DISABLE,ENABLE  
////parameter   integer PMA_CH2_REG_RX_SIGDET_LONG_CHK_WINDOW = 25,          //
parameter   integer PMA_CH2_REG_RX_SIGDET_IC_I          = 10,            //
parameter           PMA_CH2_REG_RX_OOB_DETECTOR_RESET_N_OW = "DISABLE",  //DISABLE,ENABLE
parameter           PMA_CH2_REG_RX_OOB_DETECTOR_RESET_N = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high  
parameter           PMA_CH2_REG_RX_OOB_DETECTOR_PD_OW   = "DISABLE",     //DISABLE,ENABLE  
parameter           PMA_CH2_REG_RX_OOB_DETECTOR_PD      = "ON",          //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_CH2_REG_RX_TERM_CM_CTRL         = "5DIV7",       //"5DIV7","2DIV3","5DIV6","4DIV5"
//PMA LANE Rx end   
//PMA LANE Tx begin 
parameter           PMA_CH2_REG_TX_PD                   = "ON",         //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_CH2_REG_TX_PD_OW                = "DISABLE",     //DISABLE,ENABLE       
parameter           PMA_CH2_REG_TX_CLKPATH_PD           = "ON",         //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_CH2_REG_TX_CLKPATH_PD_OW        = "DISABLE",     //DISABLE,ENABLE
parameter   integer PMA_CH2_REG_TX_BEACON_TIMER_SEL     = 0,            // 
parameter           PMA_CH2_REG_TX_RXDET_REQ_OW         = "DISABLE",    //DISABLE,ENABLE
parameter           PMA_CH2_REG_TX_RXDET_REQ            = "FALSE",      //FALSE,TRUE FALSE=low, TRUE=high
parameter           PMA_CH2_REG_TX_BEACON_EN_OW         = "DISABLE",     //DISABLE,ENABLE      
parameter           PMA_CH2_REG_TX_BEACON_EN            = "FALSE",      //FALSE,TRUE
parameter           PMA_CH2_REG_TX_EI_EN_OW             = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH2_REG_TX_EI_EN                = "FALSE",      //FALSE,TRUE
parameter           PMA_CH2_REG_TX_RES_CAL_EN           = "FALSE",      //FALSE,TRUE
parameter   integer PMA_CH2_REG_TX_RES_CAL              = 51,           // 
parameter           PMA_CH2_REG_TX_BIAS_CAL_EN          = "FALSE",      //FALSE,TRUE
parameter   integer PMA_CH2_REG_TX_BIAS_CTRL            = 48,           //
parameter           PMA_CH2_REG_TX_RXDET_TIMER_SEL      = "12CYCLE",     //"3CYCLE","12CYCLE","24CYCLE","36CYCLE"
parameter           PMA_CH2_REG_TX_SYNC_OW              = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH2_REG_TX_SYNC                 = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH2_REG_TX_PD_POST              = "OFF",        //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_CH2_REG_TX_PD_POST_OW           = "DISABLE",      //DISABLE,ENABLE
parameter           PMA_CH2_REG_TX_RESET_N_OW           = "DISABLE",     //DISABLE,ENABLE     
parameter           PMA_CH2_REG_TX_RESET_N              = "TRUE",       //FALSE,TRUE FALSE=low, TRUE=high 
parameter           PMA_CH2_REG_TX_DCC_RESET_N_OW       = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH2_REG_TX_DCC_RESET_N          = "TRUE",       //FALSE,TRUE FALSE=low, TRUE=high
parameter           PMA_CH2_REG_TX_BUSWIDTH_OW          = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH2_REG_TX_BUSWIDTH             = "20BIT",      //"8BIT","10BIT","16BIT","20BIT"
parameter           PMA_CH2_REG_PLL_READY_OW            = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH2_REG_PLL_READY               = "TRUE",       //FALSE,TRUE FALSE=low, TRUE=high 
parameter           PMA_CH2_REG_TX_PCLK_SW_OW           = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH2_REG_TX_PCLK_SW              = "TRUE",        //FALSE,TRUE FALSE=low, TRUE=high 
parameter   integer PMA_CH2_REG_EI_PCLK_DELAY_SEL       = 0,             //
parameter   integer PMA_CH2_REG_TX_DRV01_DAC0           = 0,             //
parameter   integer PMA_CH2_REG_TX_DRV01_DAC1           = 10,            //
parameter   integer PMA_CH2_REG_TX_DRV01_DAC2           = 16,            //
parameter   integer PMA_CH2_REG_TX_DRV00_DAC0           = 63,            //
parameter   integer PMA_CH2_REG_TX_DRV00_DAC1           = 53,            //
parameter   integer PMA_CH2_REG_TX_DRV00_DAC2           = 48,            //
parameter   integer PMA_CH2_REG_TX_AMP0                 = 8,             //
parameter   integer PMA_CH2_REG_TX_AMP1                 = 16,            //
parameter   integer PMA_CH2_REG_TX_AMP2                 = 32,            //
parameter   integer PMA_CH2_REG_TX_AMP3                 = 48,            //
parameter   integer PMA_CH2_REG_TX_AMP4                 = 56,            //
parameter   integer PMA_CH2_REG_TX_MARGIN               = 0,             // 
parameter           PMA_CH2_REG_TX_MARGIN_OW            = "DISABLE",     //DISABLE,ENABLE
parameter   integer PMA_CH2_REG_TX_DEEMP                = 0,             // 
parameter           PMA_CH2_REG_TX_DEEMP_OW             = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH2_REG_TX_SWING                = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high
parameter           PMA_CH2_REG_TX_SWING_OW             = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH2_REG_TX_RXDET_THRESHOLD      = "100MV",       //"50MV","75MV","100MV","125MV"
parameter   integer PMA_CH2_REG_TX_BEACON_OSC_CTRL      = 4,             //
parameter   integer PMA_CH2_REG_TX_PREDRV_DAC           = 1,             //
parameter   integer PMA_CH2_REG_TX_PREDRV_CM_CTRL       = 1,             //
parameter           PMA_CH2_REG_TX_TX2RX_SLPBACK_EN     = "FALSE",      //FALSE,TRUE
parameter           PMA_CH2_REG_TX_PCLK_EDGE_SEL        = "POS_EDGE",    //"NEG_EDGE","POS_EDGE"
parameter           PMA_CH2_REG_TX_RXDET_STATUS_OW      = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH2_REG_TX_RXDET_STATUS         = "TRUE",        //FALSE,TRUE FALSE=low, TRUE=high 
parameter           PMA_CH2_REG_TX_PRBS_GEN_EN          = "FALSE",      //FALSE,TRUE    
parameter           PMA_CH2_REG_TX_PRBS_GEN_WIDTH_SEL   = "20BIT",       //"8BIT","10BIT","16BIT","20BIT"
parameter           PMA_CH2_REG_TX_PRBS_SEL             = "PRBS7",       //"PRBS7","PRBS15","PRBS23","PRBS31"
parameter   integer PMA_CH2_REG_TX_UDP_DATA             = 256773,        //
parameter           PMA_CH2_REG_TX_FIFO_RST_N           = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high 
parameter   integer PMA_CH2_REG_TX_FIFO_WP_CTRL         = 2,             //
parameter           PMA_CH2_REG_TX_FIFO_EN              = "FALSE",      //FALSE,TRUE         
parameter   integer PMA_CH2_REG_TX_DATA_MUX_SEL         = 2,             //
parameter           PMA_CH2_REG_TX_ERR_INSERT           = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high 
parameter           PMA_CH2_REG_TX_SATA_EN              = "FALSE",       //FALSE,TRUE                  
parameter           PMA_CH2_REG_RATE_CHANGE_TXPCLK_ON_OW = "DISABLE",    //DISABLE,ENABLE 
parameter           PMA_CH2_REG_RATE_CHANGE_TXPCLK_ON   = "ENABLE",      //DISABLE,ENABLE 
parameter   integer PMA_CH2_REG_TX_PULLUP_DAC0          = 8,            //
parameter   integer PMA_CH2_REG_TX_PULLUP_DAC1          = 8,            //
parameter   integer PMA_CH2_REG_TX_PULLUP_DAC2          = 8,            //
parameter   integer PMA_CH2_REG_TX_PULLUP_DAC3          = 8,            //
parameter   integer PMA_CH2_REG_TX_OOB_DELAY_SEL        = 0,            //
parameter           PMA_CH2_REG_TX_POLARITY             = "NORMAL",      //"NORMAL","REVERSE"
parameter   integer PMA_CH2_REG_TX_SLPBK_AMP            = 1,             //
parameter           PMA_CH2_REG_TX_LS_MODE_EN           = "FALSE",       //FALSE,TRUE   
parameter           PMA_CH2_REG_TX_JTAG_MODE_EN_OW      = "DISABLE",     //DISABLE,ENABLE 
parameter           PMA_CH2_REG_TX_JTAG_MODE_EN         = "FALSE",       //FALSE,TRUE
parameter           PMA_CH2_REG_RX_JTAG_MODE_EN_OW      = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH2_REG_RX_JTAG_MODE_EN         = "FALSE",       //FALSE,TRUE
parameter           PMA_CH2_REG_RX_JTAG_OE              = "DISABLE",     //DISABLE,ENABLE 
parameter   integer PMA_CH2_REG_RX_ACJTAG_VHYSTSE       = 0,             //
parameter           PMA_CH2_REG_TX_FBCLK_FAR_EN         = "FALSE",       //FALSE,TRUE
parameter   integer PMA_CH2_REG_RX_TERM_MODE_CTRL       = 6,             //
parameter           PMA_CH2_REG_PLPBK_TXPCLK_EN         = "TRUE",        //FALSE,TRUE
//PMA LANE Tx end   
//PMA LANE CFG begin
parameter           PMA_CH2_CFG_LANE_POWERUP            = "OFF",         //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_CH2_CFG_PMA_POR_N               = "FALSE",      //FALSE,TRUE FALSE=low, TRUE=high    
parameter           PMA_CH2_CFG_RX_LANE_POWERUP         = "OFF",       //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_CH2_CFG_RX_PMA_RSTN             = "FALSE",      //FALSE,TRUE FALSE=low, TRUE=high   
parameter           PMA_CH2_CFG_TX_LANE_POWERUP         = "OFF",       //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_CH2_CFG_TX_PMA_RSTN             = "FALSE",      //FALSE,TRUE FALSE=low, TRUE=high
//PMA LANE CFG end  
////reserved reg    
parameter   integer PMA_CH2_REG_RESERVED_48_45          = 0,             //  
parameter   integer PMA_CH2_REG_RESERVED_69             = 0,             //
parameter   integer PMA_CH2_REG_RESERVED_77_76          = 0,             //
parameter   integer PMA_CH2_REG_RESERVED_171_164        = 0,             //
parameter   integer PMA_CH2_REG_RESERVED_175_172        = 0,             //
parameter   integer PMA_CH2_REG_RESERVED_190            = 0,             //
parameter   integer PMA_CH2_REG_RESERVED_233_232        = 0,             //
parameter   integer PMA_CH2_REG_RESERVED_235_234        = 0,             //
parameter   integer PMA_CH2_REG_RESERVED_241_240        = 0,             //
parameter   integer PMA_CH2_REG_RESERVED_285_283        = 0,             //
parameter   integer PMA_CH2_REG_RESERVED_286            = 0,             //
parameter   integer PMA_CH2_REG_RESERVED_295            = 0,             //
parameter   integer PMA_CH2_REG_RESERVED_298            = 0,             //
parameter   integer PMA_CH2_REG_RESERVED_332_325        = 0,             //
parameter   integer PMA_CH2_REG_RESERVED_340_333        = 0,             //
parameter   integer PMA_CH2_REG_RESERVED_348_341        = 0,             //
parameter   integer PMA_CH2_REG_RESERVED_354_349        = 0,             //
parameter   integer PMA_CH2_REG_RESERVED_373            = 0,             //
parameter   integer PMA_CH2_REG_RESERVED_376            = 0,             //
parameter   integer PMA_CH2_REG_RESERVED_452            = 0,             //
parameter   integer PMA_CH2_REG_RESERVED_502_499        = 0,             //
//parameter   integer PMA_CH2_REG_RESERVED_503            = 0,             // 
parameter   integer PMA_CH2_REG_RESERVED_506_505        = 0,             //
parameter   integer PMA_CH2_REG_RESERVED_550_549        = 0,             //
parameter   integer PMA_CH2_REG_RESERVED_556_552        = 0,             //
////reserved end    
//PMA LANE2 end     
                    
//PMA LANE3 begin   
//PMA LANE Rx begin 
parameter           PMA_CH3_REG_RX_PD                   = "ON",         //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_CH3_REG_RX_PD_EN                = "FALSE",      //FALSE,TRUE  
parameter           PMA_CH3_REG_RX_CLKPATH_PD           = "ON",         //ON,OFF   ON=poweron,OFF= powerdown,reserved
parameter           PMA_CH3_REG_RX_CLKPATH_PD_EN        = "FALSE",      //FALSE,TRUE  ,reserved
parameter           PMA_CH3_REG_RX_DATAPATH_PD          = "ON",         //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_CH3_REG_RX_DATAPATH_PD_EN       = "FALSE",      //FALSE,TRUE
parameter           PMA_CH3_REG_RX_SIGDET_PD            = "ON",         //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_CH3_REG_RX_SIGDET_PD_EN         = "FALSE",      //FALSE,TRUE
parameter           PMA_CH3_REG_RX_DCC_RST_N            = "TRUE",       //FALSE,TRUE  FALSE=low, TRUE=high
parameter           PMA_CH3_REG_RX_DCC_RST_N_EN         = "FALSE",       //FALSE,TRUE
parameter           PMA_CH3_REG_RX_CDR_RST_N            = "TRUE",       //FALSE,TRUE  FALSE=low, TRUE=high
parameter           PMA_CH3_REG_RX_CDR_RST_N_EN         = "FALSE",       //FALSE,TRUE
parameter           PMA_CH3_REG_RX_SIGDET_RST_N         = "TRUE",       //FALSE,TRUE  FALSE=low, TRUE=high
parameter           PMA_CH3_REG_RX_SIGDET_RST_N_EN      = "FALSE",       //FALSE,TRUE
parameter           PMA_CH3_REG_RXPCLK_SLIP             = "FALSE",      //FALSE,TRUE
parameter           PMA_CH3_REG_RXPCLK_SLIP_OW          = "DISABLE",    //DISABLE,ENABLE
parameter           PMA_CH3_REG_RX_PCLKSWITCH_RST_N     = "TRUE",       //FALSE,TRUE  FALSE=low, TRUE=high
parameter           PMA_CH3_REG_RX_PCLKSWITCH_RST_N_EN  = "FALSE",       //FALSE,TRUE
parameter           PMA_CH3_REG_RX_PCLKSWITCH           = "FALSE",      //FALSE,TRUE
parameter           PMA_CH3_REG_RX_PCLKSWITCH_EN        = "FALSE",       //FALSE,TRUE
parameter           PMA_CH3_REG_RX_HIGHZ                = "FALSE",      //FALSE,TRUE
parameter           PMA_CH3_REG_RX_HIGHZ_EN             = "FALSE",       //FALSE,TRUE
parameter   integer PMA_CH3_REG_RX_EQ_C_SET             = 8,            // 
parameter   integer PMA_CH3_REG_RX_EQ_R_SET             = 8,            // 
parameter           PMA_CH3_REG_RX_BUSWIDTH             = "20BIT",       //"8BIT","10BIT","16BIT","20BIT" 
parameter           PMA_CH3_REG_RX_BUSWIDTH_EN          = "FALSE",       //FALSE,TRUE
parameter           PMA_CH3_REG_RX_RATE                 = "DIV1",       //"DIV8","DIV4","DIV2","DIV1"           
parameter           PMA_CH3_REG_RX_RATE_EN              = "FALSE",       //FALSE,TRUE
parameter   integer PMA_CH3_REG_RX_RES_TRIM             = 51,           //
parameter           PMA_CH3_REG_RX_RES_TRIM_EN          = "FALSE",       //FALSE,TRUE
parameter           PMA_CH3_REG_RX_EQ_OFF               = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high
parameter   integer PMA_CH3_REG_RX_PREAMP_IC            = 1367,          //
parameter           PMA_CH3_REG_RX_PCLK_EDGE_SEL        = "POS_EDGE",    //"POS_EDGE","NEG_EDGE"
parameter   integer PMA_CH3_REG_RX_PIBUF_IC             = 2,             //
parameter   integer PMA_CH3_REG_RX_DCC_IC_RX            = 3,             //
parameter   integer PMA_CH3_REG_RX_DCC_IC_TX            = 3,             //
parameter           PMA_CH3_REG_RX_ICTRL_TRX            = "100PCT",      //"87_5PCT","100PCT","112_5PCT","125PCT" 
////parameter           PMA_CH3_REG_RX_ICTRL_SIGDET         = "100PCT",      //"87_5PCT","100PCT","112_5PCT","125PCT"  
parameter   integer PMA_CH3_REG_RX_ICTRL_SIGDET         = 5,
parameter           PMA_CH3_REG_RX_ICTRL_PREAMP         = "100PCT",      //"87_5PCT","100PCT","112_5PCT","125PCT"  
parameter           PMA_CH3_REG_RX_ICTRL_SLICER         = "100PCT",      //"87_5PCT","100PCT","112_5PCT","125PCT"  
parameter           PMA_CH3_REG_RX_ICTRL_PIBUF          = "100PCT",      //"87_5PCT","100PCT","112_5PCT","125PCT" 
parameter           PMA_CH3_REG_RX_ICTRL_PI             = "100PCT",      //"87_5PCT","100PCT","112_5PCT","125PCT" 
parameter           PMA_CH3_REG_RX_ICTRL_DCC            = "100PCT",      //"87_5PCT","100PCT","112_5PCT","125PCT"
parameter           PMA_CH3_REG_RX_ICTRL_PREDRV         = "100PCT",      //"87_5PCT","100PCT","112_5PCT","125PCT"
parameter           PMA_CH3_REG_TX_RATE                 = "DIV1",        //"DIV8","DIV4","DIV2","DIV1"  
parameter           PMA_CH3_REG_TX_RATE_EN              = "FALSE",       //FALSE,TRUE
parameter           PMA_CH3_REG_RX_TX2RX_PLPBK_RST_N    = "TRUE",       //FALSE,TRUE  FALSE=low, TRUE=high
parameter           PMA_CH3_REG_RX_TX2RX_PLPBK_RST_N_EN = "FALSE",       //FALSE,TRUE
parameter           PMA_CH3_REG_RX_TX2RX_PLPBK_EN       = "FALSE",       //FALSE,TRUE
parameter           PMA_CH3_REG_TXCLK_SEL               = "PLL",        //"PLL","RXCLK"
parameter           PMA_CH3_REG_RX_DATA_POLARITY        = "NORMAL",     //"NORMAL","REVERSE"
parameter           PMA_CH3_REG_RX_ERR_INSERT           = "FALSE",      //FALSE,TRUE FALSE=low, TRUE=high
parameter           PMA_CH3_REG_UDP_CHK_EN              = "FALSE",       //FALSE,TRUE
parameter           PMA_CH3_REG_PRBS_SEL                = "PRBS7",      //"PRBS7","PRBS15","PRBS23","PRBS31"
parameter           PMA_CH3_REG_PRBS_CHK_EN             = "FALSE",       //FALSE,TRUE
parameter           PMA_CH3_REG_PRBS_CHK_WIDTH_SEL      = "20BIT",      //"8BIT","10BIT","16BIT","20BIT"
parameter           PMA_CH3_REG_BIST_CHK_PAT_SEL        = "PRBS",       //"PRBS","CONSTANT"
parameter           PMA_CH3_REG_LOAD_ERR_CNT            = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH3_REG_CHK_COUNTER_EN          = "FALSE",       //FALSE,TRUE 
parameter   integer PMA_CH3_REG_CDR_PROP_GAIN           = 2,             //
parameter   integer PMA_CH3_REG_CDR_PROP_TURBO_GAIN     = 6,             //
parameter   integer PMA_CH3_REG_CDR_INT_GAIN            = 2,             //
parameter   integer PMA_CH3_REG_CDR_INT_TURBO_GAIN      = 6,             //      
parameter   integer PMA_CH3_REG_CDR_INT_SAT_MAX         = 992,          //
parameter   integer PMA_CH3_REG_CDR_INT_SAT_MIN         = 32,            //
parameter           PMA_CH3_REG_CDR_INT_RST             = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high
parameter           PMA_CH3_REG_CDR_INT_RST_OW          = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH3_REG_CDR_PROP_RST            = "FALSE",      //FALSE,TRUE FALSE=low, TRUE=high 
parameter           PMA_CH3_REG_CDR_PROP_RST_OW         = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH3_REG_CDR_LOCK_RST            = "FALSE",      //FALSE,TRUE FALSE=low, TRUE=high 
parameter           PMA_CH3_REG_CDR_LOCK_RST_OW         = "DISABLE",    //DISABLE,ENABLE
parameter   integer PMA_CH3_REG_CDR_RX_PI_FORCE_SEL     = 0,             //
parameter   integer PMA_CH3_REG_CDR_RX_PI_FORCE_D       = 0,             //
parameter           PMA_CH3_REG_CDR_LOCK_TIMER          = "1_2U",        //"0_8U","1_2U","1_6U","2_4U","3_2U","4_8U","12_8U","25_6U"
parameter   integer PMA_CH3_REG_CDR_TURBO_MODE_TIMER    = 1,             //  
parameter           PMA_CH3_REG_CDR_LOCK_VAL            = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high 
parameter           PMA_CH3_REG_CDR_LOCK_OW             = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH3_REG_CDR_INT_SAT_DET_EN      = "TRUE",       //FALSE,TRUE
parameter           PMA_CH3_REG_CDR_SAT_DET_STATUS_EN   = "FALSE",       //FALSE,TRUE
parameter           PMA_CH3_REG_CDR_SAT_DET_STATUS_RESET_EN = "FALSE",       //FALSE,TRUE
parameter           PMA_CH3_REG_CDR_PI_CTRL_RST         = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high 
parameter           PMA_CH3_REG_CDR_PI_CTRL_RST_OW      = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH3_REG_CDR_SAT_DET_RST         = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high 
parameter           PMA_CH3_REG_CDR_SAT_DET_RST_OW      = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH3_REG_CDR_SAT_DET_STICKY_RST  = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high
parameter           PMA_CH3_REG_CDR_SAT_DET_STICKY_RST_OW = "DISABLE",   //DISABLE,ENABLE
parameter           PMA_CH3_REG_CDR_SIGDET_STATUS_DIS   = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high
parameter   integer PMA_CH3_REG_CDR_SAT_DET_TIMER       = 2,             //
parameter           PMA_CH3_REG_CDR_SAT_DET_STATUS_VAL  = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high
parameter           PMA_CH3_REG_CDR_SAT_DET_STATUS_OW   = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH3_REG_CDR_TURBO_MODE_EN       = "TRUE",       //FALSE,TRUE   
parameter   integer PMA_CH3_REG_CDR_STATUS_RADDR_INIT   = 0,             //
parameter           PMA_CH3_REG_CDR_STATUS_FIFO_EN      = "TRUE",       //FALSE,TRUE
parameter   integer PMA_CH3_REG_PMA_TEST_SEL            = 0,             //
parameter   integer PMA_CH3_REG_OOB_COMWAKE_GAP_MIN     = 3,             //
parameter   integer PMA_CH3_REG_OOB_COMWAKE_GAP_MAX     = 11,            //
parameter   integer PMA_CH3_REG_OOB_COMINIT_GAP_MIN     = 15,            //
parameter   integer PMA_CH3_REG_OOB_COMINIT_GAP_MAX     = 35,            //
parameter   integer PMA_CH3_REG_RX_PIBUF_IC_TX          = 1,             //
parameter   integer PMA_CH3_REG_COMWAKE_STATUS_CLEAR    = 0,             //
parameter   integer PMA_CH3_REG_COMINIT_STATUS_CLEAR    = 0,             //
parameter           PMA_CH3_REG_RX_SYNC_RST_N_EN        = "FALSE",       //FALSE,TRUE
parameter           PMA_CH3_REG_RX_SYNC_RST_N           = "TRUE",       //FALSE,TRUE  FALSE=low, TRUE=high           
parameter           PMA_CH3_REG_RX_SATA_COMINIT_OW      = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH3_REG_RX_SATA_COMINIT         = "FALSE",      //FALSE,TRUE FALSE=low, TRUE=high    
parameter           PMA_CH3_REG_RX_SATA_COMWAKE_OW      = "DISABLE",     //DISABLE,ENABLE      
parameter           PMA_CH3_REG_RX_SATA_COMWAKE         = "FALSE",      //FALSE,TRUE FALSE=low, TRUE=high          
parameter           PMA_CH3_REG_RX_DCC_DISABLE          = "ENABLE",     //DISABLE,ENABLE   
parameter           PMA_CH3_REG_TX_DCC_DISABLE          = "ENABLE",     //DISABLE,ENABLE  
parameter           PMA_CH3_REG_RX_SLIP_SEL_EN          = "FALSE",       //FALSE,TRUE 
parameter   integer PMA_CH3_REG_RX_SLIP_SEL             = 0,             //
parameter           PMA_CH3_REG_RX_SLIP_EN              = "FALSE",       //FALSE,TRUE 
parameter   integer PMA_CH3_REG_RX_SIGDET_STATUS_SEL    = 5,             //
parameter           PMA_CH3_REG_RX_SIGDET_FSM_RST_N     = "TRUE",        //FALSE,TRUE  FALSE=low, TRUE=high     
parameter           PMA_CH3_REG_RX_SIGDET_STATUS_OW     = "DISABLE",     //DISABLE,ENABLE    
parameter           PMA_CH3_REG_RX_SIGDET_STATUS        = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high         
parameter           PMA_CH3_REG_RX_SIGDET_VTH           = "50MV",        //"12_5MV","25MV","37_5MV","50MV","62_5MV","75MV","87_5MV","100MV"
parameter   integer PMA_CH3_REG_RX_SIGDET_GRM           = 0,             // 
parameter           PMA_CH3_REG_RX_SIGDET_PULSE_EXT     = "DISABLE",     //DISABLE,ENABLE  
parameter   integer PMA_CH3_REG_RX_SIGDET_CH2_SEL       = 0,             // 
parameter   integer PMA_CH3_REG_RX_SIGDET_CH2_CHK_WINDOW =3,             //
parameter           PMA_CH3_REG_RX_SIGDET_CHK_WINDOW_EN = "TRUE",       //FALSE,TRUE
parameter   integer PMA_CH3_REG_RX_SIGDET_NOSIG_COUNT_SETTING = 4,       //
parameter   integer PMA_CH3_REG_RX_SIGDET_OOB_DET_COUNT_VAL= 0,             //
parameter           PMA_CH3_REG_SLIP_FIFO_INV_EN        = "FALSE",       //FALSE,TRUE
parameter           PMA_CH3_REG_SLIP_FIFO_INV           = "POS_EDGE",    //POS_EDGE,NEG_EDGE
parameter   integer PMA_CH3_REG_RX_SIGDET_4OOB_DET_SEL   =7,             //
////parameter   integer PMA_CH3_REG_RX_SIGDET_CHK_WINDOW    = 5,             //
////parameter   integer PMA_CH3_REG_RX_SIGDET_CHK_WINDOW_COUNT =3,             //
////parameter          PMA_CH3_REG_RX_SIGDET_LONG_CHK_WINDOW_EN = "DISABLE",  //DISABLE,ENABLE  
////parameter   integer PMA_CH3_REG_RX_SIGDET_LONG_CHK_WINDOW = 25,          //
parameter   integer PMA_CH3_REG_RX_SIGDET_IC_I          = 10,            //
parameter           PMA_CH3_REG_RX_OOB_DETECTOR_RESET_N_OW = "DISABLE",  //DISABLE,ENABLE
parameter           PMA_CH3_REG_RX_OOB_DETECTOR_RESET_N = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high  
parameter           PMA_CH3_REG_RX_OOB_DETECTOR_PD_OW   = "DISABLE",     //DISABLE,ENABLE  
parameter           PMA_CH3_REG_RX_OOB_DETECTOR_PD      = "ON",          //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_CH3_REG_RX_TERM_CM_CTRL         = "5DIV7",       //"5DIV7","2DIV3","5DIV6","4DIV5"
//PMA LANE Rx end   
//PMA LANE Tx begin  
parameter           PMA_CH3_REG_TX_PD                   = "ON",          //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_CH3_REG_TX_PD_OW                = "DISABLE",     //DISABLE,ENABLE       
parameter           PMA_CH3_REG_TX_CLKPATH_PD           = "ON",         //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_CH3_REG_TX_CLKPATH_PD_OW        = "DISABLE",     //DISABLE,ENABLE
parameter   integer PMA_CH3_REG_TX_BEACON_TIMER_SEL     = 0,            // 
parameter           PMA_CH3_REG_TX_RXDET_REQ_OW         = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH3_REG_TX_RXDET_REQ            = "FALSE",      //FALSE,TRUE FALSE=low, TRUE=high
parameter           PMA_CH3_REG_TX_BEACON_EN_OW         = "DISABLE",     //DISABLE,ENABLE         
parameter           PMA_CH3_REG_TX_BEACON_EN            = "FALSE",      //FALSE,TRUE
parameter           PMA_CH3_REG_TX_EI_EN_OW             = "DISABLE",    //DISABLE,ENABLE
parameter           PMA_CH3_REG_TX_EI_EN                = "FALSE",      //FALSE,TRUE
parameter           PMA_CH3_REG_TX_RES_CAL_EN           = "FALSE",      //FALSE,TRUE
parameter   integer PMA_CH3_REG_TX_RES_CAL              = 51,           // 
parameter           PMA_CH3_REG_TX_BIAS_CAL_EN          = "FALSE",      //FALSE,TRUE
parameter   integer PMA_CH3_REG_TX_BIAS_CTRL            = 48,           //
parameter           PMA_CH3_REG_TX_RXDET_TIMER_SEL      = "12CYCLE",    //"3CYCLE","12CYCLE","24CYCLE","36CYCLE"
parameter           PMA_CH3_REG_TX_SYNC_OW              = "DISABLE",    //DISABLE,ENABLE
parameter           PMA_CH3_REG_TX_SYNC                 = "DISABLE",    //DISABLE,ENABLE
parameter           PMA_CH3_REG_TX_PD_POST              = "OFF",        //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_CH3_REG_TX_PD_POST_OW           = "DISABLE",      //DISABLE,ENABLE
parameter           PMA_CH3_REG_TX_RESET_N_OW           = "DISABLE",     //DISABLE,ENABLE     
parameter           PMA_CH3_REG_TX_RESET_N              = "TRUE",       //FALSE,TRUE FALSE=low, TRUE=high 
parameter           PMA_CH3_REG_TX_DCC_RESET_N_OW       = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH3_REG_TX_DCC_RESET_N          = "TRUE",       //FALSE,TRUE FALSE=low, TRUE=high
parameter           PMA_CH3_REG_TX_BUSWIDTH_OW          = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH3_REG_TX_BUSWIDTH             = "20BIT",      //"8BIT","10BIT","16BIT","20BIT"
parameter           PMA_CH3_REG_PLL_READY_OW            = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH3_REG_PLL_READY               = "TRUE",       //FALSE,TRUE FALSE=low, TRUE=high 
parameter           PMA_CH3_REG_TX_PCLK_SW_OW           = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH3_REG_TX_PCLK_SW              = "TRUE",        //FALSE,TRUE FALSE=low, TRUE=high 
parameter   integer PMA_CH3_REG_EI_PCLK_DELAY_SEL       = 0,             //
parameter   integer PMA_CH3_REG_TX_DRV01_DAC0           = 0,             //
parameter   integer PMA_CH3_REG_TX_DRV01_DAC1           = 10,            //
parameter   integer PMA_CH3_REG_TX_DRV01_DAC2           = 16,            //
parameter   integer PMA_CH3_REG_TX_DRV00_DAC0           = 63,            //
parameter   integer PMA_CH3_REG_TX_DRV00_DAC1           = 53,            //
parameter   integer PMA_CH3_REG_TX_DRV00_DAC2           = 48,            //
parameter   integer PMA_CH3_REG_TX_AMP0                 = 8,             //
parameter   integer PMA_CH3_REG_TX_AMP1                 = 16,            //
parameter   integer PMA_CH3_REG_TX_AMP2                 = 32,            //
parameter   integer PMA_CH3_REG_TX_AMP3                 = 48,            //
parameter   integer PMA_CH3_REG_TX_AMP4                 = 56,            //
parameter   integer PMA_CH3_REG_TX_MARGIN               = 0,             // 
parameter           PMA_CH3_REG_TX_MARGIN_OW            = "DISABLE",     //DISABLE,ENABLE
parameter   integer PMA_CH3_REG_TX_DEEMP                = 0,             // 
parameter           PMA_CH3_REG_TX_DEEMP_OW             = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH3_REG_TX_SWING                = "FALSE",      //FALSE,TRUE FALSE=low, TRUE=high
parameter           PMA_CH3_REG_TX_SWING_OW             = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH3_REG_TX_RXDET_THRESHOLD      = "100MV",       //"50MV","75MV","100MV","125MV"
parameter   integer PMA_CH3_REG_TX_BEACON_OSC_CTRL      = 4,             //
parameter   integer PMA_CH3_REG_TX_PREDRV_DAC           = 1,             //
parameter   integer PMA_CH3_REG_TX_PREDRV_CM_CTRL       = 1,             //
parameter           PMA_CH3_REG_TX_TX2RX_SLPBACK_EN     = "FALSE",      //FALSE,TRUE
parameter           PMA_CH3_REG_TX_PCLK_EDGE_SEL        = "POS_EDGE",    //"NEG_EDGE","POS_EDGE"
parameter           PMA_CH3_REG_TX_RXDET_STATUS_OW      = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH3_REG_TX_RXDET_STATUS         = "TRUE",        //FALSE,TRUE FALSE=low, TRUE=high 
parameter           PMA_CH3_REG_TX_PRBS_GEN_EN          = "FALSE",      //FALSE,TRUE     
parameter           PMA_CH3_REG_TX_PRBS_GEN_WIDTH_SEL   = "20BIT",       //"8BIT","10BIT","16BIT","20BIT"
parameter           PMA_CH3_REG_TX_PRBS_SEL             = "PRBS7",       //"PRBS7","PRBS15","PRBS23","PRBS31"
parameter   integer PMA_CH3_REG_TX_UDP_DATA             = 256773,        //
parameter           PMA_CH3_REG_TX_FIFO_RST_N           = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high 
parameter   integer PMA_CH3_REG_TX_FIFO_WP_CTRL         = 2,             //
parameter           PMA_CH3_REG_TX_FIFO_EN              = "FALSE",      //FALSE,TRUE         
parameter   integer PMA_CH3_REG_TX_DATA_MUX_SEL         = 2,             //
parameter           PMA_CH3_REG_TX_ERR_INSERT           = "FALSE",       //FALSE,TRUE FALSE=low, TRUE=high 
parameter           PMA_CH3_REG_TX_SATA_EN              = "FALSE",       //FALSE,TRUE                   
parameter           PMA_CH3_REG_RATE_CHANGE_TXPCLK_ON_OW = "DISABLE",    //DISABLE,ENABLE 
parameter           PMA_CH3_REG_RATE_CHANGE_TXPCLK_ON   = "ENABLE",      //DISABLE,ENABLE 
parameter   integer PMA_CH3_REG_TX_PULLUP_DAC0          = 8,            //
parameter   integer PMA_CH3_REG_TX_PULLUP_DAC1          = 8,            //
parameter   integer PMA_CH3_REG_TX_PULLUP_DAC2          = 8,            //
parameter   integer PMA_CH3_REG_TX_PULLUP_DAC3          = 8,            //
parameter   integer PMA_CH3_REG_TX_OOB_DELAY_SEL        = 0,            //
parameter           PMA_CH3_REG_TX_POLARITY             = "NORMAL",      //"NORMAL","REVERSE"
parameter   integer PMA_CH3_REG_TX_SLPBK_AMP            = 1,             //
parameter           PMA_CH3_REG_TX_LS_MODE_EN           = "FALSE",       //FALSE,TRUE   
parameter           PMA_CH3_REG_TX_JTAG_MODE_EN_OW      = "DISABLE",     //DISABLE,ENABLE 
parameter           PMA_CH3_REG_TX_JTAG_MODE_EN         = "FALSE",       //FALSE,TRUE
parameter           PMA_CH3_REG_RX_JTAG_MODE_EN_OW      = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_CH3_REG_RX_JTAG_MODE_EN         = "FALSE",       //FALSE,TRUE
parameter           PMA_CH3_REG_RX_JTAG_OE              = "DISABLE",     //DISABLE,ENABLE 
parameter   integer PMA_CH3_REG_RX_ACJTAG_VHYSTSE       = 0,             //
parameter           PMA_CH3_REG_TX_FBCLK_FAR_EN         = "FALSE",       //FALSE,TRUE
parameter   integer PMA_CH3_REG_RX_TERM_MODE_CTRL       = 6,             //
parameter           PMA_CH3_REG_PLPBK_TXPCLK_EN         = "TRUE",        //FALSE,TRUE
//PMA LANE Tx end   
//PMA LANE CFG begin
parameter           PMA_CH3_CFG_LANE_POWERUP            = "OFF",         //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_CH3_CFG_PMA_POR_N               = "FALSE",      //FALSE,TRUE FALSE=low, TRUE=high    
parameter           PMA_CH3_CFG_RX_LANE_POWERUP         = "OFF",       //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_CH3_CFG_RX_PMA_RSTN             = "FALSE",      //FALSE,TRUE FALSE=low, TRUE=high   
parameter           PMA_CH3_CFG_TX_LANE_POWERUP         = "OFF",       //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_CH3_CFG_TX_PMA_RSTN             = "FALSE",      //FALSE,TRUE FALSE=low, TRUE=high
//PMA LANE CFG end  
////reserved reg    
parameter   integer PMA_CH3_REG_RESERVED_48_45          = 0,             //  
parameter   integer PMA_CH3_REG_RESERVED_69             = 0,             //
parameter   integer PMA_CH3_REG_RESERVED_77_76          = 0,             //
parameter   integer PMA_CH3_REG_RESERVED_171_164        = 0,             //
parameter   integer PMA_CH3_REG_RESERVED_175_172        = 0,             //
parameter   integer PMA_CH3_REG_RESERVED_190            = 0,             //
parameter   integer PMA_CH3_REG_RESERVED_233_232        = 0,             //
parameter   integer PMA_CH3_REG_RESERVED_235_234        = 0,             //
parameter   integer PMA_CH3_REG_RESERVED_241_240        = 0,             //
parameter   integer PMA_CH3_REG_RESERVED_285_283        = 0,             //
parameter   integer PMA_CH3_REG_RESERVED_286            = 0,             //
parameter   integer PMA_CH3_REG_RESERVED_295            = 0,             //
parameter   integer PMA_CH3_REG_RESERVED_298            = 0,             //
parameter   integer PMA_CH3_REG_RESERVED_332_325        = 0,             //
parameter   integer PMA_CH3_REG_RESERVED_340_333        = 0,             //
parameter   integer PMA_CH3_REG_RESERVED_348_341        = 0,             //
parameter   integer PMA_CH3_REG_RESERVED_354_349        = 0,             //
parameter   integer PMA_CH3_REG_RESERVED_373            = 0,             //
parameter   integer PMA_CH3_REG_RESERVED_376            = 0,             //
parameter   integer PMA_CH3_REG_RESERVED_452            = 0,             //
parameter   integer PMA_CH3_REG_RESERVED_502_499        = 0,             //
//parameter   integer PMA_CH3_REG_RESERVED_503            = 0,             // 
parameter   integer PMA_CH3_REG_RESERVED_506_505        = 0,             //
parameter   integer PMA_CH3_REG_RESERVED_550_549        = 0,             //
parameter   integer PMA_CH3_REG_RESERVED_556_552        = 0,             //
////reserved end    
//PMA LANE3 end     
                    
//PMA PLL begin     
parameter           PMA_PLL0_REG_PLL_POWERDOWN_OW       = "DISABLE",     //DISABLE,ENABLE  enable REG_PLL_POWERDOWN
parameter           PMA_PLL0_REG_PLL_POWERDOWN          = "ON",         //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_PLL0_REG_PLL_RESET_N_OW         = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_PLL0_REG_PLL_RESET_N            = "TRUE",       //FALSE,TRUE  FALSE=low, TRUE=high
parameter           PMA_PLL0_REG_PLL_READY_OW           = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_PLL0_REG_PLL_READY              = "FALSE",      //FALSE,TRUE
parameter           PMA_PLL0_REG_LANE_SYNC_OW           = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_PLL0_REG_LANE_SYNC              = "FALSE",       //FALSE,TRUE
////parameter           PMA_PLL0_REG_RESCAL_ENABLE_OW      = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_PLL0_REG_LOCKDET_REPEAT         = "DISABLE",    //DISABLE,ENABLE
////parameter           PMA_PLL0_REG_RESCAL_ENABLE         = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_PLL0_REG_RESCAL_I_CODE_PMA      = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_PLL0_REG_RESCAL_RESET_N_OW      = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_PLL0_REG_RESCAL_RESET_N         = "FALSE",       //FALSE,TRUE  FALSE=low, TRUE=high
parameter           PMA_PLL0_REG_RESCAL_DONE_OW         = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_PLL0_REG_RESCAL_DONE            = "FALSE",      //FALSE,TRUE
parameter           PMA_PLL0_REG_RESCAL_CODE_OW         = "DISABLE",     //DISABLE,ENABLE
////parameter   integer PMA_PLL0_REG_RESCAL_I_OFFSET       = 1,             // 
parameter   integer PMA_PLL0_REG_LDO_VREF_SEL           = 2,
parameter   integer PMA_PLL0_REG_BIAS_VCOREP_C          = 1,
////parameter   integer PMA_PLL0_REG_RESCAL_R_OFFSET       = 14,            // 
parameter   integer PMA_PLL0_REG_RESCAL_I_CODE          = 32,
parameter           PMA_PLL0_REG_RESCAL_ONCHIP_SMALL_OW = "DISABLE",     //DISABLE,ENABLE
parameter   integer PMA_PLL0_REG_RESCAL_ONCHIP_SMALL    = 0,             // 
////parameter   integer PMA_PLL0_REG_RESCAL_ITER           = 0,             // 
parameter           PMA_PLL0_REG_JTAG_OE                = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_PLL0_REG_JTAG_AC_MODE           = "DISABLE",     //DISABLE,ENABLE
////parameter           PMA_PLL0_REG_RESCAL_REPEAT_EN      = "DISABLE";     //DISABLE,ENABLE
////parameter   integer PMA_PLL0_REG_RESCAL_TIMEOUT        = 0,             // 
parameter   integer PMA_PLL0_REG_JTAG_VHYSTSEL          = 0,
parameter           PMA_PLL0_REG_PLL_LOCKDET_EN_OW      = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_PLL0_REG_PLL_LOCKDET_EN         = "FALSE",       //FALSE,TRUE
parameter           PMA_PLL0_REG_PLL_LOCKDET_RESET_N_OW = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_PLL0_REG_PLL_LOCKDET_RESET_N    = "FALSE",       //FALSE,TRUE  FALSE=low, TRUE=high
parameter           PMA_PLL0_REG_PLL_LOCKED_OW          = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_PLL0_REG_PLL_LOCKED             = "FALSE",       //FALSE,TRUE
parameter           PMA_PLL0_REG_PLL_LOCKED_STICKY_CLEAR = "FALSE",       //FALSE,TRUE
parameter           PMA_PLL0_REG_PLL_UNLOCKED_STICKY_CLEAR = "FALSE",      //FALSE,TRUE
parameter           PMA_PLL0_REG_NOFBCLK_STICKY_CLEAR   = "FALSE",       //FALSE,TRUE
parameter   integer PMA_PLL0_REG_PLL_LOCKDET_REFCT      = 7,             // 
parameter   integer PMA_PLL0_REG_PLL_LOCKDET_FBCT       = 7,             // 
parameter   integer PMA_PLL0_REG_PLL_LOCKDET_LOCKCT     = 4,             // 
parameter   integer PMA_PLL0_REG_PLL_LOCKDET_ITER       = 3,             // 
parameter   integer PMA_PLL0_REG_PLL_UNLOCKDET_ITER     = 2,             //
parameter           PMA_PLL0_REG_PD_VCO                 = "ON",          //ON,OFF   ON=poweron,OFF= powerdown   
parameter           PMA_PLL0_REG_FBCLK_TEST_EN          = "FALSE",       //FALSE,TRUE
parameter           PMA_PLL0_REG_REFCLK_TEST_EN         = "FALSE",       //FALSE,TRUE
parameter   integer PMA_PLL0_REG_TEST_SEL               = 0,             // 
parameter           PMA_PLL0_REG_TEST_V_EN              = "FALSE",       //FALSE,TRUE
parameter           PMA_PLL0_REG_TEST_SIG_HALF_EN       = "FALSE",       //FALSE,TRUE
parameter   integer PMA_PLL0_REG_TEST_FSM               = 0,             // 
parameter           PMA_PLL0_REG_REFCLK_OUT_PD          = "OFF",         //ON,OFF   ON=poweron,OFF= powerdown 
parameter           PMA_PLL0_REG_BGR_STARTUP_EN         = "FALSE",       //FALSE,TRUE
parameter           PMA_PLL0_REG_BGR_STARTUP            = "FALSE",       //FALSE,TRUE
parameter           PMA_PLL0_REG_PD_BGR                 = "ON",          //ON,OFF   ON=poweron,OFF= powerdown  
parameter           PMA_PLL0_REG_REFCLK_TERM_VCM_EN     = "TRUE",        //FALSE,TRUE
parameter           PMA_PLL0_REG_FBDIVA_5_EN            = "TRUE",        //FALSE,TRUE
parameter   integer PMA_PLL0_REG_FBDIVB                 = 1,             //  
parameter           PMA_PLL0_REG_RESET_N_PFDQP_OW       = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_PLL0_REG_RESET_N_PFDQP          = "FALSE",       //FALSE,TRUE  FALSE=low, TRUE=high
parameter   integer PMA_PLL0_REG_QPCURRENT              = 12,            //  
parameter           PMA_PLL0_REG_VC_FORCE_EN            = "FALSE",       //FALSE,TRUE
parameter   integer PMA_PLL0_REG_VCRESET_C_RING         = 24,            //  
parameter   integer PMA_PLL0_REG_LPF_R_C                = 0,             // 
parameter   integer PMA_PLL0_REG_LPF_TR_C               = 2,             //
parameter           PMA_PLL0_REG_PD_BIAS                = "ON",          //ON,OFF   ON=poweron,OFF= powerdown  
parameter   integer PMA_PLL0_REG_ICTRL_PLL              = 1,            //  
parameter   integer PMA_PLL0_REG_BIAS_QP                = 1,            //  
parameter   integer PMA_PLL0_REG_BIAS_LANE_SYNC         = 1,            //  
parameter   integer PMA_PLL0_REG_BIAS_CLKBUFS1          = 1,            //
////parameter   integer PMA_PLL0_REG_BIAS_CLKBUFS2          = 1,             //
parameter   integer PMA_PLL0_REG_TXPCLK_SEL             = 0,             //2018_7_17
parameter   integer PMA_PLL0_REG_BIAS_CLKBUFS3          = 1,             //
////parameter   integer PMA_PLL0_REG_BIAS_CLKBUFS4          = 1,             //
parameter           PMA_PLL0_REG_LANE_SYNC_EN           = "FALSE",       //FALSE,TRUE
parameter           PMA_PLL0_REG_LANE_SYNC_EN_OW        = "DISABLE",       //DISABLE,ENABLE,2018_7_17
parameter   integer PMA_PLL0_REG_BIAS_D2S               = 1,             //
parameter   integer PMA_PLL0_REG_BIAS_REFD2S_C          = 1,             //
parameter   integer PMA_PLL0_REG_BIAS_VCRST_C           = 1,             //
parameter   integer PMA_PLL0_REG_BIAS_REFBUF_C          = 1,             //
parameter   integer PMA_PLL0_REG_CLKBUFS1_C             = 1,             //
parameter   integer PMA_PLL0_REG_CLKBUFS2_C             = 6,             //
parameter   integer PMA_PLL0_REG_CLKBUFS3_C             = 6,             //
parameter   integer PMA_PLL0_REG_CLKBUFS4_C             = 1,             //
////parameter   integer PMA_PLL0_REG_D2S_C                  = 3,             //
parameter   integer PMA_PLL0_REG_PLL_REFCLK_CML_SEL     = 0,             //
parameter           PMA_PLL0_REG_REFCLK_SEL             = "FALSE",       //FALSE,TRUE 
parameter           PMA_PLL0_REG_RESCAL_R_CODE_SIGN     = "TRUE",        //FALSE,TRUE
parameter           PMA_PLL0_REG_PLL_UNLOCKED_OW        = "DISABLE",     //DISABLE,ENABLE  
parameter           PMA_PLL0_REG_PLL_UNLOCKED           = "FALSE",       //FALSE,TRUE    
parameter           PMA_PLL0_REG_PLL_LOCKDET_MODE       = "FALSE",       //FALSE,TRUE 
parameter           PMA_PLL0_REG_PLL_CLKBUF_PD_LEFT     = "ON",          //ON,OFF   ON=poweron,OFF= powerdown  
parameter           PMA_PLL0_REG_PLL_CLKBUF_PD_RIGHT    = "ON",          //ON,OFF   ON=poweron,OFF= powerdown 
////parameter   integer PMA_PLL0_REG_REFCLK_CML_SEL         = 0,             //
parameter           PMA_PLL0_REG_RESCAL_EN              = "FALSE",       //FALSE,TRUE
parameter   integer PMA_PLL0_REG_RESCAL_I_CODE_VAL      = 0,             //
////parameter           PMA_PLL0_REG_LANE_SYNC_PD_LEFT      = "ON",          //ON,OFF   ON=poweron,OFF= powerdown  
////parameter           PMA_PLL0_REG_LANE_SYNC_PD_RIGHT     = "ON",          //ON,OFF   ON=poweron,OFF= powerdown 
////parameter           PMA_PLL0_REG_TXPCLK_ON_PD_LEFT      = "ON",          //ON,OFF   ON=poweron,OFF= powerdown
////parameter           PMA_PLL0_REG_TXPCLK_ON_PD_RIGHT     = "ON",          //ON,OFF   ON=poweron,OFF= powerdown
parameter   integer PMA_PLL0_REG_RESCAL_I_CODE_OW       = 0,             //
parameter   integer PMA_PLL0_REG_RESCAL_ITER_VALID_SEL  = 0,             //
parameter   integer PMA_PLL0_REG_RESCAL_WAIT_SEL        = 0,             //
parameter   integer PMA_PLL0_REG_I_CTRL_MAX             = 45,            //
parameter   integer PMA_PLL0_REG_I_CTRL_MIN             = 19,            //
//                  
parameter           PARM_CFG_HSST_RSTN                  = "FALSE",       //FALSE,TRUE  FALSE=low, TRUE=high
parameter           PARM_PLL0_POWERUP                   = "OFF",         //ON,OFF   ON=poweron,OFF= powerdown
parameter           PARM_PLL0_RSTN                      = "FALSE",       //FALSE,TRUE  FALSE=low, TRUE=high
//pll0 end          
//pll1              
parameter           PMA_PLL1_REG_PLL_POWERDOWN_OW       = "DISABLE",     //DISABLE,ENABLE  enable REG_PLL_POWERDOWN
parameter           PMA_PLL1_REG_PLL_POWERDOWN          = "ON",         //ON,OFF   ON=poweron,OFF= powerdown
parameter           PMA_PLL1_REG_PLL_RESET_N_OW         = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_PLL1_REG_PLL_RESET_N            = "TRUE",       //FALSE,TRUE  FALSE=low, TRUE=high
parameter           PMA_PLL1_REG_PLL_READY_OW           = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_PLL1_REG_PLL_READY              = "FALSE",      //FALSE,TRUE
parameter           PMA_PLL1_REG_LANE_SYNC_OW           = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_PLL1_REG_LANE_SYNC              = "FALSE",       //FALSE,TRUE
////parameter           PMA_PLL1_REG_RESCAL_ENABLE_OW       = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_PLL1_REG_LOCKDET_REPEAT         = "DISABLE",     //DISABLE,ENABLE
////parameter           PMA_PLL1_REG_RESCAL_ENABLE          = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_PLL1_REG_RESCAL_I_CODE_PMA      = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_PLL1_REG_RESCAL_RESET_N_OW      = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_PLL1_REG_RESCAL_RESET_N         = "FALSE",       //FALSE,TRUE  FALSE=low, TRUE=high
parameter           PMA_PLL1_REG_RESCAL_DONE_OW         = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_PLL1_REG_RESCAL_DONE            = "FALSE",       //FALSE,TRUE
parameter           PMA_PLL1_REG_RESCAL_CODE_OW         = "DISABLE",     //DISABLE,ENABLE
////parameter   integer PMA_PLL1_REG_RESCAL_I_OFFSET        = 1,             // 
parameter   integer PMA_PLL1_REG_LDO_VREF_SEL           = 2,
parameter   integer PMA_PLL1_REG_BIAS_VCOREP_C          = 1,
////parameter   integer PMA_PLL1_REG_RESCAL_R_OFFSET        = 14,            // 
parameter   integer PMA_PLL1_REG_RESCAL_I_CODE          = 32,
parameter           PMA_PLL1_REG_RESCAL_ONCHIP_SMALL_OW = "DISABLE",     //DISABLE,ENABLE
parameter   integer PMA_PLL1_REG_RESCAL_ONCHIP_SMALL    = 0,            // 
////parameter   integer PMA_PLL1_REG_RESCAL_ITER            = 0,            // 
parameter           PMA_PLL1_REG_JTAG_OE                = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_PLL1_REG_JTAG_AC_MODE           = "DISABLE",     //DISABLE,ENABLE
////parameter           PMA_PLL1_REG_RESCAL_REPEAT_EN       = "DISABLE",     //DISABLE,ENABLE
////parameter   integer PMA_PLL1_REG_RESCAL_TIMEOUT         = 0,             // 
parameter   integer PMA_PLL1_REG_JTAG_VHYSTSEL          = 0,
parameter           PMA_PLL1_REG_PLL_LOCKDET_EN_OW      = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_PLL1_REG_PLL_LOCKDET_EN         = "FALSE",       //FALSE,TRUE
parameter           PMA_PLL1_REG_PLL_LOCKDET_RESET_N_OW = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_PLL1_REG_PLL_LOCKDET_RESET_N    = "FALSE",       //FALSE,TRUE  FALSE=low, TRUE=high
parameter           PMA_PLL1_REG_PLL_LOCKED_OW          = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_PLL1_REG_PLL_LOCKED             = "FALSE",       //FALSE,TRUE
parameter           PMA_PLL1_REG_PLL_LOCKED_STICKY_CLEAR= "FALSE",       //FALSE,TRUE
parameter           PMA_PLL1_REG_PLL_UNLOCKED_STICKY_CLEAR= "FALSE",       //FALSE,TRUE
parameter           PMA_PLL1_REG_NOFBCLK_STICKY_CLEAR   = "FALSE",       //FALSE,TRUE
parameter   integer PMA_PLL1_REG_PLL_LOCKDET_REFCT      = 7,             // 
parameter   integer PMA_PLL1_REG_PLL_LOCKDET_FBCT       = 7,             // 
parameter   integer PMA_PLL1_REG_PLL_LOCKDET_LOCKCT     = 4,             // 
parameter   integer PMA_PLL1_REG_PLL_LOCKDET_ITER       = 3,             // 
parameter   integer PMA_PLL1_REG_PLL_UNLOCKDET_ITER     = 2,             //
parameter           PMA_PLL1_REG_PD_VCO                 = "ON",          //ON,OFF   ON=poweron,OFF= powerdown   
parameter           PMA_PLL1_REG_FBCLK_TEST_EN          = "FALSE",       //FALSE,TRUE
parameter           PMA_PLL1_REG_REFCLK_TEST_EN         = "FALSE",       //FALSE,TRUE
parameter   integer PMA_PLL1_REG_TEST_SEL               = 0,            // 
parameter           PMA_PLL1_REG_TEST_V_EN              = "FALSE",       //FALSE,TRUE
parameter           PMA_PLL1_REG_TEST_SIG_HALF_EN       = "FALSE",       //FALSE,TRUE
parameter   integer PMA_PLL1_REG_TEST_FSM               = 0,             // 
parameter           PMA_PLL1_REG_REFCLK_OUT_PD          = "OFF",         //ON,OFF   ON=poweron,OFF= powerdown 
parameter           PMA_PLL1_REG_BGR_STARTUP_EN         = "FALSE",       //FALSE,TRUE
parameter           PMA_PLL1_REG_BGR_STARTUP            = "FALSE",       //FALSE,TRUE
parameter           PMA_PLL1_REG_PD_BGR                 = "ON",          //ON,OFF   ON=poweron,OFF= powerdown  
parameter           PMA_PLL1_REG_REFCLK_TERM_VCM_EN     = "TRUE",        //FALSE,TRUE
parameter           PMA_PLL1_REG_FBDIVA_5_EN            = "TRUE",        //FALSE,TRUE
parameter   integer PMA_PLL1_REG_FBDIVB                 = 1,             //  
parameter           PMA_PLL1_REG_RESET_N_PFDQP_OW       = "DISABLE",     //DISABLE,ENABLE
parameter           PMA_PLL1_REG_RESET_N_PFDQP          = "FALSE",       //FALSE,TRUE  FALSE=low, TRUE=high
parameter   integer PMA_PLL1_REG_QPCURRENT              = 12,            //  
parameter           PMA_PLL1_REG_VC_FORCE_EN            = "FALSE",       //FALSE,TRUE
parameter   integer PMA_PLL1_REG_VCRESET_C_RING         = 24,            //  
parameter   integer PMA_PLL1_REG_LPF_R_C                = 0,            // 
parameter   integer PMA_PLL1_REG_LPF_TR_C               = 2,            //
parameter           PMA_PLL1_REG_PD_BIAS                = "ON",          //ON,OFF   ON=poweron,OFF= powerdown  
parameter   integer PMA_PLL1_REG_ICTRL_PLL              = 1,             //  
parameter   integer PMA_PLL1_REG_BIAS_QP                = 1,             //  
parameter   integer PMA_PLL1_REG_BIAS_LANE_SYNC         = 1,             //  
parameter   integer PMA_PLL1_REG_BIAS_CLKBUFS1          = 1,             //
////parameter   integer PMA_PLL1_REG_BIAS_CLKBUFS2          = 1,             //
parameter   integer PMA_PLL1_REG_TXPCLK_SEL             = 0,             //2018_7_17
parameter   integer PMA_PLL1_REG_BIAS_CLKBUFS3          = 1,             //
////parameter   integer PMA_PLL1_REG_BIAS_CLKBUFS4          = 1,             //
parameter           PMA_PLL1_REG_LANE_SYNC_EN           = "FALSE",       //FALSE,TRUE
parameter           PMA_PLL1_REG_LANE_SYNC_EN_OW        = "DISABLE",       //DISABLE,ENABLE,2018_7_17
parameter   integer PMA_PLL1_REG_BIAS_D2S               = 1,             //
parameter   integer PMA_PLL1_REG_BIAS_REFD2S_C          = 1,             //
parameter   integer PMA_PLL1_REG_BIAS_VCRST_C           = 1,             //
parameter   integer PMA_PLL1_REG_BIAS_REFBUF_C          = 1,             //
parameter   integer PMA_PLL1_REG_CLKBUFS1_C             = 1,             //
parameter   integer PMA_PLL1_REG_CLKBUFS2_C             = 6,             //
parameter   integer PMA_PLL1_REG_CLKBUFS3_C             = 6,             //
parameter   integer PMA_PLL1_REG_CLKBUFS4_C             = 1,             //
////parameter   integer PMA_PLL1_REG_D2S_C                  = 3,             //
parameter   integer PMA_PLL1_REG_PLL_REFCLK_CML_SEL     = 0,             //
parameter           PMA_PLL1_REG_REFCLK_SEL             = "FALSE",       //FALSE,TRUE 
parameter           PMA_PLL1_REG_RESCAL_R_CODE_SIGN     = "TRUE",        //FALSE,TRUE
parameter           PMA_PLL1_REG_PLL_UNLOCKED_OW        = "DISABLE",     //DISABLE,ENABLE  
parameter           PMA_PLL1_REG_PLL_UNLOCKED           = "FALSE",      //FALSE,TRUE    
parameter           PMA_PLL1_REG_PLL_LOCKDET_MODE       = "FALSE",      //FALSE,TRUE 
parameter           PMA_PLL1_REG_PLL_CLKBUF_PD_LEFT     = "ON",          //ON,OFF   ON=poweron,OFF= powerdown  
parameter           PMA_PLL1_REG_PLL_CLKBUF_PD_RIGHT    = "ON",          //ON,OFF   ON=poweron,OFF= powerdown 
////parameter   integer PMA_PLL1_REG_REFCLK_CML_SEL         = 0,             //
parameter           PMA_PLL1_REG_RESCAL_EN              = "FALSE",       //FALSE,TRUE
parameter   integer PMA_PLL1_REG_RESCAL_I_CODE_VAL      = 0,             //
////parameter           PMA_PLL1_REG_LANE_SYNC_PD_LEFT      = "ON",          //ON,OFF   ON=poweron,OFF= powerdown  
////parameter           PMA_PLL1_REG_LANE_SYNC_PD_RIGHT     = "ON",          //ON,OFF   ON=poweron,OFF= powerdown 
////parameter           PMA_PLL1_REG_TXPCLK_ON_PD_LEFT      = "ON",          //ON,OFF   ON=poweron,OFF= powerdown
////parameter           PMA_PLL1_REG_TXPCLK_ON_PD_RIGHT     = "ON",          //ON,OFF   ON=poweron,OFF= powerdown
parameter   integer PMA_PLL1_REG_RESCAL_I_CODE_OW       = 0,             //
parameter   integer PMA_PLL1_REG_RESCAL_ITER_VALID_SEL  = 0,             //
parameter   integer PMA_PLL1_REG_RESCAL_WAIT_SEL        = 0,             //
parameter   integer PMA_PLL1_REG_I_CTRL_MAX             = 45,            //
parameter   integer PMA_PLL1_REG_I_CTRL_MIN             = 19,            //
//                  
parameter           PARM_PLL1_POWERUP                   = "OFF",          //ON,OFF   ON=poweron,OFF= powerdown
parameter           PARM_PLL1_RSTN                      = "FALSE",       //FALSE,TRUE  FALSE=low, TRUE=high
//PMA PLL end       
parameter           PARM_GRSN_DIS                       = "FALSE",       //FALSE,TRUE  FALSE=low, TRUE=high
parameter           PARM_CFG_RSTN                       = "FALSE"       //FALSE,TRUE  FALSE=low, TRUE=high

)
(
///////////////////////////
/////PORT DECLARATIONS/////
///////////////////////////
        //if with port
input                P_REFCLKP_0,
input                P_REFCLKN_0,
output               P_PLL_TEST_0,
input                P_REFCLKP_1,       
input                P_REFCLKN_1,            
output               P_PLL_TEST_1,
input                P_RX_SDP0,     
input                P_RX_SDN0,        
output               P_TX_SDP0,
output               P_TX_SDN0,
input                P_RX_SDP1,                                
input                P_RX_SDN1,        
output               P_TX_SDP1,
output               P_TX_SDN1,        
input                P_RX_SDP2,                                
input                P_RX_SDN2,        
output               P_TX_SDP2,
output               P_TX_SDN2,  
input                P_RX_SDP3,                                
input                P_RX_SDN3,        
output               P_TX_SDP3,
output               P_TX_SDN3,  
        //if with user logic
input                P_RX0_CLK_FR_CORE,       
input                P_RX1_CLK_FR_CORE,         
input                P_RX2_CLK_FR_CORE,         
input                P_RX3_CLK_FR_CORE,         
input                P_TX0_CLK_FR_CORE,       
input                P_TX1_CLK_FR_CORE,         
input                P_TX2_CLK_FR_CORE,         
input                P_TX3_CLK_FR_CORE, 
input                P_HSST_RST,
input                P_PCS_RX_RST_0,
input                P_PCS_RX_RST_1,        
input                P_PCS_RX_RST_2,
input                P_PCS_RX_RST_3,        
input                P_PCS_TX_RST_0,
input                P_PCS_TX_RST_1,        
input                P_PCS_TX_RST_2,        
input                P_PCS_TX_RST_3,
input                P_CFG_CLK,
input                P_CFG_RST,
input                P_CFG_ENABLE,
input                P_CFG_WRITE,
input    [15:0]      P_CFG_ADDR,
input    [7:0]       P_CFG_WDATA,
input    [44:0]      P_TDATA_0,
input    [44:0]      P_TDATA_1,
input    [44:0]      P_TDATA_2,
input    [44:0]      P_TDATA_3,
input    [3:0]       P_PCS_WORD_ALIGN_EN,
input    [3:0]       P_RX_POLARITY_INVERT,
input    [3:0]       P_CEB_ADETECT_EN,
input    [3:0]       P_PCS_MCB_EXT_EN,
input    [3:0]       P_PCS_NEAREND_LOOP,
input    [3:0]       P_PCS_FAREND_LOOP,
output               P_CFG_READY,
output   [7:0]       P_CFG_RDATA,
output               P_CFG_INT,
output   [3:0]       P_PCS_RX_MCB_STATUS,
output   [3:0]       P_PCS_LSM_SYNCED,
output   [46:0]      P_RDATA_0,
output   [46:0]      P_RDATA_1,
output   [46:0]      P_RDATA_2,
output   [46:0]      P_RDATA_3,
output   [3:0]       P_RCLK2FABRIC,
output   [3:0]       P_TCLK2FABRIC,
input                P_RESCAL_RST_I,       
input    [5:0]       P_RESCAL_I_CODE_I,   
output   [5:0]       P_RESCAL_I_CODE_O,
output               P_REFCK2CORE_0,
input                P_PLL_REF_CLK_0,
input                P_PLL_RST_0,
input                P_PLLPOWERDOWN_0,
output               P_PLL_READY_0,
input                P_LANE_SYNC_0,
input                P_LANE_SYNC_EN_0,
input                P_RATE_CHANGE_TCLK_ON_0,
output               P_REFCK2CORE_1,
input                P_PLL_REF_CLK_1,
input                P_PLL_RST_1,
input                P_PLLPOWERDOWN_1,
output               P_PLL_READY_1,
input                P_LANE_SYNC_1,
input                P_LANE_SYNC_EN_1,
input                P_RATE_CHANGE_TCLK_ON_1,
//Lanes
input                P_LANE_PD_0,
input                P_LANE_RST_0,
input                P_RX_LANE_PD_0,
input                P_RX_PMA_RST_0,
output               P_RX_SIGDET_STATUS_0,
output               P_RX_SATA_COMINIT_0,
output               P_RX_SATA_COMWAKE_0,
output               P_RX_LS_DATA_0,
output               P_RX_READY_0,
output   [19:0]      P_TEST_STATUS_0,
input    [1:0]       P_TX_DEEMP_0,
input                P_TX_LS_DATA_0,
input                P_TX_BEACON_EN_0,
input                P_TX_SWING_0,
input                P_TX_RXDET_REQ_0,
input    [2:0]       P_TX_RATE_0,
input    [2:0]       P_TX_BUSWIDTH_0,
input    [2:0]       P_TX_MARGIN_0,
output               P_TX_RXDET_STATUS_0,
input                P_TX_PMA_RST_0,
input                P_TX_LANE_PD_0,
input    [2:0]       P_RX_RATE_0,
input    [2:0]       P_RX_BUSWIDTH_0,
input                P_RX_HIGHZ_0,
output   [3:0]       P_CA_ALIGN_RX,
output   [3:0]       P_CA_ALIGN_TX,
input    [7:0]       P_CIM_CLK_ALIGNER_RX0,
input    [7:0]       P_CIM_CLK_ALIGNER_TX0,
input                P_CIM_DYN_DLY_SEL_RX0,
input                P_CIM_DYN_DLY_SEL_TX0,
input                P_CIM_START_ALIGN_RX0,
input                P_CIM_START_ALIGN_TX0,
input                P_LANE_PD_1,
input                P_LANE_RST_1,
input                P_RX_LANE_PD_1,
input                P_RX_PMA_RST_1,
output               P_RX_SIGDET_STATUS_1,
output               P_RX_SATA_COMINIT_1,
output               P_RX_SATA_COMWAKE_1,
output               P_RX_LS_DATA_1,
output               P_RX_READY_1,
output   [19:0]      P_TEST_STATUS_1,
input    [1:0]       P_TX_DEEMP_1,
input                P_TX_LS_DATA_1,
input                P_TX_BEACON_EN_1,
input                P_TX_SWING_1,
input                P_TX_RXDET_REQ_1,
input    [2:0]       P_TX_RATE_1,
input    [2:0]       P_TX_BUSWIDTH_1,
input    [2:0]       P_TX_MARGIN_1,
output               P_TX_RXDET_STATUS_1,
input                P_TX_PMA_RST_1,
input                P_TX_LANE_PD_1,
input    [2:0]       P_RX_RATE_1,
input    [2:0]       P_RX_BUSWIDTH_1,
input                P_RX_HIGHZ_1,
input    [7:0]       P_CIM_CLK_ALIGNER_RX1,
input    [7:0]       P_CIM_CLK_ALIGNER_TX1,
input                P_CIM_DYN_DLY_SEL_RX1,
input                P_CIM_DYN_DLY_SEL_TX1,
input                P_CIM_START_ALIGN_RX1,
input                P_CIM_START_ALIGN_TX1,
input                P_LANE_PD_2,
input                P_LANE_RST_2,
input                P_RX_LANE_PD_2,
input                P_RX_PMA_RST_2,
output               P_RX_SIGDET_STATUS_2,
output               P_RX_SATA_COMINIT_2,
output               P_RX_SATA_COMWAKE_2,
output               P_RX_LS_DATA_2,
output               P_RX_READY_2,
output   [19:0]      P_TEST_STATUS_2,
input    [1:0]       P_TX_DEEMP_2,
input                P_TX_LS_DATA_2,
input                P_TX_BEACON_EN_2,
input                P_TX_SWING_2,
input                P_TX_RXDET_REQ_2,
input    [2:0]       P_TX_RATE_2,
input    [2:0]       P_TX_BUSWIDTH_2,
input    [2:0]       P_TX_MARGIN_2,
output               P_TX_RXDET_STATUS_2,
input                P_TX_PMA_RST_2,
input                P_TX_LANE_PD_2,
input    [2:0]       P_RX_RATE_2,
input    [2:0]       P_RX_BUSWIDTH_2,
input                P_RX_HIGHZ_2,
input    [7:0]       P_CIM_CLK_ALIGNER_RX2,
input    [7:0]       P_CIM_CLK_ALIGNER_TX2,
input                P_CIM_DYN_DLY_SEL_RX2,
input                P_CIM_DYN_DLY_SEL_TX2,
input                P_CIM_START_ALIGN_RX2,
input                P_CIM_START_ALIGN_TX2,
input                P_LANE_PD_3,
input                P_LANE_RST_3,
input                P_RX_LANE_PD_3,
input                P_RX_PMA_RST_3,
output               P_RX_SIGDET_STATUS_3,
output               P_RX_SATA_COMINIT_3,
output               P_RX_SATA_COMWAKE_3,
output               P_RX_LS_DATA_3,
output               P_RX_READY_3,
output   [19:0]      P_TEST_STATUS_3,
input    [1:0]       P_TX_DEEMP_3,
input                P_TX_LS_DATA_3,
input                P_TX_BEACON_EN_3,
input                P_TX_SWING_3,
input                P_TX_RXDET_REQ_3,
input    [2:0]       P_TX_RATE_3,
input    [2:0]       P_TX_BUSWIDTH_3,
input    [2:0]       P_TX_MARGIN_3,
output               P_TX_RXDET_STATUS_3,
input                P_TX_PMA_RST_3,
input                P_TX_LANE_PD_3,
input    [2:0]       P_RX_RATE_3,
input    [2:0]       P_RX_BUSWIDTH_3,
input                P_RX_HIGHZ_3,
input    [7:0]       P_CIM_CLK_ALIGNER_RX3,
input    [7:0]       P_CIM_CLK_ALIGNER_TX3,
input                P_CIM_DYN_DLY_SEL_RX3,
input                P_CIM_DYN_DLY_SEL_TX3,
input                P_CIM_START_ALIGN_RX3,
input                P_CIM_START_ALIGN_TX3

);


HSST 
#(
    .CP_PCS_CH0_BYPASS_WORD_ALIGN                (PCS_CH0_BYPASS_WORD_ALIGN),    
    .CP_PCS_CH0_BYPASS_DENC                      (PCS_CH0_BYPASS_DENC),         
    .CP_PCS_CH0_BYPASS_BONDING                   (PCS_CH0_BYPASS_BONDING),      
    .CP_PCS_CH0_BYPASS_CTC                       (PCS_CH0_BYPASS_CTC),          
    .CP_PCS_CH0_BYPASS_GEAR                      (PCS_CH0_BYPASS_GEAR),         
    .CP_PCS_CH0_BYPASS_BRIDGE                    (PCS_CH0_BYPASS_BRIDGE),       
    .CP_PCS_CH0_DATA_MODE                        (PCS_CH0_DATA_MODE),           
    .CP_PCS_CH0_RX_POLARITY_INV                  (PCS_CH0_RX_POLARITY_INV),     
    .CP_PCS_CH0_ALIGN_MODE                       (PCS_CH0_ALIGN_MODE),          
    .CP_PCS_CH0_SAMP_16B                         (PCS_CH0_SAMP_16B),            
    .CP_PCS_CH0_COMMA_REG0                       (PCS_CH0_COMMA_REG0),          
    .CP_PCS_CH0_COMMA_MASK                       (PCS_CH0_COMMA_MASK),          
    .CP_PCS_CH0_CEB_MODE                         (PCS_CH0_CEB_MODE),            
    .CP_PCS_CH0_CTC_MODE                         (PCS_CH0_CTC_MODE),            
    .CP_PCS_CH0_A_REG                            (PCS_CH0_A_REG),               
    .CP_PCS_CH0_GE_AUTO_EN                       (PCS_CH0_GE_AUTO_EN),          
    .CP_PCS_CH0_SKIP_REG0                        (PCS_CH0_SKIP_REG0),           
    .CP_PCS_CH0_SKIP_REG1                        (PCS_CH0_SKIP_REG1),           
    .CP_PCS_CH0_SKIP_REG2                        (PCS_CH0_SKIP_REG2),           
    .CP_PCS_CH0_SKIP_REG3                        (PCS_CH0_SKIP_REG3),           
    .CP_PCS_CH0_DEC_DUAL                         (PCS_CH0_DEC_DUAL),             
    .CP_PCS_CH0_SPLIT                            (PCS_CH0_SPLIT),                
    .CP_PCS_CH0_FIFOFLAG_CTC                     (PCS_CH0_FIFOFLAG_CTC),         
    .CP_PCS_CH0_COMMA_DET_MODE                   (PCS_CH0_COMMA_DET_MODE),       
    .CP_PCS_CH0_ERRDETECT_SILENCE                (PCS_CH0_ERRDETECT_SILENCE),    
    .CP_PCS_CH0_PMA_RCLK_POLINV                  (PCS_CH0_PMA_RCLK_POLINV),      
    .CP_PCS_CH0_PCS_RCLK_SEL                     (PCS_CH0_PCS_RCLK_SEL),         
    .CP_PCS_CH0_MCB_RCLK_POLINV                  (PCS_CH0_MCB_RCLK_POLINV),      
    .CP_PCS_CH0_CB_RCLK_SEL                      (PCS_CH0_CB_RCLK_SEL),           
    .CP_PCS_CH0_AFTER_CTC_RCLK_SEL               (PCS_CH0_AFTER_CTC_RCLK_SEL),    
    .CP_PCS_CH0_RCLK_POLINV                      (PCS_CH0_RCLK_POLINV),              
    .CP_PCS_CH0_BRIDGE_RCLK_SEL                  (PCS_CH0_BRIDGE_RCLK_SEL),          
    .CP_PCS_CH0_PCS_RCLK_EN                      (PCS_CH0_PCS_RCLK_EN),              
    .CP_PCS_CH0_CB_RCLK_EN                       (PCS_CH0_CB_RCLK_EN),               
    .CP_PCS_CH0_AFTER_CTC_RCLK_EN                (PCS_CH0_AFTER_CTC_RCLK_EN),        
    .CP_PCS_CH0_AFTER_CTC_RCLK_EN_GB             (PCS_CH0_AFTER_CTC_RCLK_EN_GB),     
    .CP_PCS_CH0_BRIDGE_RCLK_EN                   (PCS_CH0_BRIDGE_RCLK_EN),           
    .CP_PCS_CH0_PCS_RX_RSTN                      (PCS_CH0_PCS_RX_RSTN),              
    .CP_PCS_CH0_SLAVE                            (PCS_CH0_SLAVE),                    
    .CP_PCS_CH0_PCIE_SLAVE                       (PCS_CH0_PCIE_SLAVE),                
    .CP_PCS_CH0_PCS_CB_RSTN                      (PCS_CH0_PCS_CB_RSTN),               
    .CP_PCS_CH0_TX_BYPASS_BRIDGE_UINT            (PCS_CH0_TX_BYPASS_BRIDGE_UINT),     
    .CP_PCS_CH0_TX_BYPASS_GEAR                   (PCS_CH0_TX_BYPASS_GEAR),            
    .CP_PCS_CH0_TX_BYPASS_ENC                    (PCS_CH0_TX_BYPASS_ENC),             
    .CP_PCS_CH0_TX_BYPASS_BIT_SLIP               (PCS_CH0_TX_BYPASS_BIT_SLIP),        
    .CP_PCS_CH0_TX_GEAR_SPLIT                    (PCS_CH0_TX_GEAR_SPLIT),             
    .CP_PCS_CH0_TX_DRIVE_REG_MODE                (PCS_CH0_TX_DRIVE_REG_MODE),          
    .CP_PCS_CH0_TX_BIT_SLIP_CYCLES               (PCS_CH0_TX_BIT_SLIP_CYCLES),         
    .CP_PCS_CH0_INT_TX_MASK_0                    (PCS_CH0_INT_TX_MASK_0),              
    .CP_PCS_CH0_INT_TX_MASK_1                    (PCS_CH0_INT_TX_MASK_1),              
    .CP_PCS_CH0_INT_TX_MASK_2                    (PCS_CH0_INT_TX_MASK_2),              
    .CP_PCS_CH0_INT_TX_CLR_0                     (PCS_CH0_INT_TX_CLR_0),               
    .CP_PCS_CH0_INT_TX_CLR_1                     (PCS_CH0_INT_TX_CLR_1),               
    .CP_PCS_CH0_INT_TX_CLR_2                     (PCS_CH0_INT_TX_CLR_2),               
    .CP_PCS_CH0_TX_PMA_TCLK_POLINV               (PCS_CH0_TX_PMA_TCLK_POLINV),           
    .CP_PCS_CH0_TX_PCS_CLK_EN_SEL                (PCS_CH0_TX_PCS_CLK_EN_SEL),            
    .CP_PCS_CH0_TX_BRIDGE_TCLK_SEL               (PCS_CH0_TX_BRIDGE_TCLK_SEL),           
    .CP_PCS_CH0_TX_TCLK_POLINV                   (PCS_CH0_TX_TCLK_POLINV),               
    .CP_PCS_CH0_TX_PCS_TX_RSTN                   (PCS_CH0_TX_PCS_TX_RSTN),               
    .CP_PCS_CH0_TX_SLAVE                         (PCS_CH0_TX_SLAVE),                     
    .CP_PCS_CH0_TX_BRIDGE_CLK_EN_SEL             (PCS_CH0_TX_BRIDGE_CLK_EN_SEL),         
    .CP_PCS_CH0_DATA_WIDTH_MODE                  (PCS_CH0_DATA_WIDTH_MODE),              
    .CP_PCS_CH0_TX_TCLK2FABRIC_SEL               (PCS_CH0_TX_TCLK2FABRIC_SEL),           
    .CP_PCS_CH0_TX_OUTZZ                         (PCS_CH0_TX_OUTZZ),                     
    .CP_PCS_CH0_ENC_DUAL                         (PCS_CH0_ENC_DUAL),             
    .CP_PCS_CH0_TX_BITSLIP_DATA_MODE             (PCS_CH0_TX_BITSLIP_DATA_MODE), 
    .CP_PCS_CH0_COMMA_REG1                       (PCS_CH0_COMMA_REG1),           
    .CP_PCS_CH0_RAPID_IMAX                       (PCS_CH0_RAPID_IMAX),           
    .CP_PCS_CH0_RAPID_VMIN_1                     (PCS_CH0_RAPID_VMIN_1),         
    .CP_PCS_CH0_RAPID_VMIN_2                     (PCS_CH0_RAPID_VMIN_2),            
    .CP_PCS_CH0_RX_PRBS_MODE                     (PCS_CH0_RX_PRBS_MODE),            
    .CP_PCS_CH0_RX_ERRCNT_CLR                    (PCS_CH0_RX_ERRCNT_CLR),           
    .CP_PCS_CH0_TX_PRBS_MODE                     (PCS_CH0_TX_PRBS_MODE),            
    .CP_PCS_CH0_TX_INSERT_ER                     (PCS_CH0_TX_INSERT_ER),            
    .CP_PCS_CH0_ENABLE_PRBS_GEN                  (PCS_CH0_ENABLE_PRBS_GEN),      
    .CP_PCS_CH0_ERR_CNT                          (PCS_CH0_ERR_CNT),              
    .CP_PCS_CH0_DEFAULT_RADDR                    (PCS_CH0_DEFAULT_RADDR),        
    .CP_PCS_CH0_MASTER_CHECK_OFFSET              (PCS_CH0_MASTER_CHECK_OFFSET),  
    .CP_PCS_CH0_DELAY_SET                        (PCS_CH0_DELAY_SET),            
    .CP_PCS_CH0_SEACH_OFFSET                     (PCS_CH0_SEACH_OFFSET),         
    .CP_PCS_CH0_CEB_RAPIDLS_MMAX                 (PCS_CH0_CEB_RAPIDLS_MMAX),     
    .CP_PCS_CH0_CTC_AFULL                        (PCS_CH0_CTC_AFULL),            
    .CP_PCS_CH0_CTC_AEMPTY                       (PCS_CH0_CTC_AEMPTY),           
    .CP_PCS_CH0_CTC_CONTI_SKP_SET                (PCS_CH0_CTC_CONTI_SKP_SET),      
    .CP_PCS_CH0_FAR_LOOP                         (PCS_CH0_FAR_LOOP),               
    .CP_PCS_CH0_NEAR_LOOP                        (PCS_CH0_NEAR_LOOP),              
    .CP_PCS_CH0_INT_RX_MASK_0                    (PCS_CH0_INT_RX_MASK_0),          
    .CP_PCS_CH0_INT_RX_MASK_1                    (PCS_CH0_INT_RX_MASK_1),          
    .CP_PCS_CH0_INT_RX_MASK_2                    (PCS_CH0_INT_RX_MASK_2),          
    .CP_PCS_CH0_INT_RX_MASK_3                    (PCS_CH0_INT_RX_MASK_3),          
    .CP_PCS_CH0_INT_RX_MASK_4                    (PCS_CH0_INT_RX_MASK_4),          
    .CP_PCS_CH0_INT_RX_MASK_5                    (PCS_CH0_INT_RX_MASK_5),          
    .CP_PCS_CH0_INT_RX_MASK_6                    (PCS_CH0_INT_RX_MASK_6),          
    .CP_PCS_CH0_INT_RX_MASK_7                    (PCS_CH0_INT_RX_MASK_7),          
    .CP_PCS_CH0_INT_RX_CLR_0                     (PCS_CH0_INT_RX_CLR_0),             
    .CP_PCS_CH0_INT_RX_CLR_1                     (PCS_CH0_INT_RX_CLR_1),             
    .CP_PCS_CH0_INT_RX_CLR_2                     (PCS_CH0_INT_RX_CLR_2),             
    .CP_PCS_CH0_INT_RX_CLR_3                     (PCS_CH0_INT_RX_CLR_3),             
    .CP_PCS_CH0_INT_RX_CLR_4                     (PCS_CH0_INT_RX_CLR_4),           
    .CP_PCS_CH0_INT_RX_CLR_5                     (PCS_CH0_INT_RX_CLR_5),           
    .CP_PCS_CH0_INT_RX_CLR_6                     (PCS_CH0_INT_RX_CLR_6),           
    .CP_PCS_CH0_INT_RX_CLR_7                     (PCS_CH0_INT_RX_CLR_7),            
    .CP_PCS_CH0_CA_RX                            (PCS_CH0_CA_RX),                  
    .CP_PCS_CH1_CA_RX                            (PCS_CH1_CA_RX),                  
    .CP_PCS_CH2_CA_RX                            (PCS_CH2_CA_RX),                  
    .CP_PCS_CH3_CA_RX                            (PCS_CH3_CA_RX),                  
    .CP_PCS_CH0_CA_TX                            (PCS_CH0_CA_TX),                    
    .CP_PCS_CH1_CA_TX                            (PCS_CH1_CA_TX),                    
    .CP_PCS_CH2_CA_TX                            (PCS_CH2_CA_TX),                    
    .CP_PCS_CH3_CA_TX                            (PCS_CH3_CA_TX),                    
    .CP_PCS_CH0_CA_DYN_DLY_EN_RX                 (PCS_CH0_CA_DYN_DLY_EN_RX),         
    .CP_PCS_CH1_CA_DYN_DLY_EN_RX                 (PCS_CH1_CA_DYN_DLY_EN_RX),         
    .CP_PCS_CH2_CA_DYN_DLY_EN_RX                 (PCS_CH2_CA_DYN_DLY_EN_RX),         
    .CP_PCS_CH3_CA_DYN_DLY_EN_RX                 (PCS_CH3_CA_DYN_DLY_EN_RX),         
    .CP_PCS_CH0_CA_DYN_DLY_EN_TX                 (PCS_CH0_CA_DYN_DLY_EN_TX),         
    .CP_PCS_CH1_CA_DYN_DLY_EN_TX                 (PCS_CH1_CA_DYN_DLY_EN_TX),         
    .CP_PCS_CH2_CA_DYN_DLY_EN_TX                 (PCS_CH2_CA_DYN_DLY_EN_TX),         
    .CP_PCS_CH3_CA_DYN_DLY_EN_TX                 (PCS_CH3_CA_DYN_DLY_EN_TX),         
    .CP_PCS_CH0_CA_DYN_DLY_SEL_RX                (PCS_CH0_CA_DYN_DLY_SEL_RX),        
    .CP_PCS_CH1_CA_DYN_DLY_SEL_RX                (PCS_CH1_CA_DYN_DLY_SEL_RX),        
    .CP_PCS_CH2_CA_DYN_DLY_SEL_RX                (PCS_CH2_CA_DYN_DLY_SEL_RX),        
    .CP_PCS_CH3_CA_DYN_DLY_SEL_RX                (PCS_CH3_CA_DYN_DLY_SEL_RX),           
    .CP_PCS_CH0_CA_DYN_DLY_SEL_TX                (PCS_CH0_CA_DYN_DLY_SEL_TX),           
    .CP_PCS_CH1_CA_DYN_DLY_SEL_TX                (PCS_CH1_CA_DYN_DLY_SEL_TX),           
    .CP_PCS_CH2_CA_DYN_DLY_SEL_TX                (PCS_CH2_CA_DYN_DLY_SEL_TX),           
    .CP_PCS_CH3_CA_DYN_DLY_SEL_TX                (PCS_CH3_CA_DYN_DLY_SEL_TX),           
    .CP_PCS_CH0_CA_RSTN_RX                       (PCS_CH0_CA_RSTN_RX),                  
    .CP_PCS_CH1_CA_RSTN_RX                       (PCS_CH1_CA_RSTN_RX),                  
    .CP_PCS_CH2_CA_RSTN_RX                       (PCS_CH2_CA_RSTN_RX),                  
    .CP_PCS_CH3_CA_RSTN_RX                       (PCS_CH3_CA_RSTN_RX),                  
    .CP_PCS_CH0_CA_RSTN_TX                       (PCS_CH0_CA_RSTN_TX),                  
    .CP_PCS_CH1_CA_RSTN_TX                       (PCS_CH1_CA_RSTN_TX),                  
    .CP_PCS_CH2_CA_RSTN_TX                       (PCS_CH2_CA_RSTN_TX),                  
    .CP_PCS_CH3_CA_RSTN_TX                       (PCS_CH3_CA_RSTN_TX),                  
    .CP_PCS_CH1_BYPASS_WORD_ALIGN                (PCS_CH1_BYPASS_WORD_ALIGN),           
    .CP_PCS_CH1_BYPASS_DENC                      (PCS_CH1_BYPASS_DENC),                
    .CP_PCS_CH1_BYPASS_BONDING                   (PCS_CH1_BYPASS_BONDING),           
    .CP_PCS_CH1_BYPASS_CTC                       (PCS_CH1_BYPASS_CTC),               
    .CP_PCS_CH1_BYPASS_GEAR                      (PCS_CH1_BYPASS_GEAR),              
    .CP_PCS_CH1_BYPASS_BRIDGE                    (PCS_CH1_BYPASS_BRIDGE),            
    .CP_PCS_CH1_DATA_MODE                        (PCS_CH1_DATA_MODE),                
    .CP_PCS_CH1_RX_POLARITY_INV                  (PCS_CH1_RX_POLARITY_INV),          
    .CP_PCS_CH1_ALIGN_MODE                       (PCS_CH1_ALIGN_MODE),               
    .CP_PCS_CH1_SAMP_16B                         (PCS_CH1_SAMP_16B),                 
    .CP_PCS_CH1_COMMA_REG0                       (PCS_CH1_COMMA_REG0),               
    .CP_PCS_CH1_COMMA_MASK                       (PCS_CH1_COMMA_MASK),               
    .CP_PCS_CH1_CEB_MODE                         (PCS_CH1_CEB_MODE),                 
    .CP_PCS_CH1_CTC_MODE                         (PCS_CH1_CTC_MODE),                 
    .CP_PCS_CH1_A_REG                            (PCS_CH1_A_REG),                  
    .CP_PCS_CH1_GE_AUTO_EN                       (PCS_CH1_GE_AUTO_EN),             
    .CP_PCS_CH1_SKIP_REG0                        (PCS_CH1_SKIP_REG0),              
    .CP_PCS_CH1_SKIP_REG1                        (PCS_CH1_SKIP_REG1),              
    .CP_PCS_CH1_SKIP_REG2                        (PCS_CH1_SKIP_REG2),              
    .CP_PCS_CH1_SKIP_REG3                        (PCS_CH1_SKIP_REG3),              
    .CP_PCS_CH1_DEC_DUAL                         (PCS_CH1_DEC_DUAL),               
    .CP_PCS_CH1_SPLIT                            (PCS_CH1_SPLIT),                  
    .CP_PCS_CH1_FIFOFLAG_CTC                     (PCS_CH1_FIFOFLAG_CTC),           
    .CP_PCS_CH1_COMMA_DET_MODE                   (PCS_CH1_COMMA_DET_MODE),         
    .CP_PCS_CH1_ERRDETECT_SILENCE                (PCS_CH1_ERRDETECT_SILENCE),      
    .CP_PCS_CH1_PMA_RCLK_POLINV                  (PCS_CH1_PMA_RCLK_POLINV),        
    .CP_PCS_CH1_PCS_RCLK_SEL                     (PCS_CH1_PCS_RCLK_SEL),           
    .CP_PCS_CH1_MCB_RCLK_POLINV                  (PCS_CH1_MCB_RCLK_POLINV),        
    .CP_PCS_CH1_CB_RCLK_SEL                      (PCS_CH1_CB_RCLK_SEL),            
    .CP_PCS_CH1_AFTER_CTC_RCLK_SEL               (PCS_CH1_AFTER_CTC_RCLK_SEL),     
    .CP_PCS_CH1_RCLK_POLINV                      (PCS_CH1_RCLK_POLINV),            
    .CP_PCS_CH1_BRIDGE_RCLK_SEL                  (PCS_CH1_BRIDGE_RCLK_SEL),        
    .CP_PCS_CH1_PCS_RCLK_EN                      (PCS_CH1_PCS_RCLK_EN),            
    .CP_PCS_CH1_CB_RCLK_EN                       (PCS_CH1_CB_RCLK_EN),             
    .CP_PCS_CH1_AFTER_CTC_RCLK_EN                (PCS_CH1_AFTER_CTC_RCLK_EN),      
    .CP_PCS_CH1_AFTER_CTC_RCLK_EN_GB             (PCS_CH1_AFTER_CTC_RCLK_EN_GB),   
    .CP_PCS_CH1_BRIDGE_RCLK_EN                   (PCS_CH1_BRIDGE_RCLK_EN),          
    .CP_PCS_CH1_PCS_RX_RSTN                      (PCS_CH1_PCS_RX_RSTN),             
    .CP_PCS_CH1_SLAVE                            (PCS_CH1_SLAVE),                   
    .CP_PCS_CH1_PCIE_SLAVE                       (PCS_CH1_PCIE_SLAVE),              
    .CP_PCS_CH1_PCS_CB_RSTN                      (PCS_CH1_PCS_CB_RSTN),             
    .CP_PCS_CH1_TX_BYPASS_BRIDGE_UINT            (PCS_CH1_TX_BYPASS_BRIDGE_UINT),   
    .CP_PCS_CH1_TX_BYPASS_GEAR                   (PCS_CH1_TX_BYPASS_GEAR),          
    .CP_PCS_CH1_TX_BYPASS_ENC                    (PCS_CH1_TX_BYPASS_ENC),           
    .CP_PCS_CH1_TX_BYPASS_BIT_SLIP               (PCS_CH1_TX_BYPASS_BIT_SLIP),      
    .CP_PCS_CH1_TX_GEAR_SPLIT                    (PCS_CH1_TX_GEAR_SPLIT),           
    .CP_PCS_CH1_TX_DRIVE_REG_MODE                (PCS_CH1_TX_DRIVE_REG_MODE),       
    .CP_PCS_CH1_TX_BIT_SLIP_CYCLES               (PCS_CH1_TX_BIT_SLIP_CYCLES),      
    .CP_PCS_CH1_INT_TX_MASK_0                    (PCS_CH1_INT_TX_MASK_0),           
    .CP_PCS_CH1_INT_TX_MASK_1                    (PCS_CH1_INT_TX_MASK_1),           
    .CP_PCS_CH1_INT_TX_MASK_2                    (PCS_CH1_INT_TX_MASK_2),           
    .CP_PCS_CH1_INT_TX_CLR_0                     (PCS_CH1_INT_TX_CLR_0),            
    .CP_PCS_CH1_INT_TX_CLR_1                     (PCS_CH1_INT_TX_CLR_1),            
    .CP_PCS_CH1_INT_TX_CLR_2                     (PCS_CH1_INT_TX_CLR_2),            
    .CP_PCS_CH1_TX_PMA_TCLK_POLINV               (PCS_CH1_TX_PMA_TCLK_POLINV),      
    .CP_PCS_CH1_TX_PCS_CLK_EN_SEL                (PCS_CH1_TX_PCS_CLK_EN_SEL),        
    .CP_PCS_CH1_TX_BRIDGE_TCLK_SEL               (PCS_CH1_TX_BRIDGE_TCLK_SEL),       
    .CP_PCS_CH1_TX_TCLK_POLINV                   (PCS_CH1_TX_TCLK_POLINV),           
    .CP_PCS_CH1_TX_PCS_TX_RSTN                   (PCS_CH1_TX_PCS_TX_RSTN),           
    .CP_PCS_CH1_TX_SLAVE                         (PCS_CH1_TX_SLAVE),                 
    .CP_PCS_CH1_TX_BRIDGE_CLK_EN_SEL             (PCS_CH1_TX_BRIDGE_CLK_EN_SEL),     
    .CP_PCS_CH1_DATA_WIDTH_MODE                  (PCS_CH1_DATA_WIDTH_MODE),          
    .CP_PCS_CH1_TX_TCLK2FABRIC_SEL               (PCS_CH1_TX_TCLK2FABRIC_SEL),       
    .CP_PCS_CH1_TX_OUTZZ                         (PCS_CH1_TX_OUTZZ),                 
    .CP_PCS_CH1_ENC_DUAL                         (PCS_CH1_ENC_DUAL),                 
    .CP_PCS_CH1_TX_BITSLIP_DATA_MODE             (PCS_CH1_TX_BITSLIP_DATA_MODE),     
    .CP_PCS_CH1_COMMA_REG1                       (PCS_CH1_COMMA_REG1),               
    .CP_PCS_CH1_RAPID_IMAX                       (PCS_CH1_RAPID_IMAX),               
    .CP_PCS_CH1_RAPID_VMIN_1                     (PCS_CH1_RAPID_VMIN_1),             
    .CP_PCS_CH1_RAPID_VMIN_2                     (PCS_CH1_RAPID_VMIN_2),             
    .CP_PCS_CH1_RX_PRBS_MODE                     (PCS_CH1_RX_PRBS_MODE),             
    .CP_PCS_CH1_RX_ERRCNT_CLR                    (PCS_CH1_RX_ERRCNT_CLR),            
    .CP_PCS_CH1_TX_PRBS_MODE                     (PCS_CH1_TX_PRBS_MODE),             
    .CP_PCS_CH1_TX_INSERT_ER                     (PCS_CH1_TX_INSERT_ER),             
    .CP_PCS_CH1_ENABLE_PRBS_GEN                  (PCS_CH1_ENABLE_PRBS_GEN),          
    .CP_PCS_CH1_ERR_CNT                          (PCS_CH1_ERR_CNT),                  
    .CP_PCS_CH1_DEFAULT_RADDR                    (PCS_CH1_DEFAULT_RADDR),            
    .CP_PCS_CH1_MASTER_CHECK_OFFSET              (PCS_CH1_MASTER_CHECK_OFFSET),      
    .CP_PCS_CH1_DELAY_SET                        (PCS_CH1_DELAY_SET),                
    .CP_PCS_CH1_SEACH_OFFSET                     (PCS_CH1_SEACH_OFFSET),             
    .CP_PCS_CH1_CEB_RAPIDLS_MMAX                 (PCS_CH1_CEB_RAPIDLS_MMAX),         
    .CP_PCS_CH1_CTC_AFULL                        (PCS_CH1_CTC_AFULL),                
    .CP_PCS_CH1_CTC_AEMPTY                       (PCS_CH1_CTC_AEMPTY),               
    .CP_PCS_CH1_CTC_CONTI_SKP_SET                (PCS_CH1_CTC_CONTI_SKP_SET),        
    .CP_PCS_CH1_FAR_LOOP                         (PCS_CH1_FAR_LOOP),                 
    .CP_PCS_CH1_NEAR_LOOP                        (PCS_CH1_NEAR_LOOP),                
    .CP_PCS_CH1_INT_RX_MASK_0                    (PCS_CH1_INT_RX_MASK_0),         
    .CP_PCS_CH1_INT_RX_MASK_1                    (PCS_CH1_INT_RX_MASK_1),         
    .CP_PCS_CH1_INT_RX_MASK_2                    (PCS_CH1_INT_RX_MASK_2),         
    .CP_PCS_CH1_INT_RX_MASK_3                    (PCS_CH1_INT_RX_MASK_3),         
    .CP_PCS_CH1_INT_RX_MASK_4                    (PCS_CH1_INT_RX_MASK_4),         
    .CP_PCS_CH1_INT_RX_MASK_5                    (PCS_CH1_INT_RX_MASK_5),         
    .CP_PCS_CH1_INT_RX_MASK_6                    (PCS_CH1_INT_RX_MASK_6),         
    .CP_PCS_CH1_INT_RX_MASK_7                    (PCS_CH1_INT_RX_MASK_7),         
    .CP_PCS_CH1_INT_RX_CLR_0                     (PCS_CH1_INT_RX_CLR_0),          
    .CP_PCS_CH1_INT_RX_CLR_1                     (PCS_CH1_INT_RX_CLR_1),          
    .CP_PCS_CH1_INT_RX_CLR_2                     (PCS_CH1_INT_RX_CLR_2),          
    .CP_PCS_CH1_INT_RX_CLR_3                     (PCS_CH1_INT_RX_CLR_3),          
    .CP_PCS_CH1_INT_RX_CLR_4                     (PCS_CH1_INT_RX_CLR_4),          
    .CP_PCS_CH1_INT_RX_CLR_5                     (PCS_CH1_INT_RX_CLR_5),          
    .CP_PCS_CH1_INT_RX_CLR_6                     (PCS_CH1_INT_RX_CLR_6),          
    .CP_PCS_CH1_INT_RX_CLR_7                     (PCS_CH1_INT_RX_CLR_7),          
    .CP_PCS_CH2_BYPASS_WORD_ALIGN                (PCS_CH2_BYPASS_WORD_ALIGN),    
    .CP_PCS_CH2_BYPASS_DENC                      (PCS_CH2_BYPASS_DENC),          
    .CP_PCS_CH2_BYPASS_BONDING                   (PCS_CH2_BYPASS_BONDING),       
    .CP_PCS_CH2_BYPASS_CTC                       (PCS_CH2_BYPASS_CTC),           
    .CP_PCS_CH2_BYPASS_GEAR                      (PCS_CH2_BYPASS_GEAR),          
    .CP_PCS_CH2_BYPASS_BRIDGE                    (PCS_CH2_BYPASS_BRIDGE),        
    .CP_PCS_CH2_DATA_MODE                        (PCS_CH2_DATA_MODE),            
    .CP_PCS_CH2_RX_POLARITY_INV                  (PCS_CH2_RX_POLARITY_INV),      
    .CP_PCS_CH2_ALIGN_MODE                       (PCS_CH2_ALIGN_MODE),           
    .CP_PCS_CH2_SAMP_16B                         (PCS_CH2_SAMP_16B),             
    .CP_PCS_CH2_COMMA_REG0                       (PCS_CH2_COMMA_REG0),           
    .CP_PCS_CH2_COMMA_MASK                       (PCS_CH2_COMMA_MASK),           
    .CP_PCS_CH2_CEB_MODE                         (PCS_CH2_CEB_MODE),             
    .CP_PCS_CH2_CTC_MODE                         (PCS_CH2_CTC_MODE),             
    .CP_PCS_CH2_A_REG                            (PCS_CH2_A_REG),                
    .CP_PCS_CH2_GE_AUTO_EN                       (PCS_CH2_GE_AUTO_EN),           
    .CP_PCS_CH2_SKIP_REG0                        (PCS_CH2_SKIP_REG0),            
    .CP_PCS_CH2_SKIP_REG1                        (PCS_CH2_SKIP_REG1),            
    .CP_PCS_CH2_SKIP_REG2                        (PCS_CH2_SKIP_REG2),            
    .CP_PCS_CH2_SKIP_REG3                        (PCS_CH2_SKIP_REG3),            
    .CP_PCS_CH2_DEC_DUAL                         (PCS_CH2_DEC_DUAL),             
    .CP_PCS_CH2_SPLIT                            (PCS_CH2_SPLIT),                
    .CP_PCS_CH2_FIFOFLAG_CTC                     (PCS_CH2_FIFOFLAG_CTC),         
    .CP_PCS_CH2_COMMA_DET_MODE                   (PCS_CH2_COMMA_DET_MODE),       
    .CP_PCS_CH2_ERRDETECT_SILENCE                (PCS_CH2_ERRDETECT_SILENCE),    
    .CP_PCS_CH2_PMA_RCLK_POLINV                  (PCS_CH2_PMA_RCLK_POLINV),      
    .CP_PCS_CH2_PCS_RCLK_SEL                     (PCS_CH2_PCS_RCLK_SEL),         
    .CP_PCS_CH2_MCB_RCLK_POLINV                  (PCS_CH2_MCB_RCLK_POLINV),        
    .CP_PCS_CH2_CB_RCLK_SEL                      (PCS_CH2_CB_RCLK_SEL),            
    .CP_PCS_CH2_AFTER_CTC_RCLK_SEL               (PCS_CH2_AFTER_CTC_RCLK_SEL),   
    .CP_PCS_CH2_RCLK_POLINV                      (PCS_CH2_RCLK_POLINV),          
    .CP_PCS_CH2_BRIDGE_RCLK_SEL                  (PCS_CH2_BRIDGE_RCLK_SEL),      
    .CP_PCS_CH2_PCS_RCLK_EN                      (PCS_CH2_PCS_RCLK_EN),          
    .CP_PCS_CH2_CB_RCLK_EN                       (PCS_CH2_CB_RCLK_EN),           
    .CP_PCS_CH2_AFTER_CTC_RCLK_EN                (PCS_CH2_AFTER_CTC_RCLK_EN),    
    .CP_PCS_CH2_AFTER_CTC_RCLK_EN_GB             (PCS_CH2_AFTER_CTC_RCLK_EN_GB), 
    .CP_PCS_CH2_BRIDGE_RCLK_EN                   (PCS_CH2_BRIDGE_RCLK_EN),       
    .CP_PCS_CH2_PCS_RX_RSTN                      (PCS_CH2_PCS_RX_RSTN),          
    .CP_PCS_CH2_SLAVE                            (PCS_CH2_SLAVE),                
    .CP_PCS_CH2_PCIE_SLAVE                       (PCS_CH2_PCIE_SLAVE),           
    .CP_PCS_CH2_PCS_CB_RSTN                      (PCS_CH2_PCS_CB_RSTN),          
    .CP_PCS_CH2_TX_BYPASS_BRIDGE_UINT            (PCS_CH2_TX_BYPASS_BRIDGE_UINT),
    .CP_PCS_CH2_TX_BYPASS_GEAR                   (PCS_CH2_TX_BYPASS_GEAR),       
    .CP_PCS_CH2_TX_BYPASS_ENC                    (PCS_CH2_TX_BYPASS_ENC),        
    .CP_PCS_CH2_TX_BYPASS_BIT_SLIP               (PCS_CH2_TX_BYPASS_BIT_SLIP),   
    .CP_PCS_CH2_TX_GEAR_SPLIT                    (PCS_CH2_TX_GEAR_SPLIT),        
    .CP_PCS_CH2_TX_DRIVE_REG_MODE                (PCS_CH2_TX_DRIVE_REG_MODE),    
    .CP_PCS_CH2_TX_BIT_SLIP_CYCLES               (PCS_CH2_TX_BIT_SLIP_CYCLES),   
    .CP_PCS_CH2_INT_TX_MASK_0                    (PCS_CH2_INT_TX_MASK_0),        
    .CP_PCS_CH2_INT_TX_MASK_1                    (PCS_CH2_INT_TX_MASK_1),        
    .CP_PCS_CH2_INT_TX_MASK_2                    (PCS_CH2_INT_TX_MASK_2),          
    .CP_PCS_CH2_INT_TX_CLR_0                     (PCS_CH2_INT_TX_CLR_0),           
    .CP_PCS_CH2_INT_TX_CLR_1                     (PCS_CH2_INT_TX_CLR_1),           
    .CP_PCS_CH2_INT_TX_CLR_2                     (PCS_CH2_INT_TX_CLR_2),                
    .CP_PCS_CH2_TX_PMA_TCLK_POLINV               (PCS_CH2_TX_PMA_TCLK_POLINV),     
    .CP_PCS_CH2_TX_PCS_CLK_EN_SEL                (PCS_CH2_TX_PCS_CLK_EN_SEL),        
    .CP_PCS_CH2_TX_BRIDGE_TCLK_SEL               (PCS_CH2_TX_BRIDGE_TCLK_SEL),         
    .CP_PCS_CH2_TX_TCLK_POLINV                   (PCS_CH2_TX_TCLK_POLINV),           
    .CP_PCS_CH2_TX_PCS_TX_RSTN                   (PCS_CH2_TX_PCS_TX_RSTN),         
    .CP_PCS_CH2_TX_SLAVE                         (PCS_CH2_TX_SLAVE),               
    .CP_PCS_CH2_TX_BRIDGE_CLK_EN_SEL             (PCS_CH2_TX_BRIDGE_CLK_EN_SEL),     
    .CP_PCS_CH2_DATA_WIDTH_MODE                  (PCS_CH2_DATA_WIDTH_MODE),        
    .CP_PCS_CH2_TX_TCLK2FABRIC_SEL               (PCS_CH2_TX_TCLK2FABRIC_SEL),      
    .CP_PCS_CH2_TX_OUTZZ                         (PCS_CH2_TX_OUTZZ),                
    .CP_PCS_CH2_ENC_DUAL                         (PCS_CH2_ENC_DUAL),                 
    .CP_PCS_CH2_TX_BITSLIP_DATA_MODE             (PCS_CH2_TX_BITSLIP_DATA_MODE),      
    .CP_PCS_CH2_COMMA_REG1                       (PCS_CH2_COMMA_REG1),                
    .CP_PCS_CH2_RAPID_IMAX                       (PCS_CH2_RAPID_IMAX),               
    .CP_PCS_CH2_RAPID_VMIN_1                     (PCS_CH2_RAPID_VMIN_1),              
    .CP_PCS_CH2_RAPID_VMIN_2                     (PCS_CH2_RAPID_VMIN_2),             
    .CP_PCS_CH2_RX_PRBS_MODE                     (PCS_CH2_RX_PRBS_MODE),            
    .CP_PCS_CH2_RX_ERRCNT_CLR                    (PCS_CH2_RX_ERRCNT_CLR),           
    .CP_PCS_CH2_TX_PRBS_MODE                     (PCS_CH2_TX_PRBS_MODE),             
    .CP_PCS_CH2_TX_INSERT_ER                     (PCS_CH2_TX_INSERT_ER),            
    .CP_PCS_CH2_ENABLE_PRBS_GEN                  (PCS_CH2_ENABLE_PRBS_GEN),          
    .CP_PCS_CH2_ERR_CNT                          (PCS_CH2_ERR_CNT),                 
    .CP_PCS_CH2_DEFAULT_RADDR                    (PCS_CH2_DEFAULT_RADDR),            
    .CP_PCS_CH2_MASTER_CHECK_OFFSET              (PCS_CH2_MASTER_CHECK_OFFSET),       
    .CP_PCS_CH2_DELAY_SET                        (PCS_CH2_DELAY_SET),               
    .CP_PCS_CH2_SEACH_OFFSET                     (PCS_CH2_SEACH_OFFSET),          
    .CP_PCS_CH2_CEB_RAPIDLS_MMAX                 (PCS_CH2_CEB_RAPIDLS_MMAX),            
    .CP_PCS_CH2_CTC_AFULL                        (PCS_CH2_CTC_AFULL),            
    .CP_PCS_CH2_CTC_AEMPTY                       (PCS_CH2_CTC_AEMPTY),            
    .CP_PCS_CH2_CTC_CONTI_SKP_SET                (PCS_CH2_CTC_CONTI_SKP_SET),      
    .CP_PCS_CH2_FAR_LOOP                         (PCS_CH2_FAR_LOOP),                        
    .CP_PCS_CH2_NEAR_LOOP                        (PCS_CH2_NEAR_LOOP),              
    .CP_PCS_CH2_INT_RX_MASK_0                    (PCS_CH2_INT_RX_MASK_0),         
    .CP_PCS_CH2_INT_RX_MASK_1                    (PCS_CH2_INT_RX_MASK_1),          
    .CP_PCS_CH2_INT_RX_MASK_2                    (PCS_CH2_INT_RX_MASK_2),         
    .CP_PCS_CH2_INT_RX_MASK_3                    (PCS_CH2_INT_RX_MASK_3),        
    .CP_PCS_CH2_INT_RX_MASK_4                    (PCS_CH2_INT_RX_MASK_4),             
    .CP_PCS_CH2_INT_RX_MASK_5                    (PCS_CH2_INT_RX_MASK_5),             
    .CP_PCS_CH2_INT_RX_MASK_6                    (PCS_CH2_INT_RX_MASK_6),             
    .CP_PCS_CH2_INT_RX_MASK_7                    (PCS_CH2_INT_RX_MASK_7),                 
    .CP_PCS_CH2_INT_RX_CLR_0                     (PCS_CH2_INT_RX_CLR_0),           
    .CP_PCS_CH2_INT_RX_CLR_1                     (PCS_CH2_INT_RX_CLR_1),               
    .CP_PCS_CH2_INT_RX_CLR_2                     (PCS_CH2_INT_RX_CLR_2),          
    .CP_PCS_CH2_INT_RX_CLR_3                     (PCS_CH2_INT_RX_CLR_3),         
    .CP_PCS_CH2_INT_RX_CLR_4                     (PCS_CH2_INT_RX_CLR_4),         
    .CP_PCS_CH2_INT_RX_CLR_5                     (PCS_CH2_INT_RX_CLR_5),             
    .CP_PCS_CH2_INT_RX_CLR_6                     (PCS_CH2_INT_RX_CLR_6),             
    .CP_PCS_CH2_INT_RX_CLR_7                     (PCS_CH2_INT_RX_CLR_7),            
    .CP_PCS_CH3_BYPASS_WORD_ALIGN                (PCS_CH3_BYPASS_WORD_ALIGN),     
    .CP_PCS_CH3_BYPASS_DENC                      (PCS_CH3_BYPASS_DENC),            
    .CP_PCS_CH3_BYPASS_BONDING                   (PCS_CH3_BYPASS_BONDING),          
    .CP_PCS_CH3_BYPASS_CTC                       (PCS_CH3_BYPASS_CTC),            
    .CP_PCS_CH3_BYPASS_GEAR                      (PCS_CH3_BYPASS_GEAR),                   
    .CP_PCS_CH3_BYPASS_BRIDGE                    (PCS_CH3_BYPASS_BRIDGE),          
    .CP_PCS_CH3_DATA_MODE                        (PCS_CH3_DATA_MODE),               
    .CP_PCS_CH3_RX_POLARITY_INV                  (PCS_CH3_RX_POLARITY_INV),       
    .CP_PCS_CH3_ALIGN_MODE                       (PCS_CH3_ALIGN_MODE),              
    .CP_PCS_CH3_SAMP_16B                         (PCS_CH3_SAMP_16B),                
    .CP_PCS_CH3_COMMA_REG0                       (PCS_CH3_COMMA_REG0),            
    .CP_PCS_CH3_COMMA_MASK                       (PCS_CH3_COMMA_MASK),              
    .CP_PCS_CH3_CEB_MODE                         (PCS_CH3_CEB_MODE),             
    .CP_PCS_CH3_CTC_MODE                         (PCS_CH3_CTC_MODE),              
    .CP_PCS_CH3_A_REG                            (PCS_CH3_A_REG),                  
    .CP_PCS_CH3_GE_AUTO_EN                       (PCS_CH3_GE_AUTO_EN),            
    .CP_PCS_CH3_SKIP_REG0                        (PCS_CH3_SKIP_REG0),            
    .CP_PCS_CH3_SKIP_REG1                        (PCS_CH3_SKIP_REG1),            
    .CP_PCS_CH3_SKIP_REG2                        (PCS_CH3_SKIP_REG2),            
    .CP_PCS_CH3_SKIP_REG3                        (PCS_CH3_SKIP_REG3),               
    .CP_PCS_CH3_DEC_DUAL                         (PCS_CH3_DEC_DUAL),               
    .CP_PCS_CH3_SPLIT                            (PCS_CH3_SPLIT),                  
    .CP_PCS_CH3_FIFOFLAG_CTC                     (PCS_CH3_FIFOFLAG_CTC),         
    .CP_PCS_CH3_COMMA_DET_MODE                   (PCS_CH3_COMMA_DET_MODE),               
    .CP_PCS_CH3_ERRDETECT_SILENCE                (PCS_CH3_ERRDETECT_SILENCE),       
    .CP_PCS_CH3_PMA_RCLK_POLINV                  (PCS_CH3_PMA_RCLK_POLINV),          
    .CP_PCS_CH3_PCS_RCLK_SEL                     (PCS_CH3_PCS_RCLK_SEL),         
    .CP_PCS_CH3_MCB_RCLK_POLINV                  (PCS_CH3_MCB_RCLK_POLINV),       
    .CP_PCS_CH3_CB_RCLK_SEL                      (PCS_CH3_CB_RCLK_SEL),            
    .CP_PCS_CH3_AFTER_CTC_RCLK_SEL               (PCS_CH3_AFTER_CTC_RCLK_SEL),      
    .CP_PCS_CH3_RCLK_POLINV                      (PCS_CH3_RCLK_POLINV),           
    .CP_PCS_CH3_BRIDGE_RCLK_SEL                  (PCS_CH3_BRIDGE_RCLK_SEL),       
    .CP_PCS_CH3_PCS_RCLK_EN                      (PCS_CH3_PCS_RCLK_EN),           
    .CP_PCS_CH3_CB_RCLK_EN                       (PCS_CH3_CB_RCLK_EN),            
    .CP_PCS_CH3_AFTER_CTC_RCLK_EN                (PCS_CH3_AFTER_CTC_RCLK_EN),         
    .CP_PCS_CH3_AFTER_CTC_RCLK_EN_GB             (PCS_CH3_AFTER_CTC_RCLK_EN_GB),      
    .CP_PCS_CH3_BRIDGE_RCLK_EN                   (PCS_CH3_BRIDGE_RCLK_EN),           
    .CP_PCS_CH3_PCS_RX_RSTN                      (PCS_CH3_PCS_RX_RSTN),             
    .CP_PCS_CH3_SLAVE                            (PCS_CH3_SLAVE),                    
    .CP_PCS_CH3_PCIE_SLAVE                       (PCS_CH3_PCIE_SLAVE),              
    .CP_PCS_CH3_PCS_CB_RSTN                      (PCS_CH3_PCS_CB_RSTN),           
    .CP_PCS_CH3_TX_BYPASS_BRIDGE_UINT            (PCS_CH3_TX_BYPASS_BRIDGE_UINT),  
    .CP_PCS_CH3_TX_BYPASS_GEAR                   (PCS_CH3_TX_BYPASS_GEAR),        
    .CP_PCS_CH3_TX_BYPASS_ENC                    (PCS_CH3_TX_BYPASS_ENC),            
    .CP_PCS_CH3_TX_BYPASS_BIT_SLIP               (PCS_CH3_TX_BYPASS_BIT_SLIP),       
    .CP_PCS_CH3_TX_GEAR_SPLIT                    (PCS_CH3_TX_GEAR_SPLIT),                    
    .CP_PCS_CH3_TX_DRIVE_REG_MODE                (PCS_CH3_TX_DRIVE_REG_MODE),         
    .CP_PCS_CH3_TX_BIT_SLIP_CYCLES               (PCS_CH3_TX_BIT_SLIP_CYCLES),      
    .CP_PCS_CH3_INT_TX_MASK_0                    (PCS_CH3_INT_TX_MASK_0),        
    .CP_PCS_CH3_INT_TX_MASK_1                    (PCS_CH3_INT_TX_MASK_1),        
    .CP_PCS_CH3_INT_TX_MASK_2                    (PCS_CH3_INT_TX_MASK_2),        
    .CP_PCS_CH3_INT_TX_CLR_0                     (PCS_CH3_INT_TX_CLR_0),         
    .CP_PCS_CH3_INT_TX_CLR_1                     (PCS_CH3_INT_TX_CLR_1),         
    .CP_PCS_CH3_INT_TX_CLR_2                     (PCS_CH3_INT_TX_CLR_2),         
    .CP_PCS_CH3_TX_PMA_TCLK_POLINV               (PCS_CH3_TX_PMA_TCLK_POLINV),        
    .CP_PCS_CH3_TX_PCS_CLK_EN_SEL                (PCS_CH3_TX_PCS_CLK_EN_SEL),         
    .CP_PCS_CH3_TX_BRIDGE_TCLK_SEL               (PCS_CH3_TX_BRIDGE_TCLK_SEL),        
    .CP_PCS_CH3_TX_TCLK_POLINV                   (PCS_CH3_TX_TCLK_POLINV),            
    .CP_PCS_CH3_TX_PCS_TX_RSTN                   (PCS_CH3_TX_PCS_TX_RSTN),            
    .CP_PCS_CH3_TX_SLAVE                         (PCS_CH3_TX_SLAVE),                  
    .CP_PCS_CH3_TX_BRIDGE_CLK_EN_SEL             (PCS_CH3_TX_BRIDGE_CLK_EN_SEL),      
    .CP_PCS_CH3_DATA_WIDTH_MODE                  (PCS_CH3_DATA_WIDTH_MODE),           
    .CP_PCS_CH3_TX_TCLK2FABRIC_SEL               (PCS_CH3_TX_TCLK2FABRIC_SEL),        
    .CP_PCS_CH3_TX_OUTZZ                         (PCS_CH3_TX_OUTZZ),                  
    .CP_PCS_CH3_ENC_DUAL                         (PCS_CH3_ENC_DUAL),                  
    .CP_PCS_CH3_TX_BITSLIP_DATA_MODE             (PCS_CH3_TX_BITSLIP_DATA_MODE),      
    .CP_PCS_CH3_COMMA_REG1                       (PCS_CH3_COMMA_REG1),                
    .CP_PCS_CH3_RAPID_IMAX                       (PCS_CH3_RAPID_IMAX),               
    .CP_PCS_CH3_RAPID_VMIN_1                     (PCS_CH3_RAPID_VMIN_1),             
    .CP_PCS_CH3_RAPID_VMIN_2                     (PCS_CH3_RAPID_VMIN_2),             
    .CP_PCS_CH3_RX_PRBS_MODE                     (PCS_CH3_RX_PRBS_MODE),             
    .CP_PCS_CH3_RX_ERRCNT_CLR                    (PCS_CH3_RX_ERRCNT_CLR),            
    .CP_PCS_CH3_TX_PRBS_MODE                     (PCS_CH3_TX_PRBS_MODE),             
    .CP_PCS_CH3_TX_INSERT_ER                     (PCS_CH3_TX_INSERT_ER),             
    .CP_PCS_CH3_ENABLE_PRBS_GEN                  (PCS_CH3_ENABLE_PRBS_GEN),          
    .CP_PCS_CH3_ERR_CNT                          (PCS_CH3_ERR_CNT),                  
    .CP_PCS_CH3_DEFAULT_RADDR                    (PCS_CH3_DEFAULT_RADDR),             
    .CP_PCS_CH3_MASTER_CHECK_OFFSET              (PCS_CH3_MASTER_CHECK_OFFSET),       
    .CP_PCS_CH3_DELAY_SET                        (PCS_CH3_DELAY_SET),                 
    .CP_PCS_CH3_SEACH_OFFSET                     (PCS_CH3_SEACH_OFFSET),              
    .CP_PCS_CH3_CEB_RAPIDLS_MMAX                 (PCS_CH3_CEB_RAPIDLS_MMAX),          
    .CP_PCS_CH3_CTC_AFULL                        (PCS_CH3_CTC_AFULL),                 
    .CP_PCS_CH3_CTC_AEMPTY                       (PCS_CH3_CTC_AEMPTY),                
    .CP_PCS_CH3_CTC_CONTI_SKP_SET                (PCS_CH3_CTC_CONTI_SKP_SET),         
    .CP_PCS_CH3_FAR_LOOP                         (PCS_CH3_FAR_LOOP),                  
    .CP_PCS_CH3_NEAR_LOOP                        (PCS_CH3_NEAR_LOOP),                 
    .CP_PCS_CH3_INT_RX_MASK_0                    (PCS_CH3_INT_RX_MASK_0),             
    .CP_PCS_CH3_INT_RX_MASK_1                    (PCS_CH3_INT_RX_MASK_1),             
    .CP_PCS_CH3_INT_RX_MASK_2                    (PCS_CH3_INT_RX_MASK_2),             
    .CP_PCS_CH3_INT_RX_MASK_3                    (PCS_CH3_INT_RX_MASK_3),             
    .CP_PCS_CH3_INT_RX_MASK_4                    (PCS_CH3_INT_RX_MASK_4),             
    .CP_PCS_CH3_INT_RX_MASK_5                    (PCS_CH3_INT_RX_MASK_5),             
    .CP_PCS_CH3_INT_RX_MASK_6                    (PCS_CH3_INT_RX_MASK_6),             
    .CP_PCS_CH3_INT_RX_MASK_7                    (PCS_CH3_INT_RX_MASK_7),             
    .CP_PCS_CH3_INT_RX_CLR_0                     (PCS_CH3_INT_RX_CLR_0),              
    .CP_PCS_CH3_INT_RX_CLR_1                     (PCS_CH3_INT_RX_CLR_1),              
    .CP_PCS_CH3_INT_RX_CLR_2                     (PCS_CH3_INT_RX_CLR_2),              
    .CP_PCS_CH3_INT_RX_CLR_3                     (PCS_CH3_INT_RX_CLR_3),              
    .CP_PCS_CH3_INT_RX_CLR_4                     (PCS_CH3_INT_RX_CLR_4),              
    .CP_PCS_CH3_INT_RX_CLR_5                     (PCS_CH3_INT_RX_CLR_5),              
    .CP_PCS_CH3_INT_RX_CLR_6                     (PCS_CH3_INT_RX_CLR_6),              
    .CP_PCS_CH3_INT_RX_CLR_7                     (PCS_CH3_INT_RX_CLR_7),              
    .CP_PMA_CH0_REG_RX_PD                        (PMA_CH0_REG_RX_PD),                  
    .CP_PMA_CH0_REG_RX_PD_EN                     (PMA_CH0_REG_RX_PD_EN),              
    .CP_PMA_CH0_REG_RX_CLKPATH_PD                (PMA_CH0_REG_RX_CLKPATH_PD),         
    .CP_PMA_CH0_REG_RX_CLKPATH_PD_EN             (PMA_CH0_REG_RX_CLKPATH_PD_EN),      
    .CP_PMA_CH0_REG_RX_DATAPATH_PD               (PMA_CH0_REG_RX_DATAPATH_PD),        
    .CP_PMA_CH0_REG_RX_DATAPATH_PD_EN            (PMA_CH0_REG_RX_DATAPATH_PD_EN),     
    .CP_PMA_CH0_REG_RX_SIGDET_PD                 (PMA_CH0_REG_RX_SIGDET_PD),          
    .CP_PMA_CH0_REG_RX_SIGDET_PD_EN              (PMA_CH0_REG_RX_SIGDET_PD_EN),       
    .CP_PMA_CH0_REG_RX_DCC_RST_N                 (PMA_CH0_REG_RX_DCC_RST_N),          
    .CP_PMA_CH0_REG_RX_DCC_RST_N_EN              (PMA_CH0_REG_RX_DCC_RST_N_EN),       
    .CP_PMA_CH0_REG_RX_CDR_RST_N                 (PMA_CH0_REG_RX_CDR_RST_N),          
    .CP_PMA_CH0_REG_RX_CDR_RST_N_EN              (PMA_CH0_REG_RX_CDR_RST_N_EN),       
    .CP_PMA_CH0_REG_RX_SIGDET_RST_N              (PMA_CH0_REG_RX_SIGDET_RST_N),       
    .CP_PMA_CH0_REG_RX_SIGDET_RST_N_EN           (PMA_CH0_REG_RX_SIGDET_RST_N_EN),    
    .CP_PMA_CH0_REG_RXPCLK_SLIP                  (PMA_CH0_REG_RXPCLK_SLIP),           
    .CP_PMA_CH0_REG_RXPCLK_SLIP_OW               (PMA_CH0_REG_RXPCLK_SLIP_OW),        
    .CP_PMA_CH0_REG_RX_PCLKSWITCH_RST_N          (PMA_CH0_REG_RX_PCLKSWITCH_RST_N),   
    .CP_PMA_CH0_REG_RX_PCLKSWITCH_RST_N_EN       (PMA_CH0_REG_RX_PCLKSWITCH_RST_N_EN),
    .CP_PMA_CH0_REG_RX_PCLKSWITCH                (PMA_CH0_REG_RX_PCLKSWITCH),          
    .CP_PMA_CH0_REG_RX_PCLKSWITCH_EN             (PMA_CH0_REG_RX_PCLKSWITCH_EN),       
    .CP_PMA_CH0_REG_RX_HIGHZ                     (PMA_CH0_REG_RX_HIGHZ),               
    .CP_PMA_CH0_REG_RX_HIGHZ_EN                  (PMA_CH0_REG_RX_HIGHZ_EN),            
    .CP_PMA_CH0_REG_RX_EQ_C_SET                  (PMA_CH0_REG_RX_EQ_C_SET),            
    .CP_PMA_CH0_REG_RX_EQ_R_SET                  (PMA_CH0_REG_RX_EQ_R_SET),            
    .CP_PMA_CH0_REG_RX_BUSWIDTH                  (PMA_CH0_REG_RX_BUSWIDTH),            
    .CP_PMA_CH0_REG_RX_BUSWIDTH_EN               (PMA_CH0_REG_RX_BUSWIDTH_EN),         
    .CP_PMA_CH0_REG_RX_RATE                      (PMA_CH0_REG_RX_RATE),                
    .CP_PMA_CH0_REG_RX_RATE_EN                   (PMA_CH0_REG_RX_RATE_EN),             
    .CP_PMA_CH0_REG_RX_RES_TRIM                  (PMA_CH0_REG_RX_RES_TRIM),            
    .CP_PMA_CH0_REG_RX_RES_TRIM_EN               (PMA_CH0_REG_RX_RES_TRIM_EN),         
    .CP_PMA_CH0_REG_RX_EQ_OFF                    (PMA_CH0_REG_RX_EQ_OFF),              
    .CP_PMA_CH0_REG_RX_PREAMP_IC                 (PMA_CH0_REG_RX_PREAMP_IC),           
    .CP_PMA_CH0_REG_RX_PCLK_EDGE_SEL             (PMA_CH0_REG_RX_PCLK_EDGE_SEL),       
    .CP_PMA_CH0_REG_RX_PIBUF_IC                  (PMA_CH0_REG_RX_PIBUF_IC),            
    .CP_PMA_CH0_REG_RX_DCC_IC_RX                 (PMA_CH0_REG_RX_DCC_IC_RX),           
    .CP_PMA_CH0_REG_RX_DCC_IC_TX                 (PMA_CH0_REG_RX_DCC_IC_TX),           
    .CP_PMA_CH0_REG_RX_ICTRL_TRX                 (PMA_CH0_REG_RX_ICTRL_TRX),           
    .CP_PMA_CH0_REG_RX_ICTRL_SIGDET              (PMA_CH0_REG_RX_ICTRL_SIGDET),        
    .CP_PMA_CH0_REG_RX_ICTRL_PREAMP              (PMA_CH0_REG_RX_ICTRL_PREAMP),        
    .CP_PMA_CH0_REG_RX_ICTRL_SLICER              (PMA_CH0_REG_RX_ICTRL_SLICER),        
    .CP_PMA_CH0_REG_RX_ICTRL_PIBUF               (PMA_CH0_REG_RX_ICTRL_PIBUF),         
    .CP_PMA_CH0_REG_RX_ICTRL_PI                  (PMA_CH0_REG_RX_ICTRL_PI),            
    .CP_PMA_CH0_REG_RX_ICTRL_DCC                 (PMA_CH0_REG_RX_ICTRL_DCC),           
    .CP_PMA_CH0_REG_RX_ICTRL_PREDRV              (PMA_CH0_REG_RX_ICTRL_PREDRV),        
    .CP_PMA_CH0_REG_TX_RATE                      (PMA_CH0_REG_TX_RATE),                
    .CP_PMA_CH0_REG_TX_RATE_EN                   (PMA_CH0_REG_TX_RATE_EN),             
    .CP_PMA_CH0_REG_RX_TX2RX_PLPBK_RST_N         (PMA_CH0_REG_RX_TX2RX_PLPBK_RST_N),   
    .CP_PMA_CH0_REG_RX_TX2RX_PLPBK_RST_N_EN      (PMA_CH0_REG_RX_TX2RX_PLPBK_RST_N_EN),
    .CP_PMA_CH0_REG_RX_TX2RX_PLPBK_EN            (PMA_CH0_REG_RX_TX2RX_PLPBK_EN),          
    .CP_PMA_CH0_REG_TXCLK_SEL                    (PMA_CH0_REG_TXCLK_SEL),                  
    .CP_PMA_CH0_REG_RX_DATA_POLARITY             (PMA_CH0_REG_RX_DATA_POLARITY),           
    .CP_PMA_CH0_REG_RX_ERR_INSERT                (PMA_CH0_REG_RX_ERR_INSERT),             
    .CP_PMA_CH0_REG_UDP_CHK_EN                   (PMA_CH0_REG_UDP_CHK_EN),                 
    .CP_PMA_CH0_REG_PRBS_SEL                     (PMA_CH0_REG_PRBS_SEL),                   
    .CP_PMA_CH0_REG_PRBS_CHK_EN                  (PMA_CH0_REG_PRBS_CHK_EN),                
    .CP_PMA_CH0_REG_PRBS_CHK_WIDTH_SEL           (PMA_CH0_REG_PRBS_CHK_WIDTH_SEL),         
    .CP_PMA_CH0_REG_BIST_CHK_PAT_SEL             (PMA_CH0_REG_BIST_CHK_PAT_SEL),           
    .CP_PMA_CH0_REG_LOAD_ERR_CNT                 (PMA_CH0_REG_LOAD_ERR_CNT),               
    .CP_PMA_CH0_REG_CHK_COUNTER_EN               (PMA_CH0_REG_CHK_COUNTER_EN),             
    .CP_PMA_CH0_REG_CDR_PROP_GAIN                (PMA_CH0_REG_CDR_PROP_GAIN),              
    .CP_PMA_CH0_REG_CDR_PROP_TURBO_GAIN          (PMA_CH0_REG_CDR_PROP_TURBO_GAIN),        
    .CP_PMA_CH0_REG_CDR_INT_GAIN                 (PMA_CH0_REG_CDR_INT_GAIN),               
    .CP_PMA_CH0_REG_CDR_INT_TURBO_GAIN           (PMA_CH0_REG_CDR_INT_TURBO_GAIN),         
    .CP_PMA_CH0_REG_CDR_INT_SAT_MAX              (PMA_CH0_REG_CDR_INT_SAT_MAX),            
    .CP_PMA_CH0_REG_CDR_INT_SAT_MIN              (PMA_CH0_REG_CDR_INT_SAT_MIN),            
    .CP_PMA_CH0_REG_CDR_INT_RST                  (PMA_CH0_REG_CDR_INT_RST),                
    .CP_PMA_CH0_REG_CDR_INT_RST_OW               (PMA_CH0_REG_CDR_INT_RST_OW),             
    .CP_PMA_CH0_REG_CDR_PROP_RST                 (PMA_CH0_REG_CDR_PROP_RST),               
    .CP_PMA_CH0_REG_CDR_PROP_RST_OW              (PMA_CH0_REG_CDR_PROP_RST_OW),            
    .CP_PMA_CH0_REG_CDR_LOCK_RST                 (PMA_CH0_REG_CDR_LOCK_RST),               
    .CP_PMA_CH0_REG_CDR_LOCK_RST_OW              (PMA_CH0_REG_CDR_LOCK_RST_OW),            
    .CP_PMA_CH0_REG_CDR_RX_PI_FORCE_SEL          (PMA_CH0_REG_CDR_RX_PI_FORCE_SEL),        
    .CP_PMA_CH0_REG_CDR_RX_PI_FORCE_D            (PMA_CH0_REG_CDR_RX_PI_FORCE_D),          
    .CP_PMA_CH0_REG_CDR_LOCK_TIMER               (PMA_CH0_REG_CDR_LOCK_TIMER),             
    .CP_PMA_CH0_REG_CDR_TURBO_MODE_TIMER         (PMA_CH0_REG_CDR_TURBO_MODE_TIMER),       
    .CP_PMA_CH0_REG_CDR_LOCK_VAL                 (PMA_CH0_REG_CDR_LOCK_VAL),               
    .CP_PMA_CH0_REG_CDR_LOCK_OW                  (PMA_CH0_REG_CDR_LOCK_OW),                
    .CP_PMA_CH0_REG_CDR_INT_SAT_DET_EN           (PMA_CH0_REG_CDR_INT_SAT_DET_EN),         
    .CP_PMA_CH0_REG_CDR_SAT_DET_STATUS_EN        (PMA_CH0_REG_CDR_SAT_DET_STATUS_EN),      
    .CP_PMA_CH0_REG_CDR_SAT_DET_STATUS_RESET_EN  (PMA_CH0_REG_CDR_SAT_DET_STATUS_RESET_EN),
    .CP_PMA_CH0_REG_CDR_PI_CTRL_RST              (PMA_CH0_REG_CDR_PI_CTRL_RST),              
    .CP_PMA_CH0_REG_CDR_PI_CTRL_RST_OW           (PMA_CH0_REG_CDR_PI_CTRL_RST_OW),           
    .CP_PMA_CH0_REG_CDR_SAT_DET_RST              (PMA_CH0_REG_CDR_SAT_DET_RST),              
    .CP_PMA_CH0_REG_CDR_SAT_DET_RST_OW           (PMA_CH0_REG_CDR_SAT_DET_RST_OW),           
    .CP_PMA_CH0_REG_CDR_SAT_DET_STICKY_RST       (PMA_CH0_REG_CDR_SAT_DET_STICKY_RST),       
    .CP_PMA_CH0_REG_CDR_SAT_DET_STICKY_RST_OW    (PMA_CH0_REG_CDR_SAT_DET_STICKY_RST_OW),    
    .CP_PMA_CH0_REG_CDR_SIGDET_STATUS_DIS        (PMA_CH0_REG_CDR_SIGDET_STATUS_DIS),        
    .CP_PMA_CH0_REG_CDR_SAT_DET_TIMER            (PMA_CH0_REG_CDR_SAT_DET_TIMER),            
    .CP_PMA_CH0_REG_CDR_SAT_DET_STATUS_VAL       (PMA_CH0_REG_CDR_SAT_DET_STATUS_VAL),       
    .CP_PMA_CH0_REG_CDR_SAT_DET_STATUS_OW        (PMA_CH0_REG_CDR_SAT_DET_STATUS_OW),        
    .CP_PMA_CH0_REG_CDR_TURBO_MODE_EN            (PMA_CH0_REG_CDR_TURBO_MODE_EN),            
    .CP_PMA_CH0_REG_CDR_STATUS_RADDR_INIT        (PMA_CH0_REG_CDR_STATUS_RADDR_INIT),        
    .CP_PMA_CH0_REG_CDR_STATUS_FIFO_EN           (PMA_CH0_REG_CDR_STATUS_FIFO_EN),           
    .CP_PMA_CH0_REG_PMA_TEST_SEL                 (PMA_CH0_REG_PMA_TEST_SEL),                 
    .CP_PMA_CH0_REG_OOB_COMWAKE_GAP_MIN          (PMA_CH0_REG_OOB_COMWAKE_GAP_MIN),          
    .CP_PMA_CH0_REG_OOB_COMWAKE_GAP_MAX          (PMA_CH0_REG_OOB_COMWAKE_GAP_MAX),          
    .CP_PMA_CH0_REG_OOB_COMINIT_GAP_MIN          (PMA_CH0_REG_OOB_COMINIT_GAP_MIN),          
    .CP_PMA_CH0_REG_OOB_COMINIT_GAP_MAX          (PMA_CH0_REG_OOB_COMINIT_GAP_MAX),          
    .CP_PMA_CH0_REG_RX_PIBUF_IC_TX               (PMA_CH0_REG_RX_PIBUF_IC_TX),               
    .CP_PMA_CH0_REG_COMWAKE_STATUS_CLEAR         (PMA_CH0_REG_COMWAKE_STATUS_CLEAR),         
    .CP_PMA_CH0_REG_COMINIT_STATUS_CLEAR         (PMA_CH0_REG_COMINIT_STATUS_CLEAR),         
    .CP_PMA_CH0_REG_RX_SYNC_RST_N_EN             (PMA_CH0_REG_RX_SYNC_RST_N_EN),             
    .CP_PMA_CH0_REG_RX_SYNC_RST_N                (PMA_CH0_REG_RX_SYNC_RST_N),                
    .CP_PMA_CH0_REG_RX_SATA_COMINIT_OW           (PMA_CH0_REG_RX_SATA_COMINIT_OW),           
    .CP_PMA_CH0_REG_RX_SATA_COMINIT              (PMA_CH0_REG_RX_SATA_COMINIT),              
    .CP_PMA_CH0_REG_RX_SATA_COMWAKE_OW           (PMA_CH0_REG_RX_SATA_COMWAKE_OW),           
    .CP_PMA_CH0_REG_RX_SATA_COMWAKE              (PMA_CH0_REG_RX_SATA_COMWAKE),              
    .CP_PMA_CH0_REG_RX_DCC_DISABLE               (PMA_CH0_REG_RX_DCC_DISABLE),               
    .CP_PMA_CH0_REG_TX_DCC_DISABLE               (PMA_CH0_REG_TX_DCC_DISABLE),               
    .CP_PMA_CH0_REG_RX_SLIP_SEL_EN               (PMA_CH0_REG_RX_SLIP_SEL_EN),               
    .CP_PMA_CH0_REG_RX_SLIP_SEL                  (PMA_CH0_REG_RX_SLIP_SEL),                  
    .CP_PMA_CH0_REG_RX_SLIP_EN                   (PMA_CH0_REG_RX_SLIP_EN),                   
    .CP_PMA_CH0_REG_RX_SIGDET_STATUS_SEL         (PMA_CH0_REG_RX_SIGDET_STATUS_SEL),         
    .CP_PMA_CH0_REG_RX_SIGDET_FSM_RST_N          (PMA_CH0_REG_RX_SIGDET_FSM_RST_N),          
    .CP_PMA_CH0_REG_RX_SIGDET_STATUS_OW          (PMA_CH0_REG_RX_SIGDET_STATUS_OW),          
    .CP_PMA_CH0_REG_RX_SIGDET_STATUS             (PMA_CH0_REG_RX_SIGDET_STATUS),             
    .CP_PMA_CH0_REG_RX_SIGDET_VTH                (PMA_CH0_REG_RX_SIGDET_VTH),                
    .CP_PMA_CH0_REG_RX_SIGDET_GRM                (PMA_CH0_REG_RX_SIGDET_GRM),                
    .CP_PMA_CH0_REG_RX_SIGDET_PULSE_EXT          (PMA_CH0_REG_RX_SIGDET_PULSE_EXT),          
    .CP_PMA_CH0_REG_RX_SIGDET_CH2_SEL            (PMA_CH0_REG_RX_SIGDET_CH2_SEL),            
    .CP_PMA_CH0_REG_RX_SIGDET_CH2_CHK_WINDOW     (PMA_CH0_REG_RX_SIGDET_CH2_CHK_WINDOW),     
    .CP_PMA_CH0_REG_RX_SIGDET_CHK_WINDOW_EN      (PMA_CH0_REG_RX_SIGDET_CHK_WINDOW_EN),      
    .CP_PMA_CH0_REG_RX_SIGDET_NOSIG_COUNT_SETTING(PMA_CH0_REG_RX_SIGDET_NOSIG_COUNT_SETTING),
    .CP_PMA_CH0_REG_RX_SIGDET_OOB_DET_COUNT_VAL  (PMA_CH0_REG_RX_SIGDET_OOB_DET_COUNT_VAL),  
    .CP_PMA_CH0_REG_SLIP_FIFO_INV_EN             (PMA_CH0_REG_SLIP_FIFO_INV_EN),             
    .CP_PMA_CH0_REG_SLIP_FIFO_INV                (PMA_CH0_REG_SLIP_FIFO_INV),                
    .CP_PMA_CH0_REG_RX_SIGDET_4OOB_DET_SEL       (PMA_CH0_REG_RX_SIGDET_4OOB_DET_SEL),       
    .CP_PMA_CH0_REG_RX_SIGDET_IC_I               (PMA_CH0_REG_RX_SIGDET_IC_I),               
    .CP_PMA_CH0_REG_RX_OOB_DETECTOR_RESET_N_OW   (PMA_CH0_REG_RX_OOB_DETECTOR_RESET_N_OW),   
    .CP_PMA_CH0_REG_RX_OOB_DETECTOR_RESET_N      (PMA_CH0_REG_RX_OOB_DETECTOR_RESET_N),      
    .CP_PMA_CH0_REG_RX_OOB_DETECTOR_PD_OW        (PMA_CH0_REG_RX_OOB_DETECTOR_PD_OW),        
    .CP_PMA_CH0_REG_RX_OOB_DETECTOR_PD           (PMA_CH0_REG_RX_OOB_DETECTOR_PD),           
    .CP_PMA_CH0_REG_RX_TERM_CM_CTRL              (PMA_CH0_REG_RX_TERM_CM_CTRL),              
    .CP_PMA_CH0_REG_TX_PD                        (PMA_CH0_REG_TX_PD),                        
    .CP_PMA_CH0_REG_TX_PD_OW                     (PMA_CH0_REG_TX_PD_OW),                     
    .CP_PMA_CH0_REG_TX_CLKPATH_PD                (PMA_CH0_REG_TX_CLKPATH_PD),                
    .CP_PMA_CH0_REG_TX_CLKPATH_PD_OW             (PMA_CH0_REG_TX_CLKPATH_PD_OW),             
    .CP_PMA_CH0_REG_TX_BEACON_TIMER_SEL          (PMA_CH0_REG_TX_BEACON_TIMER_SEL),          
    .CP_PMA_CH0_REG_TX_RXDET_REQ_OW              (PMA_CH0_REG_TX_RXDET_REQ_OW),              
    .CP_PMA_CH0_REG_TX_RXDET_REQ                 (PMA_CH0_REG_TX_RXDET_REQ),                 
    .CP_PMA_CH0_REG_TX_BEACON_EN_OW              (PMA_CH0_REG_TX_BEACON_EN_OW),              
    .CP_PMA_CH0_REG_TX_BEACON_EN                 (PMA_CH0_REG_TX_BEACON_EN),                 
    .CP_PMA_CH0_REG_TX_EI_EN_OW                  (PMA_CH0_REG_TX_EI_EN_OW),                  
    .CP_PMA_CH0_REG_TX_EI_EN                     (PMA_CH0_REG_TX_EI_EN),                     
    .CP_PMA_CH0_REG_TX_RES_CAL_EN                (PMA_CH0_REG_TX_RES_CAL_EN),                
    .CP_PMA_CH0_REG_TX_RES_CAL                   (PMA_CH0_REG_TX_RES_CAL),                   
    .CP_PMA_CH0_REG_TX_BIAS_CAL_EN               (PMA_CH0_REG_TX_BIAS_CAL_EN),               
    .CP_PMA_CH0_REG_TX_BIAS_CTRL                 (PMA_CH0_REG_TX_BIAS_CTRL),                 
    .CP_PMA_CH0_REG_TX_RXDET_TIMER_SEL           (PMA_CH0_REG_TX_RXDET_TIMER_SEL),           
    .CP_PMA_CH0_REG_TX_SYNC_OW                   (PMA_CH0_REG_TX_SYNC_OW),                   
    .CP_PMA_CH0_REG_TX_SYNC                      (PMA_CH0_REG_TX_SYNC),                      
    .CP_PMA_CH0_REG_TX_PD_POST                   (PMA_CH0_REG_TX_PD_POST),                   
    .CP_PMA_CH0_REG_TX_PD_POST_OW                (PMA_CH0_REG_TX_PD_POST_OW),                
    .CP_PMA_CH0_REG_TX_RESET_N_OW                (PMA_CH0_REG_TX_RESET_N_OW),                
    .CP_PMA_CH0_REG_TX_RESET_N                   (PMA_CH0_REG_TX_RESET_N),                   
    .CP_PMA_CH0_REG_TX_DCC_RESET_N_OW            (PMA_CH0_REG_TX_DCC_RESET_N_OW),            
    .CP_PMA_CH0_REG_TX_DCC_RESET_N               (PMA_CH0_REG_TX_DCC_RESET_N),               
    .CP_PMA_CH0_REG_TX_BUSWIDTH_OW               (PMA_CH0_REG_TX_BUSWIDTH_OW),               
    .CP_PMA_CH0_REG_TX_BUSWIDTH                  (PMA_CH0_REG_TX_BUSWIDTH),                  
    .CP_PMA_CH0_REG_PLL_READY_OW                 (PMA_CH0_REG_PLL_READY_OW),                 
    .CP_PMA_CH0_REG_PLL_READY                    (PMA_CH0_REG_PLL_READY),                    
    .CP_PMA_CH0_REG_TX_PCLK_SW_OW                (PMA_CH0_REG_TX_PCLK_SW_OW),                
    .CP_PMA_CH0_REG_TX_PCLK_SW                   (PMA_CH0_REG_TX_PCLK_SW),                   
    .CP_PMA_CH0_REG_EI_PCLK_DELAY_SEL            (PMA_CH0_REG_EI_PCLK_DELAY_SEL),            
    .CP_PMA_CH0_REG_TX_DRV01_DAC0                (PMA_CH0_REG_TX_DRV01_DAC0),                
    .CP_PMA_CH0_REG_TX_DRV01_DAC1                (PMA_CH0_REG_TX_DRV01_DAC1),                
    .CP_PMA_CH0_REG_TX_DRV01_DAC2                (PMA_CH0_REG_TX_DRV01_DAC2),                
    .CP_PMA_CH0_REG_TX_DRV00_DAC0                (PMA_CH0_REG_TX_DRV00_DAC0),                
    .CP_PMA_CH0_REG_TX_DRV00_DAC1                (PMA_CH0_REG_TX_DRV00_DAC1),                
    .CP_PMA_CH0_REG_TX_DRV00_DAC2                (PMA_CH0_REG_TX_DRV00_DAC2),                
    .CP_PMA_CH0_REG_TX_AMP0                      (PMA_CH0_REG_TX_AMP0),                      
    .CP_PMA_CH0_REG_TX_AMP1                      (PMA_CH0_REG_TX_AMP1),                      
    .CP_PMA_CH0_REG_TX_AMP2                      (PMA_CH0_REG_TX_AMP2),                      
    .CP_PMA_CH0_REG_TX_AMP3                      (PMA_CH0_REG_TX_AMP3),                      
    .CP_PMA_CH0_REG_TX_AMP4                      (PMA_CH0_REG_TX_AMP4),                      
    .CP_PMA_CH0_REG_TX_MARGIN                    (PMA_CH0_REG_TX_MARGIN),                    
    .CP_PMA_CH0_REG_TX_MARGIN_OW                 (PMA_CH0_REG_TX_MARGIN_OW),                 
    .CP_PMA_CH0_REG_TX_DEEMP                     (PMA_CH0_REG_TX_DEEMP),                     
    .CP_PMA_CH0_REG_TX_DEEMP_OW                  (PMA_CH0_REG_TX_DEEMP_OW),                  
    .CP_PMA_CH0_REG_TX_SWING                     (PMA_CH0_REG_TX_SWING),                     
    .CP_PMA_CH0_REG_TX_SWING_OW                  (PMA_CH0_REG_TX_SWING_OW),                  
    .CP_PMA_CH0_REG_TX_RXDET_THRESHOLD           (PMA_CH0_REG_TX_RXDET_THRESHOLD),           
    .CP_PMA_CH0_REG_TX_BEACON_OSC_CTRL           (PMA_CH0_REG_TX_BEACON_OSC_CTRL),           
    .CP_PMA_CH0_REG_TX_PREDRV_DAC                (PMA_CH0_REG_TX_PREDRV_DAC),                
    .CP_PMA_CH0_REG_TX_PREDRV_CM_CTRL            (PMA_CH0_REG_TX_PREDRV_CM_CTRL),            
    .CP_PMA_CH0_REG_TX_TX2RX_SLPBACK_EN          (PMA_CH0_REG_TX_TX2RX_SLPBACK_EN),          
    .CP_PMA_CH0_REG_TX_PCLK_EDGE_SEL             (PMA_CH0_REG_TX_PCLK_EDGE_SEL),             
    .CP_PMA_CH0_REG_TX_RXDET_STATUS_OW           (PMA_CH0_REG_TX_RXDET_STATUS_OW),           
    .CP_PMA_CH0_REG_TX_RXDET_STATUS              (PMA_CH0_REG_TX_RXDET_STATUS),              
    .CP_PMA_CH0_REG_TX_PRBS_GEN_EN               (PMA_CH0_REG_TX_PRBS_GEN_EN),               
    .CP_PMA_CH0_REG_TX_PRBS_GEN_WIDTH_SEL        (PMA_CH0_REG_TX_PRBS_GEN_WIDTH_SEL),        
    .CP_PMA_CH0_REG_TX_PRBS_SEL                  (PMA_CH0_REG_TX_PRBS_SEL),                  
    .CP_PMA_CH0_REG_TX_UDP_DATA                  (PMA_CH0_REG_TX_UDP_DATA),                  
    .CP_PMA_CH0_REG_TX_FIFO_RST_N                (PMA_CH0_REG_TX_FIFO_RST_N),                
    .CP_PMA_CH0_REG_TX_FIFO_WP_CTRL              (PMA_CH0_REG_TX_FIFO_WP_CTRL),              
    .CP_PMA_CH0_REG_TX_FIFO_EN                   (PMA_CH0_REG_TX_FIFO_EN),                   
    .CP_PMA_CH0_REG_TX_DATA_MUX_SEL              (PMA_CH0_REG_TX_DATA_MUX_SEL),              
    .CP_PMA_CH0_REG_TX_ERR_INSERT                (PMA_CH0_REG_TX_ERR_INSERT),                
    .CP_PMA_CH0_REG_TX_SATA_EN                   (PMA_CH0_REG_TX_SATA_EN),                   
    .CP_PMA_CH0_REG_RATE_CHANGE_TXPCLK_ON_OW     (PMA_CH0_REG_RATE_CHANGE_TXPCLK_ON_OW),     
    .CP_PMA_CH0_REG_RATE_CHANGE_TXPCLK_ON        (PMA_CH0_REG_RATE_CHANGE_TXPCLK_ON),        
    .CP_PMA_CH0_REG_TX_PULLUP_DAC0               (PMA_CH0_REG_TX_PULLUP_DAC0),               
    .CP_PMA_CH0_REG_TX_PULLUP_DAC1               (PMA_CH0_REG_TX_PULLUP_DAC1),               
    .CP_PMA_CH0_REG_TX_PULLUP_DAC2               (PMA_CH0_REG_TX_PULLUP_DAC2),               
    .CP_PMA_CH0_REG_TX_PULLUP_DAC3               (PMA_CH0_REG_TX_PULLUP_DAC3),               
    .CP_PMA_CH0_REG_TX_OOB_DELAY_SEL             (PMA_CH0_REG_TX_OOB_DELAY_SEL),             
    .CP_PMA_CH0_REG_TX_POLARITY                  (PMA_CH0_REG_TX_POLARITY),                  
    .CP_PMA_CH0_REG_TX_SLPBK_AMP                 (PMA_CH0_REG_TX_SLPBK_AMP),                 
    .CP_PMA_CH0_REG_TX_LS_MODE_EN                (PMA_CH0_REG_TX_LS_MODE_EN),                
    .CP_PMA_CH0_REG_TX_JTAG_MODE_EN_OW           (PMA_CH0_REG_TX_JTAG_MODE_EN_OW),           
    .CP_PMA_CH0_REG_TX_JTAG_MODE_EN              (PMA_CH0_REG_TX_JTAG_MODE_EN),              
    .CP_PMA_CH0_REG_RX_JTAG_MODE_EN_OW           (PMA_CH0_REG_RX_JTAG_MODE_EN_OW),           
    .CP_PMA_CH0_REG_RX_JTAG_MODE_EN              (PMA_CH0_REG_RX_JTAG_MODE_EN),              
    .CP_PMA_CH0_REG_RX_JTAG_OE                   (PMA_CH0_REG_RX_JTAG_OE),                   
    .CP_PMA_CH0_REG_RX_ACJTAG_VHYSTSE            (PMA_CH0_REG_RX_ACJTAG_VHYSTSE),            
    .CP_PMA_CH0_REG_TX_FBCLK_FAR_EN              (PMA_CH0_REG_TX_FBCLK_FAR_EN),              
    .CP_PMA_CH0_REG_RX_TERM_MODE_CTRL            (PMA_CH0_REG_RX_TERM_MODE_CTRL),            
    .CP_PMA_CH0_REG_PLPBK_TXPCLK_EN              (PMA_CH0_REG_PLPBK_TXPCLK_EN),              
    .CP_PMA_CH0_CFG_LANE_POWERUP                 (PMA_CH0_CFG_LANE_POWERUP),                 
    .CP_PMA_CH0_CFG_PMA_POR_N                    (PMA_CH0_CFG_PMA_POR_N),                    
    .CP_PMA_CH0_CFG_RX_LANE_POWERUP              (PMA_CH0_CFG_RX_LANE_POWERUP),              
    .CP_PMA_CH0_CFG_RX_PMA_RSTN                  (PMA_CH0_CFG_RX_PMA_RSTN),                  
    .CP_PMA_CH0_CFG_TX_LANE_POWERUP              (PMA_CH0_CFG_TX_LANE_POWERUP),              
    .CP_PMA_CH0_CFG_TX_PMA_RSTN                  (PMA_CH0_CFG_TX_PMA_RSTN),                  
    .CP_PMA_CH0_REG_RESERVED_48_45               (PMA_CH0_REG_RESERVED_48_45),               
    .CP_PMA_CH0_REG_RESERVED_69                  (PMA_CH0_REG_RESERVED_69),                  
    .CP_PMA_CH0_REG_RESERVED_77_76               (PMA_CH0_REG_RESERVED_77_76),               
    .CP_PMA_CH0_REG_RESERVED_171_164             (PMA_CH0_REG_RESERVED_171_164),             
    .CP_PMA_CH0_REG_RESERVED_175_172             (PMA_CH0_REG_RESERVED_175_172),             
    .CP_PMA_CH0_REG_RESERVED_190                 (PMA_CH0_REG_RESERVED_190),                 
    .CP_PMA_CH0_REG_RESERVED_233_232             (PMA_CH0_REG_RESERVED_233_232),             
    .CP_PMA_CH0_REG_RESERVED_235_234             (PMA_CH0_REG_RESERVED_235_234),             
    .CP_PMA_CH0_REG_RESERVED_241_240             (PMA_CH0_REG_RESERVED_241_240),             
    .CP_PMA_CH0_REG_RESERVED_285_283             (PMA_CH0_REG_RESERVED_285_283),             
    .CP_PMA_CH0_REG_RESERVED_286                 (PMA_CH0_REG_RESERVED_286),                 
    .CP_PMA_CH0_REG_RESERVED_295                 (PMA_CH0_REG_RESERVED_295),                 
    .CP_PMA_CH0_REG_RESERVED_298                 (PMA_CH0_REG_RESERVED_298),                 
    .CP_PMA_CH0_REG_RESERVED_332_325             (PMA_CH0_REG_RESERVED_332_325),             
    .CP_PMA_CH0_REG_RESERVED_340_333             (PMA_CH0_REG_RESERVED_340_333),             
    .CP_PMA_CH0_REG_RESERVED_348_341             (PMA_CH0_REG_RESERVED_348_341),             
    .CP_PMA_CH0_REG_RESERVED_354_349             (PMA_CH0_REG_RESERVED_354_349),             
    .CP_PMA_CH0_REG_RESERVED_373                 (PMA_CH0_REG_RESERVED_373),                 
    .CP_PMA_CH0_REG_RESERVED_376                 (PMA_CH0_REG_RESERVED_376),                 
    .CP_PMA_CH0_REG_RESERVED_452                 (PMA_CH0_REG_RESERVED_452),                 
    .CP_PMA_CH0_REG_RESERVED_502_499             (PMA_CH0_REG_RESERVED_502_499),             
    .CP_PMA_CH0_REG_RESERVED_506_505             (PMA_CH0_REG_RESERVED_506_505),             
    .CP_PMA_CH0_REG_RESERVED_550_549             (PMA_CH0_REG_RESERVED_550_549),             
    .CP_PMA_CH0_REG_RESERVED_556_552             (PMA_CH0_REG_RESERVED_556_552),             
    .CP_PMA_CH1_REG_RX_PD                        (PMA_CH1_REG_RX_PD),                        
    .CP_PMA_CH1_REG_RX_PD_EN                     (PMA_CH1_REG_RX_PD_EN),                     
    .CP_PMA_CH1_REG_RX_CLKPATH_PD                (PMA_CH1_REG_RX_CLKPATH_PD),                
    .CP_PMA_CH1_REG_RX_CLKPATH_PD_EN             (PMA_CH1_REG_RX_CLKPATH_PD_EN),             
    .CP_PMA_CH1_REG_RX_DATAPATH_PD               (PMA_CH1_REG_RX_DATAPATH_PD),               
    .CP_PMA_CH1_REG_RX_DATAPATH_PD_EN            (PMA_CH1_REG_RX_DATAPATH_PD_EN),            
    .CP_PMA_CH1_REG_RX_SIGDET_PD                 (PMA_CH1_REG_RX_SIGDET_PD),                 
    .CP_PMA_CH1_REG_RX_SIGDET_PD_EN              (PMA_CH1_REG_RX_SIGDET_PD_EN),              
    .CP_PMA_CH1_REG_RX_DCC_RST_N                 (PMA_CH1_REG_RX_DCC_RST_N),                 
    .CP_PMA_CH1_REG_RX_DCC_RST_N_EN              (PMA_CH1_REG_RX_DCC_RST_N_EN),              
    .CP_PMA_CH1_REG_RX_CDR_RST_N                 (PMA_CH1_REG_RX_CDR_RST_N),                 
    .CP_PMA_CH1_REG_RX_CDR_RST_N_EN              (PMA_CH1_REG_RX_CDR_RST_N_EN),              
    .CP_PMA_CH1_REG_RX_SIGDET_RST_N              (PMA_CH1_REG_RX_SIGDET_RST_N),              
    .CP_PMA_CH1_REG_RX_SIGDET_RST_N_EN           (PMA_CH1_REG_RX_SIGDET_RST_N_EN),           
    .CP_PMA_CH1_REG_RXPCLK_SLIP                  (PMA_CH1_REG_RXPCLK_SLIP),                  
    .CP_PMA_CH1_REG_RXPCLK_SLIP_OW               (PMA_CH1_REG_RXPCLK_SLIP_OW),               
    .CP_PMA_CH1_REG_RX_PCLKSWITCH_RST_N          (PMA_CH1_REG_RX_PCLKSWITCH_RST_N),          
    .CP_PMA_CH1_REG_RX_PCLKSWITCH_RST_N_EN       (PMA_CH1_REG_RX_PCLKSWITCH_RST_N_EN),       
    .CP_PMA_CH1_REG_RX_PCLKSWITCH                (PMA_CH1_REG_RX_PCLKSWITCH),                
    .CP_PMA_CH1_REG_RX_PCLKSWITCH_EN             (PMA_CH1_REG_RX_PCLKSWITCH_EN),             
    .CP_PMA_CH1_REG_RX_HIGHZ                     (PMA_CH1_REG_RX_HIGHZ),                     
    .CP_PMA_CH1_REG_RX_HIGHZ_EN                  (PMA_CH1_REG_RX_HIGHZ_EN),                  
    .CP_PMA_CH1_REG_RX_EQ_C_SET                  (PMA_CH1_REG_RX_EQ_C_SET),                  
    .CP_PMA_CH1_REG_RX_EQ_R_SET                  (PMA_CH1_REG_RX_EQ_R_SET),                  
    .CP_PMA_CH1_REG_RX_BUSWIDTH                  (PMA_CH1_REG_RX_BUSWIDTH),                  
    .CP_PMA_CH1_REG_RX_BUSWIDTH_EN               (PMA_CH1_REG_RX_BUSWIDTH_EN),               
    .CP_PMA_CH1_REG_RX_RATE                      (PMA_CH1_REG_RX_RATE),                      
    .CP_PMA_CH1_REG_RX_RATE_EN                   (PMA_CH1_REG_RX_RATE_EN),                   
    .CP_PMA_CH1_REG_RX_RES_TRIM                  (PMA_CH1_REG_RX_RES_TRIM),                  
    .CP_PMA_CH1_REG_RX_RES_TRIM_EN               (PMA_CH1_REG_RX_RES_TRIM_EN),               
    .CP_PMA_CH1_REG_RX_EQ_OFF                    (PMA_CH1_REG_RX_EQ_OFF),                    
    .CP_PMA_CH1_REG_RX_PREAMP_IC                 (PMA_CH1_REG_RX_PREAMP_IC),                 
    .CP_PMA_CH1_REG_RX_PCLK_EDGE_SEL             (PMA_CH1_REG_RX_PCLK_EDGE_SEL),             
    .CP_PMA_CH1_REG_RX_PIBUF_IC                  (PMA_CH1_REG_RX_PIBUF_IC),                  
    .CP_PMA_CH1_REG_RX_DCC_IC_RX                 (PMA_CH1_REG_RX_DCC_IC_RX),                 
    .CP_PMA_CH1_REG_RX_DCC_IC_TX                 (PMA_CH1_REG_RX_DCC_IC_TX),                 
    .CP_PMA_CH1_REG_RX_ICTRL_TRX                 (PMA_CH1_REG_RX_ICTRL_TRX),                 
    .CP_PMA_CH1_REG_RX_ICTRL_SIGDET              (PMA_CH1_REG_RX_ICTRL_SIGDET),              
    .CP_PMA_CH1_REG_RX_ICTRL_PREAMP              (PMA_CH1_REG_RX_ICTRL_PREAMP),              
    .CP_PMA_CH1_REG_RX_ICTRL_SLICER              (PMA_CH1_REG_RX_ICTRL_SLICER),              
    .CP_PMA_CH1_REG_RX_ICTRL_PIBUF               (PMA_CH1_REG_RX_ICTRL_PIBUF),               
    .CP_PMA_CH1_REG_RX_ICTRL_PI                  (PMA_CH1_REG_RX_ICTRL_PI),                  
    .CP_PMA_CH1_REG_RX_ICTRL_DCC                 (PMA_CH1_REG_RX_ICTRL_DCC),                 
    .CP_PMA_CH1_REG_RX_ICTRL_PREDRV              (PMA_CH1_REG_RX_ICTRL_PREDRV),              
    .CP_PMA_CH1_REG_TX_RATE                      (PMA_CH1_REG_TX_RATE),                      
    .CP_PMA_CH1_REG_TX_RATE_EN                   (PMA_CH1_REG_TX_RATE_EN),                   
    .CP_PMA_CH1_REG_RX_TX2RX_PLPBK_RST_N         (PMA_CH1_REG_RX_TX2RX_PLPBK_RST_N),         
    .CP_PMA_CH1_REG_RX_TX2RX_PLPBK_RST_N_EN      (PMA_CH1_REG_RX_TX2RX_PLPBK_RST_N_EN),      
    .CP_PMA_CH1_REG_RX_TX2RX_PLPBK_EN            (PMA_CH1_REG_RX_TX2RX_PLPBK_EN),            
    .CP_PMA_CH1_REG_TXCLK_SEL                    (PMA_CH1_REG_TXCLK_SEL),                    
    .CP_PMA_CH1_REG_RX_DATA_POLARITY             (PMA_CH1_REG_RX_DATA_POLARITY),             
    .CP_PMA_CH1_REG_RX_ERR_INSERT                (PMA_CH1_REG_RX_ERR_INSERT),                
    .CP_PMA_CH1_REG_UDP_CHK_EN                   (PMA_CH1_REG_UDP_CHK_EN),                   
    .CP_PMA_CH1_REG_PRBS_SEL                     (PMA_CH1_REG_PRBS_SEL),                     
    .CP_PMA_CH1_REG_PRBS_CHK_EN                  (PMA_CH1_REG_PRBS_CHK_EN),                  
    .CP_PMA_CH1_REG_PRBS_CHK_WIDTH_SEL           (PMA_CH1_REG_PRBS_CHK_WIDTH_SEL),           
    .CP_PMA_CH1_REG_BIST_CHK_PAT_SEL             (PMA_CH1_REG_BIST_CHK_PAT_SEL),             
    .CP_PMA_CH1_REG_LOAD_ERR_CNT                 (PMA_CH1_REG_LOAD_ERR_CNT),                 
    .CP_PMA_CH1_REG_CHK_COUNTER_EN               (PMA_CH1_REG_CHK_COUNTER_EN),               
    .CP_PMA_CH1_REG_CDR_PROP_GAIN                (PMA_CH1_REG_CDR_PROP_GAIN),                
    .CP_PMA_CH1_REG_CDR_PROP_TURBO_GAIN          (PMA_CH1_REG_CDR_PROP_TURBO_GAIN),          
    .CP_PMA_CH1_REG_CDR_INT_GAIN                 (PMA_CH1_REG_CDR_INT_GAIN),                 
    .CP_PMA_CH1_REG_CDR_INT_TURBO_GAIN           (PMA_CH1_REG_CDR_INT_TURBO_GAIN),           
    .CP_PMA_CH1_REG_CDR_INT_SAT_MAX              (PMA_CH1_REG_CDR_INT_SAT_MAX),              
    .CP_PMA_CH1_REG_CDR_INT_SAT_MIN              (PMA_CH1_REG_CDR_INT_SAT_MIN),              
    .CP_PMA_CH1_REG_CDR_INT_RST                  (PMA_CH1_REG_CDR_INT_RST),                  
    .CP_PMA_CH1_REG_CDR_INT_RST_OW               (PMA_CH1_REG_CDR_INT_RST_OW),               
    .CP_PMA_CH1_REG_CDR_PROP_RST                 (PMA_CH1_REG_CDR_PROP_RST),                 
    .CP_PMA_CH1_REG_CDR_PROP_RST_OW              (PMA_CH1_REG_CDR_PROP_RST_OW),              
    .CP_PMA_CH1_REG_CDR_LOCK_RST                 (PMA_CH1_REG_CDR_LOCK_RST),                 
    .CP_PMA_CH1_REG_CDR_LOCK_RST_OW              (PMA_CH1_REG_CDR_LOCK_RST_OW),              
    .CP_PMA_CH1_REG_CDR_RX_PI_FORCE_SEL          (PMA_CH1_REG_CDR_RX_PI_FORCE_SEL),          
    .CP_PMA_CH1_REG_CDR_RX_PI_FORCE_D            (PMA_CH1_REG_CDR_RX_PI_FORCE_D),            
    .CP_PMA_CH1_REG_CDR_LOCK_TIMER               (PMA_CH1_REG_CDR_LOCK_TIMER),               
    .CP_PMA_CH1_REG_CDR_TURBO_MODE_TIMER         (PMA_CH1_REG_CDR_TURBO_MODE_TIMER),         
    .CP_PMA_CH1_REG_CDR_LOCK_VAL                 (PMA_CH1_REG_CDR_LOCK_VAL),                 
    .CP_PMA_CH1_REG_CDR_LOCK_OW                  (PMA_CH1_REG_CDR_LOCK_OW),                  
    .CP_PMA_CH1_REG_CDR_INT_SAT_DET_EN           (PMA_CH1_REG_CDR_INT_SAT_DET_EN),           
    .CP_PMA_CH1_REG_CDR_SAT_DET_STATUS_EN        (PMA_CH1_REG_CDR_SAT_DET_STATUS_EN),        
    .CP_PMA_CH1_REG_CDR_SAT_DET_STATUS_RESET_EN  (PMA_CH1_REG_CDR_SAT_DET_STATUS_RESET_EN),   
    .CP_PMA_CH1_REG_CDR_PI_CTRL_RST              (PMA_CH1_REG_CDR_PI_CTRL_RST),              
    .CP_PMA_CH1_REG_CDR_PI_CTRL_RST_OW           (PMA_CH1_REG_CDR_PI_CTRL_RST_OW),           
    .CP_PMA_CH1_REG_CDR_SAT_DET_RST              (PMA_CH1_REG_CDR_SAT_DET_RST),              
    .CP_PMA_CH1_REG_CDR_SAT_DET_RST_OW           (PMA_CH1_REG_CDR_SAT_DET_RST_OW),           
    .CP_PMA_CH1_REG_CDR_SAT_DET_STICKY_RST       (PMA_CH1_REG_CDR_SAT_DET_STICKY_RST),       
    .CP_PMA_CH1_REG_CDR_SAT_DET_STICKY_RST_OW    (PMA_CH1_REG_CDR_SAT_DET_STICKY_RST_OW),    
    .CP_PMA_CH1_REG_CDR_SIGDET_STATUS_DIS        (PMA_CH1_REG_CDR_SIGDET_STATUS_DIS),        
    .CP_PMA_CH1_REG_CDR_SAT_DET_TIMER            (PMA_CH1_REG_CDR_SAT_DET_TIMER),            
    .CP_PMA_CH1_REG_CDR_SAT_DET_STATUS_VAL       (PMA_CH1_REG_CDR_SAT_DET_STATUS_VAL),       
    .CP_PMA_CH1_REG_CDR_SAT_DET_STATUS_OW        (PMA_CH1_REG_CDR_SAT_DET_STATUS_OW),        
    .CP_PMA_CH1_REG_CDR_TURBO_MODE_EN            (PMA_CH1_REG_CDR_TURBO_MODE_EN),            
    .CP_PMA_CH1_REG_CDR_STATUS_RADDR_INIT        (PMA_CH1_REG_CDR_STATUS_RADDR_INIT),        
    .CP_PMA_CH1_REG_CDR_STATUS_FIFO_EN           (PMA_CH1_REG_CDR_STATUS_FIFO_EN),           
    .CP_PMA_CH1_REG_PMA_TEST_SEL                 (PMA_CH1_REG_PMA_TEST_SEL),                 
    .CP_PMA_CH1_REG_OOB_COMWAKE_GAP_MIN          (PMA_CH1_REG_OOB_COMWAKE_GAP_MIN),          
    .CP_PMA_CH1_REG_OOB_COMWAKE_GAP_MAX          (PMA_CH1_REG_OOB_COMWAKE_GAP_MAX),          
    .CP_PMA_CH1_REG_OOB_COMINIT_GAP_MIN          (PMA_CH1_REG_OOB_COMINIT_GAP_MIN),          
    .CP_PMA_CH1_REG_OOB_COMINIT_GAP_MAX          (PMA_CH1_REG_OOB_COMINIT_GAP_MAX),          
    .CP_PMA_CH1_REG_RX_PIBUF_IC_TX               (PMA_CH1_REG_RX_PIBUF_IC_TX),               
    .CP_PMA_CH1_REG_COMWAKE_STATUS_CLEAR         (PMA_CH1_REG_COMWAKE_STATUS_CLEAR),         
    .CP_PMA_CH1_REG_COMINIT_STATUS_CLEAR         (PMA_CH1_REG_COMINIT_STATUS_CLEAR),         
    .CP_PMA_CH1_REG_RX_SYNC_RST_N_EN             (PMA_CH1_REG_RX_SYNC_RST_N_EN),             
    .CP_PMA_CH1_REG_RX_SYNC_RST_N                (PMA_CH1_REG_RX_SYNC_RST_N),                
    .CP_PMA_CH1_REG_RX_SATA_COMINIT_OW           (PMA_CH1_REG_RX_SATA_COMINIT_OW),           
    .CP_PMA_CH1_REG_RX_SATA_COMINIT              (PMA_CH1_REG_RX_SATA_COMINIT),              
    .CP_PMA_CH1_REG_RX_SATA_COMWAKE_OW           (PMA_CH1_REG_RX_SATA_COMWAKE_OW),           
    .CP_PMA_CH1_REG_RX_SATA_COMWAKE              (PMA_CH1_REG_RX_SATA_COMWAKE),              
    .CP_PMA_CH1_REG_RX_DCC_DISABLE               (PMA_CH1_REG_RX_DCC_DISABLE),               
    .CP_PMA_CH1_REG_TX_DCC_DISABLE               (PMA_CH1_REG_TX_DCC_DISABLE),               
    .CP_PMA_CH1_REG_RX_SLIP_SEL_EN               (PMA_CH1_REG_RX_SLIP_SEL_EN),               
    .CP_PMA_CH1_REG_RX_SLIP_SEL                  (PMA_CH1_REG_RX_SLIP_SEL),                  
    .CP_PMA_CH1_REG_RX_SLIP_EN                   (PMA_CH1_REG_RX_SLIP_EN),                   
    .CP_PMA_CH1_REG_RX_SIGDET_STATUS_SEL         (PMA_CH1_REG_RX_SIGDET_STATUS_SEL),         
    .CP_PMA_CH1_REG_RX_SIGDET_FSM_RST_N          (PMA_CH1_REG_RX_SIGDET_FSM_RST_N),          
    .CP_PMA_CH1_REG_RX_SIGDET_STATUS_OW          (PMA_CH1_REG_RX_SIGDET_STATUS_OW),          
    .CP_PMA_CH1_REG_RX_SIGDET_STATUS             (PMA_CH1_REG_RX_SIGDET_STATUS),             
    .CP_PMA_CH1_REG_RX_SIGDET_VTH                (PMA_CH1_REG_RX_SIGDET_VTH),                
    .CP_PMA_CH1_REG_RX_SIGDET_GRM                (PMA_CH1_REG_RX_SIGDET_GRM),                
    .CP_PMA_CH1_REG_RX_SIGDET_PULSE_EXT          (PMA_CH1_REG_RX_SIGDET_PULSE_EXT),          
    .CP_PMA_CH1_REG_RX_SIGDET_CH2_SEL            (PMA_CH1_REG_RX_SIGDET_CH2_SEL),            
    .CP_PMA_CH1_REG_RX_SIGDET_CH2_CHK_WINDOW     (PMA_CH1_REG_RX_SIGDET_CH2_CHK_WINDOW),     
    .CP_PMA_CH1_REG_RX_SIGDET_CHK_WINDOW_EN      (PMA_CH1_REG_RX_SIGDET_CHK_WINDOW_EN),      
    .CP_PMA_CH1_REG_RX_SIGDET_NOSIG_COUNT_SETTING(PMA_CH1_REG_RX_SIGDET_NOSIG_COUNT_SETTING),
    .CP_PMA_CH1_REG_RX_SIGDET_OOB_DET_COUNT_VAL  (PMA_CH1_REG_RX_SIGDET_OOB_DET_COUNT_VAL),  
    .CP_PMA_CH1_REG_SLIP_FIFO_INV_EN             (PMA_CH1_REG_SLIP_FIFO_INV_EN),             
    .CP_PMA_CH1_REG_SLIP_FIFO_INV                (PMA_CH1_REG_SLIP_FIFO_INV),                
    .CP_PMA_CH1_REG_RX_SIGDET_4OOB_DET_SEL       (PMA_CH1_REG_RX_SIGDET_4OOB_DET_SEL),       
    .CP_PMA_CH1_REG_RX_SIGDET_IC_I               (PMA_CH1_REG_RX_SIGDET_IC_I),               
    .CP_PMA_CH1_REG_RX_OOB_DETECTOR_RESET_N_OW   (PMA_CH1_REG_RX_OOB_DETECTOR_RESET_N_OW),   
    .CP_PMA_CH1_REG_RX_OOB_DETECTOR_RESET_N      (PMA_CH1_REG_RX_OOB_DETECTOR_RESET_N),      
    .CP_PMA_CH1_REG_RX_OOB_DETECTOR_PD_OW        (PMA_CH1_REG_RX_OOB_DETECTOR_PD_OW),        
    .CP_PMA_CH1_REG_RX_OOB_DETECTOR_PD           (PMA_CH1_REG_RX_OOB_DETECTOR_PD),           
    .CP_PMA_CH1_REG_RX_TERM_CM_CTRL              (PMA_CH1_REG_RX_TERM_CM_CTRL),              
    .CP_PMA_CH1_REG_TX_PD                        (PMA_CH1_REG_TX_PD),                        
    .CP_PMA_CH1_REG_TX_PD_OW                     (PMA_CH1_REG_TX_PD_OW),                     
    .CP_PMA_CH1_REG_TX_CLKPATH_PD                (PMA_CH1_REG_TX_CLKPATH_PD),                
    .CP_PMA_CH1_REG_TX_CLKPATH_PD_OW             (PMA_CH1_REG_TX_CLKPATH_PD_OW),             
    .CP_PMA_CH1_REG_TX_BEACON_TIMER_SEL          (PMA_CH1_REG_TX_BEACON_TIMER_SEL),          
    .CP_PMA_CH1_REG_TX_RXDET_REQ_OW              (PMA_CH1_REG_TX_RXDET_REQ_OW),              
    .CP_PMA_CH1_REG_TX_RXDET_REQ                 (PMA_CH1_REG_TX_RXDET_REQ),                 
    .CP_PMA_CH1_REG_TX_BEACON_EN_OW              (PMA_CH1_REG_TX_BEACON_EN_OW),              
    .CP_PMA_CH1_REG_TX_BEACON_EN                 (PMA_CH1_REG_TX_BEACON_EN),                 
    .CP_PMA_CH1_REG_TX_EI_EN_OW                  (PMA_CH1_REG_TX_EI_EN_OW),                  
    .CP_PMA_CH1_REG_TX_EI_EN                     (PMA_CH1_REG_TX_EI_EN),                     
    .CP_PMA_CH1_REG_TX_RES_CAL_EN                (PMA_CH1_REG_TX_RES_CAL_EN),                
    .CP_PMA_CH1_REG_TX_RES_CAL                   (PMA_CH1_REG_TX_RES_CAL),                   
    .CP_PMA_CH1_REG_TX_BIAS_CAL_EN               (PMA_CH1_REG_TX_BIAS_CAL_EN),               
    .CP_PMA_CH1_REG_TX_BIAS_CTRL                 (PMA_CH1_REG_TX_BIAS_CTRL),                 
    .CP_PMA_CH1_REG_TX_RXDET_TIMER_SEL           (PMA_CH1_REG_TX_RXDET_TIMER_SEL),           
    .CP_PMA_CH1_REG_TX_SYNC_OW                   (PMA_CH1_REG_TX_SYNC_OW),                   
    .CP_PMA_CH1_REG_TX_SYNC                      (PMA_CH1_REG_TX_SYNC),                      
    .CP_PMA_CH1_REG_TX_PD_POST                   (PMA_CH1_REG_TX_PD_POST),                   
    .CP_PMA_CH1_REG_TX_PD_POST_OW                (PMA_CH1_REG_TX_PD_POST_OW),               
    .CP_PMA_CH1_REG_TX_RESET_N_OW                (PMA_CH1_REG_TX_RESET_N_OW),                
    .CP_PMA_CH1_REG_TX_RESET_N                   (PMA_CH1_REG_TX_RESET_N),                   
    .CP_PMA_CH1_REG_TX_DCC_RESET_N_OW            (PMA_CH1_REG_TX_DCC_RESET_N_OW),            
    .CP_PMA_CH1_REG_TX_DCC_RESET_N               (PMA_CH1_REG_TX_DCC_RESET_N),               
    .CP_PMA_CH1_REG_TX_BUSWIDTH_OW               (PMA_CH1_REG_TX_BUSWIDTH_OW),               
    .CP_PMA_CH1_REG_TX_BUSWIDTH                  (PMA_CH1_REG_TX_BUSWIDTH),                  
    .CP_PMA_CH1_REG_PLL_READY_OW                 (PMA_CH1_REG_PLL_READY_OW),                 
    .CP_PMA_CH1_REG_PLL_READY                    (PMA_CH1_REG_PLL_READY),                    
    .CP_PMA_CH1_REG_TX_PCLK_SW_OW                (PMA_CH1_REG_TX_PCLK_SW_OW),                
    .CP_PMA_CH1_REG_TX_PCLK_SW                   (PMA_CH1_REG_TX_PCLK_SW),                   
    .CP_PMA_CH1_REG_EI_PCLK_DELAY_SEL            (PMA_CH1_REG_EI_PCLK_DELAY_SEL),            
    .CP_PMA_CH1_REG_TX_DRV01_DAC0                (PMA_CH1_REG_TX_DRV01_DAC0),                
    .CP_PMA_CH1_REG_TX_DRV01_DAC1                (PMA_CH1_REG_TX_DRV01_DAC1),                
    .CP_PMA_CH1_REG_TX_DRV01_DAC2                (PMA_CH1_REG_TX_DRV01_DAC2),                
    .CP_PMA_CH1_REG_TX_DRV00_DAC0                (PMA_CH1_REG_TX_DRV00_DAC0),                
    .CP_PMA_CH1_REG_TX_DRV00_DAC1                (PMA_CH1_REG_TX_DRV00_DAC1),                
    .CP_PMA_CH1_REG_TX_DRV00_DAC2                (PMA_CH1_REG_TX_DRV00_DAC2),                
    .CP_PMA_CH1_REG_TX_AMP0                      (PMA_CH1_REG_TX_AMP0),                      
    .CP_PMA_CH1_REG_TX_AMP1                      (PMA_CH1_REG_TX_AMP1),                      
    .CP_PMA_CH1_REG_TX_AMP2                      (PMA_CH1_REG_TX_AMP2),                      
    .CP_PMA_CH1_REG_TX_AMP3                      (PMA_CH1_REG_TX_AMP3),                      
    .CP_PMA_CH1_REG_TX_AMP4                      (PMA_CH1_REG_TX_AMP4),                      
    .CP_PMA_CH1_REG_TX_MARGIN                    (PMA_CH1_REG_TX_MARGIN),                    
    .CP_PMA_CH1_REG_TX_MARGIN_OW                 (PMA_CH1_REG_TX_MARGIN_OW),                 
    .CP_PMA_CH1_REG_TX_DEEMP                     (PMA_CH1_REG_TX_DEEMP),                     
    .CP_PMA_CH1_REG_TX_DEEMP_OW                  (PMA_CH1_REG_TX_DEEMP_OW),                  
    .CP_PMA_CH1_REG_TX_SWING                     (PMA_CH1_REG_TX_SWING),                     
    .CP_PMA_CH1_REG_TX_SWING_OW                  (PMA_CH1_REG_TX_SWING_OW),                  
    .CP_PMA_CH1_REG_TX_RXDET_THRESHOLD           (PMA_CH1_REG_TX_RXDET_THRESHOLD),           
    .CP_PMA_CH1_REG_TX_BEACON_OSC_CTRL           (PMA_CH1_REG_TX_BEACON_OSC_CTRL),           
    .CP_PMA_CH1_REG_TX_PREDRV_DAC                (PMA_CH1_REG_TX_PREDRV_DAC),                
    .CP_PMA_CH1_REG_TX_PREDRV_CM_CTRL            (PMA_CH1_REG_TX_PREDRV_CM_CTRL),            
    .CP_PMA_CH1_REG_TX_TX2RX_SLPBACK_EN          (PMA_CH1_REG_TX_TX2RX_SLPBACK_EN),          
    .CP_PMA_CH1_REG_TX_PCLK_EDGE_SEL             (PMA_CH1_REG_TX_PCLK_EDGE_SEL),             
    .CP_PMA_CH1_REG_TX_RXDET_STATUS_OW           (PMA_CH1_REG_TX_RXDET_STATUS_OW),           
    .CP_PMA_CH1_REG_TX_RXDET_STATUS              (PMA_CH1_REG_TX_RXDET_STATUS),              
    .CP_PMA_CH1_REG_TX_PRBS_GEN_EN               (PMA_CH1_REG_TX_PRBS_GEN_EN),               
    .CP_PMA_CH1_REG_TX_PRBS_GEN_WIDTH_SEL        (PMA_CH1_REG_TX_PRBS_GEN_WIDTH_SEL),        
    .CP_PMA_CH1_REG_TX_PRBS_SEL                  (PMA_CH1_REG_TX_PRBS_SEL),                  
    .CP_PMA_CH1_REG_TX_UDP_DATA                  (PMA_CH1_REG_TX_UDP_DATA),                  
    .CP_PMA_CH1_REG_TX_FIFO_RST_N                (PMA_CH1_REG_TX_FIFO_RST_N),                
    .CP_PMA_CH1_REG_TX_FIFO_WP_CTRL              (PMA_CH1_REG_TX_FIFO_WP_CTRL),              
    .CP_PMA_CH1_REG_TX_FIFO_EN                   (PMA_CH1_REG_TX_FIFO_EN),                   
    .CP_PMA_CH1_REG_TX_DATA_MUX_SEL              (PMA_CH1_REG_TX_DATA_MUX_SEL),              
    .CP_PMA_CH1_REG_TX_ERR_INSERT                (PMA_CH1_REG_TX_ERR_INSERT),                
    .CP_PMA_CH1_REG_TX_SATA_EN                   (PMA_CH1_REG_TX_SATA_EN),                   
    .CP_PMA_CH1_REG_RATE_CHANGE_TXPCLK_ON_OW     (PMA_CH1_REG_RATE_CHANGE_TXPCLK_ON_OW),     
    .CP_PMA_CH1_REG_RATE_CHANGE_TXPCLK_ON        (PMA_CH1_REG_RATE_CHANGE_TXPCLK_ON),        
    .CP_PMA_CH1_REG_TX_PULLUP_DAC0               (PMA_CH1_REG_TX_PULLUP_DAC0),               
    .CP_PMA_CH1_REG_TX_PULLUP_DAC1               (PMA_CH1_REG_TX_PULLUP_DAC1),               
    .CP_PMA_CH1_REG_TX_PULLUP_DAC2               (PMA_CH1_REG_TX_PULLUP_DAC2),               
    .CP_PMA_CH1_REG_TX_PULLUP_DAC3               (PMA_CH1_REG_TX_PULLUP_DAC3),               
    .CP_PMA_CH1_REG_TX_OOB_DELAY_SEL             (PMA_CH1_REG_TX_OOB_DELAY_SEL),             
    .CP_PMA_CH1_REG_TX_POLARITY                  (PMA_CH1_REG_TX_POLARITY),                  
    .CP_PMA_CH1_REG_TX_SLPBK_AMP                 (PMA_CH1_REG_TX_SLPBK_AMP),                 
    .CP_PMA_CH1_REG_TX_LS_MODE_EN                (PMA_CH1_REG_TX_LS_MODE_EN),                
    .CP_PMA_CH1_REG_TX_JTAG_MODE_EN_OW           (PMA_CH1_REG_TX_JTAG_MODE_EN_OW),           
    .CP_PMA_CH1_REG_TX_JTAG_MODE_EN              (PMA_CH1_REG_TX_JTAG_MODE_EN),              
    .CP_PMA_CH1_REG_RX_JTAG_MODE_EN_OW           (PMA_CH1_REG_RX_JTAG_MODE_EN_OW),           
    .CP_PMA_CH1_REG_RX_JTAG_MODE_EN              (PMA_CH1_REG_RX_JTAG_MODE_EN),              
    .CP_PMA_CH1_REG_RX_JTAG_OE                   (PMA_CH1_REG_RX_JTAG_OE),                   
    .CP_PMA_CH1_REG_RX_ACJTAG_VHYSTSE            (PMA_CH1_REG_RX_ACJTAG_VHYSTSE),            
    .CP_PMA_CH1_REG_TX_FBCLK_FAR_EN              (PMA_CH1_REG_TX_FBCLK_FAR_EN),              
    .CP_PMA_CH1_REG_RX_TERM_MODE_CTRL            (PMA_CH1_REG_RX_TERM_MODE_CTRL),            
    .CP_PMA_CH1_REG_PLPBK_TXPCLK_EN              (PMA_CH1_REG_PLPBK_TXPCLK_EN),              
    .CP_PMA_CH1_CFG_LANE_POWERUP                 (PMA_CH1_CFG_LANE_POWERUP),                 
    .CP_PMA_CH1_CFG_PMA_POR_N                    (PMA_CH1_CFG_PMA_POR_N),                    
    .CP_PMA_CH1_CFG_RX_LANE_POWERUP              (PMA_CH1_CFG_RX_LANE_POWERUP),              
    .CP_PMA_CH1_CFG_RX_PMA_RSTN                  (PMA_CH1_CFG_RX_PMA_RSTN),                  
    .CP_PMA_CH1_CFG_TX_LANE_POWERUP              (PMA_CH1_CFG_TX_LANE_POWERUP),              
    .CP_PMA_CH1_CFG_TX_PMA_RSTN                  (PMA_CH1_CFG_TX_PMA_RSTN),                  
    .CP_PMA_CH1_REG_RESERVED_48_45               (PMA_CH1_REG_RESERVED_48_45),               
    .CP_PMA_CH1_REG_RESERVED_69                  (PMA_CH1_REG_RESERVED_69),                  
    .CP_PMA_CH1_REG_RESERVED_77_76               (PMA_CH1_REG_RESERVED_77_76),               
    .CP_PMA_CH1_REG_RESERVED_171_164             (PMA_CH1_REG_RESERVED_171_164),             
    .CP_PMA_CH1_REG_RESERVED_175_172             (PMA_CH1_REG_RESERVED_175_172),             
    .CP_PMA_CH1_REG_RESERVED_190                 (PMA_CH1_REG_RESERVED_190),                 
    .CP_PMA_CH1_REG_RESERVED_233_232             (PMA_CH1_REG_RESERVED_233_232),             
    .CP_PMA_CH1_REG_RESERVED_235_234             (PMA_CH1_REG_RESERVED_235_234),             
    .CP_PMA_CH1_REG_RESERVED_241_240             (PMA_CH1_REG_RESERVED_241_240),             
    .CP_PMA_CH1_REG_RESERVED_285_283             (PMA_CH1_REG_RESERVED_285_283),             
    .CP_PMA_CH1_REG_RESERVED_286                 (PMA_CH1_REG_RESERVED_286),                 
    .CP_PMA_CH1_REG_RESERVED_295                 (PMA_CH1_REG_RESERVED_295),                 
    .CP_PMA_CH1_REG_RESERVED_298                 (PMA_CH1_REG_RESERVED_298),                 
    .CP_PMA_CH1_REG_RESERVED_332_325             (PMA_CH1_REG_RESERVED_332_325),             
    .CP_PMA_CH1_REG_RESERVED_340_333             (PMA_CH1_REG_RESERVED_340_333),             
    .CP_PMA_CH1_REG_RESERVED_348_341             (PMA_CH1_REG_RESERVED_348_341),             
    .CP_PMA_CH1_REG_RESERVED_354_349             (PMA_CH1_REG_RESERVED_354_349),             
    .CP_PMA_CH1_REG_RESERVED_373                 (PMA_CH1_REG_RESERVED_373),                 
    .CP_PMA_CH1_REG_RESERVED_376                 (PMA_CH1_REG_RESERVED_376),                 
    .CP_PMA_CH1_REG_RESERVED_452                 (PMA_CH1_REG_RESERVED_452),                 
    .CP_PMA_CH1_REG_RESERVED_502_499             (PMA_CH1_REG_RESERVED_502_499),             
    .CP_PMA_CH1_REG_RESERVED_506_505             (PMA_CH1_REG_RESERVED_506_505),             
    .CP_PMA_CH1_REG_RESERVED_550_549             (PMA_CH1_REG_RESERVED_550_549),             
    .CP_PMA_CH1_REG_RESERVED_556_552             (PMA_CH1_REG_RESERVED_556_552),             
    .CP_PMA_CH2_REG_RX_PD                        (PMA_CH2_REG_RX_PD),                        
    .CP_PMA_CH2_REG_RX_PD_EN                     (PMA_CH2_REG_RX_PD_EN),                     
    .CP_PMA_CH2_REG_RX_CLKPATH_PD                (PMA_CH2_REG_RX_CLKPATH_PD),                
    .CP_PMA_CH2_REG_RX_CLKPATH_PD_EN             (PMA_CH2_REG_RX_CLKPATH_PD_EN),             
    .CP_PMA_CH2_REG_RX_DATAPATH_PD               (PMA_CH2_REG_RX_DATAPATH_PD),               
    .CP_PMA_CH2_REG_RX_DATAPATH_PD_EN            (PMA_CH2_REG_RX_DATAPATH_PD_EN),            
    .CP_PMA_CH2_REG_RX_SIGDET_PD                 (PMA_CH2_REG_RX_SIGDET_PD),                 
    .CP_PMA_CH2_REG_RX_SIGDET_PD_EN              (PMA_CH2_REG_RX_SIGDET_PD_EN),              
    .CP_PMA_CH2_REG_RX_DCC_RST_N                 (PMA_CH2_REG_RX_DCC_RST_N),                 
    .CP_PMA_CH2_REG_RX_DCC_RST_N_EN              (PMA_CH2_REG_RX_DCC_RST_N_EN),              
    .CP_PMA_CH2_REG_RX_CDR_RST_N                 (PMA_CH2_REG_RX_CDR_RST_N),                 
    .CP_PMA_CH2_REG_RX_CDR_RST_N_EN              (PMA_CH2_REG_RX_CDR_RST_N_EN),              
    .CP_PMA_CH2_REG_RX_SIGDET_RST_N              (PMA_CH2_REG_RX_SIGDET_RST_N),              
    .CP_PMA_CH2_REG_RX_SIGDET_RST_N_EN           (PMA_CH2_REG_RX_SIGDET_RST_N_EN),           
    .CP_PMA_CH2_REG_RXPCLK_SLIP                  (PMA_CH2_REG_RXPCLK_SLIP),                  
    .CP_PMA_CH2_REG_RXPCLK_SLIP_OW               (PMA_CH2_REG_RXPCLK_SLIP_OW),               
    .CP_PMA_CH2_REG_RX_PCLKSWITCH_RST_N          (PMA_CH2_REG_RX_PCLKSWITCH_RST_N),          
    .CP_PMA_CH2_REG_RX_PCLKSWITCH_RST_N_EN       (PMA_CH2_REG_RX_PCLKSWITCH_RST_N_EN),       
    .CP_PMA_CH2_REG_RX_PCLKSWITCH                (PMA_CH2_REG_RX_PCLKSWITCH),                
    .CP_PMA_CH2_REG_RX_PCLKSWITCH_EN             (PMA_CH2_REG_RX_PCLKSWITCH_EN),             
    .CP_PMA_CH2_REG_RX_HIGHZ                     (PMA_CH2_REG_RX_HIGHZ),                     
    .CP_PMA_CH2_REG_RX_HIGHZ_EN                  (PMA_CH2_REG_RX_HIGHZ_EN),                  
    .CP_PMA_CH2_REG_RX_EQ_C_SET                  (PMA_CH2_REG_RX_EQ_C_SET),                  
    .CP_PMA_CH2_REG_RX_EQ_R_SET                  (PMA_CH2_REG_RX_EQ_R_SET),                  
    .CP_PMA_CH2_REG_RX_BUSWIDTH                  (PMA_CH2_REG_RX_BUSWIDTH),                  
    .CP_PMA_CH2_REG_RX_BUSWIDTH_EN               (PMA_CH2_REG_RX_BUSWIDTH_EN),              
    .CP_PMA_CH2_REG_RX_RATE                      (PMA_CH2_REG_RX_RATE),                      
    .CP_PMA_CH2_REG_RX_RATE_EN                   (PMA_CH2_REG_RX_RATE_EN),                   
    .CP_PMA_CH2_REG_RX_RES_TRIM                  (PMA_CH2_REG_RX_RES_TRIM),                  
    .CP_PMA_CH2_REG_RX_RES_TRIM_EN               (PMA_CH2_REG_RX_RES_TRIM_EN),               
    .CP_PMA_CH2_REG_RX_EQ_OFF                    (PMA_CH2_REG_RX_EQ_OFF),                    
    .CP_PMA_CH2_REG_RX_PREAMP_IC                 (PMA_CH2_REG_RX_PREAMP_IC),                 
    .CP_PMA_CH2_REG_RX_PCLK_EDGE_SEL             (PMA_CH2_REG_RX_PCLK_EDGE_SEL),             
    .CP_PMA_CH2_REG_RX_PIBUF_IC                  (PMA_CH2_REG_RX_PIBUF_IC),                  
    .CP_PMA_CH2_REG_RX_DCC_IC_RX                 (PMA_CH2_REG_RX_DCC_IC_RX),                 
    .CP_PMA_CH2_REG_RX_DCC_IC_TX                 (PMA_CH2_REG_RX_DCC_IC_TX),                 
    .CP_PMA_CH2_REG_RX_ICTRL_TRX                 (PMA_CH2_REG_RX_ICTRL_TRX),                 
    .CP_PMA_CH2_REG_RX_ICTRL_SIGDET              (PMA_CH2_REG_RX_ICTRL_SIGDET),              
    .CP_PMA_CH2_REG_RX_ICTRL_PREAMP              (PMA_CH2_REG_RX_ICTRL_PREAMP),              
    .CP_PMA_CH2_REG_RX_ICTRL_SLICER              (PMA_CH2_REG_RX_ICTRL_SLICER),              
    .CP_PMA_CH2_REG_RX_ICTRL_PIBUF               (PMA_CH2_REG_RX_ICTRL_PIBUF),               
    .CP_PMA_CH2_REG_RX_ICTRL_PI                  (PMA_CH2_REG_RX_ICTRL_PI),                  
    .CP_PMA_CH2_REG_RX_ICTRL_DCC                 (PMA_CH2_REG_RX_ICTRL_DCC),                 
    .CP_PMA_CH2_REG_RX_ICTRL_PREDRV              (PMA_CH2_REG_RX_ICTRL_PREDRV),              
    .CP_PMA_CH2_REG_TX_RATE                      (PMA_CH2_REG_TX_RATE),                      
    .CP_PMA_CH2_REG_TX_RATE_EN                   (PMA_CH2_REG_TX_RATE_EN),                   
    .CP_PMA_CH2_REG_RX_TX2RX_PLPBK_RST_N         (PMA_CH2_REG_RX_TX2RX_PLPBK_RST_N),         
    .CP_PMA_CH2_REG_RX_TX2RX_PLPBK_RST_N_EN      (PMA_CH2_REG_RX_TX2RX_PLPBK_RST_N_EN),      
    .CP_PMA_CH2_REG_RX_TX2RX_PLPBK_EN            (PMA_CH2_REG_RX_TX2RX_PLPBK_EN),            
    .CP_PMA_CH2_REG_TXCLK_SEL                    (PMA_CH2_REG_TXCLK_SEL),                    
    .CP_PMA_CH2_REG_RX_DATA_POLARITY             (PMA_CH2_REG_RX_DATA_POLARITY),             
    .CP_PMA_CH2_REG_RX_ERR_INSERT                (PMA_CH2_REG_RX_ERR_INSERT),                
    .CP_PMA_CH2_REG_UDP_CHK_EN                   (PMA_CH2_REG_UDP_CHK_EN),                   
    .CP_PMA_CH2_REG_PRBS_SEL                     (PMA_CH2_REG_PRBS_SEL),                     
    .CP_PMA_CH2_REG_PRBS_CHK_EN                  (PMA_CH2_REG_PRBS_CHK_EN),                  
    .CP_PMA_CH2_REG_PRBS_CHK_WIDTH_SEL           (PMA_CH2_REG_PRBS_CHK_WIDTH_SEL),           
    .CP_PMA_CH2_REG_BIST_CHK_PAT_SEL             (PMA_CH2_REG_BIST_CHK_PAT_SEL),             
    .CP_PMA_CH2_REG_LOAD_ERR_CNT                 (PMA_CH2_REG_LOAD_ERR_CNT),                 
    .CP_PMA_CH2_REG_CHK_COUNTER_EN               (PMA_CH2_REG_CHK_COUNTER_EN),               
    .CP_PMA_CH2_REG_CDR_PROP_GAIN                (PMA_CH2_REG_CDR_PROP_GAIN),                
    .CP_PMA_CH2_REG_CDR_PROP_TURBO_GAIN          (PMA_CH2_REG_CDR_PROP_TURBO_GAIN),          
    .CP_PMA_CH2_REG_CDR_INT_GAIN                 (PMA_CH2_REG_CDR_INT_GAIN),                 
    .CP_PMA_CH2_REG_CDR_INT_TURBO_GAIN           (PMA_CH2_REG_CDR_INT_TURBO_GAIN),           
    .CP_PMA_CH2_REG_CDR_INT_SAT_MAX              (PMA_CH2_REG_CDR_INT_SAT_MAX),              
    .CP_PMA_CH2_REG_CDR_INT_SAT_MIN              (PMA_CH2_REG_CDR_INT_SAT_MIN),              
    .CP_PMA_CH2_REG_CDR_INT_RST                  (PMA_CH2_REG_CDR_INT_RST),                  
    .CP_PMA_CH2_REG_CDR_INT_RST_OW               (PMA_CH2_REG_CDR_INT_RST_OW),               
    .CP_PMA_CH2_REG_CDR_PROP_RST                 (PMA_CH2_REG_CDR_PROP_RST),                 
    .CP_PMA_CH2_REG_CDR_PROP_RST_OW              (PMA_CH2_REG_CDR_PROP_RST_OW),              
    .CP_PMA_CH2_REG_CDR_LOCK_RST                 (PMA_CH2_REG_CDR_LOCK_RST),                 
    .CP_PMA_CH2_REG_CDR_LOCK_RST_OW              (PMA_CH2_REG_CDR_LOCK_RST_OW),              
    .CP_PMA_CH2_REG_CDR_RX_PI_FORCE_SEL          (PMA_CH2_REG_CDR_RX_PI_FORCE_SEL),          
    .CP_PMA_CH2_REG_CDR_RX_PI_FORCE_D            (PMA_CH2_REG_CDR_RX_PI_FORCE_D),            
    .CP_PMA_CH2_REG_CDR_LOCK_TIMER               (PMA_CH2_REG_CDR_LOCK_TIMER),               
    .CP_PMA_CH2_REG_CDR_TURBO_MODE_TIMER         (PMA_CH2_REG_CDR_TURBO_MODE_TIMER),         
    .CP_PMA_CH2_REG_CDR_LOCK_VAL                 (PMA_CH2_REG_CDR_LOCK_VAL),                 
    .CP_PMA_CH2_REG_CDR_LOCK_OW                  (PMA_CH2_REG_CDR_LOCK_OW),                  
    .CP_PMA_CH2_REG_CDR_INT_SAT_DET_EN           (PMA_CH2_REG_CDR_INT_SAT_DET_EN),           
    .CP_PMA_CH2_REG_CDR_SAT_DET_STATUS_EN        (PMA_CH2_REG_CDR_SAT_DET_STATUS_EN),        
    .CP_PMA_CH2_REG_CDR_SAT_DET_STATUS_RESET_EN  (PMA_CH2_REG_CDR_SAT_DET_STATUS_RESET_EN),  
    .CP_PMA_CH2_REG_CDR_PI_CTRL_RST              (PMA_CH2_REG_CDR_PI_CTRL_RST),              
    .CP_PMA_CH2_REG_CDR_PI_CTRL_RST_OW           (PMA_CH2_REG_CDR_PI_CTRL_RST_OW),           
    .CP_PMA_CH2_REG_CDR_SAT_DET_RST              (PMA_CH2_REG_CDR_SAT_DET_RST),              
    .CP_PMA_CH2_REG_CDR_SAT_DET_RST_OW           (PMA_CH2_REG_CDR_SAT_DET_RST_OW),           
    .CP_PMA_CH2_REG_CDR_SAT_DET_STICKY_RST       (PMA_CH2_REG_CDR_SAT_DET_STICKY_RST),       
    .CP_PMA_CH2_REG_CDR_SAT_DET_STICKY_RST_OW    (PMA_CH2_REG_CDR_SAT_DET_STICKY_RST_OW),    
    .CP_PMA_CH2_REG_CDR_SIGDET_STATUS_DIS        (PMA_CH2_REG_CDR_SIGDET_STATUS_DIS),        
    .CP_PMA_CH2_REG_CDR_SAT_DET_TIMER            (PMA_CH2_REG_CDR_SAT_DET_TIMER),            
    .CP_PMA_CH2_REG_CDR_SAT_DET_STATUS_VAL       (PMA_CH2_REG_CDR_SAT_DET_STATUS_VAL),       
    .CP_PMA_CH2_REG_CDR_SAT_DET_STATUS_OW        (PMA_CH2_REG_CDR_SAT_DET_STATUS_OW),        
    .CP_PMA_CH2_REG_CDR_TURBO_MODE_EN            (PMA_CH2_REG_CDR_TURBO_MODE_EN),            
    .CP_PMA_CH2_REG_CDR_STATUS_RADDR_INIT        (PMA_CH2_REG_CDR_STATUS_RADDR_INIT),        
    .CP_PMA_CH2_REG_CDR_STATUS_FIFO_EN           (PMA_CH2_REG_CDR_STATUS_FIFO_EN),           
    .CP_PMA_CH2_REG_PMA_TEST_SEL                 (PMA_CH2_REG_PMA_TEST_SEL),                 
    .CP_PMA_CH2_REG_OOB_COMWAKE_GAP_MIN          (PMA_CH2_REG_OOB_COMWAKE_GAP_MIN),          
    .CP_PMA_CH2_REG_OOB_COMWAKE_GAP_MAX          (PMA_CH2_REG_OOB_COMWAKE_GAP_MAX),          
    .CP_PMA_CH2_REG_OOB_COMINIT_GAP_MIN          (PMA_CH2_REG_OOB_COMINIT_GAP_MIN),          
    .CP_PMA_CH2_REG_OOB_COMINIT_GAP_MAX          (PMA_CH2_REG_OOB_COMINIT_GAP_MAX),          
    .CP_PMA_CH2_REG_RX_PIBUF_IC_TX               (PMA_CH2_REG_RX_PIBUF_IC_TX),               
    .CP_PMA_CH2_REG_COMWAKE_STATUS_CLEAR         (PMA_CH2_REG_COMWAKE_STATUS_CLEAR),         
    .CP_PMA_CH2_REG_COMINIT_STATUS_CLEAR         (PMA_CH2_REG_COMINIT_STATUS_CLEAR),         
    .CP_PMA_CH2_REG_RX_SYNC_RST_N_EN             (PMA_CH2_REG_RX_SYNC_RST_N_EN),             
    .CP_PMA_CH2_REG_RX_SYNC_RST_N                (PMA_CH2_REG_RX_SYNC_RST_N),                
    .CP_PMA_CH2_REG_RX_SATA_COMINIT_OW           (PMA_CH2_REG_RX_SATA_COMINIT_OW),           
    .CP_PMA_CH2_REG_RX_SATA_COMINIT              (PMA_CH2_REG_RX_SATA_COMINIT),              
    .CP_PMA_CH2_REG_RX_SATA_COMWAKE_OW           (PMA_CH2_REG_RX_SATA_COMWAKE_OW),           
    .CP_PMA_CH2_REG_RX_SATA_COMWAKE              (PMA_CH2_REG_RX_SATA_COMWAKE),              
    .CP_PMA_CH2_REG_RX_DCC_DISABLE               (PMA_CH2_REG_RX_DCC_DISABLE),               
    .CP_PMA_CH2_REG_TX_DCC_DISABLE               (PMA_CH2_REG_TX_DCC_DISABLE),               
    .CP_PMA_CH2_REG_RX_SLIP_SEL_EN               (PMA_CH2_REG_RX_SLIP_SEL_EN),               
    .CP_PMA_CH2_REG_RX_SLIP_SEL                  (PMA_CH2_REG_RX_SLIP_SEL),                  
    .CP_PMA_CH2_REG_RX_SLIP_EN                   (PMA_CH2_REG_RX_SLIP_EN),                   
    .CP_PMA_CH2_REG_RX_SIGDET_STATUS_SEL         (PMA_CH2_REG_RX_SIGDET_STATUS_SEL),         
    .CP_PMA_CH2_REG_RX_SIGDET_FSM_RST_N          (PMA_CH2_REG_RX_SIGDET_FSM_RST_N),          
    .CP_PMA_CH2_REG_RX_SIGDET_STATUS_OW          (PMA_CH2_REG_RX_SIGDET_STATUS_OW),          
    .CP_PMA_CH2_REG_RX_SIGDET_STATUS             (PMA_CH2_REG_RX_SIGDET_STATUS),             
    .CP_PMA_CH2_REG_RX_SIGDET_VTH                (PMA_CH2_REG_RX_SIGDET_VTH),                
    .CP_PMA_CH2_REG_RX_SIGDET_GRM                (PMA_CH2_REG_RX_SIGDET_GRM),                
    .CP_PMA_CH2_REG_RX_SIGDET_PULSE_EXT          (PMA_CH2_REG_RX_SIGDET_PULSE_EXT),          
    .CP_PMA_CH2_REG_RX_SIGDET_CH2_SEL            (PMA_CH2_REG_RX_SIGDET_CH2_SEL),            
    .CP_PMA_CH2_REG_RX_SIGDET_CH2_CHK_WINDOW     (PMA_CH2_REG_RX_SIGDET_CH2_CHK_WINDOW),     
    .CP_PMA_CH2_REG_RX_SIGDET_CHK_WINDOW_EN      (PMA_CH2_REG_RX_SIGDET_CHK_WINDOW_EN),      
    .CP_PMA_CH2_REG_RX_SIGDET_NOSIG_COUNT_SETTING(PMA_CH2_REG_RX_SIGDET_NOSIG_COUNT_SETTING),
    .CP_PMA_CH2_REG_RX_SIGDET_OOB_DET_COUNT_VAL  (PMA_CH2_REG_RX_SIGDET_OOB_DET_COUNT_VAL),  
    .CP_PMA_CH2_REG_SLIP_FIFO_INV_EN             (PMA_CH2_REG_SLIP_FIFO_INV_EN),             
    .CP_PMA_CH2_REG_SLIP_FIFO_INV                (PMA_CH2_REG_SLIP_FIFO_INV),                
    .CP_PMA_CH2_REG_RX_SIGDET_4OOB_DET_SEL       (PMA_CH2_REG_RX_SIGDET_4OOB_DET_SEL),       
    .CP_PMA_CH2_REG_RX_SIGDET_IC_I               (PMA_CH2_REG_RX_SIGDET_IC_I),               
    .CP_PMA_CH2_REG_RX_OOB_DETECTOR_RESET_N_OW   (PMA_CH2_REG_RX_OOB_DETECTOR_RESET_N_OW),   
    .CP_PMA_CH2_REG_RX_OOB_DETECTOR_RESET_N      (PMA_CH2_REG_RX_OOB_DETECTOR_RESET_N),      
    .CP_PMA_CH2_REG_RX_OOB_DETECTOR_PD_OW        (PMA_CH2_REG_RX_OOB_DETECTOR_PD_OW),        
    .CP_PMA_CH2_REG_RX_OOB_DETECTOR_PD           (PMA_CH2_REG_RX_OOB_DETECTOR_PD),           
    .CP_PMA_CH2_REG_RX_TERM_CM_CTRL              (PMA_CH2_REG_RX_TERM_CM_CTRL),              
    .CP_PMA_CH2_REG_TX_PD                        (PMA_CH2_REG_TX_PD),                        
    .CP_PMA_CH2_REG_TX_PD_OW                     (PMA_CH2_REG_TX_PD_OW),                     
    .CP_PMA_CH2_REG_TX_CLKPATH_PD                (PMA_CH2_REG_TX_CLKPATH_PD),                
    .CP_PMA_CH2_REG_TX_CLKPATH_PD_OW             (PMA_CH2_REG_TX_CLKPATH_PD_OW),             
    .CP_PMA_CH2_REG_TX_BEACON_TIMER_SEL          (PMA_CH2_REG_TX_BEACON_TIMER_SEL),          
    .CP_PMA_CH2_REG_TX_RXDET_REQ_OW              (PMA_CH2_REG_TX_RXDET_REQ_OW),              
    .CP_PMA_CH2_REG_TX_RXDET_REQ                 (PMA_CH2_REG_TX_RXDET_REQ),                 
    .CP_PMA_CH2_REG_TX_BEACON_EN_OW              (PMA_CH2_REG_TX_BEACON_EN_OW),              
    .CP_PMA_CH2_REG_TX_BEACON_EN                 (PMA_CH2_REG_TX_BEACON_EN),                 
    .CP_PMA_CH2_REG_TX_EI_EN_OW                  (PMA_CH2_REG_TX_EI_EN_OW),                  
    .CP_PMA_CH2_REG_TX_EI_EN                     (PMA_CH2_REG_TX_EI_EN),                     
    .CP_PMA_CH2_REG_TX_RES_CAL_EN                (PMA_CH2_REG_TX_RES_CAL_EN),                
    .CP_PMA_CH2_REG_TX_RES_CAL                   (PMA_CH2_REG_TX_RES_CAL),                   
    .CP_PMA_CH2_REG_TX_BIAS_CAL_EN               (PMA_CH2_REG_TX_BIAS_CAL_EN),               
    .CP_PMA_CH2_REG_TX_BIAS_CTRL                 (PMA_CH2_REG_TX_BIAS_CTRL),                 
    .CP_PMA_CH2_REG_TX_RXDET_TIMER_SEL           (PMA_CH2_REG_TX_RXDET_TIMER_SEL),           
    .CP_PMA_CH2_REG_TX_SYNC_OW                   (PMA_CH2_REG_TX_SYNC_OW),                   
    .CP_PMA_CH2_REG_TX_SYNC                      (PMA_CH2_REG_TX_SYNC),                      
    .CP_PMA_CH2_REG_TX_PD_POST                   (PMA_CH2_REG_TX_PD_POST),                   
    .CP_PMA_CH2_REG_TX_PD_POST_OW                (PMA_CH2_REG_TX_PD_POST_OW),                
    .CP_PMA_CH2_REG_TX_RESET_N_OW                (PMA_CH2_REG_TX_RESET_N_OW),                
    .CP_PMA_CH2_REG_TX_RESET_N                   (PMA_CH2_REG_TX_RESET_N),                   
    .CP_PMA_CH2_REG_TX_DCC_RESET_N_OW            (PMA_CH2_REG_TX_DCC_RESET_N_OW),            
    .CP_PMA_CH2_REG_TX_DCC_RESET_N               (PMA_CH2_REG_TX_DCC_RESET_N),               
    .CP_PMA_CH2_REG_TX_BUSWIDTH_OW               (PMA_CH2_REG_TX_BUSWIDTH_OW),               
    .CP_PMA_CH2_REG_TX_BUSWIDTH                  (PMA_CH2_REG_TX_BUSWIDTH),                  
    .CP_PMA_CH2_REG_PLL_READY_OW                 (PMA_CH2_REG_PLL_READY_OW),                 
    .CP_PMA_CH2_REG_PLL_READY                    (PMA_CH2_REG_PLL_READY),                    
    .CP_PMA_CH2_REG_TX_PCLK_SW_OW                (PMA_CH2_REG_TX_PCLK_SW_OW),                
    .CP_PMA_CH2_REG_TX_PCLK_SW                   (PMA_CH2_REG_TX_PCLK_SW),                   
    .CP_PMA_CH2_REG_EI_PCLK_DELAY_SEL            (PMA_CH2_REG_EI_PCLK_DELAY_SEL),            
    .CP_PMA_CH2_REG_TX_DRV01_DAC0                (PMA_CH2_REG_TX_DRV01_DAC0),                
    .CP_PMA_CH2_REG_TX_DRV01_DAC1                (PMA_CH2_REG_TX_DRV01_DAC1),                
    .CP_PMA_CH2_REG_TX_DRV01_DAC2                (PMA_CH2_REG_TX_DRV01_DAC2),                
    .CP_PMA_CH2_REG_TX_DRV00_DAC0                (PMA_CH2_REG_TX_DRV00_DAC0),                
    .CP_PMA_CH2_REG_TX_DRV00_DAC1                (PMA_CH2_REG_TX_DRV00_DAC1),                
    .CP_PMA_CH2_REG_TX_DRV00_DAC2                (PMA_CH2_REG_TX_DRV00_DAC2),                
    .CP_PMA_CH2_REG_TX_AMP0                      (PMA_CH2_REG_TX_AMP0),                      
    .CP_PMA_CH2_REG_TX_AMP1                      (PMA_CH2_REG_TX_AMP1),                      
    .CP_PMA_CH2_REG_TX_AMP2                      (PMA_CH2_REG_TX_AMP2),                      
    .CP_PMA_CH2_REG_TX_AMP3                      (PMA_CH2_REG_TX_AMP3),                      
    .CP_PMA_CH2_REG_TX_AMP4                      (PMA_CH2_REG_TX_AMP4),                      
    .CP_PMA_CH2_REG_TX_MARGIN                    (PMA_CH2_REG_TX_MARGIN),                    
    .CP_PMA_CH2_REG_TX_MARGIN_OW                 (PMA_CH2_REG_TX_MARGIN_OW),                 
    .CP_PMA_CH2_REG_TX_DEEMP                     (PMA_CH2_REG_TX_DEEMP),                     
    .CP_PMA_CH2_REG_TX_DEEMP_OW                  (PMA_CH2_REG_TX_DEEMP_OW),                  
    .CP_PMA_CH2_REG_TX_SWING                     (PMA_CH2_REG_TX_SWING),                     
    .CP_PMA_CH2_REG_TX_SWING_OW                  (PMA_CH2_REG_TX_SWING_OW),                  
    .CP_PMA_CH2_REG_TX_RXDET_THRESHOLD           (PMA_CH2_REG_TX_RXDET_THRESHOLD),           
    .CP_PMA_CH2_REG_TX_BEACON_OSC_CTRL           (PMA_CH2_REG_TX_BEACON_OSC_CTRL),           
    .CP_PMA_CH2_REG_TX_PREDRV_DAC                (PMA_CH2_REG_TX_PREDRV_DAC),                
    .CP_PMA_CH2_REG_TX_PREDRV_CM_CTRL            (PMA_CH2_REG_TX_PREDRV_CM_CTRL),            
    .CP_PMA_CH2_REG_TX_TX2RX_SLPBACK_EN          (PMA_CH2_REG_TX_TX2RX_SLPBACK_EN),          
    .CP_PMA_CH2_REG_TX_PCLK_EDGE_SEL             (PMA_CH2_REG_TX_PCLK_EDGE_SEL),             
    .CP_PMA_CH2_REG_TX_RXDET_STATUS_OW           (PMA_CH2_REG_TX_RXDET_STATUS_OW),           
    .CP_PMA_CH2_REG_TX_RXDET_STATUS              (PMA_CH2_REG_TX_RXDET_STATUS),              
    .CP_PMA_CH2_REG_TX_PRBS_GEN_EN               (PMA_CH2_REG_TX_PRBS_GEN_EN),               
    .CP_PMA_CH2_REG_TX_PRBS_GEN_WIDTH_SEL        (PMA_CH2_REG_TX_PRBS_GEN_WIDTH_SEL),        
    .CP_PMA_CH2_REG_TX_PRBS_SEL                  (PMA_CH2_REG_TX_PRBS_SEL),                  
    .CP_PMA_CH2_REG_TX_UDP_DATA                  (PMA_CH2_REG_TX_UDP_DATA),                  
    .CP_PMA_CH2_REG_TX_FIFO_RST_N                (PMA_CH2_REG_TX_FIFO_RST_N),                
    .CP_PMA_CH2_REG_TX_FIFO_WP_CTRL              (PMA_CH2_REG_TX_FIFO_WP_CTRL),              
    .CP_PMA_CH2_REG_TX_FIFO_EN                   (PMA_CH2_REG_TX_FIFO_EN),                   
    .CP_PMA_CH2_REG_TX_DATA_MUX_SEL              (PMA_CH2_REG_TX_DATA_MUX_SEL),              
    .CP_PMA_CH2_REG_TX_ERR_INSERT                (PMA_CH2_REG_TX_ERR_INSERT),                
    .CP_PMA_CH2_REG_TX_SATA_EN                   (PMA_CH2_REG_TX_SATA_EN),                             
    .CP_PMA_CH2_REG_RATE_CHANGE_TXPCLK_ON_OW     (PMA_CH2_REG_RATE_CHANGE_TXPCLK_ON_OW),     
    .CP_PMA_CH2_REG_RATE_CHANGE_TXPCLK_ON        (PMA_CH2_REG_RATE_CHANGE_TXPCLK_ON),        
    .CP_PMA_CH2_REG_TX_PULLUP_DAC0               (PMA_CH2_REG_TX_PULLUP_DAC0),               
    .CP_PMA_CH2_REG_TX_PULLUP_DAC1               (PMA_CH2_REG_TX_PULLUP_DAC1),               
    .CP_PMA_CH2_REG_TX_PULLUP_DAC2               (PMA_CH2_REG_TX_PULLUP_DAC2),               
    .CP_PMA_CH2_REG_TX_PULLUP_DAC3               (PMA_CH2_REG_TX_PULLUP_DAC3),               
    .CP_PMA_CH2_REG_TX_OOB_DELAY_SEL             (PMA_CH2_REG_TX_OOB_DELAY_SEL),             
    .CP_PMA_CH2_REG_TX_POLARITY                  (PMA_CH2_REG_TX_POLARITY),                  
    .CP_PMA_CH2_REG_TX_SLPBK_AMP                 (PMA_CH2_REG_TX_SLPBK_AMP),                 
    .CP_PMA_CH2_REG_TX_LS_MODE_EN                (PMA_CH2_REG_TX_LS_MODE_EN),                
    .CP_PMA_CH2_REG_TX_JTAG_MODE_EN_OW           (PMA_CH2_REG_TX_JTAG_MODE_EN_OW),           
    .CP_PMA_CH2_REG_TX_JTAG_MODE_EN              (PMA_CH2_REG_TX_JTAG_MODE_EN),              
    .CP_PMA_CH2_REG_RX_JTAG_MODE_EN_OW           (PMA_CH2_REG_RX_JTAG_MODE_EN_OW),           
    .CP_PMA_CH2_REG_RX_JTAG_MODE_EN              (PMA_CH2_REG_RX_JTAG_MODE_EN),              
    .CP_PMA_CH2_REG_RX_JTAG_OE                   (PMA_CH2_REG_RX_JTAG_OE),                   
    .CP_PMA_CH2_REG_RX_ACJTAG_VHYSTSE            (PMA_CH2_REG_RX_ACJTAG_VHYSTSE),            
    .CP_PMA_CH2_REG_TX_FBCLK_FAR_EN              (PMA_CH2_REG_TX_FBCLK_FAR_EN),              
    .CP_PMA_CH2_REG_RX_TERM_MODE_CTRL            (PMA_CH2_REG_RX_TERM_MODE_CTRL),            
    .CP_PMA_CH2_REG_PLPBK_TXPCLK_EN              (PMA_CH2_REG_PLPBK_TXPCLK_EN),              
    .CP_PMA_CH2_CFG_LANE_POWERUP                 (PMA_CH2_CFG_LANE_POWERUP),                 
    .CP_PMA_CH2_CFG_PMA_POR_N                    (PMA_CH2_CFG_PMA_POR_N),                    
    .CP_PMA_CH2_CFG_RX_LANE_POWERUP              (PMA_CH2_CFG_RX_LANE_POWERUP),              
    .CP_PMA_CH2_CFG_RX_PMA_RSTN                  (PMA_CH2_CFG_RX_PMA_RSTN),                  
    .CP_PMA_CH2_CFG_TX_LANE_POWERUP              (PMA_CH2_CFG_TX_LANE_POWERUP),              
    .CP_PMA_CH2_CFG_TX_PMA_RSTN                  (PMA_CH2_CFG_TX_PMA_RSTN),                  
    .CP_PMA_CH2_REG_RESERVED_48_45               (PMA_CH2_REG_RESERVED_48_45),               
    .CP_PMA_CH2_REG_RESERVED_69                  (PMA_CH2_REG_RESERVED_69),                  
    .CP_PMA_CH2_REG_RESERVED_77_76               (PMA_CH2_REG_RESERVED_77_76),               
    .CP_PMA_CH2_REG_RESERVED_171_164             (PMA_CH2_REG_RESERVED_171_164),             
    .CP_PMA_CH2_REG_RESERVED_175_172             (PMA_CH2_REG_RESERVED_175_172),             
    .CP_PMA_CH2_REG_RESERVED_190                 (PMA_CH2_REG_RESERVED_190),                 
    .CP_PMA_CH2_REG_RESERVED_233_232             (PMA_CH2_REG_RESERVED_233_232),             
    .CP_PMA_CH2_REG_RESERVED_235_234             (PMA_CH2_REG_RESERVED_235_234),             
    .CP_PMA_CH2_REG_RESERVED_241_240             (PMA_CH2_REG_RESERVED_241_240),             
    .CP_PMA_CH2_REG_RESERVED_285_283             (PMA_CH2_REG_RESERVED_285_283),             
    .CP_PMA_CH2_REG_RESERVED_286                 (PMA_CH2_REG_RESERVED_286),                 
    .CP_PMA_CH2_REG_RESERVED_295                 (PMA_CH2_REG_RESERVED_295),                 
    .CP_PMA_CH2_REG_RESERVED_298                 (PMA_CH2_REG_RESERVED_298),                 
    .CP_PMA_CH2_REG_RESERVED_332_325             (PMA_CH2_REG_RESERVED_332_325),             
    .CP_PMA_CH2_REG_RESERVED_340_333             (PMA_CH2_REG_RESERVED_340_333),             
    .CP_PMA_CH2_REG_RESERVED_348_341             (PMA_CH2_REG_RESERVED_348_341),             
    .CP_PMA_CH2_REG_RESERVED_354_349             (PMA_CH2_REG_RESERVED_354_349),             
    .CP_PMA_CH2_REG_RESERVED_373                 (PMA_CH2_REG_RESERVED_373),                 
    .CP_PMA_CH2_REG_RESERVED_376                 (PMA_CH2_REG_RESERVED_376),                 
    .CP_PMA_CH2_REG_RESERVED_452                 (PMA_CH2_REG_RESERVED_452),                 
    .CP_PMA_CH2_REG_RESERVED_502_499             (PMA_CH2_REG_RESERVED_502_499),             
    .CP_PMA_CH2_REG_RESERVED_506_505             (PMA_CH2_REG_RESERVED_506_505),             
    .CP_PMA_CH2_REG_RESERVED_550_549             (PMA_CH2_REG_RESERVED_550_549),             
    .CP_PMA_CH2_REG_RESERVED_556_552             (PMA_CH2_REG_RESERVED_556_552),             
    .CP_PMA_CH3_REG_RX_PD                        (PMA_CH3_REG_RX_PD),                        
    .CP_PMA_CH3_REG_RX_PD_EN                     (PMA_CH3_REG_RX_PD_EN),                     
    .CP_PMA_CH3_REG_RX_CLKPATH_PD                (PMA_CH3_REG_RX_CLKPATH_PD),                
    .CP_PMA_CH3_REG_RX_CLKPATH_PD_EN             (PMA_CH3_REG_RX_CLKPATH_PD_EN),             
    .CP_PMA_CH3_REG_RX_DATAPATH_PD               (PMA_CH3_REG_RX_DATAPATH_PD),               
    .CP_PMA_CH3_REG_RX_DATAPATH_PD_EN            (PMA_CH3_REG_RX_DATAPATH_PD_EN),            
    .CP_PMA_CH3_REG_RX_SIGDET_PD                 (PMA_CH3_REG_RX_SIGDET_PD),                 
    .CP_PMA_CH3_REG_RX_SIGDET_PD_EN              (PMA_CH3_REG_RX_SIGDET_PD_EN),              
    .CP_PMA_CH3_REG_RX_DCC_RST_N                 (PMA_CH3_REG_RX_DCC_RST_N),                 
    .CP_PMA_CH3_REG_RX_DCC_RST_N_EN              (PMA_CH3_REG_RX_DCC_RST_N_EN),              
    .CP_PMA_CH3_REG_RX_CDR_RST_N                 (PMA_CH3_REG_RX_CDR_RST_N),                 
    .CP_PMA_CH3_REG_RX_CDR_RST_N_EN              (PMA_CH3_REG_RX_CDR_RST_N_EN),              
    .CP_PMA_CH3_REG_RX_SIGDET_RST_N              (PMA_CH3_REG_RX_SIGDET_RST_N),              
    .CP_PMA_CH3_REG_RX_SIGDET_RST_N_EN           (PMA_CH3_REG_RX_SIGDET_RST_N_EN),           
    .CP_PMA_CH3_REG_RXPCLK_SLIP                  (PMA_CH3_REG_RXPCLK_SLIP),                  
    .CP_PMA_CH3_REG_RXPCLK_SLIP_OW               (PMA_CH3_REG_RXPCLK_SLIP_OW),               
    .CP_PMA_CH3_REG_RX_PCLKSWITCH_RST_N          (PMA_CH3_REG_RX_PCLKSWITCH_RST_N),          
    .CP_PMA_CH3_REG_RX_PCLKSWITCH_RST_N_EN       (PMA_CH3_REG_RX_PCLKSWITCH_RST_N_EN),       
    .CP_PMA_CH3_REG_RX_PCLKSWITCH                (PMA_CH3_REG_RX_PCLKSWITCH),                
    .CP_PMA_CH3_REG_RX_PCLKSWITCH_EN             (PMA_CH3_REG_RX_PCLKSWITCH_EN),             
    .CP_PMA_CH3_REG_RX_HIGHZ                     (PMA_CH3_REG_RX_HIGHZ),                     
    .CP_PMA_CH3_REG_RX_HIGHZ_EN                  (PMA_CH3_REG_RX_HIGHZ_EN),                  
    .CP_PMA_CH3_REG_RX_EQ_C_SET                  (PMA_CH3_REG_RX_EQ_C_SET),                  
    .CP_PMA_CH3_REG_RX_EQ_R_SET                  (PMA_CH3_REG_RX_EQ_R_SET),                  
    .CP_PMA_CH3_REG_RX_BUSWIDTH                  (PMA_CH3_REG_RX_BUSWIDTH),                  
    .CP_PMA_CH3_REG_RX_BUSWIDTH_EN               (PMA_CH3_REG_RX_BUSWIDTH_EN),               
    .CP_PMA_CH3_REG_RX_RATE                      (PMA_CH3_REG_RX_RATE),                      
    .CP_PMA_CH3_REG_RX_RATE_EN                   (PMA_CH3_REG_RX_RATE_EN),                   
    .CP_PMA_CH3_REG_RX_RES_TRIM                  (PMA_CH3_REG_RX_RES_TRIM),                  
    .CP_PMA_CH3_REG_RX_RES_TRIM_EN               (PMA_CH3_REG_RX_RES_TRIM_EN),               
    .CP_PMA_CH3_REG_RX_EQ_OFF                    (PMA_CH3_REG_RX_EQ_OFF),                    
    .CP_PMA_CH3_REG_RX_PREAMP_IC                 (PMA_CH3_REG_RX_PREAMP_IC),                 
    .CP_PMA_CH3_REG_RX_PCLK_EDGE_SEL             (PMA_CH3_REG_RX_PCLK_EDGE_SEL),             
    .CP_PMA_CH3_REG_RX_PIBUF_IC                  (PMA_CH3_REG_RX_PIBUF_IC),                  
    .CP_PMA_CH3_REG_RX_DCC_IC_RX                 (PMA_CH3_REG_RX_DCC_IC_RX),                 
    .CP_PMA_CH3_REG_RX_DCC_IC_TX                 (PMA_CH3_REG_RX_DCC_IC_TX),                 
    .CP_PMA_CH3_REG_RX_ICTRL_TRX                 (PMA_CH3_REG_RX_ICTRL_TRX),                 
    .CP_PMA_CH3_REG_RX_ICTRL_SIGDET              (PMA_CH3_REG_RX_ICTRL_SIGDET),              
    .CP_PMA_CH3_REG_RX_ICTRL_PREAMP              (PMA_CH3_REG_RX_ICTRL_PREAMP),              
    .CP_PMA_CH3_REG_RX_ICTRL_SLICER              (PMA_CH3_REG_RX_ICTRL_SLICER),              
    .CP_PMA_CH3_REG_RX_ICTRL_PIBUF               (PMA_CH3_REG_RX_ICTRL_PIBUF),               
    .CP_PMA_CH3_REG_RX_ICTRL_PI                  (PMA_CH3_REG_RX_ICTRL_PI),                  
    .CP_PMA_CH3_REG_RX_ICTRL_DCC                 (PMA_CH3_REG_RX_ICTRL_DCC),                 
    .CP_PMA_CH3_REG_RX_ICTRL_PREDRV              (PMA_CH3_REG_RX_ICTRL_PREDRV),              
    .CP_PMA_CH3_REG_TX_RATE                      (PMA_CH3_REG_TX_RATE),                      
    .CP_PMA_CH3_REG_TX_RATE_EN                   (PMA_CH3_REG_TX_RATE_EN),                   
    .CP_PMA_CH3_REG_RX_TX2RX_PLPBK_RST_N         (PMA_CH3_REG_RX_TX2RX_PLPBK_RST_N),         
    .CP_PMA_CH3_REG_RX_TX2RX_PLPBK_RST_N_EN      (PMA_CH3_REG_RX_TX2RX_PLPBK_RST_N_EN),      
    .CP_PMA_CH3_REG_RX_TX2RX_PLPBK_EN            (PMA_CH3_REG_RX_TX2RX_PLPBK_EN),            
    .CP_PMA_CH3_REG_TXCLK_SEL                    (PMA_CH3_REG_TXCLK_SEL),                    
    .CP_PMA_CH3_REG_RX_DATA_POLARITY             (PMA_CH3_REG_RX_DATA_POLARITY),             
    .CP_PMA_CH3_REG_RX_ERR_INSERT                (PMA_CH3_REG_RX_ERR_INSERT),                
    .CP_PMA_CH3_REG_UDP_CHK_EN                   (PMA_CH3_REG_UDP_CHK_EN),                   
    .CP_PMA_CH3_REG_PRBS_SEL                     (PMA_CH3_REG_PRBS_SEL),                     
    .CP_PMA_CH3_REG_PRBS_CHK_EN                  (PMA_CH3_REG_PRBS_CHK_EN),                  
    .CP_PMA_CH3_REG_PRBS_CHK_WIDTH_SEL           (PMA_CH3_REG_PRBS_CHK_WIDTH_SEL),           
    .CP_PMA_CH3_REG_BIST_CHK_PAT_SEL             (PMA_CH3_REG_BIST_CHK_PAT_SEL),             
    .CP_PMA_CH3_REG_LOAD_ERR_CNT                 (PMA_CH3_REG_LOAD_ERR_CNT),                 
    .CP_PMA_CH3_REG_CHK_COUNTER_EN               (PMA_CH3_REG_CHK_COUNTER_EN),               
    .CP_PMA_CH3_REG_CDR_PROP_GAIN                (PMA_CH3_REG_CDR_PROP_GAIN),                
    .CP_PMA_CH3_REG_CDR_PROP_TURBO_GAIN          (PMA_CH3_REG_CDR_PROP_TURBO_GAIN),          
    .CP_PMA_CH3_REG_CDR_INT_GAIN                 (PMA_CH3_REG_CDR_INT_GAIN),                 
    .CP_PMA_CH3_REG_CDR_INT_TURBO_GAIN           (PMA_CH3_REG_CDR_INT_TURBO_GAIN),           
    .CP_PMA_CH3_REG_CDR_INT_SAT_MAX              (PMA_CH3_REG_CDR_INT_SAT_MAX),              
    .CP_PMA_CH3_REG_CDR_INT_SAT_MIN              (PMA_CH3_REG_CDR_INT_SAT_MIN),              
    .CP_PMA_CH3_REG_CDR_INT_RST                  (PMA_CH3_REG_CDR_INT_RST),                  
    .CP_PMA_CH3_REG_CDR_INT_RST_OW               (PMA_CH3_REG_CDR_INT_RST_OW),               
    .CP_PMA_CH3_REG_CDR_PROP_RST                 (PMA_CH3_REG_CDR_PROP_RST),                 
    .CP_PMA_CH3_REG_CDR_PROP_RST_OW              (PMA_CH3_REG_CDR_PROP_RST_OW),              
    .CP_PMA_CH3_REG_CDR_LOCK_RST                 (PMA_CH3_REG_CDR_LOCK_RST),                 
    .CP_PMA_CH3_REG_CDR_LOCK_RST_OW              (PMA_CH3_REG_CDR_LOCK_RST_OW),              
    .CP_PMA_CH3_REG_CDR_RX_PI_FORCE_SEL          (PMA_CH3_REG_CDR_RX_PI_FORCE_SEL),          
    .CP_PMA_CH3_REG_CDR_RX_PI_FORCE_D            (PMA_CH3_REG_CDR_RX_PI_FORCE_D),            
    .CP_PMA_CH3_REG_CDR_LOCK_TIMER               (PMA_CH3_REG_CDR_LOCK_TIMER),               
    .CP_PMA_CH3_REG_CDR_TURBO_MODE_TIMER         (PMA_CH3_REG_CDR_TURBO_MODE_TIMER),         
    .CP_PMA_CH3_REG_CDR_LOCK_VAL                 (PMA_CH3_REG_CDR_LOCK_VAL),                 
    .CP_PMA_CH3_REG_CDR_LOCK_OW                  (PMA_CH3_REG_CDR_LOCK_OW),                  
    .CP_PMA_CH3_REG_CDR_INT_SAT_DET_EN           (PMA_CH3_REG_CDR_INT_SAT_DET_EN),           
    .CP_PMA_CH3_REG_CDR_SAT_DET_STATUS_EN        (PMA_CH3_REG_CDR_SAT_DET_STATUS_EN),        
    .CP_PMA_CH3_REG_CDR_SAT_DET_STATUS_RESET_EN  (PMA_CH3_REG_CDR_SAT_DET_STATUS_RESET_EN),  
    .CP_PMA_CH3_REG_CDR_PI_CTRL_RST              (PMA_CH3_REG_CDR_PI_CTRL_RST),              
    .CP_PMA_CH3_REG_CDR_PI_CTRL_RST_OW           (PMA_CH3_REG_CDR_PI_CTRL_RST_OW),           
    .CP_PMA_CH3_REG_CDR_SAT_DET_RST              (PMA_CH3_REG_CDR_SAT_DET_RST),              
    .CP_PMA_CH3_REG_CDR_SAT_DET_RST_OW           (PMA_CH3_REG_CDR_SAT_DET_RST_OW),           
    .CP_PMA_CH3_REG_CDR_SAT_DET_STICKY_RST       (PMA_CH3_REG_CDR_SAT_DET_STICKY_RST),       
    .CP_PMA_CH3_REG_CDR_SAT_DET_STICKY_RST_OW    (PMA_CH3_REG_CDR_SAT_DET_STICKY_RST_OW),    
    .CP_PMA_CH3_REG_CDR_SIGDET_STATUS_DIS        (PMA_CH3_REG_CDR_SIGDET_STATUS_DIS),        
    .CP_PMA_CH3_REG_CDR_SAT_DET_TIMER            (PMA_CH3_REG_CDR_SAT_DET_TIMER),            
    .CP_PMA_CH3_REG_CDR_SAT_DET_STATUS_VAL       (PMA_CH3_REG_CDR_SAT_DET_STATUS_VAL),       
    .CP_PMA_CH3_REG_CDR_SAT_DET_STATUS_OW        (PMA_CH3_REG_CDR_SAT_DET_STATUS_OW),       
    .CP_PMA_CH3_REG_CDR_TURBO_MODE_EN            (PMA_CH3_REG_CDR_TURBO_MODE_EN),            
    .CP_PMA_CH3_REG_CDR_STATUS_RADDR_INIT        (PMA_CH3_REG_CDR_STATUS_RADDR_INIT),        
    .CP_PMA_CH3_REG_CDR_STATUS_FIFO_EN           (PMA_CH3_REG_CDR_STATUS_FIFO_EN),           
    .CP_PMA_CH3_REG_PMA_TEST_SEL                 (PMA_CH3_REG_PMA_TEST_SEL),                 
    .CP_PMA_CH3_REG_OOB_COMWAKE_GAP_MIN          (PMA_CH3_REG_OOB_COMWAKE_GAP_MIN),          
    .CP_PMA_CH3_REG_OOB_COMWAKE_GAP_MAX          (PMA_CH3_REG_OOB_COMWAKE_GAP_MAX),          
    .CP_PMA_CH3_REG_OOB_COMINIT_GAP_MIN          (PMA_CH3_REG_OOB_COMINIT_GAP_MIN),          
    .CP_PMA_CH3_REG_OOB_COMINIT_GAP_MAX          (PMA_CH3_REG_OOB_COMINIT_GAP_MAX),          
    .CP_PMA_CH3_REG_RX_PIBUF_IC_TX               (PMA_CH3_REG_RX_PIBUF_IC_TX),               
    .CP_PMA_CH3_REG_COMWAKE_STATUS_CLEAR         (PMA_CH3_REG_COMWAKE_STATUS_CLEAR),         
    .CP_PMA_CH3_REG_COMINIT_STATUS_CLEAR         (PMA_CH3_REG_COMINIT_STATUS_CLEAR),         
    .CP_PMA_CH3_REG_RX_SYNC_RST_N_EN             (PMA_CH3_REG_RX_SYNC_RST_N_EN),             
    .CP_PMA_CH3_REG_RX_SYNC_RST_N                (PMA_CH3_REG_RX_SYNC_RST_N),                
    .CP_PMA_CH3_REG_RX_SATA_COMINIT_OW           (PMA_CH3_REG_RX_SATA_COMINIT_OW),           
    .CP_PMA_CH3_REG_RX_SATA_COMINIT              (PMA_CH3_REG_RX_SATA_COMINIT),              
    .CP_PMA_CH3_REG_RX_SATA_COMWAKE_OW           (PMA_CH3_REG_RX_SATA_COMWAKE_OW),           
    .CP_PMA_CH3_REG_RX_SATA_COMWAKE              (PMA_CH3_REG_RX_SATA_COMWAKE),              
    .CP_PMA_CH3_REG_RX_DCC_DISABLE               (PMA_CH3_REG_RX_DCC_DISABLE),               
    .CP_PMA_CH3_REG_TX_DCC_DISABLE               (PMA_CH3_REG_TX_DCC_DISABLE),               
    .CP_PMA_CH3_REG_RX_SLIP_SEL_EN               (PMA_CH3_REG_RX_SLIP_SEL_EN),               
    .CP_PMA_CH3_REG_RX_SLIP_SEL                  (PMA_CH3_REG_RX_SLIP_SEL),                  
    .CP_PMA_CH3_REG_RX_SLIP_EN                   (PMA_CH3_REG_RX_SLIP_EN),                   
    .CP_PMA_CH3_REG_RX_SIGDET_STATUS_SEL         (PMA_CH3_REG_RX_SIGDET_STATUS_SEL),         
    .CP_PMA_CH3_REG_RX_SIGDET_FSM_RST_N          (PMA_CH3_REG_RX_SIGDET_FSM_RST_N),          
    .CP_PMA_CH3_REG_RX_SIGDET_STATUS_OW          (PMA_CH3_REG_RX_SIGDET_STATUS_OW),          
    .CP_PMA_CH3_REG_RX_SIGDET_STATUS             (PMA_CH3_REG_RX_SIGDET_STATUS),             
    .CP_PMA_CH3_REG_RX_SIGDET_VTH                (PMA_CH3_REG_RX_SIGDET_VTH),                
    .CP_PMA_CH3_REG_RX_SIGDET_GRM                (PMA_CH3_REG_RX_SIGDET_GRM),                
    .CP_PMA_CH3_REG_RX_SIGDET_PULSE_EXT          (PMA_CH3_REG_RX_SIGDET_PULSE_EXT),          
    .CP_PMA_CH3_REG_RX_SIGDET_CH2_SEL            (PMA_CH3_REG_RX_SIGDET_CH2_SEL),            
    .CP_PMA_CH3_REG_RX_SIGDET_CH2_CHK_WINDOW     (PMA_CH3_REG_RX_SIGDET_CH2_CHK_WINDOW),     
    .CP_PMA_CH3_REG_RX_SIGDET_CHK_WINDOW_EN      (PMA_CH3_REG_RX_SIGDET_CHK_WINDOW_EN),      
    .CP_PMA_CH3_REG_RX_SIGDET_NOSIG_COUNT_SETTING(PMA_CH3_REG_RX_SIGDET_NOSIG_COUNT_SETTING),
    .CP_PMA_CH3_REG_RX_SIGDET_OOB_DET_COUNT_VAL  (PMA_CH3_REG_RX_SIGDET_OOB_DET_COUNT_VAL),
    .CP_PMA_CH3_REG_SLIP_FIFO_INV_EN             (PMA_CH3_REG_SLIP_FIFO_INV_EN),          
    .CP_PMA_CH3_REG_SLIP_FIFO_INV                (PMA_CH3_REG_SLIP_FIFO_INV),             
    .CP_PMA_CH3_REG_RX_SIGDET_4OOB_DET_SEL       (PMA_CH3_REG_RX_SIGDET_4OOB_DET_SEL),    
    .CP_PMA_CH3_REG_RX_SIGDET_IC_I               (PMA_CH3_REG_RX_SIGDET_IC_I),            
    .CP_PMA_CH3_REG_RX_OOB_DETECTOR_RESET_N_OW   (PMA_CH3_REG_RX_OOB_DETECTOR_RESET_N_OW),
    .CP_PMA_CH3_REG_RX_OOB_DETECTOR_RESET_N      (PMA_CH3_REG_RX_OOB_DETECTOR_RESET_N),   
    .CP_PMA_CH3_REG_RX_OOB_DETECTOR_PD_OW        (PMA_CH3_REG_RX_OOB_DETECTOR_PD_OW),     
    .CP_PMA_CH3_REG_RX_OOB_DETECTOR_PD           (PMA_CH3_REG_RX_OOB_DETECTOR_PD),        
    .CP_PMA_CH3_REG_RX_TERM_CM_CTRL              (PMA_CH3_REG_RX_TERM_CM_CTRL),           
    .CP_PMA_CH3_REG_TX_PD                        (PMA_CH3_REG_TX_PD),                     
    .CP_PMA_CH3_REG_TX_PD_OW                     (PMA_CH3_REG_TX_PD_OW),                  
    .CP_PMA_CH3_REG_TX_CLKPATH_PD                (PMA_CH3_REG_TX_CLKPATH_PD),             
    .CP_PMA_CH3_REG_TX_CLKPATH_PD_OW             (PMA_CH3_REG_TX_CLKPATH_PD_OW),          
    .CP_PMA_CH3_REG_TX_BEACON_TIMER_SEL          (PMA_CH3_REG_TX_BEACON_TIMER_SEL),       
    .CP_PMA_CH3_REG_TX_RXDET_REQ_OW              (PMA_CH3_REG_TX_RXDET_REQ_OW),           
    .CP_PMA_CH3_REG_TX_RXDET_REQ                 (PMA_CH3_REG_TX_RXDET_REQ),              
    .CP_PMA_CH3_REG_TX_BEACON_EN_OW              (PMA_CH3_REG_TX_BEACON_EN_OW),           
    .CP_PMA_CH3_REG_TX_BEACON_EN                 (PMA_CH3_REG_TX_BEACON_EN),              
    .CP_PMA_CH3_REG_TX_EI_EN_OW                  (PMA_CH3_REG_TX_EI_EN_OW),               
    .CP_PMA_CH3_REG_TX_EI_EN                     (PMA_CH3_REG_TX_EI_EN),                  
    .CP_PMA_CH3_REG_TX_RES_CAL_EN                (PMA_CH3_REG_TX_RES_CAL_EN),             
    .CP_PMA_CH3_REG_TX_RES_CAL                   (PMA_CH3_REG_TX_RES_CAL),                
    .CP_PMA_CH3_REG_TX_BIAS_CAL_EN               (PMA_CH3_REG_TX_BIAS_CAL_EN),            
    .CP_PMA_CH3_REG_TX_BIAS_CTRL                 (PMA_CH3_REG_TX_BIAS_CTRL),              
    .CP_PMA_CH3_REG_TX_RXDET_TIMER_SEL           (PMA_CH3_REG_TX_RXDET_TIMER_SEL),        
    .CP_PMA_CH3_REG_TX_SYNC_OW                   (PMA_CH3_REG_TX_SYNC_OW),                
    .CP_PMA_CH3_REG_TX_SYNC                      (PMA_CH3_REG_TX_SYNC),                   
    .CP_PMA_CH3_REG_TX_PD_POST                   (PMA_CH3_REG_TX_PD_POST),                
    .CP_PMA_CH3_REG_TX_PD_POST_OW                (PMA_CH3_REG_TX_PD_POST_OW),             
    .CP_PMA_CH3_REG_TX_RESET_N_OW                (PMA_CH3_REG_TX_RESET_N_OW),             
    .CP_PMA_CH3_REG_TX_RESET_N                   (PMA_CH3_REG_TX_RESET_N),                
    .CP_PMA_CH3_REG_TX_DCC_RESET_N_OW            (PMA_CH3_REG_TX_DCC_RESET_N_OW),         
    .CP_PMA_CH3_REG_TX_DCC_RESET_N               (PMA_CH3_REG_TX_DCC_RESET_N),            
    .CP_PMA_CH3_REG_TX_BUSWIDTH_OW               (PMA_CH3_REG_TX_BUSWIDTH_OW),            
    .CP_PMA_CH3_REG_TX_BUSWIDTH                  (PMA_CH3_REG_TX_BUSWIDTH),               
    .CP_PMA_CH3_REG_PLL_READY_OW                 (PMA_CH3_REG_PLL_READY_OW),              
    .CP_PMA_CH3_REG_PLL_READY                    (PMA_CH3_REG_PLL_READY),                 
    .CP_PMA_CH3_REG_TX_PCLK_SW_OW                (PMA_CH3_REG_TX_PCLK_SW_OW),             
    .CP_PMA_CH3_REG_TX_PCLK_SW                   (PMA_CH3_REG_TX_PCLK_SW),                
    .CP_PMA_CH3_REG_EI_PCLK_DELAY_SEL            (PMA_CH3_REG_EI_PCLK_DELAY_SEL),         
    .CP_PMA_CH3_REG_TX_DRV01_DAC0                (PMA_CH3_REG_TX_DRV01_DAC0),             
    .CP_PMA_CH3_REG_TX_DRV01_DAC1                (PMA_CH3_REG_TX_DRV01_DAC1),             
    .CP_PMA_CH3_REG_TX_DRV01_DAC2                (PMA_CH3_REG_TX_DRV01_DAC2),             
    .CP_PMA_CH3_REG_TX_DRV00_DAC0                (PMA_CH3_REG_TX_DRV00_DAC0),             
    .CP_PMA_CH3_REG_TX_DRV00_DAC1                (PMA_CH3_REG_TX_DRV00_DAC1),             
    .CP_PMA_CH3_REG_TX_DRV00_DAC2                (PMA_CH3_REG_TX_DRV00_DAC2),             
    .CP_PMA_CH3_REG_TX_AMP0                      (PMA_CH3_REG_TX_AMP0),                   
    .CP_PMA_CH3_REG_TX_AMP1                      (PMA_CH3_REG_TX_AMP1),                   
    .CP_PMA_CH3_REG_TX_AMP2                      (PMA_CH3_REG_TX_AMP2),                   
    .CP_PMA_CH3_REG_TX_AMP3                      (PMA_CH3_REG_TX_AMP3),                   
    .CP_PMA_CH3_REG_TX_AMP4                      (PMA_CH3_REG_TX_AMP4),                   
    .CP_PMA_CH3_REG_TX_MARGIN                    (PMA_CH3_REG_TX_MARGIN),                 
    .CP_PMA_CH3_REG_TX_MARGIN_OW                 (PMA_CH3_REG_TX_MARGIN_OW),              
    .CP_PMA_CH3_REG_TX_DEEMP                     (PMA_CH3_REG_TX_DEEMP),                  
    .CP_PMA_CH3_REG_TX_DEEMP_OW                  (PMA_CH3_REG_TX_DEEMP_OW),               
    .CP_PMA_CH3_REG_TX_SWING                     (PMA_CH3_REG_TX_SWING),                  
    .CP_PMA_CH3_REG_TX_SWING_OW                  (PMA_CH3_REG_TX_SWING_OW),               
    .CP_PMA_CH3_REG_TX_RXDET_THRESHOLD           (PMA_CH3_REG_TX_RXDET_THRESHOLD),        
    .CP_PMA_CH3_REG_TX_BEACON_OSC_CTRL           (PMA_CH3_REG_TX_BEACON_OSC_CTRL),        
    .CP_PMA_CH3_REG_TX_PREDRV_DAC                (PMA_CH3_REG_TX_PREDRV_DAC),             
    .CP_PMA_CH3_REG_TX_PREDRV_CM_CTRL            (PMA_CH3_REG_TX_PREDRV_CM_CTRL),         
    .CP_PMA_CH3_REG_TX_TX2RX_SLPBACK_EN          (PMA_CH3_REG_TX_TX2RX_SLPBACK_EN),       
    .CP_PMA_CH3_REG_TX_PCLK_EDGE_SEL             (PMA_CH3_REG_TX_PCLK_EDGE_SEL),          
    .CP_PMA_CH3_REG_TX_RXDET_STATUS_OW           (PMA_CH3_REG_TX_RXDET_STATUS_OW),        
    .CP_PMA_CH3_REG_TX_RXDET_STATUS              (PMA_CH3_REG_TX_RXDET_STATUS),           
    .CP_PMA_CH3_REG_TX_PRBS_GEN_EN               (PMA_CH3_REG_TX_PRBS_GEN_EN),            
    .CP_PMA_CH3_REG_TX_PRBS_GEN_WIDTH_SEL        (PMA_CH3_REG_TX_PRBS_GEN_WIDTH_SEL),     
    .CP_PMA_CH3_REG_TX_PRBS_SEL                  (PMA_CH3_REG_TX_PRBS_SEL),               
    .CP_PMA_CH3_REG_TX_UDP_DATA                  (PMA_CH3_REG_TX_UDP_DATA),               
    .CP_PMA_CH3_REG_TX_FIFO_RST_N                (PMA_CH3_REG_TX_FIFO_RST_N),             
    .CP_PMA_CH3_REG_TX_FIFO_WP_CTRL              (PMA_CH3_REG_TX_FIFO_WP_CTRL),           
    .CP_PMA_CH3_REG_TX_FIFO_EN                   (PMA_CH3_REG_TX_FIFO_EN),                
    .CP_PMA_CH3_REG_TX_DATA_MUX_SEL              (PMA_CH3_REG_TX_DATA_MUX_SEL),           
    .CP_PMA_CH3_REG_TX_ERR_INSERT                (PMA_CH3_REG_TX_ERR_INSERT),             
    .CP_PMA_CH3_REG_TX_SATA_EN                   (PMA_CH3_REG_TX_SATA_EN),                
    .CP_PMA_CH3_REG_RATE_CHANGE_TXPCLK_ON_OW     (PMA_CH3_REG_RATE_CHANGE_TXPCLK_ON_OW),  
    .CP_PMA_CH3_REG_RATE_CHANGE_TXPCLK_ON        (PMA_CH3_REG_RATE_CHANGE_TXPCLK_ON),     
    .CP_PMA_CH3_REG_TX_PULLUP_DAC0               (PMA_CH3_REG_TX_PULLUP_DAC0),            
    .CP_PMA_CH3_REG_TX_PULLUP_DAC1               (PMA_CH3_REG_TX_PULLUP_DAC1),            
    .CP_PMA_CH3_REG_TX_PULLUP_DAC2               (PMA_CH3_REG_TX_PULLUP_DAC2),            
    .CP_PMA_CH3_REG_TX_PULLUP_DAC3               (PMA_CH3_REG_TX_PULLUP_DAC3),            
    .CP_PMA_CH3_REG_TX_OOB_DELAY_SEL             (PMA_CH3_REG_TX_OOB_DELAY_SEL),          
    .CP_PMA_CH3_REG_TX_POLARITY                  (PMA_CH3_REG_TX_POLARITY),               
    .CP_PMA_CH3_REG_TX_SLPBK_AMP                 (PMA_CH3_REG_TX_SLPBK_AMP),              
    .CP_PMA_CH3_REG_TX_LS_MODE_EN                (PMA_CH3_REG_TX_LS_MODE_EN),             
    .CP_PMA_CH3_REG_TX_JTAG_MODE_EN_OW           (PMA_CH3_REG_TX_JTAG_MODE_EN_OW),        
    .CP_PMA_CH3_REG_TX_JTAG_MODE_EN              (PMA_CH3_REG_TX_JTAG_MODE_EN),           
    .CP_PMA_CH3_REG_RX_JTAG_MODE_EN_OW           (PMA_CH3_REG_RX_JTAG_MODE_EN_OW),        
    .CP_PMA_CH3_REG_RX_JTAG_MODE_EN              (PMA_CH3_REG_RX_JTAG_MODE_EN),           
    .CP_PMA_CH3_REG_RX_JTAG_OE                   (PMA_CH3_REG_RX_JTAG_OE),                
    .CP_PMA_CH3_REG_RX_ACJTAG_VHYSTSE            (PMA_CH3_REG_RX_ACJTAG_VHYSTSE),         
    .CP_PMA_CH3_REG_TX_FBCLK_FAR_EN              (PMA_CH3_REG_TX_FBCLK_FAR_EN),           
    .CP_PMA_CH3_REG_RX_TERM_MODE_CTRL            (PMA_CH3_REG_RX_TERM_MODE_CTRL),         
    .CP_PMA_CH3_REG_PLPBK_TXPCLK_EN              (PMA_CH3_REG_PLPBK_TXPCLK_EN),           
    .CP_PMA_CH3_CFG_LANE_POWERUP                 (PMA_CH3_CFG_LANE_POWERUP),              
    .CP_PMA_CH3_CFG_PMA_POR_N                    (PMA_CH3_CFG_PMA_POR_N),                 
    .CP_PMA_CH3_CFG_RX_LANE_POWERUP              (PMA_CH3_CFG_RX_LANE_POWERUP),           
    .CP_PMA_CH3_CFG_RX_PMA_RSTN                  (PMA_CH3_CFG_RX_PMA_RSTN),               
    .CP_PMA_CH3_CFG_TX_LANE_POWERUP              (PMA_CH3_CFG_TX_LANE_POWERUP),           
    .CP_PMA_CH3_CFG_TX_PMA_RSTN                  (PMA_CH3_CFG_TX_PMA_RSTN),               
    .CP_PMA_CH3_REG_RESERVED_48_45               (PMA_CH3_REG_RESERVED_48_45),            
    .CP_PMA_CH3_REG_RESERVED_69                  (PMA_CH3_REG_RESERVED_69),               
    .CP_PMA_CH3_REG_RESERVED_77_76               (PMA_CH3_REG_RESERVED_77_76),            
    .CP_PMA_CH3_REG_RESERVED_171_164             (PMA_CH3_REG_RESERVED_171_164),          
    .CP_PMA_CH3_REG_RESERVED_175_172             (PMA_CH3_REG_RESERVED_175_172),          
    .CP_PMA_CH3_REG_RESERVED_190                 (PMA_CH3_REG_RESERVED_190),              
    .CP_PMA_CH3_REG_RESERVED_233_232             (PMA_CH3_REG_RESERVED_233_232),          
    .CP_PMA_CH3_REG_RESERVED_235_234             (PMA_CH3_REG_RESERVED_235_234),          
    .CP_PMA_CH3_REG_RESERVED_241_240             (PMA_CH3_REG_RESERVED_241_240),          
    .CP_PMA_CH3_REG_RESERVED_285_283             (PMA_CH3_REG_RESERVED_285_283),          
    .CP_PMA_CH3_REG_RESERVED_286                 (PMA_CH3_REG_RESERVED_286),              
    .CP_PMA_CH3_REG_RESERVED_295                 (PMA_CH3_REG_RESERVED_295),              
    .CP_PMA_CH3_REG_RESERVED_298                 (PMA_CH3_REG_RESERVED_298),              
    .CP_PMA_CH3_REG_RESERVED_332_325             (PMA_CH3_REG_RESERVED_332_325),          
    .CP_PMA_CH3_REG_RESERVED_340_333             (PMA_CH3_REG_RESERVED_340_333),          
    .CP_PMA_CH3_REG_RESERVED_348_341             (PMA_CH3_REG_RESERVED_348_341),          
    .CP_PMA_CH3_REG_RESERVED_354_349             (PMA_CH3_REG_RESERVED_354_349),          
    .CP_PMA_CH3_REG_RESERVED_373                 (PMA_CH3_REG_RESERVED_373),              
    .CP_PMA_CH3_REG_RESERVED_376                 (PMA_CH3_REG_RESERVED_376),              
    .CP_PMA_CH3_REG_RESERVED_452                 (PMA_CH3_REG_RESERVED_452),              
    .CP_PMA_CH3_REG_RESERVED_502_499             (PMA_CH3_REG_RESERVED_502_499),          
    .CP_PMA_CH3_REG_RESERVED_506_505             (PMA_CH3_REG_RESERVED_506_505),          
    .CP_PMA_CH3_REG_RESERVED_550_549             (PMA_CH3_REG_RESERVED_550_549),          
    .CP_PMA_CH3_REG_RESERVED_556_552             (PMA_CH3_REG_RESERVED_556_552),          
    .CP_PMA_PLL0_REG_PLL_POWERDOWN_OW            (PMA_PLL0_REG_PLL_POWERDOWN_OW),         
    .CP_PMA_PLL0_REG_PLL_POWERDOWN               (PMA_PLL0_REG_PLL_POWERDOWN),            
    .CP_PMA_PLL0_REG_PLL_RESET_N_OW              (PMA_PLL0_REG_PLL_RESET_N_OW),           
    .CP_PMA_PLL0_REG_PLL_RESET_N                 (PMA_PLL0_REG_PLL_RESET_N),              
    .CP_PMA_PLL0_REG_PLL_READY_OW                (PMA_PLL0_REG_PLL_READY_OW),             
    .CP_PMA_PLL0_REG_PLL_READY                   (PMA_PLL0_REG_PLL_READY),                
    .CP_PMA_PLL0_REG_LANE_SYNC_OW                (PMA_PLL0_REG_LANE_SYNC_OW),             
    .CP_PMA_PLL0_REG_LANE_SYNC                   (PMA_PLL0_REG_LANE_SYNC),                
    .CP_PMA_PLL0_REG_LOCKDET_REPEAT              (PMA_PLL0_REG_LOCKDET_REPEAT),           
    .CP_PMA_PLL0_REG_RESCAL_I_CODE_PMA           (PMA_PLL0_REG_RESCAL_I_CODE_PMA),        
    .CP_PMA_PLL0_REG_RESCAL_RESET_N_OW           (PMA_PLL0_REG_RESCAL_RESET_N_OW),        
    .CP_PMA_PLL0_REG_RESCAL_RESET_N              (PMA_PLL0_REG_RESCAL_RESET_N),           
    .CP_PMA_PLL0_REG_RESCAL_DONE_OW              (PMA_PLL0_REG_RESCAL_DONE_OW),           
    .CP_PMA_PLL0_REG_RESCAL_DONE                 (PMA_PLL0_REG_RESCAL_DONE),              
    .CP_PMA_PLL0_REG_RESCAL_CODE_OW              (PMA_PLL0_REG_RESCAL_CODE_OW),           
    .CP_PMA_PLL0_REG_LDO_VREF_SEL                (PMA_PLL0_REG_LDO_VREF_SEL),             
    .CP_PMA_PLL0_REG_BIAS_VCOREP_C               (PMA_PLL0_REG_BIAS_VCOREP_C),            
    .CP_PMA_PLL0_REG_RESCAL_I_CODE               (PMA_PLL0_REG_RESCAL_I_CODE),            
    .CP_PMA_PLL0_REG_RESCAL_ONCHIP_SMALL_OW      (PMA_PLL0_REG_RESCAL_ONCHIP_SMALL_OW),   
    .CP_PMA_PLL0_REG_RESCAL_ONCHIP_SMALL         (PMA_PLL0_REG_RESCAL_ONCHIP_SMALL),      
    .CP_PMA_PLL0_REG_JTAG_OE                     (PMA_PLL0_REG_JTAG_OE),                  
    .CP_PMA_PLL0_REG_JTAG_AC_MODE                (PMA_PLL0_REG_JTAG_AC_MODE),             
    .CP_PMA_PLL0_REG_JTAG_VHYSTSEL               (PMA_PLL0_REG_JTAG_VHYSTSEL),            
    .CP_PMA_PLL0_REG_PLL_LOCKDET_EN_OW           (PMA_PLL0_REG_PLL_LOCKDET_EN_OW),        
    .CP_PMA_PLL0_REG_PLL_LOCKDET_EN              (PMA_PLL0_REG_PLL_LOCKDET_EN),           
    .CP_PMA_PLL0_REG_PLL_LOCKDET_RESET_N_OW      (PMA_PLL0_REG_PLL_LOCKDET_RESET_N_OW),   
    .CP_PMA_PLL0_REG_PLL_LOCKDET_RESET_N         (PMA_PLL0_REG_PLL_LOCKDET_RESET_N),      
    .CP_PMA_PLL0_REG_PLL_LOCKED_OW               (PMA_PLL0_REG_PLL_LOCKED_OW),            
    .CP_PMA_PLL0_REG_PLL_LOCKED                  (PMA_PLL0_REG_PLL_LOCKED),               
    .CP_PMA_PLL0_REG_PLL_LOCKED_STICKY_CLEAR     (PMA_PLL0_REG_PLL_LOCKED_STICKY_CLEAR),  
    .CP_PMA_PLL0_REG_PLL_UNLOCKED_STICKY_CLEAR   (PMA_PLL0_REG_PLL_UNLOCKED_STICKY_CLEAR),
    .CP_PMA_PLL0_REG_NOFBCLK_STICKY_CLEAR        (PMA_PLL0_REG_NOFBCLK_STICKY_CLEAR),     
    .CP_PMA_PLL0_REG_PLL_LOCKDET_REFCT           (PMA_PLL0_REG_PLL_LOCKDET_REFCT),        
    .CP_PMA_PLL0_REG_PLL_LOCKDET_FBCT            (PMA_PLL0_REG_PLL_LOCKDET_FBCT),         
    .CP_PMA_PLL0_REG_PLL_LOCKDET_LOCKCT          (PMA_PLL0_REG_PLL_LOCKDET_LOCKCT),       
    .CP_PMA_PLL0_REG_PLL_LOCKDET_ITER            (PMA_PLL0_REG_PLL_LOCKDET_ITER),         
    .CP_PMA_PLL0_REG_PLL_UNLOCKDET_ITER          (PMA_PLL0_REG_PLL_UNLOCKDET_ITER),       
    .CP_PMA_PLL0_REG_PD_VCO                      (PMA_PLL0_REG_PD_VCO),                   
    .CP_PMA_PLL0_REG_FBCLK_TEST_EN               (PMA_PLL0_REG_FBCLK_TEST_EN),            
    .CP_PMA_PLL0_REG_REFCLK_TEST_EN              (PMA_PLL0_REG_REFCLK_TEST_EN),           
    .CP_PMA_PLL0_REG_TEST_SEL                    (PMA_PLL0_REG_TEST_SEL),                 
    .CP_PMA_PLL0_REG_TEST_V_EN                   (PMA_PLL0_REG_TEST_V_EN),                
    .CP_PMA_PLL0_REG_TEST_SIG_HALF_EN            (PMA_PLL0_REG_TEST_SIG_HALF_EN),         
    .CP_PMA_PLL0_REG_TEST_FSM                    (PMA_PLL0_REG_TEST_FSM),                 
    .CP_PMA_PLL0_REG_REFCLK_OUT_PD               (PMA_PLL0_REG_REFCLK_OUT_PD),            
    .CP_PMA_PLL0_REG_BGR_STARTUP_EN              (PMA_PLL0_REG_BGR_STARTUP_EN),           
    .CP_PMA_PLL0_REG_BGR_STARTUP                 (PMA_PLL0_REG_BGR_STARTUP),              
    .CP_PMA_PLL0_REG_PD_BGR                      (PMA_PLL0_REG_PD_BGR),                   
    .CP_PMA_PLL0_REG_REFCLK_TERM_VCM_EN          (PMA_PLL0_REG_REFCLK_TERM_VCM_EN),       
    .CP_PMA_PLL0_REG_FBDIVA_5_EN                 (PMA_PLL0_REG_FBDIVA_5_EN),              
    .CP_PMA_PLL0_REG_FBDIVB                      (PMA_PLL0_REG_FBDIVB),                   
    .CP_PMA_PLL0_REG_RESET_N_PFDQP_OW            (PMA_PLL0_REG_RESET_N_PFDQP_OW),         
    .CP_PMA_PLL0_REG_RESET_N_PFDQP               (PMA_PLL0_REG_RESET_N_PFDQP),            
    .CP_PMA_PLL0_REG_QPCURRENT                   (PMA_PLL0_REG_QPCURRENT),                
    .CP_PMA_PLL0_REG_VC_FORCE_EN                 (PMA_PLL0_REG_VC_FORCE_EN),              
    .CP_PMA_PLL0_REG_VCRESET_C_RING              (PMA_PLL0_REG_VCRESET_C_RING),           
    .CP_PMA_PLL0_REG_LPF_R_C                     (PMA_PLL0_REG_LPF_R_C),                  
    .CP_PMA_PLL0_REG_LPF_TR_C                    (PMA_PLL0_REG_LPF_TR_C),                 
    .CP_PMA_PLL0_REG_PD_BIAS                     (PMA_PLL0_REG_PD_BIAS),                  
    .CP_PMA_PLL0_REG_ICTRL_PLL                   (PMA_PLL0_REG_ICTRL_PLL),                
    .CP_PMA_PLL0_REG_BIAS_QP                     (PMA_PLL0_REG_BIAS_QP),                  
    .CP_PMA_PLL0_REG_BIAS_LANE_SYNC              (PMA_PLL0_REG_BIAS_LANE_SYNC),           
    .CP_PMA_PLL0_REG_BIAS_CLKBUFS1               (PMA_PLL0_REG_BIAS_CLKBUFS1),            
    .CP_PMA_PLL0_REG_TXPCLK_SEL                  (PMA_PLL0_REG_TXPCLK_SEL),               
    .CP_PMA_PLL0_REG_BIAS_CLKBUFS3               (PMA_PLL0_REG_BIAS_CLKBUFS3),            
    .CP_PMA_PLL0_REG_LANE_SYNC_EN                (PMA_PLL0_REG_LANE_SYNC_EN),             
    .CP_PMA_PLL0_REG_LANE_SYNC_EN_OW             (PMA_PLL0_REG_LANE_SYNC_EN_OW),          
    .CP_PMA_PLL0_REG_BIAS_D2S                    (PMA_PLL0_REG_BIAS_D2S),                 
    .CP_PMA_PLL0_REG_BIAS_REFD2S_C               (PMA_PLL0_REG_BIAS_REFD2S_C),            
    .CP_PMA_PLL0_REG_BIAS_VCRST_C                (PMA_PLL0_REG_BIAS_VCRST_C),             
    .CP_PMA_PLL0_REG_BIAS_REFBUF_C               (PMA_PLL0_REG_BIAS_REFBUF_C),            
    .CP_PMA_PLL0_REG_CLKBUFS1_C                  (PMA_PLL0_REG_CLKBUFS1_C),               
    .CP_PMA_PLL0_REG_CLKBUFS2_C                  (PMA_PLL0_REG_CLKBUFS2_C),               
    .CP_PMA_PLL0_REG_CLKBUFS3_C                  (PMA_PLL0_REG_CLKBUFS3_C),               
    .CP_PMA_PLL0_REG_CLKBUFS4_C                  (PMA_PLL0_REG_CLKBUFS4_C),               
    .CP_PMA_PLL0_REG_PLL_REFCLK_CML_SEL          (PMA_PLL0_REG_PLL_REFCLK_CML_SEL),      
    .CP_PMA_PLL0_REG_REFCLK_SEL                  (PMA_PLL0_REG_REFCLK_SEL),               
    .CP_PMA_PLL0_REG_RESCAL_R_CODE_SIGN          (PMA_PLL0_REG_RESCAL_R_CODE_SIGN),       
    .CP_PMA_PLL0_REG_PLL_UNLOCKED_OW             (PMA_PLL0_REG_PLL_UNLOCKED_OW),          
    .CP_PMA_PLL0_REG_PLL_UNLOCKED                (PMA_PLL0_REG_PLL_UNLOCKED),             
    .CP_PMA_PLL0_REG_PLL_LOCKDET_MODE            (PMA_PLL0_REG_PLL_LOCKDET_MODE),         
    .CP_PMA_PLL0_REG_PLL_CLKBUF_PD_LEFT          (PMA_PLL0_REG_PLL_CLKBUF_PD_LEFT),       
    .CP_PMA_PLL0_REG_PLL_CLKBUF_PD_RIGHT         (PMA_PLL0_REG_PLL_CLKBUF_PD_RIGHT),      
    .CP_PMA_PLL0_REG_RESCAL_EN                   (PMA_PLL0_REG_RESCAL_EN),                
    .CP_PMA_PLL0_REG_RESCAL_I_CODE_VAL           (PMA_PLL0_REG_RESCAL_I_CODE_VAL),        
    .CP_PMA_PLL0_REG_RESCAL_I_CODE_OW            (PMA_PLL0_REG_RESCAL_I_CODE_OW),         
    .CP_PMA_PLL0_REG_RESCAL_ITER_VALID_SEL       (PMA_PLL0_REG_RESCAL_ITER_VALID_SEL),    
    .CP_PMA_PLL0_REG_RESCAL_WAIT_SEL             (PMA_PLL0_REG_RESCAL_WAIT_SEL),          
    .CP_PMA_PLL0_REG_I_CTRL_MAX                  (PMA_PLL0_REG_I_CTRL_MAX),               
    .CP_PMA_PLL0_REG_I_CTRL_MIN                  (PMA_PLL0_REG_I_CTRL_MIN),               
    .CP_PARM_CFG_HSST_RSTN                       (PARM_CFG_HSST_RSTN),                    
    .CP_PARM_PLL0_POWERUP                        (PARM_PLL0_POWERUP),                     
    .CP_PARM_PLL0_RSTN                           (PARM_PLL0_RSTN),                        
    .CP_PMA_PLL1_REG_PLL_POWERDOWN_OW            (PMA_PLL1_REG_PLL_POWERDOWN_OW),         
    .CP_PMA_PLL1_REG_PLL_POWERDOWN               (PMA_PLL1_REG_PLL_POWERDOWN),            
    .CP_PMA_PLL1_REG_PLL_RESET_N_OW              (PMA_PLL1_REG_PLL_RESET_N_OW),           
    .CP_PMA_PLL1_REG_PLL_RESET_N                 (PMA_PLL1_REG_PLL_RESET_N),              
    .CP_PMA_PLL1_REG_PLL_READY_OW                (PMA_PLL1_REG_PLL_READY_OW),             
    .CP_PMA_PLL1_REG_PLL_READY                   (PMA_PLL1_REG_PLL_READY),                
    .CP_PMA_PLL1_REG_LANE_SYNC_OW                (PMA_PLL1_REG_LANE_SYNC_OW),             
    .CP_PMA_PLL1_REG_LANE_SYNC                   (PMA_PLL1_REG_LANE_SYNC),                
    .CP_PMA_PLL1_REG_LOCKDET_REPEAT              (PMA_PLL1_REG_LOCKDET_REPEAT),           
    .CP_PMA_PLL1_REG_RESCAL_I_CODE_PMA           (PMA_PLL1_REG_RESCAL_I_CODE_PMA),        
    .CP_PMA_PLL1_REG_RESCAL_RESET_N_OW           (PMA_PLL1_REG_RESCAL_RESET_N_OW),        
    .CP_PMA_PLL1_REG_RESCAL_RESET_N              (PMA_PLL1_REG_RESCAL_RESET_N),           
    .CP_PMA_PLL1_REG_RESCAL_DONE_OW              (PMA_PLL1_REG_RESCAL_DONE_OW),           
    .CP_PMA_PLL1_REG_RESCAL_DONE                 (PMA_PLL1_REG_RESCAL_DONE),              
    .CP_PMA_PLL1_REG_RESCAL_CODE_OW              (PMA_PLL1_REG_RESCAL_CODE_OW),           
    .CP_PMA_PLL1_REG_LDO_VREF_SEL                (PMA_PLL1_REG_LDO_VREF_SEL),             
    .CP_PMA_PLL1_REG_BIAS_VCOREP_C               (PMA_PLL1_REG_BIAS_VCOREP_C),            
    .CP_PMA_PLL1_REG_RESCAL_I_CODE               (PMA_PLL1_REG_RESCAL_I_CODE),            
    .CP_PMA_PLL1_REG_RESCAL_ONCHIP_SMALL_OW      (PMA_PLL1_REG_RESCAL_ONCHIP_SMALL_OW),  
    .CP_PMA_PLL1_REG_RESCAL_ONCHIP_SMALL         (PMA_PLL1_REG_RESCAL_ONCHIP_SMALL),      
    .CP_PMA_PLL1_REG_JTAG_OE                     (PMA_PLL1_REG_JTAG_OE),                  
    .CP_PMA_PLL1_REG_JTAG_AC_MODE                (PMA_PLL1_REG_JTAG_AC_MODE),             
    .CP_PMA_PLL1_REG_JTAG_VHYSTSEL               (PMA_PLL1_REG_JTAG_VHYSTSEL),            
    .CP_PMA_PLL1_REG_PLL_LOCKDET_EN_OW           (PMA_PLL1_REG_PLL_LOCKDET_EN_OW),        
    .CP_PMA_PLL1_REG_PLL_LOCKDET_EN              (PMA_PLL1_REG_PLL_LOCKDET_EN),           
    .CP_PMA_PLL1_REG_PLL_LOCKDET_RESET_N_OW      (PMA_PLL1_REG_PLL_LOCKDET_RESET_N_OW),   
    .CP_PMA_PLL1_REG_PLL_LOCKDET_RESET_N         (PMA_PLL1_REG_PLL_LOCKDET_RESET_N),      
    .CP_PMA_PLL1_REG_PLL_LOCKED_OW               (PMA_PLL1_REG_PLL_LOCKED_OW),            
    .CP_PMA_PLL1_REG_PLL_LOCKED                  (PMA_PLL1_REG_PLL_LOCKED),               
    .CP_PMA_PLL1_REG_PLL_LOCKED_STICKY_CLEAR     (PMA_PLL1_REG_PLL_LOCKED_STICKY_CLEAR),  
    .CP_PMA_PLL1_REG_PLL_UNLOCKED_STICKY_CLEAR   (PMA_PLL1_REG_PLL_UNLOCKED_STICKY_CLEAR),
    .CP_PMA_PLL1_REG_NOFBCLK_STICKY_CLEAR        (PMA_PLL1_REG_NOFBCLK_STICKY_CLEAR),     
    .CP_PMA_PLL1_REG_PLL_LOCKDET_REFCT           (PMA_PLL1_REG_PLL_LOCKDET_REFCT),        
    .CP_PMA_PLL1_REG_PLL_LOCKDET_FBCT            (PMA_PLL1_REG_PLL_LOCKDET_FBCT),         
    .CP_PMA_PLL1_REG_PLL_LOCKDET_LOCKCT          (PMA_PLL1_REG_PLL_LOCKDET_LOCKCT),       
    .CP_PMA_PLL1_REG_PLL_LOCKDET_ITER            (PMA_PLL1_REG_PLL_LOCKDET_ITER),         
    .CP_PMA_PLL1_REG_PLL_UNLOCKDET_ITER          (PMA_PLL1_REG_PLL_UNLOCKDET_ITER),       
    .CP_PMA_PLL1_REG_PD_VCO                      (PMA_PLL1_REG_PD_VCO),                   
    .CP_PMA_PLL1_REG_FBCLK_TEST_EN               (PMA_PLL1_REG_FBCLK_TEST_EN),            
    .CP_PMA_PLL1_REG_REFCLK_TEST_EN              (PMA_PLL1_REG_REFCLK_TEST_EN),           
    .CP_PMA_PLL1_REG_TEST_SEL                    (PMA_PLL1_REG_TEST_SEL),                 
    .CP_PMA_PLL1_REG_TEST_V_EN                   (PMA_PLL1_REG_TEST_V_EN),                
    .CP_PMA_PLL1_REG_TEST_SIG_HALF_EN            (PMA_PLL1_REG_TEST_SIG_HALF_EN),         
    .CP_PMA_PLL1_REG_TEST_FSM                    (PMA_PLL1_REG_TEST_FSM),                 
    .CP_PMA_PLL1_REG_REFCLK_OUT_PD               (PMA_PLL1_REG_REFCLK_OUT_PD),            
    .CP_PMA_PLL1_REG_BGR_STARTUP_EN              (PMA_PLL1_REG_BGR_STARTUP_EN),           
    .CP_PMA_PLL1_REG_BGR_STARTUP                 (PMA_PLL1_REG_BGR_STARTUP),              
    .CP_PMA_PLL1_REG_PD_BGR                      (PMA_PLL1_REG_PD_BGR),                   
    .CP_PMA_PLL1_REG_REFCLK_TERM_VCM_EN          (PMA_PLL1_REG_REFCLK_TERM_VCM_EN),       
    .CP_PMA_PLL1_REG_FBDIVA_5_EN                 (PMA_PLL1_REG_FBDIVA_5_EN),              
    .CP_PMA_PLL1_REG_FBDIVB                      (PMA_PLL1_REG_FBDIVB),                   
    .CP_PMA_PLL1_REG_RESET_N_PFDQP_OW            (PMA_PLL1_REG_RESET_N_PFDQP_OW),         
    .CP_PMA_PLL1_REG_RESET_N_PFDQP               (PMA_PLL1_REG_RESET_N_PFDQP),            
    .CP_PMA_PLL1_REG_QPCURRENT                   (PMA_PLL1_REG_QPCURRENT),                
    .CP_PMA_PLL1_REG_VC_FORCE_EN                 (PMA_PLL1_REG_VC_FORCE_EN),              
    .CP_PMA_PLL1_REG_VCRESET_C_RING              (PMA_PLL1_REG_VCRESET_C_RING),           
    .CP_PMA_PLL1_REG_LPF_R_C                     (PMA_PLL1_REG_LPF_R_C),                  
    .CP_PMA_PLL1_REG_LPF_TR_C                    (PMA_PLL1_REG_LPF_TR_C),                 
    .CP_PMA_PLL1_REG_PD_BIAS                     (PMA_PLL1_REG_PD_BIAS),                  
    .CP_PMA_PLL1_REG_ICTRL_PLL                   (PMA_PLL1_REG_ICTRL_PLL),                
    .CP_PMA_PLL1_REG_BIAS_QP                     (PMA_PLL1_REG_BIAS_QP),                  
    .CP_PMA_PLL1_REG_BIAS_LANE_SYNC              (PMA_PLL1_REG_BIAS_LANE_SYNC),           
    .CP_PMA_PLL1_REG_BIAS_CLKBUFS1               (PMA_PLL1_REG_BIAS_CLKBUFS1),            
    .CP_PMA_PLL1_REG_TXPCLK_SEL                  (PMA_PLL1_REG_TXPCLK_SEL),               
    .CP_PMA_PLL1_REG_BIAS_CLKBUFS3               (PMA_PLL1_REG_BIAS_CLKBUFS3),            
    .CP_PMA_PLL1_REG_LANE_SYNC_EN                (PMA_PLL1_REG_LANE_SYNC_EN),             
    .CP_PMA_PLL1_REG_LANE_SYNC_EN_OW             (PMA_PLL1_REG_LANE_SYNC_EN_OW),          
    .CP_PMA_PLL1_REG_BIAS_D2S                    (PMA_PLL1_REG_BIAS_D2S),                 
    .CP_PMA_PLL1_REG_BIAS_REFD2S_C               (PMA_PLL1_REG_BIAS_REFD2S_C),            
    .CP_PMA_PLL1_REG_BIAS_VCRST_C                (PMA_PLL1_REG_BIAS_VCRST_C),             
    .CP_PMA_PLL1_REG_BIAS_REFBUF_C               (PMA_PLL1_REG_BIAS_REFBUF_C),            
    .CP_PMA_PLL1_REG_CLKBUFS1_C                  (PMA_PLL1_REG_CLKBUFS1_C),               
    .CP_PMA_PLL1_REG_CLKBUFS2_C                  (PMA_PLL1_REG_CLKBUFS2_C),               
    .CP_PMA_PLL1_REG_CLKBUFS3_C                  (PMA_PLL1_REG_CLKBUFS3_C),               
    .CP_PMA_PLL1_REG_CLKBUFS4_C                  (PMA_PLL1_REG_CLKBUFS4_C),               
    .CP_PMA_PLL1_REG_PLL_REFCLK_CML_SEL          (PMA_PLL1_REG_PLL_REFCLK_CML_SEL),       
    .CP_PMA_PLL1_REG_REFCLK_SEL                  (PMA_PLL1_REG_REFCLK_SEL),               
    .CP_PMA_PLL1_REG_RESCAL_R_CODE_SIGN          (PMA_PLL1_REG_RESCAL_R_CODE_SIGN),       
    .CP_PMA_PLL1_REG_PLL_UNLOCKED_OW             (PMA_PLL1_REG_PLL_UNLOCKED_OW),          
    .CP_PMA_PLL1_REG_PLL_UNLOCKED                (PMA_PLL1_REG_PLL_UNLOCKED),             
    .CP_PMA_PLL1_REG_PLL_LOCKDET_MODE            (PMA_PLL1_REG_PLL_LOCKDET_MODE),         
    .CP_PMA_PLL1_REG_PLL_CLKBUF_PD_LEFT          (PMA_PLL1_REG_PLL_CLKBUF_PD_LEFT),       
    .CP_PMA_PLL1_REG_PLL_CLKBUF_PD_RIGHT         (PMA_PLL1_REG_PLL_CLKBUF_PD_RIGHT),      
    .CP_PMA_PLL1_REG_RESCAL_EN                   (PMA_PLL1_REG_RESCAL_EN),                
    .CP_PMA_PLL1_REG_RESCAL_I_CODE_VAL           (PMA_PLL1_REG_RESCAL_I_CODE_VAL),        
    .CP_PMA_PLL1_REG_RESCAL_I_CODE_OW            (PMA_PLL1_REG_RESCAL_I_CODE_OW),         
    .CP_PMA_PLL1_REG_RESCAL_ITER_VALID_SEL       (PMA_PLL1_REG_RESCAL_ITER_VALID_SEL),    
    .CP_PMA_PLL1_REG_RESCAL_WAIT_SEL             (PMA_PLL1_REG_RESCAL_WAIT_SEL),          
    .CP_PMA_PLL1_REG_I_CTRL_MAX                  (PMA_PLL1_REG_I_CTRL_MAX),               
    .CP_PMA_PLL1_REG_I_CTRL_MIN                  (PMA_PLL1_REG_I_CTRL_MIN),               
    .CP_PARM_PLL1_POWERUP                        (PARM_PLL1_POWERUP),                     
    .CP_PARM_PLL1_RSTN                           (PARM_PLL1_RSTN),                        
    .CP_PARM_GRSN_DIS                            (PARM_GRSN_DIS),                         
    .CP_PARM_CFG_RSTN                            (PARM_CFG_RSTN)                         
)  
gtp_hsst_wrap
(
    .PAD_REFCLKP_0                      (P_REFCLKP_0), 
    .PAD_REFCLKN_0                      (P_REFCLKN_0), 
    .PAD_PLL_TEST_0                     (P_PLL_TEST_0),
    .PAD_REFCLKP_1                      (P_REFCLKP_1),        
    .PAD_REFCLKN_1                      (P_REFCLKN_1),             
    .PAD_PLL_TEST_1                     (P_PLL_TEST_1),
    .PAD_RX_SDP0                        (P_RX_SDP0),        
    .PAD_RX_SDN0                        (P_RX_SDN0),           
    .PAD_TX_SDP0                        (P_TX_SDP0),   
    .PAD_TX_SDN0                        (P_TX_SDN0),   
    .PAD_RX_SDP1                        (P_RX_SDP1),                                   
    .PAD_RX_SDN1                        (P_RX_SDN1),           
    .PAD_TX_SDP1                        (P_TX_SDP1),   
    .PAD_TX_SDN1                        (P_TX_SDN1),           
    .PAD_RX_SDP2                        (P_RX_SDP2),                                   
    .PAD_RX_SDN2                        (P_RX_SDN2),           
    .PAD_TX_SDP2                        (P_TX_SDP2),   
    .PAD_TX_SDN2                        (P_TX_SDN2),     
    .PAD_RX_SDP3                        (P_RX_SDP3),                                   
    .PAD_RX_SDN3                        (P_RX_SDN3),           
    .PAD_TX_SDP3                        (P_TX_SDP3),   
    .PAD_TX_SDN3                        (P_TX_SDN3),     
    .RX0_CLK_FR_CORE                    (P_RX0_CLK_FR_CORE),       
    .RX1_CLK_FR_CORE                    (P_RX1_CLK_FR_CORE),         
    .RX2_CLK_FR_CORE                    (P_RX2_CLK_FR_CORE),         
    .RX3_CLK_FR_CORE                    (P_RX3_CLK_FR_CORE),         
    .TX0_CLK_FR_CORE                    (P_TX0_CLK_FR_CORE),       
    .TX1_CLK_FR_CORE                    (P_TX1_CLK_FR_CORE),         
    .TX2_CLK_FR_CORE                    (P_TX2_CLK_FR_CORE),         
    .TX3_CLK_FR_CORE                    (P_TX3_CLK_FR_CORE), 
    .HSST_RST                           (P_HSST_RST),
    .PCS_RX_RST_0                       (P_PCS_RX_RST_0),
    .PCS_RX_RST_1                       (P_PCS_RX_RST_1),        
    .PCS_RX_RST_2                       (P_PCS_RX_RST_2),
    .PCS_RX_RST_3                       (P_PCS_RX_RST_3),        
    .PCS_TX_RST_0                       (P_PCS_TX_RST_0),
    .PCS_TX_RST_1                       (P_PCS_TX_RST_1),        
    .PCS_TX_RST_2                       (P_PCS_TX_RST_2),        
    .PCS_TX_RST_3                       (P_PCS_TX_RST_3),
    .CFG_CLK                            (P_CFG_CLK),   
    .CFG_RST                            (P_CFG_RST),   
    .CFG_ENABLE                         (P_CFG_ENABLE),
    .CFG_WRITE                          (P_CFG_WRITE), 
    .CFG_ADDR                           (P_CFG_ADDR),  
    .CFG_WDATA                          (P_CFG_WDATA), 
    .TDATA_0                            (P_TDATA_0),
    .TDATA_1                            (P_TDATA_1),
    .TDATA_2                            (P_TDATA_2),
    .TDATA_3                            (P_TDATA_3),
    .PCS_WORD_ALIGN_EN                  (P_PCS_WORD_ALIGN_EN), 
    .RX_POLARITY_INVERT                 (P_RX_POLARITY_INVERT),
    .CEB_ADETECT_EN                     (P_CEB_ADETECT_EN),    
    .PCS_MCB_EXT_EN                     (P_PCS_MCB_EXT_EN),    
    .PCS_NEAREND_LOOP                   (P_PCS_NEAREND_LOOP),  
    .PCS_FAREND_LOOP                    (P_PCS_FAREND_LOOP),   
    .CFG_READY                          (P_CFG_READY),         
    .CFG_RDATA                          (P_CFG_RDATA),         
    .CFG_INT                            (P_CFG_INT),           
    .PCS_RX_MCB_STATUS                  (P_PCS_RX_MCB_STATUS), 
    .PCS_LSM_SYNCED                     (P_PCS_LSM_SYNCED),    
    .RDATA_0                            (P_RDATA_0),
    .RDATA_1                            (P_RDATA_1),
    .RDATA_2                            (P_RDATA_2),
    .RDATA_3                            (P_RDATA_3),
    .RCLK2FABRIC                        (P_RCLK2FABRIC),    
    .TCLK2FABRIC                        (P_TCLK2FABRIC),    
    .RESCAL_RST_I                       (P_RESCAL_RST_I),          
    .RESCAL_I_CODE_I                    (P_RESCAL_I_CODE_I),   
    .RESCAL_I_CODE_O                    (P_RESCAL_I_CODE_O),
    .REFCK2CORE_0                       (P_REFCK2CORE_0),         
    .PLL_REF_CLK_0                      (P_PLL_REF_CLK_0),        
    .PLL_RST_0                          (P_PLL_RST_0), 
    .PLLPOWERDOWN_0                     (P_PLLPOWERDOWN_0),
    .PLL_READY_0                        (P_PLL_READY_0),          
    .LANE_SYNC_0                        (P_LANE_SYNC_0),          
    .LANE_SYNC_EN_0                     (P_LANE_SYNC_EN_0),       
    .RATE_CHANGE_TCLK_ON_0              (P_RATE_CHANGE_TCLK_ON_0),
    .REFCK2CORE_1                       (P_REFCK2CORE_1),         
    .PLL_REF_CLK_1                      (P_PLL_REF_CLK_1),        
    .PLL_RST_1                          (P_PLL_RST_1),            
    .PLLPOWERDOWN_1                     (P_PLLPOWERDOWN_1),       
    .PLL_READY_1                        (P_PLL_READY_1),          
    .LANE_SYNC_1                        (P_LANE_SYNC_1),          
    .LANE_SYNC_EN_1                     (P_LANE_SYNC_EN_1),       
    .RATE_CHANGE_TCLK_ON_1              (P_RATE_CHANGE_TCLK_ON_1),
    .LANE_PD_0                          (P_LANE_PD_0),         
    .LANE_RST_0                         (P_LANE_RST_0),        
    .RX_LANE_PD_0                       (P_RX_LANE_PD_0),      
    .RX_PMA_RST_0                       (P_RX_PMA_RST_0),      
    .RX_SIGDET_STATUS_0                 (P_RX_SIGDET_STATUS_0),
    .RX_SATA_COMINIT_0                  (P_RX_SATA_COMINIT_0), 
    .RX_SATA_COMWAKE_0                  (P_RX_SATA_COMWAKE_0), 
    .RX_LS_DATA_0                       (P_RX_LS_DATA_0),      
    .RX_READY_0                         (P_RX_READY_0),        
    .TEST_STATUS_0                      (P_TEST_STATUS_0),     
    .TX_DEEMP_0                         (P_TX_DEEMP_0),        
    .TX_LS_DATA_0                       (P_TX_LS_DATA_0),      
    .TX_BEACON_EN_0                     (P_TX_BEACON_EN_0),    
    .TX_SWING_0                         (P_TX_SWING_0),        
    .TX_RXDET_REQ_0                     (P_TX_RXDET_REQ_0),    
    .TX_RATE_0                          (P_TX_RATE_0),         
    .TX_BUSWIDTH_0                      (P_TX_BUSWIDTH_0),     
    .TX_MARGIN_0                        (P_TX_MARGIN_0),       
    .TX_RXDET_STATUS_0                  (P_TX_RXDET_STATUS_0), 
    .TX_PMA_RST_0                       (P_TX_PMA_RST_0),      
    .TX_LANE_PD_0                       (P_TX_LANE_PD_0),      
    .RX_RATE_0                          (P_RX_RATE_0),         
    .RX_BUSWIDTH_0                      (P_RX_BUSWIDTH_0),     
    .RX_HIGHZ_0                         (P_RX_HIGHZ_0),        
    .CA_ALIGN_RX                        (P_CA_ALIGN_RX),       
    .CA_ALIGN_TX                        (P_CA_ALIGN_TX),       
    .CIM_CLK_ALIGNER_RX0                (P_CIM_CLK_ALIGNER_RX0),
    .CIM_CLK_ALIGNER_TX0                (P_CIM_CLK_ALIGNER_TX0),
    .CIM_DYN_DLY_SEL_RX0                (P_CIM_DYN_DLY_SEL_RX0),
    .CIM_DYN_DLY_SEL_TX0                (P_CIM_DYN_DLY_SEL_TX0),
    .CIM_START_ALIGN_RX0                (P_CIM_START_ALIGN_RX0),
    .CIM_START_ALIGN_TX0                (P_CIM_START_ALIGN_TX0),
    .LANE_PD_1                          (P_LANE_PD_1),         
    .LANE_RST_1                         (P_LANE_RST_1),        
    .RX_LANE_PD_1                       (P_RX_LANE_PD_1),      
    .RX_PMA_RST_1                       (P_RX_PMA_RST_1),      
    .RX_SIGDET_STATUS_1                 (P_RX_SIGDET_STATUS_1),
    .RX_SATA_COMINIT_1                  (P_RX_SATA_COMINIT_1), 
    .RX_SATA_COMWAKE_1                  (P_RX_SATA_COMWAKE_1), 
    .RX_LS_DATA_1                       (P_RX_LS_DATA_1),      
    .RX_READY_1                         (P_RX_READY_1),        
    .TEST_STATUS_1                      (P_TEST_STATUS_1),     
    .TX_DEEMP_1                         (P_TX_DEEMP_1),        
    .TX_LS_DATA_1                       (P_TX_LS_DATA_1),      
    .TX_BEACON_EN_1                     (P_TX_BEACON_EN_1),    
    .TX_SWING_1                         (P_TX_SWING_1),        
    .TX_RXDET_REQ_1                     (P_TX_RXDET_REQ_1),    
    .TX_RATE_1                          (P_TX_RATE_1),         
    .TX_BUSWIDTH_1                      (P_TX_BUSWIDTH_1),     
    .TX_MARGIN_1                        (P_TX_MARGIN_1),       
    .TX_RXDET_STATUS_1                  (P_TX_RXDET_STATUS_1), 
    .TX_PMA_RST_1                       (P_TX_PMA_RST_1),      
    .TX_LANE_PD_1                       (P_TX_LANE_PD_1),      
    .RX_RATE_1                          (P_RX_RATE_1),         
    .RX_BUSWIDTH_1                      (P_RX_BUSWIDTH_1),     
    .RX_HIGHZ_1                         (P_RX_HIGHZ_1),        
    .CIM_CLK_ALIGNER_RX1                (P_CIM_CLK_ALIGNER_RX1),
    .CIM_CLK_ALIGNER_TX1                (P_CIM_CLK_ALIGNER_TX1),
    .CIM_DYN_DLY_SEL_RX1                (P_CIM_DYN_DLY_SEL_RX1),
    .CIM_DYN_DLY_SEL_TX1                (P_CIM_DYN_DLY_SEL_TX1),
    .CIM_START_ALIGN_RX1                (P_CIM_START_ALIGN_RX1),
    .CIM_START_ALIGN_TX1                (P_CIM_START_ALIGN_TX1),
    .LANE_PD_2                          (P_LANE_PD_2),         
    .LANE_RST_2                         (P_LANE_RST_2),        
    .RX_LANE_PD_2                       (P_RX_LANE_PD_2),      
    .RX_PMA_RST_2                       (P_RX_PMA_RST_2),      
    .RX_SIGDET_STATUS_2                 (P_RX_SIGDET_STATUS_2),
    .RX_SATA_COMINIT_2                  (P_RX_SATA_COMINIT_2), 
    .RX_SATA_COMWAKE_2                  (P_RX_SATA_COMWAKE_2), 
    .RX_LS_DATA_2                       (P_RX_LS_DATA_2),      
    .RX_READY_2                         (P_RX_READY_2),        
    .TEST_STATUS_2                      (P_TEST_STATUS_2),     
    .TX_DEEMP_2                         (P_TX_DEEMP_2),        
    .TX_LS_DATA_2                       (P_TX_LS_DATA_2),      
    .TX_BEACON_EN_2                     (P_TX_BEACON_EN_2),    
    .TX_SWING_2                         (P_TX_SWING_2),        
    .TX_RXDET_REQ_2                     (P_TX_RXDET_REQ_2),    
    .TX_RATE_2                          (P_TX_RATE_2),         
    .TX_BUSWIDTH_2                      (P_TX_BUSWIDTH_2),     
    .TX_MARGIN_2                        (P_TX_MARGIN_2),       
    .TX_RXDET_STATUS_2                  (P_TX_RXDET_STATUS_2), 
    .TX_PMA_RST_2                       (P_TX_PMA_RST_2),      
    .TX_LANE_PD_2                       (P_TX_LANE_PD_2),      
    .RX_RATE_2                          (P_RX_RATE_2),         
    .RX_BUSWIDTH_2                      (P_RX_BUSWIDTH_2),     
    .RX_HIGHZ_2                         (P_RX_HIGHZ_2),        
    .CIM_CLK_ALIGNER_RX2                (P_CIM_CLK_ALIGNER_RX2),
    .CIM_CLK_ALIGNER_TX2                (P_CIM_CLK_ALIGNER_TX2),
    .CIM_DYN_DLY_SEL_RX2                (P_CIM_DYN_DLY_SEL_RX2),
    .CIM_DYN_DLY_SEL_TX2                (P_CIM_DYN_DLY_SEL_TX2),
    .CIM_START_ALIGN_RX2                (P_CIM_START_ALIGN_RX2),
    .CIM_START_ALIGN_TX2                (P_CIM_START_ALIGN_TX2),
    .LANE_PD_3                          (P_LANE_PD_3),         
    .LANE_RST_3                         (P_LANE_RST_3),        
    .RX_LANE_PD_3                       (P_RX_LANE_PD_3),      
    .RX_PMA_RST_3                       (P_RX_PMA_RST_3),      
    .RX_SIGDET_STATUS_3                 (P_RX_SIGDET_STATUS_3),
    .RX_SATA_COMINIT_3                  (P_RX_SATA_COMINIT_3), 
    .RX_SATA_COMWAKE_3                  (P_RX_SATA_COMWAKE_3), 
    .RX_LS_DATA_3                       (P_RX_LS_DATA_3),      
    .RX_READY_3                         (P_RX_READY_3),        
    .TEST_STATUS_3                      (P_TEST_STATUS_3),     
    .TX_DEEMP_3                         (P_TX_DEEMP_3),        
    .TX_LS_DATA_3                       (P_TX_LS_DATA_3),      
    .TX_BEACON_EN_3                     (P_TX_BEACON_EN_3),    
    .TX_SWING_3                         (P_TX_SWING_3),        
    .TX_RXDET_REQ_3                     (P_TX_RXDET_REQ_3),    
    .TX_RATE_3                          (P_TX_RATE_3),         
    .TX_BUSWIDTH_3                      (P_TX_BUSWIDTH_3),     
    .TX_MARGIN_3                        (P_TX_MARGIN_3),       
    .TX_RXDET_STATUS_3                  (P_TX_RXDET_STATUS_3), 
    .TX_PMA_RST_3                       (P_TX_PMA_RST_3),      
    .TX_LANE_PD_3                       (P_TX_LANE_PD_3),      
    .RX_RATE_3                          (P_RX_RATE_3),         
    .RX_BUSWIDTH_3                      (P_RX_BUSWIDTH_3),     
    .RX_HIGHZ_3                         (P_RX_HIGHZ_3),        
    .CIM_CLK_ALIGNER_RX3                (P_CIM_CLK_ALIGNER_RX3),
    .CIM_CLK_ALIGNER_TX3                (P_CIM_CLK_ALIGNER_TX3),
    .CIM_DYN_DLY_SEL_RX3                (P_CIM_DYN_DLY_SEL_RX3),
    .CIM_DYN_DLY_SEL_TX3                (P_CIM_DYN_DLY_SEL_TX3),
    .CIM_START_ALIGN_RX3                (P_CIM_START_ALIGN_RX3),
    .CIM_START_ALIGN_TX3                (P_CIM_START_ALIGN_TX3),
    .TEST_SI0                           (),
    .TEST_SI1                           (),
    .TEST_SI2                           (),
    .TEST_SI3                           (),
    .TEST_SI4                           (),
    .TEST_SI5                           (),
    .TEST_SI6                           (),
    .TEST_SI7                           (),
    .TEST_SE_N                          (),
    .TEST_MODE_N                        (1'b1),
    .TEST_CLK                           (),
    .TEST_RSTN                          (1'b1),
    .COMPRESSION_MODE                   (),
    .PLL_BYPASS                         (),
    .PLL_RESET                          (),
    .TEST_SO0                           (),
    .TEST_SO1                           (),
    .TEST_SO2                           (),
    .TEST_SO3                           (),
    .TEST_SO4                           (),
    .TEST_SO5                           (),
    .TEST_SO6                           (),
    .TEST_SO7                           ()
);

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_SCANCHAIN.v
//
// Functional description: JTAG TAP Controller simulation model
//
// Parameter description:
//      
//
// Port description:
//      
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale  1 ns / 1 ps

module GTP_SCANCHAIN
#(
    parameter [31:0] IDCODE = 32'haaaa5555, //dr idcode
    parameter   CHAIN_NUM = 1 //1 2 3 4 available
)
(
    input      TCK      ,//JTAG signals
    input      TDI      ,
    input      TMS      ,
    output reg TDO      ,
    
    output reg CAPDR    ,//scanchain signals
    output     JCLK     ,
    output reg RST      ,
    output reg FLG_USER ,
    output reg SHFTDR   ,
    output     TDI_USER ,
    output reg UPDR     ,
    input      TDO_USER 
);

wire           flg_capture_ir  ;
wire           flg_shift_ir    ;
wire           flg_update_ir   ;
wire           flg_capture_dr  ;
wire           flg_shift_dr    ;
wire           flg_update_dr   ;
wire           flg_idcode      ;
wire           flg_bypass      ;
wire           flg_bypass_highz;

wire           irq             ;
wire           drq_bypass      ;
wire           drq_idcode      ;
wire	       flg_user        ;

reg    [3:0]   s               ;
reg    [3:0]   ns              ;

reg            flg_jclk        ;
reg    [9:0]   USER	       ;
reg    [9:0]   shift_ir        ;
reg    [9:0]   update          ;

wire           flg_highz       ;


//////////JTAG signals///////////
reg            JTAG_USER = 1'bz;

localparam TEST_LOGIC_RESET  =  4'd0 ,
           RUN_TEST_IDLE     =  4'd1 ,
           SELECT_IR_SCAN    =  4'd2 ,
           CAPTURE_IR        =  4'd3 ,
           SHIFT_IR          =  4'd4 ,
           EXIT1_IR          =  4'd5 ,
           PAUSE_IR          =  4'd6 ,
           EXIT2_IR          =  4'd7 ,
           UPDATE_IR         =  4'd8 ,
           SELECT_DR_SCAN    =  4'd9 ,
           CAPTURE_DR        =  4'd10,
           SHIFT_DR          =  4'd11,
           EXIT1_DR          =  4'd12,
           PAUSE_DR          =  4'd13,
           EXIT2_DR          =  4'd14,
           UPDATE_DR         =  4'd15;

localparam USER1                =  10'b10_1000_0110, // Access user-defined register 1
           USER2                =  10'b10_1000_0111, // Access user-defined register 2
           USER3                =  10'b10_1000_1000, // Access user-defined register 3
           USER4                =  10'b10_1000_1001, // Access user-defined register 4
           ID_CODE               =  10'b10_1000_0011, // Enables shifting out of ID code
           HIGHZ                =  10'b10_1000_0101, // 3-state output pins while enabling
           BYPASS               =  10'b11_1111_1111; // Enables BYPASS


                    
initial 
     begin
       case (CHAIN_NUM)
           1: USER <= USER1;
           2: USER <= USER2;
           3: USER <= USER3;
           4: USER <= USER4;
     default: 
            $display("Error: CHAIN_NUM is not available");
endcase
end
           


/*always @(posedge TCK)
       begin
          scanchain <= SCANCHAIN;
end
*/
always @(posedge TCK)
    begin
        s <= ns;
    end

always @(*)
    begin
        case(s)
            TEST_LOGIC_RESET:
                begin
                    if(TMS)
                        ns = TEST_LOGIC_RESET;
                    else
                        ns = RUN_TEST_IDLE;
                end

            RUN_TEST_IDLE:
                begin
                    if(TMS)
                        ns = SELECT_DR_SCAN;
                    else
                        ns = RUN_TEST_IDLE;
                end

            SELECT_IR_SCAN:
                begin
                    if(TMS)
                        ns = TEST_LOGIC_RESET;
                    else
                        ns = CAPTURE_IR;
                end

            CAPTURE_IR, SHIFT_IR:
                begin
                    if(TMS)
                        ns = EXIT1_IR;
                    else
                        ns = SHIFT_IR;
                end
            
            EXIT1_IR:
                begin
                    if(TMS)
                        ns = UPDATE_IR;
                    else
                        ns = PAUSE_IR;
                end

            PAUSE_IR:
                begin
                    if(TMS)
                        ns = EXIT2_IR;
                    else
                        ns = PAUSE_IR;
                end

            EXIT2_IR:
                begin
                    if(TMS)
                        ns = UPDATE_IR;
                    else
                        ns = SHIFT_IR;
                end

            UPDATE_IR, UPDATE_DR:
                begin
                    if(TMS)
                        ns = SELECT_DR_SCAN;
                    else
                        ns = RUN_TEST_IDLE;
                end

            SELECT_DR_SCAN:
                begin
                    if(TMS)
                        ns = SELECT_IR_SCAN;
                    else
                        ns = CAPTURE_DR;
                end

            CAPTURE_DR, SHIFT_DR:
                begin
                    if(TMS)
                        ns = EXIT1_DR;
                    else
                        ns = SHIFT_DR;
                end

            EXIT1_DR:
                begin
                    if(TMS)
                        ns = UPDATE_DR;
                    else
                        ns = PAUSE_DR;
                end

            PAUSE_DR:
                begin
                    if(TMS)
                        ns = EXIT2_DR;
                    else
                        ns = PAUSE_DR;
                end

            EXIT2_DR:
                begin
                    if(TMS)
                        ns = UPDATE_DR;
                    else
                        ns = SHIFT_DR;
                end
        default: 
               ns = TEST_LOGIC_RESET;
        endcase
    end

always @(negedge TCK)
    begin
        if(s == TEST_LOGIC_RESET)
            RST <= 1'b1;
        else
            RST <= 1'b0;
    end
       
assign flg_capture_ir = (s == CAPTURE_IR);
assign flg_shift_ir   = (s == SHIFT_IR  );
assign flg_update_ir  = (s == UPDATE_IR );
assign flg_capture_dr = (s == CAPTURE_DR);
assign flg_shift_dr   = (s == SHIFT_DR  );
assign flg_update_dr  = (s == UPDATE_DR );

/*always@(negedge RST)
    begin

     case (scanchain)
        3'd1:
    	    USER = USER1;
        3'd2:
            USER = USER2;
        3'd3:
            USER = USER3;
        3'd4:
            USER = USER4; 
       default:
            $display("Error: SCANCHAIN mismatched");

endcase
end
*/
always @(posedge TCK)
    begin
        if(RST)
            shift_ir <= 10'd0;
        else if(flg_capture_ir)
            shift_ir <= 10'd0;
        else if(flg_shift_ir)
            shift_ir <= {TDI, shift_ir[9:1]};
    end

assign irq = shift_ir[0];

always @(negedge TCK)
    begin
        if(RST)
            update <= ID_CODE;//ir idcode
        else if(flg_update_ir)
            update <= shift_ir;
    end

assign flg_user                 =  (update == USER );
assign flg_idcode               =  (update == ID_CODE);
assign flg_bypass               =  (update == BYPASS);
assign flg_highz                =  (update == HIGHZ );
assign flg_bypass_highz         =  flg_bypass | flg_highz;

reg    shift_bypass;
assign drq_bypass = shift_bypass;

always @(posedge TCK)
    begin
        if(RST)
            shift_bypass <= 1'b0;
        else if(flg_bypass_highz)
            begin
                if(flg_capture_dr)
                    shift_bypass <= 1'b0;
                else if(flg_shift_dr)
                    shift_bypass <= TDI;
            end
    end


reg    [31:0]    shift_id;
assign drq_idcode = shift_id[0];

always @(posedge TCK)
    begin
        if(RST)
            shift_id <= 32'd0;
        else if(flg_idcode)
            begin
                if(flg_capture_dr)
                    shift_id <= IDCODE;//dr idcode
                else if(flg_shift_dr)
                    shift_id <= {TDI, shift_id[31:1]};
                else
                    shift_id <= 32'd0;
            end
        else
            shift_id <= 32'd0;
    end


always @(negedge TCK)
    begin
        if(RST)
            begin
                CAPDR  <= 1'b0;
                SHFTDR <= 1'b0;
                UPDR   <= 1'b0;
            end
        else
            begin
                CAPDR  <= flg_capture_dr;
                SHFTDR <= flg_shift_dr  ;
                UPDR   <= flg_update_dr ;
            end
    end

always @(negedge TCK)
    begin
        if(RST)
            flg_jclk <= 1'b0;
        else if(CAPDR)
            flg_jclk <= 1'b1;
        else if(UPDR)
            flg_jclk <= 1'b0;
    end

assign JCLK = flg_user & (CAPDR | flg_jclk) & TCK;

always @(negedge TCK)
    begin
        if(RST)
            TDO <= 1'b0;
        else if(flg_shift_ir)
            TDO <= irq;
        else if(flg_shift_dr)
            case({flg_bypass_highz, flg_idcode, flg_user})
                3'b10_0: TDO <= drq_bypass;
                3'b01_0: TDO <= drq_idcode;
                3'b00_1: TDO <= TDO_USER;
                default: TDO <= 1'b0;
            endcase
    end
always@(*)

	begin 
		FLG_USER <= flg_user;
	end
////////////////////user tdo//////////
always@(*)
	begin
		JTAG_USER <= TDO_USER;
end
assign TDI_USER = TDI;

endmodule









//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_I2C.v
//
// Functional description: I2C Circuit
//
// Parameter description:
//      
//
// Port description:
//      
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////


`timescale 1 ns / 1 ps
module GTP_I2C
#(
    parameter   I2C_NUM = 0 //0 1 available
)
(
input         SCL_I,
output        SCL_O,
input         SDA_I,
output        SDA_O,
output        IRQ
);

assign  GTP_GRS.i2c0_scl_i = (I2C_NUM == 0) ? SCL_I : 1'bz;
assign  GTP_GRS.i2c0_sda_i = (I2C_NUM == 0) ? SDA_I : 1'bz;
assign  GTP_GRS.i2c1_scl_i = (I2C_NUM == 1) ? SCL_I : 1'bz;
assign  GTP_GRS.i2c1_sda_i = (I2C_NUM == 1) ? SDA_I : 1'bz;
assign  SCL_O = (I2C_NUM == 0) ? GTP_GRS.i2c0_scl_o : ((I2C_NUM == 1) ? GTP_GRS.i2c1_scl_o : 1'bz);
assign  SDA_O = (I2C_NUM == 0) ? GTP_GRS.i2c0_sda_o : ((I2C_NUM == 1) ? GTP_GRS.i2c1_sda_o : 1'bz);
assign  IRQ   = (I2C_NUM == 0) ? GTP_GRS.irq_i2c0   : ((I2C_NUM == 1) ? GTP_GRS.irq_i2c1   : 1'bz);

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2016 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_LUT6D.v
//
// Functional description: 6-input Look-Up-Table with double output
//
// Parameter description:
//      INIT: init value
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_LUT6D
#(
    parameter [63:0] INIT = 64'h0000_0000_0000_0000
) (
    output wire Z, Z5,
    input wire I0, I1, I2, I3, I4, I5
);

    wire z5a, z5b;

    GTP_LUT5 #(.INIT(INIT[31:0]))
        l5a (.I0(I0), .I1(I1), .I2(I2), .I3(I3), .I4(I4), .Z(z5a));

    GTP_LUT5 #(.INIT(INIT[63:32]))
        l5b (.I0(I0), .I1(I1), .I2(I2), .I3(I3), .I4(I4), .Z(z5b));

    GTP_MUX2LUT6 mxl6 (.I0(z5a), .I1(z5b), .S(I5), .Z(Z));
    buf (Z5, z5a);

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_DRM9K.v
//
// Functional description:
//
// Parameter  description:
//
// Port description:
//
// Revision history:
//   2017/05/23: Copy from GTP_DRM9K, Remve WW conflict feature, Size change
//               to be 9K.
//   2018/01/09: Update display informations.
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_DRM9K
#(
    parameter GRS_EN = "TRUE",
    //parameter [2:0] CSA_MASK = 3'b000,
    //parameter [2:0] CSB_MASK = 3'b000,
    parameter integer DATA_WIDTH_A = 18,
    parameter integer DATA_WIDTH_B = 18,
    parameter WRITE_MODE_A = "NORMAL_WRITE",
    parameter WRITE_MODE_B = "NORMAL_WRITE",
    parameter integer DOA_REG = 0,
    parameter integer DOB_REG = 0,
    parameter integer DOA_REG_CLKINV = 0,
    parameter integer DOB_REG_CLKINV = 0,
    parameter RST_TYPE = "SYNC",
    parameter RAM_MODE = "TRUE_DUAL_PORT",
    parameter SIM_DEVICE = "LOGOS",
    parameter [287:0] INIT_00 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_01 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_02 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_03 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_04 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_05 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_06 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_07 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_08 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_09 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_10 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_11 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_12 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_13 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_14 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_15 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_16 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_17 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_18 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_19 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_FILE = "NONE",
    parameter integer BLOCK_X = 0,
    parameter integer BLOCK_Y = 0,
    parameter integer RAM_DATA_WIDTH = 9,
    parameter integer RAM_ADDR_WIDTH = 10,
    parameter INIT_FORMAT = "BIN"
) (
    output [17:0] DOA,
    output [17:0] DOB,
    input [17:0] DIA,
    input [17:0] DIB,
    input [12:0] ADDRA,
    input ADDRA_HOLD,
    input [12:0] ADDRB,
    input ADDRB_HOLD,
    //input [2:0] CSA,
    //input [2:0] CSB,
    input CLKA,
    input CLKB,
    input CEA,
    input CEB,
    input WEA,
    input WEB,
    input ORCEA,
    input ORCEB,
    input RSTA,
    input RSTB
);

    localparam  BLOCK_DEPTH = 2**(DATA_WIDTH_A == 1 ? 13 :    // block type 8k*1
                                  DATA_WIDTH_A == 2 ? 12 :    // block type 4k*2
                                  DATA_WIDTH_A == 4 ? 11 :    // block type 2k*4
                                  DATA_WIDTH_A <= 9 ? 10 :    // block type 1k*8 or 1k*9
                                 DATA_WIDTH_A <= 18 ? 9 : 8); // block type 256*36 or 256*32     block memory address width

    localparam  BLOCK_WIDTH =   DATA_WIDTH_A;             //block memory data width
//end add for initialization

    localparam MEM_SIZE = 9216;
    localparam width_a = (DATA_WIDTH_A == 32) ? 16 : (DATA_WIDTH_A == 36) ? 18 : DATA_WIDTH_A;
    localparam width_b = (DATA_WIDTH_B == 32) ? 16 : (DATA_WIDTH_B == 36) ? 18 : DATA_WIDTH_B;

    integer  cnt;
    reg [9-1:0] mem [MEM_SIZE/9-1:0];

    //reg [2:0] csa_reg = 3'b0, csb_reg = 3'b0;
    reg [12:0] ada_reg = 13'b0, adb_reg = 13'b0;
    reg [17:0] da_reg = 18'b0, db_reg = 18'b0;
    reg wea_reg = 1'b0, web_reg = 1'b0;
    wire [3:0] bea_reg;   // modify for byte_write_enable bug
    wire [1:0] beb_reg;
    wire write_en_a, write_en_b, read_en_a, read_en_b;

    reg [17:0] a_out = 18'b0, a_out_reg = 18'b0;
    //reg [17:0] a_out_reg_sync = 18'b0, a_out_reg_async = 18'b0, a_out_reg_async_sy = 18'b0;
    reg [17:0] b_out = 18'b0, b_out_reg = 18'b0;
    //reg [17:0] b_out_reg_sync = 18'b0, b_out_reg_async = 18'b0, b_out_reg_async_sy = 18'b0;

    wire grs, rsta_grs, rstb_grs;
    reg rsta_async_sy = 1'b0, rstb_async_sy = 1'b0;
    wire rsta_grs_sync;
    wire rstb_grs_sync;
    wire rsta_grs_async;
    wire rstb_grs_async;
    wire rsta_async_synrel;
    wire rstb_async_synrel;
    wire rsta_int;
    wire rstb_int;
    
    reg [17:0] doa;
    reg [17:0] dob;

    initial begin
        doa = 0;
        dob = 0;
    end

// synthesis translate_off
// add for memory initialization 2014/7/2 10:59:37    1) add ini_mem reg array to load init.dat
//                                                    2) init_file contain all the initial data of cascaded DRMS
   reg [RAM_DATA_WIDTH-1:0] ini_mem [2**RAM_ADDR_WIDTH-1:0];
   integer p;
   initial
   begin
      if(INIT_FILE != "NONE")
      begin
          if(INIT_FORMAT == "BIN")
              $readmemb(INIT_FILE,ini_mem);
          else
              $readmemh(INIT_FILE,ini_mem);
          for(p=0;p<20;p=p+1)
              $display("ini_mem[%d] = %b",p,ini_mem[p]);
      end
   end
//end  add
///////////////////
// parameter check
///////////////////
    initial begin
        case (DATA_WIDTH_A)
            1, 2, 4, 8, 16, 32: begin
                case (DATA_WIDTH_B)
                    1, 2, 4, 8, 16, 32:  ; //null
                    default: begin
                        $display("ERROR: GTP_DRM9K instance %m parameter DATA_WIDTH_B:%d is illegal. The legal values are 1,2,4,8,16 or 32.",DATA_WIDTH_B);
                        $finish;
                    end
                endcase
            end
            9, 18, 36: begin
                case (DATA_WIDTH_B)
                    9, 18, 36:    ; //null
                    default: begin
                        $display("ERROR: GTP_DRM9K instance %m parameter DATA_WIDTH_B:%d is illegal. The legal values are 9,18 or 36.",DATA_WIDTH_B);
                        $finish;
                    end
                endcase
            end
            default: begin
                $display("ERROR: GTP_DRM9K instance %m parameter DATA_WIDTH_A:%d is illegal. The legal values are 1,2,4,8,9,16,18,32 or 36.",DATA_WIDTH_A);
                $finish;
            end
        endcase

        case (WRITE_MODE_A)
            "NORMAL_WRITE",
            "TRANSPARENT_WRITE",
            "READ_BEFORE_WRITE":    ; //null 
            default: begin
                $display("ERROR: GTP_DRM9K instance %m parameter WRITE_MODE_A: %s is illegal. The legal values are NORMAL_WRITE,TRANSPARENT_WRITE or READ_BEFORE_WRITE.", WRITE_MODE_A);
                $finish;
            end
        endcase

        case (WRITE_MODE_B)
            "NORMAL_WRITE",
            "TRANSPARENT_WRITE",
            "READ_BEFORE_WRITE":    ; //null  
            default: begin
                $display("ERROR: GTP_DRM9K instance %m parameter WRITE_MODE_B: %s is illegal. The legal values are NORMAL_WRITE,TRANSPARENT_WRITE or READ_BEFORE_WRITE.", WRITE_MODE_B);
                $finish;
            end
        endcase

        case (RST_TYPE)
            "ASYNC",
            "ASYNC_SYNC_RELEASE",
            "SYNC":     ;//null
            default: begin
                $display("ERROR: GTP_DRM9K instance %m parameter RST_TYPE: %s is illegal. The legal values are ASYNC,ASYNC_SYNC_RELEASE or SYNC.", RST_TYPE);
                $finish;
            end
        endcase

        case (RAM_MODE)
            "ROM",
            "SINGLE_PORT","SIMPLE_DUAL_PORT":     ;//null
            "TRUE_DUAL_PORT": begin
                if (DATA_WIDTH_A > 18 || DATA_WIDTH_B > 18) begin
                    $display("ERROR: GTP_DRM9K instance %m parameter DATA_WIDTH_A and DATA_WIDTH_B in TRUE_DUAL_PORT MODE:%d,%d is illegal. The legal values are 1,2,4,8,9,16 or 18.",DATA_WIDTH_A,DATA_WIDTH_B);
                    $finish;
                end
            end
            default: begin
                $display("ERROR: GTP_DRM9K instance %m parameter RAM_MODE value: %s is illegal. The legal values are ROM or SINGLE_PORT or SIMPLE_DUAL_PORT or TRUE_DUAL_PORT.", RAM_MODE);
                $finish;
            end
        endcase

        case (SIM_DEVICE)
            "LOGOS","PGL22G":    ;//null
            default: begin
                   $display("ERROR: GTP_DRM9K instance %m parameter SIM_DEVICE value: %s is illegal. The legal values are LOGOS or PGL22G.", SIM_DEVICE);
                   $finish;
            end
        endcase

    end

/////////////////=
// initialization
/////////////////=

    initial begin
        if (INIT_FILE == "NONE") begin
            for (cnt = 0; cnt < 32; cnt = cnt + 1) begin
                mem[32*0 + cnt] = INIT_00[cnt*9 +: 9];
                mem[32*1 + cnt] = INIT_01[cnt*9 +: 9];
                mem[32*2 + cnt] = INIT_02[cnt*9 +: 9];
                mem[32*3 + cnt] = INIT_03[cnt*9 +: 9];
                mem[32*4 + cnt] = INIT_04[cnt*9 +: 9];
                mem[32*5 + cnt] = INIT_05[cnt*9 +: 9];
                mem[32*6 + cnt] = INIT_06[cnt*9 +: 9];
                mem[32*7 + cnt] = INIT_07[cnt*9 +: 9];
                mem[32*8 + cnt] = INIT_08[cnt*9 +: 9];
                mem[32*9 + cnt] = INIT_09[cnt*9 +: 9];
                mem[32*10 + cnt] = INIT_0A[cnt*9 +: 9];
                mem[32*11 + cnt] = INIT_0B[cnt*9 +: 9];
                mem[32*12 + cnt] = INIT_0C[cnt*9 +: 9];
                mem[32*13 + cnt] = INIT_0D[cnt*9 +: 9];
                mem[32*14 + cnt] = INIT_0E[cnt*9 +: 9];
                mem[32*15 + cnt] = INIT_0F[cnt*9 +: 9];
                mem[32*16 + cnt] = INIT_10[cnt*9 +: 9];
                mem[32*17 + cnt] = INIT_11[cnt*9 +: 9];
                mem[32*18 + cnt] = INIT_12[cnt*9 +: 9];
                mem[32*19 + cnt] = INIT_13[cnt*9 +: 9];
                mem[32*20 + cnt] = INIT_14[cnt*9 +: 9];
                mem[32*21 + cnt] = INIT_15[cnt*9 +: 9];
                mem[32*22 + cnt] = INIT_16[cnt*9 +: 9];
                mem[32*23 + cnt] = INIT_17[cnt*9 +: 9];
                mem[32*24 + cnt] = INIT_18[cnt*9 +: 9];
                mem[32*25 + cnt] = INIT_19[cnt*9 +: 9];
                mem[32*26 + cnt] = INIT_1A[cnt*9 +: 9];
                mem[32*27 + cnt] = INIT_1B[cnt*9 +: 9];
                mem[32*28 + cnt] = INIT_1C[cnt*9 +: 9];
                mem[32*29 + cnt] = INIT_1D[cnt*9 +: 9];
                mem[32*30 + cnt] = INIT_1E[cnt*9 +: 9];
                mem[32*31 + cnt] = INIT_1F[cnt*9 +: 9];
            end
        end
        else  begin      // INIT_FILE 
//add for initialization RAM     1) load initial data from ini_mem to every mem block  when  cascaded with DRMS
// 2) the ini_mem contain  the whole data of init_file  3) distribute the initdata to every mem in cascaded DRMs
            case(DATA_WIDTH_A)
                1: begin  //DRM TYPE 8K*1
                   for(cnt=0; cnt<1024;cnt = cnt+1)
                       mem[cnt][7:0] = {ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*8+7][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*8+6][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*8+5][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*8+4][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*8+3][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*8+2][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*8+1][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*8][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH]};
                end
                2: begin //DRM TYPE 4K*2
                   for(cnt=0; cnt<1024;cnt = cnt+1)
                       mem[cnt][7:0] = {ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*4+3][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*4+2][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*4+1][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*4][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH]};
                end
                4: begin //DRM TYPE 2K*4
                   for(cnt=0; cnt<1024;cnt = cnt+1)
                       {mem[cnt][7:0]} = {ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*2+1][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                          ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*2][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH]};
                end
                8: begin //DRM TYPE 1K*8
                   for(cnt=0; cnt<1024;cnt = cnt+1)
                       mem[cnt][7:0] = ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH];
                end
                9: begin //DRM TYPE 1K*9
                   for(cnt=0; cnt<1024;cnt = cnt+1)
                       mem[cnt] = ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH];
                end
                16:begin //DRM TYPE 512*16
                   for(cnt=0; cnt<512;cnt = cnt+1)
                       {mem[cnt*2+1][7:0], mem[cnt*2][7:0]} = ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH];
                end
                18:begin //DRM TYPE 512*18
                   for(cnt=0; cnt<512;cnt = cnt+1)
                       {mem[cnt*2+1], mem[cnt*2]} = ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH];
                end
                32:begin //DRM TYPE 256*32
                   for(cnt=0; cnt<256;cnt = cnt+1)
                       {mem[cnt*4+3][7:0],mem[cnt*4+2][7:0],mem[cnt*4+1][7:0],mem[cnt*4][7:0]} = ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH];
                end
                36:begin //DRM TYPE 256*36
                   for(cnt=0; cnt<256;cnt = cnt+1)
                       {mem[cnt*4+3],mem[cnt*4+2],mem[cnt*4+1],mem[cnt*4]} = ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH];
                end
            endcase
        end
    end

    //always @(posedge CLKA) begin
    //    if (CEA)
    //        csa_reg <= CSA;
    //end
    always @(posedge CLKA) begin
        if (CEA) begin
            // high to hold the address
            if (ADDRA_HOLD == 1'b0) begin
                ada_reg <= ADDRA;
            end
            da_reg[17:0] <= DIA[17:0];
            wea_reg <= WEA;
        end
    end
    //always @(posedge CLKB) begin
    //    if (CEB)
    //        csb_reg <= CSB;
    //end
    always @(posedge CLKB) begin
        if (CEB) begin
            // high to hold the address
            if (ADDRB_HOLD == 1'b0) begin
                adb_reg <= ADDRB;
            end
                web_reg <= WEB;
        end
    end
    // byte write enable
    assign bea_reg = ada_reg[3:0];   // modify for byte_write_enable bug
    assign beb_reg = adb_reg[1:0];

    ///////////////////
    // task & function
    ///////////////////

    function [DATA_WIDTH_A-1:0] mem_read_a;
        input [12:0]  addr;
    begin
        case (DATA_WIDTH_A)
            1: mem_read_a = mem[addr[12:3]][addr[2:0]];
            2: mem_read_a = mem[addr[12:3]][addr[2:1]*2 +: 2];
            4: mem_read_a = mem[addr[12:3]][addr[2]*4 +: 4];
            8: mem_read_a = mem[addr[12:3]][7:0];
            9: mem_read_a = mem[addr[12:3]];
            16: mem_read_a = {mem[addr[12:4]*2+1][7:0], mem[addr[12:4]*2][7:0]};
            18: mem_read_a = {mem[addr[12:4]*2+1],      mem[addr[12:4]*2]};
            32: mem_read_a = {mem[addr[12:5]*4+3][7:0], mem[addr[12:5]*4+2][7:0],
                              mem[addr[12:5]*4+1][7:0], mem[addr[12:5]*4][7:0]};
            36: mem_read_a = {mem[addr[12:5]*4+3],      mem[addr[12:5]*4+2],
                              mem[addr[12:5]*4+1],      mem[addr[12:5]*4]};
            default:      ;//null 
        endcase
    end
    endfunction

    function [DATA_WIDTH_B-1:0] mem_read_b;
        input [12:0] addr;
    begin
        case (DATA_WIDTH_B)
            1: mem_read_b = mem[addr[12:3]][addr[2:0]];
            2: mem_read_b = mem[addr[12:3]][addr[2:1]*2 +: 2];
            4: mem_read_b = mem[addr[12:3]][addr[2]*4 +: 4];
            8: mem_read_b = mem[addr[12:3]][7:0];
            9: mem_read_b = mem[addr[12:3]];
            16: mem_read_b = {mem[addr[12:4]*2+1][7:0], mem[addr[12:4]*2][7:0]};
            18: mem_read_b = {mem[addr[12:4]*2+1],      mem[addr[12:4]*2]};
            32: mem_read_b = {mem[addr[12:5]*4+3][7:0], mem[addr[12:5]*4+2][7:0],
                              mem[addr[12:5]*4+1][7:0], mem[addr[12:5]*4][7:0]};
            36: mem_read_b = {mem[addr[12:5]*4+3],      mem[addr[12:5]*4+2],
                              mem[addr[12:5]*4+1],      mem[addr[12:5]*4]};
            default:      ;//null
        endcase
    end
    endfunction

    task mem_write_a;
        input [12:0] addr;
        input [35:0] data;
        input [3:0]  byte_en;
    begin
        case (DATA_WIDTH_A)
            1: mem[addr[12:3]][addr[2:0]] = data[0];
            2: mem[addr[12:3]][addr[2:1]*2 +: 2] = data[1:0];
            4: mem[addr[12:3]][addr[2]*4 +: 4] = data[3:0];
            8: mem[addr[12:3]][7:0] = data[7:0];
            9: mem[addr[12:3]] = data[8:0];
            16: begin
                if (byte_en[1])
                    mem[addr[12:4]*2+1][7:0] = data[16:9];
                if (byte_en[0])
                    mem[addr[12:4]*2][7:0]   = data[7:0];
            end
            18: begin
                if (byte_en[1])
                    mem[addr[12:4]*2+1] = data[17:9];
                if (byte_en[0])
                    mem[addr[12:4]*2]   = data[8:0];
            end
            32: begin
                if (byte_en[3])
                    mem[addr[12:5]*4+3][7:0] = data[34:27];
                if (byte_en[2])
                    mem[addr[12:5]*4+2][7:0] = data[25:18];
                if (byte_en[1])
                    mem[addr[12:5]*4+1][7:0] = data[16:9];
                if (byte_en[0])
                    mem[addr[12:5]*4][7:0]   = data[7:0];
            end
            36: begin
                if (byte_en[3])
                    mem[addr[12:5]*4+3] = data[35:27];
                if (byte_en[2])
                    mem[addr[12:5]*4+2] = data[26:18];
                if (byte_en[1])
                    mem[addr[12:5]*4+1] = data[17:9];
                if (byte_en[0])
                    mem[addr[12:5]*4]   = data[8:0];
            end
            default:     ;//null
        endcase
    end
    endtask

    task mem_write_b;
        input [12:0] addr;
        input [17:0] data;
        input [3:0]  byte_en;
    begin
        case (DATA_WIDTH_B)
            1: mem[addr[12:3]][addr[2:0]] = data[0];
            2: mem[addr[12:3]][addr[2:1]*2 +: 2] = data[1:0];
            4: mem[addr[12:3]][addr[2]*4 +: 4] = data[3:0];
            8: mem[addr[12:3]][7:0] = data[7:0];
            9: mem[addr[12:3]] = data[8:0];
            16: begin
                if (byte_en[1])
                    mem[addr[12:4]*2+1][7:0] = data[16:9];
                if (byte_en[0])
                    mem[addr[12:4]*2][7:0]   = data[7:0];
            end
            18: begin
                if (byte_en[1])
                    mem[addr[12:4]*2+1] = data[17:9];
                if (byte_en[0])
                    mem[addr[12:4]*2]   = data[8:0];
            end
            default:     ;//null
        endcase
    end
    endtask

    ///////////////
    // memory core
    ///////////////
reg CLKA_active;
reg CLKB_active;
initial begin
  CLKA_active = 1'b0;
  CLKB_active = 1'b0;
end
always @(posedge CLKA) begin
   if (CEA) begin
      CLKA_active <= 1'b1;
      #0.2 CLKA_active = 1'b0;
   end
   else
      CLKA_active <= 1'b0;
end
always @(posedge CLKB) begin
   if (CEB) begin
      CLKB_active <= 1'b1;
      #0.2 CLKB_active = 1'b0;
   end
   else
      CLKB_active <= 1'b0;
end

generate
////////////////////////////////////////////////////////////////////////////////////////////
// ROM or SINGLE_PORT 
////////////////////////////////////////////////////////////////////////////////////////////
if(RAM_MODE == "ROM" || RAM_MODE == "SINGLE_PORT") begin:ROMorSP_MODE  //1 no clock region switch  2 no mix width

    always @(posedge CLKA) begin    //modify for db_reg syn with CLKA
        if (CEA)
            db_reg[17:0] <= DIB[17:0];
    end
    if (DATA_WIDTH_A >= 32 || DATA_WIDTH_B >= 32) begin

        assign write_en_a = (wea_reg == 1'b1);
        assign read_en_b  = (web_reg == 1'b0);
        // Port A operations
        always @(negedge CLKA_active) begin
            if (write_en_a) begin  // write
                mem_write_a(ada_reg, {db_reg[17:0], da_reg[17:0]}, bea_reg[3:0]);
            end
        end
        always@(negedge CLKB_active or posedge rstb_int) begin
            if (rstb_int)
               {b_out[width_b-1:0], a_out[width_b-1:0]} = 'b0;
            else if(read_en_b)
               {b_out[width_b-1:0], a_out[width_b-1:0]} = mem_read_b(adb_reg);
        end

    end
    else  begin   //x1 x2 x4 x8 x9 x16 x18 

        assign write_en_a = (wea_reg == 1'b1);
        assign read_en_a  = (wea_reg == 1'b0);
        always @(negedge CLKA_active) begin
            if (write_en_a)  begin  // write
               // read during write
               if (WRITE_MODE_A == "TRANSPARENT_WRITE") begin
                   a_out[width_a-1:0] = mem_read_a(ada_reg);

                   if(DATA_WIDTH_A == 16) begin
                       if(bea_reg[0])
                           a_out[7:0] = da_reg[7:0];
                       else
                           a_out[7:0] = a_out[7:0];

                       if(bea_reg[1])
                           a_out[15:8] = da_reg[16:9];
                       else
                           a_out[15:8] = a_out[15:8];
                   end
                   else if(DATA_WIDTH_A == 18) begin
                        if(bea_reg[0])
                            a_out[8:0] = da_reg[8:0];
                        else
                            a_out[8:0] = a_out[8:0];

                        if(bea_reg[1])
                            a_out[17:9] = da_reg[17:9];
                        else
                            a_out[17:9] = a_out[17:9];
                   end
                   else begin
                      a_out[width_a-1:0] = da_reg[width_a-1:0];
                   end
               end
               else if (WRITE_MODE_A == "READ_BEFORE_WRITE")
                   a_out[width_a-1:0] = mem_read_a(ada_reg);

               mem_write_a(ada_reg, da_reg[17:0], {2'b0,bea_reg[1:0]});
            end
        end
        always @(negedge CLKA_active or posedge rsta_int) begin
            if (rsta_int)
               a_out[width_a-1:0] = 'b0;
            else if (read_en_a)          // read 
               a_out[width_a-1:0] = mem_read_a(ada_reg);
        end
        // Port B operations

    end
end
////////////////////////////////////////////////////////////////////////////////////////////
//SIMPLE_DUAL_PORT
////////////////////////////////////////////////////////////////////////////////////////////
else if(RAM_MODE == "SIMPLE_DUAL_PORT")begin:SDP_MODE  //1 clock region switch 2 mix width
    //port_A operation: only write in SDP MODE
    if (DATA_WIDTH_A >= 32) begin:PORTA

        assign write_en_a = (wea_reg == 1'b1);

        always @(posedge CLKA) begin
           if (CEA)
              db_reg[17:0]  <= DIB[17:0];   //the valid width of db_reg is equal to da_reg
        end
        always @(negedge CLKA_active) begin
           if (write_en_a)    // write 
              mem_write_a(ada_reg, {db_reg[17:0], da_reg[17:0]},bea_reg[3:0]);
        end
    end
    else  begin:PORTA    //  x1 x2 x4 x8 x9 x16 x18 

        assign write_en_a = (wea_reg == 1'b1);

        always @(negedge CLKA_active) begin
           if (write_en_a)     // write 
              mem_write_a(ada_reg, da_reg[17:0], {2'b0,bea_reg[1:0]});
        end
    end
    //port_B operation:only read in SDP MODE
    if (DATA_WIDTH_B >= 32) begin:PORTB
// SIMPLE_DUAL_PORT 
        assign read_en_b  = (web_reg == 1'b0);

        always @(negedge CLKB_active or posedge rstb_int) begin
           if (rstb_int)
              {b_out[width_b-1 : 0], a_out[width_b-1 : 0]} = 'b0;
           else if (read_en_b)       // read 
              {b_out[width_b-1 : 0], a_out[width_b-1 : 0]} = mem_read_b(adb_reg);
        end
    end
    else  begin:PORTB  //  x1 x2 x4 x8 x9 x16 x18 

        assign read_en_b  = (web_reg == 1'b0);

        always @(negedge CLKB_active or posedge rstb_int) begin
           if (rstb_int)
              b_out[width_b-1 : 0] = 'b0;
           else if (read_en_b)   //  read 
              b_out[width_b-1 : 0] = mem_read_b(adb_reg);
        end
    end
end
////////////////////////////////////////////////////////////////////////////////////////////
//DP_MODE
////////////////////////////////////////////////////////////////////////////////////////////
else   begin:DP_MODE   //  --x1 x2 x4 x8 x9 x16 x18--    1) no clock region switch   2)mix width
    assign write_en_a = (wea_reg == 1'b1) ;
    assign read_en_a  = (wea_reg == 1'b0) ;
    assign write_en_b = (web_reg == 1'b1) ;
    assign read_en_b  = (web_reg == 1'b0) ;
    // Port A operations
    always @(negedge CLKA_active ) begin
        if (write_en_a)  begin  // write
            // read during write
            if (WRITE_MODE_A == "TRANSPARENT_WRITE") begin
               a_out[width_a-1:0] = mem_read_a(ada_reg);

               if(DATA_WIDTH_A == 16) begin
                   if(bea_reg[0])
                       a_out[7:0] = da_reg[7:0];
                   else
                       a_out[7:0] = a_out[7:0];

                   if(bea_reg[1])
                       a_out[15:8] = da_reg[16:9];
                   else
                       a_out[15:8] = a_out[15:8];
               end
               else if(DATA_WIDTH_A == 18) begin
                    if(bea_reg[0])
                        a_out[8:0] = da_reg[8:0];
                    else
                        a_out[8:0] = a_out[8:0];

                    if(bea_reg[1])
                        a_out[17:9] = da_reg[17:9];
                    else
                        a_out[17:9] = a_out[17:9];
               end
               else begin
                  a_out[width_a-1:0] = da_reg[width_a-1:0];
               end
            end
            else if (WRITE_MODE_A == "READ_BEFORE_WRITE")
                a_out[width_a-1 : 0] = mem_read_a(ada_reg);

            mem_write_a(ada_reg, da_reg[17:0], {2'b0,bea_reg[1:0]});
        end
    end
    always @(negedge CLKA_active or posedge rsta_int) begin
        if (rsta_int)
           a_out[width_a-1 : 0] = 'b0;
        else if (read_en_a)
           a_out[width_a-1 : 0] = mem_read_a(ada_reg);
    end
    // Port B operations
    always @(posedge CLKB) begin  // modify for db_reg syn with CLKB
         if (CEB)
            db_reg[17:0] <= DIB[17:0];
    end

    always @(negedge CLKB_active ) begin
        if (write_en_b)  begin  // write
            // read during write
            if (WRITE_MODE_B == "TRANSPARENT_WRITE") begin

                b_out[width_b-1:0] = mem_read_b(adb_reg);

                if(DATA_WIDTH_B == 16) begin
                    if(beb_reg[0])
                        b_out[7:0] = db_reg[7:0];
                    else
                        b_out[7:0] = b_out[7:0];

                    if(beb_reg[1])
                        b_out[15:8] = db_reg[16:9];
                    else
                        b_out[15:8] = b_out[15:8];
                end
                else if(DATA_WIDTH_B == 18) begin
                    if(beb_reg[0])
                        b_out[8:0] = db_reg[8:0];
                    else
                        b_out[8:0] = b_out[8:0];

                    if(beb_reg[1])
                        b_out[17:9] = db_reg[17:9];
                    else
                        b_out[17:9] = b_out[17:9];
                end
                else begin
                   b_out[width_b-1:0] = db_reg[width_b-1:0];
                end
            end
            else if (WRITE_MODE_B == "READ_BEFORE_WRITE")
                b_out[width_b-1 : 0] = mem_read_b(adb_reg);

            mem_write_b(adb_reg, db_reg[17:0], {2'b0,beb_reg[1:0]});
        end
    end
    always @(negedge CLKB_active or posedge rstb_int) begin
        if (rstb_int)
           b_out[width_b-1 : 0] = 'b0;
        else if (read_en_b)
           b_out[width_b-1 : 0] = mem_read_b(adb_reg);
    end
end

endgenerate

    //////////////
    // core latch
    //////////////
    assign grsn =  (GRS_EN == "TRUE") ? GRS_INST.GRSNET : 1'b1;
    assign grs =  ~grsn;
    or (rsta_grs, grs, RSTA);
    or (rstb_grs, grs, RSTB);

wire CLKA_for_or,CLKB_for_or;
    // async reset
reg rsta_grsn_d;

    always @(posedge CLKA_for_or ) begin
        if (RSTA) begin
            rsta_grsn_d   <= 1'b1;
        end
        else begin
            rsta_grsn_d   <= 1'b0;
        end
    end

    always @(posedge CLKA_for_or or posedge RSTA) begin
        if (RSTA) begin
            rsta_async_sy <= 1'b1;
        end
        else begin
            rsta_async_sy <= rsta_grsn_d;
        end
    end

reg rstb_grsn_d;
    always @(posedge CLKB_for_or) begin
        if (RSTB) begin
            rstb_grsn_d   <= 1'b1;
        end
        else begin
            rstb_grsn_d   <= 1'b0;
        end
    end

    always @(posedge CLKB_for_or or posedge RSTB) begin
        if (RSTB) begin
            rstb_async_sy <= 1'b1;
        end
        else begin
            rstb_async_sy <= rstb_grsn_d;
        end
    end

initial begin
    rsta_grsn_d = 1'b1;
    rsta_async_sy = 1'b1;
    rstb_grsn_d = 1'b1;
    rstb_async_sy = 1'b1;
end

assign rsta_grs_sync  = (RST_TYPE == "SYNC") ? rsta_grsn_d : 1'b0; //register to match with CLKA_ative falling edge
assign rstb_grs_sync  = (RST_TYPE == "SYNC") ? rstb_grsn_d : 1'b0; //register to match with CLKA_ative falling edge
assign rsta_grs_async = (RST_TYPE == "ASYNC") ? rsta_grs : grs;
assign rstb_grs_async = (RST_TYPE == "ASYNC") ? rstb_grs : grs;
assign rsta_async_synrel = rsta_grs | rsta_async_sy;
assign rstb_async_synrel = rstb_grs | rstb_async_sy;
assign rsta_int = (RST_TYPE == "ASYNC_SYNC_RELEASE") ? rsta_async_synrel : rsta_grs_sync | rsta_grs_async;
assign rstb_int = (RST_TYPE == "ASYNC_SYNC_RELEASE") ? rstb_async_synrel : rstb_grs_sync | rstb_grs_async;
/////////////////////////////////////////////////////////////////////
//port out
assign CLKA_for_or = (DOA_REG_CLKINV == 1) ? ~CLKA : CLKA;
assign CLKB_for_or = (DOB_REG_CLKINV == 1) ? ~CLKB : CLKB;
generate
if (DATA_WIDTH_B >= 32) begin:FAKE_DP_OUT
    ///////////////////
    // output register
    ///////////////////
    always @(posedge CLKB_for_or or posedge rstb_int) begin
        if (rstb_int)
            a_out_reg <= 0;
        else if (ORCEB)
            a_out_reg[width_b-1 : 0] <= a_out[width_b-1 : 0];
    end
    //doa combination logic
    always @(*) begin
        if (DOB_REG == 0)
        begin
            case(DATA_WIDTH_B)
                32: {doa[16:9],doa[7:0]} = {a_out[15:8],a_out[7:0]};
                36:  doa[width_b-1:0] = a_out[width_b-1:0]        ;
            endcase
        end
        else
        begin
            case(DATA_WIDTH_B)
                32: {doa[16:9],doa[7:0]} = {a_out_reg[15:8],a_out_reg[7:0]};
                36:  doa[width_b-1:0] = a_out_reg[width_b-1 : 0];
            endcase
        end
    end

    //port_B output
    always @(posedge CLKB_for_or or posedge rstb_int) begin
        if (rstb_int)
            b_out_reg <= 0;
        else if (ORCEB)
            b_out_reg[width_b-1 : 0] <= b_out[width_b-1 : 0];
    end
    //dob combination logic
    always @(*) begin
        if (DOB_REG == 0)
        begin
            case(DATA_WIDTH_B)
                32:{dob[16:9],dob[7:0]} = {b_out[15:8],b_out[7:0]};
                36: dob[width_b-1:0] = b_out[width_b-1 : 0];
            endcase
        end
        else
        begin
            case(DATA_WIDTH_B)
                32:{dob[16:9],dob[7:0]} = {b_out_reg[15:8],b_out_reg[7:0]};
                36: dob[width_b-1:0] = b_out_reg[width_b-1 : 0];
            endcase
        end
    end
end
else  begin:TRUE_DP_OUT   // x1 x2 x4 x8 x9 x16 x18    

    //port_A output
    always @(posedge CLKA_for_or or posedge rsta_int) begin
        if (rsta_int)
            a_out_reg <= 0;
        else if (ORCEA)
            a_out_reg[width_a-1 : 0] <= a_out[width_a-1 : 0];
    end
    //doa combination logic
    always @(*) begin
        if (DOA_REG == 0)
        begin
            case(DATA_WIDTH_A)
               1: {doa[16:9],doa[7:0]} = {16{a_out[width_a-1:0]}};
               2: {doa[16:9],doa[7:0]} = { 8{a_out[width_a-1:0]}};
               4: {doa[16:9],doa[7:0]} = { 4{a_out[width_a-1:0]}};
               8: {doa[16:9],doa[7:0]} = { 2{a_out[width_a-1:0]}};
               9: {doa[17:9],doa[8:0]} = { 2{a_out[width_a-1:0]}};
               16:{doa[16:9],doa[7:0]} =     a_out[width_a-1:0]  ;
               18: doa[17:0]          =     a_out[width_a-1:0]  ;
            endcase
        end
        else
        begin
            case(DATA_WIDTH_A)
               1: {doa[16:9],doa[7:0]} = {16{a_out_reg[width_a-1:0]}};
               2: {doa[16:9],doa[7:0]} = { 8{a_out_reg[width_a-1:0]}};
               4: {doa[16:9],doa[7:0]} = { 4{a_out_reg[width_a-1:0]}};
               8: {doa[16:9],doa[7:0]} = { 2{a_out_reg[width_a-1:0]}};
               9: {doa[17:9],doa[8:0]} = { 2{a_out_reg[width_a-1:0]}};
               16:{doa[16:9],doa[7:0]} =     a_out_reg[width_a-1:0] ;
               18: doa[17:0]          =     a_out_reg[width_a-1:0] ;
            endcase
        end
    end

    //port_B output
    always @(posedge CLKB_for_or or posedge rstb_int) begin
        if (rstb_int)
            b_out_reg <= 0;
        else if (ORCEB)
            b_out_reg[width_b-1 : 0] <= b_out[width_b-1 : 0];
    end
    //dob combination logic
    always @(*) begin
        if (DOB_REG == 0)
        begin
            case(DATA_WIDTH_B)
               1: {dob[16:9],dob[7:0]} = {16{b_out[width_b-1:0]}};
               2: {dob[16:9],dob[7:0]} = { 8{b_out[width_b-1:0]}};
               4: {dob[16:9],dob[7:0]} = { 4{b_out[width_b-1:0]}};
               8: {dob[16:9],dob[7:0]} = { 2{b_out[width_b-1:0]}};
               9: {dob[17:9],dob[8:0]} = { 2{b_out[width_b-1:0]}};
               16:{dob[16:9],dob[7:0]} =     b_out[width_b-1:0] ;
               18: dob[17:0]          =     b_out[width_b-1:0] ;
            endcase
        end
        else
            case(DATA_WIDTH_B)
               1: {dob[16:9],dob[7:0]} = {16{b_out_reg[width_b-1:0]}};
               2: {dob[16:9],dob[7:0]} = { 8{b_out_reg[width_b-1:0]}};
               4: {dob[16:9],dob[7:0]} = { 4{b_out_reg[width_b-1:0]}};
               8: {dob[16:9],dob[7:0]} = { 2{b_out_reg[width_b-1:0]}};
               9: {dob[17:9],dob[8:0]} = { 2{b_out_reg[width_b-1:0]}};
               16:{dob[16:9],dob[7:0]} =     b_out_reg[width_b-1:0] ;
               18: dob[17:0]          =     b_out_reg[width_b-1:0] ;
            endcase
    end
end

endgenerate
assign DOA = doa;
assign DOB = dob;

// synthesis translate_on
endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2016 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_ADC_E2.v
//
// Functional description: ADC_E2
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////
`timescale 1 ns / 1 ps



module GTP_ADC_E2
#(
    parameter [15:0] CREG_00H = 16'h0001,
    parameter [15:0] CREG_01H = 16'hC83F,
    parameter [15:0] CREG_02H = 16'h0009,
    parameter [13:0] CREG_31H = 14'h0000,
    parameter [15:0] CREG_03H = 16'h0000,
    parameter [15:0] CREG_04H = 16'h0000,
    parameter [15:0] CREG_0AH = 16'h0000,
    parameter [15:0] CREG_05H = 16'h0000,
    parameter [15:0] CREG_06H = 16'h0000,
    parameter [15:0] CREG_0CH = 16'h0000,
    parameter [15:0] CREG_07H = 16'h0000,
    parameter [15:0] CREG_08H = 16'h0000,
    parameter [15:0] CREG_0EH = 16'h0000,
    parameter [11:0] CREG_20H = 12'h000,//TEMP_SENSOR_HIGH
    parameter [11:0] CREG_21H = 12'h000,//TEMP_SENSOR_LOW
    parameter [11:0] CREG_22H = 12'h000,//VCC_HIGH
    parameter [11:0] CREG_23H = 12'h000,//VCC_LOW
    parameter [11:0] CREG_24H = 12'h000,//VCCA_HIGH
    parameter [11:0] CREG_25H = 12'h000,//VCCA_LOW
    parameter [11:0] CREG_26H = 12'h000,//VCC_DRM_HIGH
    parameter [11:0] CREG_27H = 12'h000,//VCC_DRM_LOW
    parameter [11:0] CREG_28H = 12'h000,//VCC_CRAM_HIGH
    parameter [11:0] CREG_29H = 12'h000,//VCC_CRAM_LOW
    parameter [11:0] CREG_2AH = 12'hCC2,//OVER_TEMP_LIMIT
    parameter [11:0] CREG_2BH = 12'hA5B//OVER_TEMP_RESET
    //parameter        ADC_EN = "FALSE"
)(
    //Analog Input
    input [1:0]VA, //0:N, 1:P
    input [31:0] VAUX, //even:N, odd:P

    //APB
    input DCLK, //PCLK,
    input [7:0] DADDR, //PADDR,
    input DEN, //PSEL,
    input SECEN, //PENABLE
    input DWE, //PWRITE,
    input [15:0] DI, //PWDATA,
    output [15:0] DO, //PRDATA,
    output DRDY, //PREADY,

    //SRB
    input           CONVST, //EVENT_DRV,
    input           RST_N,
    input           LOADSC_N,//LOAD_SC_N,
    output          OVER_TEMP,
    output          LOGIC_DONE_A,
    output          LOGIC_DONE_B,
    output          ADC_CLK_OUT,
    output          DMODIFIED, //PMODIFIED,
    output [4:0]    ALARM   
);
//synthesis translate_off
    
      
    
    //Analog Input
    reg I10U_BG     ;
    reg VREF_INT    ;
    reg POR_N_1P8V  ;
    reg VREFADC_P   ;
    reg VREFADC_N   ;
    //reg TSDP        ;
    //reg TSDN        ;
    //JTAG
    reg TCK      ;
    reg CLOCKDR  ;
    reg SHIFTDR  ;
    reg TDI      ;
    reg UPDATEDR ;
    reg FLG_JTAG ;
    reg CAPTUREDR;

    reg           GWEN          ;
    reg           GLOGEN        ;
    reg           POR_N         ;
    reg           CLK_OSC       ;
    reg           AD_TRIM_MODE  ;
    reg [11:0]    AD_TEMP_OFFSET;
    
    initial
    begin
    
    //Analog Input
        I10U_BG      = 1'b1;
        VREF_INT     = 1'b0;
        POR_N_1P8V   = 1'b0;
        VREFADC_P    = 1'b1;
        VREFADC_N    = 1'b0;
    //JTAG
        TCK       = 1'b0;
        CLOCKDR   = 1'b0;
        SHIFTDR   = 1'b0;
        TDI       = 1'b0;
        UPDATEDR  = 1'b0;
        FLG_JTAG  = 1'b0;
        CAPTUREDR = 1'b0;
        CLK_OSC   = 1'b0;

        GWEN           = 1'b0;
        GLOGEN         = 1'b0;
        POR_N          = 1'b0;
        AD_TRIM_MODE   = 1'b0;
        AD_TEMP_OFFSET = 0;
        #500
        POR_N          = 1'b1;
        POR_N_1P8V   = 1'b1;
        #22500
        GWEN           = 1'b1;
        GLOGEN         = 1'b1;
    end

    always #9.615 CLK_OSC = ~CLK_OSC;//2019/12/05,update
    
    wire [15:0] SC_CREG_00H;
    wire [15:0] SC_CREG_01H;
    wire [15:0] SC_CREG_02H;
    wire [13:0] SC_CREG_31H;
    wire [15:0] SC_SEQ_03H;
    wire [15:0] SC_SEQ_04H;
    wire [15:0] SC_SEQ_05H;
    wire [15:0] SC_SEQ_06H;
    wire [15:0] SC_SEQ_07H;
    wire [15:0] SC_SEQ_08H;
    wire [15:0] SC_SEQ_0AH;
    wire [15:0] SC_SEQ_0CH;
    wire [15:0] SC_SEQ_0EH;
    wire [11:0] SC_ALM_20H;
    wire [11:0] SC_ALM_21H;
    wire [11:0] SC_ALM_22H;
    wire [11:0] SC_ALM_23H;
    wire [11:0] SC_ALM_24H;
    wire [11:0] SC_ALM_25H;
    wire [11:0] SC_ALM_26H;
    wire [11:0] SC_ALM_27H;
    wire [11:0] SC_ALM_28H;
    wire [11:0] SC_ALM_29H;
    wire [11:0] SC_ALM_2AH;
    wire [11:0] SC_ALM_2BH;
    //wire        SC_ADC_EN;
    
    assign SC_CREG_00H = CREG_00H;
    assign SC_CREG_01H = CREG_01H;
    assign SC_CREG_02H = CREG_02H;
    assign SC_CREG_31H = CREG_31H;
    assign SC_SEQ_03H  = CREG_03H;
    assign SC_SEQ_04H  = CREG_04H;
    assign SC_SEQ_0AH  = CREG_0AH;
    assign SC_SEQ_05H  = CREG_05H;
    assign SC_SEQ_06H  = CREG_06H;
    assign SC_SEQ_0CH  = CREG_0CH;
    assign SC_SEQ_07H  = CREG_07H;
    assign SC_SEQ_08H  = CREG_08H;
    assign SC_SEQ_0EH  = CREG_0EH;
    assign SC_ALM_20H  = CREG_20H;
    assign SC_ALM_21H  = CREG_21H;
    assign SC_ALM_22H  = CREG_22H;
    assign SC_ALM_23H  = CREG_23H;
    assign SC_ALM_24H  = CREG_24H;
    assign SC_ALM_25H  = CREG_25H;
    assign SC_ALM_26H  = CREG_26H;
    assign SC_ALM_27H  = CREG_27H;
    assign SC_ALM_28H  = CREG_28H;
    assign SC_ALM_29H  = CREG_29H;
    assign SC_ALM_2AH  = CREG_2AH;
    assign SC_ALM_2BH  = CREG_2BH;
    //assign SC_ADC_EN   =(ADC_EN == "FALSE") ? 1'b0 : 1'b1; 

    /////signal begin/////
    wire           temps_clk_en           ; 
    wire           temps_rstn             ; 
    wire           adc_clk                ; 
    wire           adc_rstn_a             ; 
    wire           adc_rstn_b             ; 
    wire [1:0]     adc_pd                 ; 
    wire [13:0]    ibias_ctrl             ; 
    wire [1:0]     scale_ctrl             ; 
    wire [1:0]     vcm_ctrl               ; 
    wire           vref_type_sel          ; 
    wire           adc_bipolar_en_a       ; 
    wire           adc_clk_en_a           ; 
    wire [3:0]     vaa_chsel_a            ; 
    wire [3:0]     input_chsel_a          ; 
    wire [1:0]     input_res_vaach_ctrl_a ; 
    wire           adc_bipolar_en_b       ; 
    wire           adc_clk_en_b           ; 
    wire [3:0]     vaa_chsel_b            ; 
    wire [3:0]     input_chsel_b          ; 
    wire [1:0]     input_res_vaach_ctrl_b ; 
    wire           adca_sh_outp           ; 
    wire           adca_sh_outn           ; 
    wire  [11:0]   adca_data              ; 
    wire           adca_done              ; 
    wire           adcb_sh_outp           ; 
    wire           adcb_sh_outn           ; 
    wire  [11:0]   adcb_data              ; 
    wire           adcb_done              ; 



    ////instance/////
    adc_e2_logic_top   adc_logic_top
     (
///////////////////////////////////////////////////////////////////////
    .ad_temp_clk_en            (temps_clk_en            ) ,
    .ad_temp_rstn              (temps_rstn              ) ,
    .ad_clk                    (adc_clk                 ) ,
    .ad_rstn_a                 (adc_rstn_a                ) ,
    .ad_rstn_b                 (adc_rstn_b) ,
    .ad_bias_pd                (adc_pd                  ) ,
    .ad_ibias_ctrl             (ibias_ctrl              ) ,
    .ad_scale_ctrl             (scale_ctrl              ) ,
    .ad_vcm_in                 (vcm_ctrl                ) ,
    .ad_vref_sel               (vref_type_sel           ) ,
    .ad_bipolar_en_a           (adc_bipolar_en_a        ) ,
    .ad_clk_en_a               (adc_clk_en_a            ) ,
    .ad_vaa_chsel_a            (vaa_chsel_a             ) ,
    .ad_input_chsel_a          (input_chsel_a           ) ,
    .ad_input_res_vaach_ctrl_a (input_res_vaach_ctrl_a  ) ,
    .ad_bipolar_en_b           (adc_bipolar_en_b        ) ,
    .ad_clk_en_b               (adc_clk_en_b            ) ,
    .ad_vaa_chsel_b            (vaa_chsel_b             ) ,
    .ad_input_chsel_b          (input_chsel_b           ) ,
    .ad_input_res_vaach_ctrl_b (input_res_vaach_ctrl_b  ) ,

    .ad_dat_a                  (adca_data               ) ,
    .ad_done_a                 (adca_done               ) ,
    .ad_dat_b                  (adcb_data               ) ,
    .ad_done_b                 (adcb_done               ) ,
    .logic_done_a              (LOGIC_DONE_A            ) ,
    .logic_done_b              (LOGIC_DONE_B            ) ,

///////////////////////////////////////////////////////////////////////////
    .pclk               (DCLK             ) ,
    .psel               (DEN             ) ,
    .pwrite             (DWE              ) ,
    .paddr              (DADDR            ) ,
    .pwdata             (DI               ) ,
    .prdata             (DO               ) ,
    .penable            (SECEN              ) ,
    .pready             (DRDY             ) ,
    .pmodified          (DMODIFIED        ) ,

    .tck                (TCK              ) ,
    .flg_jtag           (FLG_JTAG         ) ,
    .tdi                (TDI              ) ,
    .tdo                (                 ) ,
    .clockdr            (CLOCKDR          ) ,
    .capturedr          (CAPTUREDR        ) ,
    .shiftdr            (SHIFTDR          ) ,
    .updatedr           (UPDATEDR         ) ,
    
    .sc_creg_00h        (SC_CREG_00H      ) ,
    .sc_creg_01h        (SC_CREG_01H      ) ,
    .sc_creg_02h        (SC_CREG_02H      ) ,
    .sc_creg_31h        (SC_CREG_31H      ) ,
    .sc_seq_03h         (SC_SEQ_03H       ) ,
    .sc_seq_04h         (SC_SEQ_04H       ) ,
    .sc_seq_05h         (SC_SEQ_05H       ) ,
    .sc_seq_06h         (SC_SEQ_06H       ) ,
    .sc_seq_07h         (SC_SEQ_07H       ) ,
    .sc_seq_08h         (SC_SEQ_08H       ) ,
    .sc_seq_0Ah         (SC_SEQ_0AH       ) ,
    .sc_seq_0Ch         (SC_SEQ_0CH       ) ,
    .sc_seq_0Eh         (SC_SEQ_0EH       ) ,
    .sc_alm_20h         (SC_ALM_20H       ) ,
    .sc_alm_21h         (SC_ALM_21H       ) ,
    .sc_alm_22h         (SC_ALM_22H       ) ,
    .sc_alm_23h         (SC_ALM_23H       ) ,
    .sc_alm_24h         (SC_ALM_24H       ) ,
    .sc_alm_25h         (SC_ALM_25H       ) ,
    .sc_alm_26h         (SC_ALM_26H       ) ,
    .sc_alm_27h         (SC_ALM_27H       ) ,
    .sc_alm_28h         (SC_ALM_28H       ) ,
    .sc_alm_29h         (SC_ALM_29H       ) ,
    .sc_alm_2Ah         (SC_ALM_2AH       ) ,
    .sc_alm_2Bh         (SC_ALM_2BH       ) ,
    .sc_adc_en          (1'b1             ) ,//SC_ADC_EN

    .event_drv          (CONVST           ) ,
    .load_sc_n          (LOADSC_N         ) ,
    .rst_n              (RST_N            ) ,
    .gwen               (GWEN             ) ,
    .ad_trim_mode       (AD_TRIM_MODE     ) ,
    .ad_temp_offset     (AD_TEMP_OFFSET   ) ,
    .alarm              (ALARM            ) ,
    .over_temp          (OVER_TEMP        ) ,
    .clk_out            (ADC_CLK_OUT      ) ,
    .glogen             (GLOGEN           ) ,
    .por_n              (POR_N            ) ,
    .over_temp_ccs      (                 ) ,
    .clk_osc            (CLK_OSC          ) ,
    .osc_turn_on        (                 ) ,
    .test_si_0          (1'b1   ) ,
    .test_si_1          (1'b1   ) ,
    .test_si_2          (1'b1   ) ,
    .test_si_3          (1'b1   ) ,
    .test_so_0          (       ) ,
    .test_so_1          (       ) ,
    .test_so_2          (       ) ,
    .test_so_3          (       ) ,
    .test_clk           (1'b1   ) ,
    .test_rst_n         (1'b1   ) ,
    .test_mode_n        (1'b1   ) ,
    .test_scan_en_n     (1'b1   )  
    );

/////instance/////
adc_e2_analog_top ADC_ANALOG_TOP
    (
    .VCCADC                  () ,
    .VCCAUX                  () ,
    .VSSADC                  () ,
    .VSSAUX                  () ,
    .VCC_SENSOR_P            () ,
    .VCC_SENSOR_N            () ,
    .VCCA_SENSOR_P           () ,
    .VCCA_SENSOR_N           () ,
    .VCC_CRAM_SENSOR_P       () ,
    .VCC_CRAM_SENSOR_N       () ,
    .VCC_DRM_SENSOR_P        () ,
    .VCC_DRM_SENSOR_N        () ,
    //.I10U_BG                 (I10U_BG  ) ,
    //.VREF_INT                (VREF_INT ) ,
    .VREFADC_P               (VREFADC_P   ) ,
    .VREFADC_N               (VREFADC_N   ) ,
    .VAADC_P                 (VA[1]          ) ,
    .VAADC_N                 (VA[0]       ) ,
    .VAAP                    ({VAUX[31],VAUX[29],VAUX[27],VAUX[25],VAUX[23],VAUX[21],VAUX[19],VAUX[17],VAUX[15],VAUX[13],VAUX[11],VAUX[9],VAUX[7],VAUX[5],VAUX[3],VAUX[1]}) ,
    .VAAN                    ({VAUX[30],VAUX[28],VAUX[26],VAUX[24],VAUX[22],VAUX[20],VAUX[18],VAUX[16],VAUX[14],VAUX[12],VAUX[10],VAUX[8],VAUX[6],VAUX[4],VAUX[2],VAUX[0]}) ,
    .TBD_P                   () ,
    .TBD_N                   () ,
    .TEMPS_CLK_EN            (temps_clk_en          ) ,
    .TEMPS_RSTN              (temps_rstn            ) ,
    .ADC_CLK                 (adc_clk               ) ,
    .ADC_RSTN_A              (adc_rstn_a            ) ,
    .ADC_RSTN_B              (adc_rstn_b            ) ,
    .ADC_PD                  (adc_pd                ) ,
    .IBIAS_CTRL              (ibias_ctrl            ) ,
    .SCALE_CTRL              (scale_ctrl            ) ,
    .VCM_CTRL                (vcm_ctrl              ) ,
    .VREF_TYPE_SEL           (vref_type_sel         ) ,
    .ADC_BIPOLAR_EN_A        (adc_bipolar_en_a      ) ,
    .ADC_CLK_EN_A            (adc_clk_en_a          ) ,
    .VAA_CHSEL_A             (vaa_chsel_a           ) ,
    .INPUT_CHSEL_A           (input_chsel_a         ) ,
    .INPUT_RES_VAACH_CTRL_A  (input_res_vaach_ctrl_a) ,
    .ADC_BIPOLAR_EN_B        (adc_bipolar_en_b      ) ,
    .ADC_CLK_EN_B            (adc_clk_en_b          ) ,
    .VAA_CHSEL_B             (vaa_chsel_b           ) ,
    .INPUT_CHSEL_B           (input_chsel_b         ) ,
    .INPUT_RES_VAACH_CTRL_B  (input_res_vaach_ctrl_b) ,
    .ADCA_DATA               (adca_data             ) ,
    .ADCA_DONE               (adca_done             ) ,
    .ADCB_DATA               (adcb_data             ) ,
    .ADCB_DONE               (adcb_done             ) ,
    .ADC_VREFP_CP            (                      ) ,
    .TSDP                    (                      ) ,
    .TSDN                    (                      )     
    );

//synthesis translate_on
endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_MULT18.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

//P=A*B
module GTP_MULT18 #(
    parameter GRS_EN    = "TRUE", //"TRUE"; "FALSE"
    parameter SYNC_RST  = "FALSE", //"TRUE"; "FALSE"
    parameter INREG_EN  = "FALSE", //"TRUE"; "FALSE"
    parameter OUTREG_EN = "FALSE"  //"TRUE"; "FALSE"
) (
    output  [36-1:0] P,
    input   CE,
    input   RST,
    input   CLK,
    input   A_SIGNED,
    input   [18-1:0] A,
    input   B_SIGNED,
    input   [18-1:0] B
);


    INT_PREADD_MULT #(
        .GRS_EN(GRS_EN),
        .SYNC_RST(SYNC_RST),
        .INREG_EN(INREG_EN),
        .OUTREG_EN(OUTREG_EN),
        .ASIZE(18),
        .BSIZE(18),
        .PREADD_EN(0)
    ) U_INT_MULT (
        .CE(CE),
        .RST(RST),
        .CLK(CLK),
        .A_SIGNED(A_SIGNED),
        .A(A),
        .B_SIGNED(B_SIGNED),
        .B(B),
        .C_SIGNED(B_SIGNED),
        .C(18'b0),
        .PREADDSUB(1'b0),
        .P(P)
    );

endmodule






//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_APB.v
//
// Functional description: APB Circuit
//
// Parameter description:
//      
//
// Port description:
//      
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////
`timescale 1 ns / 1 ps

module GTP_APB
#(
    parameter [31:0] IDCODE = 32'haaaa5555,
    parameter [31:0] USERCODE = 32'h0
)
(
input         CLK,
input         RST_N,
input  [4:0]  ADDR,
input         SEL_CCS,
input         SEL_SPI,
input         SEL_I2C0,
input         SEL_I2C1,
input         SEL_TIMER,
input         SEL_PLL0,
input         SEL_PLL1,
input         EN,
input         WR,
input  [7:0]  WDATA,
output [7:0]  RDATA,
output        RDY,
output        IRQ,
output        IRQ_CCS
);

wire            init_complete;
wire            done;
wire            efb_rstb;
wire            efb_en;

wire    [1:0]   U_Seq;
wire    [2:0]   U_Ndac2;
wire    [2:0]   U_Ndac3;
wire    [1:0]   U_Slope;
wire    [2:0]   U_Bdac;
wire    [3:0]   U_Idac, U_Itim;
wire    [3:0]   U_Mode;
wire   [31:0]   U_Din;
wire   [31:0]   dout;
wire            dout_en;
wire   [31:0]   doutg;
wire    [4:0]   U_Ndacp, U_Pdacp, U_Ndace, U_Pdace, U_Rdac;
wire    [5:0]   U_Ca, U_Pa;
wire   [10:0]   U_Ra;
wire            U_Aclk;
wire            U_Axa;
wire            U_Pd1,U_Pd2,U_Sleep,U_Oe;
wire            U_Pe;
wire            U_Pw;
wire            U_Reset;

wire    [1:0]   F_Seq;
wire    [1:0]   F_Wmod, F_Wbytesel, F_Rmod,F_Rbytesel;        
wire    [2:0]   F_Ndac2;
wire    [2:0]   F_Ndac3;
wire    [2:0]   F_Slope;
wire    [3:0]   F_Bdac;
wire    [3:0]   F_Idac, F_Itim;
wire    [3:0]   F_Mode;
wire   [10:0]   F_Tm_reserved;
wire            F_Tm_daa,
                F_Tm_disneg,
                F_Tm_dispos,
                F_Tm_isa,
                F_Tm_itim,    
                F_Pnb;
wire            F_Tm_vhl;    
wire            F_Tm_disrow;
wire            F_Tm_rdhvpl;
wire    [3:0]   F_Tm;
wire   [31:0]   F_Din;
wire    [4:0]   F_Ndacp, F_Pdacp, F_Ndace, F_Pdace,F_Rdac;
 
wire    [6:0]   F_Ca, F_Pa;

wire    [9:0]   F_Ra;
wire            F_Aclk;
wire            F_Axa;
wire            F_Pd1,F_Pd2,F_Sleep,F_Oe;
wire            F_Pe;
wire            F_Pw;
wire            F_Reset;
wire            F_Turbo;

wire            fpclkg;

reg clk;
reg fpclk;
reg rstn;

initial 
    begin
        clk = 1'b0;
        fpclk = 1'b0;
        rstn = 1'b0;
        #10;
        rstn = 1'b1;
    end

always #24.438 clk = ~clk;
always #17 fpclk = ~fpclk;

INT_APB_CCS  INT_APB_CCS (

.idcode               (IDCODE),
.usercode             (USERCODE),

.por_n                (rstn),
.rst_n                (rstn),

.init_n               (init_complete),
.init_complete        (init_complete),

.done_i               (done),
.done                 (done),

.fpclk                (fpclk),
.fpclkg               (fpclkg),

.efb_rstb             (efb_rstb),
.efb_en               (efb_en),

.axa                  (U_Axa),
.ra                   (U_Ra),
.ca                   (U_Ca),
.pa                   (U_Pa),
.mode                 (U_Mode),
.seq                  (U_Seq),
.aclk                 (U_Aclk),
.din                  (U_Din),
.dout                 (dout),
.dout_en              (dout_en),
.pw                   (U_Pw),
.pe                   (U_Pe),
.oe                   (U_Oe),
.pd1                  (U_Pd1),
.pd2                  (U_Pd2),
.reset                (U_Reset),
.sleep                (U_Sleep),

.itim                 (U_Itim),
.idac                 (U_Idac),
.slope                (U_Slope),
.bdac                 (U_Bdac),
.pdace                (U_Pdace),
.pdacp                (U_Pdacp),
.ndace                (U_Ndace),
.ndacp                (U_Ndacp),
.ndac2                (U_Ndac2),
.ndac3                (U_Ndac3),
.rdac                 (U_Rdac),

.glogen_fb            (glogen),
.glogen               (glogen),

.clk                  (clk),

.pctlr_clk            (clk_pctl),
.rstn_pctl            (rstn_pctl),

.pclk                 (CLK),
.presetn              (RST_N),
.paddr                (ADDR),
.psel_ccs             (SEL_CCS),
.psel_spi             (SEL_SPI),
.psel_i2c0            (SEL_I2C0),
.psel_i2c1            (SEL_I2C1),
.psel_timer           (SEL_TIMER),
.psel_pll0            (SEL_PLL0),
.psel_pll1            (SEL_PLL1),
.penable              (EN),
.pwrite               (WR),
.pwdata               (WDATA),
.prdata               (RDATA),
.pready               (RDY),

.irq                  (IRQ),
.irq_ccs              (IRQ_CCS),

.pll0_prdata          (GTP_GRS.pll0_prdata),
.pll0_pready          (GTP_GRS.pll0_pready),

.pll1_prdata          (8'h0),
.pll1_pready          (1'b0),

.rbcrc_clk            (1'b1),
.rbcrc_rst            (1'b1),
.rbcrc_start          (1'b1),
.rbcrc_err            (),
.rbcrc_valid          (),

.spi_ss_i_n           (GTP_GRS.spi_ss_i_n   ),
.spi_ss_o_n           (GTP_GRS.spi_ss_o_n   ),
.spi_sck_oe_n         (GTP_GRS.spi_sck_oe_n ),
.spi_sck_i            (GTP_GRS.spi_sck_i    ),
.spi_sck_o            (GTP_GRS.spi_sck_o    ),
.spi_mosi_oe_n        (GTP_GRS.spi_mosi_oe_n),
.spi_mosi_i           (GTP_GRS.spi_mosi_i   ),
.spi_mosi_o           (GTP_GRS.spi_mosi_o   ),
.spi_miso_oe_n        (GTP_GRS.spi_miso_oe_n),
.spi_miso_i           (GTP_GRS.spi_miso_i   ),
.spi_miso_o           (GTP_GRS.spi_miso_o   ),
.irq_spi              (GTP_GRS.irq_spi      ),
.spi_wakeup           (GTP_GRS.spi_wakeup_pctl),

.i2c0_scl_i           (GTP_GRS.i2c0_scl_i),
.i2c0_scl_o           (GTP_GRS.i2c0_scl_o),
.i2c0_sda_i           (GTP_GRS.i2c0_sda_i),
.i2c0_sda_o           (GTP_GRS.i2c0_sda_o),
.irq_i2c0             (GTP_GRS.irq_i2c0  ),
.i2c0_wakeup          (GTP_GRS.i2c0_wakeup_pctl),

.i2c1_scl_i           (GTP_GRS.i2c1_scl_i),
.i2c1_scl_o           (GTP_GRS.i2c1_scl_o),
.i2c1_sda_i           (GTP_GRS.i2c1_sda_i),
.i2c1_sda_o           (GTP_GRS.i2c1_sda_o),
.irq_i2c1             (GTP_GRS.irq_i2c1  ),
.i2c1_wakeup          (GTP_GRS.i2c1_wakeup_pctl),

.timer_rstn           (GTP_GRS.timer_rstn ),
.timer_clk            (GTP_GRS.timer_clk  ),
.timer_stamp          (GTP_GRS.timer_stamp),
.timer_pwm            (GTP_GRS.timer_pwm  ),
.irq_timer            (GTP_GRS.irq_timer  )

);

HL55LEFBISTV01  efbist (

.F_Aclk               (F_Aclk        ),
.F_Axa                (F_Axa         ),
.F_Ba                 (),
.F_Bdac               (F_Bdac        ),
.F_Ca                 (F_Ca          ),
.F_Din                (F_Din         ),
.F_Dout               (dout),
.F_Idac               (F_Idac        ),
.F_Itim               (F_Itim        ),
.F_Mode               (F_Mode        ),
.F_Ndac2              (F_Ndac2       ),
.F_Ndac3              (F_Ndac3       ),
.F_Ndace              (F_Ndace       ),
.F_Ndacp              (F_Ndacp       ),
.F_Oe                 (F_Oe          ),
.F_Pa                 (F_Pa          ),
.F_Pd1                (F_Pd1         ),
.F_Pd2                (F_Pd2         ),
.F_Pdace              (F_Pdace       ),
.F_Pdacp              (F_Pdacp       ),
.F_Pe                 (F_Pe          ),
.F_Pnb                (F_Pnb         ),
.F_Pw                 (F_Pw          ),
.F_Ra                 (F_Ra          ),
.F_Rbytesel           (F_Rbytesel    ),
.F_Rdac               (F_Rdac        ),
.F_Reset              (F_Reset       ),
.F_Rmod               (F_Rmod        ),
.F_Seq                (F_Seq         ),
.F_Sleep              (F_Sleep       ),
.F_Slope              (F_Slope       ),
.F_Tm                 (F_Tm          ),
.F_Tm_daa             (F_Tm_daa      ),
.F_Tm_disneg          (F_Tm_disneg   ),
.F_Tm_dispos          (F_Tm_dispos   ),
.F_Tm_disrow          (F_Tm_disrow   ),
.F_Tm_isa             (F_Tm_isa      ),
.F_Tm_itim            (F_Tm_itim     ),
.F_Tm_rdhvpl          (F_Tm_rdhvpl   ),
.F_Tm_reserved        (F_Tm_reserved ),
.F_Tm_vhl             (F_Tm_vhl      ),
.IP_Trim              (),
.F_Turbo              (F_Turbo       ),
.F_Wbytesel           (F_Wbytesel    ),
.F_Wmod               (F_Wmod        ),
.Tck                  (1'b1),
.Tdi                  (1'b1),
.Tdo                  (),
.Ten                  (efb_en        ),
.Toe                  (),
.Trstb                (efb_rstb      ),
.Tstr                 (1'b1),
.U_Aclk               (U_Aclk        ),
.U_Axa                (U_Axa         ),
.U_Ba                 (4'd0),
.U_Bdac               ({1'b0, U_Bdac}),
.U_Ca                 ({1'b0, U_Ca}  ),
.U_Din                (U_Din         ),
.U_Idac               (U_Idac        ),
.U_Itim               (U_Itim        ),
.U_Mode               (U_Mode        ),
.U_Ndac2              (U_Ndac2       ),
.U_Ndac3              (U_Ndac3       ),
.U_Ndace              (U_Ndace       ),
.U_Ndacp              (U_Ndacp       ),
.U_Oe                 (U_Oe          ),
.U_Pa                 ({1'b0, U_Pa}  ),
.U_Pd1                (U_Pd1         ),
.U_Pd2                (U_Pd2         ),
.U_Pdace              (U_Pdace       ),
.U_Pdacp              (U_Pdacp       ),
.U_Pe                 (U_Pe          ),
.U_Pw                 (U_Pw          ),
.U_Ra                 (U_Ra[9:0]),
.U_Rbytesel           (2'b00),
.U_Rdac               (U_Rdac        ),
.U_Reset              (U_Reset       ),
.U_Rmod               (2'b11),
.U_Seq                (U_Seq         ),
.U_Sleep              (U_Sleep       ),
.U_Slope              ({1'b0, U_Slope}),
.U_Trim               (18'd0),
.U_Turbo              (1'b0),
.U_Wbytesel           (2'b00),
.U_Wmod               (2'b11),
.Vgnd                 (1'b0),
.Vpwr                 (1'b1)

);

HL55FGEF21248X32GSA01  eflash (

.Aclk             (F_Aclk        ),
.Pclk             (fpclkg        ),
.Pw               (F_Pw          ),
.Reset            (F_Reset       ),
.Sleep            (F_Sleep       ),
.Itim             (F_Itim        ),
.Idac             (F_Idac        ),
.Slope            (F_Slope[1:0]  ),
.Mode             (F_Mode        ),
.Seq              (F_Seq         ),
.Turbo            (F_Turbo       ),
.Vref             (1'b1),
.Iref             (1'b1),
.Pd1              (F_Pd1         ),
.Pd2              (F_Pd2         ),
.Pe               (F_Pe          ),
.Pdace            (F_Pdace       ),
.Pdacp            (F_Pdacp       ),
.Rdac             (F_Rdac        ),
.Ndace            (F_Ndace       ),
.Ndacp            (F_Ndacp       ),
.Ndac2            (F_Ndac2       ),
.Ndac3            (F_Ndac3       ),
.Bdac             (F_Bdac[2:0]),
.Axa              (F_Axa         ),
.Ra               (F_Ra[8:0]     ),
.Ca               (F_Ca[5:0]     ),
.Wmod             (F_Wmod        ),
.Wbytesel         (F_Wbytesel    ),
.Pa               (F_Pa[5:0]     ),
.Din              (F_Din         ),
.Rmod             (F_Rmod        ),
.Rbytesel         (F_Rbytesel    ),
.Dout             (dout),
.Oe               (1'b1          ),
.Tp               (F_Tp          ),
.Tp_bias          (F_Tp_bias     ),
.Tm               (F_Tm          ),
.Tm_isa           (F_Tm_isa      ),
.Tm_itim          (F_Tm_itim     ),
.Pnb              (F_Pnb         ),
.Tm_rdhvpl        (F_Tm_rdhvpl   ),
.Tm_daa           (F_Tm_daa      ),
.Tm_vhl           (F_Tm_vhl      ),
.Tm_disrow        (F_Tm_disrow   ),
.Tm_dispos        (F_Tm_dispos   ),
.Tm_disneg        (F_Tm_disneg   )

);
endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_DFF_C.v
//
// Functional description: D-type flip-flop with async clear
//
// Parameter description:
//      INIT: init value
//
// Port description:
//      C : asynchronous clear
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_DFF_C
#(
    parameter GRS_EN = "TRUE",
    parameter INIT = 1'b0
) (
    output reg Q,
    input wire D,
    input wire CLK, C
);

    wire grs_n;
    wire grs, RS;

    tri1 grsnet = GRS_INST.GRSNET;
    assign grs_n=(GRS_EN=="TRUE")?grsnet:1'b1;
 
    not (grs, grs_n);
    or (RS, grs, C);

    initial Q = 1'bx;

    always @(posedge CLK or posedge RS) begin
        if (RS)
            Q <= 1'b0;
        else
            Q <= D;
    end

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_MULTACC18.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

//P = MAC + A*B
module GTP_MULTACC18 #(
    parameter GRS_EN              = "TRUE", //"TRUE"; "FALSE"
    parameter SYNC_RST            = "FALSE", //"TRUE"; "FALSE"
    parameter INREG_EN            = "FALSE",  //"TRUE"; "FALSE"
    parameter PIPEREG_EN          = "FALSE",   //"TRUE"; "FALSE"
    parameter ACC_ADDSUB_OP       = 0,
    parameter DYN_ACC_ADDSUB_OP   = 1,     //Select parameter ADDSUB or input ADDSUB
    parameter OVERFLOW_MASK       = 64'h0, //PSIZE = 64 OVERflow setting =  'h8000_0000_0000_00XX , bit width = PSIZE
    parameter PATTERN             = 64'h0, //compare pattern
    parameter MASKPAT             = 64'h0, //mask pattern
    parameter DYN_ACC_INIT        = 0,   //acc init value dynamic input
    parameter ACC_INIT_VALUE      = 64'h0  //acc init value parameter
) (
    output  [63:0] P,
    output  OVER,
    output  UNDER,
    output  EQZ,
    output  EQZM,
    output  EQOM,
    output  EQPAT,
    output  EQPATN,

    input   CE,
    input   RST,
    input   CLK,
    input   [17:0] A,
    input   [17:0] B,
    input   A_SIGNED,
    input   B_SIGNED,
    input   [63:0] ACC_INIT,
    input   ACC_ADDSUB,
    input   RELOAD
);

    wire [63:0] R;

    INT_PREADD_MULTACC #(
        . GRS_EN(GRS_EN),     
        . SYNC_RST(SYNC_RST),   
        . INREG_EN(INREG_EN),   
        . PIPEREG_EN(PIPEREG_EN), 
        . ACCUMADDSUB_OP(ACC_ADDSUB_OP), 
        . DYN_OP_SEL(DYN_ACC_ADDSUB_OP),     
        . ASIZE(18),    
        . BSIZE(18),    
        . PSIZE(64),    
        . PREADD_EN(0),
        . MASK(OVERFLOW_MASK),      
        . DYN_ACC_INIT(DYN_ACC_INIT),
        . ACC_INIT_VALUE(ACC_INIT_VALUE)
    ) U_MACC (
        .CE(CE),
        .RST(RST),
        .CLK(CLK),
        .A(A),
        .B(B),
        .A_SIGNED(A_SIGNED),
        .B_SIGNED(B_SIGNED),
        .C_SIGNED(B_SIGNED),
        .C(18'b0),
        .PREADDSUB(1'b0),
        .ACCUM_INIT(ACC_INIT),
        .ACCUMADDSUB(ACC_ADDSUB),
        .RELOAD(RELOAD),
        .P(P),
        .OVER(OVER),
        .UNDER(UNDER),
        .R(R)     
    );

    INT_FLAG #(
        . GRS_EN(GRS_EN),
        . SYNC_RST(SYNC_RST),
        . PSIZE(64),
        . PATSIZE(64),
        . MASKPATSIZE(64),
        . OUTREG_EN("TRUE")
    ) U_FLAG (
        . CE(CE),
        . RST(RST),
        . CLK(CLK),
        . P(P),
        . PATTERN(PATTERN),
        . MASKPAT(MASKPAT),
        . OVERFLOW_MASK(OVERFLOW_MASK),
        . R(R),
        . eqz(EQZ),
        . eqzm(EQZM),
        . eqom(EQOM),
        . eqpat(EQPAT),
        . eqpatn(EQPATN)
    );

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_DFF_R.v
//
// Functional description: D-type flip-flop with sync clear
//
// Parameter description:
//      INIT: init value
//
// Port description:
//      R: synchronous clear
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_DFF_R
#(
    parameter GRS_EN = "TRUE",
    parameter INIT = 1'b0
) (
    output reg Q,
    input wire D,
    input wire CLK, R
);

    wire grs_n;
    wire RS;

    tri1 grsnet = GRS_INST.GRSNET;
    assign grs_n=(GRS_EN=="TRUE")?grsnet:1'b1;

    not (RS, grs_n);

    initial Q = 1'bx;

    always @(posedge CLK or posedge RS) begin
        if (RS)
            Q <= 1'b0;
        else if (R)
            Q <= 1'b0;
        else
            Q <= D;
    end

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_MUX2LUT7.v
//
// Functional description: 2-to-1 MUX to generate LUT7 func
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_MUX2LUT7
(
    output wire Z,
    input wire I0, I1, S
);

    INT_LUTMUX2_UDP (Z, S, I1, I0);

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2016 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_CLKBUFGMUX_E2.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_CLKBUFGMUX_E2
#(
    parameter TRIGGER_MODE = "NEGEDGE",//"POSEDGE","NEGEDGE"
    parameter INIT_SEL = "CLK0"//"CLK0","CLK1"
) (
    output CLKOUT,
    input CLKIN0,
    input CLKIN1,
    input DETECT_CLK0,
    input DETECT_CLK1,
    input SEL
);

//synthesis translate_off

    initial begin
        if(TRIGGER_MODE != "POSEDGE" && TRIGGER_MODE != "NEGEDGE") begin
            $display("ERROR: The attribute TRIGGER_MODE on instance %m is %s. Legal value are POSEDGE or NEGEDGE.", TRIGGER_MODE);
            $finish;
        end
        if(INIT_SEL != "CLK0" && INIT_SEL != "CLK1") begin
            $display("ERROR: The attribute INIT_SEL on instance %m is %s. Legal value are CLK0 or CLK1.", INIT_SEL);
            $finish;
        end        
    end

///////////////////////////////////////initialization//////////////////////////////////////////////
    reg  clk_out_init_enable;
    
    initial begin
        clk_out_init_enable = 1;
        #0.1 clk_out_init_enable = 0;
    end   

//////////////////////////////////////////////dynamic control/////////////////////////////////////////
    wire clk_detect0_pos;
    wire clk_detect0_neg;
    wire clk_detect1_pos;
    wire clk_detect1_neg;
    wire dis0_rstn;
    wire dis0_setn;
    wire dis1_rstn;
    wire dis1_setn;

    reg clk_detect0_syn_pos;
    reg clk_detect0_syn_neg;
    reg clk_detect1_syn_pos;
    reg clk_detect1_syn_neg;
    reg clk_detect0_syn_pos_temp;
    reg clk_detect0_syn_neg_temp;
    reg clk_detect1_syn_pos_temp;
    reg clk_detect1_syn_neg_temp;
    reg clk_out_syn;
    reg clk_out_asyn;
    reg clk_out;

    initial begin
        if(INIT_SEL == "CLK0") begin
            //#0.1 ;
            clk_detect0_syn_pos <= 1;
            clk_detect0_syn_neg <= 1;
            clk_detect1_syn_pos <= 0;
            clk_detect1_syn_neg <= 0;
            clk_detect0_syn_pos_temp <= 1;
            clk_detect0_syn_neg_temp <= 1;
            clk_detect1_syn_pos_temp <= 0;
            clk_detect1_syn_neg_temp <= 0;
        end
        else begin
            //#0.1 ;
            clk_detect0_syn_pos <= 0;
            clk_detect0_syn_neg <= 0;
            clk_detect1_syn_pos <= 1;
            clk_detect1_syn_neg <= 1;
            clk_detect0_syn_pos_temp <= 0;
            clk_detect0_syn_neg_temp <= 0;
            clk_detect1_syn_pos_temp <= 1;
            clk_detect1_syn_neg_temp <= 1;
        end
    end
    
    assign clk_detect0_pos = (SEL == 0 && clk_detect1_syn_pos == 0) ? 1 : 0;
    assign clk_detect0_neg = (SEL == 0 && clk_detect1_syn_neg == 0) ? 1 : 0;
    assign clk_detect1_pos = (SEL == 1 && clk_detect0_syn_pos == 0) ? 1 : 0;
    assign clk_detect1_neg = (SEL == 1 && clk_detect0_syn_neg == 0) ? 1 : 0;
    assign dis0_rstn  = (DETECT_CLK0 == 1'b0) ? ~SEL : 1'b1;
    assign dis0_setn  = (DETECT_CLK0 == 1'b0) ?  SEL : 1'b1;
    assign dis1_rstn  = (DETECT_CLK1 == 1'b0) ?  SEL : 1'b1;
    assign dis1_setn  = (DETECT_CLK1 == 1'b0) ? ~SEL : 1'b1;

    always @(posedge CLKIN0 or negedge dis0_rstn or negedge dis0_setn) begin
        if(!clk_out_init_enable) begin
            if(!dis0_rstn) begin
                clk_detect0_syn_pos <= 0;
                clk_detect0_syn_pos_temp <= 0;
            end
            else if(!dis0_setn) begin
                clk_detect0_syn_pos <= 1;
                clk_detect0_syn_pos_temp <= 1;
            end
            else begin
                clk_detect0_syn_pos <= clk_detect0_syn_pos_temp;
                clk_detect0_syn_pos_temp <= clk_detect0_pos;
            end
        end
    end    
    
    always @(negedge CLKIN0 or negedge dis0_rstn or negedge dis0_setn) begin
        if(!clk_out_init_enable) begin
            if(!dis0_rstn) begin
                clk_detect0_syn_neg <= 0;
                clk_detect0_syn_neg_temp <= 0;
            end
            else if(!dis0_setn) begin
                clk_detect0_syn_neg <= 1;
                clk_detect0_syn_neg_temp <= 1;
            end
            else begin
                clk_detect0_syn_neg <= clk_detect0_syn_neg_temp;
                clk_detect0_syn_neg_temp <= clk_detect0_neg;
            end
        end
    end    
    
    always @(posedge CLKIN1 or negedge dis1_rstn or negedge dis1_setn) begin
        if(!clk_out_init_enable) begin
            if(!dis1_rstn) begin
                clk_detect1_syn_pos <= 0;
                clk_detect1_syn_pos_temp <= 0;
            end
            else if(!dis1_setn) begin
                clk_detect1_syn_pos <= 1;
                clk_detect1_syn_pos_temp <= 1;
            end
            else begin
                clk_detect1_syn_pos <= clk_detect1_syn_pos_temp;
                clk_detect1_syn_pos_temp <= clk_detect1_pos;
            end
        end
    end    
    
    always @(negedge CLKIN1 or negedge dis1_rstn or negedge dis1_setn) begin
        if(!clk_out_init_enable) begin
            if(!dis1_rstn) begin
                clk_detect1_syn_neg <= 0;
                clk_detect1_syn_neg_temp <= 0;
            end
            else if(!dis1_setn) begin
                clk_detect1_syn_neg <= 1;
                clk_detect1_syn_neg_temp <= 1;
            end 
            else begin
                clk_detect1_syn_neg <= clk_detect1_syn_neg_temp;
                clk_detect1_syn_neg_temp <= clk_detect1_neg;
            end
        end
    end    
    

    always@(*) begin
        if(TRIGGER_MODE == "POSEDGE") begin
            if(clk_detect0_syn_pos && DETECT_CLK0) begin
                clk_out_syn = CLKIN0; 
            end
            else if(clk_detect1_syn_pos && DETECT_CLK1) begin
                clk_out_syn = CLKIN1;
            end
            else begin
                clk_out_syn = 1;
            end
        end
        else begin
            if(clk_detect0_syn_neg && DETECT_CLK0) begin
                clk_out_syn = CLKIN0; 
            end
            else if(clk_detect1_syn_neg && DETECT_CLK1) begin
                clk_out_syn = CLKIN1;
            end
            else begin
                clk_out_syn = 0;
            end
        end
    end

    always@(*) begin
        if(!SEL) begin
            clk_out_asyn = CLKIN0;
        end
        else begin
            clk_out_asyn = CLKIN1;
        end
    end

/////////////////////////////output///////////////////////////////////

    assign CLKOUT = clk_out;

    always@(*)begin
        if(clk_out_init_enable) begin
            if(INIT_SEL == "CLK1") begin
                clk_out = CLKIN1;
            end
            else if(INIT_SEL == "CLK0")begin
                clk_out = CLKIN0;
            end
        end
        else begin
            if(DETECT_CLK0 || DETECT_CLK1) begin
                clk_out = clk_out_syn;
            end
            else begin
                clk_out = clk_out_asyn;
            end
        end
    end

//synthesis translate_on

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_OUTBUFCO.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_OUTBUFCO #(
    parameter IOSTANDARD = "DEFAULT"
)(
    output O,
    output OB,
    input I
) /* synthesis syn_black_box */ ;
  
  initial begin
    case (IOSTANDARD)
    "SSTL18D_I", "SSTL18D_II", "SSTL15D_I", "SSTL15D_II", "HSTL15D_I", "SSTL25D_I", "SSTL25D_II", "SSTL15D_I_CAL", "SSTL15D_II_CAL", "HSTL15D_I_CAL","LVPECL",
    "LVCMOS25D", "LVCMOS33D", "RSDS", "PPDS","BLVDS", "LVDS25E", "DEFAULT" :;
    default : begin
           $display("Attribute Syntax Error : The attribute IOSTANDARD on GTP_OUTBUFCO instance %m is set to %s.", IOSTANDARD);
           $finish;
              end
    endcase
    end 

    buf (O, I);
    not (OB, I);

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_MULTADDSUM9.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

//P = (A0*B0 +/- A1*B1) +- (A2*B2 +/- A3*B3)
module GTP_MULTADDSUM9  #(
    parameter GRS_EN            = "TRUE", //"TRUE"; "FALSE"
    parameter SYNC_RST          = "FALSE", //"TRUE"; "FALSE"
    parameter INREG_EN          = "FALSE",  //"TRUE"; "FALSE"
    parameter PIPEREG_EN        = "FALSE",  //"TRUE"; "FALSE"
    parameter OUTREG_EN         = "FALSE",   //"TRUE"; "FALSE"
    parameter ADDSUB_OP         = 2'b00 ,
    parameter SUM_ADDSUB_OP     = 0 ,
    parameter DYN_ADDSUB_OP     = 2'b11,
    parameter DYN_SUM_ADDSUB_OP = 1
)(
    output  [20-1:0] P,
    input   CE,
    input   RST,
    input   CLK,
    input   [1:0] A_SIGNED,
    input   [9-1:0] A0,
    input   [9-1:0] A1,
    input   [9-1:0] A2,
    input   [9-1:0] A3,
    input   [1:0] B_SIGNED,
    input   [9-1:0] B0,
    input   [9-1:0] B1,
    input   [9-1:0] B2,
    input   [9-1:0] B3,
    input   [1:0] ADDSUB,
    input   SUM_ADDSUB
);

    INT_MULTADDSUM #(
        . GRS_EN(GRS_EN),    
        . SYNC_RST(SYNC_RST),  
        . INREG_EN(INREG_EN),  
        . PIPEREG_EN(PIPEREG_EN),
        . OUTREG_EN(OUTREG_EN), 
        . ADDSUB_OP01(ADDSUB_OP[0]),  
        . ADDSUB_OP23(ADDSUB_OP[1]),  
        . ADDSUBSUM_OP(SUM_ADDSUB_OP), 
        . DYN_OP_SEL0(DYN_ADDSUB_OP[0]),
        . DYN_OP_SEL1(DYN_ADDSUB_OP[1]),
        . DYN_OP_SEL2(DYN_SUM_ADDSUB_OP),
        . ASIZE(9),
        . BSIZE(9)
    ) U_INT_MULTADDSUM (
        . CE(CE),
        . RST(RST),
        . CLK(CLK),
        . A_SIGNED01(A_SIGNED[0]),
        . A_SIGNED23(A_SIGNED[1]),
        . A0(A0),
        . A1(A1),
        . A2(A2),
        . A3(A3),
        . B_SIGNED01(B_SIGNED[0]),
        . B_SIGNED23(B_SIGNED[1]), 
        . B0(B0),
        . B1(B1),
        . B2(B2),
        . B3(B3),
        . ADDSUB01(ADDSUB[0]),
        . ADDSUB23(ADDSUB[1]),
        . ADDSUBSUM(SUM_ADDSUB),
        . P(P)
    );               


endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////

//P = MAC + (A*(B+C))
`timescale 1 ns / 1 ps

module INT_PREADD_MULTACC
#(
    parameter GRS_EN      = "FALSE", //"TRUE"; "FALSE"
    parameter SYNC_RST    = "FALSE", //"TRUE"; "FALSE"
    parameter INREG_EN    = "FALSE",  //"TRUE"; "FALSE"
    parameter PREREG_EN   = "FALSE",  //"TRUE"; "FALSE"
    parameter PIPEREG_EN  = "FALSE",   //"TRUE"; "FALSE"
    parameter ACCUMADDSUB_OP = 0,
    parameter DYN_OP_SEL  = 1,     //Select parameter ADDSUB or input ADDSUB
    parameter integer ASIZE = 9,   // LEGAL ASIZE = 9,18,27,36
    parameter integer BSIZE = 8,   //LEGAL BSIZE = 8,18,26,18
    parameter integer PSIZE = 32,  // LEGAL PSIZE for 9x9 = 32;
                                   // LEGAL PSIZE for other mode = 64
    parameter [PSIZE-1:0] MASK = 'h0,   //PSIZE = 64 OVERflow setting= 'h8000_0000_0000_0000, bit width = PSIZE
    parameter DYN_ACC_INIT   = 0,   //acc init value dynamic input
    parameter [PSIZE-1:0] ACC_INIT_VALUE = 'b0, //acc init value parameter
    parameter [ASIZE-2:0] SC_PSE_A = 'b0, //SC_PSE = 0, disable PSE,  bit width = ASIZE-1
    parameter [BSIZE-2:0] SC_PSE_B = 'b0, //SC_PSE = 0, disable PSE,  bit width = BSIZE-1
    parameter [BSIZE-2:0] SC_PSE_C = 'b0, //SC_PSE = 0, disable PSE,  bit width = BSIZE-1
    parameter integer PREADD_EN = 1
) (
    input   CE,
    input   RST,
    input   CLK,
    input   [ASIZE-1:0] A,
    input   [BSIZE-1:0] B,
    input   A_SIGNED,
    input   B_SIGNED,
    input   C_SIGNED,
    input   [BSIZE-1:0] C,
    input   PREADDSUB,
    input   [PSIZE-1:0] ACCUM_INIT,
    input   ACCUMADDSUB,
    input   RELOAD,
    output  [PSIZE-1:0] P,
    output  reg OVER,
    output  reg UNDER,
    output  [PSIZE-1:0] R
);

initial begin
    if ((PREADD_EN != 0) && (PREADD_EN != 1))
    begin
        $finish;
    end
    case (ASIZE)
        9:  if ((BSIZE + PREADD_EN) != 9 || PSIZE != 32)
            begin
                $finish;
            end
        18, 36: if (BSIZE != 18 || PSIZE != 64)
            begin
                $finish;
            end
        27: if ((BSIZE + PREADD_EN) != 27 || PSIZE != 64)
            begin
                $finish;
            end
        default :
            $finish;
    endcase
    //$display (" INT_PREADD_MULTACC error :illegal ASIZE or BSIZE or PSIZE");

    if ((GRS_EN != "TRUE") && (GRS_EN != "FALSE")) begin
        $display("GRS_EN error");
        $finish;
    end
    if ((SYNC_RST != "TRUE") && (SYNC_RST != "FALSE")) begin
        $display("SYNC_RST error");
        $finish;
    end

    if ((INREG_EN != "TRUE") && (INREG_EN != "FALSE")) begin
        $display("INREG_EN error");
        $finish;
    end
    if ((PREREG_EN != "TRUE") && (PREREG_EN != "FALSE")) begin
        $display("PREREG_EN error");
        $finish;
    end
    if ((PIPEREG_EN != "TRUE") && (PIPEREG_EN != "FALSE")) begin
        $display("PIPEREG_EN error");
        $finish;
    end
end    

localparam Psize = ASIZE + BSIZE + PREADD_EN;
localparam BIT_EXT = PSIZE - Psize;

wire [ASIZE-1:0] A_PSE;
wire [BSIZE-1:0] B_PSE;
wire [BSIZE-1:0] C_PSE;

reg  [ASIZE-1:0] a_ireg;
reg  [BSIZE-1:0] b_ireg;
reg  [BSIZE-1:0] c_ireg;
reg  asign_ireg, bsign_ireg, csign_ireg;
reg  preaddsub_ireg;
reg  [PSIZE-1:0] acc_init_ireg;
reg  reload_ireg, acc_addsub_ireg;
reg  reload_preg, acc_addsub_preg;

wire [ASIZE-1:0] a_in;
wire [BSIZE-1:0] b_in;
wire [BSIZE-1:0] c_in;
wire asign_in, bsign_in, csign_in;
wire preaddsub_in;
wire [PSIZE-1:0] acc_init_value;
wire [PSIZE-1:0] acc_init_in;
wire reload_in, acc_addsub_in;
wire reload_real, acc_addsub_real;

wire [BSIZE:0] b2prad;
wire [BSIZE:0] c2prad;
wire [BSIZE:0] prad_sum;
wire [BSIZE:0] b_inmux;
wire prad_sign, bsign_inmux;

reg  [ASIZE-1:0] a_pareg;
reg  [BSIZE:0]   b_pareg;
reg  asign_pareg, bsign_pareg;

wire [ASIZE-1:0] a_mult;
wire [BSIZE:0]   b_mult;
wire asign_mult, bsign_mult;

wire [Psize-1:0] a_mext;
wire [Psize-1:0] b_mext;
wire [Psize-1:0] PRODUCT;
wire         PSIGN1; 

reg  [PSIZE-1:0] PRODUCT_reg;
wire [PSIZE-1:0] PRODUCT_out;

reg  [PSIZE-1:0] DPO_reg;
wire global_rstn, RST_sync, RST_async, rst_asyncomb;

assign global_rstn = GRS_EN == "TRUE" ? GRS_INST.GRSNET : 1'b1;
assign RST_sync = (SYNC_RST == "TRUE") ? RST : 1'b0;
assign RST_async = (SYNC_RST == "FALSE") ? RST : 1'b0;
assign rst_asyncomb = RST_async | (~global_rstn);

assign acc_init_value = DYN_ACC_INIT ? ACCUM_INIT : ACC_INIT_VALUE;

INT_PSE #(.ASIZE(ASIZE), .SC_PSE(SC_PSE_A)) U1_PSE (.A(A), .SIGN(A_SIGNED), .A_PSE(A_PSE));
INT_PSE #(.ASIZE(BSIZE), .SC_PSE(SC_PSE_B)) U2_PSE (.A(B), .SIGN(B_SIGNED), .A_PSE(B_PSE));
INT_PSE #(.ASIZE(BSIZE), .SC_PSE(SC_PSE_C)) U3_PSE (.A(C), .SIGN(C_SIGNED), .A_PSE(C_PSE));

initial begin
    {asign_ireg, a_ireg} = 'b0;
    {bsign_ireg, b_ireg} = 'b0;
    {csign_ireg, c_ireg} = 'b0;
     preaddsub_ireg = 'b0;
     acc_init_ireg  = 'b0;
     reload_ireg    = 'b0;
     acc_addsub_ireg = 'b0;
     PRODUCT_reg = 'b0;
     DPO_reg    = 'b0;
end
always @(posedge CLK or posedge rst_asyncomb)
    if (rst_asyncomb || RST_sync) begin
        {asign_ireg, a_ireg} <= 'b0;
        {bsign_ireg, b_ireg} <= 'b0;
        {csign_ireg, c_ireg} <= 'b0;
         preaddsub_ireg   <= 'b0;
         acc_init_ireg    <= 'b0;
         reload_ireg      <= 'b0;
         acc_addsub_ireg  <= 'b0;
    end
    else if (CE) begin
        {asign_ireg, a_ireg} <= {A_SIGNED, A_PSE};
        {bsign_ireg, b_ireg} <= {B_SIGNED, B_PSE};
        {csign_ireg, c_ireg} <= {C_SIGNED, C_PSE};
         preaddsub_ireg   <= PREADDSUB;
         acc_init_ireg    <= acc_init_value;
         reload_ireg      <= RELOAD;
         acc_addsub_ireg  <= (DYN_OP_SEL == 1'b1)?ACCUMADDSUB :ACCUMADDSUB_OP;
    end

assign {asign_in, a_in} = (INREG_EN == "TRUE") ? {asign_ireg, a_ireg} : {A_SIGNED, A_PSE};
assign {bsign_in, b_in} = (INREG_EN == "TRUE") ? {bsign_ireg, b_ireg} : {B_SIGNED, B_PSE};
assign {csign_in, c_in} = (INREG_EN == "TRUE") ? {csign_ireg, c_ireg} : {C_SIGNED, C_PSE};
assign  preaddsub_in    = (INREG_EN == "TRUE") ?  preaddsub_ireg      :  PREADDSUB;

assign b2prad = {(bsign_in & b_in[BSIZE-1]), b_in};
assign c2prad = {(csign_in & c_in[BSIZE-1]), c_in};
assign prad_sum  = preaddsub_in ? (b2prad - c2prad) : (b2prad + c2prad);
assign prad_sign = bsign_in | csign_in;


reg preadd_over_flag;
always @(*)begin
  if(preaddsub_in==1'b0 && PREADD_EN==1)begin
    if((bsign_in==1'b1 && b_in[BSIZE-1]==1'b0 && csign_in==1'b0 && prad_sum[BSIZE]==1'b1) || (bsign_in==1'b0 && csign_in==1'b1 && c_in[BSIZE-1]==1'b0 && prad_sum[BSIZE]==1'b1))begin
      preadd_over_flag = 1'b1;
    end
    else begin
      preadd_over_flag = 1'b0;
    end
  end
  else if(preaddsub_in==1'b1 && PREADD_EN==1)begin
    if((bsign_in==1'b1 && b_in[BSIZE-1]==1'b1 && csign_in==1'b0 && prad_sum[BSIZE]==1'b0) || (bsign_in==1'b0 && csign_in==1'b1 && c_in[BSIZE-1]==1'b1 && prad_sum[BSIZE]==1'b1) ||
      (bsign_in ==1'b0 && csign_in==1'b0 && (b_in<c_in)))begin
      preadd_over_flag = 1'b1;
    end
    else begin
      preadd_over_flag = 1'b0;
    end
  end
end

always @(preadd_over_flag) begin
    if (preadd_over_flag==1 && PREADD_EN==1)
    $display("Error: PREADD result is overflow!");
end

always @(*) begin
    if (PREADD_EN && (BSIZE == 26) && (prad_sign == 1'b0))
        if ((preaddsub_in == 1'b1) && (prad_sum[BSIZE] == 1'b1)) begin
            $display("PG30-ERROR: Unexpected function mismatch.");
        end
end

assign acc_init_in   = (INREG_EN == "TRUE") ? acc_init_ireg   : acc_init_value;
assign reload_in     = (INREG_EN == "TRUE") ? reload_ireg     : RELOAD;
assign acc_addsub_in = (INREG_EN == "TRUE") ? acc_addsub_ireg :(DYN_OP_SEL == 1'b1)?ACCUMADDSUB :ACCUMADDSUB_OP; 

assign b_inmux     = PREADD_EN ? prad_sum : {1'b0, b_in};
assign bsign_inmux = PREADD_EN ? prad_sign : bsign_in;
always @(posedge CLK or posedge rst_asyncomb)
    if (rst_asyncomb || RST_sync) begin
        {asign_pareg, a_pareg} <= 'b0;
        {bsign_pareg, b_pareg} <= 'b0;
    end
    else if (CE) begin
        {asign_pareg, a_pareg} <= {asign_in, a_in};
        {bsign_pareg, b_pareg} <= {bsign_inmux, b_inmux};
    end

assign {asign_mult, a_mult} = (PREREG_EN == "TRUE") ? {asign_pareg, a_pareg} : {asign_in, a_in};
assign {bsign_mult, b_mult} = (PREREG_EN == "TRUE") ? {bsign_pareg, b_pareg} : {bsign_inmux, b_inmux};

assign a_mext = {{(Psize-ASIZE){asign_mult & a_mult[ASIZE-1]}}, a_mult};
assign b_mext = {{(Psize-BSIZE-PREADD_EN){bsign_mult & b_mult[BSIZE+PREADD_EN-1]}}, b_mult[BSIZE+PREADD_EN-1:0]};
assign PRODUCT = a_mext * b_mext;
assign PSIGN1  = asign_mult | bsign_mult;

always @(posedge CLK or posedge rst_asyncomb)
    if (rst_asyncomb || RST_sync) begin
        PRODUCT_reg <= 0;
        reload_preg <= 0;
        acc_addsub_preg <= 0;
    end
    else if (CE) begin
        PRODUCT_reg <= {{(PSIZE-Psize){PSIGN1&PRODUCT[Psize-1]}},PRODUCT};
        reload_preg <= reload_in;
        acc_addsub_preg <= acc_addsub_in;
    end

assign reload_real = (PIPEREG_EN == "TRUE") ? reload_preg : reload_in; 
assign acc_addsub_real = (PIPEREG_EN == "TRUE") ? acc_addsub_preg : acc_addsub_in; 
assign PRODUCT_out = (PIPEREG_EN == "TRUE") ? PRODUCT_reg : {{(PSIZE-Psize){PSIGN1&PRODUCT[Psize-1]}},PRODUCT};

assign R = reload_real ? acc_init_in
                     : (acc_addsub_real? DPO_reg - PRODUCT_out : DPO_reg + PRODUCT_out);

always @(posedge CLK or posedge rst_asyncomb)
    if (rst_asyncomb || RST_sync) begin
        DPO_reg <= 'b0;
    end
    else if (CE) begin
        DPO_reg <= R;
    end
   
assign P =  DPO_reg;

wire eqzero;
wire eqone;
reg eqzero_d;
reg eqone_d;
wire eqzero_one;
wire over;
wire under;

assign eqzero = &(~R | MASK);
assign eqone  = &( R | MASK);
assign eqzero_one = ~(eqzero|eqone);

always @ (posedge CLK or posedge rst_asyncomb)
    if (rst_asyncomb || RST_sync) begin
        eqzero_d  <= 0;
        eqone_d   <= 0;
        OVER      <= 0;
        UNDER     <= 0;
    end
    else if (CE) begin
        eqzero_d  <= eqzero;
        eqone_d   <= eqone;
        OVER      <= over;
        UNDER     <= under;
    end

assign over = eqzero_d & eqzero_one;
assign under = eqone_d & eqzero_one;

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_IGDES10.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_IGDES10 #(
parameter GRS_EN = "TRUE", //"TRUE"; "FALSE"
parameter LRS_EN = "TRUE",  //"TRUE"; "FALSE"
parameter DPI_EN = "FALSE"  //"TRUE"; "FALSE"
)(
output [9:0] Q,
output [1:0] DPI_STS,
input [1:0] DPI_CTRL,
input DPI_STS_CLR_N,
input PADI,
input DESCLK,
input RCLK,
input RST
);

//synthesis translate_off
wire [7:0] PADI_D;
reg DPI_P;
reg [1:0] DPI_STS_R;
reg DPI_N_reg;
wire COMP_BEFORE;
wire COMP_AFTER;
wire COMP_BEFORE_D;
wire COMP_AFTER_D;
wire PD_BEFORE;
wire PD_AFTER;
wire DPI_BEFORE_POS_REG_T;
wire DPI_AFTER_POS_REG_T;
wire DPI_BEFORE_NEG_REG_T;
wire DPI_AFTER_NEG_REG_T;
wire AFTER_POS;
wire BEFORE_POS;
wire AFTER_NEG;
wire BEFORE_NEG;
reg DPI_BEFORE;
reg DPI_AFTER;
reg DPI_BEFORE_POS_REG;
reg DPI_BEFORE_NEG_REG;
reg DPI_AFTER_POS_REG;
reg DPI_AFTER_NEG_REG;
reg [9:0] shift_reg;
reg [9:0] capture_reg;
reg [2:0] cnt;
wire capture_en;
reg [9:0] Q_reg;

initial begin
DPI_P        = 0;
DPI_STS_R    = 0;
DPI_N_reg    = 0;
DPI_BEFORE   = 0;
DPI_AFTER    = 0;
DPI_BEFORE_POS_REG = 0;
DPI_BEFORE_NEG_REG = 0;
DPI_AFTER_POS_REG  = 0;
DPI_AFTER_NEG_REG  = 0;
shift_reg   = 0;
capture_reg = 0;
cnt         = 0;
Q_reg       = 0;  
end
assign global_rstn = (GRS_EN == "TRUE") ? GRS_INST.GRSNET : 1'b1;
assign lsr_rstn = LRS_EN == "TRUE" ? (~RST) : 1'b1;


assign  #0.05 PADI_D[0] =  PADI;
assign  #0.05 PADI_D[1] =  PADI_D[0];
assign  #0.05 PADI_D[2] =  PADI_D[1];
assign  #0.05 PADI_D[3] =  PADI_D[2];
assign  #0.05 PADI_D[4] =  PADI_D[3];
assign  #0.05 PADI_D[5] =  PADI_D[4];
assign  #0.05 PADI_D[6] =  PADI_D[5];
assign  #0.05 PADI_D[7] =  PADI_D[6];

assign PADI_SAMPLE = (DPI_EN == "TRUE") ? PADI_D[3] : PADI;

always @(posedge DESCLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_P <= 0;
   else if (!lsr_rstn)
      DPI_P <= 0;
   else
      DPI_P <= PADI_SAMPLE;
end

always @(negedge DESCLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_N_reg <= 0;
   else if (!lsr_rstn)
      DPI_N_reg <= 0;
   else 
      DPI_N_reg <= PADI_SAMPLE;
end

always @(*) begin
   case (DPI_CTRL[1:0])
      2'd0:    begin DPI_BEFORE = PADI_D[2];  DPI_AFTER = PADI_D[4]; end
      2'd1:    begin DPI_BEFORE = PADI_D[1];  DPI_AFTER = PADI_D[5]; end
      2'd2:    begin DPI_BEFORE = PADI_D[0];  DPI_AFTER = PADI_D[6]; end
      default: begin DPI_BEFORE = PADI;       DPI_AFTER = PADI_D[7]; end
   endcase
end

always @(posedge DESCLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_BEFORE_POS_REG <= 0;
   else if (!lsr_rstn)
      DPI_BEFORE_POS_REG <= 0;
   else   
      DPI_BEFORE_POS_REG <= DPI_BEFORE;
end

always @(negedge DESCLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_BEFORE_NEG_REG <= 0;
   else if (!lsr_rstn)
      DPI_BEFORE_NEG_REG <= 0;
   else     
      DPI_BEFORE_NEG_REG <= DPI_BEFORE;
end


always @(posedge DESCLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_AFTER_POS_REG <= 0;
   else if (!lsr_rstn)
      DPI_AFTER_POS_REG <= 0;
   else   
      DPI_AFTER_POS_REG <= DPI_AFTER;
end


always @(negedge DESCLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_AFTER_NEG_REG <= 0;
   else if (!lsr_rstn)
      DPI_AFTER_NEG_REG <= 0;
   else     
      DPI_AFTER_NEG_REG <= DPI_AFTER;
end


assign BEFORE_POS = DPI_BEFORE_POS_REG_T ^ DPI_P;
assign DPI_BEFORE_POS_REG_T = (DPI_EN == "TRUE") ? DPI_BEFORE_POS_REG : 0;

assign AFTER_POS = DPI_AFTER_POS_REG_T ^ DPI_P;
assign DPI_AFTER_POS_REG_T = (DPI_EN == "TRUE") ? DPI_AFTER_POS_REG : 0;

assign BEFORE_NEG = DPI_BEFORE_NEG_REG_T ^ DPI_N_reg;
assign DPI_BEFORE_NEG_REG_T = (DPI_EN == "TRUE") ? DPI_BEFORE_NEG_REG : 0;

assign AFTER_NEG = DPI_AFTER_NEG_REG_T ^ DPI_N_reg;
assign DPI_AFTER_NEG_REG_T = (DPI_EN == "TRUE") ? DPI_AFTER_NEG_REG : 0;


assign COMP_BEFORE = BEFORE_POS || BEFORE_NEG;
assign COMP_AFTER = AFTER_POS || AFTER_NEG;

assign #0.1 COMP_BEFORE_D = COMP_BEFORE;
assign #0.1 COMP_AFTER_D = COMP_AFTER;

assign PD_BEFORE = COMP_BEFORE && COMP_BEFORE_D;
assign PD_AFTER = COMP_AFTER && COMP_AFTER_D;


always @(posedge DPI_STS_CLR_N or negedge global_rstn or negedge lsr_rstn or posedge PD_BEFORE) begin
   if (!global_rstn)
      DPI_STS_R[0] <= 0;
   else if (!lsr_rstn)
      DPI_STS_R[0] <= 0;
   else if (PD_BEFORE)     
      DPI_STS_R[0] <= 1'b1;
   else
      DPI_STS_R[0] <= 1'b0;
end

always @(posedge DPI_STS_CLR_N or negedge global_rstn or negedge lsr_rstn or posedge PD_AFTER) begin
   if (!global_rstn)
      DPI_STS_R[1] <= 0;
   else if (!lsr_rstn)
      DPI_STS_R[1] <= 0;
   else if (PD_AFTER)     
      DPI_STS_R[1] <= 1'b1;
   else
      DPI_STS_R[1] <= 1'b0;
end

assign DPI_STS[0] = DPI_STS_R[0];
assign DPI_STS[1] = DPI_STS_R[1];

always @(posedge DESCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      shift_reg <= 0;
   else if (!lsr_rstn)
      shift_reg <= 0;
   else
      shift_reg <= {DPI_N_reg, DPI_P, shift_reg[9:2]};

always @(posedge DESCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      cnt <= 0;
   else if (!lsr_rstn)
      cnt <= 0;
   else if (cnt == 4)
      cnt <= 0;
   else   
      cnt <= cnt + 1;

assign capture_en = cnt == 4;

always @(posedge DESCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      capture_reg <= 0;
   else if (!lsr_rstn)
      capture_reg <= 0;
   else if (capture_en)
      capture_reg <= shift_reg;
      
always @(posedge RCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      Q_reg <= 0;
   else if (!lsr_rstn)
      Q_reg <= 0;
   else
      Q_reg <= capture_reg;      

assign Q = Q_reg;

//synthesis translate_on

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2016 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_LUT6CARRY.v
//
// Functional description: LUT6 and CARRY
//
// Parameter description:
//      I5_TO_CARRY : 'TRUE'  I5    to Carry-mux(I0)
//                    'FALSE' LUT5B to Carry-mux(I0)
//      I5_TO_LUT   : 'TRUE'  I5  to muxL6.Sel
//                    'FALSE' CIN to muxL6.Sel
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_LUT6CARRY
#(
    parameter [63:0] INIT = 64'h0000_0000_0000_0000,
    parameter I5_TO_CARRY = "TRUE",
    parameter I5_TO_LUT = "FALSE"
) (
    output COUT, 
    output Z,
    input CIN, 
    input I0,
    input I1,
    input I2,
    input I3,
    input I4,
    input I5
);

    initial
    begin
        if (I5_TO_LUT != "TRUE" && I5_TO_LUT != "FALSE")
        begin
            $display("ERROR: The attribute I5_TO_LUT on instance %m is %s. Legal values are TRUE or FALSE.", I5_TO_LUT);
            $finish;
        end

        if (I5_TO_CARRY != "TRUE" && I5_TO_CARRY != "FALSE")
        begin
            $display("ERROR: The attribute I5_TO_CARRY on instance %m is %s. Legal values are TRUE or FALSE.", I5_TO_CARRY);
            $finish;
        end
    end

    wire c0_int;
    wire i5_int;
    wire z5a, z5b;

    assign c0_int = (I5_TO_CARRY == "TRUE") ? I5 : z5b;
    assign i5_int = (I5_TO_LUT == "FALSE") ? CIN : I5;

    GTP_LUT5 #(.INIT(INIT[31:0]))
        l5a (.I0(I0), .I1(I1), .I2(I2), .I3(I3), .I4(I4), .Z(z5a));

    GTP_LUT5 #(.INIT(INIT[63:32]))
        l5b (.I0(I0), .I1(I1), .I2(I2), .I3(I3), .I4(I4), .Z(z5b));

    INT_LUTMUX2_UDP (Z,    i5_int, z5b, z5a);
    INT_LUTMUX2_UDP (COUT, z5a,    CIN, c0_int);

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_MULTADDACC9.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

//P = MAC + (A0*B0 + A1*B1)
module GTP_MULTADDACC9 #(
    parameter  GRS_EN             = "TRUE", //"TRUE"; "FALSE"
    parameter  SYNC_RST           = "FALSE", //"TRUE"; "FALSE"
    parameter  INREG_EN           = "FALSE",  //"TRUE"; "FALSE"
    parameter  PIPEREG_EN         = "FALSE",//"TRUE"; "FALSE"
    parameter  ADDSUB_OP          = 0 ,
    parameter  ACC_ADDSUB_OP      = 0,
    parameter  DYN_ADDSUB_OP      = 1,
    parameter  DYN_ACC_ADDSUB_OP  = 1,
    parameter  OVERFLOW_MASK      = 32'h0, //PSZIE = 32 OVERflow setting = 'h1_0000_0000, bit width = PSIZE
    parameter  PATTERN            = 32'h0, //compare pattern
    parameter  MASKPAT            = 32'h0, //pattern mask
    parameter  DYN_ACC_INIT       = 0,     //acc init value dynamic input
    parameter  ACC_INIT_VALUE     = 32'h0  //acc init value parameter
) (
    output  [31:0] P,
    output  OVER,
    output  UNDER,
    output  EQZ,
    output  EQZM,
    output  EQOM,
    output  EQPAT,
    output  EQPATN,

    input   CE,
    input   RST,
    input   CLK,
    input   A_SIGNED,
    input   [8:0] A0,
    input   [8:0] A1,
    input   B_SIGNED,
    input   [8:0] B0,
    input   [8:0] B1,
    input   [31:0] ACC_INIT,
    input   ADDSUB,
    input   ACC_ADDSUB,
    input   RELOAD
);

    wire [31:0] R;

    INT_PREADD_MULTADDACC #(
        . GRS_EN(GRS_EN),     
        . SYNC_RST(SYNC_RST),   
        . INREG_EN(INREG_EN),   
        . PIPEREG_EN(PIPEREG_EN), 
        . ADDSUB_OP(ADDSUB_OP),    
        . ACCUMADDSUB_OP(ACC_ADDSUB_OP),
        . DYN_OP_ADDSUB(DYN_ADDSUB_OP),   
        . DYN_OP_ACC(DYN_ACC_ADDSUB_OP),  
        . ASIZE(9), 
        . BSIZE(9), 
        . PSIZE(32), 
        . PREADD_EN(0),
        . MASK(OVERFLOW_MASK), 
        . DYN_ACC_INIT(DYN_ACC_INIT),
        . ACC_INIT_VALUE(ACC_INIT_VALUE)
    ) U_MACC (
        . CE(CE),
        . RST(RST),
        . CLK(CLK),
        . A_SIGNED(A_SIGNED),
        . A0(A0),
        . A1(A1),
        . B_SIGNED(B_SIGNED),
        . B0(B0),
        . B1(B1),
        . C_SIGNED(B_SIGNED),
        . C0(9'b0),
        . C1(9'b0),
        . PREADDSUB(2'b0),
        . ACCUM_INIT(ACC_INIT),
        . ADDSUB(ADDSUB),
        . ACCUMADDSUB(ACC_ADDSUB),
        . RELOAD(RELOAD),
        . P(P),
        . OVER(OVER),
        . UNDER(UNDER),
        . R(R) 
    );

    INT_FLAG #(
        . GRS_EN(GRS_EN),
        . SYNC_RST(SYNC_RST),
        . PSIZE(32),
        . PATSIZE(32),
        . MASKPATSIZE(32),
        . OUTREG_EN("TRUE")
    ) U_FLAG (
        . CE(CE),
        . RST(RST),
        . CLK(CLK),
        . P(P),
        . PATTERN(PATTERN),
        . MASKPAT(MASKPAT),
        . OVERFLOW_MASK(OVERFLOW_MASK),
        . R(R),
        . eqz(EQZ),
        . eqzm(EQZM),
        . eqom(EQOM),
        . eqpat(EQPAT),
        . eqpatn(EQPATN)
    );

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_DFF_CE.v
//
// Functional description: D-type flip-flop with async clear and enable
//
// Parameter description:
//      INIT: init value
//
// Port description:
//      C : asynchronous clear
//      CE   : enable
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_DFF_CE
#(
    parameter GRS_EN = "TRUE",
    parameter INIT = 1'b0
) (
    output reg Q,
    input wire D,
    input wire CLK, C, CE
);

    wire grs_n;
    wire grs, RS;

    tri1 grsnet = GRS_INST.GRSNET;
    assign grs_n=(GRS_EN=="TRUE")?grsnet:1'b1;

    not (grs, grs_n);
    or (RS, grs, C);

    initial Q = 1'bx;

    always @(posedge CLK or posedge RS) begin
        if (RS)
            Q <= 1'b0;
        else if (CE)
            Q <= D;
    end

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_IOBUFEDS.v
//
// Functional description: Differential Signaling Input/Output Buffer
//
// Parameter description:
//
// Port description:
//
// Revision:
//    06/18/14 - Initial version.
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_IOBUFEDS #(
    parameter IOSTANDARD = "DEFAULT",
    parameter TERM_DIFF = "ON"
)(
    output reg O,
    inout IO,
    inout IOB,
    input I,
    input EN,                    // 1: enable inbuf, normal mode; 0: disable inbuf, standby mode.
    input T
) /* synthesis syn_black_box */ ;
  
  initial begin
    case (IOSTANDARD)
    "LVDS", "MINI-LVDS", "SUB-LVDS", "TMDS", "DEFAULT" :;
    default : begin
           $display("Attribute Syntax Error : The attribute IOSTANDARD on GTP_IOBUFEDS instance %m is set to %s.", IOSTANDARD);
           $finish;
              end
    endcase

    case (TERM_DIFF)
    "ON", "OFF" :;
    default : begin
           $display("Attribute Syntax Error : The attribute TERM_DIFF on GTP_IOBUFEDS instance %m is set to %s.", TERM_DIFF);
           $finish;
              end
    endcase
    end


    bufif0 (IO, I, T);
    notif0 (IOB, I, T);

  always @(*)
    begin
      if (EN == 1'b1)
        begin
        if (IO == 1'b1 && IOB == 1'b0)
            O = IO;
        else if (IO == 1'b0 && IOB == 1'b1)
            O = IO;
        else
            O = 1'bx;
        end
     else
            O = 1'b1;
    end

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_CLKBUFG.v
//
// Functional description: Global Clock Buffer
//
// Parameter description:
//
// Port description:
//
// Revision:
//    06/18/14 - Initial version.
//    05/11/14 - 
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_CLKBUFG
(
    output CLKOUT,
    input CLKIN
);

    assign CLKOUT = CLKIN;

endmodule




 //////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2016 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library:
// Filename: GTP_DDRPHY.v
//
// Functional description:DDR_PHY
//
// Parameter description:
//
// Port description:
//
// Revision:1.0(initial)
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1ns/1ps

module GTP_DDRPHY #(   
    parameter     [31:0]      TEST_PATTERN2             =32'h0000_0000,								
    parameter     [31:0]      TEST_PATTERN3             =32'h0000_0000,
    parameter     integer     T200US                    =54000,        //0~131071
    parameter     [15:0]      MR0_DDR3                  =16'h1108,
    parameter     [15:0]      MR1_DDR3                  =16'h0001,
    parameter     [15:0]      MR2_DDR3                  =16'h0000,
    parameter     [15:0]      MR3_DDR3                  =16'h0000,
    parameter     [15:0]      MR_DDR2                   =16'h0100,
    parameter     [15:0]      EMR1_DDR2                 =16'h0401,
    parameter     [15:0]      EMR2_DDR2                 =16'h0000,
    parameter     [15:0]      EMR3_DDR2                 =16'h0000,
    parameter     [15:0]      MR_LPDDR                  =16'h0003,
    parameter     [15:0]      EMR_LPDDR                 =16'h0000,
    parameter     integer     TMRD                      =0,        //0~3		
    parameter     integer     TMOD                      =0,        //0~7 	
    parameter     integer     TZQINIT                   =0,        //0~1023	
    parameter     integer     TXPR                      =0,        //0~15			
    parameter     integer     TRP                       =0,        //0~7
    parameter     integer     TRFC                      =0,        //0~255		
    parameter                 WL_EN                     ="FALSE",   //"TRUE" or  "FALSE"
    parameter                 DDR_TYPE                  ="DDR3",   //"DDR3" ,"DDR2", "LPDDR"   
    parameter                 DATA_WIDTH                ="16BIT",  //"16BIT","8BIT"	
    parameter     [1:0]       DQS_GATE_MODE             =2'b00,    //2'b00~2'b11	
    parameter                 WRDATA_PATH_ADJ           ="FALSE",   //"TRUE" or  "FALSE"
    parameter                 CTRL_PATH_ADJ             ="FALSE",   //"TRUE" or  "FALSE" 
    parameter     [7:0]       WL_MAX_STEP               =8'h00,
    parameter     [4:0]       WL_MAX_CHECK              =5'h0,
    parameter                 MAN_WRLVL_DQS_L           = "FALSE",   //"TRUE" or  "FALSE"
    parameter                 MAN_WRLVL_DQS_H           = "FALSE",   //"TRUE" or  "FALSE"
    parameter     [2:0]       WL_CTRL_L                 = 3'h0,
    parameter     [2:0]       WL_CTRL_H                 = 3'h0,
    parameter     [1:0]       INIT_READ_CLK_CTRL        = 2'b00,
    parameter     [1:0]       INIT_READ_CLK_CTRL_H      = 2'b00,
    parameter     [3:0]       INIT_SLIP_STEP            = 4'h0,
    parameter     [3:0]       INIT_SLIP_STEP_H          = 4'h0,
    parameter                 FORCE_READ_CLK_CTRL_L     ="FALSE",   //"TRUE" or  "FALSE"
    parameter                 FORCE_READ_CLK_CTRL_H     ="FALSE",   //"TRUE" or  "FALSE"
    parameter                 STOP_WITH_ERROR           = "TRUE",   //"TRUE" or  "FALSE"
    parameter                 DQGT_DEBUG                = 1'b0,
    parameter                 WRITE_DEBUG               = 1'b0,
    parameter     [4:0]       RDEL_ADJ_MAX_RANG         = 5'h0,
    parameter     [3:0]       MIN_DQSI_WIN              = 4'h0,
    parameter     [7:0]       INIT_SAMP_POSITION        = 8'h0,
    parameter     [7:0]       INIT_SAMP_POSITION_H      = 8'h0,
    parameter                 FORCE_SAMP_POSITION_L     ="FALSE",   //"TRUE" or  "FALSE"
    parameter                 FORCE_SAMP_POSITION_H     ="FALSE",  //"TRUE" or  "FALSE"
    parameter     [18:0]      RDEL_RD_CNT               = 19'h0,
    parameter     integer     T400NS                    = 0,      //0~127 
    parameter     [8:0]       T_LPDDR                   = 9'h0,
    parameter     [7:0]       REF_CNT                   = 8'h0,
    parameter                 APB_VLD                   = "FALSE",  //"TRUE" or  "FALSE"
    parameter     [127:0]     TEST_PATTERN1             = 128'h0000ffff0000ffff0000ffff0000ffff,
    parameter                 TRAIN_RST_TYPE            ="FALSE",  //"TRUE" or  "FALSE"
    parameter     [7:0]       TXS                       =8'h0 ,
    parameter                 WL_SETTING                =1'b1 ,
    parameter                 WCLK_DEL_SEL              =1'b0 ,
    parameter     [7:0]       INIT_WRLVL_STEP_L         =8'h0 ,
    parameter     [7:0]       INIT_WRLVL_STEP_H         =8'h0
	)(
    //---------------------------Clock and reset---------------------
    input         [1:0]      DDRPHY_UPDATE_TYPE,
    input         [1:0]      DDRPHY_UPDATE_COMP_VAL_L,
    input                    DDRPHY_UPDATE_COMP_DIR_L,
    input         [1:0]      DDRPHY_UPDATE_COMP_VAL_H,
    input                    DDRPHY_UPDATE_COMP_DIR_H,
    input                    DDRPHY_CLKIN, 
    input                    DDRPHY_RST,     
    output                   DDRPHY_RST_REQ,   
    input                    DDRPHY_RST_ACK,   
    input                    DDRPHY_UPDATE,
    output                   DDRPHY_UPDATE_DONE,

    //---------------------------APB interface-------------------------                          	
    input                    PCLK,
    input                    PRESET,
    input  [11:0]            PADDR,
    input  [31:0]            PWDATA,
    input                    PWRITE,
    input                    PSEL,
    input                    PENABLE,
    output                   PREADY,
    output [31:0]            PRDATA,

   

	//-----------------------Cmd and data ------------------------
    output                   DDRPHY_GATEI_H  ,
    output                   DDRPHY_GATEI_L  ,
    input  [7:0]             DDRPHY_DQ_L     ,
    input  [7:0]             DDRPHY_DQ_H     ,
    input                    DLL_UPDATE_ACK  ,
    output                   DLL_UPDATE_REQ  ,   
    output [7:0]             DDRPHY_WL_STEP_L, 
    output [2:0]             DDRPHY_WL_CTRL_L,
    output [2:0]             DDRPHY_RDQS_STEP_L,
    output [1:0]             DDRPHY_DQS_GATE_CTRL_L,
    output [2:0]             DDRPHY_READ_CLK_CTRL_L,
    input                    DDRPHY_WL_OV_L,   
    input                    DDRPHY_DGTS_L,
    input                    DDRPHY_READ_VALID_L, 
    input [7:0]              DDRPHY_DLL_STEP,
    input                    DDRPHY_RDEL_OV_L,
    input [31:0]             DDRPHY_RDATA_L,
    output [15:0]            DDRPHY_WEN_L,
    output [31:0]            DDRPHY_WDATA_L,
    output [3:0]             DDRPHY_WDQS_L,
    output [1:0]             DDRPHY_WDQS_EN_L,
    output [3:0]             DDRPHY_DM_L,
	
	
    output [7:0]             DDRPHY_WL_STEP_H, 
    output [2:0]             DDRPHY_WL_CTRL_H,
    output [2:0]             DDRPHY_RDQS_STEP_H,
    output [1:0]             DDRPHY_DQS_GATE_CTRL_H,
    output [2:0]             DDRPHY_READ_CLK_CTRL_H, 
	
    input                    DDRPHY_WL_OV_H,
    input                    DDRPHY_DGTS_H,
    input                    DDRPHY_READ_VALID_H,
    input                    DDRPHY_RDEL_OV_H,
    output [15:0]            DDRPHY_WEN_H,
	
    input  [31:0]            DDRPHY_RDATA_H, 
    output [31:0]            DDRPHY_WDATA_H,
    output [3:0]             DDRPHY_WDQS_H,
    output [3:0]             DDRPHY_DM_H,
    output [1:0]             DDRPHY_WDQS_EN_H,
	
	//----------------Command address-------------------------------
    output[59:0]             IOL_CE,                                                             
    output[59:0]             IOL_CLK_SYS,                                                       
    output[59:0]             IOL_LRS,                                                   
    output                   RST_DLL,                                                           
    output                   UPDATE_N,                                                                                                                             
    output                   DLL_CLK_INPUT,                                                    
    output                   DLL_FREEZE,                                                                                
    output[4:0]              DQS_RST,                                               
    output[4:0]              DQS_RST_TRAINING_N,                                       
    output[4:0]              DQS_CLK_REGIONAL,                                
    output[2:0]              DQS_GATEI,                                                 
    output[23:0]             DQS_WL_STEP,                                                     
    output[8:0]              DQS_WL_CTRL,                                            
    output[11:0]             DQS_DQS_GATE_CTRL,                                              
    output[3:0]              DQS_DQS_GATE_CTRL_TF2,                                                 
    output[8:0]              DQS_READ_CLK_CTRL,                                                     
    output[8:0]              DQS_RDEL_CTRL,                                                             
    output[103:0]            IOL_TX_DATA_TF8,                                                          
    output[183:0]            IOL_TX_DATA_TF4,                                                       
    output[6:0]              IOL_TX_DATA_TF7,                                                                                                            
    output[179:0]            IOL_IODLY_CTRL,                                                                     
    output[59:0]             IOL_MIPI_SW_DYN_I,                                                                    
    output[51:0]             IOL_TS_CTRL_TF4,                                                     
    output[91:0]             IOL_TS_CTRL_TF2,                                                                                   
    output[2:0]              IOL_TS_CTRL_TF3, 
    output                   MEM_RST_EN,
    input                    SRB_RST_DLL,
    input                    DLL_UPDATE_N,
    input                    SRB_DLL_FREEZE,
    input                    SRB_IOL_RST,
    input                    SRB_DQS_RST,
    input                    SRB_DQS_RST_TRAINING,    
    output [55:0]            DDRPHY_CA_EN,                        
    output [63:0]            DDRPHY_ADDR,
    output [11:0]            DDRPHY_BA,
    output [3:0]             DDRPHY_CK,
    output [3:0]             DDRPHY_CKE,
    output [3:0]             DDRPHY_CS_N,
    output [3:0]             DDRPHY_RAS_N,
    output [3:0]             DDRPHY_CAS_N,
    output [3:0]             DDRPHY_WE_N,
    output [3:0]             DDRPHY_ODT,
    output                   DDRPHY_MEM_RST,
                        
	//---------------DFI Interface--------------------------------
    output[63:0]             DFI_RDDATA, 
    output[3:0]              DFI_RDDATA_VALID,
    output                   DFI_CTRLUPD_ACK,           // THIS ACk is from PHY 
    output                   DFI_INIT_COMPLETE, 
    output                   DFI_PHYUPD_REQ,     // dfi phy UPDATE request 
    output [1:0]             DFI_PHYUPD_TYPE,    // dfi phy UPDATE type 
    output                   DFI_LP_ACK,         // dfi lp ACKNOWLEdge
    output                   DFI_ERROR,            
    output[2:0]              DFI_ERROR_INFO ,

    input [31:0]             DFI_ADDRESS             ,  
    input [5:0]              DFI_BANK                ,  
    input [1:0]              DFI_CAS_N               ,  
    input [1:0]              DFI_RAS_N               ,  
    input [1:0]              DFI_WE_N                ,  
    input [1:0]              DFI_CKE                 ,  
    input [1:0]              DFI_CS                  ,  
    input [1:0]              DFI_ODT                 ,  
    input [1:0]              DFI_RESET_N             ,  
    input [63:0]             DFI_WRDATA              ,  
    input [7:0]              DFI_WRDATA_MASK         ,  
    input [3:0]              DFI_WRDATA_EN           ,  
    input [3:0]              DFI_RDDATA_EN           ,  
    input                    DFI_CTRLUPD_REQ         , 
    input                    DFI_DRAM_CLK_DISABLE    ,  
    input                    DFI_INIT_START          ,  
    input [4:0]              DFI_FREQUENCY           ,  
    input                    DFI_PHYUPD_ACK          ,  
    input                    DFI_LP_REQ              ,  
    input [3:0]              DFI_LP_WAKEUP           
	);
    //synthesis translate_off 
	ddrphy_gtp_wrap #(
        .TEST_PATTERN2          (TEST_PATTERN2        ),  	
        .TEST_PATTERN3          (TEST_PATTERN3        ),
        .T200US                 (T200US               ),
        .MR0_DDR3               (MR0_DDR3             ),
        .MR1_DDR3               (MR1_DDR3             ),
        .MR2_DDR3               (MR2_DDR3             ),
        .MR3_DDR3               (MR3_DDR3             ),
        .MR_DDR2                (MR_DDR2              ),
        .EMR1_DDR2              (EMR1_DDR2            ),
        .EMR2_DDR2              (EMR2_DDR2            ),
        .EMR3_DDR2              (EMR3_DDR2            ),
        .MR_LPDDR               (MR_LPDDR             ),
        .EMR_LPDDR              (EMR_LPDDR            ),
        .TMRD                   (TMRD                 ),
        .TMOD                   (TMOD                 ),
        .TZQINIT                (TZQINIT              ),
        .TXPR                   (TXPR                 ),
        .TRP                    (TRP                  ),
        .TRFC                   (TRFC                 ),
        .WL_EN                  (WL_EN                ),
        .DDR_TYPE               (DDR_TYPE             ),
        .DATA_WIDTH             (DATA_WIDTH           ),
        .DQS_GATE_MODE          (DQS_GATE_MODE        ),
        .WRDATA_PATH_ADJ        (WRDATA_PATH_ADJ      ),
        .CTRL_PATH_ADJ          (CTRL_PATH_ADJ        ),
        .WL_MAX_STEP            (WL_MAX_STEP          ),
        .WL_MAX_CHECK           (WL_MAX_CHECK         ),
        .MAN_WRLVL_DQS_L        (MAN_WRLVL_DQS_L      ),
        .MAN_WRLVL_DQS_H        (MAN_WRLVL_DQS_H      ),
        .WL_CTRL_L              (WL_CTRL_L            ),
        .WL_CTRL_H              (WL_CTRL_H            ),
        .INIT_READ_CLK_CTRL     (INIT_READ_CLK_CTRL   ),
        .INIT_READ_CLK_CTRL_H   (INIT_READ_CLK_CTRL_H ),
        .INIT_SLIP_STEP         (INIT_SLIP_STEP       ),
        .INIT_SLIP_STEP_H       (INIT_SLIP_STEP_H     ),
        .FORCE_READ_CLK_CTRL_L  (FORCE_READ_CLK_CTRL_L),
        .FORCE_READ_CLK_CTRL_H  (FORCE_READ_CLK_CTRL_H),
        .STOP_WITH_ERROR        (STOP_WITH_ERROR      ),
        .DQGT_DEBUG             (DQGT_DEBUG           ),
        .WRITE_DEBUG            (WRITE_DEBUG          ),
        .RDEL_ADJ_MAX_RANG      (RDEL_ADJ_MAX_RANG    ),
        .MIN_DQSI_WIN           (MIN_DQSI_WIN         ),
        .INIT_SAMP_POSITION     (INIT_SAMP_POSITION   ),
        .INIT_SAMP_POSITION_H   (INIT_SAMP_POSITION_H ),
        .FORCE_SAMP_POSITION_L  (FORCE_SAMP_POSITION_L),
        .FORCE_SAMP_POSITION_H  (FORCE_SAMP_POSITION_H),
        .RDEL_RD_CNT            (RDEL_RD_CNT          ),
        .T400NS                 (T400NS               ),
        .T_LPDDR                (T_LPDDR              ),
        .REF_CNT                (REF_CNT              ),
        .APB_VLD                (APB_VLD              ),
        .TEST_PATTERN1          (TEST_PATTERN1        ),
        .TRAIN_RST_TYPE         (TRAIN_RST_TYPE       ),    
        .TXS                    (TXS                  ),
        .WL_SETTING             (WL_SETTING           ),
        .WCLK_DEL_SEL           (WCLK_DEL_SEL         ),
        .INIT_WRLVL_STEP_L      (INIT_WRLVL_STEP_L    ),
        .INIT_WRLVL_STEP_H      (INIT_WRLVL_STEP_H    )
   	 )    
	GTP_DDRPHY_WRAP(
    .mode_sel_dbg               (1'b0                ),
    .ddrphy_dbg                 (                    ),
    .srb_rst_dll                (SRB_RST_DLL         ),
    .dll_update_n               (DLL_UPDATE_N        ),
    .srb_dll_freeze             (SRB_DLL_FREEZE      ),
    .srb_iol_rst                (SRB_IOL_RST           ),
    .srb_dqs_rst                (SRB_DQS_RST           ),
    .srb_dqs_rst_training       (SRB_DQS_RST_TRAINING),
    .iol_ce                      (IOL_CE               ),                                  
    .iol_clk_sys                 (IOL_CLK_SYS          ),                                       
    .iol_lrs                     (IOL_LRS              ),                           
    .rst_dll                     (RST_DLL              ),                                   
    .update_n                    (UPDATE_N             ),                                                                                                       
    .dll_clk_input               (DLL_CLK_INPUT        ),                                       
    .dll_freeze                  (DLL_FREEZE           ),                                                             
    .dqs_rst                     (DQS_RST              ),                      
    .dqs_rst_training_n          (DQS_RST_TRAINING_N   ),                                   
    .dqs_clk_regional            (DQS_CLK_REGIONAL     ),                       
    .dqs_gatei                   (DQS_GATEI            ),                          
    .dqs_wl_step                 (DQS_WL_STEP          ),                                   
    .dqs_wl_ctrl                 (DQS_WL_CTRL          ),                          
    .dqs_dqs_gate_ctrl           (DQS_DQS_GATE_CTRL    ),                                       
    .dqs_dqs_gate_ctrl_tf2       (DQS_DQS_GATE_CTRL_TF2),                                                 
    .dqs_read_clk_ctrl           (DQS_READ_CLK_CTRL    ),                                            
    .dqs_rdel_ctrl               (DQS_RDEL_CTRL        ),                                            
    .iol_tx_data_tf8             (IOL_TX_DATA_TF8      ),                                              
    .iol_tx_data_tf4             (IOL_TX_DATA_TF4      ),                                           
    .iol_tx_data_tf7             (IOL_TX_DATA_TF7      ),                                                                                                 
    .iol_iodly_ctrl              (IOL_IODLY_CTRL       ),                                                       
    .iol_mipi_sw_dyn_i           (IOL_MIPI_SW_DYN_I    ),                                                             
    .iol_ts_ctrl_tf4             (IOL_TS_CTRL_TF4      ),                                          
    .iol_ts_ctrl_tf2             (IOL_TS_CTRL_TF2      ),                                                                       
    .iol_ts_ctrl_tf3             (IOL_TS_CTRL_TF3      ),                                                                                                 
    .mem_rst_en                  (MEM_RST_EN           ),                             
    .update_type                 (DDRPHY_UPDATE_TYPE),
    .update_comp_val_l           (DDRPHY_UPDATE_COMP_VAL_L),
    .update_comp_dir_l           (DDRPHY_UPDATE_COMP_DIR_L),
    .update_comp_val_h           (DDRPHY_UPDATE_COMP_VAL_H),
    .update_comp_dir_h           (DDRPHY_UPDATE_COMP_DIR_H),
    .ddrphy_clkin                (DDRPHY_CLKIN           ),
	.ddrphy_rst                  (DDRPHY_RST           ),
	.ddrphy_rst_req              (DDRPHY_RST_REQ         ),
	.ddrphy_rst_ack              (DDRPHY_RST_ACK         ),
	.ddrphy_update               (DDRPHY_UPDATE          ),
	.ddrphy_update_done          (DDRPHY_UPDATE_DONE     ),
	.pclk                        (PCLK                   ),
	.preset                      (PRESET                ),
	.paddr                       (PADDR                  ),
	.pwdata                      (PWDATA                 ),
	.pwrite                      (PWRITE                 ),
	.psel                        (PSEL                   ),
	.penable                     (PENABLE                ),
	.pready                      (PREADY                 ),
	.prdata                      (PRDATA                 ),
	.ddrphy_wl_step_l            (DDRPHY_WL_STEP_L       ),
	.ddrphy_wl_ctrl_l            (DDRPHY_WL_CTRL_L       ),
	.ddrphy_rdqs_step_l          (DDRPHY_RDQS_STEP_L     ),
	.ddrphy_dqs_gate_ctrl_l      (DDRPHY_DQS_GATE_CTRL_L ),
	.ddrphy_read_clk_ctrl_l      (DDRPHY_READ_CLK_CTRL_L ),
	.ddrphy_wl_ov_l              (DDRPHY_WL_OV_L         ),
	.ddrphy_dgts_l               (DDRPHY_DGTS_L          ),
	.ddrphy_read_valid_l         (DDRPHY_READ_VALID_L    ),
	.ddrphy_dll_step             (DDRPHY_DLL_STEP      ),
	.ddrphy_rdel_ov_l            (DDRPHY_RDEL_OV_L       ),
	.ddrphy_rdata_l              (DDRPHY_RDATA_L         ),
	.ddrphy_wen_l                (DDRPHY_WEN_L           ),
	.ddrphy_wdata_l              (DDRPHY_WDATA_L         ),
	.ddrphy_wdqs_l               (DDRPHY_WDQS_L          ),
	.ddrphy_wdqs_en_l            (DDRPHY_WDQS_EN_L       ),
	.ddrphy_dm_l                 (DDRPHY_DM_L            ),
    .ddrphy_wl_step_h            (DDRPHY_WL_STEP_H       ),
	.ddrphy_wl_ctrl_h            (DDRPHY_WL_CTRL_H       ),
	.ddrphy_rdqs_step_h          (DDRPHY_RDQS_STEP_H     ),
	.ddrphy_dqs_gate_ctrl_h      (DDRPHY_DQS_GATE_CTRL_H ),
	.ddrphy_read_clk_ctrl_h      (DDRPHY_READ_CLK_CTRL_H ),
	.ddrphy_wl_ov_h              (DDRPHY_WL_OV_H         ),
	.ddrphy_dgts_h               (DDRPHY_DGTS_H          ),
	.ddrphy_read_valid_h         (DDRPHY_READ_VALID_H    ),
	.ddrphy_rdel_ov_h            (DDRPHY_RDEL_OV_H       ),
	.ddrphy_wen_h                (DDRPHY_WEN_H           ),
	.ddrphy_rdata_h              (DDRPHY_RDATA_H         ),
	.ddrphy_wdata_h              (DDRPHY_WDATA_H         ),
	.ddrphy_wdqs_h               (DDRPHY_WDQS_H          ),
	.ddrphy_dm_h                 (DDRPHY_DM_H            ),
	.ddrphy_wdqs_en_h            (DDRPHY_WDQS_EN_H       ),
	.ddrphy_ca_en                (DDRPHY_CA_EN           ),
	.ddrphy_addr                 (DDRPHY_ADDR            ),
	.ddrphy_ba                   (DDRPHY_BA              ),
	.ddrphy_ck                   (DDRPHY_CK              ),
	.ddrphy_cke                  (DDRPHY_CKE             ),
	.ddrphy_cs_n                 (DDRPHY_CS_N            ),
	.ddrphy_ras_n                (DDRPHY_RAS_N           ),
	.ddrphy_cas_n                (DDRPHY_CAS_N           ),
	.ddrphy_we_n                 (DDRPHY_WE_N            ),
	.ddrphy_odt                  (DDRPHY_ODT             ),
	.ddrphy_mem_rst              (DDRPHY_MEM_RST     ),
	.dfi_rddata                  (DFI_RDDATA             ),
	.dfi_rddata_valid            (DFI_RDDATA_VALID       ),
	.dfi_ctrlupd_ack             (DFI_CTRLUPD_ACK        ),
    .dfi_init_complete           (DFI_INIT_COMPLETE      ),
	.dfi_phyupd_req              (DFI_PHYUPD_REQ         ),
	.dfi_phyupd_type             (DFI_PHYUPD_TYPE        ),
	.dfi_lp_ack                  (DFI_LP_ACK             ),
	.dfi_error                   (DFI_ERROR              ),
	.dfi_error_info              (DFI_ERROR_INFO         ),
	.dfi_address                   (DFI_ADDRESS          ), 
	.dfi_bank                      (DFI_BANK             ),
	.dfi_cas_n                     (DFI_CAS_N            ),
	.dfi_ras_n                     (DFI_RAS_N            ),
	.dfi_we_n                      (DFI_WE_N             ),
	.dfi_cke                       (DFI_CKE              ),
	.dfi_cs                        (DFI_CS               ),
	.dfi_odt                       (DFI_ODT              ),
	.dfi_reset_n                   (DFI_RESET_N          ),
	.dfi_wrdata                    (DFI_WRDATA           ),
	.dfi_wrdata_mask               (DFI_WRDATA_MASK      ),
	.dfi_wrdata_en                 (DFI_WRDATA_EN        ),
	.dfi_rddata_en                 (DFI_RDDATA_EN        ),
	.dfi_ctrlupd_req               (DFI_CTRLUPD_REQ      ),
	.dfi_dram_clk_disable          (DFI_DRAM_CLK_DISABLE ),
	.dfi_init_start                (DFI_INIT_START       ),
	.dfi_frequency                 (DFI_FREQUENCY        ),
	.dfi_phyupd_ack                (DFI_PHYUPD_ACK       ),
	.dfi_lp_req                    (DFI_LP_REQ           ),
	.dfi_lp_wakeup                 (DFI_LP_WAKEUP        ),
    .ddrphy_gatei_h                (DDRPHY_GATEI_H       ),
    .ddrphy_gatei_l                (DDRPHY_GATEI_L       ),
    .ddrphy_dq_l                   (DDRPHY_DQ_L),
    .ddrphy_dq_h                   (DDRPHY_DQ_H),
    .dll_update_ack                (DLL_UPDATE_ACK),
    .dll_update_req                (DLL_UPDATE_REQ)
	);
	//synthesis translate_on
	
endmodule
	
	
	
	
	
	
	






//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_MULT9.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

//P=A*B
module GTP_MULT9 #(
    parameter GRS_EN    = "TRUE",  //"TRUE"; "FALSE"
    parameter SYNC_RST  = "FALSE",  //"TRUE"; "FALSE"
    parameter INREG_EN  = "FALSE",  //"TRUE"; "FALSE"
    parameter OUTREG_EN = "FALSE"   //"TRUE"; "FALSE"
) (
    output  [18-1:0] P,
    input   CE,
    input   RST,
    input   CLK,
    input   A_SIGNED,
    input   [9-1:0] A,
    input   B_SIGNED,
    input   [9-1:0] B
);


    INT_PREADD_MULT #(
        .GRS_EN(GRS_EN),
        .SYNC_RST(SYNC_RST),
        .INREG_EN(INREG_EN),
        .OUTREG_EN(OUTREG_EN),
        .ASIZE(9),
        .BSIZE(9),
        .PREADD_EN(0)
    ) U_INT_MULT (
        .CE(CE),
        .RST(RST),
        .CLK(CLK),
        .A_SIGNED(A_SIGNED),
        .A(A),
        .B_SIGNED(B_SIGNED),
        .B(B),
        .C_SIGNED(B_SIGNED),
        .C(9'b0),
        .PREADDSUB(1'b0),
        .P(P)
    );

endmodule






//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_PREADD_MULT18.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

//P = A*(B+C)
`timescale 1 ns / 1 ps

module GTP_PREADD_MULT18 #(
    parameter GRS_EN      = "TRUE", //"TRUE"; "FALSE"
    parameter SYNC_RST    = "FALSE", //"TRUE"; "FALSE"
    parameter INREG_EN    = "FALSE", //"TRUE"; "FALSE"
    parameter PREREG_EN   = "FALSE", //"TRUE"; "FALSE"
    parameter OUTREG_EN   = "FALSE"  //"TRUE"; "FALSE"
)(
    output  [37-1:0] P,
    input   CE,
    input   RST,
    input   CLK,
    input   A_SIGNED,
    input   [18-1:0] A,
    input   B_SIGNED,
    input   [18-1:0] B,
    input   C_SIGNED,
    input   [18-1:0] C,
    input   PREADDSUB
);

    INT_PREADD_MULT  #(.GRS_EN(GRS_EN),
         .SYNC_RST(SYNC_RST),    
         .INREG_EN(INREG_EN),    
         .PREREG_EN(PREREG_EN),    
         .OUTREG_EN(OUTREG_EN),   
         .ASIZE(18),
         .BSIZE(18)
    )  U_INT_PREADD_MULT (
        .CE(CE),
        .RST(RST),
        .CLK(CLK),
        .A_SIGNED(A_SIGNED),
        .A(A),
        .B_SIGNED(B_SIGNED),
        .B(B),
        .C_SIGNED(C_SIGNED),
        .C(C),
        .PREADDSUB(PREADDSUB),
        .P(P)
    );

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2016 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_CLKBUFXCE.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_CLKBUFXCE
#(
    parameter TRIGGER_MODE = "POSEDGE",
    parameter CE_TYPE = "SYNC",
    parameter CE_INV = "FALSE"

) (
    output CLKOUT,
    input CLKIN,
    input CE
);

//synthesis translate_off

    initial begin
        if(CE_TYPE != "SYNC" && CE_TYPE != "ASYNC") begin
            $display("ERROR: The attribute CE_TYPE on instance %m is %s. Legal value are SYNC or ASYNC.", CE_TYPE);
            $finish;
        end
        if(TRIGGER_MODE != "POSEDGE" && TRIGGER_MODE != "NEGEDGE") begin
            $display("ERROR: The attribute TRIGGER_MODE on instance %m is %s. Legal value are POSEDGE or NEGEDGE.", TRIGGER_MODE);
            $finish;
        end
        if(CE_INV != "TRUE" && CE_INV != "FALSE") begin
            $display("ERROR: The attribute CE_INV on instance %m is %s. Legal value are TRUE or FALSE.", CE_INV);
            $finish;
        end        
    end

    wire ce;
    wire outs;
    wire outps;
    wire outns;
    wire outa;
    wire outpa;
    wire outna;
    
    reg flag1;
    reg flag2;
    reg mid1;
    reg mid2;

    initial begin
        flag1 = 0;
        flag2 = 0;
        mid1 = 0;
        mid2 = 0;
        #0.1 ;
        flag1 = 0;
        flag2 = 0;
        mid1 = 0;
        mid2 = 0;
    end

    assign ce = (CE_INV == "FALSE")? CE : !CE;
    assign CLKOUT = (CE_TYPE == "SYNC")? outs : outa;
    assign outs = (TRIGGER_MODE == "POSEDGE")? outps : outns;
    assign outps = flag1? CLKIN : 1'b1;
    assign outns = flag2? CLKIN : 1'b0;
    assign outa = (TRIGGER_MODE == "POSEDGE")? outpa : outna;
    assign outpa = ce? CLKIN : 1'b1;
    assign outna = ce? CLKIN : 1'b0;

    always@(posedge CLKIN) begin
        if(ce) begin
            flag1 <= mid1;
            mid1 <= 1;
        end        
        else begin
            flag1 <= mid1;
            mid1 <= 0;
        end
    end

    always@(negedge CLKIN) begin
        if(ce) begin
            flag2 <= mid2;
            mid2 <= 1;
    
        end
        else begin
            flag2 <= mid2;
            mid2 <= 0;
        end        
    end


//synthesis translate_on

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2016 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_CFGCLK
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_CFGCLK
#(

) (
    input CLKIN,
    input CE_N
);

//synthesis translate_off


//synthesis translate_on
endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_START_E1.v
//
// Functional description: startup Logic Control Circuit
//
// Parameter description:
//      
//
// Port description:
//      
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps 

module GTP_START_E1
(
    input           CLK    ,          //start signals
    input tri0      GOE,
    input tri0      GRS_N  ,
    input tri0      GWE  ,
    output reg      WAKEUP_OVER
);

wire        GOUTEN     ;
wire        GRSN       ;
wire        GWEN       ;

assign GOUTEN = GOE;
assign GRSN   = GRS_N  ;
assign GWEN   = GWE  ;

initial begin
    WAKEUP_OVER = 1'b1;
#50000
    WAKEUP_OVER = 1'b0;
end

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_ROM64X1.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_ROM64X1
#(
    parameter [63:0] INIT = 64'h0000_0000_0000_0000
) (
    output Z,
    input I0, I1, I2, I3, I4, I5
);

   reg [63:0] mem;
   wire [5:0] addr;

   initial mem = INIT;

   assign addr = {I5, I4, I3, I2, I1, I0};
   //assign Z = mem[addr];
   assign Z = INIT[addr];

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_PREADD_MULT36.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

//P = A*(B+C)
`timescale 1 ns / 1 ps

module GTP_PREADD_MULT36 #(
    parameter GRS_EN      = "TRUE", //"TRUE"; "FALSE"
    parameter SYNC_RST    = "FALSE", //"TRUE"; "FALSE"
    parameter INREG_EN    = "FALSE",  //"TRUE"; "FALSE"
    parameter PREREG_EN   = "FALSE",  //"TRUE"; "FALSE"
    parameter OUTREG_EN   = "FALSE"    //"TRUE"; "FALSE"
)(
    output  [55-1:0] P,
    input   CE,
    input   RST,
    input   CLK,
    input   A_SIGNED,
    input   [36-1:0] A,
    input   B_SIGNED,
    input   [18-1:0] B,
    input   C_SIGNED,
    input   [18-1:0] C,
    input   PREADDSUB
);

    INT_PREADD_MULT  #(.GRS_EN(GRS_EN),
        .SYNC_RST(SYNC_RST),    
        .INREG_EN(INREG_EN),    
        .PREREG_EN(PREREG_EN),    
        .OUTREG_EN(OUTREG_EN),   
        .ASIZE(36),  
        .BSIZE(18)
    ) U_INT_PREADD_MULT (
        .CE(CE),
        .RST(RST),
        .CLK(CLK),
        .A_SIGNED(A_SIGNED),
        .A(A),
        .B_SIGNED(B_SIGNED),
        .B(B),
        .C_SIGNED(C_SIGNED),
        .C(C),
        .PREADDSUB(PREADDSUB),
        .P(P)
    );

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2016 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_RAM64X1DP.v
//
// Functional description: simple-dual-port 64x1 distributed ram
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_RAM64X1DP
#(
    parameter [63:0] INIT = 64'h0000_0000_0000_0000
) (
    output  DO,
    input   DI,
    input [5:0] RADDR,
    input [5:0] WADDR,
    input WCLK,
    input WE
);
//synthesis translate_off
    reg [63:0] mem ;

    initial begin
        mem = INIT;
    end

    always @(posedge WCLK) begin
        if (WE == 1'b1) begin
            mem[WADDR] <= DI;
        end
    end

    assign DO = mem[RADDR];
//synthesis translate_on
endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_DDC_E1.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_DDC_E1 #(
parameter GRS_EN = "TRUE",             //"TRUE"; "FALSE"
parameter DDC_MODE = "FULL_RATE", //"FULL_RATE"; "HALF_RATE"; "QUAD_RATE"
parameter IFIFO_GENERIC  ="FALSE",       //"TRUE"; "FALSE"
parameter WCLK_DELAY_OFFSET = 9'd0,          //0~255 for posedge adjust; 256~511 for negedge adjust; bit[8] used as signed flag
parameter DQSI_DELAY_OFFSET = 9'd0,          //0~255 for posedge adjust; 256~511 for negedge adjust; bit[8] used as signed flag
parameter CLKA_GATE_EN = "FALSE",
parameter R_DELAY_STEP_EN = "TRUE", //"TRUE"; "FALSE"
parameter R_MOVE_EN = "FALSE", //"TRUE"; "FALSE"
parameter W_MOVE_EN = "FALSE", //"TRUE"; "FALSE"
parameter R_EXTEND = "FALSE", //"TRUE"; "FALSE"
parameter GATE_SEL = "FALSE",   //"TRUE"; "FALSE"
parameter WCLK_DELAY_SEL = "FALSE", //"TRUE"; "FALSE"
parameter RCLK_SEL = "FALSE", //"TRUE"; "FALSE"
parameter RADDR_INIT = 3'd0
)(
    //output
    output WDELAY_OB,
    output WCLK,
    output WCLK_DELAY,
    output RCLK,
    output RDELAY_OB,
    output DQSI_DELAY,
    output DGTS,
    output READ_VALID,
    output GATE_OUT,
    output [2:0] IFIFO_WADDR,
    output [2:0] IFIFO_RADDR,
    output [1:0] DQS_DRIFT,
    output DRIFT_DETECT_ERR,
    output DQS_DRIFT_STATUS,
    //input
    input RST,
    input CLKB,
    input CLKA,
    input CLKA_GATE,
    input [7:0] DELAY_STEP1,
    input [7:0] DELAY_STEP0,
    input       W_DIRECTION,
    input       W_MOVE,
    input       W_LOAD_N,
    input [3:0] DQS_GATE_CTRL,
    input [2:0] READ_CLK_CTRL,
    input DQSI,
    input GATE_IN,
    input      R_DIRECTION,
    input      R_MOVE,
    input      R_LOAD_N,
    input      RST_TRAINING_N
)/* synthesis syn_black_box */;

//synthesis translate_off
    //reg statement
    reg wclk_source_dly;
    reg wclk_del_source_dly;
    reg dqsin_gated_dly;
    reg [1:0] DQS_GATE_CTRL_gate_d;
    reg [1:0] DQS_GATE_CTRL_gate_dd;
    reg [3:0] DQS_GATE_CTRL_d1;
    reg [3:0] DQS_GATE_CTRL_d2;
    reg [3:0] DQS_GATE_CTRL_d3;
    reg gate_st;
    reg [3:0] DQS_GATE_CTRL_d4;
    reg DQS_GATE_CTRL_d5;
    reg DQS_GATE_CTRL_d6;
    reg sel_gate_clk;
    reg DQS_GATE_CTRL_gate;
    reg DQS_GATE_CTRL_comb_d1;
    reg DQS_GATE_CTRL_comb_d2;
    reg [1:0] DQS_GATE_CTRL_comb_and_d;
    reg start_wr;
    reg [2:0] WADDR_reg;
    reg [2:0] IFIFO_WADDR_reg;
    reg start_rd;
    reg [2:0] RADDR_reg;
    reg RDVALID_reg;
    reg DQSIN_gated_reg;
    reg [7:0] adj_dly_wclk_del;
    reg [7:0] adj_dly_dqsi;
    reg read_enable_tmp;
    reg new_st;
    reg new_transfer_d;
    reg read_enable_d1;
    reg read_enable_d2;
    reg [1:0] cnt;
    reg [1:0] gate_cnt;
    reg [1:0] new_cnt;
    reg [2:0] gate_d;
    reg [1:0] cnt_gate;
    reg [2:0] WADDR_reg_d1;
    reg [2:0] WADDR_reg_d2;
    reg [2:0] RADDR_reg_plus1;
    reg new_rd_en_reg;
    reg new_cnt_reg;
    reg [3:0] q;
    reg [1:0] dqs_drift_reg;
    reg       drift_detect_err_reg;
    reg w_move_enable;
    reg r_move_enable;
    reg out;
    //wire statement
    wire saout;
    wire saout_b;
    wire drift_status_0;
    wire drift_status_1;
    wire dqs_drift_status;

    wire DQSIN_gated;
    wire new_transfer;
    
    wire DQS_GATE_CTRL_d2_d;
    wire DQS_GATE_CTRL_d2_dd;
    wire[3:0] DQS_GATE_CTRL_d3_d;
    wire DQS_GATE_CTRL_d5_d;
    wire DQS_GATE_CTRL_d6_d;
    wire set_en;
    wire DQS_GATE_CTRL_gate_dly;

initial 
begin
    if ((GRS_EN == "TRUE")  || (GRS_EN == "FALSE")) 
    begin
    end
    else
    begin
        $display (" GTP_DDC_E1 error: illegal setting for GRS_EN"); 
    end
    if ((DDC_MODE == "FULL_RATE") || (DDC_MODE == "HALF_RATE")  || (DDC_MODE == "QUAD_RATE")) 
    begin
    end
    else 
    begin
        $display (" GTP_DDC_E1 error: illegal setting for DDC_MODE");
    end
    if ((IFIFO_GENERIC == "TRUE") || (IFIFO_GENERIC == "FALSE")) 
    begin
    end
    else
    begin
       $display (" GTP_DDC_E1 error: illegal setting for IFIFO_GENERIC");
    end
    if ((CLKA_GATE_EN == "TRUE")   || (CLKA_GATE_EN == "FALSE")) 
    begin
    end
    else
    begin
        $display (" GTP_DDC_E1 error: illegal setting for CLKA_GATE_EN");
    end
    if ((R_DELAY_STEP_EN == "TRUE")   || (R_DELAY_STEP_EN == "FALSE")) 
    begin
    end
    else
    begin
        $display (" GTP_DDC_E1 error: illegal setting for R_DELAY_STEP_EN");
    end
    if ((R_MOVE_EN == "TRUE")   || (R_MOVE_EN == "FALSE")) 
    begin
    end
    else
    begin
        $display (" GTP_DDC_E1 error: illegal setting for R_MOVE_EN");
    end
    if ((W_MOVE_EN == "TRUE")   || (W_MOVE_EN == "FALSE")) 
    begin
    end
    else
    begin
        $display (" GTP_DDC_E1 error: illegal setting for W_MOVE_EN");
    end
    if ((R_EXTEND == "TRUE")   || (R_EXTEND == "FALSE")) 
    begin
    end
    else
    begin
        $display (" GTP_DDC_E1 error: illegal setting for R_EXTEND");
    end

    if ((GATE_SEL == "TRUE")   || (GATE_SEL == "FALSE"))
    begin
    end
    else
    begin
        $display (" GTP_DDC_E1 error: illegal setting for GATE_SEL");
    end

    if ((RCLK_SEL == "TRUE")   || (RCLK_SEL == "FALSE"))
    begin
    end
    else
    begin
        $display (" GTP_DDC_E1 error: illegal setting for RCLK_SEL");
    end

    if ((WCLK_DELAY_SEL == "TRUE")   || (WCLK_DELAY_SEL == "FALSE"))
    begin
    end
    else
    begin
        $display (" GTP_DDC_E1 error: illegal setting for WCLK_DELAY_SEL");
    end

    DQSIN_gated_reg = 1'b0;  
    DQS_GATE_CTRL_gate_d = 0;
    DQS_GATE_CTRL_gate_dd = 0;
    DQS_GATE_CTRL_d1 = 0;
    DQS_GATE_CTRL_d2 = 0;
    DQS_GATE_CTRL_d3 = 0;
    gate_st          = 0;
    DQS_GATE_CTRL_d4 = 0;
    DQS_GATE_CTRL_d5 = 0;
    DQS_GATE_CTRL_d6 = 0;
    sel_gate_clk = 0;
    DQS_GATE_CTRL_gate = 0;
    DQS_GATE_CTRL_comb_d1 = 0;
    DQS_GATE_CTRL_comb_d2 = 0;
    DQS_GATE_CTRL_comb_and_d = 0;
    start_wr  = 0;
    WADDR_reg = 0;
    IFIFO_WADDR_reg = 0;
    start_rd  = 0;
    RADDR_reg = RADDR_INIT;
    RDVALID_reg = 0;
    DQSIN_gated_reg = 0;
    adj_dly_wclk_del = 0;
    adj_dly_dqsi = 0;
    read_enable_tmp = 0;
    new_st = 0;
    new_transfer_d = 0;
    read_enable_d1 = 0;
    read_enable_d2 = 0;
    cnt = 0;
    gate_cnt = 0;
    new_cnt = 0;  
    gate_d = 0;
    WADDR_reg_d1 = 0;
    WADDR_reg_d2 = 0;
    RADDR_reg_plus1 = 0;
    new_rd_en_reg = 0;
    new_cnt_reg = 0;
    cnt_gate = 2'b0;
    q = 4'b0;
    dqs_drift_reg = 2'b0;
    drift_detect_err_reg = 1'b0;
    dqsin_gated_dly = 1'b0;
    wclk_source_dly = 1'b0;
    wclk_del_source_dly = 1'b0;
    out = 1'b0;
    w_move_enable = 1'b0;
    r_move_enable = 1'b0; 
end

assign global_rstn = GRS_EN == "TRUE" ? GRS_INST.GRSNET : 1'b1;
assign lsr_rstn = ~RST;

wire [1:0] cnt_gate_next;
wire global_rstn_cgn;
wire lsr_rstn_cgn;
wire gatein;

wire rst_transfer_n;

assign gatein = CLKA_GATE_EN == "TRUE" ? (~CLKA_GATE) : 1'b1;

assign rstn_fifo = (lsr_rstn & global_rstn) & gatein & RST_TRAINING_N;

assign rst_start_rd = start_rd & rstn_fifo;

assign rst_transfer_n = lsr_rstn & global_rstn;

always @(negedge CLKA or posedge RST)
begin
    if (RST) 
    begin
        gate_d <= 3'd0;
    end
    else if (CLKA_GATE_EN == "TRUE")
        gate_d <= {gate_d[1:0], CLKA_GATE};
    else
        gate_d <= 3'd0;
end

always @(negedge CLKA or posedge RST)
begin
   if (RST)
   begin
       cnt_gate <= 2'b0;
   end
   else if((gate_d[2]==1'b1)||(cnt_gate!=2'b0))
       cnt_gate <= cnt_gate_next;
end

assign cnt_gate_next[0] = ~cnt_gate[0];
assign cnt_gate_next[1] = cnt_gate[0] ? ~cnt_gate[1] : cnt_gate[1];

assign ioclk_gated = (gate_d[2]==1'b1)||(cnt_gate!=2'b0) ? 0 : CLKA;

wire [255:0] wclk_delay_chain;
wire wclk_source;

assign wclk_source = (DDC_MODE == "FULL_RATE") ? CLKB : ioclk_gated;

always @(*)
begin
    wclk_source_dly <= #0.2 wclk_source;
end

assign wclk_delay_chain[0] =  wclk_source_dly;
genvar gen_i;
generate  
    for(gen_i=1;gen_i<256;gen_i=gen_i+1) 
    begin
        assign #0.025 wclk_delay_chain[gen_i] =  wclk_delay_chain[gen_i-1];
    end
endgenerate

assign WCLK_comb = DELAY_STEP0[7] ? wclk_delay_chain[127] :  wclk_delay_chain[DELAY_STEP0];

assign WCLK = WCLK_comb;

wire clk_r0;

assign clk_r0 = wclk_delay_chain[0];

assign RCLK = (RCLK_SEL == "TRUE") ? clk_r0 : (~clk_r0);

assign WL_CTRL_b0_tmp = W_MOVE_EN == "TRUE" ? W_LOAD_N : 1'b1;
wire [8:0]  WCLK_DEL_OFFSET_tmp = WCLK_DELAY_OFFSET;

//wire [7:0] DLL_STEP_PLUS_WCLK_DEL_OFFSET = WCLK_DEL_OFFSET_tmp[8] ? (DLL_STEP - WCLK_DEL_OFFSET_tmp[7:0]) : (DLL_STEP + WCLK_DEL_OFFSET_tmp[7:0]);
wire [7:0] DLL_STEP_PLUS_WCLK_DEL_OFFSET = DELAY_STEP1 + WCLK_DEL_OFFSET_tmp[7:0];

wire DLL_STEP_PLUS_WCLK_DEL_OFFSET_co_0 = DELAY_STEP1[0] && WCLK_DEL_OFFSET_tmp[0];
wire DLL_STEP_PLUS_WCLK_DEL_OFFSET_co_1 = (DELAY_STEP1[1] && WCLK_DEL_OFFSET_tmp[1]) || ((DELAY_STEP1[1] || WCLK_DEL_OFFSET_tmp[1]) && DLL_STEP_PLUS_WCLK_DEL_OFFSET_co_0);
wire DLL_STEP_PLUS_WCLK_DEL_OFFSET_co_2 = (DELAY_STEP1[2] && WCLK_DEL_OFFSET_tmp[2]) || ((DELAY_STEP1[2] || WCLK_DEL_OFFSET_tmp[2]) && DLL_STEP_PLUS_WCLK_DEL_OFFSET_co_1);
wire DLL_STEP_PLUS_WCLK_DEL_OFFSET_co_3 = (DELAY_STEP1[3] && WCLK_DEL_OFFSET_tmp[3]) || ((DELAY_STEP1[3] || WCLK_DEL_OFFSET_tmp[3]) && DLL_STEP_PLUS_WCLK_DEL_OFFSET_co_2);
wire DLL_STEP_PLUS_WCLK_DEL_OFFSET_co_4 = (DELAY_STEP1[4] && WCLK_DEL_OFFSET_tmp[4]) || ((DELAY_STEP1[4] || WCLK_DEL_OFFSET_tmp[4]) && DLL_STEP_PLUS_WCLK_DEL_OFFSET_co_3);
wire DLL_STEP_PLUS_WCLK_DEL_OFFSET_co_5 = (DELAY_STEP1[5] && WCLK_DEL_OFFSET_tmp[5]) || ((DELAY_STEP1[5] || WCLK_DEL_OFFSET_tmp[5]) && DLL_STEP_PLUS_WCLK_DEL_OFFSET_co_4);
wire DLL_STEP_PLUS_WCLK_DEL_OFFSET_co_6 = (DELAY_STEP1[6] && WCLK_DEL_OFFSET_tmp[6]) || ((DELAY_STEP1[6] || WCLK_DEL_OFFSET_tmp[6]) && DLL_STEP_PLUS_WCLK_DEL_OFFSET_co_5);
wire DLL_STEP_PLUS_WCLK_DEL_OFFSET_co_7 = (DELAY_STEP1[7] && WCLK_DEL_OFFSET_tmp[7]) || ((DELAY_STEP1[7] || WCLK_DEL_OFFSET_tmp[7]) && DLL_STEP_PLUS_WCLK_DEL_OFFSET_co_6);


assign DLL_STEP_PLUS_WCLK_DEL_OFFSET_sel= ~(WCLK_DEL_OFFSET_tmp[8] ^ DLL_STEP_PLUS_WCLK_DEL_OFFSET_co_7);


wire [7:0] DLL_STEP_WCLK_DEL = WCLK_DEL_OFFSET_tmp[8] ? (DLL_STEP_PLUS_WCLK_DEL_OFFSET_sel ? DLL_STEP_PLUS_WCLK_DEL_OFFSET[7:0] : 8'd0) :
                              (DLL_STEP_PLUS_WCLK_DEL_OFFSET_sel ? DLL_STEP_PLUS_WCLK_DEL_OFFSET[7:0] : 8'd255);

wire [7:0] WL_STEP_24 = (DDC_MODE == "FULL_RATE") ? 8'd0 : DELAY_STEP0; 

wire [7:0] adj_dly_wclk_del_9b = DLL_STEP_WCLK_DEL + WL_STEP_24;

wire DLL_STEP_PLUS_WCLK_DEL_OFFSET2_co_0 = DLL_STEP_WCLK_DEL[0] && WL_STEP_24[0];
wire DLL_STEP_PLUS_WCLK_DEL_OFFSET2_co_1 = (DLL_STEP_WCLK_DEL[1] && WL_STEP_24[1]) || ((DLL_STEP_WCLK_DEL[1] || WL_STEP_24[1]) && DLL_STEP_PLUS_WCLK_DEL_OFFSET2_co_0);
wire DLL_STEP_PLUS_WCLK_DEL_OFFSET2_co_2 = (DLL_STEP_WCLK_DEL[2] && WL_STEP_24[2]) || ((DLL_STEP_WCLK_DEL[2] || WL_STEP_24[2]) && DLL_STEP_PLUS_WCLK_DEL_OFFSET2_co_1);
wire DLL_STEP_PLUS_WCLK_DEL_OFFSET2_co_3 = (DLL_STEP_WCLK_DEL[3] && WL_STEP_24[3]) || ((DLL_STEP_WCLK_DEL[3] || WL_STEP_24[3]) && DLL_STEP_PLUS_WCLK_DEL_OFFSET2_co_2);
wire DLL_STEP_PLUS_WCLK_DEL_OFFSET2_co_4 = (DLL_STEP_WCLK_DEL[4] && WL_STEP_24[4]) || ((DLL_STEP_WCLK_DEL[4] || WL_STEP_24[4]) && DLL_STEP_PLUS_WCLK_DEL_OFFSET2_co_3);
wire DLL_STEP_PLUS_WCLK_DEL_OFFSET2_co_5 = (DLL_STEP_WCLK_DEL[5] && WL_STEP_24[5]) || ((DLL_STEP_WCLK_DEL[5] || WL_STEP_24[5]) && DLL_STEP_PLUS_WCLK_DEL_OFFSET2_co_4);
wire DLL_STEP_PLUS_WCLK_DEL_OFFSET2_co_6 = (DLL_STEP_WCLK_DEL[6] && WL_STEP_24[6]) || ((DLL_STEP_WCLK_DEL[6] || WL_STEP_24[6]) && DLL_STEP_PLUS_WCLK_DEL_OFFSET2_co_5);
wire DLL_STEP_PLUS_WCLK_DEL_OFFSET2_co_7 = (DLL_STEP_WCLK_DEL[7] && WL_STEP_24[7]) || ((DLL_STEP_WCLK_DEL[7] || WL_STEP_24[7]) && DLL_STEP_PLUS_WCLK_DEL_OFFSET2_co_6);

assign DLL_STEP_PLUS_WCLK_DEL_OFFSET_sel2= ~(1'b0 ^ DLL_STEP_PLUS_WCLK_DEL_OFFSET2_co_7);

wire [7:0] adj_dly_wclk_del_init = DLL_STEP_PLUS_WCLK_DEL_OFFSET_sel2 ? adj_dly_wclk_del_9b[7:0] : 8'd255;



always @(WL_CTRL_b0_tmp or adj_dly_wclk_del_init) 
begin
    if (WL_CTRL_b0_tmp) 
        adj_dly_wclk_del <= adj_dly_wclk_del_init;    
end
always @(*)
begin
    w_move_enable <= #3 W_MOVE&(~WDELAY_OB);
end
      
always @(negedge W_MOVE) 
begin
    if (WL_CTRL_b0_tmp)
        adj_dly_wclk_del <= adj_dly_wclk_del_init;
    else if(w_move_enable)
    begin
        if (W_DIRECTION && (adj_dly_wclk_del != 8'd0))
            adj_dly_wclk_del <= adj_dly_wclk_del - 1;
        else if ((~W_DIRECTION) && (adj_dly_wclk_del[6:0] != 7'd127)&&(~adj_dly_wclk_del[7]))
            adj_dly_wclk_del <= adj_dly_wclk_del + 1;
    end
end


assign WDELAY_OB = (W_DIRECTION && (adj_dly_wclk_del == 8'd0)) || ((~W_DIRECTION) && ((adj_dly_wclk_del[6:0] == 7'd127)||(adj_dly_wclk_del[7])));

wire [255:0] wclk_del_delay_chain;
wire wclk_del_source;

assign wclk_del_source = (DDC_MODE == "FULL_RATE") ? CLKB : ioclk_gated;

always @(*)
begin
    wclk_del_source_dly <= #0.2 wclk_del_source;
end 
    
assign wclk_del_delay_chain[0] = wclk_del_source_dly;
genvar gen_j;
generate  
    for(gen_j=1;gen_j<256;gen_j=gen_j+1) 
    begin
        assign #0.025 wclk_del_delay_chain[gen_j] =  wclk_del_delay_chain[gen_j-1];
    end
endgenerate

assign WCLK_DEL_TMP = ~(adj_dly_wclk_del[7] ?  wclk_del_delay_chain[127] : wclk_del_delay_chain[adj_dly_wclk_del]);
assign WCLK_DELAY = (WCLK_DELAY_SEL == "TRUE") ? ~WCLK_DEL_TMP : WCLK_DEL_TMP;

wire clk_r270;

assign clk_r270 = ~(DLL_STEP_WCLK_DEL[7] ? wclk_del_delay_chain[127] : wclk_del_delay_chain[DLL_STEP_WCLK_DEL]);

always @(posedge CLKB or negedge global_rstn or negedge lsr_rstn)
begin
    if (!global_rstn) 
    begin
        DQS_GATE_CTRL_d1 <= 0;
        DQS_GATE_CTRL_d2 <= 0;
    end
    else if (!lsr_rstn) 
    begin
        DQS_GATE_CTRL_d1 <= 0;
        DQS_GATE_CTRL_d2 <= 0;
    end
    else 
    begin
        if (DDC_MODE == "QUAD_RATE")
            DQS_GATE_CTRL_d2 <= DQS_GATE_CTRL;
        else 
        begin
            DQS_GATE_CTRL_d1 <= DQS_GATE_CTRL;
            DQS_GATE_CTRL_d2 <= DQS_GATE_CTRL_d1;   
        end
    end
end
assign WCLK_sel = (DDC_MODE == "FULL_RATE") ? CLKB :  clk_r0;

always @(posedge WCLK_sel or negedge global_rstn or negedge lsr_rstn)
begin
    if (!global_rstn) 
    begin
        cnt <= 0;
    end
    else if (!lsr_rstn) 
    begin
        cnt <= 0;
    end
    else 
    begin
      cnt <= cnt + 1;
    end
end

assign capture = (DDC_MODE == "HALF_RATE") ? (~cnt[0]) : cnt == 3;

always @(posedge WCLK_sel or negedge global_rstn or negedge lsr_rstn)
begin
    if (!global_rstn)
        DQS_GATE_CTRL_d3 <= 0;
    else if (!lsr_rstn)
        DQS_GATE_CTRL_d3 <= 0;
    else if (capture)
        DQS_GATE_CTRL_d3 <= DQS_GATE_CTRL_d2;
end
assign #0.2 DQS_GATE_CTRL_d3_d = DQS_GATE_CTRL_d3;
assign #0.2 DQS_GATE_CTRL_d2_d = DQS_GATE_CTRL_d2[0];

always @(posedge WCLK_sel or negedge global_rstn or negedge lsr_rstn)
begin
    if (!global_rstn) 
    begin
        gate_st       <= 0;
        gate_cnt      <= 0;
    end
    else if (!lsr_rstn) 
    begin
        gate_st       <= 0;
        gate_cnt      <= 0;
    end
    else 
    begin
        gate_st       <= 1;
        if (gate_st)
            gate_cnt   <= gate_cnt + 1;
    end
end

assign shift = R_EXTEND == "TRUE" ? ((DDC_MODE == "HALF_RATE") ? gate_cnt[0] : (gate_cnt == 2)) :
                 ((DDC_MODE == "HALF_RATE") ? ~gate_cnt[0] : (gate_cnt == 1));

always @(posedge WCLK_sel or negedge global_rstn or negedge lsr_rstn)
begin
    if (!global_rstn)
        DQS_GATE_CTRL_d4 <= 0;
    else if (!lsr_rstn)
        DQS_GATE_CTRL_d4 <= 0;
    else if (shift)
        DQS_GATE_CTRL_d4 <= DQS_GATE_CTRL_d3_d;     
    else
        DQS_GATE_CTRL_d4 <= {1'b0, DQS_GATE_CTRL_d4[3:1]};
end

always @(posedge WCLK_sel or negedge global_rstn or negedge lsr_rstn)
begin
    if (!global_rstn) 
    begin
        DQS_GATE_CTRL_d5 <= 0;
        DQS_GATE_CTRL_d6 <= 0;
    end
    else if (!lsr_rstn) 
    begin
        DQS_GATE_CTRL_d5 <= 0;
        DQS_GATE_CTRL_d6 <= 0;
    end   
    else 
    begin     
        DQS_GATE_CTRL_d5 <= DQS_GATE_CTRL_d4[0];
        if (DDC_MODE == "FULL_RATE")
            DQS_GATE_CTRL_d6 <= DQS_GATE_CTRL_d2_d;
        else
            DQS_GATE_CTRL_d6 <= DQS_GATE_CTRL_d5;
    end
end

always @(READ_CLK_CTRL or WCLK_sel or clk_r270) 
begin
    case (READ_CLK_CTRL[1:0])
        2'd0: sel_gate_clk = ~clk_r270;
        2'd1: sel_gate_clk = ~ WCLK_sel;
        2'd2: sel_gate_clk = clk_r270;
        2'd3: sel_gate_clk = WCLK_sel;
    endcase
end
assign #0.2 DQS_GATE_CTRL_d6_d = DQS_GATE_CTRL_d6;
assign #0.4 DQS_GATE_CTRL_d2_dd = DQS_GATE_CTRL_d2[0];
assign #0.2 DQS_GATE_CTRL_d5_d = DQS_GATE_CTRL_d5;

always @(posedge sel_gate_clk or negedge global_rstn or negedge lsr_rstn)
begin
    if (!global_rstn)
        DQS_GATE_CTRL_comb_d1 <= 0;
    else if (!lsr_rstn)
        DQS_GATE_CTRL_comb_d1 <= 0;
    else 
    begin
        if (READ_CLK_CTRL[2])
            DQS_GATE_CTRL_comb_d1 <= DQS_GATE_CTRL_d6_d;
        else if (DDC_MODE == "FULL_RATE")
            DQS_GATE_CTRL_comb_d1 <= DQS_GATE_CTRL_d2_dd;
        else   
            DQS_GATE_CTRL_comb_d1 <= DQS_GATE_CTRL_d5_d;
    end
end

always @(negedge sel_gate_clk or negedge global_rstn or negedge lsr_rstn)
begin
    if (!global_rstn)
        DQS_GATE_CTRL_comb_d2 <= 0;
    else if (!lsr_rstn)
        DQS_GATE_CTRL_comb_d2 <= 0;
    else
        DQS_GATE_CTRL_comb_d2 <= DQS_GATE_CTRL_comb_d1;
end

assign dqs_gate_ctrl_comb = (GATE_SEL=="TRUE")? DQS_GATE_CTRL_comb_d1 & DQS_GATE_CTRL_comb_d2 : GATE_IN;
assign GATE_OUT = DQS_GATE_CTRL_comb_d1 & DQS_GATE_CTRL_comb_d2;

assign set_en = lsr_rstn&RST_TRAINING_N&dqs_gate_ctrl_comb;

always @(negedge DQSIN_gated or negedge global_rstn or negedge lsr_rstn or negedge RST_TRAINING_N or posedge set_en)
begin
    if (!global_rstn)
        DQS_GATE_CTRL_gate <= 1'b0;
    else if (!lsr_rstn)
        DQS_GATE_CTRL_gate <= 1'b0;
    else if (!RST_TRAINING_N)
        DQS_GATE_CTRL_gate <= 1'b0;
    else if (set_en)
        DQS_GATE_CTRL_gate <= 1'b1;
    else
        DQS_GATE_CTRL_gate <= 1'b0;
end

assign DQSIN_gated = DQS_GATE_CTRL_gate & DQSI;

assign saout   = dqs_gate_ctrl_comb ? out : 1'b1;
assign saout_b = dqs_gate_ctrl_comb ? ~out: 1'b1;

always@(posedge dqs_gate_ctrl_comb)
begin
    if(dqs_gate_ctrl_comb)
    begin
        case ({DQSI,~DQSI})
            2'b10 : out = 1'b1;
            2'b01 : out = 1'b0;
            2'b11 : out = 1'bx;
            default : out = 1'bx;
        endcase
    end else
        out = 1'bz;
end

assign drift_status_0 = ~(saout&lsr_rstn&global_rstn&drift_status_1);
assign drift_status_1 = ~(saout_b&lsr_rstn&global_rstn&drift_status_0);
assign dqs_drift_status = ~drift_status_0;

assign DQS_DRIFT_STATUS = dqs_drift_status;

always @(posedge DQSIN_gated or negedge global_rstn or negedge lsr_rstn)
begin
    if(!global_rstn)
        q <= 4'b0;
    else if(!lsr_rstn)
        q <= 4'b0;
    else
        q <= {~clk_r270, ~WCLK_sel, clk_r270, WCLK_sel};
end

always @(posedge DQSIN_gated or negedge global_rstn or negedge lsr_rstn)
begin
    if(!global_rstn)
    begin
        dqs_drift_reg <= 2'b0;
        drift_detect_err_reg <= 1'b0;
    end
    else if(!lsr_rstn)
    begin
        dqs_drift_reg <= 2'b0;
        drift_detect_err_reg <= 1'b0;
    end
    else if((q == 4'b0001)||(q == 4'b1001)||(q == 4'b1101))
    begin
        dqs_drift_reg <= 2'b00;
        drift_detect_err_reg <= 1'b0;
    end
    else if((q == 4'b1100)||(q == 4'b1110)||(q == 4'b1000))
    begin
        dqs_drift_reg <= 2'b01;
        drift_detect_err_reg <= 1'b0;
    end
    else if((q == 4'b0100)||(q == 4'b0110)||(q == 4'b0111))
    begin
        dqs_drift_reg <= 2'b11;
        drift_detect_err_reg <= 1'b0;
    end
    else if((q == 4'b0011)||(q == 4'b0010)||(q == 4'b1011))
    begin
        dqs_drift_reg <= 2'b10;
        drift_detect_err_reg <= 1'b0;
    end
    else if(q == 4'b0000)
    begin
        dqs_drift_reg <= dqs_drift_reg;
        drift_detect_err_reg <= 1'b0;
    end
    else
        drift_detect_err_reg <= 1'b1;
end

assign DQS_DRIFT = dqs_drift_reg;
assign DRIFT_DETECT_ERR = drift_detect_err_reg;

wire [7:0] DLL_STEP_tmp = R_DELAY_STEP_EN == "TRUE" ? DELAY_STEP1 :8'd0;
wire RDEL_CTRL_b0_tmp = R_MOVE_EN == "TRUE" ? R_LOAD_N : 1'b1;

wire [8:0] DQSI_DEL_OFFSET_tmp = DQSI_DELAY_OFFSET;

//wire [7:0] tmp_dqsi_del = DQSI_DEL_OFFSET_tmp[8] ? (DLL_STEP_tmp - DQSI_DEL_OFFSET_tmp[7:0]) : (DLL_STEP_tmp + DQSI_DEL_OFFSET_tmp[7:0]);
wire [7:0] tmp_dqsi_del = (DLL_STEP_tmp + DQSI_DEL_OFFSET_tmp[7:0]);

wire tmp_dqsi_del_co_0 = DLL_STEP_tmp[0] && DQSI_DEL_OFFSET_tmp[0];
wire tmp_dqsi_del_co_1 = (DLL_STEP_tmp[1] && DQSI_DEL_OFFSET_tmp[1]) || ((DLL_STEP_tmp[1] || DQSI_DEL_OFFSET_tmp[1]) && tmp_dqsi_del_co_0);
wire tmp_dqsi_del_co_2 = (DLL_STEP_tmp[2] && DQSI_DEL_OFFSET_tmp[2]) || ((DLL_STEP_tmp[2] || DQSI_DEL_OFFSET_tmp[2]) && tmp_dqsi_del_co_1);
wire tmp_dqsi_del_co_3 = (DLL_STEP_tmp[3] && DQSI_DEL_OFFSET_tmp[3]) || ((DLL_STEP_tmp[3] || DQSI_DEL_OFFSET_tmp[3]) && tmp_dqsi_del_co_2);
wire tmp_dqsi_del_co_4 = (DLL_STEP_tmp[4] && DQSI_DEL_OFFSET_tmp[4]) || ((DLL_STEP_tmp[4] || DQSI_DEL_OFFSET_tmp[4]) && tmp_dqsi_del_co_3); 
wire tmp_dqsi_del_co_5 = (DLL_STEP_tmp[5] && DQSI_DEL_OFFSET_tmp[5]) || ((DLL_STEP_tmp[5] || DQSI_DEL_OFFSET_tmp[5]) && tmp_dqsi_del_co_4);
wire tmp_dqsi_del_co_6 = (DLL_STEP_tmp[6] && DQSI_DEL_OFFSET_tmp[6]) || ((DLL_STEP_tmp[6] || DQSI_DEL_OFFSET_tmp[6]) && tmp_dqsi_del_co_5);
wire tmp_dqsi_del_co_7 = (DLL_STEP_tmp[7] && DQSI_DEL_OFFSET_tmp[7]) || ((DLL_STEP_tmp[7] || DQSI_DEL_OFFSET_tmp[7]) && tmp_dqsi_del_co_6);


assign tmp_dqsi_del_sel= ~(DQSI_DEL_OFFSET_tmp[8] ^ tmp_dqsi_del_co_7);
wire [7:0] adj_dly_dqsi_tmp = DQSI_DEL_OFFSET_tmp[8] ? (tmp_dqsi_del_sel ?  tmp_dqsi_del[7:0] : 8'd0) :
                              (tmp_dqsi_del_sel ? tmp_dqsi_del[7:0] : 8'd255);

always @(*) 
begin
    if (RDEL_CTRL_b0_tmp)
        adj_dly_dqsi <= adj_dly_dqsi_tmp;
end

always @(*)
begin
    r_move_enable <= #3 R_MOVE&(~RDELAY_OB);
end

always @(negedge R_MOVE)
begin
    if (RDEL_CTRL_b0_tmp)
        adj_dly_dqsi <= adj_dly_dqsi_tmp;
    else if(r_move_enable)
    begin 
        if (R_DIRECTION && (adj_dly_dqsi != 8'd0))
            adj_dly_dqsi <= adj_dly_dqsi - 1;
        else if ((~R_DIRECTION) && (adj_dly_dqsi[6:0] != 7'd127)&&(~adj_dly_dqsi[7]))
            adj_dly_dqsi <= adj_dly_dqsi + 1;
    end
end

assign RDELAY_OB = (R_DIRECTION && (adj_dly_dqsi == 8'd0)) || ((~R_DIRECTION) && ((adj_dly_dqsi[6:0] == 7'd127)||(adj_dly_dqsi[7])));

wire [255:0] dqsi_delay_chain;

always @(*)
begin
    dqsin_gated_dly <= #0.2 DQSIN_gated;
end

assign dqsi_delay_chain[0] = dqsin_gated_dly;
genvar gen_k;
generate  
    for(gen_k=1;gen_k<256;gen_k=gen_k+1) 
    begin
        assign #0.025 dqsi_delay_chain[gen_k] =  dqsi_delay_chain[gen_k-1];
    end
endgenerate

assign DQSI_DELAY = adj_dly_dqsi[7] ? dqsi_delay_chain[127] : dqsi_delay_chain[adj_dly_dqsi];


assign #0.2 DQS_GATE_CTRL_comb_d1_dly = DQS_GATE_CTRL_comb_d1;
assign DQS_GATE_CTRL_comb_d1_rising = DQS_GATE_CTRL_comb_d1 & (~DQS_GATE_CTRL_comb_d1_dly);
assign #0.1 DQS_GATE_CTRL_gate_dly = DQS_GATE_CTRL_gate;

always @(posedge DQSIN_gated or posedge DQS_GATE_CTRL_comb_d1_rising or negedge global_rstn or negedge lsr_rstn or negedge RST_TRAINING_N)
begin
    if (!global_rstn)
        DQS_GATE_CTRL_gate_d <= 2'b0;
    else if (!lsr_rstn)
        DQS_GATE_CTRL_gate_d <= 2'b0;
    else if (!RST_TRAINING_N)
        DQS_GATE_CTRL_gate_d <= 2'b0;
    else if (DQS_GATE_CTRL_comb_d1_rising)
        DQS_GATE_CTRL_gate_d <= 2'b0;
    else if (DQS_GATE_CTRL_gate_dly) 
    begin
        DQS_GATE_CTRL_gate_d <= DQS_GATE_CTRL_gate_d + 1;
    end
end

always @(negedge DQSIN_gated or posedge DQS_GATE_CTRL_comb_d1_rising or negedge global_rstn or negedge lsr_rstn or negedge RST_TRAINING_N)
begin
    if (!global_rstn)
        DQS_GATE_CTRL_gate_dd <= 2'b0;
    else if (!lsr_rstn)
        DQS_GATE_CTRL_gate_dd <= 2'b0;
    else if (!RST_TRAINING_N)
        DQS_GATE_CTRL_gate_dd <= 2'b0;
    else if (DQS_GATE_CTRL_comb_d1_rising)
        DQS_GATE_CTRL_gate_dd <= 2'b0;
    else
    begin
        DQS_GATE_CTRL_gate_dd <= DQS_GATE_CTRL_gate_dd + 1;
    end
end

always @(negedge DQSIN_gated or posedge DQS_GATE_CTRL_comb_d1_rising or negedge global_rstn or negedge lsr_rstn or negedge RST_TRAINING_N)
begin
    if (!global_rstn)
        DQS_GATE_CTRL_comb_and_d <= 2'b0;
    else if (!lsr_rstn)
        DQS_GATE_CTRL_comb_and_d <= 2'b0;
    else if (!RST_TRAINING_N)
        DQS_GATE_CTRL_comb_and_d <= 2'b0;
    else if (DQS_GATE_CTRL_comb_d1_rising)
        DQS_GATE_CTRL_comb_and_d <= 2'b0;
    else if (dqs_gate_ctrl_comb) 
    begin
        DQS_GATE_CTRL_comb_and_d <= DQS_GATE_CTRL_comb_and_d + 1;
    end
end

assign DGTS_a = (~DQS_GATE_CTRL_gate_dly) && (DQS_GATE_CTRL_gate_d == 2'b00);
assign DGTS_b = (DQS_GATE_CTRL_gate_dd == 2'b00) &&  (DQS_GATE_CTRL_comb_and_d == 2'b11);

assign DGTS = DGTS_a & DGTS_b;


always @(posedge DQSI_DELAY or negedge rstn_fifo)
begin
    if (!rstn_fifo)
        start_wr <= 0;
    else
        start_wr <= rstn_fifo;
end

assign start_wr_comb = (IFIFO_GENERIC == "TRUE") ?  start_wr : rstn_fifo;

always @(posedge DQSI_DELAY or negedge start_wr_comb)
begin
    if (!start_wr_comb)
        WADDR_reg <= 0;
    else 
    begin
        case (WADDR_reg)
            3'b000: WADDR_reg <= 3'b001;
            3'b001: WADDR_reg <= 3'b011;
            3'b011: WADDR_reg <= 3'b010;
            3'b010: WADDR_reg <= 3'b110;
            3'b110: WADDR_reg <= 3'b111;
            3'b111: WADDR_reg <= 3'b101;
            3'b101: WADDR_reg <= 3'b100;
            3'b100: WADDR_reg <= 3'b000;
        endcase
    end
end

always @(negedge DQSI_DELAY or negedge start_wr_comb)
begin
    if (!start_wr_comb)
        IFIFO_WADDR_reg <= 0;
    else
        IFIFO_WADDR_reg <= WADDR_reg;
end

assign IFIFO_WADDR = IFIFO_WADDR_reg;

assign rd_clk = (DDC_MODE == "FULL_RATE") ? CLKB : CLKA;

always @(posedge rd_clk or negedge rstn_fifo)
begin
    if (!rstn_fifo)
        start_rd <= 0;
    else
        start_rd <= rstn_fifo;
end

always @(posedge rd_clk or negedge rst_start_rd)
begin
    if (!rst_start_rd)
        WADDR_reg_d1 <= 3'd0;
    else
        WADDR_reg_d1 <= WADDR_reg;
end

always @(posedge rd_clk or negedge rst_start_rd)
begin
    if (!rst_start_rd)
        WADDR_reg_d2 <= 3'd0;
    else
        WADDR_reg_d2 <= WADDR_reg_d1;
end

assign buffer_empty = WADDR_reg_d2 == RADDR_reg;
assign buffer_almost_empty = WADDR_reg_d2 == RADDR_reg_plus1;


always @(posedge rd_clk or negedge rst_transfer_n)
begin
    if (!rst_transfer_n) 
    begin
        new_st         <= 0;
        new_cnt        <= 0;
        new_transfer_d <= 0;
    end
    else 
    begin
        new_st       <= 1;
        if (new_st)
            new_cnt      <= new_cnt + 1;
            new_transfer_d <= new_transfer;
    end
end

always @(posedge rd_clk or negedge rst_transfer_n)
begin
    if (!rst_transfer_n)
    begin
        new_cnt_reg <= 1'b0;
    end
    else
    begin
        new_cnt_reg <= new_cnt[0];
    end
end

assign  new_transfer =  (DDC_MODE == "HALF_RATE") ? new_cnt_reg : (new_cnt == 2);

always @(posedge rd_clk or negedge rst_start_rd)
begin
    if (!rst_start_rd) 
    begin
        new_rd_en_reg <= 0;
    end
    else if ((DDC_MODE == "FULL_RATE") || new_transfer) 
    begin //sel port
        if (new_rd_en_reg) 
        begin
            if (buffer_almost_empty)
                new_rd_en_reg <= 1'b0;
        end
        else 
        begin
            if (~buffer_empty)
                new_rd_en_reg <= 1'b1;
        end
    end
end

wire read_enable = (new_rd_en_reg && (~buffer_empty)) || (IFIFO_GENERIC == "TRUE");

wire start_generic_read = (IFIFO_GENERIC == "TRUE") ? new_st : (~buffer_empty);


always @(posedge rd_clk or negedge rst_start_rd)
begin
    if (!rst_start_rd)
        RADDR_reg <= RADDR_INIT;
    else if (read_enable && start_generic_read) 
    begin
        case (RADDR_reg)
            3'b000: RADDR_reg <= 3'b001;
            3'b001: RADDR_reg <= 3'b011;
            3'b011: RADDR_reg <= 3'b010;
            3'b010: RADDR_reg <= 3'b110;
            3'b110: RADDR_reg <= 3'b111;
            3'b111: RADDR_reg <= 3'b101;
            3'b101: RADDR_reg <= 3'b100;
            3'b100: RADDR_reg <= 3'b000;
        endcase
    end
end

always @(*) 
begin
    case (RADDR_reg)
        3'b000: RADDR_reg_plus1 <= 3'b001;
        3'b001: RADDR_reg_plus1 <= 3'b011;
        3'b011: RADDR_reg_plus1 <= 3'b010;
        3'b010: RADDR_reg_plus1 <= 3'b110;
        3'b110: RADDR_reg_plus1 <= 3'b111;
        3'b111: RADDR_reg_plus1 <= 3'b101;
        3'b101: RADDR_reg_plus1 <= 3'b100;
        3'b100: RADDR_reg_plus1 <= 3'b000;
    endcase
end

assign IFIFO_RADDR = RADDR_reg;

always @(posedge rd_clk or negedge rst_start_rd)
begin
    if (!rst_start_rd) 
    begin
        read_enable_d1 <= 0;
        read_enable_d2 <= 0;
    end
    else 
    begin
        read_enable_d1 <= (new_rd_en_reg && (~buffer_empty));
        if (new_transfer_d)
            read_enable_d2 <= read_enable_d1;
    end
end

always @(posedge CLKB or negedge rst_start_rd)
begin
    if (!rst_start_rd)
        RDVALID_reg <= 0;
    else if (DDC_MODE == "FULL_RATE") 
    begin
        if (IFIFO_GENERIC == "TRUE")
            RDVALID_reg <= 1'b1;
        else
            RDVALID_reg <=  (new_rd_en_reg && (~buffer_empty));
    end
    else 
        RDVALID_reg <= read_enable_d2;
end

assign READ_VALID = RDVALID_reg;
//synthesis translate_on

endmodule





































//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_PREADD_MULTACC9.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

//P = MAC + (A*(B+C))
`timescale 1 ns / 1 ps

module GTP_PREADD_MULTACC9 #(
    parameter GRS_EN            = "TRUE", //"TRUE"; "FALSE"
    parameter SYNC_RST          = "FALSE", //"TRUE"; "FALSE"
    parameter INREG_EN          = "FALSE",  //"TRUE"; "FALSE"
    parameter PREREG_EN         = "FALSE",  //"TRUE"; "FALSE"
    parameter PIPEREG_EN        = "FALSE",   //"TRUE"; "FALSE"
    parameter ACC_ADDSUB_OP     = 0,
    parameter DYN_ACC_ADDSUB_OP = 1,     //Select parameter ADDSUB or input ADDSUB
    parameter OVERFLOW_MASK     = 32'h0, //32 OVERflow setting= 'h1_0000_0000, bit width = 32
    parameter PATTERN           = 32'h0, //compare pattern
    parameter MASKPAT           = 32'h0, //pattern mask
    parameter ACC_INIT_VALUE    = 32'h0  //ACC_INIT_VALUE value
) (
    output  [31:0] P,
    output  OVER,
    output  UNDER,
    output  EQZ,
    output  EQZM,
    output  EQOM,
    output  EQPAT,
    output  EQPATN,

    input   CE,
    input   RST,
    input   CLK,
    input   [8:0] A,
    input   [7:0] B,
    input   A_SIGNED,
    input   B_SIGNED,
    input   C_SIGNED,
    input   [7:0] C,
    input   PREADDSUB,
    input   ACC_ADDSUB,
    input   RELOAD
);

    wire [31:0] R;

    INT_PREADD_MULTACC #(
        . GRS_EN(GRS_EN),      
        . SYNC_RST(SYNC_RST),    
        . INREG_EN(INREG_EN),    
        . PREREG_EN(PREREG_EN),    
        . PIPEREG_EN(PIPEREG_EN),  
        . ACCUMADDSUB_OP(ACC_ADDSUB_OP), 
        . DYN_OP_SEL(DYN_ACC_ADDSUB_OP),    
        . ASIZE(9), 
        . BSIZE(8), 
        . PSIZE(32), 
        . MASK(OVERFLOW_MASK),     
        . DYN_ACC_INIT(0),
        . ACC_INIT_VALUE(ACC_INIT_VALUE)
    ) U_MACC (
        . CE(CE),
        . RST(RST),
        . CLK(CLK),
        . A(A),
        . B(B),
        . A_SIGNED(A_SIGNED),
        . B_SIGNED(B_SIGNED),
        . C_SIGNED(C_SIGNED),
        . C(C),
        . PREADDSUB(PREADDSUB),
        . ACCUM_INIT(32'b0),
        . ACCUMADDSUB(ACC_ADDSUB),
        . RELOAD(RELOAD),
        . P(P),
        . OVER(OVER),
        . UNDER(UNDER),
        . R(R)
    );

    INT_FLAG #(
        . GRS_EN(GRS_EN),
        . SYNC_RST(SYNC_RST),
        . PSIZE(32),
        . PATSIZE(32),
        . MASKPATSIZE(32),
        . OUTREG_EN("TRUE")
    ) U_FLAG (
        . CE(CE),
        . RST(RST),
        . CLK(CLK),
        . P(P),
        . PATTERN(PATTERN),
        . MASKPAT(MASKPAT),
        . OVERFLOW_MASK(OVERFLOW_MASK),
        . R(R),
        . eqz(EQZ),
        . eqzm(EQZM),
        . eqom(EQOM),
        . eqpat(EQPAT),
        . eqpatn(EQPATN)
    );

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_ODDR.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//2017/12/21 : initial version
//2018/01/02 : update due to software feedback
//2018/04/09 : change SYNC_RS to RS_TYPE
//2018/04/24 : change default value of GRS_EN to "TRUE"
/////////////////////////////////////////////////////////////////////////////
module GTP_ODDR #(
parameter GRS_EN   = "TRUE",        //"FALSE", "TRUE"
parameter RS_TYPE  = "ASYNC_SET"      //"ASYNC_SET", "ASYNC_RESET", "SYNC_SET", "SYNC_RESET"
) (

output Q,
input  D0,
input  D1,
input  CE,
input  RS,
input  CLK
); /* synthesis syn_black_box */

//synthesis translate_off

reg ce_reg;
reg q_reg0;
reg q_reg1;
reg q_reg2;

wire global_rsn;
wire global_rstn;
wire global_setn;
wire local_rst_async;
wire local_set_async; 
wire local_rst_sync;
wire local_set_sync; 
wire rstn_async;
wire setn_async;
wire rstn_sync;
wire setn_sync;
wire clk_gated;

initial begin
    if(GRS_EN != "TRUE" && GRS_EN != "FALSE")
    begin
      $display("GTP_IDDR Error: Illegal setting of GRS_EN %s",GRS_EN);
      $finish;
    end
    if(RS_TYPE != "ASYNC_SET" && RS_TYPE != "ASYNC_RESET" && RS_TYPE != "SYNC_SET" && RS_TYPE != "SYNC_RESET")
    begin
      $display("GTP_IDDR Error: Illegal setting of RS_TYPE %s",RS_TYPE);
      $finish;
    end
    ce_reg = 1'b0;
    q_reg0 = 1'b0;
    q_reg1 = 1'b0;
    q_reg2 = 1'b0;
end

//////////////////////////////////////////////////////////////////////
assign global_rsn  = (GRS_EN == "TRUE")    ? GRS_INST.GRSNET : 1'b1;

assign global_rstn = (RS_TYPE == "SYNC_SET" || RS_TYPE == "ASYNC_SET")   ? 1'b1 : global_rsn;
assign global_setn = (RS_TYPE == "SYNC_RESET" || RS_TYPE == "ASYNC_RESET") ? 1'b1 : global_rsn;


assign local_rst_async = (RS_TYPE == "ASYNC_RESET") ? RS : 1'b0;
assign local_set_async = (RS_TYPE == "ASYNC_SET")   ? RS : 1'b0;

assign local_rst_sync  = (RS_TYPE == "ASYNC_RESET" || RS_TYPE == "SYNC_RESET") ? RS : 1'b0;
assign local_set_sync  = (RS_TYPE == "ASYNC_SET" || RS_TYPE == "SYNC_SET")     ? RS : 1'b0;


assign rstn_async = global_rstn&(~local_rst_async);
assign setn_async = global_setn&(~local_set_async);

assign rstn_sync  = global_rstn&(~local_rst_sync);
assign setn_sync  = global_setn&(~local_set_sync);


always @(negedge CLK or negedge global_rsn)
begin
    if(!global_rsn)
        ce_reg <= 1'b0;
    else
        ce_reg <= CE;
end

assign clk_gated = ce_reg&CLK;

always @(posedge clk_gated or negedge setn_async or negedge rstn_async)
begin
    if(!(rstn_async&rstn_sync))
        q_reg0 <= 1'b0;
    else if(!(setn_async&setn_sync))
        q_reg0 <= 1'b1;
    else
        q_reg0 <= D0;
end

always @(posedge clk_gated or negedge setn_async or negedge rstn_async)
begin
    if(!(rstn_async&rstn_sync))
        q_reg1 <= 1'b0;
    else if(!(setn_async&setn_sync))
        q_reg1 <= 1'b1;    
    else
        q_reg1 <= D1;
end

always @(negedge clk_gated or negedge setn_async or negedge rstn_async)
begin
    if(!(rstn_async&rstn_sync))
        q_reg2 <= 1'b0;
    else if(!(setn_async&setn_sync))
        q_reg2 <= 1'b1;
    else
        q_reg2 <= q_reg1; 
end 

assign Q = clk_gated ? q_reg2 : q_reg0;

//synthesis translate_on
endmodule




































//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_RAM16X4DP.v
//
// Functional description: simple-dual-port 16x4 distributed ram
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_RAM16X4DP
#(
    parameter [15:0] INIT_0 = 16'h0000,
    parameter [15:0] INIT_1 = 16'h0000,
    parameter [15:0] INIT_2 = 16'h0000,
    parameter [15:0] INIT_3 = 16'h0000
) (
    output [3:0] DO,
    input [3:0] DI,
    input [3:0] RADDR, WADDR,
    input WCLK, WE
);

    reg [15:0] mem [3:0];

    initial begin
        mem[0] = INIT_0;
        mem[1] = INIT_1;
        mem[2] = INIT_2;
        mem[3] = INIT_3;
    end

    always @(posedge WCLK) begin
        if (WE == 1'b1) begin
            mem[0][WADDR] <= DI[0];
            mem[1][WADDR] <= DI[1];
            mem[2][WADDR] <= DI[2];
            mem[3][WADDR] <= DI[3];
        end
    end

    assign DO[0] = mem[0][RADDR];
    assign DO[1] = mem[1][RADDR];
    assign DO[2] = mem[2][RADDR];
    assign DO[3] = mem[3][RADDR];

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_PREADD_MULTACC36.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

//P = MAC + (A*(B+C))
`timescale 1 ns / 1 ps

module GTP_PREADD_MULTACC36 #(
    parameter GRS_EN            = "TRUE", //"TRUE"; "FALSE"
    parameter SYNC_RST          = "FALSE", //"TRUE"; "FALSE"
    parameter INREG_EN          = "FALSE",  //"TRUE"; "FALSE"
    parameter PREREG_EN         = "FALSE",  //"TRUE"; "FALSE"
    parameter PIPEREG_EN        = "FALSE",   //"TRUE"; "FALSE"
    parameter ACC_ADDSUB_OP     = 0,
    parameter DYN_ACC_ADDSUB_OP = 1,     //Select parameter ADDSUB or input ADDSUB
    parameter OVERFLOW_MASK     = 64'h0, //PSIZE = 64 OVERflow setting= 'h8000_0000_0000_0000, bit width = PSIZE
    parameter PATTERN           = 64'h0, //compare pattern
    parameter MASKPAT           = 64'h0, //pattern mask
    parameter ACC_INIT_VALUE    = 64'h0  //ACC_INIT_VALUE value
) (
    output  [63:0] P,
    output  OVER,
    output  UNDER,
    output  EQZ,
    output  EQZM,
    output  EQOM,
    output  EQPAT,
    output  EQPATN,

    input   CE,
    input   RST,
    input   CLK,
    input   [35:0] A,
    input   [17:0] B,
    input   A_SIGNED,
    input   B_SIGNED,
    input   C_SIGNED,
    input   [17:0] C,
    input   PREADDSUB,
    input   ACC_ADDSUB,
    input   RELOAD
);

    wire [63:0] R;

    INT_PREADD_MULTACC #(
        . GRS_EN(GRS_EN),      
        . SYNC_RST(SYNC_RST),    
        . INREG_EN(INREG_EN),    
        . PREREG_EN(PREREG_EN),    
        . PIPEREG_EN(PIPEREG_EN),  
        . ACCUMADDSUB_OP(ACC_ADDSUB_OP), 
        . DYN_OP_SEL(DYN_ACC_ADDSUB_OP),    
        . ASIZE(36), 
        . BSIZE(18), 
        . PSIZE(64), 
        . MASK(OVERFLOW_MASK),     
        . DYN_ACC_INIT(0),
        . ACC_INIT_VALUE(ACC_INIT_VALUE)
    ) U_MACC (
        . CE(CE),
        . RST(RST),
        . CLK(CLK),
        . A(A),
        . B(B),
        . A_SIGNED(A_SIGNED),
        . B_SIGNED(B_SIGNED),
        . C_SIGNED(C_SIGNED),
        . C(C),
        . PREADDSUB(PREADDSUB),
        . ACCUM_INIT(64'b0),
        . ACCUMADDSUB(ACC_ADDSUB),
        . RELOAD(RELOAD),
        . P(P),
        . OVER(OVER),
        . UNDER(UNDER),
        . R(R)
    );

    INT_FLAG #(
        . GRS_EN(GRS_EN),
        . SYNC_RST(SYNC_RST),
        . PSIZE(64),
        . PATSIZE(64),
        . MASKPATSIZE(64),
        . OUTREG_EN("TRUE")
    ) U_FLAG (
        . CE(CE),
        . RST(RST),
        . CLK(CLK),
        . P(P),
        . PATTERN(PATTERN),
        . MASKPAT(MASKPAT),
        . OVERFLOW_MASK(OVERFLOW_MASK),
        . R(R),
        . eqz(EQZ),
        . eqzm(EQZM),
        . eqom(EQOM),
        . eqpat(EQPAT),
        . eqpatn(EQPATN)
    );

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2016 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_RAM64X1SP.v
//
// Functional description: single-port 64x1 distributed ram
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_RAM64X1SP
#(
    parameter [63:0] INIT = 64'h0000_0000_0000_0000
) (
    output  DO,
    input   DI,
    input [5:0] ADDR,
    input WCLK, WE
);
//synthesis translate_off
    reg [63:0] mem ;

    initial begin
        mem = INIT;
    end

    always @(posedge WCLK) begin
        if (WE == 1'b1) begin
            mem[ADDR] <= DI;
        end
    end

    assign DO = mem[ADDR];
//synthesis translate_on
endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2016 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_IOCLKDIV_E2.v
//
// Functional description:
//
// Parameter description: DIV_FACTOR
//
// Port description:
//
// Revision:
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_IOCLKDIV_E2
#(
    parameter DIV_FACTOR = "BYPASS" //1, 2, 3, 4, 5, 6, 7, 8, BYPASS
) (
    output CLKDIVOUT,
    input CLKIN,
    input RST_N,
    input CE
);

//synthesis translate_off

    initial begin
        if (DIV_FACTOR != "BYPASS" && DIV_FACTOR != "1" && DIV_FACTOR != "2" && DIV_FACTOR != "3" && DIV_FACTOR != "4" && DIV_FACTOR != "5" && DIV_FACTOR != "6" && DIV_FACTOR != "7" && DIV_FACTOR != "8") begin
            $display("ERROR: The attribute DIV_FACTOR on instance %m is %s. Legal values are BYPASS or 1 or 2 or 3 or 4 or 5 or 6 or 7 or 8.", DIV_FACTOR);
            $finish;
        end
    end

    reg [3:0] div_mode;
    initial
    begin
        if(DIV_FACTOR == "BYPASS")
            div_mode=4'h0;
        else if(DIV_FACTOR == "1")
            div_mode=4'h1;
        else if(DIV_FACTOR == "2")
            div_mode=4'h2;
        else if(DIV_FACTOR == "3")
            div_mode=4'h3;
        else if(DIV_FACTOR == "4")
            div_mode=4'h4;
        else if(DIV_FACTOR == "5")
            div_mode=4'h5;
        else if(DIV_FACTOR == "6")
            div_mode=4'h6;
        else if(DIV_FACTOR == "7")
            div_mode=4'h7;
        else if(DIV_FACTOR == "8")
            div_mode=4'h8;
        else 
            div_mode=4'hx;
    end

    wire [3:0] idivider;
    wire div1;
    wire [3:0] duty_ctrl;
    wire clk_out_div;
    wire clk_out_mode;
    wire rst_n;
    reg rstn_idiv;
    reg [3:0] counter;
    reg clkdivr;
    reg div1_en;
    wire clk_in_div;
    
    assign idivider = div_mode;
    assign div1 = (idivider == 4'h1)?1:0;
    assign duty_ctrl = (idivider[0] == 1)?(idivider-1)>>1:idivider>>1;
    assign clk_out_div = (div1_en==1'b1)? clk_in_div:clkdivr;
    assign clk_out_mode = (idivider == 4'h0)? CLKIN:clk_out_div;
    assign CLKDIVOUT = clk_out_mode;
    assign rst_n = RST_N;
    assign clk_in_div  = CLKIN & CE;

    always @(posedge clk_in_div or negedge rst_n)
    begin
        if(!rst_n)
            rstn_idiv <= 1'b0;
        else
            rstn_idiv <= 1'b1;
    end 

    always @(posedge clk_in_div or negedge rstn_idiv)
    begin
        if(!rstn_idiv)
            counter <= 4'h0;
        else
        begin
            if(counter == idivider-1)
                counter <= 4'h0;
            else
                counter <= counter+1;
        end
    end

    always @(posedge clk_in_div or negedge rstn_idiv)
    begin
        if(!rstn_idiv)
            clkdivr <= 0;
        else
        begin
            if(counter < duty_ctrl)
                clkdivr <= 1;
            else 
                clkdivr <= 0;
        end
    end

    always @(posedge clk_in_div or negedge rstn_idiv)
    begin
        if(!rstn_idiv)
            div1_en <= 1'b0;
        else
        begin
            if(div1)
                div1_en <= 1'b1;
            else
                div1_en <= 1'b0;
        end
    end

      
//synthesis translate_on
endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_LUT3.v
//
// Functional description: 3-input Look-Up-Table
//
// Parameter description:
//      INIT: init value
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_LUT3
#(
    parameter [7:0] INIT = 8'h00
) (
    output wire Z,
    input wire I0, I1, I2
);

    wire x1, x0;

    INT_LUTMUX4_UDP (x1, I1, I0, INIT[7], INIT[6], INIT[5], INIT[4]);
    INT_LUTMUX4_UDP (x0, I1, I0, INIT[3], INIT[2], INIT[1], INIT[0]);
    INT_LUTMUX2_UDP (Z, I2, x1, x0);

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_PREADD_MULTACC27.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

//P = MAC + (A*(B+C))
`timescale 1 ns / 1 ps

module GTP_PREADD_MULTACC27 #(
    parameter GRS_EN            = "TRUE", //"TRUE"; "FALSE"
    parameter SYNC_RST          = "FALSE", //"TRUE"; "FALSE"
    parameter INREG_EN          = "FALSE",  //"TRUE"; "FALSE"
    parameter PREREG_EN         = "FALSE",  //"TRUE"; "FALSE"
    parameter PIPEREG_EN        = "FALSE",   //"TRUE"; "FALSE"
    parameter ACC_ADDSUB_OP     = 0,
    parameter DYN_ACC_ADDSUB_OP = 1,     //Select parameter ADDSUB or input ADDSUB
    parameter OVERFLOW_MASK     = 64'h0, //PSIZE = 64 OVERflow setting= 'h8000_0000_0000_0000, bit width = PSIZE
    parameter PATTERN           = 64'h0, //compare pattern
    parameter MASKPAT           = 64'h0, //pattern mask
    parameter ACC_INIT_VALUE    = 64'h0  //ACC_INIT_VALUE value
) (
    output  [63:0] P,
    output  OVER,
    output  UNDER,
    output  EQZ,
    output  EQZM,
    output  EQOM,
    output  EQPAT,
    output  EQPATN,

    input   CE,
    input   RST,
    input   CLK,
    input   [26:0] A,
    input   [25:0] B,
    input   A_SIGNED,
    input   B_SIGNED,
    input   C_SIGNED,
    input   [25:0] C,
    input   PREADDSUB,
    input   ACC_ADDSUB,
    input   RELOAD
);

    wire [63:0] R;

    INT_PREADD_MULTACC #(
        . GRS_EN(GRS_EN),      
        . SYNC_RST(SYNC_RST),    
        . INREG_EN(INREG_EN),    
        . PREREG_EN(PREREG_EN),    
        . PIPEREG_EN(PIPEREG_EN),  
        . ACCUMADDSUB_OP(ACC_ADDSUB_OP), 
        . DYN_OP_SEL(DYN_ACC_ADDSUB_OP),    
        . ASIZE(27), 
        . BSIZE(26), 
        . PSIZE(64), 
        . MASK(OVERFLOW_MASK),     
        . DYN_ACC_INIT(0),
        . ACC_INIT_VALUE(ACC_INIT_VALUE)
    ) U_MACC (
        . CE(CE),
        . RST(RST),
        . CLK(CLK),
        . A(A),
        . B(B),
        . A_SIGNED(A_SIGNED),
        . B_SIGNED(B_SIGNED),
        . C_SIGNED(C_SIGNED),
        . C(C),
        . PREADDSUB(PREADDSUB),
        . ACCUM_INIT(64'b0),
        . ACCUMADDSUB(ACC_ADDSUB),
        . RELOAD(RELOAD),
        . P(P),
        . OVER(OVER),
        . UNDER(UNDER),
        . R(R)
    );

    INT_FLAG #(
        . GRS_EN(GRS_EN),
        . SYNC_RST(SYNC_RST),
        . PSIZE(64),
        . PATSIZE(64),
        . MASKPATSIZE(64),
        . OUTREG_EN("TRUE")
    ) U_FLAG (
        . CE(CE),
        . RST(RST),
        . CLK(CLK),
        . P(P),
        . PATTERN(PATTERN),
        . MASKPAT(MASKPAT),
        . OVERFLOW_MASK(OVERFLOW_MASK),
        . R(R),
        . eqz(EQZ),
        . eqzm(EQZM),
        . eqom(EQOM),
        . eqpat(EQPAT),
        . eqpatn(EQPATN)
    );

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_PREADD_MULTADDSUM18.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

//P = (A0*(B0+/-C0) +/- A1*(B1 +/-C1)) +- (A2*(B2+/-C2) +/- A3*(B3+/-C3))
`timescale 1 ns / 1 ps

module GTP_PREADD_MULTADDSUM18  #(
    parameter GRS_EN             = "TRUE", //"TRUE"; "FALSE"
    parameter SYNC_RST           = "FALSE", //"TRUE"; "FALSE"
    parameter INREG_EN           = "FALSE",  //"TRUE"; "FALSE"
    parameter PREREG_EN          = "FALSE",  //"TRUE"; "FALSE"
    parameter PIPEREG_EN         = "FALSE",  //"TRUE"; "FALSE"
    parameter OUTREG_EN          = "FALSE",   //"TRUE"; "FALSE"
    parameter ADDSUB_OP          = 2'b00 ,
    parameter SUM_ADDSUB_OP      = 0 ,
    parameter DYN_ADDSUB_OP      = 2'b11,
    parameter DYN_SUM_ADDSUB_OP  = 1
)(
    output  [39-1:0] P,
    input   CE,
    input   RST,
    input   CLK,
    input   [1:0] A_SIGNED,
    input   [18-1:0] A0,
    input   [18-1:0] A1,
    input   [18-1:0] A2,
    input   [18-1:0] A3,
    input   [1:0] B_SIGNED,
    input   [1:0] C_SIGNED,
    input   [18-1:0] B0,
    input   [18-1:0] B1,
    input   [18-1:0] B2,
    input   [18-1:0] B3,
    input   [18-1:0] C0,
    input   [18-1:0] C1,
    input   [18-1:0] C2,
    input   [18-1:0] C3,
    input   [3:0] PREADDSUB,
    input   [1:0] ADDSUB,
    input   SUM_ADDSUB
);

    INT_PREADD_MULTADDSUM #(
        . GRS_EN(GRS_EN),    
        . SYNC_RST(SYNC_RST),  
        . INREG_EN(INREG_EN),  
        . PREREG_EN(PREREG_EN),
        . PIPEREG_EN(PIPEREG_EN),
        . OUTREG_EN(OUTREG_EN), 
        . ADDSUB_OP01(ADDSUB_OP[0]),  
        . ADDSUB_OP23(ADDSUB_OP[1]),  
        . ADDSUBSUM_OP(SUM_ADDSUB_OP), 
        . DYN_OP_SEL0(DYN_ADDSUB_OP[0]),
        . DYN_OP_SEL1(DYN_ADDSUB_OP[1]),
        . DYN_OP_SEL2(DYN_SUM_ADDSUB_OP),
        . ASIZE(18),
        . BSIZE(18)
    ) U_INT_PREADD_MULTADDSUM18 (
        . CE(CE),
        . RST(RST),
        . CLK(CLK),
        . A_SIGNED01(A_SIGNED[0]),
        . A_SIGNED23(A_SIGNED[1]),
        . A0(A0),
        . A1(A1),
        . A2(A2),
        . A3(A3),
        . B_SIGNED01(B_SIGNED[0]),
        . B_SIGNED23(B_SIGNED[1]), 
        . C_SIGNED01(C_SIGNED[0]),
        . C_SIGNED23(C_SIGNED[1]), 
        . B0(B0),
        . B1(B1),
        . B2(B2),
        . B3(B3),
        . C0(C0),
        . C1(C1),
        . C2(C2),
        . C3(C3),
        . PREADDSUB01(PREADDSUB[1:0]),
        . PREADDSUB23(PREADDSUB[3:2]),
        . ADDSUB01(ADDSUB[0]),
        . ADDSUB23(ADDSUB[1]),
        . ADDSUBSUM(SUM_ADDSUB),
        . P(P)
    );               

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_RAM16X4SP.v
//
// Functional description: single-port 16x4 distributed ram
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_RAM16X4SP
#(
    parameter [15:0] INIT_0 = 16'h0000,
    parameter [15:0] INIT_1 = 16'h0000,
    parameter [15:0] INIT_2 = 16'h0000,
    parameter [15:0] INIT_3 = 16'h0000
) (
    output [3:0] DO,
    input [3:0] DI,
    input [3:0] ADDR,
    input WCLK, WE
);

    reg [15:0] mem [3:0];

    initial begin
        mem[0] = INIT_0;
        mem[1] = INIT_1;
        mem[2] = INIT_2;
        mem[3] = INIT_3;
    end

    always @(posedge WCLK) begin
        if (WE == 1'b1) begin
            mem[0][ADDR] <= DI[0];
            mem[1][ADDR] <= DI[1];
            mem[2][ADDR] <= DI[2];
            mem[3][ADDR] <= DI[3];
        end
    end

    assign DO[0] = mem[0][ADDR];
    assign DO[1] = mem[1][ADDR];
    assign DO[2] = mem[2][ADDR];
    assign DO[3] = mem[3][ADDR];

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2017 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_OSC_E2.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1ns/10fs
module GTP_OSC_E2 #(
    parameter USER_DIV_EN  = "TRUE", // "TRUE", "FALSE"
    parameter CLK_DIV = 0       // 0~127
    )(

    input EN_N,
    output CLKOUT,
    output CLKCRC

    );

    // pragma translate_off
    reg user_en; 
    reg clk_532_reg; 
    reg [6:0] user_div_reg;
    reg [1:0] en_user;
    reg [6:0] cnt_user_reg;
    reg clk_out_reg;


    reg [1:0] en_sed;
    reg [6:0] cnt_sed_reg;
    reg clk_sed_reg;

    wire[6:0] div_ratio_user;

    initial
    begin


        if(USER_DIV_EN == "FALSE")
            user_en = 1'b0;
        else if(USER_DIV_EN == "TRUE")
            user_en = 1'b1;

        clk_532_reg = 1'b0;

        user_div_reg = CLK_DIV;
        en_user      = 2'b00;
        cnt_user_reg = 7'b000_0000;
        clk_out_reg = 1'b0;

        en_sed      = 2'b00;
        cnt_sed_reg = 7'b000_0000;
        clk_sed_reg = 1'b0;

    end
    ////////////////////////////////////////////////////////
    ////OSC_Analog_Core/////////////////////////////////////
    assign oscen = ~EN_N | en_user | en_sed[1];

    always begin
        wait (oscen == 1'b1)
        begin
            clk_532_reg = 1'b0;
            #0.94;
            clk_532_reg = 1'b1;
            #0.94;
        end
    end

    always begin
        wait (oscen != 1'b1)
        begin
            force clk_532_reg = 1'b0;
            #2 release clk_532_reg;
        end
    end
    ////////////////////////////////////////////////////////
    ////OSC_USER_DIVIDER////////////////////////////////////
    always @(negedge clk_out_reg)
    begin
        en_user <= {en_user[0], (~EN_N) & user_en};
    end

    assign rstn_user = ((~EN_N) & user_en) | en_user[1];

   assign div_ratio_user = (user_div_reg == 7'd1) ? 7'd2 : user_div_reg;

    always @(posedge clk_532_reg or negedge rstn_user)
    begin
        if (!rstn_user)
        begin
            cnt_user_reg <= 7'b000_0000;
            clk_out_reg <= 1'b0;
        end
        else 
            if(cnt_user_reg == div_ratio_user - 7'b1)
            begin
                cnt_user_reg <= 7'b000000;
                clk_out_reg <= ~clk_out_reg;
            end
            else
            begin
                cnt_user_reg <= cnt_user_reg + 1'b1;
                clk_out_reg <= clk_out_reg;
        end
    end

    assign CLKOUT = clk_out_reg;

    ////////////////////////////////////////////////////////
    ////OSC_SED_DIVIDER/////////////////////////////////////
    always @(negedge clk_sed_reg)
    begin
        en_sed <= {en_sed[0], ~EN_N};
    end

    assign rstn_sed = ~EN_N | en_sed[1];

    always @(posedge clk_532_reg or negedge rstn_sed)
    begin
        if (!rstn_sed)
        begin
            cnt_sed_reg <= 7'b000_0000;
            clk_sed_reg <= 1'b0;
        end
        else 
            if(cnt_sed_reg == 7'b111_1111)
            begin
                cnt_sed_reg <= 7'b000000;
                clk_sed_reg <= ~clk_sed_reg;
            end
            else
            begin
                cnt_sed_reg <= cnt_sed_reg + 1'b1;
                clk_sed_reg <= clk_sed_reg;
        end
    end

    assign CLKCRC = clk_sed_reg;

    // pragma translate_on
endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2016 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_IPAL_E1.v
//
// Functional description: the simulation model of configuration and readback
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_IPAL_E1
#(
    parameter     [31:0] IDCODE = 32'haaaa5555,
    parameter            DATA_WIDTH = "X8", //X8, X16, X32, Ipal data width select
    parameter            SIM_DEVICE = "PGL25G"
) (
    output        [31:0] DO,//Ipal data out
    output               RBCRC_ERR,//readback CRC error flag
    output               RBCRC_VALID,//readback CRC result valid
    output               ECC_VALID,//SEU result valid
    output        [11:0] ECC_INDEX,//address of single error bit
    output               SERROR,//single-bit error flag
    output               DERROR,//double-bit error flag
    output               BUSY,

    input                RST_N,
    input                CLK,// 50M system clock
    input                CS_N,// chip select to enable the pal data bus, active low
    input                RW_SEL,//Ipal rdw, 0: write, 1: read
    input        [31:0]  DI//Ipal data in
 
);

//synthesis translate_off

/////////////////////////////  Extra features //////////////////////


  reg        [7:0]  SEU_FRAME_ADDR;//current frame address of SEU
  reg        [7:0]  SEU_COLUMN_ADDR;//current column address of SEU
  reg        [4:0]  SEU_REGION_ADDR;//current region address of SEU
  reg    [7:0]  SEU_FRAME_NADDR;//next frame address of SEU
  reg    [7:0]  SEU_COLUMN_NADDR;//next column address of SEU
  reg    [4:0]  SEU_REGION_NADDR;//next region address of SEU
  wire               PRCFG_OVER;// Partial reconfiguration over pulse
  wire               PRCFG_ERR;// Partial reconfiguration error flag
  wire               DRCFG_OVER;
  wire               DRCFG_ERR;


////////////////////////////////////////////////////////////////////

    localparam          MEM_DEPTH = (SIM_DEVICE == "PGL25G") ? 3500 : 1616;
    localparam          HEADER       =  1'b0;
    localparam          DAT          =  1'b1;

    wire    [31:0]  data; //aligned 32-bit input data
    wire            data_valid;
    wire            flg_rcmem;
    wire            flg_read_tmp;
    wire            flg_write_tmp;
    wire            flg_type1;
    wire            flg_type2;
    wire    [26:0]  word_count_tmp;
    wire            flg_desync;
    wire            flg_prcfgen;
    wire            flg_prcfgdis;
    wire            flg_drcfgen;
    wire            flg_drcfgdis;
    wire            flg_rbcrc;
    wire            flg_rrbcrc;
    wire            rbcrc_en;
    wire            seu_en;
    wire            re_rb;
    wire            we;
    wire            flg_rb_reg;
    wire    [1:0]   cmemtype;
    wire    [4:0]   addr_region;
    wire    [7:0]   addr_column;
    wire    [7:0]   addr_frame;
    wire            region0;
    wire            region1;
    wire            region2;
    wire            region3;
    wire            serror;
    wire            derror;
    wire    [11:0]  index; 
    wire            cmemclk;
    wire            crc_err;
    wire            flg_rstcrc;
    wire            prcfg_err;
    wire            drcfg_err;
    


    reg     [31:0]  data_rb;
    reg     [1:0]   ipal_m;
    reg     [4:0]   regaddr;
    reg             flg_write;
    reg             flg_rb_cmem;
    reg             flg_rb_cmem_d;
    reg             s;
    reg             ns;
    reg     [26:0]  word_count;
    reg     [26:0]  word_count_rb;
    reg             prcfg_en;
    reg             prcfg_en_d;
    reg             prcfg_over;
    reg             drcfg_en; 
    reg             drcfg_en_d;   
    reg             drcfg_over;
    
    reg     [4:0]   reg_cmd;
    reg     [31:0]  data_rb_reg;  
    reg             serror_d;
    reg             derror_d;
  //  reg     [3231:0]cmem [0:7999];   
    reg      [2175:0] cmem [0:MEM_DEPTH-1]; // 2176:Number of bits in a frame  3500:The number of all frames 
    reg             [13:0] addr_row;
    reg             [13:0] naddr_row;
    reg             [6:0] addr_word;
    reg             flg_region_end;
    reg             flg_column_end;
    reg             flg_frame_end;


    reg     [31:0]  reg_crcr;
    reg     [31:0]  reg_idr;
    reg     [31:0]  reg_cmdr;
    reg     [31:0]  reg_ctrl0r;
    reg     [31:0]  reg_ctrl1r;
    reg     [31:0]  reg_cmemir;
    reg     [31:0]  reg_mfwriter;
    reg     [95:0]  reg_ivr;
    reg     [31:0]  reg_chainr;
    reg     [31:0]  reg_adrr;
    reg     [31:0]  reg_sbpir;
    reg     [31:0]  reg_seur;
    reg     [31:0]  reg_irstctrlr;
    reg     [31:0]  reg_irstadrr;
    reg     [31:0]  reg_watchdogr;
    reg     [31:0]  reg_cmaskr;
    reg     [255:0]  reg_keyr;
    reg     [31:0]  reg_option0r;
    reg     [31:0]  reg_option1r;
    reg     [31:0]  reg_rcrr;
    reg     [8383:0]  reg_autr;
    reg     [31:0]  reg_seuaddr;
    reg     [31:0]  reg_seunaddr;

    reg     [31:0]  reg_cmemor;
    reg     [31:0]  reg_statusr;
    reg     [31:0]  reg_seustatusr;
    reg     [31:0]  reg_hstatusr;
    reg     [31:0]  reg_adrr_seu;

    integer         i;

    //     read-write switch delay
    reg rws_flg;
    reg [7:0]rws_cnt;


///////////////////////////////////////////////////ISPAL/////////////////////////////////////////////////////////////

    initial begin
        case(DATA_WIDTH)
            "X8"  :  ipal_m = 2'd0;
            "X16" :  ipal_m = 2'd1;
            "X32" :  ipal_m = 2'd2;
          default :  begin
                     ipal_m = 2'd0;
                     $display("Setting Error : The DATA_WIDTH is set to %s. Legal values is X8,X16,X32",DATA_WIDTH);
                     $finish;                  
          end
        endcase
    end

   initial begin
        $readmemb("cmem.txt", cmem);  // read cmem.txt
   end


    ipal_e1_if_ispal CCS_IF_ISPAL (

        .rstn               (RST_N),
        .clk                (CLK), 
        .en                 (1'b1), 
        .m                  (ipal_m), 
        .din                (DI), 
        .cs_n               (CS_N), 
        .rdwr_n             (RW_SEL), 
        .flg_desync         (flg_desync),
        .data_rb            (data_rb), 
        .empty              (1'b0),

        .dout               (DO),
        .rws_flg            (rws_flg),  
        .data               (data), 
        .data_valid         (data_valid), 
        .re_rb              (re_rb));


/////////////////////////////////////// frame interval delay //////////////////////////////////////////

localparam FRAME_CNT_MAX = 68;
localparam DELAY_CNT_MAX = 8;
reg [7:0] frame_cnt;  //read back count: 0~67
reg [7:0] delay_cnt;  // frame interval delay: 8 CLK
reg       delay_flg;  // delay flag
reg [26:0]word_count_tmp_reg;  // latch number of write/read data

//    word_count_tmp_reg
always@(posedge CLK or negedge RST_N)
begin
    if(RST_N==0)
        word_count_tmp_reg <= 27'd0;
    else if(flg_type1==1&&flg_read_tmp==1)
        word_count_tmp_reg <= data[21:0];
    else if(flg_type2==1&&flg_read_tmp==1)
        word_count_tmp_reg <= data[26:0];
end

//    frame_flg
//always@(posedge CLK or negedge RST_N)
//begin
//    if(RST_N==0)
//        frame_flg <= 0;
//    else if(word_count_tmp_reg<FRAME_CNT_MAX)
//        frame_flg <= 0;
//    else if(word_count_tmp_reg>=FRAME_CNT_MAX) // a frame number
//        frame_flg <= 1;
//end

assign frame_flg = (word_count_tmp_reg>68)?1:0;
//    frame_cnt 
always@(posedge CLK or negedge RST_N)
begin
    if(RST_N==0)
        frame_cnt <= 8'd0;
    else if(delay_flg==1'b1) // frame interval delay
        frame_cnt <= frame_cnt;
    else if(frame_cnt == FRAME_CNT_MAX-1'b1&&flg_rb_cmem && re_rb)  // read back a frame
        frame_cnt <= 8'd0;
    else if(frame_flg==1&&rws_flg==0)  
        begin
            if(flg_rb_cmem==0)  // read back end
                frame_cnt <= 0;
            else if(flg_rb_cmem && re_rb) // continue read back start
                frame_cnt <= frame_cnt + 1'b1;
        end
end

//    delay_flg
always@(posedge CLK or negedge RST_N)
begin
    if(RST_N==0)
        delay_flg <= 1'b0;  
    else if(delay_cnt == DELAY_CNT_MAX-1'b1&&delay_flg==1'b1)  //delay 8 CLK
        delay_flg <= 1'b0;
    else if(frame_cnt == FRAME_CNT_MAX-1'b1&&flg_rb_cmem && re_rb) // 
        delay_flg <= 1'b1;
end

//    delay_cnt
always@(posedge CLK or negedge RST_N)
begin
    if(RST_N==0)
        delay_cnt <= 8'd0;
    else if(delay_cnt==DELAY_CNT_MAX-1'b1&&delay_flg==1'b1)
        delay_cnt <= 8'd0;
    else if(delay_flg==1'b1)
        delay_cnt <= delay_cnt + 1'b1;
end


//////////////////////////////////// BUSY  ///////////////////////////////////////

assign BUSY = (delay_flg==1||rws_flg==1)?1:0;


///////////////////////////// read-write switch delay ////////////////////////

localparam RWS_CNT_MAX = 16;

//reg rw_sel_reg; // latch RW_SEL
//always@(posedge CLK or negedge RST_N)
//begin
//    if(RST_N==0)
//       rw_sel_reg <= 0;
//    else if(CS_N==0)
//       rw_sel_reg <= RW_SEL; 
//end

//always@(posedge CLK or negedge RST_N)
//begin
//    if(RST_N==0)
//        rws_flg <= 0;
//    else if(rws_cnt==RWS_CNT_MAX-1&&rws_flg==1)
//        rws_flg <= 0;
//    else if((CS_N==1&&RW_SEL==1&&flg_rb_cmem==1)||(CS_N==0&&RW_SEL==1&&flg_rb_cmem==1))
//        rws_flg <= 1;
//end
reg data_valid_r;
always@(posedge CLK or negedge RST_N)
begin
    if(RST_N==0)
        data_valid_r <= 0;
    else 
        data_valid_r <= data_valid;
end
always@(*)
begin
    if(RST_N==0)
        rws_flg <= 0;
    else if(rws_cnt==RWS_CNT_MAX)
        rws_flg <= 0;
   // else if((word_count_rb==word_count_tmp-1)&&RW_SEL==1&&flg_rb_cmem==1&&CS_N==0)
   // else if((word_count_rb==word_count_tmp-1)&&RW_SEL==1&&flg_rb_cmem==1)
   // else if((word_count_rb==word_count_tmp-1)&&flg_type2==1)
      else if((word_count_rb==word_count_tmp-1)&&data_valid_r==1&&flg_type2==1&&flg_read_tmp==1) // package 2
        rws_flg <= 1;
end

//always@(posedge CLK or negedge RST_N)
//begin
//    if(RST_N==0)
//        rws_flg <= 0;
//    else if(rws_cnt==RWS_CNT_MAX-1)
//        rws_flg <= 0;
//    else if(data_valid==1&&flg_type2==1&&flg_read_tmp==1)
//        rws_flg <= 1;
//end

//  delay

//always@(posedge CLK or negedge RST_N)
//begin
//    if(RST_N==0)
//        rws_cnt <= 0;
//    else if(RW_SEL==0)
//        rws_cnt <= 0;
//    else if(rws_cnt==RWS_CNT_MAX)
//        rws_cnt <= rws_cnt;
//    else if(rws_flg==1)
//        rws_cnt <= rws_cnt + 1;
//end

always@(posedge CLK or negedge RST_N)
begin
    if(RST_N==0)
        rws_cnt <= 0;
    else if(rws_flg==0&&rws_cnt==RWS_CNT_MAX)
        rws_cnt <= 0;
//    else if(rws_cnt==RWS_CNT_MAX)
//        rws_cnt <= rws_cnt;
    else if(rws_flg==1)
        rws_cnt <= rws_cnt + 1;
end





////////////////////// data_rb ////////////////////


    always@(*) begin
        if(RW_SEL&&!CS_N) begin
            if(flg_rb_reg && !flg_rb_cmem)
                data_rb = data_rb_reg;
            else if(BUSY==1)
                data_rb = 32'hFFFF_FFFF;
            else if(flg_rb_cmem && !flg_rb_reg)
                data_rb = reg_cmemor;
            else 
                data_rb = 32'hFFFF_FFFF;
        end
        else begin
            data_rb = 32'hFFFF_FFFF;
        end
    end



///////////////////////////////packet processor////////////////////////////////////////

    assign flg_read_tmp   = (data_valid==1)?(data[28:27] == 2'b10):flg_read_tmp;
    assign flg_write_tmp  = (data_valid==1)?(data[28:27] == 2'b01):flg_write_tmp;
    assign flg_type1      = (data_valid==1)?(data[31:29] == 3'b101):flg_type1;
    assign flg_type2      = (data_valid==1)?(data[31:29] == 3'b010):flg_type2;
    assign word_count_tmp = (flg_type1==1&&data_valid==1)?{5'd0, data[21:0]} : data[26:0]; 
    assign flg_rb_reg = ~CS_N & RW_SEL & (~flg_rb_cmem);

//State machine to indicate HEADER or DATA for current data
    always @(posedge CLK or negedge RST_N)begin
        if(RST_N == 1'b0)
            s <= HEADER;
        else if(data_valid||re_rb)
            s <= ns;
    end

    always @(*) begin
        case(s)
            HEADER: begin
                if(((flg_type1 || flg_type2) && (flg_read_tmp || flg_write_tmp)) && (word_count_tmp != 27'd0))
                    ns = DAT;
                else
                    ns = HEADER;
            end

            DAT:  begin
                if((data_valid && (word_count == 27'd0)) || (re_rb && (word_count_rb == 27'd0)))
                    ns = HEADER;
                else
                    ns = DAT;
            end
        endcase
    end

//get address
    always @(posedge CLK or negedge RST_N) begin
        if(RST_N == 1'b0)
            regaddr <= 5'd0;
        else if((data_valid || re_rb) && (s == HEADER) && flg_type1 && (flg_read_tmp || flg_write_tmp))
            regaddr <= data[26:22];
    end

//write flag
    always @(posedge CLK or negedge RST_N) begin
        if(RST_N == 1'b0)
            flg_write <= 1'b0;
        else if(data_valid) begin
            if((s == HEADER) && (flg_type1 || flg_type2) && flg_write_tmp && (word_count_tmp != 27'd0))
                flg_write <= 1'b1;
            else if(word_count == 27'd0)
                flg_write <= 1'b0;
        end
    end

//write operation count
    always @(posedge CLK or negedge RST_N) begin
        if(RST_N == 1'b0)
            word_count <= 27'd0;
        else if(data_valid) begin
            if((s == HEADER) && (flg_type1 || flg_type2) && flg_write_tmp && (word_count_tmp != 27'd0))
                word_count <= word_count_tmp - 1'b1;
            else if((s == DAT) && (word_count != 27'd0))
                word_count <= word_count - 1'b1;
            else
                word_count <= 27'd0;
        end
    end

//cmem readback count
    always @(posedge CLK or negedge RST_N) begin   
        if(RST_N == 1'b0)
            word_count_rb <= 27'd0;
        else if(delay_flg==1)     // delay 8 CLK
            word_count_rb <= word_count_rb;
     //   else if(/*re_rb && */(s == HEADER) && (flg_type1 || flg_type2) && flg_read_tmp && (word_count_tmp != 27'd0) && flg_rcmem)
        else if(/*re_rb && */(s == HEADER) && (flg_type1 || flg_type2) && flg_read_tmp && (word_count_tmp != 27'd0) && flg_rcmem&&data_valid==1)

            word_count_rb <= word_count_tmp - 1;
        else if(rws_flg==0)
            begin
                if((re_rb || flg_rb_reg) && (word_count_rb != 27'd0))
                    word_count_rb <= word_count_rb - 1'b1;
            end 
    end

//cmem readback flag

    assign flg_rcmem   = (reg_cmd == 5'b00110);//read cmem, 
    always @(posedge CLK or negedge RST_N) begin
        if(RST_N == 1'b0)
            flg_rb_cmem <= 1'b0;
        else if(RW_SEL) begin
            if((flg_type1 || flg_type2) && flg_read_tmp && (word_count_rb != 27'd0) && flg_rcmem && (regaddr == 5'b0_0111))
                flg_rb_cmem <= 1'b1;
            //else if(word_count_rb == 27'd0)
                //flg_rb_cmem <= 1'b0;
            else if((re_rb || flg_rb_reg) && (word_count_rb == 27'd0))
                flg_rb_cmem <= 1'b0;
        end
        else begin
            flg_rb_cmem <= 1'b0;
        end
    end

    always @(posedge CLK or negedge RST_N) begin
        if(RST_N == 1'b0)
            flg_rb_cmem_d <= 1'b0;
        else 
            flg_rb_cmem_d <= flg_rb_cmem;
    end

    wire flg_rb_cmem_seu;
    assign flg_rb_cmem_seu = !flg_rb_cmem_d&flg_rb_cmem;

//command
    always@(*) begin
        if(!RST_N)
            reg_cmd = 0;
        else if(data_valid && flg_write && regaddr == 5'b00010)
            reg_cmd <= data[4:0];
    end

    assign flg_desync  = (reg_cmd == 5'b01011);//DESYNC


//////////////////////////////////////////////////reg array////////////////////////////////////////////////////////////////////

    always@(*) begin
        if(!RST_N) begin
            reg_crcr <= 0;
            reg_idr <= 0;
            reg_cmdr <= 0;
            reg_ctrl0r <= 0;
            reg_ctrl1r <= 0;
            reg_cmemir <= 0;
            reg_mfwriter <= 0;
            reg_ivr <= 0;
            reg_chainr <= 0;
            reg_adrr <= 0;
            reg_sbpir <= 0;
            reg_seur <= 0;
            reg_irstctrlr <= 0;
            reg_irstadrr <= 0;
            reg_watchdogr <= 0;
            reg_cmaskr <= 0;
            reg_keyr <= 0;
            reg_option0r <= 0;
            reg_option1r <= 0;
            reg_rcrr <= 0;
            reg_autr <= 0;
            reg_cmemor <= 32'hFFFF_FFFF;
            reg_seustatusr <= 0;
            reg_seuaddr <= 0;
            reg_seunaddr <= 0;
        end
        else begin
            if(data_valid && flg_write) begin
                case(regaddr)
                5'b00000 : reg_crcr <= data;          //
                5'b00001 : reg_idr <= IDCODE;         //
                5'b00010 : reg_cmdr <= data;          //
                5'b00011 : reg_ctrl0r <= data;        //
                5'b00100 : reg_ctrl1r <= data;        //
                5'b00101 : reg_cmemir <= data;        //
                5'b00110 : reg_mfwriter <= data;      //
                5'b01000 : reg_ivr <= data;           //
                5'b01010 : reg_chainr <= data;        //
                5'b01011 : begin                      //
                                reg_adrr <= data;     
                                reg_adrr_seu <= data;  
                           end
                5'b01100 : reg_sbpir <= data;         //
                5'b01101 : reg_seur <= data;          //
                5'b01111 : reg_irstctrlr <= data;     //
                5'b10000 : reg_irstadrr <= data;      //
                5'b10001 : reg_watchdogr <= data;     //
                5'b10111 : reg_cmaskr <= data;        //
                5'b11000 : reg_keyr <= data;          //
                5'b11001 : reg_option0r <= data;      //
                5'b11010 : reg_option1r <= data;      //
                5'b11011 : reg_rcrr <= data;          //
                5'b11110 : reg_autr <= data;          
                endcase
            end
            else if(!CS_N && flg_rb_reg) begin
                case(regaddr)
                5'b00000 : data_rb_reg <= reg_crcr;
                5'b00001 : data_rb_reg <= IDCODE;
                5'b00010 : data_rb_reg <= reg_cmdr;
                5'b00011 : data_rb_reg <= 32'h0000_0010;//reg_ctrl0r;
                5'b00100 : data_rb_reg <= reg_ctrl1r;
                5'b00111 : data_rb_reg <= reg_cmemor;
                5'b01001 : data_rb_reg <= reg_statusr;
                5'b01011 : data_rb_reg <= reg_adrr;
                5'b01100 : data_rb_reg <= reg_sbpir;
                5'b01101 : data_rb_reg <= reg_seur;
                5'b01110 : data_rb_reg <= reg_seustatusr;
                5'b01111 : data_rb_reg <= reg_irstctrlr;
                5'b10000 : data_rb_reg <= reg_irstadrr;
                5'b10001 : data_rb_reg <= 32'h3FFF_FFFF;//reg_watchdogr;
                5'b10010 : data_rb_reg <= reg_hstatusr;
                5'b10111 : data_rb_reg <= reg_cmaskr;
                5'b11001 : data_rb_reg <= reg_option0r;
                5'b11010 : data_rb_reg <= reg_option1r;
                5'b11011 : data_rb_reg <= 32'h0360_0000;//reg_rcrr;
                5'b11110 : data_rb_reg <= reg_autr;
                5'b11101 : data_rb_reg <= reg_seuaddr;
                5'b11111 : data_rb_reg <= reg_seunaddr;
                default  : data_rb_reg <= 32'hFFFF_FFFF;
                endcase                
            end
        end                    
    end

////////////////////////////////////////////////cmem_e1////////////////////////////////////////////////


    assign cmemclk = CLK && (data_valid || re_rb);
    assign we = (flg_write == 1 && regaddr == 5'b00101 && reg_cmd == 5'b00100) ? 1'b1 : 1'b0;
    assign cmemtype = reg_adrr[26:25];
    assign addr_region = reg_adrr[24:20];
    assign addr_column = reg_adrr[17:10];
    assign addr_frame = reg_adrr[7:0];
    assign region0 = (addr_region == 5'd0) ? 1 : 0;
    assign region1 = (addr_region == 5'd1) ? 1 : 0;
    assign region2 = (addr_region == 5'd2) ? 1 : 0;
    assign region3 = (addr_region == 5'd3) ? 1 : 0;


//    always@(posedge CLK or negedge RST_N) begin
//        if(!RST_N) begin
//            addr_word <= 0; 
//            flg_frame_end <= 0;
//            flg_column_end <= 0;
//            flg_region_end <= 0;
//         end
//        else if((we && data_valid) || (flg_rb_cmem && re_rb)) begin
//            addr_word <= addr_word + 1;
//            if(addr_word == 67) begin
//                addr_word <= 0;   
//                flg_frame_end <= 1;
//                reg_adrr[7:0] <= reg_adrr[7:0] + 1;//addr_frame + 1
//            end
//            else
//                flg_frame_end <= 0;
//        end
//    end


always@(posedge CLK or negedge RST_N)
begin
    if(RST_N==0)
        begin
            addr_word <= 0; 
            flg_frame_end <= 0;
            flg_column_end <= 0;
            flg_region_end <= 0;
        end
    else if(delay_flg==1)    // delay 10 CLK    
        addr_word <= addr_word;
    else if(we&&data_valid)  //write data to cmem
        begin
            addr_word <= addr_word + 1;
            if(addr_word == 67)  // number of a frame
                begin
                   addr_word <= 0;
                   flg_frame_end <= 1;
                   reg_adrr[7:0] <= reg_adrr[7:0] + 1;//addr_frame + 1
                end
            else 
                flg_frame_end <= 0;
        end
  //  else if(rws_flg==0)
      else if(rws_flg==0&&CS_N==0)
      begin
         if(flg_rb_cmem && re_rb) // read data from cmem
           begin
             addr_word <= addr_word + 1;
            if(addr_word == 67)
               begin
                  addr_word <= 0;
                  flg_frame_end <= 1;
                  reg_adrr[7:0] <= reg_adrr[7:0] + 1;//addr_frame + 1
               end
            else 
               flg_frame_end <= 0;               
        end
     end
end





    always@(posedge flg_rcmem) begin
        if(seu_en)
            flg_frame_end = 1;
    end


    always@(negedge CLK) begin//CLK
            if(we && data_valid) begin
                    cmem[addr_row][(67 - addr_word)*32] <= reg_cmemir[0];
                    cmem[addr_row][(67 - addr_word)*32 + 1] <= reg_cmemir[1];
                    cmem[addr_row][(67 - addr_word)*32 + 2] <= reg_cmemir[2];
                    cmem[addr_row][(67 - addr_word)*32 + 3] <= reg_cmemir[3];
                    cmem[addr_row][(67 - addr_word)*32 + 4] <= reg_cmemir[4];
                    cmem[addr_row][(67 - addr_word)*32 + 5] <= reg_cmemir[5];
                    cmem[addr_row][(67 - addr_word)*32 + 6] <= reg_cmemir[6];
                    cmem[addr_row][(67 - addr_word)*32 + 7] <= reg_cmemir[7];
                    cmem[addr_row][(67 - addr_word)*32 + 8] <= reg_cmemir[8];
                    cmem[addr_row][(67 - addr_word)*32 + 9] <= reg_cmemir[9];
                    cmem[addr_row][(67 - addr_word)*32 + 10] <= reg_cmemir[10];
                    cmem[addr_row][(67 - addr_word)*32 + 11] <= reg_cmemir[11];
                    cmem[addr_row][(67 - addr_word)*32 + 12] <= reg_cmemir[12];
                    cmem[addr_row][(67 - addr_word)*32 + 13] <= reg_cmemir[13];
                    cmem[addr_row][(67 - addr_word)*32 + 14] <= reg_cmemir[14];
                    cmem[addr_row][(67 - addr_word)*32 + 15] <= reg_cmemir[15];
                    cmem[addr_row][(67 - addr_word)*32 + 16] <= reg_cmemir[16];
                    cmem[addr_row][(67 - addr_word)*32 + 17] <= reg_cmemir[17];
                    cmem[addr_row][(67 - addr_word)*32 + 18] <= reg_cmemir[18];
                    cmem[addr_row][(67 - addr_word)*32 + 19] <= reg_cmemir[19];
                    cmem[addr_row][(67 - addr_word)*32 + 20] <= reg_cmemir[20];
                    cmem[addr_row][(67 - addr_word)*32 + 21] <= reg_cmemir[21];
                    cmem[addr_row][(67 - addr_word)*32 + 22] <= reg_cmemir[22];
                    cmem[addr_row][(67 - addr_word)*32 + 23] <= reg_cmemir[23];
                    cmem[addr_row][(67 - addr_word)*32 + 24] <= reg_cmemir[24];
                    cmem[addr_row][(67 - addr_word)*32 + 25] <= reg_cmemir[25];
                    cmem[addr_row][(67 - addr_word)*32 + 26] <= reg_cmemir[26];
                    cmem[addr_row][(67 - addr_word)*32 + 27] <= reg_cmemir[27];
                    cmem[addr_row][(67 - addr_word)*32 + 28] <= reg_cmemir[28];
                    cmem[addr_row][(67 - addr_word)*32 + 29] <= reg_cmemir[29];
                    cmem[addr_row][(67 - addr_word)*32 + 30] <= reg_cmemir[30];
                    cmem[addr_row][(67 - addr_word)*32 + 31] <= reg_cmemir[31];
                end
        end
        always@(*) begin
                if(flg_rb_cmem && !CS_N) begin
                    reg_cmemor[0] <= cmem[addr_row][(67 - addr_word)*32];
                    reg_cmemor[1] <= cmem[addr_row][(67 - addr_word)*32 + 1];
                    reg_cmemor[2] <= cmem[addr_row][(67 - addr_word)*32 + 2];
                    reg_cmemor[3] <= cmem[addr_row][(67 - addr_word)*32 + 3];
                    reg_cmemor[4] <= cmem[addr_row][(67 - addr_word)*32 + 4];
                    reg_cmemor[5] <= cmem[addr_row][(67 - addr_word)*32 + 5];
                    reg_cmemor[6] <= cmem[addr_row][(67 - addr_word)*32 + 6];
                    reg_cmemor[7] <= cmem[addr_row][(67 - addr_word)*32 + 7];
                    reg_cmemor[8] <= cmem[addr_row][(67 - addr_word)*32 + 8];
                    reg_cmemor[9] <= cmem[addr_row][(67 - addr_word)*32 + 9];
                    reg_cmemor[10] <= cmem[addr_row][(67 - addr_word)*32 + 10];
                    reg_cmemor[11] <= cmem[addr_row][(67 - addr_word)*32 + 11];
                    reg_cmemor[12] <= cmem[addr_row][(67 - addr_word)*32 + 12];
                    reg_cmemor[13] <= cmem[addr_row][(67 - addr_word)*32 + 13];
                    reg_cmemor[14] <= cmem[addr_row][(67 - addr_word)*32 + 14];
                    reg_cmemor[15] <= cmem[addr_row][(67 - addr_word)*32 + 15];
                    reg_cmemor[16] <= cmem[addr_row][(67 - addr_word)*32 + 16];
                    reg_cmemor[17] <= cmem[addr_row][(67 - addr_word)*32 + 17];
                    reg_cmemor[18] <= cmem[addr_row][(67 - addr_word)*32 + 18];
                    reg_cmemor[19] <= cmem[addr_row][(67 - addr_word)*32 + 19];
                    reg_cmemor[20] <= cmem[addr_row][(67 - addr_word)*32 + 20];
                    reg_cmemor[21] <= cmem[addr_row][(67 - addr_word)*32 + 21];
                    reg_cmemor[22] <= cmem[addr_row][(67 - addr_word)*32 + 22];
                    reg_cmemor[23] <= cmem[addr_row][(67 - addr_word)*32 + 23];
                    reg_cmemor[24] <= cmem[addr_row][(67 - addr_word)*32 + 24];
                    reg_cmemor[25] <= cmem[addr_row][(67 - addr_word)*32 + 25];
                    reg_cmemor[26] <= cmem[addr_row][(67 - addr_word)*32 + 26];
                    reg_cmemor[27] <= cmem[addr_row][(67 - addr_word)*32 + 27];
                    reg_cmemor[28] <= cmem[addr_row][(67 - addr_word)*32 + 28];
                    reg_cmemor[29] <= cmem[addr_row][(67 - addr_word)*32 + 29];
                    reg_cmemor[30] <= cmem[addr_row][(67 - addr_word)*32 + 30];
                    reg_cmemor[31] <= cmem[addr_row][(67 - addr_word)*32 + 31];
                end
    end



    //always@(posedge flg_rb_cmem) begin
    //    $readmemb("cmem.txt", cmem);  
    //end

    always@(negedge flg_rb_cmem) begin
        addr_word <= 0;
        reg_cmemor <= 32'hFFFF_FFFF;
    end


    always@(*)begin
        case(addr_region)
            0:  case (addr_column)
                    2, 3, 4, 5, 6, 7, 9, 10, 11, 12, 14, 15, 16, 17, 18, 19, 21, 22, 23, 24, 26, 27, 28, 29: begin //CLM
                        if(addr_frame < 28) begin
                            addr_row = 0 + 28* addr_column + addr_frame;
                            if(addr_frame == 27) begin
                                if(addr_column == 29)begin
                                   flg_column_end = 1;
                                   flg_region_end = 1; 
                                end                               
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 1;
                            end
                        end
                        else begin
                                flg_region_end = 0;
                                flg_column_end = 0;
                             end
                         end
                        else if(addr_frame == 28) begin 
                             if(addr_column == 29)begin
                                reg_adrr[7:0] = 0;
                                reg_adrr[17:10] =0;
                                reg_adrr[24:20] = 1;
                        end
                        else begin 
                                reg_adrr[7:0] = 0;
                                reg_adrr[17:10] = reg_adrr[17:10] + 1;
                         end
                       end
                    end
                    8, 13, 25: begin // DRM
                        if(addr_frame < 23) begin
                            addr_row = 0 + 28*addr_column + addr_frame;
                            if(addr_frame == 22) begin
                                flg_column_end = 1;
                                flg_region_end = 0;
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0;
                            end
                        end
                        else if(addr_frame == 23) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end    
                    20: begin //APM
                        if(addr_frame < 24) begin
                            addr_row = 0 + 28*addr_column + addr_frame;
                            if(addr_frame == 23) begin
                                flg_column_end = 1;
                                flg_region_end = 0;                
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0;
                            end
                        end
                        else if(addr_frame == 24) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;                        
                        end
                    end  
                    1: begin //IOL
                        if(addr_frame < 24) begin
                            addr_row = 0 + 28*addr_column + addr_frame;
                            if(addr_frame == 23) begin
                                flg_column_end = 1;
                                flg_region_end = 0;  
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0;
                            end
                        end
                        else if(addr_frame == 24) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end 
                    0: begin //IOB
                        if(addr_frame < 2) begin
                            addr_row = 0 + 28*addr_column + addr_frame;
                            if(addr_frame == 1) begin
                                flg_column_end = 1;
                                flg_region_end = 0;  
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0;
                            end
                        end
                        else if(addr_frame == 2) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;

                        end
                    end 
                   endcase
            1:  case(addr_column)
                 0, 1, 2, 3, 5, 6, 7, 8, 9, 10, 12, 13, 14, 15, 16, 17, 18, 19, 21, 22, 23, 24, 25, 26, 27:begin //CLM
                        if(addr_frame < 28) begin
                            addr_row = 28*30 + 28*addr_column + addr_frame;
                            if(addr_frame == 27) begin
                                flg_region_end = 0;
                                flg_column_end = 1;
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0;
                            end
                        end
                        else if(addr_frame == 28)begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end
                    4, 20: begin //DRM
                        if(addr_frame < 23) begin
                            addr_row = 28*30 + 28*addr_column + addr_frame;
                            if(addr_frame == 22) begin
                                flg_region_end = 0;
                                flg_column_end = 1;   
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0;     
                            end                       
                        end
                        else if(addr_frame == 23) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;                         
                        end
                    end
                    11 : begin //APM
                        if(addr_frame < 24) begin
                            addr_row = 28*30 + 28*addr_column + addr_frame;
                            if(addr_frame == 23) begin
                                flg_region_end = 0;
                                flg_column_end = 1;    
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0;  
                            end

                        end
                        else if(addr_frame == 24) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;                      
                        end
                    end
                    28: begin //IOL
                        if(addr_frame < 24) begin
                            addr_row = 28*30 + 28*addr_column + addr_frame;
                            if(addr_frame == 23) begin
                                flg_region_end = 0;
                                flg_column_end = 1;  
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0;  
                            end
                        end
                        else if(addr_frame == 24)begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1; 
                        end
                    end
                    29 : begin //IOB
                        if(addr_frame < 2) begin
                            addr_row = 28*30 + 28*addr_column + addr_frame;
                            if(addr_frame == 1) begin
                                    flg_region_end = 1;
                                    flg_column_end = 1;  
                                end
                                else begin
                                    flg_region_end = 0;
                                    flg_column_end = 0;  
                                end
                            end
                        else if(addr_frame == 2) begin
                                reg_adrr[7:0] = 0;
                                reg_adrr[17:10] = 0;
                                reg_adrr[24:20] = 2;
                            end
                         end              
                endcase
            2:  case(addr_column)
                    2, 3, 4, 5, 6, 7, 9, 10, 11, 12, 14, 15, 16, 17, 18, 19, 21, 22, 23, 24, 26, 27, 28, 29 :begin //CLM
                        if(addr_frame < 28) begin
                            addr_row = 28*(30 + 30) + 28*addr_column + addr_frame;
                            if(addr_frame == 27) begin
                               if(addr_column == 29)begin
                                flg_region_end = 1;
                                flg_column_end = 1;
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 1;
                            end
                        end
                        else begin 
                                flg_region_end = 0;
                                flg_column_end = 0;
                             end
                         end
                        else if(addr_frame == 28)begin
                           if(addr_column == 29)begin
                              reg_adrr[7:0] = 0;
                              reg_adrr[17:10] = 0;
                              reg_adrr[24:20] = 3;
                            end
                            else begin
                              reg_adrr[7:0] = 0;
                              reg_adrr[17:10] = reg_adrr[17:10] + 1;
                            end
                        end
                    end
                    8, 13, 25: begin //DRM
                        if(addr_frame < 23) begin
                            addr_row = 28*(30 + 30) + 28*addr_column + addr_frame;
                            if(addr_frame == 22) begin
                                flg_region_end = 0;
                                flg_column_end = 1; 
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0;    
                            end                        
                        end
                        else if(addr_frame == 23) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;                           
                        end
                    end
                    20: begin //APM
                            if(addr_frame < 24) begin
                            addr_row = 28*(30 + 30) + 28*addr_column + addr_frame;
                            if(addr_frame == 23) begin
                                flg_region_end = 0;
                                flg_column_end = 1;  
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0; 
                            end
                        end
                        else if(addr_frame == 24) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;                        
                        end
                    end
                    1: begin //IOL
                        if(addr_frame < 24) begin
                            addr_row = 28*(30 + 30) + 28*addr_column + addr_frame;
                            if(addr_frame == 23) begin
                                flg_region_end = 0;
                                flg_column_end = 1;   
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0;  
                            end
                        end
                        else if(addr_frame == 24)begin
                                reg_adrr[7:0] = 0;
                                reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end
                    0: begin //IOB
                        if(addr_frame < 2) begin
                            addr_row = 28*(30 + 30) + 28*addr_column + addr_frame;
                            if(addr_frame == 1) begin
                                 flg_region_end = 0;
                                 flg_column_end = 1;  
                                end
                             else begin
                                flg_region_end = 0;
                                flg_column_end = 0;  
                            end
                        end
                        else if(addr_frame == 2) begin
                                reg_adrr[7:0] = 0;
                                reg_adrr[17:10] = reg_adrr[17:10] + 1;
                            end
                    end                     
                endcase

            3:  case (addr_column)
                  0, 1, 2, 3, 5, 6, 7, 8, 9, 10, 12, 13, 14, 15, 16, 17, 18, 19, 21, 22, 23, 24, 25, 26, 27: begin //CLM
                        if(addr_frame < 28) begin
                            addr_row = 28*(30 + 30 + 30) + 28* addr_column + addr_frame;
                            if(addr_frame == 27) begin
                                flg_column_end = 1;
                                flg_region_end = 0;
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0;
                            end
                        end
                        else if(addr_frame == 28) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end
                    4, 20: begin // DRM
                        if(addr_frame < 23) begin
                            addr_row = 28*(30 + 30 + 30) + 28*addr_column + addr_frame;
                            if(addr_frame == 22) begin
                                flg_column_end = 1;
                                flg_region_end = 0;
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0;
                            end
                        end
                        else if(addr_frame == 23) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end    
                    11: begin //APM
                        if(addr_frame < 24) begin
                            addr_row = 28*(30 + 30 + 30) + 28*addr_column + addr_frame;
                            if(addr_frame == 23) begin
                                flg_column_end = 1;
                                flg_region_end = 0;  
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0;
                            end
                        end
                        else if(addr_frame == 24) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;                          
                        end
                    end  
                    28: begin //IOL
                        if(addr_frame < 24) begin
                            addr_row = 28*(30 + 30 + 30) + 30*addr_column + addr_frame;
                            if(addr_frame == 23) begin
                                flg_column_end = 1;
                                flg_region_end = 0;  
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0;
                            end
                        end
                        else if(addr_frame == 24) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end 
                    29: begin //IOB
                        if(addr_frame < 2) begin
                            addr_row = 28*(30 + 30 + 30) + 28*addr_column + addr_frame;
                            if(addr_frame == 1) begin
                                flg_column_end = 1;
                                flg_region_end = 1;  
                            end
                            else begin
                                flg_region_end = 0;
                                flg_column_end = 0;
                            end
                        end
                        else if(addr_frame == 2) begin
                                reg_adrr[7:0] = 0;
                                reg_adrr[17:10] = 0;
                                reg_adrr[24:20] = 0;
                             end
                          end
                    endcase
        endcase
    end    

///////////////////////////////////////////rb_crc///////////////////////////////////////////////////
    assign rbcrc_en = reg_seur[0];
    assign seu_en = (cmemtype == 2'b00) ? reg_seur[1] : 0;
    assign flg_rrbcrc = (rbcrc_en && (reg_cmd == 5'b01101)) ? 1 : 0;//reset readback CRC
    assign flg_rbcrc = (rbcrc_en && (reg_cmd == 5'b01110)) ? 1 : 0;//readback CRC

    ipal_e1_rbcrc CCS_RBCRC(

        .rstn               (RST_N),
        .clk                (CLK & (re_rb | data_valid)),
        .rbcrc_en           (rbcrc_en),
        .data               (reg_cmemor),
        .data_valid         (flg_rb_cmem),//
        .flg_rrbcrc         (flg_rrbcrc),
        .flg_rbcrc          (flg_rbcrc),
        .irstn              (RST_N),
        .iclk               (CLK & (re_rb | data_valid)),

        .rbcrc_err          (RBCRC_ERR),
        .rbcrc_valid        (RBCRC_VALID)
    );

///////////////////////////////////////seu///////////////////////////////////////////////////////////


    wire seu_we;
    wire ecc_valid_tmp;
    wire seu_clk;
    wire [31:0] seu_din;
    wire [6:0] seu_addr;
    reg  seu_we_d;
    reg  seu_we_d2;
    //reg  [6:0] addr_word_d;
    reg re_rb_d;
    reg re_rb_d2;
    reg re_rb_d3;
    reg re_rb_d4;
    wire clk_div;
    always@(posedge CLK or negedge RST_N) begin
        if(!RST_N) begin
            re_rb_d <= 0;
            re_rb_d2 <= 0;
            re_rb_d3 <= 0;
            re_rb_d4 <= 0;
        end
        else begin
            re_rb_d <= re_rb;
            re_rb_d2 <= re_rb_d;
            re_rb_d3 <= re_rb_d2;
            re_rb_d4 <= re_rb_d3;
        end
    end
    assign clk_div = (DATA_WIDTH == "X16") ? (re_rb | re_rb_d2) : (re_rb | re_rb_d4);
    assign seu_we = (DATA_WIDTH == "X32") ? flg_rb_cmem : re_rb;    
    assign seu_clk = (DATA_WIDTH == "X32") ? CLK : flg_rb_cmem ? clk_div : CLK;
    always@(negedge RST_N or posedge ECC_VALID or negedge CS_N) begin
        if(!RST_N) begin
            seu_we_d <= 0;
        end
        else if(ECC_VALID)
            seu_we_d <= 0;
        else begin
            if(!CS_N && RW_SEL && addr_word == 0 && seu_en)
                #0.1 seu_we_d <= 1;//seu_we;
            //else
                //seu_we_d <= 0;

            //addr_word_d <= addr_word;
        end
    end


    assign #0.1 seu_addr = addr_word;
    assign #0.1 seu_din = reg_cmemor;

    ipal_e1_secded CCS_SECDED (
        .rstn               (RST_N),
        .clk                (seu_clk),//seu_clk
        .en                 (seu_en),
        .addr               (seu_addr),//addr_word_d
        .we                 (seu_we_d),
        .din                (seu_din),//reg_cmemor

        .flg_ecc_over       (ecc_valid_tmp),
        .flg_sec            (serror),
        .flg_ded            (derror),
        .index              (ECC_INDEX)
    );
    reg ecc_valid_tmp_d;
    wire ecc_valid_tmp_p;
    always@(posedge CLK or negedge RST_N) begin
        if(!RST_N)
            ecc_valid_tmp_d <= 0;
        else
            ecc_valid_tmp_d <= ecc_valid_tmp;
    end
    assign ecc_valid_tmp_p = !ecc_valid_tmp_d&ecc_valid_tmp;
    assign ECC_VALID = ecc_valid_tmp_p&flg_rcmem; 

    always@(posedge CLK or negedge RST_N) begin
        if(!RST_N) begin
            serror_d <= 0;
            derror_d <= 0;
        end
        else begin
            serror_d <= serror;
            derror_d <= derror;
        end
    end

    assign SERROR = serror; //(!serror_d && serror) ? 1 : 0;
    assign DERROR = derror; //(!derror_d && derror) ? 1 : 0;



    
    reg serror_reg;
    reg derror_reg;
    reg [11:0]ecc_index_reg;
    reg ecc_valid_reg;

    always@(posedge ECC_VALID or negedge RST_N) begin
        if(!RST_N) begin
            serror_reg <= 0;
            derror_reg <= 0;
            ecc_index_reg <= 0;
            ecc_valid_reg <= 0;
        end
        else begin
            serror_reg <= SERROR;
            derror_reg <= DERROR;
            ecc_index_reg <= ECC_INDEX;
            ecc_valid_reg <= 1'b1;
        end
    end

    reg drcfg_over_reg;
    reg drcfg_err_reg;

    always@(posedge DRCFG_OVER or negedge RST_N) begin
        if(!RST_N) begin
            drcfg_over_reg <= 0;
            drcfg_err_reg <= 0;
        end
        else begin
            drcfg_over_reg <= DRCFG_OVER;
            drcfg_err_reg <= DRCFG_ERR;
        end
    end


    always@(*) begin
        if(RST_N) begin
            reg_seustatusr[31:17] = 0;
            reg_seustatusr[16] = drcfg_over_reg;
            reg_seustatusr[15] = drcfg_err_reg;
            reg_seustatusr[14:3] = ecc_index_reg;
            reg_seustatusr[2] = derror_reg;
            reg_seustatusr[1] = serror_reg;
            reg_seustatusr[0] = ecc_valid_reg;
        end
    end

/////////////////////////////////////////prcfg and drcfg/////////////////////////////////////////


    assign flg_prcfgen    = (reg_cmd == 5'b10100);
    assign flg_prcfgdis   = (reg_cmd == 5'b10101);
    assign flg_drcfgen    = (reg_cmd == 5'b10110);
    assign flg_drcfgdis   = (reg_cmd == 5'b10111);
    assign flg_rstcrc     = (reg_cmd == 5'b00001);
 
    assign PRCFG_OVER     = prcfg_over;
    assign PRCFG_ERR      = PRCFG_OVER ? prcfg_err : 0;
    assign DRCFG_OVER     = drcfg_over;
    assign DRCFG_ERR      = DRCFG_OVER ? drcfg_err : 0;

    always @(posedge CLK or negedge RST_N) begin
        if(RST_N == 1'b0)
            prcfg_en <= 1'b0;
        else if(flg_prcfgen)
            prcfg_en <= 1'b1;
        else if(flg_prcfgdis)
            prcfg_en <= 1'b0;
    end

    always@(posedge CLK or negedge RST_N) begin
        if(!RST_N)
            drcfg_en <= 0;
        else if(flg_drcfgen)
            drcfg_en <= 1;
        else if(flg_drcfgdis)
            drcfg_en <= 0;
    end

    always @(posedge CLK or negedge RST_N) begin
        if(RST_N == 1'b0)
            prcfg_en_d <= 1'b0;
        else
            prcfg_en_d <= prcfg_en;
    end

    always@(posedge CLK or negedge RST_N) begin
        if(!RST_N)
            drcfg_en_d <= 0;
        else
            drcfg_en_d <= drcfg_en;
    end

    always @(posedge CLK or negedge RST_N) begin
        if(RST_N == 1'b0)
            prcfg_over <= 1'b0;
        else if(!prcfg_en && prcfg_en_d)
            prcfg_over <= 1'b1;
        else
            prcfg_over <= 1'b0;
    end

    always@(posedge CLK or negedge RST_N) begin
        if(!RST_N)
            drcfg_over <= 0;
        else if(!drcfg_en && drcfg_en_d)
            drcfg_over <= 1;
        else 
            drcfg_over <= 0;
    end



 //   ipal_e1_crc  crc (

 //       .rstn                   (RST_N),
 //       .clk                    (CLK),
        
 //       .regaddr                (regaddr),
 //       .id_err                 (1'b0),
 //       .crc_disable            (reg_option1r[0]),//
 //       .data                   (data),
 //       .data_valid             (data_valid),
 //       .flg_write              (flg_write),
 //       .flg_rstcrc             (flg_rstcrc),//
//        .reg_crc                (reg_crcr),
//        .prcfg_en               (prcfg_en),
//        .prcfg_err              (prcfg_err),
//        .drcfg_en               (drcfg_en),
//        .drcfg_err              (drcfg_err),
//        .crc_err                (crc_err)//floating

//);
/////////////////////////////////////////FRAME\COLUMN\REGION/////////////////////////////////////////
    reg [7:0] addr_frame_seu;
    reg [7:0] addr_column_seu;
    reg [4:0] addr_region_seu;
    initial begin
        addr_frame_seu <= 0;
        addr_column_seu <= 0;
        addr_region_seu <= 0;
        reg_adrr_seu <= 0;
    end
    always@(reg_adrr) begin
        if(seu_en) begin
            addr_frame_seu <= reg_adrr_seu[7:0];
            addr_column_seu <= reg_adrr_seu[17:10];
            addr_region_seu <= reg_adrr_seu[24:20];
        end
    end

    //assign SEU_FRAME_ADDR = seu_en ? reg_adrr_seu[7:0] : 0;
    //assign SEU_COLUMN_ADDR = seu_en ? reg_adrr_seu[17:10] : 0;
    //assign SEU_REGION_ADDR = seu_en ? reg_adrr_seu[24:20] : 0;


    //assign SEU_FRAME_NADDR = seu_en ? (flg_column_end ? 0: SEU_FRAME_ADDR + flg_frame_end) : 0;
    //assign SEU_COLUMN_NADDR = seu_en ? (flg_region_end ? 0: SEU_COLUMN_ADDR + flg_column_end) : 0;
    //assign SEU_REGION_NADDR = seu_en ? (SEU_REGION_ADDR != 3 ? SEU_REGION_ADDR + flg_region_end : 0) : 0;


    initial begin
        SEU_REGION_ADDR = 0;
        SEU_COLUMN_ADDR = 0;
        SEU_FRAME_ADDR = 0;
        SEU_REGION_NADDR = 0;
        SEU_COLUMN_NADDR = 0;
        SEU_FRAME_NADDR = 0;   
    end

    always@(posedge CLK or negedge RST_N) begin
        if(!RST_N) begin
            SEU_REGION_ADDR = 0;
            SEU_COLUMN_ADDR = 0;
            SEU_FRAME_ADDR = 0;

            SEU_REGION_NADDR = 0;
            SEU_COLUMN_NADDR = 0;
            SEU_FRAME_NADDR = 0;
        end
        else if(flg_rb_cmem_seu && addr_word == 0)begin
            SEU_FRAME_ADDR = seu_en ? reg_adrr[7:0] : 0;
            SEU_COLUMN_ADDR = seu_en ? reg_adrr[17:10] : 0;
            SEU_REGION_ADDR = seu_en ? reg_adrr[24:20] : 0;

            SEU_FRAME_NADDR = seu_en ? (flg_column_end ? 0: SEU_FRAME_ADDR + flg_frame_end) : 0;
            SEU_COLUMN_NADDR = seu_en ? (flg_region_end ? 0: SEU_COLUMN_ADDR + flg_column_end) : 0;
            SEU_REGION_NADDR[1:0] = seu_en ? SEU_REGION_ADDR + flg_region_end : 0;  
        end
    end

    always@(*) begin
        reg_seuaddr <= {10'b0, SEU_REGION_ADDR, SEU_COLUMN_ADDR, SEU_FRAME_ADDR};
        reg_seunaddr <= {10'b0, SEU_REGION_NADDR, SEU_COLUMN_NADDR, SEU_FRAME_NADDR};
    end
//synthesis translate_on
endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: Internal simulation model
// Filename: INT_RAM144K.v
//
// Functional description: internal RAM block simulation model
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module INT_RAM144K
#(
    parameter GRS_EN = "TRUE",
    parameter integer DATA_WIDTH_A = 18,  /* 1 2 4 8 16 32 ; 9 18 36 */
    parameter integer DATA_WIDTH_B = 18,  /* 1 2 4 8 16 32 ; 9 18 36 */
    parameter CLEAR_TYPE   = "SYNC", /* ASYNC */
    parameter OUTPUT_REG_A = 0, /* ENABLE */
    parameter OUTPUT_REG_B = 0,
    parameter WRITE_MODE_A = "NORMAL_WRITE", /* TRANSPARENT_WRITE|READ_BEFORE_WRITE */
    parameter WRITE_MODE_B = "NORMAL_WRITE",
    parameter WRITE_COLLISION_ARBITER = "NULL", /* PORTA PORTB */
    parameter INIT_FILE = "NONE",
    parameter INIT_000 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_001 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_002 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_003 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_004 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_005 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_006 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_007 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_008 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_009 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_00A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_00B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_00C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_00D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_00E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_00F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_010 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_011 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_012 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_013 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_014 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_015 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_016 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_017 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_018 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_019 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_01A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_01B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_01C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_01D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_01E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_01F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_020 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_021 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_022 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_023 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_024 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_025 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_026 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_027 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_028 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_029 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_02A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_02B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_02C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_02D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_02E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_02F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_030 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_031 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_032 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_033 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_034 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_035 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_036 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_037 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_038 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_039 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_03A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_03B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_03C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_03D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_03E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_03F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_040 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_041 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_042 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_043 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_044 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_045 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_046 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_047 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_048 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_049 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_04A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_04B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_04C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_04D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_04E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_04F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_050 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_051 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_052 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_053 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_054 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_055 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_056 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_057 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_058 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_059 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_05A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_05B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_05C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_05D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_05E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_05F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_060 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_061 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_062 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_063 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_064 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_065 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_066 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_067 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_068 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_069 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_06A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_06B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_06C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_06D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_06E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_06F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_070 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_071 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_072 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_073 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_074 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_075 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_076 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_077 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_078 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_079 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_07A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_07B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_07C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_07D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_07E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_07F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_080 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_081 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_082 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_083 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_084 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_085 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_086 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_087 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_088 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_089 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_08A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_08B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_08C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_08D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_08E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_08F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_090 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_091 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_092 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_093 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_094 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_095 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_096 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_097 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_098 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_099 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_09A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_09B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_09C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_09D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_09E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_09F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0A0 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0A1 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0A2 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0A3 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0A4 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0A5 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0A6 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0A7 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0A8 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0A9 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0AA = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0AB = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0AC = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0AD = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0AE = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0AF = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0B0 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0B1 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0B2 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0B3 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0B4 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0B5 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0B6 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0B7 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0B8 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0B9 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0BA = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0BB = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0BC = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0BD = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0BE = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0BF = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0C0 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0C1 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0C2 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0C3 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0C4 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0C5 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0C6 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0C7 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0C8 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0C9 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0CA = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0CB = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0CC = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0CD = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0CE = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0CF = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0D0 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0D1 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0D2 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0D3 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0D4 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0D5 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0D6 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0D7 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0D8 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0D9 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0DA = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0DB = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0DC = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0DD = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0DE = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0DF = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0E0 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0E1 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0E2 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0E3 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0E4 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0E5 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0E6 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0E7 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0E8 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0E9 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0EA = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0EB = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0EC = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0ED = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0EE = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0EF = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0F0 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0F1 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0F2 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0F3 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0F4 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0F5 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0F6 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0F7 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0F8 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0F9 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0FA = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0FB = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0FC = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0FD = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0FE = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0FF = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_100 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_101 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_102 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_103 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_104 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_105 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_106 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_107 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_108 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_109 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_10A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_10B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_10C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_10D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_10E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_10F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_110 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_111 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_112 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_113 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_114 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_115 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_116 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_117 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_118 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_119 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_11A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_11B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_11C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_11D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_11E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_11F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_120 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_121 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_122 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_123 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_124 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_125 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_126 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_127 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_128 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_129 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_12A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_12B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_12C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_12D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_12E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_12F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_130 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_131 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_132 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_133 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_134 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_135 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_136 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_137 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_138 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_139 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_13A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_13B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_13C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_13D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_13E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_13F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_140 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_141 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_142 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_143 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_144 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_145 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_146 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_147 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_148 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_149 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_14A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_14B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_14C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_14D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_14E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_14F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_150 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_151 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_152 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_153 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_154 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_155 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_156 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_157 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_158 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_159 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_15A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_15B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_15C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_15D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_15E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_15F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_160 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_161 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_162 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_163 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_164 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_165 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_166 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_167 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_168 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_169 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_16A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_16B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_16C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_16D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_16E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_16F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_170 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_171 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_172 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_173 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_174 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_175 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_176 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_177 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_178 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_179 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_17A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_17B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_17C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_17D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_17E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_17F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_180 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_181 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_182 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_183 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_184 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_185 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_186 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_187 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_188 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_189 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_18A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_18B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_18C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_18D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_18E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_18F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_190 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_191 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_192 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_193 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_194 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_195 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_196 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_197 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_198 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_199 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_19A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_19B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_19C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_19D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_19E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_19F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1A0 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1A1 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1A2 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1A3 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1A4 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1A5 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1A6 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1A7 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1A8 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1A9 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1AA = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1AB = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1AC = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1AD = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1AE = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1AF = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1B0 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1B1 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1B2 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1B3 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1B4 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1B5 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1B6 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1B7 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1B8 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1B9 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1BA = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1BB = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1BC = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1BD = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1BE = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1BF = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1C0 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1C1 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1C2 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1C3 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1C4 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1C5 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1C6 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1C7 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1C8 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1C9 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1CA = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1CB = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1CC = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1CD = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1CE = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1CF = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1D0 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1D1 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1D2 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1D3 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1D4 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1D5 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1D6 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1D7 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1D8 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1D9 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1DA = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1DB = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1DC = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1DD = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1DE = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1DF = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1E0 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1E1 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1E2 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1E3 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1E4 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1E5 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1E6 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1E7 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1E8 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1E9 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1EA = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1EB = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1EC = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1ED = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1EE = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1EF = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1F0 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1F1 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1F2 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1F3 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1F4 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1F5 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1F6 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1F7 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1F8 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1F9 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1FA = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1FB = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1FC = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1FD = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1FE = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1FF = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter RAM_MODE = "TRUE_DUAL_PORT"
) (
    input wire CLKA, CEA,
    input wire WEA,
    input wire [3:0] BEA, /* byte write enable */
    input wire [16:0] ADDRA,
    input wire [35:0] DIA,
    input wire ORCEA, /* output reg clock enable*/
    input wire CLRA,  /* async/sync clear */
    output [35:0] DOA,
    //output reg [35:0] DOA,

    input wire CLKB, CEB,
    input wire WEB,
    input wire [3:0] BEB,
    input wire [16:0] ADDRB,
    input wire [35:0] DIB,
    input wire ORCEB, /* output reg clock enable*/
    input wire CLRB,  /* async/sync clear */
    output [35:0] DOB
    //output reg [35:0] DOB
);

    localparam MEM_WORDS = 16384;

    reg [8:0] mem [MEM_WORDS-1:0];

    integer cnt;
    reg [9*MEM_WORDS-1:0] init_value;

    reg [35:0] doa_buf = 'b0, doa_out = 'b0, doa_reg = 'b0;
    reg [35:0] dob_buf = 'b0, dob_out = 'b0, dob_reg = 'b0;

    assign grs =  (GRS_EN == "TRUE") ? ~GRS_INST.GRSNET : 1'b0;

    wire aclr_a = (CLEAR_TYPE == "ASYNC") ? (CLRA | grs): grs;
    wire sclr_a = (CLEAR_TYPE == "ASYNC") ? 1'b0 : CLRA;
    wire aclr_b = (CLEAR_TYPE == "ASYNC") ? (CLRB | grs): grs;
    wire sclr_b = (CLEAR_TYPE == "ASYNC") ? 1'b0 : CLRB;

    initial
    begin
        init_value = {
            INIT_1FF, INIT_1FE, INIT_1FD, INIT_1FC, INIT_1FB, INIT_1FA, INIT_1F9, INIT_1F8, INIT_1F7, INIT_1F6, INIT_1F5, INIT_1F4, INIT_1F3, INIT_1F2, INIT_1F1, INIT_1F0,
            INIT_1EF, INIT_1EE, INIT_1ED, INIT_1EC, INIT_1EB, INIT_1EA, INIT_1E9, INIT_1E8, INIT_1E7, INIT_1E6, INIT_1E5, INIT_1E4, INIT_1E3, INIT_1E2, INIT_1E1, INIT_1E0,
            INIT_1DF, INIT_1DE, INIT_1DD, INIT_1DC, INIT_1DB, INIT_1DA, INIT_1D9, INIT_1D8, INIT_1D7, INIT_1D6, INIT_1D5, INIT_1D4, INIT_1D3, INIT_1D2, INIT_1D1, INIT_1D0,
            INIT_1CF, INIT_1CE, INIT_1CD, INIT_1CC, INIT_1CB, INIT_1CA, INIT_1C9, INIT_1C8, INIT_1C7, INIT_1C6, INIT_1C5, INIT_1C4, INIT_1C3, INIT_1C2, INIT_1C1, INIT_1C0,
            INIT_1BF, INIT_1BE, INIT_1BD, INIT_1BC, INIT_1BB, INIT_1BA, INIT_1B9, INIT_1B8, INIT_1B7, INIT_1B6, INIT_1B5, INIT_1B4, INIT_1B3, INIT_1B2, INIT_1B1, INIT_1B0,
            INIT_1AF, INIT_1AE, INIT_1AD, INIT_1AC, INIT_1AB, INIT_1AA, INIT_1A9, INIT_1A8, INIT_1A7, INIT_1A6, INIT_1A5, INIT_1A4, INIT_1A3, INIT_1A2, INIT_1A1, INIT_1A0,
            INIT_19F, INIT_19E, INIT_19D, INIT_19C, INIT_19B, INIT_19A, INIT_199, INIT_198, INIT_197, INIT_196, INIT_195, INIT_194, INIT_193, INIT_192, INIT_191, INIT_190,
            INIT_18F, INIT_18E, INIT_18D, INIT_18C, INIT_18B, INIT_18A, INIT_189, INIT_188, INIT_187, INIT_186, INIT_185, INIT_184, INIT_183, INIT_182, INIT_181, INIT_180,
            INIT_17F, INIT_17E, INIT_17D, INIT_17C, INIT_17B, INIT_17A, INIT_179, INIT_178, INIT_177, INIT_176, INIT_175, INIT_174, INIT_173, INIT_172, INIT_171, INIT_170,
            INIT_16F, INIT_16E, INIT_16D, INIT_16C, INIT_16B, INIT_16A, INIT_169, INIT_168, INIT_167, INIT_166, INIT_165, INIT_164, INIT_163, INIT_162, INIT_161, INIT_160,
            INIT_15F, INIT_15E, INIT_15D, INIT_15C, INIT_15B, INIT_15A, INIT_159, INIT_158, INIT_157, INIT_156, INIT_155, INIT_154, INIT_153, INIT_152, INIT_151, INIT_150,
            INIT_14F, INIT_14E, INIT_14D, INIT_14C, INIT_14B, INIT_14A, INIT_149, INIT_148, INIT_147, INIT_146, INIT_145, INIT_144, INIT_143, INIT_142, INIT_141, INIT_140,
            INIT_13F, INIT_13E, INIT_13D, INIT_13C, INIT_13B, INIT_13A, INIT_139, INIT_138, INIT_137, INIT_136, INIT_135, INIT_134, INIT_133, INIT_132, INIT_131, INIT_130,
            INIT_12F, INIT_12E, INIT_12D, INIT_12C, INIT_12B, INIT_12A, INIT_129, INIT_128, INIT_127, INIT_126, INIT_125, INIT_124, INIT_123, INIT_122, INIT_121, INIT_120,
            INIT_11F, INIT_11E, INIT_11D, INIT_11C, INIT_11B, INIT_11A, INIT_119, INIT_118, INIT_117, INIT_116, INIT_115, INIT_114, INIT_113, INIT_112, INIT_111, INIT_110,
            INIT_10F, INIT_10E, INIT_10D, INIT_10C, INIT_10B, INIT_10A, INIT_109, INIT_108, INIT_107, INIT_106, INIT_105, INIT_104, INIT_103, INIT_102, INIT_101, INIT_100,
            INIT_0FF, INIT_0FE, INIT_0FD, INIT_0FC, INIT_0FB, INIT_0FA, INIT_0F9, INIT_0F8, INIT_0F7, INIT_0F6, INIT_0F5, INIT_0F4, INIT_0F3, INIT_0F2, INIT_0F1, INIT_0F0,
            INIT_0EF, INIT_0EE, INIT_0ED, INIT_0EC, INIT_0EB, INIT_0EA, INIT_0E9, INIT_0E8, INIT_0E7, INIT_0E6, INIT_0E5, INIT_0E4, INIT_0E3, INIT_0E2, INIT_0E1, INIT_0E0,
            INIT_0DF, INIT_0DE, INIT_0DD, INIT_0DC, INIT_0DB, INIT_0DA, INIT_0D9, INIT_0D8, INIT_0D7, INIT_0D6, INIT_0D5, INIT_0D4, INIT_0D3, INIT_0D2, INIT_0D1, INIT_0D0,
            INIT_0CF, INIT_0CE, INIT_0CD, INIT_0CC, INIT_0CB, INIT_0CA, INIT_0C9, INIT_0C8, INIT_0C7, INIT_0C6, INIT_0C5, INIT_0C4, INIT_0C3, INIT_0C2, INIT_0C1, INIT_0C0,
            INIT_0BF, INIT_0BE, INIT_0BD, INIT_0BC, INIT_0BB, INIT_0BA, INIT_0B9, INIT_0B8, INIT_0B7, INIT_0B6, INIT_0B5, INIT_0B4, INIT_0B3, INIT_0B2, INIT_0B1, INIT_0B0,
            INIT_0AF, INIT_0AE, INIT_0AD, INIT_0AC, INIT_0AB, INIT_0AA, INIT_0A9, INIT_0A8, INIT_0A7, INIT_0A6, INIT_0A5, INIT_0A4, INIT_0A3, INIT_0A2, INIT_0A1, INIT_0A0,
            INIT_09F, INIT_09E, INIT_09D, INIT_09C, INIT_09B, INIT_09A, INIT_099, INIT_098, INIT_097, INIT_096, INIT_095, INIT_094, INIT_093, INIT_092, INIT_091, INIT_090,
            INIT_08F, INIT_08E, INIT_08D, INIT_08C, INIT_08B, INIT_08A, INIT_089, INIT_088, INIT_087, INIT_086, INIT_085, INIT_084, INIT_083, INIT_082, INIT_081, INIT_080,
            INIT_07F, INIT_07E, INIT_07D, INIT_07C, INIT_07B, INIT_07A, INIT_079, INIT_078, INIT_077, INIT_076, INIT_075, INIT_074, INIT_073, INIT_072, INIT_071, INIT_070,
            INIT_06F, INIT_06E, INIT_06D, INIT_06C, INIT_06B, INIT_06A, INIT_069, INIT_068, INIT_067, INIT_066, INIT_065, INIT_064, INIT_063, INIT_062, INIT_061, INIT_060,
            INIT_05F, INIT_05E, INIT_05D, INIT_05C, INIT_05B, INIT_05A, INIT_059, INIT_058, INIT_057, INIT_056, INIT_055, INIT_054, INIT_053, INIT_052, INIT_051, INIT_050,
            INIT_04F, INIT_04E, INIT_04D, INIT_04C, INIT_04B, INIT_04A, INIT_049, INIT_048, INIT_047, INIT_046, INIT_045, INIT_044, INIT_043, INIT_042, INIT_041, INIT_040,
            INIT_03F, INIT_03E, INIT_03D, INIT_03C, INIT_03B, INIT_03A, INIT_039, INIT_038, INIT_037, INIT_036, INIT_035, INIT_034, INIT_033, INIT_032, INIT_031, INIT_030,
            INIT_02F, INIT_02E, INIT_02D, INIT_02C, INIT_02B, INIT_02A, INIT_029, INIT_028, INIT_027, INIT_026, INIT_025, INIT_024, INIT_023, INIT_022, INIT_021, INIT_020,
            INIT_01F, INIT_01E, INIT_01D, INIT_01C, INIT_01B, INIT_01A, INIT_019, INIT_018, INIT_017, INIT_016, INIT_015, INIT_014, INIT_013, INIT_012, INIT_011, INIT_010,
            INIT_00F, INIT_00E, INIT_00D, INIT_00C, INIT_00B, INIT_00A, INIT_009, INIT_008, INIT_007, INIT_006, INIT_005, INIT_004, INIT_003, INIT_002, INIT_001, INIT_000
            };
        if (INIT_FILE == "NONE")
        begin
            for (cnt = 0; cnt < MEM_WORDS; cnt = cnt + 1)
            begin
                mem[cnt] = init_value[cnt*9 +: 9];
            end
        end
        else
        begin
            $display("INIT_FILE do not support now.");
            $finish;
        end
    end

    //
    // input registers
    //=================
    //  ADDRA
    //  DIA
    //  WEA
    //  BEA
    //
    //  ADDRB
    //  DIB
    //  WEB
    //  BEB
    //

    //
    // task & function 
    //

    function [35:0] read_mem_a;
        input [16:0] addr;
    begin
        case (DATA_WIDTH_A)
            1: read_mem_a[0] = mem[addr[16:3]][addr[2:0]];
            2: read_mem_a[1:0] = mem[addr[16:3]][addr[2:1]*2 +: 2];
            4: read_mem_a[3:0] = mem[addr[16:3]][addr[2]*4 +: 4];
            8: read_mem_a[7:0] = mem[addr[16:3]][7:0];
            9: read_mem_a[8:0] = mem[addr[16:3]];
            16,
            18: read_mem_a[17:0] = {mem[addr[16:4]*2+1], mem[addr[16:4]*2]};
            32,
            36: read_mem_a = {mem[addr[16:5]*4+3], mem[addr[16:5]*4+2],
                              mem[addr[16:5]*4+1], mem[addr[16:5]*4]};
            default: /* null */ ;
        endcase
    end
    endfunction

    function [35:0] read_mem_b;
        input [16:0] addr;
    begin
        case (DATA_WIDTH_B)
            1: read_mem_b[0] = mem[addr[16:3]][addr[2:0]];
            2: read_mem_b[1:0] = mem[addr[16:3]][addr[2:1]*2 +: 2];
            4: read_mem_b[3:0] = mem[addr[16:3]][addr[2]*4 +: 4];
            8: read_mem_b[7:0] = mem[addr[16:3]][7:0];
            9: read_mem_b[8:0] = mem[addr[16:3]];
            16,
            18: read_mem_b[17:0] = {mem[addr[16:4]*2+1], mem[addr[16:4]*2]};
            32,
            36: read_mem_b = {mem[addr[16:5]*4+3], mem[addr[16:5]*4+2],
                              mem[addr[16:5]*4+1], mem[addr[16:5]*4]};
            default: /* null */ ;
        endcase
    end
    endfunction

    task write_mem_a;
        input [16:0] addr;
        input [35:0] data;
        input [3:0] byte_en;
    begin
        case (DATA_WIDTH_A)
            1: mem[addr[16:3]][addr[2:0]] = data[0];
            2: mem[addr[16:3]][addr[2:1]*2 +: 2] = data[1:0];
            4: mem[addr[16:3]][addr[2]*4 +: 4] = data[3:0];
            8: mem[addr[16:3]][7:0] = data[7:0];
            9: mem[addr[16:3]] = data[8:0];
            16: begin
                if (byte_en[1])
                    mem[addr[16:4]*2+1][7:0] = data[16:9];
                if (byte_en[0])
                    mem[addr[16:4]*2][7:0]   = data[7:0];
            end
            18: begin
                if (byte_en[1])
                    mem[addr[16:4]*2+1] = data[17:9];
                if (byte_en[0])
                    mem[addr[16:4]*2]   = data[8:0];
            end
            32: begin
                if (byte_en[3])
                    mem[addr[16:5]*4+3][7:0] = data[34:27];
                if (byte_en[2])
                    mem[addr[16:5]*4+2][7:0] = data[25:18];
                if (byte_en[1])
                    mem[addr[16:5]*4+1][7:0] = data[16:9];
                if (byte_en[0])
                    mem[addr[16:5]*4][7:0]   = data[7:0];
            end
            36: begin
                if (byte_en[3])
                    mem[addr[16:5]*4+3] = data[35:27];
                if (byte_en[2])
                    mem[addr[16:5]*4+2] = data[26:18];
                if (byte_en[1])
                    mem[addr[16:5]*4+1] = data[17:9];
                if (byte_en[0])
                    mem[addr[16:5]*4]   = data[8:0];
            end
            default: /* null */ ;
        endcase
    end
    endtask

    task write_mem_b;
        input [16:0] addr;
        input [35:0] data;
        input [3:0] byte_en;
    begin
        case (DATA_WIDTH_B)
            1: mem[addr[16:3]][addr[2:0]] = data[0];
            2: mem[addr[16:3]][addr[2:1]*2 +: 2] = data[1:0];
            4: mem[addr[16:3]][addr[2]*4 +: 4] = data[3:0];
            8: mem[addr[16:3]][7:0] = data[7:0];
            9: mem[addr[16:3]] = data[8:0];
            16: begin
                if (byte_en[1])
                    mem[addr[16:4]*2+1][7:0] = data[16:9];
                if (byte_en[0])
                    mem[addr[16:4]*2][7:0]   = data[7:0];
            end
            18: begin
                if (byte_en[1])
                    mem[addr[16:4]*2+1] = data[17:9];
                if (byte_en[0])
                    mem[addr[16:4]*2]   = data[8:0];
            end
            32: begin
                if (byte_en[3])
                    mem[addr[16:5]*4+3][7:0] = data[34:27];
                if (byte_en[2])
                    mem[addr[16:5]*4+2][7:0] = data[25:18];
                if (byte_en[1])
                    mem[addr[16:5]*4+1][7:0] = data[16:9];
                if (byte_en[0])
                    mem[addr[16:5]*4][7:0]   = data[7:0];
            end
            36: begin
                if (byte_en[3])
                    mem[addr[16:5]*4+3] = data[35:27];
                if (byte_en[2])
                    mem[addr[16:5]*4+2] = data[26:18];
                if (byte_en[1])
                    mem[addr[16:5]*4+1] = data[17:9];
                if (byte_en[0])
                    mem[addr[16:5]*4]   = data[8:0];
            end
            default: /* null */ ;
        endcase
    end
    endtask

    //
    // memory core
    //

    always @(posedge CLKA or posedge aclr_a)
    begin
        if (aclr_a == 1'b1 || sclr_a == 1'b1)
        begin
            doa_out <= 'b0;
        end

        if (CEA == 1'b1)
        begin
            if (aclr_a == 1'b1 || sclr_a == 1'b1)
            begin
                doa_buf = 'b0;
//                doa_out <= 'b0;
            end

            if (aclr_a == 1'b0 && sclr_a == 1'b0)
            begin
                if (WRITE_MODE_A == "READ_BEFORE_WRITE")
                    doa_buf = read_mem_a(ADDRA);
            end

            if (WEA == 1'b1)
            begin
                //if (CEB && WEB && (ADDRA == ADDRB) && (BEA == BEB) && sclr_a == 1'b0)
                ////if (CEB && WEB && (ADDRA == ADDRB) && sclr_a == 1'b0)
                //begin
                //    $display("RAM write collision at time %.3f ns (addr: %h)", $time/1000.0, ADDRA);
                //    if (WRITE_COLLISION_ARBITER == "PORTB")
                //        $display(" => WRITE_COLLISION_ARBITER is \"PORTB\", ignore port-A write");
                //    else
                //        write_mem_a(ADDRA, DIA, BEA);

                ////    if (WRITE_MODE_A == "READ_BEFORE_WRITE")
                ////        doa_buf = 'bx;
                //end
                //else
                    write_mem_a(ADDRA, DIA, BEA);
            end

            if (aclr_a == 1'b0 && sclr_a == 1'b0)
            begin /* read */
                if (WRITE_MODE_A != "READ_BEFORE_WRITE")
                    doa_buf = read_mem_a(ADDRA);

                // (Port A)read-write(Port B) collision
                //if (WEA == 1'b0 && CEB && WEB && ADDRA == ADDRB)
                //    if (WRITE_MODE_A == "READ_BEFORE_WRITE")
                //begin
                //    $display("RAM read(port-A) write(port-B) collision at time %.3f ns (addr: %h), force to 'X' output", $time/1000.0, ADDRA);
                //    doa_buf = 'bx;
                //end

                if (WEA == 1'b0 || WRITE_MODE_A != "NORMAL_WRITE")
                    doa_out <= doa_buf;
            end
        end
    end

    always @(posedge CLKB or posedge aclr_b)
    begin
        if (aclr_b == 1'b1 || sclr_b == 1'b1)
begin
        dob_out <= 'b0;
end
        if (CEB == 1'b1)
        begin
            if (aclr_b == 1'b1 || sclr_b == 1'b1)
            begin
                dob_buf = 'b0;
  //              dob_out <= 'b0;
            end

            if (aclr_b == 1'b0 && sclr_b == 1'b0)
            begin
                if (WRITE_MODE_B == "READ_BEFORE_WRITE")
                    dob_buf = read_mem_b(ADDRB);
            end

            if (WEB == 1'b1)
            begin
                //if (CEA && WEA && (ADDRA == ADDRB) && (BEA == BEB) && sclr_b == 1'b0)
                //begin
                //    $display("RAM write collision at time %.3f ns (addr: %h)", $time/1000.0, ADDRB);
                //    if (WRITE_COLLISION_ARBITER == "PORTA")
                //        $display(" => WRITE_COLLISION_ARBITER is \"PORTA\", ignore port-B write");
                //    else
                //        write_mem_b(ADDRB, DIB, BEB);

                //    //if (WRITE_MODE_B == "READ_BEFORE_WRITE")
                //    //    dob_buf = 'bx;
                //end
                //else
                    write_mem_b(ADDRB, DIB, BEB);
            end

            if (aclr_b == 1'b0 && sclr_b == 1'b0)
            begin /* read */
                if (WRITE_MODE_B != "READ_BEFORE_WRITE")
                    dob_buf = read_mem_b(ADDRB);

                // (Port B)read-write(Port A) collision
                //if (WEB == 1'b0 && CEA && WEA && ADDRA == ADDRB)
                //    if (WRITE_MODE_B == "READ_BEFORE_WRITE")
                //begin
                //    $display("RAM read(port-B) write(port-A) collision at time %.3f ns (addr: %h), force to 'X' output", $time/1000.0, ADDRB);
                //    dob_buf = 'bx;
                //end

                if (WEB == 1'b0 || WRITE_MODE_B != "NORMAL_WRITE")
                    dob_out <= dob_buf;
            end
        end
    end

    //
    // output register
    //

    always @(posedge CLKA or posedge aclr_a)
    begin
        if (OUTPUT_REG_A != 0)
        begin
            if (aclr_a == 1'b1 || sclr_a == 1'b1)
                doa_reg <= 'b0;
            else if (aclr_a == 1'b0 && sclr_a == 1'b0 && ORCEA == 1'b1)
                doa_reg <= doa_out;
        end
    end

    always @(posedge CLKB or posedge aclr_b)
    begin
        if (OUTPUT_REG_B != 0)
        begin
            if (aclr_b == 1'b1 || sclr_b == 1'b1)
                dob_reg <= 'b0;
            else if (aclr_b == 1'b0 && sclr_b == 1'b0 && ORCEB == 1'b1)
                dob_reg <= dob_out;
        end
    end

    assign DOA = ((OUTPUT_REG_A == 0) && (DATA_WIDTH_A == 1)) ? {19'b0,{8{doa_out[0]}},1'b0,{8{doa_out[0]}}} :
                 ((OUTPUT_REG_A == 0) && (DATA_WIDTH_A == 2)) ? {19'b0,{4{doa_out[1:0]}},1'b0,{4{doa_out[1:0]}}} :
                 ((OUTPUT_REG_A == 0) && (DATA_WIDTH_A == 4)) ? {19'b0,{2{doa_out[3:0]}},1'b0,{2{doa_out[3:0]}}} :
                 ((OUTPUT_REG_A == 0) && (DATA_WIDTH_A == 8)) ? {19'b0,doa_out[7:0],1'b0,doa_out[7:0]} :
                 ((OUTPUT_REG_A == 0) && (DATA_WIDTH_A == 9)) ? {18'b0,{2{doa_out[8:0]}}} :
                 ((OUTPUT_REG_A == 0) && (DATA_WIDTH_A == 16)) ? {19'b0,doa_out[16:9],1'b0,doa_out[7:0]} :
                 ((OUTPUT_REG_A == 0) && (DATA_WIDTH_A == 18)) ? {18'b0,doa_out[17:0]} :
                 ((OUTPUT_REG_A == 0) && ((DATA_WIDTH_A == 32) || (DATA_WIDTH_A == 36))) ? doa_out :
                 ((OUTPUT_REG_A == 1) && (DATA_WIDTH_A == 1)) ? {19'b0,{8{doa_reg[0]}},1'b0,{8{doa_reg[0]}}} :
                 ((OUTPUT_REG_A == 1) && (DATA_WIDTH_A == 2)) ? {19'b0,{4{doa_reg[1:0]}},1'b0,{4{doa_reg[1:0]}}} :
                 ((OUTPUT_REG_A == 1) && (DATA_WIDTH_A == 4)) ? {19'b0,{2{doa_reg[3:0]}},1'b0,{2{doa_reg[3:0]}}} :
                 ((OUTPUT_REG_A == 1) && (DATA_WIDTH_A == 8)) ? {19'b0,doa_reg[7:0],1'b0,doa_reg[7:0]} :
                 ((OUTPUT_REG_A == 1) && (DATA_WIDTH_A == 9)) ? {18'b0,{2{doa_reg[8:0]}}} :
                 ((OUTPUT_REG_A == 1) && (DATA_WIDTH_A == 16)) ? {19'b0,doa_reg[16:9],1'b0,doa_reg[7:0]} :
                 ((OUTPUT_REG_A == 1) && (DATA_WIDTH_A == 18)) ? {18'b0,doa_reg[17:0]} :
                 ((OUTPUT_REG_A == 1) && ((DATA_WIDTH_A == 32) || (DATA_WIDTH_A == 36))) ? doa_reg : 36'bx;

//    always @(*)
//    begin
//        if (OUTPUT_REG_A == 0)
//        begin
//            case (DATA_WIDTH_A)
//                1: DOA[35:0] = {19'b0,{8{doa_out[0]}},1'b0,{8{doa_out[0]}}};
//                2: DOA[35:0] = {19'b0,{4{doa_out[1:0]}},1'b0,{4{doa_out[1:0]}}};
//                4: DOA[35:0] = {19'b0,{2{doa_out[3:0]}},1'b0,{2{doa_out[3:0]}}};
//                8: DOA[35:0] = {19'b0,doa_out[7:0],1'b0,doa_out[7:0]};
//                9:  DOA[35:0]           = {18'b0,{2{doa_out[8:0]}}};
//                16:DOA[35:0] = {19'b0,doa_out[16:9],1'b0,doa_out[7:0]};
//                18: DOA[35:0] = {18'b0,doa_out[17:0]};
//                default: DOA = doa_out;
//            endcase
//        end
//        else
//        begin
//            case (DATA_WIDTH_A)
//                1: DOA[35:0] = {19'b0,{8{doa_reg[0]}},1'b0,{8{doa_reg[0]}}};
//                2: DOA[35:0] = {19'b0,{4{doa_reg[1:0]}},1'b0,{4{doa_reg[1:0]}}};
//                4: DOA[35:0] = {19'b0,{2{doa_reg[3:0]}},1'b0,{2{doa_reg[3:0]}}};
//                8: DOA[35:0] = {19'b0,doa_reg[7:0],1'b0,doa_reg[7:0]};
//                9:  DOA[35:0]           = {18'b0,{2{doa_reg[8:0]}}};
//                16:DOA[35:0] = {19'b0,doa_reg[16:9],1'b0,doa_reg[7:0]};
//                18: DOA[35:0] = {18'b0,doa_reg[17:0]};
//                default: DOA = doa_reg;
//            endcase
//        end
//    end

    assign DOB = ((OUTPUT_REG_B == 0) && (DATA_WIDTH_B == 1)) ? {19'b0,{8{dob_out[0]}},1'b0,{8{dob_out[0]}}} :
                 ((OUTPUT_REG_B == 0) && (DATA_WIDTH_B == 2)) ? {19'b0,{4{dob_out[1:0]}},1'b0,{4{dob_out[1:0]}}} :
                 ((OUTPUT_REG_B == 0) && (DATA_WIDTH_B == 4)) ? {19'b0,{2{dob_out[3:0]}},1'b0,{2{dob_out[3:0]}}} :
                 ((OUTPUT_REG_B == 0) && (DATA_WIDTH_B == 8)) ? {19'b0,dob_out[7:0],1'b0,dob_out[7:0]} :
                 ((OUTPUT_REG_B == 0) && (DATA_WIDTH_B == 9)) ? {18'b0,{2{dob_out[8:0]}}} :
                 ((OUTPUT_REG_B == 0) && (DATA_WIDTH_B == 16)) ? {19'b0,dob_out[16:9],1'b0,dob_out[7:0]} :
                 ((OUTPUT_REG_B == 0) && (DATA_WIDTH_B == 18)) ? {18'b0,dob_out[17:0]} :
                 ((OUTPUT_REG_B == 0) && ((DATA_WIDTH_B == 32) || (DATA_WIDTH_B == 36))) ? dob_out :
                 ((OUTPUT_REG_B == 1) && (DATA_WIDTH_B == 1)) ? {19'b0,{8{dob_reg[0]}},1'b0,{8{dob_reg[0]}}} :
                 ((OUTPUT_REG_B == 1) && (DATA_WIDTH_B == 2)) ? {19'b0,{4{dob_reg[1:0]}},1'b0,{4{dob_reg[1:0]}}} :
                 ((OUTPUT_REG_B == 1) && (DATA_WIDTH_B == 4)) ? {19'b0,{2{dob_reg[3:0]}},1'b0,{2{dob_reg[3:0]}}} :
                 ((OUTPUT_REG_B == 1) && (DATA_WIDTH_B == 8)) ? {19'b0,dob_reg[7:0],1'b0,dob_reg[7:0]} :
                 ((OUTPUT_REG_B == 1) && (DATA_WIDTH_B == 9)) ? {18'b0,{2{dob_reg[8:0]}}} :
                 ((OUTPUT_REG_B == 1) && (DATA_WIDTH_B == 16)) ? {19'b0,dob_reg[16:9],1'b0,dob_reg[7:0]} :
                 ((OUTPUT_REG_B == 1) && (DATA_WIDTH_B == 18)) ? {18'b0,dob_reg[17:0]} :
                 ((OUTPUT_REG_B == 1) && ((DATA_WIDTH_B == 32) || (DATA_WIDTH_B == 36))) ? dob_reg : 36'bx;
//    always @(*)
//    begin
//        if (OUTPUT_REG_B == 0)
//        begin
//            case (DATA_WIDTH_B)
//                1: DOB[35:0] = {19'b0,{8{dob_out[0]}},1'b0,{8{dob_out[0]}}};
//                2: DOB[35:0] = {19'b0,{4{dob_out[1:0]}},1'b0,{4{dob_out[1:0]}}};
//                4: DOB[35:0] = {19'b0,{2{dob_out[3:0]}},1'b0,{2{dob_out[3:0]}}};
//                8: DOB[35:0] = {19'b0,dob_out[7:0],1'b0,dob_out[7:0]};
//                9:  DOB[35:0]           = {18'b0,{2{dob_out[8:0]}}};
//                16:DOB[35:0] = {19'b0,dob_out[16:9],1'b0,dob_out[7:0]};
//                18: DOB[35:0] = {18'b0,dob_out[17:0]};
//                default: DOB = dob_out;
//            endcase
//        end
//        else
//        begin
//            case (DATA_WIDTH_B)
//                1: DOB[35:0] = {19'b0,{8{dob_reg[0]}},1'b0,{8{dob_reg[0]}}};
//                2: DOB[35:0] = {19'b0,{4{dob_reg[1:0]}},1'b0,{4{dob_reg[1:0]}}};
//                4: DOB[35:0] = {19'b0,{2{dob_reg[3:0]}},1'b0,{2{dob_reg[3:0]}}};
//                8: DOB[35:0] = {19'b0,dob_reg[7:0],1'b0,dob_reg[7:0]};
//                9:  DOB[35:0]           = {18'b0,{2{dob_reg[8:0]}}};
//                16:DOB[35:0] = {19'b0,dob_reg[16:9],1'b0,dob_reg[7:0]};
//                18: DOB[35:0] = {18'b0,dob_reg[17:0]};
//                default: DOB = dob_reg;
//            endcase
//        end
//    end

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_MULTADDSUM18.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

//P = (A0*B0 +/- A1*B1) +- (A2*B2 +/- A3*B3)
module GTP_MULTADDSUM18  #(
    parameter GRS_EN            = "TRUE", //"TRUE"; "FALSE"
    parameter SYNC_RST          = "FALSE", //"TRUE"; "FALSE"
    parameter INREG_EN          = "FALSE",  //"TRUE"; "FALSE"
    parameter PIPEREG_EN        = "FALSE",  //"TRUE"; "FALSE"
    parameter OUTREG_EN         = "FALSE",   //"TRUE"; "FALSE"
    parameter ADDSUB_OP         =2'b00 ,
    parameter SUM_ADDSUB_OP     = 0 ,
    parameter DYN_ADDSUB_OP     = 2'b11,
    parameter DYN_SUM_ADDSUB_OP = 1
)(
    output  [38-1:0] P,
    input   CE,
    input   RST,
    input   CLK,
    input   [1:0] A_SIGNED,
    input   [18-1:0] A0,
    input   [18-1:0] A1,
    input   [18-1:0] A2,
    input   [18-1:0] A3,
    input   [1:0] B_SIGNED,
    input   [18-1:0] B0,
    input   [18-1:0] B1,
    input   [18-1:0] B2,
    input   [18-1:0] B3,
    input   [1:0] ADDSUB,
    input   SUM_ADDSUB
);

    INT_MULTADDSUM #(
        . GRS_EN(GRS_EN),    
        . SYNC_RST(SYNC_RST),  
        . INREG_EN(INREG_EN),  
        . PIPEREG_EN(PIPEREG_EN),
        . OUTREG_EN(OUTREG_EN), 
        . ADDSUB_OP01(ADDSUB_OP[0]),  
        . ADDSUB_OP23(ADDSUB_OP[1]),  
        . ADDSUBSUM_OP(SUM_ADDSUB_OP), 
        . DYN_OP_SEL0(DYN_ADDSUB_OP[0]),
        . DYN_OP_SEL1(DYN_ADDSUB_OP[1]),
        . DYN_OP_SEL2(DYN_SUM_ADDSUB_OP),
        . ASIZE(18),
        . BSIZE(18)
    ) U_INT_MULTADDSUM (
        . CE(CE),
        . RST(RST),
        . CLK(CLK),
        . A_SIGNED01(A_SIGNED[0]),
        . A_SIGNED23(A_SIGNED[1]),
        . A0(A0),
        . A1(A1),
        . A2(A2),
        . A3(A3),
        . B_SIGNED01(B_SIGNED[0]),
        . B_SIGNED23(B_SIGNED[1]), 
        . B0(B0),
        . B1(B1),
        . B2(B2),
        . B3(B3),
        . ADDSUB01(ADDSUB[0]),
        . ADDSUB23(ADDSUB[1]),
        . ADDSUBSUM(SUM_ADDSUB),
        . P(P)
    );               

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////

//P = (A0*B0 +/- A1*B1) +- (A2*B2 +/- A3*B3)
`timescale 1 ns / 1 ps

module INT_MULTADDSUM  #(
parameter GRS_EN      = "FALSE", //"TRUE"; "FALSE"
parameter SYNC_RST    = "FALSE", //"TRUE"; "FALSE"
parameter SIB1_EN     = "FALSE", //"TRUE"; "FALSE"
parameter SIB2_EN     = "FALSE", //"TRUE"; "FALSE"
parameter SIB3_EN     = "FALSE", //"TRUE"; "FALSE"
parameter INREG_EN    = "FALSE",  //"TRUE"; "FALSE"
parameter PIPEREG_EN  = "FALSE",  //"TRUE"; "FALSE"
parameter OUTREG_EN   = "FALSE",   //"TRUE"; "FALSE"
parameter ADDSUB_OP01     = 1 ,
parameter ADDSUB_OP23     = 1 ,
parameter ADDSUBSUM_OP     = 1 ,
parameter SC_PSE_A0 = 0, //SC_PSE = 0, disable PSE, bit width = ASIZE-1
parameter SC_PSE_A1 = 0, //SC_PSE = 0, disable PSE, bit width = ASIZE-1  
parameter SC_PSE_A2 = 0, //SC_PSE = 0, disable PSE, bit width = ASIZE-1
parameter SC_PSE_A3 = 0, //SC_PSE = 0, disable PSE, bit width = ASIZE-1
parameter SC_PSE_B0 = 0, //SC_PSE = 0, disable PSE, bit width = BSIZE-1  
parameter SC_PSE_B1 = 0, //SC_PSE = 0, disable PSE, bit width = BSIZE-1
parameter SC_PSE_B2 = 0, //SC_PSE = 0, disable PSE, bit width = BSIZE-1
parameter SC_PSE_B3 = 0, //SC_PSE = 0, disable PSE, bit width = BSIZE-1
parameter DYN_OP_SEL0  = 1,
parameter DYN_OP_SEL1  = 1,
parameter DYN_OP_SEL2  = 1,
parameter ASIZE = 9,               //LEGAL ASIZE = 9, 18
parameter BSIZE = 9,               //LEGAL BSIZE = 9, 18
parameter PSIZE = ASIZE +BSIZE +1
)(
input   CE,
input   RST,
input   CLK,
input   A_SIGNED01,
input   A_SIGNED23,
input   [ASIZE-1:0] A0,
input   [ASIZE-1:0] A1,
input   [ASIZE-1:0] A2,
input   [ASIZE-1:0] A3,
input   B_SIGNED01,
input   B_SIGNED23,
input   [BSIZE-1:0] B0,
input   [BSIZE-1:0] B1,
input   [BSIZE-1:0] B2,
input   [BSIZE-1:0] B3,
input   ADDSUB01,
input   ADDSUB23,
input   ADDSUBSUM,
output  [PSIZE:0] P
);
parameter PRODUCT_SIZE = (ASIZE + BSIZE) *2;
parameter P_EXT  = ASIZE +3;
initial begin
    if ((ASIZE == 9 && BSIZE == 9) || (ASIZE == 18 && BSIZE == 18))
    begin 
    end
    else
        $display (" INT_MULTADDSUM error: illegal setting of ASIZE or BSIZE ");

    if (SIB1_EN != "FALSE" || SIB2_EN != "FALSE" || SIB3_EN != "FALSE") begin
        $display("DRC error");
        $finish;
    end
end      


reg  [ASIZE-1:0] P1_reg_A0;
reg  [ASIZE-1:0] P1_reg_A1;
reg  [ASIZE-1:0] P1_reg_A2;
reg  [ASIZE-1:0] P1_reg_A3;
reg  P1_reg_A_SIGNED01;
reg  P1_reg_A_SIGNED23;
reg  [BSIZE-1:0] P1_reg_B0;
reg  [BSIZE-1:0] P1_reg_B1;
reg  [BSIZE-1:0] P1_reg_B2;
reg  [BSIZE-1:0] P1_reg_B3;
reg  P1_reg_B_SIGNED01;
reg  P1_reg_B_SIGNED23;
reg  P1_reg_ADDSUB01;
reg  P1_reg_ADDSUB23;
reg  P1_reg_ADDSUBSUM;
wire [ASIZE-1:0] P1_reg_A0_comb;
wire [ASIZE-1:0] P1_reg_A1_comb;
wire [ASIZE-1:0] P1_reg_A2_comb;
wire [ASIZE-1:0] P1_reg_A3_comb;
wire P1_reg_A_SIGNED01_comb;
wire P1_reg_A_SIGNED23_comb;
wire [BSIZE-1:0] P1_reg_B0_comb;
wire [BSIZE-1:0] P1_reg_B1_comb;
wire [BSIZE-1:0] P1_reg_B2_comb;
wire [BSIZE-1:0] P1_reg_B3_comb;
wire P1_reg_B_SIGNED01_comb;
wire P1_reg_B_SIGNED23_comb;
reg  [PSIZE+1:0] P1_reg_A0_comb_ext;
reg  [PSIZE+1:0] P1_reg_A1_comb_ext;
reg  [PSIZE+1:0] P1_reg_A2_comb_ext;
reg  [PSIZE+1:0] P1_reg_A3_comb_ext;
reg  [PSIZE+1:0] P1_reg_B0_comb_ext;
reg  [PSIZE+1:0] P1_reg_B1_comb_ext;
reg  [PSIZE+1:0] P1_reg_B2_comb_ext;
reg  [PSIZE+1:0] P1_reg_B3_comb_ext;
wire [PRODUCT_SIZE-1:0] PRODUCT_0;
wire [PRODUCT_SIZE-1:0] PRODUCT_1;
wire [PRODUCT_SIZE-1:0] PRODUCT_2;
wire [PRODUCT_SIZE-1:0] PRODUCT_3;
wire  PRODUCT0_signed;
wire  PRODUCT1_signed;
wire  PRODUCT2_signed;
wire  PRODUCT3_signed;

reg  [PSIZE:0] P2_reg_PRODUCT_0;
reg  [PSIZE:0] P2_reg_PRODUCT_1;
reg  [PSIZE:0] P2_reg_PRODUCT_2;
reg  [PSIZE:0] P2_reg_PRODUCT_3;
reg  P2_reg_ADDSUB01;
wire P2_reg_ADDSUB01_comb;
reg  P2_reg_ADDSUB23;
wire P2_reg_ADDSUB23_comb;
reg  P2_reg_ADDSUBSUM;
wire P2_reg_ADDSUBSUM_comb;
wire [PSIZE:0] P2_reg_PRODUCT_0_comb;
wire [PSIZE:0] P2_reg_PRODUCT_1_comb;
wire [PSIZE:0] P2_reg_PRODUCT_2_comb;
wire [PSIZE:0] P2_reg_PRODUCT_3_comb;
wire [PSIZE:0] sum01;
wire [PSIZE:0] sum23;
wire [PSIZE:0] sum;
reg  [PSIZE:0] P_reg;
wire [ASIZE-1:0]  A1_comb;
wire [BSIZE-1:0]  B1_comb;
wire [ASIZE-1:0]  A2_comb;
wire [BSIZE-1:0]  B2_comb;
wire [ASIZE-1:0]  A3_comb;
wire [BSIZE-1:0]  B3_comb;
wire P1_reg_ADDSUB01_comb;
wire P1_reg_ADDSUB23_comb;
wire P1_reg_ADDSUBSUM_comb;
wire [ASIZE-1:0] A0_PSE;
wire [ASIZE-1:0] A1_PSE;
wire [ASIZE-1:0] A2_PSE;
wire [ASIZE-1:0] A3_PSE;
wire [BSIZE-1:0] B0_PSE;
wire [BSIZE-1:0] B1_PSE;
wire [BSIZE-1:0] B2_PSE;
wire [BSIZE-1:0] B3_PSE;

wire global_rstn, RST_sync, RST_async, rst_asyncomb;

assign global_rstn = GRS_EN == "TRUE" ? GRS_INST.GRSNET : 1'b1;
assign RST_sync = (SYNC_RST == "TRUE") ? RST : 1'b0;
assign RST_async = (SYNC_RST == "FALSE") ? RST : 1'b0;
assign rst_asyncomb = RST_async | (~global_rstn);

assign A1_comb = A1_PSE;
assign B1_comb = (SIB1_EN == "TRUE") ?  P1_reg_B0_comb :  B1_PSE;
assign A2_comb = A2_PSE;
assign B2_comb = (SIB2_EN == "TRUE") ?  P1_reg_B1_comb :  B2_PSE;
assign A3_comb = A3_PSE;
assign B3_comb = (SIB3_EN == "TRUE") ?  P1_reg_B2_comb :  B3_PSE;

INT_PSE #(.ASIZE(ASIZE),.SC_PSE(SC_PSE_A0)) U1_PSE(.A(A0), .SIGN(A_SIGNED01), .A_PSE(A0_PSE));
INT_PSE #(.ASIZE(ASIZE),.SC_PSE(SC_PSE_A1)) U2_PSE(.A(A1), .SIGN(A_SIGNED01), .A_PSE(A1_PSE));
INT_PSE #(.ASIZE(ASIZE),.SC_PSE(SC_PSE_A2)) U3_PSE(.A(A2), .SIGN(A_SIGNED23), .A_PSE(A2_PSE));
INT_PSE #(.ASIZE(ASIZE),.SC_PSE(SC_PSE_A3)) U4_PSE(.A(A3), .SIGN(A_SIGNED23), .A_PSE(A3_PSE));

INT_PSE #(.ASIZE(BSIZE),.SC_PSE(SC_PSE_B0)) U5_PSE(.A(B0), .SIGN(B_SIGNED01), .A_PSE(B0_PSE));
INT_PSE #(.ASIZE(BSIZE),.SC_PSE(SC_PSE_B1)) U6_PSE(.A(B1), .SIGN(B_SIGNED01), .A_PSE(B1_PSE));
INT_PSE #(.ASIZE(BSIZE),.SC_PSE(SC_PSE_B2)) U7_PSE(.A(B2), .SIGN(B_SIGNED23), .A_PSE(B2_PSE));
INT_PSE #(.ASIZE(BSIZE),.SC_PSE(SC_PSE_B3)) U8_PSE(.A(B3), .SIGN(B_SIGNED23), .A_PSE(B3_PSE));

initial begin
      P1_reg_A0        = 0;
      P1_reg_A1        = 0;
      P1_reg_A2        = 0;
      P1_reg_A3        = 0;      
      P1_reg_A_SIGNED01 = 0;
      P1_reg_A_SIGNED23 = 0;
      P1_reg_B0        = 0;
      P1_reg_B1        = 0;
      P1_reg_B2        = 0;
      P1_reg_B3        = 0;      
      P1_reg_B_SIGNED01 = 0;
      P1_reg_B_SIGNED23 = 0;
      P1_reg_ADDSUB01 = 0;
      P1_reg_ADDSUB23 = 0;
      P1_reg_ADDSUBSUM = 0;
      P2_reg_PRODUCT_0 = 0;
      P2_reg_PRODUCT_1 = 0;
      P2_reg_PRODUCT_2 = 0;
      P2_reg_PRODUCT_3 = 0;         
      P2_reg_ADDSUB01 = 0;
      P2_reg_ADDSUB23 = 0;
      P2_reg_ADDSUBSUM = 0;
      P_reg    = 0;
end

always @(posedge CLK or posedge rst_asyncomb)
   if (rst_asyncomb || RST_sync) begin
      P1_reg_A0        <= 0;
      P1_reg_A1        <= 0;
      P1_reg_A2        <= 0;
      P1_reg_A3        <= 0;      
      P1_reg_A_SIGNED01 <= 0;
      P1_reg_A_SIGNED23 <= 0;
      P1_reg_B0        <= 0;
      P1_reg_B1        <= 0;
      P1_reg_B2        <= 0;
      P1_reg_B3        <= 0;      
      P1_reg_B_SIGNED01 <= 0;
      P1_reg_B_SIGNED23 <= 0;
      P1_reg_ADDSUB01 <= 0;
      P1_reg_ADDSUB23 <= 0;
      P1_reg_ADDSUBSUM <= 0;
   end
      else if (CE) begin
         P1_reg_A0        <= A0_PSE;
         P1_reg_A1        <= A1_comb;
         P1_reg_A2        <= A2_comb;
         P1_reg_A3        <= A3_comb;
         P1_reg_A_SIGNED01 <= A_SIGNED01;
         P1_reg_A_SIGNED23 <= A_SIGNED23;
         P1_reg_B0        <= B0_PSE;
         P1_reg_B1        <= B1_comb;
         P1_reg_B2        <= B2_comb;         
         P1_reg_B3        <= B3_comb;         
         P1_reg_B_SIGNED01 <= B_SIGNED01;
         P1_reg_B_SIGNED23 <= B_SIGNED23;
         P1_reg_ADDSUB01 <= (DYN_OP_SEL0 == 1'b1)? ADDSUB01 : ADDSUB_OP01;
         P1_reg_ADDSUB23 <= (DYN_OP_SEL1 == 1'b1)? ADDSUB23 : ADDSUB_OP23;
         P1_reg_ADDSUBSUM <= (DYN_OP_SEL2 == 1'b1)? ADDSUBSUM:ADDSUBSUM_OP;
   end
   
assign P1_reg_A0_comb        = (INREG_EN == "TRUE") ? P1_reg_A0        : A0_PSE;
assign P1_reg_A1_comb        = (INREG_EN == "TRUE") ? P1_reg_A1        : A1_comb;
assign P1_reg_A2_comb        = (INREG_EN == "TRUE") ? P1_reg_A2        : A2_comb;
assign P1_reg_A3_comb        = (INREG_EN == "TRUE") ? P1_reg_A3        : A3_comb;
assign P1_reg_A_SIGNED01_comb = (INREG_EN == "TRUE") ? P1_reg_A_SIGNED01 : A_SIGNED01;
assign P1_reg_A_SIGNED23_comb = (INREG_EN == "TRUE") ? P1_reg_A_SIGNED23 : A_SIGNED23;
assign P1_reg_B0_comb        = (INREG_EN == "TRUE") ? P1_reg_B0        : B0_PSE;
assign P1_reg_B1_comb        = (INREG_EN == "TRUE") ? P1_reg_B1        : B1_comb;
assign P1_reg_B2_comb        = (INREG_EN == "TRUE") ? P1_reg_B2        : B2_comb;
assign P1_reg_B3_comb        = (INREG_EN == "TRUE") ? P1_reg_B3        : B3_comb;
assign P1_reg_B_SIGNED01_comb = (INREG_EN == "TRUE") ? P1_reg_B_SIGNED01 : B_SIGNED01;
assign P1_reg_B_SIGNED23_comb = (INREG_EN == "TRUE") ? P1_reg_B_SIGNED23 : B_SIGNED23;
assign P1_reg_ADDSUB01_comb = (INREG_EN == "TRUE") ? P1_reg_ADDSUB01 : (DYN_OP_SEL0 == 1'b1)? ADDSUB01 : ADDSUB_OP01;
assign P1_reg_ADDSUB23_comb = (INREG_EN == "TRUE") ? P1_reg_ADDSUB23 : (DYN_OP_SEL1 == 1'b1)? ADDSUB23 : ADDSUB_OP23;
assign P1_reg_ADDSUBSUM_comb = (INREG_EN == "TRUE") ? P1_reg_ADDSUBSUM :(DYN_OP_SEL2 == 1'b1)? ADDSUBSUM:ADDSUBSUM_OP ;


always @(*) begin
   if (P1_reg_A_SIGNED01_comb) begin
      P1_reg_A0_comb_ext = {{P_EXT{P1_reg_A0_comb[ASIZE-1]}}, P1_reg_A0_comb};
      P1_reg_A1_comb_ext = {{P_EXT{P1_reg_A1_comb[ASIZE-1]}}, P1_reg_A1_comb};
   end
   else begin
      P1_reg_A0_comb_ext = {{P_EXT{1'd0}}, P1_reg_A0_comb};
      P1_reg_A1_comb_ext = {{P_EXT{1'd0}}, P1_reg_A1_comb};
   end
end

always @(*) begin
   if (P1_reg_A_SIGNED23_comb) begin
      P1_reg_A2_comb_ext = {{P_EXT{P1_reg_A2_comb[ASIZE-1]}}, P1_reg_A2_comb};
      P1_reg_A3_comb_ext = {{P_EXT{P1_reg_A3_comb[ASIZE-1]}}, P1_reg_A3_comb};
   end
   else begin
      P1_reg_A2_comb_ext = {{P_EXT{1'd0}}, P1_reg_A2_comb};
      P1_reg_A3_comb_ext = {{P_EXT{1'd0}}, P1_reg_A3_comb};
   end
end

always @(*) begin
   if (P1_reg_B_SIGNED01_comb) begin
      P1_reg_B0_comb_ext = {{P_EXT{P1_reg_B0_comb[BSIZE-1]}}, P1_reg_B0_comb};
      P1_reg_B1_comb_ext = {{P_EXT{P1_reg_B1_comb[BSIZE-1]}}, P1_reg_B1_comb};
   end
   else begin
      P1_reg_B0_comb_ext = {{P_EXT{1'd0}}, P1_reg_B0_comb};
      P1_reg_B1_comb_ext = {{P_EXT{1'd0}}, P1_reg_B1_comb};
   end
end

always @(*) begin
   if (P1_reg_B_SIGNED23_comb) begin
      P1_reg_B2_comb_ext = {{P_EXT{P1_reg_B2_comb[BSIZE-1]}}, P1_reg_B2_comb};
      P1_reg_B3_comb_ext = {{P_EXT{P1_reg_B3_comb[BSIZE-1]}}, P1_reg_B3_comb};
   end
   else begin
      P1_reg_B2_comb_ext = {{P_EXT{1'd0}}, P1_reg_B2_comb};
      P1_reg_B3_comb_ext = {{P_EXT{1'd0}}, P1_reg_B3_comb};
   end
end

assign PRODUCT_0 = P1_reg_A0_comb_ext * P1_reg_B0_comb_ext;
assign PRODUCT_1 = P1_reg_A1_comb_ext * P1_reg_B1_comb_ext;
assign PRODUCT_2 = P1_reg_A2_comb_ext * P1_reg_B2_comb_ext;
assign PRODUCT_3 = P1_reg_A3_comb_ext * P1_reg_B3_comb_ext;
assign PRODUCT0_signed = P1_reg_A_SIGNED01_comb | P1_reg_B_SIGNED01_comb;
assign PRODUCT1_signed = P1_reg_A_SIGNED01_comb | P1_reg_B_SIGNED01_comb;
assign PRODUCT2_signed = P1_reg_A_SIGNED23_comb | P1_reg_B_SIGNED23_comb;
assign PRODUCT3_signed = P1_reg_A_SIGNED23_comb | P1_reg_B_SIGNED23_comb;

always @(posedge CLK or posedge rst_asyncomb)
   if (rst_asyncomb || RST_sync) begin
         P2_reg_PRODUCT_0 <= 0;
         P2_reg_PRODUCT_1 <= 0;
         P2_reg_PRODUCT_2 <= 0;
         P2_reg_PRODUCT_3 <= 0;         
         P2_reg_ADDSUB01 <= 0;
         P2_reg_ADDSUB23 <= 0;
         P2_reg_ADDSUBSUM <= 0;
   end
         else if (CE) begin
            P2_reg_PRODUCT_0 <= PRODUCT_0[PSIZE:0];
            P2_reg_PRODUCT_1 <= PRODUCT_1[PSIZE:0];
            P2_reg_PRODUCT_2 <= PRODUCT_2[PSIZE:0];
            P2_reg_PRODUCT_3 <= PRODUCT_3[PSIZE:0];
            P2_reg_ADDSUB01 <= P1_reg_ADDSUB01_comb;
            P2_reg_ADDSUB23 <= P1_reg_ADDSUB23_comb;
            P2_reg_ADDSUBSUM <= P1_reg_ADDSUBSUM_comb;
   end


assign P2_reg_PRODUCT_0_comb = (PIPEREG_EN == "TRUE") ? P2_reg_PRODUCT_0 : PRODUCT_0[PSIZE:0];
assign P2_reg_PRODUCT_1_comb = (PIPEREG_EN == "TRUE") ? P2_reg_PRODUCT_1 : PRODUCT_1[PSIZE:0];
assign P2_reg_PRODUCT_2_comb = (PIPEREG_EN == "TRUE") ? P2_reg_PRODUCT_2 : PRODUCT_2[PSIZE:0];
assign P2_reg_PRODUCT_3_comb = (PIPEREG_EN == "TRUE") ? P2_reg_PRODUCT_3 : PRODUCT_3[PSIZE:0];
assign P2_reg_ADDSUB01_comb = (PIPEREG_EN == "TRUE") ? P2_reg_ADDSUB01 : P1_reg_ADDSUB01_comb;
assign P2_reg_ADDSUB23_comb = (PIPEREG_EN == "TRUE") ? P2_reg_ADDSUB23 : P1_reg_ADDSUB23_comb;
assign P2_reg_ADDSUBSUM_comb = (PIPEREG_EN == "TRUE") ? P2_reg_ADDSUBSUM : P1_reg_ADDSUBSUM_comb;

assign sum01 = (P2_reg_ADDSUB01_comb == 0) ? (P2_reg_PRODUCT_0_comb + P2_reg_PRODUCT_1_comb) : 
                                       (P2_reg_PRODUCT_0_comb - P2_reg_PRODUCT_1_comb);
assign sum23 = (P2_reg_ADDSUB23_comb == 0) ? (P2_reg_PRODUCT_2_comb + P2_reg_PRODUCT_3_comb) : 
                                       (P2_reg_PRODUCT_2_comb - P2_reg_PRODUCT_3_comb);                                       
assign sum =   (P2_reg_ADDSUBSUM_comb == 0)? (sum01 + sum23) : (sum01 - sum23);

always @(posedge CLK or posedge rst_asyncomb)
   if (rst_asyncomb || RST_sync) begin
         P_reg    <= 0;
   end
         else if (CE) begin
         P_reg    <= sum;             
   end
   
assign P = (OUTREG_EN == "TRUE") ? P_reg : sum;

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2016 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_JTAGIF.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_JTAGIF
#(
    parameter USERCODE = 32'hFFFF_FFFF,
    parameter IDCODE = 32'h5555_AAAA
) (
    output      TDO,//user JTAG Test Data Out

    input       TCK,//50M user JTAG Test Clock
    input       TMS,//user JTAG Test Mode Select. determining the sequence of states through the tap controller on the rising edge of tck
    input       TDI//user JTAG Test Data In. the serial input to all JTAG instruction and data registers on the rising edge of tck
);
//synthesis translate_off

    localparam  TEST_LOGIC_RESET  =  4'd0;
    localparam  RUN_TEST_IDLE     =  4'd1;
    localparam  SELECT_IR_SCAN    =  4'd2;
    localparam  CAPTURE_IR        =  4'd3;
    localparam  SHIFT_IR          =  4'd4;
    localparam  EXIT1_IR          =  4'd5;
    localparam  PAUSE_IR          =  4'd6;
    localparam  EXIT2_IR          =  4'd7;
    localparam  UPDATE_IR         =  4'd8;
    localparam  SELECT_DR_SCAN    =  4'd9;
    localparam  CAPTURE_DR        =  4'd10;
    localparam  SHIFT_DR          =  4'd11;
    localparam  EXIT1_DR          =  4'd12;
    localparam  PAUSE_DR          =  4'd13;
    localparam  EXIT2_DR          =  4'd14;
    localparam  UPDATE_DR         =  4'd15;    




    reg [3:0] s;
    reg [3:0] ns;
    reg  jrst;
    reg  rti;
    reg [9:0] shift_ir;
    reg [9:0] update;
    reg capturedr;
    reg shiftdr;
    reg updatedr;
    reg exit1dr;
    reg exit2dr;
    reg shiftir;

    wire rst;
    wire flg_rti;
    wire flg_capture_ir;
    wire flg_shift_ir;
    wire flg_update_ir;
    wire flg_captre_dr;
    wire flg_shift_dr;
    wire flg_update_dr;
    wire flg_exit1_dr;
    wire flg_exit2_dr;
    wire tdo_ir;

//////////////////////////////////////////////////////tap control///////////////////////////////////////////////////////////////////////

    initial begin
        s <= 0;
        ns <= 0;
    end    

    always @(posedge TCK) begin
        s <= ns;
    end

    always @(*) begin
        case(s)

            TEST_LOGIC_RESET:
                begin
                    if(TMS)
                        ns = TEST_LOGIC_RESET;
                    else
                        ns = RUN_TEST_IDLE;
                end

            RUN_TEST_IDLE:
                begin
                    if(TMS)
                        ns = SELECT_DR_SCAN;
                    else
                        ns = RUN_TEST_IDLE;
                end

            SELECT_IR_SCAN:
                begin
                    if(TMS)
                        ns = TEST_LOGIC_RESET;
                    else
                        ns = CAPTURE_IR;
                end

            CAPTURE_IR, SHIFT_IR:
                begin
                    if(TMS)
                        ns = EXIT1_IR;
                    else
                        ns = SHIFT_IR;
                end
            
            EXIT1_IR:
                begin
                    if(TMS)
                        ns = UPDATE_IR;
                    else
                        ns = PAUSE_IR;
                end

            PAUSE_IR:
                begin
                    if(TMS)
                        ns = EXIT2_IR;
                    else
                        ns = PAUSE_IR;
                end

            EXIT2_IR:
                begin
                    if(TMS)
                        ns = UPDATE_IR;
                    else
                        ns = SHIFT_IR;
                end

            UPDATE_IR, UPDATE_DR:
                begin
                    if(TMS)
                        ns = SELECT_DR_SCAN;
                    else
                        ns = RUN_TEST_IDLE;
                end

            SELECT_DR_SCAN:
                begin
                    if(TMS)
                        ns = SELECT_IR_SCAN;
                    else
                        ns = CAPTURE_DR;
                end

            CAPTURE_DR, SHIFT_DR:
                begin
                    if(TMS)
                        ns = EXIT1_DR;
                    else
                        ns = SHIFT_DR;
                end

            EXIT1_DR:
                begin
                    if(TMS)
                        ns = UPDATE_DR;
                    else
                        ns = PAUSE_DR;
                end

            PAUSE_DR:
                begin
                    if(TMS)
                        ns = EXIT2_DR;
                    else
                        ns = PAUSE_DR;
                end

            EXIT2_DR:
                begin
                    if(TMS)
                        ns = UPDATE_DR;
                    else
                        ns = SHIFT_DR;
                end

        endcase
    end

    always @(negedge TCK) begin
        if(s == TEST_LOGIC_RESET)
            jrst <= 1'b1;
        else
            jrst <= 1'b0;
    end

    always @(negedge TCK) begin
        if(flg_rti)
            rti <= 1'b1;
        else
            rti <= 1'b0;
    end

    assign rst = (s == TEST_LOGIC_RESET);
    assign flg_rti = (s == RUN_TEST_IDLE);
    assign flg_capture_ir = (s == CAPTURE_IR);
    assign flg_shift_ir = (s == SHIFT_IR);
    assign flg_update_ir = (s == UPDATE_IR);
    assign flg_capture_dr = (s == CAPTURE_DR);
    assign flg_shift_dr = (s == SHIFT_DR);
    assign flg_update_dr = (s == UPDATE_DR);
    assign flg_exit1_dr = (s == EXIT1_DR);
    assign flg_exit2_dr = (s == EXIT2_DR);


//////////////////////////////////////////////////////////////////////IR///////////////////////////////////////////////////////
    localparam INS_IDCODE = 10'b10_1000_0011;

    always @(posedge TCK) begin
        if(rst)
            shift_ir <= 10'd0;
        else if(flg_capture_ir)
            shift_ir <= 10'b0;
        else if(flg_shift_ir)
            shift_ir <= {TDI, shift_ir[9:1]};
    end

    assign tdo_ir = shift_ir[0];

    always @(negedge TCK) begin
        if(rst)
            update <= INS_IDCODE;
        else if(flg_update_ir)
            update <= shift_ir;
    end


///////////////////////////////////////////////////////////////DR////////////////////////////////////////////////////////////
    always @(negedge TCK) begin
        if(rst)
            begin
                capturedr <= 1'b0;
                shiftdr <= 1'b0;
                updatedr <= 1'b0;
                exit1dr <= 1'b0;
                exit2dr <= 1'b0;
                shiftir <= 1'b0;
            end
        else
            begin
                capturedr <= flg_capture_dr;
                shiftdr <= flg_shift_dr;
                updatedr <= flg_update_dr;
                exit1dr <= flg_exit1_dr;
                exit2dr <= flg_exit2_dr;
                shiftir <= flg_shift_ir;
            end
    end

    reg tdo_tmp;
    always @(negedge TCK) begin
        if(rst)
            tdo_tmp <= 1'b0;
        else if(flg_shift_ir)
            tdo_tmp <= tdo_ir;
    end


    reg utdo;
    always @(*) begin
        if(shiftdr) begin
            //if(flg_read_flash)
                //utdo = tdo_flash;
            //else
                utdo = tdo_tmp;
        end
        else
            utdo = tdo_tmp;
    end

    assign TDO = (shiftir || shiftdr) ? utdo : 1'bz;


////////////////////////////////////////////////////////////////////////////////////////////////////

//bypass and highz and isc_enable and isc_disable and isc_noop and jrst and cfgi and jwakeup and jwakedown and program_flash and read_flash
    wire        tdo_bypass;
    wire        flg_bypass;
    wire        flg_highz;
    wire        flg_isc_enable;
    wire        flg_isc_disable;
    wire        flg_isc_noop;
    wire        flg_jrst;
    wire        flg_cfgi;
    wire        flg_jwakeup;
    wire        flg_jwakedown;
    wire        flg_program_flash;
    wire        flg_read_flash;

    reg         shift_bypass;

    localparam BYPASS = 10'b11_1111_1111;
    localparam HIGHZ = 10'b10_1000_0101;
    localparam ISC_ENABLE = 10'b01_0100_0000;
    localparam ISC_DISABLE = 10'b01_0100_0001;
    localparam ISC_NOOP = 10'b01_0100_0010;
    localparam JRST = 10'b10_1000_1010;
    localparam CFGI = 10'b10_1000_1011;
    localparam JWAKEUP = 10'b10_1000_1101;
    localparam JWAKEDOWN = 10'b10_1000_1110;
    localparam PROGRAM_FLASH = 10'b01_0100_1111;


    assign flg_bypass = (update == BYPASS);
    assign flg_highz = (update == HIGHZ);
    assign flg_isc_enable = (update == ISC_ENABLE);
    assign flg_isc_disable = (update == ISC_DISABLE);
    assign flg_isc_noop = (update == ISC_NOOP);
    assign flg_jrst = (update == JRST);
    assign flg_cfgi = (update == CFGI);
    assign flg_jwakeup = (update == JWAKEUP);
    assign flg_jwakedown = (update == JWAKEDOWN);
    assign flg_program_flash = (update == PROGRAM_FLASH);



    always@(posedge TCK) begin
        if(rst)
            shift_bypass <= 0;
        else if(capturedr)
            shift_bypass <= 0;
        else if((flg_bypass || flg_highz || flg_isc_enable || flg_isc_disable || flg_isc_noop ||flg_jrst || flg_cfgi || flg_jwakeup || flg_jwakedown || flg_program_flash) && shiftdr)
            shift_bypass <= TDI;
    end

    assign tdo_bypass = shift_bypass;

    always@(negedge TCK)begin
        if((flg_shift_dr) && (flg_bypass || flg_highz || flg_isc_enable || flg_isc_disable || flg_isc_noop ||flg_jrst || flg_cfgi || flg_jwakeup || flg_jwakedown || flg_program_flash))
        tdo_tmp <= tdo_bypass;
    end

//sample

    wire        tdo_sample;
    wire        flg_sample;
    
    reg [1:0]   shift_sample;

    localparam SAMPLE = 10'b10_1000_0000;

    assign flg_sample = (update == SAMPLE);

    always@(posedge TCK)begin
        if(rst)
            shift_sample <= 0;
        else if(flg_sample)begin
            if(capturedr) ;
            else if(shiftdr)
                shift_sample <= {TDI, shift_sample[1]};
            else if(updatedr) ;
        end
    end

    assign tdo_sample = shift_sample[0];

    always@(negedge TCK)begin
        if(flg_shift_dr && flg_sample)
            tdo_tmp <= tdo_sample;
    end

//idcode

    wire        tdo_idcode;
    wire        flg_idcode;

    reg [31:0]  shift_idcode;
    reg [31:0]  reg_idcode = 32'haaaa5555;

    assign flg_idcode = (update == INS_IDCODE);

    always@(posedge TCK) begin
        if(rst)
            shift_idcode <= 0;
        else if(flg_idcode)begin
            if(capturedr) 
                shift_idcode <= IDCODE;
            else if(shiftdr)
                shift_idcode <= {TDI, shift_idcode[31:1]};
        end
    end

    assign tdo_idcode = shift_idcode[0];

    always@(negedge TCK)begin
        if(flg_shift_dr && flg_idcode)
            tdo_tmp <= tdo_idcode;
    end

    
//usercode

    wire        tdo_usercode;
    wire        flg_usercode;

    reg [31:0]  shift_usercode;

    localparam USERCODEIR = 10'b10_1000_0100;

    assign flg_usercode = (update == USERCODEIR);
    
    always@(posedge TCK) begin
        if(rst)
            shift_usercode <= 0;
        else if(flg_usercode) begin
            if(capturedr) 
                shift_usercode <= USERCODE;
            else if(shiftdr)
                shift_usercode <= {TDI, shift_usercode[31:1]};
        end
    end

    assign tdo_usercode = shift_usercode[0];

    always@(negedge TCK)begin
        if(flg_shift_dr && flg_usercode)
            tdo_tmp <= tdo_usercode;
    end

//isc_program and isc_read

    wire        tdo_isc_program;
    wire        flg_isc_program;
    wire        flg_isc_read;

    reg [31:0]  shift_isc_program;

    localparam ISC_PROGRAM = 10'b01_0100_0011;
    localparam ISC_READ = 10'b01_0100_0100;

    assign flg_isc_program = (update == ISC_PROGRAM);
    assign flg_isc_read = (update == ISC_READ);

    always@(posedge TCK) begin
        if(rst)
            shift_isc_program <= 0;
        else if(flg_isc_program) begin
            if(shiftdr)
                shift_isc_program <= {shift_isc_program[30:0], TDI};
        end
        else if(flg_isc_read) begin
            if(shiftdr)
                shift_isc_program <= {shift_isc_program[30:0], TDI};
            else if(flg_rti) ;     
        end        
    end

    assign tdo_isc_program = shift_isc_program[31];

    always@(negedge TCK)begin
        if(flg_shift_dr &&(flg_isc_program || flg_isc_read))
            tdo_tmp <= tdo_isc_program;
    end

//userdr

//cfgo
    wire        flg_cfgo;
    wire        tdo_cfgo;

    reg [31:0]  shift_cfgo;
    reg [31:0]  shift_cfgo2;
    reg [31:0]  data_rb;
    reg         flg_rb_cmem;
    
    localparam CFGO = 10'b10_1000_1100;

    assign flg_cfgo = (update == CFGO);

    always@(posedge TCK)begin
        if(rst) begin
            shift_cfgo <= 0;
            shift_cfgo2 <= 0;
        end
        else if(flg_cfgo)begin
            if(capturedr) begin
                shift_cfgo  <= data_rb;
                shift_cfgo2 <= data_rb;
            end
            else if(shiftdr) begin
                if(flg_rb_cmem)
                    shift_cfgo2 <= {shift_cfgo2[30:0],TDI};
                else
                    shift_cfgo <= {shift_cfgo[30:0],TDI};
            end
        end
    end

    assign tdo_cfgo = flg_rb_cmem ? shift_cfgo2[31] : shift_cfgo[31];

    always@(negedge TCK)begin
        if(flg_shift_dr && flg_cfgo)
            tdo_tmp <= tdo_cfgo;
    end

//rdsr
    wire            tdo_rdsr;
    wire            flg_rdsr;

    reg     [31:0]  shift_rdsr;
    reg     [31:0]  reg_statusr;

    localparam RDSR = 10'b01_0101_1001;

    assign flg_rdsr = (update == RDSR);
    
    always@(posedge TCK) begin
        if(rst)
            shift_rdsr <= 0;
        else if(flg_rdsr) begin
            if(capturedr) 
                shift_rdsr <= reg_statusr;
            else if(shiftdr)
                shift_rdsr <= {TDI, shift_rdsr[31:1]};
        end        
    end

    assign tdo_rdsr = shift_rdsr[0];

    always@(negedge TCK)begin
        if(flg_shift_dr && flg_rdsr)
            tdo_tmp <= tdo_rdsr;
    end

//jdrp

    wire        tdo_jdrp;
    wire        flg_jdrp;
    reg [31:0]  shift_jdrp;
    reg [31:0]  update_jdrp;

    localparam JDRP = 10'b10_1000_1111;

    assign flg_jdrp = (update == JDRP);

    always@(posedge TCK) begin
        if(rst)
            shift_jdrp <= 0;
        else if(flg_jdrp) begin
            if(capturedr) 
                shift_jdrp <= 0;//{16'h0, ADC_register}
            else if(shiftdr)
                shift_jdrp <= {TDI, shift_jdrp[31:1]};
        end        
    end

    always@(negedge TCK) begin
        if(updatedr) 
            update_jdrp <= shift_jdrp;
    end

    assign tdo_jdrp = shift_jdrp[0];

    always@(negedge TCK)begin
        if(flg_shift_dr && flg_jdrp)
            tdo_tmp <= tdo_jdrp;
    end


//program_key and read_key
    wire        tdo_key;
    wire        flg_program_key;
    wire        flg_read_key;

    reg [255:0] shift_key;
    reg [255:0] capture_key;
    reg [255:0] update_key;
    reg         shift_keylock = 0;


    localparam PROGRAM_KEY = 10'b01_0100_0101;
    localparam READ_KEY = 10'b01_0100_0110;

    assign flg_program_key = (update == PROGRAM_KEY);
    assign flg_read_key = (update == READ_KEY);

    always@(posedge TCK) begin
        if(rst) begin
            shift_key <= 0;
            update_key <= 0;
        end
        else if(flg_program_key || flg_read_key)begin
            if(capturedr && !shift_keylock) 
                shift_key <= capture_key;
            else if(shiftdr)            
                shift_key <= {TDI, shift_key[255:1]};
        end
        else 
            shift_key <= shift_key;
    end

    always@(negedge TCK)begin
        if((flg_program_key || flg_read_key) && updatedr)
            update_key <= shift_key;
    end

    assign tdo_key = shift_key[0];

    always@(negedge TCK)begin
        if(flg_shift_dr && (flg_program_key || flg_read_key))
            tdo_tmp <= tdo_key;
    end

//program_keylock and read_keylock
    wire        tdo_keylock;
    wire        flg_program_keylock;
    wire        flg_read_keylock;

    //reg         shift_keylock = 0;
    reg         capture_keylock;
    reg         update_keylock;

    localparam PROGRAM_KEYLOCK = 10'b01_0100_0111;
    localparam READ_KEYLOCK = 10'b01_0100_1000;

    assign flg_program_keylock = (update == PROGRAM_KEYLOCK);
    assign flg_read_keylock = (update == READ_KEYLOCK);

    always@(posedge TCK) begin
        if(rst)
            shift_keylock <= 0;
        else if(flg_program_keylock) begin// || flg_read_keylock) && shiftdr)
            if(capturedr)
                shift_keylock <= capture_keylock;//from eFuse
            else if(shiftdr)
                shift_keylock <= TDI;
            else if(flg_rti)
                update_keylock <= shift_keylock;// to eFuse
        end
        else if(flg_read_keylock) begin
            if(capturedr)
                shift_keylock <= capture_keylock;//from eFuse
            else if(shiftdr)
                shift_keylock <= TDI;
        end
        else 
            shift_keylock <= shift_keylock;
    end

    assign tdo_keylock = shift_keylock;

    always@(negedge TCK) begin
        if(flg_shift_dr && (flg_program_keylock || flg_read_keylock))
            tdo_tmp <= tdo_keylock; 
    end

//program_fuse and read_fuse
    wire        tdo_fuse;
    wire        flg_program_fuse;
    wire        flg_read_fuse;

    reg [31:0]   shift_fuse;

    localparam PROGRAM_FUSE = 10'b01_0100_1001;
    localparam READ_FUSE = 10'b01_0100_1010;

    assign flg_program_fuse = (update == PROGRAM_FUSE);
    assign flg_read_fuse = (update == READ_FUSE);

    always@(posedge TCK) begin
        if(rst)
            shift_fuse <= 0;
        else if((flg_program_fuse || flg_read_fuse) && shiftdr)
            shift_fuse <= {TDI, shift_fuse[31:1]};
        else 
            shift_fuse <= shift_fuse;
    end

    assign tdo_fuse = shift_fuse[0];

    always@(negedge TCK)begin
        if(flg_shift_dr && (flg_program_fuse || flg_read_fuse))
            tdo_tmp <= tdo_fuse;
    end

//program_uid and read_uid
    wire        tdo_uid;
    wire        flg_program_uid;
    wire        flg_read_uid;

    reg [95:0]   shift_uid;

    localparam PROGRAM_UID = 10'b01_0100_1011;
    localparam READ_UID = 10'b01_0100_1100;

    assign flg_program_uid = (update == PROGRAM_UID);
    assign flg_read_uid = (update == READ_UID);

    always@(posedge TCK) begin
        if(rst)
            shift_uid <= 0;
        else if((flg_program_uid || flg_read_uid) && shiftdr)
            shift_uid <= {TDI, shift_uid[95:1]};
        else 
            shift_uid <= shift_uid;
    end

    assign tdo_uid = shift_uid[0];

    always@(negedge TCK) begin
        if(flg_shift_dr && (flg_program_uid || flg_read_uid))
            tdo_tmp <= tdo_uid;
    end

//program_tkey and read_tkey
    wire        tdo_tkey;
    wire        flg_program_tkey;
    wire        flg_read_tkey;

    reg [255:0]   shift_tkey;

    localparam PROGRAM_TKEY = 10'b01_0100_1101;
    localparam READ_TKEY = 10'b01_0100_1110;

    assign flg_program_tkey = (update == PROGRAM_TKEY);
    assign flg_read_tkey = (update == READ_TKEY);

    always@(posedge TCK) begin
        if(rst)
            shift_tkey <= 0;
        else if((flg_program_tkey || flg_read_tkey) && shiftdr)
            shift_tkey <= {TDI, shift_tkey[255:1]};
        else 
            shift_tkey <= shift_tkey;
    end

    assign tdo_tkey = shift_tkey[0];

    always@(negedge TCK)begin
        if(flg_shift_dr && (flg_program_tkey || flg_read_tkey))
            tdo_tmp <= tdo_tkey;
    end

//program_uidplock and read_uidplock
    wire        tdo_uidplock;
    wire        flg_program_uidplock;
    wire        flg_read_uidplock;

    reg         shift_uidplock;

    localparam PROGRAM_UIDPLOCK = 10'b01_0101_0101;
    localparam READ_UIDPLOCK = 10'b01_0101_0110;

    assign flg_program_uidplock = (update == PROGRAM_UIDPLOCK);
    assign flg_read_uidplock = (update == READ_UIDPLOCK);

    always@(posedge TCK) begin
        if(rst)
            shift_uidplock <= 0;
        else if((flg_program_uidplock || flg_read_uidplock) && shiftdr)
            shift_uidplock <= TDI;
        else 
            shift_uidplock <= shift_uidplock;
    end

    assign tdo_uidplock = shift_uidplock;

    always@(negedge TCK) begin
        if(flg_shift_dr && (flg_program_uidplock || flg_read_uidplock))
            tdo_tmp <= tdo_uidplock;
    end

//program_fuseplock and read_fuseplock
    wire        tdo_fuseplock;
    wire        flg_program_fuseplock;
    wire        flg_read_fuseplock;

    reg         shift_fuseplock;

    localparam PROGRAM_FUSEPLOCK = 10'b01_0101_0111;
    localparam READ_FUSEPLOCK = 10'b01_0101_1000;

    assign flg_program_fuseplock = (update == PROGRAM_FUSEPLOCK);
    assign flg_read_fuseplock = (update == READ_FUSEPLOCK);

    always@(posedge TCK) begin
        if(rst)
            shift_fuseplock <= 0;
        else if((flg_program_fuseplock || flg_read_fuseplock) && shiftdr)
            shift_fuseplock <= TDI;
        else 
            shift_fuseplock <= shift_fuseplock;
    end

    assign tdo_fuseplock = shift_fuseplock;

    always@(negedge TCK)begin
        if(flg_shift_dr && (flg_program_fuseplock || flg_read_fuseplock))
            tdo_tmp <= tdo_fuseplock;
    end

//program_ed and read_ed
    wire        tdo_ed;
    wire        flg_program_ed;
    wire        flg_read_ed;

    reg [383:0] shift_ed;

    localparam PROGRAM_ED = 10'b01_1000_0100;
    localparam READ_ED = 10'b01_1000_0101;

    assign flg_program_ed = (update == PROGRAM_ED);
    assign flg_read_ed = (update == READ_ED);

    always@(posedge TCK) begin
        if(rst)
            shift_ed <= 0;
        else if((flg_program_ed || flg_read_ed) && shiftdr)
            shift_ed <= {TDI, shift_ed[383:1]};
        else 
            shift_ed <= shift_ed;
    end

    assign tdo_ed = shift_ed[0];

    always@(negedge TCK)begin
        if(flg_shift_dr && (flg_program_ed || flg_read_ed))
            tdo_tmp <= tdo_ed;
    end

//program_ted and read_ted
    wire        tdo_ted;
    wire        flg_program_ted;
    wire        flg_read_ted;

    reg [383:0] shift_ted;

    localparam PROGRAM_TED = 10'b01_1000_0110;
    localparam READ_TED = 10'b01_1000_0111;
    
    assign flg_program_ted = (update == PROGRAM_TED);
    assign flg_read_ted = (update == READ_TED);

    always@(posedge TCK) begin
        if(rst)
            shift_ted <= 0;
        else if((flg_program_ted || flg_read_ted) && shiftdr)
            shift_ted <= {TDI, shift_ted[383:1]};
        else 
            shift_ted <= shift_ted;
    end

    assign tdo_ted = shift_ted[0];

    always@(negedge TCK)begin
        if(flg_shift_dr && (flg_program_ted || flg_read_ted))
            tdo_tmp <= tdo_ted;
    end

//program_edlock and read_edlock
    wire        tdo_edlock;
    wire        flg_program_edlock;
    wire        flg_read_edlock;

    reg         shift_edlock;

    localparam PROGRAM_EDLOCK = 10'b01_1000_1000;
    localparam READ_EDLOCK = 10'b01_1000_1001;

    assign flg_program_edlock = (update == PROGRAM_EDLOCK);
    assign flg_read_edlock = (update == READ_EDLOCK);

    always@(posedge TCK) begin
        if(rst)
            shift_edlock <= 0;
        else if((flg_program_edlock || flg_read_edlock) && shiftdr)
            shift_edlock <= TDI;
        else 
            shift_edlock <= shift_edlock;
    end

    assign tdo_edlock = shift_edlock;

    always@(negedge TCK) begin
        if(flg_shift_dr && (flg_program_edlock || flg_read_edlock))
            tdo_tmp <= tdo_edlock;
    end

//program_aut and read_aut
    wire        tdo_aut;
    wire        flg_program_aut;
    wire        flg_read_aut;

    reg         shift_aut;

    localparam PROGRAM_AUT = 10'b01_1000_1010;
    localparam READ_AUT = 10'b01_1000_1011;

    assign flg_program_aut = (update == PROGRAM_AUT);
    assign flg_read_aut = (update == READ_AUT);

    always@(posedge TCK) begin
        if(rst)
            shift_aut <= 0;
        else if((flg_program_aut || flg_read_aut) && shiftdr)
            shift_aut <= TDI;
        else 
            shift_aut <= shift_aut;
    end

    assign tdo_aut = shift_aut;

    always@(negedge TCK)begin
        if(flg_shift_dr && (flg_program_aut || flg_read_aut))
            tdo_tmp <= tdo_aut;
    end

//program_dpa and read_dpa
    wire        tdo_dpa;
    wire        flg_program_dpa;
    wire        flg_read_dpa;

    reg         shift_dpa;

    localparam PROGRAM_DPA = 10'b01_1000_1100;
    localparam READ_DPA = 10'b01_1000_1101;

    assign flg_program_dpa = (update == PROGRAM_DPA);
    assign flg_read_dpa = (update == READ_DPA);

    always@(posedge TCK) begin
        if(rst)
            shift_dpa <= 0;
        else if((flg_program_dpa || flg_read_dpa) && shiftdr)
            shift_dpa <= TDI;
        else 
            shift_dpa <= shift_dpa;
    end

    assign tdo_dpa = shift_dpa;

    always@(negedge TCK) begin
        if(flg_shift_dr && (flg_program_dpa || flg_read_dpa))
            tdo_tmp <= tdo_dpa;
    end

//program_tag and read_tag
    wire        tdo_tag;
    wire        flg_program_tag;
    wire        flg_read_tag;

    reg [127:0]   shift_tag;

    localparam PROGRAM_TAG = 10'b01_1000_1110;
    localparam READ_TAG = 10'b01_1000_1111;

    assign flg_program_tag = (update == PROGRAM_TAG);
    assign flg_read_tag = (update == READ_TAG);

    always@(posedge TCK) begin
        if(rst)
            shift_tag <= 0;
        else if((flg_program_tag || flg_read_tag) && shiftdr)
            shift_tag <= {TDI, shift_tag[127:1]};
        else 
            shift_tag <= shift_tag;
    end

    assign tdo_tag = shift_tag[0];

    always@(negedge TCK)begin
        if(flg_shift_dr && (flg_program_tag || flg_read_tag))
            tdo_tmp <= tdo_tag;
    end

//program_ttag and read_ttag
    wire        tdo_ttag;
    wire        flg_program_ttag;
    wire        flg_read_ttag;

    reg [127:0]   shift_ttag;

    localparam PROGRAM_TTAG = 10'b01_1001_0000;
    localparam READ_TTAG = 10'b01_1001_0001;

    assign flg_program_ttag = (update == PROGRAM_TTAG);
    assign flg_read_ttag = (update == READ_TTAG);

    always@(posedge TCK) begin
        if(rst)
            shift_ttag <= 0;
        else if((flg_program_ttag || flg_read_ttag) && shiftdr)
            shift_ttag <= {TDI, shift_ttag[127:1]};
        else 
            shift_ttag <= shift_ttag;
    end

    assign tdo_ttag = shift_ttag[0];
    
    always@(negedge TCK)begin
        if(flg_shift_dr && (flg_program_ttag || flg_read_ttag))
            tdo_tmp <= tdo_ttag;
    end

//program_obfus and read_obfus
    wire        tdo_obfus;
    wire        flg_program_obfus;
    wire        flg_read_obfus;

    reg         shift_obfus;

    localparam PROGRAM_OBFUS = 10'b01_1001_0010;
    localparam READ_OBFUS = 10'b01_1001_0011;

    assign flg_program_obfus = (update == PROGRAM_OBFUS);
    assign flg_read_obfus = (update == READ_OBFUS);
    
    always@(posedge TCK) begin
        if(rst)
            shift_obfus <= 0;
        else if((flg_program_obfus || flg_read_obfus) && shiftdr)
            shift_obfus <= TDI;
        else 
            shift_obfus <= shift_obfus;
    end

    assign tdo_obfus = shift_obfus;

    always@(negedge TCK)begin
        if(flg_shift_dr && (flg_program_obfus || flg_read_obfus))
            tdo_tmp <= tdo_obfus;
    end

//program_fuselock and read_fuselock
    wire        tdo_fuselock;
    wire        flg_program_fuselock;
    wire        flg_read_fuselock;

    reg         shift_fuselock;

    localparam PROGRAM_FUSELOCK = 10'b01_1001_0100;
    localparam READ_FUSELOCK = 10'b01_1001_0101;

    assign flg_program_fuselock = (update == PROGRAM_FUSELOCK);
    assign flg_read_fuselock = (update == READ_FUSELOCK);
    
    always@(posedge TCK) begin
        if(rst)
            shift_fuselock <= 0;
        else if((flg_program_fuselock || flg_read_fuselock) && shiftdr)
            shift_fuselock <= TDI;
        else 
            shift_fuselock <= shift_fuselock;
    end

    assign tdo_fuselock = shift_fuselock;

    always@(negedge TCK) begin
        if(flg_shift_dr && (flg_program_fuselock || flg_read_fuselock))
            tdo_tmp <= tdo_fuselock;
    end

//program_efuseclk and read_efuseclk
    wire        tdo_efuseclk;
    wire        flg_program_efuseclk;
    wire        flg_read_efuseclk;

    reg [9:0]   shift_efuseclk;
    reg [9:0]   update_efuseclk;

    localparam PROGRAM_EFUSECLK = 10'b01_1001_0110;
    localparam READ_EFUSECLK = 10'b01_1001_0111;

    assign flg_program_efuseclk = (update == PROGRAM_EFUSECLK);
    assign flg_read_efuseclk = (update == READ_EFUSECLK);

    always@(posedge TCK) begin
        if(rst) begin
            shift_efuseclk <= 0;
            update_efuseclk <= 0;
        end
        else if((flg_program_efuseclk || flg_read_efuseclk))begin
            if(capturedr)
                shift_efuseclk <= update_efuseclk;
            else if(shiftdr)   
                shift_efuseclk <= {TDI, shift_efuseclk[9:1]};
        end
        else 
            shift_efuseclk <= shift_efuseclk;
    end

    always@(negedge TCK)begin
        if((flg_program_efuseclk || flg_read_efuseclk) && updatedr)
            update_efuseclk <= shift_efuseclk;
    end

    assign tdo_efuseclk = shift_efuseclk[0];

    always@(negedge TCK) begin
        if(flg_shift_dr && (flg_program_efuseclk || flg_read_efuseclk))
            tdo_tmp <= tdo_efuseclk;
    end

//program_drmdpa and read_drmdpa
    wire        tdo_drmdpa;
    wire        flg_program_drmdpa;
    wire        flg_read_drmdpa;

    reg         shift_drmdpa;

    localparam PROGRAM_DRMDPA = 10'b01_1001_1000;
    localparam READ_DRMDPA = 10'b01_1001_1001;

    assign flg_program_drmdpa = (update == PROGRAM_DRMDPA);
    assign flg_read_drmdpa = (update == READ_DRMDPA);

    always@(posedge TCK) begin
        if(rst)
            shift_drmdpa <= 0;
        else if((flg_program_drmdpa || flg_read_drmdpa) && shiftdr)
            shift_drmdpa <= TDI;
        else 
            shift_drmdpa <= shift_drmdpa;
    end

    assign tdo_drmdpa = shift_drmdpa;

    always@(negedge TCK)begin
        if(flg_shift_dr && (flg_program_drmdpa || flg_read_drmdpa))
            tdo_tmp <= tdo_drmdpa;
    end

//program_taglock and read_taglock
    wire        tdo_taglock;
    wire        flg_program_taglock;
    wire        flg_read_taglock;

    reg         shift_taglock;

    localparam PROGRAM_TAGLOCK = 10'b01_1001_1010;
    localparam READ_TAGLOCK = 10'b01_1001_1011;
    
    assign flg_program_taglock = (update == PROGRAM_TAGLOCK);
    assign flg_read_taglock = (update == READ_TAGLOCK);

    always@(posedge TCK) begin
        if(rst)
            shift_taglock <= 0;
        else if((flg_program_taglock || flg_read_taglock) && shiftdr)
            shift_taglock <= TDI;
        else 
            shift_taglock <= shift_taglock;
    end

    assign tdo_taglock = shift_taglock;

    always@(negedge TCK)begin
        if(flg_shift_dr && (flg_program_taglock || flg_read_taglock))
            tdo_tmp <= tdo_taglock;
    end

//program_obfuslock and read_obfuslock
    wire        tdo_obfuslock;
    wire        flg_program_obfuslock;
    wire        flg_read_obfuslock;

    reg         shift_obfuslock;

    localparam PROGRAM_OBFUSLOCK = 10'b01_1001_1100;
    localparam READ_OBFUSLOCK = 10'b01_1001_1101;

    assign flg_program_obfuslock = (update == PROGRAM_OBFUSLOCK);
    assign flg_read_obfuslock = (update == READ_OBFUSLOCK);

    always@(posedge TCK) begin
        if(rst)
            shift_obfuslock <= 0;
        else if((flg_program_obfuslock || flg_read_obfuslock) && shiftdr)
            shift_obfuslock <= TDI;
        else 
            shift_obfuslock <= shift_obfuslock;
    end

    assign tdo_obfuslock = shift_obfuslock;

    always@(negedge TCK)begin
        if(flg_shift_dr && (flg_program_obfuslock || flg_read_obfuslock))
            tdo_tmp <= tdo_obfuslock;
    end

//program_autlock and read_autlock
    wire        tdo_autlock;
    wire        flg_program_autlock;
    wire        flg_read_autlock;

    reg         shift_autlock;

    localparam PROGRAM_AUTLOCK = 10'b01_1001_1110;
    localparam READ_AUTLOCK = 10'b01_1001_1111;

    assign flg_program_autlock = (update == PROGRAM_AUTLOCK);
    assign flg_read_autlock = (update == READ_AUTLOCK);

    always@(posedge TCK) begin
        if(rst)
            shift_autlock <= 0;
        else if((flg_program_autlock || flg_read_autlock) && shiftdr)
            shift_autlock <= TDI;
        else 
            shift_autlock <= shift_autlock;
    end

    assign tdo_autlock = shift_autlock;

    always@(negedge TCK) begin
        if(flg_shift_dr && (flg_program_autlock || flg_read_autlock))
            tdo_tmp <= tdo_autlock;
    end

//program_dpalock and read_dpalock
    wire        tdo_dpalock;
    wire        flg_program_dpalock;
    wire        flg_read_dpalock;

    reg         shift_dpalock;

    localparam PROGRAM_DPALOCK = 10'b01_1010_0000;
    localparam READ_DPALOCK = 10'b01_1010_0001;

    assign flg_program_dpalock = (update == PROGRAM_DPALOCK);
    assign flg_read_dpalock = (update == READ_DPALOCK);

    always@(posedge TCK) begin
        if(rst)
            shift_dpalock <= 0;
        else if((flg_program_dpalock || flg_read_dpalock) && shiftdr)
            shift_dpalock <= TDI;
        else 
            shift_dpalock <= shift_dpalock;
    end

    assign tdo_dpalock = shift_dpalock;

    always@(negedge TCK)begin
        if(flg_shift_dr && (flg_program_dpalock || flg_read_dpalock))
            tdo_tmp <= tdo_dpalock;
    end

//program_drmdpalock and read_drmdpalock
    wire        tdo_drmdpalock;
    wire        flg_program_drmdpalock;
    wire        flg_read_drmdpalock;

    reg         shift_drmdpalock;

    localparam PROGRAM_DRMDPALOCK = 10'b01_1010_0010;
    localparam READ_DRMDPALOCK = 10'b01_1010_0011;
    
    assign flg_program_drmdpalock = (update == PROGRAM_DRMDPALOCK);
    assign flg_read_drmdpalock = (update == READ_DRMDPALOCK);

    always@(posedge TCK) begin
        if(rst)
            shift_drmdpalock <= 0;
        else if((flg_program_drmdpalock || flg_read_drmdpalock) && shiftdr)
            shift_drmdpalock <= TDI;
        else 
            shift_drmdpalock <= shift_drmdpalock;
    end

    assign tdo_drmdpalock = shift_drmdpalock;

    always@(negedge TCK)begin
        if(flg_shift_dr && (flg_program_drmdpalock || flg_read_drmdpalock))
            tdo_tmp <= tdo_drmdpalock;
    end

//program_tdec and read_tdec
    wire        tdo_tdec;
    wire        flg_program_tdec;
    wire        flg_read_tdec;

    reg         shift_tdec;

    localparam PROGRAM_TDEC = 10'b01_1010_0100;
    localparam READ_TDEC = 10'b01_1010_0101;

    assign flg_program_tdec = (update == PROGRAM_TDEC);
    assign flg_read_tdec = (update == READ_TDEC);

    always@(posedge TCK) begin
        if(rst)
            shift_tdec <= 0;
        else if((flg_program_tdec || flg_read_tdec) && shiftdr)
            shift_tdec <= TDI;
        else 
            shift_tdec <= shift_tdec;
    end

    assign tdo_tdec = shift_tdec;

    always@(negedge TCK)begin
        if(flg_shift_dr && (flg_program_tdec || flg_read_tdec))
            tdo_tmp <= tdo_tdec;
    end

//program_tobfus and read_tobfus
    wire        tdo_tobfus;
    wire        flg_program_tobfus;
    wire        flg_read_tobfus;

    reg         shift_tobfus;

    localparam PROGRAM_TOBFUS = 10'b01_1010_0110;
    localparam READ_TOBFUS = 10'b01_1010_0111;

    assign flg_program_tobfus = (update == PROGRAM_TOBFUS);
    assign flg_read_tobfus = (update == READ_TOBFUS);

    always@(posedge TCK) begin
        if(rst)
            shift_tobfus <= 0;
        else if((flg_program_tobfus || flg_read_tobfus) && shiftdr)
            shift_tobfus <= TDI;
        else 
            shift_tobfus <= shift_tobfus;
    end

    assign tdo_tobfus = shift_tobfus;

    always@(negedge TCK)begin
        if(flg_shift_dr && (flg_program_tobfus || flg_read_tobfus))
            tdo_tmp <= tdo_tobfus;
    end

//program_taut and read_taut
    wire        tdo_taut;
    wire        flg_program_taut;
    wire        flg_read_taut;

    reg         shift_taut;

    localparam PROGRAM_TAUT = 10'b01_1010_1000;
    localparam READ_TAUT = 10'b01_1010_1001;

    assign flg_program_taut = (update == PROGRAM_TAUT);
    assign flg_read_taut = (update == READ_TAUT);

    always@(posedge TCK) begin
        if(rst)
            shift_taut <= 0;
        else if((flg_program_taut || flg_read_taut) && shiftdr)
            shift_taut <= TDI;
        else 
            shift_taut <= shift_taut;
    end

    assign tdo_taut = shift_taut;

    always@(negedge TCK)begin
        if(flg_shift_dr && (flg_program_taut || flg_read_taut))
            tdo_tmp <= tdo_taut;
    end

//program_tdpa and read_tdpa
    wire        tdo_tdpa;
    wire        flg_program_tdpa;
    wire        flg_read_tdpa;

    reg         shift_tdpa;

    localparam PROGRAM_TDPA = 10'b01_1010_1010;
    localparam READ_TDPA = 10'b01_1010_1011;

    assign flg_program_tdpa = (update == PROGRAM_TDPA);
    assign flg_read_tdpa = (update == READ_TDPA);

    always@(posedge TCK) begin
        if(rst)
            shift_tdpa <= 0;
        else if((flg_program_tdpa || flg_read_tdpa) && shiftdr)
            shift_tdpa <= TDI;
        else 
            shift_tdpa <= shift_tdpa;
    end

    assign tdo_tdpa = shift_tdpa;

    always@(negedge TCK)begin
        if(flg_shift_dr && (flg_program_tdpa || flg_read_tdpa))
            tdo_tmp <= tdo_tdpa;
    end

//program_tdrmdpa and read_tdrmdpa
    wire        tdo_tdrmdpa;
    wire        flg_program_tdrmdpa;
    wire        flg_read_tdrmdpa;

    reg         shift_tdrmdpa;

    localparam PROGRAM_TDRMDPA = 10'b01_1010_1100;
    localparam READ_TDRMDPA = 10'b01_1010_1101;

    assign flg_program_tdrmdpa = (update == PROGRAM_TDRMDPA);
    assign flg_read_tdrmdpa = (update == READ_TDRMDPA);

    always@(posedge TCK) begin
        if(rst)
            shift_tdrmdpa <= 0;
        else if((flg_program_tdrmdpa || flg_read_tdrmdpa) && shiftdr)
            shift_tdrmdpa <= TDI;
        else 
            shift_tdrmdpa <= shift_tdrmdpa;
    end

    assign tdo_tdrmdpa = shift_tdrmdpa;

    always@(negedge TCK)begin
        if(flg_shift_dr && (flg_program_tdrmdpa || flg_read_tdrmdpa))
            tdo_tmp <= tdo_tdrmdpa;
    end

//program_dec and read_dec
    wire        tdo_dec;
    wire        flg_program_dec;
    wire        flg_read_dec;

    reg         shift_dec;

    localparam PROGRAM_DEC = 10'b01_1010_1110;
    localparam READ_DEC = 10'b01_1010_1111;

    assign flg_program_dec = (update == PROGRAM_DEC);
    assign flg_read_dec = (update == READ_DEC);

    always@(posedge TCK) begin
        if(rst)
            shift_dec <= 0;
        else if((flg_program_dec || flg_read_dec) && shiftdr)
            shift_dec <= TDI;
        else 
            shift_dec <= shift_dec;
    end

    assign tdo_dec = shift_dec;

    always@(negedge TCK)begin
        if(flg_shift_dr && (flg_program_dec || flg_read_dec))
            tdo_tmp <= tdo_dec;
    end

//program_declock and read_declock
    wire        tdo_declock;
    wire        flg_program_declock;
    wire        flg_read_declock;

    reg         shift_declock;

    localparam PROGRAM_DECLOCK = 10'b01_1011_0000;
    localparam READ_DECLOCK = 10'b01_1011_0001;

    assign flg_program_declock = (update == PROGRAM_DECLOCK);
    assign flg_read_declock = (update == READ_DECLOCK);

    always@(posedge TCK) begin
        if(rst)
            shift_declock <= 0;
        else if((flg_program_declock || flg_read_declock) && shiftdr)
            shift_declock <= TDI;
        else 
            shift_declock <= shift_declock;
    end

    assign tdo_declock = shift_declock;

    always@(negedge TCK)begin
        if(flg_shift_dr && (flg_program_declock || flg_read_declock))
            tdo_tmp <= tdo_declock;
    end

//program_bbkey and read_bbkey
    wire        tdo_bbkey;
    wire        flg_program_bbkey;
    wire        flg_read_bbkey;

    reg [255:0] shift_bbkey;

    localparam PROGRAM_BBKEY = 10'b01_1011_0010;
    localparam READ_BBKEY = 10'b01_1011_0011;

    assign flg_program_bbkey = (update == PROGRAM_BBKEY);
    assign flg_read_bbkey = (update == READ_BBKEY);

    always@(posedge TCK) begin
        if(rst) 
            shift_bbkey <= 0;
        else if((flg_program_bbkey || flg_read_bbkey) && shiftdr)
            shift_bbkey <= {TDI, shift_bbkey[255:1]};
        else 
            shift_bbkey <= shift_bbkey;
    end

    assign tdo_bbkey = shift_bbkey[0];

    always@(negedge TCK)begin
        if(flg_shift_dr && (flg_program_bbkey || flg_read_bbkey))
            tdo_tmp <= tdo_bbkey;
    end

//peogram_bbkeylock and read_bbkeylock
    wire        tdo_bbkeylock;
    wire        flg_program_bbkeylock;
    wire        flg_read_bbkeylock;

    reg         shift_bbkeylock;

    localparam PROGRAM_BBKEYLOCK = 10'b01_1011_0100;
    localparam READ_BBKEYLOCK = 10'b01_1011_0101;
    
    assign flg_program_bbkeylock = (update == PROGRAM_BBKEYLOCK);
    assign flg_read_bbkeylock = (update == READ_BBKEYLOCK);

    always@(posedge TCK) begin
        if(rst)
            shift_bbkeylock <= 0;
        else if((flg_program_bbkeylock || flg_read_bbkeylock) && shiftdr)
            shift_bbkeylock <= TDI;
        else 
            shift_bbkeylock <= shift_bbkeylock;
    end

    assign tdo_bbkeylock = shift_bbkeylock;

    always@(negedge TCK)begin
        if(flg_shift_dr && (flg_program_bbkeylock || flg_read_bbkeylock))
            tdo_tmp <= tdo_bbkeylock;
    end

//program_keyen and read_keyen
    wire        tdo_keyen;
    wire        flg_program_keyen;
    wire        flg_read_keyen;

    reg         shift_keyen;

    localparam PROGRAM_KEYEN = 10'b01_1011_0110;
    localparam READ_KEYEN = 10'b01_1011_0111;

    assign flg_program_keyen = (update == PROGRAM_KEYEN);
    assign flg_read_keyen = (update == READ_KEYEN);

    always@(posedge TCK) begin
        if(rst)
            shift_keyen <= 0;
        else if((flg_program_keyen || flg_read_keyen) && shiftdr)
            shift_keyen <= TDI;
        else 
            shift_keyen <= shift_keyen;
    end

    assign tdo_keyen = shift_keyen;

    always@(negedge TCK)begin
        if(flg_shift_dr && (flg_program_keyen || flg_read_keyen))
            tdo_tmp <= tdo_keyen;
    end

//program_keyenlock and read_keyenlock
    wire        tdo_keyenlock;
    wire        flg_program_keyenlock;
    wire        flg_read_keyenlock;

    reg         shift_keyenlock;

    localparam PROGRAM_KEYENLOCK = 10'b01_1011_1000;
    localparam READ_KEYENLOCK = 10'b01_1011_1001;

    assign flg_program_keyenlock = (update == PROGRAM_KEYENLOCK);
    assign flg_read_keyenlock = (update == READ_KEYENLOCK);

    always@(posedge TCK) begin
        if(rst)
            shift_keyenlock <= 0;
        else if((flg_program_keyenlock || flg_read_keyenlock) && shiftdr)
            shift_keyenlock <= TDI;
        else 
            shift_keyenlock <= shift_keyenlock;
    end

    assign tdo_keyenlock = shift_keyenlock;

    always@(negedge TCK)begin
        if(flg_shift_dr && (flg_program_keyenlock || flg_read_keyenlock))
            tdo_tmp <= tdo_keyenlock;
    end

//program_jtagdis and read_jtagdis
    wire        tdo_jtagdis;
    wire        flg_program_jtagdis;
    wire        flg_read_jtagdis;

    reg         shift_jtagdis;

    localparam PROGRAM_JTAGDIS = 10'b01_1011_1010;
    localparam READ_JTAGDIS = 10'b01_1011_1011;

    assign flg_program_jtagdis = (update == PROGRAM_JTAGDIS);
    assign flg_read_jtagdis = (update == READ_JTAGDIS);

    always@(posedge TCK) begin
        if(rst)
            shift_jtagdis <= 0;
        else if((flg_program_jtagdis || flg_read_jtagdis) && shiftdr)
            shift_jtagdis <= TDI;
        else 
            shift_jtagdis <= shift_jtagdis;
    end

    assign tdo_jtagdis = shift_jtagdis;

    always@(negedge TCK)begin
        if(flg_shift_dr && (flg_program_jtagdis || flg_read_jtagdis))
            tdo_tmp <= tdo_jtagdis;
    end

//program_jtaglock and read_jtaglock
    wire        tdo_jtaglock;
    wire        flg_program_jtaglock;
    wire        flg_read_jtaglock;

    reg         shift_jtaglock;

    localparam PROGRAM_JTAGLOCK = 10'b01_1011_1100;
    localparam READ_JTAGLOCK = 10'b01_1011_1101;

    assign flg_program_jtaglock = (update == PROGRAM_JTAGLOCK);
    assign flg_read_jtaglock = (update == READ_JTAGLOCK);

    always@(posedge TCK) begin
        if(rst)
            shift_jtaglock <= 0;
        else if((flg_program_jtaglock || flg_read_jtaglock) && shiftdr)
            shift_jtaglock <= TDI;
        else 
            shift_jtaglock <= shift_jtaglock;
    end

    assign tdo_jtaglock = shift_jtaglock;

    always@(negedge TCK)begin
        if(flg_shift_dr && (flg_program_jtaglock || flg_read_jtaglock))
            tdo_tmp <= tdo_jtaglock;
    end

//program_scandis and read_scandis
    wire        tdo_scandis;
    wire        flg_program_scandis;
    wire        flg_read_scandis;

    reg         shift_scandis;

    localparam PROGRAM_SCANDIS = 10'b01_1011_1110;
    localparam READ_SCANDIS = 10'b01_1011_1111;

    assign flg_program_scandis = (update == PROGRAM_SCANDIS);
    assign flg_read_scandis = (update == READ_SCANDIS);

    always@(posedge TCK) begin
        if(rst)
            shift_scandis <= 0;
        else if((flg_program_scandis || flg_read_scandis) && shiftdr)
            shift_scandis <= TDI;
        else 
            shift_scandis <= shift_scandis;
    end

    assign tdo_scandis = shift_scandis;

    always@(negedge TCK)begin
        if(flg_shift_dr && (flg_program_scandis || flg_read_scandis))
            tdo_tmp <= tdo_scandis;
    end

//program_scanlock and read_scanlock
    wire        tdo_scanlock;
    wire        flg_program_scanlock;
    wire        flg_read_scanlock;

    reg         shift_scanlock;

    localparam PROGRAM_SCANLOCK = 10'b01_1100_0000;
    localparam READ_SCANLOCK = 10'b01_1100_0001;

    assign flg_program_scanlock = (update == PROGRAM_SCANLOCK);
    assign flg_read_scanlock = (update == READ_SCANLOCK);

    always@(posedge TCK) begin
        if(rst)
            shift_scanlock <= 0;
        else if((flg_program_scanlock || flg_read_scanlock) && shiftdr)
            shift_scanlock <= TDI;
        else 
            shift_scanlock <= shift_scanlock;
    end

    assign tdo_scanlock = shift_scanlock;

    always@(negedge TCK)begin
        if(flg_shift_dr &&(flg_program_scanlock || flg_read_scanlock))
            tdo_tmp <= tdo_scanlock;
    end

//program_efuseen and read_efuseen
    wire        tdo_efuseen;
    wire        flg_program_efuseen;
    wire        flg_read_efuseen;

    reg         shift_efuseen;

    localparam PROGRAM_EFUSEEN = 10'b01_1100_0010;
    localparam READ_EFUSEEN = 10'b01_1100_0011;

    assign flg_program_efuseen = (update == PROGRAM_EFUSEEN);
    assign flg_read_efuseen = (update == READ_EFUSEEN);

    always@(posedge TCK) begin
        if(rst)
            shift_efuseen <= 0;
        else if((flg_program_efuseen || flg_read_efuseen) && shiftdr)
            shift_efuseen <= TDI;
        else 
            shift_efuseen <= shift_efuseen;
    end

    assign tdo_efuseen = shift_efuseen;

    always@(negedge TCK)begin
        if(flg_shift_dr && (flg_program_efuseen || flg_read_efuseen))
            tdo_tmp <= tdo_efuseen;
    end

//program_efuselock and read_efuselock
    wire        tdo_efuselock;
    wire        flg_program_efuselock;
    wire        flg_read_efuselock;

    reg         shift_efuselock;

    localparam PROGRAM_EFUSELOCK = 10'b01_1100_0100;
    localparam READ_EFUSELOCK = 10'b01_1100_0101;

    assign flg_program_efuselock = (update == PROGRAM_EFUSELOCK);
    assign flg_read_efuselock = (update == READ_EFUSELOCK);

    always@(posedge TCK) begin
        if(rst)
            shift_efuselock <= 0;
        else if((flg_program_efuselock || flg_read_efuselock) && shiftdr)
            shift_efuselock <= TDI;
        else 
            shift_efuselock <= shift_efuselock;
    end

    assign tdo_efuselock = shift_efuselock;
    
    always@(negedge TCK) begin
        if(flg_shift_dr && (flg_program_efuselock || flg_read_efuselock))
            tdo_tmp <= tdo_efuselock;
    end

//program_id
    wire        tdo_id;
    wire        flg_program_id;

    reg [1:0]   shift_id;

    localparam PROGRAM_ID = 10'b01_1100_0110;

    assign flg_program_id = (update == PROGRAM_ID);

    always@(posedge TCK) begin
        if(rst)
            shift_id <= 0;
        else if(flg_program_id && shiftdr)
            shift_id <= {TDI, shift_id[1]};
        else 
            shift_id <= shift_id;
    end

    assign tdo_id = shift_id[0];

    always@(negedge TCK)begin
        if(flg_shift_dr && flg_program_id)
            tdo_tmp <= tdo_id;
    end

//program_idlock and read idlock
    wire        tdo_idlock;
    wire        flg_program_idlock;
    wire        flg_read_idlock;

    reg         shift_idlock;

    localparam PROGRAM_IDLOCK = 10'b01_1100_0111;
    localparam READ_IDLOCK = 10'b01_1100_1000;

    assign flg_program_idlock = (update == PROGRAM_IDLOCK);
    assign flg_read_idlock = (update == READ_IDLOCK);

    always@(posedge TCK) begin
        if(rst)
            shift_idlock <= 0;
        else if((flg_program_idlock || flg_read_idlock) && shiftdr)
            shift_idlock <= TDI;
        else 
            shift_idlock <= shift_idlock;
    end

    assign tdo_idlock = shift_idlock;

    always@(negedge TCK)begin
        if(flg_shift_dr && (flg_program_idlock || flg_read_idlock))
            tdo_tmp <= tdo_idlock;
    end

/////////////////////////////////////////////aligned 32-bit data///////////////////////////////////////////////////////

    reg [31:0]  data;
    reg [4:0]   count;
    reg         data_valid; 
    reg [4:0]   reg_cmd;
    reg         flg_desync_d;
    reg         flg_syn_reg;
    reg         flg_syn_d;
    reg         flg_syn_d2;
    reg         rstn;

    wire        flg_syn_start;
    wire        flg_desync;
    wire        desync_rose;
    wire        flg_syn;
    wire        flg_wcmemdis;
    wire        flg_rcmemdis;
    wire        cmemclk;


    always@(posedge TCK or negedge rstn)begin
        if(!rstn)begin
            data <= 0;
            data_rb <= 0;
            count <= 0;
        end
        else if(flg_cfgi && shiftdr) begin
            data = {data[30:0],TDI};
            if(flg_syn_d2)begin
                count = count + 1;
                if(count == 5'b11111)
                    data_valid = 1;
                else 
                    data_valid = 0;
            end
            else
                data_valid <= 0;
        end
        else 
            data_valid <= 0;
    end

    assign flg_syn_start = (data == 32'h0133_2d94);
    assign flg_desync = (reg_cmd == 5'b01011);
    assign flg_wcmemdis = (reg_cmd == 5'b10000);
    assign flg_rcmemdis = (reg_cmd == 5'b10001);

    always@(posedge TCK or negedge rstn)begin
        if(!rstn) begin
            reg_cmd <= 0;
            flg_desync_d <= 0;
        end
        else
            flg_desync_d <= flg_desync;
    end

    assign desync_rose = ~flg_desync_d & flg_desync;

    always@(posedge TCK or rstn) begin
        if(!rstn)
            flg_syn_reg <= 0;
        else if(flg_syn_start)
            flg_syn_reg <= 1;
        else if(desync_rose)
            flg_syn_reg <= 0;
    end

    assign flg_syn = flg_syn_start | flg_syn_reg;

    always@(posedge TCK or negedge rstn) begin
        if(!rstn)begin
            flg_syn_d <= 0;
            flg_syn_d2 <= 0;
        end
        else begin
            flg_syn_d <= flg_syn; 
            flg_syn_d2 <= flg_syn_d;
        end
    end


///////////////////////////////packet processor////////////////////////////////////////

    localparam  HEADER = 1'b0;
    localparam  DAT = 1'b1;

    wire        flg_read_tmp;
    wire        flg_write_tmp;
    wire        flg_type1;
    wire        flg_type2;
    wire [26:0] word_count_tmp;
    wire        flg_rb_reg;

    reg         s2;
    reg         ns2;
    reg [4:0]   regaddr;
    reg [26:0]  word_count;
    reg [26:0]  word_count_rb;
    reg [31:0]  data_rb_reg;
    reg         flg_write;

    initial begin
           rstn = 0;
        #2 rstn = 1;
    end
    
    assign flg_read_tmp   = ((data[28:27] == 2'b10) && data_valid && (s2 == HEADER) && flg_cfgi) | ((data[28:27] == 2'b10) && flg_cfgo);    
    assign flg_write_tmp  = ((data[28:27] == 2'b01) && data_valid && (s2 == HEADER) && flg_cfgi) |((data[28:27] == 2'b01 && flg_cfgo));
    assign flg_type1      = ((data[31:29] == 3'b101) && data_valid && (s2 == HEADER) && flg_cfgi) | ((data[31:29] == 3'b101) && flg_cfgo);
    assign flg_type2      = ((data[31:29] == 3'b010) && data_valid && (s2 == HEADER) && flg_cfgi) | ((data[31:29] == 3'b010) && flg_cfgo);
    assign word_count_tmp = (data_valid && s2 == HEADER) ? (flg_type1 ? {5'd0, data[21:0]} : data[26:0]) : word_count_tmp;

    assign flg_rb_reg = flg_cfgo & (~flg_rb_cmem);

//command
    always@(*) begin
        if(rst)
            reg_cmd = 0;
        else if(data_valid && flg_write) begin
            case(regaddr)
                5'b00010: reg_cmd <= data[4:0];
            endcase
        end
    end


//State machine to indicate HEADER or DATA for current data

    initial begin
        s2 = 0;
        ns2 = 0;
    end

    always @(posedge TCK or negedge rstn)begin
        if(!rstn)
            s2 <= HEADER;
        else if(data_valid || flg_cfgo)
            s2 <= ns2;
    end

    always @(*) begin
        if(data_valid)begin
        case(s2)
            HEADER: begin
                if(((flg_type1 || flg_type2) && (flg_read_tmp || flg_write_tmp)) && (word_count_tmp != 27'd0))
                    ns2 = DAT;
                else
                    ns2 = HEADER;
            end

            DAT:  begin
                if((data_valid && (word_count == 27'd0)) || (flg_cfgo && (word_count_rb == 27'd0)))
                    ns2 = HEADER;
                else
                    ns2 = DAT;
            end
        endcase
        end
    end

//get address
    always @(negedge TCK or negedge rstn) begin
        if(!rstn)
            regaddr <= 5'd0;
        else if((data_valid || flg_cfgi) && (s2 == HEADER) && flg_type1 && (flg_read_tmp || flg_write_tmp))
            regaddr <= data[26:22];
    end

//write flag
    always @(negedge TCK or negedge rstn) begin
        if(!rstn)
            flg_write <= 1'b0;
        else if(data_valid) begin
            if((s2 == HEADER) && (flg_type1 || flg_type2) && flg_write_tmp && (word_count_tmp != 27'd0))
                flg_write <= 1'b1;
            else if(word_count == 27'd0)
                flg_write <= 1'b0;
        end
    end

//write operation count
    always @(negedge TCK or negedge rstn) begin
        if(!rstn)
            word_count <= 27'd0;
        else if(data_valid) begin
            if((s2 == HEADER) && (flg_type1 || flg_type2) && flg_write_tmp && (word_count_tmp != 27'd0))begin
                if(regaddr == 5'b00101 && reg_cmd == 5'b00100)
                    word_count <= word_count_tmp;
                else
                    word_count <= word_count_tmp - 1'b1;
            end
            else if((s2 == DAT) && (word_count != 27'd0))
                word_count <= word_count - 1'b1;
            else
                word_count <= 27'd0;
        end
    end

////////////////////////////////////////////////////////readback cmem/////////////////////////////////////////////////////

    wire        flg_rcmem;


//cmem readback count
    always @(posedge TCK or negedge rstn) begin
        if(!rstn)
            word_count_rb <= 27'd0;
        else if(flg_cfgi && (s2 == HEADER) && (flg_type1 || flg_type2) && flg_read_tmp && (word_count_tmp != 27'd0) && flg_rcmem)
            word_count_rb <= word_count_tmp - 1'b1;
        else if((flg_cfgo || flg_rb_reg) && (word_count_rb != 27'd0))
            word_count_rb <= word_count_rb - 1'b1;
    end

//cmem readback flag

    assign flg_rcmem   = (reg_cmd == 5'b00110);//read cmem, 
    always @(posedge TCK or negedge rstn) begin
        if(!rstn)
            flg_rb_cmem <= 1'b0;
        else if(flg_cfgi) begin
                if((s2 == HEADER) && (flg_type1 || flg_type2) && flg_read_tmp && (word_count_tmp != 27'd0) && flg_rcmem && (regaddr == 5'b0_0111))
                    flg_rb_cmem <= 1'b1;
                else if(word_count_rb == 27'd0)
                    flg_rb_cmem <= 1'b0;
        end
    end


    reg     [31:0]  reg_cmemor;

    always@(*) begin
        if(flg_cfgo) begin
            if(flg_rb_reg && !flg_rb_cmem)
                data_rb = data_rb_reg;
            else if(flg_rb_cmem && !flg_rb_reg)
                data_rb = reg_cmemor;
            else 
                data_rb = 32'hFFFF_FFFF;
        end
        else begin
            data_rb = 32'hFFFF_FFFF;
        end
    end

//////////////////////////////////////////////////reg array////////////////////////////////////////////////////////////////////

    reg     [31:0]  reg_idr;
    reg     [31:0]  reg_cmdr;
    reg     [31:0]  reg_cmemir;
    reg     [31:0]  reg_adrr;


    always@(*) begin
        if(!rstn) begin 
            reg_idr <= 0;
            reg_cmdr <= 0;
            reg_cmemir <= 0;
            reg_adrr <= 0;
            reg_cmemor <= 0;
        end
        else begin
            if(data_valid && flg_write && (s2 == DAT)) begin
                case(regaddr)
                5'b00010 : reg_cmdr <= data;
                5'b00101 : reg_cmemir <= data;
                5'b01011 : reg_adrr <= data;
                endcase
            end
            else if(flg_cfgo && flg_rb_reg) begin
                case(regaddr)
                5'b00001 : data_rb_reg <= IDCODE;
                5'b00010 : data_rb_reg <= reg_cmdr;
                5'b00111 : data_rb_reg <= reg_cmemor;
                5'b01011 : data_rb_reg <= reg_adrr;
                default  : data_rb_reg <= 32'hFFFF_FFFF;
                endcase                
            end
        end                    
    end

////////////////////////////////////////////////cmem///////////////////////////////////////////////

    wire            we;
    wire    [1:0]   cmemtype;
    wire    [4:0]   addr_region;
    wire    [7:0]   addr_column;
    wire    [7:0]   addr_frame;
    reg     [5:0]   count32;
    reg             flg_count32;

    assign cmemclk = (flg_cfgi & data_valid) | (flg_cfgo & flg_count32);
    assign we = (flg_write == 1 && regaddr == 5'b00101 && reg_cmd == 5'b00100 && s2 == DAT) ? 1'b1 : 1'b0;
    assign cmemtype = reg_adrr[26:25];
    assign addr_region = reg_adrr[24:20];
    assign addr_column = reg_adrr[17:10];
    assign addr_frame = reg_adrr[7:0];


////////////////////////////////////////////////cmem_e2////////////////////////////////////////////////

    integer i;
    reg [3231:0] cmem [0:7327];
    reg [13:0] addr_row;
    reg [13:0] naddr_row;
    reg [6:0] addr_word;
    always@(posedge TCK or negedge rstn) begin
        if(!rstn) begin
            count32 <= 0;
            flg_count32 <= 0;
        end
        else if(flg_rb_cmem && flg_cfgo && shiftdr) begin
            count32 = count32 + 1;
            if(count32 == 32) begin
                flg_count32 <= 1;
                count32 <= 0;
            end
            else 
                flg_count32 <= 0;
        end

    end

    always@(negedge shiftdr) begin
        count32 <= 0;
        flg_count32 <= 0;
    end

    always@(*) begin
        if(flg_count32)
            shift_cfgo2 <= data_rb;
    end

    always@(posedge cmemclk or negedge rstn) begin
        if(!rstn) begin
            addr_word <= 0; 
            for(i = 0; i < 7328; i = i + 1)
                cmem[i] <= 0;
        end
        else if(we || (flg_rb_cmem && flg_cfgo && shiftdr)) begin
            addr_word <= addr_word + 1;
            if(addr_word == 100) begin
                addr_word <= 0; 
                reg_adrr[7:0] <= reg_adrr[7:0] + 1;//addr_frame + 1
            end
        end
        else
            addr_word <= 0;
    end


    always@(negedge TCK) begin
            if(we && data_valid) begin
                    cmem[addr_row][addr_word*32] <= reg_cmemir[0];
                    cmem[addr_row][addr_word*32 + 1] <= reg_cmemir[1];
                    cmem[addr_row][addr_word*32 + 2] <= reg_cmemir[2];
                    cmem[addr_row][addr_word*32 + 3] <= reg_cmemir[3];
                    cmem[addr_row][addr_word*32 + 4] <= reg_cmemir[4];
                    cmem[addr_row][addr_word*32 + 5] <= reg_cmemir[5];
                    cmem[addr_row][addr_word*32 + 6] <= reg_cmemir[6];
                    cmem[addr_row][addr_word*32 + 7] <= reg_cmemir[7];
                    cmem[addr_row][addr_word*32 + 8] <= reg_cmemir[8];
                    cmem[addr_row][addr_word*32 + 9] <= reg_cmemir[9];
                    cmem[addr_row][addr_word*32 + 10] <= reg_cmemir[10];
                    cmem[addr_row][addr_word*32 + 11] <= reg_cmemir[11];
                    cmem[addr_row][addr_word*32 + 12] <= reg_cmemir[12];
                    cmem[addr_row][addr_word*32 + 13] <= reg_cmemir[13];
                    cmem[addr_row][addr_word*32 + 14] <= reg_cmemir[14];
                    cmem[addr_row][addr_word*32 + 15] <= reg_cmemir[15];
                    cmem[addr_row][addr_word*32 + 16] <= reg_cmemir[16];
                    cmem[addr_row][addr_word*32 + 17] <= reg_cmemir[17];
                    cmem[addr_row][addr_word*32 + 18] <= reg_cmemir[18];
                    cmem[addr_row][addr_word*32 + 19] <= reg_cmemir[19];
                    cmem[addr_row][addr_word*32 + 20] <= reg_cmemir[20];
                    cmem[addr_row][addr_word*32 + 21] <= reg_cmemir[21];
                    cmem[addr_row][addr_word*32 + 22] <= reg_cmemir[22];
                    cmem[addr_row][addr_word*32 + 23] <= reg_cmemir[23];
                    cmem[addr_row][addr_word*32 + 24] <= reg_cmemir[24];
                    cmem[addr_row][addr_word*32 + 25] <= reg_cmemir[25];
                    cmem[addr_row][addr_word*32 + 26] <= reg_cmemir[26];
                    cmem[addr_row][addr_word*32 + 27] <= reg_cmemir[27];
                    cmem[addr_row][addr_word*32 + 28] <= reg_cmemir[28];
                    cmem[addr_row][addr_word*32 + 29] <= reg_cmemir[29];
                    cmem[addr_row][addr_word*32 + 30] <= reg_cmemir[30];
                    cmem[addr_row][addr_word*32 + 31] <= reg_cmemir[31];
                end
                else if(flg_rcmem && cmemclk && shiftdr) begin//flg_rb_cmem
                    reg_cmemor[0] <=  cmem[addr_row][addr_word*32];
                    reg_cmemor[1] <=  cmem[addr_row][addr_word*32 + 1];
                    reg_cmemor[2] <=  cmem[addr_row][addr_word*32 + 2];
                    reg_cmemor[3] <=  cmem[addr_row][addr_word*32 + 3];
                    reg_cmemor[4] <=  cmem[addr_row][addr_word*32 + 4];
                    reg_cmemor[5] <=  cmem[addr_row][addr_word*32 + 5];
                    reg_cmemor[6] <=  cmem[addr_row][addr_word*32 + 6];
                    reg_cmemor[7] <=  cmem[addr_row][addr_word*32 + 7];
                    reg_cmemor[8] <=  cmem[addr_row][addr_word*32 + 8];
                    reg_cmemor[9] <=  cmem[addr_row][addr_word*32 + 9];
                    reg_cmemor[10] <= cmem[addr_row][addr_word*32 + 10];
                    reg_cmemor[11] <= cmem[addr_row][addr_word*32 + 11];
                    reg_cmemor[12] <= cmem[addr_row][addr_word*32 + 12];
                    reg_cmemor[13] <= cmem[addr_row][addr_word*32 + 13];
                    reg_cmemor[14] <= cmem[addr_row][addr_word*32 + 14];
                    reg_cmemor[15] <= cmem[addr_row][addr_word*32 + 15];
                    reg_cmemor[16] <= cmem[addr_row][addr_word*32 + 16];
                    reg_cmemor[17] <= cmem[addr_row][addr_word*32 + 17];
                    reg_cmemor[18] <= cmem[addr_row][addr_word*32 + 18];
                    reg_cmemor[19] <= cmem[addr_row][addr_word*32 + 19];
                    reg_cmemor[20] <= cmem[addr_row][addr_word*32 + 20];
                    reg_cmemor[21] <= cmem[addr_row][addr_word*32 + 21];
                    reg_cmemor[22] <= cmem[addr_row][addr_word*32 + 22];
                    reg_cmemor[23] <= cmem[addr_row][addr_word*32 + 23];
                    reg_cmemor[24] <= cmem[addr_row][addr_word*32 + 24];
                    reg_cmemor[25] <= cmem[addr_row][addr_word*32 + 25];
                    reg_cmemor[26] <= cmem[addr_row][addr_word*32 + 26];
                    reg_cmemor[27] <= cmem[addr_row][addr_word*32 + 27];
                    reg_cmemor[28] <= cmem[addr_row][addr_word*32 + 28];
                    reg_cmemor[29] <= cmem[addr_row][addr_word*32 + 29];
                    reg_cmemor[30] <= cmem[addr_row][addr_word*32 + 30];
                    reg_cmemor[31] <= cmem[addr_row][addr_word*32 + 31];
                end
                else 
                    ;        
    end

    always@(posedge we) begin
        addr_word <= 0;
    end

    always@(negedge we) begin
        $writememb("cmem.txt", cmem);
    end

    always@(posedge flg_rb_cmem) begin
        $readmemb("cmem.txt", cmem);  
        addr_word <= 0;
    end
    

    always@(*)begin
        case(addr_region)
            0:  case (addr_column)
                    0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46: begin
                        if(addr_frame < 36)
                            addr_row = 0 + 36* addr_column + addr_frame;
                        else if(addr_frame == 36) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end
                    47, 48, 49, 50: begin
                        if(addr_frame < 28)
                            naddr_row = 0 + 36*47 + 28*(addr_column - 47) + addr_frame - 1;
                        else if(addr_frame == 28) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end    
                    51, 52, 53: begin
                        if(addr_frame < 28)
                            addr_row = 0 + 36*47 + 28*4 + 28*(addr_column - 51) + addr_frame - 1;
                        else if(addr_frame == 28) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end  
                    54: begin
                        if(addr_frame < 34)
                            addr_row = 0 + 36*47 + 28*4 + 28*3 + 34*(addr_column - 54) + addr_frame - 1;
                        else if(addr_frame == 34) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end 
                    55: begin
                        if(addr_frame < 2)
                            addr_row = 0 + 36*47 + 28*4 + 28*3 + 34*1 + 2*(addr_column - 55) + addr_frame - 1;
                        else if(addr_frame == 2) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end 

                    56, 57: begin
                        if(addr_frame < 28)
                            addr_row = 0 + 36*47 + 28*4 + 28*3 + 34*1 + 2*1 + 28*(addr_column - 56) + addr_frame - 1;
                        else if(addr_frame == 28) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end 
                    58: begin
                        if(addr_frame < 28)
                            addr_row = 0 + 36*47 + 28*4 + 28*3 + 34*1 + 2*1 + 28*2 + 28*(addr_column - 58) + addr_frame - 1;
                        else if(addr_frame == 28) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = 0;
                            reg_adrr[24:20] = 1;
                        end
                    end 
                endcase
            1:  case(addr_column)
                    0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36:begin
                        if(addr_frame < 36)
                            addr_row = 2008 + 36*addr_column + addr_frame;
                        else if(addr_frame == 36)begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end
                    37, 38, 39, 40: begin
                        if(addr_frame < 28)
                            addr_row = 2008 + 36*37 + 28*(addr_column - 37) + addr_frame - 1;
                        else if(addr_frame == 28) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end
                    41, 42, 43: begin
                        if(addr_frame < 28)
                            addr_row = 2008 + 36*37 + 28*4 + 28*(addr_column - 41) + addr_frame - 1;
                        else if(addr_frame == 28) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end
                    44, 45: begin
                        if(addr_frame < 34)
                            addr_row = 2008 + 36*37 + 28*4 + 28*3 + 34*(addr_column - 44) + addr_frame - 1;
                        else if(addr_frame == 34)begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end
                    46, 47: begin
                        if(addr_frame < 2)
                            addr_row = 2008 + 36*37 + 28*4 + 28*3 + 34*2 + 2*(addr_column - 46) + addr_frame - 1;
                        else if(addr_frame == 2) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end
                    48, 49: begin 
                        if(addr_frame < 28)
                            addr_row = 2008 + 36*37 + 28*4 + 28*3 + 34*2 + 2*2 + 28*(addr_column - 48) + addr_frame - 1;
                        else if(addr_frame == 28) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                            if(addr_column == 49) begin
                                reg_adrr[17:10] = 0;
                                reg_adrr[24:20] = 2;
                            end
                        end   
                    end             
                endcase
            2:  case(addr_column)
                    0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36:begin
                        if(addr_frame < 36)
                            addr_row = 3664 + 36*addr_column + addr_frame;
                        else if(addr_frame == 36)begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end
                    37, 38, 39, 40: begin
                        if(addr_frame < 28)
                            addr_row = 3664 + 36*37 + 28*(addr_column - 37) + addr_frame - 1;
                        else if(addr_frame == 28) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end
                    41, 42, 43: begin
                        if(addr_frame < 28)
                            addr_row = 3664 + 36*37 + 28*4 + 28*(addr_column - 41) + addr_frame - 1;
                        else if(addr_frame == 28) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end
                    44, 45: begin
                        if(addr_frame < 34)
                            addr_row = 3664 + 36*37 + 28*4 + 28*3 + 34*(addr_column - 44) + addr_frame - 1;
                        else if(addr_frame == 34)begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end
                    46, 47: begin
                        if(addr_frame < 2)
                            addr_row = 3664 + 36*37 + 28*4 + 28*3 + 34*2 + 2*(addr_column - 46) + addr_frame - 1;
                        else if(addr_frame == 2) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end
                    48, 49: begin 
                        if(addr_frame < 28)
                            addr_row = 3664 + 36*37 + 28*4 + 28*3 + 34*2 + 2*2 + 28*(addr_column - 48) + addr_frame - 1;
                        else if(addr_frame == 28) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                            if(addr_column == 49) begin
                                reg_adrr[17:10] = 0;
                                reg_adrr[24:20] = 3;
                            end
                        end   
                    end             
                endcase

            3:  case (addr_column)
                    0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46: begin
                        if(addr_frame < 36)
                            addr_row = 5320 + 36* addr_column + addr_frame;
                        else if(addr_frame == 36) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end
                    47, 48, 49, 50: begin
                        if(addr_frame < 28)
                            addr_row = 5320 + 36*47 + 28*(addr_column - 47) + addr_frame - 1;
                        else if(addr_frame == 28) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end    
                    51, 52, 53: begin
                        if(addr_frame < 28)
                            addr_row = 5320 + 36*47 + 28*4 + 28*(addr_column - 51) + addr_frame - 1;
                        else if(addr_frame == 28) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end  
                    54: begin
                        if(addr_frame < 34)
                            addr_row = 5320 + 36*47 + 28*4 + 28*3 + 34*(addr_column - 54) + addr_frame - 1;
                        else if(addr_frame == 34) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end 
                    55: begin
                        if(addr_frame < 2)
                            addr_row = 5320 + 36*47 + 28*4 + 28*3 + 34*1 + 2*(addr_column - 55) + addr_frame - 1;
                        else if(addr_frame == 2) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end 

                    56, 57: begin
                        if(addr_frame < 28)
                            addr_row = 5320 + 36*47 + 28*4 + 28*3 + 34*1 + 2*1 + 28*(addr_column - 56) + addr_frame - 1;
                        else if(addr_frame == 28) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = reg_adrr[17:10] + 1;
                        end
                    end 
                    58: begin
                        if(addr_frame < 28)
                            addr_row = 5320 + 36*47 + 28*4 + 28*3 + 34*1 + 2*1 + 28*2 + 28*(addr_column - 58) + addr_frame - 1;
                        else if(addr_frame == 28) begin
                            reg_adrr[7:0] = 0;
                            reg_adrr[17:10] = 0;
                        end
                    end 
                endcase

        endcase
    end


//synthesis translate_on
endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2018 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_PLL_E3.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1ns/10fs
module GTP_PLL_E3 #(
    parameter real CLKIN_FREQ = 50.0,
    parameter PFDEN_EN        = "FALSE", //"TRUE"; "FALSE"
    parameter VCOCLK_DIV2     = 1'b0,    //1'b0~1'b1
    parameter DYNAMIC_RATIOI_EN = "FALSE", //"TRUE"; "FALSE"
    parameter DYNAMIC_RATIOM_EN = "FALSE", //"TRUE"; "FALSE"
    parameter DYNAMIC_RATIO0_EN = "FALSE", //"TRUE"; "FALSE"
    parameter DYNAMIC_RATIO1_EN = "FALSE", //"TRUE"; "FALSE"
    parameter DYNAMIC_RATIO2_EN = "FALSE", //"TRUE"; "FALSE"
    parameter DYNAMIC_RATIO3_EN = "FALSE", //"TRUE"; "FALSE"
    parameter DYNAMIC_RATIO4_EN = "FALSE", //"TRUE"; "FALSE"
    parameter DYNAMIC_RATIOF_EN = "FALSE", //"TRUE"; "FALSE"
    parameter integer STATIC_RATIOI = 1, //1~512
    parameter integer STATIC_RATIOM = 1, //1~64
    parameter integer STATIC_RATIO0 = 1, //1~512
    parameter integer STATIC_RATIO1 = 1, //1~512
    parameter integer STATIC_RATIO2 = 1, //1~512
    parameter integer STATIC_RATIO3 = 1, //1~512
    parameter integer STATIC_RATIO4 = 1, //1~512
    parameter integer STATIC_RATIOF = 1, //1~512
    parameter DYNAMIC_DUTY0_EN = "FALSE", //"TRUE"; "FALSE"
    parameter DYNAMIC_DUTY1_EN = "FALSE", //"TRUE"; "FALSE"
    parameter DYNAMIC_DUTY2_EN = "FALSE", //"TRUE"; "FALSE"
    parameter DYNAMIC_DUTY3_EN = "FALSE", //"TRUE"; "FALSE"
    parameter DYNAMIC_DUTY4_EN = "FALSE", //"TRUE"; "FALSE"
    parameter integer STATIC_DUTY0 = 2, //2<=STATIC_DUTY0<=2*STATIC_RATIO0-2
    parameter integer STATIC_DUTY1 = 2, //2<=STATIC_DUTY1<=2*STATIC_RATIO1-2
    parameter integer STATIC_DUTY2 = 2, //2<=STATIC_DUTY2<=2*STATIC_RATIO2-2
    parameter integer STATIC_DUTY3 = 2, //2<=STATIC_DUTY3<=2*STATIC_RATIO3-2
    parameter integer STATIC_DUTY4 = 2, //2<=STATIC_DUTY4<=2*STATIC_RATIO4-2
    parameter integer STATIC_PHASE0  = 0, //0~7
    parameter integer STATIC_PHASE1  = 0, //0~7
    parameter integer STATIC_PHASE2  = 0, //0~7
    parameter integer STATIC_PHASE3  = 0, //0~7
    parameter integer STATIC_PHASE4  = 0, //0~7
    parameter integer STATIC_PHASEF  = 0, //0~7
    parameter integer STATIC_CPHASE0 = 0, //0~511
    parameter integer STATIC_CPHASE1 = 0, //0~511
    parameter integer STATIC_CPHASE2 = 0, //0~511
    parameter integer STATIC_CPHASE3 = 0, //0~511
    parameter integer STATIC_CPHASE4 = 0, //0~511
    parameter integer STATIC_CPHASEF = 0, //0~511
    parameter CLK_CAS1_EN = "FALSE", //"TRUE"; "FALSE"
    parameter CLK_CAS2_EN = "FALSE", //"TRUE"; "FALSE"
    parameter CLK_CAS3_EN = "FALSE", //"TRUE"; "FALSE"
    parameter CLK_CAS4_EN = "FALSE", //"TRUE"; "FALSE"
    parameter integer CLKOUT5_SEL = 0, //0~4
    parameter CLKIN_BYPASS_EN     = "FALSE", //"TRUE"; "FALSE"
    parameter CLKOUT0_SYN_EN      = "FALSE", //"TRUE"; "FALSE"
    parameter CLKOUT0_EXT_SYN_EN  = "FALSE", //"TRUE"; "FALSE"
    parameter CLKOUT1_SYN_EN      = "FALSE", //"TRUE"; "FALSE"
    parameter CLKOUT2_SYN_EN      = "FALSE", //"TRUE"; "FALSE"
    parameter CLKOUT3_SYN_EN      = "FALSE", //"TRUE"; "FALSE"
    parameter CLKOUT4_SYN_EN      = "FALSE", //"TRUE"; "FALSE"
    parameter CLKOUT5_SYN_EN      = "FALSE", //"TRUE"; "FALSE"
    parameter INTERNAL_FB = "ENABLE",  //"ENABLE"; "DISABLE"
    parameter EXTERNAL_FB = "DISABLE", //"CLKOUT0"; "CLKOUT1"; "CLKOUT2"; "CLKOUT3"; "CLKOUT4"; "DISABLE";
    parameter DYNAMIC_LOOP_EN = "FALSE", //"TRUE"; "FALSE"
    parameter LOOP_MAPPING_EN = "FALSE", //"TRUE"; "FALSE"
    parameter BANDWIDTH = "OPTIMIZED"    //"LOW"; "OPTIMIZED"; "HIGH"
    )(
    output CLKOUT0,
    output CLKOUT0_EXT,
    output CLKOUT1,
    output CLKOUT2,
    output CLKOUT3,
    output CLKOUT4,
    output CLKOUT5,
    output CLKSWITCH_FLAG,
    output LOCK,
    input CLKIN1,
    input CLKIN2,
    input CLKFB,
    input CLKIN_SEL,
    input CLKIN_SEL_EN,
    input PFDEN,
    input ICP_BASE,
    input [3:0] ICP_SEL,
    input [2:0] LPFRES_SEL,
    input CRIPPLE_SEL,
    input [2:0] PHASE_SEL,
    input PHASE_DIR,
    input PHASE_STEP_N,
    input LOAD_PHASE,
    input [9:0] RATIOI,
    input [6:0] RATIOM,
    input [9:0] RATIO0,
    input [9:0] RATIO1,
    input [9:0] RATIO2,
    input [9:0] RATIO3,
    input [9:0] RATIO4,
    input [9:0] RATIOF,
    input [9:0] DUTY0,
    input [9:0] DUTY1,
    input [9:0] DUTY2,
    input [9:0] DUTY3,
    input [9:0] DUTY4,
    input CLKOUT0_SYN,
    input CLKOUT0_EXT_SYN,
    input CLKOUT1_SYN,
    input CLKOUT2_SYN,
    input CLKOUT3_SYN,
    input CLKOUT4_SYN,
    input CLKOUT5_SYN,
    input PLL_PWD,
    input RST,
    input RSTODIV
    )/* synthesis syn_black_box */;

    initial
    begin
        if((PFDEN_EN == "TRUE") || (PFDEN_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E3 error: illegal setting for PFDEN_EN");

        if((DYNAMIC_RATIOI_EN == "TRUE") || (DYNAMIC_RATIOI_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E3 error: illegal setting for DYNAMIC_RATIOI_EN");

        if((DYNAMIC_RATIOM_EN == "TRUE") || (DYNAMIC_RATIOM_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E3 error: illegal setting for DYNAMIC_RATIOM_EN");

        if((DYNAMIC_RATIO0_EN == "TRUE") || (DYNAMIC_RATIO0_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E3 error: illegal setting for DYNAMIC_RATIO0_EN");

        if((DYNAMIC_RATIO1_EN == "TRUE") || (DYNAMIC_RATIO1_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E3 error: illegal setting for DYNAMIC_RATIO1_EN");

        if((DYNAMIC_RATIO2_EN == "TRUE") || (DYNAMIC_RATIO2_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E3 error: illegal setting for DYNAMIC_RATIO2_EN");

        if((DYNAMIC_RATIO3_EN == "TRUE") || (DYNAMIC_RATIO3_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E3 error: illegal setting for DYNAMIC_RATIO3_EN");

        if((DYNAMIC_RATIO4_EN == "TRUE") || (DYNAMIC_RATIO4_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E3 error: illegal setting for DYNAMIC_RATIO4_EN");

        if((DYNAMIC_RATIOF_EN == "TRUE") || (DYNAMIC_RATIOF_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E3 error: illegal setting for DYNAMIC_RATIOF_EN");

        if((DYNAMIC_DUTY0_EN == "TRUE") || (DYNAMIC_DUTY0_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E3 error: illegal setting for DYNAMIC_DUTY0_EN");

        if((DYNAMIC_DUTY1_EN == "TRUE") || (DYNAMIC_DUTY1_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E3 error: illegal setting for DYNAMIC_DUTY1_EN");

        if((DYNAMIC_DUTY2_EN == "TRUE") || (DYNAMIC_DUTY2_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E3 error: illegal setting for DYNAMIC_DUTY2_EN");

        if((DYNAMIC_DUTY3_EN == "TRUE") || (DYNAMIC_DUTY3_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E3 error: illegal setting for DYNAMIC_DUTY3_EN");

        if((DYNAMIC_DUTY4_EN == "TRUE") || (DYNAMIC_DUTY4_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E3 error: illegal setting for DYNAMIC_DUTY4_EN");

        if((CLK_CAS1_EN == "TRUE") || (CLK_CAS1_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E3 error: illegal setting for CLK_CAS1_EN");

        if((CLK_CAS2_EN == "TRUE") || (CLK_CAS2_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E3 error: illegal setting for CLK_CAS2_EN");

        if((CLK_CAS3_EN == "TRUE") || (CLK_CAS3_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E3 error: illegal setting for CLK_CAS3_EN");

        if((CLK_CAS4_EN == "TRUE") || (CLK_CAS4_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E3 error: illegal setting for CLK_CAS4_EN");

        if((CLKIN_BYPASS_EN == "TRUE") || (CLKIN_BYPASS_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E3 error: illegal setting for CLKIN_BYPASS_EN");

        if((CLKOUT0_SYN_EN == "TRUE") || (CLKOUT0_SYN_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E3 error: illegal setting for CLKOUT0_SYN_EN");

        if((CLKOUT0_EXT_SYN_EN == "TRUE") || (CLKOUT0_EXT_SYN_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E3 error: illegal setting for CLKOUT0_EXT_SYN_EN");

        if((CLKOUT1_SYN_EN == "TRUE") || (CLKOUT1_SYN_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E3 error: illegal setting for CLKOUT1_SYN_EN");

        if((CLKOUT2_SYN_EN == "TRUE") || (CLKOUT2_SYN_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E3 error: illegal setting for CLKOUT2_SYN_EN");

        if((CLKOUT3_SYN_EN == "TRUE") || (CLKOUT3_SYN_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E3 error: illegal setting for CLKOUT3_SYN_EN");

        if((CLKOUT4_SYN_EN == "TRUE") || (CLKOUT4_SYN_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E3 error: illegal setting for CLKOUT4_SYN_EN");

        if((CLKOUT5_SYN_EN == "TRUE") || (CLKOUT5_SYN_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E3 error: illegal setting for CLKOUT5_SYN_EN");

        if((INTERNAL_FB == "ENABLE") || (INTERNAL_FB == "DISABLE"))
        begin
        end
        else
            $display ("GTP_PLL_E3 error: illegal setting for INTERNAL_FB");

        if((EXTERNAL_FB == "CLKOUT0") || (EXTERNAL_FB == "CLKOUT1") || (EXTERNAL_FB == "CLKOUT2") || (EXTERNAL_FB == "CLKOUT3") || (EXTERNAL_FB == "CLKOUT4") || (EXTERNAL_FB == "DISABLE"))
        begin
        end
        else
            $display ("GTP_PLL_E3 error: illegal setting for EXTERNAL_FB");

        if((BANDWIDTH == "LOW") || (BANDWIDTH == "OPTIMIZED") || (BANDWIDTH == "HIGH"))
        begin
        end
        else
            $display ("GTP_PLL_E3 error: illegal setting for BANDWIDTH");

        if((DYNAMIC_LOOP_EN == "TRUE") || (DYNAMIC_LOOP_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E3 error: illegal setting for DYNAMIC_LOOP_EN");

        if((LOOP_MAPPING_EN == "TRUE") || (LOOP_MAPPING_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E3 error: illegal setting for LOOP_MAPPING_EN");
    end
///////////////////////////////////////////////////////
    wire rst_n, rstodiv_n;
///////////////////////////////////////////////////////
    wire clk_sel, clk_in, clk0, clk1, rstclksw_n;
    reg [1:0] cnt0, cnt1;
    reg dynauto_clkin;
///////////////////////////////////////////////////////
    reg clk_in_first_time, clk_fb_first_time;
    realtime clk_in_first_edge, clk_fb_first_edge;
    reg adjust;
    realtime fb_route_delay, virtual_delay1;
    integer tmp_ratio;
    realtime tmp_delay, real_delay;
///////////////////////////////////////////////////////
    wire pfden;
    reg [1:0] pfd_en_reg;
    reg clk_pfd, vcolow;
    integer cnt;

    reg clk_test, clkwo;
    realtime clk_test_time1 , clk_test_time2, clk_test_time3;
///////////////////////////////////////////////////////
    wire [9:0] idivider, divider0, divider1, divider2, divider3, divider4, fdivider;
    wire [6:0] mdivider;
    real fsdiv_set_int, fbdiv_set_int;
    reg [5:0] fbdiv_sel;
    integer prop;

    wire rstanalog_n;
    realtime clkin_rtime_last, clkin_rtime_next;
    realtime clkin_time, clkin_time1, clkin_time2, clkin_time3;
    reg clkout_lock;
    realtime vcoclk_period, vcoclk_period_half;
    realtime clkout0_time, clkout1_time, clkout2_time, clkout3_time, clkout4_time;
    integer  vcoclk_period_amp;
    realtime vcoclk_period_real, vcoclk_period_dev;

    reg done;
    integer idiv_set;
    integer fdiv_set;
    integer swap_set;
    integer fdiv_int;
    realtime offset;

    real cnt_fdiv;
    reg clk_gate, inner_clk;
    reg vcoclk;
    reg clk_vcodiv2;
    wire clkout;
///////////////////////////////////////////////////////
    wire clk_lock;
    reg [2:0] cnt_clkfb;
    reg start_clk;
    reg [10:0] cnt_lock;
    reg lock_reg;
///////////////////////////////////////////////////////
    wire clk_sel0, clk_sel1, clk_sel2, clk_sel3, clk_sel4;
    wire odiv0_rstn, odiv1_rstn, odiv2_rstn, odiv3_rstn, odiv4_rstn;
    wire [9:0] odiv0_duty, odiv1_duty, odiv2_duty, odiv3_duty, odiv4_duty;
    wire [9:0] odiv0_duty_ctrl, odiv1_duty_ctrl, odiv2_duty_ctrl, odiv3_duty_ctrl, odiv4_duty_ctrl;
    reg [2:0] enclk0, enclk1, enclk2, enclk3, enclk4;
    wire clk_en0, clk_en1, clk_en2, clk_en3, clk_en4;
    reg [9:0] odiv0_counter, odiv1_counter, odiv2_counter, odiv3_counter, odiv4_counter;
    reg odiv0_clkdivr, odiv1_clkdivr, odiv2_clkdivr, odiv3_clkdivr, odiv4_clkdivr;
    reg odiv0_set, odiv1_set, odiv2_set, odiv3_set, odiv4_set;
    wire odiv0_out, odiv1_out, odiv2_out, odiv3_out, odiv4_out;
///////////////////////////////////////////////////////
    reg fphase_step, last_fphase_step;
    integer step_odiv0, step_odiv1, step_odiv2, step_odiv3, step_odiv4;
    integer step_odiv0_1, step_odiv1_1, step_odiv2_1, step_odiv3_1, step_odiv4_1;
    integer step_odiv0_2, step_odiv1_2, step_odiv2_2, step_odiv3_2, step_odiv4_2;
    integer step_odiv0_3, step_odiv1_3, step_odiv2_3, step_odiv3_3, step_odiv4_3;
    integer step_odiv0_4, step_odiv1_4, step_odiv2_4, step_odiv3_4, step_odiv4_4;
    integer step_odiv0_5, step_odiv1_5, step_odiv2_5, step_odiv3_5, step_odiv4_5;

    realtime vco_fphase_delay0, vco_fphase_delay1, vco_fphase_delay2, vco_fphase_delay3, vco_fphase_delay4;
    integer phase0, phase1, phase2, phase3, phase4;
    realtime cphase_delay0, cphase_delay1, cphase_delay2, cphase_delay3, cphase_delay4;
    reg odiv0_out_delay1, odiv1_out_delay1, odiv2_out_delay1, odiv3_out_delay1, odiv4_out_delay1;
    reg odiv0_out_delay, odiv1_out_delay, odiv2_out_delay, odiv3_out_delay, odiv4_out_delay;
///////////////////////////////////////////////////////
    reg [2:0] clk_out0_gate, clk_out0_ext_gate, clk_out1_gate, clk_out2_gate, clk_out3_gate, clk_out4_gate, clk_out5_gate;
    reg clk_out5_reg;
    wire clkout0_en, clkout0_ext_en, clkout1_en, clkout1_adc_en, clkout2_en, clkout3_en, clkout4_en, clkout5_en, clkout4_sel;
    reg inner_rstn;
///////////////////////////////////////////////////////
    initial
    begin
        cnt0 = 2'b00;
        cnt1 = 2'b00;
        dynauto_clkin = 1'b0;
        clk_in_first_time = 1'b0;
        clk_fb_first_time = 1'b0;
        clk_in_first_edge = 0.0;
        clk_fb_first_edge = 0.0;
        fb_route_delay = 0.0;
        tmp_ratio = 0;
        tmp_delay = 0.0;
        real_delay = 0.0;
        clk_pfd  = 1'b0;
        clk_test = 1'b0;
        fsdiv_set_int = 0;
        fbdiv_set_int = 0;
        fbdiv_sel     = 6'b000001;
        done = 1'b0;
        idiv_set = 0;
        fdiv_set = 0;
        swap_set = 0;
        fdiv_int = 0;
        offset = 0;
        cnt_fdiv  = 0;
        clk_gate  = 1'b1;
        inner_clk = 1'b0;
        vcoclk    = 1'b0;
        fphase_step = 1'b0;
        last_fphase_step = 1'b0;
        step_odiv0 = 0;
        step_odiv1 = 0;
        step_odiv2 = 0;
        step_odiv3 = 0;
        step_odiv4 = 0;
        step_odiv0_1 = STATIC_PHASE0;
        step_odiv1_1 = STATIC_PHASE1;
        step_odiv2_1 = STATIC_PHASE2;
        step_odiv3_1 = STATIC_PHASE3;
        step_odiv4_1 = STATIC_PHASE4;
        step_odiv0_2 = STATIC_PHASE0;
        step_odiv1_2 = STATIC_PHASE1;
        step_odiv2_2 = STATIC_PHASE2;
        step_odiv3_2 = STATIC_PHASE3;
        step_odiv4_2 = STATIC_PHASE4;
        step_odiv0_3 = STATIC_PHASE0;
        step_odiv1_3 = STATIC_PHASE1;
        step_odiv2_3 = STATIC_PHASE2;
        step_odiv3_3 = STATIC_PHASE3;
        step_odiv4_3 = STATIC_PHASE4;
        step_odiv0_4 = STATIC_PHASE0;
        step_odiv1_4 = STATIC_PHASE1;
        step_odiv2_4 = STATIC_PHASE2;
        step_odiv3_4 = STATIC_PHASE3;
        step_odiv4_4 = STATIC_PHASE4;
        vco_fphase_delay0 = 0.0;
        vco_fphase_delay1 = 0.0;
        vco_fphase_delay2 = 0.0;
        vco_fphase_delay3 = 0.0;
        vco_fphase_delay4 = 0.0;
        cphase_delay0 = 0.0;
        cphase_delay1 = 0.0;
        cphase_delay2 = 0.0;
        cphase_delay3 = 0.0;
        cphase_delay4 = 0.0;
        odiv0_out_delay1 = 1'b0;
        odiv1_out_delay1 = 1'b0;
        odiv2_out_delay1 = 1'b0;
        odiv3_out_delay1 = 1'b0;
        odiv4_out_delay1 = 1'b0;
        odiv0_out_delay = 1'b0;
        odiv1_out_delay = 1'b0;
        odiv2_out_delay = 1'b0;
        odiv3_out_delay = 1'b0;
        odiv4_out_delay = 1'b0;
        clk_out0_gate = 3'b000;
        clk_out0_ext_gate = 3'b000;
        clk_out1_gate = 3'b000;
        clk_out2_gate = 3'b000;
        clk_out3_gate = 3'b000;
        clk_out4_gate = 3'b000;
        clk_out5_gate = 3'b000;
        clk_out5_reg  = 1'b0;
        inner_rstn = 1'b0;
        #1;
        inner_rstn = 1'b1;
        clk_in_first_time = 1'b1;
        clk_fb_first_time = 1'b1;
    end
///////////////////////////////////////////////////////
////RESET//////////////////////////////////////////////
    assign rst_n     = ~(PLL_PWD | RST) & inner_rstn;
    assign rstodiv_n = rst_n & (~RSTODIV);
///////////////////////////////////////////////////////
////INPUT_CLK_SEL//////////////////////////////////////
    assign clk_sel = (CLKIN_SEL_EN == 1'b0) ? dynauto_clkin : CLKIN_SEL;
    assign clk_in  = (clk_sel == 1'b0) ? CLKIN1 : CLKIN2;

    assign clk0 = CLKIN1 & (~CLKIN_SEL_EN);
    assign clk1 = CLKIN2 & (~CLKIN_SEL_EN);

    assign rstclksw_n = ~PLL_PWD & (~CLKIN_SEL_EN) & (~(cnt0[0] & cnt1[0] & (cnt0[1] | cnt1[1]))) & (~((cnt0[1]^cnt0[0]) & (cnt1[1]^cnt1[0])));

    always @(posedge clk0 or negedge rstclksw_n)
    begin
        if(!rstclksw_n)
            cnt0 <= 2'b00;
        else
            cnt0 <= cnt0+1;
    end

    always @(posedge clk1 or negedge rstclksw_n)
    begin
        if(!rstclksw_n)
            cnt1 <= 2'b00;
        else
            cnt1 <= cnt1+1;
    end

    always @(*)
    begin
        if(cnt0 == 2'b11)
            dynauto_clkin <= 1'b0;
        else
            if(cnt1 == 2'b11)
                dynauto_clkin <= 1'b1;
            else
                dynauto_clkin <= dynauto_clkin;
    end

    assign CLKSWITCH_FLAG = dynauto_clkin;
///////////////////////////////////////////////////////
////FBCK_DELAY/////////////////////////////////////////
    always @(posedge clk_in or negedge rst_n)
    begin
        if(!rst_n)
        begin
            clk_in_first_time = 1'b1;
            clk_in_first_edge = 0.0;
        end
        else
        begin
            if(clk_in_first_time == 1'b1)
                clk_in_first_edge = $realtime;
            clk_in_first_time = 1'b0;
        end
    end

    always @(posedge CLKFB or negedge rst_n)
    begin
        if(!rst_n)
        begin
            clk_fb_first_time = 1'b1;
            clk_fb_first_edge = 0.0;
        end
        else
        begin
            if(clk_fb_first_time == 1'b1)
                clk_fb_first_edge = $realtime;
            clk_fb_first_time = 1'b0;
        end
    end
///////////////////////////////////////////////////////
////PFD_ENABLE/////////////////////////////////////////
    assign pfden = (PFDEN_EN == "TRUE") ? PFDEN : 1'b1;

    always # 0.5 clk_pfd = ~clk_pfd;

    always @(posedge clk_in or negedge rst_n)
    begin
        if(!rst_n)
            pfd_en_reg <= 2'b11;
        else
            pfd_en_reg <= {pfd_en_reg[0], pfden};
    end

    always @(posedge clk_pfd or negedge rst_n)
    begin
        if(!rst_n)
        begin
            vcolow <= 0;
            cnt = 0;
        end
        else
            if(pfd_en_reg[1])
            begin
                vcolow <= 0;
                cnt = 0;
            end
            else
            begin
                cnt = cnt + 1;
                if(cnt == 500000)
                    vcolow <= 1;
            end
    end

    always #200 clk_test = ~clk_test;

    always @(posedge clk_test or negedge rst_n)
    begin
        if(!rst_n)
        begin
            clkwo <= 1'b0;
            clk_test_time1 = 0;
            clk_test_time2 = 0;
            clk_test_time3 = 0;

        end
        else
        begin
            clk_test_time3 = clk_test_time2;
            clk_test_time2 = clk_test_time1;
            clk_test_time1 = clkin_rtime_next;
            if(clk_test_time3 == clk_test_time1)
                clkwo <= 1'b1;
            else
                clkwo <= 1'b0;
        end
    end
///////////////////////////////////////////////////////
////PLL_ANALOG/////////////////////////////////////////
////FEEDBACK_DIVIDER_CAL///////////////////////////////
    assign idivider = (DYNAMIC_RATIOI_EN == "TRUE") ? RATIOI : STATIC_RATIOI;
    assign divider0 = (DYNAMIC_RATIO0_EN == "TRUE") ? RATIO0 : STATIC_RATIO0;
    assign divider1 = (DYNAMIC_RATIO1_EN == "TRUE") ? RATIO1 : STATIC_RATIO1;
    assign divider2 = (DYNAMIC_RATIO2_EN == "TRUE") ? RATIO2 : STATIC_RATIO2;
    assign divider3 = (DYNAMIC_RATIO3_EN == "TRUE") ? RATIO3 : STATIC_RATIO3;
    assign divider4 = (DYNAMIC_RATIO4_EN == "TRUE") ? RATIO4 : STATIC_RATIO4;
    assign fdivider = (DYNAMIC_RATIOF_EN == "TRUE") ? RATIOF : STATIC_RATIOF;
    assign mdivider = (DYNAMIC_RATIOM_EN == "TRUE") ? RATIOM : STATIC_RATIOM;

    always @(*)
    begin
        if(INTERNAL_FB == "ENABLE")
        begin
            fsdiv_set_int = fdivider;
            fbdiv_sel = 6'b000001;
        end
        else
            case(EXTERNAL_FB)
                "CLKOUT0": begin
                             fsdiv_set_int = divider0;
                             fbdiv_sel = 6'b000010;
                         end
                "CLKOUT1": begin
                             fsdiv_set_int = divider1;
                             fbdiv_sel = 6'b000100;
                         end
                "CLKOUT2": begin
                             fsdiv_set_int = divider2;
                             fbdiv_sel = 6'b001000;
                         end
                "CLKOUT3": begin
                             fsdiv_set_int = divider3;
                             fbdiv_sel = 6'b010000;
                         end
                "CLKOUT4": begin
                             fsdiv_set_int = divider4;
                             fbdiv_sel = 6'b100000;
                         end
            endcase
    end

    always @(*)
    begin
        if(VCOCLK_DIV2 == 1'b1)
        begin
            fbdiv_set_int = mdivider * fsdiv_set_int * 2;
            prop = 2;
        end
        else
        begin
            fbdiv_set_int = mdivider * fsdiv_set_int;
            prop = 1;
        end
    end
////PLL_VCO_CAL////////////////////////////////////////
    assign rstanalog_n = rst_n & ~vcolow;

    always @(posedge clk_in or negedge rstanalog_n)
    begin
        if(!rstanalog_n)
        begin
            clkin_rtime_last = 0.0;
            clkin_rtime_next = 0.0;
            clkin_time  <= 0.0;
            clkin_time1 <= 0.0;
            clkin_time2 <= 0.0;
            clkin_time3 <= 0.0;
            clkout_lock <= 0.0;
            vcoclk_period <= 1'b0;
            vcoclk_period_half <= 0.0;
            clkout0_time       <= 0.0;
            clkout1_time       <= 0.0;
            clkout2_time       <= 0.0;
            clkout3_time       <= 0.0;
            clkout4_time       <= 0.0;
            vcoclk_period_amp  <= 0.0;
            vcoclk_period_real <= 0.0;
            vcoclk_period_dev  <= 0.0;
        end
        else
        begin
            clkin_rtime_last = clkin_rtime_next;
            clkin_rtime_next = $realtime;
            if(clkin_rtime_last > 0)
            begin
                clkin_time  <= clkin_rtime_next-clkin_rtime_last;
                clkin_time1 <= clkin_time;
                clkin_time2 <= clkin_time1;
                clkin_time3 <= clkin_time2;
            end
            if(clkin_time > 0)
            begin
                clkout_lock <= (clkin_time  > 0) &&
                               (clkin_time1 > 0) &&
                               (clkin_time2 > 0) &&
                               (clkin_time3 > 0) &&
                               ((clkin_time - clkin_time1)  < 0.0001) &&
                               ((clkin_time1 - clkin_time)  < 0.0001) &&
                               ((clkin_time1 - clkin_time2) < 0.0001) &&
                               ((clkin_time2 - clkin_time1) < 0.0001) &&
                               ((clkin_time2 - clkin_time3) < 0.0001) &&
                               ((clkin_time3 - clkin_time2) < 0.0001);
            end
            if(clkin_time > 0)
            begin
                vcoclk_period      = (clkin_time * idivider) / fbdiv_set_int;
                vcoclk_period_half = vcoclk_period / 2;
                clkout0_time       = vcoclk_period * divider0 * prop;
                clkout1_time       = vcoclk_period * divider1 * prop;
                clkout2_time       = vcoclk_period * divider2 * prop;
                clkout3_time       = vcoclk_period * divider3 * prop;
                clkout4_time       = vcoclk_period * divider4 * prop;
                vcoclk_period_amp  = vcoclk_period_half * 100000;
                vcoclk_period_real = vcoclk_period_amp / 100000.0;
                vcoclk_period_dev  = (clkin_time - (vcoclk_period_real * 2 * fbdiv_set_int) / idivider) / 2;
            end
        end
    end

    always @(*)
    begin
        if(!rst_n)
        begin
            done = 1'b0;
            idiv_set = 0;
            fdiv_set = 0;
            swap_set = 0;
            fdiv_int = 0;
            offset = 0;
        end
        else
        begin
            idiv_set = idivider;
            fdiv_set = fbdiv_set_int;
            while(!done)
            begin
                if(idiv_set < fdiv_set)
                begin
                    swap_set = idiv_set;
                    idiv_set = fdiv_set;
                    fdiv_set = swap_set;
                end
                else
                    if(fdiv_set != 0)
                        idiv_set = idiv_set - fdiv_set;
                    else
                        done = 1;
            end
            fdiv_int = idiv_set;
            offset = vcoclk_period_dev * idivider/fdiv_int;
        end
    end

    always @(clkout_lock or inner_clk or clkwo)
    begin
        if(clkout_lock == 1'b0 || clkwo == 1'b1)
        begin
            inner_clk <= 1'b0;
            clk_gate  <= 1'b1;
            cnt_fdiv   = 0;
        end
        else
            if(clk_gate == 1)
            begin
                inner_clk <= 1'b1;
                clk_gate  <= 1'b0;
                cnt_fdiv   = 0;
            end
            else
            begin
                cnt_fdiv = cnt_fdiv + 1;
                if(cnt_fdiv == fbdiv_set_int/fdiv_int)
                begin
                    inner_clk <= #(vcoclk_period_half + offset) ~inner_clk;
                    cnt_fdiv = 0;
                end
                else
                    inner_clk <= #vcoclk_period_half ~inner_clk;
            end
    end

    always @(clk_in or CLKFB or negedge rst_n)
    begin
        if(!rst_n)
        begin
            adjust <= 1'b1;
            fb_route_delay = 0.0;
            tmp_ratio  = 0;
            tmp_delay  = 0.0;
            real_delay = 0.0;
        end
        else
            if(adjust == 1'b1)
            begin
                fb_route_delay = clk_fb_first_edge - clk_in_first_edge;
                if((clkin_time > 0) && (fb_route_delay > 0))
                begin
                    tmp_ratio  = fb_route_delay / clkin_time;
                    tmp_delay  = fb_route_delay - (clkin_time * tmp_ratio);
                    real_delay = clkin_time - tmp_delay;
                    adjust <= 1'b0;
                end
            end
    end

    always @(inner_clk)
    begin
        if(EXTERNAL_FB == "CLKOUT0" || EXTERNAL_FB == "CLKOUT1" || EXTERNAL_FB == "CLKOUT2" || EXTERNAL_FB == "CLKOUT3" || EXTERNAL_FB == "CLKOUT4")
            vcoclk <= #real_delay inner_clk;
        else
            vcoclk <= inner_clk;
    end
////VCO_CLK_DIV2///////////////////////////////////////
    always @(posedge vcoclk or negedge rst_n)
    begin
        if(!rst_n)
            clk_vcodiv2 <= 1'b0;
        else
            if(VCOCLK_DIV2)
                clk_vcodiv2 <= ~clk_vcodiv2;
            else
                clk_vcodiv2 <= 1'b0;
    end

    assign clkout = (VCOCLK_DIV2 == 1'b0) ? vcoclk : clk_vcodiv2;
///////////////////////////////////////////////////////
////PLL_LOCK///////////////////////////////////////////
    assign clk_lock = (INTERNAL_FB == "ENABLE") ? clk_in : CLKFB;

    always @(posedge clk_lock or negedge rstanalog_n)
    begin
        if(!rstanalog_n)
        begin
            start_clk <= 1'b0;
            cnt_clkfb <= 2'b00;
        end
        else
            if(cnt_clkfb == 3)
                start_clk = 1'b1;
            else
                cnt_clkfb = cnt_clkfb + 1;
    end

    always @(posedge clk_in or negedge rstanalog_n or clk_gate)
    begin
        if(!rstanalog_n)
        begin
            cnt_lock <= 11'b000_0000_0001;
            lock_reg <= 1'b0;
        end
        else
            if(!clk_gate && start_clk)
                if(cnt_lock == idivider * 3)
                    lock_reg <= 1'b1;
                else
                    cnt_lock <= cnt_lock+1;
            else
            begin
                cnt_lock <= 11'b000_0000_0001;
                lock_reg <= 1'b0;
            end
    end

    assign LOCK = lock_reg;
///////////////////////////////////////////////////////
////PLL_ODIV///////////////////////////////////////////
////ODIV0//////////////////////////////////////////////
    assign clk_sel0   = clkout;
    assign odiv0_rstn = rst_n & (fbdiv_sel[1] | rstodiv_n);

    assign odiv0_duty      = (DYNAMIC_DUTY0_EN  == "TRUE") ? DUTY0 : STATIC_DUTY0;
    assign odiv0_duty_ctrl = (odiv0_duty[0] == 1'b1) ? (odiv0_duty+1'b1) >> 1 : odiv0_duty >> 1;

    always @(negedge clk_sel0 or negedge odiv0_rstn)
    begin
        if(!odiv0_rstn)
            enclk0 <= 3'b000;
        else
            enclk0 <= {enclk0[1:0],1'b1};
    end

    assign clk_en0 = clk_sel0 & enclk0[2];

    always @(posedge clk_en0 or negedge odiv0_rstn)
    begin
        if(!odiv0_rstn)
            odiv0_counter <= 10'b00_0000_0000;
        else
            if(odiv0_counter == divider0 - 1'b1)
                odiv0_counter <= 10'b00_0000_0000;
            else
                odiv0_counter <= odiv0_counter + 1'b1;
    end

    always @(posedge clk_en0 or negedge odiv0_rstn)
    begin
        if(!odiv0_rstn)
            odiv0_clkdivr <= 1'b0;
        else
            if(odiv0_counter < odiv0_duty_ctrl)
                odiv0_clkdivr <= 1'b1;
            else
                odiv0_clkdivr <= 1'b0;
    end

    always @(negedge clk_en0 or negedge odiv0_rstn)
    begin
        if(!odiv0_rstn)
            odiv0_set <= 1'b0;
        else
            if(odiv0_counter == odiv0_duty_ctrl)
                odiv0_set <= odiv0_duty[0];
            else
                odiv0_set <= 1'b0;
    end

    assign odiv0_out = (divider0 == 10'b00_0000_0001) ? clk_en0 & enclk0[2] : odiv0_clkdivr & (~odiv0_set);
////ODIV1//////////////////////////////////////////////
    assign clk_sel1   = (CLK_CAS1_EN == "TRUE") ? odiv0_out : clkout;
    assign odiv1_rstn = rst_n & (fbdiv_sel[2] | rstodiv_n);

    assign odiv1_duty      = (DYNAMIC_DUTY1_EN  == "TRUE") ? DUTY1 : STATIC_DUTY1;
    assign odiv1_duty_ctrl = (odiv1_duty[0] == 1'b1) ? (odiv1_duty+1'b1) >> 1 : odiv1_duty >> 1;

    always @(negedge clk_sel1 or negedge odiv1_rstn)
    begin
        if(!odiv1_rstn)
            enclk1 <= 3'b000;
        else
            enclk1 <= {enclk1[1:0],1'b1};
    end

    assign clk_en1 = clk_sel1 & enclk1[2];

    always @(posedge clk_en1 or negedge odiv1_rstn)
    begin
        if(!odiv1_rstn)
            odiv1_counter <= 10'b00_0000_0000;
        else
            if(odiv1_counter == divider1 - 1'b1)
                odiv1_counter <= 10'b00_0000_0000;
            else
                odiv1_counter <= odiv1_counter + 1'b1;
    end

    always @(posedge clk_en1 or negedge odiv1_rstn)
    begin
        if(!odiv1_rstn)
            odiv1_clkdivr <= 1'b0;
        else
            if(odiv1_counter < odiv1_duty_ctrl)
                odiv1_clkdivr <= 1'b1;
            else
                odiv1_clkdivr <= 1'b0;
    end

    always @(negedge clk_en1 or negedge odiv1_rstn)
    begin
        if(!odiv1_rstn)
            odiv1_set <= 1'b0;
        else
            if(odiv1_counter == odiv1_duty_ctrl)
                odiv1_set <= odiv1_duty[0];
            else
                odiv1_set <= 1'b0;
    end

    assign odiv1_out = (divider1 == 10'b00_0000_0001) ? clk_en1 & enclk1[2] : odiv1_clkdivr & (~odiv1_set);
////ODIV2//////////////////////////////////////////////
    assign clk_sel2   = (CLK_CAS2_EN == "TRUE") ? odiv1_out : clkout;
    assign odiv2_rstn = rst_n & (fbdiv_sel[3] | rstodiv_n);

    assign odiv2_duty      = (DYNAMIC_DUTY2_EN  == "TRUE") ? DUTY2 : STATIC_DUTY2;
    assign odiv2_duty_ctrl = (odiv2_duty[0] == 1'b1) ? (odiv2_duty+1'b1) >> 1 : odiv2_duty >> 1;

    always @(negedge clk_sel2 or negedge odiv2_rstn)
    begin
        if(!odiv2_rstn)
            enclk2 <= 3'b000;
        else
            enclk2 <= {enclk2[1:0],1'b1};
    end

    assign clk_en2 = clk_sel2 & enclk2[2];

    always @(posedge clk_en2 or negedge odiv2_rstn)
    begin
        if(!odiv2_rstn)
            odiv2_counter <= 10'b00_0000_0000;
        else
            if(odiv2_counter == divider2 - 1'b1)
                odiv2_counter <= 10'b00_0000_0000;
            else
                odiv2_counter <= odiv2_counter + 1'b1;
    end

    always @(posedge clk_en2 or negedge odiv2_rstn)
    begin
        if(!odiv2_rstn)
            odiv2_clkdivr <= 1'b0;
        else
            if(odiv2_counter < odiv2_duty_ctrl)
                odiv2_clkdivr <= 1'b1;
            else
                odiv2_clkdivr <= 1'b0;
    end

    always @(negedge clk_en2 or negedge odiv2_rstn)
    begin
        if(!odiv2_rstn)
            odiv2_set <= 1'b0;
        else
            if(odiv2_counter == odiv2_duty_ctrl)
                odiv2_set <= odiv2_duty[0];
            else
                odiv2_set <= 1'b0;
    end

    assign odiv2_out = (divider2 == 10'b00_0000_0001) ? clk_en2 & enclk2[2] : odiv2_clkdivr & (~odiv2_set);
////ODIV3//////////////////////////////////////////////
    assign clk_sel3   = (CLK_CAS3_EN == "TRUE") ? odiv2_out : clkout;
    assign odiv3_rstn = rst_n & (fbdiv_sel[4] | rstodiv_n);

    assign odiv3_duty      = (DYNAMIC_DUTY3_EN  == "TRUE") ? DUTY3 : STATIC_DUTY3;
    assign odiv3_duty_ctrl = (odiv3_duty[0] == 1'b1) ? (odiv3_duty+1'b1) >> 1 : odiv3_duty >> 1;

    always @(negedge clk_sel3 or negedge odiv3_rstn)
    begin
        if(!odiv3_rstn)
            enclk3 <= 3'b000;
        else
            enclk3 <= {enclk3[1:0],1'b1};
    end

    assign clk_en3 = clk_sel3 & enclk3[2];

    always @(posedge clk_en3 or negedge odiv3_rstn)
    begin
        if(!odiv3_rstn)
            odiv3_counter <= 10'b00_0000_0000;
        else
            if(odiv3_counter == divider3 - 1'b1)
                odiv3_counter <= 10'b00_0000_0000;
            else
                odiv3_counter <= odiv3_counter + 1'b1;
    end

    always @(posedge clk_en3 or negedge odiv3_rstn)
    begin
        if(!odiv3_rstn)
            odiv3_clkdivr <= 1'b0;
        else
            if(odiv3_counter < odiv3_duty_ctrl)
                odiv3_clkdivr <= 1'b1;
            else
                odiv3_clkdivr <= 1'b0;
    end

    always @(negedge clk_en3 or negedge odiv3_rstn)
    begin
        if(!odiv3_rstn)
            odiv3_set <= 1'b0;
        else
            if(odiv3_counter == odiv3_duty_ctrl)
                odiv3_set <= odiv3_duty[0];
            else
                odiv3_set <= 1'b0;
    end

    assign odiv3_out = (divider3 == 10'b00_0000_0001) ? clk_en3 & enclk3[2] : odiv3_clkdivr & (~odiv3_set);
////ODIV4//////////////////////////////////////////////
    assign clk_sel4   = (CLK_CAS4_EN == "TRUE") ? odiv3_out : clkout;
    assign odiv4_rstn = rst_n & (fbdiv_sel[5] | rstodiv_n);

    assign odiv4_duty      = (DYNAMIC_DUTY4_EN  == "TRUE") ? DUTY4 : STATIC_DUTY4;
    assign odiv4_duty_ctrl = (odiv4_duty[0] == 1'b1) ? (odiv4_duty+1'b1) >> 1 : odiv4_duty >> 1;

    always @(negedge clk_sel4 or negedge odiv4_rstn)
    begin
        if(!odiv4_rstn)
            enclk4 <= 3'b000;
        else
            enclk4 <= {enclk4[1:0],1'b1};
    end

    assign clk_en4 = clk_sel4 & enclk4[2];

    always @(posedge clk_en4 or negedge odiv4_rstn)
    begin
        if(!odiv4_rstn)
            odiv4_counter <= 10'b00_0000_0000;
        else
            if(odiv4_counter == divider4 - 1'b1)
                odiv4_counter <= 10'b00_0000_0000;
            else
                odiv4_counter <= odiv4_counter + 1'b1;
    end

    always @(posedge clk_en4 or negedge odiv4_rstn)
    begin
        if(!odiv4_rstn)
            odiv4_clkdivr <= 1'b0;
        else
            if(odiv4_counter < odiv4_duty_ctrl)
                odiv4_clkdivr <= 1'b1;
            else
                odiv4_clkdivr <= 1'b0;
    end

    always @(negedge clk_en4 or negedge odiv4_rstn)
    begin
        if(!odiv4_rstn)
            odiv4_set <= 1'b0;
        else
            if(odiv4_counter == odiv4_duty_ctrl)
                odiv4_set <= odiv4_duty[0];
            else
                odiv4_set <= 1'b0;
    end

    assign odiv4_out = (divider4 == 10'b00_0000_0001) ? clk_en4 & enclk4[2] : odiv4_clkdivr & (~odiv4_set);
///////////////////////////////////////////////////////
////PHASE_SHIFT////////////////////////////////////////
    always @(*)
    begin
        fphase_step = PHASE_STEP_N;
    end

    always @(fphase_step)
    begin
        last_fphase_step <= fphase_step;
    end

    always @(*)
    begin
        if(LOAD_PHASE == 1'b1)
        begin
            step_odiv0 = step_odiv0_1;
            step_odiv1 = step_odiv1_1;
            step_odiv2 = step_odiv2_1;
            step_odiv3 = step_odiv3_1;
            step_odiv4 = step_odiv4_1;
        end
        else
            if(PHASE_SEL == 3'b000)
            begin
                if(fphase_step === 1'b0 && last_fphase_step === 1'b1)
                    if(PHASE_DIR == 1'b0)
                        step_odiv0 <= step_odiv0 + 1;
                    else
                        step_odiv0 <= step_odiv0 - 1;
            end
            else if(PHASE_SEL == 3'b001)
            begin
                if(fphase_step === 1'b0 && last_fphase_step === 1'b1)
                    if(PHASE_DIR == 1'b0)
                        step_odiv1 <= step_odiv1 + 1;
                    else
                        step_odiv1 <= step_odiv1 - 1;
            end
            else if(PHASE_SEL == 3'b010)
            begin
                if(fphase_step === 1'b0 && last_fphase_step === 1'b1)
                    if(PHASE_DIR == 1'b0)
                        step_odiv2 <= step_odiv2 + 1;
                    else
                        step_odiv2 <= step_odiv2 - 1;
            end
            else if(PHASE_SEL == 3'b011)
            begin
                if(fphase_step === 1'b0 && last_fphase_step === 1'b1)
                    if(PHASE_DIR == 1'b0)
                        step_odiv3 <= step_odiv3 + 1;
                    else
                        step_odiv3 <= step_odiv3 - 1;
            end
            else if(PHASE_SEL == 3'b100)
            begin
                if(fphase_step === 1'b0 && last_fphase_step === 1'b1)
                    if(PHASE_DIR == 1'b0)
                        step_odiv4 <= step_odiv4 + 1;
                    else
                        step_odiv4 <= step_odiv4 - 1;
            end
    end

    always @(posedge last_fphase_step or negedge rst_n)
    begin
        if(!rst_n)
        begin
            step_odiv0_1 <= STATIC_PHASE0;
            step_odiv1_1 <= STATIC_PHASE1;
            step_odiv2_1 <= STATIC_PHASE2;
            step_odiv3_1 <= STATIC_PHASE3;
            step_odiv4_1 <= STATIC_PHASE4;
        end
        else
        begin
            step_odiv0_1 <= step_odiv0;
            step_odiv1_1 <= step_odiv1;
            step_odiv2_1 <= step_odiv2;
            step_odiv3_1 <= step_odiv3;
            step_odiv4_1 <= step_odiv4;
        end
    end

    always @(posedge inner_clk)
    begin
        step_odiv0_2 <= step_odiv0_1;
        step_odiv0_3 <= step_odiv0_2;
        step_odiv1_2 <= step_odiv1_1;
        step_odiv1_3 <= step_odiv1_2;
        step_odiv2_2 <= step_odiv2_1;
        step_odiv2_3 <= step_odiv2_2;
        step_odiv3_2 <= step_odiv3_1;
        step_odiv3_3 <= step_odiv3_2;
        step_odiv4_2 <= step_odiv4_1;
        step_odiv4_3 <= step_odiv4_2;
    end

    always @(negedge inner_clk)
    begin
        step_odiv0_4 <= step_odiv0_3;
        step_odiv1_4 <= step_odiv1_3;
        step_odiv2_4 <= step_odiv2_3;
        step_odiv3_4 <= step_odiv3_3;
        step_odiv4_4 <= step_odiv4_3;
    end
////PHASE_SHIFT_CAL////////////////////////////////////
    always @(*)
    begin
        if(step_odiv0_4 >= 0)
            step_odiv0_5 <= step_odiv0_4;
        else
            step_odiv0_5 <= step_odiv0_4 + (~step_odiv0_4/(8*divider0))*8*divider0;

        if(step_odiv1_4 >= 0)
            step_odiv1_5 <= step_odiv1_4;
        else
            step_odiv1_5 <= step_odiv1_4 + (~step_odiv1_4/(8*divider1))*8*divider1;

        if(step_odiv2_4 >= 0)
            step_odiv2_5 <= step_odiv2_4;
        else
            step_odiv2_5 <= step_odiv2_4 + (~step_odiv2_4/(8*divider2))*8*divider2;

        if(step_odiv3_4 >= 0)
            step_odiv3_5 <= step_odiv3_4;
        else
            step_odiv3_5 <= step_odiv3_4 + (~step_odiv3_4/(8*divider3))*8*divider3;

        if(step_odiv4_4 >= 0)
            step_odiv4_5 <= step_odiv4_4;
        else
            step_odiv4_5 <= step_odiv4_4 + (~step_odiv4_4/(8*divider4))*8*divider4;
    end

    always @(*)
    begin
        if(clkout0_time > 0)
            if(step_odiv0_5 >= 0)
                vco_fphase_delay0 <= (step_odiv0_5 * clkout0_time) / (8 * prop * divider0);
            else
                vco_fphase_delay0 <= clkout0_time + (step_odiv0_5 * clkout0_time) / (8 * prop * divider0);

        if(clkout1_time > 0)
            if(step_odiv1_5 >= 0)
                vco_fphase_delay1 <= (step_odiv1_5 * clkout1_time) / (8 * prop * divider1);
            else
                vco_fphase_delay1 <= clkout1_time + (step_odiv1_5 * clkout1_time) / (8 * prop * divider1);

        if(clkout2_time > 0)
            if(step_odiv2_5 >= 0)
                vco_fphase_delay2 <= (step_odiv2_5 * clkout2_time) / (8 * prop * divider2);
            else
                vco_fphase_delay2 <= clkout2_time + (step_odiv2_5 * clkout2_time) / (8 * prop * divider2);

        if(clkout3_time > 0)
            if(step_odiv3_5 >= 0)
                vco_fphase_delay3 <= (step_odiv3_5 * clkout3_time) / (8 * prop * divider3);
            else
                vco_fphase_delay3 <= clkout3_time + (step_odiv3_5 * clkout3_time) / (8 * prop * divider3);

        if(clkout4_time > 0)
            if(step_odiv4_5 >= 0)
                vco_fphase_delay4 <= (step_odiv4_5 * clkout4_time) / (8 * prop * divider4);
            else
                vco_fphase_delay4 <= clkout4_time + (step_odiv4_5 * clkout4_time) / (8 * prop * divider4);
    end

    always @(*)
    begin
        if(divider0 > STATIC_CPHASE0)
            phase0 = STATIC_CPHASE0;
        else
            phase0 = STATIC_CPHASE0 - (STATIC_CPHASE0/divider0)*divider0;

        if(divider1 > STATIC_CPHASE1)
            phase1 = STATIC_CPHASE1;
        else
            phase1 = STATIC_CPHASE1 - (STATIC_CPHASE1/divider1)*divider1;

        if(divider2 > STATIC_CPHASE2)
            phase2 = STATIC_CPHASE2;
        else
            phase2 = STATIC_CPHASE2 - (STATIC_CPHASE2/divider2)*divider2;

        if(divider3 > STATIC_CPHASE3)
            phase3 = STATIC_CPHASE3;
        else
            phase3 = STATIC_CPHASE3 - (STATIC_CPHASE3/divider3)*divider3;

        if(divider4 > STATIC_CPHASE4)
            phase4 = STATIC_CPHASE4;
        else
            phase4 = STATIC_CPHASE4 - (STATIC_CPHASE4/divider4)*divider4;
    end

    always @(*)
    begin
        if(clkout0_time > 0)
            cphase_delay0 <= clkout0_time - (((divider0 - phase0) * clkout0_time) / divider0);
        else
            cphase_delay0 <= 0.0;

        if(clkout1_time > 0)
            cphase_delay1 <= clkout1_time - (((divider1 - phase1) * clkout1_time) / divider1);
        else
            cphase_delay1 <= 0.0;

        if(clkout2_time > 0)
            cphase_delay2 <= clkout2_time - (((divider2 - phase2) * clkout2_time) / divider2);
        else
            cphase_delay2 <= 0.0;

        if(clkout3_time > 0)
            cphase_delay3 <= clkout3_time - (((divider3 - phase3) * clkout3_time) / divider3);
        else
            cphase_delay3 <= 0.0;

        if(clkout4_time > 0)
            cphase_delay4 <= clkout4_time - (((divider4 - phase4) * clkout4_time) / divider4);
        else
            cphase_delay4 <= 0.0;
    end
////PHASE_SHIFT_DLY////////////////////////////////////
    always @(odiv0_out)
    begin
        odiv0_out_delay1 <= #vco_fphase_delay0 odiv0_out;
    end

    always @(odiv0_out_delay1)
    begin
        odiv0_out_delay <= #cphase_delay0 odiv0_out_delay1;
    end

    always @(odiv1_out)
    begin
        odiv1_out_delay1 <= #vco_fphase_delay1 odiv1_out;
    end

    always @(odiv1_out_delay1)
    begin
        odiv1_out_delay <= #cphase_delay1 odiv1_out_delay1;
    end

    always @(odiv2_out)
    begin
        odiv2_out_delay1 <= #vco_fphase_delay2 odiv2_out;
    end

    always @(odiv2_out_delay1)
    begin
        odiv2_out_delay <= #cphase_delay2 odiv2_out_delay1;
    end

    always @(odiv3_out)
    begin
        odiv3_out_delay1 <= #vco_fphase_delay3 odiv3_out;
    end

    always @(odiv3_out_delay1)
    begin
        odiv3_out_delay <= #cphase_delay3 odiv3_out_delay1;
    end

    always @(odiv4_out)
    begin
        odiv4_out_delay1 <= #vco_fphase_delay4 odiv4_out;
    end

    always @(odiv4_out_delay1)
    begin
        odiv4_out_delay <= #cphase_delay4 odiv4_out_delay1;
    end
///////////////////////////////////////////////////////
////PLL_GATE///////////////////////////////////////////
    always @(negedge odiv0_out_delay or negedge inner_rstn)
    begin
        if(!inner_rstn)
            clk_out0_gate <= 3'b000;
        else
            clk_out0_gate <= {clk_out0_gate[1:0],~CLKOUT0_SYN};
    end

    assign clkout0_gate = (CLKOUT0_SYN_EN == "TRUE") ? clk_out0_gate[2] : 1'b1;
    assign CLKOUT0      = odiv0_out_delay & clkout0_gate;

    always @(negedge odiv0_out_delay or negedge inner_rstn)
    begin
        if(!inner_rstn)
            clk_out0_ext_gate <= 3'b000;
        else
            clk_out0_ext_gate <= {clk_out0_ext_gate[1:0],~CLKOUT0_EXT_SYN};
    end

    assign clkout0_ext_gate = (CLKOUT0_EXT_SYN_EN == "TRUE") ? clk_out0_ext_gate[2] : 1'b1;
    assign CLKOUT0_EXT      = odiv0_out_delay & clkout0_ext_gate;

    always @(negedge odiv1_out_delay or negedge inner_rstn)
    begin
        if(!inner_rstn)
            clk_out1_gate <= 3'b000;
        else
            clk_out1_gate <= {clk_out1_gate[1:0],~CLKOUT1_SYN};
    end

    assign clkout1_gate = (CLKOUT1_SYN_EN == "TRUE") ? clk_out1_gate[2] : 1'b1;
    assign CLKOUT1      = odiv1_out_delay & clkout1_gate;

    always @(negedge odiv2_out_delay or negedge inner_rstn)
    begin
        if(!inner_rstn)
            clk_out2_gate <= 3'b000;
        else
            clk_out2_gate <= {clk_out2_gate[1:0],~CLKOUT2_SYN};
    end

    assign clkout2_gate = (CLKOUT2_SYN_EN == "TRUE") ? clk_out2_gate[2] : 1'b1;
    assign CLKOUT2      = odiv2_out_delay & clkout2_gate;

    always @(negedge odiv3_out_delay or negedge inner_rstn)
    begin
        if(!inner_rstn)
            clk_out3_gate <= 3'b000;
        else
            clk_out3_gate <= {clk_out3_gate[1:0],~CLKOUT3_SYN};
    end

    assign clkout3_gate = (CLKOUT3_SYN_EN == "TRUE") ? clk_out3_gate[2] : 1'b1;
    assign CLKOUT3      = odiv3_out_delay & clkout3_gate;

    assign clkout4_sel = (CLKIN_BYPASS_EN == "TRUE") ? clk_in : odiv4_out_delay;

    always @(negedge clkout4_sel or negedge inner_rstn)
    begin
        if(!inner_rstn)
            clk_out4_gate <= 3'b000;
        else
            clk_out4_gate <= {clk_out4_gate[1:0],~CLKOUT4_SYN};
    end

    assign clkout4_gate = (CLKOUT4_SYN_EN == "TRUE") ? clk_out4_gate[2] : 1'b1;
    assign CLKOUT4      = clkout4_sel & clkout4_gate;

    always @(*)
    begin
        case(CLKOUT5_SEL)
            0: clk_out5_reg = odiv0_out_delay;
            1: clk_out5_reg = odiv1_out_delay;
            2: clk_out5_reg = odiv2_out_delay;
            3: clk_out5_reg = odiv3_out_delay;
            4: clk_out5_reg = odiv4_out_delay;
            default: clk_out5_reg = odiv0_out_delay;
        endcase
    end

    assign clkout5_synen = (CLKOUT5_SYN_EN == "TRUE") ? 1'b1 : 1'b0;

    always @(negedge clk_out5_reg or negedge inner_rstn)
    begin
        if(!inner_rstn)
            clk_out5_gate <= 3'b000;
        else
            clk_out5_gate <= {clk_out5_gate[1:0],~CLKOUT5_SYN};
    end

    assign clkout5_gate = (CLKOUT5_SYN_EN == "TRUE") ? clk_out5_gate[2] : 1'b1;
    assign CLKOUT5      = clk_out5_reg & clkout5_gate;
endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_RAM16X1SP.v
//
// Functional description: single-port 16x1 distributed ram
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_RAM16X1SP
#(
    parameter [15:0] INIT = 16'h0000
) (
    output  DO,
    input   DI,
    input [3:0] ADDR,
    input WCLK, WE
);

    reg [15:0] mem ;

    initial begin
        mem = INIT;
    end

    always @(posedge WCLK) begin
        if (WE == 1'b1) begin
            mem[ADDR] <= DI;
        end
    end

    assign DO = mem[ADDR];

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_ISERDES.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//2017/12/20 : initial version
//2018/01/02 : change DELAY_STEP to DELAY_STEP_VALUE;
//             change DYN_CTRL_EN to DELAY_STEP_SEL;
//             change DELAY_CTRL to DELAY_STEP;
//2018/03/20 : fix bug XA-30
//2018/04/13 : delete parameter DELAY_EN
/////////////////////////////////////////////////////////////////////////////
`timescale 1 ns / 1 ps

module GTP_IODELAY_E1 #(
parameter [4:0] DELAY_STEP_VALUE = 5'h00, //5'h00 ~ 5'h1F
parameter DELAY_STEP_SEL   = "PARAMETER"   //"PARAMETER", "PORT"
)(
output      DO,
input       DI,
input [4:0] DELAY_STEP
); /* synthesis syn_black_box */ 

//synthesis translate_off
///////////////////////////////////////////////////////////////////////////

initial 
begin
    if(DELAY_STEP_SEL != "PARAMETER" && DELAY_STEP_SEL != "PORT")
    begin
      $display("GTP_IODELAY_E1 Error: Illegal setting of DELAY_STEP_SEL %s",DELAY_STEP_SEL);
      $finish;
    end

    if(DELAY_STEP_VALUE > 5'd31 || DELAY_STEP_VALUE < 0)
    begin
      $display("GTP_IODELAY_E1 Error: Illegal setting of DELAY_STEP_VALUE %s",DELAY_STEP_VALUE);
      $finish;
    end
end

wire [4:0] ioldly_step;
assign ioldly_step = (DELAY_STEP_SEL == "PORT") ? DELAY_STEP : DELAY_STEP_VALUE;

wire [31:0] ioldly;
assign ioldly[0] = DI;

genvar i;
generate
    for(i=1;i<4;i=i+1)begin
      assign #0.22 ioldly[i] = ioldly[i-1];
    end
endgenerate

assign #0.22 ioldly[4]  = (ioldly_step[4]||ioldly_step[3]) ? ioldly[3]  : 1'b0;
genvar j;
generate
    for(j=5;j<8;j=j+1)begin
      assign #0.22 ioldly[j] = ioldly[j-1];
    end
endgenerate

assign #0.22 ioldly[8] = ioldly_step[4] ? ioldly[7] : 1'b0;
genvar k;
generate
    for(k=9;k<12;k=k+1)begin
      assign #0.22 ioldly[k] = ioldly[k-1];
    end
endgenerate

assign #0.22 ioldly[12] = (ioldly_step[4]&&ioldly_step[3]) ? ioldly[11] : 1'b0;
genvar l;
generate
    for(l=13;l<16;l=l+1)begin
      assign #0.22 ioldly[l] = ioldly[l-1];
    end
endgenerate

wire ioldly_out_even;
wire ioldly_out_odd;

assign ioldly_out_even = ioldly[ioldly_step[4:1]];
assign #0.11 ioldly_out_odd  = ioldly_out_even;

wire ioldly_out;
assign ioldly_out = ioldly_step[0] ? ioldly_out_odd : ioldly_out_even;

assign DO = ioldly_out;

//synthesis translate_on

endmodule

























//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_OGSER8.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_OGSER8 #(
parameter GRS_EN = "TRUE", //"TRUE"; "FALSE" 
parameter LRS_EN = "TRUE"   //"TRUE"; "FALSE" 
)(
output  PADO,
output  PADT,
input [7:0] D,
input [3:0] T,
input RCLK,
input SERCLK,
input RST
);

//synthesis translate_off
reg [7:0] d_rclk;
reg [3:0] t_rclk;
reg [1:0] cnt;
reg [7:0] capture_d_reg;
reg [3:0] capture_t_reg;
reg [7:0] shift_d_reg;
reg [3:0] shift_t_reg;
wire capture_en;
reg PADO_POS;
reg PADT_reg;
reg PADO_NEG;

initial begin
d_rclk        = 0;
t_rclk        = 0;
cnt           = 0;
capture_d_reg = 0;
capture_t_reg = 0;
shift_d_reg   = 0;
shift_t_reg   = 0;
PADO_POS      = 0;
PADT_reg      = 0;
PADO_NEG      = 0;
end

assign global_rstn = (GRS_EN == "TRUE") ? GRS_INST.GRSNET : 1'b1;
assign lsr_rstn = LRS_EN == "TRUE" ? (~RST) : 1'b1;

always @(posedge RCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn) begin
      d_rclk <= 0;
      t_rclk <= 0;
   end
   else if (!lsr_rstn) begin
      d_rclk <= 0;
      t_rclk <= 0;
   end   
   else begin
      d_rclk <= D;
      t_rclk <= T;    
   end
   
always @(posedge SERCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      cnt <= 0;
   else if (!lsr_rstn)
      cnt <= 0;
   else
      cnt <= cnt + 1;

assign capture_en = cnt == 3;      
assign shift_en = cnt == 2;

always @(posedge SERCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn) begin
      capture_d_reg <= 0;
      capture_t_reg <= 0;
   end   
   else if (!lsr_rstn) begin
      capture_d_reg <= 0;
      capture_t_reg <= 0;
   end   
   else if (capture_en) begin
      capture_d_reg <= d_rclk;
      capture_t_reg <= t_rclk;
   end
   
always @(posedge SERCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn) begin
      shift_d_reg <= 0;
      shift_t_reg <= 0;
   end   
   else if (!lsr_rstn) begin
      shift_d_reg <= 0;
      capture_t_reg <= 0;
   end   
   else if (shift_en) begin
      shift_d_reg <= capture_d_reg;
      shift_t_reg <= capture_t_reg;
   end
   else begin
      shift_d_reg <= {2'd0, shift_d_reg[7:2]};
      shift_t_reg <= {1'b0, shift_t_reg[3:1]};    
   end      
   
always @(posedge SERCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn) begin
      PADO_POS <= 0;
      PADT_reg <= 0;
   end
   else if (!lsr_rstn) begin
      PADO_POS <= 0;
      PADT_reg <= 0;
   end
   else begin
      PADO_POS <= shift_d_reg[1];
      PADT_reg <= shift_t_reg[0];     
   end           
   
always @(negedge SERCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn) begin
      PADO_NEG <= 0;
   end
   else if (!lsr_rstn) begin
      PADO_NEG <= 0;
   end
   else begin
      PADO_NEG <= shift_d_reg[0];
   end           
   
assign PADO =  SERCLK ? PADO_NEG : PADO_POS;
assign PADT = PADT_reg;
   
//synthesis translate_on

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_FIR_B.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_FIR_B
#(
    parameter GRS_EN    = "TRUE", //"TRUE"; "FALSE"
    parameter SYNC_RST  = "FALSE", //"TRUE"; "FALSE"
    parameter INREG_EN  = "TRUE",
    parameter OUTREG_EN = "TRUE",
    parameter INPUT_OP    = 1'b1,
    parameter DYN_OP_SEL  = 1'b1,
    parameter OPCD_DYN_SEL = 1'b0,
    parameter OPCD_CPI_SEL = 1'b0
) (
    output  [26:0] CYO,
    output         CYO_SIGNED,
    output [63:0] CPO,                  //p
    output        CPO_SIGNED,
    output [63:0] P,

    input   CE,
    input   RST,
    input   CLK,
    input [26:0] CYI,
    input        CYI_SIGNED,
    input [26:0] Y0,                  //y0 ,DYIB,DYIA
    input        Y0_SIGNED,
    input [26:0] H0,                  //h0 ,DXIB,DXIA
    input        H0_SIGNED,
    input [63:0] CPI,
    input        CPI_SIGNED,
    input        S0,
    input        OPCD_CPI_DYN
);

//PSE parameter
localparam [25:0] SC_PSE_Y0 = 26'b0;  //SC_PSE = 0, disable PSE, parameter bit width=26
localparam [25:0] SC_PSE_H0 = 26'b0;  //SC_PSE = 0, disable PSE, parameter bit width=26

initial begin
    if ((GRS_EN != "TRUE") && (GRS_EN != "FALSE")) begin
        $display("GRS_EN error");
        $finish;
    end
    if ((SYNC_RST != "TRUE") && (SYNC_RST != "FALSE")) begin
        $display("SYNC_RST error");
        $finish;
    end
end

reg [26:0] h0_d;
reg        h0_signed_d;
reg [26:0] y0_d;
reg        y0_signed_d;

wire [26:0] y0_sel;
wire        y0_signed_sel;

wire        s0_d_sel, s0_sel;
wire [26:0] y0_d_sel;
wire        y0_signed_d_sel;
wire [26:0] h0_d_sel;
wire        h0_signed_d_sel;

wire INPUT_OP_CODE;

wire [53:0] mult1_in1;
wire [53:0] mult1_in2;

wire [53:0] mult1;
wire        mult1_signed;

wire [63:0] sum;
wire        sum_signed;
reg  [63:0] sum_d;
reg         sum_signed_d;

reg  [26:0] cyo_d;
reg         cyo_signed_d;
wire [26:0] cyo;
wire        cyo_signed;

wire global_rstn ;
wire RST_sync ;
wire RST_async;
wire rst_asyncomb ;

wire [26:0] Y0_PSE;
wire [26:0] H0_PSE;

wire [63:0] CPI_SEL;
wire        OPCD_SEL;

assign OPCD_SEL = (OPCD_DYN_SEL == 1'b1)?OPCD_CPI_DYN :OPCD_CPI_SEL;
assign CPI_SEL  = (OPCD_SEL == 1'b1)? 64'b0 : CPI;

assign global_rstn = GRS_EN == "TRUE" ? GRS_INST.GRSNET : 1'b1;
assign RST_sync = (SYNC_RST == "TRUE") ? RST : 1'b0;
assign RST_async = (SYNC_RST == "FALSE") ? RST : 1'b0;
assign rst_asyncomb = RST_async | (~global_rstn);

INT_PSE #(.ASIZE(27),.SC_PSE(SC_PSE_Y0)) U1_PSE(.A(y0_sel),.SIGN(y0_signed_sel),.A_PSE(Y0_PSE));
INT_PSE #(.ASIZE(27),.SC_PSE(SC_PSE_H0)) U2_PSE(.A(H0),    .SIGN(H0_SIGNED),    .A_PSE(H0_PSE));

initial begin
    {h0_signed_d, h0_d} = 'b0;
    {y0_signed_d, y0_d} = 'b0;
end

INT_REG #(.SIZE(1)) USEL (.Q(s0_d_sel),
    .BYPASS(INREG_EN == "TRUE" ? 1'b0 : 1'b1),
    .D(S0),
    .CLK(CLK), .CE(CE), .ARST(rst_asyncomb), .SRST(RST_sync));
assign s0_sel = (DYN_OP_SEL == 1'b1) ? s0_d_sel : INPUT_OP[0];

always @(posedge CLK or posedge rst_asyncomb)
    if (rst_asyncomb || RST_sync) begin
        {h0_signed_d, h0_d} <= 'b0;
        {y0_signed_d, y0_d} <= 'b0;
    end
    else if (CE) begin
        {h0_signed_d, h0_d} <= {H0_SIGNED, H0_PSE};
        {y0_signed_d, y0_d} <= {y0_signed_sel, Y0_PSE};
    end

assign {h0_signed_d_sel, h0_d_sel} = (INREG_EN == "TRUE")? {h0_signed_d, h0_d} : {H0_SIGNED, H0_PSE};
assign {y0_signed_d_sel, y0_d_sel} = (INREG_EN == "TRUE")? {y0_signed_d, y0_d} : {y0_signed_sel, Y0_PSE};

assign {y0_signed_sel, y0_sel} = (s0_sel == 1'b1)? {CYI_SIGNED, CYI} : {Y0_SIGNED, Y0}; // default S0 = 1 

assign {cyo_signed, cyo} = {y0_signed_d_sel, y0_d_sel};


assign mult1_in1 = {{27{y0_signed_d_sel & y0_d_sel[26]}},y0_d_sel};
assign mult1_in2 = {{27{h0_signed_d_sel & h0_d_sel[26]}},h0_d_sel}; 

assign mult1 = mult1_in1 * mult1_in2;
assign mult1_signed = y0_signed_d_sel | h0_signed_d_sel;

assign sum = {{10{mult1_signed & mult1[53]}},mult1} + CPI_SEL;
assign sum_signed = mult1_signed | CPI_SIGNED;


always @(posedge CLK or posedge rst_asyncomb)
    if (rst_asyncomb || RST_sync) begin
        {cyo_signed_d, cyo_d} <= 'b0;
        {sum_signed_d, sum_d} <= 65'b0;
    end
    else if (CE) begin
        {cyo_signed_d, cyo_d} <= {cyo_signed, cyo};
        {sum_signed_d, sum_d} <= {sum_signed, sum};
    end

assign {CYO_SIGNED, CYO} = (OUTREG_EN == "TRUE")? {cyo_signed_d, cyo_d}: {cyo_signed, cyo};
assign {CPO_SIGNED, CPO} = (OUTREG_EN == "TRUE")? {sum_signed_d, sum_d}: {sum_signed, sum};
assign P = CPO;

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_INBUFGDS.v
//
// Functional description: Differential Signaling Input Clock Buffer
//
// Parameter description:
//
// Port description:
//
// Revision:
//    06/18/14 - Initial version.
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_INBUFGDS #(
    parameter IOSTANDARD = "DEFAULT",
    parameter TERM_DIFF = "ON"
)(
    output reg O,
    input I,
    input IB
) /* synthesis syn_black_box */ ;

  
  initial begin
    case (IOSTANDARD)
    "LVDS", "MINI-LVDS", "LVPECL", "SUB-LVDS", "SSTL18D_I", "SSTL18D_II", "SSTL15D_I", "SSTL15D_II", "HSTL18D_I", "HSTL18D_II", "HSTL15D_I", "SSTL25D_I", "RSDS", "PPDS", "TMDS", "SSTL25D_II", "BLVDS", "SSTL15D_I_CAL", "SSTL15D_II_CAL", "HSTL15D_I_CAL", "DEFAULT" :;
    default : begin
           $display("Attribute Syntax Error : The attribute IOSTANDARD on GTP_INBUFGDS instance %m is set to %s.", IOSTANDARD);
           $finish;
              end
    endcase

    case (TERM_DIFF)
    "ON", "OFF" :;
    default : begin
           $display("Attribute Syntax Error : The attribute TERM_DIFF on GTP_INBUFGDS instance %m is set to %s.", TERM_DIFF);
           $finish;
              end
    endcase
    end
   
    always @(*)
    begin
        if (I == 1'b1 && IB == 1'b0)
            O = I;
        else if (I == 1'b0 && IB == 1'b1)
            O = I;
        else
            O = 1'bx;
    end

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_PREADD_MULTADD36.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

//P = A0*(B0+-C0) +/- A1*(B1+-C1)
`timescale 1 ns / 1 ps

module GTP_PREADD_MULTADD36 #(
    parameter GRS_EN           = "TRUE", //"TRUE"; "FALSE"
    parameter SYNC_RST         = "FALSE", //"TRUE"; "FALSE"  
    parameter INREG_EN         = "FALSE", //"TRUE"; "FALSE"
    parameter PREREG_EN        = "FALSE", //"TRUE"; "FALSE"
    parameter PIPEREG_EN       = "FALSE", //"TRUE"; "FALSE"
    parameter OUTREG_EN        = "FALSE", //"TRUE"; "FALSE"
    parameter ADDSUB_OP        = 0 ,
    parameter DYN_ADDSUB_OP    = 1
)(
    output  [56-1:0] P,
    input   CE,
    input   RST,
    input   CLK,
    input   [36-1:0] A0,
    input   [36-1:0] A1,
    input   [18-1:0] B0,
    input   [18-1:0] B1,
    input   [18-1:0] C0,
    input   [18-1:0] C1,
    input   A_SIGNED,
    input   B_SIGNED,
    input   C_SIGNED,
    input   [1:0] PREADDSUB,
    input   ADDSUB
);


    INT_PREADD_MULTADD #(
        . GRS_EN(GRS_EN),    
        . SYNC_RST(SYNC_RST),  
        . INREG_EN(INREG_EN), 
        . PREREG_EN(PREREG_EN), 
        . PIPEREG_EN(PIPEREG_EN),
        . OUTREG_EN(OUTREG_EN), 
        . ADDSUB_OP(ADDSUB_OP),   
        . DYN_OP_ADDSUB(DYN_ADDSUB_OP),
        . ASIZE(36), 
        . BSIZE(18)
    ) U_INT_PREADD_MULTADD(
        . CE(CE),
        . RST(RST),
        . CLK(CLK),
        . A0(A0),
        . A1(A1),
        . B0(B0),
        . B1(B1),
        . C0(C0),
        . C1(C1),
        . A_SIGNED(A_SIGNED),
        . B_SIGNED(B_SIGNED),
        . C_SIGNED(C_SIGNED),
        . PREADDSUB(PREADDSUB),
        . ADDSUB(ADDSUB),
        . P(P)
    );   

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_INBUFDS.v
//
// Functional description: Differential Signaling Input Buffer
//
// Parameter description:
//
// Port description:
//
// Revision:
//    06/18/14 - Initial version.
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_INBUFDS #(
    parameter IOSTANDARD = "DEFAULT",
    parameter TERM_DIFF = "ON"
)(
    output reg O,
    input I,
    input IB
) /* synthesis syn_black_box */ ;
  
  initial begin
    case (IOSTANDARD)
    "LVDS", "MINI-LVDS", "LVPECL", "SUB-LVDS", "SSTL18D_I", "SSTL18D_II", "SSTL15D_I", "SSTL15D_II", "HSTL18D_I", "HSTL18D_II", "HSTL15D_I", "SSTL25D_I", "RSDS", "PPDS", "TMDS", "SSTL25D_II", "BLVDS", "SSTL15D_I_CAL", "SSTL15D_II_CAL", "HSTL15D_I_CAL", "DEFAULT" :;
    default : begin
           $display("Attribute Syntax Error : The attribute IOSTANDARD on GTP_INBUFDS instance %m is set to %s.", IOSTANDARD);
           $finish;
              end
    endcase

    case (TERM_DIFF)
    "ON", "OFF" :;
    default : begin
           $display("Attribute Syntax Error : The attribute TERM_DIFF on GTP_INBUFDS instance %m is set to %s.", TERM_DIFF);
           $finish;
              end
    endcase
    end

    always @(*)
    begin
        if (I == 1'b1 && IB == 1'b0)
            O = I;
        else if (I == 1'b0 && IB == 1'b1)
            O = I;
        else
            O = 1'bx;
    end

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2019 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_IOCLKDIV_E3.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//////////////////////////////////////////////////////////////////////////////
//
`timescale 1 ns / 1 ps
module GTP_IOCLKDIV_E3
#(
parameter  DIV_FACTOR ="8",       //"4":quater frequency;"8":eighth frequency;
parameter  PHASE_SHIFT ="0"   //PHASE_SHIFT add 1 = CLKDIVOUT delays for 1 CLKIN cycle;
)(
input  RST,
input  CLKIN,
output CLKDIVOUT
); // synthesis syn_black_box

//synthesis translate_off

reg [2:0] INI_CNT;
reg [2:0] SC_DIV_FACTOR;
reg [2:0] clk_cnt;
reg clk_out_reg;
wire [2:0] cnt_div2;
wire rst_n;

initial
begin
    if ((DIV_FACTOR == "4") || (DIV_FACTOR == "8")) begin
    end
    else
        $display (" GTP_IOCLKDIV_E3 error: illegal setting for DIV_FACTOR");

    if ((PHASE_SHIFT == "0") || (PHASE_SHIFT == "1") || (PHASE_SHIFT == "2") || (PHASE_SHIFT == "3") || (PHASE_SHIFT == "4") || (PHASE_SHIFT == "5") || (PHASE_SHIFT == "6") || (PHASE_SHIFT == "7")) begin
    end
    else
        $display (" GTP_IOCLKDIV_E3 error: illegal setting for PHASE_SHIFT");

    case(DIV_FACTOR)
    "4"      :SC_DIV_FACTOR=3'b011;
    "8"      :SC_DIV_FACTOR=3'b111;
     default: SC_DIV_FACTOR=3'b111;
    endcase

    if(DIV_FACTOR == "8")
     begin
       case(PHASE_SHIFT)
       "0"      :INI_CNT=3'b100;
       "1"      :INI_CNT=3'b011;
       "2"      :INI_CNT=3'b010;
       "3"      :INI_CNT=3'b001;
       "4"      :INI_CNT=3'b000;
       "5"      :INI_CNT=3'b111;
       "6"      :INI_CNT=3'b110;
       "7"      :INI_CNT=3'b101;
       default:  INI_CNT=3'b100;
       endcase
     end
    else
     begin
       case(PHASE_SHIFT)
       "0"      :INI_CNT=3'b010;
       "1"      :INI_CNT=3'b001;
       "2"      :INI_CNT=3'b000;
       "3"      :INI_CNT=3'b011;
       default:  INI_CNT=3'b010;
       endcase
     end
   
        if (INI_CNT < SC_DIV_FACTOR) begin
    end
    else
        $display (" GTP_IOCLKDIV_E3 error: illegal setting for PHASE_SHIFT");
end

assign rst_n = ~RST;
assign cnt_div2 = {1'b0,SC_DIV_FACTOR[2:1]} + 1;

always @(posedge CLKIN or negedge rst_n)
begin
    if(!rst_n)
    clk_cnt <= INI_CNT;
    else if(clk_cnt < SC_DIV_FACTOR)
    clk_cnt <= clk_cnt + 3'd1;
    else
    clk_cnt <= 3'd0;
end

always @(posedge CLKIN or negedge rst_n)
begin
    if(!rst_n)
    clk_out_reg <= 0;
    else if(clk_cnt == 3'd0)
    clk_out_reg <= 0;
    else if(clk_cnt == cnt_div2)
    clk_out_reg <= 1;
end

assign CLKDIVOUT = clk_out_reg;
//synthesis translate_on
endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_IMDDR.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_IMDDR #(
parameter GRS_EN = "TRUE", //"TRUE"; "FALSE"
parameter LRS_EN = "TRUE",  //"TRUE"; "FALSE"
parameter DPI_EN = "FALSE"  //"TRUE"; "FALSE"
)(
output  [1:0] Q,
output [1:0] DPI_STS,
input [1:0] DPI_CTRL,
input DPI_STS_CLR_N,
input PADI,
input ICLK,
input RCLK,
input [2:0] IFIFO_WADDR,
input [2:0] IFIFO_RADDR,
input RST
);

//synthesis translate_off
wire [7:0] PADI_D;
reg DPI_P;
reg [1:0] DPI_STS_R;
reg DPI_N_reg;
wire COMP_BEFORE;
wire COMP_AFTER;
wire COMP_BEFORE_D;
wire COMP_AFTER_D;
wire PD_BEFORE;
wire PD_AFTER;
wire DPI_BEFORE_POS_REG_T;
wire DPI_AFTER_POS_REG_T;
wire DPI_BEFORE_NEG_REG_T;
wire DPI_AFTER_NEG_REG_T;
wire AFTER_POS;
wire BEFORE_POS;
wire AFTER_NEG;
wire BEFORE_NEG;
reg DPI_BEFORE;
reg DPI_AFTER;
reg DPI_BEFORE_POS_REG;
reg DPI_BEFORE_NEG_REG;
reg DPI_AFTER_POS_REG;
reg DPI_AFTER_NEG_REG;
reg [7:0] PADI_POS_fifo;
reg [7:0] PADI_NEG_fifo;
reg [1:0] Q_reg;

initial begin
DPI_P              = 0;
DPI_STS_R          = 0;
DPI_N_reg          = 0;
DPI_BEFORE         = 0;
DPI_AFTER          = 0;
DPI_BEFORE_POS_REG = 0;
DPI_BEFORE_NEG_REG = 0;
DPI_AFTER_POS_REG  = 0;
DPI_AFTER_NEG_REG  = 0;
PADI_POS_fifo      = 0;
PADI_NEG_fifo      = 0;
Q_reg              = 0;
end

assign global_rstn = (GRS_EN == "TRUE") ? GRS_INST.GRSNET : 1'b1;
assign lsr_rstn = LRS_EN == "TRUE" ? (~RST) : 1'b1;



assign  #0.05 PADI_D[0] =  PADI;
assign  #0.05 PADI_D[1] =  PADI_D[0];
assign  #0.05 PADI_D[2] =  PADI_D[1];
assign  #0.05 PADI_D[3] =  PADI_D[2];
assign  #0.05 PADI_D[4] =  PADI_D[3];
assign  #0.05 PADI_D[5] =  PADI_D[4];
assign  #0.05 PADI_D[6] =  PADI_D[5];
assign  #0.05 PADI_D[7] =  PADI_D[6];

assign PADI_SAMPLE = (DPI_EN == "TRUE") ? PADI_D[3] : PADI;

always @(posedge ICLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_P <= 0;
   else if (!lsr_rstn)
      DPI_P <= 0;
   else
      DPI_P <= PADI_SAMPLE;
end

always @(negedge ICLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_N_reg <= 0;
   else if (!lsr_rstn)
      DPI_N_reg <= 0;
   else 
      DPI_N_reg <= PADI_SAMPLE;
end

always @(*) begin
   case (DPI_CTRL[1:0])
      2'd0:    begin DPI_BEFORE = PADI_D[2];  DPI_AFTER = PADI_D[4]; end
      2'd1:    begin DPI_BEFORE = PADI_D[1];  DPI_AFTER = PADI_D[5]; end
      2'd2:    begin DPI_BEFORE = PADI_D[0];  DPI_AFTER = PADI_D[6]; end
      default: begin DPI_BEFORE = PADI;       DPI_AFTER = PADI_D[7]; end
   endcase
end

always @(posedge ICLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_BEFORE_POS_REG <= 0;
   else if (!lsr_rstn)
      DPI_BEFORE_POS_REG <= 0;
   else   
      DPI_BEFORE_POS_REG <= DPI_BEFORE;
end

always @(negedge ICLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_BEFORE_NEG_REG <= 0;
   else if (!lsr_rstn)
      DPI_BEFORE_NEG_REG <= 0;
   else     
      DPI_BEFORE_NEG_REG <= DPI_BEFORE;
end


always @(posedge ICLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_AFTER_POS_REG <= 0;
   else if (!lsr_rstn)
      DPI_AFTER_POS_REG <= 0;
   else   
      DPI_AFTER_POS_REG <= DPI_AFTER;
end


always @(negedge ICLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_AFTER_NEG_REG <= 0;
   else if (!lsr_rstn)
      DPI_AFTER_NEG_REG <= 0;
   else     
      DPI_AFTER_NEG_REG <= DPI_AFTER;
end

assign BEFORE_POS = DPI_BEFORE_POS_REG_T ^ DPI_P;
assign DPI_BEFORE_POS_REG_T = (DPI_EN == "TRUE") ? DPI_BEFORE_POS_REG : 0;

assign AFTER_POS = DPI_AFTER_POS_REG_T ^ DPI_P;
assign DPI_AFTER_POS_REG_T = (DPI_EN == "TRUE") ? DPI_AFTER_POS_REG : 0;

assign BEFORE_NEG = DPI_BEFORE_NEG_REG_T ^ DPI_N_reg;
assign DPI_BEFORE_NEG_REG_T = (DPI_EN == "TRUE") ? DPI_BEFORE_NEG_REG : 0;

assign AFTER_NEG = DPI_AFTER_NEG_REG_T ^ DPI_N_reg;
assign DPI_AFTER_NEG_REG_T = (DPI_EN == "TRUE") ? DPI_AFTER_NEG_REG : 0;


assign COMP_BEFORE = BEFORE_POS || BEFORE_NEG;
assign COMP_AFTER = AFTER_POS || AFTER_NEG;

assign #0.1 COMP_BEFORE_D = COMP_BEFORE;
assign #0.1 COMP_AFTER_D = COMP_AFTER;

assign PD_BEFORE = COMP_BEFORE && COMP_BEFORE_D;
assign PD_AFTER = COMP_AFTER && COMP_AFTER_D;


always @(posedge DPI_STS_CLR_N or negedge global_rstn or negedge lsr_rstn or posedge PD_BEFORE) begin
   if (!global_rstn)
      DPI_STS_R[0] <= 0;
   else if (!lsr_rstn)
      DPI_STS_R[0] <= 0;
   else if (PD_BEFORE)     
      DPI_STS_R[0] <= 1'b1;
   else
      DPI_STS_R[0] <= 1'b0;
end

always @(posedge DPI_STS_CLR_N or negedge global_rstn or negedge lsr_rstn or posedge PD_AFTER) begin
   if (!global_rstn)
      DPI_STS_R[1] <= 0;
   else if (!lsr_rstn)
      DPI_STS_R[1] <= 0;
   else if (PD_AFTER)     
      DPI_STS_R[1] <= 1'b1;
   else
      DPI_STS_R[1] <= 1'b0;
end

assign DPI_STS[0] = DPI_STS_R[0];
assign DPI_STS[1] = DPI_STS_R[1];

      
always @(negedge ICLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      PADI_POS_fifo <= 0;
   else if (!lsr_rstn)
      PADI_POS_fifo <= 0;
   else
      PADI_POS_fifo[IFIFO_WADDR] <= DPI_P;

always @(negedge ICLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      PADI_NEG_fifo <= 0;
   else if (!lsr_rstn)
      PADI_NEG_fifo <= 0;
   else
      PADI_NEG_fifo[IFIFO_WADDR] <= PADI_SAMPLE;      
      
always @(posedge RCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      Q_reg <= 0;
   else if (!lsr_rstn)
      Q_reg <= 0;
   else
      Q_reg <= {PADI_NEG_fifo[IFIFO_RADDR], PADI_POS_fifo[IFIFO_RADDR]};      

assign Q = Q_reg;      
//synthesis translate_on

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2019 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_CLKPD.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//////////////////////////////////////////////////////////////////////////////
//
`timescale 1 ns / 1 ps

module GTP_CLKPD (
    //output
    output FLAG_PD,
    output LOCK,
    //input
    input RST,
    input CLK_SAMPLE,
    input CLK_CTRL,
    input CLK_PHY,
    input DONE
)/* synthesis syn_black_box */;

//synthesis translate_off
   //reg statement
    reg cpd_up_reg;
   //wire statement
    wire  dff_clk;
    wire  dff_din;
    reg   SC_CPD_EN;
    reg   cpd_lock;
    
    
    initial
       begin
          SC_CPD_EN = 1'b1;
       end
    

    assign dff_din = CLK_CTRL;
    assign dff_clk = CLK_PHY;
    assign FLAG_PD = cpd_up_reg;
    
    always @(posedge dff_clk or negedge RST)
    begin
       if(!RST)
       begin
          cpd_up_reg <= 1'b1;
       end
       else
       begin
          cpd_up_reg <= dff_din;
       end
    end

reg d0, d1, ioclk, en;
reg [2:0] acc;
wire clk_int, clk_int2, x;

//clock gating, save power
assign clk_int = SC_CPD_EN? CLK_SAMPLE : 1'b0;

always @ (DONE or clk_int)
begin
  if (~clk_int)
    en=~DONE;
end

assign clk_int2 = en & clk_int;
  
//clock divided by 2
always @ (posedge clk_int2 or negedge RST)
begin
if (~RST)
  ioclk <= 1'b0;
else
  ioclk <= ~ioclk;
end

  always @ (posedge ioclk or negedge RST)
    if(~RST) begin
      d0 <= 1'b0;
      d1 <= 1'b0;
    end
    else begin
      d0 <= FLAG_PD;
      d1 <= d0;
    end

assign x = d0 ^ d1;

  always @ (posedge ioclk or negedge RST) begin
    if(~RST) 
      acc <= 3'b000;
    else 
    if(x)
      acc <= acc+ 1'b1;
    else
      acc <= acc;
  end

assign y = d0 & d1;

  always @ (posedge ioclk or negedge RST) begin
    if(~RST)
      cpd_lock<=0;
    else if (acc==3'b100 && y==1'b0)
           cpd_lock <=1;
  end
assign LOCK = cpd_lock;
    //synthesis translate_on
endmodule






//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2016 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_IODELAY_E2.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
/////////////////////////////////////////////////////////////////////////////
`timescale 1 ps / 1 ps

module GTP_IODELAY_E2 #(
parameter       DELAY_STEP_SEL   = "PARAMETER",   // "PARAMETER", "PORT"
parameter [7:0] DELAY_STEP_VALUE = 8'h00          // 8'h00 ~ 8'hF7
)(
output      DO,
input       DI,
input       DELAY_SEL,
input [7:0] DELAY_STEP                       // 8'h00 ~ 8'hF7 

); /* synthesis syn_black_box */ 

//synthesis translate_off
///////////////////////////////////////////////////////////////////////////


wire [7:0]  gray_code;

reg  [61:0] data0_0;
reg  [3:0]  data0_1;
reg  [61:0] data1_0;
reg  [3:0]  data1_1;

reg         gray_code_bit3;
reg  [63:0] therm_code;


initial begin
    if(DELAY_STEP_SEL != "PARAMETER" && DELAY_STEP_SEL != "PORT")
    begin
      $display("Error: Illegal setting DELAY_STEP_SEL of %s",DELAY_STEP_SEL);
      $finish;
    end

    if(DELAY_STEP_VALUE > 8'hF7 || DELAY_STEP_VALUE < 8'h00)    //  248 cases 
    begin
      $display("Error: Illegal setting DELAY_STEP_VALUE of %b",DELAY_STEP_VALUE);
      $finish;
    end
end        


    initial 
    begin
       data0_0 = 62'h0000000000000000;
       data1_0 = 62'h0000000000000000;
       data0_1 = 4'b0000;
       data1_1 = 4'b0000;
    end


    genvar i;
    generate
        always@(*) data0_0[0] <= DI;
        for (i=1; i<=61; i=i+1)
        begin
           always@(*) data0_0[i]  <= #20.0 data0_0[i-1];
        end
    endgenerate

    wire data0_0_out;
    assign data0_0_out = (therm_code[63:3] == 61'h0000000000000000) ? data0_0[0]   : 
                         (therm_code[63:3] == 61'h0000000000000001) ? data0_0[1]   :
                         (therm_code[63:3] == 61'h0000000000000003) ? data0_0[2]   : 
                         (therm_code[63:3] == 61'h0000000000000007) ? data0_0[3]   : 
                         (therm_code[63:3] == 61'h000000000000000F) ? data0_0[4]   :
                         (therm_code[63:3] == 61'h000000000000001F) ? data0_0[5]   :
                         (therm_code[63:3] == 61'h000000000000003F) ? data0_0[6]   : 
                         (therm_code[63:3] == 61'h000000000000007F) ? data0_0[7]   :
                         (therm_code[63:3] == 61'h00000000000000FF) ? data0_0[8]   :
                         (therm_code[63:3] == 61'h00000000000001FF) ? data0_0[9]   : 
                         (therm_code[63:3] == 61'h00000000000003FF) ? data0_0[10]  :
                         (therm_code[63:3] == 61'h00000000000007FF) ? data0_0[11]  :
                         (therm_code[63:3] == 61'h0000000000000FFF) ? data0_0[12]  : 
                         (therm_code[63:3] == 61'h0000000000001FFF) ? data0_0[13]  :
                         (therm_code[63:3] == 61'h0000000000003FFF) ? data0_0[14]  :
                         (therm_code[63:3] == 61'h0000000000007FFF) ? data0_0[15]  : 
                         (therm_code[63:3] == 61'h000000000000FFFF) ? data0_0[16]  :
                         (therm_code[63:3] == 61'h000000000001FFFF) ? data0_0[17]  : 
                         (therm_code[63:3] == 61'h000000000003FFFF) ? data0_0[18]  : 
                         (therm_code[63:3] == 61'h000000000007FFFF) ? data0_0[19]  :
                         (therm_code[63:3] == 61'h00000000000FFFFF) ? data0_0[20]  :
                         (therm_code[63:3] == 61'h00000000001FFFFF) ? data0_0[21]  : 
                         (therm_code[63:3] == 61'h00000000003FFFFF) ? data0_0[22]  :
                         (therm_code[63:3] == 61'h00000000007FFFFF) ? data0_0[23]  :
                         (therm_code[63:3] == 61'h0000000000FFFFFF) ? data0_0[24]  : 
                         (therm_code[63:3] == 61'h0000000001FFFFFF) ? data0_0[25]  :
                         (therm_code[63:3] == 61'h0000000003FFFFFF) ? data0_0[26]  :
                         (therm_code[63:3] == 61'h0000000007FFFFFF) ? data0_0[27]  : 
                         (therm_code[63:3] == 61'h000000000FFFFFFF) ? data0_0[28]  :
                         (therm_code[63:3] == 61'h000000001FFFFFFF) ? data0_0[29]  :
                         (therm_code[63:3] == 61'h000000003FFFFFFF) ? data0_0[30]  :  
                         (therm_code[63:3] == 61'h000000007FFFFFFF) ? data0_0[31]  :
                         (therm_code[63:3] == 61'h00000000FFFFFFFF) ? data0_0[32]  : 
                         (therm_code[63:3] == 61'h00000001FFFFFFFF) ? data0_0[33]  :
                         (therm_code[63:3] == 61'h00000003FFFFFFFF) ? data0_0[34]  : 
                         (therm_code[63:3] == 61'h00000007FFFFFFFF) ? data0_0[35]  : 
                         (therm_code[63:3] == 61'h0000000FFFFFFFFF) ? data0_0[36]  :
                         (therm_code[63:3] == 61'h0000001FFFFFFFFF) ? data0_0[37]  :
                         (therm_code[63:3] == 61'h0000003FFFFFFFFF) ? data0_0[38]  : 
                         (therm_code[63:3] == 61'h0000007FFFFFFFFF) ? data0_0[39]  : 
                         (therm_code[63:3] == 61'h000000FFFFFFFFFF) ? data0_0[40]  :
                         (therm_code[63:3] == 61'h000001FFFFFFFFFF) ? data0_0[41]  : 
                         (therm_code[63:3] == 61'h000003FFFFFFFFFF) ? data0_0[42]  :
                         (therm_code[63:3] == 61'h000007FFFFFFFFFF) ? data0_0[43]  :
                         (therm_code[63:3] == 61'h00000FFFFFFFFFFF) ? data0_0[44]  : 
                         (therm_code[63:3] == 61'h00001FFFFFFFFFFF) ? data0_0[45]  :
                         (therm_code[63:3] == 61'h00003FFFFFFFFFFF) ? data0_0[46]  :
                         (therm_code[63:3] == 61'h00007FFFFFFFFFFF) ? data0_0[47]  : 
                         (therm_code[63:3] == 61'h0000FFFFFFFFFFFF) ? data0_0[48]  :
                         (therm_code[63:3] == 61'h0001FFFFFFFFFFFF) ? data0_0[49]  : 
                         (therm_code[63:3] == 61'h0003FFFFFFFFFFFF) ? data0_0[50]  : 
                         (therm_code[63:3] == 61'h0007FFFFFFFFFFFF) ? data0_0[51]  :
                         (therm_code[63:3] == 61'h000FFFFFFFFFFFFF) ? data0_0[52]  :
                         (therm_code[63:3] == 61'h001FFFFFFFFFFFFF) ? data0_0[53]  : 
                         (therm_code[63:3] == 61'h003FFFFFFFFFFFFF) ? data0_0[54]  : 
                         (therm_code[63:3] == 61'h007FFFFFFFFFFFFF) ? data0_0[55]  :
                         (therm_code[63:3] == 61'h00FFFFFFFFFFFFFF) ? data0_0[56]  : 
                         (therm_code[63:3] == 61'h01FFFFFFFFFFFFFF) ? data0_0[57]  :
                         (therm_code[63:3] == 61'h03FFFFFFFFFFFFFF) ? data0_0[58]  :
                         (therm_code[63:3] == 61'h07FFFFFFFFFFFFFF) ? data0_0[59]  : 
                         (therm_code[63:3] == 61'h0FFFFFFFFFFFFFFF) ? data0_0[60]  : data0_0[61];
                

    wire    data0_1_out;
    genvar j;
    generate
        always@(*) data0_1[0]  <=  data0_0_out;
        for (j=1; j<4; j=j+1)
        begin
           always@(*) data0_1[j]  <= #5.0 data0_1[j-1];
        end
    endgenerate
    assign data0_1_out =  (therm_code[2:0]==3'b000) ? data0_1[0]   :
                        (therm_code[2:0]==3'b001) ? data0_1[1]   :
                        (therm_code[2:0]==3'b011) ? data0_1[2]   : data0_1[3];

   //2X

    genvar m;
    generate 
        always@(*) data1_0[0] <= data0_1_out;
        for (m=1; m<=61; m=m+1)
        begin
           always@(*) data1_0[m]  <= #20.0 data1_0[m-1];
        end
    endgenerate


    wire data1_0_out;
    assign data1_0_out = (therm_code[63:3] == 61'h0000000000000000) ? data1_0[0]   : 
                         (therm_code[63:3] == 61'h0000000000000001) ? data1_0[1]   :
                         (therm_code[63:3] == 61'h0000000000000003) ? data1_0[2]   : 
                         (therm_code[63:3] == 61'h0000000000000007) ? data1_0[3]   : 
                         (therm_code[63:3] == 61'h000000000000000F) ? data1_0[4]   :
                         (therm_code[63:3] == 61'h000000000000001F) ? data1_0[5]   :
                         (therm_code[63:3] == 61'h000000000000003F) ? data1_0[6]   : 
                         (therm_code[63:3] == 61'h000000000000007F) ? data1_0[7]   :
                         (therm_code[63:3] == 61'h00000000000000FF) ? data1_0[8]   :
                         (therm_code[63:3] == 61'h00000000000001FF) ? data1_0[9]   : 
                         (therm_code[63:3] == 61'h00000000000003FF) ? data1_0[10]  :
                         (therm_code[63:3] == 61'h00000000000007FF) ? data1_0[11]  :
                         (therm_code[63:3] == 61'h0000000000000FFF) ? data1_0[12]  : 
                         (therm_code[63:3] == 61'h0000000000001FFF) ? data1_0[13]  :
                         (therm_code[63:3] == 61'h0000000000003FFF) ? data1_0[14]  :
                         (therm_code[63:3] == 61'h0000000000007FFF) ? data1_0[15]  : 
                         (therm_code[63:3] == 61'h000000000000FFFF) ? data1_0[16]  :
                         (therm_code[63:3] == 61'h000000000001FFFF) ? data1_0[17]  : 
                         (therm_code[63:3] == 61'h000000000003FFFF) ? data1_0[18]  : 
                         (therm_code[63:3] == 61'h000000000007FFFF) ? data1_0[19]  :
                         (therm_code[63:3] == 61'h00000000000FFFFF) ? data1_0[20]  :
                         (therm_code[63:3] == 61'h00000000001FFFFF) ? data1_0[21]  : 
                         (therm_code[63:3] == 61'h00000000003FFFFF) ? data1_0[22]  :
                         (therm_code[63:3] == 61'h00000000007FFFFF) ? data1_0[23]  :
                         (therm_code[63:3] == 61'h0000000000FFFFFF) ? data1_0[24]  : 
                         (therm_code[63:3] == 61'h0000000001FFFFFF) ? data1_0[25]  :
                         (therm_code[63:3] == 61'h0000000003FFFFFF) ? data1_0[26]  :
                         (therm_code[63:3] == 61'h0000000007FFFFFF) ? data1_0[27]  : 
                         (therm_code[63:3] == 61'h000000000FFFFFFF) ? data1_0[28]  :
                         (therm_code[63:3] == 61'h000000001FFFFFFF) ? data1_0[29]  :
                         (therm_code[63:3] == 61'h000000003FFFFFFF) ? data1_0[30]  :  
                         (therm_code[63:3] == 61'h000000007FFFFFFF) ? data1_0[31]  :
                         (therm_code[63:3] == 61'h00000000FFFFFFFF) ? data1_0[32]  : 
                         (therm_code[63:3] == 61'h00000001FFFFFFFF) ? data1_0[33]  :
                         (therm_code[63:3] == 61'h00000003FFFFFFFF) ? data1_0[34]  : 
                         (therm_code[63:3] == 61'h00000007FFFFFFFF) ? data1_0[35]  : 
                         (therm_code[63:3] == 61'h0000000FFFFFFFFF) ? data1_0[36]  :
                         (therm_code[63:3] == 61'h0000001FFFFFFFFF) ? data1_0[37]  :
                         (therm_code[63:3] == 61'h0000003FFFFFFFFF) ? data1_0[38]  : 
                         (therm_code[63:3] == 61'h0000007FFFFFFFFF) ? data1_0[39]  : 
                         (therm_code[63:3] == 61'h000000FFFFFFFFFF) ? data1_0[40]  :
                         (therm_code[63:3] == 61'h000001FFFFFFFFFF) ? data1_0[41]  : 
                         (therm_code[63:3] == 61'h000003FFFFFFFFFF) ? data1_0[42]  :
                         (therm_code[63:3] == 61'h000007FFFFFFFFFF) ? data1_0[43]  :
                         (therm_code[63:3] == 61'h00000FFFFFFFFFFF) ? data1_0[44]  : 
                         (therm_code[63:3] == 61'h00001FFFFFFFFFFF) ? data1_0[45]  :
                         (therm_code[63:3] == 61'h00003FFFFFFFFFFF) ? data1_0[46]  :
                         (therm_code[63:3] == 61'h00007FFFFFFFFFFF) ? data1_0[47]  : 
                         (therm_code[63:3] == 61'h0000FFFFFFFFFFFF) ? data1_0[48]  :
                         (therm_code[63:3] == 61'h0001FFFFFFFFFFFF) ? data1_0[49]  : 
                         (therm_code[63:3] == 61'h0003FFFFFFFFFFFF) ? data1_0[50]  : 
                         (therm_code[63:3] == 61'h0007FFFFFFFFFFFF) ? data1_0[51]  :
                         (therm_code[63:3] == 61'h000FFFFFFFFFFFFF) ? data1_0[52]  :
                         (therm_code[63:3] == 61'h001FFFFFFFFFFFFF) ? data1_0[53]  : 
                         (therm_code[63:3] == 61'h003FFFFFFFFFFFFF) ? data1_0[54]  : 
                         (therm_code[63:3] == 61'h007FFFFFFFFFFFFF) ? data1_0[55]  :
                         (therm_code[63:3] == 61'h00FFFFFFFFFFFFFF) ? data1_0[56]  : 
                         (therm_code[63:3] == 61'h01FFFFFFFFFFFFFF) ? data1_0[57]  :
                         (therm_code[63:3] == 61'h03FFFFFFFFFFFFFF) ? data1_0[58]  :
                         (therm_code[63:3] == 61'h07FFFFFFFFFFFFFF) ? data1_0[59]  : 
                         (therm_code[63:3] == 61'h0FFFFFFFFFFFFFFF) ? data1_0[60]  : data1_0[61];
                

    wire    data1_1_out;
    genvar n;
    generate 
        always@(*) data1_1[0]  <=  data1_0_out;
        for (n=1; n<4; n=n+1)
        begin
           always@(*) data1_1[n]  <= #5.0 data1_1[n-1];
        end
    endgenerate
    assign data1_1_out =  (therm_code[2:0]==3'b000) ? data1_1[0]   :
                          (therm_code[2:0]==3'b001) ? data1_1[1]   :
                          (therm_code[2:0]==3'b011) ? data1_1[2]   : data1_1[3];
    assign  DO   =  DELAY_SEL ? data1_1_out : data0_1_out;



assign gray_code = (DELAY_STEP_SEL == "PORT") ? DELAY_STEP : DELAY_STEP_VALUE;

always@(*)
    case(gray_code[7:4])
	4'h0: gray_code_bit3 =  gray_code[3];
	4'h1: gray_code_bit3 =  ~gray_code[3];
	4'h3: gray_code_bit3 =  gray_code[3];
	4'h2: gray_code_bit3 =  ~gray_code[3];
	4'h6: gray_code_bit3 =  gray_code[3];
	4'h7: gray_code_bit3 =  ~gray_code[3];
	4'h5: gray_code_bit3 =  gray_code[3]; 
	4'h4: gray_code_bit3 =  ~gray_code[3];
	4'hc: gray_code_bit3 =  gray_code[3];
	4'hd: gray_code_bit3 =  ~gray_code[3];
	4'hf: gray_code_bit3 =  gray_code[3];
	4'he: gray_code_bit3 =  ~gray_code[3];
	4'ha: gray_code_bit3 =  gray_code[3];
	4'hb: gray_code_bit3 =  ~gray_code[3];
	4'h9: gray_code_bit3 =  gray_code[3];
	4'h8: gray_code_bit3 =  ~gray_code[3];
    endcase

always@(*)
    if(gray_code[7:3] == 5'b10000 )
        therm_code[2:0] = 3'd7       ;
    else
    case({gray_code_bit3, gray_code[2:0]})
        4'h0 : therm_code[2:0] = 3'd0;
	    4'h1 : therm_code[2:0] = 3'd1;
	    4'h3 : therm_code[2:0] = 3'd3;
	    4'h2 : therm_code[2:0] = 3'd7;
	    4'h6 : therm_code[2:0] = 3'd0;
	    4'h7 : therm_code[2:0] = 3'd1;
	    4'h5 : therm_code[2:0] = 3'd3;
	    4'h4 : therm_code[2:0] = 3'd7;
	    4'hc : therm_code[2:0] = 3'd0;
	    4'hd : therm_code[2:0] = 3'd1;
	    4'hf : therm_code[2:0] = 3'd3;
	    4'he : therm_code[2:0] = 3'd7;
	    4'ha : therm_code[2:0] = 3'd0;
	    4'hb : therm_code[2:0] = 3'd1;
	    4'h9 : therm_code[2:0] = 3'd3;
	    4'h8 : therm_code[2:0] = 3'd7;
    endcase

always@(*)
    case(gray_code[7:2])
        6'h0 : therm_code[63:3] = 61'h0                ;
	    6'h1 : therm_code[63:3] = 61'h1                ;
	    6'h3 : therm_code[63:3] = 61'h3                ;
	    6'h2 : therm_code[63:3] = 61'h7                ;
	    6'h6 : therm_code[63:3] = 61'hf                ;
	    6'h7 : therm_code[63:3] = 61'h1f               ;
	    6'h5 : therm_code[63:3] = 61'h3f               ;
	    6'h4 : therm_code[63:3] = 61'h7f               ;
	    6'hc : therm_code[63:3] = 61'hff               ;
	    6'hd : therm_code[63:3] = 61'h1ff              ;
	    6'hf : therm_code[63:3] = 61'h3ff              ;
	    6'he : therm_code[63:3] = 61'h7ff              ;
	    6'ha : therm_code[63:3] = 61'hfff              ;
	    6'hb : therm_code[63:3] = 61'h1fff             ;
	    6'h9 : therm_code[63:3] = 61'h3fff             ;
	    6'h8 : therm_code[63:3] = 61'h7fff             ;
	    6'h18: therm_code[63:3] = 61'hffff             ;
	    6'h19: therm_code[63:3] = 61'h1ffff            ;
	    6'h1b: therm_code[63:3] = 61'h3ffff            ;
	    6'h1a: therm_code[63:3] = 61'h7ffff            ;
	    6'h1e: therm_code[63:3] = 61'hfffff            ;
	    6'h1f: therm_code[63:3] = 61'h1fffff           ;
	    6'h1d: therm_code[63:3] = 61'h3fffff           ;
	    6'h1c: therm_code[63:3] = 61'h7fffff           ;
	    6'h14: therm_code[63:3] = 61'hffffff           ;
	    6'h15: therm_code[63:3] = 61'h1ffffff          ;
	    6'h17: therm_code[63:3] = 61'h3ffffff          ;
	    6'h16: therm_code[63:3] = 61'h7ffffff          ;
	    6'h12: therm_code[63:3] = 61'hfffffff          ;
	    6'h13: therm_code[63:3] = 61'h1fffffff         ;
	    6'h11: therm_code[63:3] = 61'h3fffffff         ;
	    6'h10: therm_code[63:3] = 61'h7fffffff         ;
        6'h30: therm_code[63:3] = 61'hffffffff         ; 
        6'h31: therm_code[63:3] = 61'h1ffffffff        ; 
        6'h33: therm_code[63:3] = 61'h3ffffffff        ; 
	    6'h32: therm_code[63:3] = 61'h7ffffffff        ; 		  
        6'h36: therm_code[63:3] = 61'hfffffffff        ; 
        6'h37: therm_code[63:3] = 61'h1fffffffff       ; 
        6'h35: therm_code[63:3] = 61'h3fffffffff       ; 
        6'h34: therm_code[63:3] = 61'h7fffffffff       ; 
        6'h3c: therm_code[63:3] = 61'hffffffffff       ; 
        6'h3d: therm_code[63:3] = 61'h1ffffffffff      ; 
        6'h3f: therm_code[63:3] = 61'h3ffffffffff      ; 
        6'h3e: therm_code[63:3] = 61'h7ffffffffff      ; 
        6'h3a: therm_code[63:3] = 61'hfffffffffff      ; 
        6'h3b: therm_code[63:3] = 61'h1fffffffffff     ; 
        6'h39: therm_code[63:3] = 61'h3fffffffffff     ; 
        6'h38: therm_code[63:3] = 61'h7fffffffffff     ; 
        6'h28: therm_code[63:3] = 61'hffffffffffff     ; 
        6'h29: therm_code[63:3] = 61'h1ffffffffffff    ;
        6'h2b: therm_code[63:3] = 61'h3ffffffffffff    ;
        6'h2a: therm_code[63:3] = 61'h7ffffffffffff    ;
        6'h2e: therm_code[63:3] = 61'hfffffffffffff    ;
        6'h2f: therm_code[63:3] = 61'h1fffffffffffff   ;
        6'h2d: therm_code[63:3] = 61'h3fffffffffffff   ;
        6'h2c: therm_code[63:3] = 61'h7fffffffffffff   ;
        6'h24: therm_code[63:3] = 61'hffffffffffffff   ; 
        6'h25: therm_code[63:3] = 61'h1ffffffffffffff  ;
	    6'h27: therm_code[63:3] = 61'h3ffffffffffffff  ;
        6'h26: therm_code[63:3] = 61'h7ffffffffffffff  ;
        6'h22: therm_code[63:3] = 61'hfffffffffffffff  ;
        6'h23: therm_code[63:3] = 61'h1fffffffffffffff ;
	default    therm_code[63:3] = 61'h1fffffffffffffff ;
    endcase


//synthesis translate_on      

endmodule                                                                                                    




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_DLL.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//2018/01/09 update code to fix bug 2299
//2018/01/10 fix dv err
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_DLL #(
parameter GRS_EN = "TRUE", //TRUE, FALSE;
parameter FAST_LOCK = "TRUE", //FALSE, TRUE
parameter DELAY_STEP_OFFSET = 0  //-4, -3,-2, -1, 0, 1, 2, 3, 4
)(
output [7:0] DELAY_STEP,
output LOCK,
input CLKIN,
input UPDATE_N,
input RST,
input PWD
)/* synthesis syn_black_box */;

//synthesis translate_off
reg        false_clk;
reg [1:0] pwd_clkin_en;
reg [1:0] pwd_falseclk_en;
reg [10:0] cnt_div;
reg [1:0]  clkin_div_d;
reg [11:0] cnt;
reg [1:0]  state_q;
reg [2:0]  stop_q;
reg        carry_q0;
reg        carry_q1;
reg [7:0]  sample_cnt_reg0;
reg        dll_lock;
reg [7:0]  delay_step_reg;
reg [1:0]  next_state;

wire counter_rst;
wire check_carry;
wire act_carry;
wire update;
wire carry_d;
wire [11:0] cnt_scaled;
wire [8:0] sample_cnt_tmp;
wire [7:0]  sample_cnt;
wire false_clk_tmp;
wire clkin_tmp;
wire clkin_div;


assign global_rstn =  (GRS_EN == "TRUE") ? GRS_INST.GRSNET : 1'b1;
assign lsr_rstn    = ~RST ;

initial 
begin
    if ((GRS_EN == "TRUE")  || (GRS_EN == "FALSE")) begin
    end
    else
        $display (" GTP_DLL error: illegal setting for GRS_EN"); 
    
    if ((FAST_LOCK == "TRUE")  || (FAST_LOCK == "FALSE")) begin
    end
    else
        $display (" GTP_DLL error: illegal setting for FAST_LOCK");

    if ((DELAY_STEP_OFFSET == -4)  || (DELAY_STEP_OFFSET == -3) || (DELAY_STEP_OFFSET == -2)  || (DELAY_STEP_OFFSET == -1) ||(DELAY_STEP_OFFSET == 0)  || (DELAY_STEP_OFFSET == 1) ||(DELAY_STEP_OFFSET == 2)  || (DELAY_STEP_OFFSET == 3) ||(DELAY_STEP_OFFSET == 4)) begin
    end
    else
        $display (" GTP_DLL error: illegal setting for DELAY_STEP_OFFSET");

    false_clk = 0;
    pwd_falseclk_en = 2'b0;
    pwd_clkin_en = 2'b0;
    cnt_div = 11'b0;
    clkin_div_d = 2'b0;
    cnt = 12'b0;
    state_q = 2'b0;
    stop_q = 3'b0;
    carry_q0 = 1'b0;
    carry_q1 = 1'b0;
    sample_cnt_reg0 = 8'b0;
    dll_lock = 1'b0;
    delay_step_reg = 8'b0;
    next_state = 2'b0;
end

always #6.4 false_clk = ~ false_clk;

always @(negedge false_clk or negedge global_rstn or negedge lsr_rstn)
begin
    if(!global_rstn)
    pwd_falseclk_en <= 2'b0;
    else if(!lsr_rstn)
    pwd_falseclk_en <= 2'b0;
    else
    begin
        pwd_falseclk_en[0] <= PWD;
        pwd_falseclk_en[1] <= pwd_falseclk_en[0];
    end
end

always @(negedge CLKIN or negedge global_rstn or negedge lsr_rstn)
begin
    if(!global_rstn)
    pwd_clkin_en <= 2'b0;
    else if(!lsr_rstn)
    pwd_clkin_en <= 2'b0;
    else
    begin
        pwd_clkin_en[0] <= PWD;
        pwd_clkin_en[1] <= pwd_clkin_en[0];
    end
end

assign false_clk_tmp = (~pwd_falseclk_en[1])&&false_clk;

assign clkin_tmp = (~pwd_clkin_en[1])&&CLKIN;

always @(negedge clkin_tmp or negedge global_rstn or negedge lsr_rstn)
begin
    if (!global_rstn)
        cnt_div <= 0;
    else if (!lsr_rstn)
        cnt_div <= 0;
    else
        cnt_div <= cnt_div + 1;
end

assign clkin_div = cnt_div[10];

always @(negedge false_clk_tmp or negedge global_rstn or negedge lsr_rstn)
begin
    if (!global_rstn)
        clkin_div_d <= 0; 
    else if (!lsr_rstn)
        clkin_div_d <= 0; 
    else
        clkin_div_d <= {clkin_div_d[0], clkin_div};
end

always @(posedge false_clk_tmp or negedge global_rstn or negedge lsr_rstn or posedge counter_rst)
begin
    if (!global_rstn)
        cnt <= 1; 
    else if (!lsr_rstn)
        cnt <= 1;
    else if (counter_rst)
        cnt <= 1;
    else if (clkin_div_d[1])
        cnt <= cnt + 1;
    else
        cnt <= cnt;
end

always @(posedge false_clk_tmp or negedge global_rstn or negedge lsr_rstn)
begin
    if (!global_rstn)
        state_q <= 2'b00;
    else if (!lsr_rstn)
        state_q <= 2'b00;
    else 
        state_q <= next_state;
end

always @(state_q or clkin_div_d[1] or stop_q)
begin
    case(state_q)
        2'b00: if(clkin_div_d[1])
                next_state = 2'b01;
            else
                next_state = 2'b00;
        2'b01: if(~clkin_div_d[1])
                next_state = 2'b10;
            else
                next_state = 2'b01;
        2'b10: if(clkin_div_d[1] == 1'b0 && stop_q == 3'h7)
                next_state = 2'b11;
            else
                next_state = 2'b10;
        2'b11: begin
                next_state = 2'b00;
            end
    endcase
end

always @(posedge false_clk_tmp or negedge global_rstn or negedge lsr_rstn)
begin
    if(!global_rstn)
        stop_q <= 3'b0;
    else if(!lsr_rstn)
        stop_q <= 3'b0;
    else if(state_q == 2'b10)
        stop_q <= stop_q + 1;
    else
        stop_q <= 3'b0;
end

assign counter_rst = (state_q == 2'b11) ? 1'b1 : 1'b0;

assign check_carry = ((state_q == 2'b10)&&(stop_q == 3'b0)) ? 1'b1 : 1'b0;

assign act_carry = ((stop_q == 3'b010)||(stop_q == 3'b011)) ? 1'b1 : 1'b0;

always @(posedge false_clk_tmp or negedge global_rstn or negedge lsr_rstn)
begin
    if (!global_rstn)
        carry_q0 <= 1'b0;
    else if (!lsr_rstn)
        carry_q0 <= 1'b0;
    else if (check_carry)
        carry_q0 <= carry_d;
end

always @(posedge act_carry or negedge global_rstn or negedge lsr_rstn or posedge counter_rst)
begin
    if (!global_rstn)
        carry_q1 <= 1'b0;
    else if (!lsr_rstn)
        carry_q1 <= 1'b0;
    else 
        carry_q1 <= carry_q0;
end

assign cnt_scaled = cnt[10:0] * (8 + DELAY_STEP_OFFSET)/8;


assign carry_d = carry_q0 ? (cnt_scaled[2]||cnt_scaled[1]) : cnt_scaled[2]&&cnt_scaled[1];

assign sample_cnt_tmp = cnt_scaled[10:3] + carry_q1;

assign sample_cnt = (cnt[11]|cnt_scaled[11]|sample_cnt_tmp[8]) ? 8'b11111111 : sample_cnt_tmp[7:0];

always @(posedge false_clk_tmp or negedge global_rstn or negedge lsr_rstn)
begin
    if (!global_rstn)
        sample_cnt_reg0 <= 0; 
    else if (!lsr_rstn)
        sample_cnt_reg0 <= 0;
    else if (stop_q == 3'b110)
        sample_cnt_reg0 <= sample_cnt;
end

always @(posedge false_clk_tmp or negedge global_rstn or negedge lsr_rstn)
begin
    if (!global_rstn)
        dll_lock <= 1'b0;
    else if (!lsr_rstn)
        dll_lock <= 1'b0;
    else if (stop_q == 3'b110)
        dll_lock <= 1'b1;
end

always @(UPDATE_N or sample_cnt_reg0 or global_rstn or lsr_rstn) 
begin
    if(!global_rstn)
        delay_step_reg = 8'b0;
    else if(!lsr_rstn)
        delay_step_reg = 8'b0;
    else if (~UPDATE_N)
        delay_step_reg = sample_cnt_reg0;
end

assign DELAY_STEP = delay_step_reg;
assign LOCK = dll_lock;

//synthesis translate_on

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////

//P = A*(B+C)
`timescale 1 ns / 1 ps

module INT_PREADD_MULT
#(
    parameter GRS_EN    = "FALSE",  //"TRUE"; "FALSE"
    parameter SYNC_RST  = "FALSE",  //"TRUE"; "FALSE"
    parameter INREG_EN  = "FALSE",  //"TRUE"; "FALSE"
    parameter PREREG_EN = "FALSE",  //"TRUE"; "FALSE"
    parameter OUTREG_EN = "FALSE",  //"TRUE"; "FALSE"
    parameter integer ASIZE = 18,   //LEGAL ASIZE = 9,   18, 27,    36
    parameter integer BSIZE = 18,   //LEGAL BSIZE = 9/8, 18, 27/26, 18
    //PSE parameters
    parameter [ASIZE-2:0] SC_PSE_A = 'b0, //SC_PSE = 0, disable PSE, parameter bit width = ASIZE-1
    parameter [BSIZE-2:0] SC_PSE_B = 'b0, //SC_PSE = 0, disable PSE, parameter bit width = BSIZE-1
    parameter [BSIZE-2:0] SC_PSE_C = 'b0, //SC_PSE = 0, disable PSE, parameter bit width = BSIZE-1
    parameter integer PREADD_EN = 1,
    parameter integer PSIZE = ASIZE + BSIZE + PREADD_EN
) (
    input   CE,
    input   CLK,
    input   RST,
    input   A_SIGNED,
    input   [ASIZE-1:0] A,
    input   B_SIGNED,
    input   [BSIZE-1:0] B,
    input   C_SIGNED,
    input   [BSIZE-1:0] C,
    input   PREADDSUB,
    output  [PSIZE-1:0] P
);

initial begin
    if ((PREADD_EN != 0) && (PREADD_EN != 1))
    begin
        $finish;
    end
    case (ASIZE)
        9:  if ((BSIZE + PREADD_EN) != 9)
            begin
                $finish;
            end
        18, 36: if (BSIZE != 18)
            begin
                $finish;
            end
        27: if ((BSIZE + PREADD_EN) != 27)
            begin
                $finish;
            end
        default :
            $finish;
    endcase
    //$display (" INT_PREADD_MULT error :illegal setting of ASIZE or BSIZE");

    if ((GRS_EN != "TRUE") && (GRS_EN != "FALSE")) begin
        $display("GRS_EN error");
        $finish;
    end
    if ((SYNC_RST != "TRUE") && (SYNC_RST != "FALSE")) begin
        $display("SYNC_RST error");
        $finish;
    end

    if ((INREG_EN != "TRUE") && (INREG_EN != "FALSE")) begin
        $display("INREG_EN error");
        $finish;
    end
    if ((PREREG_EN != "TRUE") && (PREREG_EN != "FALSE")) begin
        $display("PREREG_EN error");
        $finish;
    end
    if ((OUTREG_EN != "TRUE") && (OUTREG_EN != "FALSE")) begin
        $display("OUTREG_EN error");
        $finish;
    end
end      

wire [ASIZE-1:0] A_PSE;
wire [BSIZE-1:0] B_PSE;
wire [BSIZE-1:0] C_PSE;

wire [PSIZE-1:0] P_OUT;
wire [PSIZE-1:0] P_ROUND;

reg  [ASIZE-1:0] a_ireg;
reg  [BSIZE-1:0] b_ireg;
reg  [BSIZE-1:0] c_ireg;
reg  asign_ireg, bsign_ireg, csign_ireg;
reg  preaddsub_ireg;

wire [ASIZE-1:0] a_in;
wire [BSIZE-1:0] b_in;
wire [BSIZE-1:0] c_in;
wire asign_in, bsign_in, csign_in;
wire preaddsub_in;

wire [BSIZE:0] b2prad;
wire [BSIZE:0] c2prad;
wire [BSIZE:0] prad_sum;
wire [BSIZE:0] b_inmux;
wire prad_sign, bsign_inmux;

reg  [ASIZE-1:0] a_pareg;
reg  [BSIZE:0]   b_pareg;
reg  asign_pareg, bsign_pareg;

wire [ASIZE-1:0] a_mult;
wire [BSIZE:0]   b_mult;
wire asign_mult, bsign_mult;

wire [PSIZE-1:0] a_mext;
wire [PSIZE-1:0] b_mext;
wire [PSIZE-1:0] PRODUCT;
reg  [PSIZE-1:0] P_reg;

wire global_rstn, RST_sync, RST_async, rst_asyncomb;

assign global_rstn = (GRS_EN == "FALSE") ? 1'b1 : GRS_INST.GRSNET;
assign RST_sync  = (SYNC_RST == "FALSE") ? 1'b0 : RST;
assign RST_async = (SYNC_RST == "FALSE") ? RST : 1'b0;
assign rst_asyncomb = RST_async | (~global_rstn);

INT_PSE #(.ASIZE(ASIZE), .SC_PSE(SC_PSE_A)) U1_PSE (.A(A), .SIGN(A_SIGNED), .A_PSE(A_PSE));
INT_PSE #(.ASIZE(BSIZE), .SC_PSE(SC_PSE_B)) U2_PSE (.A(B), .SIGN(B_SIGNED), .A_PSE(B_PSE));
INT_PSE #(.ASIZE(BSIZE), .SC_PSE(SC_PSE_C)) U3_PSE (.A(C), .SIGN(C_SIGNED), .A_PSE(C_PSE));

initial begin
    a_ireg = 'b0;
    b_ireg = 'b0;
    c_ireg = 'b0;
    preaddsub_ireg = 1'b0;
    P_reg   = 'b0;
end

always @(posedge CLK or posedge rst_asyncomb)
    if (rst_asyncomb) begin
        {asign_ireg, a_ireg} <= 'b0;
        {bsign_ireg, b_ireg} <= 'b0;
        {csign_ireg, c_ireg} <= 'b0;
        preaddsub_ireg       <= 1'b0;
    end
    else if (RST_sync) begin
        {asign_ireg, a_ireg} <= 'b0;
        {bsign_ireg, b_ireg} <= 'b0;
        {csign_ireg, c_ireg} <= 'b0;
        preaddsub_ireg       <= 1'b0;
    end
    else if (CE) begin
        {asign_ireg, a_ireg} <= {A_SIGNED, A_PSE};
        {bsign_ireg, b_ireg} <= {B_SIGNED, B_PSE};
        {csign_ireg, c_ireg} <= {C_SIGNED, C_PSE};
        preaddsub_ireg       <= PREADDSUB;
    end

assign {asign_in, a_in} = (INREG_EN == "TRUE") ? {asign_ireg, a_ireg} : {A_SIGNED, A_PSE};
assign {bsign_in, b_in} = (INREG_EN == "TRUE") ? {bsign_ireg, b_ireg} : {B_SIGNED, B_PSE};
assign {csign_in, c_in} = (INREG_EN == "TRUE") ? {csign_ireg, c_ireg} : {C_SIGNED, C_PSE};
assign  preaddsub_in    = (INREG_EN == "TRUE") ?  preaddsub_ireg      : PREADDSUB;

assign b2prad = {(bsign_in & b_in[BSIZE-1]), b_in};
assign c2prad = {(csign_in & c_in[BSIZE-1]), c_in};
assign prad_sum  = preaddsub_in ? (b2prad - c2prad) : (b2prad + c2prad);
assign prad_sign = bsign_in | csign_in;


reg preadd_over_flag;
always @(*)begin
  if(preaddsub_in==1'b0 && PREADD_EN==1)begin
    if((bsign_in==1'b1 && b_in[BSIZE-1]==1'b0 && csign_in==1'b0 && prad_sum[BSIZE]==1'b1) || (bsign_in==1'b0 && csign_in==1'b1 && c_in[BSIZE-1]==1'b0 && prad_sum[BSIZE]==1'b1))begin
      preadd_over_flag = 1'b1;
    end
    else begin
      preadd_over_flag = 1'b0;
    end
  end
  else if(preaddsub_in==1'b1 && PREADD_EN==1)begin
    if((bsign_in==1'b1 && b_in[BSIZE-1]==1'b1 && csign_in==1'b0 && prad_sum[BSIZE]==1'b0) || (bsign_in==1'b0 && csign_in==1'b1 && c_in[BSIZE-1]==1'b1 && prad_sum[BSIZE]==1'b1) ||
      (bsign_in ==1'b0 && csign_in==1'b0 && (b_in<c_in)))begin
      preadd_over_flag = 1'b1;
    end
    else begin
      preadd_over_flag = 1'b0;
    end
  end
end

always @(preadd_over_flag) begin
    if (preadd_over_flag==1 && PREADD_EN==1)
    $display("Error: PREADD result is overflow!");
end

always @(*) begin
    if (PREADD_EN && (BSIZE == 26) && (prad_sign == 1'b0))
        if ((preaddsub_in == 1'b1) && (prad_sum[BSIZE] == 1'b1)) begin
            $display("PG30-ERROR: Unexpected function mismatch.");
        end
end

assign b_inmux     = PREADD_EN ? prad_sum : {1'b0, b_in};
assign bsign_inmux = PREADD_EN ? prad_sign : bsign_in;
always @(posedge CLK or posedge rst_asyncomb)
    if (rst_asyncomb) begin
        {asign_pareg, a_pareg} <= 'b0;
        {bsign_pareg, b_pareg} <= 'b0;
    end
    else if (RST_sync) begin
        {asign_pareg, a_pareg} <= 'b0;
        {bsign_pareg, b_pareg} <= 'b0;
    end
    else if (CE) begin
        {asign_pareg, a_pareg} <= {asign_in, a_in};
        {bsign_pareg, b_pareg} <= {bsign_inmux, b_inmux};
    end

assign {asign_mult, a_mult} = (PREREG_EN == "TRUE") ? {asign_pareg, a_pareg} : {asign_in, a_in};
assign {bsign_mult, b_mult} = (PREREG_EN == "TRUE") ? {bsign_pareg, b_pareg} : {bsign_inmux, b_inmux};

assign a_mext = {{(PSIZE-ASIZE){asign_mult & a_mult[ASIZE-1]}}, a_mult};
assign b_mext = {{(PSIZE-BSIZE-PREADD_EN){bsign_mult & b_mult[BSIZE+PREADD_EN-1]}}, b_mult[BSIZE+PREADD_EN-1:0]};
assign PRODUCT = a_mext * b_mext;

always @(posedge CLK or posedge rst_asyncomb)
    if (rst_asyncomb) begin
        P_reg <= 'b0;
    end
    else if (RST_sync) begin
        P_reg <= 'b0;
    end
    else if (CE) begin
        P_reg <= PRODUCT;
    end
   
assign P_OUT = (OUTREG_EN == "TRUE") ? P_reg : PRODUCT;

assign P = P_OUT;

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_OGSER4.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_OGSER4 #(
parameter GRS_EN = "TRUE", //"TRUE"; "FALSE" 
parameter LRS_EN = "TRUE"   //"TRUE"; "FALSE" 
)(
output PADO,
output PADT,
input [3:0] D,
input [1:0] T,
input RCLK,
input SERCLK,
input RST
);


//synthesis translate_off
reg [3:0] d_rclk;
reg [1:0] t_rclk;
reg [3:0] capture_d_reg;
reg [1:0] capture_t_reg;
reg [3:0] shift_d_reg;
reg [1:0] shift_t_reg;
reg rstn_dly;
reg capture_en;
reg shift_en;
reg PADO_POS;
reg PADT_reg;
reg PADO_NEG;

initial begin
d_rclk        = 0;
t_rclk        = 0;
capture_d_reg = 0;
capture_t_reg = 0;
shift_d_reg   = 0;
shift_t_reg   = 0;
rstn_dly      = 0;
capture_en      = 0;
PADO_POS      = 0;
PADT_reg      = 0;
PADO_NEG      = 0;  
shift_en      = 0;
end

assign global_rstn = (GRS_EN == "TRUE") ? GRS_INST.GRSNET : 1'b1;
assign lsr_rstn = LRS_EN == "TRUE" ? (~RST) : 1'b1;

always @(posedge RCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn) begin
      d_rclk <= 0;
      t_rclk <= 0;
   end
   else if (!lsr_rstn) begin
      d_rclk <= 0;
      t_rclk <= 0;
   end   
   else begin
      d_rclk <= D;
      t_rclk <= T;    
   end   

always @(posedge SERCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn) begin
      rstn_dly       <= 0;
      capture_en <= 0;
   end
   else if (!lsr_rstn) begin
      rstn_dly       <= 0;
      capture_en <= 0;
   end   
   else begin
      rstn_dly       <= 1;
      if (rstn_dly)
        capture_en <= ~ capture_en;     
      
      shift_en <= capture_en;  
   end
   
always @(posedge SERCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn) begin
      capture_d_reg <= 0;
      capture_t_reg <= 0;
   end
   else if (!lsr_rstn) begin
      capture_d_reg <= 0;
      capture_t_reg <= 0;
   end   
   else begin
      if (capture_en) begin
         capture_d_reg <= d_rclk;
         capture_t_reg <= t_rclk;     
      end
   end 
   
always @(posedge SERCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn) begin
      shift_d_reg <= 0;
      shift_t_reg <= 0;
   end
   else if (!lsr_rstn) begin
      shift_d_reg <= 0;
      shift_t_reg <= 0;
   end   
   else begin
      if (shift_en) begin
         shift_d_reg <= capture_d_reg;
         shift_t_reg <= capture_t_reg;    
      end
      else begin
         shift_d_reg <= {2'd0, shift_d_reg[3:2]};
         shift_t_reg <= {1'b0, shift_t_reg[1]};             
      end
   end
   
always @(posedge SERCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn) begin
      PADO_POS <= 0;
      PADT_reg <= 0;
   end
   else if (!lsr_rstn) begin
      PADO_POS <= 0;
      PADT_reg <= 0;
   end
   else begin
      PADO_POS <= shift_d_reg[1];
      PADT_reg <= shift_t_reg[0];     
   end           
   
always @(negedge SERCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn) begin
      PADO_NEG <= 0;
   end
   else if (!lsr_rstn) begin
      PADO_NEG <= 0;
   end
   else begin
      PADO_NEG <= shift_d_reg[0];
   end           
   
assign PADO =  SERCLK ? PADO_NEG : PADO_POS;
assign PADT = PADT_reg;
//synthesis translate_on

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_MULTADD27.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

//P = A0*B0 +/- A1*B1
module GTP_MULTADD27 #(
    parameter GRS_EN        = "TRUE", //"TRUE"; "FALSE"
    parameter SYNC_RST      = "FALSE", //"TRUE"; "FALSE"
    parameter INREG_EN      = "FALSE", //"TRUE"; "FALSE"
    parameter PIPEREG_EN    = "FALSE", //"TRUE"; "FALSE"
    parameter OUTREG_EN     = "FALSE", //"TRUE"; "FALSE"
    parameter ADDSUB_OP     = 0 ,
    parameter DYN_ADDSUB_OP = 1
)(
    output  [55-1:0] P,          //product
    input   CE,
    input   RST,
    input   CLK,
    input   A_SIGNED,
    input   [27-1:0] A0,
    input   [27-1:0] A1,
    input   B_SIGNED,
    input   [27-1:0] B0,
    input   [27-1:0] B1,
    input   ADDSUB
);

    INT_PREADD_MULTADD #(
        . GRS_EN(GRS_EN),
        . SYNC_RST(SYNC_RST),   
        . INREG_EN(INREG_EN),   
        . PIPEREG_EN(PIPEREG_EN), 
        . OUTREG_EN(OUTREG_EN),  
        . ADDSUB_OP(ADDSUB_OP),  
        . DYN_OP_ADDSUB(DYN_ADDSUB_OP), 
        . ASIZE(27), 
        . BSIZE(27),
        . PREADD_EN(0)
    ) U_MULTADD27 (
        . CE(CE),
        . RST(RST),
        . CLK(CLK),
        . A_SIGNED(A_SIGNED),
        . A0(A0),
        . A1(A1),
        . B_SIGNED(B_SIGNED),
        . B0(B0),
        . B1(B1),
        . C_SIGNED(B_SIGNED),
        . C0(27'b0),
        . C1(27'b0),
        . PREADDSUB(2'b0),
        . ADDSUB(ADDSUB),
        . P(P)
    );

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_DFF_P.v
//
// Functional description: D-type flip-flop with async set
//
// Parameter description:
//      INIT: init value
//
// Port description:
//      P: asynchronous set
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_DFF_P
#(
    parameter GRS_EN = "TRUE",
    parameter INIT = 1'b1
) (
    output reg Q,
    input wire D,
    input wire CLK, P
);

    wire grs_n;
    wire grs, RS;

    tri1 grsnet = GRS_INST.GRSNET;
    assign grs_n=(GRS_EN=="TRUE")?grsnet:1'b1;

    not (grs, grs_n);
    or (RS, grs, P);

    initial Q = 1'bx;

    always @(posedge CLK or posedge RS) begin
        if (RS)
            Q <= 1'b1;
        else
            Q <= D;
    end

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: Internal simulation model
// Filename: GTP_OUTBUFT.v
//
// Functional description: output buffer with tri-state
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_OUTBUFT #(
    parameter IOSTANDARD = "DEFAULT",
    parameter SLEW_RATE = "SLOW",
    parameter DRIVE_STRENGTH = "8"
)(
    output O,
    input I,
    input T
) /* synthesis syn_black_box */ ;

  initial begin
    case (IOSTANDARD)
    "LVTTL33", "PCI33", "LVCMOS33", "LVCMOS25", "LVCMOS18", "LVCMOS15", "LVCMOS12", "SSTL25_I", "SSTL25_II", "SSTL18_I", "SSTL18_II", "SSTL15_I", "SSTL15_II", "HSTL18_I", "HSTL18_II", "HSTL15_I", "SSTL15_I_CAL", "SSTL15_II_CAL", "HSTL15_I_CAL", "DEFAULT" :;
    default : begin
           $display("Attribute Syntax Error : The attribute IOSTANDARD on GTP_OUTBUFT instance %m is set to %s.", IOSTANDARD);
           $finish;
              end
    endcase

    case (SLEW_RATE)
    "FAST", "SLOW":;
    default : begin
           $display("Attribute Syntax Error : The attribute SLEW_RATE on GTP_OUTBUFT instance %m is set to %s.", SLEW_RATE);
           $finish;
              end
    endcase

    case (DRIVE_STRENGTH)
    "2", "4", "6", "8", "12", "16", "24":;
    default : begin
           $display("Attribute Syntax Error : The attribute DRIVE_STRENGTH on GTP_OUTBUFT instance %m is set to %s.", DRIVE_STRENGTH);
           $finish;
              end
    endcase
    end
    bufif0 (O, I, T);

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library:
// Filename: GTP_IOCLKDIV.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_IOCLKDIV #(
parameter DIV_FACTOR = "2", //"2"; "3.5"; "4"; "5"; 
parameter GRS_EN = "TRUE" //"TRUE"; "FALSE"
)(
output CLKDIVOUT,
input CLKIN,
input RST_N
);                        // synthesis syn_black_box

//synthesis translate_off
assign global_rstn = ((GRS_EN == "TRUE" )? GRS_INST.GRSNET : 1'b1);

reg rstn_dly;
reg [3:0] cnt;
reg CLKI_div2;
reg CLKI_DIV_reg;
reg CLKI_DIV_reg_neg;


initial begin
// parameter check
if ((DIV_FACTOR == "2") || (DIV_FACTOR == "3.5") ||  (DIV_FACTOR == "4") || (DIV_FACTOR == "5")) begin
end
else
   $display (" GTP_IOCLKDIV error: illegal setting for DIV_FACTOR");

if ((GRS_EN == "TRUE")  || (GRS_EN == "FALSE")) begin
end
else
   $display (" GTP_IOCLKDIV error: illegal setting for GRS_EN");

rstn_dly          = 0;
cnt               = 0;
CLKI_div2         = 0;
CLKI_DIV_reg      = 0;
CLKI_DIV_reg_neg  = 0;
end


always @(posedge CLKIN or negedge global_rstn or negedge RST_N)
   if (!global_rstn)
      rstn_dly <= 1'b0;
   else if (!RST_N)   
      rstn_dly <= 1'b0;
   else
      rstn_dly <= 1'b1;

always @(posedge CLKIN or negedge rstn_dly)
   if (!rstn_dly)
      CLKI_div2 <= 0;
   else
      CLKI_div2 <= ~ CLKI_div2;

always @(posedge CLKIN or negedge global_rstn or negedge RST_N)
   if (!global_rstn)
      cnt <= 0;
   else if (!RST_N)
      cnt <= 0;
   else if ((DIV_FACTOR == "3.5") && (cnt == 6))
      cnt <= 0;
   else if ((DIV_FACTOR == "4") && (cnt == 7))
      cnt <= 0;
   else if ((DIV_FACTOR == "5") && (cnt == 9))
      cnt <= 0;
   else   
      cnt <= cnt + 1;

always @(posedge CLKIN or negedge global_rstn or negedge RST_N)
   if (!global_rstn)
      CLKI_DIV_reg <= 1'b0;
   else if (!RST_N)
      CLKI_DIV_reg <= 1'b0;
   else if (DIV_FACTOR == "3.5") begin
      if (cnt == 1)
         CLKI_DIV_reg <= 1'b1;
      else if (cnt == 3)   
         CLKI_DIV_reg <= 1'b0;
   end      
   else if (DIV_FACTOR == "4") begin
      if (cnt == 1)
         CLKI_DIV_reg <= 1'b1;
      else if (cnt == 3)   
         CLKI_DIV_reg <= 1'b0;
      else if (cnt == 5)   
         CLKI_DIV_reg <= 1'b1;
      else if (cnt == 7)
         CLKI_DIV_reg <= 1'b0;      
   end
   else if (DIV_FACTOR == "5") begin
      if (cnt == 1)
         CLKI_DIV_reg <= 1'b1;
      else if (cnt == 4)   
         CLKI_DIV_reg <= 1'b0;
      else if (cnt == 6)   
         CLKI_DIV_reg <= 1'b1;
      else if (cnt == 9)
         CLKI_DIV_reg <= 1'b0;          
   end        

always @(negedge CLKIN or negedge global_rstn or negedge RST_N)
   if (!global_rstn)
      CLKI_DIV_reg_neg <= 1'b0;
   else if (!RST_N)
      CLKI_DIV_reg_neg <= 1'b0;     
   else if (DIV_FACTOR == "3.5") begin
      if (cnt == 5)
         CLKI_DIV_reg_neg <= 1'b1;
      else if (cnt == 0)   
         CLKI_DIV_reg_neg <= 1'b0;
   end
      
assign CLKDIVOUT = ((DIV_FACTOR == "2") ? CLKI_div2 : (CLKI_DIV_reg_neg | CLKI_DIV_reg));       
//synthesis translate_on


endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_IGDDR.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_IGDDR #(
parameter GRS_EN = "TRUE", //"TRUE"; "FALSE"
parameter LRS_EN = "TRUE",  //"TRUE"; "FALSE"
parameter DPI_EN = "FALSE"  //"TRUE"; "FALSE"
)(
output  [1:0] Q,
output [1:0] DPI_STS,
input [1:0] DPI_CTRL,
input DPI_STS_CLR_N,
input PADI,
input RCLK,
input RST
);
//synthesis translate_off
wire [7:0] PADI_D;
reg DPI_P;
reg [1:0] DPI_STS_R;
reg DPI_N_reg;
wire COMP_BEFORE;
wire COMP_AFTER;
wire COMP_BEFORE_D;
wire COMP_AFTER_D;
wire PD_BEFORE;
wire PD_AFTER;
wire DPI_BEFORE_POS_REG_T;
wire DPI_AFTER_POS_REG_T;
wire DPI_BEFORE_NEG_REG_T;
wire DPI_AFTER_NEG_REG_T;
wire AFTER_POS;
wire BEFORE_POS;
wire AFTER_NEG;
wire BEFORE_NEG;
reg DPI_BEFORE;
reg DPI_AFTER;
reg DPI_BEFORE_POS_REG;
reg DPI_BEFORE_NEG_REG;
reg DPI_AFTER_POS_REG;
reg DPI_AFTER_NEG_REG;
reg [1:0] Q_reg;

initial begin
   DPI_P              = 0;
   DPI_STS_R          = 0;
   DPI_N_reg          = 0;
   DPI_BEFORE         = 0;
   DPI_AFTER          = 0;
   DPI_BEFORE_POS_REG = 0;
   DPI_BEFORE_NEG_REG = 0;
   DPI_AFTER_POS_REG  = 0;
   DPI_AFTER_NEG_REG  = 0;
   Q_reg              = 0;  
end

assign global_rstn = (GRS_EN == "TRUE") ? GRS_INST.GRSNET : 1'b1;
assign lsr_rstn = LRS_EN == "TRUE" ? (~RST) : 1'b1;

assign  #0.05 PADI_D[0] =  PADI;
assign  #0.05 PADI_D[1] =  PADI_D[0];
assign  #0.05 PADI_D[2] =  PADI_D[1];
assign  #0.05 PADI_D[3] =  PADI_D[2];
assign  #0.05 PADI_D[4] =  PADI_D[3];
assign  #0.05 PADI_D[5] =  PADI_D[4];
assign  #0.05 PADI_D[6] =  PADI_D[5];
assign  #0.05 PADI_D[7] =  PADI_D[6];

assign PADI_SAMPLE = (DPI_EN == "TRUE") ? PADI_D[3] : PADI;

always @(posedge RCLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_P <= 0;
   else if (!lsr_rstn)
      DPI_P <= 0;
   else
      DPI_P <= PADI_SAMPLE;
end

always @(negedge RCLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_N_reg <= 0;
   else if (!lsr_rstn)
      DPI_N_reg <= 0;
   else 
      DPI_N_reg <= PADI_SAMPLE;
end

always @(*) begin
   case (DPI_CTRL[1:0])
      2'd0:    begin DPI_BEFORE = PADI_D[2];  DPI_AFTER = PADI_D[4]; end
      2'd1:    begin DPI_BEFORE = PADI_D[1];  DPI_AFTER = PADI_D[5]; end
      2'd2:    begin DPI_BEFORE = PADI_D[0];  DPI_AFTER = PADI_D[6]; end
      default: begin DPI_BEFORE = PADI;       DPI_AFTER = PADI_D[7]; end
   endcase
end

always @(posedge RCLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_BEFORE_POS_REG <= 0;
   else if (!lsr_rstn)
      DPI_BEFORE_POS_REG <= 0;
   else   
      DPI_BEFORE_POS_REG <= DPI_BEFORE;
end

always @(negedge RCLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_BEFORE_NEG_REG <= 0;
   else if (!lsr_rstn)
      DPI_BEFORE_NEG_REG <= 0;
   else     
      DPI_BEFORE_NEG_REG <= DPI_BEFORE;
end


always @(posedge RCLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_AFTER_POS_REG <= 0;
   else if (!lsr_rstn)
      DPI_AFTER_POS_REG <= 0;
   else   
      DPI_AFTER_POS_REG <= DPI_AFTER;
end


always @(negedge RCLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_AFTER_NEG_REG <= 0;
   else if (!lsr_rstn)
      DPI_AFTER_NEG_REG <= 0;
   else     
      DPI_AFTER_NEG_REG <= DPI_AFTER;
end


assign BEFORE_POS = DPI_BEFORE_POS_REG_T ^ DPI_P;
assign DPI_BEFORE_POS_REG_T = (DPI_EN == "TRUE") ? DPI_BEFORE_POS_REG : 0;

assign AFTER_POS = DPI_AFTER_POS_REG_T ^ DPI_P;
assign DPI_AFTER_POS_REG_T = (DPI_EN == "TRUE") ? DPI_AFTER_POS_REG : 0;

assign BEFORE_NEG = DPI_BEFORE_NEG_REG_T ^ DPI_N_reg;
assign DPI_BEFORE_NEG_REG_T = (DPI_EN == "TRUE") ? DPI_BEFORE_NEG_REG : 0;

assign AFTER_NEG = DPI_AFTER_NEG_REG_T ^ DPI_N_reg;
assign DPI_AFTER_NEG_REG_T = (DPI_EN == "TRUE") ? DPI_AFTER_NEG_REG : 0;


assign COMP_BEFORE = BEFORE_POS || BEFORE_NEG;
assign COMP_AFTER = AFTER_POS || AFTER_NEG;

assign #0.1 COMP_BEFORE_D = COMP_BEFORE;
assign #0.1 COMP_AFTER_D = COMP_AFTER;

assign PD_BEFORE = COMP_BEFORE && COMP_BEFORE_D;
assign PD_AFTER = COMP_AFTER && COMP_AFTER_D;


always @(posedge DPI_STS_CLR_N or negedge global_rstn or negedge lsr_rstn or posedge PD_BEFORE) begin
   if (!global_rstn)
      DPI_STS_R[0] <= 0;
   else if (!lsr_rstn)
      DPI_STS_R[0] <= 0;
   else if (PD_BEFORE)     
      DPI_STS_R[0] <= 1'b1;
   else
      DPI_STS_R[0] <= 1'b0;
end

always @(posedge DPI_STS_CLR_N or negedge global_rstn or negedge lsr_rstn or posedge PD_AFTER) begin
   if (!global_rstn)
      DPI_STS_R[1] <= 0;
   else if (!lsr_rstn)
      DPI_STS_R[1] <= 0;
   else if (PD_AFTER)     
      DPI_STS_R[1] <= 1'b1;
   else
      DPI_STS_R[1] <= 1'b0;
end

assign DPI_STS[0] = DPI_STS_R[0];
assign DPI_STS[1] = DPI_STS_R[1];

always @(posedge RCLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      Q_reg <= 0;
   else if (!lsr_rstn)
      Q_reg <= 0;
   else
      Q_reg <= {DPI_N_reg, DPI_P};      
end

assign Q = Q_reg;      
//synthesis translate_on

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2016 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General Technology Primitive
// Filename: GTP_OSC_E3.v
//
// Functional description: oscillator
//
// Parameter description:
// CLK_DIV:    CLKOUT frequency setting( f = 200MHz/CLK_DIV )[f=200MHz/128, when CLK_DIV=0]
//
// Port description:
// inputs:
// EN_N:           OSC enable
// RST_N:        Reset clock divider
//
// outputs:
// CLKOUT:    100MHz(default)
//
// Revision: V1.0
//
//////////////////////////////////////////////////////////////////////////////
`timescale 1ns/1ps

module GTP_OSC_E3
   #(
     parameter integer CLK_DIV = 2
     )
    (
     output CLKOUT,
    
     input  EN_N,
     input  RST_N
     )/* synthesis syn_black_box */;

    //synthesis translate_off
    wire    rst_wire;
    wire    oscen_wire;
    reg     clk_400_reg; // intrinsic frequency
    reg [6:0] div_reg;
    reg [6:0] count_reg;
    reg       clk_user_reg;
    reg       rst_reg;

    initial 
    begin
        // parameter check
        if ( (CLK_DIV >= 0) && (CLK_DIV <= 127) )
        begin
            div_reg = CLK_DIV;
        end
        else
        begin
            $display ("GTP_OSC_E3 error: illegal setting for CLK_DIV(0 ~ 127)");
        end

        // analog //
        clk_400_reg = 1'b0;

        // divider //
        count_reg = 7'b0000000;
        clk_user_reg = 1'b0;
        rst_reg = 1'b0;
    end
    
    assign rst_wire = !RST_N || EN_N;
    assign oscen_wire = !EN_N;
    assign CLKOUT = clk_user_reg;
    
    // osc_analog //
    always
    begin
        wait (oscen_wire == 1'b1)
           begin
               clk_400_reg = 1'b0;
               #1.25;
               clk_400_reg = 1'b1;
               #1.25;
           end
    end

    always
    begin
        wait (oscen_wire != 1'b1)
           begin
               force clk_400_reg = 1'b0;
               #2 release clk_400_reg;
           end
    end
    // end of osc_analog //
    
    // osc_divider_128 //
    always @ (posedge clk_400_reg or posedge rst_wire)
    begin
        if (rst_wire)
        begin
            clk_user_reg <= 1'b0;
            count_reg <= 7'b000_0000;
            rst_reg <= 1'b1;
        end
        else if (rst_reg)
        begin
            rst_reg <= 1'b0;
            clk_user_reg <= 1'b1;
            count_reg <= 7'b000_0000;
        end
        else if (count_reg == div_reg-7'b1)
        begin
            clk_user_reg <= ~clk_user_reg;
            count_reg <= 7'b000000;
        end
        else
        begin
            clk_user_reg <= clk_user_reg;
            count_reg <= count_reg + 1'b1;
        end
    end
    // end of osc_divider_128 //
    
    //synthesis translate_on
endmodule // GTP_OSC_E3




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_PREADD_FIR_A.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_PREADD_FIR_A
#(
    parameter GRS_EN    = "TRUE", //"TRUE"; "FALSE"
    parameter SYNC_RST  = "FALSE", //"TRUE"; "FALSE"
    parameter INREG_EN  = "TRUE",
    parameter INREG_Z1_EN  = "TRUE",
    parameter OUTREG_EN = "TRUE",
    parameter INPUT_OP    = 8'b11000110,
    parameter DYN_OP_SEL  = 8'b11111111,
    parameter OPCD_DYN_SEL = 1'b0,
    parameter OPCD_CPI_SEL = 1'b0
) (
    output  [17:0] CYO,
    output        CYO_SIGNED,
    output  [63:0] CPO,                  //p
    output         CPO_SIGNED,
    output [17:0] CZO,
    output        CZO_SIGNED,
    output  [63:0] P,                  //p

    input   CE,
    input   RST,
    input   CLK,
    input [17:0] CYI,
    input        CYI_SIGNED,
    input [17:0] Y0,                  //y0 ,DYIA
    input        Y0_SIGNED,
    input [17:0] Z0,                  //z0 ,DZIA
    input        Z0_SIGNED,            
    input [17:0] H0,                  //h0 ,DXIA
    input        H0_SIGNED,
    input [17:0] H1,                  //h1 ,DXIB
    input        H1_SIGNED,
    input [17:0] Y1,                  //y1 ,DYIB
    input        Y1_SIGNED,
    input [17:0] Z1,                  //z1, DZIB
    input        Z1_SIGNED,
    input [17:0] CZI,
    input        CZI_SIGNED,
    input [63:0] CPI,
    input        CPI_SIGNED,
    input        S0,
    input        S1,
    input [5:0]  DYN_OP,
    input        OPCD_CPI_DYN
);

//PSE parameters
localparam [16:0] SC_PSE_Y0 = 17'b0;  //SC_PSE = 0, disable PSE, parameter bit width=17
localparam [16:0] SC_PSE_Y1 = 17'b0;  //SC_PSE = 0, disable PSE, parameter bit width=17
localparam [16:0] SC_PSE_Z0 = 17'b0;  //SC_PSE = 0, disable PSE, parameter bit width=17
localparam [16:0] SC_PSE_Z1 = 17'b0;  //SC_PSE = 0, disable PSE, parameter bit width=17
localparam [16:0] SC_PSE_H0 = 17'b0;  //SC_PSE = 0, disable PSE, parameter bit width=17
localparam [16:0] SC_PSE_H1 = 17'b0;  //SC_PSE = 0, disable PSE, parameter bit width=17

initial begin
    if ((GRS_EN != "TRUE") && (GRS_EN != "FALSE")) begin
        $display("GRS_EN error");
        $finish;
    end
    if ((SYNC_RST != "TRUE") && (SYNC_RST != "FALSE")) begin
        $display("SYNC_RST error");
        $finish;
    end

    if (DYN_OP_SEL[5:3] != 3'b111) begin
        $display("DRC ERROR");
        $finish;
    end
end

wire [7:0] dyn_op;
reg [17:0] h0_d;
reg        h0_signed_d;
wire [17:0] h0_d_sel;
wire        h0_signed_d_sel;
reg [17:0] y0_d;
reg        y0_signed_d;
wire [17:0] y0_d_sel;
wire        y0_signed_d_sel;

wire [17:0] y0_sel;
wire        y0_signed_sel;

reg [17:0] z0_d;
reg        z0_signed_d;

wire [17:0] z0_sel;
wire        z0_signed_sel;

reg [17:0] h1_d;
reg        h1_signed_d;
wire [17:0] h1_d_sel;
wire        h1_signed_d_sel;
reg [17:0] y1_d;
reg        y1_signed_d;
wire [17:0] y1_d_sel;
wire        y1_signed_d_sel;
reg [17:0] z1_d;
reg        z1_signed_d;
wire [17:0] z1_d_sel;
wire        z1_signed_d_sel;

wire [17:0] y1_sel;
wire        y1_signed_sel;
wire [17:0] z1_sel;
wire        z1_signed_sel;

wire [17:0] czi_sel;
wire        czi_sel_signed;

wire [18:0] preadd_1;
wire        preadd_1_signed;
wire [18:0] preadd_2;
wire        preadd_2_signed;

wire [36:0] mult1_in1;
wire [36:0] mult2_in1;
wire [36:0] mult1_in2;
wire [36:0] mult2_in2;

wire [36:0] mult1;
wire        mult1_signed;
wire [36:0] mult2;
wire        mult2_signed;

wire [63:0] ma, mb;
wire [63:0] sum;
wire        sum_signed;

wire [7:0] INPUT_OP_CODE;

wire [17:0] cyo;
wire        cyo_signed;

wire global_rstn ;
wire RST_sync ;
wire RST_async;
wire rst_asyncomb ;

reg [63:0]  CPO_d ;
reg [17:0]  CYO_d ;
reg  CPO_SIGNED_d ;
reg  CYO_SIGNED_d ;

wire [17:0] Y0_PSE; 
wire [17:0] Y1_PSE; 
wire [17:0] H0_PSE;
wire [17:0] H1_PSE;
wire [17:0] Z0_PSE;
wire [17:0] Z1_PSE;

wire [63:0] CPI_SEL;
wire        OPCD_SEL;

assign global_rstn = GRS_EN == "TRUE" ? GRS_INST.GRSNET : 1'b1;
assign RST_sync = (SYNC_RST == "TRUE") ? RST : 1'b0;
assign RST_async = (SYNC_RST == "FALSE") ? RST : 1'b0;
assign rst_asyncomb = RST_async | (~global_rstn);

assign OPCD_SEL = (OPCD_DYN_SEL == 1'b1)?OPCD_CPI_DYN :OPCD_CPI_SEL;
assign CPI_SEL  = (OPCD_SEL == 1'b1)? 64'b0 : CPI;

INT_REG #(.SIZE(8)) USEL (.Q(dyn_op),
    .BYPASS(INREG_EN == "TRUE" ? 1'b0 : 1'b1),
    .D({S0, S1, DYN_OP}),
    .CLK(CLK), .CE(CE), .ARST(rst_asyncomb), .SRST(RST_sync)
);
assign INPUT_OP_CODE[7] = (DYN_OP_SEL[7]) ? dyn_op[7] : INPUT_OP[7]; //ir_op[0]
assign INPUT_OP_CODE[6] = (DYN_OP_SEL[6]) ? dyn_op[6] : INPUT_OP[6]; //ir_op[3]
assign INPUT_OP_CODE[5] = (DYN_OP_SEL[5]) ? dyn_op[5] : INPUT_OP[5]; //ir_op[6]
assign INPUT_OP_CODE[4] = (DYN_OP_SEL[4]) ? dyn_op[4] : INPUT_OP[4]; //ir_op[5]
assign INPUT_OP_CODE[3] = (DYN_OP_SEL[3]) ? dyn_op[3] : INPUT_OP[3]; //ir_op[4]
assign INPUT_OP_CODE[2] = (DYN_OP_SEL[2]) ? dyn_op[2] : INPUT_OP[2]; //ir_op[7]
assign INPUT_OP_CODE[1] = (DYN_OP_SEL[1]) ? dyn_op[1] : INPUT_OP[1]; //ir_op[1]
assign INPUT_OP_CODE[0] = (DYN_OP_SEL[0]) ? dyn_op[0] : INPUT_OP[0]; //ir_op[2]

INT_PSE #(.ASIZE(18),.SC_PSE(SC_PSE_Y0)) U1_PSE(.A(y0_sel),.SIGN(y0_signed_sel),.A_PSE(Y0_PSE));
INT_PSE #(.ASIZE(18),.SC_PSE(SC_PSE_Y1)) U2_PSE(.A(y1_sel),.SIGN(y1_signed_sel),.A_PSE(Y1_PSE));
INT_PSE #(.ASIZE(18),.SC_PSE(SC_PSE_Z0)) U3_PSE(.A(z0_sel),.SIGN(z0_signed_sel),.A_PSE(Z0_PSE));
INT_PSE #(.ASIZE(18),.SC_PSE(SC_PSE_Z1)) U4_PSE(.A(z1_sel),.SIGN(z1_signed_sel),.A_PSE(Z1_PSE));
INT_PSE #(.ASIZE(18),.SC_PSE(SC_PSE_H0)) U5_PSE(.A(H0),    .SIGN(H0_SIGNED),    .A_PSE(H0_PSE));
INT_PSE #(.ASIZE(18),.SC_PSE(SC_PSE_H1)) U6_PSE(.A(H1),    .SIGN(H1_SIGNED),    .A_PSE(H1_PSE));

always @(posedge CLK or posedge rst_asyncomb)
   if (rst_asyncomb || RST_sync) begin
       {h0_signed_d, h0_d} <= 'b0;
       {y0_signed_d, y0_d} <= 'b0;
       {z0_signed_d, z0_d} <= 'b0;
   end
      else if (CE) begin
       {h0_signed_d, h0_d} <= {H0_SIGNED, H0_PSE};
       {y0_signed_d, y0_d} <= {y0_signed_sel, Y0_PSE};
       {z0_signed_d, z0_d} <= {z0_signed_sel, Z0_PSE};
   end

always @(posedge CLK or posedge rst_asyncomb)
   if (rst_asyncomb || RST_sync) begin
       {h1_signed_d, h1_d} <= 'b0;
       {y1_signed_d, y1_d} <= 'b0;
       {z1_signed_d, z1_d} <= 'b0;
   end
      else if (CE) begin
       {h1_signed_d, h1_d} <= {H1_SIGNED, H1_PSE};
       {y1_signed_d, y1_d} <= {y1_signed_sel, Y1_PSE};
       {z1_signed_d, z1_d} <= {z1_signed_sel, Z1_PSE};
   end

assign {h0_signed_d_sel, h0_d_sel} = (INREG_EN == "TRUE")? {h0_signed_d, h0_d} : {H0_SIGNED, H0_PSE};
assign {y0_signed_d_sel, y0_d_sel} = (INREG_EN == "TRUE")? {y0_signed_d, y0_d} : {y0_signed_sel, Y0_PSE};

assign {h1_signed_d_sel, h1_d_sel} = (INREG_EN == "TRUE")? {h1_signed_d, h1_d} : {H1_SIGNED, H1_PSE};
assign {y1_signed_d_sel, y1_d_sel} = (INREG_EN == "TRUE")? {y1_signed_d, y1_d} : {y1_signed_sel, Y1_PSE};
assign {z1_signed_d_sel, z1_d_sel} = (INREG_Z1_EN == "TRUE")? {z1_signed_d, z1_d} : {z1_signed_sel, Z1_PSE};

assign {y1_signed_sel, y1_sel} = (INPUT_OP_CODE[6] == 1'b1)? {y0_signed_d_sel, y0_d_sel} : {Y1_SIGNED, Y1}; //default ir_op[3] = 1, S1            
assign {y0_signed_sel, y0_sel} = (INPUT_OP_CODE[7] == 1'b1)? {CYI_SIGNED     , CYI     } : {Y0_SIGNED, Y0}; //default ir_op[0] = 1, S0
assign {z1_signed_sel, z1_sel} = (INPUT_OP_CODE[2] == 1'b1)? {czi_sel_signed, czi_sel} : {Z1_SIGNED, Z1}; //default ir_op[7] = 1
assign {z0_signed_sel, z0_sel} = (INPUT_OP_CODE[1] == 1'b1)? {czi_sel_signed, czi_sel} : {Z0_SIGNED, Z0}; //default ir_op[1] = 1  

assign {czi_sel_signed, czi_sel} = (INPUT_OP_CODE[5] == 1'b0)? {CZI_SIGNED, CZI} : {CYO_SIGNED, CYO};

assign {cyo_signed, cyo} = (INPUT_OP_CODE[3] == 1'b0)? {y1_signed_d_sel, y1_d_sel} : {y0_signed_d_sel, y0_d_sel}; //default ir_op[4] = 0
assign {CZO_SIGNED, CZO} = (INPUT_OP_CODE[0] == 1'b0)? {z0_signed_d    , z0_d    } : {z0_signed_sel, Z0_PSE};     //default ir_op[2] = 0


assign preadd_1 = {y0_d_sel[17]&y0_signed_d_sel,y0_d_sel} + {CZO[17]&CZO_SIGNED, CZO}; 
assign preadd_1_signed = y0_signed_d_sel | CZO_SIGNED;
assign preadd_2 = {y1_d_sel[17]&y1_signed_d_sel,y1_d_sel} + {z1_d_sel[17]&z1_signed_d_sel, z1_d_sel}; 
assign preadd_2_signed = y1_signed_d_sel | z1_signed_d_sel;

reg preadd_over_flag0;
always @(*)begin
    if((y0_signed_d_sel==1'b1 && y0_d_sel[17]==1'b0 && CZO_SIGNED==1'b0 && preadd_1[18]==1'b1) || (y0_signed_d_sel==1'b0 && CZO_SIGNED==1'b1 && CZO[17]==1'b0 && preadd_1[18]==1'b1))begin
      preadd_over_flag0 = 1'b1;
    end
    else begin
      preadd_over_flag0 = 1'b0;
    end
  end

reg preadd_over_flag1;
always @(*)begin
    if((y1_signed_d_sel==1'b1 && y1_d_sel[17]==1'b0 && z1_signed_d_sel==1'b0 && preadd_2[18]==1'b1) || (y1_signed_d_sel==1'b0 && z1_signed_d_sel==1'b1 && z1_d_sel[17]==1'b0 && preadd_2[18]==1'b1))begin
      preadd_over_flag1 = 1'b1;
    end
    else begin
      preadd_over_flag1 = 1'b0;
    end
  end

always @(preadd_over_flag0 or preadd_over_flag1) begin
    if (preadd_over_flag0==1 || preadd_over_flag1==1)
    $display("Error: PREADD result is overflow!");
end

assign mult1_in1 = {{18{preadd_1_signed & preadd_1[18]}},preadd_1};
assign mult2_in1 = {{18{preadd_2_signed & preadd_2[18]}},preadd_2}; 

assign mult1_in2 = {{19{h0_signed_d_sel & h0_d_sel[17]}},h0_d_sel}; 
assign mult2_in2 = {{19{h1_signed_d_sel & h1_d_sel[17]}},h1_d_sel};

assign mult1 = mult1_in1 * mult1_in2;
assign mult1_signed = preadd_1_signed | h0_signed_d_sel;
assign mult2 = mult2_in1 * mult2_in2;
assign mult2_signed = preadd_2_signed | h1_signed_d_sel;

assign ma = {{27{mult1_signed&mult1[36]}},mult1};
assign mb = {{27{mult2_signed&mult2[36]}},mult2};
assign sum = ma + mb + CPI_SEL;
assign sum_signed = mult1_signed | mult2_signed | CPI_SIGNED;

initial begin
    {h0_signed_d, h0_d} = 'b0;
    {y0_signed_d, y0_d} = 'b0;
    {z0_signed_d, z0_d} = 'b0;
    {CYO_SIGNED_d, CYO_d} = 19'b0;
    {CPO_SIGNED_d, CPO_d} = 65'b0;
end

always @(posedge CLK or posedge rst_asyncomb)
    if (rst_asyncomb || RST_sync) begin
        {CYO_SIGNED_d, CYO_d} <= 19'b0;
        {CPO_SIGNED_d, CPO_d} <= 65'b0;
    end
    else if (CE) begin
        {CYO_SIGNED_d, CYO_d} <= {cyo_signed, cyo};
        {CPO_SIGNED_d, CPO_d} <= {sum_signed, sum};
    end

assign {CYO_SIGNED, CYO} = (INPUT_OP_CODE[4] == 1'b0)? {CYO_SIGNED_d, CYO_d} : {cyo_signed, cyo}; // ir_op[5]
assign {CPO_SIGNED, CPO} = (OUTREG_EN == "TRUE")     ? {CPO_SIGNED_d, CPO_d} : {sum_signed, sum};
assign P= CPO;
endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library:
// Filename: GTP_IOCLKBUF.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_IOCLKBUF
#(
    parameter GATE_EN = "FALSE"   //FALSE; TRUE
) 
(
output CLKOUT,
input CLKIN,
input DI
);       //synthesis syn_black_box 

reg reg1, reg2,reg3;

initial 
begin
  reg1 = 1'b0;
  reg2 = 1'b0;
end


initial 
begin
  if(GATE_EN=="FALSE")
    reg3 =1'b1;
  else
    if(GATE_EN=="TRUE")
       reg3 = 1'b0;
    else 
       $display ("GTP_IOCLKBUF error : illegal setting for GATE_EN");
end



always @(negedge CLKIN) begin
   if(reg3 == 1'b0) 
      begin
         reg2 <= reg1;
         reg1 <= DI;
      end
   else
      begin
        reg2 <= 1'b0;
        reg1 <= 1'b0;
      end
end

assign CLKOUT = (reg2 | reg3) & CLKIN;

endmodule








//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2016 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
//
// GTP model of APML device
//
//
//////////////////////////////////////////////////////////////////////////////
`timescale 1 ns / 1 ps

`define assert(condition, message) \
        if (!(condition)) begin \
            $display($realtime, "ERROR: ASSERTION FAILED in %s, line %d: %s", `__FILE__, `__LINE__, message); \
            $finish; \
        end

// module declaration 
module GTP_APM_E1 #(

    parameter GRS_EN = "TRUE",  //"TRUE","FALSE",enable global reset
    parameter X_SIGNED = 0, //signedness of X. X[17:9] and X[8:0] share the same signedness in mult9x9 mode
    parameter Y_SIGNED = 0, //signedness of Y. Y[17:9] and Y[8:0] share the same signedness in mult9x9 mode

    parameter USE_POSTADD = 0, //enable postadder 0/1
    parameter USE_PREADD = 0,  //enable preadder 0/1
    parameter PREADD_REG = 0,  //preadder reg 0/1

    parameter X_REG = 0,  //X input reg 0/1
    parameter CXO_REG = 0, //X cascade out reg latency, 0/1/2/3
    parameter Y_REG = 0,  //Y input reg 0/1
    parameter Z_REG = 0,  //Z input reg 0/1
    parameter MULT_REG = 0,  //multiplier reg 0/1
    parameter P_REG = 0,  //post adder reg 0/1
    parameter MODEX_REG = 0,  //MODEX reg
    parameter MODEY_REG = 0,  //MODEY reg
    parameter MODEZ_REG = 0,  //MODEZ reg

    parameter X_SEL = 0,  // mult X input select X/CXI
    parameter XB_SEL = 0, //X back propagate mux select. 0/1/2/3
    parameter ASYNC_RST = 0,  // RST is sync/async
    parameter USE_SIMD = 0,   // single addsub18_mult18_add48 / dual addsub9_mult9_add24
    parameter [47:0] Z_INIT = {48{1'b0}},  //Z constant input (RTI parameter in APM of PG family)

    parameter CPO_REG = 0, // CPO,COUT use register output
    parameter USE_ACCLOW = 0, // accumulator use lower 18-bit feedback only
    parameter CIN_SEL = 0 // select CIN for postadder carry in

)(

    output [47:0] P,  //Postadder resout
    output [47:0] CPO, //P cascade out
    output COUT,         //Postadder carry out
    output [17:0] CXO, //X cascade out
    output [17:0] CXBO, //X backward cascade out

    input [17:0] X,
    input [17:0] CXI, //X cascade in
    input [17:0] CXBI, //X backward cascade in
    input [17:0] Y,
    input [47:0] Z,
    input [47:0] CPI, //P cascade in
    input CIN,          //Postadder carry in
    input       MODEX,  // preadder add/sub, 0/1
    input [2:0] MODEY,
// MODEY encoding: 0/1
// [0]     produce all-0 input to post adder / enable P register feedback. MODEY[1] needs to be 1 for MODEY[0] to take effect.
// [1]     enable/disable mult input for post adder
// [2]     +/- (mult-mux output polarity)

    input [3:0] MODEZ,
// MODEZ encoding: 0/1
// [0]     CPI / (CPI >>> 18) (select shift or non-shift CPI)
// [2:1]   Z_INIT/P/Z/CPI (zmux input select)
// [3]     +/- (zmux output polarity)       


    input CLK,

    input RSTX,
    input RSTY,
    input RSTZ,
    input RSTM,
    input RSTP,
    input RSTPRE,
    input RSTMODEX,
    input RSTMODEY,
    input RSTMODEZ,

    input CEX,
    input CEY,
    input CEZ,
    input CEM,
    input CEP,
    input CEPRE,
    input CEMODEX,
    input CEMODEY,
    input CEMODEZ

);

    wire grs;
    assign grs = (GRS_EN == "TRUE") ? !GRS_INST.GRSNET : 1'b0;


// prepare intermediate array  
    wire mode_ce [2:0];
    wire mode_rst [2:0];

    assign mode_ce[0] = CEMODEZ;
    assign mode_ce[1] = CEMODEY;
    assign mode_ce[2] = CEMODEX;

    assign mode_rst[0] = RSTMODEZ;
    assign mode_rst[1] = RSTMODEY;
    assign mode_rst[2] = RSTMODEX;

    wire [1:0] mode_group_idx [7:0]; //lookup table, each MODE register bit belongs to 1 of 3 groups

    assign mode_group_idx[0] = 0;
    assign mode_group_idx[1] = 0;
    assign mode_group_idx[2] = 0;
    assign mode_group_idx[3] = 0;
    assign mode_group_idx[4] = 1;
    assign mode_group_idx[5] = 1;
    assign mode_group_idx[6] = 1;
    assign mode_group_idx[7] = 2;

    genvar i;

    wire [7:0] MODE = {MODEX, MODEY, MODEZ};
    wire [2:0] MODEREG = {MODEX_REG[0], MODEY_REG[0], MODEZ_REG[0]};

    wire [17:0] Xv = X;
    wire [17:0] Yv = Y;
    wire [47:0] Zv = Z;
    wire [7:0] MODEv = MODE;

// registers 

    wire [17:0] X1; // X register (latency == 1)
// X cascade output bus
    localparam XREG_WIDTH = 18;
    localparam XREG_DEPTH = 3;
    wire [XREG_WIDTH-1:0] xreg_d; 
    assign xreg_d = X_SEL ? CXI : Xv;
    assign xreg_rsta = (ASYNC_RST == 1'b1) ? (RSTX | grs) : grs;
    assign xreg_rsts = (ASYNC_RST == 1'b1) ? 1'b0 : RSTX;

    reg [XREG_WIDTH-1:0] xreg_qarr[XREG_DEPTH:0];
    always @(*) begin
        // pragma translate_off
        if (CXO_REG < 0 || CXO_REG > XREG_DEPTH) begin
            $display("ERROR: GTP_APM_E1 instance %m parameter CXO_REG = %d is illegal. The legal values are 0,1,2,3.", CXO_REG);
            $finish;
        end
        // pragma translate_on
        xreg_qarr[0] = xreg_d ;
    end

    integer j;
    always @(posedge CLK or posedge xreg_rsta) begin
        for (j = 1; j <= XREG_DEPTH; j = j + 1) begin
            if (xreg_rsta == 1'b1) begin
                xreg_qarr[j] <= {XREG_WIDTH{1'b0}};
            end else if (xreg_rsts == 1'b1) begin
                xreg_qarr[j] <= {XREG_WIDTH{1'b0}};
            end else if (CEX == 1'b1) begin
                xreg_qarr[j] <= xreg_qarr[j - 1];
            end
        end
    end

    assign CXO = xreg_qarr[CXO_REG];
    assign X1 = xreg_qarr[1];


    wire [17:0] Xi; //registered (optional) X internal bus
    assign Xi = X_REG ? X1 : (X_SEL ? CXI : Xv);

    wire [17:0] Yi; //registered (optional) Y internal
    localparam YREG_WIDTH = 18;
    localparam YREG_DEPTH = 1;
    wire [YREG_WIDTH-1:0] yreg_d; 
    assign yreg_d = Yv;
    assign yreg_rsta = (ASYNC_RST == 1'b1) ? (RSTY | grs) : grs;
    assign yreg_rsts = (ASYNC_RST == 1'b1) ? 1'b0 : RSTY;

    reg [YREG_WIDTH-1:0] yreg_qarr[YREG_DEPTH:0];
    always @(*) begin
        // pragma translate_off
        if (Y_REG < 0 || Y_REG > YREG_DEPTH) begin
            $display("ERROR: GTP_APM_E1 instance %m parameter Y_REG = %d is illegal. The legal value is 0,1.", Y_REG);
            $finish;
        end
        // pragma translate_on
        yreg_qarr[0] = yreg_d ;
    end

    always @(posedge CLK or posedge yreg_rsta) begin
        for (j = 1; j <= YREG_DEPTH; j = j + 1) begin
            if (yreg_rsta == 1'b1) begin
                yreg_qarr[j] <= {YREG_WIDTH{1'b0}};
            end else if (yreg_rsts == 1'b1) begin
                yreg_qarr[j] <= {YREG_WIDTH{1'b0}};
            end else if (CEY == 1'b1) begin
                yreg_qarr[j] <= yreg_qarr[j - 1];
            end
        end
    end

    assign Yi = yreg_qarr[Y_REG];

    wire [47:0] Zi; //registered (optional) Z internal
    localparam ZREG_WIDTH = 48;
    localparam ZREG_DEPTH = 1;
    wire [ZREG_WIDTH-1:0] zreg_d; 
    assign zreg_d = Zv;
    assign zreg_rsta = (ASYNC_RST == 1'b1) ? (RSTZ | grs) : grs;
    assign zreg_rsts = (ASYNC_RST == 1'b1) ? 1'b0 : RSTZ;

    reg [ZREG_WIDTH-1:0] zreg_qarr[ZREG_DEPTH:0];
    always @(*) begin
        // pragma translate_off
        if (Z_REG < 0 || Z_REG > ZREG_DEPTH) begin
            $display("ERROR: GTP_APM_E1 instance %m parameter Z_REG = %d is illegal. The legal value is 0,1.", Z_REG);
            $finish;
        end
        // pragma translate_on
        zreg_qarr[0] = zreg_d ;
    end

    always @(posedge CLK or posedge zreg_rsta) begin
        for (j = 1; j <= ZREG_DEPTH; j = j + 1) begin
            if (zreg_rsta == 1'b1) begin
                zreg_qarr[j] <= {ZREG_WIDTH{1'b0}};
            end else if (zreg_rsts == 1'b1) begin
                zreg_qarr[j] <= {ZREG_WIDTH{1'b0}};
            end else if (CEZ == 1'b1) begin
                zreg_qarr[j] <= zreg_qarr[j - 1];
            end
        end
    end

    assign Zi = zreg_qarr[Z_REG];

    wire [7:0] MODEi; //registered (optional) MODE internal

    generate
    for (i = 0; i < 8; i = i + 1) begin
    localparam MODEREG_WIDTH = 1;
    localparam MODEREG_DEPTH = 1;
    wire [MODEREG_WIDTH-1:0] modereg_d; 
    assign modereg_d = MODEv[i];
    assign modereg_rsta = (ASYNC_RST == 1'b1) ? (mode_rst[mode_group_idx[i]] | grs) : grs;
    assign modereg_rsts = (ASYNC_RST == 1'b1) ? 1'b0 : mode_rst[mode_group_idx[i]];

    reg [MODEREG_WIDTH-1:0] modereg_qarr[MODEREG_DEPTH:0];
    always @(*) begin
        // pragma translate_off
        if (MODEREG[mode_group_idx[i]] < 0 || MODEREG[mode_group_idx[i]] > MODEREG_DEPTH) begin
            $display("ERROR: GTP_APM_E1 instance %m parameter MODE_REG = %d is illegal. The legal value is 0,1.", MODEREG[mode_group_idx[i]]);
            $finish;
        end
        // pragma translate_on
        modereg_qarr[0] = modereg_d ;
    end

    always @(posedge CLK or posedge modereg_rsta) begin
        for (j = 1; j <= MODEREG_DEPTH; j = j + 1) begin
            if (modereg_rsta == 1'b1) begin
                modereg_qarr[j] <= {MODEREG_WIDTH{1'b0}};
            end else if (modereg_rsts == 1'b1) begin
                modereg_qarr[j] <= {MODEREG_WIDTH{1'b0}};
            end else if (mode_ce[mode_group_idx[i]] == 1'b1) begin
                modereg_qarr[j] <= modereg_qarr[j - 1];
            end
        end
    end

    assign MODEi[i] = modereg_qarr[MODEREG[mode_group_idx[i]]];
    end
    endgenerate

// preadder
    wire [17:0] XBr; //registered CXBI
    localparam XBREG_WIDTH = 18;
    localparam XBREG_DEPTH = 1;
    wire [XBREG_WIDTH-1:0] xbreg_d; 
    assign xbreg_d = CXBI;
    assign xbreg_rsta = (ASYNC_RST == 1'b1) ? (RSTZ | grs) : grs;
    assign xbreg_rsts = (ASYNC_RST == 1'b1) ? 1'b0 : RSTZ;

    reg [XBREG_WIDTH-1:0] xbreg_qarr[XBREG_DEPTH:0];
    always @(*) begin
        xbreg_qarr[0] = xbreg_d ;
    end

    always @(posedge CLK or posedge xbreg_rsta) begin
        for (j = 1; j <= XBREG_DEPTH; j = j + 1) begin
            if (xbreg_rsta == 1'b1) begin
                xbreg_qarr[j] <= {XBREG_WIDTH{1'b0}};
            end else if (xbreg_rsts == 1'b1) begin
                xbreg_qarr[j] <= {XBREG_WIDTH{1'b0}};
            end else if (CEZ == 1'b1) begin
                xbreg_qarr[j] <= xbreg_qarr[j - 1];
            end
        end
    end

    assign XBr = xbreg_qarr[1];

    reg [17:0] XBi;
    always @(*) begin
        case (XB_SEL)
            2'b00 : XBi = Zi[47:30];
            2'b01 : XBi = CXBI;
            2'b10 : XBi = XBr;
            2'b11 : XBi = CXO;
        endcase
    end
    assign CXBO = XBi;

    //
    // PRE add/sub with SIMD feature
    //
    wire [17:0] PREc; //combinational preadder output
    localparam PREADD_WIDTH = 18;
    wire preadd_sub;
    wire [PREADD_WIDTH-1:0] preadd_S;
    wire [PREADD_WIDTH/2-1:0] preadd_A_hi, preadd_A_lo;
    wire [PREADD_WIDTH/2-1:0] preadd_B_hi, preadd_B_lo;
    wire [PREADD_WIDTH/2-1:0] preadd_S_hi, preadd_S_lo;
    assign preadd_sub = MODEi[7];
    assign preadd_A_hi = Xi[PREADD_WIDTH - 1 : PREADD_WIDTH/2];
    assign preadd_B_hi = XBi[PREADD_WIDTH - 1 : PREADD_WIDTH/2];
    assign preadd_A_lo = Xi[PREADD_WIDTH/2 - 1 : 0];
    assign preadd_B_lo = XBi[PREADD_WIDTH/2 - 1 : 0];
    // 18-bit addsub
    assign preadd_S = preadd_sub ? Xi - XBi : Xi + XBi;
    // dual 9-bit addsub
    assign preadd_S_hi = preadd_sub ? preadd_A_hi - preadd_B_hi : preadd_A_hi + preadd_B_hi;
    assign preadd_S_lo = preadd_sub ? preadd_A_lo - preadd_B_lo : preadd_A_lo + preadd_B_lo;
    //
    assign PREc = (USE_SIMD == 1'b1)? {preadd_S_hi, preadd_S_lo} : preadd_S;

    wire [17:0] PREi; //registered (optional) preadder output
    localparam PREREG_WIDTH = 18;
    localparam PREREG_DEPTH = 1;
    wire [PREREG_WIDTH-1:0] prereg_d; 
    assign prereg_d = PREc;
    assign prereg_rsta = (ASYNC_RST == 1'b1) ? (RSTPRE | grs) : grs;
    assign prereg_rsts = (ASYNC_RST == 1'b1) ? 1'b0 : RSTPRE;

    reg [PREREG_WIDTH-1:0] prereg_qarr[PREREG_DEPTH:0];
    always @(*) begin
        // pragma translate_off
        if (PREADD_REG < 0 || PREADD_REG > PREREG_DEPTH) begin
            $display("ERROR: GTP_APM_E1 instance %m parameter PREADD_REG = %d is illegal. The legal value is 0,1.", PREADD_REG);
            $finish;
        end
        // pragma translate_on
        prereg_qarr[0] = prereg_d ;
    end

    always @(posedge CLK or posedge prereg_rsta) begin
        for (j = 1; j <= PREREG_DEPTH; j = j + 1) begin
            if (prereg_rsta == 1'b1) begin
                prereg_qarr[j] <= {PREREG_WIDTH{1'b0}};
            end else if (prereg_rsts == 1'b1) begin
                prereg_qarr[j] <= {PREREG_WIDTH{1'b0}};
            end else if (CEPRE == 1'b1) begin
                prereg_qarr[j] <= prereg_qarr[j - 1];
            end
        end
    end

    assign PREi = prereg_qarr[PREADD_REG];

// multiplier
    wire [47:0] Mc; //mult combinational output
    wire [17:0] mult_x;
    wire [17:0] mult_y;
    assign mult_x = USE_PREADD ? PREi : Xi;
    assign mult_y = Yi;
    localparam MULT_IWIDTH = 18;
    localparam MULT_OWIDTH = 48;
    wire [MULT_OWIDTH-1:0] mult_p0;
    wire [MULT_OWIDTH-1:0] mult_p1;
    // mult18
    wire multp0_sign_x;
    wire multp0_sign_y;
    assign multp0_sign_x = X_SIGNED ? mult_x[MULT_IWIDTH-1] : 1'b0;
    assign multp0_sign_y = Y_SIGNED ? mult_y[MULT_IWIDTH-1] : 1'b0;
    wire [MULT_OWIDTH-1:0] multp0_Xi;
    wire [MULT_OWIDTH-1:0] multp0_Yi;
    assign multp0_Xi = {{(MULT_OWIDTH-MULT_IWIDTH){multp0_sign_x}},mult_x};
    assign multp0_Yi = {{(MULT_OWIDTH-MULT_IWIDTH){multp0_sign_y}},mult_y};
    assign mult_p0 = multp0_Xi * multp0_Yi;
    //mult9_0
    wire multp1_0_sign_x;
    wire multp1_0_sign_y;
    assign multp1_0_sign_x = X_SIGNED ? mult_x[MULT_IWIDTH/2-1] : 1'b0;
    //assign multp1_0_sign_y = Y_SIGNED ? mult_y[MULT_IWIDTH/2-1] : 1'b0;
    assign multp1_0_sign_y = Y_SIGNED ? mult_y[8] : 1'b0;
    wire [MULT_OWIDTH/2-1:0] multp1_0_Xi;
    wire [MULT_OWIDTH/2-1:0] multp1_0_Yi;
    assign multp1_0_Xi = {{(MULT_OWIDTH/2-MULT_IWIDTH/2){multp1_0_sign_x}},mult_x[MULT_IWIDTH/2-1:0]};
    assign multp1_0_Yi = {{(MULT_OWIDTH/2-MULT_IWIDTH/2){multp1_0_sign_y}},mult_y[MULT_IWIDTH/2-1:0]};
    assign mult_p1[MULT_OWIDTH/2-1:0] = multp1_0_Xi * multp1_0_Yi;
    //mult9_1
    wire multp1_1_sign_x;
    wire multp1_1_sign_y;
    assign multp1_1_sign_x = X_SIGNED ? mult_x[MULT_IWIDTH-1] : 1'b0;
    assign multp1_1_sign_y = Y_SIGNED ? mult_y[MULT_IWIDTH-1] : 1'b0;
    wire [MULT_OWIDTH-1:MULT_OWIDTH/2] multp1_1_Xi;
    wire [MULT_OWIDTH-1:MULT_OWIDTH/2] multp1_1_Yi;
    assign multp1_1_Xi = {{(MULT_OWIDTH/2-MULT_IWIDTH/2){multp1_1_sign_x}},mult_x[MULT_IWIDTH-1:MULT_IWIDTH/2]};
    assign multp1_1_Yi = {{(MULT_OWIDTH/2-MULT_IWIDTH/2){multp1_1_sign_y}},mult_y[MULT_IWIDTH-1:MULT_IWIDTH/2]};
    assign mult_p1[MULT_OWIDTH-1:MULT_OWIDTH/2] = multp1_1_Xi * multp1_1_Yi;

    assign Mc = (USE_SIMD == 1'b1) ? mult_p1 : mult_p0;

    wire [47:0] Mi; //registered (optional) mult internal output
    localparam MREG_WIDTH = 48;
    localparam MREG_DEPTH = 1;
    wire [MREG_WIDTH-1:0] mreg_d; 
    assign mreg_d = Mc;
    assign mreg_rsta = (ASYNC_RST == 1'b1) ? (RSTM | grs) : grs;
    assign mreg_rsts = (ASYNC_RST == 1'b1) ? 1'b0 : RSTM;

    reg [MREG_WIDTH-1:0] mreg_qarr[MREG_DEPTH:0];
    always @(*) begin
        // pragma translate_off
        if (MULT_REG < 0 || MULT_REG > MREG_DEPTH) begin
            $display("ERROR: GTP_APM_E1 instance %m parameter MULT_REG = %d is illegal. The legal value is 0,1.", MULT_REG);
            $finish;
        end
        // pragma translate_on
        mreg_qarr[0] = mreg_d ;
    end

    always @(posedge CLK or posedge mreg_rsta) begin
        for (j = 1; j <= MREG_DEPTH; j = j + 1) begin
            if (mreg_rsta == 1'b1) begin
                mreg_qarr[j] <= {MREG_WIDTH{1'b0}};
            end else if (mreg_rsts == 1'b1) begin
                mreg_qarr[j] <= {MREG_WIDTH{1'b0}};
            end else if (CEM == 1'b1) begin
                mreg_qarr[j] <= mreg_qarr[j - 1];
            end
        end
    end

    assign Mi = mreg_qarr[MULT_REG];

// post adder 
    reg  [47:0] Pai; // post adder input a before inverter
    wire [47:0] Pa = MODEi[6] ? ~Pai : Pai; // post adder input a after inverter
    reg  [47:0] Pbi; // post adder input b before inverter
    wire [47:0] Pb = MODEi[3] ? ~Pbi : Pbi; // post adder input b after inverter

    wire [47:0] Pc; // post adder combinational output
    wire [47:0] Pr; // post adder regstered feedback
    wire [47:0] Pri =  USE_ACCLOW ? { {30{1'b0}}, Pr[17:0] } : Pr; //post adder lower portion feedback

    always @ (*) begin
        case(MODEi[5])
            1'b0 : Pai = Mi;
            1'b1 : Pai = Pri & {48{MODEi[4]}};
        endcase
    end

    always @(*) begin
        case(MODEi[2:1])
            2'b00 : Pbi = Z_INIT;
            2'b01 : Pbi = Pri;
            2'b10 : Pbi = Zi;
            2'b11 : Pbi = MODEi[0] ? ($signed(CPI) >>> 18) : $signed(CPI); //both branch need $signed
        endcase
    end

    //
    // adder with SIMD feature
    //
    localparam ADD48_WIDTH = 48;
    wire add48_CO, add48_CI;
    wire [ADD48_WIDTH-1:0] add48_S;
    wire [ADD48_WIDTH/2-1:0] add48_A_hi, add48_A_lo;
    wire [ADD48_WIDTH/2-1:0] add48_B_hi, add48_B_lo;
    wire [ADD48_WIDTH/2-1:0] add48_S_hi, add48_S_lo;
    assign add48_CI = CIN_SEL ? CIN : (MODEi[6] | MODEi[3]);
    assign add48_A_hi = Pa[ADD48_WIDTH - 1 : ADD48_WIDTH/2];
    assign add48_B_hi = Pb[ADD48_WIDTH - 1 : ADD48_WIDTH/2];
    assign add48_A_lo = Pa[ADD48_WIDTH/2 - 1 : 0];
    assign add48_B_lo = Pb[ADD48_WIDTH/2 - 1 : 0];
    // 48-bit adder
    assign {add48_CO, add48_S} = Pa + Pb + add48_CI;
    // dual 24-bit adders with identical CI
    assign add48_S_hi = add48_A_hi + add48_B_hi + add48_CI;
    assign add48_S_lo = add48_A_lo + add48_B_lo + add48_CI;
    //
    assign Pc = (USE_SIMD == 1'b1) ? {add48_S_hi, add48_S_lo} : add48_S;

    wire [47:0] Pi;
    localparam PREG_WIDTH = 48;
    localparam PREG_DEPTH = 1;
    wire [PREG_WIDTH-1:0] preg_d; 
    assign preg_d = Pc;
    assign preg_rsta = (ASYNC_RST == 1'b1) ? (RSTP | grs) : grs;
    assign preg_rsts = (ASYNC_RST == 1'b1) ? 1'b0 : RSTP;

    reg [PREG_WIDTH-1:0] preg_qarr[PREG_DEPTH:0];
    always @(*) begin
        // pragma translate_off
        if (P_REG < 0 || P_REG > PREG_DEPTH) begin
            $display("ERROR: GTP_APM_E1 instance %m parameter P_REG = %d is illegal. The legal value is 0,1.", P_REG);
            $finish;
        end
        // pragma translate_on
        preg_qarr[0] = preg_d ;
    end

    always @(posedge CLK or posedge preg_rsta) begin
        for (j = 1; j <= PREG_DEPTH; j = j + 1) begin
            if (preg_rsta == 1'b1) begin
                preg_qarr[j] <= {PREG_WIDTH{1'b0}};
            end else if (preg_rsts == 1'b1) begin
                preg_qarr[j] <= {PREG_WIDTH{1'b0}};
            end else if (CEP == 1'b1) begin
                preg_qarr[j] <= preg_qarr[j - 1];
            end
        end
    end

    assign Pi = preg_qarr[P_REG];
    assign Pr = preg_qarr[1];

    assign P = USE_POSTADD ? Pi : Mi;
    assign CPO = USE_POSTADD? (CPO_REG ? Pr : Pc) : Mi;

    wire PCOr;
    localparam PCOREG_WIDTH = 1;
    localparam PCOREG_DEPTH = 1;
    wire [PCOREG_WIDTH-1:0] pcoreg_d; 
    assign pcoreg_d = add48_CO;
    assign pcoreg_rsta = (ASYNC_RST == 1'b1) ? (RSTP | grs) : grs;
    assign pcoreg_rsts = (ASYNC_RST == 1'b1) ? 1'b0 : RSTP;

    reg [PCOREG_WIDTH-1:0] pcoreg_qarr[PCOREG_DEPTH:0];
    always @(*) begin
        pcoreg_qarr[0] = pcoreg_d ;
    end

    always @(posedge CLK or posedge pcoreg_rsta) begin
        for (j = 1; j <= PCOREG_DEPTH; j = j + 1) begin
            if (pcoreg_rsta == 1'b1) begin
                pcoreg_qarr[j] <= {PCOREG_WIDTH{1'b0}};
            end else if (pcoreg_rsts == 1'b1) begin
                pcoreg_qarr[j] <= {PCOREG_WIDTH{1'b0}};
            end else if (CEP == 1'b1) begin
                pcoreg_qarr[j] <= pcoreg_qarr[j - 1];
            end
        end
    end

    assign PCOr = pcoreg_qarr[1];
    assign COUT = CPO_REG ? PCOr : add48_CO;

// DRC check
// pragma translate_off
    initial begin
        `assert(X_REG <= 1, "X_REG <= 1")
        `assert(XB_SEL != 3 || CXO_REG >=  X_REG, "X_REG <= CXO_REG in back-propogation mode")
        `assert(CXO_REG <= 3, "CXO_REG <= 3")
        `assert(Y_REG <= 1, "Y_REG <= 1")
        `assert(Z_REG <= 1, "Z_REG <= 1")
        `assert(MULT_REG <= 1, "MULT_REG <= 1")
        `assert(P_REG <= 1, "P_REG <= 1")
        `assert(PREADD_REG <= 1, "PREADD_REG <= 1")
        `assert(MODEX_REG <= 1, "MODEX_REG <= 1")
        `assert(MODEY_REG <= 1, "MODEY_REG <= 1")
        `assert(MODEZ_REG <= 1, "MODEZ_REG <= 1")
    end
// pragma translate_on

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2016 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_CLKBUFM.v
//
// Functional description: CLOCK BUFFER
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_CLKBUFM
(
    output CLKOUT,
    input CLKIN
);

//synthesis translate_off

    assign CLKOUT = CLKIN;

//synthesis translate_on
endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_RAM32X2SP.v
//
// Functional description: single-port 32x2 distributed ram
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_RAM32X2SP
#(
    parameter [31:0] INIT_0 = 32'h00000000 ,
    parameter [31:0] INIT_1 = 32'h00000000
) (
    output [1:0] DO,
    input  [1:0] DI,
    input [4:0] ADDR,
    input WCLK, WE
);

    reg [31:0] mem [1:0];

    initial begin
        mem[0] = INIT_0;
        mem[1] = INIT_1;
    end

    always @(posedge WCLK) begin
        if (WE == 1'b1) begin
            mem[0][ADDR] <= DI[0];
            mem[1][ADDR] <= DI[1];
        end
    end

    assign DO[0] = mem[0][ADDR];
    assign DO[1] = mem[1][ADDR];

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_SPI.v
//
// Functional description: SPI Circuit
//
// Parameter description:
//      
//
// Port description:
//      
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////


`timescale 1 ns / 1 ps
module GTP_SPI
(
output        SCK_OE_N,
input         SCK_I,
output        SCK_O,
output  [7:0] SS_O_N,
input         SS_I_N,
output        MISO_OE_N,
input         MISO_I,
output        MISO_O,
output        MOSI_OE_N,
input         MOSI_I,
output        MOSI_O,
output        IRQ
);

assign  GTP_GRS.spi_sck_i    = SCK_I;
assign  GTP_GRS.spi_ss_i_n   = SS_I_N;
assign  GTP_GRS.spi_miso_i   = MISO_I;
assign  GTP_GRS.spi_mosi_i   = MOSI_I;
assign  SS_O_N = GTP_GRS.spi_ss_o_n    ;
assign  SCK_OE_N = GTP_GRS.spi_sck_oe_n  ;
assign  SCK_O = GTP_GRS.spi_sck_o     ;
assign  MOSI_OE_N = GTP_GRS.spi_mosi_oe_n ;
assign  MOSI_O = GTP_GRS.spi_mosi_o    ;
assign  MISO_OE_N = GTP_GRS.spi_miso_oe_n ;
assign  MISO_O = GTP_GRS.spi_miso_o    ;
assign  IRQ = GTP_GRS.irq_spi       ;

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_PREADD_MULTADDACC9.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

//P = MAC + (A0*(B0+C0) + A1*(B1+C1))
`timescale 1 ns / 1 ps

module GTP_PREADD_MULTADDACC9 #(
    parameter GRS_EN            = "TRUE", //"TRUE"; "FALSE"
    parameter SYNC_RST          = "FALSE", //"TRUE"; "FALSE"
    parameter INREG_EN          = "FALSE",  //"TRUE"; "FALSE"
    parameter PREREG_EN         = "FALSE",  //"TRUE"; "FALSE"
    parameter PIPEREG_EN        = "FALSE",//"TRUE"; "FALSE"
    parameter ADDSUB_OP         = 0 ,
    parameter ACC_ADDSUB_OP     = 0,
    parameter DYN_ADDSUB_OP     = 1,
    parameter DYN_ACC_ADDSUB_OP = 1,
    parameter OVERFLOW_MASK     = 32'h0,  //PSIZE = 32 OVERflow setting = 'h1_0000_0000 , bit width = PSIZE
    parameter PATTERN           = 32'h0,  //compare pattern
    parameter MASKPAT           = 32'h0,  //pattern mask
    parameter ACC_INIT_VALUE    = 32'h0   //ACC_INIT_VALUE value
) (
    output  [31:0] P,
    output  OVER,
    output  UNDER,
    output  EQZ,
    output  EQZM,
    output  EQOM,
    output  EQPAT,
    output  EQPATN,

    input   CE,
    input   RST,
    input   CLK,
    input   A_SIGNED,
    input   [8:0] A0,
    input   [8:0] A1,
    input   B_SIGNED,
    input   [7:0] B0,
    input   [7:0] B1,
    input   C_SIGNED,
    input   [7:0] C0,
    input   [7:0] C1,
    input   [1:0] PREADDSUB,
    input   ADDSUB,
    input   ACC_ADDSUB,
    input   RELOAD
);

    wire [31:0] R;

    INT_PREADD_MULTADDACC #(
        . GRS_EN(GRS_EN),      
        . SYNC_RST(SYNC_RST),    
        . INREG_EN(INREG_EN),    
        . PREREG_EN(PREREG_EN),    
        . PIPEREG_EN(PIPEREG_EN),  
        . ADDSUB_OP(ADDSUB_OP),     
        . ACCUMADDSUB_OP(ACC_ADDSUB_OP),
        . DYN_OP_ADDSUB(DYN_ADDSUB_OP),   
        . DYN_OP_ACC(DYN_ACC_ADDSUB_OP),   
        . ASIZE(9),
        . BSIZE(8),
        . PSIZE(32),
        . DYN_ACC_INIT(0),
        . ACC_INIT_VALUE(ACC_INIT_VALUE),
        . MASK(OVERFLOW_MASK)
    ) U_MACC (
        . CE(CE),
        . RST(RST),
        . CLK(CLK),
        . A_SIGNED(A_SIGNED),
        . A0(A0),
        . A1(A1),
        . B_SIGNED(B_SIGNED),
        . B0(B0),
        . B1(B1),
        . C_SIGNED(C_SIGNED),
        . C0(C0),
        . C1(C1),
        . PREADDSUB(PREADDSUB),
        . ACCUM_INIT(32'b0),
        . ADDSUB(ADDSUB),
        . ACCUMADDSUB(ACC_ADDSUB),
        . RELOAD(RELOAD),
        . P(P),
        . OVER(OVER),
        . UNDER(UNDER),
        . R(R) 
    );     

    INT_FLAG #(
        . GRS_EN(GRS_EN),
        . SYNC_RST(SYNC_RST),
        . PSIZE(32),
        . PATSIZE(32),
        . MASKPATSIZE(32),
        . OUTREG_EN("TRUE")
    ) U_FLAG (
        . CE(CE),
        . RST(RST),
        . CLK(CLK),
        . P(P),
        . PATTERN(PATTERN),
        . MASKPAT(MASKPAT),
        . OVERFLOW_MASK(OVERFLOW_MASK),
        . R(R),
        . eqz(EQZ),
        . eqzm(EQZM),
        . eqom(EQOM),
        . eqpat(EQPAT),
        . eqpatn(EQPATN)
    );

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_IOBUFECO.v
//
// Functional description: Differential Signaling Input/Output Buffer
//
// Parameter description:
//
// Port description:
//
// Revision:
//    06/18/14 - Initial version.
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_IOBUFECO #(
    parameter IOSTANDARD = "DEFAULT",
    parameter TERM_DDR = "ON"
)(
    output reg O,
    inout IO,
    inout IOB,
    input I,
    input EN,                    // 1: enable inbuf, normal mode; 0: disable inbuf, standby mode.
    input T
) /* synthesis syn_black_box */ ;
  
  initial begin
    case (IOSTANDARD)
    "SSTL18D_I", "SSTL18D_II", "SSTL15D_I", "SSTL15D_II", "HSTL15D_I", "SSTL25D_I", "SSTL25D_II", "SSTL15D_I_CAL", "SSTL15D_II_CAL", "HSTL15D_I_CAL", "LVPECL", "RSDS", "PPDS", "BLVDS", "LVCMOS25D", "LVCMOS33D","LVDS25E", "DEFAULT":;
    default : begin
           $display("Attribute Syntax Error : The attribute IOSTANDARD on GTP_IOBUFECO instance %m is set to %s.", IOSTANDARD);
           $finish;
              end
    endcase

    case (TERM_DDR)
    "ON", "OFF" :;
    default : begin
           $display("Attribute Syntax Error : The attribute TERM_DDR on GTP_IOBUFECO instance %m is set to %s.", TERM_DDR);
           $finish;
              end
    endcase
    end 
    bufif0 (IO, I, T);
    notif0 (IOB, I, T);

  always @(*)
    begin
      if (EN == 1'b1)
        begin
        if (IO == 1'b1 && IOB == 1'b0)
            O = IO;
        else if (IO == 1'b0 && IOB == 1'b1)
            O = IO;
        else
            O = 1'bx;
        end
     else
            O = 1'b1;
    end

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_CLKBUFR.v
//
// Functional description: Regional Clock Buffer
//
// Parameter description:
//
// Port description:
//
// Revision:
//    06/30/16 - Initial version.
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_CLKBUFR
(
    output CLKOUT,
    input CLKIN
);

    assign CLKOUT = CLKIN;

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_IOBUF_RX_MIPI.v
//
// Functional description: Input Buffer For MIPI Protocol
//
// Parameter description:
//
// Port description:
//
// Revision:
//    05/18/18 - Initial version.
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_IOBUF_RX_MIPI 
#(
  parameter IOSTANDARD  ="DEFAULT",
  parameter SLEW_RATE = "SLOW",
  parameter DRIVE_STRENGTH = "6",
  parameter TERM_DIFF = "ON"
) (
    output wire O_LP,
    output wire OB_LP,
    output reg  O_HS,
    inout  wire IO,
    inout  wire IOB,
    input  wire I_LP,
    input  wire IB_LP,
    input  wire T,
    input  wire TB,
    input  wire M
);

    reg [23:0]  STR_I, STR_IB;
    
    always @(*)
      begin
         $sformat(STR_I, "%v", IO);
         $sformat(STR_IB, "%v", IOB);
      end

    initial   begin
         case(IOSTANDARD) 
           "MIPI", "DEFAULT" : ;
           default:  begin
             $display("Attribute ERROR: Illegal IOSTANDARD value %s.", IOSTANDARD);
             $finish;
             end
         endcase

    case (TERM_DIFF)
    "ON", "OFF" :;
    default : begin
           $display("Attribute Syntax Error : The attribute TERM_DIFF on instance %m is set to %s.", TERM_DIFF);
           $finish;
              end
    endcase

    case (SLEW_RATE)
    "FAST", "SLOW":;
    default : begin
           $display("Attribute Syntax Error : The attribute SLEW_RATE on instance %m is set to %s.", SLEW_RATE);
           $finish;
              end
    endcase

    case (DRIVE_STRENGTH)
    "2", "4", "6" :;
    default : begin
           $display("Attribute Syntax Error : The attribute DRIVE_STRENGTH on GTP_IOBUF_RX_MIPI instance %m is set to %s.", DRIVE_STRENGTH);
           $finish;
              end
    endcase

     end

// low power input

    assign O_LP  = (T == 1'b0) ? 1'b1 : 
                   (T == 1'b1) ? ((STR_I[23:16] == "S" && STR_IB[23:16] == "S") ? IO : 1'b0)
                               : 1'bx;
    assign OB_LP = (TB == 1'b0) ? IOB : 
                   (TB == 1'b1) ? ((STR_I[23:16] == "S" && STR_IB[23:16] == "S") ? IOB : 1'b0)
                               : 1'bx;

// low power output

    assign T_LP = M || T;
    assign TB_LP = M || TB;
 
    bufif0 (IO, I_LP, T_LP);
    bufif0 (IOB, IB_LP, TB_LP);

    always @(*)
    begin
// high speed input 
        if(M == 1)
        begin
           if (IO == 1'b1 && IOB == 1'b0)
             begin
               O_HS = 1'b1;
             end
           else if (IO == 1'b0 && IOB == 1'b1)
             begin
               O_HS = 0;
             end
           else
             begin
              O_HS = 1'bx;
             end
        end
// low power mode
        else if(M == 0) 
        begin
           O_HS = 1'b1;
        end           
    end
    
endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_ISERDES.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//2017/12/21 : initial version
//2018/01/02 : update dut to software feedback
//2018/04/09 : change SYNC_RS to RS_TYPE
//2018/04/24 : change default value of GRS_N to "TRUE"
/////////////////////////////////////////////////////////////////////////////
module GTP_IDDR #(
parameter RS_TYPE  = "ASYNC_SET",     //"ASYNC_SET", "ASYNC_RESET", "SYNC_SET", "SYNC_RESET"
parameter GRS_EN    = "TRUE"         //"FALSE", "TRUE"
) (
output Q0,
output Q1,
input D,
input CE,
input RS,
input CLK
); /* synthesis syn_black_box */

//synthesis translate_off

reg ce_reg;
reg q_reg0;
reg q_reg1;
reg q_reg2;
reg q_reg3;

wire global_rsn;
wire global_rstn;
wire global_setn;
wire local_rst_async;
wire local_set_async; 
wire local_rst_sync;
wire local_set_sync; 
wire rstn_async;
wire setn_async;
wire rstn_sync;
wire setn_sync;
wire clk_gated;

initial begin
    if(GRS_EN != "TRUE" && GRS_EN != "FALSE")
    begin
      $display("GTP_IDDR Error: Illegal setting of GRS_EN %s",GRS_EN);
      $finish;
    end
    if(RS_TYPE != "ASYNC_SET" && RS_TYPE != "ASYNC_RESET" && RS_TYPE != "SYNC_SET" && RS_TYPE != "SYNC_RESET")
    begin
      $display("GTP_IDDR Error: Illegal setting of RS_TYPE %s",RS_TYPE);
      $finish;
    end

    ce_reg = 1'b0;
    q_reg0 = 1'b0;
    q_reg1 = 1'b0;
    q_reg2 = 1'b0;
    q_reg3 = 1'b0;
end

//////////////////////////////////////////////////////////////////////
assign global_rsn  = (GRS_EN == "TRUE")    ? GRS_INST.GRSNET : 1'b1;

assign global_rstn = (RS_TYPE == "SYNC_SET" || RS_TYPE == "ASYNC_SET")   ? 1'b1 : global_rsn;
assign global_setn = (RS_TYPE == "SYNC_RESET" || RS_TYPE == "ASYNC_RESET") ? 1'b1 : global_rsn;


assign local_rst_async = (RS_TYPE == "ASYNC_RESET") ? RS : 1'b0;
assign local_set_async = (RS_TYPE == "ASYNC_SET")   ? RS : 1'b0;

assign local_rst_sync  = (RS_TYPE == "ASYNC_RESET" || RS_TYPE == "SYNC_RESET") ? RS : 1'b0;
assign local_set_sync  = (RS_TYPE == "ASYNC_SET" || RS_TYPE == "SYNC_SET")     ? RS : 1'b0;


assign rstn_async = global_rstn&(~local_rst_async);
assign setn_async = global_setn&(~local_set_async);

assign rstn_sync  = global_rstn&(~local_rst_sync);
assign setn_sync  = global_setn&(~local_set_sync);


always @(negedge CLK or negedge global_rsn)
begin
    if(!global_rsn)
        ce_reg <= 1'b0;
    else
        ce_reg <= CE;
end

assign clk_gated = ce_reg&CLK;

always @(negedge clk_gated or negedge setn_async or negedge rstn_async)
begin
    if(!(rstn_async&rstn_sync))
        q_reg0 <= 1'b0;
    else if(!(setn_async&setn_sync))
        q_reg0 <= 1'b1;
    else
        q_reg0 <= D;
end

always @(posedge clk_gated or negedge setn_async or negedge rstn_async)
begin
    if(!(rstn_async&rstn_sync))
        q_reg1 <= 1'b0;
    else if(!(setn_async&setn_sync))
        q_reg1 <= 1'b1;    
    else
        q_reg1 <= q_reg0;
end

always @(posedge clk_gated or negedge setn_async or negedge rstn_async)
begin
    if(!(rstn_async&rstn_sync))
        q_reg2 <= 1'b0;
    else if(!(setn_async&setn_sync))
        q_reg2 <= 1'b1;
    else
        q_reg2 <= D; 
end 

always @(posedge clk_gated or negedge setn_async or negedge rstn_async)
begin
    if(!(rstn_async&rstn_sync))
        q_reg3 <= 1'b0;
    else if(!(setn_async&setn_sync))
        q_reg3 <= 1'b1;
    else
        q_reg3 <= q_reg2; 
end 

assign Q1 = q_reg1;
assign Q0 = q_reg3;

//synthesis translate_on
endmodule




































//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_IMDES4.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_IMDES4 #(
parameter GRS_EN = "TRUE", //"TRUE"; "FALSE"
parameter LRS_EN = "TRUE",  //"TRUE"; "FALSE"
parameter DPI_EN = "FALSE"  //"TRUE"; "FALSE"
)(
output  [3:0] Q,
output [1:0] DPI_STS,
input [1:0] DPI_CTRL,
input DPI_STS_CLR_N, 
input PADI,
input ICLK,
input DESCLK,
input RCLK,
input [2:0] IFIFO_WADDR,
input [2:0] IFIFO_RADDR,
input RST
);

//synthesis translate_off


wire [7:0] PADI_D;
reg DPI_P;
reg [1:0] DPI_STS_R;
reg DPI_N_reg;
wire COMP_BEFORE;
wire COMP_AFTER;
wire COMP_BEFORE_D;
wire COMP_AFTER_D;
wire PD_BEFORE;
wire PD_AFTER;
wire DPI_BEFORE_POS_REG_T;
wire DPI_AFTER_POS_REG_T;
wire DPI_BEFORE_NEG_REG_T;
wire DPI_AFTER_NEG_REG_T;
wire AFTER_POS;
wire BEFORE_POS;
wire AFTER_NEG;
wire BEFORE_NEG;
reg DPI_BEFORE;
reg DPI_AFTER;
reg DPI_BEFORE_POS_REG;
reg DPI_BEFORE_NEG_REG;
reg DPI_AFTER_POS_REG;
reg DPI_AFTER_NEG_REG;
reg [7:0] PADI_POS_fifo;
reg [7:0] PADI_NEG_fifo;
reg [3:0] Q_reg;
reg [3:0] shift_reg;
reg capture_en_b;
reg capture_en;
reg [3:0] capture_reg;

initial begin
DPI_P      = 0;
DPI_STS_R  = 0;
DPI_N_reg  = 0;
DPI_BEFORE = 0;
DPI_AFTER  = 0;
DPI_BEFORE_POS_REG = 0;
DPI_BEFORE_NEG_REG = 0;
DPI_AFTER_POS_REG  = 0;
DPI_AFTER_NEG_REG  = 0;
PADI_POS_fifo = 0;
PADI_NEG_fifo = 0;
Q_reg = 0;
shift_reg= 0;
capture_en_b = 0;
capture_en   = 0;
capture_reg  = 0;
end
assign global_rstn = (GRS_EN == "TRUE") ? GRS_INST.GRSNET : 1'b1;
assign lsr_rstn = LRS_EN == "TRUE" ? (~RST) : 1'b1;

assign  #0.05 PADI_D[0] =  PADI;
assign  #0.05 PADI_D[1] =  PADI_D[0];
assign  #0.05 PADI_D[2] =  PADI_D[1];
assign  #0.05 PADI_D[3] =  PADI_D[2];
assign  #0.05 PADI_D[4] =  PADI_D[3];
assign  #0.05 PADI_D[5] =  PADI_D[4];
assign  #0.05 PADI_D[6] =  PADI_D[5];
assign  #0.05 PADI_D[7] =  PADI_D[6];

assign PADI_SAMPLE = (DPI_EN == "TRUE") ? PADI_D[3] : PADI;

always @(posedge ICLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_P <= 0;
   else if (!lsr_rstn)
      DPI_P <= 0;
   else
      DPI_P <= PADI_SAMPLE;
end

always @(negedge ICLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_N_reg <= 0;
   else if (!lsr_rstn)
      DPI_N_reg <= 0;
   else 
      DPI_N_reg <= PADI_SAMPLE;
end

always @(*) begin
   case (DPI_CTRL[1:0])
      2'd0:    begin DPI_BEFORE = PADI_D[2];  DPI_AFTER = PADI_D[4]; end
      2'd1:    begin DPI_BEFORE = PADI_D[1];  DPI_AFTER = PADI_D[5]; end
      2'd2:    begin DPI_BEFORE = PADI_D[0];  DPI_AFTER = PADI_D[6]; end
      default: begin DPI_BEFORE = PADI;       DPI_AFTER = PADI_D[7]; end
   endcase
end

always @(posedge ICLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_BEFORE_POS_REG <= 0;
   else if (!lsr_rstn)
      DPI_BEFORE_POS_REG <= 0;
   else   
      DPI_BEFORE_POS_REG <= DPI_BEFORE;
end

always @(negedge ICLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_BEFORE_NEG_REG <= 0;
   else if (!lsr_rstn)
      DPI_BEFORE_NEG_REG <= 0;
   else     
      DPI_BEFORE_NEG_REG <= DPI_BEFORE;
end


always @(posedge ICLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_AFTER_POS_REG <= 0;
   else if (!lsr_rstn)
      DPI_AFTER_POS_REG <= 0;
   else   
      DPI_AFTER_POS_REG <= DPI_AFTER;
end


always @(negedge ICLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_AFTER_NEG_REG <= 0;
   else if (!lsr_rstn)
      DPI_AFTER_NEG_REG <= 0;
   else     
      DPI_AFTER_NEG_REG <= DPI_AFTER;
end


assign BEFORE_POS = DPI_BEFORE_POS_REG_T ^ DPI_P;
assign DPI_BEFORE_POS_REG_T = (DPI_EN == "TRUE") ? DPI_BEFORE_POS_REG : 0;

assign AFTER_POS = DPI_AFTER_POS_REG_T ^ DPI_P;
assign DPI_AFTER_POS_REG_T = (DPI_EN == "TRUE") ? DPI_AFTER_POS_REG : 0;

assign BEFORE_NEG = DPI_BEFORE_NEG_REG_T ^ DPI_N_reg;
assign DPI_BEFORE_NEG_REG_T = (DPI_EN == "TRUE") ? DPI_BEFORE_NEG_REG : 0;

assign AFTER_NEG = DPI_AFTER_NEG_REG_T ^ DPI_N_reg;
assign DPI_AFTER_NEG_REG_T = (DPI_EN == "TRUE") ? DPI_AFTER_NEG_REG : 0;


assign COMP_BEFORE = BEFORE_POS || BEFORE_NEG;
assign COMP_AFTER = AFTER_POS || AFTER_NEG;

assign #0.1 COMP_BEFORE_D = COMP_BEFORE;
assign #0.1 COMP_AFTER_D = COMP_AFTER;

assign PD_BEFORE = COMP_BEFORE && COMP_BEFORE_D;
assign PD_AFTER = COMP_AFTER && COMP_AFTER_D;


always @(posedge DPI_STS_CLR_N or negedge global_rstn or negedge lsr_rstn or posedge PD_BEFORE) begin
   if (!global_rstn)
      DPI_STS_R[0] <= 0;
   else if (!lsr_rstn)
      DPI_STS_R[0] <= 0;
   else if (PD_BEFORE)     
      DPI_STS_R[0] <= 1'b1;
   else
      DPI_STS_R[0] <= 1'b0;
end

always @(posedge DPI_STS_CLR_N or negedge global_rstn or negedge lsr_rstn or posedge PD_AFTER) begin
   if (!global_rstn)
      DPI_STS_R[1] <= 0;
   else if (!lsr_rstn)
      DPI_STS_R[1] <= 0;
   else if (PD_AFTER)     
      DPI_STS_R[1] <= 1'b1;
   else
      DPI_STS_R[1] <= 1'b0;
end

assign DPI_STS[0] = DPI_STS_R[0];
assign DPI_STS[1] = DPI_STS_R[1];
     
always @(negedge ICLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      PADI_POS_fifo <= 0;
   else if (!lsr_rstn)
      PADI_POS_fifo <= 0;
   else
      PADI_POS_fifo[IFIFO_WADDR] <= DPI_P;

always @(negedge ICLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      PADI_NEG_fifo <= 0;
   else if (!lsr_rstn)
      PADI_NEG_fifo <= 0;
   else
      PADI_NEG_fifo[IFIFO_WADDR] <= PADI_SAMPLE;   
         
always @(posedge DESCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      shift_reg <= 0;
   else if (!lsr_rstn)
      shift_reg <= 0;
   else
      shift_reg <= {PADI_NEG_fifo[IFIFO_RADDR], PADI_POS_fifo[IFIFO_RADDR], shift_reg[3:2]};

always @(posedge DESCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn) begin
      capture_en_b <= 0;
      capture_en   <= 0;
   end   
   else if (!lsr_rstn) begin
      capture_en_b <= 0;
      capture_en   <= 0;      
   end
   else begin
      capture_en_b <= ~ capture_en_b;
      capture_en   <= capture_en_b;            
   end   

always @(posedge DESCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      capture_reg <= 0;
   else if (!lsr_rstn)
      capture_reg <= 0;
   else if (capture_en)
      capture_reg <= shift_reg;
      
always @(posedge RCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      Q_reg <= 0;
   else if (!lsr_rstn)
      Q_reg <= 0;
   else
      Q_reg <= capture_reg;      

assign Q = Q_reg;      
 

//synthesis translate_on

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2016 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_CLKBUFGMUX_E1.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_CLKBUFGMUX_E1
#(
    parameter TRIGGER_MODE = "NEGEDGE",
    parameter INIT_SEL = "CLK0"
) (
    output CLKOUT,
    input CLKIN0,
    input CLKIN1,
    input SEL,
    input EN
);

//synthesis translate_off

    initial begin
        if(TRIGGER_MODE != "POSEDGE" && TRIGGER_MODE != "NEGEDGE") begin
            $display("ERROR: The attribute TRIGGER_MODE on instance %m is %s. Legal value are POSEDGE or NEGEDGE.", TRIGGER_MODE);
            $finish;
        end
        if(INIT_SEL != "CLK0" && INIT_SEL != "CLK1") begin
            $display("ERROR: The attribute INIT_SEL on instance %m is %s. Legal value are CLK0 or CLK1.", INIT_SEL);
            $finish;
        end        
    end


///////////////////////////////////////initialization//////////////////////////////////////////////
    reg  clk_out_init_enable;
    
    initial begin
        clk_out_init_enable = 1;
        #0.1 clk_out_init_enable = 0;
    end



////////////////////////////////////////dynamic control///////////////////////////////////////////////
    wire clk0_pos;
    wire clk0_neg;
    wire clk1_pos;
    wire clk1_neg;

    reg clk0_syn_pos;
    reg clk0_syn_neg;
    reg clk1_syn_pos;
    reg clk1_syn_neg;
    reg clk0_syn_pos_temp;
    reg clk0_syn_neg_temp;
    reg clk1_syn_pos_temp;
    reg clk1_syn_neg_temp;
    reg clk_out_syn;
    reg clk_out;

    initial fork
        if(INIT_SEL == "CLK0") fork
            #0.1 clk0_syn_pos <= 1;
            #0.1 clk0_syn_neg <= 1;
            #0.1 clk1_syn_pos <= 0;
            #0.1 clk1_syn_neg <= 0;
            #0.1 clk0_syn_pos_temp <= 1;
            #0.1 clk0_syn_neg_temp <= 1;
            #0.1 clk1_syn_pos_temp <= 0;
            #0.1 clk1_syn_neg_temp <= 0;

        join
        else fork
            #0.1 clk0_syn_pos <= 0;
            #0.1 clk0_syn_neg <= 0;
            #0.1 clk1_syn_pos <= 1;
            #0.1 clk1_syn_neg <= 1;
            #0.1 clk0_syn_pos_temp <= 0;
            #0.1 clk0_syn_neg_temp <= 0;
            #0.1 clk1_syn_pos_temp <= 1;
            #0.1 clk1_syn_neg_temp <= 1;
        join
    join


    assign clk0_pos = (TRIGGER_MODE == "POSEDGE" && SEL == 0 && clk1_syn_pos == 0 && EN == 1) ? 1 : 0;
    assign clk0_neg = (TRIGGER_MODE == "NEGEDGE" && SEL == 0 && clk1_syn_neg == 0 && EN == 1) ? 1 : 0;
    assign clk1_pos = (TRIGGER_MODE == "POSEDGE" && SEL == 1 && clk0_syn_pos == 0 && EN == 1) ? 1 : 0;
    assign clk1_neg = (TRIGGER_MODE == "NEGEDGE" && SEL == 1 && clk0_syn_neg == 0 && EN == 1) ? 1 : 0;

    always @(posedge CLKIN0) begin
        if(!clk_out_init_enable)begin
            if(clk0_pos) begin
                clk0_syn_pos <= clk0_syn_pos_temp;
                clk0_syn_pos_temp <= 1'b1;
            end
            else begin
                clk0_syn_pos <= clk0_syn_pos_temp;
                clk0_syn_pos_temp <= 1'b0;
            end
        end
    end    
    
    always @(negedge CLKIN0) begin
        if(!clk_out_init_enable) begin
            if(clk0_neg) begin
                clk0_syn_neg <= clk0_syn_neg_temp;
                clk0_syn_neg_temp <= 1'b1;
            end
            else begin
                clk0_syn_neg <= clk0_syn_neg_temp;
                clk0_syn_neg_temp <= 1'b0;
            end
        end
    end    
    
    always @(posedge CLKIN1) begin
        if(!clk_out_init_enable) begin
            if(clk1_pos) begin
                clk1_syn_pos <= clk1_syn_pos_temp;
                clk1_syn_pos_temp <= 1'b1;
            end
            else begin
                clk1_syn_pos <= clk1_syn_pos_temp;
                clk1_syn_pos_temp <= 1'b0;
            end
        end
    end    
    
    always @(negedge CLKIN1) begin
        if(!clk_out_init_enable) begin
            if(clk1_neg) begin
                clk1_syn_neg <= clk1_syn_neg_temp;
                clk1_syn_neg_temp <= 1'b1;
            end
            else begin
                clk1_syn_neg <= clk1_syn_neg_temp;
                clk1_syn_neg_temp <= 1'b0;
            end
        end
    end    
    

    always@(*) begin
        if(TRIGGER_MODE == "POSEDGE") begin
            if(clk0_syn_pos) begin
                clk_out_syn = CLKIN0; 
            end
            else if(clk1_syn_pos) begin
                clk_out_syn = CLKIN1;
            end
            else begin
                clk_out_syn = 1;
            end
        end
        else begin
            if(clk0_syn_neg) begin
                clk_out_syn = CLKIN0; 
            end
            else if(clk1_syn_neg) begin
                clk_out_syn = CLKIN1;
            end
            else begin
                clk_out_syn = 0;
            end
        end
    end



///////////////////////////////////////////output/////////////////////////////////////////////

    assign CLKOUT = clk_out;

    always@(*)begin
        if(clk_out_init_enable) begin
            if(INIT_SEL == "CLK1") begin
                clk_out = CLKIN1;
            end
            else if(INIT_SEL == "CLK0")begin
                clk_out = CLKIN0;
            end
        end
        else begin
            clk_out = clk_out_syn;
        end
    end

//synthesis translate_on

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2015 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_FIFO36K_E1.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps
 
module  GTP_FIFO36K_E1
#(
    parameter GRS_EN = "TRUE",
    parameter integer DATA_WIDTH = 18,
    parameter integer DO_REG = 0,
    parameter ECC_WRITE_EN = "FALSE",
    parameter ECC_READ_EN = "FALSE",
    parameter [14:0]  ALMOST_FULL_OFFSET  = 15'h0000,
    parameter [14:0]  ALMOST_EMPTY_OFFSET = 15'h0000,
    parameter [71:0]  RST_VAL = 72'b0,
    parameter integer USE_EMPTY = 0,
    parameter integer USE_FULL = 0,
    parameter SYNC_FIFO = "FALSE"
)(
    output        ALMOST_EMPTY,
    output        ALMOST_FULL,
    output        EMPTY,
    output        FULL,
    output [71:0] DO,
    input  [71:0] DI,
    input         WCLK,
    input         RCLK,
    input         WCE,
    input         RCE,
    input         ORCE,
    input         RST,
    input         INJECT_SBITERR,
    input         INJECT_DBITERR,
    output        ECC_SBITERR,
    output        ECC_DBITERR
);
//synthesis translate_off
    reg  [15:0]   rd_binary;
    reg  [15:0]   wr_binary;
    reg  [14:0]   wcnt;
    reg  [14:0]   rcnt;
    reg  [15:0]   wr_binary_next;
    reg  [15:0]   rd_binary_next;
    reg           empty_reg;
    reg           full_reg;
    reg            full_val;
    reg           almost_full_reg;
    reg           almost_empty_reg;
    reg           flagempty_en;
    reg           flagfull_en;
    reg           dout_reg_en;
    reg           sync_fifo;
    reg           grs_en;
    reg              ecc_wren;
    reg              ecc_rden;
    reg  [71:0]   dout;
    reg  [71:0]   dout_reg;

    wire [71:0]   din_ecc;
    wire [71:0]   data_dec;
    wire [15:0]   wptr_next;
    wire [15:0]   rptr_next;
    reg  [15:0]   wptr_rclk;
    reg  [15:0]   rptr_wclk;
    wire [15:0]   wptr_next_gray;
    reg  [15:0]   wdata_buf;
    reg  [15:0]   wdata_buf_d1;
    reg  [15:0]   wdata_buf_d2;
    wire [15:0]   rptr_next_gray;
    reg  [15:0]   rdata_buf;
    reg  [15:0]   rdata_buf_d1;
    reg  [15:0]   rdata_buf_d2;
    wire          wclk,rclk;
    wire          wr_en,rd_en;
    wire          rstw,rstr;
    wire          full,empty;
    wire [71:0]   din;
    wire [71:0]   dout_ecc;
    wire [71:0]   dout_int;
    wire          almost_empty,almost_full;
    wire          global_rstn;
    wire [15:0]   rd_binary_inc;


//////////////////////////////////////////////////////////////////////////////
    reg  [(DATA_WIDTH-1):0] mem [(1<<15)-1 : 0];

    initial   
    begin
        case(SYNC_FIFO)
            "FALSE" : sync_fifo = 0;
            "TRUE"  : sync_fifo = 1;
            default : begin
                $display ("ERROR: GTP_FIFO36K_E1 instance %m parameter SYNC_FIFO:%s, The legal values are FALSE or TRUE.",SYNC_FIFO);
                $finish;
            end
        endcase
        
        case(USE_EMPTY)
            1'b0 : flagempty_en = 0;
            1'b1 : flagempty_en = 1;
            default : begin
                $display ("ERROR: GTP_FIFO36K_E1 instance %m parameter USE_EMPTY:%d, The legal values are 0 or 1.",USE_EMPTY);
                $finish;
            end
        endcase
        
        case(USE_FULL)
            1'b0 : flagfull_en = 0;
            1'b1 : flagfull_en = 1;
            default : begin
                $display ("ERROR: GTP_FIFO36K_E1 instance %m parameter USE_FULL:%d, The legal values are 0 or 1.",USE_FULL);
                $finish;
            end
        endcase
        
        case(DO_REG)
            1'b0 : dout_reg_en = 0;
            1'b1 : dout_reg_en = 1;
            default : begin
                $display ("ERROR: GTP_FIFO36K_E1 instance %m parameter DO_REG:%d, The legal values are 0 or 1.",DO_REG);
                $finish;
            end
        endcase
    
        case(GRS_EN)
            "FALSE" : grs_en = 0;
            "TRUE"  : grs_en = 1;
            default : begin
                $display ("ERROR: GTP_FIFO36K_E1 instance %m parameter GRS_EN:%s, The legal values are FALSE or TRUE.",GRS_EN);
                $finish;
            end
        endcase

        case(ECC_WRITE_EN)
            "FALSE" : ecc_wren = 0;
            "TRUE"  : begin 
                ecc_wren = 1;
                if(DATA_WIDTH != 72) begin
                    $display ("ERROR: GTP_FIFO36K_E1 instance %m parameter DATA_WIDTH:%s not supported when ECC_WRITE_EN = TRUE.",DATA_WIDTH);
                    $finish;
                end
            end
            default : begin
                $display ("ERROR: GTP_FIFO36K_E1 instance %m parameter ECC_WRITE_EN:%s, The legal values are FALSE or TRUE.",ECC_WRITE_EN);
                $finish;
            end
        endcase

        case(ECC_READ_EN)
            "FALSE" : ecc_rden = 0;
            "TRUE"  : begin
                ecc_rden = 1;
                if(DATA_WIDTH != 72) begin
                    $display ("ERROR: GTP_FIFO36K_E1 instance %m parameter DATA_WIDTH:%s not supported when ECC_READ_EN = TRUE.",DATA_WIDTH);
                    $finish;
                end
            end
            default : begin
                $display ("ERROR: GTP_FIFO36K_E1 instance %m parameter ECC_READ_EN:%s, The legal values are FALSE or TRUE.",ECC_READ_EN);
                $finish;
            end
        endcase

        dout_reg ='b0;
    end
//////////////////////////////////////////////////////////////////////////////////////
    assign orce_in = ORCE;
    assign din = din_ecc;
    assign wclk = WCLK;
    assign rclk = RCLK;
    assign wr_en = WCE;
    assign rd_en = RCE;
    assign rstw = ~RST & global_rstn;
    assign rstr = ~RST & global_rstn;
    assign EMPTY = empty;
    assign FULL  = full;
    assign ALMOST_EMPTY = almost_empty;
    assign ALMOST_FULL = almost_full;
    assign WCNT = wcnt;
    assign RCNT = rcnt;
    
    always @(posedge rclk or negedge rstr )
    begin
        if(rstr == 1'b0)
            dout_reg <= RST_VAL;
        else if(orce_in)
            dout_reg <= dout_int;
    end    
    
    assign DO = dout_reg_en ? dout_reg : dout_int;
    
    assign global_rstn = grs_en ? GRS_INST.GRSNET : 1'b1;
//////////////////////////////////////////////////////////////////////////////////////
    always @ (posedge wclk or negedge rstw )  //////wr binary addr
    begin
        if (rstw == 1'b0)
             wr_binary <= 0;
        else
             wr_binary <= wr_binary_next;
    end
    
    always @ (*)
    begin
        if (full == 1'b0)
             wr_binary_next = wr_binary + wr_en;
        else
             wr_binary_next = wr_binary;
    end
    
    assign wptr_next = wr_binary_next;
//////////////////////////////////////////////////////////////////////////////////////
    always @ (*) begin
        case(DATA_WIDTH)
        1: begin
             full_val = (wr_binary_next[15:0] == {~rptr_wclk[15],rptr_wclk[14:0]});
        end
        2: begin
             full_val = (wr_binary_next[14:0] == {~rptr_wclk[14],rptr_wclk[13:0]});
        end
        4: begin
             full_val = (wr_binary_next[13:0] == {~rptr_wclk[13],rptr_wclk[12:0]});
        end
        8: begin
             full_val = (wr_binary_next[12:0] == {~rptr_wclk[12],rptr_wclk[11:0]});
        end
        9: begin
             full_val = (wr_binary_next[12:0] == {~rptr_wclk[12],rptr_wclk[11:0]});
        end
        16: begin
             full_val = (wr_binary_next[11:0] == {~rptr_wclk[11],rptr_wclk[10:0]});
        end
        18: begin
             full_val = (wr_binary_next[11:0] == {~rptr_wclk[11],rptr_wclk[10:0]});
        end
        32,36: begin
             full_val = (wr_binary_next[10:0] == {~rptr_wclk[10],rptr_wclk[9:0]});
        end
        64,72: begin
             full_val = (wr_binary_next[9:0] == {~rptr_wclk[9],rptr_wclk[8:0]});
        end
        default: begin  //default x18
             full_val = (wr_binary_next[11:0] == {~rptr_wclk[11],rptr_wclk[10:0]});
        end
        endcase
    end
    
    always @ (posedge wclk or negedge rstw) begin //////write full flag
        if (rstw == 1'b0)
             full_reg <= 1'b0;
        else
             full_reg <= full_val;
    end
    
    assign full = flagfull_en & full_reg;
    
    always @ (posedge wclk or negedge rstw) begin //////write almost_full flag
        if (rstw == 1'b0)
             almost_full_reg <= 1'b0;
        else
             almost_full_reg <= (wr_binary_next- rptr_wclk) >= ALMOST_FULL_OFFSET;
    end
    
    assign almost_full = flagfull_en & almost_full_reg;
//////////////////////////////////////////////////////////////////////////////////////
    always @ (posedge rclk or negedge rstr) begin
        if(rstr == 1'b0)
             rd_binary <= 0;
        else
             rd_binary <= rd_binary_next;
    end


    always @ (*) begin
          if ((~empty_reg) & rd_en)
             rd_binary_next = rd_binary + 1;
          else
             rd_binary_next = rd_binary;
    end
    
    assign rptr_next = rd_binary_next;

    always @ (posedge rclk or negedge rstr) begin
          if (rstr == 1'b0) begin
              empty_reg <= 1'b1;
          end
          else begin
              empty_reg <= wptr_rclk == rd_binary_next;
          end
    end
    
    assign empty = ~flagempty_en |empty_reg;
    
    always @ (posedge rclk or negedge rstr) begin
          if (rstr == 1'b0) begin
              almost_empty_reg <= 1'b1;
          end
          else begin
              almost_empty_reg <= (wptr_rclk - rd_binary_next) <= ALMOST_EMPTY_OFFSET;
          end
    end
    
    assign almost_empty = ~flagempty_en |almost_empty_reg;
//////////////////////////////////////////////////////////////////////////////////////
    always @ (wr_binary) begin
        case(DATA_WIDTH)
             1:     wcnt <=  wr_binary[14:0];
             2:     wcnt <= {wr_binary[13:0],1'b1};
             4:     wcnt <= {wr_binary[12:0],2'b11};
             8:     wcnt <= {wr_binary[11:0],3'b111};
             9:     wcnt <= {wr_binary[11:0],3'b111};
             16:    wcnt <= {wr_binary[10:0],4'b1111};
             18:    wcnt <= {wr_binary[10:0],4'b1111};
             32:    wcnt <= {wr_binary[9:0],5'b1111};
             36:    wcnt <= {wr_binary[9:0],5'b1111};
             64:    wcnt <= {wr_binary[8:0],5'b1111};
             72:    wcnt <= {wr_binary[8:0],5'b1111};
             default:
                    wcnt <= 15'b0;
        endcase
    end
    
    always @ (rd_binary) begin
        case(DATA_WIDTH)
             1:     rcnt <=  rd_binary[14:0];
             2:     rcnt <= {rd_binary[13:0],1'b1};
             4:     rcnt <= {rd_binary[12:0],2'b11};
             8:     rcnt <= {rd_binary[11:0],3'b111};
             9:     rcnt <= {rd_binary[11:0],3'b111};
             16:    rcnt <= {rd_binary[10:0],4'b1111};
             18:    rcnt <= {rd_binary[10:0],4'b1111};
             32:    rcnt <= {rd_binary[9:0],5'b1111};
             36:    rcnt <= {rd_binary[9:0],5'b1111};
             64:    rcnt <= {rd_binary[8:0],5'b1111};
             72:    rcnt <= {rd_binary[8:0],5'b1111};
             default:
                    rcnt <= 15'b0;
        endcase
    end
//////////////////////////////////////////////////////////////////////////////////////
    assign wptr_next_gray = (wptr_next>>1)^wptr_next;
    assign rptr_next_gray = (rptr_next>>1)^rptr_next;
    
    always @(posedge wclk or negedge rstw)
    begin
        if(rstw == 1'b0)
        begin 
            wdata_buf <= 0;
            rdata_buf_d1 <= 0;
            rdata_buf_d2 <= 0;
        end else begin
            wdata_buf <= wptr_next_gray;
            rdata_buf_d1 <= rdata_buf;
            if(sync_fifo)
                rdata_buf_d2 <= rptr_next_gray;
            else
                rdata_buf_d2 <= rdata_buf_d1;
        end
    end
    
    always @(posedge rclk or negedge rstr)
    begin
        if(rstr == 1'b0)
        begin
            wdata_buf_d1 <= 0;
            wdata_buf_d2 <= 0;
            rdata_buf <= 0;
        end else begin
            wdata_buf_d1 <= wdata_buf;
            rdata_buf <= rptr_next_gray;
            if(sync_fifo)
                wdata_buf_d2 <= wptr_next_gray;
            else
                wdata_buf_d2 <= wdata_buf_d1;
        end
    end
    
    integer i,j,k;
    
    always @(wdata_buf_d2) begin
       for (i=0; i< 16;i=i+1)
           wptr_rclk[i] = ^(wdata_buf_d2>>i);
    end
    
    always @(rdata_buf_d2) begin
       for (j=0; j< 16;j=j+1)
           rptr_wclk[j] = ^(rdata_buf_d2>>j);
    end
//////////////////////////////////////////////////////////////////////////////////////
    initial
    begin
        for(k=0;k<(1<<15);k=k+1)
            mem[k] <= {DATA_WIDTH{1'b0}};
    end
    
    always @(posedge rclk or negedge rstr)
    begin
        if(rstr == 1'b0)
            dout <= RST_VAL;
        else if(rd_en)
            dout <= mem[rcnt];
    end

    assign dout_int = ecc_rden ? data_dec : dout;


    always @(posedge wclk)
    begin
        if(wr_en && !full_reg)
            mem[wcnt] <= din;
    end


//////////////////////////////////////////ecc/////////////////////////////////////////

    wire clkqb0;
    reg rst_ecc;
    assign clkqb0 = RCLK&ORCE;
    initial begin
        rst_ecc = 1;
        #0.1 rst_ecc = 0;
    end


wire        SC_ECC_WREN;
wire [63:0] WD;
wire [7:0]  ADD_DATA;
wire        ECC_INJ_SBITERR;
wire        ECC_INJ_DBITERR;
wire [71:0] DATA_TO_SDP;
wire [7:0]  ECC_PARTY;
wire        SC_ECC_RDEN;
wire [71:0] DATA_FROM_SDP;
wire [71:0] RD;
wire        SC_ORCE;
wire        rst;
wire [8:0]  ecc_rdaddr;
wire [8:0]  ECC_RDADDR;
wire        porn_int;
wire        pcka;
wire        pcea;
wire        ckqb;

assign SC_ECC_WREN = ecc_wren;
assign WD = {DI[70:63], DI[61:54], DI[52:45], DI[43:36], DI[34:27], DI[25:18], DI[16:9], DI[7:0]};
assign ADD_DATA = {DI[71], DI[62], DI[53], DI[44], DI[35], DI[26],DI[17], DI[8]};
assign ECC_INJ_SBITERR = INJECT_SBITERR;
assign ECC_INJ_DBITERR = INJECT_DBITERR;
assign din_ecc = DATA_TO_SDP;
assign SC_ECC_RDEN = ecc_rden;
assign DATA_FROM_SDP = dout;
assign data_dec = RD;
assign SC_OREB = dout_reg_en;
assign rst = rst_ecc;
assign porn_int = 1'b0;
assign pcka = 1'b1;
assign pcea = 1'b1;
assign ckqb = clkqb0;


//ECC Encoder
wire          ERR30bit;
wire          ERR62bit;
wire  [63:0]  data_enc63;
wire  [71:0]  DATA_no_enc;
wire  [71:0]  DATA_enc72;
wire  [7:0]   ecc_parity;

assign ecc_parity[7] = (WD[63]) ^ (WD[60]) ^ (^WD[58:56]) ^ (WD[53]) ^ (^WD[51:50]) ^ (^WD[47:46]) ^ (WD[44]) ^ (WD[41]) ^ (^WD[39:38]) ^ (WD[36]) ^ (^WD[33:32]) ^ (WD[29]) ^ (^WD[27:26]) ^ (^WD[24:23]) ^ (WD[21]) ^ (^WD[18:17]) ^ (WD[14]) ^ (^WD[12:10]) ^ WD[7] ^ (^WD[5:4]) ^ (^WD[2:0]);
assign ecc_parity[6] = ^WD[63:57];
assign ecc_parity[5] = ^WD[56:26];
assign ecc_parity[4] = ( ^WD[56:41] ) ^ ( ^WD[25:11] );
assign ecc_parity[3] = ( ^WD[56:49] ) ^ ( ^WD[40:33] ) ^ ( ^WD[25:18] ) ^ ( ^WD[10:4] );
assign ecc_parity[2] = ( ^WD[63:60] ) ^ ( ^WD[56:53] ) ^ ( ^WD[48:45] ) ^ ( ^WD[40:37] ) ^ ( ^WD[32:29] ) ^ ( ^WD[25:22] ) ^ ( ^WD[17:14] ) ^ ( ^WD[10:7] ) ^ ( ^WD[3:1] );
assign ecc_parity[1] = ( ^WD[63:62] ) ^ ( ^WD[59:58] ) ^ ( ^WD[56:55] ) ^ ( ^WD[52:51] ) ^ ( ^WD[48:47] ) ^ ( ^WD[44:43] ) ^ ( ^WD[40:39] ) ^ ( ^WD[36:35] ) ^ ( ^WD[32:31] ) ^ ( ^WD[28:27] ) ^ ( ^WD[25:24] ) ^ ( ^WD[21:20] ) ^( ^WD[17:16] )^( ^WD[13:12] ) ^ ( ^WD[10:9] ) ^ ( ^WD[6:5] ) ^ ( ^WD[3:2] ) ^ WD[0] ;
assign ecc_parity[0] = WD[63] ^ WD[61] ^ WD[59] ^ ( ^WD[57:56] ) ^ WD[54] ^ WD[52] ^ WD[50] ^ WD[48] ^ WD[46] ^ WD[44] ^ WD[42] ^ WD[40] ^ WD[38] ^ WD[36] ^ WD[34] ^ WD[32] ^ WD[30] ^ WD[28] ^ ( ^WD[26:25] ) ^ WD[23] ^ WD[21] ^ WD[19] ^ WD[17] ^ WD[15] ^ WD[13] ^ ( ^WD[11:10] ) ^ WD[8] ^ WD[6] ^ ( ^WD[4:3] ) ^ ( ^WD[1:0] ) ;



assign ERR30bit = (ECC_INJ_SBITERR || ECC_INJ_DBITERR) ? ~WD[30] : WD[30];
assign ERR62bit = ECC_INJ_DBITERR ? ~WD[62] : WD[62];
assign data_enc63 = {WD[63],ERR62bit,WD[61:31],ERR30bit,WD[29:0]};


assign DATA_no_enc = {ADD_DATA[7],WD[63:56],ADD_DATA[6],WD[55:48],
    ADD_DATA[5],WD[47:40],ADD_DATA[4],WD[39:32],ADD_DATA[3],WD[31:24],
    ADD_DATA[2],WD[23:16],ADD_DATA[1],WD[15:8],ADD_DATA[0],WD[7:0]}; 

assign DATA_enc72 = {ecc_parity[7],data_enc63[63:56],ecc_parity[6],data_enc63[55:48],
    ecc_parity[5],data_enc63[47:40],ecc_parity[4],data_enc63[39:32],ecc_parity[3],data_enc63[31:24],
    ecc_parity[2],data_enc63[23:16],ecc_parity[1],data_enc63[15:8],ecc_parity[0],data_enc63[7:0]}; 

assign DATA_TO_SDP = SC_ECC_WREN ? DATA_enc72 : DATA_no_enc;








//ECC Decoder
wire  [71:0]  data_dec1;
wire          ecc_sbiterr;
wire          ecc_dbiterr;
wire  [63:0]  DO1;
wire  [7:0]   DOP;
wire  [7:0]   dec_syndrome;
wire          ecc_err;
wire  [6:0]   err_pos;
reg   [71:0]  ecc_corrected;

assign DO1 = {DATA_FROM_SDP[70:63],DATA_FROM_SDP[61:54],DATA_FROM_SDP[52:45],DATA_FROM_SDP[43:36],DATA_FROM_SDP[34:27],DATA_FROM_SDP[25:18],DATA_FROM_SDP[16:9],DATA_FROM_SDP[7:0]};
assign DOP = {DATA_FROM_SDP[71],DATA_FROM_SDP[62],DATA_FROM_SDP[53],DATA_FROM_SDP[44],DATA_FROM_SDP[35],DATA_FROM_SDP[26],DATA_FROM_SDP[17],DATA_FROM_SDP[8]};


assign dec_syndrome[7] = ((DO1[63]) ^ (DO1[60]) ^ (^DO1[58:56]) ^ (DO1[53]) ^ (^DO1[51:50]) ^ (^DO1[47:46]) ^ (DO1[44]) ^ (DO1[41]) ^ (^DO1[39:38]) ^ (DO1[36]) ^ (^DO1[33:32]) ^ (DO1[29]) ^ (^DO1[27:26]) ^ (^DO1[24:23]) ^ (DO1[21]) ^ (^DO1[18:17]) ^ (DO1[14]) ^ (^DO1[12:10]) ^ DO1[7] ^ (^DO1[5:4]) ^ (^DO1[2:0]))^DOP[7];  
assign dec_syndrome[6] = (^DO1[63:57])^DOP[6];
assign dec_syndrome[5] = (^DO1[56:26])^DOP[5];
assign dec_syndrome[4] = (^DO1[56:41])^(^DO1[25:11])^DOP[4];
assign dec_syndrome[3] = (^DO1[56:49])^(^DO1[40:33])^(^DO1[25:18])^(^DO1[10:4])^DOP[3];
assign dec_syndrome[2] = (^DO1[63:60])^(^DO1[56:53])^(^DO1[48:45])^(^DO1[40:37])^(^DO1[32:29])^(^DO1[25:22])^(^DO1[17:14])^(^DO1[10:7])^(^DO1[3:1])^DOP[2];
assign dec_syndrome[1] = (^DO1[63:62])^(^DO1[59:58])^(^DO1[56:55])^(^DO1[52:51])^(^DO1[48:47])^(^DO1[44:43])^(^DO1[40:39])^(^DO1[36:35])^(^DO1[32:31])^(^DO1[28:27])^(^DO1[25:24])^(^DO1[21:20])^(^DO1[17:16])^(^DO1[13:12])^(^DO1[10:9])^(^DO1[6:5])^(^DO1[3:2])^DO1[0]^DOP[1];
assign dec_syndrome[0] = DO1[63]^DO1[61]^DO1[59]^(^DO1[57:56])^DO1[54]^DO1[52]^DO1[50]^DO1[48]^DO1[46]^DO1[44]^DO1[42]^DO1[40]^DO1[38]^DO1[36]^DO1[34]^DO1[32]^DO1[30]^DO1[28]^(^DO1[26:25])^DO1[23]^DO1[21]^DO1[19]^DO1[17]^DO1[15]^DO1[13]^(^DO1[11:10])^DO1[8]^DO1[6]^(^DO1[4:3])^(^DO1[1:0])^DOP[0];

assign	ecc_err = |dec_syndrome[6:0];	//dec_syndrome != 0;
assign 	err_pos = dec_syndrome[6:0];

assign ecc_sbiterr = ^dec_syndrome;
assign ecc_dbiterr = ecc_err && ~(^dec_syndrome);

always @(*) begin
    ecc_corrected = {DO1[63:57], DOP[6], DO1[56:26], DOP[5], DO1[25:11], DOP[4], DO1[10:4], DOP[3], DO1[3:1], DOP[2], DO1[0], DOP[1:0], DOP[7]};

    ecc_corrected[err_pos] = ~ecc_corrected[err_pos];
end
assign data_dec1 = {ecc_corrected[0],ecc_corrected[71:65],ecc_corrected[63],ecc_corrected[64],ecc_corrected[62:55],ecc_corrected[32],ecc_corrected[54:47],ecc_corrected[16],ecc_corrected[46:39],ecc_corrected[8],ecc_corrected[38:33],ecc_corrected[31:30],ecc_corrected[4],ecc_corrected[29:22],ecc_corrected[2],ecc_corrected[21:17],ecc_corrected[15:13],ecc_corrected[1],ecc_corrected[12:9],ecc_corrected[7:5],ecc_corrected[3]};
assign RD = (SC_ECC_RDEN && ecc_sbiterr) ? data_dec1 : DATA_FROM_SDP; 





//OR
reg  [8:0]    ecc_rdaddr_reg;
reg           ecc_sbiterr_reg;
reg           ecc_dbiterr_reg;
reg  [7:0]    ecc_parity_reg;

initial begin
    ecc_sbiterr_reg <= 1'b0;
    ecc_dbiterr_reg <= 1'b0;
end

always @(posedge ckqb or posedge rst)
begin
    if (rst) 
    begin
        ecc_rdaddr_reg <= 9'b0;
        ecc_sbiterr_reg <= 1'b0;
        ecc_dbiterr_reg <= 1'b0;
    end
    else 
    begin
        ecc_rdaddr_reg <= ecc_rdaddr;
        ecc_sbiterr_reg <= ecc_sbiterr;
        ecc_dbiterr_reg <= ecc_dbiterr;
    end
end

always @(posedge pcka or negedge porn_int)
begin
    if (!porn_int) 
    begin
        ecc_parity_reg <= 8'b0;
    end
    else if (pcea) 
    begin
        ecc_parity_reg <= ecc_parity;
    end
end

assign ECC_RDADDR =  (SC_ECC_RDEN == 1'b0) ? 9'h1ff : (SC_OREB ? ecc_rdaddr_reg : ecc_rdaddr);
assign ECC_SBITERR = (SC_ECC_RDEN == 1'b0) ? 1'b1 : (SC_OREB ? ecc_sbiterr_reg : ecc_sbiterr);
assign ECC_DBITERR = (SC_ECC_RDEN == 1'b0) ? 1'b1 : (SC_OREB ? ecc_dbiterr_reg : ecc_dbiterr);
assign ECC_PARITY = (SC_ECC_WREN == 1'b0) ? 8'hff : ecc_parity_reg;

// synthesis translate_on
endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_ROM128X1.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_ROM128X1
#(
    parameter [127:0] INIT = 128'h00000000_00000000_00000000_00000000
) (
    output Z,
    input I0, I1, I2, I3, I4, I5, I6
);

   reg [127:0] mem;
   wire [7:0] addr;

   initial mem = INIT;

   assign addr = {I6, I5, I4, I3, I2, I1, I0};
   //assign Z = mem[addr];
   assign Z = INIT[addr];

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_INBUFEDS.v
//
// Functional description: Differential Signaling Input Buffer
//
// Parameter description:
//
// Port description:
//
// Revision:
//    06/18/14 - Initial version.
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_INBUFEDS #(
    parameter IOSTANDARD = "DEFAULT",
    parameter TERM_DIFF = "ON"
)(
    output reg O,
    input EN,                    // 1: enable inbuf, normal mode; 0: disable inbuf, standby mode.
    input I,
    input IB
) /* synthesis syn_black_box */ ;
  
  initial begin
    case (IOSTANDARD)
    "LVDS", "MINI-LVDS", "LVPECL", "SUB-LVDS", "SSTL18D_I", "SSTL18D_II", "SSTL15D_I", "SSTL15D_II", "HSTL18D_I", "HSTL18D_II", "HSTL15D_I", "SSTL25D_I", "RSDS", "PPDS", "TMDS", "SSTL25D_II", "BLVDS", "SSTL15D_I_CAL", "SSTL15D_II_CAL", "HSTL15D_I_CAL", "DEFAULT" :;
    default : begin
           $display("Attribute Syntax Error : The attribute IOSTANDARD on GTP_INBUFDS instance %m is set to %s.", IOSTANDARD);
           $finish;
              end
    endcase

    case (TERM_DIFF)
    "ON", "OFF" :;
    default : begin
           $display("Attribute Syntax Error : The attribute TERM_DIFF on GTP_INBUFDS instance %m is set to %s.", TERM_DIFF);
           $finish;
              end
    endcase
    end

    always @(*)
    begin
        if (EN == 1'b1)
            O = I && ~IB;
        else
            O = 1'b1;
    end

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_PREADD_MULTADDACC18.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

//P = MAC + (A0*(B0+C0) + A1*(B1+C1))
`timescale 1 ns / 1 ps

module GTP_PREADD_MULTADDACC18 #(
    parameter GRS_EN            = "TRUE", //"TRUE"; "FALSE"
    parameter SYNC_RST          = "FALSE", //"TRUE"; "FALSE"
    parameter INREG_EN          = "FALSE",  //"TRUE"; "FALSE"
    parameter PREREG_EN         = "FALSE",  //"TRUE"; "FALSE"
    parameter PIPEREG_EN        = "FALSE",//"TRUE"; "FALSE"
    parameter ADDSUB_OP         = 0 ,
    parameter ACC_ADDSUB_OP     = 0,
    parameter DYN_ADDSUB_OP     = 1,
    parameter DYN_ACC_ADDSUB_OP = 1,
    parameter OVERFLOW_MASK     = 64'h0,  //PSIZE = 64 OVERflow setting = 'h10000_0000_0000_0000 , bit width = PSIZE
    parameter PATTERN           = 64'h0,  //compare pattern
    parameter MASKPAT           = 64'h0,  //pattern mask
    parameter ACC_INIT_VALUE    = 64'h0   //ACC_INIT_VALUE value
) (
    output  [63:0] P,
    output  OVER,
    output  UNDER,
    output  EQZ,
    output  EQZM,
    output  EQOM,
    output  EQPAT,
    output  EQPATN,

    input   CE,
    input   RST,
    input   CLK,
    input   A_SIGNED,
    input   [17:0] A0,
    input   [17:0] A1,
    input   B_SIGNED,
    input   [17:0] B0,
    input   [17:0] B1,
    input   C_SIGNED,
    input   [17:0] C0,
    input   [17:0] C1,
    input   [1:0] PREADDSUB,
    input   ADDSUB,
    input   ACC_ADDSUB,
    input   RELOAD
);

    wire [63:0] R;

    INT_PREADD_MULTADDACC #(
        . GRS_EN(GRS_EN),      
        . SYNC_RST(SYNC_RST),    
        . INREG_EN(INREG_EN),    
        . PREREG_EN(PREREG_EN),    
        . PIPEREG_EN(PIPEREG_EN),  
        . ADDSUB_OP(ADDSUB_OP),     
        . ACCUMADDSUB_OP(ACC_ADDSUB_OP),
        . DYN_OP_ADDSUB(DYN_ADDSUB_OP),   
        . DYN_OP_ACC(DYN_ACC_ADDSUB_OP),   
        . ASIZE(18),
        . BSIZE(18),
        . PSIZE(64),
        . DYN_ACC_INIT(0),
        . ACC_INIT_VALUE(ACC_INIT_VALUE),
        . MASK(OVERFLOW_MASK)
    ) U_MACC (
        . CE(CE),
        . RST(RST),
        . CLK(CLK),
        . A_SIGNED(A_SIGNED),
        . A0(A0),
        . A1(A1),
        . B_SIGNED(B_SIGNED),
        . B0(B0),
        . B1(B1),
        . C_SIGNED(C_SIGNED),
        . C0(C0),
        . C1(C1),
        . PREADDSUB(PREADDSUB),
        . ACCUM_INIT(64'b0),
        . ADDSUB(ADDSUB),
        . ACCUMADDSUB(ACC_ADDSUB),
        . RELOAD(RELOAD),
        . P(P),
        . OVER(OVER),
        . UNDER(UNDER),
        . R(R) 
    );     

    INT_FLAG #(
        . GRS_EN(GRS_EN),
        . SYNC_RST(SYNC_RST),
        . PSIZE(64),
        . PATSIZE(64),
        . MASKPATSIZE(64),
        . OUTREG_EN("TRUE")
    ) U_FLAG (
        . CE(CE),
        . RST(RST),
        . CLK(CLK),
        . P(P),
        . PATTERN(PATTERN),
        . MASKPAT(MASKPAT),
        . OVERFLOW_MASK(OVERFLOW_MASK),
        . R(R),
        . eqz(EQZ),
        . eqzm(EQZM),
        . eqom(EQOM),
        . eqpat(EQPAT),
        . eqpatn(EQPATN)
    );

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module INT_PSE #(
    parameter   ASIZE = 9,
    parameter  [ASIZE-2:0] SC_PSE = 0
) (
    input      [ASIZE-1:0] A,
    input                  SIGN,
    output reg [ASIZE-1:0] A_PSE
);

localparam SC_SIGNED_EN = (ASIZE == 26 || ASIZE == 27) ? 1'b1 : 1'b0;
         
integer i;
always @ (*) begin
    // ((|SC_PSE)==1'b1) means PSE enabled
    A_PSE[ASIZE-1] = ((|SC_PSE)==1'b1) ? A[ASIZE-1] & (~SC_SIGNED_EN | SIGN) : A[ASIZE-1];
    for (i=0; i <= ASIZE-2; i=i+1) begin
        A_PSE[i] = A[i] | (SC_PSE[i] & A[ASIZE-1] & (~SC_SIGNED_EN | SIGN));
    end
end  
endmodule


module INT_REG #(
    parameter SIZE = 1
) (
    input [SIZE-1:0] D,
    input BYPASS,
    input CLK, CE,
    input ARST, SRST,
    output [SIZE-1:0] Q
);
reg  [SIZE-1:0] qout;
initial qout = {SIZE{1'b0}};
always @(posedge CLK or posedge ARST) begin
    if (ARST == 1'b1)
        qout <= {SIZE{1'b0}};
    else if (SRST == 1'b1)
        qout <= {SIZE{1'b0}};
    else if (CE == 1'b1)
        qout <= D;
end
assign Q = (BYPASS == 1'b1) ? D : qout;
endmodule


module INT_REG2D #(
    parameter SIZE = 1
) (
    input DSEL,
    input [SIZE-1:0] D0,
    input [SIZE-1:0] D1,
    input BYPASS,
    input CLK, CE,
    input ARST, SRST,
    output [SIZE-1:0] Q
);
reg  [SIZE-1:0] qout;
wire [SIZE-1:0] din;
initial qout = {SIZE{1'b0}};
assign din = (DSEL == 1'b0) ? D0 : D1;
always @(posedge CLK or posedge ARST) begin
    if (ARST == 1'b1)
        qout <= {SIZE{1'b0}};
    else if (SRST == 1'b1)
        qout <= {SIZE{1'b0}};
    else if (CE == 1'b1)
        qout <= din;
end
assign Q = (BYPASS == 1'b1) ? din : qout;
endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2016 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library:
// Filename: GTP_DDRC.v
//
// Functional description:DDR Controller
//
// Parameter description:
//
// Port description:
//
// Revision:1.1
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1ns/1ps

module GTP_DDRC (
    input                                CORE_DDRC_CORE_CLK,
    input                                CORE_DDRC_RST,

    //----------------------------------------------- 
    // AXI Interface
    //-----------------------------------------------
    // AXI Port 0 Global Signals (clock, reset, low-power)
    input                                ARESET_0,
    input                                ACLK_0,
    // AXI Port 0 Write Address Channel
    input[7:0]                           AWID_0,
    input[31:0]                          AWADDR_0,
    input[7:0]                           AWLEN_0,
    input[2:0]                           AWSIZE_0,
    input[1:0]                           AWBURST_0,
    input                                AWLOCK_0,
    
    
    input                                AWVALID_0,
    output                               AWREADY_0,
    input                                AWURGENT_0,
    input                                AWPOISON_0,
        
    
    // AXI Port 0 Write Data Channel
    input[127:0]                         WDATA_0,
    input[15:0]                          WSTRB_0,
    input                                WLAST_0,
    input                                WVALID_0,
    output                               WREADY_0,
    
    // AXI Port 0 Write Response Channel
    output[7:0]                          BID_0,
    output[1:0]                          BRESP_0,
    output                               BVALID_0,
    input                                BREADY_0,
    
    // AXI Port 0 Read Address Channel
    input[7:0]                           ARID_0,
    input[31:0]                          ARADDR_0,
    input[7:0]                           ARLEN_0,
    input[2:0]                           ARSIZE_0,
    input[1:0]                           ARBURST_0,
    input                                ARLOCK_0,
    
    input                                ARVALID_0,
    output                               ARREADY_0,
    input                                ARPOISON_0,
       
    // AXI Port 0 Read Data Channel
    output[7:0]                          RID_0,
    output[127:0]                        RDATA_0,
    output[1:0]                          RRESP_0,
    output                               RLAST_0,
    output                               RVALID_0,
    input                                RREADY_0,
    input                                ARURGENT_0,
    output                               RAQ_PUSH_0,
    output                               RAQ_SPLIT_0,                                       
    output                               WAQ_PUSH_0,
    output                               WAQ_SPLIT_0,

          
    // AXI Port 1 Global Signals (clock, reset, low-power)
    input                                ARESET_1,
    input                                ACLK_1,
    // AXI Port 1 Write Address Channel
    input[7:0]                           AWID_1,
    input[31:0]                          AWADDR_1,
    input[7:0]                           AWLEN_1,
    input[2:0]                           AWSIZE_1,
    input[1:0]                           AWBURST_1,
    input                                AWLOCK_1,
    
    input                                AWVALID_1,
    output                               AWREADY_1,
    input                                AWURGENT_1,
    input                                AWPOISON_1,
          
    // AXI Port 1 Write Data Channel
    input[63:0]                          WDATA_1,
    input[7:0]                           WSTRB_1,
    input                                WLAST_1,
    input                                WVALID_1,
    output                               WREADY_1,
    
    // AXI Port 1 Write Response Channel
    output[7:0]                          BID_1,
    output[1:0]                          BRESP_1,
    output                               BVALID_1,
    input                                BREADY_1,
    
    // AXI Port 1 Read Address Channel
    input[7:0]                           ARID_1,
    input[31:0]                          ARADDR_1,
    input[7:0]                           ARLEN_1,
    input[2:0]                           ARSIZE_1,
    input[1:0]                           ARBURST_1,
    input                                ARLOCK_1,
    
    input                                ARVALID_1,
    output                               ARREADY_1,
    input                                ARPOISON_1,
          
    // AXI Port 1 Read Data Channel
    output[7:0]                          RID_1,
    output[63:0]                         RDATA_1,
    output[1:0]                          RRESP_1,
    output                               RLAST_1,
    output                               RVALID_1,
    input                                RREADY_1,
                                        
    input                                ARURGENT_1,
    output                               RAQ_PUSH_1,
    output                               RAQ_SPLIT_1,                                       
    output                               WAQ_PUSH_1,
    output                               WAQ_SPLIT_1,
    
    // AXI Port 2 Global Signals (clock, reset, low-power)
    input                                ARESET_2,
    input                                ACLK_2,
    // AXI Port 2 Write Address Channel
    input[7:0]                           AWID_2,
    input[31:0]                          AWADDR_2,
    input[7:0]                           AWLEN_2,
    input[2:0]                           AWSIZE_2,
    input[1:0]                           AWBURST_2,
    input                                AWLOCK_2,
    
    input                                AWVALID_2,
    output                               AWREADY_2,
    input                                AWURGENT_2,
    input                                AWPOISON_2,
    
       
    // AXI Port 2 Write Data Channel
    input[63:0]                          WDATA_2,
    input[7:0]                           WSTRB_2,
    input                                WLAST_2,
    input                                WVALID_2,
    output                               WREADY_2,
    
    // AXI Port 2 Write Response Channel
    output[7:0]                          BID_2,
    output[1:0]                          BRESP_2,
    output                               BVALID_2,
    input                                BREADY_2,
    
    // AXI Port 2 Read Address Channel
    input[7:0]                           ARID_2,
    input[31:0]                          ARADDR_2,
    input[7:0]                           ARLEN_2,
    input[2:0]                           ARSIZE_2,
    input[1:0]                           ARBURST_2,
    input                                ARLOCK_2,
    
    input                                ARVALID_2,
    output                               ARREADY_2,
    input                                ARPOISON_2,
    
    // AXI Port 2 Read Data Channel
    output[7:0]                          RID_2,
    output[63:0]                         RDATA_2,
    output[1:0]                          RRESP_2,
    output                               RLAST_2,
    output                               RVALID_2,
    input                                RREADY_2,
    
    input                                ARURGENT_2,
    output                               RAQ_PUSH_2,
    output                               RAQ_SPLIT_2,                              
    output                               WAQ_PUSH_2,
    output                               WAQ_SPLIT_2,
    // QOS
    input[3:0]                           AWQOS_0,
    input[3:0]                           ARQOS_0,
    input[3:0]                           AWQOS_1,
    input[3:0]                           ARQOS_1,
    input[3:0]                           AWQOS_2,
    input[3:0]                           ARQOS_2,
    //-----------------------------------------------
    //DDRC Low Power Interface
    //-----------------------------------------------	
    input                                CSYSREQ_0,
    output                               CSYSACK_0,
    output                               CACTIVE_0,
    input                                CSYSREQ_1,
    output                               CSYSACK_1,
    output                               CACTIVE_1,
    input                                CSYSREQ_2,
    output                               CSYSACK_2,
    output                               CACTIVE_2,
                                        
    input                                CSYSREQ_DDRC,
    output                               CSYSACK_DDRC,
    output                               CACTIVE_DDRC,
    input[2:0]                           PA_RMASK,
    input[2:0]                           PA_WMASK,

   
    //----------------------------------------------- 
    // DFI Interface 
    //-----------------------------------------------  

    output[31:0]                         DFI_ADDRESS,
    output[5:0]                          DFI_BANK,
    output[1:0]                          DFI_CAS_N,
    output[1:0]                          DFI_RAS_N,
    output[1:0]                          DFI_WE_N,
    output[1:0]                          DFI_CKE,
    output[1:0]                          DFI_CS,
    output[1:0]                          DFI_ODT,
    output[1:0]                          DFI_RESET_N,
    output[63:0]                         DFI_WRDATA,
    output[7:0]                          DFI_WRDATA_MASK,
    output[3:0]                          DFI_WRDATA_EN,
    input[63:0]                          DFI_RDDATA,
    output[3:0]                          DFI_RDDATA_EN,
    input[3:0]                           DFI_RDDATA_VALID,
    input                                DFI_CTRLUPD_ACK,          
    output                               DFI_CTRLUPD_REQ,
    output                               DFI_DRAM_CLK_DISABLE, 
    input                                DFI_INIT_COMPLETE,    
    output                               DFI_INIT_START,
    output[4:0]                          DFI_FREQUENCY,
    input                                DFI_PHYUPD_REQ,    // DFI PHY update request 
    input[1:0]                           DFI_PHYUPD_TYPE,   // DFI PHY update type 
    output                               DFI_PHYUPD_ACK,   // DFI PHY update acknowledge 
    output                               DFI_LP_REQ,         // DFI LP request
    output[3:0]                          DFI_LP_WAKEUP,     // DFI LP wakeup
    input                                DFI_LP_ACK,        // DFI LP acknowledge
    input                                PCLK,
    input                                PRESET,
    input[11:0]                          PADDR,
    input[31:0]                          PWDATA,
    input                                PWRITE,
    input                                PSEL,
    input                                PENABLE,
    output                               PREADY,
    output[31:0]                         PRDATA,
    output                               PSLVERR
    );
   //synthesis translate_off 
    ddrc_gtp_wrap  GTP_DDRC_WRAP(
    .core_ddrc_core_clk(CORE_DDRC_CORE_CLK),    
    .core_ddrc_rst     (CORE_DDRC_RST),
    .areset_0          (ARESET_0),
    .aclk_0            (ACLK_0),
    .awid_0            (AWID_0),
    .awaddr_0          (AWADDR_0),
    .awlen_0           (AWLEN_0),
    .awsize_0          (AWSIZE_0),
    .awburst_0         (AWBURST_0),
    .awlock_0          (AWLOCK_0),
    .awvalid_0         (AWVALID_0),
    .awready_0         (AWREADY_0),
    .awurgent_0        (AWURGENT_0),
    .awpoison_0        (AWPOISON_0),
    .awpoison_intr_0   (),
    .waq_push_0        (WAQ_PUSH_0),
    .waq_split_0       (WAQ_SPLIT_0),
    .wdata_0           (WDATA_0),
    .wstrb_0           (WSTRB_0),
    .wlast_0           (WLAST_0),
    .wvalid_0          (WVALID_0),
    .wready_0          (WREADY_0),
    .bid_0             (BID_0),
    .bresp_0           (BRESP_0),
    .bvalid_0          (BVALID_0),
    .bready_0          (BREADY_0),
    .arid_0            (ARID_0),
    .araddr_0          (ARADDR_0),
    .arlen_0           (ARLEN_0),
    .arsize_0          (ARSIZE_0),
    .arburst_0         (ARBURST_0),
    .arlock_0          (ARLOCK_0),
    .arvalid_0         (ARVALID_0),
    .arready_0         (ARREADY_0),
    .arpoison_0        (ARPOISON_0),
    .arpoison_intr_0   (),
    .arurgent_0        (ARURGENT_0),
    .raq_push_0        (RAQ_PUSH_0),
    .raq_split_0       (RAQ_SPLIT_0),
    .rid_0             (RID_0),
    .rdata_0           (RDATA_0),
    .rresp_0           (RRESP_0),
    .rlast_0           (RLAST_0),
    .rvalid_0          (RVALID_0),
    .rready_0          (RREADY_0),
    .areset_1          (ARESET_1),
    .aclk_1            (ACLK_1),
    .awid_1            (AWID_1),
    .awaddr_1          (AWADDR_1),
    .awlen_1           (AWLEN_1),
    .awsize_1          (AWSIZE_1),
    .awburst_1         (AWBURST_1),
    .awlock_1          (AWLOCK_1),
    .awvalid_1         (AWVALID_1),
    .awready_1         (AWREADY_1),
    .awurgent_1        (AWURGENT_1),
    .awpoison_1        (AWPOISON_1),
    .awpoison_intr_1   (),
    .waq_push_1        (WAQ_PUSH_1),
    .waq_split_1       (WAQ_SPLIT_1),
    .wdata_1           (WDATA_1),
    .wstrb_1           (WSTRB_1),
    .wlast_1           (WLAST_1),
    .wvalid_1          (WVALID_1),
    .wready_1          (WREADY_1),
    .bid_1             (BID_1),
    .bresp_1           (BRESP_1),
    .bvalid_1          (BVALID_1),
    .bready_1          (BREADY_1),
    .arid_1            (ARID_1),
    .araddr_1          (ARADDR_1),
    .arlen_1           (ARLEN_1),
    .arsize_1          (ARSIZE_1),
    .arburst_1         (ARBURST_1),
    .arlock_1          (ARLOCK_1),
    .arvalid_1         (ARVALID_1),
    .arready_1         (ARREADY_1),
    .arpoison_1        (ARPOISON_1),
    .arpoison_intr_1   (),
    .arurgent_1        (ARURGENT_1),
    .raq_push_1        (RAQ_PUSH_1),
    .raq_split_1       (RAQ_SPLIT_1),
    .rid_1             (RID_1),
    .rdata_1           (RDATA_1),
    .rresp_1           (RRESP_1),
    .rlast_1           (RLAST_1),
    .rvalid_1          (RVALID_1),
    .rready_1          (RREADY_1),
    .areset_2          (ARESET_2),
    .aclk_2            (ACLK_2),
    .awid_2            (AWID_2),
    .awaddr_2          (AWADDR_2),
    .awlen_2           (AWLEN_2),
    .awsize_2          (AWSIZE_2),
    .awburst_2         (AWBURST_2),
    .awlock_2          (AWLOCK_2),
    .awvalid_2         (AWVALID_2),
    .awready_2         (AWREADY_2),
    .awurgent_2        (AWURGENT_2),
    .awpoison_2        (AWPOISON_2),
    .awpoison_intr_2   (),
    .waq_push_2        (WAQ_PUSH_2),
    .waq_split_2       (WAQ_SPLIT_2),
    .wdata_2           (WDATA_2),
    .wstrb_2           (WSTRB_2),
    .wlast_2           (WLAST_2),
    .wvalid_2          (WVALID_2),
    .wready_2          (WREADY_2),
    .bid_2             (BID_2),
    .bresp_2           (BRESP_2),
    .bvalid_2          (BVALID_2),
    .bready_2          (BREADY_2),
    .arid_2            (ARID_2),
    .araddr_2          (ARADDR_2),
    .arlen_2           (ARLEN_2),
    .arsize_2          (ARSIZE_2),
    .arburst_2         (ARBURST_2),
    .arlock_2          (ARLOCK_2),
    .arvalid_2         (ARVALID_2),
    .arready_2         (ARREADY_2),
    .arpoison_2        (ARPOISON_2),
    .arpoison_intr_2   (),
    .arurgent_2        (ARURGENT_2),
    .raq_push_2        (RAQ_PUSH_2),
    .raq_split_2       (RAQ_SPLIT_2),
    .rid_2             (RID_2),
    .rdata_2           (RDATA_2),
    .rresp_2           (RRESP_2),
    .rlast_2           (RLAST_2),
    .rvalid_2          (RVALID_2),
    .rready_2          (RREADY_2),
    .csysreq_0          (CSYSREQ_0),
    .csysack_0          (CSYSACK_0),
    .cactive_0          (CACTIVE_0),
    .csysreq_1          (CSYSREQ_1),
    .csysack_1          (CSYSACK_1),
    .cactive_1          (CACTIVE_1),
    .csysreq_2          (CSYSREQ_2),
    .csysack_2          (CSYSACK_2),
    .cactive_2          (CACTIVE_2),
    .csysreq_ddrc       (CSYSREQ_DDRC),
    .csysack_ddrc       (CSYSACK_DDRC),
    .cactive_ddrc       (CACTIVE_DDRC),
    .pa_rmask           (PA_RMASK),
    .pa_wmask                            (PA_WMASK),
    .dfi_address                         (DFI_ADDRESS),
    .dfi_bank                            (DFI_BANK),
    .dfi_cas_n                           (DFI_CAS_N),
    .dfi_cke                             (DFI_CKE),
    .dfi_cs                              (DFI_CS),
    .dfi_odt                             (DFI_ODT),
    .dfi_ras_n                           (DFI_RAS_N),
    .dfi_reset_n                         (DFI_RESET_N),
    .dfi_we_n                            (DFI_WE_N),
    .dfi_wrdata                          (DFI_WRDATA),
    .dfi_wrdata_en                       (DFI_WRDATA_EN),
    .dfi_wrdata_mask                     (DFI_WRDATA_MASK),
    .dfi_rddata                          (DFI_RDDATA),
    .dfi_rddata_en                       (DFI_RDDATA_EN),
    .dfi_rddata_valid                    (DFI_RDDATA_VALID),
    .dfi_ctrlupd_req                     (DFI_CTRLUPD_REQ),
    .dfi_ctrlupd_ack                     (DFI_CTRLUPD_ACK),
    .dfi_dram_clk_disable                (DFI_DRAM_CLK_DISABLE),
    .dfi_init_complete                   (DFI_INIT_COMPLETE),
    .dfi_init_start                      (DFI_INIT_START),
    .dfi_frequency                       (DFI_FREQUENCY),
    .dfi_phyupd_req                      (DFI_PHYUPD_REQ),
    .dfi_phyupd_type                     (DFI_PHYUPD_TYPE),
    .dfi_phyupd_ack                      (DFI_PHYUPD_ACK),
    .dfi_lp_req                          (DFI_LP_REQ),
    .dfi_lp_wakeup                       (DFI_LP_WAKEUP),
    .dfi_lp_ack                          (DFI_LP_ACK),
    .pclk                                (PCLK),
    .preset                              (PRESET),
    .paddr                               (PADDR),
    .pwdata                              (PWDATA),
    .pwrite                              (PWRITE),
    .psel                                (PSEL),
    .penable                             (PENABLE),
    .pready                              (PREADY),
    .prdata                              (PRDATA),
    .pslverr                             (PSLVERR),
    .awqos_0                             (AWQOS_0),
    .arqos_0                             (ARQOS_0),
    .awqos_1                             (AWQOS_1),
    .arqos_1                             (ARQOS_1),
    .awqos_2                             (AWQOS_2),
    .arqos_2                             (ARQOS_2),
    .raq_wcount_0                        ()                              ,
     .raq_pop_0                          ()                               ,
     .waq_wcount_0                       ()                               ,
     .waq_pop_0                          ()                               ,
     .raq_wcount_1                       ()                               ,
     .raq_pop_1                          ()                               ,
     .waq_wcount_1                       ()                               ,
     .waq_pop_1                          ()                               ,
     .raq_wcount_2                       ()                               ,
     .raq_pop_2                          ()                               ,
     .waq_wcount_2                       ()                               ,
     .waq_pop_2                          ()                               ,
     .stat_ddrc_reg_selfref_type         ()                               ,
     .perf_hif_rd_or_wr                  ()                               ,
     .perf_hif_wr                        ()                               ,
     .perf_hif_rd                        ()                               ,
     .perf_hif_rmw                       ()                               ,
     .perf_hif_hi_pri_rd                 ()                               ,
     .perf_dfi_wr_data_cycles            ()                               ,
     .perf_dfi_rd_data_cycles            ()                               ,
     .perf_hpr_xact_when_critical        ()                               ,
     .perf_lpr_xact_when_critical        ()                               ,
     .perf_wr_xact_when_critical         ()                               ,
     .perf_op_is_activate                ()                               ,
     .perf_op_is_rd_or_wr                ()                               ,
     .perf_op_is_rd_activate             ()                               ,
     .perf_op_is_rd                      ()                               ,
     .perf_op_is_wr                      ()                               ,
     .perf_op_is_precharge               ()                               ,
     .perf_precharge_for_rdwr            ()                               ,
     .perf_precharge_for_other           ()                               ,
     .perf_rdwr_transitions              ()                               ,
     .perf_write_combine                 ()                               ,
     .perf_war_hazard                    ()                               ,
     .perf_raw_hazard                    ()                               ,
     .perf_waw_hazard                    ()                               ,
     .perf_op_is_enter_selfref           ()                               ,
     .perf_op_is_enter_powerdown         ()                               ,
     .perf_op_is_enter_deeppowerdown     ()                               ,
     .perf_selfref_mode                  ()                               ,
     .perf_op_is_refresh                 ()                               ,
     .perf_op_is_load_mode               ()                               ,
     .perf_op_is_zqcl                    ()                               ,
     .perf_op_is_zqcs                    ()                               ,
     .perf_bank                          ()                               ,
     .perf_hpr_req_with_nocredit         ()                               ,
     .perf_lpr_req_with_nocredit         ()                               ,
     .lpr_credit_cnt                     ()                               ,
     .hpr_credit_cnt                     ()                               ,
     .wr_credit_cnt                      ()                               ,
     .scanmode_n                         (1'b1)                               , 
     .scan_reset                         (1'b1)                                  
);
//synthesis translate_on	
endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_RAM16X1DP.v
//
// Functional description: simple-dual-port 16x1 distributed ram
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_RAM16X1DP
#(
    parameter [15:0] INIT = 16'h0000
) (
    output  DO,
    input   DI,
    input [3:0] RADDR, WADDR,
    input WCLK, WE
);

    reg [15:0] mem ;

    initial begin
        mem = INIT;
    end

    always @(posedge WCLK) begin
        if (WE == 1'b1) begin
            mem[WADDR] <= DI;
        end
    end

    assign DO = mem[RADDR];

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2016 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_ZEROHOLDDELAY.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
/////////////////////////////////////////////////////////////////////////////
`timescale 1 ps / 1 ps

module GTP_ZEROHOLDDELAY #(
parameter        ZHOLD_SET  = "NODELAY"    //  "NODELAY","100ps","200ps","300ps","400ps","500ps","600ps","700ps","800ps","900ps","1000ps","1100ps","1200ps","1300ps","1400ps","1500ps"
)(
output      DO,
input       DI
); /* synthesis syn_black_box */ 

//synthesis translate_off
///////////////////////////////////////////////////////////////////////////

reg  [14:0] therm_code;
wire [15:0]  data;


initial begin
    if(ZHOLD_SET != "NODELAY" && ZHOLD_SET != "100ps" && ZHOLD_SET != "200ps" && ZHOLD_SET != "300ps" && ZHOLD_SET != "400ps" && ZHOLD_SET != "500ps" && ZHOLD_SET != "600ps" && ZHOLD_SET != "700ps" && ZHOLD_SET != "800ps" && ZHOLD_SET != "900ps" && ZHOLD_SET != "1000ps" && ZHOLD_SET != "1100ps" && ZHOLD_SET != "1200ps" && ZHOLD_SET != "1300ps" && ZHOLD_SET != "1400ps" && ZHOLD_SET != "1500ps")    //  16 kinds
    begin
      $display("Error: Illegal setting ZHOLD_SET of %s",ZHOLD_SET);
      $finish;
    end
end             

initial begin
    case(ZHOLD_SET)
    "NODELAY": therm_code = 15'h0000;
    "100ps"  : therm_code = 15'h0001;
    "200ps"  : therm_code = 15'h0003;
    "300ps"  : therm_code = 15'h0007;
    "400ps"  : therm_code = 15'h000F;
    "500ps"  : therm_code = 15'h001F;
    "600ps"  : therm_code = 15'h003F;
    "700ps"  : therm_code = 15'h007F;
    "800ps"  : therm_code = 15'h00FF;
    "900ps"  : therm_code = 15'h01FF;
    "1000ps" : therm_code = 15'h03FF;
    "1100ps" : therm_code = 15'h07FF;
    "1200ps" : therm_code = 15'h0FFF;
    "1300ps" : therm_code = 15'h1FFF;
    "1400ps" : therm_code = 15'h3FFF;
    "1500ps" : therm_code = 15'h7FFF;
    default  : therm_code = 15'h0000;
    endcase
end

assign   data[0] = DI;

genvar i;
generate 
    for (i=1; i<=15; i=i+1)
    begin
       assign #100  data[i]  = data[i-1];
    end
endgenerate

assign DO  =    (therm_code  == 15'h0000) ? data[0]   : 
                (therm_code  == 15'h0001) ? data[1]   :
                (therm_code  == 15'h0003) ? data[2]   : 
                (therm_code  == 15'h0007) ? data[3]   : 
                (therm_code  == 15'h000F) ? data[4]   :
                (therm_code  == 15'h001F) ? data[5]   :
                (therm_code  == 15'h003F) ? data[6]   : 
                (therm_code  == 15'h007F) ? data[7]   :
                (therm_code  == 15'h00FF) ? data[8]   :
                (therm_code  == 15'h01FF) ? data[9]   : 
                (therm_code  == 15'h03FF) ? data[10]  :
                (therm_code  == 15'h07FF) ? data[11]  :
                (therm_code  == 15'h0FFF) ? data[12]  : 
                (therm_code  == 15'h1FFF) ? data[13]  :
                (therm_code  == 15'h3FFF) ? data[14]  :  data[15];

//synthesis translate_on 

endmodule                                                                                                    




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_DLATCH.v
//
// Functional description: D-type latch
//
// Parameter description:
//      INIT: init value
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_DLATCH
#(
    parameter GRS_EN = "TRUE",
    parameter INIT = 1'b0
) (
    output reg Q,
    input wire D,
    input wire G
);

    wire grs_n;
    wire RS;

    tri1 grsnet = GRS_INST.GRSNET;
    assign grs_n=(GRS_EN=="TRUE")?grsnet:1'b1;
 
    not (RS, grs_n);

    initial Q = 1'bx;

    always @(D or G or RS) begin
        if (RS)
            Q <= 1'b0;
        else if (G)
            Q <= D;
    end

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_START.v
//
// Functional description: startup Logic Control Circuit
//
// Parameter description:
//      
//
// Port description:
//      
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps 

module GTP_START
(
    input        CLK    ,          //start signals
    input tri0   GOE,
    input tri0   GRS_N  ,
    input tri0   GWE   
);

wire        GOUTEN     ;
wire        GRSN       ;
wire        GWEN       ;

assign GOUTEN = GOE;
assign GRSN   = GRS_N  ;
assign GWEN   = GWE  ;


endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_LUT4.v
//
// Functional description: 4-input Look-Up-Table
//
// Parameter description:
//      INIT: init value
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_LUT4
#(
    parameter [15:0] INIT = 16'h0000
) (
    output wire Z,
    input wire I0, I1, I2, I3
);

    wire x3, x2, x1, x0;

    INT_LUTMUX4_UDP (x3, I1, I0, INIT[15], INIT[14], INIT[13], INIT[12]);
    INT_LUTMUX4_UDP (x2, I1, I0, INIT[11], INIT[10], INIT[9], INIT[8]);
    INT_LUTMUX4_UDP (x1, I1, I0, INIT[7], INIT[6], INIT[5], INIT[4]);
    INT_LUTMUX4_UDP (x0, I1, I0, INIT[3], INIT[2], INIT[1], INIT[0]);
    INT_LUTMUX4_UDP (Z, I3, I2, x3, x2, x1, x0);

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_IOBUF_TX_MIPI.v
//
// Functional description: Input Buffer For MIPI Protocol
//
// Parameter description:
//
// Port description:
//
// Revision:
//    05/18/18 - Initial version.
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_IOBUF_TX_MIPI 
#(
  parameter IOSTANDARD  ="DEFAULT",
  parameter SLEW_RATE = "SLOW",
  parameter DRIVE_STRENGTH = "6",
  parameter TERM_DIFF = "ON"
) (
    output wire O_LP,
    output wire OB_LP,
    inout  wire IO,
    inout  wire IOB,
    input  wire I_HS,
    input  wire I_LP,
    input  wire IB_LP,
    input  wire T,
    input  wire TB,
    input  wire M
);

    reg [23:0]  STR_I, STR_IB;
    reg         O_LP_reg;
    reg         OB_LP_reg; 

    wire  I;

    assign I = (M == 1'b1) ? I_HS : I_LP;
     
    always @(*)
      begin
         $sformat(STR_I, "%v", IO);
         $sformat(STR_IB, "%v", IOB);
      end

    initial   begin
         case(IOSTANDARD) 
           "MIPI", "DEFAULT" : ;
           default:  begin
             $display("Attribute ERROR: Illegal IOSTANDARD value %s.", IOSTANDARD);
             $finish;
             end
         endcase

    case (TERM_DIFF)
    "ON", "OFF" :;
    default : begin
           $display("Attribute Syntax Error : The attribute TERM_DIFF on instance %m is set to %s.", TERM_DIFF);
           $finish;
              end
    endcase

    case (SLEW_RATE)
    "FAST", "SLOW":;
    default : begin
           $display("Attribute Syntax Error : The attribute SLEW_RATE on instance %m is set to %s.", SLEW_RATE);
           $finish;
              end
    endcase

    case (DRIVE_STRENGTH)
    "2", "4", "6" :;
    default : begin
           $display("Attribute Syntax Error : The attribute DRIVE_STRENGTH on GTP_IOBUF_TX_MIPI instance %m is set to %s.", DRIVE_STRENGTH);
           $finish;
              end
    endcase

     end

//    assign O_LP = O_LP_reg;
//    assign OB_LP = OB_LP_reg;


    assign TS_HS = !T && M;
    assign TS_LP = T || M;
    assign TS_LP_B = TB || M;

//high speed output

    bufif1 bufd_hs  (IO, I, TS_HS);
    notif1 bufdb_hs (IOB, I, TS_HS);

//low power output

    bufif0 buf_lp   (IO, I, TS_LP);
    bufif0 bufb_lp  (IOB, IB_LP, TS_LP_B);
   
//lower power input

    buf ibuf_lp (O_LP, O_LP_reg);
    buf ibufb_lp (OB_LP, OB_LP_reg);

    always @(*)
       if(M == 1'b0) 
             if(T == 1'b1 && TB == 1'b1)
                begin
                  O_LP_reg  <= IO;
                  OB_LP_reg <= IOB;
                end
             else if ( T == 1'b0 && TB == 1'b0 )
                begin
                   O_LP_reg <= 1'b1;
                   OB_LP_reg <= 1'b1;
                end 
             else
                begin
                   O_LP_reg  <= 1'bx;
                   OB_LP_reg <= 1'bx;
                end
       else if ( M == 1'b1 )
            begin
               O_LP_reg  <= 1'b1;
               OB_LP_reg <= 1'b1;
            end
       else
            begin
              O_LP_reg   <= 1'bx;
              OB_LP_reg  <= 1'bx; 
            end
    
endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_PREADD_MULTADDSUM9.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

//P = (A0*(B0+/-C0) +/- A1*(B1 +/-C1)) +- (A2*(B2+/-C2) +/- A3*(B3+/-C3))
`timescale 1 ns / 1 ps

module GTP_PREADD_MULTADDSUM9  #(
    parameter GRS_EN             = "TRUE", //"TRUE"; "FALSE"
    parameter SYNC_RST           = "FALSE", //"TRUE"; "FALSE"
    parameter INREG_EN           = "FALSE",  //"TRUE"; "FALSE"
    parameter PREREG_EN          = "FALSE",  //"TRUE"; "FALSE"
    parameter PIPEREG_EN         = "FALSE",  //"TRUE"; "FALSE"
    parameter OUTREG_EN          = "FALSE",   //"TRUE"; "FALSE"
    parameter ADDSUB_OP          = 2'b00 ,
    parameter SUM_ADDSUB_OP      = 0 ,
    parameter DYN_ADDSUB_OP      = 2'b11,
    parameter DYN_SUM_ADDSUB_OP  = 1
)(
    output  [20-1:0] P,
    input   CE,
    input   RST,
    input   CLK,
    input   [1:0] A_SIGNED,
    input   [9-1:0] A0,
    input   [9-1:0] A1,
    input   [9-1:0] A2,
    input   [9-1:0] A3,
    input   [1:0] B_SIGNED,
    input   [1:0] C_SIGNED,
    input   [8-1:0] B0,
    input   [8-1:0] B1,
    input   [8-1:0] B2,
    input   [8-1:0] B3,
    input   [8-1:0] C0,
    input   [8-1:0] C1,
    input   [8-1:0] C2,
    input   [8-1:0] C3,
    input   [3:0] PREADDSUB,
    input   [1:0] ADDSUB,
    input   SUM_ADDSUB
);

    INT_PREADD_MULTADDSUM #(
        . GRS_EN(GRS_EN),    
        . SYNC_RST(SYNC_RST),  
        . INREG_EN(INREG_EN),  
        . PREREG_EN(PREREG_EN),  
        . PIPEREG_EN(PIPEREG_EN),
        . OUTREG_EN(OUTREG_EN), 
        . ADDSUB_OP01(ADDSUB_OP[0]),  
        . ADDSUB_OP23(ADDSUB_OP[1]),  
        . ADDSUBSUM_OP(SUM_ADDSUB_OP), 
        . DYN_OP_SEL0(DYN_ADDSUB_OP[0]),
        . DYN_OP_SEL1(DYN_ADDSUB_OP[1]),
        . DYN_OP_SEL2(DYN_SUM_ADDSUB_OP),
        . ASIZE(9),
        . BSIZE(8)
    ) U_INT_PREADD_MULTADDSUM (
        . CE(CE),
        . RST(RST),
        . CLK(CLK),
        . A_SIGNED01(A_SIGNED[0]),
        . A_SIGNED23(A_SIGNED[1]),
        . A0(A0),
        . A1(A1),
        . A2(A2),
        . A3(A3),
        . B_SIGNED01(B_SIGNED[0]),
        . B_SIGNED23(B_SIGNED[1]), 
        . C_SIGNED01(C_SIGNED[0]),
        . C_SIGNED23(C_SIGNED[1]), 
        . B0(B0),
        . B1(B1),
        . B2(B2),
        . B3(B3),
        . C0(C0),
        . C1(C1),
        . C2(C2),
        . C3(C3),
        . PREADDSUB01(PREADDSUB[1:0]),
        . PREADDSUB23(PREADDSUB[3:2]),
        . ADDSUB01(ADDSUB[0]),
        . ADDSUB23(ADDSUB[1]),
        . ADDSUBSUM(SUM_ADDSUB),
        . P(P)
    );               

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_BUF.v
//
// Functional description: 1-bit Buffer
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_BUF
(
    output wire Z,
    input wire I
);

    buf (Z, I);

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2016 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General Technology Primitive
// Filename: GTP_OSC_E1.v
//
// Functional description: oscillator
//
// Parameter description:
// CLK_DIV:    CLKOUT frequency setting( f = 200MHz/CLK_DIV )[f=200MHz/128, when CLK_DIV=0]
//
// Port description:
// inputs:
// EN:           OSC enable
// RST_N:        Reset clock divider
//
// outputs:
// CLKOUT:    100MHz(default)
//
// Revision: V1.0
//
//////////////////////////////////////////////////////////////////////////////
`timescale 1ns/1ps

module GTP_OSC_E1
   #(
     parameter integer CLK_DIV = 2
     )
    (
     output CLKOUT,
    
     input  EN,
     input  RST_N
     )/* synthesis syn_black_box */;

    //synthesis translate_off
    wire    rst_wire;
    wire    oscen_wire;
    reg     clk_400_reg; // intrinsic frequency
    reg [6:0] div_reg;
    reg [6:0] count_reg;
    reg       clk_user_reg;
    reg       rst_reg;

    initial 
    begin
        // parameter check
        if ( (CLK_DIV >= 0) && (CLK_DIV <= 127) )
        begin
            div_reg = CLK_DIV;
        end
        else
        begin
            $display ("GTP_OSC_E1 error: illegal setting for CLK_DIV(0 ~ 127)");
        end

        // analog //
        clk_400_reg = 1'b0;

        // divider //
        count_reg = 7'b0000000;
        clk_user_reg = 1'b0;
        rst_reg = 1'b0;
    end
    
    assign rst_wire = !RST_N || !EN;
    assign oscen_wire = EN;
    assign CLKOUT = clk_user_reg;
    
    // osc_analog //
    always
    begin
        wait (oscen_wire == 1'b1)
           begin
               clk_400_reg = 1'b0;
               #1.25;
               clk_400_reg = 1'b1;
               #1.25;
           end
    end

    always
    begin
        wait (oscen_wire != 1'b1)
           begin
               force clk_400_reg = 1'b0;
               #2 release clk_400_reg;
           end
    end
    // end of osc_analog //
    
    // osc_divider_128 //
    always @ (posedge clk_400_reg or posedge rst_wire)
    begin
        if (rst_wire)
        begin
            clk_user_reg <= 1'b0;
            count_reg <= 7'b000_0000;
            rst_reg <= 1'b1;
        end
        else if (rst_reg)
        begin
            rst_reg <= 1'b0;
            clk_user_reg <= 1'b1;
            count_reg <= 7'b000_0000;
        end
        else if (count_reg == div_reg-7'b1)
        begin
            clk_user_reg <= ~clk_user_reg;
            count_reg <= 7'b000000;
        end
        else
        begin
            clk_user_reg <= clk_user_reg;
            count_reg <= count_reg + 1'b1;
        end
    end
    // end of osc_divider_128 //
    
    //synthesis translate_on
endmodule // GTP_OSC_E1



//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_LUT5CARRY.v
//
// Functional description: LUT5 and CARRY
//
// Parameter description:
//      ID_TO_LUT   : 'TRUE'  ID to LUT.I0
//                    'FALSE' I0 to LUT.I0
//      CIN_TO_LUT  : 'TRUE' CIN to LUT.I0
//                    'FALSE' I0 to LUT.I0
//      I4_TO_CARRY : 'TRUE'  I4 to I0
//                    'FALSE' LUT to CARRY
//      I4_TO_LUT   : 'TRUE'
//                    'FALSE'
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_LUT5CARRY
#(
    parameter [31:0] INIT = 32'h0000_0000,
    parameter ID_TO_LUT = "FALSE",
    parameter CIN_TO_LUT = "TRUE",
    parameter I4_TO_CARRY = "TRUE",
    parameter I4_TO_LUT = "FALSE"
) (
    output COUT, Z,
    input CIN, I0, ID, I1, I2, I3, I4
);

    wire i4, i3, i2, i1, ci, ci0, i00, i10;
    wire x7, x6, x5, x4, x3, x2, x1, x0;
    wire z, co, y0, y1;

    initial
    begin
        if (ID_TO_LUT != "TRUE" && ID_TO_LUT != "FALSE")
        begin
            $display("ERROR: The attribute ID_TO_LUT on instance %m is %s. Legal values are TRUE or FALSE.", ID_TO_LUT);
            $finish;
        end

        if (I4_TO_LUT != "TRUE" && I4_TO_LUT != "FALSE")
        begin
            $display("ERROR: The attribute I4_TO_LUT on instance %m is %s. Legal values are TRUE or FALSE.", I4_TO_LUT);
            $finish;
        end

        if (CIN_TO_LUT != "TRUE" && CIN_TO_LUT != "FALSE")
        begin
            $display("ERROR: The attribute CIN_TO_LUT on instance %m is %s. Legal values are TRUE or FALSE.", CIN_TO_LUT);
            $finish;
        end

        if (I4_TO_CARRY != "TRUE" && I4_TO_CARRY != "FALSE")
        begin
            $display("ERROR: The attribute I4_TO_CARRY on instance %m is %s. Legal values are TRUE or FALSE.", I4_TO_CARRY);
            $finish;
        end
    end

    buf (i3, I3);
    buf (i2, I2);
    buf (i1, I1);
    buf (ci, CIN);
    assign i00 = (ID_TO_LUT == "FALSE") ? I0 : ID;
    assign i10 = (CIN_TO_LUT == "TRUE") ? CIN : I0;
    assign ci0 = (I4_TO_CARRY == "TRUE") ? I4 : y1;
    assign i4  = (I4_TO_LUT == "FALSE") ? 1'b1 : I4;

    INT_LUTMUX4_UDP (x7, i1, i10, INIT[31], INIT[30], INIT[29], INIT[28]);
    INT_LUTMUX4_UDP (x6, i1, i10, INIT[27], INIT[26], INIT[25], INIT[24]);
    INT_LUTMUX4_UDP (x5, i1, i10, INIT[23], INIT[22], INIT[21], INIT[20]);
    INT_LUTMUX4_UDP (x4, i1, i10, INIT[19], INIT[18], INIT[17], INIT[16]);
    INT_LUTMUX4_UDP (x3, i1, i00, INIT[15], INIT[14], INIT[13], INIT[12]);
    INT_LUTMUX4_UDP (x2, i1, i00, INIT[11], INIT[10], INIT[9], INIT[8]);
    INT_LUTMUX4_UDP (x1, i1, i00, INIT[7], INIT[6], INIT[5], INIT[4]);
    INT_LUTMUX4_UDP (x0, i1, i00, INIT[3], INIT[2], INIT[1], INIT[0]);

    INT_LUTMUX4_UDP (y1, i3, i2, x7, x6, x5, x4);
    INT_LUTMUX4_UDP (y0, i3, i2, x3, x2, x1, x0);
    INT_LUTMUX2_UDP (co, y0, ci, ci0);
    INT_LUTMUX2_UDP (z, i4, y1, y0);

    buf (Z, z);
    buf (COUT, co);

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2016 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_CLKBUFX.v
//
// Functional description: CLOCK BUFFER
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_CLKBUFX
(
    output CLKOUT,
    input CLKIN
);

//synthesis translate_off

    assign CLKOUT = CLKIN;

//synthesis translate_on
endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_FLASHIF.v
//
// Functional description: FLASHIF for user
//
// Parameter description:
//      
//
// Port description:
//      
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////
`timescale 1 ns / 1 ps
module   GTP_FLASHIF  (
input             EN_N,
input             CLK ,
input             CS_N,
input    [3:0]    DIN ,
input    [2:0]    DOUT_EN_N ,
output   [3:0]    DOUT 
);


endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_DCC.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_DCC #(
parameter GRS_EN = "TRUE",  //FALSE; TRUE;
parameter SAMPLE_CLKDIV_FACTOR = "2" //"1"; "2"; "3.5"; "4"; "5"; 
)(
output SAMPLE_CLKOUT,
output PROBE_CLKOUT,
output SAMPLE_CLKDIVOUT,
input [2:0] CLKOUT_CTRL,
input  CLKIN0,
input  CLKIN1,
input RST,
input [1:0] CLK0_SEL,
input [1:0] CLK1_SEL,
input [7:0] DELAY_STEP0,
input [7:0] DELAY_STEP1
)/* synthesis syn_black_box */;

//synthesis translate_off
reg CLK0_reg;
reg CLK1_reg;
reg [1:0] DCC_CLKCTRL_b0_clk0_d;
reg [1:0] DCC_CLKCTRL_b0_clk1_d;
reg DCC_CLKCTRL_b2_d;
reg sample_clk_reg;
reg DCC_CLKCTRL_b1_d;
reg probe_clk_reg;
reg [2:0] cnt;
reg [3:0] cnt2;
reg CLKI_div2;
reg CLKI_DIV_reg;
reg CLKI_DIV_reg_neg;
reg [3:0] start_d;
reg rstn_dly;

initial 
begin
// parameter check
    if ((GRS_EN == "TRUE")  || (GRS_EN == "FALSE")) begin
    end
   else
       $display (" GTP_DCC error: illegal setting for GRS_EN"); 
   
    if ((SAMPLE_CLKDIV_FACTOR == "1") || (SAMPLE_CLKDIV_FACTOR == "2")  || (SAMPLE_CLKDIV_FACTOR == "3.5") || (SAMPLE_CLKDIV_FACTOR == "4") || (SAMPLE_CLKDIV_FACTOR == "5")) 
    begin
    end
    else
        $display (" GTP_DCC error: illegal setting for SAMPLE_CLKDIV_FACTOR");
    CLK0_reg  = 0;
    CLK1_reg  = 0;
    DCC_CLKCTRL_b0_clk0_d  = 0;
    DCC_CLKCTRL_b0_clk1_d  = 0;
    DCC_CLKCTRL_b2_d  = 0;
    sample_clk_reg  = 0;
    DCC_CLKCTRL_b1_d  = 0;
    probe_clk_reg  = 0;
    cnt  = 0;
    cnt2              = 0;
    CLKI_div2         = 0;
    CLKI_DIV_reg      = 0;
    CLKI_DIV_reg_neg  = 0;
    start_d = 0;
    rstn_dly = 0;
end

assign global_rstn = (GRS_EN == "TRUE") ? GRS_INST.GRSNET : 1'b1;
assign local_rstn =  ~RST;

always @(CLK0_SEL[1:0] or CLKIN0 or CLKIN1) 
begin
    case (CLK0_SEL[1:0])
        2'd0: CLK0_reg = CLKIN0;
        2'd1: CLK0_reg = CLKIN1;
        2'd2: CLK0_reg = ~ CLKIN0;
        2'd3: CLK0_reg = ~ CLKIN1;
    endcase
end

//
wire [255:0] clk0_delay_chain;
assign clk0_delay_chain[0] = CLK0_reg;
genvar gen_i;
generate  
    for(gen_i=1;gen_i<256;gen_i=gen_i+1) 
    begin
        assign #0.025 clk0_delay_chain[gen_i] =  clk0_delay_chain[gen_i-1];
    end
endgenerate

assign clk0_comb = clk0_delay_chain[DELAY_STEP0];

always @(CLK1_SEL[1:0] or CLKIN0 or CLKIN1) 
begin
    case (CLK1_SEL[1:0])
        2'd0: CLK1_reg = CLKIN0;
        2'd1: CLK1_reg = CLKIN1;
        2'd2: CLK1_reg = ~ CLKIN0;
        2'd3: CLK1_reg = ~ CLKIN1;
    endcase
end

wire [255:0] clk1_delay_chain;
assign clk1_delay_chain[0] = CLK1_reg;
genvar gen_j;
generate  
    for(gen_j=1;gen_j<256;gen_j=gen_j+1) 
    begin
        assign #0.025 clk1_delay_chain[gen_j] =  clk1_delay_chain[gen_j-1];
    end
endgenerate

assign clk1_comb = clk1_delay_chain[DELAY_STEP1];

always @(negedge clk0_comb or negedge global_rstn or negedge local_rstn)
begin
    if (!global_rstn)
        DCC_CLKCTRL_b0_clk0_d <= 0;
    else if (!local_rstn)
        DCC_CLKCTRL_b0_clk0_d <= 0;
    else   
        DCC_CLKCTRL_b0_clk0_d <= {DCC_CLKCTRL_b0_clk0_d[0], CLKOUT_CTRL[0]};
end

always @(negedge clk1_comb or negedge global_rstn or negedge local_rstn)
begin
    if (!global_rstn)
        DCC_CLKCTRL_b0_clk1_d <= 0;
    else if (!local_rstn)
        DCC_CLKCTRL_b0_clk1_d <= 0;
    else   
        DCC_CLKCTRL_b0_clk1_d <= {DCC_CLKCTRL_b0_clk1_d[0], CLKOUT_CTRL[0]};      
end

assign switch_clk = ~ ((~ (DCC_CLKCTRL_b0_clk0_d[1] & DCC_CLKCTRL_b0_clk1_d[1])) & (~ (clk0_comb | clk1_comb)));

always @(negedge switch_clk or negedge global_rstn or negedge local_rstn)
begin
    if (!global_rstn)
        DCC_CLKCTRL_b2_d <= 0;
    else if (!local_rstn)
        DCC_CLKCTRL_b2_d <= 0;
    else
        DCC_CLKCTRL_b2_d <= CLKOUT_CTRL[2];
end

always @(*) 
begin
    if (DCC_CLKCTRL_b2_d)
        sample_clk_reg = clk1_comb;
    else
        sample_clk_reg = clk0_comb;
end      

always @(negedge switch_clk or negedge global_rstn or negedge local_rstn)
begin
    if (!global_rstn)
        DCC_CLKCTRL_b1_d <= 0;
    else if (!local_rstn)
        DCC_CLKCTRL_b1_d <= 0;
    else
        DCC_CLKCTRL_b1_d <= CLKOUT_CTRL[1];
end

always @(*) 
begin
    if (DCC_CLKCTRL_b1_d)
        probe_clk_reg = clk0_comb;
    else
        probe_clk_reg = clk1_comb;
end    

always @(negedge sample_clk_reg)
begin
    if (!global_rstn)
        start_d[0] <= 0;
    else if (!local_rstn)
        start_d[0] <= 0;
    else
        start_d[0] <= 1;
end

always @(negedge sample_clk_reg)
begin
    start_d[3:1] <= start_d[2:0];
end

assign SAMPLE_CLKOUT = sample_clk_reg & start_d[3];
assign PROBE_CLKOUT = probe_clk_reg & start_d[3];


always @(posedge SAMPLE_CLKOUT or negedge start_d[3])
begin
    if (!start_d[3])
        rstn_dly <= 0;
    else
        rstn_dly <= 1'b1;
end

always @(posedge SAMPLE_CLKOUT or negedge rstn_dly)
begin
    if (!rstn_dly)
        CLKI_div2 <= 0;
    else
        CLKI_div2 <= ~ CLKI_div2;
end

always @(posedge SAMPLE_CLKOUT or negedge rstn_dly)
begin
    if (!rstn_dly)
        cnt2 <= 0;
    else if ((SAMPLE_CLKDIV_FACTOR == "3.5") && (cnt2 == 6))
        cnt2 <= 0;
    else if ((SAMPLE_CLKDIV_FACTOR == "4") && (cnt2 == 7))
        cnt2 <= 0;
    else if ((SAMPLE_CLKDIV_FACTOR == "5") && (cnt2 == 9))
        cnt2 <= 0;
    else   
        cnt2 <= cnt2 + 1;
end
always @(posedge SAMPLE_CLKOUT or negedge rstn_dly)
begin
    if (!rstn_dly)
        CLKI_DIV_reg <= 1'b0;
    else if (SAMPLE_CLKDIV_FACTOR == "3.5") 
    begin
        if (cnt2 == 0)
            CLKI_DIV_reg <= 1'b1;
        else if (cnt2 == 2)   
            CLKI_DIV_reg <= 1'b0;
    end      
    else if (SAMPLE_CLKDIV_FACTOR == "4") 
    begin
        if (cnt2 == 0)
            CLKI_DIV_reg <= 1'b1;
        else if (cnt2 == 2)   
            CLKI_DIV_reg <= 1'b0;
        else if (cnt2 == 4)   
            CLKI_DIV_reg <= 1'b1;
        else if (cnt2 == 6)
            CLKI_DIV_reg <= 1'b0;      
    end
    else if (SAMPLE_CLKDIV_FACTOR == "5") 
    begin
        if (cnt2 == 0)
            CLKI_DIV_reg <= 1'b1;
        else if (cnt2 == 3)   
            CLKI_DIV_reg <= 1'b0;
        else if (cnt2 == 5)   
            CLKI_DIV_reg <= 1'b1;
        else if (cnt2 == 8)
            CLKI_DIV_reg <= 1'b0;          
    end        
end

always @(negedge SAMPLE_CLKOUT or negedge rstn_dly)
begin
    if (!rstn_dly)
        CLKI_DIV_reg_neg <= 1'b0;     
    else if (SAMPLE_CLKDIV_FACTOR == "3.5") 
    begin
        if (cnt2 == 4)
            CLKI_DIV_reg_neg <= 1'b1;
        else if (cnt2 == 6)   
            CLKI_DIV_reg_neg <= 1'b0;
    end               
end
  
assign SAMPLE_CLKDIVOUT = (SAMPLE_CLKDIV_FACTOR == "1") ? SAMPLE_CLKOUT : ((SAMPLE_CLKDIV_FACTOR == "2") ? CLKI_div2 : (CLKI_DIV_reg_neg | CLKI_DIV_reg));   
     
//synthesis translate_on

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_MUX2LUT6.v
//
// Functional description: 2-to-1 MUX to generate LUT6 func
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_MUX2LUT6
(
    output wire Z,
    input wire I0, I1, S
);

    INT_LUTMUX2_UDP (Z, S, I1, I0);

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_INBUFG.v
//
// Functional description: Input Clock Buffer
//
// Parameter description:
//
// Port description:
//
// Revision:
//    06/18/14 - Initial version.
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_INBUFG #(
    parameter IOSTANDARD = "DEFAULT",
    parameter TERM_DDR = "ON"
)(
    output O,
    input I
) /* synthesis syn_black_box */ ;

  
  initial begin
    case (IOSTANDARD)
    "LVCMOS33", "LVCMOS25", "LVCMOS18", "LVCMOS15", "LVCMOS12", "SSTL25_I", "SSTL25_II", "SSTL18_I", "SSTL18_II", "SSTL15_I", "SSTL15_II", "HSTL18_I", "HSTL18_II", "HSTL15_I", "SSTL15_I_CAL", "SSTL15_II_CAL", "HSTL15_I_CAL", "DEFAULT" :;
    default : begin
           $display("Attribute Syntax Error : The attribute IOSTANDARD on GTP_INBUFG instance %m is set to %s.", IOSTANDARD);
           $finish;
              end
    endcase

    case (TERM_DDR)
    "ON", "OFF" :;
    default : begin
           $display("Attribute Syntax Error : The attribute TERM_DDR on GTP_INBUFG instance %m is set to %s.", TERM_DDR);
           $finish;
              end
    endcase
    end

    buf (O, I);

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2016 PANGO MICROSYSTEMS, INC
// ALL RIGHTS REVERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
//Library:
//FileName:
//
//Functional description:
//GTP for HSSTLP_LANE of PGL2 HSSTLP.
//Parameter description:
//
//Port description:
//
//Author:Gan Linghao
//Revision:
//  2019/08/28: Initial Version.
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1ns/1ps 
module GTP_HSSTLP_LANE
#(
    parameter    integer    MUX_BIAS = 2,//Only listed, default value:3'b010
    parameter    integer    PD_CLK = 0,//Only listed, default value:1'b0
    parameter    integer    REG_SYNC = 0,
    parameter    integer    REG_SYNC_OW = 0,
    parameter    integer    PLL_LOCK_OW = 0,
    parameter    integer    PLL_LOCK_OW_EN = 0,

    //pcs
    parameter    integer    PCS_SLAVE = 0,//Altered in 2019.12.05, should be configured by user, software only checks corresponding connection of clock

    parameter               PCS_BYPASS_WORD_ALIGN = "FALSE",          
    parameter               PCS_BYPASS_DENC = "FALSE",           
    parameter               PCS_BYPASS_BONDING = "FALSE", 
    parameter               PCS_BYPASS_CTC = "FALSE", 
    parameter               PCS_BYPASS_GEAR = "FALSE", 
    parameter               PCS_BYPASS_BRIDGE = "FALSE", 
    parameter               PCS_BYPASS_BRIDGE_FIFO = "FALSE", 
    parameter               PCS_DATA_MODE = "X8", 
    parameter               PCS_RX_POLARITY_INV = "DELAY", 
    parameter               PCS_ALIGN_MODE = "1GB", 
    parameter               PCS_SAMP_16B = "X20",          
    parameter               PCS_FARLP_PWR_REDUCTION = "FALSE",           
    parameter    integer    PCS_COMMA_REG0 = 0, 
    parameter    integer    PCS_COMMA_MASK = 0, 
    parameter               PCS_CEB_MODE = "10GB", 
    parameter               PCS_CTC_MODE = "1SKIP", 
    parameter    integer    PCS_A_REG = 0, 
    parameter               PCS_GE_AUTO_EN = "FALSE", 
    parameter    integer    PCS_SKIP_REG0 = 0, 
    parameter    integer    PCS_SKIP_REG1 = 0, 
    parameter    integer    PCS_SKIP_REG2 = 0,          
    parameter    integer    PCS_SKIP_REG3 = 0,           
    parameter               PCS_DEC_DUAL = "FALSE", 
    parameter               PCS_SPLIT = "FALSE", 
    parameter               PCS_FIFOFLAG_CTC = "FALSE", 
    parameter               PCS_COMMA_DET_MODE = "COMMA_PATTERN", 
    parameter               PCS_ERRDETECT_SILENCE = "FALSE", 
    parameter               PCS_PMA_RCLK_POLINV = "PMA_RCLK", 
    parameter               PCS_PCS_RCLK_SEL = "PMA_RCLK", 
    parameter               PCS_CB_RCLK_SEL = "PMA_RCLK", 
    parameter               PCS_AFTER_CTC_RCLK_SEL = "PMA_RCLK",           
    parameter               PCS_RCLK_POLINV = "RCLK", 
    parameter               PCS_BRIDGE_RCLK_SEL = "PMA_RCLK", 
    parameter               PCS_PCS_RCLK_EN = "FALSE",
    parameter               PCS_CB_RCLK_EN = "FALSE",
    parameter               PCS_AFTER_CTC_RCLK_EN = "FALSE",
    parameter               PCS_AFTER_CTC_RCLK_EN_GB = "FALSE",
    parameter               PCS_PCS_RX_RSTN = "FALSE",
    parameter               PCS_PCIE_SLAVE = "MASTER",
    parameter               PCS_RX_64B66B_67B = "NORMAL",
    parameter               PCS_RX_BRIDGE_CLK_POLINV = "RX_BRIDGE_CLK",
    parameter               PCS_PCS_CB_RSTN = "FALSE",
    parameter               PCS_TX_BRIDGE_GEAR_SEL = "FALSE",
    parameter               PCS_TX_BYPASS_BRIDGE_UINT = "FALSE",
    parameter               PCS_TX_BYPASS_BRIDGE_FIFO = "FALSE",
    parameter               PCS_TX_BYPASS_GEAR = "FALSE",
    parameter               PCS_TX_BYPASS_ENC = "FALSE",
    parameter               PCS_TX_BYPASS_BIT_SLIP = "FALSE",
    parameter               PCS_TX_GEAR_SPLIT = "FALSE",
    parameter               PCS_TX_DRIVE_REG_MODE = "NO_CHANGE",
    parameter    integer    PCS_TX_BIT_SLIP_CYCLES = 0,
    parameter               PCS_INT_TX_MASK_0 = "FALSE",
    parameter               PCS_INT_TX_MASK_1 = "FALSE",
    parameter               PCS_INT_TX_MASK_2 = "FALSE",
    parameter               PCS_INT_TX_CLR_0 = "FALSE",
    parameter               PCS_INT_TX_CLR_1 = "FALSE",
    parameter               PCS_INT_TX_CLR_2 = "FALSE",
    parameter               PCS_TX_PMA_TCLK_POLINV = "PMA_TCLK",
    parameter               PCS_TX_PCS_CLK_EN_SEL = "FALSE",
    parameter               PCS_TX_BRIDGE_TCLK_SEL = "TCLK",
    parameter               PCS_TX_TCLK_POLINV = "TCLK",
    parameter               PCS_PCS_TCLK_SEL= "PMA_TCLK",
    parameter               PCS_TX_PCS_TX_RSTN = "FALSE",
    parameter               PCS_TX_SLAVE = "MASTER",
    parameter               PCS_TX_GEAR_CLK_EN_SEL = "FALSE",
    parameter               PCS_DATA_WIDTH_MODE = "X20",
    parameter               PCS_TX_64B66B_67B = "NORMAL",
    parameter               PCS_GEAR_TCLK_SEL = "PMA_TCLK",
    parameter               PCS_TX_TCLK2FABRIC_SEL = "FALSE",
    parameter               PCS_TX_OUTZZ = "FALSE",
    parameter               PCS_ENC_DUAL = "FALSE",
    parameter               PCS_TX_BITSLIP_DATA_MODE = "X10",
    parameter               PCS_TX_BRIDGE_CLK_POLINV = "TX_BRIDGE_CLK",
    parameter    integer    PCS_COMMA_REG1 = 0,
    parameter    integer    PCS_RAPID_IMAX = 0,
    parameter    integer    PCS_RAPID_VMIN_1 = 0,
    parameter    integer    PCS_RAPID_VMIN_2 = 0,
    parameter               PCS_RX_PRBS_MODE = "DISABLE",
    parameter               PCS_RX_ERRCNT_CLR = "FALSE",
    parameter               PCS_PRBS_ERR_LPBK = "FALSE",
    parameter               PCS_TX_PRBS_MODE = "DISABLE",
    parameter               PCS_TX_INSERT_ER = "FALSE",
    parameter               PCS_ENABLE_PRBS_GEN = "FALSE",
    parameter    integer    PCS_DEFAULT_RADDR = 0,
    parameter    integer    PCS_MASTER_CHECK_OFFSET = 0,
    parameter    integer    PCS_DELAY_SET = 0,
    parameter               PCS_SEACH_OFFSET = "20BIT",
    parameter    integer    PCS_CEB_RAPIDLS_MMAX = 0,
    parameter    integer    PCS_CTC_AFULL = 20,
    parameter    integer    PCS_CTC_AEMPTY = 12,
    parameter    integer    PCS_CTC_CONTI_SKP_SET = 0,
    parameter               PCS_FAR_LOOP = "FALSE",
    parameter               PCS_NEAR_LOOP = "FALSE",
    parameter               PCS_PMA_TX2RX_PLOOP_EN = "FALSE",
    parameter               PCS_PMA_TX2RX_SLOOP_EN = "FALSE",
    parameter               PCS_PMA_RX2TX_PLOOP_EN = "FALSE",
    parameter               PCS_INT_RX_MASK_0 = "FALSE",
    parameter               PCS_INT_RX_MASK_1 = "FALSE",
    parameter               PCS_INT_RX_MASK_2 = "FALSE",
    parameter               PCS_INT_RX_MASK_3 = "FALSE",
    parameter               PCS_INT_RX_MASK_4 = "FALSE",
    parameter               PCS_INT_RX_MASK_5 = "FALSE",
    parameter               PCS_INT_RX_MASK_6 = "FALSE",
    parameter               PCS_INT_RX_MASK_7 = "FALSE",
    parameter               PCS_INT_RX_CLR_0 = "FALSE",
    parameter               PCS_INT_RX_CLR_1 = "FALSE",
    parameter               PCS_INT_RX_CLR_2 = "FALSE",
    parameter               PCS_INT_RX_CLR_3 = "FALSE",
    parameter               PCS_INT_RX_CLR_4 = "FALSE",
    parameter               PCS_INT_RX_CLR_5 = "FALSE",
    parameter               PCS_INT_RX_CLR_6 = "FALSE",
    parameter               PCS_INT_RX_CLR_7 = "FALSE",
    parameter               PCS_CA_RSTN_RX = "FALSE",
    parameter               PCS_CA_DYN_DLY_EN_RX = "FALSE",
    parameter               PCS_CA_DYN_DLY_SEL_RX = "FALSE",
    parameter    integer    PCS_CA_RX = 0,
    parameter               PCS_CA_RSTN_TX = "FALSE",
    parameter               PCS_CA_DYN_DLY_EN_TX = "FALSE",
    parameter               PCS_CA_DYN_DLY_SEL_TX = "FALSE",
    parameter    integer    PCS_CA_TX = 0,
    parameter               PCS_RXPRBS_PWR_REDUCTION = "NORMAL",
    parameter               PCS_WDALIGN_PWR_REDUCTION = "NORMAL",
    parameter               PCS_RXDEC_PWR_REDUCTION = "NORMAL",
    parameter               PCS_RXCB_PWR_REDUCTION = "NORMAL",
    parameter               PCS_RXCTC_PWR_REDUCTION = "NORMAL",
    parameter               PCS_RXGEAR_PWR_REDUCTION = "NORMAL",
    parameter               PCS_RXBRG_PWR_REDUCTION = "NORMAL",
    parameter               PCS_RXTEST_PWR_REDUCTION = "NORMAL",
    parameter               PCS_TXBRG_PWR_REDUCTION = "NORMAL",
    parameter               PCS_TXGEAR_PWR_REDUCTION = "NORMAL",
    parameter               PCS_TXENC_PWR_REDUCTION = "NORMAL",
    parameter               PCS_TXBSLP_PWR_REDUCTION = "NORMAL",
    parameter               PCS_TXPRBS_PWR_REDUCTION = "NORMAL",

    //pma_rx 
    parameter               PMA_REG_RX_PD = "ON",
    parameter               PMA_REG_RX_PD_EN = "FALSE",
    parameter               PMA_REG_RX_RESERVED_2 = "FALSE",
    parameter               PMA_REG_RX_RESERVED_3 = "FALSE",
    parameter               PMA_REG_RX_DATAPATH_PD = "ON",
    parameter               PMA_REG_RX_DATAPATH_PD_EN = "FALSE",
    parameter               PMA_REG_RX_SIGDET_PD = "ON",
    parameter               PMA_REG_RX_SIGDET_PD_EN = "FALSE",
    parameter               PMA_REG_RX_DCC_RST_N = "TRUE",
    parameter               PMA_REG_RX_DCC_RST_N_EN = "FALSE",
    parameter               PMA_REG_RX_CDR_RST_N = "TRUE",
    parameter               PMA_REG_RX_CDR_RST_N_EN = "FALSE",
    parameter               PMA_REG_RX_SIGDET_RST_N = "TRUE",
    parameter               PMA_REG_RX_SIGDET_RST_N_EN = "FALSE",
    parameter               PMA_REG_RXPCLK_SLIP = "FALSE",
    parameter               PMA_REG_RXPCLK_SLIP_OW = "FALSE",
    parameter               PMA_REG_RX_PCLKSWITCH_RST_N = "TRUE",
    parameter               PMA_REG_RX_PCLKSWITCH_RST_N_EN = "FALSE",
    parameter               PMA_REG_RX_PCLKSWITCH = "FALSE",
    parameter               PMA_REG_RX_PCLKSWITCH_EN = "FALSE",
    parameter               PMA_REG_RX_HIGHZ = "FALSE",
    parameter               PMA_REG_RX_HIGHZ_EN = "FALSE",
    parameter               PMA_REG_RX_SIGDET_CLK_WINDOW = "FALSE",
    parameter               PMA_REG_RX_SIGDET_CLK_WINDOW_OW = "FALSE",
    parameter               PMA_REG_RX_PD_BIAS_RX = "FALSE",
    parameter               PMA_REG_RX_PD_BIAS_RX_OW = "FALSE",
    parameter               PMA_REG_RX_RESET_N = "FALSE",
    parameter               PMA_REG_RX_RESET_N_OW = "FALSE",
    parameter    integer    PMA_REG_RX_RESERVED_29_28 = 0,
    parameter               PMA_REG_RX_BUSWIDTH = "20BIT",
    parameter               PMA_REG_RX_BUSWIDTH_EN = "FALSE",
    parameter               PMA_REG_RX_RATE = "DIV1",
    parameter               PMA_REG_RX_RESERVED_36 = "FALSE",
    parameter               PMA_REG_RX_RATE_EN = "FALSE",
    parameter    integer    PMA_REG_RX_RES_TRIM = 46,
    parameter               PMA_REG_RX_RESERVED_44 = "FALSE",
    parameter               PMA_REG_RX_RESERVED_45 = "FALSE",
    parameter               PMA_REG_RX_SIGDET_STATUS_EN = "FALSE",
    parameter    integer    PMA_REG_RX_RESERVED_48_47 = 0,
    parameter    integer    PMA_REG_RX_ICTRL_SIGDET = 5,
    parameter    integer    PMA_REG_CDR_READY_THD = 2734,
    parameter               PMA_REG_RX_RESERVED_65 = "FALSE",
    parameter               PMA_REG_RX_PCLK_EDGE_SEL = "POS_EDGE",
    parameter    integer    PMA_REG_RX_PIBUF_IC = 1,
    parameter               PMA_REG_RX_RESERVED_69 = "FALSE",
    parameter    integer    PMA_REG_RX_DCC_IC_RX = 1,
    parameter    integer    PMA_REG_CDR_READY_CHECK_CTRL = 0,
    parameter               PMA_REG_RX_ICTRL_TRX = "100PCT",
    parameter    integer    PMA_REG_RX_RESERVED_77_76 = 0,
    parameter    integer    PMA_REG_RX_RESERVED_79_78 = 1,
    parameter    integer    PMA_REG_RX_RESERVED_81_80 = 1,
    parameter               PMA_REG_RX_ICTRL_PIBUF = "100PCT",
    parameter               PMA_REG_RX_ICTRL_PI = "100PCT",
    parameter               PMA_REG_RX_ICTRL_DCC = "100PCT",
    parameter    integer    PMA_REG_RX_RESERVED_89_88 = 1,
    parameter               PMA_REG_TX_RATE = "DIV1",
    parameter               PMA_REG_RX_RESERVED_92 = "FALSE",
    parameter               PMA_REG_TX_RATE_EN = "FALSE",
    parameter               PMA_REG_RX_TX2RX_PLPBK_RST_N = "TRUE",
    parameter               PMA_REG_RX_TX2RX_PLPBK_RST_N_EN = "FALSE",
    parameter               PMA_REG_RX_TX2RX_PLPBK_EN = "FALSE",
    parameter               PMA_REG_TXCLK_SEL = "PLL",
    parameter               PMA_REG_RX_DATA_POLARITY = "NORMAL",
    parameter               PMA_REG_RX_ERR_INSERT = "FALSE",
    parameter               PMA_REG_UDP_CHK_EN = "FALSE",
    parameter               PMA_REG_PRBS_SEL = "PRBS7",
    parameter               PMA_REG_PRBS_CHK_EN = "FALSE",
    parameter               PMA_REG_PRBS_CHK_WIDTH_SEL = "20BIT",
    parameter               PMA_REG_BIST_CHK_PAT_SEL = "PRBS",
    parameter               PMA_REG_LOAD_ERR_CNT = "FALSE",
    parameter               PMA_REG_CHK_COUNTER_EN = "FALSE",
    parameter    integer    PMA_REG_CDR_PROP_GAIN = 7,
    parameter    integer    PMA_REG_CDR_PROP_TURBO_GAIN = 5,
    parameter    integer    PMA_REG_CDR_INT_GAIN = 7,
    parameter    integer    PMA_REG_CDR_INT_TURBO_GAIN = 5,
    parameter    integer    PMA_REG_CDR_INT_SAT_MAX = 768,
    parameter    integer    PMA_REG_CDR_INT_SAT_MIN = 255,
    parameter               PMA_REG_CDR_INT_RST = "FALSE",
    parameter               PMA_REG_CDR_INT_RST_OW = "FALSE",
    parameter               PMA_REG_CDR_PROP_RST = "FALSE",
    parameter               PMA_REG_CDR_PROP_RST_OW = "FALSE",
    parameter               PMA_REG_CDR_LOCK_RST = "FALSE",
    parameter               PMA_REG_CDR_LOCK_RST_OW = "FALSE",
    parameter    integer    PMA_REG_CDR_RX_PI_FORCE_SEL = 0,
    parameter    integer    PMA_REG_CDR_RX_PI_FORCE_D = 0,
    parameter               PMA_REG_CDR_LOCK_TIMER = "1_2U",
    parameter    integer    PMA_REG_CDR_TURBO_MODE_TIMER = 1,
    parameter               PMA_REG_CDR_LOCK_VAL = "FALSE",
    parameter               PMA_REG_CDR_LOCK_OW = "FALSE",
    parameter               PMA_REG_CDR_INT_SAT_DET_EN = "TRUE",
    parameter               PMA_REG_CDR_SAT_AUTO_DIS = "TRUE",
    parameter               PMA_REG_CDR_GAIN_AUTO = "FALSE",
    parameter               PMA_REG_CDR_TURBO_GAIN_AUTO = "FALSE",
    parameter    integer    PMA_REG_RX_RESERVED_171_167 = 0,
    parameter    integer    PMA_REG_RX_RESERVED_175_172 = 0,
    parameter               PMA_REG_CDR_SAT_DET_STATUS_EN = "FALSE",
    parameter               PMA_REG_CDR_SAT_DET_STATUS_RESET_EN = "FALSE",
    parameter               PMA_REG_CDR_PI_CTRL_RST = "FALSE",
    parameter               PMA_REG_CDR_PI_CTRL_RST_OW = "FALSE",
    parameter               PMA_REG_CDR_SAT_DET_RST = "FALSE",
    parameter               PMA_REG_CDR_SAT_DET_RST_OW = "FALSE",
    parameter               PMA_REG_CDR_SAT_DET_STICKY_RST = "FALSE",
    parameter               PMA_REG_CDR_SAT_DET_STICKY_RST_OW = "FALSE",
    parameter               PMA_REG_CDR_SIGDET_STATUS_DIS = "FALSE",
    parameter    integer    PMA_REG_CDR_SAT_DET_TIMER = 2,
    parameter               PMA_REG_CDR_SAT_DET_STATUS_VAL = "FALSE",
    parameter               PMA_REG_CDR_SAT_DET_STATUS_OW = "FALSE",
    parameter               PMA_REG_CDR_TURBO_MODE_EN = "TRUE",
    parameter               PMA_REG_RX_RESERVED_190 = "FALSE",
    parameter    integer    PMA_REG_RX_RESERVED_193_191 = 0,
    parameter               PMA_REG_CDR_STATUS_FIFO_EN = "TRUE",
    parameter    integer    PMA_REG_PMA_TEST_SEL = 0,
    parameter    integer    PMA_REG_OOB_COMWAKE_GAP_MIN = 3,
    parameter    integer    PMA_REG_OOB_COMWAKE_GAP_MAX = 11,
    parameter    integer    PMA_REG_OOB_COMINIT_GAP_MIN = 15,
    parameter    integer    PMA_REG_OOB_COMINIT_GAP_MAX = 35,
    parameter    integer    PMA_REG_RX_RESERVED_227_226 = 1,
    parameter    integer    PMA_REG_COMWAKE_STATUS_CLEAR = 0,
    parameter    integer    PMA_REG_COMINIT_STATUS_CLEAR = 0,
    parameter               PMA_REG_RX_SYNC_RST_N_EN = "FALSE",
    parameter               PMA_REG_RX_SYNC_RST_N = "TRUE",
    parameter    integer    PMA_REG_RX_RESERVED_233_232 = 0,
    parameter    integer    PMA_REG_RX_RESERVED_235_234 = 0,
    parameter               PMA_REG_RX_SATA_COMINIT_OW = "FALSE",
    parameter               PMA_REG_RX_SATA_COMINIT = "FALSE",
    parameter               PMA_REG_RX_SATA_COMWAKE_OW = "FALSE",
    parameter               PMA_REG_RX_SATA_COMWAKE = "FALSE",
    parameter    integer    PMA_REG_RX_RESERVED_241_240 = 0,
    parameter               PMA_REG_RX_DCC_DISABLE = "FALSE",
    parameter               PMA_REG_RX_RESERVED_243 = "FALSE",
    parameter               PMA_REG_RX_SLIP_SEL_EN = "FALSE",
    parameter    integer    PMA_REG_RX_SLIP_SEL = 0,
    parameter               PMA_REG_RX_SLIP_EN = "FALSE",
    parameter    integer    PMA_REG_RX_SIGDET_STATUS_SEL = 5,
    parameter               PMA_REG_RX_SIGDET_FSM_RST_N = "TRUE",
    parameter               PMA_REG_RX_RESERVED_254 = "FALSE",
    parameter               PMA_REG_RX_SIGDET_STATUS = "FALSE",
    parameter               PMA_REG_RX_SIGDET_VTH = "27MV",
    parameter    integer    PMA_REG_RX_SIGDET_GRM = 0,
    parameter               PMA_REG_RX_SIGDET_PULSE_EXT = "FALSE",
    parameter    integer    PMA_REG_RX_SIGDET_CH2_SEL = 0,
    parameter    integer    PMA_REG_RX_SIGDET_CH2_CHK_WINDOW = 3,
    parameter               PMA_REG_RX_SIGDET_CHK_WINDOW_EN = "TRUE",
    parameter    integer    PMA_REG_RX_SIGDET_NOSIG_COUNT_SETTING = 4,
    parameter               PMA_REG_SLIP_FIFO_INV_EN = "FALSE",
    parameter               PMA_REG_SLIP_FIFO_INV = "POS_EDGE",
    parameter    integer    PMA_REG_RX_SIGDET_OOB_DET_COUNT_VAL = 0,
    parameter    integer    PMA_REG_RX_SIGDET_4OOB_DET_SEL = 7,
    parameter    integer    PMA_REG_RX_RESERVED_285_283 = 0,
    parameter               PMA_REG_RX_RESERVED_286 = "FALSE",
    parameter    integer    PMA_REG_RX_SIGDET_IC_I = 10,
    parameter               PMA_REG_RX_OOB_DETECTOR_RESET_N_OW = "FALSE",
    parameter               PMA_REG_RX_OOB_DETECTOR_RESET_N = "FALSE",
    parameter               PMA_REG_RX_OOB_DETECTOR_PD_OW = "FALSE",
    parameter               PMA_REG_RX_OOB_DETECTOR_PD = "ON",
    parameter               PMA_REG_RX_LS_MODE_EN = "FALSE",
    parameter               PMA_REG_ANA_RX_EQ1_R_SET_FB_O_SEL = "FALSE",
    parameter               PMA_REG_ANA_RX_EQ2_R_SET_FB_O_SEL = "FALSE",
    parameter    integer    PMA_REG_RX_EQ1_R_SET_TOP = 0,
    parameter    integer    PMA_REG_RX_EQ1_R_SET_FB = 0,
    parameter    integer    PMA_REG_RX_EQ1_C_SET_FB = 0,
    parameter               PMA_REG_RX_EQ1_OFF = "FALSE",
    parameter    integer    PMA_REG_RX_EQ2_R_SET_TOP = 0,
    parameter    integer    PMA_REG_RX_EQ2_R_SET_FB = 0,
    parameter    integer    PMA_REG_RX_EQ2_C_SET_FB = 0,
    parameter               PMA_REG_RX_EQ2_OFF = "FALSE",
    parameter    integer    PMA_REG_EQ_DAC = 0,
    parameter    integer    PMA_REG_RX_ICTRL_EQ = 2,
    parameter               PMA_REG_EQ_DC_CALIB_EN = "FALSE",
    parameter               PMA_REG_EQ_DC_CALIB_SEL = "FALSE",
    parameter    integer    PMA_REG_RX_RESERVED_337_330 = 0,
    parameter    integer    PMA_REG_RX_RESERVED_345_338 = 0,
    parameter    integer    PMA_REG_RX_RESERVED_353_346 = 0,
    parameter    integer    PMA_REG_RX_RESERVED_361_354 = 0,
    parameter    integer    PMA_CTLE_CTRL_REG_I = 0,
    parameter               PMA_CTLE_REG_FORCE_SEL_I = "FALSE",
    parameter               PMA_CTLE_REG_HOLD_I = "FALSE",
    parameter    integer    PMA_CTLE_REG_INIT_DAC_I = 0,
    parameter               PMA_CTLE_REG_POLARITY_I = "FALSE",
    parameter    integer    PMA_CTLE_REG_SHIFTER_GAIN_I = 0,        
    parameter    integer    PMA_CTLE_REG_THRESHOLD_I = 0,
    parameter               PMA_REG_RX_RES_TRIM_EN = "FALSE",
    parameter    integer    PMA_REG_RX_RESERVED_393_389 = 0,
    parameter               PMA_CFG_RX_LANE_POWERUP = "OFF",
    parameter               PMA_CFG_RX_PMA_RSTN = "FALSE",
    parameter               PMA_INT_PMA_RX_MASK_0 = "FALSE",
    parameter               PMA_INT_PMA_RX_CLR_0 = "FALSE",
    parameter               PMA_CFG_CTLE_ADP_RSTN = "TRUE",
 
    //pma_tx
    parameter               PMA_REG_TX_PD = "ON",  
    parameter               PMA_REG_TX_PD_OW = "TRUE",
    parameter               PMA_REG_TX_MAIN_PRE_Z = "FALSE",
    parameter               PMA_REG_TX_MAIN_PRE_Z_OW = "FALSE",
    parameter    integer    PMA_REG_TX_BEACON_TIMER_SEL = 0,
    parameter               PMA_REG_TX_RXDET_REQ_OW = "FALSE",
    parameter               PMA_REG_TX_RXDET_REQ = "FALSE",
    parameter               PMA_REG_TX_BEACON_EN_OW = "FALSE",
    parameter               PMA_REG_TX_BEACON_EN = "FALSE",
    parameter               PMA_REG_TX_EI_EN_OW = "FALSE",
    parameter               PMA_REG_TX_EI_EN = "FALSE",
    parameter               PMA_REG_TX_BIT_CONV = "FALSE",
    parameter    integer    PMA_REG_TX_RES_CAL = 50,
    parameter               PMA_REG_TX_RESERVED_19 = "FALSE",
    parameter    integer    PMA_REG_TX_RESERVED_25_20 = 32,
    parameter    integer    PMA_REG_TX_RESERVED_33_26 = 0,
    parameter    integer    PMA_REG_TX_RESERVED_41_34 = 0,
    parameter    integer    PMA_REG_TX_RESERVED_49_42 = 0,
    parameter    integer    PMA_REG_TX_RESERVED_57_50 = 0,
    parameter               PMA_REG_TX_SYNC_OW = "FALSE",
    parameter               PMA_REG_TX_SYNC = "FALSE",
    parameter               PMA_REG_TX_PD_POST = "OFF",
    parameter               PMA_REG_TX_PD_POST_OW = "TRUE",
    parameter               PMA_REG_TX_RESET_N_OW = "FALSE",
    parameter               PMA_REG_TX_RESET_N = "TRUE",
    parameter               PMA_REG_TX_RESERVED_64 = "FALSE",
    parameter               PMA_REG_TX_RESERVED_65 = "TRUE",
    parameter               PMA_REG_TX_BUSWIDTH_OW = "FALSE",
    parameter               PMA_REG_TX_BUSWIDTH = "20BIT",
    parameter               PMA_REG_PLL_READY_OW = "FALSE",
    parameter               PMA_REG_PLL_READY = "TRUE",
    parameter               PMA_REG_TX_RESERVED_72 = "FALSE",
    parameter               PMA_REG_TX_RESERVED_73 = "FALSE",
    parameter               PMA_REG_TX_RESERVED_74 = "FALSE",
    parameter    integer    PMA_REG_EI_PCLK_DELAY_SEL = 0,
    parameter               PMA_REG_TX_RESERVED_77 = "FALSE",
    parameter    integer    PMA_REG_TX_RESERVED_83_78 = 0,
    parameter    integer    PMA_REG_TX_RESERVED_89_84 = 0,
    parameter    integer    PMA_REG_TX_RESERVED_95_90 = 0,
    parameter    integer    PMA_REG_TX_RESERVED_101_96 = 0,
    parameter    integer    PMA_REG_TX_RESERVED_107_102 = 0,
    parameter    integer    PMA_REG_TX_RESERVED_113_108 = 0,
    parameter    integer    PMA_REG_TX_AMP_DAC0 = 25,
    parameter    integer    PMA_REG_TX_AMP_DAC1 = 19,
    parameter    integer    PMA_REG_TX_AMP_DAC2 = 14,
    parameter    integer    PMA_REG_TX_AMP_DAC3 = 9,
    parameter    integer    PMA_REG_TX_RESERVED_143_138 = 5,
    parameter    integer    PMA_REG_TX_MARGIN = 0,
    parameter               PMA_REG_TX_MARGIN_OW = "FALSE",
    parameter    integer    PMA_REG_TX_RESERVED_149_148 = 0,
    parameter               PMA_REG_TX_RESERVED_150 = "FALSE",
    parameter               PMA_REG_TX_SWING = "FALSE",
    parameter               PMA_REG_TX_SWING_OW = "FALSE",
    parameter               PMA_REG_TX_RESERVED_153 = "FALSE",
    parameter               PMA_REG_TX_RXDET_THRESHOLD = "84MV",
    parameter    integer    PMA_REG_TX_RESERVED_157_156 = 0,
    parameter               PMA_REG_TX_BEACON_OSC_CTRL = "FALSE",
    parameter    integer    PMA_REG_TX_RESERVED_160_159 = 0,
    parameter    integer    PMA_REG_TX_RESERVED_162_161 = 0,
    parameter               PMA_REG_TX_TX2RX_SLPBACK_EN = "FALSE",
    parameter               PMA_REG_TX_PCLK_EDGE_SEL = "FALSE",
    parameter               PMA_REG_TX_RXDET_STATUS_OW = "FALSE",
    parameter               PMA_REG_TX_RXDET_STATUS = "TRUE",
    parameter               PMA_REG_TX_PRBS_GEN_EN = "FALSE",
    parameter               PMA_REG_TX_PRBS_GEN_WIDTH_SEL = "20BIT",
    parameter               PMA_REG_TX_PRBS_SEL = "PRBS7",
    parameter    integer    PMA_REG_TX_UDP_DATA_7_TO_0 = 5,
    parameter    integer    PMA_REG_TX_UDP_DATA_15_TO_8 = 235,
    parameter    integer    PMA_REG_TX_UDP_DATA_19_TO_16 = 3,
    parameter               PMA_REG_TX_RESERVED_192 = "FALSE",
    parameter    integer    PMA_REG_TX_FIFO_WP_CTRL = 4,
    parameter               PMA_REG_TX_FIFO_EN = "FALSE",
    parameter    integer    PMA_REG_TX_DATA_MUX_SEL = 0,
    parameter               PMA_REG_TX_ERR_INSERT = "FALSE",
    parameter    integer    PMA_REG_TX_RESERVED_203_200 = 0,
    parameter               PMA_REG_TX_RESERVED_204 = "FALSE",
    parameter               PMA_REG_TX_SATA_EN = "FALSE",
    parameter    integer    PMA_REG_TX_RESERVED_207_206 = 0,
    parameter               PMA_REG_RATE_CHANGE_TXPCLK_ON_OW = "FALSE",
    parameter               PMA_REG_RATE_CHANGE_TXPCLK_ON = "TRUE",
    parameter    integer    PMA_REG_TX_CFG_POST1 = 0,
    parameter    integer    PMA_REG_TX_CFG_POST2 = 0,
    parameter    integer    PMA_REG_TX_DEEMP = 0,
    parameter               PMA_REG_TX_DEEMP_OW = "FALSE",
    parameter    integer    PMA_REG_TX_RESERVED_224_223 = 0,
    parameter               PMA_REG_TX_RESERVED_225 = "FALSE",
    parameter    integer    PMA_REG_TX_RESERVED_229_226 = 0,
    parameter    integer    PMA_REG_TX_OOB_DELAY_SEL = 0,
    parameter               PMA_REG_TX_POLARITY = "NORMAL",
    parameter               PMA_REG_ANA_TX_JTAG_DATA_O_SEL = "FALSE",
    parameter               PMA_REG_TX_RESERVED_236 = "FALSE",
    parameter               PMA_REG_TX_LS_MODE_EN = "FALSE",
    parameter               PMA_REG_TX_JTAG_MODE_EN_OW = "FALSE",
    parameter               PMA_REG_TX_JTAG_MODE_EN = "FALSE",
    parameter               PMA_REG_RX_JTAG_MODE_EN_OW = "FALSE",
    parameter               PMA_REG_RX_JTAG_MODE_EN = "FALSE",
    parameter               PMA_REG_RX_JTAG_OE = "TRUE",
    parameter    integer    PMA_REG_RX_ACJTAG_VHYSTSEL = 0,
    parameter               PMA_REG_TX_RES_CAL_EN = "FALSE",
    parameter    integer    PMA_REG_RX_TERM_MODE_CTRL = 4,
    parameter    integer    PMA_REG_TX_RESERVED_251_250 = 0,
    parameter               PMA_REG_PLPBK_TXPCLK_EN = "FALSE",
    parameter               PMA_REG_TX_RESERVED_253 = "FALSE",
    parameter               PMA_REG_TX_RESERVED_254 = "FALSE",
    parameter               PMA_REG_TX_RESERVED_255 = "FALSE",
    parameter               PMA_REG_TX_RESERVED_256 = "FALSE",
    parameter               PMA_REG_TX_RESERVED_257 = "FALSE",
    parameter    integer    PMA_REG_TX_PH_SEL = 1,
    parameter    integer    PMA_REG_TX_CFG_PRE = 0, 
    parameter    integer    PMA_REG_TX_CFG_MAIN = 0,
    parameter    integer    PMA_REG_CFG_POST = 0,
    parameter               PMA_REG_PD_MAIN = "TRUE",
    parameter               PMA_REG_PD_PRE = "TRUE",
    parameter               PMA_REG_TX_LS_DATA = "FALSE",
    parameter    integer    PMA_REG_TX_DCC_BUF_SZ_SEL = 0,
    parameter    integer    PMA_REG_TX_DCC_CAL_CUR_TUNE = 0,
    parameter               PMA_REG_TX_DCC_CAL_EN = "FALSE",
    parameter    integer    PMA_REG_TX_DCC_CUR_SS = 0,
    parameter               PMA_REG_TX_DCC_FA_CTRL = "FALSE",
    parameter               PMA_REG_TX_DCC_RI_CTRL = "FALSE",
    parameter    integer    PMA_REG_ATB_SEL_2_TO_0 = 0,
    parameter    integer    PMA_REG_ATB_SEL_9_TO_3 = 0,
    parameter    integer    PMA_REG_TX_CFG_7_TO_0 = 0,
    parameter    integer    PMA_REG_TX_CFG_15_TO_8 = 0,
    parameter    integer    PMA_REG_TX_CFG_23_TO_16 = 0,
    parameter    integer    PMA_REG_TX_CFG_31_TO_24 = 0,
    parameter               PMA_REG_TX_OOB_EI_EN = "FALSE",
    parameter               PMA_REG_TX_OOB_EI_EN_OW = "FALSE",
    parameter               PMA_REG_TX_BEACON_EN_DELAYED = "FALSE",
    parameter               PMA_REG_TX_BEACON_EN_DELAYED_OW = "FALSE",
    parameter               PMA_REG_TX_JTAG_DATA = "FALSE",
    parameter    integer    PMA_REG_TX_RXDET_TIMER_SEL = 87,
    parameter    integer    PMA_REG_TX_CFG1_7_0 = 0,
    parameter    integer    PMA_REG_TX_CFG1_15_8 = 0,
    parameter    integer    PMA_REG_TX_CFG1_23_16 = 0,
    parameter    integer    PMA_REG_TX_CFG1_31_24 = 0,
    parameter               PMA_REG_CFG_LANE_POWERUP = "OFF",
    //parameter               PMA_REG_CFG_PMA_POR_N = "TRUE",
    parameter               PMA_REG_CFG_TX_LANE_POWERUP_CLKPATH = "FALSE",
    parameter               PMA_REG_CFG_TX_LANE_POWERUP_PISO = "FALSE",
    parameter               PMA_REG_CFG_TX_LANE_POWERUP_DRIVER = "FALSE"
    //parameter               PMA_REG_CFG_TX_PMA_RSTN = "TRUE"
    
)(

//////////Output/////////////////////////////////////////////////////////
    //PAD
    output              P_TX_SDN,  
    output              P_TX_SDP,

    //SRB related
    output              P_PCS_RX_MCB_STATUS, 
    output              P_PCS_LSM_SYNCED, 
    output              P_CFG_READY,
    output [7:0]        P_CFG_RDATA, 
    output              P_CFG_INT, 
    output [46:0]       P_RDATA, 
    output              P_RCLK2FABRIC, 
    output              P_TCLK2FABRIC, 

    output              P_RX_SIGDET_STATUS, 
    output              P_RX_SATA_COMINIT, 
    output              P_RX_SATA_COMWAKE, 
    output              P_RX_LS_DATA, 
    output              P_RX_READY, 
    output [19:0]       P_TEST_STATUS, 
    output              P_TX_RXDET_STATUS, 
    output              P_CA_ALIGN_RX, 
    output              P_CA_ALIGN_TX, 

    //New Added
    output              PMA_RCLK,

    //cin and cout
    output [18:0]       LANE_COUT_BUS_FORWARD,

    //output              RFIFO_EN_CB_COUT, 
    //output              RFIFO_EN_AFTER_CTC_COUT, 
    //output              RFIFO_EN_AFTER_CTC_GB_COUT, 
    //output              RFIFO_EN_BRIDGE_COUT, 
    //output              TFIFO_EN_PCS_TX_COUT, 
    //output              TFIFO_EN_BRIDGE_COUT, 
    //output              PCS_TCLK_EN_COUT, 
    //output              GEAR_TCLK_EN_COUT, 
    //output              APATTERN_MATCH_LSB_COUT, 
    //output              APATTERN_MATCH_MSB_COUT, 
    //output              APATTERN_SEACHING_PROC_COUT, 
    //output              CB_RCLK_EN_COUT, 
    //output              AFTER_CTC_RCLK_EN_COUT, 
    //output              AFTER_CTC_RCLK_EN_GB_COUT, 
    //output              SKIP_ADD_MCB_COUT, 
    //output              SKIP_DEL_MCB_COUT, 
    //output              SKIP_DEL_LSB_MCB_COUT, 
    //output              SKIP_ADD_LSB_MCB_COUT, 
    //output              CTC_RD_FIFO_COUT, 

    output              APATTERN_STATUS_COUT, //Backword

    //out
    output              TXPCLK_PLL,

//////////Input/////////////////////////////////////////////////////////
    //PAD
    input               P_RX_SDN,
    input               P_RX_SDP,

    //SRB related
    input               P_RX_CLK_FR_CORE,
    input               P_RCLK2_FR_CORE,
    input               P_TX_CLK_FR_CORE,
    input               P_TCLK2_FR_CORE,
    input               P_PCS_TX_RST,
    input               P_PCS_RX_RST,
    input               P_PCS_CB_RST,
    input               P_RXGEAR_SLIP,
    input               P_CFG_CLK,
    input               P_CFG_RST,
    input               P_CFG_PSEL,
    input               P_CFG_ENABLE,
    input               P_CFG_WRITE,
    input [11:0]        P_CFG_ADDR,
    input [7:0]         P_CFG_WDATA,
    input [45:0]        P_TDATA,
    input               P_PCS_WORD_ALIGN_EN,
    input               P_RX_POLARITY_INVERT,
    input               P_CEB_ADETECT_EN,
    input               P_PCS_MCB_EXT_EN,
    input               P_PCS_NEAREND_LOOP,
    input               P_PCS_FAREND_LOOP,
    input               P_PMA_NEAREND_PLOOP,
    input               P_PMA_NEAREND_SLOOP,
    input               P_PMA_FAREND_PLOOP,

    input               P_LANE_PD,
    input               P_LANE_RST,
    input               P_RX_LANE_PD,
    input               P_RX_PMA_RST,
    input               P_CTLE_ADP_RST,
    input [1:0]         P_TX_DEEMP,
    input               P_TX_LS_DATA,
    input               P_TX_BEACON_EN,
    input               P_TX_SWING,
    input               P_TX_RXDET_REQ,
    input [2:0]         P_TX_RATE,
    input [2:0]         P_TX_BUSWIDTH,
    input [2:0]         P_TX_MARGIN,
    input               P_TX_PMA_RST,
    input               P_TX_LANE_PD_CLKPATH,
    input               P_TX_LANE_PD_PISO,
    input               P_TX_LANE_PD_DRIVER,
    input [2:0]         P_RX_RATE,
    input [2:0]         P_RX_BUSWIDTH,
    input               P_RX_HIGHZ,
    input [7:0]         P_CIM_CLK_ALIGNER_RX,
    input [7:0]         P_CIM_CLK_ALIGNER_TX,
    input               P_CIM_DYN_DLY_SEL_RX,
    input               P_CIM_DYN_DLY_SEL_TX,
    input               P_CIM_START_ALIGN_RX,
    input               P_CIM_START_ALIGN_TX,

    //New Added
    input               MCB_RCLK,
    input               SYNC,
    input               RATE_CHANGE,
    input               PLL_LOCK_SEL,

    //cin and cout 
    input [18:0]        LANE_CIN_BUS_FORWARD,

    //input               RFIFO_EN_CB_CIN,
    //input               RFIFO_EN_AFTER_CTC_CIN,
    //input               RFIFO_EN_AFTER_CTC_GB_CIN,
    //input               RFIFO_EN_BRIDGE_CIN,
    //input               TFIFO_EN_PCS_TX_CIN,
    //input               TFIFO_EN_BRIDGE_CIN,
    //input               PCS_TCLK_EN_CIN,
    //input               GEAR_TCLK_EN_CIN,
    //input               APATTERN_MATCH_LSB_CIN,
    //input               APATTERN_MATCH_MSB_CIN,
    //input               APATTERN_SEACHING_PROC_CIN,
    //input               CB_RCLK_EN_CIN,
    //input               AFTER_CTC_RCLK_EN_CIN,
    //input               AFTER_CTC_RCLK_EN_GB_CIN,
    //input               SKIP_ADD_MCB_CIN,
    //input               SKIP_DEL_MCB_CIN,
    //input               SKIP_DEL_LSB_MCB_CIN,
    //input               SKIP_ADD_LSB_MCB_CIN,
    //input               CTC_RD_FIFO_CIN,

    input               APATTERN_STATUS_CIN,//Backward

    //From PLL
    input               CLK_TXP,
    input               CLK_TXN,
    input               CLK_RX0,
    input               CLK_RX90,
    input               CLK_RX180,
    input               CLK_RX270,

    input               PLL_PD_I,
    input               PLL_RESET_I,
    input               PLL_REFCLK_I,
    input [5:0]         PLL_RES_TRIM_I

);

HSSTLP_LANE
#(

    .CP_MUX_BIAS                                    (MUX_BIAS),
    .CP_PD_CLK                                      (PD_CLK),
    .CP_REG_SYNC                                    (REG_SYNC),
    .CP_REG_SYNC_OW                                 (REG_SYNC_OW),
    .CP_PLL_LOCK_OW                                 (PLL_LOCK_OW),
    .CP_PLL_LOCK_OW_EN                              (PLL_LOCK_OW_EN),

    //pcs
    .CP_PCS_SLAVE                                   (PCS_SLAVE),

    .CP_PCS_BYPASS_WORD_ALIGN                       (PCS_BYPASS_WORD_ALIGN),          
    .CP_PCS_BYPASS_DENC                             (PCS_BYPASS_DENC),           
    .CP_PCS_BYPASS_BONDING                          (PCS_BYPASS_BONDING), 
    .CP_PCS_BYPASS_CTC                              (PCS_BYPASS_CTC), 
    .CP_PCS_BYPASS_GEAR                             (PCS_BYPASS_GEAR), 
    .CP_PCS_BYPASS_BRIDGE                           (PCS_BYPASS_BRIDGE), 
    .CP_PCS_BYPASS_BRIDGE_FIFO                      (PCS_BYPASS_BRIDGE_FIFO), 
    .CP_PCS_DATA_MODE                               (PCS_DATA_MODE), 
    .CP_PCS_RX_POLARITY_INV                         (PCS_RX_POLARITY_INV), 
    .CP_PCS_ALIGN_MODE                              (PCS_ALIGN_MODE), 
    .CP_PCS_SAMP_16B                                (PCS_SAMP_16B),          
    .CP_PCS_FARLP_PWR_REDUCTION                     (PCS_FARLP_PWR_REDUCTION),           
    .CP_PCS_COMMA_REG0                              (PCS_COMMA_REG0), 
    .CP_PCS_COMMA_MASK                              (PCS_COMMA_MASK), 
    .CP_PCS_CEB_MODE                                (PCS_CEB_MODE), 
    .CP_PCS_CTC_MODE                                (PCS_CTC_MODE), 
    .CP_PCS_A_REG                                   (PCS_A_REG), 
    .CP_PCS_GE_AUTO_EN                              (PCS_GE_AUTO_EN), 
    .CP_PCS_SKIP_REG0                               (PCS_SKIP_REG0), 
    .CP_PCS_SKIP_REG1                               (PCS_SKIP_REG1), 
    .CP_PCS_SKIP_REG2                               (PCS_SKIP_REG2),          
    .CP_PCS_SKIP_REG3                               (PCS_SKIP_REG3),           
    .CP_PCS_DEC_DUAL                                (PCS_DEC_DUAL), 
    .CP_PCS_SPLIT                                   (PCS_SPLIT), 
    .CP_PCS_FIFOFLAG_CTC                            (PCS_FIFOFLAG_CTC), 
    .CP_PCS_COMMA_DET_MODE                          (PCS_COMMA_DET_MODE), 
    .CP_PCS_ERRDETECT_SILENCE                       (PCS_ERRDETECT_SILENCE), 
    .CP_PCS_PMA_RCLK_POLINV                         (PCS_PMA_RCLK_POLINV), 
    .CP_PCS_PCS_RCLK_SEL                            (PCS_PCS_RCLK_SEL), 
    .CP_PCS_CB_RCLK_SEL                             (PCS_CB_RCLK_SEL),  
    .CP_PCS_AFTER_CTC_RCLK_SEL                      (PCS_AFTER_CTC_RCLK_SEL),           
    .CP_PCS_RCLK_POLINV                             (PCS_RCLK_POLINV), 
    .CP_PCS_BRIDGE_RCLK_SEL                         (PCS_BRIDGE_RCLK_SEL), 
    .CP_PCS_PCS_RCLK_EN                             (PCS_PCS_RCLK_EN),
    .CP_PCS_CB_RCLK_EN                              (PCS_CB_RCLK_EN),
    .CP_PCS_AFTER_CTC_RCLK_EN                       (PCS_AFTER_CTC_RCLK_EN),
    .CP_PCS_AFTER_CTC_RCLK_EN_GB                    (PCS_AFTER_CTC_RCLK_EN_GB),
    .CP_PCS_PCS_RX_RSTN                             (PCS_PCS_RX_RSTN),
    .CP_PCS_PCIE_SLAVE                              (PCS_PCIE_SLAVE),
    .CP_PCS_RX_64B66B_67B                           (PCS_RX_64B66B_67B),
    .CP_PCS_RX_BRIDGE_CLK_POLINV                    (PCS_RX_BRIDGE_CLK_POLINV),
    .CP_PCS_PCS_CB_RSTN                             (PCS_PCS_CB_RSTN),
    .CP_PCS_TX_BRIDGE_GEAR_SEL                      (PCS_TX_BRIDGE_GEAR_SEL),
    .CP_PCS_TX_BYPASS_BRIDGE_UINT                   (PCS_TX_BYPASS_BRIDGE_UINT),
    .CP_PCS_TX_BYPASS_BRIDGE_FIFO                   (PCS_TX_BYPASS_BRIDGE_FIFO),
    .CP_PCS_TX_BYPASS_GEAR                          (PCS_TX_BYPASS_GEAR),
    .CP_PCS_TX_BYPASS_ENC                           (PCS_TX_BYPASS_ENC),
    .CP_PCS_TX_BYPASS_BIT_SLIP                      (PCS_TX_BYPASS_BIT_SLIP),
    .CP_PCS_TX_GEAR_SPLIT                           (PCS_TX_GEAR_SPLIT),
    .CP_PCS_TX_DRIVE_REG_MODE                       (PCS_TX_DRIVE_REG_MODE),
    .CP_PCS_TX_BIT_SLIP_CYCLES                      (PCS_TX_BIT_SLIP_CYCLES),
    .CP_PCS_INT_TX_MASK_0                           (PCS_INT_TX_MASK_0),
    .CP_PCS_INT_TX_MASK_1                           (PCS_INT_TX_MASK_1),
    .CP_PCS_INT_TX_MASK_2                           (PCS_INT_TX_MASK_2),
    .CP_PCS_INT_TX_CLR_0                            (PCS_INT_TX_CLR_0),
    .CP_PCS_INT_TX_CLR_1                            (PCS_INT_TX_CLR_1),
    .CP_PCS_INT_TX_CLR_2                            (PCS_INT_TX_CLR_2),
    .CP_PCS_TX_PMA_TCLK_POLINV                      (PCS_TX_PMA_TCLK_POLINV),
    .CP_PCS_TX_PCS_CLK_EN_SEL                       (PCS_TX_PCS_CLK_EN_SEL),
    .CP_PCS_TX_BRIDGE_TCLK_SEL                      (PCS_TX_BRIDGE_TCLK_SEL),
    .CP_PCS_TX_TCLK_POLINV                          (PCS_TX_TCLK_POLINV),
    .CP_PCS_PCS_TCLK_SEL                            (PCS_PCS_TCLK_SEL),
    .CP_PCS_TX_PCS_TX_RSTN                          (PCS_TX_PCS_TX_RSTN),
    .CP_PCS_TX_SLAVE                                (PCS_TX_SLAVE),
    .CP_PCS_TX_GEAR_CLK_EN_SEL                      (PCS_TX_GEAR_CLK_EN_SEL),
    .CP_PCS_DATA_WIDTH_MODE                         (PCS_DATA_WIDTH_MODE),
    .CP_PCS_TX_64B66B_67B                           (PCS_TX_64B66B_67B),
    .CP_PCS_GEAR_TCLK_SEL                           (PCS_GEAR_TCLK_SEL),
    .CP_PCS_TX_TCLK2FABRIC_SEL                      (PCS_TX_TCLK2FABRIC_SEL),
    .CP_PCS_TX_OUTZZ                                (PCS_TX_OUTZZ),
    .CP_PCS_ENC_DUAL                                (PCS_ENC_DUAL),
    .CP_PCS_TX_BITSLIP_DATA_MODE                    (PCS_TX_BITSLIP_DATA_MODE),
    .CP_PCS_TX_BRIDGE_CLK_POLINV                    (PCS_TX_BRIDGE_CLK_POLINV),
    .CP_PCS_COMMA_REG1                              (PCS_COMMA_REG1),
    .CP_PCS_RAPID_IMAX                              (PCS_RAPID_IMAX),
    .CP_PCS_RAPID_VMIN_1                            (PCS_RAPID_VMIN_1),
    .CP_PCS_RAPID_VMIN_2                            (PCS_RAPID_VMIN_2),
    .CP_PCS_RX_PRBS_MODE                            (PCS_RX_PRBS_MODE),
    .CP_PCS_RX_ERRCNT_CLR                           (PCS_RX_ERRCNT_CLR),
    .CP_PCS_PRBS_ERR_LPBK                           (PCS_PRBS_ERR_LPBK),
    .CP_PCS_TX_PRBS_MODE                            (PCS_TX_PRBS_MODE),
    .CP_PCS_TX_INSERT_ER                            (PCS_TX_INSERT_ER),
    .CP_PCS_ENABLE_PRBS_GEN                         (PCS_ENABLE_PRBS_GEN),
    .CP_PCS_DEFAULT_RADDR                           (PCS_DEFAULT_RADDR),
    .CP_PCS_MASTER_CHECK_OFFSET                     (PCS_MASTER_CHECK_OFFSET),
    .CP_PCS_DELAY_SET                               (PCS_DELAY_SET),
    .CP_PCS_SEACH_OFFSET                            (PCS_SEACH_OFFSET),
    .CP_PCS_CEB_RAPIDLS_MMAX                        (PCS_CEB_RAPIDLS_MMAX),
    .CP_PCS_CTC_AFULL                               (PCS_CTC_AFULL),
    .CP_PCS_CTC_AEMPTY                              (PCS_CTC_AEMPTY),
    .CP_PCS_CTC_CONTI_SKP_SET                       (PCS_CTC_CONTI_SKP_SET),
    .CP_PCS_FAR_LOOP                                (PCS_FAR_LOOP),
    .CP_PCS_NEAR_LOOP                               (PCS_NEAR_LOOP),
    .CP_PCS_PMA_TX2RX_PLOOP_EN                      (PCS_PMA_TX2RX_PLOOP_EN),
    .CP_PCS_PMA_TX2RX_SLOOP_EN                      (PCS_PMA_TX2RX_SLOOP_EN),
    .CP_PCS_PMA_RX2TX_PLOOP_EN                      (PCS_PMA_RX2TX_PLOOP_EN),
    .CP_PCS_INT_RX_MASK_0                           (PCS_INT_RX_MASK_0),
    .CP_PCS_INT_RX_MASK_1                           (PCS_INT_RX_MASK_1),
    .CP_PCS_INT_RX_MASK_2                           (PCS_INT_RX_MASK_2),
    .CP_PCS_INT_RX_MASK_3                           (PCS_INT_RX_MASK_3),
    .CP_PCS_INT_RX_MASK_4                           (PCS_INT_RX_MASK_4),
    .CP_PCS_INT_RX_MASK_5                           (PCS_INT_RX_MASK_5),
    .CP_PCS_INT_RX_MASK_6                           (PCS_INT_RX_MASK_6),
    .CP_PCS_INT_RX_MASK_7                           (PCS_INT_RX_MASK_7),
    .CP_PCS_INT_RX_CLR_0                            (PCS_INT_RX_CLR_0),
    .CP_PCS_INT_RX_CLR_1                            (PCS_INT_RX_CLR_1),
    .CP_PCS_INT_RX_CLR_2                            (PCS_INT_RX_CLR_2),
    .CP_PCS_INT_RX_CLR_3                            (PCS_INT_RX_CLR_3),
    .CP_PCS_INT_RX_CLR_4                            (PCS_INT_RX_CLR_4),
    .CP_PCS_INT_RX_CLR_5                            (PCS_INT_RX_CLR_5),
    .CP_PCS_INT_RX_CLR_6                            (PCS_INT_RX_CLR_6),
    .CP_PCS_INT_RX_CLR_7                            (PCS_INT_RX_CLR_7),
    .CP_PCS_CA_RSTN_RX                              (PCS_CA_RSTN_RX),
    .CP_PCS_CA_DYN_DLY_EN_RX                        (PCS_CA_DYN_DLY_EN_RX),
    .CP_PCS_CA_DYN_DLY_SEL_RX                       (PCS_CA_DYN_DLY_SEL_RX),
    .CP_PCS_CA_RX                                   (PCS_CA_RX),
    .CP_PCS_CA_RSTN_TX                              (PCS_CA_RSTN_TX),
    .CP_PCS_CA_DYN_DLY_EN_TX                        (PCS_CA_DYN_DLY_EN_TX),
    .CP_PCS_CA_DYN_DLY_SEL_TX                       (PCS_CA_DYN_DLY_SEL_TX),
    .CP_PCS_CA_TX                                   (PCS_CA_TX),
    .CP_PCS_RXPRBS_PWR_REDUCTION                    (PCS_RXPRBS_PWR_REDUCTION),
    .CP_PCS_WDALIGN_PWR_REDUCTION                   (PCS_WDALIGN_PWR_REDUCTION),
    .CP_PCS_RXDEC_PWR_REDUCTION                     (PCS_RXDEC_PWR_REDUCTION),
    .CP_PCS_RXCB_PWR_REDUCTION                      (PCS_RXCB_PWR_REDUCTION),
    .CP_PCS_RXCTC_PWR_REDUCTION                     (PCS_RXCTC_PWR_REDUCTION),
    .CP_PCS_RXGEAR_PWR_REDUCTION                    (PCS_RXGEAR_PWR_REDUCTION),
    .CP_PCS_RXBRG_PWR_REDUCTION                     (PCS_RXBRG_PWR_REDUCTION),
    .CP_PCS_RXTEST_PWR_REDUCTION                    (PCS_RXTEST_PWR_REDUCTION),
    .CP_PCS_TXBRG_PWR_REDUCTION                     (PCS_TXBRG_PWR_REDUCTION),
    .CP_PCS_TXGEAR_PWR_REDUCTION                    (PCS_TXGEAR_PWR_REDUCTION),
    .CP_PCS_TXENC_PWR_REDUCTION                     (PCS_TXENC_PWR_REDUCTION),
    .CP_PCS_TXBSLP_PWR_REDUCTION                    (PCS_TXBSLP_PWR_REDUCTION),
    .CP_PCS_TXPRBS_PWR_REDUCTION                    (PCS_TXPRBS_PWR_REDUCTION),

    //pma_rx 
    .CP_PMA_REG_RX_PD                               (PMA_REG_RX_PD),
    .CP_PMA_REG_RX_PD_EN                            (PMA_REG_RX_PD_EN),
    .CP_PMA_REG_RX_RESERVED_2                       (PMA_REG_RX_RESERVED_2),
    .CP_PMA_REG_RX_RESERVED_3                       (PMA_REG_RX_RESERVED_3),
    .CP_PMA_REG_RX_DATAPATH_PD                      (PMA_REG_RX_DATAPATH_PD),
    .CP_PMA_REG_RX_DATAPATH_PD_EN                   (PMA_REG_RX_DATAPATH_PD_EN),
    .CP_PMA_REG_RX_SIGDET_PD                        (PMA_REG_RX_SIGDET_PD),
    .CP_PMA_REG_RX_SIGDET_PD_EN                     (PMA_REG_RX_SIGDET_PD_EN),
    .CP_PMA_REG_RX_DCC_RST_N                        (PMA_REG_RX_DCC_RST_N),
    .CP_PMA_REG_RX_DCC_RST_N_EN                     (PMA_REG_RX_DCC_RST_N_EN),
    .CP_PMA_REG_RX_CDR_RST_N                        (PMA_REG_RX_CDR_RST_N),
    .CP_PMA_REG_RX_CDR_RST_N_EN                     (PMA_REG_RX_CDR_RST_N_EN),
    .CP_PMA_REG_RX_SIGDET_RST_N                     (PMA_REG_RX_SIGDET_RST_N),
    .CP_PMA_REG_RX_SIGDET_RST_N_EN                  (PMA_REG_RX_SIGDET_RST_N_EN),
    .CP_PMA_REG_RXPCLK_SLIP                         (PMA_REG_RXPCLK_SLIP),
    .CP_PMA_REG_RXPCLK_SLIP_OW                      (PMA_REG_RXPCLK_SLIP_OW),
    .CP_PMA_REG_RX_PCLKSWITCH_RST_N                 (PMA_REG_RX_PCLKSWITCH_RST_N),
    .CP_PMA_REG_RX_PCLKSWITCH_RST_N_EN              (PMA_REG_RX_PCLKSWITCH_RST_N_EN),
    .CP_PMA_REG_RX_PCLKSWITCH                       (PMA_REG_RX_PCLKSWITCH),
    .CP_PMA_REG_RX_PCLKSWITCH_EN                    (PMA_REG_RX_PCLKSWITCH_EN),
    .CP_PMA_REG_RX_HIGHZ                            (PMA_REG_RX_HIGHZ),
    .CP_PMA_REG_RX_HIGHZ_EN                         (PMA_REG_RX_HIGHZ_EN),
    .CP_PMA_REG_RX_SIGDET_CLK_WINDOW                (PMA_REG_RX_SIGDET_CLK_WINDOW),
    .CP_PMA_REG_RX_SIGDET_CLK_WINDOW_OW             (PMA_REG_RX_SIGDET_CLK_WINDOW_OW),
    .CP_PMA_REG_RX_PD_BIAS_RX                       (PMA_REG_RX_PD_BIAS_RX),
    .CP_PMA_REG_RX_PD_BIAS_RX_OW                    (PMA_REG_RX_PD_BIAS_RX_OW),
    .CP_PMA_REG_RX_RESET_N                          (PMA_REG_RX_RESET_N),
    .CP_PMA_REG_RX_RESET_N_OW                       (PMA_REG_RX_RESET_N_OW),
    .CP_PMA_REG_RX_RESERVED_29_28                   (PMA_REG_RX_RESERVED_29_28),
    .CP_PMA_REG_RX_BUSWIDTH                         (PMA_REG_RX_BUSWIDTH),
    .CP_PMA_REG_RX_BUSWIDTH_EN                      (PMA_REG_RX_BUSWIDTH_EN),
    .CP_PMA_REG_RX_RATE                             (PMA_REG_RX_RATE),
    .CP_PMA_REG_RX_RESERVED_36                      (PMA_REG_RX_RESERVED_36),
    .CP_PMA_REG_RX_RATE_EN                          (PMA_REG_RX_RATE_EN),
    .CP_PMA_REG_RX_RES_TRIM                         (PMA_REG_RX_RES_TRIM),
    .CP_PMA_REG_RX_RESERVED_44                      (PMA_REG_RX_RESERVED_44),
    .CP_PMA_REG_RX_RESERVED_45                      (PMA_REG_RX_RESERVED_45),
    .CP_PMA_REG_RX_SIGDET_STATUS_EN                 (PMA_REG_RX_SIGDET_STATUS_EN),
    .CP_PMA_REG_RX_RESERVED_48_47                   (PMA_REG_RX_RESERVED_48_47),
    .CP_PMA_REG_RX_ICTRL_SIGDET                     (PMA_REG_RX_ICTRL_SIGDET),
    .CP_PMA_REG_CDR_READY_THD                       (PMA_REG_CDR_READY_THD),
    .CP_PMA_REG_RX_RESERVED_65                      (PMA_REG_RX_RESERVED_65),
    .CP_PMA_REG_RX_PCLK_EDGE_SEL                    (PMA_REG_RX_PCLK_EDGE_SEL),
    .CP_PMA_REG_RX_PIBUF_IC                         (PMA_REG_RX_PIBUF_IC),
    .CP_PMA_REG_RX_RESERVED_69                      (PMA_REG_RX_RESERVED_69),
    .CP_PMA_REG_RX_DCC_IC_RX                        (PMA_REG_RX_DCC_IC_RX),
    .CP_PMA_REG_CDR_READY_CHECK_CTRL                (PMA_REG_CDR_READY_CHECK_CTRL),
    .CP_PMA_REG_RX_ICTRL_TRX                        (PMA_REG_RX_ICTRL_TRX),
    .CP_PMA_REG_RX_RESERVED_77_76                   (PMA_REG_RX_RESERVED_77_76),
    .CP_PMA_REG_RX_RESERVED_79_78                   (PMA_REG_RX_RESERVED_79_78),
    .CP_PMA_REG_RX_RESERVED_81_80                   (PMA_REG_RX_RESERVED_81_80),
    .CP_PMA_REG_RX_ICTRL_PIBUF                      (PMA_REG_RX_ICTRL_PIBUF),
    .CP_PMA_REG_RX_ICTRL_PI                         (PMA_REG_RX_ICTRL_PI),
    .CP_PMA_REG_RX_ICTRL_DCC                        (PMA_REG_RX_ICTRL_DCC),
    .CP_PMA_REG_RX_RESERVED_89_88                   (PMA_REG_RX_RESERVED_89_88),
    .CP_PMA_REG_TX_RATE                             (PMA_REG_TX_RATE),
    .CP_PMA_REG_RX_RESERVED_92                      (PMA_REG_RX_RESERVED_92),
    .CP_PMA_REG_TX_RATE_EN                          (PMA_REG_TX_RATE_EN),
    .CP_PMA_REG_RX_TX2RX_PLPBK_RST_N                (PMA_REG_RX_TX2RX_PLPBK_RST_N),
    .CP_PMA_REG_RX_TX2RX_PLPBK_RST_N_EN             (PMA_REG_RX_TX2RX_PLPBK_RST_N_EN),
    .CP_PMA_REG_RX_TX2RX_PLPBK_EN                   (PMA_REG_RX_TX2RX_PLPBK_EN),
    .CP_PMA_REG_TXCLK_SEL                           (PMA_REG_TXCLK_SEL),
    .CP_PMA_REG_RX_DATA_POLARITY                    (PMA_REG_RX_DATA_POLARITY),
    .CP_PMA_REG_RX_ERR_INSERT                       (PMA_REG_RX_ERR_INSERT),
    .CP_PMA_REG_UDP_CHK_EN                          (PMA_REG_UDP_CHK_EN),
    .CP_PMA_REG_PRBS_SEL                            (PMA_REG_PRBS_SEL),
    .CP_PMA_REG_PRBS_CHK_EN                         (PMA_REG_PRBS_CHK_EN),
    .CP_PMA_REG_PRBS_CHK_WIDTH_SEL                  (PMA_REG_PRBS_CHK_WIDTH_SEL),
    .CP_PMA_REG_BIST_CHK_PAT_SEL                    (PMA_REG_BIST_CHK_PAT_SEL),
    .CP_PMA_REG_LOAD_ERR_CNT                        (PMA_REG_LOAD_ERR_CNT),
    .CP_PMA_REG_CHK_COUNTER_EN                      (PMA_REG_CHK_COUNTER_EN),
    .CP_PMA_REG_CDR_PROP_GAIN                       (PMA_REG_CDR_PROP_GAIN),
    .CP_PMA_REG_CDR_PROP_TURBO_GAIN                 (PMA_REG_CDR_PROP_TURBO_GAIN),
    .CP_PMA_REG_CDR_INT_GAIN                        (PMA_REG_CDR_INT_GAIN),
    .CP_PMA_REG_CDR_INT_TURBO_GAIN                  (PMA_REG_CDR_INT_TURBO_GAIN),
    .CP_PMA_REG_CDR_INT_SAT_MAX                     (PMA_REG_CDR_INT_SAT_MAX),
    .CP_PMA_REG_CDR_INT_SAT_MIN                     (PMA_REG_CDR_INT_SAT_MIN),
    .CP_PMA_REG_CDR_INT_RST                         (PMA_REG_CDR_INT_RST),
    .CP_PMA_REG_CDR_INT_RST_OW                      (PMA_REG_CDR_INT_RST_OW),
    .CP_PMA_REG_CDR_PROP_RST                        (PMA_REG_CDR_PROP_RST),
    .CP_PMA_REG_CDR_PROP_RST_OW                     (PMA_REG_CDR_PROP_RST_OW),
    .CP_PMA_REG_CDR_LOCK_RST                        (PMA_REG_CDR_LOCK_RST),
    .CP_PMA_REG_CDR_LOCK_RST_OW                     (PMA_REG_CDR_LOCK_RST_OW),
    .CP_PMA_REG_CDR_RX_PI_FORCE_SEL                 (PMA_REG_CDR_RX_PI_FORCE_SEL),
    .CP_PMA_REG_CDR_RX_PI_FORCE_D                   (PMA_REG_CDR_RX_PI_FORCE_D),
    .CP_PMA_REG_CDR_LOCK_TIMER                      (PMA_REG_CDR_LOCK_TIMER),
    .CP_PMA_REG_CDR_TURBO_MODE_TIMER                (PMA_REG_CDR_TURBO_MODE_TIMER),
    .CP_PMA_REG_CDR_LOCK_VAL                        (PMA_REG_CDR_LOCK_VAL),
    .CP_PMA_REG_CDR_LOCK_OW                         (PMA_REG_CDR_LOCK_OW),
    .CP_PMA_REG_CDR_INT_SAT_DET_EN                  (PMA_REG_CDR_INT_SAT_DET_EN),
    .CP_PMA_REG_CDR_SAT_AUTO_DIS                    (PMA_REG_CDR_SAT_AUTO_DIS),
    .CP_PMA_REG_CDR_GAIN_AUTO                       (PMA_REG_CDR_GAIN_AUTO),
    .CP_PMA_REG_CDR_TURBO_GAIN_AUTO                 (PMA_REG_CDR_TURBO_GAIN_AUTO),
    .CP_PMA_REG_RX_RESERVED_171_167                 (PMA_REG_RX_RESERVED_171_167),
    .CP_PMA_REG_RX_RESERVED_175_172                 (PMA_REG_RX_RESERVED_175_172),
    .CP_PMA_REG_CDR_SAT_DET_STATUS_EN               (PMA_REG_CDR_SAT_DET_STATUS_EN),
    .CP_PMA_REG_CDR_SAT_DET_STATUS_RESET_EN         (PMA_REG_CDR_SAT_DET_STATUS_RESET_EN),
    .CP_PMA_REG_CDR_PI_CTRL_RST                     (PMA_REG_CDR_PI_CTRL_RST),
    .CP_PMA_REG_CDR_PI_CTRL_RST_OW                  (PMA_REG_CDR_PI_CTRL_RST_OW),
    .CP_PMA_REG_CDR_SAT_DET_RST                     (PMA_REG_CDR_SAT_DET_RST),
    .CP_PMA_REG_CDR_SAT_DET_RST_OW                  (PMA_REG_CDR_SAT_DET_RST_OW),
    .CP_PMA_REG_CDR_SAT_DET_STICKY_RST              (PMA_REG_CDR_SAT_DET_STICKY_RST),
    .CP_PMA_REG_CDR_SAT_DET_STICKY_RST_OW           (PMA_REG_CDR_SAT_DET_STICKY_RST_OW),
    .CP_PMA_REG_CDR_SIGDET_STATUS_DIS               (PMA_REG_CDR_SIGDET_STATUS_DIS),
    .CP_PMA_REG_CDR_SAT_DET_TIMER                   (PMA_REG_CDR_SAT_DET_TIMER),
    .CP_PMA_REG_CDR_SAT_DET_STATUS_VAL              (PMA_REG_CDR_SAT_DET_STATUS_VAL),
    .CP_PMA_REG_CDR_SAT_DET_STATUS_OW               (PMA_REG_CDR_SAT_DET_STATUS_OW),
    .CP_PMA_REG_CDR_TURBO_MODE_EN                   (PMA_REG_CDR_TURBO_MODE_EN),
    .CP_PMA_REG_RX_RESERVED_190                     (PMA_REG_RX_RESERVED_190),
    .CP_PMA_REG_RX_RESERVED_193_191                 (PMA_REG_RX_RESERVED_193_191),
    .CP_PMA_REG_CDR_STATUS_FIFO_EN                  (PMA_REG_CDR_STATUS_FIFO_EN),
    .CP_PMA_REG_PMA_TEST_SEL                        (PMA_REG_PMA_TEST_SEL),
    .CP_PMA_REG_OOB_COMWAKE_GAP_MIN                 (PMA_REG_OOB_COMWAKE_GAP_MIN),
    .CP_PMA_REG_OOB_COMWAKE_GAP_MAX                 (PMA_REG_OOB_COMWAKE_GAP_MAX),
    .CP_PMA_REG_OOB_COMINIT_GAP_MIN                 (PMA_REG_OOB_COMINIT_GAP_MIN),
    .CP_PMA_REG_OOB_COMINIT_GAP_MAX                 (PMA_REG_OOB_COMINIT_GAP_MAX),
    .CP_PMA_REG_RX_RESERVED_227_226                 (PMA_REG_RX_RESERVED_227_226),
    .CP_PMA_REG_COMWAKE_STATUS_CLEAR                (PMA_REG_COMWAKE_STATUS_CLEAR),
    .CP_PMA_REG_COMINIT_STATUS_CLEAR                (PMA_REG_COMINIT_STATUS_CLEAR),
    .CP_PMA_REG_RX_SYNC_RST_N_EN                    (PMA_REG_RX_SYNC_RST_N_EN),
    .CP_PMA_REG_RX_SYNC_RST_N                       (PMA_REG_RX_SYNC_RST_N),
    .CP_PMA_REG_RX_RESERVED_233_232                 (PMA_REG_RX_RESERVED_233_232),
    .CP_PMA_REG_RX_RESERVED_235_234                 (PMA_REG_RX_RESERVED_235_234),
    .CP_PMA_REG_RX_SATA_COMINIT_OW                  (PMA_REG_RX_SATA_COMINIT_OW),
    .CP_PMA_REG_RX_SATA_COMINIT                     (PMA_REG_RX_SATA_COMINIT),
    .CP_PMA_REG_RX_SATA_COMWAKE_OW                  (PMA_REG_RX_SATA_COMWAKE_OW),
    .CP_PMA_REG_RX_SATA_COMWAKE                     (PMA_REG_RX_SATA_COMWAKE),
    .CP_PMA_REG_RX_RESERVED_241_240                 (PMA_REG_RX_RESERVED_241_240),
    .CP_PMA_REG_RX_DCC_DISABLE                      (PMA_REG_RX_DCC_DISABLE),
    .CP_PMA_REG_RX_RESERVED_243                     (PMA_REG_RX_RESERVED_243),
    .CP_PMA_REG_RX_SLIP_SEL_EN                      (PMA_REG_RX_SLIP_SEL_EN),
    .CP_PMA_REG_RX_SLIP_SEL                         (PMA_REG_RX_SLIP_SEL),
    .CP_PMA_REG_RX_SLIP_EN                          (PMA_REG_RX_SLIP_EN),
    .CP_PMA_REG_RX_SIGDET_STATUS_SEL                (PMA_REG_RX_SIGDET_STATUS_SEL),
    .CP_PMA_REG_RX_SIGDET_FSM_RST_N                 (PMA_REG_RX_SIGDET_FSM_RST_N),
    .CP_PMA_REG_RX_RESERVED_254                     (PMA_REG_RX_RESERVED_254),
    .CP_PMA_REG_RX_SIGDET_STATUS                    (PMA_REG_RX_SIGDET_STATUS),
    .CP_PMA_REG_RX_SIGDET_VTH                       (PMA_REG_RX_SIGDET_VTH),
    .CP_PMA_REG_RX_SIGDET_GRM                       (PMA_REG_RX_SIGDET_GRM),
    .CP_PMA_REG_RX_SIGDET_PULSE_EXT                 (PMA_REG_RX_SIGDET_PULSE_EXT),
    .CP_PMA_REG_RX_SIGDET_CH2_SEL                   (PMA_REG_RX_SIGDET_CH2_SEL),
    .CP_PMA_REG_RX_SIGDET_CH2_CHK_WINDOW            (PMA_REG_RX_SIGDET_CH2_CHK_WINDOW),
    .CP_PMA_REG_RX_SIGDET_CHK_WINDOW_EN             (PMA_REG_RX_SIGDET_CHK_WINDOW_EN),
    .CP_PMA_REG_RX_SIGDET_NOSIG_COUNT_SETTING       (PMA_REG_RX_SIGDET_NOSIG_COUNT_SETTING),
    .CP_PMA_REG_SLIP_FIFO_INV_EN                    (PMA_REG_SLIP_FIFO_INV_EN),
    .CP_PMA_REG_SLIP_FIFO_INV                       (PMA_REG_SLIP_FIFO_INV),
    .CP_PMA_REG_RX_SIGDET_OOB_DET_COUNT_VAL         (PMA_REG_RX_SIGDET_OOB_DET_COUNT_VAL),
    .CP_PMA_REG_RX_SIGDET_4OOB_DET_SEL              (PMA_REG_RX_SIGDET_4OOB_DET_SEL),
    .CP_PMA_REG_RX_RESERVED_285_283                 (PMA_REG_RX_RESERVED_285_283),
    .CP_PMA_REG_RX_RESERVED_286                     (PMA_REG_RX_RESERVED_286),
    .CP_PMA_REG_RX_SIGDET_IC_I                      (PMA_REG_RX_SIGDET_IC_I),
    .CP_PMA_REG_RX_OOB_DETECTOR_RESET_N_OW          (PMA_REG_RX_OOB_DETECTOR_RESET_N_OW),
    .CP_PMA_REG_RX_OOB_DETECTOR_RESET_N             (PMA_REG_RX_OOB_DETECTOR_RESET_N),
    .CP_PMA_REG_RX_OOB_DETECTOR_PD_OW               (PMA_REG_RX_OOB_DETECTOR_PD_OW),
    .CP_PMA_REG_RX_OOB_DETECTOR_PD                  (PMA_REG_RX_OOB_DETECTOR_PD),
    .CP_PMA_REG_RX_LS_MODE_EN                       (PMA_REG_RX_LS_MODE_EN),
    .CP_PMA_REG_ANA_RX_EQ1_R_SET_FB_O_SEL           (PMA_REG_ANA_RX_EQ1_R_SET_FB_O_SEL),
    .CP_PMA_REG_ANA_RX_EQ2_R_SET_FB_O_SEL           (PMA_REG_ANA_RX_EQ2_R_SET_FB_O_SEL),
    .CP_PMA_REG_RX_EQ1_R_SET_TOP                    (PMA_REG_RX_EQ1_R_SET_TOP),
    .CP_PMA_REG_RX_EQ1_R_SET_FB                     (PMA_REG_RX_EQ1_R_SET_FB),
    .CP_PMA_REG_RX_EQ1_C_SET_FB                     (PMA_REG_RX_EQ1_C_SET_FB),
    .CP_PMA_REG_RX_EQ1_OFF                          (PMA_REG_RX_EQ1_OFF),
    .CP_PMA_REG_RX_EQ2_R_SET_TOP                    (PMA_REG_RX_EQ2_R_SET_TOP),
    .CP_PMA_REG_RX_EQ2_R_SET_FB                     (PMA_REG_RX_EQ2_R_SET_FB),
    .CP_PMA_REG_RX_EQ2_C_SET_FB                     (PMA_REG_RX_EQ2_C_SET_FB),
    .CP_PMA_REG_RX_EQ2_OFF                          (PMA_REG_RX_EQ2_OFF),
    .CP_PMA_REG_EQ_DAC                              (PMA_REG_EQ_DAC),
    .CP_PMA_REG_RX_ICTRL_EQ                         (PMA_REG_RX_ICTRL_EQ),
    .CP_PMA_REG_EQ_DC_CALIB_EN                      (PMA_REG_EQ_DC_CALIB_EN),
    .CP_PMA_REG_EQ_DC_CALIB_SEL                     (PMA_REG_EQ_DC_CALIB_SEL),
    .CP_PMA_REG_RX_RESERVED_337_330                 (PMA_REG_RX_RESERVED_337_330),
    .CP_PMA_REG_RX_RESERVED_345_338                 (PMA_REG_RX_RESERVED_345_338),
    .CP_PMA_REG_RX_RESERVED_353_346                 (PMA_REG_RX_RESERVED_353_346),
    .CP_PMA_REG_RX_RESERVED_361_354                 (PMA_REG_RX_RESERVED_361_354),
    .CP_PMA_CTLE_CTRL_REG_I                         (PMA_CTLE_CTRL_REG_I),
    .CP_PMA_CTLE_REG_FORCE_SEL_I                    (PMA_CTLE_REG_FORCE_SEL_I),
    .CP_PMA_CTLE_REG_HOLD_I                         (PMA_CTLE_REG_HOLD_I),
    .CP_PMA_CTLE_REG_INIT_DAC_I                     (PMA_CTLE_REG_INIT_DAC_I),
    .CP_PMA_CTLE_REG_POLARITY_I                     (PMA_CTLE_REG_POLARITY_I),
    .CP_PMA_CTLE_REG_SHIFTER_GAIN_I                 (PMA_CTLE_REG_SHIFTER_GAIN_I),        
    .CP_PMA_CTLE_REG_THRESHOLD_I                    (PMA_CTLE_REG_THRESHOLD_I),
    .CP_PMA_REG_RX_RES_TRIM_EN                      (PMA_REG_RX_RES_TRIM_EN),
    .CP_PMA_REG_RX_RESERVED_393_389                 (PMA_REG_RX_RESERVED_393_389),
    .CP_PMA_CFG_RX_LANE_POWERUP                     (PMA_CFG_RX_LANE_POWERUP),
    .CP_PMA_CFG_RX_PMA_RSTN                         (PMA_CFG_RX_PMA_RSTN),
    .CP_PMA_INT_PMA_RX_MASK_0                       (PMA_INT_PMA_RX_MASK_0),
    .CP_PMA_INT_PMA_RX_CLR_0                        (PMA_INT_PMA_RX_CLR_0),
    .CP_PMA_CFG_CTLE_ADP_RSTN                       (PMA_CFG_CTLE_ADP_RSTN),
 
    //pma_tx
    .CP_PMA_REG_TX_PD                               (PMA_REG_TX_PD),  
    .CP_PMA_REG_TX_PD_OW                            (PMA_REG_TX_PD_OW),
    .CP_PMA_REG_TX_MAIN_PRE_Z                       (PMA_REG_TX_MAIN_PRE_Z),
    .CP_PMA_REG_TX_MAIN_PRE_Z_OW                    (PMA_REG_TX_MAIN_PRE_Z_OW),
    .CP_PMA_REG_TX_BEACON_TIMER_SEL                 (PMA_REG_TX_BEACON_TIMER_SEL),
    .CP_PMA_REG_TX_RXDET_REQ_OW                     (PMA_REG_TX_RXDET_REQ_OW),
    .CP_PMA_REG_TX_RXDET_REQ                        (PMA_REG_TX_RXDET_REQ),
    .CP_PMA_REG_TX_BEACON_EN_OW                     (PMA_REG_TX_BEACON_EN_OW),
    .CP_PMA_REG_TX_BEACON_EN                        (PMA_REG_TX_BEACON_EN),
    .CP_PMA_REG_TX_EI_EN_OW                         (PMA_REG_TX_EI_EN_OW),
    .CP_PMA_REG_TX_EI_EN                            (PMA_REG_TX_EI_EN),
    .CP_PMA_REG_TX_BIT_CONV                         (PMA_REG_TX_BIT_CONV),
    .CP_PMA_REG_TX_RES_CAL                          (PMA_REG_TX_RES_CAL),
    .CP_PMA_REG_TX_RESERVED_19                      (PMA_REG_TX_RESERVED_19),
    .CP_PMA_REG_TX_RESERVED_25_20                   (PMA_REG_TX_RESERVED_25_20),
    .CP_PMA_REG_TX_RESERVED_33_26                   (PMA_REG_TX_RESERVED_33_26),
    .CP_PMA_REG_TX_RESERVED_41_34                   (PMA_REG_TX_RESERVED_41_34),
    .CP_PMA_REG_TX_RESERVED_49_42                   (PMA_REG_TX_RESERVED_49_42),
    .CP_PMA_REG_TX_RESERVED_57_50                   (PMA_REG_TX_RESERVED_57_50),
    .CP_PMA_REG_TX_SYNC_OW                          (PMA_REG_TX_SYNC_OW),
    .CP_PMA_REG_TX_SYNC                             (PMA_REG_TX_SYNC),
    .CP_PMA_REG_TX_PD_POST                          (PMA_REG_TX_PD_POST),
    .CP_PMA_REG_TX_PD_POST_OW                       (PMA_REG_TX_PD_POST_OW),
    .CP_PMA_REG_TX_RESET_N_OW                       (PMA_REG_TX_RESET_N_OW),
    .CP_PMA_REG_TX_RESET_N                          (PMA_REG_TX_RESET_N),
    .CP_PMA_REG_TX_RESERVED_64                      (PMA_REG_TX_RESERVED_64),
    .CP_PMA_REG_TX_RESERVED_65                      (PMA_REG_TX_RESERVED_65),
    .CP_PMA_REG_TX_BUSWIDTH_OW                      (PMA_REG_TX_BUSWIDTH_OW),
    .CP_PMA_REG_TX_BUSWIDTH                         (PMA_REG_TX_BUSWIDTH),
    .CP_PMA_REG_PLL_READY_OW                        (PMA_REG_PLL_READY_OW),
    .CP_PMA_REG_PLL_READY                           (PMA_REG_PLL_READY),
    .CP_PMA_REG_TX_RESERVED_72                      (PMA_REG_TX_RESERVED_72),
    .CP_PMA_REG_TX_RESERVED_73                      (PMA_REG_TX_RESERVED_73),
    .CP_PMA_REG_TX_RESERVED_74                      (PMA_REG_TX_RESERVED_74),
    .CP_PMA_REG_EI_PCLK_DELAY_SEL                   (PMA_REG_EI_PCLK_DELAY_SEL),
    .CP_PMA_REG_TX_RESERVED_77                      (PMA_REG_TX_RESERVED_77),
    .CP_PMA_REG_TX_RESERVED_83_78                   (PMA_REG_TX_RESERVED_83_78),
    .CP_PMA_REG_TX_RESERVED_89_84                   (PMA_REG_TX_RESERVED_89_84),
    .CP_PMA_REG_TX_RESERVED_95_90                   (PMA_REG_TX_RESERVED_95_90),
    .CP_PMA_REG_TX_RESERVED_101_96                  (PMA_REG_TX_RESERVED_101_96),
    .CP_PMA_REG_TX_RESERVED_107_102                 (PMA_REG_TX_RESERVED_107_102),
    .CP_PMA_REG_TX_RESERVED_113_108                 (PMA_REG_TX_RESERVED_113_108),
    .CP_PMA_REG_TX_AMP_DAC0                         (PMA_REG_TX_AMP_DAC0),
    .CP_PMA_REG_TX_AMP_DAC1                         (PMA_REG_TX_AMP_DAC1),
    .CP_PMA_REG_TX_AMP_DAC2                         (PMA_REG_TX_AMP_DAC2),
    .CP_PMA_REG_TX_AMP_DAC3                         (PMA_REG_TX_AMP_DAC3),
    .CP_PMA_REG_TX_RESERVED_143_138                 (PMA_REG_TX_RESERVED_143_138),
    .CP_PMA_REG_TX_MARGIN                           (PMA_REG_TX_MARGIN),
    .CP_PMA_REG_TX_MARGIN_OW                        (PMA_REG_TX_MARGIN_OW),
    .CP_PMA_REG_TX_RESERVED_149_148                 (PMA_REG_TX_RESERVED_149_148),
    .CP_PMA_REG_TX_RESERVED_150                     (PMA_REG_TX_RESERVED_150),
    .CP_PMA_REG_TX_SWING                            (PMA_REG_TX_SWING),
    .CP_PMA_REG_TX_SWING_OW                         (PMA_REG_TX_SWING_OW),
    .CP_PMA_REG_TX_RESERVED_153                     (PMA_REG_TX_RESERVED_153),
    .CP_PMA_REG_TX_RXDET_THRESHOLD                  (PMA_REG_TX_RXDET_THRESHOLD),
    .CP_PMA_REG_TX_RESERVED_157_156                 (PMA_REG_TX_RESERVED_157_156),
    .CP_PMA_REG_TX_BEACON_OSC_CTRL                  (PMA_REG_TX_BEACON_OSC_CTRL),
    .CP_PMA_REG_TX_RESERVED_160_159                 (PMA_REG_TX_RESERVED_160_159),
    .CP_PMA_REG_TX_RESERVED_162_161                 (PMA_REG_TX_RESERVED_162_161),
    .CP_PMA_REG_TX_TX2RX_SLPBACK_EN                 (PMA_REG_TX_TX2RX_SLPBACK_EN),
    .CP_PMA_REG_TX_PCLK_EDGE_SEL                    (PMA_REG_TX_PCLK_EDGE_SEL),
    .CP_PMA_REG_TX_RXDET_STATUS_OW                  (PMA_REG_TX_RXDET_STATUS_OW),
    .CP_PMA_REG_TX_RXDET_STATUS                     (PMA_REG_TX_RXDET_STATUS),
    .CP_PMA_REG_TX_PRBS_GEN_EN                      (PMA_REG_TX_PRBS_GEN_EN),
    .CP_PMA_REG_TX_PRBS_GEN_WIDTH_SEL               (PMA_REG_TX_PRBS_GEN_WIDTH_SEL),
    .CP_PMA_REG_TX_PRBS_SEL                         (PMA_REG_TX_PRBS_SEL),
    .CP_PMA_REG_TX_UDP_DATA_7_TO_0                  (PMA_REG_TX_UDP_DATA_7_TO_0),
    .CP_PMA_REG_TX_UDP_DATA_15_TO_8                 (PMA_REG_TX_UDP_DATA_15_TO_8),
    .CP_PMA_REG_TX_UDP_DATA_19_TO_16                (PMA_REG_TX_UDP_DATA_19_TO_16),
    .CP_PMA_REG_TX_RESERVED_192                     (PMA_REG_TX_RESERVED_192),
    .CP_PMA_REG_TX_FIFO_WP_CTRL                     (PMA_REG_TX_FIFO_WP_CTRL),
    .CP_PMA_REG_TX_FIFO_EN                          (PMA_REG_TX_FIFO_EN),
    .CP_PMA_REG_TX_DATA_MUX_SEL                     (PMA_REG_TX_DATA_MUX_SEL),
    .CP_PMA_REG_TX_ERR_INSERT                       (PMA_REG_TX_ERR_INSERT),
    .CP_PMA_REG_TX_RESERVED_203_200                 (PMA_REG_TX_RESERVED_203_200),
    .CP_PMA_REG_TX_RESERVED_204                     (PMA_REG_TX_RESERVED_204),
    .CP_PMA_REG_TX_SATA_EN                          (PMA_REG_TX_SATA_EN),
    .CP_PMA_REG_TX_RESERVED_207_206                 (PMA_REG_TX_RESERVED_207_206),
    .CP_PMA_REG_RATE_CHANGE_TXPCLK_ON_OW            (PMA_REG_RATE_CHANGE_TXPCLK_ON_OW),
    .CP_PMA_REG_RATE_CHANGE_TXPCLK_ON               (PMA_REG_RATE_CHANGE_TXPCLK_ON),
    .CP_PMA_REG_TX_CFG_POST1                        (PMA_REG_TX_CFG_POST1),
    .CP_PMA_REG_TX_CFG_POST2                        (PMA_REG_TX_CFG_POST2),
    .CP_PMA_REG_TX_DEEMP                            (PMA_REG_TX_DEEMP),
    .CP_PMA_REG_TX_DEEMP_OW                         (PMA_REG_TX_DEEMP_OW),
    .CP_PMA_REG_TX_RESERVED_224_223                 (PMA_REG_TX_RESERVED_224_223),
    .CP_PMA_REG_TX_RESERVED_225                     (PMA_REG_TX_RESERVED_225),
    .CP_PMA_REG_TX_RESERVED_229_226                 (PMA_REG_TX_RESERVED_229_226),
    .CP_PMA_REG_TX_OOB_DELAY_SEL                    (PMA_REG_TX_OOB_DELAY_SEL),
    .CP_PMA_REG_TX_POLARITY                         (PMA_REG_TX_POLARITY),
    .CP_PMA_REG_ANA_TX_JTAG_DATA_O_SEL              (PMA_REG_ANA_TX_JTAG_DATA_O_SEL),
    .CP_PMA_REG_TX_RESERVED_236                     (PMA_REG_TX_RESERVED_236),
    .CP_PMA_REG_TX_LS_MODE_EN                       (PMA_REG_TX_LS_MODE_EN),
    .CP_PMA_REG_TX_JTAG_MODE_EN_OW                  (PMA_REG_TX_JTAG_MODE_EN_OW),
    .CP_PMA_REG_TX_JTAG_MODE_EN                     (PMA_REG_TX_JTAG_MODE_EN),
    .CP_PMA_REG_RX_JTAG_MODE_EN_OW                  (PMA_REG_RX_JTAG_MODE_EN_OW),
    .CP_PMA_REG_RX_JTAG_MODE_EN                     (PMA_REG_RX_JTAG_MODE_EN),
    .CP_PMA_REG_RX_JTAG_OE                          (PMA_REG_RX_JTAG_OE),
    .CP_PMA_REG_RX_ACJTAG_VHYSTSEL                  (PMA_REG_RX_ACJTAG_VHYSTSEL),
    .CP_PMA_REG_TX_RES_CAL_EN                       (PMA_REG_TX_RES_CAL_EN),
    .CP_PMA_REG_RX_TERM_MODE_CTRL                   (PMA_REG_RX_TERM_MODE_CTRL),
    .CP_PMA_REG_TX_RESERVED_251_250                 (PMA_REG_TX_RESERVED_251_250),
    .CP_PMA_REG_PLPBK_TXPCLK_EN                     (PMA_REG_PLPBK_TXPCLK_EN),
    .CP_PMA_REG_TX_RESERVED_253                     (PMA_REG_TX_RESERVED_253),
    .CP_PMA_REG_TX_RESERVED_254                     (PMA_REG_TX_RESERVED_254),
    .CP_PMA_REG_TX_RESERVED_255                     (PMA_REG_TX_RESERVED_255),
    .CP_PMA_REG_TX_RESERVED_256                     (PMA_REG_TX_RESERVED_256),
    .CP_PMA_REG_TX_RESERVED_257                     (PMA_REG_TX_RESERVED_257),
    .CP_PMA_REG_TX_PH_SEL                           (PMA_REG_TX_PH_SEL),
    .CP_PMA_REG_TX_CFG_PRE                          (PMA_REG_TX_CFG_PRE), 
    .CP_PMA_REG_TX_CFG_MAIN                         (PMA_REG_TX_CFG_MAIN),
    .CP_PMA_REG_CFG_POST                            (PMA_REG_CFG_POST),
    .CP_PMA_REG_PD_MAIN                             (PMA_REG_PD_MAIN),
    .CP_PMA_REG_PD_PRE                              (PMA_REG_PD_PRE),
    .CP_PMA_REG_TX_LS_DATA                          (PMA_REG_TX_LS_DATA),
    .CP_PMA_REG_TX_DCC_BUF_SZ_SEL                   (PMA_REG_TX_DCC_BUF_SZ_SEL),
    .CP_PMA_REG_TX_DCC_CAL_CUR_TUNE                 (PMA_REG_TX_DCC_CAL_CUR_TUNE),
    .CP_PMA_REG_TX_DCC_CAL_EN                       (PMA_REG_TX_DCC_CAL_EN),
    .CP_PMA_REG_TX_DCC_CUR_SS                       (PMA_REG_TX_DCC_CUR_SS),
    .CP_PMA_REG_TX_DCC_FA_CTRL                      (PMA_REG_TX_DCC_FA_CTRL),
    .CP_PMA_REG_TX_DCC_RI_CTRL                      (PMA_REG_TX_DCC_RI_CTRL),
    .CP_PMA_REG_ATB_SEL_2_TO_0                      (PMA_REG_ATB_SEL_2_TO_0),
    .CP_PMA_REG_ATB_SEL_9_TO_3                      (PMA_REG_ATB_SEL_9_TO_3),
    .CP_PMA_REG_TX_CFG_7_TO_0                       (PMA_REG_TX_CFG_7_TO_0),
    .CP_PMA_REG_TX_CFG_15_TO_8                      (PMA_REG_TX_CFG_15_TO_8),
    .CP_PMA_REG_TX_CFG_23_TO_16                     (PMA_REG_TX_CFG_23_TO_16),
    .CP_PMA_REG_TX_CFG_31_TO_24                     (PMA_REG_TX_CFG_31_TO_24),
    .CP_PMA_REG_TX_OOB_EI_EN                        (PMA_REG_TX_OOB_EI_EN),
    .CP_PMA_REG_TX_OOB_EI_EN_OW                     (PMA_REG_TX_OOB_EI_EN_OW),
    .CP_PMA_REG_TX_BEACON_EN_DELAYED                (PMA_REG_TX_BEACON_EN_DELAYED),
    .CP_PMA_REG_TX_BEACON_EN_DELAYED_OW             (PMA_REG_TX_BEACON_EN_DELAYED_OW),
    .CP_PMA_REG_TX_JTAG_DATA                        (PMA_REG_TX_JTAG_DATA),
    .CP_PMA_REG_TX_RXDET_TIMER_SEL                  (PMA_REG_TX_RXDET_TIMER_SEL),
    .CP_PMA_REG_TX_CFG1_7_0                         (PMA_REG_TX_CFG1_7_0),
    .CP_PMA_REG_TX_CFG1_15_8                        (PMA_REG_TX_CFG1_15_8),
    .CP_PMA_REG_TX_CFG1_23_16                       (PMA_REG_TX_CFG1_23_16),
    .CP_PMA_REG_TX_CFG1_31_24                       (PMA_REG_TX_CFG1_31_24),
    .CP_PMA_REG_CFG_LANE_POWERUP                    (PMA_REG_CFG_LANE_POWERUP),
    .CP_PMA_REG_CFG_PMA_POR_N                       ("TRUE"),
    .CP_PMA_REG_CFG_TX_LANE_POWERUP_CLKPATH         (PMA_REG_CFG_TX_LANE_POWERUP_CLKPATH),
    .CP_PMA_REG_CFG_TX_LANE_POWERUP_PISO            (PMA_REG_CFG_TX_LANE_POWERUP_PISO),
    .CP_PMA_REG_CFG_TX_LANE_POWERUP_DRIVER          (PMA_REG_CFG_TX_LANE_POWERUP_DRIVER),
    .CP_PMA_REG_CFG_TX_PMA_RSTN                     ("TRUE"),
    
    //global
    .CP_GRSN_DIS                                    ("FALSE"),
    .CP_HSST_EN                                     ("TRUE"),
    .CP_CFG_RSTN                                    ("TRUE")

) U0_HSSTLP_LANE (
//////////PAD/////////////////////////////////////////////////////////
    //output
    .PAD_TX_SDN                                     (P_TX_SDN),  
    .PAD_TX_SDP                                     (P_TX_SDP),    

    //input
    .PAD_RX_SDN                                     (P_RX_SDN),
    .PAD_RX_SDP                                     (P_RX_SDP),

//////////SRB related/////////////////////////////////////////////////////////
    //output
    .PCS_RX_MCB_STATUS                              (P_PCS_RX_MCB_STATUS), 
    .PCS_LSM_SYNCED                                 (P_PCS_LSM_SYNCED),
    .CFG_READY                                      (P_CFG_READY),
    .CFG_RDATA                                      (P_CFG_RDATA), 
    .CFG_INT                                        (P_CFG_INT),  
    .RDATA                                          (P_RDATA), 
    .RCLK2FABRIC                                    (P_RCLK2FABRIC), 
    .TCLK2FABRIC                                    (P_TCLK2FABRIC), 

    .RX_SIGDET_STATUS                               (P_RX_SIGDET_STATUS), 
    .RX_SATA_COMINIT                                (P_RX_SATA_COMINIT), 
    .RX_SATA_COMWAKE                                (P_RX_SATA_COMWAKE), 
    .RX_LS_DATA                                     (P_RX_LS_DATA), 
    .RX_READY                                       (P_RX_READY), 
    .TEST_STATUS                                    (P_TEST_STATUS), 
    .TX_RXDET_STATUS                                (P_TX_RXDET_STATUS), 
    .CA_ALIGN_RX                                    (P_CA_ALIGN_RX), 
    .CA_ALIGN_TX                                    (P_CA_ALIGN_TX), 

    //input
    .RX_CLK_FR_CORE                                 (P_RX_CLK_FR_CORE),
    .RCLK2_FR_CORE                                  (P_RCLK2_FR_CORE),
    .TX_CLK_FR_CORE                                 (P_TX_CLK_FR_CORE),
    .TCLK2_FR_CORE                                  (P_TCLK2_FR_CORE),
    .HSST_RST                                       (1'b0),
    .PCS_TX_RST                                     (P_PCS_TX_RST),
    .PCS_RX_RST                                     (P_PCS_RX_RST),
    .PCS_CB_RST                                     (P_PCS_CB_RST),
    .RXGEAR_SLIP                                    (P_RXGEAR_SLIP),
    .CFG_CLK                                        (P_CFG_CLK),
    .CFG_RST                                        (P_CFG_RST),
    .CFG_PSEL                                       (P_CFG_PSEL),
    .CFG_ENABLE                                     (P_CFG_ENABLE),
    .CFG_WRITE                                      (P_CFG_WRITE),
    .CFG_ADDR                                       (P_CFG_ADDR),
    .CFG_WDATA                                      (P_CFG_WDATA),
    .TDATA                                          (P_TDATA),
    .PCS_WORD_ALIGN_EN                              (P_PCS_WORD_ALIGN_EN),
    .RX_POLARITY_INVERT                             (P_RX_POLARITY_INVERT),
    .CEB_ADETECT_EN                                 (P_CEB_ADETECT_EN),
    .PCS_MCB_EXT_EN                                 (P_PCS_MCB_EXT_EN),
    .PCS_NEAREND_LOOP                               (P_PCS_NEAREND_LOOP),
    .PCS_FAREND_LOOP                                (P_PCS_FAREND_LOOP),
    .PMA_NEAREND_PLOOP                              (P_PMA_NEAREND_PLOOP),
    .PMA_NEAREND_SLOOP                              (P_PMA_NEAREND_SLOOP),
    .PMA_FAREND_PLOOP                               (P_PMA_FAREND_PLOOP),

    .LANE_PD                                        (P_LANE_PD),
    .LANE_RST                                       (P_LANE_RST),
    .RX_LANE_PD                                     (P_RX_LANE_PD),
    .RX_PMA_RST                                     (P_RX_PMA_RST),
    .CTLE_ADP_RST                                   (P_CTLE_ADP_RST),
    .TX_DEEMP                                       (P_TX_DEEMP),
    .TX_LS_DATA                                     (P_TX_LS_DATA),
    .TX_BEACON_EN                                   (P_TX_BEACON_EN),
    .TX_SWING                                       (P_TX_SWING),
    .TX_RXDET_REQ                                   (P_TX_RXDET_REQ),
    .TX_RATE                                        (P_TX_RATE),
    .TX_BUSWIDTH                                    (P_TX_BUSWIDTH),
    .TX_MARGIN                                      (P_TX_MARGIN),
    .TX_PMA_RST                                     (P_TX_PMA_RST),
    .TX_LANE_PD_CLKPATH                             (P_TX_LANE_PD_CLKPATH),
    .TX_LANE_PD_PISO                                (P_TX_LANE_PD_PISO),
    .TX_LANE_PD_DRIVER                              (P_TX_LANE_PD_DRIVER),
    .RX_RATE                                        (P_RX_RATE),
    .RX_BUSWIDTH                                    (P_RX_BUSWIDTH),
    .RX_HIGHZ                                       (P_RX_HIGHZ),
    .CIM_CLK_ALIGNER_RX                             (P_CIM_CLK_ALIGNER_RX),
    .CIM_CLK_ALIGNER_TX                             (P_CIM_CLK_ALIGNER_TX),
    .CIM_DYN_DLY_SEL_RX                             (P_CIM_DYN_DLY_SEL_RX),
    .CIM_DYN_DLY_SEL_TX                             (P_CIM_DYN_DLY_SEL_TX),
    .CIM_START_ALIGN_RX                             (P_CIM_START_ALIGN_RX),
    .CIM_START_ALIGN_TX                             (P_CIM_START_ALIGN_TX),

//////////New Added/////////////////////////////////////////////////////////
    //output
    .PMA_RCLK                                       (PMA_RCLK),

    //input
    .MCB_RCLK                                       (MCB_RCLK),
    .SYNC                                           (SYNC),
    .RATE_CHANGE                                    (RATE_CHANGE),
    .PLL_LOCK_SEL                                   (PLL_LOCK_SEL),

//////////cin and cout/////////////////////////////////////////////////////////
    //output
    .RFIFO_EN_CB_COUT                               (LANE_COUT_BUS_FORWARD[18]), 
    .RFIFO_EN_AFTER_CTC_COUT                        (LANE_COUT_BUS_FORWARD[17]), 
    .RFIFO_EN_AFTER_CTC_GB_COUT                     (LANE_COUT_BUS_FORWARD[16]), 
    .RFIFO_EN_BRIDGE_COUT                           (LANE_COUT_BUS_FORWARD[15]), 
    .TFIFO_EN_PCS_TX_COUT                           (LANE_COUT_BUS_FORWARD[14]), 
    .TFIFO_EN_BRIDGE_COUT                           (LANE_COUT_BUS_FORWARD[13]), 
    .PCS_TCLK_EN_COUT                               (LANE_COUT_BUS_FORWARD[12]), 
    .GEAR_TCLK_EN_COUT                              (LANE_COUT_BUS_FORWARD[11]), 
    .APATTERN_MATCH_LSB_COUT                        (LANE_COUT_BUS_FORWARD[10]), 
    .APATTERN_MATCH_MSB_COUT                        (LANE_COUT_BUS_FORWARD[9]), 
    .APATTERN_SEACHING_PROC_COUT                    (LANE_COUT_BUS_FORWARD[8]), 
    .CB_RCLK_EN_COUT                                (LANE_COUT_BUS_FORWARD[7]), 
    .AFTER_CTC_RCLK_EN_COUT                         (LANE_COUT_BUS_FORWARD[6]), 
    .AFTER_CTC_RCLK_EN_GB_COUT                      (LANE_COUT_BUS_FORWARD[5]), 
    .SKIP_ADD_MCB_COUT                              (LANE_COUT_BUS_FORWARD[4]), 
    .SKIP_DEL_MCB_COUT                              (LANE_COUT_BUS_FORWARD[3]), 
    .SKIP_DEL_LSB_MCB_COUT                          (LANE_COUT_BUS_FORWARD[2]), 
    .SKIP_ADD_LSB_MCB_COUT                          (LANE_COUT_BUS_FORWARD[1]), 
    .CTC_RD_FIFO_COUT                               (LANE_COUT_BUS_FORWARD[0]), 

    .APATTERN_STATUS_COUT                           (APATTERN_STATUS_COUT), 

    //input
    .RFIFO_EN_CB_CIN                                (LANE_CIN_BUS_FORWARD[18]),
    .RFIFO_EN_AFTER_CTC_CIN                         (LANE_CIN_BUS_FORWARD[17]),
    .RFIFO_EN_AFTER_CTC_GB_CIN                      (LANE_CIN_BUS_FORWARD[16]),
    .RFIFO_EN_BRIDGE_CIN                            (LANE_CIN_BUS_FORWARD[15]),
    .TFIFO_EN_PCS_TX_CIN                            (LANE_CIN_BUS_FORWARD[14]),
    .TFIFO_EN_BRIDGE_CIN                            (LANE_CIN_BUS_FORWARD[13]),
    .PCS_TCLK_EN_CIN                                (LANE_CIN_BUS_FORWARD[12]),
    .GEAR_TCLK_EN_CIN                               (LANE_CIN_BUS_FORWARD[11]),
    .APATTERN_MATCH_LSB_CIN                         (LANE_CIN_BUS_FORWARD[10]),
    .APATTERN_MATCH_MSB_CIN                         (LANE_CIN_BUS_FORWARD[9]),
    .APATTERN_SEACHING_PROC_CIN                     (LANE_CIN_BUS_FORWARD[8]),
    .CB_RCLK_EN_CIN                                 (LANE_CIN_BUS_FORWARD[7]),
    .AFTER_CTC_RCLK_EN_CIN                          (LANE_CIN_BUS_FORWARD[6]),
    .AFTER_CTC_RCLK_EN_GB_CIN                       (LANE_CIN_BUS_FORWARD[5]),
    .SKIP_ADD_MCB_CIN                               (LANE_CIN_BUS_FORWARD[4]),
    .SKIP_DEL_MCB_CIN                               (LANE_CIN_BUS_FORWARD[3]),
    .SKIP_DEL_LSB_MCB_CIN                           (LANE_CIN_BUS_FORWARD[2]),
    .SKIP_ADD_LSB_MCB_CIN                           (LANE_CIN_BUS_FORWARD[1]),
    .CTC_RD_FIFO_CIN                                (LANE_CIN_BUS_FORWARD[0]),

    .APATTERN_STATUS_CIN                            (APATTERN_STATUS_CIN),

//////////From PLL/////////////////////////////////////////////////////////
    .CLK_TXP                                        (CLK_TXP),
    .CLK_TXN                                        (CLK_TXN),
    .CLK_RX0                                        (CLK_RX0),
    .CLK_RX90                                       (CLK_RX90),
    .CLK_RX180                                      (CLK_RX180),
    .CLK_RX270                                      (CLK_RX270),

    .PLL_PD_I                                       (PLL_PD_I),
    .PLL_RESET_I                                    (PLL_RESET_I),
    .PLL_REFCLK_I                                   (PLL_REFCLK_I),
    .PLL_RES_TRIM_I                                 (PLL_RES_TRIM_I),

//////////out/////////////////////////////////////////////////////////
    .TXPCLK_PLL                                     (TXPCLK_PLL),

//////////DFT/////////////////////////////////////////////////////////
    .TEST_SO0                                       (),
    .TEST_SO1                                       (),
    .TEST_SO2                                       (),
    .TEST_SO3                                       (),
    .TEST_SO4                                       (),
    .TEST_SE_N                                      (1'b1),
    .TEST_MODE_N                                    (1'b1),
    .TEST_RSTN                                      (),
    .TEST_SI0                                       (),
    .TEST_SI1                                       (),
    .TEST_SI2                                       (),
    .TEST_SI3                                       (),
    .TEST_SI4                                       (),
    
    .FOR_PMA_TEST_SO                                (),
    .FOR_PMA_TEST_MODE_N                            (1'b1),
    .FOR_PMA_TEST_SE_N                              (2'b11),
    .FOR_PMA_TEST_CLK                               (),
    .FOR_PMA_TEST_RSTN                              (),
    .FOR_PMA_TEST_SI                                ()

);

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_INV.v
//
// Functional description: 1-bit Inverter
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_INV
(
    output wire Z,
    input wire I
);

    not (Z, I);

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_DRM36K_E1.v
//
// Functional description:
// Fake module
//
// Parameter  description:
//
// Port description:
//
// Revision history:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_DRM36K_E1
#(
    parameter GRS_EN = "TRUE",
    parameter [2:0] CSA_MASK = 3'b000,
    parameter [2:0] CSB_MASK = 3'b000,
    parameter integer DATA_WIDTH_A = 18,
    parameter integer DATA_WIDTH_B = 18,
    parameter WRITE_MODE_A = "NORMAL_WRITE",
    parameter WRITE_MODE_B = "NORMAL_WRITE",
    parameter integer DOA_REG = 0,
    parameter integer DOB_REG = 0,
    parameter integer DOA_REG_CLKINV = 0,
    parameter integer DOB_REG_CLKINV = 0,
    parameter [35:0] RSTA_VAL = 36'b0,
    parameter [35:0] RSTB_VAL = 36'b0,
    parameter RST_TYPE = "SYNC",
    parameter RAM_MODE = "TRUE_DUAL_PORT",
    parameter RAM_CASCADE = "NONE",
    parameter ECC_WRITE_EN = "FALSE",
    parameter ECC_READ_EN = "FALSE",
    parameter [287:0] INIT_00 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_01 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_02 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_03 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_04 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_05 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_06 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_07 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_08 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_09 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_10 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_11 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_12 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_13 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_14 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_15 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_16 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_17 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_18 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_19 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_20 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_21 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_22 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_23 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_24 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_25 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_26 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_27 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_28 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_29 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_2A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_2B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_2C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_2D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_2E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_2F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_30 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_31 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_32 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_33 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_34 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_35 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_36 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_37 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_38 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_39 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_3A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_3B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_3C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_3D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_3E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_3F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_40 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_41 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_42 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_43 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_44 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_45 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_46 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_47 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_48 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_49 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_4A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_4B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_4C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_4D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_4E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_4F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_50 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_51 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_52 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_53 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_54 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_55 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_56 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_57 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_58 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_59 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_5A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_5B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_5C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_5D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_5E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_5F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_60 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_61 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_62 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_63 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_64 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_65 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_66 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_67 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_68 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_69 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_6A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_6B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_6C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_6D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_6E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_6F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_70 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_71 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_72 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_73 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_74 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_75 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_76 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_77 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_78 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_79 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_7A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_7B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_7C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_7D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_7E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_7F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_FILE = "NONE",
    parameter integer BLOCK_X = 0,
    parameter integer BLOCK_Y = 0,
    parameter integer RAM_DATA_WIDTH = 18,
    parameter integer RAM_ADDR_WIDTH = 11,
    parameter INIT_FORMAT = "BIN"
) (
    output [35:0] DOA,
    output [35:0] DOB,
    input  [35:0] DIA,
    input  [35:0] DIB,
    input  [15:0] ADDRA,
    input  [15:0] ADDRB,
    input  ADDRA_HOLD,
    input  ADDRB_HOLD,
    input  [2:0] CSA,
    input  [2:0] CSB,
    input  [7:0] BWEA,
    input  [3:0] BWEB,
    input  CLKA,
    input  CLKB,
    input  CEA,
    input  CEB,
    input  WEA,
    input  WEB,
    input  ORCEA,
    input  ORCEB,
    input  RSTA,
    input  RSTB,
    input  CINA,
    input  CINB,
    input  INJECT_SBITERR,
    input  INJECT_DBITERR,
    output ECC_SBITERR,
    output ECC_DBITERR,
    output [8:0] ECC_RDADDR,
    output [7:0] ECC_PARITY,
    output COUTA,
    output COUTB
);
// synthesis translate_off


    localparam  BLOCK_DEPTH = 2**(DATA_WIDTH_A == 1 ? 15 :      // block type 32k*1
                                  DATA_WIDTH_A == 2 ? 14 :      // block type 16k*2
                                  DATA_WIDTH_A == 4 ? 13 :      // block type 8k*4
                                  DATA_WIDTH_A <= 9 ? 12 :      // block type 4k*8 or 4k*9
                                  DATA_WIDTH_A <= 18 ? 11 :     // block type 1k*36 or 1k*32
                                  DATA_WIDTH_A <= 36 ? 10 : 9); // block type 512*72 or 512*64     block memory address width

    localparam  BLOCK_WIDTH =   DATA_WIDTH_A;             //block memory data width

    localparam MEM_SIZE = 36864;
    localparam width_a = (DATA_WIDTH_A == 72) ? 36 : (DATA_WIDTH_A == 64) ? 32 : DATA_WIDTH_A;
    localparam width_b = (DATA_WIDTH_B == 72) ? 36 : (DATA_WIDTH_B == 64) ? 32 : DATA_WIDTH_B;

    integer  cnt;
    reg [9-1:0] mem [MEM_SIZE/9-1:0];

    reg csa_reg = 1'b0, csb_reg = 1'b0;
    reg [15:0] ada_reg = 16'b0, adb_reg = 16'b0;
    reg [35:0] da_reg = 36'b0, db_reg = 36'b0;
    reg wea_reg = 1'b0, web_reg = 1'b0;
    reg [7:0] bea_reg;
    reg [3:0] beb_reg;
    wire write_en_a, write_en_b, read_en_a, read_en_b;
    reg [35:0] DIA_int,DIB_int;
    reg ecc_wren,ecc_rden;
    wire ecc_sbiterr_int,ecc_dbiterr_int;
    reg ecc_sbiterr,ecc_dbiterr,ecc_sbiterr_reg,ecc_dbiterr_reg;
    reg [8:0] ecc_rdaddr,ecc_rdaddr_reg;
    reg [35:0] a_out_ecc,b_out_ecc;

    wire [7:0] ecc_p_enc,ecc_p_dec,ecc_p_out;
    wire [63:0] ecc_d_dec;
    wire [63:0] ecc_d_in;
    wire [63:0] ecc_d_out;
    wire [71:0] d_out_ecc;
    reg  [71:0] ecc_corrected;
    reg  [7:0] ecc_p_reg;

    reg [35:0] a_out;
    reg [35:0] a_out_reg;
    reg [35:0] b_out;
    reg [35:0] b_out_reg;

    wire grs, rsta_grs, rstb_grs;
    wire rsta_grs_sync;
    wire rstb_grs_sync;
    wire rsta_grs_async;
    wire rstb_grs_async;
    
    reg [35:0] doa, doa_mux, doa_reg;
    reg [35:0] dob, dob_mux, dob_reg;

    reg [1:0] cas_en;
    wire cas_inta, cas_intb;
    reg  cas_sela=1'b1, cas_selb=1'b1;
    wire [35:0] a_out_mux;
    wire [35:0] b_out_mux;
    wire CLKA_for_or, CLKB_for_or;
    wire rsta_int, rstb_int;

    wire [35:0] rsta_val_int;
    wire [35:0] rstb_val_int;

// synthesis translate_off

    assign rsta_val_int = ((DATA_WIDTH_A == 16 | DATA_WIDTH_A == 32) & DATA_WIDTH_B !=64) ? {4'h0,RSTA_VAL[34:27],RSTA_VAL[25:18],RSTA_VAL[16:9],RSTA_VAL[7:0]}:RSTA_VAL;
    assign rstb_val_int =  (DATA_WIDTH_B == 16 | DATA_WIDTH_B == 32) ? {4'h0,RSTB_VAL[34:27],RSTB_VAL[25:18],RSTB_VAL[16:9],RSTB_VAL[7:0]}:RSTB_VAL;

    initial begin
        #1;
        a_out = rsta_val_int;
        a_out_reg = rsta_val_int;
        b_out = rstb_val_int;
        b_out_reg = rstb_val_int;
        doa = RSTA_VAL;
        dob = RSTB_VAL;
        doa_mux = RSTA_VAL;
        dob_mux = RSTB_VAL;
    end

   reg [RAM_DATA_WIDTH-1:0] ini_mem [2**RAM_ADDR_WIDTH-1:0];
   integer p;
   initial
   begin
      if(INIT_FILE != "NONE")
      begin
          if(INIT_FORMAT == "BIN")
              $readmemb(INIT_FILE,ini_mem);
          else
              $readmemh(INIT_FILE,ini_mem);
          for(p=0;p<20;p=p+1)
              $display("ini_mem[%d] = %b",p,ini_mem[p]);
      end
   end
///////////////////
// parameter check
///////////////////
    initial begin
        case (DATA_WIDTH_A)
            1, 2, 4, 8, 16, 32, 64: begin
                case (DATA_WIDTH_B)
                    1, 2, 4, 8, 16, 32, 64:  ; //null
                    default: begin
                        $display("ERROR: GTP_DRM36K_E1 instance %m parameter DATA_WIDTH_B:%d is illegal. The legal values are 1,2,4,8,16,32 or 64.",DATA_WIDTH_B);
                        $finish;
                    end
                endcase
            end
            9, 18, 36, 72: begin
                case (DATA_WIDTH_B)
                    9, 18, 36, 72:    ; //null
                    default: begin
                        $display("ERROR: GTP_DRM36K_E1 instance %m parameter DATA_WIDTH_B:%d is illegal. The legal values are 9,18,32 or 72.",DATA_WIDTH_B);
                        $finish;
                    end
                endcase
            end
            default: begin
                $display("ERROR: GTP_DRM36K_E1 instance %m parameter DATA_WIDTH_A:%d is illegal. The legal values are 1,2,4,8,9,16,18,32,36,64 or 72.",DATA_WIDTH_A);
                $finish;
            end
        endcase

        case (WRITE_MODE_A)
            "NORMAL_WRITE",
            "TRANSPARENT_WRITE",
            "READ_BEFORE_WRITE":    ; //null 
            default: begin
                $display("ERROR: GTP_DRM36K_E1 instance %m parameter WRITE_MODE_A: %s is illegal. The legal values are NORMAL_WRITE,TRANSPARENT_WRITE or READ_BEFORE_WRITE.", WRITE_MODE_A);
                $finish;
            end
        endcase

        case (WRITE_MODE_B)
            "NORMAL_WRITE",
            "TRANSPARENT_WRITE",
            "READ_BEFORE_WRITE":    ; //null  
            default: begin
                $display("ERROR: GTP_DRM36K_E1 instance %m parameter WRITE_MODE_B: %s is illegal. The legal values are NORMAL_WRITE,TRANSPARENT_WRITE or READ_BEFORE_WRITE.", WRITE_MODE_B);
                $finish;
            end
        endcase

        case (DOA_REG)
            0,1:     ;//null
            default: begin
                $display("ERROR: GTP_DRM36K_E1 instance %m parameter DOA_REG: %s is illegal. The legal values are 0 or 1.", DOA_REG);
                $finish;
            end
        endcase

        case (DOB_REG)
            0,1:     ;//null
            default: begin
                $display("ERROR: GTP_DRM36K_E1 instance %m parameter DOB_REG: %s is illegal. The legal values are 0 or 1.", DOB_REG);
                $finish;
            end
        endcase

        case (DOA_REG_CLKINV)
            0,1:     ;//null
            default: begin
                $display("ERROR: GTP_DRM36K_E1 instance %m parameter DOA_REG_CLKINV: %s is illegal. The legal values are 0 or 1.", DOA_REG_CLKINV);
                $finish;
            end
        endcase

        case (DOB_REG_CLKINV)
            0,1:     ;//null
            default: begin
                $display("ERROR: GTP_DRM36K_E1 instance %m parameter DOB_REG_CLKINV: %s is illegal. The legal values are 0 or 1.", DOB_REG_CLKINV);
                $finish;
            end
        endcase

        case (RST_TYPE)
            "ASYNC",
            "SYNC":     ;//null
            default: begin
                $display("ERROR: GTP_DRM36K_E1 instance %m parameter RST_TYPE: %s is illegal. The legal values are ASYNC or SYNC.", RST_TYPE);
                $finish;
            end
        endcase

        case (RAM_MODE)
            "ROM",
            "SINGLE_PORT":      ;//null
            "SIMPLE_DUAL_PORT": begin
                if (DATA_WIDTH_A <= 36 && WRITE_MODE_A != "NORMAL_WRITE") begin
                    $display("Warrning: GTP_DRM36K_E1 instance %m suggest to use TRUE_DUAL_PORT RAM_MODE if DATA_WIDTH_A and WRITE_MODE_A: %d,%s.",DATA_WIDTH_A,WRITE_MODE_A);
                end
            end
            "TRUE_DUAL_PORT": begin
                if (DATA_WIDTH_A > 36 || DATA_WIDTH_B > 36) begin
                    $display("ERROR: GTP_DRM36K_E1 instance %m parameter DATA_WIDTH_A and DATA_WIDTH_B in TRUE_DUAL_PORT MODE:%d,%d is illegal. The legal values are 1,2,4,8,9,16 or 18.",DATA_WIDTH_A,DATA_WIDTH_B);
                    $finish;
                end
            end
            default: begin
                $display("ERROR: GTP_DRM36K_E1 instance %m parameter RAM_MODE value: %s is illegal. The legal values are ROM or SINGLE_PORT, SIMPLE_DUAL_PORT or TRUE_DUAL_PORT.", RAM_MODE);
                $finish;
            end
        endcase
        
        case (RAM_CASCADE)
            "NONE": begin
                cas_en = 2'b00;
            end
            "LOWER": begin
                if (DATA_WIDTH_A != 1 || DATA_WIDTH_B != 1) begin
                    $display("ERROR: GTP_DRM36K_E1 instance %m parameter DATA_WIDTH_A and DATA_WIDTH_B:%s,%s in CASCADING MODE:%s are illegal, then DATA_WIDTH_A and DATA_WIDTH_B have to be set to 1.",DATA_WIDTH_A,DATA_WIDTH_B,RAM_CASCADE);
                    $finish;
                end
                cas_en = 2'b01;
            end
            "UPPER": begin
                if (DATA_WIDTH_A != 1 || DATA_WIDTH_B != 1) begin
                    $display("ERROR: GTP_DRM36K_E1 instance %m parameter DATA_WIDTH_A and DATA_WIDTH_B:%s,%s in CASCADING MODE:%s are illegal, then DATA_WIDTH_A and DATA_WIDTH_B have to be set to 1.",DATA_WIDTH_A,DATA_WIDTH_B,RAM_CASCADE);
                    $finish;
                end
                cas_en = 2'b11;
            end
            default: begin
                $display("ERROR: GTP_DRM36K_E1 instance %m parameter RAM_CASCADE: %s is illegal, the legal values are NONE,LOWER or UPPER", RAM_CASCADE);
                $finish;
            end
        endcase

        case (ECC_WRITE_EN)
            "FALSE": ecc_wren = 1'b0;
            "TRUE" : begin
                ecc_wren = 1'b1;
                if (DATA_WIDTH_A != 72 || DATA_WIDTH_B != 72) begin
                    $display("ERROR: ECCWR_ERROR GTP_DRM36K_E1 instance %m parameter DATA_WIDTH_A and DATA_WIDTH_B:%s,%s in ECC MODE:%s are illegal, then DATA_WIDTH_A and DATA_WIDTH_B have to be set to 72.",DATA_WIDTH_A,DATA_WIDTH_B,ECC_WRITE_EN);
                    $finish;
                end
            end
            default: begin
                    $display("ERROR: ECCWR_ERROR GTP_DRM36K_E1 instance %m parameter ECC_WRITE_EN:%s is illegal, the lecal values are TRUE or FALSE.",ECC_WRITE_EN);
                    $finish;
            end
        endcase

        case (ECC_READ_EN)
            "FALSE": ecc_rden = 1'b0;
            "TRUE" : begin
                ecc_rden = 1'b1;
                if (DATA_WIDTH_A != 72 || DATA_WIDTH_B != 72) begin
                    $display("ERROR: ECCRD_ERROR GTP_DRM36K_E1 instance %m parameter DATA_WIDTH_A and DATA_WIDTH_B:%s,%s in ECC MODE:%s are illegal, then DATA_WIDTH_A and DATA_WIDTH_B have to be set to 72.",DATA_WIDTH_A,DATA_WIDTH_B,ECC_READ_EN);
                    $finish;
                end
            end
            default: begin
                    $display("ERROR: ECCRD_ERROR GTP_DRM36K_E1 instance %m parameter ECC_READ_EN:%s is illegal, the lecal values are TRUE or FALSE.",ECC_READ_EN);
                    $finish;
            end
        endcase
    end

/////////////////
// initialization
/////////////////

    initial begin
        if (INIT_FILE == "NONE") begin
            for (cnt = 0; cnt < 32; cnt = cnt + 1) begin
                mem[32*0 + cnt] = INIT_00[cnt*9 +: 9];
                mem[32*1 + cnt] = INIT_01[cnt*9 +: 9];
                mem[32*2 + cnt] = INIT_02[cnt*9 +: 9];
                mem[32*3 + cnt] = INIT_03[cnt*9 +: 9];
                mem[32*4 + cnt] = INIT_04[cnt*9 +: 9];
                mem[32*5 + cnt] = INIT_05[cnt*9 +: 9];
                mem[32*6 + cnt] = INIT_06[cnt*9 +: 9];
                mem[32*7 + cnt] = INIT_07[cnt*9 +: 9];
                mem[32*8 + cnt] = INIT_08[cnt*9 +: 9];
                mem[32*9 + cnt] = INIT_09[cnt*9 +: 9];
                mem[32*10 + cnt] = INIT_0A[cnt*9 +: 9];
                mem[32*11 + cnt] = INIT_0B[cnt*9 +: 9];
                mem[32*12 + cnt] = INIT_0C[cnt*9 +: 9];
                mem[32*13 + cnt] = INIT_0D[cnt*9 +: 9];
                mem[32*14 + cnt] = INIT_0E[cnt*9 +: 9];
                mem[32*15 + cnt] = INIT_0F[cnt*9 +: 9];
                mem[32*16 + cnt] = INIT_10[cnt*9 +: 9];
                mem[32*17 + cnt] = INIT_11[cnt*9 +: 9];
                mem[32*18 + cnt] = INIT_12[cnt*9 +: 9];
                mem[32*19 + cnt] = INIT_13[cnt*9 +: 9];
                mem[32*20 + cnt] = INIT_14[cnt*9 +: 9];
                mem[32*21 + cnt] = INIT_15[cnt*9 +: 9];
                mem[32*22 + cnt] = INIT_16[cnt*9 +: 9];
                mem[32*23 + cnt] = INIT_17[cnt*9 +: 9];
                mem[32*24 + cnt] = INIT_18[cnt*9 +: 9];
                mem[32*25 + cnt] = INIT_19[cnt*9 +: 9];
                mem[32*26 + cnt] = INIT_1A[cnt*9 +: 9];
                mem[32*27 + cnt] = INIT_1B[cnt*9 +: 9];
                mem[32*28 + cnt] = INIT_1C[cnt*9 +: 9];
                mem[32*29 + cnt] = INIT_1D[cnt*9 +: 9];
                mem[32*30 + cnt] = INIT_1E[cnt*9 +: 9];
                mem[32*31 + cnt] = INIT_1F[cnt*9 +: 9];
                mem[32*32 + cnt] = INIT_20[cnt*9 +: 9];
                mem[32*33 + cnt] = INIT_21[cnt*9 +: 9];
                mem[32*34 + cnt] = INIT_22[cnt*9 +: 9];
                mem[32*35 + cnt] = INIT_23[cnt*9 +: 9];
                mem[32*36 + cnt] = INIT_24[cnt*9 +: 9];
                mem[32*37 + cnt] = INIT_25[cnt*9 +: 9];
                mem[32*38 + cnt] = INIT_26[cnt*9 +: 9];
                mem[32*39 + cnt] = INIT_27[cnt*9 +: 9];
                mem[32*40 + cnt] = INIT_28[cnt*9 +: 9];
                mem[32*41 + cnt] = INIT_29[cnt*9 +: 9];
                mem[32*42 + cnt] = INIT_2A[cnt*9 +: 9];
                mem[32*43 + cnt] = INIT_2B[cnt*9 +: 9];
                mem[32*44 + cnt] = INIT_2C[cnt*9 +: 9];
                mem[32*45 + cnt] = INIT_2D[cnt*9 +: 9];
                mem[32*46 + cnt] = INIT_2E[cnt*9 +: 9];
                mem[32*47 + cnt] = INIT_2F[cnt*9 +: 9];
                mem[32*48 + cnt] = INIT_30[cnt*9 +: 9];
                mem[32*49 + cnt] = INIT_31[cnt*9 +: 9];
                mem[32*50 + cnt] = INIT_32[cnt*9 +: 9];
                mem[32*51 + cnt] = INIT_33[cnt*9 +: 9];
                mem[32*52 + cnt] = INIT_34[cnt*9 +: 9];
                mem[32*53 + cnt] = INIT_35[cnt*9 +: 9];
                mem[32*54 + cnt] = INIT_36[cnt*9 +: 9];
                mem[32*55 + cnt] = INIT_37[cnt*9 +: 9];
                mem[32*56 + cnt] = INIT_38[cnt*9 +: 9];
                mem[32*57 + cnt] = INIT_39[cnt*9 +: 9];
                mem[32*58 + cnt] = INIT_3A[cnt*9 +: 9];
                mem[32*59 + cnt] = INIT_3B[cnt*9 +: 9];
                mem[32*60 + cnt] = INIT_3C[cnt*9 +: 9];
                mem[32*61 + cnt] = INIT_3D[cnt*9 +: 9];
                mem[32*62 + cnt] = INIT_3E[cnt*9 +: 9];
                mem[32*63 + cnt] = INIT_3F[cnt*9 +: 9];
                mem[32*64 + cnt] = INIT_40[cnt*9 +: 9];
                mem[32*65 + cnt] = INIT_41[cnt*9 +: 9];
                mem[32*66 + cnt] = INIT_42[cnt*9 +: 9];
                mem[32*67 + cnt] = INIT_43[cnt*9 +: 9];
                mem[32*68 + cnt] = INIT_44[cnt*9 +: 9];
                mem[32*69 + cnt] = INIT_45[cnt*9 +: 9];
                mem[32*70 + cnt] = INIT_46[cnt*9 +: 9];
                mem[32*71 + cnt] = INIT_47[cnt*9 +: 9];
                mem[32*72 + cnt] = INIT_48[cnt*9 +: 9];
                mem[32*73 + cnt] = INIT_49[cnt*9 +: 9];
                mem[32*74 + cnt] = INIT_4A[cnt*9 +: 9];
                mem[32*75 + cnt] = INIT_4B[cnt*9 +: 9];
                mem[32*76 + cnt] = INIT_4C[cnt*9 +: 9];
                mem[32*77 + cnt] = INIT_4D[cnt*9 +: 9];
                mem[32*78 + cnt] = INIT_4E[cnt*9 +: 9];
                mem[32*79 + cnt] = INIT_4F[cnt*9 +: 9];
                mem[32*80 + cnt] = INIT_50[cnt*9 +: 9];
                mem[32*81 + cnt] = INIT_51[cnt*9 +: 9];
                mem[32*82 + cnt] = INIT_52[cnt*9 +: 9];
                mem[32*83 + cnt] = INIT_53[cnt*9 +: 9];
                mem[32*84 + cnt] = INIT_54[cnt*9 +: 9];
                mem[32*85 + cnt] = INIT_55[cnt*9 +: 9];
                mem[32*86 + cnt] = INIT_56[cnt*9 +: 9];
                mem[32*87 + cnt] = INIT_57[cnt*9 +: 9];
                mem[32*88 + cnt] = INIT_58[cnt*9 +: 9];
                mem[32*89 + cnt] = INIT_59[cnt*9 +: 9];
                mem[32*90 + cnt] = INIT_5A[cnt*9 +: 9];
                mem[32*91 + cnt] = INIT_5B[cnt*9 +: 9];
                mem[32*92 + cnt] = INIT_5C[cnt*9 +: 9];
                mem[32*93 + cnt] = INIT_5D[cnt*9 +: 9];
                mem[32*94 + cnt] = INIT_5E[cnt*9 +: 9];
                mem[32*95 + cnt] = INIT_5F[cnt*9 +: 9];
                mem[32*96 + cnt] = INIT_60[cnt*9 +: 9];
                mem[32*97 + cnt] = INIT_61[cnt*9 +: 9];
                mem[32*98 + cnt] = INIT_62[cnt*9 +: 9];
                mem[32*99 + cnt] = INIT_63[cnt*9 +: 9];
                mem[32*100 + cnt] = INIT_64[cnt*9 +: 9];
                mem[32*101 + cnt] = INIT_65[cnt*9 +: 9];
                mem[32*102 + cnt] = INIT_66[cnt*9 +: 9];
                mem[32*103 + cnt] = INIT_67[cnt*9 +: 9];
                mem[32*104 + cnt] = INIT_68[cnt*9 +: 9];
                mem[32*105 + cnt] = INIT_69[cnt*9 +: 9];
                mem[32*106 + cnt] = INIT_6A[cnt*9 +: 9];
                mem[32*107 + cnt] = INIT_6B[cnt*9 +: 9];
                mem[32*108 + cnt] = INIT_6C[cnt*9 +: 9];
                mem[32*109 + cnt] = INIT_6D[cnt*9 +: 9];
                mem[32*110 + cnt] = INIT_6E[cnt*9 +: 9];
                mem[32*111 + cnt] = INIT_6F[cnt*9 +: 9];
                mem[32*112 + cnt] = INIT_70[cnt*9 +: 9];
                mem[32*113 + cnt] = INIT_71[cnt*9 +: 9];
                mem[32*114 + cnt] = INIT_72[cnt*9 +: 9];
                mem[32*115 + cnt] = INIT_73[cnt*9 +: 9];
                mem[32*116 + cnt] = INIT_74[cnt*9 +: 9];
                mem[32*117 + cnt] = INIT_75[cnt*9 +: 9];
                mem[32*118 + cnt] = INIT_76[cnt*9 +: 9];
                mem[32*119 + cnt] = INIT_77[cnt*9 +: 9];
                mem[32*120 + cnt] = INIT_78[cnt*9 +: 9];
                mem[32*121 + cnt] = INIT_79[cnt*9 +: 9];
                mem[32*122 + cnt] = INIT_7A[cnt*9 +: 9];
                mem[32*123 + cnt] = INIT_7B[cnt*9 +: 9];
                mem[32*124 + cnt] = INIT_7C[cnt*9 +: 9];
                mem[32*125 + cnt] = INIT_7D[cnt*9 +: 9];
                mem[32*126 + cnt] = INIT_7E[cnt*9 +: 9];
                mem[32*127 + cnt] = INIT_7F[cnt*9 +: 9];
            end
        end
        else  begin      // INIT_FILE 
            case(DATA_WIDTH_A)
                1: begin  //DRM TYPE 32K*1
                   for(cnt=0; cnt<4*1024;cnt = cnt+1)
                       mem[cnt][7:0] = {ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*8+7][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*8+6][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*8+5][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*8+4][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*8+3][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*8+2][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*8+1][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*8][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH]};
                end
                2: begin //DRM TYPE 16K*2
                   for(cnt=0; cnt<4*1024;cnt = cnt+1)
                       mem[cnt][7:0] = {ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*4+3][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*4+2][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*4+1][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*4][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH]};
                end
                4: begin //DRM TYPE 8K*4
                   for(cnt=0; cnt<4*1024;cnt = cnt+1)
                       {mem[cnt][7:0]} = {ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*2+1][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                          ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*2][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH]};
                end
                8: begin //DRM TYPE 4K*8
                   for(cnt=0; cnt<4*1024;cnt = cnt+1)
                       mem[cnt][7:0] = ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH];
                end
                9: begin //DRM TYPE 4K*9
                   for(cnt=0; cnt<4*1024;cnt = cnt+1)
                       mem[cnt] = ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH];
                end
                16:begin //DRM TYPE 2k*16
                   for(cnt=0; cnt<2*1024;cnt = cnt+1)
                       {mem[cnt*2+1][7:0], mem[cnt*2][7:0]} = ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH];
                end
                18:begin //DRM TYPE 2k*18
                   for(cnt=0; cnt<2*1024;cnt = cnt+1)
                       {mem[cnt*2+1], mem[cnt*2]} = ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH];
                end
                32:begin //DRM TYPE 1k*32
                   for(cnt=0; cnt<1024;cnt = cnt+1)
                       {mem[cnt*4+3][7:0],mem[cnt*4+2][7:0],mem[cnt*4+1][7:0],mem[cnt*4][7:0]} = ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH];
                end
                36:begin //DRM TYPE 1k*36
                   for(cnt=0; cnt<1024;cnt = cnt+1)
                       {mem[cnt*4+3],mem[cnt*4+2],mem[cnt*4+1],mem[cnt*4]} = ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH];
                end
                64:begin //DRM TYPE 512*64
                   for(cnt=0; cnt<512;cnt = cnt+1)
                       {mem[cnt*8+7][7:0],mem[cnt*8+6][7:0],mem[cnt*8+5][7:0],mem[cnt*8+4][7:0],
                        mem[cnt*8+3][7:0],mem[cnt*8+2][7:0],mem[cnt*8+1][7:0],mem[cnt*8][7:0]} = ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH];
                end
                72:begin //DRM TYPE 512*72
                   for(cnt=0; cnt<512;cnt = cnt+1)
                       {mem[cnt*8+7],mem[cnt*8+6],mem[cnt*8+5],mem[cnt*8+4],
                        mem[cnt*8+3],mem[cnt*8+2],mem[cnt*8+1],mem[cnt*8]} = ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH];
                end
            endcase
        end
    end

    always @(*) begin
        DIB_int = ecc_wren ? {ecc_p_enc[7],DIB[34:27],ecc_p_enc[6],DIB[25:18],ecc_p_enc[3],DIB[16:9],ecc_p_enc[2],DIB[7:0]} : DIB;
        DIA_int = ecc_wren ? {ecc_p_enc[5],DIA[34:27],ecc_p_enc[4],DIA[25:18],ecc_p_enc[1],DIA[16:9],ecc_p_enc[0],DIA[7:0]} : DIA;
        if(ecc_wren && (INJECT_SBITERR || INJECT_DBITERR)) begin
            DIB_int[15] = ~ DIB_int[15];
        end
        if(ecc_wren && INJECT_DBITERR) begin
            DIB_int[33] = ~ DIB_int[33];
        end
    end

    always @(posedge CLKA) begin
        if (CEA) begin
            // high to hold the address
            if (ADDRA_HOLD == 1'b0) begin
                if(CSA == CSA_MASK) begin
                    ada_reg <= ADDRA;
                end
                csa_reg <= (CSA == CSA_MASK);
            end
            da_reg <= DIA_int;
            wea_reg <= WEA;
            bea_reg <= BWEA;
            ecc_p_reg <= ecc_p_enc;
        end
    end

    always @(posedge CLKB) begin
        if (CEB) begin
            // high to hold the address
            if (ADDRB_HOLD == 1'b0) begin
                if(CSB == CSB_MASK) begin
                   adb_reg <= ADDRB;
                end
                csb_reg <= (CSB == CSB_MASK);
            end
          //db_reg <= DIB_int;
            web_reg <= WEB;
            beb_reg <= BWEB;
        end
    end

    ///////////////////
    // task & function
    ///////////////////

    function [DATA_WIDTH_A-1:0] mem_read_a;
        input [14:0]  addr;
    begin
        case (DATA_WIDTH_A)
            1: mem_read_a = mem[addr[14:3]][addr[2:0]];
            2: mem_read_a = mem[addr[14:3]][addr[2:1]*2 +: 2];
            4: mem_read_a = mem[addr[14:3]][addr[2]*4 +: 4];
            8: mem_read_a = mem[addr[14:3]][7:0];
            9: mem_read_a = mem[addr[14:3]];
            16: mem_read_a = {mem[addr[14:4]*2+1][7:0], mem[addr[14:4]*2][7:0]};
            18: mem_read_a = {mem[addr[14:4]*2+1]     , mem[addr[14:4]*2]};
            32: mem_read_a = {mem[addr[14:5]*4+3][7:0], mem[addr[14:5]*4+2][7:0], mem[addr[14:5]*4+1][7:0], mem[addr[14:5]*4][7:0]};
            36: mem_read_a = {mem[addr[14:5]*4+3]     , mem[addr[14:5]*4+2]     , mem[addr[14:5]*4+1]     , mem[addr[14:5]*4]};
            default:      ;//null 
        endcase
    end
    endfunction

    function [DATA_WIDTH_B-1:0] mem_read_b;
        input [14:0]  addr;
    begin
        case (DATA_WIDTH_B)
            1: mem_read_b = mem[addr[14:3]][addr[2:0]];
            2: mem_read_b = mem[addr[14:3]][addr[2:1]*2 +: 2];
            4: mem_read_b = mem[addr[14:3]][addr[2]*4 +: 4];
            8: mem_read_b = mem[addr[14:3]][7:0];
            9: mem_read_b = mem[addr[14:3]];
            16: mem_read_b = {mem[addr[14:4]*2+1][7:0], mem[addr[14:4]*2][7:0]};
            18: mem_read_b = {mem[addr[14:4]*2+1]     , mem[addr[14:4]*2]};
            32: mem_read_b = {mem[addr[14:5]*4+3][7:0], mem[addr[14:5]*4+2][7:0], mem[addr[14:5]*4+1][7:0], mem[addr[14:5]*4][7:0]};
            36: mem_read_b = {mem[addr[14:5]*4+3]     , mem[addr[14:5]*4+2]     , mem[addr[14:5]*4+1]     , mem[addr[14:5]*4]};
            64: mem_read_b = {mem[addr[14:6]*8+7][7:0], mem[addr[14:6]*8+6][7:0], mem[addr[14:6]*8+5][7:0], mem[addr[14:6]*8+4][7:0],
                              mem[addr[14:6]*8+3][7:0], mem[addr[14:6]*8+2][7:0], mem[addr[14:6]*8+1][7:0], mem[addr[14:6]*8][7:0]};
            72: mem_read_b = {mem[addr[14:6]*8+7], mem[addr[14:6]*8+6], mem[addr[14:6]*8+5], mem[addr[14:6]*8+4],
                              mem[addr[14:6]*8+3], mem[addr[14:6]*8+2], mem[addr[14:6]*8+1], mem[addr[14:6]*8]};
            default:      ;//null 
        endcase
    end
    endfunction

    task mem_write_a;
        input [14:0] addr;
        input [71:0] data;
        input [7:0]  byte_en;
    begin
        case (DATA_WIDTH_A)
            1: mem[addr[14:3]][addr[2:0]] = data[0];
            2: mem[addr[14:3]][addr[2:1]*2 +: 2] = data[1:0];
            4: mem[addr[14:3]][addr[2]*4 +: 4] = data[3:0];
            8: mem[addr[14:3]][7:0] = data[7:0];
            9: mem[addr[14:3]] = data[8:0];
            16: begin
                if (byte_en[1])
                    mem[addr[14:4]*2+1][7:0] = data[16:9];
                if (byte_en[0])
                    mem[addr[14:4]*2][7:0]   = data[7:0];
            end
            18: begin
                if (byte_en[1])
                    mem[addr[14:4]*2+1] = data[17:9];
                if (byte_en[0])
                    mem[addr[14:4]*2]   = data[8:0];
            end
            32: begin
                if (byte_en[3])
                    mem[addr[14:5]*4+3][7:0] = data[34:27];
                if (byte_en[2])
                    mem[addr[14:5]*4+2][7:0] = data[25:18];
                if (byte_en[1])
                    mem[addr[14:5]*4+1][7:0] = data[16:9];
                if (byte_en[0])
                    mem[addr[14:5]*4][7:0]   = data[7:0];
            end
            36: begin
                if (byte_en[3])
                    mem[addr[14:5]*4+3] = data[35:27];
                if (byte_en[2])
                    mem[addr[14:5]*4+2] = data[26:18];
                if (byte_en[1])
                    mem[addr[14:5]*4+1] = data[17:9];
                if (byte_en[0])
                    mem[addr[14:5]*4]   = data[8:0];
            end
            64: begin
                if (byte_en[7])
                    mem[addr[14:6]*8+7][7:0] = data[70:63];
                if (byte_en[6])
                    mem[addr[14:6]*8+6][7:0] = data[61:54];
                if (byte_en[5])
                    mem[addr[14:6]*8+5][7:0] = data[52:45];
                if (byte_en[4])
                    mem[addr[14:6]*8+4][7:0] = data[43:36];
                if (byte_en[3])
                    mem[addr[14:6]*8+3][7:0] = data[34:27];
                if (byte_en[2])
                    mem[addr[14:6]*8+2][7:0] = data[25:18];
                if (byte_en[1])
                    mem[addr[14:6]*8+1][7:0] = data[16:9];
                if (byte_en[0])
                    mem[addr[14:6]*8][7:0]   = data[7:0];
            end
            72: begin
                if (byte_en[7])
                    mem[addr[14:6]*8+7] = data[71:63];
                if (byte_en[6])
                    mem[addr[14:6]*8+6] = data[62:54];
                if (byte_en[5])
                    mem[addr[14:6]*8+5] = data[53:45];
                if (byte_en[4])
                    mem[addr[14:6]*8+4] = data[44:36];
                if (byte_en[3])
                    mem[addr[14:6]*8+3] = data[35:27];
                if (byte_en[2])
                    mem[addr[14:6]*8+2] = data[26:18];
                if (byte_en[1])
                    mem[addr[14:6]*8+1] = data[17:9];
                if (byte_en[0])
                    mem[addr[14:6]*8]   = data[8:0];
            end
            default:     ;//null
        endcase
    end
    endtask

    task mem_write_b;
        input [14:0] addr;
        input [35:0] data;
        input [3:0]  byte_en;
    begin
        case (DATA_WIDTH_B)
            1: mem[addr[14:3]][addr[2:0]] = data[0];
            2: mem[addr[14:3]][addr[2:1]*2 +: 2] = data[1:0];
            4: mem[addr[14:3]][addr[2]*4 +: 4] = data[3:0];
            8: mem[addr[14:3]][7:0] = data[7:0];
            9: mem[addr[14:3]] = data[8:0];
            16: begin
                if (byte_en[1])
                    mem[addr[14:4]*2+1][7:0] = data[16:9];
                if (byte_en[0])
                    mem[addr[14:4]*2][7:0]   = data[7:0];
            end
            18: begin
                if (byte_en[1])
                    mem[addr[14:4]*2+1] = data[17:9];
                if (byte_en[0])
                    mem[addr[14:4]*2]   = data[8:0];
            end
            32: begin
                if (byte_en[3])
                    mem[addr[14:5]*4+3][7:0] = data[34:27];
                if (byte_en[2])
                    mem[addr[14:5]*4+2][7:0] = data[25:18];
                if (byte_en[1])
                    mem[addr[14:5]*4+1][7:0] = data[16:9];
                if (byte_en[0])
                    mem[addr[14:5]*4][7:0]   = data[7:0];
            end
            36: begin
                if (byte_en[3])
                    mem[addr[14:5]*4+3] = data[35:27];
                if (byte_en[2])
                    mem[addr[14:5]*4+2] = data[26:18];
                if (byte_en[1])
                    mem[addr[14:5]*4+1] = data[17:9];
                if (byte_en[0])
                    mem[addr[14:5]*4]   = data[8:0];
            end
            default:     ;//null
        endcase
    end
    endtask

    function [7:0] func_ecc;
        input [63:0] ecc_din;
    begin
        func_ecc[0] = ecc_din[0]^ecc_din[1]^ecc_din[3]^ecc_din[4]^ecc_din[6]^ecc_din[8]
                         ^ecc_din[10]^ecc_din[11]^ecc_din[13]^ecc_din[15]^ecc_din[17]^ecc_din[19]
                         ^ecc_din[21]^ecc_din[23]^ecc_din[25]^ecc_din[26]^ecc_din[28]^ecc_din[30]
                         ^ecc_din[32]^ecc_din[34]^ecc_din[36]^ecc_din[38]^ecc_din[40]^ecc_din[42]
                         ^ecc_din[44]^ecc_din[46]^ecc_din[48]^ecc_din[50]^ecc_din[52]^ecc_din[54]
                         ^ecc_din[56]^ecc_din[57]^ecc_din[59]^ecc_din[61]^ecc_din[63];
        func_ecc[1] = ecc_din[0]^ecc_din[2]^ecc_din[3]^ecc_din[5]^ecc_din[6]^ecc_din[9]
                         ^ecc_din[10]^ecc_din[12]^ecc_din[13]^ecc_din[16]^ecc_din[17]^ecc_din[20]
                         ^ecc_din[21]^ecc_din[24]^ecc_din[25]^ecc_din[27]^ecc_din[28]^ecc_din[31]
                         ^ecc_din[32]^ecc_din[35]^ecc_din[36]^ecc_din[39]^ecc_din[40]^ecc_din[43]
                         ^ecc_din[44]^ecc_din[47]^ecc_din[48]^ecc_din[51]^ecc_din[52]^ecc_din[55]
                         ^ecc_din[56]^ecc_din[58]^ecc_din[59]^ecc_din[62]^ecc_din[63];
        func_ecc[2] = ecc_din[1]^ecc_din[2]^ecc_din[3]^ecc_din[7]^ecc_din[8]^ecc_din[9]
                         ^ecc_din[10]^ecc_din[14]^ecc_din[15]^ecc_din[16]^ecc_din[17]^ecc_din[22]
                         ^ecc_din[23]^ecc_din[24]^ecc_din[25]^ecc_din[29]^ecc_din[30]^ecc_din[31]
                         ^ecc_din[32]^ecc_din[37]^ecc_din[38]^ecc_din[39]^ecc_din[40]^ecc_din[45]
                         ^ecc_din[46]^ecc_din[47]^ecc_din[48]^ecc_din[53]^ecc_din[54]^ecc_din[55]
                         ^ecc_din[56]^ecc_din[60]^ecc_din[61]^ecc_din[62]^ecc_din[63];
        func_ecc[3] = ecc_din[4]^ecc_din[5]^ecc_din[6]^ecc_din[7]^ecc_din[8]^ecc_din[9]
                         ^ecc_din[10]^ecc_din[18]^ecc_din[19]^ecc_din[20]^ecc_din[21]^ecc_din[22]
                         ^ecc_din[23]^ecc_din[24]^ecc_din[25]^ecc_din[33]^ecc_din[34]^ecc_din[35]
                         ^ecc_din[36]^ecc_din[37]^ecc_din[38]^ecc_din[39]^ecc_din[40]^ecc_din[49]
                         ^ecc_din[50]^ecc_din[51]^ecc_din[52]^ecc_din[53]^ecc_din[54]^ecc_din[55]^ecc_din[56];
        func_ecc[4] = ecc_din[11]^ecc_din[12]^ecc_din[13]^ecc_din[14]^ecc_din[15]^ecc_din[16]
                         ^ecc_din[17]^ecc_din[18]^ecc_din[19]^ecc_din[20]^ecc_din[21]^ecc_din[22]
                         ^ecc_din[23]^ecc_din[24]^ecc_din[25]^ecc_din[41]^ecc_din[42]^ecc_din[43]
                         ^ecc_din[44]^ecc_din[45]^ecc_din[46]^ecc_din[47]^ecc_din[48]^ecc_din[49]
                         ^ecc_din[50]^ecc_din[51]^ecc_din[52]^ecc_din[53]^ecc_din[54]^ecc_din[55]^ecc_din[56];
        func_ecc[5] = ecc_din[26]^ecc_din[27]^ecc_din[28]^ecc_din[29]^ecc_din[30]^ecc_din[31]
                         ^ecc_din[32]^ecc_din[33]^ecc_din[34]^ecc_din[35]^ecc_din[36]^ecc_din[37]
                         ^ecc_din[38]^ecc_din[39]^ecc_din[40]^ecc_din[41]^ecc_din[42]^ecc_din[43]
                         ^ecc_din[44]^ecc_din[45]^ecc_din[46]^ecc_din[47]^ecc_din[48]^ecc_din[49]
                         ^ecc_din[50]^ecc_din[51]^ecc_din[52]^ecc_din[53]^ecc_din[54]^ecc_din[55]^ecc_din[56];
        func_ecc[6] = ecc_din[57]^ecc_din[58]^ecc_din[59]^ecc_din[60]^ecc_din[61]^ecc_din[62]^ecc_din[63];
        
        func_ecc[7] = ecc_din[0]^ecc_din[1]^ecc_din[2]^ecc_din[4]^ecc_din[5]^ecc_din[7]
                         ^ecc_din[10]^ecc_din[11]^ecc_din[12]^ecc_din[14]^ecc_din[17]^ecc_din[18]
                         ^ecc_din[21]^ecc_din[23]^ecc_din[24]^ecc_din[26]^ecc_din[27]^ecc_din[29]
                         ^ecc_din[32]^ecc_din[33]^ecc_din[36]^ecc_din[38]^ecc_din[39]^ecc_din[41]
                         ^ecc_din[44]^ecc_din[46]^ecc_din[47]^ecc_din[50]^ecc_din[51]^ecc_din[53]
                         ^ecc_din[56]^ecc_din[57]^ecc_din[58]^ecc_din[60]^ecc_din[63];
    end
    endfunction

    ///////////////
    // memory core
    ///////////////
reg CLKA_active;
reg CLKB_active;
initial begin
  CLKA_active = 1'b0;
  CLKB_active = 1'b0;
end
always @(posedge CLKA) begin
   if (CEA) begin
      CLKA_active <= 1'b1;
      #0.2 CLKA_active = 1'b0;
   end
   else
      CLKA_active <= 1'b0;
end
always @(posedge CLKB) begin
   if (CEB) begin
      CLKB_active <= 1'b1;
      #0.2 CLKB_active = 1'b0;
   end
   else
      CLKB_active <= 1'b0;
end

////////////////////////////////////////////////////////////////////////////////////////////
assign cas_inta = cas_en[1] ? ~ada_reg[15] : ada_reg[15];
assign cas_intb = cas_en[1] ? ~adb_reg[15] : adb_reg[15];

always @(*) begin
    if(WRITE_MODE_A == "NORMAL_WRITE" && wea_reg == 1'b1 || ~csa_reg) begin
        cas_sela = cas_sela;
    end else begin
        cas_sela = cas_inta;
    end
end
always @(*) begin
    if(WRITE_MODE_B == "NORMAL_WRITE" && web_reg == 1'b1 || ~csb_reg) begin
        cas_selb = cas_selb;
    end else begin
        cas_selb = cas_intb;
    end
end

assign a_out_mux[0] = ((cas_sela == 1'b0) && cas_en == 2'b11) ? CINA : a_out[0];
assign a_out_mux[35:1] = a_out[35:1];
assign b_out_mux[0] = ((cas_selb == 1'b0) && cas_en == 2'b11) ? CINB : b_out[0];
assign b_out_mux[35:1] = b_out[35:1];

assign COUTA = a_out[0];
assign COUTB = b_out[0];

generate
////////////////////////////////////////////////////////////////////////////////////////////
// ROM or SINGLE_PORT 
////////////////////////////////////////////////////////////////////////////////////////////
if(RAM_MODE == "ROM" || RAM_MODE == "SINGLE_PORT") begin:ROMorSP_MODE

    always @(posedge CLKA) begin
        if (CEA)
            db_reg <= DIB_int;
    end

    if (DATA_WIDTH_A > 36 || DATA_WIDTH_B > 36) begin

        assign write_en_a = csa_reg && cas_inta && (wea_reg == 1'b1);
        assign read_en_b  = csb_reg && cas_intb && (web_reg == 1'b0);
        // Port A (wirte) operations
        always @(negedge CLKA_active)
        begin
            if (write_en_a) begin  // write
              mem_write_a(ada_reg[14:0], {db_reg[35:0], da_reg[35:0]}, bea_reg);
            end
        end
        // Port B (read) operations
        always @(negedge CLKB_active or posedge rstb_int)
        begin
            if (rstb_int)
               {b_out, a_out} = {rstb_val_int, rsta_val_int};
            else if(read_en_b)begin
              if(DATA_WIDTH_B == 64)begin
                  {b_out[34:27],b_out[25:18],b_out[16:9],b_out[7:0],a_out[34:27],a_out[25:18],a_out[16:9],a_out[7:0]} = mem_read_b(adb_reg[14:0]);
              end
              else begin
                  {b_out[35:0],a_out[35:0]} = mem_read_b(adb_reg[14:0]);
              end
            end
        end

    end
    else  begin   //x1 x2 x4 x8 x9 x16 x18 x32 x36

        assign write_en_a = csa_reg && cas_inta && (wea_reg == 1'b1);
        assign read_en_a  = csa_reg && cas_inta && (wea_reg == 1'b0);
        // Port A operations
        always @(negedge CLKA_active)
        begin
            if (write_en_a)  begin  // write
               // read during write
               if (WRITE_MODE_A == "TRANSPARENT_WRITE") begin
                   a_out[width_a-1:0] = mem_read_a(ada_reg);

                   if(DATA_WIDTH_A == 16) begin
                       if(bea_reg[0])
                           a_out[7:0] = da_reg[7:0];
                       else
                           a_out[7:0] = a_out[7:0];

                       if(bea_reg[1])
                           a_out[15:8] = da_reg[16:9];
                       else
                           a_out[15:8] = a_out[15:8];
                   end
                   else if(DATA_WIDTH_A == 18) begin
                        if(bea_reg[0])
                            a_out[8:0] = da_reg[8:0];
                        else
                            a_out[8:0] = a_out[8:0];

                        if(bea_reg[1])
                            a_out[17:9] = da_reg[17:9];
                        else
                            a_out[17:9] = a_out[17:9];
                   end
                   else if(DATA_WIDTH_A == 32) begin
                       if(bea_reg[0])
                           a_out[7:0] = da_reg[7:0];
                       else
                           a_out[7:0] = a_out[7:0];

                       if(bea_reg[1])
                           a_out[15:8] = da_reg[16:9];
                       else
                           a_out[15:8] = a_out[15:8];

                       if(bea_reg[2])
                           a_out[23:16] = da_reg[25:18];
                       else
                           a_out[23:16] = a_out[23:16];

                       if(bea_reg[3])
                           a_out[31:24] = da_reg[34:27];
                       else
                           a_out[31:24] = a_out[31:24];
                   end
                   else if(DATA_WIDTH_A == 36) begin
                        if(bea_reg[0])
                            a_out[8:0] = da_reg[8:0];
                        else
                            a_out[8:0] = a_out[8:0];

                        if(bea_reg[1])
                            a_out[17:9] = da_reg[17:9];
                        else
                            a_out[17:9] = a_out[17:9];

                        if(bea_reg[2])
                            a_out[26:18] = da_reg[26:18];
                        else
                            a_out[26:18] = a_out[26:18];

                        if(bea_reg[3])
                            a_out[35:27] = da_reg[35:27];
                        else
                            a_out[35:27] = a_out[35:27];
                   end
                   else begin
                        a_out[width_a-1:0] = da_reg[width_a-1:0];
                   end
               end
               else if (WRITE_MODE_A == "READ_BEFORE_WRITE")
                   a_out[width_a-1:0] = mem_read_a(ada_reg[14:0]);

               mem_write_a(ada_reg[14:0], {36'b0, da_reg}, bea_reg);
            end
        end

        always @(negedge CLKA_active or posedge rsta_int)
        begin
            if (rsta_int)
               a_out = rsta_val_int;
            else if (read_en_a)          // read 
               a_out[width_a-1:0] = mem_read_a(ada_reg[14:0]);
        end
    end
end
////////////////////////////////////////////////////////////////////////////////////////////
//SIMPLE_DUAL_PORT
////////////////////////////////////////////////////////////////////////////////////////////
else if(RAM_MODE == "SIMPLE_DUAL_PORT")begin:SDP_MODE
    //port_A operation: only write in SDP MODE
    if (DATA_WIDTH_A > 36) begin:PORTA

        assign write_en_a = csa_reg && cas_inta && (wea_reg == 1'b1);

        always @(posedge CLKA) begin
           if (CEA)
              db_reg  <= DIB_int;
        end
        always @(negedge CLKA_active) begin
           if (write_en_a)    // write 
              mem_write_a(ada_reg[14:0], {db_reg[35:0], da_reg[35:0]}, bea_reg);
        end
    end
    else  begin:PORTA    //  x1 x2 x4 x8 x9 x16 x18 x32 x36

        assign write_en_a = csa_reg && cas_inta && (wea_reg == 1'b1);
        assign read_en_a  = csa_reg && cas_inta && (wea_reg == 1'b0) ;

        always @(negedge CLKA_active) begin
           if (write_en_a)     // write
           begin
              mem_write_a(ada_reg[14:0], {36'b0, da_reg}, bea_reg);
           end
        end
        if(DATA_WIDTH_B <= 36) begin
           always @(negedge CLKA_active or posedge rsta_int)
           begin
               if (rsta_int)
                  a_out = rsta_val_int;
               else if (read_en_a)
                  a_out[width_a-1 : 0] = mem_read_a(ada_reg[14:0]);
           end
        end
    end
    //port_B operation:only read in SDP MODE
    if (DATA_WIDTH_B > 36) begin:PORTB
    // SIMPLE_DUAL_PORT 
        assign read_en_b  = csb_reg && cas_intb && (web_reg == 1'b0);

        always @(negedge CLKB_active or posedge rstb_int)
        begin
           if (rstb_int)
              {b_out, a_out} = {rstb_val_int, rsta_val_int};
           else if (read_en_b)       // read 
                if(DATA_WIDTH_B == 64)begin
                  {b_out[34:27],b_out[25:18],b_out[16:9],b_out[7:0],a_out[34:27],a_out[25:18],a_out[16:9],a_out[7:0]} = mem_read_b(adb_reg[14:0]);
              end
              else begin
                  {b_out[35:0],a_out[35:0]} = mem_read_b(adb_reg[14:0]);
              end
        end
    end
    else  begin:PORTB  //  x1 x2 x4 x8 x9

        assign read_en_b  = csb_reg && cas_intb && (web_reg == 1'b0);

        always @(negedge CLKB_active or posedge rstb_int)
        begin
           if (rstb_int)
              b_out = rstb_val_int;
           else if (read_en_b)   //  read 
              b_out[width_b-1 : 0] = mem_read_b(adb_reg[14:0]);
        end
    end
end
////////////////////////////////////////////////////////////////////////////////////////////
//DP_MODE
////////////////////////////////////////////////////////////////////////////////////////////
else   begin:DP_MODE   //  --x1 x2 x4 x8 x9 x16 x18 x32 x36
    assign write_en_a = csa_reg && cas_inta && (wea_reg == 1'b1) ;
    assign read_en_a  = csa_reg && cas_inta && (wea_reg == 1'b0) ;
    assign write_en_b = csb_reg && cas_intb && (web_reg == 1'b1) ;
    assign read_en_b  = csb_reg && cas_intb && (web_reg == 1'b0) ;
    // Port A operations
    always @(negedge CLKA_active)
    begin
        if (write_en_a)  begin  // write
            // read during write
            if (WRITE_MODE_A == "TRANSPARENT_WRITE")
            begin
               a_out[width_a-1:0] = mem_read_a(ada_reg);

               if(DATA_WIDTH_A == 16) begin
                   if(bea_reg[0])
                       a_out[7:0] = da_reg[7:0];
                   else
                       a_out[7:0] = a_out[7:0];

                   if(bea_reg[1])
                       a_out[15:8] = da_reg[16:9];
                   else
                       a_out[15:8] = a_out[15:8];
               end
               else if(DATA_WIDTH_A == 18) begin
                    if(bea_reg[0])
                        a_out[8:0] = da_reg[8:0];
                    else
                        a_out[8:0] = a_out[8:0];

                    if(bea_reg[1])
                        a_out[17:9] = da_reg[17:9];
                    else
                        a_out[17:9] = a_out[17:9];
               end
               else if(DATA_WIDTH_A == 32) begin
                   if(bea_reg[0])
                       a_out[7:0] = da_reg[7:0];
                   else
                       a_out[7:0] = a_out[7:0];

                   if(bea_reg[1])
                       a_out[15:8] = da_reg[16:9];
                   else
                       a_out[15:8] = a_out[15:8];

                   if(bea_reg[2])
                       a_out[23:16] = da_reg[25:18];
                   else
                       a_out[23:16] = a_out[23:16];

                   if(bea_reg[3])
                       a_out[31:24] = da_reg[34:27];
                   else
                       a_out[31:24] = a_out[31:24];
               end
               else if(DATA_WIDTH_A == 36) begin
                    if(bea_reg[0])
                        a_out[8:0] = da_reg[8:0];
                    else
                        a_out[8:0] = a_out[8:0];

                    if(bea_reg[1])
                        a_out[17:9] = da_reg[17:9];
                    else
                        a_out[17:9] = a_out[17:9];

                    if(bea_reg[2])
                        a_out[26:18] = da_reg[26:18];
                    else
                        a_out[26:18] = a_out[26:18];

                    if(bea_reg[3])
                        a_out[35:27] = da_reg[35:27];
                    else
                        a_out[35:27] = a_out[35:27];
               end
               else begin
                    a_out[width_a-1:0] = da_reg[width_a-1:0];
               end
            end
            else if (WRITE_MODE_A == "READ_BEFORE_WRITE")
               a_out[width_a-1:0] = mem_read_a(ada_reg[14:0]);

            mem_write_a(ada_reg[14:0], {36'b0, da_reg}, bea_reg);
        end
    end

    always @(negedge CLKA_active or posedge rsta_int)
    begin
        if (rsta_int)
           a_out = rsta_val_int;
        else if (read_en_a)
           a_out[width_a-1 : 0] = mem_read_a(ada_reg[14:0]);
    end
    // Port B operations
    always @(posedge CLKB) begin
         if (CEB)
            db_reg <= DIB_int;
    end

    always @(negedge CLKB_active)
    begin
        if (write_en_b)  begin  // write
            // read during write
            if (WRITE_MODE_B == "TRANSPARENT_WRITE")
            begin
                b_out[width_b-1:0] = mem_read_b(adb_reg);

                if(DATA_WIDTH_B == 16) begin
                    if(beb_reg[0])
                        b_out[7:0] = db_reg[7:0];
                    else
                        b_out[7:0] = b_out[7:0];

                    if(beb_reg[1])
                        b_out[15:8] = db_reg[16:9];
                    else
                        b_out[15:8] = b_out[15:8];
                end
                else if(DATA_WIDTH_B == 18) begin
                    if(beb_reg[0])
                        b_out[8:0] = db_reg[8:0];
                    else
                        b_out[8:0] = b_out[8:0];

                    if(beb_reg[1])
                        b_out[17:9] = db_reg[17:9];
                    else
                        b_out[17:9] = b_out[17:9];
                end
                else if(DATA_WIDTH_B == 32) begin
                    if(beb_reg[0])
                        b_out[7:0] = db_reg[7:0];
                    else
                        b_out[7:0] = b_out[7:0];

                    if(beb_reg[1])
                        b_out[15:8] = db_reg[16:9];
                    else
                        b_out[15:8] = b_out[15:8];

                    if(beb_reg[2])
                        b_out[23:16] = db_reg[25:18];
                    else
                        b_out[23:16] = b_out[23:16];

                    if(beb_reg[3])
                        b_out[31:24] = db_reg[34:27];
                    else
                        b_out[31:24] = b_out[31:24];
                end
                else if(DATA_WIDTH_B == 36) begin
                     if(beb_reg[0])
                         b_out[8:0] = db_reg[8:0];
                     else
                         b_out[8:0] = b_out[8:0];

                     if(beb_reg[1])
                         b_out[17:9] = db_reg[17:9];
                     else
                         b_out[17:9] = b_out[17:9];

                     if(beb_reg[2])
                         b_out[26:18] = db_reg[26:18];
                     else
                         b_out[26:18] = b_out[26:18];

                     if(beb_reg[3])
                         b_out[35:27] = db_reg[35:27];
                     else
                         b_out[35:27] = b_out[35:27];
                end
                else begin
                    b_out[width_b-1:0] = db_reg[width_b-1:0];
                end
            end
            else if (WRITE_MODE_B == "READ_BEFORE_WRITE")
                b_out[width_b-1:0] = mem_read_b(adb_reg[14:0]);

            mem_write_b(adb_reg[14:0], db_reg, beb_reg);
        end
    end

    always @(negedge CLKB_active or posedge rstb_int)
    begin
        if (rstb_int)
           b_out = rstb_val_int;
        else if (read_en_b)
           b_out[width_b-1 : 0] = mem_read_b(adb_reg[14:0]);
    end
end
////////////////////////////////////////////////////////////////////////////////////////////
endgenerate


//////////////
// core latch
//////////////
assign grsn =  (GRS_EN == "TRUE") ? GRS_INST.GRSNET : 1'b1;
assign grs =  ~grsn;
or (rsta_grs, grs, RSTA);
or (rstb_grs, grs, RSTB);

reg rsta_grsn_d;

    always @(posedge CLKA_for_or) begin
        if (RSTA) begin
            rsta_grsn_d   <= 1'b1;
        end
        else begin
            rsta_grsn_d   <= 1'b0;
        end
    end

reg rstb_grsn_d;
    
    always @(posedge CLKB_for_or) begin
        if (RSTB) begin
            rstb_grsn_d   <= 1'b1;
        end
        else begin
            rstb_grsn_d   <= 1'b0;
        end
    end

initial begin
    rsta_grsn_d = 1'b1;
    rstb_grsn_d = 1'b1;
end

assign rsta_grs_sync  = (RST_TYPE == "SYNC") ? rsta_grsn_d : 1'b0;
assign rstb_grs_sync  = (RST_TYPE == "SYNC") ? rstb_grsn_d : 1'b0;
assign rsta_grs_async = (RST_TYPE == "ASYNC") ? rsta_grs : grs;
assign rstb_grs_async = (RST_TYPE == "ASYNC") ? rstb_grs : grs;

assign rsta_int = rsta_grs_sync | rsta_grs_async;
assign rstb_int = rstb_grs_sync | rstb_grs_async;
/////////////////////////////////////////////////////////////////////
//port out
assign CLKA_for_or = (DOA_REG_CLKINV == 1) ? ~CLKA : CLKA;
assign CLKB_for_or = (DOB_REG_CLKINV == 1) ? ~CLKB : CLKB;


generate
////////////////////////////////////////////////////////////////////////////////////////////
assign ecc_d_in  = {DIB[34:27],DIB[25:18],DIB[16:9],DIB[7:0],DIA[34:27],DIA[25:18],DIA[16:9],DIA[7:0]};
assign ecc_p_enc = func_ecc (ecc_d_in);
assign ecc_d_dec = {b_out_mux[34:27],b_out_mux[25:18],b_out_mux[16:9],b_out_mux[7:0],a_out_mux[34:27],a_out_mux[25:18],a_out_mux[16:9],a_out_mux[7:0]};
assign ecc_p_out = {b_out_mux[35],b_out_mux[26],b_out_mux[17],b_out_mux[8],a_out_mux[35],a_out_mux[26],a_out_mux[17],a_out_mux[8]};
assign ecc_d_out = {b_out_mux[34:27],b_out_mux[25:18],b_out_mux[16:9],b_out_mux[7:0],a_out_mux[34:27],a_out_mux[25:18],a_out_mux[16:9],a_out_mux[7:0]};
assign ecc_p_dec = func_ecc (ecc_d_out) ^ ecc_p_out;

assign ecc_sbiterr_int = ^ecc_p_dec;
assign ecc_dbiterr_int = (|ecc_p_dec[6:0]) & ~ecc_sbiterr_int;
always @(*) begin
    ecc_corrected = {ecc_d_dec[63:57], ecc_p_out[6], ecc_d_dec[56:26], ecc_p_out[5], ecc_d_dec[25:11], ecc_p_out[4], ecc_d_dec[10:4], ecc_p_out[3], ecc_d_dec[3:1], ecc_p_out[2], ecc_d_dec[0], ecc_p_out[1:0], ecc_p_out[7]};
    ecc_corrected[ecc_p_dec[6:0]] = ecc_sbiterr_int ^ecc_corrected[ecc_p_dec[6:0]];
end
assign d_out_ecc = {ecc_corrected[0],ecc_corrected[71:65],ecc_corrected[63],ecc_corrected[64],ecc_corrected[62:55],ecc_corrected[32],ecc_corrected[54:47],ecc_corrected[16],ecc_corrected[46:39],ecc_corrected[8],ecc_corrected[38:33],ecc_corrected[31:30],ecc_corrected[4],ecc_corrected[29:22],ecc_corrected[2],ecc_corrected[21:17],ecc_corrected[15:13],ecc_corrected[1],ecc_corrected[12:9],ecc_corrected[7:5],ecc_corrected[3]};
////////////////////////////////////////////////////////////////////////////////////////////
if (DATA_WIDTH_B > 36)
begin:FAKE_DP_OUT
    //port_A output
    always @(posedge CLKB_for_or or posedge rstb_int)
    begin
        if (rstb_int) begin
            a_out_reg <= RSTA_VAL;
        end else if (ORCEB) begin
            a_out_reg <= ecc_rden ? d_out_ecc[35:0] : a_out;
        end
    end

    //doa combination logic
    always @(*)
    begin
        if (DOB_REG == 0)
        begin
            case(DATA_WIDTH_B)
                64: doa_mux = a_out_mux;
                72: doa_mux = ecc_rden ? d_out_ecc[35:0] : a_out_mux;
            endcase
        end
        else
        begin
            case(DATA_WIDTH_B)
                64: doa_mux = a_out_reg;
                72: doa_mux = a_out_reg;
            endcase
        end
    end

    always @(posedge CLKB_for_or or posedge rstb_int)
    begin
        if (rstb_int) begin
            b_out_reg <= RSTB_VAL;
            ecc_sbiterr_reg <= 1'b0;
            ecc_dbiterr_reg <= 1'b0;
            ecc_rdaddr_reg <= 9'h0;
        end else if (ORCEB) begin
            b_out_reg <= ecc_rden ? d_out_ecc[71:36] : b_out;
            ecc_sbiterr_reg <= ecc_sbiterr_int;
            ecc_dbiterr_reg <= ecc_dbiterr_int;
            ecc_rdaddr_reg <= adb_reg[14:6];
        end
    end

    //dob combination logic
    always @(*)
    begin
        if (DOB_REG == 0)
        begin
            case(DATA_WIDTH_B)
                64: dob_mux = b_out_mux;
                72: dob_mux = ecc_rden ? d_out_ecc[71:36] : b_out_mux;
            endcase
            ecc_sbiterr = ecc_sbiterr_int;
            ecc_dbiterr = ecc_dbiterr_int;
            ecc_rdaddr = adb_reg[14:6];
        end
        else
        begin
            case(DATA_WIDTH_B)
                64: dob_mux = b_out_reg;
                72: dob_mux = b_out_reg;
            endcase
            ecc_sbiterr = ecc_sbiterr_reg;
            ecc_dbiterr = ecc_dbiterr_reg;
            ecc_rdaddr = ecc_rdaddr_reg;
        end
    end
end
////////////////////////////////////////////////////////////////////////////////////////////
else
begin:TRUE_DP_OUT
    //port_A output

    always @(posedge CLKA_for_or or posedge rsta_int)
    begin
        if (rsta_int)
            doa_reg <= RSTA_VAL;
        else if (ORCEA)
            doa_reg <= doa;
    end

    //doa combination logic
    always @(a_out_mux)
    begin
       case(DATA_WIDTH_A)
          1: {doa[16:9],doa[7:0]} = {16{a_out_mux[width_a-1:0]}};
          2: {doa[16:9],doa[7:0]} = { 8{a_out_mux[width_a-1:0]}};
          4: {doa[16:9],doa[7:0]} = { 4{a_out_mux[width_a-1:0]}};
          8: {doa[16:9],doa[7:0]} = { 2{a_out_mux[width_a-1:0]}};
          9: {doa[17:9],doa[8:0]} = { 2{a_out_mux[width_a-1:0]}};
          16:{doa[16:9],doa[7:0]} =     a_out_mux[width_a-1:0]  ;
          18: doa[17:0]           =     a_out_mux[width_a-1:0]  ;
          32:{doa[34:27],doa[25:18],doa[16:9],doa[7:0]} = a_out_mux[width_a-1:0]  ;
          36: doa = a_out_mux;
       endcase
    end

    always @(doa or doa_reg)
    begin
        if (DOA_REG == 0)
            doa_mux = doa;
        else
            doa_mux = doa_reg;
    end

    //port_B output

    always @(posedge CLKB_for_or or posedge rstb_int)
    begin
        if (rstb_int)
            dob_reg <= RSTB_VAL;
        else if (ORCEB)
            dob_reg <= dob;
    end

    //dob combination logic
    always @(b_out_mux)
    begin
        case(DATA_WIDTH_B)  
           1: {dob[16:9],dob[7:0]} = {16{b_out_mux[width_b-1:0]}};
           2: {dob[16:9],dob[7:0]} = { 8{b_out_mux[width_b-1:0]}};
           4: {dob[16:9],dob[7:0]} = { 4{b_out_mux[width_b-1:0]}};
           8: {dob[16:9],dob[7:0]} = { 2{b_out_mux[width_b-1:0]}};
           9: {dob[17:9],dob[8:0]} = { 2{b_out_mux[width_b-1:0]}};
           16:{dob[16:9],dob[7:0]} =     b_out_mux[width_b-1:0]  ;
           18: dob[17:0]           =     b_out_mux[width_b-1:0]  ;
           32:{dob[34:27],dob[25:18],dob[16:9],dob[7:0]} = b_out_mux[width_b-1:0]  ;
           36: dob = b_out_mux;
        endcase
    end

    always @(dob or dob_reg)
    begin
        if (DOB_REG == 0)
            dob_mux = dob;
        else
            dob_mux = dob_reg;
    end

end
////////////////////////////////////////////////////////////////////////////////////////////
endgenerate

assign DOA = doa_mux;
assign DOB = dob_mux;
assign ECC_PARITY = ecc_p_reg;
assign ECC_RDADDR = ecc_rdaddr;
assign ECC_SBITERR = ecc_sbiterr;
assign ECC_DBITERR = ecc_dbiterr;
// synthesis translate_on
endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_ONE.v
//
// Functional description: constant one
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_ONE
(
    output wire Z
);

    supply1 VSS;
    buf (Z, VSS);

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_RAM144K.v
//
// Functional description: (true) Dual-Port 144K-bit RAM block
//
// Parameter description:
//      DATA_WIDTH_A : data width of input/output of Port A
//      DATA_WIDTH_B : data width of input/output of Port B
//      RST_TYPE     : async or sync clear of Port A/B outputs
//      DOA_REG      : disable or enable output register of Port A
//      DOB_REG      : disable or enable output register of Port B
//      WRITE_MODE_A : read during write mode of Port A
//      WRITE_MODE_B : read during write mode of Port B
//      INIT_FILE  : RAM content initialization
//
// Port description:
//      CLKA : clock of Port A
//      CEA  : clock enable of Port A
//      WEA  : write enable of Port A
//      BEA  : byte write enable of Port A
//      ADDRA: address of Port A
//      DIA  : write data in of Port A
//      ORCEA: output register clock enable of Port A
//      RSTA : output async/sync clear of Port A
//      DOA  : read data out of Port A
//
// Revision:
//      2018/01/09: Update display informations.
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_RAM144K
#(
    parameter GRS_EN = "TRUE",
    parameter integer DATA_WIDTH_A = 18,
    parameter integer DATA_WIDTH_B = 18,
    parameter integer DOA_REG = 0,
    parameter integer DOB_REG = 0,
    parameter RST_TYPE = "SYNC",
    parameter WRITE_MODE_A = "NORMAL_WRITE",
    parameter WRITE_MODE_B = "NORMAL_WRITE",
    parameter WRITE_COLLISION_ARBITER = "NULL",
    parameter integer DRM18K_NUMBER = 8,
    parameter INIT_000 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_001 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_002 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_003 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_004 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_005 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_006 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_007 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_008 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_009 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_00A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_00B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_00C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_00D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_00E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_00F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_010 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_011 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_012 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_013 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_014 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_015 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_016 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_017 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_018 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_019 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_01A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_01B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_01C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_01D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_01E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_01F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_020 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_021 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_022 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_023 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_024 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_025 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_026 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_027 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_028 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_029 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_02A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_02B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_02C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_02D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_02E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_02F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_030 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_031 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_032 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_033 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_034 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_035 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_036 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_037 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_038 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_039 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_03A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_03B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_03C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_03D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_03E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_03F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_040 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_041 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_042 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_043 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_044 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_045 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_046 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_047 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_048 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_049 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_04A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_04B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_04C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_04D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_04E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_04F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_050 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_051 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_052 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_053 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_054 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_055 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_056 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_057 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_058 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_059 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_05A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_05B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_05C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_05D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_05E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_05F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_060 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_061 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_062 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_063 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_064 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_065 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_066 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_067 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_068 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_069 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_06A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_06B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_06C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_06D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_06E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_06F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_070 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_071 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_072 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_073 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_074 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_075 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_076 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_077 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_078 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_079 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_07A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_07B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_07C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_07D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_07E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_07F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_080 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_081 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_082 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_083 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_084 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_085 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_086 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_087 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_088 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_089 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_08A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_08B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_08C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_08D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_08E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_08F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_090 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_091 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_092 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_093 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_094 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_095 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_096 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_097 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_098 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_099 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_09A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_09B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_09C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_09D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_09E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_09F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0A0 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0A1 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0A2 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0A3 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0A4 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0A5 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0A6 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0A7 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0A8 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0A9 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0AA = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0AB = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0AC = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0AD = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0AE = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0AF = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0B0 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0B1 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0B2 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0B3 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0B4 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0B5 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0B6 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0B7 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0B8 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0B9 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0BA = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0BB = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0BC = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0BD = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0BE = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0BF = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0C0 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0C1 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0C2 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0C3 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0C4 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0C5 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0C6 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0C7 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0C8 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0C9 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0CA = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0CB = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0CC = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0CD = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0CE = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0CF = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0D0 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0D1 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0D2 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0D3 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0D4 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0D5 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0D6 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0D7 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0D8 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0D9 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0DA = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0DB = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0DC = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0DD = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0DE = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0DF = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0E0 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0E1 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0E2 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0E3 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0E4 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0E5 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0E6 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0E7 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0E8 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0E9 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0EA = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0EB = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0EC = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0ED = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0EE = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0EF = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0F0 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0F1 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0F2 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0F3 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0F4 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0F5 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0F6 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0F7 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0F8 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0F9 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0FA = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0FB = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0FC = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0FD = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0FE = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0FF = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_100 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_101 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_102 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_103 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_104 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_105 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_106 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_107 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_108 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_109 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_10A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_10B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_10C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_10D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_10E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_10F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_110 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_111 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_112 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_113 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_114 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_115 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_116 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_117 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_118 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_119 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_11A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_11B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_11C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_11D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_11E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_11F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_120 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_121 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_122 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_123 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_124 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_125 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_126 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_127 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_128 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_129 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_12A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_12B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_12C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_12D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_12E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_12F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_130 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_131 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_132 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_133 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_134 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_135 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_136 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_137 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_138 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_139 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_13A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_13B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_13C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_13D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_13E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_13F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_140 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_141 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_142 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_143 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_144 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_145 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_146 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_147 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_148 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_149 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_14A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_14B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_14C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_14D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_14E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_14F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_150 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_151 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_152 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_153 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_154 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_155 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_156 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_157 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_158 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_159 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_15A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_15B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_15C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_15D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_15E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_15F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_160 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_161 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_162 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_163 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_164 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_165 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_166 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_167 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_168 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_169 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_16A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_16B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_16C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_16D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_16E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_16F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_170 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_171 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_172 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_173 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_174 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_175 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_176 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_177 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_178 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_179 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_17A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_17B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_17C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_17D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_17E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_17F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_180 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_181 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_182 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_183 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_184 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_185 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_186 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_187 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_188 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_189 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_18A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_18B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_18C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_18D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_18E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_18F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_190 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_191 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_192 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_193 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_194 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_195 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_196 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_197 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_198 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_199 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_19A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_19B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_19C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_19D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_19E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_19F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1A0 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1A1 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1A2 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1A3 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1A4 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1A5 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1A6 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1A7 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1A8 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1A9 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1AA = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1AB = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1AC = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1AD = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1AE = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1AF = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1B0 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1B1 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1B2 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1B3 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1B4 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1B5 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1B6 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1B7 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1B8 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1B9 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1BA = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1BB = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1BC = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1BD = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1BE = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1BF = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1C0 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1C1 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1C2 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1C3 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1C4 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1C5 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1C6 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1C7 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1C8 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1C9 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1CA = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1CB = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1CC = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1CD = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1CE = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1CF = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1D0 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1D1 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1D2 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1D3 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1D4 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1D5 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1D6 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1D7 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1D8 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1D9 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1DA = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1DB = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1DC = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1DD = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1DE = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1DF = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1E0 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1E1 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1E2 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1E3 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1E4 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1E5 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1E6 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1E7 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1E8 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1E9 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1EA = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1EB = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1EC = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1ED = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1EE = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1EF = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1F0 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1F1 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1F2 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1F3 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1F4 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1F5 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1F6 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1F7 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1F8 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1F9 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1FA = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1FB = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1FC = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1FD = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1FE = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1FF = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_FILE = "NONE"
) (
    output [17:0] DOA,
    output [17:0] DOB,
    input [17:0] DIA,
    input [17:0] DIB,
    input [16:0] ADDRA,
    input [16:0] ADDRB,
    input CLKA,
    input CLKB,
    input CEA,
    input CEB,
    input WEA,
    input WEB,
    input [1:0] BEA,
    input [1:0] BEB,
    input ORCEA,
    input ORCEB,
    input RSTA,
    input RSTB

);

    wire [17:0] dangle_a18, dangle_b18;

    //
    // parameter check
    //

    initial begin
        case (DATA_WIDTH_A)
            1, 2, 4, 8, 16, 9, 18: begin
                case (DATA_WIDTH_B)
                    1, 2, 4, 8, 16, 9, 18:    ; // null  
                    default: begin
                        $display("ERROR: GTP_RAM144K instance %m parameter DATA_WIDTH_B:%d is illegal. The legal values are 1,2,4,8,16,9 or 18.",DATA_WIDTH_B);
                        $finish;
                    end
                endcase
            end
            default: begin
                $display("ERROR: GTP_RAM144K instance %m parameter DATA_WIDTH_A:%d is illegal. The legal values are 1,2,4,8,16,9 or 18.",DATA_WIDTH_A);
                $finish;
            end
        endcase

        if (RST_TYPE != "ASYNC" && RST_TYPE != "SYNC") begin
            $display("ERROR: GTP_RAM144K instance %m parameter:%s is illegal. The legal values are ASYNC or SYNC.",RST_TYPE);
            $finish;
        end

        if (DOA_REG != 0 && DOA_REG != 1) begin
            $display("ERROR: GTP_RAM144K instance %m parameter: DOA_REG:%d is illegal. The legal values are 0 or 1 .",DOA_REG);
            $finish;
        end

        if (DOB_REG != 0 && DOB_REG != 1) begin
            $display("ERROR: GTP_RAM144K instance %m parameter DOB_REG:%d is illegal. The legal values are 0 or 1 .",DOB_REG);
            $finish;
        end

        case (WRITE_MODE_A)
            "NORMAL_WRITE",
            "TRANSPARENT_WRITE",
            "READ_BEFORE_WRITE":    ;// null
            default: begin
                $display("ERROR: GTP_RAM144K instance %m parameter WRITE_MODE_A:%s is illegal. The legal values are NORMAL_WRITE ,TRANSPARENT_WRITE or READ_BEFORE_WRITE .",WRITE_MODE_A);
                $finish;
            end
        endcase

        case (WRITE_MODE_B)
            "NORMAL_WRITE",
            "TRANSPARENT_WRITE",
            "READ_BEFORE_WRITE":    ;// null
            default: begin
                $display("ERROR: GTP_RAM144K instance %m parameter WRITE_MODE_B:%s is illegal. The legal values are NORMAL_WRITE ,TRANSPARENT_WRITE or READ_BEFORE_WRITE .",WRITE_MODE_B);
                $finish;
            end
        endcase

        case (WRITE_COLLISION_ARBITER)
            "NULL": ;
            //"PORTA",
            //"PORTB":     ;// null
            default: begin
                $display("ERROR: GTP_RAM144K instance %m parameter:%s is illegal. The legal values is NULL .",WRITE_COLLISION_ARBITER);
                $finish;
            end
        endcase
    end

    INT_RAM144K
    #(
        .GRS_EN(GRS_EN),
        .DATA_WIDTH_A(DATA_WIDTH_A),
        .DATA_WIDTH_B(DATA_WIDTH_B),
        .CLEAR_TYPE(RST_TYPE),
        .OUTPUT_REG_A(DOA_REG),
        .OUTPUT_REG_B(DOB_REG),
        .WRITE_MODE_A(WRITE_MODE_A),
        .WRITE_MODE_B(WRITE_MODE_B),
        .WRITE_COLLISION_ARBITER(WRITE_COLLISION_ARBITER),
        .INIT_FILE(INIT_FILE),
        .INIT_000(INIT_000),
        .INIT_001(INIT_001),
        .INIT_002(INIT_002),
        .INIT_003(INIT_003),
        .INIT_004(INIT_004),
        .INIT_005(INIT_005),
        .INIT_006(INIT_006),
        .INIT_007(INIT_007),
        .INIT_008(INIT_008),
        .INIT_009(INIT_009),
        .INIT_00A(INIT_00A),
        .INIT_00B(INIT_00B),
        .INIT_00C(INIT_00C),
        .INIT_00D(INIT_00D),
        .INIT_00E(INIT_00E),
        .INIT_00F(INIT_00F),
        .INIT_010(INIT_010),
        .INIT_011(INIT_011),
        .INIT_012(INIT_012),
        .INIT_013(INIT_013),
        .INIT_014(INIT_014),
        .INIT_015(INIT_015),
        .INIT_016(INIT_016),
        .INIT_017(INIT_017),
        .INIT_018(INIT_018),
        .INIT_019(INIT_019),
        .INIT_01A(INIT_01A),
        .INIT_01B(INIT_01B),
        .INIT_01C(INIT_01C),
        .INIT_01D(INIT_01D),
        .INIT_01E(INIT_01E),
        .INIT_01F(INIT_01F),
        .INIT_020(INIT_020),
        .INIT_021(INIT_021),
        .INIT_022(INIT_022),
        .INIT_023(INIT_023),
        .INIT_024(INIT_024),
        .INIT_025(INIT_025),
        .INIT_026(INIT_026),
        .INIT_027(INIT_027),
        .INIT_028(INIT_028),
        .INIT_029(INIT_029),
        .INIT_02A(INIT_02A),
        .INIT_02B(INIT_02B),
        .INIT_02C(INIT_02C),
        .INIT_02D(INIT_02D),
        .INIT_02E(INIT_02E),
        .INIT_02F(INIT_02F),
        .INIT_030(INIT_030),
        .INIT_031(INIT_031),
        .INIT_032(INIT_032),
        .INIT_033(INIT_033),
        .INIT_034(INIT_034),
        .INIT_035(INIT_035),
        .INIT_036(INIT_036),
        .INIT_037(INIT_037),
        .INIT_038(INIT_038),
        .INIT_039(INIT_039),
        .INIT_03A(INIT_03A),
        .INIT_03B(INIT_03B),
        .INIT_03C(INIT_03C),
        .INIT_03D(INIT_03D),
        .INIT_03E(INIT_03E),
        .INIT_03F(INIT_03F),
        .INIT_040(INIT_040),
        .INIT_041(INIT_041),
        .INIT_042(INIT_042),
        .INIT_043(INIT_043),
        .INIT_044(INIT_044),
        .INIT_045(INIT_045),
        .INIT_046(INIT_046),
        .INIT_047(INIT_047),
        .INIT_048(INIT_048),
        .INIT_049(INIT_049),
        .INIT_04A(INIT_04A),
        .INIT_04B(INIT_04B),
        .INIT_04C(INIT_04C),
        .INIT_04D(INIT_04D),
        .INIT_04E(INIT_04E),
        .INIT_04F(INIT_04F),
        .INIT_050(INIT_050),
        .INIT_051(INIT_051),
        .INIT_052(INIT_052),
        .INIT_053(INIT_053),
        .INIT_054(INIT_054),
        .INIT_055(INIT_055),
        .INIT_056(INIT_056),
        .INIT_057(INIT_057),
        .INIT_058(INIT_058),
        .INIT_059(INIT_059),
        .INIT_05A(INIT_05A),
        .INIT_05B(INIT_05B),
        .INIT_05C(INIT_05C),
        .INIT_05D(INIT_05D),
        .INIT_05E(INIT_05E),
        .INIT_05F(INIT_05F),
        .INIT_060(INIT_060),
        .INIT_061(INIT_061),
        .INIT_062(INIT_062),
        .INIT_063(INIT_063),
        .INIT_064(INIT_064),
        .INIT_065(INIT_065),
        .INIT_066(INIT_066),
        .INIT_067(INIT_067),
        .INIT_068(INIT_068),
        .INIT_069(INIT_069),
        .INIT_06A(INIT_06A),
        .INIT_06B(INIT_06B),
        .INIT_06C(INIT_06C),
        .INIT_06D(INIT_06D),
        .INIT_06E(INIT_06E),
        .INIT_06F(INIT_06F),
        .INIT_070(INIT_070),
        .INIT_071(INIT_071),
        .INIT_072(INIT_072),
        .INIT_073(INIT_073),
        .INIT_074(INIT_074),
        .INIT_075(INIT_075),
        .INIT_076(INIT_076),
        .INIT_077(INIT_077),
        .INIT_078(INIT_078),
        .INIT_079(INIT_079),
        .INIT_07A(INIT_07A),
        .INIT_07B(INIT_07B),
        .INIT_07C(INIT_07C),
        .INIT_07D(INIT_07D),
        .INIT_07E(INIT_07E),
        .INIT_07F(INIT_07F),
        .INIT_080(INIT_080),
        .INIT_081(INIT_081),
        .INIT_082(INIT_082),
        .INIT_083(INIT_083),
        .INIT_084(INIT_084),
        .INIT_085(INIT_085),
        .INIT_086(INIT_086),
        .INIT_087(INIT_087),
        .INIT_088(INIT_088),
        .INIT_089(INIT_089),
        .INIT_08A(INIT_08A),
        .INIT_08B(INIT_08B),
        .INIT_08C(INIT_08C),
        .INIT_08D(INIT_08D),
        .INIT_08E(INIT_08E),
        .INIT_08F(INIT_08F),
        .INIT_090(INIT_090),
        .INIT_091(INIT_091),
        .INIT_092(INIT_092),
        .INIT_093(INIT_093),
        .INIT_094(INIT_094),
        .INIT_095(INIT_095),
        .INIT_096(INIT_096),
        .INIT_097(INIT_097),
        .INIT_098(INIT_098),
        .INIT_099(INIT_099),
        .INIT_09A(INIT_09A),
        .INIT_09B(INIT_09B),
        .INIT_09C(INIT_09C),
        .INIT_09D(INIT_09D),
        .INIT_09E(INIT_09E),
        .INIT_09F(INIT_09F),
        .INIT_0A0(INIT_0A0),
        .INIT_0A1(INIT_0A1),
        .INIT_0A2(INIT_0A2),
        .INIT_0A3(INIT_0A3),
        .INIT_0A4(INIT_0A4),
        .INIT_0A5(INIT_0A5),
        .INIT_0A6(INIT_0A6),
        .INIT_0A7(INIT_0A7),
        .INIT_0A8(INIT_0A8),
        .INIT_0A9(INIT_0A9),
        .INIT_0AA(INIT_0AA),
        .INIT_0AB(INIT_0AB),
        .INIT_0AC(INIT_0AC),
        .INIT_0AD(INIT_0AD),
        .INIT_0AE(INIT_0AE),
        .INIT_0AF(INIT_0AF),
        .INIT_0B0(INIT_0B0),
        .INIT_0B1(INIT_0B1),
        .INIT_0B2(INIT_0B2),
        .INIT_0B3(INIT_0B3),
        .INIT_0B4(INIT_0B4),
        .INIT_0B5(INIT_0B5),
        .INIT_0B6(INIT_0B6),
        .INIT_0B7(INIT_0B7),
        .INIT_0B8(INIT_0B8),
        .INIT_0B9(INIT_0B9),
        .INIT_0BA(INIT_0BA),
        .INIT_0BB(INIT_0BB),
        .INIT_0BC(INIT_0BC),
        .INIT_0BD(INIT_0BD),
        .INIT_0BE(INIT_0BE),
        .INIT_0BF(INIT_0BF),
        .INIT_0C0(INIT_0C0),
        .INIT_0C1(INIT_0C1),
        .INIT_0C2(INIT_0C2),
        .INIT_0C3(INIT_0C3),
        .INIT_0C4(INIT_0C4),
        .INIT_0C5(INIT_0C5),
        .INIT_0C6(INIT_0C6),
        .INIT_0C7(INIT_0C7),
        .INIT_0C8(INIT_0C8),
        .INIT_0C9(INIT_0C9),
        .INIT_0CA(INIT_0CA),
        .INIT_0CB(INIT_0CB),
        .INIT_0CC(INIT_0CC),
        .INIT_0CD(INIT_0CD),
        .INIT_0CE(INIT_0CE),
        .INIT_0CF(INIT_0CF),
        .INIT_0D0(INIT_0D0),
        .INIT_0D1(INIT_0D1),
        .INIT_0D2(INIT_0D2),
        .INIT_0D3(INIT_0D3),
        .INIT_0D4(INIT_0D4),
        .INIT_0D5(INIT_0D5),
        .INIT_0D6(INIT_0D6),
        .INIT_0D7(INIT_0D7),
        .INIT_0D8(INIT_0D8),
        .INIT_0D9(INIT_0D9),
        .INIT_0DA(INIT_0DA),
        .INIT_0DB(INIT_0DB),
        .INIT_0DC(INIT_0DC),
        .INIT_0DD(INIT_0DD),
        .INIT_0DE(INIT_0DE),
        .INIT_0DF(INIT_0DF),
        .INIT_0E0(INIT_0E0),
        .INIT_0E1(INIT_0E1),
        .INIT_0E2(INIT_0E2),
        .INIT_0E3(INIT_0E3),
        .INIT_0E4(INIT_0E4),
        .INIT_0E5(INIT_0E5),
        .INIT_0E6(INIT_0E6),
        .INIT_0E7(INIT_0E7),
        .INIT_0E8(INIT_0E8),
        .INIT_0E9(INIT_0E9),
        .INIT_0EA(INIT_0EA),
        .INIT_0EB(INIT_0EB),
        .INIT_0EC(INIT_0EC),
        .INIT_0ED(INIT_0ED),
        .INIT_0EE(INIT_0EE),
        .INIT_0EF(INIT_0EF),
        .INIT_0F0(INIT_0F0),
        .INIT_0F1(INIT_0F1),
        .INIT_0F2(INIT_0F2),
        .INIT_0F3(INIT_0F3),
        .INIT_0F4(INIT_0F4),
        .INIT_0F5(INIT_0F5),
        .INIT_0F6(INIT_0F6),
        .INIT_0F7(INIT_0F7),
        .INIT_0F8(INIT_0F8),
        .INIT_0F9(INIT_0F9),
        .INIT_0FA(INIT_0FA),
        .INIT_0FB(INIT_0FB),
        .INIT_0FC(INIT_0FC),
        .INIT_0FD(INIT_0FD),
        .INIT_0FE(INIT_0FE),
        .INIT_0FF(INIT_0FF),
        .INIT_100(INIT_100),
        .INIT_101(INIT_101),
        .INIT_102(INIT_102),
        .INIT_103(INIT_103),
        .INIT_104(INIT_104),
        .INIT_105(INIT_105),
        .INIT_106(INIT_106),
        .INIT_107(INIT_107),
        .INIT_108(INIT_108),
        .INIT_109(INIT_109),
        .INIT_10A(INIT_10A),
        .INIT_10B(INIT_10B),
        .INIT_10C(INIT_10C),
        .INIT_10D(INIT_10D),
        .INIT_10E(INIT_10E),
        .INIT_10F(INIT_10F),
        .INIT_110(INIT_110),
        .INIT_111(INIT_111),
        .INIT_112(INIT_112),
        .INIT_113(INIT_113),
        .INIT_114(INIT_114),
        .INIT_115(INIT_115),
        .INIT_116(INIT_116),
        .INIT_117(INIT_117),
        .INIT_118(INIT_118),
        .INIT_119(INIT_119),
        .INIT_11A(INIT_11A),
        .INIT_11B(INIT_11B),
        .INIT_11C(INIT_11C),
        .INIT_11D(INIT_11D),
        .INIT_11E(INIT_11E),
        .INIT_11F(INIT_11F),
        .INIT_120(INIT_120),
        .INIT_121(INIT_121),
        .INIT_122(INIT_122),
        .INIT_123(INIT_123),
        .INIT_124(INIT_124),
        .INIT_125(INIT_125),
        .INIT_126(INIT_126),
        .INIT_127(INIT_127),
        .INIT_128(INIT_128),
        .INIT_129(INIT_129),
        .INIT_12A(INIT_12A),
        .INIT_12B(INIT_12B),
        .INIT_12C(INIT_12C),
        .INIT_12D(INIT_12D),
        .INIT_12E(INIT_12E),
        .INIT_12F(INIT_12F),
        .INIT_130(INIT_130),
        .INIT_131(INIT_131),
        .INIT_132(INIT_132),
        .INIT_133(INIT_133),
        .INIT_134(INIT_134),
        .INIT_135(INIT_135),
        .INIT_136(INIT_136),
        .INIT_137(INIT_137),
        .INIT_138(INIT_138),
        .INIT_139(INIT_139),
        .INIT_13A(INIT_13A),
        .INIT_13B(INIT_13B),
        .INIT_13C(INIT_13C),
        .INIT_13D(INIT_13D),
        .INIT_13E(INIT_13E),
        .INIT_13F(INIT_13F),
        .INIT_140(INIT_140),
        .INIT_141(INIT_141),
        .INIT_142(INIT_142),
        .INIT_143(INIT_143),
        .INIT_144(INIT_144),
        .INIT_145(INIT_145),
        .INIT_146(INIT_146),
        .INIT_147(INIT_147),
        .INIT_148(INIT_148),
        .INIT_149(INIT_149),
        .INIT_14A(INIT_14A),
        .INIT_14B(INIT_14B),
        .INIT_14C(INIT_14C),
        .INIT_14D(INIT_14D),
        .INIT_14E(INIT_14E),
        .INIT_14F(INIT_14F),
        .INIT_150(INIT_150),
        .INIT_151(INIT_151),
        .INIT_152(INIT_152),
        .INIT_153(INIT_153),
        .INIT_154(INIT_154),
        .INIT_155(INIT_155),
        .INIT_156(INIT_156),
        .INIT_157(INIT_157),
        .INIT_158(INIT_158),
        .INIT_159(INIT_159),
        .INIT_15A(INIT_15A),
        .INIT_15B(INIT_15B),
        .INIT_15C(INIT_15C),
        .INIT_15D(INIT_15D),
        .INIT_15E(INIT_15E),
        .INIT_15F(INIT_15F),
        .INIT_160(INIT_160),
        .INIT_161(INIT_161),
        .INIT_162(INIT_162),
        .INIT_163(INIT_163),
        .INIT_164(INIT_164),
        .INIT_165(INIT_165),
        .INIT_166(INIT_166),
        .INIT_167(INIT_167),
        .INIT_168(INIT_168),
        .INIT_169(INIT_169),
        .INIT_16A(INIT_16A),
        .INIT_16B(INIT_16B),
        .INIT_16C(INIT_16C),
        .INIT_16D(INIT_16D),
        .INIT_16E(INIT_16E),
        .INIT_16F(INIT_16F),
        .INIT_170(INIT_170),
        .INIT_171(INIT_171),
        .INIT_172(INIT_172),
        .INIT_173(INIT_173),
        .INIT_174(INIT_174),
        .INIT_175(INIT_175),
        .INIT_176(INIT_176),
        .INIT_177(INIT_177),
        .INIT_178(INIT_178),
        .INIT_179(INIT_179),
        .INIT_17A(INIT_17A),
        .INIT_17B(INIT_17B),
        .INIT_17C(INIT_17C),
        .INIT_17D(INIT_17D),
        .INIT_17E(INIT_17E),
        .INIT_17F(INIT_17F),
        .INIT_180(INIT_180),
        .INIT_181(INIT_181),
        .INIT_182(INIT_182),
        .INIT_183(INIT_183),
        .INIT_184(INIT_184),
        .INIT_185(INIT_185),
        .INIT_186(INIT_186),
        .INIT_187(INIT_187),
        .INIT_188(INIT_188),
        .INIT_189(INIT_189),
        .INIT_18A(INIT_18A),
        .INIT_18B(INIT_18B),
        .INIT_18C(INIT_18C),
        .INIT_18D(INIT_18D),
        .INIT_18E(INIT_18E),
        .INIT_18F(INIT_18F),
        .INIT_190(INIT_190),
        .INIT_191(INIT_191),
        .INIT_192(INIT_192),
        .INIT_193(INIT_193),
        .INIT_194(INIT_194),
        .INIT_195(INIT_195),
        .INIT_196(INIT_196),
        .INIT_197(INIT_197),
        .INIT_198(INIT_198),
        .INIT_199(INIT_199),
        .INIT_19A(INIT_19A),
        .INIT_19B(INIT_19B),
        .INIT_19C(INIT_19C),
        .INIT_19D(INIT_19D),
        .INIT_19E(INIT_19E),
        .INIT_19F(INIT_19F),
        .INIT_1A0(INIT_1A0),
        .INIT_1A1(INIT_1A1),
        .INIT_1A2(INIT_1A2),
        .INIT_1A3(INIT_1A3),
        .INIT_1A4(INIT_1A4),
        .INIT_1A5(INIT_1A5),
        .INIT_1A6(INIT_1A6),
        .INIT_1A7(INIT_1A7),
        .INIT_1A8(INIT_1A8),
        .INIT_1A9(INIT_1A9),
        .INIT_1AA(INIT_1AA),
        .INIT_1AB(INIT_1AB),
        .INIT_1AC(INIT_1AC),
        .INIT_1AD(INIT_1AD),
        .INIT_1AE(INIT_1AE),
        .INIT_1AF(INIT_1AF),
        .INIT_1B0(INIT_1B0),
        .INIT_1B1(INIT_1B1),
        .INIT_1B2(INIT_1B2),
        .INIT_1B3(INIT_1B3),
        .INIT_1B4(INIT_1B4),
        .INIT_1B5(INIT_1B5),
        .INIT_1B6(INIT_1B6),
        .INIT_1B7(INIT_1B7),
        .INIT_1B8(INIT_1B8),
        .INIT_1B9(INIT_1B9),
        .INIT_1BA(INIT_1BA),
        .INIT_1BB(INIT_1BB),
        .INIT_1BC(INIT_1BC),
        .INIT_1BD(INIT_1BD),
        .INIT_1BE(INIT_1BE),
        .INIT_1BF(INIT_1BF),
        .INIT_1C0(INIT_1C0),
        .INIT_1C1(INIT_1C1),
        .INIT_1C2(INIT_1C2),
        .INIT_1C3(INIT_1C3),
        .INIT_1C4(INIT_1C4),
        .INIT_1C5(INIT_1C5),
        .INIT_1C6(INIT_1C6),
        .INIT_1C7(INIT_1C7),
        .INIT_1C8(INIT_1C8),
        .INIT_1C9(INIT_1C9),
        .INIT_1CA(INIT_1CA),
        .INIT_1CB(INIT_1CB),
        .INIT_1CC(INIT_1CC),
        .INIT_1CD(INIT_1CD),
        .INIT_1CE(INIT_1CE),
        .INIT_1CF(INIT_1CF),
        .INIT_1D0(INIT_1D0),
        .INIT_1D1(INIT_1D1),
        .INIT_1D2(INIT_1D2),
        .INIT_1D3(INIT_1D3),
        .INIT_1D4(INIT_1D4),
        .INIT_1D5(INIT_1D5),
        .INIT_1D6(INIT_1D6),
        .INIT_1D7(INIT_1D7),
        .INIT_1D8(INIT_1D8),
        .INIT_1D9(INIT_1D9),
        .INIT_1DA(INIT_1DA),
        .INIT_1DB(INIT_1DB),
        .INIT_1DC(INIT_1DC),
        .INIT_1DD(INIT_1DD),
        .INIT_1DE(INIT_1DE),
        .INIT_1DF(INIT_1DF),
        .INIT_1E0(INIT_1E0),
        .INIT_1E1(INIT_1E1),
        .INIT_1E2(INIT_1E2),
        .INIT_1E3(INIT_1E3),
        .INIT_1E4(INIT_1E4),
        .INIT_1E5(INIT_1E5),
        .INIT_1E6(INIT_1E6),
        .INIT_1E7(INIT_1E7),
        .INIT_1E8(INIT_1E8),
        .INIT_1E9(INIT_1E9),
        .INIT_1EA(INIT_1EA),
        .INIT_1EB(INIT_1EB),
        .INIT_1EC(INIT_1EC),
        .INIT_1ED(INIT_1ED),
        .INIT_1EE(INIT_1EE),
        .INIT_1EF(INIT_1EF),
        .INIT_1F0(INIT_1F0),
        .INIT_1F1(INIT_1F1),
        .INIT_1F2(INIT_1F2),
        .INIT_1F3(INIT_1F3),
        .INIT_1F4(INIT_1F4),
        .INIT_1F5(INIT_1F5),
        .INIT_1F6(INIT_1F6),
        .INIT_1F7(INIT_1F7),
        .INIT_1F8(INIT_1F8),
        .INIT_1F9(INIT_1F9),
        .INIT_1FA(INIT_1FA),
        .INIT_1FB(INIT_1FB),
        .INIT_1FC(INIT_1FC),
        .INIT_1FD(INIT_1FD),
        .INIT_1FE(INIT_1FE),
        .INIT_1FF(INIT_1FF),
        .RAM_MODE("TRUE_DUAL_PORT")
    ) bram (
        .CLKA(CLKA), .CEA(CEA), .WEA(WEA), .BEA({2'b0, BEA}),
        .ADDRA(ADDRA), .DIA({18'b0, DIA}),
        .ORCEA(ORCEA), .CLRA(RSTA), .DOA({dangle_a18, DOA}),
        .CLKB(CLKB), .CEB(CEB), .WEB(WEB), .BEB({2'b0, BEB}),
        .ADDRB(ADDRB), .DIB({18'b0, DIB}),
        .ORCEB(ORCEB), .CLRB(RSTB), .DOB({dangle_b18, DOB})
    );

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_RAM32X1DP.v
//
// Functional description: simple-dual-port 32x1 distributed ram
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_RAM32X1DP
#(
    parameter [31:0] INIT = 32'h00000000
) (
    output  DO,
    input   DI,
    input [4:0] RADDR, WADDR,
    input WCLK, WE
);

    reg [31:0] mem ;

    initial begin
        mem = INIT;
    end

    always @(posedge WCLK) begin
        if (WE == 1'b1) begin
            mem[WADDR] <= DI;
        end
    end

    assign DO = mem[RADDR];

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_OMSER4.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_OMSER4 #(
parameter WL_EXTEND = "FALSE",     //"TRUE"; "FALSE"
parameter GRS_EN = "TRUE", //"TRUE"; "FALSE" 
parameter LRS_EN = "TRUE"   //"TRUE"; "FALSE" 
)(
output  PADO,
output  PADT,
input [3:0] D,
input [1:0] T,
input RCLK,
input SERCLK,
input OCLK,
input RST
);

//synthesis translate_off
reg [3:0] d_rclk;
reg [1:0] t_rclk;
reg [3:0] capture_d_reg;
reg [1:0] capture_t_reg;
reg [3:0] shift_d_reg;
reg [1:0] shift_t_reg;
reg PADO_POS;
reg PADT_reg;
reg PADO_NEG;
reg rstn_dly;
reg capture_en;
reg rstn_dly_oclk;
reg rstn_dly_oclk_d;
reg shift_en;

initial begin
d_rclk          = 0;
t_rclk          = 0;
capture_d_reg   = 0;
capture_t_reg   = 0;
shift_d_reg     = 0;
shift_t_reg     = 0;
PADO_POS        = 0;
PADT_reg        = 0;
PADO_NEG        = 0;
rstn_dly        = 0;
capture_en      = 0;
rstn_dly_oclk   = 0;
rstn_dly_oclk_d = 0;
shift_en        = 0;  
end

assign global_rstn = (GRS_EN == "TRUE") ? GRS_INST.GRSNET : 1'b1; 
assign lsr_rstn = LRS_EN == "TRUE" ? (~RST) : 1'b1;

always @(posedge RCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn) begin
      d_rclk <= 0;
      t_rclk <= 0;
   end   
   else if (!lsr_rstn) begin
      d_rclk <= 0;
      t_rclk <= 0;
   end   
   else begin
      d_rclk <= D;
      t_rclk <= T;
   end   

always @(posedge SERCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn) begin
      rstn_dly       <= 0;
      capture_en <= 0;
   end
   else if (!lsr_rstn) begin
      rstn_dly       <= 0;
      capture_en <= 0;
   end   
   else begin
      rstn_dly       <= 1;
      if (rstn_dly)
        capture_en <= ~ capture_en;     
      

   end

always @(posedge SERCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn) begin
      capture_d_reg <= 0;
      capture_t_reg <= 0;
   end
   else if (!lsr_rstn) begin
      capture_d_reg <= 0;
      capture_t_reg <= 0;
   end   
   else begin
      if (capture_en) begin
         capture_d_reg <= d_rclk;
         capture_t_reg <= t_rclk;     
      end
   end 

assign rstn_dly_oclk_tmp = (WL_EXTEND == "TRUE") ? rstn_dly_oclk : rstn_dly_oclk_d;

always @(posedge OCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn) begin
      rstn_dly_oclk       <= 0;
      rstn_dly_oclk_d     <= 0;
      shift_en <= 0;
   end
   else if (!lsr_rstn) begin
      rstn_dly_oclk       <= 0;
      rstn_dly_oclk_d     <= 0;
      shift_en <= 0;
   end   
   else begin
      rstn_dly_oclk       <= 1;
      rstn_dly_oclk_d     <= rstn_dly_oclk;
      if (rstn_dly_oclk_tmp)
        shift_en <= ~ shift_en;     
   end
   
always @(posedge OCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn) begin
      shift_d_reg <= 0;
      shift_t_reg <= 0;
   end   
   else if (!lsr_rstn) begin
      shift_d_reg <= 0;
      shift_t_reg <= 0;
   end   
   else if (shift_en) begin
      shift_d_reg <= capture_d_reg;
      shift_t_reg <= capture_t_reg;
   end
   else begin
      shift_d_reg <= {2'd0, shift_d_reg[3:2]};
      shift_t_reg <= {1'b0, shift_t_reg[1]};        
   end
   
always @(posedge OCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn) begin
      PADO_POS <= 0;
      PADT_reg <= 0;
   end
   else if (!lsr_rstn) begin
      PADO_POS <= 0;
      PADT_reg <= 0;
   end
   else begin
      PADO_POS <= shift_d_reg[1];
      PADT_reg <= shift_t_reg[0];     
   end           
   
always @(negedge OCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn) begin
      PADO_NEG <= 0;
   end
   else if (!lsr_rstn) begin
      PADO_NEG <= 0;
   end
   else begin
      PADO_NEG <= shift_d_reg[0];
   end           
   
assign PADO =  OCLK ? PADO_NEG : PADO_POS;
assign PADT = PADT_reg;

//synthesis translate_on

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: Internal simulation model
// Filename: GTP_INBUFE.v
//
// Functional description: Input Buffer
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_INBUFE #(
    parameter IOSTANDARD = "DEFAULT",
    parameter TERM_DDR = "ON"
)(
    output reg O,
    input EN,                    // 1: enable inbuf, normal mode; 0: disable inbuf, standby mode.
    input I
) /* synthesis syn_black_box */ ;
  
  initial begin
    case (IOSTANDARD)
    "LVTTL33", "PCI33", "LVCMOS33", "LVCMOS25", "LVCMOS18", "LVCMOS15", "LVCMOS12", "SSTL25_I", "SSTL25_II", "SSTL18_I", "SSTL18_II", "SSTL15_I", "SSTL15_II", "HSTL18_I", "HSTL18_II", "HSTL15_I", "SSTL15_I_CAL", "SSTL15_II_CAL", "HSTL15_I_CAL", "DEFAULT" :;
    default : begin
           $display("Attribute Syntax Error : The attribute IOSTANDARD on GTP_INBUF instance %m is set to %s.", IOSTANDARD);
           $finish;
              end
    endcase

    case (TERM_DDR)
    "ON", "OFF" :;
    default : begin
           $display("Attribute Syntax Error : The attribute TERM_DDR on GTP_INBUF instance %m is set to %s.", TERM_DDR);
           $finish;
              end
    endcase
    end

    always @(*)
    begin
        if (EN == 1'b1)
            O = I;
        else
            O = 1'b1;
    end

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_OUTBUFTCO.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_OUTBUFTCO #(
    parameter IOSTANDARD = "DEFAULT"
)(
    output O,
    output OB,
    input I,
    input T
) /* synthesis syn_black_box */ ;
  
  initial begin
    case (IOSTANDARD)
    "SSTL18D_I", "SSTL18D_II", "SSTL15D_I", "SSTL15D_II", "HSTL15D_I", "SSTL25D_I", "SSTL25D_II", "SSTL15D_I_CAL", "SSTL15D_II_CAL", "HSTL15D_I_CAL","LVPECL",
    "LVDS25E", "LVCMOS25D", "LVCMOS33D", "RSDS", "PPDS","BLVDS", "DEFAULT" :;
    default : begin
           $display("Attribute Syntax Error : The attribute IOSTANDARD on GTP_OUTBUFTCO instance %m is set to %s.", IOSTANDARD);
           $finish;
              end
    endcase
    end
    bufif0 (O, I, T);
    notif0 (OB, I, T);

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_MULT36.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

//P=A*B
module GTP_MULT36 #(
    parameter GRS_EN    = "TRUE", //"TRUE"; "FALSE"
    parameter SYNC_RST  = "FALSE", //"TRUE"; "FALSE"
    parameter INREG_EN  = "FALSE", //"TRUE"; "FALSE"
    parameter OUTREG_EN = "FALSE"  //"TRUE"; "FALSE"
) (
    output  [54-1:0] P,
    input   CE,
    input   RST,
    input   CLK,
    input   A_SIGNED,
    input   [36-1:0] A,
    input   B_SIGNED,
    input   [18-1:0] B
);


    INT_PREADD_MULT #(
        .GRS_EN(GRS_EN),
        .SYNC_RST(SYNC_RST),
        .INREG_EN(INREG_EN),
        .OUTREG_EN(OUTREG_EN),
        .ASIZE(36),
        .BSIZE(18),
        .PREADD_EN(0)
    ) U_INT_MULT (
        .CE(CE),
        .RST(RST),
        .CLK(CLK),
        .A_SIGNED(A_SIGNED),
        .A(A),
        .B_SIGNED(B_SIGNED),
        .B(B),
        .C_SIGNED(B_SIGNED),
        .C(18'b0),
        .PREADDSUB(1'b0),
        .P(P)
    );

endmodule






//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_FIR_A.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_FIR_A
#(
    parameter GRS_EN    = "TRUE", //"TRUE"; "FALSE"
    parameter SYNC_RST  = "FALSE", //"TRUE"; "FALSE"
    parameter INREG_EN  = "TRUE",
    parameter OUTREG_EN = "TRUE",
    parameter [1:0] INPUT_OP    = 2'b11,
    parameter [1:0] DYN_OP_SEL  = 2'b11,
    parameter OPCD_DYN_SEL = 1'b0,
    parameter OPCD_CPI_SEL = 1'b0
) (
    output  [17:0] CYO,
    output  CYO_SIGNED,
    output  [63:0] CPO,                  //p
    output   CPO_SIGNED,
    output  [63:0] P,

    input   CE,
    input   RST,
    input   CLK,
    input [17:0] CYI,
    input        CYI_SIGNED,
    input [17:0] Y0,                  //y0 ,DYIA
    input        Y0_SIGNED,
    input [17:0] H0,                  //h0 ,DXIA
    input        H0_SIGNED,
    input [17:0] H1,                  //h1 ,DXIB
    input        H1_SIGNED,
    input [17:0] Y1,                  //y1 ,DYIB
    input        Y1_SIGNED,
    input        OPCD_CPI_DYN,
    input [63:0] CPI,
    input        CPI_SIGNED,
    input        S0,
    input        S1
);

//PSE parameters 
localparam [16:0] SC_PSE_Y0 = 17'b0;  //SC_PSE = 0, disable PSE, parameter bit width=17
localparam [16:0] SC_PSE_Y1 = 17'b0;  //SC_PSE = 0, disable PSE, parameter bit width=17
localparam [16:0] SC_PSE_H0 = 17'b0;  //SC_PSE = 0, disable PSE, parameter bit width=17
localparam [16:0] SC_PSE_H1 = 17'b0;  //SC_PSE = 0, disable PSE, parameter bit width=17

initial begin
    if ((GRS_EN != "TRUE") && (GRS_EN != "FALSE")) begin
        $display("GRS_EN error");
        $finish;
    end
    if ((SYNC_RST != "TRUE") && (SYNC_RST != "FALSE")) begin
        $display("SYNC_RST error");
        $finish;
    end
end

wire [17:0] Y0_PSE;
wire [17:0] Y1_PSE;
wire [17:0] H0_PSE;
wire [17:0] H1_PSE;

reg [17:0] h0_d;
reg        h0_signed_d;
reg [17:0] y0_d;
reg        y0_signed_d;
wire [17:0] y0_sel;
wire        y0_signed_sel;

reg [17:0] h1_d;
reg        h1_signed_d;
reg [17:0] y1_d;
reg        y1_signed_d;
wire [17:0] y1_sel;
wire        y1_signed_sel;

wire [35:0] mult1_in1;
wire [35:0] mult2_in1;
wire [35:0] mult1_in2;
wire [35:0] mult2_in2;

wire [35:0] mult1;
wire        mult1_signed;
wire [35:0] mult2;
wire        mult2_signed;

wire [63:0] ma, mb;
wire [63:0] sum;
wire        sum_signed;
reg  [63:0] sum_d;
reg         sum_signed_d;

wire [17:0] cyo;
reg  [17:0] cyo_d;
wire        cyo_signed;
reg         cyo_signed_d;

wire [17:0] y0_d_sel;
wire [17:0] y1_d_sel;
wire [17:0] h0_d_sel;
wire [17:0] h1_d_sel;
wire  y0_signed_d_sel;
wire  y1_signed_d_sel;
wire  h0_signed_d_sel;
wire  h1_signed_d_sel;
wire  s0_d_sel, s0_sel;
wire  s1_d_sel, s1_sel;

wire global_rstn ;
wire RST_sync ;
wire RST_async;
wire rst_asyncomb ;

wire [63:0] CPI_SEL;
wire        OPCD_SEL;

assign global_rstn = GRS_EN == "TRUE" ? GRS_INST.GRSNET : 1'b1;
assign RST_sync = (SYNC_RST == "TRUE") ? RST : 1'b0;
assign RST_async = (SYNC_RST == "FALSE") ? RST : 1'b0;
assign rst_asyncomb = RST_async | (~global_rstn);

assign OPCD_SEL = (OPCD_DYN_SEL == 1'b1)?OPCD_CPI_DYN :OPCD_CPI_SEL;
assign CPI_SEL  = (OPCD_SEL == 1'b1)? 64'b0 : CPI; 

initial begin
    {h0_signed_d, h0_d} = 'b0;
    {y0_signed_d, y0_d} = 'b0;
    {h1_signed_d, h1_d} = 'b0;
    {y1_signed_d, y1_d} = 'b0;
    {cyo_signed_d, cyo_d} = 19'b0;
    {sum_signed_d, sum_d} = 65'b0;
end

INT_REG #(.SIZE(2)) USEL (.Q({s1_d_sel, s0_d_sel}),
    .BYPASS(INREG_EN == "TRUE" ? 1'b0 : 1'b1),
    .D({S1, S0}),
    .CLK(CLK), .CE(CE), .ARST(rst_asyncomb), .SRST(RST_sync));
assign s0_sel = (DYN_OP_SEL[0] == 1'b1) ? s0_d_sel : INPUT_OP[0];
assign s1_sel = (DYN_OP_SEL[1] == 1'b1) ? s1_d_sel : INPUT_OP[1];

always @(posedge CLK or posedge rst_asyncomb)
    if (rst_asyncomb || RST_sync) begin
        {h0_signed_d, h0_d} <= 'b0;
        {y0_signed_d, y0_d} <= 'b0;
    end
    else if (CE) begin
        {h0_signed_d, h0_d} <= {H0_SIGNED, H0_PSE};
        {y0_signed_d, y0_d} <= {y0_signed_sel, Y0_PSE};
    end

always @(posedge CLK or posedge rst_asyncomb)
    if (rst_asyncomb || RST_sync) begin
        {h1_signed_d, h1_d} <= 'b0;
        {y1_signed_d, y1_d} <= 'b0;
    end
    else if (CE) begin
        {h1_signed_d, h1_d} <= {H1_SIGNED, H1_PSE};
        {y1_signed_d, y1_d} <= {y1_signed_sel, Y1_PSE};
    end

INT_PSE #(.ASIZE(18),.SC_PSE(SC_PSE_Y0)) U1_PSE(.A(y0_sel),.SIGN(y0_signed_sel),.A_PSE(Y0_PSE));
INT_PSE #(.ASIZE(18),.SC_PSE(SC_PSE_Y1)) U2_PSE(.A(y1_sel),.SIGN(y1_signed_sel),.A_PSE(Y1_PSE));
INT_PSE #(.ASIZE(18),.SC_PSE(SC_PSE_H0)) U3_PSE(.A(H0),    .SIGN(H0_SIGNED),    .A_PSE(H0_PSE));
INT_PSE #(.ASIZE(18),.SC_PSE(SC_PSE_H1)) U4_PSE(.A(H1),    .SIGN(H1_SIGNED),    .A_PSE(H1_PSE));

assign {y0_signed_sel, y0_sel} = s0_sel ? {CYI_SIGNED, CYI} : {Y0_SIGNED, Y0};  // default s0  = 1
assign {y1_signed_sel, y1_sel} = s1_sel ? {y0_signed_d_sel, y0_d_sel} : {Y1_SIGNED, Y1};  //s1  = 1

assign {cyo_signed, cyo} = {y1_signed_d_sel, y1_d_sel};

assign {y0_signed_d_sel, y0_d_sel} = (INREG_EN == "TRUE")? {y0_signed_d, y0_d} : {y0_signed_sel, Y0_PSE};
assign {y1_signed_d_sel, y1_d_sel} = (INREG_EN == "TRUE")? {y1_signed_d, y1_d} : {y1_signed_sel, Y1_PSE};
assign {h0_signed_d_sel, h0_d_sel} = (INREG_EN == "TRUE")? {h0_signed_d, h0_d} : {H0_SIGNED, H0_PSE};
assign {h1_signed_d_sel, h1_d_sel} = (INREG_EN == "TRUE")? {h1_signed_d, h1_d} : {H1_SIGNED, H1_PSE};


assign mult1_in1 = {{18{y0_signed_d_sel & y0_d_sel[17]}},y0_d_sel};
assign mult2_in1 = {{18{y1_signed_d_sel & y1_d_sel[17]}},y1_d_sel};
assign mult1_in2 = {{18{h0_signed_d_sel & h0_d_sel[17]}},h0_d_sel};
assign mult2_in2 = {{18{h1_signed_d_sel & h1_d_sel[17]}},h1_d_sel};

assign mult1 = mult1_in1 * mult1_in2;
assign mult1_signed = y0_signed_d_sel | h0_signed_d_sel;
assign mult2 = mult2_in1 * mult2_in2;
assign mult2_signed = y1_signed_d_sel | h1_signed_d_sel;

assign ma = {{28{mult1_signed&mult1[35]}},mult1};
assign mb = {{28{mult2_signed&mult2[35]}},mult2};
assign sum = ma + mb + CPI_SEL;
assign sum_signed = mult1_signed | mult2_signed | CPI_SIGNED;


always @(posedge CLK or posedge rst_asyncomb)
    if (rst_asyncomb || RST_sync) begin
        {cyo_signed_d, cyo_d} <= 19'b0;
        {sum_signed_d, sum_d} <= 65'b0;
    end
    else if (CE) begin
        {cyo_signed_d, cyo_d} <= {cyo_signed, cyo};
        {sum_signed_d, sum_d} <= {sum_signed, sum};
    end

assign {CYO_SIGNED, CYO} = (OUTREG_EN == "TRUE")? {cyo_signed_d, cyo_d} : {cyo_signed, cyo};
assign {CPO_SIGNED, CPO} = (OUTREG_EN == "TRUE")? {sum_signed_d, sum_d} : {sum_signed, sum};
assign P = CPO;

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_DRM18K.v
//
// Functional description:
//
// Parameter  description:
//
// Port description:
//
// Revision history:
//   2018/01/09: Update display informations.
//   2018/04/02: Update to support LOGOS device.
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_DRM18K
#(
    parameter GRS_EN = "TRUE",
    parameter [2:0] CSA_MASK = 3'b000,
    parameter [2:0] CSB_MASK = 3'b000,
    parameter integer DATA_WIDTH_A = 18,
    parameter integer DATA_WIDTH_B = 18,
    parameter WRITE_MODE_A = "NORMAL_WRITE",
    parameter WRITE_MODE_B = "NORMAL_WRITE",
    parameter integer DOA_REG = 0,
    parameter integer DOB_REG = 0,
    parameter integer DOA_REG_CLKINV = 0,
    parameter integer DOB_REG_CLKINV = 0,
    parameter RST_TYPE = "SYNC",
    parameter RAM_MODE = "TRUE_DUAL_PORT",
    parameter WRITE_COLLISION_ARBITER = "NULL",
    parameter SIM_DEVICE = "TITAN",
    parameter [287:0] INIT_00 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_01 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_02 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_03 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_04 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_05 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_06 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_07 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_08 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_09 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_10 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_11 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_12 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_13 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_14 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_15 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_16 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_17 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_18 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_19 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_20 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_21 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_22 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_23 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_24 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_25 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_26 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_27 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_28 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_29 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_2A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_2B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_2C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_2D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_2E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_2F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_30 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_31 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_32 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_33 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_34 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_35 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_36 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_37 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_38 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_39 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_3A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_3B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_3C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_3D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_3E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_3F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_FILE = "NONE",
    parameter integer BLOCK_X = 0,
    parameter integer BLOCK_Y = 0,
    parameter integer RAM_DATA_WIDTH = 9,
    parameter integer RAM_ADDR_WIDTH = 11,
    parameter INIT_FORMAT = "BIN"
) (
    output [17:0] DOA,
    output [17:0] DOB,
    output WWCONF,
    input [17:0] DIA,
    input [17:0] DIB,
    input [13:0] ADDRA,
    input ADDRA_HOLD,
    input [13:0] ADDRB,
    input ADDRB_HOLD,
    input [2:0] CSA,
    input [2:0] CSB,
    input CLKA,
    input CLKB,
    input CEA,
    input CEB,
    input WEA,
    input WEB,
    input ORCEA,
    input ORCEB,
    input RSTA,
    input RSTB
);

    localparam  BLOCK_DEPTH = (2**(DATA_WIDTH_A == 1 ? 14 :    // block type 16k*1
                                  DATA_WIDTH_A == 2 ? 13 :    // block type 8k*2
                                  DATA_WIDTH_A == 4 ? 12 :    // block type 4k*4
                                  DATA_WIDTH_A <= 9 ? 11 :    // block type 2k*8 or 2k*9
                                 DATA_WIDTH_A <= 18 ? 10 : 9)); // block type 512*36 or 512*32     block memory address width

    localparam  BLOCK_WIDTH =   DATA_WIDTH_A;             //block memory data width
//end add for initialization

    localparam MEM_SIZE = 18432;
    localparam width_a = (DATA_WIDTH_A == 32) ? 16 : (DATA_WIDTH_A == 36) ? 18 : DATA_WIDTH_A;
    localparam width_b = (DATA_WIDTH_B == 32) ? 16 : (DATA_WIDTH_B == 36) ? 18 : DATA_WIDTH_B;

    integer  cnt;
    reg [9-1:0] mem [MEM_SIZE/9-1:0];

    //reg [2:0] csa_reg = 3'b0, csb_reg = 3'b0;
    reg csa_reg = 1'b0, csb_reg = 1'b0;
    reg [13:0] ada_reg = 14'b0, adb_reg = 14'b0;
    reg [17:0] da_reg = 18'b0, db_reg = 18'b0;
    reg wea_reg = 1'b0, web_reg = 1'b0;
    wire [3:0] bea_reg;   // modify for byte_write_enable bug
    wire [1:0] beb_reg;
    wire write_en_a, write_en_b, read_en_a, read_en_b;
    wire CEA_int,CEB_int;

    reg [17:0] a_out = 18'b0, a_out_reg = 18'b0;
    //reg [17:0] a_out_reg_sync = 18'b0, a_out_reg_async = 18'b0, a_out_reg_async_sy = 18'b0;
    reg [17:0] b_out = 18'b0, b_out_reg = 18'b0;
    //reg [17:0] b_out_reg_sync = 18'b0, b_out_reg_async = 18'b0, b_out_reg_async_sy = 18'b0;

    wire grs, rsta_grs, rstb_grs;
    reg rsta_async_sy = 1'b0, rstb_async_sy = 1'b0;
    wire rsta_grs_sync;
    wire rstb_grs_sync;
    wire rsta_grs_async;
    wire rstb_grs_async;
    wire rsta_async_synrel;
    wire rstb_async_synrel;
    wire rsta_int;
    wire rstb_int;
    
    reg [17:0] doa;
    reg [17:0] dob;

    initial begin
        doa = 0;
        dob = 0;
    end

// synthesis translate_off
// add for memory initialization 2014/7/2 10:59:37    1) add ini_mem reg array to load init.dat
//                                                    2) init_file contain all the initial data of cascaded DRMS
   reg [RAM_DATA_WIDTH-1:0] ini_mem [2**RAM_ADDR_WIDTH-1:0];
   integer p;
   initial
   begin
      if(INIT_FILE != "NONE")
      begin
          if(INIT_FORMAT == "BIN")
              $readmemb(INIT_FILE,ini_mem);
          else
              $readmemh(INIT_FILE,ini_mem);
          for(p=0;p<20;p=p+1)
              $display("ini_mem[%d] = %b",p,ini_mem[p]);
      end
   end
//end  add
///////////////////
// parameter check
///////////////////
    initial begin
        case (DATA_WIDTH_A)
            1, 2, 4, 8, 16, 32: begin
                case (DATA_WIDTH_B)
                    1, 2, 4, 8, 16, 32:  ; //null
                    default: begin
                        $display("ERROR: GTP_DRM18K instance %m parameter DATA_WIDTH_B:%d is illegal. The legal values are 1,2,4,8,16 or 32.",DATA_WIDTH_B);
                        $finish;
                    end
                endcase
            end
            9, 18, 36: begin
                case (DATA_WIDTH_B)
                    9, 18, 36:    ; //null
                    default: begin
                        $display("ERROR: GTP_DRM18K instance %m parameter DATA_WIDTH_B:%d is illegal. The legal values are 9,18 or 36.",DATA_WIDTH_B);
                        $finish;
                    end
                endcase
            end
            default: begin
                $display("ERROR: GTP_DRM18K instance %m parameter DATA_WIDTH_A:%d is illegal. The legal values are 1,2,4,8,9,16,18,32 or 36.",DATA_WIDTH_A);
                $finish;
            end
        endcase

        case (WRITE_MODE_A)
            "NORMAL_WRITE",
            "TRANSPARENT_WRITE",
            "READ_BEFORE_WRITE":    ; //null 
            default: begin
                $display("ERROR: GTP_DRM18K instance %m parameter WRITE_MODE_A: %s is illegal. The legal values are NORMAL_WRITE,TRANSPARENT_WRITE or READ_BEFORE_WRITE.", WRITE_MODE_A);
                $finish;
            end
        endcase

        case (WRITE_MODE_B)
            "NORMAL_WRITE",
            "TRANSPARENT_WRITE",
            "READ_BEFORE_WRITE":    ; //null  
            default: begin
                $display("ERROR: GTP_DRM18K instance %m parameter WRITE_MODE_B: %s is illegal. The legal values are NORMAL_WRITE,TRANSPARENT_WRITE or READ_BEFORE_WRITE.", WRITE_MODE_B);
                $finish;
            end
        endcase

        case (RST_TYPE)
            "ASYNC",
            "ASYNC_SYNC_RELEASE",
            "SYNC":     ;//null
            default: begin
                $display("ERROR: GTP_DRM18K instance %m parameter RST_TYPE: %s is illegal. The legal values are ASYNC,ASYNC_SYNC_RELEASE or SYNC.", RST_TYPE);
                $finish;
            end
        endcase

        case (RAM_MODE)
            "ROM",
            "SINGLE_PORT","SIMPLE_DUAL_PORT":     ;//null
            "TRUE_DUAL_PORT": begin
                if (DATA_WIDTH_A > 18 || DATA_WIDTH_B > 18) begin
                    $display("ERROR: GTP_DRM18K instance %m parameter DATA_WIDTH_A and DATA_WIDTH_B in TRUE_DUAL_PORT MODE:%d,%d is illegal. The legal values are 1,2,4,8,9,16 or 18.",DATA_WIDTH_A,DATA_WIDTH_B);
                    $finish;
                end
            end
            default: begin
                $display("ERROR: GTP_DRM18K instance %m parameter RAM_MODE value: %s is illegal. The legal values are ROM or SINGLE_PORT, SIMPLE_DUAL_PORT or TRUE_DUAL_PORT.", RAM_MODE);
                $finish;
            end
        endcase

        case (SIM_DEVICE)
            "TITAN","LOGOS","PGL22G":    ;//null
            default: begin
                $display("ERROR: GTP_DRM18K instance %m parameter SIM_DEVICE value: %s is illegal. The legal values are TITAN or LOGOS or PGL22G.", SIM_DEVICE);
                $finish;
            end
        endcase

        case (WRITE_COLLISION_ARBITER)
            "NULL":     ;//null
            //"PORTA", "PORTB": begin
            //    if( (DATA_WIDTH_A != DATA_WIDTH_B) && (RAM_MODE != "TRUE_DUAL_PORT") ) begin
            //        $display("DRM18K display: Illegal DATA_WIDTH_A DATA_WIDTH_B RAM_MODE value when WRITE_COLLISION_ARBITER != NULL:%s,%s,%s,%s",DATA_WIDTH_A,DATA_WIDTH_B,RAM_MODE,WRITE_COLLISION_ARBITER);
            //        $finish;
            //    end
            // end
            default: begin
                $display("ERROR: GTP_DRM18K instance %m parameter WRITE_COLLISION_ARBITER: %s is illegal. The legal values is NULL.",WRITE_COLLISION_ARBITER);
                $finish;
            end
        endcase

    end

/////////////////=
// initialization
/////////////////=

    initial begin
        if (INIT_FILE == "NONE") begin
            for (cnt = 0; cnt < 32; cnt = cnt + 1) begin
                mem[32*0 + cnt] = INIT_00[cnt*9 +: 9];
                mem[32*1 + cnt] = INIT_01[cnt*9 +: 9];
                mem[32*2 + cnt] = INIT_02[cnt*9 +: 9];
                mem[32*3 + cnt] = INIT_03[cnt*9 +: 9];
                mem[32*4 + cnt] = INIT_04[cnt*9 +: 9];
                mem[32*5 + cnt] = INIT_05[cnt*9 +: 9];
                mem[32*6 + cnt] = INIT_06[cnt*9 +: 9];
                mem[32*7 + cnt] = INIT_07[cnt*9 +: 9];
                mem[32*8 + cnt] = INIT_08[cnt*9 +: 9];
                mem[32*9 + cnt] = INIT_09[cnt*9 +: 9];
                mem[32*10 + cnt] = INIT_0A[cnt*9 +: 9];
                mem[32*11 + cnt] = INIT_0B[cnt*9 +: 9];
                mem[32*12 + cnt] = INIT_0C[cnt*9 +: 9];
                mem[32*13 + cnt] = INIT_0D[cnt*9 +: 9];
                mem[32*14 + cnt] = INIT_0E[cnt*9 +: 9];
                mem[32*15 + cnt] = INIT_0F[cnt*9 +: 9];
                mem[32*16 + cnt] = INIT_10[cnt*9 +: 9];
                mem[32*17 + cnt] = INIT_11[cnt*9 +: 9];
                mem[32*18 + cnt] = INIT_12[cnt*9 +: 9];
                mem[32*19 + cnt] = INIT_13[cnt*9 +: 9];
                mem[32*20 + cnt] = INIT_14[cnt*9 +: 9];
                mem[32*21 + cnt] = INIT_15[cnt*9 +: 9];
                mem[32*22 + cnt] = INIT_16[cnt*9 +: 9];
                mem[32*23 + cnt] = INIT_17[cnt*9 +: 9];
                mem[32*24 + cnt] = INIT_18[cnt*9 +: 9];
                mem[32*25 + cnt] = INIT_19[cnt*9 +: 9];
                mem[32*26 + cnt] = INIT_1A[cnt*9 +: 9];
                mem[32*27 + cnt] = INIT_1B[cnt*9 +: 9];
                mem[32*28 + cnt] = INIT_1C[cnt*9 +: 9];
                mem[32*29 + cnt] = INIT_1D[cnt*9 +: 9];
                mem[32*30 + cnt] = INIT_1E[cnt*9 +: 9];
                mem[32*31 + cnt] = INIT_1F[cnt*9 +: 9];
                mem[32*32 + cnt] = INIT_20[cnt*9 +: 9];
                mem[32*33 + cnt] = INIT_21[cnt*9 +: 9];
                mem[32*34 + cnt] = INIT_22[cnt*9 +: 9];
                mem[32*35 + cnt] = INIT_23[cnt*9 +: 9];
                mem[32*36 + cnt] = INIT_24[cnt*9 +: 9];
                mem[32*37 + cnt] = INIT_25[cnt*9 +: 9];
                mem[32*38 + cnt] = INIT_26[cnt*9 +: 9];
                mem[32*39 + cnt] = INIT_27[cnt*9 +: 9];
                mem[32*40 + cnt] = INIT_28[cnt*9 +: 9];
                mem[32*41 + cnt] = INIT_29[cnt*9 +: 9];
                mem[32*42 + cnt] = INIT_2A[cnt*9 +: 9];
                mem[32*43 + cnt] = INIT_2B[cnt*9 +: 9];
                mem[32*44 + cnt] = INIT_2C[cnt*9 +: 9];
                mem[32*45 + cnt] = INIT_2D[cnt*9 +: 9];
                mem[32*46 + cnt] = INIT_2E[cnt*9 +: 9];
                mem[32*47 + cnt] = INIT_2F[cnt*9 +: 9];
                mem[32*48 + cnt] = INIT_30[cnt*9 +: 9];
                mem[32*49 + cnt] = INIT_31[cnt*9 +: 9];
                mem[32*50 + cnt] = INIT_32[cnt*9 +: 9];
                mem[32*51 + cnt] = INIT_33[cnt*9 +: 9];
                mem[32*52 + cnt] = INIT_34[cnt*9 +: 9];
                mem[32*53 + cnt] = INIT_35[cnt*9 +: 9];
                mem[32*54 + cnt] = INIT_36[cnt*9 +: 9];
                mem[32*55 + cnt] = INIT_37[cnt*9 +: 9];
                mem[32*56 + cnt] = INIT_38[cnt*9 +: 9];
                mem[32*57 + cnt] = INIT_39[cnt*9 +: 9];
                mem[32*58 + cnt] = INIT_3A[cnt*9 +: 9];
                mem[32*59 + cnt] = INIT_3B[cnt*9 +: 9];
                mem[32*60 + cnt] = INIT_3C[cnt*9 +: 9];
                mem[32*61 + cnt] = INIT_3D[cnt*9 +: 9];
                mem[32*62 + cnt] = INIT_3E[cnt*9 +: 9];
                mem[32*63 + cnt] = INIT_3F[cnt*9 +: 9];
            end
        end
        else  begin      // INIT_FILE 
//add for initialization RAM     1) load initial data from ini_mem to every mem block  when  cascaded with DRMS
// 2) the ini_mem contain  the whole data of init_file  3) distribute the initdata to every mem in cascaded DRMs
            case(DATA_WIDTH_A)
                1: begin  //DRM TYPE 16K*1
                   for(cnt=0; cnt<2*1024;cnt = cnt+1)
                       mem[cnt][7:0] = {ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*8+7][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*8+6][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*8+5][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*8+4][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*8+3][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*8+2][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*8+1][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*8][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH]};
                end
                2: begin //DRM TYPE 8K*2
                   for(cnt=0; cnt<2*1024;cnt = cnt+1)
                       mem[cnt][7:0] = {ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*4+3][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*4+2][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*4+1][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*4][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH]};
                end
                4: begin //DRM TYPE 4K*4
                   for(cnt=0; cnt<2*1024;cnt = cnt+1)
                       {mem[cnt][7:0]} = {ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*2+1][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                          ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*2][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH]};
                end
                8: begin //DRM TYPE 2K*8
                   for(cnt=0; cnt<2*1024;cnt = cnt+1)
                       mem[cnt][7:0] = ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH];
                end
                9: begin //DRM TYPE 2K*9
                   for(cnt=0; cnt<2*1024;cnt = cnt+1)
                       mem[cnt] = ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH];
                end
                16:begin //DRM TYPE 1K*16
                   for(cnt=0; cnt<1024;cnt = cnt+1)
                       {mem[cnt*2+1][7:0], mem[cnt*2][7:0]} = ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH];
                end
                18:begin //DRM TYPE 1K*18
                   for(cnt=0; cnt<1024;cnt = cnt+1)
                       {mem[cnt*2+1], mem[cnt*2]} = ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH];
                end
                32:begin //DRM TYPE 512*32
                   for(cnt=0; cnt<512;cnt = cnt+1)
                       {mem[cnt*4+3][7:0],mem[cnt*4+2][7:0],mem[cnt*4+1][7:0],mem[cnt*4][7:0]} = ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH];
                end
                36:begin //DRM TYPE 512*36
                   for(cnt=0; cnt<512;cnt = cnt+1)
                       {mem[cnt*4+3],mem[cnt*4+2],mem[cnt*4+1],mem[cnt*4]} = ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH];
                end
            endcase
        end
    end

//write confilction process, only used when following conditions are matched
//DP RAM with CLKA = CLKB
//DATA_WIDTH_A=DATA_WIDTH_B
//ADDRA_HOLD&ADDRB_HOLD hardwired to 0
assign write_conflict = (CSA == CSA_MASK) && (CSB == CSB_MASK) && (ADDRA == ADDRB) && WEA && WEB; //&& (WRITE_COLLISION_ARBITER != "NULL") ;
assign wea_enable = write_conflict ? (WRITE_COLLISION_ARBITER != "PORTB") : 1'b1;
assign web_enable = write_conflict ? (WRITE_COLLISION_ARBITER != "PORTA") : 1'b1;

assign WWCONF = write_conflict;

/////////////////////////////////////////////////////
//
/////////////////////////////////////////////////////
generate
    case (SIM_DEVICE)
        "TITAN","PGL22G" : begin
            assign CEA_int = CEA & (CSA == CSA_MASK);
            assign CEB_int = CEB & (CSB == CSB_MASK);
        end
        "LOGOS" : begin
            assign CEA_int = CEA;
            assign CEB_int = CEB;
            always @(posedge CLKA) begin
                if(CEA_int && (ADDRA_HOLD == 1'b0)) csa_reg <= (CSA == CSA_MASK);
            end
            always @(posedge CLKB) begin
                if(CEB_int && (ADDRB_HOLD == 1'b0)) csb_reg <= (CSB == CSB_MASK);
            end
        end
    endcase
endgenerate

    always @(posedge CLKA) begin
        if (CEA_int) begin
            // high to hold the address
            if (ADDRA_HOLD == 1'b0) begin
                ada_reg <= ADDRA;
            end
            da_reg[17:0] <= DIA[17:0];
            wea_reg <= WEA && wea_enable;
        end
    end

    always @(posedge CLKB) begin
        if (CEB_int) begin
            // high to hold the address
            if (ADDRB_HOLD == 1'b0) begin
                adb_reg <= ADDRB;
            end
                web_reg <= WEB && web_enable;
        end
    end
    // byte write enable
    assign bea_reg = ada_reg[3:0];   // modify for byte_write_enable bug
    assign beb_reg = adb_reg[1:0];

    ///////////////////
    // task & function
    ///////////////////

    function [DATA_WIDTH_A-1:0] mem_read_a;
        input [13:0]  addr;
    begin
        case (DATA_WIDTH_A)
            1: mem_read_a = mem[addr[13:3]][addr[2:0]];
            2: mem_read_a = mem[addr[13:3]][addr[2:1]*2 +: 2];
            4: mem_read_a = mem[addr[13:3]][addr[2]*4 +: 4];
            8: mem_read_a = mem[addr[13:3]][7:0];
            9: mem_read_a = mem[addr[13:3]];
            16: mem_read_a = {mem[addr[13:4]*2+1][7:0], mem[addr[13:4]*2][7:0]};
            18: mem_read_a = {mem[addr[13:4]*2+1],      mem[addr[13:4]*2]};
            32: mem_read_a = {mem[addr[13:5]*4+3][7:0], mem[addr[13:5]*4+2][7:0],
                              mem[addr[13:5]*4+1][7:0], mem[addr[13:5]*4][7:0]};
            36: mem_read_a = {mem[addr[13:5]*4+3],      mem[addr[13:5]*4+2],
                              mem[addr[13:5]*4+1],      mem[addr[13:5]*4]};
            default:      ;//null 
        endcase
    end
    endfunction

    function [DATA_WIDTH_B-1:0] mem_read_b;
        input [13:0] addr;
    begin
        case (DATA_WIDTH_B)
            1: mem_read_b = mem[addr[13:3]][addr[2:0]];
            2: mem_read_b = mem[addr[13:3]][addr[2:1]*2 +: 2];
            4: mem_read_b = mem[addr[13:3]][addr[2]*4 +: 4];
            8: mem_read_b = mem[addr[13:3]][7:0];
            9: mem_read_b = mem[addr[13:3]];
            16: mem_read_b = {mem[addr[13:4]*2+1][7:0], mem[addr[13:4]*2][7:0]};
            18: mem_read_b = {mem[addr[13:4]*2+1],      mem[addr[13:4]*2]};
            32: mem_read_b = {mem[addr[13:5]*4+3][7:0], mem[addr[13:5]*4+2][7:0],
                              mem[addr[13:5]*4+1][7:0], mem[addr[13:5]*4][7:0]};
            36: mem_read_b = {mem[addr[13:5]*4+3],      mem[addr[13:5]*4+2],
                              mem[addr[13:5]*4+1],      mem[addr[13:5]*4]};
            default:      ;//null
        endcase
    end
    endfunction

    task mem_write_a;
        input [13:0] addr;
        input [35:0] data;
        input [3:0]  byte_en;
    begin
        case (DATA_WIDTH_A)
            1: mem[addr[13:3]][addr[2:0]] = data[0];
            2: mem[addr[13:3]][addr[2:1]*2 +: 2] = data[1:0];
            4: mem[addr[13:3]][addr[2]*4 +: 4] = data[3:0];
            8: mem[addr[13:3]][7:0] = data[7:0];
            9: mem[addr[13:3]] = data[8:0];
            16: begin
                if (byte_en[1])
                    mem[addr[13:4]*2+1][7:0] = data[16:9];
                if (byte_en[0])
                    mem[addr[13:4]*2][7:0]   = data[7:0];
            end
            18: begin
                if (byte_en[1])
                    mem[addr[13:4]*2+1] = data[17:9];
                if (byte_en[0])
                    mem[addr[13:4]*2]   = data[8:0];
            end
            32: begin
                if (byte_en[3])
                    mem[addr[13:5]*4+3][7:0] = data[34:27];
                if (byte_en[2])
                    mem[addr[13:5]*4+2][7:0] = data[25:18];
                if (byte_en[1])
                    mem[addr[13:5]*4+1][7:0] = data[16:9];
                if (byte_en[0])
                    mem[addr[13:5]*4][7:0]   = data[7:0];
            end
            36: begin
                if (byte_en[3])
                    mem[addr[13:5]*4+3] = data[35:27];
                if (byte_en[2])
                    mem[addr[13:5]*4+2] = data[26:18];
                if (byte_en[1])
                    mem[addr[13:5]*4+1] = data[17:9];
                if (byte_en[0])
                    mem[addr[13:5]*4]   = data[8:0];
            end
            default:     ;//null
        endcase
    end
    endtask

    task mem_write_b;
        input [13:0] addr;
        input [17:0] data;
        input [3:0]  byte_en;
    begin
        case (DATA_WIDTH_B)
            1: mem[addr[13:3]][addr[2:0]] = data[0];
            2: mem[addr[13:3]][addr[2:1]*2 +: 2] = data[1:0];
            4: mem[addr[13:3]][addr[2]*4 +: 4] = data[3:0];
            8: mem[addr[13:3]][7:0] = data[7:0];
            9: mem[addr[13:3]] = data[8:0];
            16: begin
                if (byte_en[1])
                    mem[addr[13:4]*2+1][7:0] = data[16:9];
                if (byte_en[0])
                    mem[addr[13:4]*2][7:0]   = data[7:0];
            end
            18: begin
                if (byte_en[1])
                    mem[addr[13:4]*2+1] = data[17:9];
                if (byte_en[0])
                    mem[addr[13:4]*2]   = data[8:0];
            end
            default:     ;//null
        endcase
    end
    endtask

    ///////////////
    // memory core
    ///////////////
reg CLKA_active;
reg CLKB_active;
initial begin
  CLKA_active = 1'b0;
  CLKB_active = 1'b0;
end
always @(posedge CLKA) begin
   if (CEA_int) begin
      CLKA_active <= 1'b1;
      #0.2 CLKA_active = 1'b0;
   end
   else
      CLKA_active <= 1'b0;
end
always @(posedge CLKB) begin
   if (CEB_int) begin
      CLKB_active <= 1'b1;
      #0.2 CLKB_active = 1'b0;
   end
   else
      CLKB_active <= 1'b0;
end

generate
////////////////////////////////////////////////////////////////////////////////////////////
// ROM or SINGLE_PORT 
////////////////////////////////////////////////////////////////////////////////////////////
if(RAM_MODE == "ROM" || RAM_MODE == "SINGLE_PORT") begin:ROMorSP_MODE  //1 no clock region switch  2 no mix width

    always @(posedge CLKA) begin    //modify for db_reg syn with CLKA
        if (CEA_int)
            db_reg[17:0] <= DIB[17:0];
    end
    if (DATA_WIDTH_A >= 32 || DATA_WIDTH_B >= 32) begin

    case(SIM_DEVICE)
        "TITAN" : begin
            assign write_en_a = 1'b1;
            assign read_en_b  = 1'b1;
        end 
        "PGL22G" : begin
            assign write_en_a = (wea_reg == 1'b1);
            assign read_en_b  = (web_reg == 1'b0);
        end
        "LOGOS" : begin
            assign write_en_a = csa_reg & (wea_reg == 1'b1);
            assign read_en_b  = csb_reg & (web_reg == 1'b0);
        end
    endcase
        // Port A operations
        always @(negedge CLKA_active) begin
            if (write_en_a) begin  // write
                mem_write_a(ada_reg, {db_reg[17:0], da_reg[17:0]}, bea_reg[3:0]);
            end
        end
        always@(negedge CLKB_active or posedge rstb_int) begin
            if (rstb_int)
               {b_out[width_b-1:0], a_out[width_b-1:0]} = 'b0;
            else if(read_en_b)
               {b_out[width_b-1:0], a_out[width_b-1:0]} = mem_read_b(adb_reg);
        end

    end
    else  begin   //x1 x2 x4 x8 x9 x16 x18 

    case(SIM_DEVICE)
        "TITAN","PGL22G": begin
            assign write_en_a = (wea_reg == 1'b1);
            assign read_en_a  = (wea_reg == 1'b0);
        end
        "LOGOS" : begin
            assign write_en_a = csa_reg & (wea_reg == 1'b1);
            assign read_en_a  = csa_reg & (wea_reg == 1'b0);
        end
     endcase
        // Port A operations
        always @(negedge CLKA_active) begin
            if (write_en_a)  begin  // write
               // read during write
               if (WRITE_MODE_A == "TRANSPARENT_WRITE") begin
                   a_out[width_a-1:0] = mem_read_a(ada_reg);

                   if(DATA_WIDTH_A == 16) begin
                       if(bea_reg[0])
                           a_out[7:0] = da_reg[7:0];
                       else
                           a_out[7:0] = a_out[7:0];

                       if(bea_reg[1])
                           a_out[15:8] = da_reg[16:9];
                       else
                           a_out[15:8] = a_out[15:8];
                   end
                   else if(DATA_WIDTH_A == 18) begin
                        if(bea_reg[0])
                            a_out[8:0] = da_reg[8:0];
                        else
                            a_out[8:0] = a_out[8:0];

                        if(bea_reg[1])
                            a_out[17:9] = da_reg[17:9];
                        else
                            a_out[17:9] = a_out[17:9];
                   end
                   else begin
                      a_out[width_a-1:0] = da_reg[width_a-1:0];
                   end
               end
               else if (WRITE_MODE_A == "READ_BEFORE_WRITE")
                   a_out[width_a-1:0] = mem_read_a(ada_reg);

               mem_write_a(ada_reg, da_reg[17:0], {2'b0,bea_reg[1:0]});
            end
        end

        always @(negedge CLKA_active or posedge rsta_int) begin
            if (rsta_int)
               a_out[width_a-1:0] = 'b0;
            else if (read_en_a)          // read 
               a_out[width_a-1:0] = mem_read_a(ada_reg);
        end
        // Port B operations

    end
end
////////////////////////////////////////////////////////////////////////////////////////////
//SIMPLE_DUAL_PORT
////////////////////////////////////////////////////////////////////////////////////////////
else if(RAM_MODE == "SIMPLE_DUAL_PORT")begin:SDP_MODE  //1 clock region switch 2 mix width
    //port_A operation: only write in SDP MODE
    if (DATA_WIDTH_A >= 32) begin:PORTA

        case(SIM_DEVICE)
            "TITAN" :  assign write_en_a = wea_enable;
            "PGL22G" : assign write_en_a = (wea_reg == 1'b1);
            "LOGOS" :  assign write_en_a = csa_reg & (wea_reg == 1'b1);
        endcase

        always @(posedge CLKA) begin
           if (CEA_int)
              db_reg[17:0]  <= DIB[17:0];   //the valid width of db_reg is equal to da_reg
        end
        always @(negedge CLKA_active) begin
           if (write_en_a)    // write 
              mem_write_a(ada_reg, {db_reg[17:0], da_reg[17:0]},bea_reg[3:0]);
        end
    end
    else  begin:PORTA    //  x1 x2 x4 x8 x9 x16 x18 

        case(SIM_DEVICE)
            "TITAN" :  assign write_en_a  = (wea_reg == 1'b1) & wea_enable;
            "PGL22G" : assign write_en_a  = (wea_reg == 1'b1);
            "LOGOS" :  assign write_en_a  = csa_reg & (wea_reg == 1'b1);
        endcase

        always @(negedge CLKA_active) begin
           if (write_en_a)     // write 
              mem_write_a(ada_reg, da_reg[17:0], {2'b0,bea_reg[1:0]});
        end
    end
    //port_B operation:only read in SDP MODE
    if (DATA_WIDTH_B >= 32) begin:PORTB
// SIMPLE_DUAL_PORT
        case(SIM_DEVICE)
            "TITAN" :  assign read_en_b  = web_enable;
            "PGL22G" : assign read_en_b  = (web_reg == 1'b0);
            "LOGOS" :  assign read_en_b  = csb_reg & (web_reg == 1'b0);
        endcase

        always @(negedge CLKB_active or posedge rstb_int) begin
           if (rstb_int)
              {b_out[width_b-1 : 0], a_out[width_b-1 : 0]} = 'b0;
           else if (read_en_b)       // read 
              {b_out[width_b-1 : 0], a_out[width_b-1 : 0]} = mem_read_b(adb_reg);
        end
    end
    else  begin:PORTB  //  x1 x2 x4 x8 x9 x16 x18 

        case(SIM_DEVICE)
            "TITAN" :  assign read_en_b  = (web_reg == 1'b0) && web_enable;
            "PGL22G" : assign read_en_b  = (web_reg == 1'b0);
            "LOGOS" :  assign read_en_b  = csb_reg & (web_reg == 1'b0);
        endcase

        always @(negedge CLKB_active or posedge rstb_int) begin
           if (rstb_int)
              b_out[width_b-1 : 0] = 'b0;
           else if (read_en_b)   //  read 
              b_out[width_b-1 : 0] = mem_read_b(adb_reg);
        end
    end
end
////////////////////////////////////////////////////////////////////////////////////////////
//DP_MODE
////////////////////////////////////////////////////////////////////////////////////////////
else   begin:DP_MODE   //  --x1 x2 x4 x8 x9 x16 x18--    1) no clock region switch   2)mix width
    
    case(SIM_DEVICE)
        "TITAN" : begin
            assign write_en_a = (wea_reg == 1'b1) & wea_enable;
            assign read_en_a  = (wea_reg == 1'b0) & wea_enable;
            assign write_en_b = (web_reg == 1'b1) & web_enable;
            assign read_en_b  = (web_reg == 1'b0) & web_enable;
        end
        "PGL22G" : begin
            assign write_en_a = (wea_reg == 1'b1) ;
            assign read_en_a  = (wea_reg == 1'b0) ;
            assign write_en_b = (web_reg == 1'b1) ;
            assign read_en_b  = (web_reg == 1'b0) ;
        end
        "LOGOS" : begin
            assign write_en_a = csa_reg & (wea_reg == 1'b1) ;
            assign read_en_a  = csa_reg & (wea_reg == 1'b0) ;
            assign write_en_b = csb_reg & (web_reg == 1'b1) ;
            assign read_en_b  = csb_reg & (web_reg == 1'b0) ;
        end
    endcase
    // Port A operations
    always @(negedge CLKA_active ) begin
        if (write_en_a)  begin  // write
            // read during write
            if (WRITE_MODE_A == "TRANSPARENT_WRITE") begin
               a_out[width_a-1:0] = mem_read_a(ada_reg);

               if(DATA_WIDTH_A == 16) begin
                   if(bea_reg[0])
                       a_out[7:0] = da_reg[7:0];
                   else
                       a_out[7:0] = a_out[7:0];

                   if(bea_reg[1])
                       a_out[15:8] = da_reg[16:9];
                   else
                       a_out[15:8] = a_out[15:8];
               end
               else if(DATA_WIDTH_A == 18) begin
                    if(bea_reg[0])
                        a_out[8:0] = da_reg[8:0];
                    else
                        a_out[8:0] = a_out[8:0];

                    if(bea_reg[1])
                        a_out[17:9] = da_reg[17:9];
                    else
                        a_out[17:9] = a_out[17:9];
               end
               else begin
                  a_out[width_a-1:0] = da_reg[width_a-1:0];
               end
            end
            else if (WRITE_MODE_A == "READ_BEFORE_WRITE")
                a_out[width_a-1 : 0] = mem_read_a(ada_reg);

            mem_write_a(ada_reg, da_reg[17:0], {2'b0,bea_reg[1:0]});
        end
    end

    always @(negedge CLKA_active or posedge rsta_int) begin
        if (rsta_int)
           a_out[width_a-1 : 0] = 'b0;
        else if (read_en_a)
           a_out[width_a-1 : 0] = mem_read_a(ada_reg);
    end
    // Port B operations
    always @(posedge CLKB) begin  // modify for db_reg syn with CLKB
         if (CEB_int)
            db_reg[17:0] <= DIB[17:0];
    end

    always @(negedge CLKB_active ) begin
        if (write_en_b)  begin  // write
            // read during write
            if (WRITE_MODE_B == "TRANSPARENT_WRITE") begin

                b_out[width_b-1:0] = mem_read_b(adb_reg);

                if(DATA_WIDTH_B == 16) begin
                    if(beb_reg[0])
                        b_out[7:0] = db_reg[7:0];
                    else
                        b_out[7:0] = b_out[7:0];

                    if(beb_reg[1])
                        b_out[15:8] = db_reg[16:9];
                    else
                        b_out[15:8] = b_out[15:8];
                end
                else if(DATA_WIDTH_B == 18) begin
                    if(beb_reg[0])
                        b_out[8:0] = db_reg[8:0];
                    else
                        b_out[8:0] = b_out[8:0];

                    if(beb_reg[1])
                        b_out[17:9] = db_reg[17:9];
                    else
                        b_out[17:9] = b_out[17:9];
                end
                else begin
                   b_out[width_b-1:0] = db_reg[width_b-1:0];
                end
            end
            else if (WRITE_MODE_B == "READ_BEFORE_WRITE")
                b_out[width_b-1 : 0] = mem_read_b(adb_reg);

            mem_write_b(adb_reg, db_reg[17:0], {2'b0,beb_reg[1:0]});
        end
    end

    always @(negedge CLKB_active or posedge rstb_int) begin
        if (rstb_int)
           b_out[width_b-1 : 0] = 'b0;
        else if (read_en_b)
           b_out[width_b-1 : 0] = mem_read_b(adb_reg);
    end
end

endgenerate

    //////////////
    // core latch
    //////////////
    assign grsn =  (GRS_EN == "TRUE") ? GRS_INST.GRSNET : 1'b1;
    assign grs =  ~grsn;
    or (rsta_grs, grs, RSTA);
    or (rstb_grs, grs, RSTB);

wire CLKA_for_or,CLKB_for_or;
wire CLKA_for_rs,CLKB_for_rs;

generate
    case(SIM_DEVICE)
        "TITAN" : begin
            assign CLKA_for_rs = CLKA;
            assign CLKB_for_rs = CLKB;
        end
        default : begin
            assign CLKA_for_rs = CLKA_for_or;
            assign CLKB_for_rs = CLKB_for_or;
        end
    endcase
endgenerate

reg rsta_grsn_d;

    always @(posedge CLKA_for_rs ) begin
        if (RSTA) begin
            rsta_grsn_d   <= 1'b1;
        end
        else begin
            rsta_grsn_d   <= 1'b0;
        end
    end

    always @(posedge CLKA_for_rs or posedge RSTA) begin
        if (RSTA) begin
            rsta_async_sy <= 1'b1;
        end
        else begin
            rsta_async_sy <= rsta_grsn_d;
        end
    end

reg rstb_grsn_d;
    always @(posedge CLKB_for_rs) begin
        if (RSTB) begin
            rstb_grsn_d   <= 1'b1;
        end
        else begin
            rstb_grsn_d   <= 1'b0;
        end
    end

    always @(posedge CLKB_for_rs or posedge RSTB) begin
        if (RSTB) begin
            rstb_async_sy <= 1'b1;
        end
        else begin
            rstb_async_sy <= rstb_grsn_d;
        end
    end

initial begin
    rsta_grsn_d = 1'b1;
    rsta_async_sy = 1'b1;
    rstb_grsn_d = 1'b1;
    rstb_async_sy = 1'b1;
end

assign rsta_grs_sync  = (RST_TYPE == "SYNC") ? rsta_grsn_d : 1'b0; //register to match with CLKA_ative falling edge
assign rstb_grs_sync  = (RST_TYPE == "SYNC") ? rstb_grsn_d : 1'b0; //register to match with CLKA_ative falling edge
assign rsta_grs_async = (RST_TYPE == "ASYNC") ? rsta_grs : grs;
assign rstb_grs_async = (RST_TYPE == "ASYNC") ? rstb_grs : grs;
assign rsta_async_synrel = rsta_async_sy | rsta_grs;
assign rstb_async_synrel = rstb_async_sy | rstb_grs;
assign rsta_int = (RST_TYPE == "ASYNC_SYNC_RELEASE") ? rsta_async_synrel : rsta_grs_sync | rsta_grs_async;
assign rstb_int = (RST_TYPE == "ASYNC_SYNC_RELEASE") ? rstb_async_synrel : rstb_grs_sync | rstb_grs_async;
/////////////////////////////////////////////////////////////////////
//port out
assign CLKA_for_or = (DOA_REG_CLKINV == 1) ? ~CLKA : CLKA;
assign CLKB_for_or = (DOB_REG_CLKINV == 1) ? ~CLKB : CLKB;
generate
if (DATA_WIDTH_B >= 32) begin:FAKE_DP_OUT
    ///////////////////
    // output register
    ///////////////////
    
    always @(posedge CLKB_for_or or posedge rstb_int) begin
        if (rstb_int)
            a_out_reg <= 0;
        else if (ORCEB)
            a_out_reg[width_b-1 : 0] <= a_out[width_b-1 : 0];
    end

    //doa combination logic
    always @(*) begin
        if (DOB_REG == 0)
        begin
            case(DATA_WIDTH_B)
                32: {doa[16:9],doa[7:0]} = {a_out[15:8],a_out[7:0]};
                36:  doa[width_b-1:0] = a_out[width_b-1:0]        ;
            endcase
        end
        else
        begin
            case(DATA_WIDTH_B)
                32: {doa[16:9],doa[7:0]} = {a_out_reg[15:8],a_out_reg[7:0]};
                36:  doa[width_b-1:0] = a_out_reg[width_b-1 : 0];
            endcase
        end
    end

    //port_B output
    
    always @(posedge CLKB_for_or or posedge rstb_int) begin
        if (rstb_int)
            b_out_reg <= 0;
        else if (ORCEB)
            b_out_reg[width_b-1 : 0] <= b_out[width_b-1 : 0];
    end

    //dob combination logic
    always @(*) begin
        if (DOB_REG == 0)
        begin
            case(DATA_WIDTH_B)
                32:{dob[16:9],dob[7:0]} = {b_out[15:8],b_out[7:0]};
                36: dob[width_b-1:0] = b_out[width_b-1 : 0];
            endcase
        end
        else
        begin
            case(DATA_WIDTH_B)
                32:{dob[16:9],dob[7:0]} = {b_out_reg[15:8],b_out_reg[7:0]};
                36: dob[width_b-1:0] = b_out_reg[width_b-1 : 0];
            endcase
        end
    end
end
else  begin:TRUE_DP_OUT   // x1 x2 x4 x8 x9 x16 x18    

    //port_A output

    always @(posedge CLKA_for_or or posedge rsta_int) begin
        if (rsta_int)
            a_out_reg <= 0;
        else if (ORCEA)
            a_out_reg[width_a-1 : 0] <= a_out[width_a-1 : 0];
	end

    //doa combination logic
    always @(*) begin
        if (DOA_REG == 0)
        begin
            case(DATA_WIDTH_A)
               1: {doa[16:9],doa[7:0]} = {16{a_out[width_a-1:0]}};
               2: {doa[16:9],doa[7:0]} = { 8{a_out[width_a-1:0]}};
               4: {doa[16:9],doa[7:0]} = { 4{a_out[width_a-1:0]}};
               8: {doa[16:9],doa[7:0]} = { 2{a_out[width_a-1:0]}};
               9: {doa[17:9],doa[8:0]} = { 2{a_out[width_a-1:0]}};
               16:{doa[16:9],doa[7:0]} =     a_out[width_a-1:0]  ;
               18: doa[17:0]          =     a_out[width_a-1:0]  ;
            endcase
        end
        else
        begin
            case(DATA_WIDTH_A)
               1: {doa[16:9],doa[7:0]} = {16{a_out_reg[width_a-1:0]}};
               2: {doa[16:9],doa[7:0]} = { 8{a_out_reg[width_a-1:0]}};
               4: {doa[16:9],doa[7:0]} = { 4{a_out_reg[width_a-1:0]}};
               8: {doa[16:9],doa[7:0]} = { 2{a_out_reg[width_a-1:0]}};
               9: {doa[17:9],doa[8:0]} = { 2{a_out_reg[width_a-1:0]}};
               16:{doa[16:9],doa[7:0]} =     a_out_reg[width_a-1:0] ;
               18: doa[17:0]          =     a_out_reg[width_a-1:0] ;
            endcase
        end
    end

    //port_B output

    always @(posedge CLKB_for_or or posedge rstb_int) begin
        if (rstb_int)
            b_out_reg <= 0;
        else if (ORCEB)
            b_out_reg[width_b-1 : 0] <= b_out[width_b-1 : 0];
	end
    //dob combination logic
    always @(*) begin

        if (DOB_REG == 0)
        begin
            case(DATA_WIDTH_B)
               1: {dob[16:9],dob[7:0]} = {16{b_out[width_b-1:0]}};
               2: {dob[16:9],dob[7:0]} = { 8{b_out[width_b-1:0]}};
               4: {dob[16:9],dob[7:0]} = { 4{b_out[width_b-1:0]}};
               8: {dob[16:9],dob[7:0]} = { 2{b_out[width_b-1:0]}};
               9: {dob[17:9],dob[8:0]} = { 2{b_out[width_b-1:0]}};
               16:{dob[16:9],dob[7:0]} =     b_out[width_b-1:0] ;
               18: dob[17:0]          =     b_out[width_b-1:0] ;
            endcase
        end
        else
            case(DATA_WIDTH_B)
               1: {dob[16:9],dob[7:0]} = {16{b_out_reg[width_b-1:0]}};
               2: {dob[16:9],dob[7:0]} = { 8{b_out_reg[width_b-1:0]}};
               4: {dob[16:9],dob[7:0]} = { 4{b_out_reg[width_b-1:0]}};
               8: {dob[16:9],dob[7:0]} = { 2{b_out_reg[width_b-1:0]}};
               9: {dob[17:9],dob[8:0]} = { 2{b_out_reg[width_b-1:0]}};
               16:{dob[16:9],dob[7:0]} =     b_out_reg[width_b-1:0] ;
               18: dob[17:0]          =     b_out_reg[width_b-1:0] ;
            endcase
    end
end

endgenerate
assign DOA = doa;
assign DOB = dob;

// synthesis translate_on
endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_LUTMUX4.v
//
// Functional description: Look-Up-Table for 4-to-1 MUX
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_LUTMUX4
(
    output wire Z,
    input wire S0, S1,
    input wire I0, I1, I2, I3
);

    INT_LUTMUX4_UDP (Z, S1, S0, I3, I2, I1, I0);

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_MULT27.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

//P=A*B
module GTP_MULT27 #(
    parameter GRS_EN    = "TRUE", //"TRUE"; "FALSE"
    parameter SYNC_RST  = "FALSE", //"TRUE"; "FALSE"
    parameter INREG_EN  = "FALSE", //"TRUE"; "FALSE"
    parameter OUTREG_EN = "FALSE"  //"TRUE"; "FALSE"
) (
    output  [54-1:0] P,
    input   CE,
    input   RST,
    input   CLK,
    input   A_SIGNED,
    input   [27-1:0] A,
    input   B_SIGNED,
    input   [27-1:0] B
);


    INT_PREADD_MULT #(
        .GRS_EN(GRS_EN),
        .SYNC_RST(SYNC_RST),
        .INREG_EN(INREG_EN),
        .OUTREG_EN(OUTREG_EN),
        .ASIZE(27),
        .BSIZE(27),
        .PREADD_EN(0)
    ) U_INT_MULT (
        .CE(CE),
        .RST(RST),
        .CLK(CLK),
        .A_SIGNED(A_SIGNED),
        .A(A),
        .B_SIGNED(B_SIGNED),
        .B(B),
        .C_SIGNED(B_SIGNED),
        .C(27'b0),
        .PREADDSUB(1'b0),
        .P(P)
    );

endmodule






//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_LUT2.v
//
// Functional description: 2-input Look-Up-Table
//
// Parameter description:
//      INIT: init value
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_LUT2
#(
    parameter [3:0] INIT = 4'h0
) (
    output wire Z,
    input wire I0, I1
);

    INT_LUTMUX4_UDP (Z, I1, I0, INIT[3], INIT[2], INIT[1], INIT[0]);

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_DLATCH_CE.v
//
// Functional description: D-type latch with clear and enable
//
// Parameter description:
//      INIT: init value
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_DLATCH_CE
#(
    parameter GRS_EN = "TRUE",
    parameter INIT = 1'b0
) (
    output reg Q,
    input wire D,
    input wire G, C, GE
);

    wire grs_n;
    wire grs, RS;

    tri1 grsnet = GRS_INST.GRSNET;
    assign grs_n=(GRS_EN=="TRUE")?grsnet:1'b1;

    not (grs, grs_n);
    or (RS, grs, C);

    initial Q = 1'bx;

    always @(D or G or RS or GE) begin
        if (RS)
            Q <= 1'b0;
        else if (G && GE)
            Q <= D;
    end

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_LUT1.v
//
// Functional description: 1-input Look-Up-Table
//
// Parameter description:
//      INIT: init value
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_LUT1
#(
    parameter [1:0] INIT = 2'h0
) (
    output wire Z,
    input wire I0
);

    assign Z = (INIT[0] == INIT[1]) ? INIT[0] : INIT[I0];

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_OMDDR.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_OMDDR #(
parameter GRS_EN = "TRUE", //"TRUE"; "FALSE" 
parameter LRS_EN = "TRUE"   //"TRUE"; "FALSE" 
)(
output  PADO,
output  PADT,
input [1:0] D,
input T,
input RCLK,
input OCLK,
input RST
);

//synthesis translate_off
reg [1:0] d_rclk;
reg t_rclk;
reg [1:0] shift_d_reg;
reg shift_t_reg;
reg PADO_POS;
reg PADT_reg;
reg PADO_NEG;


initial begin
d_rclk      = 0;
t_rclk      = 0;
shift_d_reg = 0;
shift_t_reg = 0;
PADO_POS    = 0;
PADT_reg    = 0;
PADO_NEG    = 0;  
end

assign global_rstn = (GRS_EN == "TRUE") ? GRS_INST.GRSNET : 1'b1; 
assign lsr_rstn = LRS_EN == "TRUE" ? (~RST) : 1'b1;

always @(posedge RCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn) begin
      d_rclk <= 0;
      t_rclk <= 0;
   end   
   else if (!lsr_rstn) begin
      d_rclk <= 0;
      t_rclk <= 0;
   end   
   else begin
      d_rclk <= D;
      t_rclk <= T;
   end   

always @(posedge OCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn) begin
      shift_d_reg <= 0;
      shift_t_reg <= 0;
   end   
   else if (!lsr_rstn) begin
      shift_d_reg <= 0;
      shift_t_reg <= 0;
   end   
   else begin
      shift_d_reg <= d_rclk;
      shift_t_reg <= t_rclk;
   end   
   
always @(posedge OCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn) begin
      PADO_POS <= 0;
      PADT_reg <= 0;
   end
   else if (!lsr_rstn) begin
      PADO_POS <= 0;
      PADT_reg <= 0;
   end
   else begin
      PADO_POS <= shift_d_reg[1];
      PADT_reg <= shift_t_reg;    
   end           
   
always @(negedge OCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn) begin
      PADO_NEG <= 0;
   end
   else if (!lsr_rstn) begin
      PADO_NEG <= 0;
   end
   else begin
      PADO_NEG <= shift_d_reg[0];
   end           


assign PADO =  OCLK ? PADO_NEG : PADO_POS;
assign PADT = PADT_reg;
//synthesis translate_on

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2016 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General Technology Primitive
// Filename: GTP_CRYSTAL.v
//
// Functional description: crystal
//
// Parameter description:
// CLK_EN:  Allow I/O used as crystal
//
// Port description:
// inputs:
// XTALA:       One pin of external crystal
// XTALB:       The other pint of external crystal
// EN_N:          Crystal input enable
//
// outputs:
// CLKOUT:      The clock out of XTAL
//
// Revision: V1.0
//
//////////////////////////////////////////////////////////////////////////////
`timescale 1ns/1ps

module GTP_CRYSTAL
   #(
     parameter CLK_EN = "FALSE" // "TRUE", "FALSE"
     )
    (
     output CLKOUT,

     input 	XTALA,
     input  XTALB,
     input 	EN_N
     )/* synthesis syn_black_box */;

    //synthesis translate_off
	reg 	out_reg;
	
    initial
    begin
        // parameter check
        if ( ("TRUE" == CLK_EN) || ("FALSE" == CLK_EN) )
        begin
        end
        else begin
            $display ("GTP_CRYSTAL error: illegal setting for CLK_EN");
        end

        out_reg = 1'b0;
    end

	assign CLKOUT = ((CLK_EN=="TRUE") && !EN_N) ? out_reg : 1'b0;

    always @(*) begin
        if (XTALA == ~XTALB) begin
            out_reg = XTALA;
        end
        else begin
            out_reg = 1'bx;
        end
    end

    //synthesis translate_on
endmodule // GTP_CRYSTAL




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_ISERDES_E1.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//   2017/12: Remove ISERDES_MODE parameter value "NONE"
//   2018/01/02: delete RST_EN & RSTC_EN
//               update IDDR_MODE
//   2018/03/27: change IDDR_MODE to ISERDES_MODE to follow GTP_ISERDES
//   2018/10/16: delete C part 
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_ISERDES_E1 #(
parameter ISERDES_MODE = "IDES4",   //"IDES4","IDES8","IDES7"
parameter GRS_EN = "TRUE"          //"TRUE"; "FALSE"
)(
output [7:0] DO,
input        DI,
input        ICLK,
input        RCLK,
input        ALIGNWD,
input        RST
)/* synthesis syn_black_box */;

//synthesis translate_off
wire global_rstn;
wire local_rstn;


wire qp7;
wire qp3;
wire update;
wire sel;
wire slip_rst;
wire cnt_en;
wire sel_trig;

reg [7:0] s_r;
reg [7:0] up_r;
reg [7:0] rx_data_reg;

reg       rstn_sync;
reg [2:0] slip_reg;
reg       slip_state;
reg [1:0] cnt;
reg       select_reg;
reg       update_reg;

initial begin
    if(GRS_EN != "TRUE" && GRS_EN != "FALSE")
    begin
      $display("GTP_ISERDES Error: Illegal setting of GRS_EN %s",GRS_EN);
      $finish;
    end
    if(ISERDES_MODE != "IDES4" && ISERDES_MODE != "IDES8" && ISERDES_MODE != "IDES7")
    begin
      $display("GTP_ISERDES Error: Illegal setting of ISERDES_MODE %s",ISERDES_MODE);
      $finish;
    end

    s_r          = 8'b0;
    up_r         = 8'b0;
    rx_data_reg  = 8'b0;
    rstn_sync  = 1'b0;
    slip_reg   = 3'b0;
    slip_state = 1'b0;
    cnt        = 2'b0;
    select_reg = 1'b0;
    update_reg = 1'b0;
end
///////////////////////////////////////////////////////////////////////////
assign global_rstn = (GRS_EN == "TRUE") ? GRS_INST.GRSNET : 1'b1;
assign local_rstn = ~RST;

////////////////////////////////stage 1///////////////////////////////////////////
always @(posedge ICLK or negedge global_rstn or negedge local_rstn) 
begin
   if (!global_rstn)
      {s_r[6],s_r[4],s_r[2], s_r[0]} <= 4'b0;
   else if (!local_rstn)
      {s_r[6],s_r[4],s_r[2], s_r[0]} <= 4'b0;
   else begin
        s_r[6] <= DI;
        s_r[4] <= s_r[6];
        s_r[2] <= (ISERDES_MODE == "IDES4") ? 1'b0 : s_r[4];
        s_r[0] <= s_r[2];
    end
end

always @(negedge ICLK or negedge global_rstn or negedge local_rstn)
begin
   if (!global_rstn)
      {s_r[7],s_r[5],s_r[3],s_r[1]} <= 4'b0;
   else if (!local_rstn)
      {s_r[7],s_r[5],s_r[3],s_r[1]} <= 4'b0;
   else begin
        s_r[7] <= DI;
        s_r[5] <= s_r[7];
        s_r[3] <= (ISERDES_MODE == "IDES4") ? 1'b0 : s_r[5];
        s_r[1] <= s_r[3];
    end
end

///////////////////////stage 2////////////////////////////////////////////
assign qp7 = (ISERDES_MODE == "IDES4") ? s_r[4] : s_r[0];

always @(posedge ICLK or negedge global_rstn or negedge local_rstn)
begin
   if (!global_rstn)
      up_r[7:4] <= 4'b0;
   else if (!local_rstn)
      up_r[7:4] <= 4'b0;
   else 
   begin
        if(update)
        begin
            if(sel)
                up_r[7:4] <= {qp7, s_r[7:5]};
            else
                up_r[7:4] <= s_r[7:4];
        end
    end
end

assign qp3 = (ISERDES_MODE == "IDES4") ? s_r[0] : s_r[4];

always @(posedge ICLK or negedge global_rstn or negedge local_rstn)
begin
   if (!global_rstn)
      up_r[3:0] <= 4'b0;
   else if (!local_rstn)
      up_r[3:0] <= 4'b0;
   else 
   begin
        if(update)
        begin
            if(sel)
                up_r[3:0] <= {qp3, s_r[3:1]};
            else
                up_r[3:0] <= s_r[3:0];
        end
    end
end

always @(posedge RCLK or negedge global_rstn or negedge local_rstn)
begin
   if (!global_rstn)
      rx_data_reg <= 8'b0;
   else if (!local_rstn)
      rx_data_reg <= 8'b0;
   else
      rx_data_reg <= up_r;
end

assign DO = rx_data_reg[7:0];
//////////////////////////////////////////////////////////////////////////

/////////////////////////update & sel & alignwd function part/////////
always @(posedge ICLK or negedge global_rstn or negedge local_rstn)
begin
   if (!global_rstn)
      rstn_sync <= 1'b0;
   else if(!local_rstn)
      rstn_sync <= 1'b0;
   else
      rstn_sync <= 1'b1;
end

always @(posedge ICLK or negedge rstn_sync)
begin
    if(!rstn_sync)
    begin
        slip_reg <= 3'b0;
    end
    else begin   
        slip_reg <= {slip_reg[1], slip_reg[0], ALIGNWD};
    end
end

assign slip_rst = slip_reg[1] & (~slip_reg[2]);

always @(posedge ICLK or negedge rstn_sync)
begin
    if(!rstn_sync)
         slip_state <= 1'b0;
    else 
    begin
        if(slip_rst)
        begin
            slip_state <= ~slip_state;
        end
        else
            slip_state <= slip_state;
    end
end

assign cnt_en =  (ISERDES_MODE == "IDES7") ? ~slip_rst : ~(slip_state & slip_rst);

assign sel_trig = (ISERDES_MODE == "IDES7") ? ((cnt == 2'b11) & (~select_reg))|(((cnt == 2'b10) & select_reg) & (~slip_rst)) : slip_rst;

always @(posedge ICLK or negedge rstn_sync)
begin
    if(!rstn_sync)
        cnt <= 2'b0;
    else begin
        if(cnt_en)
        begin
            if(ISERDES_MODE == "IDES4")
                cnt[0] <= cnt[0] + 1;
            else begin
                if((ISERDES_MODE == "IDES7")&& select_reg && (cnt == 2'b10))
                    cnt <= 2'b0;
                else
                    cnt <= cnt + 1;
            end
        end
        else
            cnt <= cnt;
    end
end

always @(posedge ICLK or negedge rstn_sync)
begin
    if (!rstn_sync)
        select_reg <= 0;
    else begin
        if(sel_trig == 1'b0)
            select_reg <= select_reg;
        else if(sel_trig == 1'b1)
            select_reg <= ~select_reg;
    end
end

always @(posedge ICLK or negedge rstn_sync)
begin
    if (!rstn_sync)
        update_reg <= 1'b0;
    else begin
        if(ISERDES_MODE == "IDES7")
        begin
            if(select_reg) begin
                update_reg <= (cnt == 2'b00);
            end
            else begin
                update_reg <= (cnt == 2'b01);
            end
        end
        else if(ISERDES_MODE == "IDES4")
        begin
            update_reg <= ~cnt[0];
        end
        else if(ISERDES_MODE == "IDES8")
        begin
            update_reg <= (cnt == 2'b01);
        end
    end
end

assign update = update_reg;
assign sel    = select_reg;

///////////////////////////////////////////////////////////////////////////

//synthesis translate_on

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2016 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_PLL_E1.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1ns/10fs
module GTP_PLL_E1 #(
    parameter real CLKIN_FREQ = 50.0,
    parameter PFDEN_EN        = "FALSE", //"TRUE"; "FALSE"
    parameter VCOCLK_DIV2     = 1'b0,    //1'b0~1'b1
    parameter DYNAMIC_RATIOI_EN = "FALSE", //"TRUE"; "FALSE"
    parameter DYNAMIC_RATIO0_EN = "FALSE", //"TRUE"; "FALSE"
    parameter DYNAMIC_RATIO1_EN = "FALSE", //"TRUE"; "FALSE"
    parameter DYNAMIC_RATIO2_EN = "FALSE", //"TRUE"; "FALSE"
    parameter DYNAMIC_RATIO3_EN = "FALSE", //"TRUE"; "FALSE"
    parameter DYNAMIC_RATIO4_EN = "FALSE", //"TRUE"; "FALSE"
    parameter DYNAMIC_RATIOF_EN = "FALSE", //"TRUE"; "FALSE"
    parameter integer STATIC_RATIOI = 1, //1~512
    parameter integer STATIC_RATIO0 = 1, //1~512
    parameter integer STATIC_RATIO1 = 1, //1~512
    parameter integer STATIC_RATIO2 = 1, //1~512
    parameter integer STATIC_RATIO3 = 1, //1~512
    parameter integer STATIC_RATIO4 = 1, //1~512
    parameter integer STATIC_RATIOF = 1, //1~512
    parameter DYNAMIC_DUTY0_EN = "FALSE", //"TRUE"; "FALSE"
    parameter DYNAMIC_DUTY1_EN = "FALSE", //"TRUE"; "FALSE"
    parameter DYNAMIC_DUTY2_EN = "FALSE", //"TRUE"; "FALSE"
    parameter DYNAMIC_DUTY3_EN = "FALSE", //"TRUE"; "FALSE"
    parameter DYNAMIC_DUTY4_EN = "FALSE", //"TRUE"; "FALSE"
    parameter DYNAMIC_DUTYF_EN = "FALSE", //"TRUE"; "FALSE"
    parameter integer STATIC_DUTY0 = 2, //2<=STATIC_DUTY0<=2*STATIC_RATIO0-2
    parameter integer STATIC_DUTY1 = 2, //2<=STATIC_DUTY1<=2*STATIC_RATIO1-2
    parameter integer STATIC_DUTY2 = 2, //2<=STATIC_DUTY2<=2*STATIC_RATIO2-2
    parameter integer STATIC_DUTY3 = 2, //2<=STATIC_DUTY3<=2*STATIC_RATIO3-2
    parameter integer STATIC_DUTY4 = 2, //2<=STATIC_DUTY4<=2*STATIC_RATIO4-2
    parameter integer STATIC_DUTYF = 2, //2<=STATIC_DUTYF<=2*STATIC_RATIOF-2
    parameter PHASE_ADJUST0_EN  = "FALSE", //"TRUE"; "FALSE"
    parameter PHASE_ADJUST1_EN  = "FALSE", //"TRUE"; "FALSE"
    parameter PHASE_ADJUST2_EN  = "FALSE", //"TRUE"; "FALSE"
    parameter PHASE_ADJUST3_EN  = "FALSE", //"TRUE"; "FALSE"
    parameter PHASE_ADJUST4_EN  = "FALSE", //"TRUE"; "FALSE"
    parameter DYNAMIC_PHASE0_EN = "FALSE", //"TRUE"; "FALSE"
    parameter DYNAMIC_PHASE1_EN = "FALSE", //"TRUE"; "FALSE"
    parameter DYNAMIC_PHASE2_EN = "FALSE", //"TRUE"; "FALSE"
    parameter DYNAMIC_PHASE3_EN = "FALSE", //"TRUE"; "FALSE"
    parameter DYNAMIC_PHASE4_EN = "FALSE", //"TRUE"; "FALSE"
    parameter DYNAMIC_PHASEF_EN = "FALSE", //"TRUE"; "FALSE"
    parameter integer STATIC_PHASE0  = 0, //0~7
    parameter integer STATIC_PHASE1  = 0, //0~7
    parameter integer STATIC_PHASE2  = 0, //0~7
    parameter integer STATIC_PHASE3  = 0, //0~7
    parameter integer STATIC_PHASE4  = 0, //0~7
    parameter integer STATIC_PHASEF  = 0, //0~7
    parameter integer STATIC_CPHASE0 = 2, //2~513
    parameter integer STATIC_CPHASE1 = 2, //2~513
    parameter integer STATIC_CPHASE2 = 2, //2~513
    parameter integer STATIC_CPHASE3 = 2, //2~513
    parameter integer STATIC_CPHASE4 = 2, //2~513
    parameter integer STATIC_CPHASEF = 2, //2~513
    parameter CLK_CAS0_EN = "FALSE", //"TRUE"; "FALSE"
    parameter CLK_CAS1_EN = "FALSE", //"TRUE"; "FALSE"
    parameter CLK_CAS2_EN = "FALSE", //"TRUE"; "FALSE"
    parameter CLK_CAS3_EN = "FALSE", //"TRUE"; "FALSE"
    parameter CLK_CAS4_EN = "FALSE", //"TRUE"; "FALSE"
    parameter integer CLKOUT5_SEL = 0, //0~4
    parameter CLKIN_BYPASS_EN     = "FALSE", //"TRUE"; "FALSE"
    parameter CLKOUT0_SYN_EN      = "FALSE", //"TRUE"; "FALSE"
    parameter CLKOUT0_EXT_SYN_EN  = "FALSE", //"TRUE"; "FALSE"
    parameter CLKOUT1_SYN_EN      = "FALSE", //"TRUE"; "FALSE"
    parameter CLKOUT2_SYN_EN      = "FALSE", //"TRUE"; "FALSE"
    parameter CLKOUT3_SYN_EN      = "FALSE", //"TRUE"; "FALSE"
    parameter CLKOUT4_SYN_EN      = "FALSE", //"TRUE"; "FALSE"
    parameter CLKOUT5_SYN_EN      = "FALSE", //"TRUE"; "FALSE"
    parameter INTERNAL_FB = "ENABLE",  //"ENABLE"; "DISABLE"
    parameter EXTERNAL_FB = "DISABLE", //"CLKOUT0"; "CLKOUT1"; "CLKOUT2"; "CLKOUT3"; "CLKOUT4"; "DISABLE";
    parameter BANDWIDTH   = "OPTIMIZED", //"LOW"; "OPTIMIZED"; "HIGH"
    parameter RSTODIV_PHASE_EN = "TRUE", //"TRUE"; "FALSE"
    parameter SIM_DEVICE = "PGL22G" //"PGL22G"; "PGL35ES"
    )(
    output CLKOUT0,
    output CLKOUT0_EXT,
    output CLKOUT1,
    output CLKOUT2,
    output CLKOUT3,
    output CLKOUT4,
    output CLKOUT5,
    output CLKSWITCH_FLAG,
    output LOCK,
    input CLKIN1,
    input CLKIN2,
    input CLKFB,
    input CLKIN_SEL,
    input CLKIN_SEL_EN,
    input PFDEN,
    input [9:0] RATIOI,
    input [9:0] RATIO0,
    input [9:0] RATIO1,
    input [9:0] RATIO2,
    input [9:0] RATIO3,
    input [9:0] RATIO4,
    input [9:0] RATIOF,
    input [9:0] DUTY0,
    input [9:0] DUTY1,
    input [9:0] DUTY2,
    input [9:0] DUTY3,
    input [9:0] DUTY4,
    input [9:0] DUTYF,
    input [2:0] PHASE0,
    input [2:0] PHASE1,
    input [2:0] PHASE2,
    input [2:0] PHASE3,
    input [2:0] PHASE4,
    input [2:0] PHASEF,
    input [9:0] CPHASE0,
    input [9:0] CPHASE1,
    input [9:0] CPHASE2,
    input [9:0] CPHASE3,
    input [9:0] CPHASE4,
    input [9:0] CPHASEF,
    input CLKOUT0_SYN,
    input CLKOUT0_EXT_SYN,
    input CLKOUT1_SYN,
    input CLKOUT2_SYN,
    input CLKOUT3_SYN,
    input CLKOUT4_SYN,
    input CLKOUT5_SYN,
    input PLL_PWD,
    input RST,
    input RSTODIV_PHASE
    )/* synthesis syn_black_box */;

    initial
    begin
        if((PFDEN_EN == "TRUE") || (PFDEN_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for PFDEN_EN");

        if((DYNAMIC_RATIOI_EN == "TRUE") || (DYNAMIC_RATIOI_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for DYNAMIC_RATIOI_EN");

        if((DYNAMIC_RATIO0_EN == "TRUE") || (DYNAMIC_RATIO0_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for DYNAMIC_RATIO0_EN");

        if((DYNAMIC_RATIO1_EN == "TRUE") || (DYNAMIC_RATIO1_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for DYNAMIC_RATIO1_EN");

        if((DYNAMIC_RATIO2_EN == "TRUE") || (DYNAMIC_RATIO2_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for DYNAMIC_RATIO2_EN");

        if((DYNAMIC_RATIO3_EN == "TRUE") || (DYNAMIC_RATIO3_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for DYNAMIC_RATIO3_EN");

        if((DYNAMIC_RATIO4_EN == "TRUE") || (DYNAMIC_RATIO4_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for DYNAMIC_RATIO4_EN");

        if((DYNAMIC_RATIOF_EN == "TRUE") || (DYNAMIC_RATIOF_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for DYNAMIC_RATIOF_EN");

        if((DYNAMIC_DUTY0_EN == "TRUE") || (DYNAMIC_DUTY0_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for DYNAMIC_DUTY0_EN");

        if((DYNAMIC_DUTY1_EN == "TRUE") || (DYNAMIC_DUTY1_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for DYNAMIC_DUTY1_EN");

        if((DYNAMIC_DUTY2_EN == "TRUE") || (DYNAMIC_DUTY2_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for DYNAMIC_DUTY2_EN");

        if((DYNAMIC_DUTY3_EN == "TRUE") || (DYNAMIC_DUTY3_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for DYNAMIC_DUTY3_EN");

        if((DYNAMIC_DUTY4_EN == "TRUE") || (DYNAMIC_DUTY4_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for DYNAMIC_DUTY4_EN");

        if((DYNAMIC_DUTYF_EN == "TRUE") || (DYNAMIC_DUTYF_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for DYNAMIC_DUTYF_EN");

        if((PHASE_ADJUST0_EN == "TRUE") || (PHASE_ADJUST0_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for PHASE_ADJUST0_EN");

        if((PHASE_ADJUST1_EN == "TRUE") || (PHASE_ADJUST1_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for PHASE_ADJUST1_EN");

        if((PHASE_ADJUST2_EN == "TRUE") || (PHASE_ADJUST2_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for PHASE_ADJUST2_EN");

        if((PHASE_ADJUST3_EN == "TRUE") || (PHASE_ADJUST3_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for PHASE_ADJUST3_EN");

        if((PHASE_ADJUST4_EN == "TRUE") || (PHASE_ADJUST4_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for PHASE_ADJUST4_EN");

        if((DYNAMIC_PHASE0_EN == "TRUE") || (DYNAMIC_PHASE0_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for DYNAMIC_PHASE0_EN");

        if((DYNAMIC_PHASE1_EN == "TRUE") || (DYNAMIC_PHASE1_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for DYNAMIC_PHASE1_EN");

        if((DYNAMIC_PHASE2_EN == "TRUE") || (DYNAMIC_PHASE2_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for DYNAMIC_PHASE2_EN");

        if((DYNAMIC_PHASE3_EN == "TRUE") || (DYNAMIC_PHASE3_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for DYNAMIC_PHASE3_EN");

        if((DYNAMIC_PHASE4_EN == "TRUE") || (DYNAMIC_PHASE4_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for DYNAMIC_PHASE4_EN");

        if((DYNAMIC_PHASEF_EN == "TRUE") || (DYNAMIC_PHASEF_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for DYNAMIC_PHASEF_EN");

        if((CLK_CAS0_EN == "TRUE") || (CLK_CAS0_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for CLK_CAS0_EN");

        if((CLK_CAS1_EN == "TRUE") || (CLK_CAS1_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for CLK_CAS1_EN");

        if((CLK_CAS2_EN == "TRUE") || (CLK_CAS2_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for CLK_CAS2_EN");

        if((CLK_CAS3_EN == "TRUE") || (CLK_CAS3_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for CLK_CAS3_EN");

        if((CLK_CAS4_EN == "TRUE") || (CLK_CAS4_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for CLK_CAS4_EN");

        if((CLKIN_BYPASS_EN == "TRUE") || (CLKIN_BYPASS_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for CLKIN_BYPASS_EN");

        if((CLKOUT0_SYN_EN == "TRUE") || (CLKOUT0_SYN_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for CLKOUT0_SYN_EN");

        if((CLKOUT0_EXT_SYN_EN == "TRUE") || (CLKOUT0_EXT_SYN_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for CLKOUT0_EXT_SYN_EN");

        if((CLKOUT1_SYN_EN == "TRUE") || (CLKOUT1_SYN_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for CLKOUT1_SYN_EN");

        if((CLKOUT2_SYN_EN == "TRUE") || (CLKOUT2_SYN_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for CLKOUT2_SYN_EN");

        if((CLKOUT3_SYN_EN == "TRUE") || (CLKOUT3_SYN_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for CLKOUT3_SYN_EN");

        if((CLKOUT4_SYN_EN == "TRUE") || (CLKOUT4_SYN_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for CLKOUT4_SYN_EN");

        if((CLKOUT5_SYN_EN == "TRUE") || (CLKOUT5_SYN_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for CLKOUT5_SYN_EN");

        if((INTERNAL_FB == "ENABLE") || (INTERNAL_FB == "DISABLE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for INTERNAL_FB");

        if((EXTERNAL_FB == "CLKOUT0") || (EXTERNAL_FB == "CLKOUT1") || (EXTERNAL_FB == "CLKOUT2") || (EXTERNAL_FB == "CLKOUT3") || (EXTERNAL_FB == "CLKOUT4") || (EXTERNAL_FB == "DISABLE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for EXTERNAL_FB");

        if((BANDWIDTH == "LOW") || (BANDWIDTH == "OPTIMIZED") || (BANDWIDTH == "HIGH"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for BANDWIDTH");

        if((RSTODIV_PHASE_EN == "TRUE") || (RSTODIV_PHASE_EN == "FALSE"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for RSTODIV_PHASE_EN");

        if((SIM_DEVICE == "PGL22G") || (SIM_DEVICE == "PGL35ES"))
        begin
        end
        else
            $display ("GTP_PLL_E1 error: illegal setting for SIM_DEVICE");
    end
///////////////////////////////////////////////////////
    wire rstodiv_en;
    wire rst_n, rstodiv_n;
///////////////////////////////////////////////////////
    wire clk_sel, clk_in, clk0, clk1, rstclksw_n;
    reg [1:0] cnt0, cnt1;
    reg dynauto_clkin;
///////////////////////////////////////////////////////
    reg clk_in_first_time, clk_fb_first_time;
    realtime clk_in_first_edge, clk_fb_first_edge;
    reg adjust;
    realtime fb_route_delay, virtual_delay1;
    integer tmp_ratio;
    realtime tmp_delay, real_delay;
///////////////////////////////////////////////////////
    wire pfden;
    reg clk_pfd, vcolow;
    integer cnt;

    reg clk_test, clkwo;
    realtime clk_test_time1 , clk_test_time2, clk_test_time3;
///////////////////////////////////////////////////////
    wire [9:0] idivider, divider0, divider1, divider2, divider3, divider4, fdivider;
    real fsdiv_set_int, fbdiv_set_int;
    reg [5:0] fbdiv_sel;

    wire rstanalog_n;
    realtime clkin_rtime_last, clkin_rtime_next;
    realtime clkin_time, clkin_time1, clkin_time2, clkin_time3;
    reg clkout_lock;
    realtime vcoclk_period, vcoclk_period_half;
    integer  vcoclk_period_amp;
    realtime vcoclk_period_real, vcoclk_period_dev;

    real cnt_fdiv;
    reg clk_gate, inner_clk, vco1_temp, vco2_temp, vco3_temp;
    wire [7:0] vco, clkout;
    reg  vcoclk;
    reg [7:0] vco_div2;
///////////////////////////////////////////////////////
    wire clk_lock;
    reg [2:0] cnt_clkfb;
    reg start_clk;
    reg [10:0] cnt_lock;
    reg lock_reg;
///////////////////////////////////////////////////////
    wire phase_bonding, rst_odiv_n;
    reg [1:0] rst_clk4_n;
    wire [4:0] clk_odivout, clk_cas, phase_adjust;

    wire [2:0] odiv0_fphase;
    wire [9:0] odiv0_cphase, odiv0_duty, odiv0_duty_ctrl;
    wire odiv0_div1;
    reg odiv0_clk_reg;
    reg odiv0_rst_clk0, odiv0_rst_high, odiv0_rst_low;
    reg [1:0] odiv0_rst_sel;
    reg odiv0_gate;
    reg [9:0] odiv0_cnt, odiv0_counter;
    reg odiv0_clkdivr, odiv0_set;

    wire [2:0] odiv1_fphase;
    wire [9:0] odiv1_cphase, odiv1_duty, odiv1_duty_ctrl;
    wire odiv1_div1;
    reg odiv1_clk_reg;
    reg odiv1_rst_clk0, odiv1_rst_high, odiv1_rst_low;
    reg [1:0] odiv1_rst_sel;
    reg odiv1_gate;
    reg [9:0] odiv1_cnt, odiv1_counter;
    reg odiv1_clkdivr, odiv1_set;

    wire [2:0] odiv2_fphase;
    wire [9:0] odiv2_cphase, odiv2_duty, odiv2_duty_ctrl;
    wire odiv2_div1;
    reg odiv2_clk_reg;
    reg odiv2_rst_clk0, odiv2_rst_high, odiv2_rst_low;
    reg [1:0] odiv2_rst_sel;
    reg odiv2_gate;
    reg [9:0] odiv2_cnt, odiv2_counter;
    reg odiv2_clkdivr, odiv2_set;

    wire [2:0] odiv3_fphase;
    wire [9:0] odiv3_cphase, odiv3_duty, odiv3_duty_ctrl;
    wire odiv3_div1;
    reg odiv3_clk_reg;
    reg odiv3_rst_clk0, odiv3_rst_high, odiv3_rst_low;
    reg [1:0] odiv3_rst_sel;
    reg odiv3_gate;
    reg [9:0] odiv3_cnt, odiv3_counter;
    reg odiv3_clkdivr, odiv3_set;

    wire [2:0] odiv4_fphase;
    wire [9:0] odiv4_cphase, odiv4_duty, odiv4_duty_ctrl;
    wire odiv4_div1;
    reg odiv4_clk_reg;
    reg odiv4_rst_clk0, odiv4_rst_high, odiv4_rst_low;
    reg [1:0] odiv4_rst_sel;
    reg odiv4_gate;
    reg [9:0] odiv4_cnt, odiv4_counter;
    reg odiv4_clkdivr, odiv4_set;
///////////////////////////////////////////////////////
    reg [2:0] clk_out0_gate, clk_out0_ext_gate, clk_out1_gate, clk_out2_gate, clk_out3_gate, clk_out4_gate, clk_out5_gate;
    reg clk_out5_reg;
    wire clkout0_en, clkout0_ext_en, clkout1_en, clkout1_adc_en, clkout2_en, clkout3_en, clkout4_en, clkout5_en, clkout4_sel;
    reg inner_rstn;
///////////////////////////////////////////////////////
    initial
    begin
        cnt0 = 2'b00;
        cnt1 = 2'b00;
        dynauto_clkin = 1'b0;
        clk_in_first_time = 1'b0;
        clk_fb_first_time = 1'b0;
        clk_in_first_edge = 0.0;
        clk_fb_first_edge = 0.0;
        fb_route_delay = 0.0;
        tmp_ratio = 0;
        tmp_delay = 0.0;
        real_delay = 0.0;
        clk_pfd = 1'b0; 
        vcolow  = 1'b0;
        cnt     = 0;
        clk_test  = 1'b0;
        clkwo     = 1'b0;
        clk_test_time1 = 0.0;
        clk_test_time2 = 0.0;
        clk_test_time3 = 0.0;
        fsdiv_set_int  = 0.0;
        fbdiv_set_int  = 0.0;
        fbdiv_sel      = 6'b000001;
        clkin_rtime_last = 0.0;
        clkin_rtime_next = 0.0;
        clkin_time  = 0.0;
        clkin_time1 = 0.0;
        clkin_time2 = 0.0;
        clkin_time3 = 0.0;
        clkout_lock = 1'b0;
        vcoclk_period      = 0.0;
        vcoclk_period_half = 0.0;
        vcoclk_period_amp  = 0;
        vcoclk_period_real = 0.0;
        vcoclk_period_dev  = 0.0;
        cnt_fdiv  = 0;
        clk_gate  = 1'b1;
        inner_clk = 1'b0;
        vcoclk    = 1'b0;
        vco1_temp = 1'b0;
        vco2_temp = 1'b0;
        vco3_temp = 1'b0;
        vco_div2 = 8'b0000_0000;
        cnt_clkfb = 3'b000;
        start_clk = 1'b0;
        cnt_lock = 11'b000_0000_0001;
        lock_reg = 0;
        rst_clk4_n = 2'b00;
        odiv0_clk_reg  = 1'b0;
        odiv0_rst_clk0 = 1'b0;
        odiv0_rst_high = 1'b0;
        odiv0_rst_low  = 1'b0;
        odiv0_rst_sel  = 2'b00;
        odiv0_gate    = 1'b0;
        odiv0_cnt     = 10'b00_0000_0000;
        odiv0_counter = 10'b00_0000_0000;
        odiv0_clkdivr = 1'b0;
        odiv0_set     = 1'b0;
        odiv1_clk_reg  = 1'b0;
        odiv1_rst_clk0 = 1'b0;
        odiv1_rst_high = 1'b0;
        odiv1_rst_low  = 1'b0;
        odiv1_rst_sel  = 2'b00;
        odiv1_gate    = 1'b0;
        odiv1_cnt     = 10'b00_0000_0000;
        odiv1_counter = 10'b00_0000_0000;
        odiv1_clkdivr = 1'b0;
        odiv1_set     = 1'b0;
        odiv2_clk_reg  = 1'b0;
        odiv2_rst_clk0 = 1'b0;
        odiv2_rst_high = 1'b0;
        odiv2_rst_low  = 1'b0;
        odiv2_rst_sel  = 2'b00;
        odiv2_gate    = 1'b0;
        odiv2_cnt     = 10'b00_0000_0000;
        odiv2_counter = 10'b00_0000_0000;
        odiv2_clkdivr = 1'b0;
        odiv2_set     = 1'b0;
        odiv3_clk_reg  = 1'b0;
        odiv3_rst_clk0 = 1'b0;
        odiv3_rst_high = 1'b0;
        odiv3_rst_low  = 1'b0;
        odiv3_rst_sel  = 2'b00;
        odiv3_gate    = 1'b0;
        odiv3_cnt     = 10'b00_0000_0000;
        odiv3_counter = 10'b00_0000_0000;
        odiv3_clkdivr = 1'b0;
        odiv3_set     = 1'b0;
        odiv4_clk_reg  = 1'b0;
        odiv4_rst_clk0 = 1'b0;
        odiv4_rst_high = 1'b0;
        odiv4_rst_low  = 1'b0;
        odiv4_rst_sel  = 2'b00;
        odiv4_gate    = 1'b0;
        odiv4_cnt     = 10'b00_0000_0000;
        odiv4_counter = 10'b00_0000_0000;
        odiv4_clkdivr = 1'b0;
        odiv4_set     = 1'b0;
        clk_out0_gate = 3'b000;
        clk_out0_ext_gate = 3'b000;
        clk_out1_gate = 3'b000;
        clk_out2_gate = 3'b000;
        clk_out3_gate = 3'b000;
        clk_out4_gate = 3'b000;
        clk_out5_gate = 3'b000;
        clk_out5_reg  = 1'b0;
        inner_rstn = 1'b0;
        #1;
        inner_rstn = 1'b1;
        clk_in_first_time = 1'b1;
        clk_fb_first_time = 1'b1;
    end
///////////////////////////////////////////////////////
////RESET//////////////////////////////////////////////
    assign rstodiv_en = (RSTODIV_PHASE_EN == "FALSE") ? 1'b0 : 1'b1;

    assign rst_n      = ~(PLL_PWD | RST) & inner_rstn;
    assign rstodiv_n  = rst_n & (~(RSTODIV_PHASE & rstodiv_en));
///////////////////////////////////////////////////////
////INPUT_CLK_SEL//////////////////////////////////////
    assign clk_sel = (CLKIN_SEL_EN == 1'b0) ? dynauto_clkin : CLKIN_SEL;
    assign clk_in  = (clk_sel == 1'b0) ? CLKIN1 : CLKIN2;

    assign clk0 = CLKIN1 & (~CLKIN_SEL_EN);
    assign clk1 = CLKIN2 & (~CLKIN_SEL_EN);

    assign rstclksw_n = ~PLL_PWD & (~CLKIN_SEL_EN) & (~(cnt0[0] & cnt1[0] & (cnt0[1] | cnt1[1]))) & (~((cnt0[1]^cnt0[0]) & (cnt1[1]^cnt1[0])));

    always @(clk0 or negedge rstclksw_n)
    begin
        if(!rstclksw_n)
            cnt0 <= 2'b00;
        else
            cnt0 <= cnt0+1;
    end

    always @(clk1 or negedge rstclksw_n)
    begin
        if(!rstclksw_n)
            cnt1 <= 2'b00;
        else
            cnt1 <= cnt1+1;
    end

    always @(*)
    begin
        if(cnt0 == 2'b11)
            dynauto_clkin <= 1'b0;
        else
            if(cnt1 == 2'b11)
                dynauto_clkin <= 1'b1;
            else
                dynauto_clkin <= dynauto_clkin;
    end

    assign CLKSWITCH_FLAG = dynauto_clkin;
///////////////////////////////////////////////////////
////FBCK_DELAY/////////////////////////////////////////
    always @(posedge clk_in or negedge rst_n)
    begin
        if(!rst_n)
        begin
            clk_in_first_time = 1'b1;
            clk_in_first_edge = 0.0;
        end
        else
        begin
            if(clk_in_first_time == 1'b1)
                clk_in_first_edge = $realtime;
            clk_in_first_time = 1'b0;
        end
    end

    always @(posedge CLKFB or negedge rst_n)
    begin
        if(!rst_n)
        begin
            clk_fb_first_time = 1'b1;
            clk_fb_first_edge = 0.0;
        end
        else
        begin
            if(clk_fb_first_time == 1'b1)
                clk_fb_first_edge = $realtime;
            clk_fb_first_time = 1'b0;
        end
    end
///////////////////////////////////////////////////////
////PFD_ENABLE/////////////////////////////////////////
    assign pfden = (PFDEN_EN == "TRUE") ? PFDEN : 1'b1;

    always # 0.5 clk_pfd = ~clk_pfd;

    always @(posedge clk_pfd or negedge rst_n)
    begin
        if(!rst_n)
        begin
            vcolow <= 0;
            cnt = 0;
        end
        else
            if(pfden)
            begin
                vcolow <= 0;
                cnt = 0;
            end
            else
            begin
                cnt = cnt + 1;
                if(cnt == 500000)
                vcolow <= 1;
            end
    end

    always #200 clk_test = ~clk_test;

    always @(posedge clk_test or negedge rst_n)
    begin
        if(!rst_n)
        begin
            clkwo <= 1'b0;
            clk_test_time1 = 0;
            clk_test_time2 = 0;
            clk_test_time3 = 0;

        end
        else
        begin
            clk_test_time3 = clk_test_time2;
            clk_test_time2 = clk_test_time1;
            clk_test_time1 = clkin_rtime_next;
            if(clk_test_time3 == clk_test_time1)
                clkwo <= 1'b1;
            else
                clkwo <= 1'b0;
        end
    end
///////////////////////////////////////////////////////
////PLL_ANALOG/////////////////////////////////////////
////FEEDBACK_DIVIDER_CAL///////////////////////////////
    assign idivider = (DYNAMIC_RATIOI_EN == "TRUE") ? RATIOI : STATIC_RATIOI;
    assign divider0 = (DYNAMIC_RATIO0_EN == "TRUE") ? RATIO0 : STATIC_RATIO0;
    assign divider1 = (DYNAMIC_RATIO1_EN == "TRUE") ? RATIO1 : STATIC_RATIO1;
    assign divider2 = (DYNAMIC_RATIO2_EN == "TRUE") ? RATIO2 : STATIC_RATIO2;
    assign divider3 = (DYNAMIC_RATIO3_EN == "TRUE") ? RATIO3 : STATIC_RATIO3;
    assign divider4 = (DYNAMIC_RATIO4_EN == "TRUE") ? RATIO4 : STATIC_RATIO4;
    assign fdivider = (DYNAMIC_RATIOF_EN == "TRUE") ? RATIOF : STATIC_RATIOF;

    always @(*)
    begin
        if(INTERNAL_FB == "ENABLE")
        begin
            fsdiv_set_int = fdivider;
            fbdiv_sel = 6'b000001;
        end
        else
            case(EXTERNAL_FB)
                "CLKOUT0": begin
                             fsdiv_set_int = divider0;
                             fbdiv_sel = 6'b000010;
                         end
                "CLKOUT1": begin
                             fsdiv_set_int = divider1;
                             fbdiv_sel = 6'b000100;
                         end
                "CLKOUT2": begin
                             fsdiv_set_int = divider2;
                             fbdiv_sel = 6'b001000;
                         end
                "CLKOUT3": begin
                             fsdiv_set_int = divider3;
                             fbdiv_sel = 6'b010000;
                         end
                "CLKOUT4": begin
                             fsdiv_set_int = divider4;
                             fbdiv_sel = 6'b100000;
                         end
            endcase
    end

    always @(*)
    begin
        if(VCOCLK_DIV2 == 1'b1)
            fbdiv_set_int = fsdiv_set_int * 2;
        else
            fbdiv_set_int = fsdiv_set_int;
    end
////PLL_VCO_CAL////////////////////////////////////////
    assign rstanalog_n = rst_n & ~vcolow;

    always @(posedge clk_in or negedge rstanalog_n)
    begin
        if(!rstanalog_n)
        begin
            clkin_rtime_last = 0.0;
            clkin_rtime_next = 0.0;
            clkin_time  <= 0.0;
            clkin_time1 <= 0.0;
            clkin_time2 <= 0.0;
            clkin_time3 <= 0.0;
            clkout_lock <= 0.0;
            vcoclk_period <= 1'b0;
            vcoclk_period_half <= 0.0;
            vcoclk_period_amp  <= 0.0;
            vcoclk_period_real <= 0.0;
            vcoclk_period_dev  <= 0.0;
        end
        else
        begin
            clkin_rtime_last = clkin_rtime_next;
            clkin_rtime_next = $realtime;
            if(clkin_rtime_last > 0)
            begin
                clkin_time  <= clkin_rtime_next-clkin_rtime_last;
                clkin_time1 <= clkin_time;
                clkin_time2 <= clkin_time1;
                clkin_time3 <= clkin_time2;
            end
            if(clkin_time > 0)
            begin
                clkout_lock <= (clkin_time  > 0) &&
                               (clkin_time1 > 0) &&
                               (clkin_time2 > 0) &&
                               (clkin_time3 > 0) &&
                               ((clkin_time - clkin_time1)  < 0.0001) &&
                               ((clkin_time1 - clkin_time)  < 0.0001) &&
                               ((clkin_time1 - clkin_time2) < 0.0001) &&
                               ((clkin_time2 - clkin_time1) < 0.0001) &&
                               ((clkin_time2 - clkin_time3) < 0.0001) &&
                               ((clkin_time3 - clkin_time2) < 0.0001);
            end
            if(clkin_time > 0)
            begin
                vcoclk_period      = (clkin_time * idivider) / fbdiv_set_int;
                vcoclk_period_half = vcoclk_period / 2;
                vcoclk_period_amp  = vcoclk_period_half * 100000;
                vcoclk_period_real = vcoclk_period_amp / 100000.0;
                vcoclk_period_dev  = (clkin_time - (vcoclk_period_real * 2 * fbdiv_set_int) / idivider) / 2;
            end
        end
    end

    always @(clkout_lock or inner_clk or clkwo)
    begin
        if(clkout_lock == 1'b0 || clkwo == 1'b1)
        begin
            inner_clk <= 1'b0;
            clk_gate  <= 1'b1;
            cnt_fdiv   = 0;
        end
        else
            if(clk_gate == 1)
            begin
                inner_clk <= 1'b1;
                clk_gate  <= 1'b0;
                cnt_fdiv   = 0;
            end
            else
            begin
                cnt_fdiv = cnt_fdiv + 1;
                if(cnt_fdiv  == fbdiv_set_int)
                begin
                    inner_clk <= #(vcoclk_period_half + vcoclk_period_dev) ~inner_clk;
                    cnt_fdiv = 0;
                end
                else
                    inner_clk <= #vcoclk_period_half ~inner_clk;
            end
    end

    always @(clk_in or CLKFB or negedge rst_n)
    begin
        if(!rst_n)
        begin
            adjust <= 1'b1;
            fb_route_delay = 0.0;
            tmp_ratio  = 0;
            tmp_delay  = 0.0;
            real_delay = 0.0;
        end
        else
            if(adjust == 1'b1)
            begin
                fb_route_delay = clk_fb_first_edge - clk_in_first_edge;
                if((clkin_time > 0) && (fb_route_delay > 0))
                begin
                    tmp_ratio  = fb_route_delay / clkin_time;
                    tmp_delay  = fb_route_delay - (clkin_time * tmp_ratio);
                    real_delay = clkin_time - tmp_delay;
                    adjust <= 1'b0;
                end
            end
    end

    always @(inner_clk)
    begin
        if(EXTERNAL_FB == "CLKOUT0" || EXTERNAL_FB == "CLKOUT1" || EXTERNAL_FB == "CLKOUT2" || EXTERNAL_FB == "CLKOUT3" || EXTERNAL_FB == "CLKOUT4")
            vcoclk <= #real_delay inner_clk;
        else
            vcoclk <= inner_clk;
    end

    assign vco[0] = vcoclk;
    assign #(vcoclk_period_half/4) vco[1] = vco[0];
    assign #(vcoclk_period_half/4) vco[2] = vco[1];
    assign #(vcoclk_period_half/4) vco[3] = vco[2];
    assign #(vcoclk_period_half/4) vco[4] = vco[3];
    assign #(vcoclk_period_half/4) vco[5] = vco[4];
    assign #(vcoclk_period_half/4) vco[6] = vco[5];
    assign #(vcoclk_period_half/4) vco[7] = vco[6];
////VCO_CLK_DIV2///////////////////////////////////////
    always @(posedge vco[0] or negedge rst_n)
    begin
        if(!rst_n)
            vco_div2[0] <= 1'b0;
        else
            if(VCOCLK_DIV2)
                vco_div2[0] <= ~vco_div2[0];
            else
                vco_div2[0] <= 1'b0;
    end

    always @(posedge vco[1] or negedge rst_n)
    begin
        if(!rst_n)
            vco_div2[1] <= 1'b0;
        else
            if(VCOCLK_DIV2)
                vco_div2[1] <= ~vco_div2[1];
            else
                vco_div2[1] <= 1'b0;
    end

    always @(posedge vco[2] or negedge rst_n)
    begin
        if(!rst_n)
            vco_div2[2] <= 1'b0;
        else
            if(VCOCLK_DIV2)
                vco_div2[2] <= ~vco_div2[2];
            else
                vco_div2[2] <= 1'b0;
    end

    always @(posedge vco[3] or negedge rst_n)
    begin
        if(!rst_n)
            vco_div2[3] <= 1'b0;
        else
            if(VCOCLK_DIV2)
                vco_div2[3] <= ~vco_div2[3];
            else
                vco_div2[3] <= 1'b0;
    end

    always @(posedge vco[4] or negedge rst_n)
    begin
        if(!rst_n)
            vco_div2[4] <= 1'b0;
        else
            if(VCOCLK_DIV2)
                vco_div2[4] <= ~vco_div2[4];
            else
                vco_div2[4] <= 1'b0;
    end

    always @(posedge vco[5] or negedge rst_n)
    begin
        if(!rst_n)
            vco_div2[5] <= 1'b0;
        else
            if(VCOCLK_DIV2) 
                vco_div2[5] <= ~vco_div2[5];
            else
                vco_div2[5] <= 1'b0;
    end

    always @(posedge vco[6] or negedge rst_n)
    begin
        if(!rst_n)
            vco_div2[6] <= 1'b0;
        else 
            if(VCOCLK_DIV2)
                vco_div2[6] <= ~vco_div2[6];
            else
                vco_div2[6] <= 1'b0; 
    end

    always @(posedge vco[7] or negedge rst_n)
    begin
        if(!rst_n)
            vco_div2[7] <= 1'b0;
        else
            if(VCOCLK_DIV2) 
                vco_div2[7] <= ~vco_div2[7];
            else
                vco_div2[7] <= 1'b0;
    end

    assign clkout = (VCOCLK_DIV2 == 1'b0) ? vco : vco_div2;
///////////////////////////////////////////////////////
////PLL_LOCK///////////////////////////////////////////
    assign clk_lock = (INTERNAL_FB == "ENABLE") ? clk_in : CLKFB;
    
    always @(posedge clk_lock or negedge rstanalog_n)
    begin
        if(!rstanalog_n)
        begin
            start_clk <= 1'b0;
            cnt_clkfb <= 2'b00;
        end
        else
            if(cnt_clkfb == 3)
                start_clk = 1'b1;
            else
                cnt_clkfb = cnt_clkfb + 1;
    end

    always @(posedge clk_in or negedge rstanalog_n)
    begin
        if(!rstanalog_n)
        begin
            cnt_lock <= 11'b000_0000_0001;
            lock_reg <= 1'b0;
        end
        else
            if(clkout_lock && start_clk)
                if(cnt_lock == idivider*6)
                    lock_reg <= 1'b1;
                else
                    cnt_lock <= cnt_lock+1;
            else
            begin
                cnt_lock <= 11'b000_0000_0001;
                lock_reg <= 1'b0;
            end
    end

    assign LOCK = lock_reg & ~clkwo;
///////////////////////////////////////////////////////
////PLL_ODIV///////////////////////////////////////////
    assign phase_bonding = (SIM_DEVICE == "PGL22G") ? 1'b0 : 1'b1;

    assign rst_odiv_n = (RSTODIV_PHASE_EN == "FALSE") ? ((SIM_DEVICE == "PGL22G") ? LOCK : rst_n) : rstodiv_n;

    always @(posedge clkout[4] or negedge rst_odiv_n)
    begin
        if(!rst_odiv_n)
            rst_clk4_n <= 2'b00;
        else
            rst_clk4_n <= {rst_clk4_n[0],1'b1};
    end

    assign clk_cas[1] = (CLK_CAS1_EN == "TRUE") ? 1'b1 : 1'b0;
    assign clk_cas[2] = (CLK_CAS2_EN == "TRUE") ? 1'b1 : 1'b0;
    assign clk_cas[3] = (CLK_CAS3_EN == "TRUE") ? 1'b1 : 1'b0;
    assign clk_cas[4] = (CLK_CAS4_EN == "TRUE") ? 1'b1 : 1'b0;
    assign phase_adjust[0] = (PHASE_ADJUST0_EN == "TRUE") ? 1'b1 : 1'b0;
    assign phase_adjust[1] = (PHASE_ADJUST1_EN == "TRUE") ? 1'b1 : 1'b0;
    assign phase_adjust[2] = (PHASE_ADJUST2_EN == "TRUE") ? 1'b1 : 1'b0;
    assign phase_adjust[3] = (PHASE_ADJUST3_EN == "TRUE") ? 1'b1 : 1'b0;
    assign phase_adjust[4] = (PHASE_ADJUST4_EN == "TRUE") ? 1'b1 : 1'b0;
////ODIV0//////////////////////////////////////////////
    assign odiv0_fphase = (DYNAMIC_PHASE0_EN == "TRUE") ? PHASE0  : STATIC_PHASE0;
    assign odiv0_cphase = (DYNAMIC_PHASE0_EN == "TRUE") ? CPHASE0 : STATIC_CPHASE0;
    assign odiv0_duty   = (DYNAMIC_DUTY0_EN  == "TRUE") ? DUTY0   : STATIC_DUTY0;
    assign odiv0_duty_ctrl = (odiv0_duty[0] == 1'b1) ? (odiv0_duty + 1) >> 1 : odiv0_duty >> 1;
    assign odiv0_div1   = (divider0 == 10'b00_0000_0001) ? 1'b1 : 1'b0;
////ODIV0_FINE_PHASE///////
    always @(*)
    begin
        case(odiv0_fphase)
            3'b000: odiv0_clk_reg = clkout[0];
            3'b001: odiv0_clk_reg = clkout[1];
            3'b010: odiv0_clk_reg = clkout[2];
            3'b011: odiv0_clk_reg = clkout[3];
            3'b100: odiv0_clk_reg = clkout[4];
            3'b101: odiv0_clk_reg = clkout[5];
            3'b110: odiv0_clk_reg = clkout[6];
            3'b111: odiv0_clk_reg = clkout[7];
        endcase
    end
////ODIV0_RESET////////////
    always @(posedge clkout[0] or negedge rst_n)
    begin
        if(!rst_n)
            odiv0_rst_clk0 <= 1'b0;
        else
            odiv0_rst_clk0 <= rst_clk4_n[1];
    end

    always @(posedge odiv0_clk_reg or negedge rst_n)
    begin
        if(!rst_n)
            odiv0_rst_high <= 1'b0;
        else
            odiv0_rst_high <= odiv0_rst_clk0;
    end

    always @(posedge odiv0_clk_reg or negedge rst_n)
    begin
        if(!rst_n)
            odiv0_rst_low <= 1'b0;
        else
            odiv0_rst_low <= rst_clk4_n[1];
    end

    always @(negedge odiv0_clk_reg or negedge rst_n)
    begin
        if(!rst_n)
            odiv0_rst_sel <= 2'b00;
        else
            if((~phase_bonding & fbdiv_sel[1]) || ~phase_adjust[0])
                odiv0_rst_sel <= {odiv0_rst_sel[0],1'b1};
            else
                if(odiv0_fphase[2])
                    odiv0_rst_sel <= {odiv0_rst_sel[0],odiv0_rst_high};
                else
                    odiv0_rst_sel <= {odiv0_rst_sel[0],odiv0_rst_low};
    end
////ODIV0_COARSE_PHASE/////
    always @(posedge odiv0_clk_reg or negedge odiv0_rst_sel[1])
    begin
        if(!odiv0_rst_sel[1])
        begin
            odiv0_gate <= 1'b0;
            odiv0_cnt  <= 10'b00_0000_0000;
        end
        else
            if(odiv0_cnt == odiv0_cphase-2)
                odiv0_gate <= 1'b1;
            else
            begin
                odiv0_gate <= 1'b0;
                odiv0_cnt  <= odiv0_cnt + 1'b1;
            end
    end
////ODIV0_DIVIDER_DUTY/////
    always @(posedge odiv0_clk_reg or negedge odiv0_rst_sel[1])
    begin
        if(!odiv0_rst_sel[1])
            odiv0_counter <= 10'b00_0000_0000;
        else
            if(odiv0_gate)
                if(odiv0_counter == divider0 - 1'b1)
                    odiv0_counter <= 10'b00_0000_0000;
                else
                    odiv0_counter <= odiv0_counter + 1'b1;
            else
                odiv0_counter <= 10'b00_0000_0000;
    end

    always @(posedge odiv0_clk_reg or negedge odiv0_rst_sel[1])
    begin
        if(!odiv0_rst_sel[1])
            odiv0_clkdivr <= 1'b0;
        else
            if(odiv0_gate)
                if(odiv0_counter < odiv0_duty_ctrl)
                    odiv0_clkdivr <= 1'b1;
                else
                    odiv0_clkdivr <= 1'b0;
            else
                odiv0_clkdivr <= 1'b0;
    end

    always @(negedge odiv0_clk_reg or negedge odiv0_rst_sel[1])
    begin
        if(!odiv0_rst_sel[1])
            odiv0_set <= 1'b0;
        else
            if(odiv0_gate)
                if(odiv0_counter == odiv0_duty_ctrl)
                    odiv0_set <= odiv0_duty[0];
                else
                    odiv0_set <= 1'b0;
            else
                odiv0_set <= 1'b0;
    end

    assign clk_odivout[0] = (odiv0_div1 == 1'b1) ? odiv0_clk_reg : odiv0_clkdivr & ~odiv0_set;
////ODIV1//////////////////////////////////////////////
    assign odiv1_fphase = (DYNAMIC_PHASE1_EN == "TRUE") ? PHASE1  : STATIC_PHASE1;
    assign odiv1_cphase = (DYNAMIC_PHASE1_EN == "TRUE") ? CPHASE1 : STATIC_CPHASE1;
    assign odiv1_duty   = (DYNAMIC_DUTY1_EN  == "TRUE") ? DUTY1   : STATIC_DUTY1;
    assign odiv1_duty_ctrl = (odiv1_duty[0] == 1'b1) ? (odiv1_duty + 1) >> 1 : odiv1_duty >> 1;
    assign odiv1_div1   = (divider1 == 10'b00_0000_0001) ? 1'b1 : 1'b0;
////ODIV1_FINE_PHASE///////
    always @(*)
    begin
        if(clk_cas[1])
            odiv1_clk_reg = clk_odivout[0];
        else
            case(odiv1_fphase)
                3'b000: odiv1_clk_reg = clkout[0];
                3'b001: odiv1_clk_reg = clkout[1];
                3'b010: odiv1_clk_reg = clkout[2];
                3'b011: odiv1_clk_reg = clkout[3];
                3'b100: odiv1_clk_reg = clkout[4];
                3'b101: odiv1_clk_reg = clkout[5];
                3'b110: odiv1_clk_reg = clkout[6];
                3'b111: odiv1_clk_reg = clkout[7];
            endcase
    end
////ODIV1_RESET////////////
    always @(posedge clkout[0] or negedge rst_n)
    begin
        if(!rst_n)
            odiv1_rst_clk0 <= 1'b0;
        else
            odiv1_rst_clk0 <= rst_clk4_n[1];
    end

    always @(posedge odiv1_clk_reg or negedge rst_n)
    begin
        if(!rst_n)
            odiv1_rst_high <= 1'b0;
        else
            odiv1_rst_high <= odiv1_rst_clk0;
    end

    always @(posedge odiv1_clk_reg or negedge rst_n)
    begin
        if(!rst_n)
            odiv1_rst_low <= 1'b0;
        else
            odiv1_rst_low <= rst_clk4_n[1];
    end

    always @(negedge odiv1_clk_reg or negedge rst_n)
    begin
        if(!rst_n)
            odiv1_rst_sel <= 2'b00;
        else
            if((~phase_bonding & fbdiv_sel[2]) || ~phase_adjust[1])
                odiv1_rst_sel <= {odiv1_rst_sel[0],1'b1};
            else
                if(odiv1_fphase[2])
                    odiv1_rst_sel <= {odiv1_rst_sel[0],odiv1_rst_high};
                else
                    odiv1_rst_sel <= {odiv1_rst_sel[0],odiv1_rst_low};
    end
////ODIV1_COARSE_PHASE/////
    always @(posedge odiv1_clk_reg or negedge odiv1_rst_sel[1])
    begin
        if(!odiv1_rst_sel[1])
        begin
            odiv1_gate <= 1'b0;
            odiv1_cnt  <= 10'b00_0000_0000;
        end
        else
            if(odiv1_cnt == odiv1_cphase-2)
                odiv1_gate <= 1'b1;
            else
            begin
                odiv1_gate <= 1'b0;
                odiv1_cnt  <= odiv1_cnt + 1'b1;
            end
    end
////ODIV1_DIVIDER_DUTY/////
    always @(posedge odiv1_clk_reg or negedge odiv1_rst_sel[1])
    begin
        if(!odiv1_rst_sel[1])
            odiv1_counter <= 10'b00_0000_0000;
        else
            if(odiv1_gate)
                if(odiv1_counter == divider1 - 1'b1)
                    odiv1_counter <= 10'b00_0000_0000;
                else
                    odiv1_counter <= odiv1_counter + 1'b1;
            else
                odiv1_counter <= 10'b00_0000_0000;
    end

    always @(posedge odiv1_clk_reg or negedge odiv1_rst_sel[1])
    begin
        if(!odiv1_rst_sel[1])
            odiv1_clkdivr <= 1'b0;
        else
            if(odiv1_gate)
                if(odiv1_counter < odiv1_duty_ctrl)
                    odiv1_clkdivr <= 1'b1;
                else
                    odiv1_clkdivr <= 1'b0;
            else
                odiv1_clkdivr <= 1'b0;
    end

    always @(negedge odiv1_clk_reg or negedge odiv1_rst_sel[1])
    begin
        if(!odiv1_rst_sel[1])
            odiv1_set <= 1'b0;
        else
            if(odiv1_gate)
                if(odiv1_counter == odiv1_duty_ctrl)
                    odiv1_set <= odiv1_duty[0];
                else
                    odiv1_set <= 1'b0;
            else
                odiv1_set <= 1'b0;
    end

    assign clk_odivout[1] = (odiv1_div1 == 1) ? odiv1_clk_reg : odiv1_clkdivr & ~odiv1_set;
////ODIV2//////////////////////////////////////////////
    assign odiv2_fphase = (DYNAMIC_PHASE2_EN == "TRUE") ? PHASE2  : STATIC_PHASE2;
    assign odiv2_cphase = (DYNAMIC_PHASE2_EN == "TRUE") ? CPHASE2 : STATIC_CPHASE2;
    assign odiv2_duty   = (DYNAMIC_DUTY2_EN  == "TRUE") ? DUTY2   : STATIC_DUTY2;
    assign odiv2_duty_ctrl = (odiv2_duty[0] == 1'b1) ? (odiv2_duty + 1) >> 1 : odiv2_duty >> 1;
    assign odiv2_div1   = (divider2 == 10'b00_0000_0001) ? 1'b1 : 1'b0;
////ODIV2_FINE_PHASE///////
    always @(*)
    begin
        if(clk_cas[2])
            odiv2_clk_reg = clk_odivout[1];
        else
            case(odiv2_fphase)
                3'b000: odiv2_clk_reg = clkout[0];
                3'b001: odiv2_clk_reg = clkout[1];
                3'b010: odiv2_clk_reg = clkout[2];
                3'b011: odiv2_clk_reg = clkout[3];
                3'b100: odiv2_clk_reg = clkout[4];
                3'b101: odiv2_clk_reg = clkout[5];
                3'b110: odiv2_clk_reg = clkout[6];
                3'b111: odiv2_clk_reg = clkout[7];
            endcase
    end
////ODIV2_RESET////////////
    always @(posedge clkout[0] or negedge rst_n)
    begin
        if(!rst_n)
            odiv2_rst_clk0 <= 1'b0;
        else
            odiv2_rst_clk0 <= rst_clk4_n[1];
    end

    always @(posedge odiv2_clk_reg or negedge rst_n)
    begin
        if(!rst_n)
            odiv2_rst_high <= 1'b0;
        else
            odiv2_rst_high <= odiv2_rst_clk0;
    end

    always @(posedge odiv2_clk_reg or negedge rst_n)
    begin
        if(!rst_n)
            odiv2_rst_low <= 1'b0;
        else
            odiv2_rst_low <= rst_clk4_n[1];
    end

    always @(negedge odiv2_clk_reg or negedge rst_n)
    begin
        if(!rst_n)
            odiv2_rst_sel <= 2'b00;
        else
            if((~phase_bonding & fbdiv_sel[3]) || ~phase_adjust[2])
                odiv2_rst_sel <= {odiv2_rst_sel[0],1'b1};
            else
                if(odiv2_fphase[2])
                    odiv2_rst_sel <= {odiv2_rst_sel[0],odiv2_rst_high};
                else
                    odiv2_rst_sel <= {odiv2_rst_sel[0],odiv2_rst_low};
    end
////ODIV2_COARSE_PHASE/////
    always @(posedge odiv2_clk_reg or negedge odiv2_rst_sel[1])
    begin
        if(!odiv2_rst_sel[1])
        begin
            odiv2_gate <= 1'b0;
            odiv2_cnt  <= 10'b00_0000_0000;
        end
        else
            if(odiv2_cnt == odiv2_cphase-2)
                odiv2_gate <= 1'b1;
            else
            begin
                odiv2_gate <= 1'b0;
                odiv2_cnt  <= odiv2_cnt + 1'b1;
            end
    end
////ODIV2_DIVIDER_DUTY/////
    always @(posedge odiv2_clk_reg or negedge odiv2_rst_sel[1])
    begin
        if(!odiv2_rst_sel[1])
            odiv2_counter <= 10'b00_0000_0000;
        else
            if(odiv2_gate)
                if(odiv2_counter == divider2 - 1'b1)
                    odiv2_counter <= 10'b00_0000_0000;
                else
                    odiv2_counter <= odiv2_counter + 1'b1;
            else
                odiv2_counter <= 10'b00_0000_0000;
    end

    always @(posedge odiv2_clk_reg or negedge odiv2_rst_sel[1])
    begin
        if(!odiv2_rst_sel[1])
            odiv2_clkdivr <= 1'b0;
        else
            if(odiv2_gate)
                if(odiv2_counter < odiv2_duty_ctrl)
                    odiv2_clkdivr <= 1'b1;
                else
                    odiv2_clkdivr <= 1'b0;
            else
                odiv2_clkdivr <= 1'b0;
    end

    always @(negedge odiv2_clk_reg or negedge odiv2_rst_sel[1])
    begin
        if(!odiv2_rst_sel[1])
            odiv2_set <= 1'b0; 
        else
            if(odiv2_gate)
                if(odiv2_counter == odiv2_duty_ctrl)
                    odiv2_set <= odiv2_duty[0];
                else
                    odiv2_set <= 1'b0;
            else
                odiv2_set <= 1'b0;
    end

    assign clk_odivout[2] = (odiv2_div1 == 1) ? odiv2_clk_reg : odiv2_clkdivr & ~odiv2_set;
////ODIV3//////////////////////////////////////////////
    assign odiv3_fphase = (DYNAMIC_PHASE3_EN == "TRUE") ? PHASE3  : STATIC_PHASE3;
    assign odiv3_cphase = (DYNAMIC_PHASE3_EN == "TRUE") ? CPHASE3 : STATIC_CPHASE3;
    assign odiv3_duty   = (DYNAMIC_DUTY3_EN  == "TRUE") ? DUTY3   : STATIC_DUTY3;
    assign odiv3_duty_ctrl = (odiv3_duty[0] == 1'b1) ? (odiv3_duty + 1) >> 1 : odiv3_duty >> 1;
    assign odiv3_div1   = (divider3 == 10'b00_0000_0001) ? 1'b1 : 1'b0;
////ODIV3_FINE_PHASE///////
    always @(*)
    begin
        if(clk_cas[3])
            odiv3_clk_reg = clk_odivout[2];
        else
            case(odiv3_fphase)
                3'b000: odiv3_clk_reg = clkout[0];
                3'b001: odiv3_clk_reg = clkout[1];
                3'b010: odiv3_clk_reg = clkout[2];
                3'b011: odiv3_clk_reg = clkout[3];
                3'b100: odiv3_clk_reg = clkout[4];
                3'b101: odiv3_clk_reg = clkout[5];
                3'b110: odiv3_clk_reg = clkout[6];
                3'b111: odiv3_clk_reg = clkout[7];
            endcase
    end
////ODIV3_RESET////////////
    always @(posedge clkout[0] or negedge rst_n)
    begin
        if(!rst_n)
            odiv3_rst_clk0 <= 1'b0;
        else
            odiv3_rst_clk0 <= rst_clk4_n[1];
    end

    always @(posedge odiv3_clk_reg or negedge rst_n)
    begin
        if(!rst_n)
            odiv3_rst_high <= 1'b0;
        else
            odiv3_rst_high <= odiv3_rst_clk0;
    end

    always @(posedge odiv3_clk_reg or negedge rst_n)
    begin
        if(!rst_n)
            odiv3_rst_low <= 1'b0;
        else
            odiv3_rst_low <= rst_clk4_n[1];
    end

    always @(negedge odiv3_clk_reg or negedge rst_n)
    begin
        if(!rst_n)
            odiv3_rst_sel <= 2'b00;
        else
            if((~phase_bonding & fbdiv_sel[4]) || ~phase_adjust[3])
                odiv3_rst_sel <= {odiv3_rst_sel[0],1'b1};
            else
                if(odiv3_fphase[2])
                    odiv3_rst_sel <= {odiv3_rst_sel[0],odiv3_rst_high};
                else
                    odiv3_rst_sel <= {odiv3_rst_sel[0],odiv3_rst_low};
    end
////ODIV3_COARSE_PHASE/////
    always @(posedge odiv3_clk_reg or negedge odiv3_rst_sel[1])
    begin
        if(!odiv3_rst_sel[1])
        begin
            odiv3_gate <= 1'b0;
            odiv3_cnt  <= 10'b00_0000_0000;
        end
        else
            if(odiv3_cnt == odiv3_cphase-2)
                odiv3_gate <= 1'b1;
            else
            begin
                odiv3_gate <= 1'b0;
                odiv3_cnt  <= odiv3_cnt + 1'b1;
            end
    end
////ODIV3_DIVIDER_DUTY/////
    always @(posedge odiv3_clk_reg or negedge odiv3_rst_sel[1])
    begin
        if(!odiv3_rst_sel[1])
            odiv3_counter <= 10'b00_0000_0000;
        else
            if(odiv3_gate)
                if(odiv3_counter == divider3 - 1'b1)
                    odiv3_counter <= 10'b00_0000_0000;
                else
                    odiv3_counter <= odiv3_counter + 1'b1;
            else
                odiv3_counter <= 10'b00_0000_0000;
    end

    always @(posedge odiv3_clk_reg or negedge odiv3_rst_sel[1])
    begin
        if(!odiv3_rst_sel[1])
            odiv3_clkdivr <= 1'b0;
        else
            if(odiv3_gate)
                if(odiv3_counter < odiv3_duty_ctrl)
                    odiv3_clkdivr <= 1'b1;
                else
                    odiv3_clkdivr <= 1'b0;
            else
                odiv3_clkdivr <= 1'b0;
    end

    always @(negedge odiv3_clk_reg or negedge odiv3_rst_sel[1])
    begin
        if(!odiv3_rst_sel[1])
            odiv3_set <= 1'b0;
        else
            if(odiv3_gate)
                if(odiv3_counter == odiv3_duty_ctrl)
                    odiv3_set <= odiv3_duty[0];
                else
                    odiv3_set <= 1'b0;
            else
                odiv3_set <= 1'b0;
    end

    assign clk_odivout[3] = (odiv3_div1 == 1) ? odiv3_clk_reg : odiv3_clkdivr & ~odiv3_set;
////ODIV4//////////////////////////////////////////////
    assign odiv4_fphase = (DYNAMIC_PHASE4_EN == "TRUE") ? PHASE4  : STATIC_PHASE4;
    assign odiv4_cphase = (DYNAMIC_PHASE4_EN == "TRUE") ? CPHASE4 : STATIC_CPHASE4;
    assign odiv4_duty   = (DYNAMIC_DUTY4_EN  == "TRUE") ? DUTY4   : STATIC_DUTY4;
    assign odiv4_duty_ctrl = (odiv4_duty[0] == 1'b1) ? (odiv4_duty + 1) >> 1 : odiv4_duty >> 1;
    assign odiv4_div1   = (divider4 == 10'b00_0000_0001) ? 1'b1 : 1'b0;
////ODIV4_FINE_PHASE///////
    always @(*)
    begin
        if(clk_cas[4])
            odiv4_clk_reg = clk_odivout[3];
        else
            case(odiv4_fphase)
                3'b000: odiv4_clk_reg = clkout[0];
                3'b001: odiv4_clk_reg = clkout[1];
                3'b010: odiv4_clk_reg = clkout[2];
                3'b011: odiv4_clk_reg = clkout[3];
                3'b100: odiv4_clk_reg = clkout[4];
                3'b101: odiv4_clk_reg = clkout[5];
                3'b110: odiv4_clk_reg = clkout[6];
                3'b111: odiv4_clk_reg = clkout[7];
            endcase
    end
////ODIV4_RESET////////////
    always @(posedge clkout[0] or negedge rst_n)
    begin
        if(!rst_n)
            odiv4_rst_clk0 <= 1'b0;
        else
            odiv4_rst_clk0 <= rst_clk4_n[1];
    end

    always @(posedge odiv4_clk_reg or negedge rst_n)
    begin
        if(!rst_n)
            odiv4_rst_high <= 1'b0;
        else
            odiv4_rst_high <= odiv4_rst_clk0;
    end

    always @(posedge odiv4_clk_reg or negedge rst_n)
    begin
        if(!rst_n)
            odiv4_rst_low <= 1'b0;
        else
            odiv4_rst_low <= rst_clk4_n[1];
    end

    always @(negedge odiv4_clk_reg or negedge rst_n)
    begin
        if(!rst_n)
            odiv4_rst_sel <= 2'b00;
        else
            if((~phase_bonding & fbdiv_sel[5]) || ~phase_adjust[4])
                odiv4_rst_sel <= {odiv4_rst_sel[0],1'b1};
            else
                if(odiv4_fphase[2])
                    odiv4_rst_sel <= {odiv4_rst_sel[0],odiv4_rst_high};
                else
                    odiv4_rst_sel <= {odiv4_rst_sel[0],odiv4_rst_low};
    end
////ODIV4_COARSE_PHASE/////
    always @(posedge odiv4_clk_reg or negedge odiv4_rst_sel[1])
    begin
        if(!odiv4_rst_sel[1])
        begin
            odiv4_gate <= 1'b0;
            odiv4_cnt  <= 10'b00_0000_0000;
        end
        else
            if(odiv4_cnt == odiv4_cphase-2)
                odiv4_gate <= 1'b1;
            else
            begin
                odiv4_gate <= 1'b0;
                odiv4_cnt  <= odiv4_cnt + 1'b1;
            end
    end
////ODIV4_DIVIDER_DUTY/////
    always @(posedge odiv4_clk_reg or negedge odiv4_rst_sel[1])
    begin
        if(!odiv4_rst_sel[1])
            odiv4_counter <= 10'b00_0000_0000;
        else
            if(odiv4_gate)
                if(odiv4_counter == divider4 - 1'b1)
                    odiv4_counter <= 10'b00_0000_0000;
                else
                    odiv4_counter <= odiv4_counter + 1'b1;
            else
                odiv4_counter <= 10'b00_0000_0000;
    end

    always @(posedge odiv4_clk_reg or negedge odiv4_rst_sel[1])
    begin
        if(!odiv4_rst_sel[1])
            odiv4_clkdivr <= 1'b0;
        else
            if(odiv4_gate)
                if(odiv4_counter < odiv4_duty_ctrl)
                    odiv4_clkdivr <= 1'b1;
                else
                    odiv4_clkdivr <= 1'b0;
            else
                odiv4_clkdivr <= 1'b0;
    end

    always @(negedge odiv4_clk_reg or negedge odiv4_rst_sel[1])
    begin
        if(!odiv4_rst_sel[1])
            odiv4_set <= 1'b0; 
        else
            if(odiv4_gate)
                if(odiv4_counter == odiv4_duty_ctrl)
                    odiv4_set <= odiv4_duty[0];
                else
                    odiv4_set <= 1'b0;
            else
                odiv4_set <= 1'b0;
    end

    assign clk_odivout[4] = (odiv4_div1 == 1) ? odiv4_clk_reg : odiv4_clkdivr & ~odiv4_set;
///////////////////////////////////////////////////////
////PLL_GATE///////////////////////////////////////////
    always @(negedge clk_odivout[0])
    begin
        clk_out0_gate <= {clk_out0_gate[1:0],~CLKOUT0_SYN};
    end

    assign clkout0_gate = (CLKOUT0_SYN_EN == "TRUE") ? clk_out0_gate[2] : 1'b1;
    assign CLKOUT0      = clk_odivout[0] & clkout0_gate;

    always @(negedge clk_odivout[0])
    begin
        clk_out0_ext_gate <= {clk_out0_ext_gate[1:0],~CLKOUT0_EXT_SYN};
    end

    assign clkout0_ext_gate = (CLKOUT0_EXT_SYN_EN == "TRUE") ? clk_out0_ext_gate[2] : 1'b1;
    assign CLKOUT0_EXT      = clk_odivout[0] & clkout0_ext_gate;

    always @(negedge clk_odivout[1])
    begin
        clk_out1_gate <= {clk_out1_gate[1:0],~CLKOUT1_SYN};
    end

    assign clkout1_gate = (CLKOUT1_SYN_EN == "TRUE") ? clk_out1_gate[2] : 1'b1;
    assign CLKOUT1      = clk_odivout[1] & clkout1_gate;

    always @(negedge clk_odivout[2])
    begin
        clk_out2_gate <= {clk_out2_gate[1:0],~CLKOUT2_SYN};
    end

    assign clkout2_gate = (CLKOUT2_SYN_EN == "TRUE") ? clk_out2_gate[2] : 1'b1;
    assign CLKOUT2      = clk_odivout[2] & clkout2_gate;

    always @(negedge clk_odivout[3])
    begin
        clk_out3_gate <= {clk_out3_gate[1:0],~CLKOUT3_SYN};
    end

    assign clkout3_gate = (CLKOUT3_SYN_EN == "TRUE") ? clk_out3_gate[2] : 1'b1;
    assign CLKOUT3      = clk_odivout[3] & clkout3_gate;

    assign clkout4_sel = (CLKIN_BYPASS_EN == "TRUE") ? clk_in : clk_odivout[4];

    always @(negedge clkout4_sel)
    begin
        clk_out4_gate <= {clk_out4_gate[1:0],~CLKOUT4_SYN};
    end

    assign clkout4_gate = (CLKOUT4_SYN_EN == "TRUE") ? clk_out4_gate[2] : 1'b1;
    assign CLKOUT4      = clkout4_sel & clkout4_gate;

    always @(*)
    begin
        case(CLKOUT5_SEL)
            0: clk_out5_reg = clk_odivout[0];
            1: clk_out5_reg = clk_odivout[1];
            2: clk_out5_reg = clk_odivout[2];
            3: clk_out5_reg = clk_odivout[3];
            4: clk_out5_reg = clk_odivout[4];
            default: clk_out5_reg = clk_odivout[0];
        endcase
    end

    always @(negedge clk_out5_reg)
    begin
        clk_out5_gate <= {clk_out5_gate[1:0],~CLKOUT5_SYN};
    end

    assign clkout5_gate = (CLKOUT5_SYN_EN == "TRUE") ? clk_out5_gate[2] : 1'b1;
    assign CLKOUT5      = clk_out5_reg & clkout5_gate;
endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////

//P = MAC + (A0*(B0+C0) + A1*(B1+C1))
`timescale 1 ns / 1 ps

module INT_PREADD_MULTADDACC
#(
    parameter GRS_EN      = "FALSE", //"TRUE"; "FALSE"
    parameter SYNC_RST    = "FALSE", //"TRUE"; "FALSE"
    parameter INREG_EN    = "FALSE",  //"TRUE"; "FALSE"
    parameter PREREG_EN    = "FALSE",  //"TRUE"; "FALSE"
    parameter PIPEREG_EN   = "FALSE",//"TRUE"; "FALSE"
    parameter SIB1_EN     = "FALSE",
    parameter SIC0_EN     = "FALSE", //"TRUE"; "FALSE"  
    parameter SIC1_EN     = "FALSE", //"TRUE"; "FALSE"
    parameter ADDSUB_OP     = 0 ,
    parameter ACCUMADDSUB_OP = 0,
    parameter DYN_OP_ADDSUB  = 1,
    parameter DYN_OP_ACC     = 1,
    parameter ASIZE = 18,              //LEGAL ASIZE = 9, 18
    parameter BSIZE = 18,              //LEGAL BSIZE = 8, 18
    parameter PSIZE = 64,             // LEGAL PSIZE for 18 mode = 64 
    parameter integer PREADD_EN = 1,
    parameter [PSIZE-1:0] MASK = 'h0, //PSIZE = 64 OVERflow setting = 'h8000_0000_0000_00XX , bit width = PSIZE
    parameter DYN_ACC_INIT   = 0,   //acc init value dynamic input
    parameter [PSIZE-1:0] ACC_INIT_VALUE = 'b0, //acc init value parameter
    parameter [ASIZE-2:0] SC_PSE_A0 = 0, //SC_PSE = 0, disable PSE ,parameter bit width = ASIZE - 1 
    parameter [ASIZE-2:0] SC_PSE_A1 = 0, //SC_PSE = 0, disable PSE ,parameter bit width = ASIZE - 1
    parameter [BSIZE-2:0] SC_PSE_B0 = 0, //SC_PSE = 0, disable PSE ,parameter bit width = BSIZE - 1
    parameter [BSIZE-2:0] SC_PSE_B1 = 0, //SC_PSE = 0, disable PSE ,parameter bit width = BSIZE - 1
    parameter [BSIZE-2:0] SC_PSE_C0 = 0, //SC_PSE = 0, disable PSE ,parameter bit width = BSIZE - 1
    parameter [BSIZE-2:0] SC_PSE_C1 = 0  //SC_PSE = 0, disable PSE ,parameter bit width = BSIZE - 1
) (
    input   CE,
    input   RST,
    input   CLK,
    input   A_SIGNED,
    input   [ASIZE-1:0] A0,
    input   [ASIZE-1:0] A1,
    input   B_SIGNED,
    input   [BSIZE-1:0] B0,
    input   [BSIZE-1:0] B1,
    input   C_SIGNED,
    input   [BSIZE-1:0] C0,
    input   [BSIZE-1:0] C1,
    input   [1:0] PREADDSUB,
    input   [PSIZE-1:0] ACCUM_INIT,
    input   ADDSUB,
    input   ACCUMADDSUB,
    input   RELOAD,
    output  [PSIZE-1:0] P,
    output  reg OVER,
    output  reg UNDER,
    output  [PSIZE-1:0] R
);

initial begin
    if ((PREADD_EN != 0) && (PREADD_EN != 1))
    begin
        $finish;
    end
    case (ASIZE)
        9:  if ((BSIZE + PREADD_EN) != 9 || PSIZE != 32)
            begin
                $finish;
            end
        18: if (BSIZE != 18 || PSIZE != 64)
            begin
                $finish;
            end
        default :
            $finish;
    endcase
    //  $display ("INT_PREADD_MULTADDACC  error :illegal ASIZE or BSIZE or PSIZE");

    if ((GRS_EN != "TRUE") && (GRS_EN != "FALSE")) begin
        $display("GRS_EN error");
        $finish;
    end
    if ((SYNC_RST != "TRUE") && (SYNC_RST != "FALSE")) begin
        $display("SYNC_RST error");
        $finish;
    end

    if ((INREG_EN != "TRUE") && (INREG_EN != "FALSE")) begin
        $display("INREG_EN error");
        $finish;
    end
    if ((PREREG_EN != "TRUE") && (PREREG_EN != "FALSE")) begin
        $display("PREREG_EN error");
        $finish;
    end
    if ((PIPEREG_EN != "TRUE") && (PIPEREG_EN != "FALSE")) begin
        $display("PIPEREG_EN error");
        $finish;
    end

    if (SIB1_EN != "FALSE" || SIC0_EN != "FALSE" || SIC1_EN != "FALSE") begin
        $display("DRC error");
        $finish;
    end
end

wire [ASIZE-1:0] A0_PSE;
wire [ASIZE-1:0] A1_PSE;
wire [BSIZE-1:0] B0_PSE;
wire [BSIZE-1:0] B1_PSE;
wire [BSIZE-1:0] C0_PSE;
wire [BSIZE-1:0] C1_PSE;

reg  [ASIZE-1:0] a0_ireg, a1_ireg;
reg  [BSIZE-1:0] b0_ireg, b1_ireg;
reg  [BSIZE-1:0] c0_ireg, c1_ireg;
reg  asign_ireg, bsign_ireg, csign_ireg;
reg  addsub_ireg;
reg  [1:0] preaddsub_ireg;

wire [PSIZE-1:0] acc_init_value;
reg  [PSIZE-1:0] P1_reg_ACCUM_INIT1;
reg  P1_reg_RELOAD1;
reg  P1_reg_ACCUMADDSUB1;

wire [ASIZE-1:0] a0_in, a1_in;
wire [BSIZE-1:0] b0_in, b1_in;
wire [BSIZE-1:0] c0_in, c1_in;
wire asign_in, bsign_in, csign_in;
wire addsub_in;
wire [1:0] preaddsub_in;

wire [PSIZE-1:0] P1_reg_ACCUM_INIT_comb ;
wire P1_reg_RELOAD_comb ; 
wire P1_reg_ACCUMADDSUB_comb;     

wire [BSIZE:0] prad_b0, prad_c0, prad_sum0;
wire [BSIZE:0] prad_b1, prad_c1, prad_sum1;
wire prad_sign;
wire [BSIZE:0] b0_inmux;
wire [BSIZE:0] b1_inmux;
wire bsign_inmux;

reg  [ASIZE-1:0] a1_pareg, a0_pareg;
reg  [BSIZE:0]   b1_pareg, b0_pareg;
reg  asign_pareg, bsign_pareg;
wire [ASIZE-1:0] mult_a1, mult_a0;
wire [BSIZE:0]   mult_b1, mult_b0;
wire mult_asign, mult_bsign;

wire [PSIZE-1:0] mult_a1ext, mult_a0ext;
wire [PSIZE-1:0] mult_b1ext, mult_b0ext;
wire [PSIZE-1:0] PRODUCT0;
wire [PSIZE-1:0] PRODUCT1;

reg  [PSIZE-1:0] P2_reg_PRODUCT_0;
wire [PSIZE-1:0] P2_reg_PRODUCT_0_comb;
reg  [PSIZE-1:0] P2_reg_PRODUCT_1;
wire [PSIZE-1:0] P2_reg_PRODUCT_1_comb;
reg P2_reg_RELOAD;
wire P2_reg_RELOAD_comb;
reg P2_reg_ACCUMADDSUB;
wire P2_reg_ACCUMADDSUB_comb;
reg  P2_reg_ADDSUB;
wire P2_reg_ADDSUB_comb;
wire [PSIZE-1:0] sum;
reg  [PSIZE-1:0] DPO_reg;
wire [BSIZE-1:0]  b1_mux;
wire [BSIZE-1:0]  c0_mux;
wire [BSIZE-1:0]  c1_mux;
wire        csign_mux;
wire global_rstn, RST_sync, RST_async, rst_asyncomb;

assign global_rstn = GRS_EN == "TRUE" ? GRS_INST.GRSNET : 1'b1;
assign RST_sync = (SYNC_RST == "TRUE") ? RST : 1'b0;
assign RST_async = (SYNC_RST == "FALSE") ? RST : 1'b0;
assign rst_asyncomb = RST_async | (~global_rstn);

assign b1_mux = (SIB1_EN == "TRUE") ?  b0_in :  B1_PSE;
assign c0_mux = (SIC0_EN == "TRUE") ?  b0_in :  C0_PSE;
assign c1_mux = (SIC1_EN == "TRUE") ?  c0_in :  C1_PSE; // FIXME
assign csign_mux = (SIC0_EN == "TRUE") ?  bsign_in : C_SIGNED ;

assign acc_init_value = DYN_ACC_INIT ? ACCUM_INIT : ACC_INIT_VALUE;

INT_PSE #(.ASIZE(ASIZE),.SC_PSE(SC_PSE_A0)) U1_PSE(.A(A0), .SIGN(A_SIGNED), .A_PSE(A0_PSE));
INT_PSE #(.ASIZE(ASIZE),.SC_PSE(SC_PSE_A1)) U2_PSE(.A(A1), .SIGN(A_SIGNED), .A_PSE(A1_PSE));
INT_PSE #(.ASIZE(BSIZE),.SC_PSE(SC_PSE_B0)) U3_PSE(.A(B0), .SIGN(B_SIGNED), .A_PSE(B0_PSE));
INT_PSE #(.ASIZE(BSIZE),.SC_PSE(SC_PSE_B1)) U4_PSE(.A(B1), .SIGN(B_SIGNED), .A_PSE(B1_PSE));
INT_PSE #(.ASIZE(BSIZE),.SC_PSE(SC_PSE_C0)) U5_PSE(.A(C0), .SIGN(C_SIGNED), .A_PSE(C0_PSE));
INT_PSE #(.ASIZE(BSIZE),.SC_PSE(SC_PSE_C1)) U6_PSE(.A(C1), .SIGN(C_SIGNED), .A_PSE(C1_PSE));

initial begin
    {asign_ireg, a1_ireg, a0_ireg} = 'b0;
    {bsign_ireg, b1_ireg, b0_ireg} = 'b0;
    {csign_ireg, c1_ireg, c0_ireg} = 'b0;
      addsub_ireg = 0;
      preaddsub_ireg = 0;
      P1_reg_ACCUM_INIT1 = 0;
      P1_reg_RELOAD1     = 0;
      P1_reg_ACCUMADDSUB1 = 0;
    P2_reg_PRODUCT_0 = 0;
    P2_reg_PRODUCT_1 = 0;
    P2_reg_ADDSUB   = 0;
    DPO_reg    = 0;
end

wire addsub_op, accumaddsub;
assign addsub_op = DYN_OP_ADDSUB ? ADDSUB : ADDSUB_OP;
assign accumaddsub = DYN_OP_ACC ? ACCUMADDSUB : ACCUMADDSUB_OP;

always @(posedge CLK or posedge rst_asyncomb)
    if (rst_asyncomb || RST_sync) begin
        {asign_ireg, a1_ireg, a0_ireg} <= 'b0;
        {bsign_ireg, b1_ireg, b0_ireg} <= 'b0;
        {csign_ireg, c1_ireg, c0_ireg} <= 'b0;
      addsub_ireg <= 0;
      preaddsub_ireg <= 0;
      P1_reg_ACCUM_INIT1 <= 0;
      P1_reg_RELOAD1     <= 0;
      P1_reg_ACCUMADDSUB1 <= 0;
    end
    else if (CE) begin
        {asign_ireg, a1_ireg, a0_ireg} <= {A_SIGNED, A1_PSE, A0_PSE};
        {bsign_ireg, b1_ireg, b0_ireg} <= {B_SIGNED, b1_mux, B0_PSE};
        {csign_ireg, c1_ireg, c0_ireg} <= {csign_mux, c1_mux, c0_mux};
         addsub_ireg <= addsub_op;
         P1_reg_ACCUM_INIT1 <= acc_init_value;
         P1_reg_RELOAD1     <= RELOAD;
         P1_reg_ACCUMADDSUB1 <= accumaddsub;
         preaddsub_ireg <= PREADDSUB;
    end
   
assign {asign_in, a1_in, a0_in} = (INREG_EN == "TRUE") ? {asign_ireg, a1_ireg, a0_ireg} : {A_SIGNED, A1_PSE, A0_PSE};
assign {bsign_in, b1_in, b0_in} = (INREG_EN == "TRUE") ? {bsign_ireg, b1_ireg, b0_ireg} : {B_SIGNED, b1_mux, B0_PSE};
assign {csign_in, c1_in, c0_in} = (INREG_EN == "TRUE") ? {csign_ireg, c1_ireg, c0_ireg} : {csign_mux, c1_mux, c0_mux};
assign preaddsub_in = (INREG_EN == "TRUE") ? preaddsub_ireg : PREADDSUB; 
assign addsub_in = (INREG_EN == "TRUE") ? addsub_ireg : addsub_op;
assign P1_reg_ACCUM_INIT_comb = (INREG_EN == "TRUE") ? P1_reg_ACCUM_INIT1 : acc_init_value;
assign P1_reg_RELOAD_comb     = (INREG_EN == "TRUE") ? P1_reg_RELOAD1     : RELOAD;
assign P1_reg_ACCUMADDSUB_comb    = (INREG_EN == "TRUE") ? P1_reg_ACCUMADDSUB1 : accumaddsub;   


assign prad_b0 = {(bsign_in & b0_in[BSIZE-1]), b0_in};
assign prad_c0 = {(csign_in & c0_in[BSIZE-1]), c0_in};
assign prad_b1 = {(bsign_in & b1_in[BSIZE-1]), b1_in};
assign prad_c1 = {(csign_in & c1_in[BSIZE-1]), c1_in};
assign prad_sum0 = preaddsub_in[0] ? (prad_b0 - prad_c0) : (prad_b0 + prad_c0);
assign prad_sum1 = preaddsub_in[1] ? (prad_b1 - prad_c1) : (prad_b1 + prad_c1);
assign prad_sign = bsign_in | csign_in;

reg preadd_over_flag0;
always @(*)begin
  if(preaddsub_in[0]==1'b0 && PREADD_EN==1)begin
    if((bsign_in==1'b1 && b0_in[BSIZE-1]==1'b0 && csign_in==1'b0 && prad_sum0[BSIZE]==1'b1) || (bsign_in==1'b0 && csign_in==1'b1 && c0_in[BSIZE-1]==1'b0 && prad_sum0[BSIZE]==1'b1))begin
      preadd_over_flag0 = 1'b1;
    end
    else begin
      preadd_over_flag0 = 1'b0; 
    end
  end
  else if(preaddsub_in[0]==1'b1 && PREADD_EN==1)begin
    if((bsign_in==1'b1 && b0_in[BSIZE-1]==1'b1 && csign_in==1'b0 && prad_sum0[BSIZE]==1'b0) || (bsign_in==1'b0 && csign_in==1'b1 && c0_in[BSIZE-1]==1'b1 && prad_sum0[BSIZE]==1'b1) ||
      (bsign_in ==1'b0 && csign_in==1'b0 && (b0_in<c0_in)))begin
      preadd_over_flag0 = 1'b1;
    end
    else begin
      preadd_over_flag0 = 1'b0;
    end
  end
end

reg preadd_over_flag1;
always @(*)begin
  if(preaddsub_in[1]==1'b0 && PREADD_EN==1)begin
    if((bsign_in==1'b1 && b1_in[BSIZE-1]==1'b0 && csign_in==1'b0 && prad_sum1[BSIZE]==1'b1) || (bsign_in==1'b0 && csign_in==1'b1 && c1_in[BSIZE-1]==1'b0 && prad_sum1[BSIZE]==1'b1))begin
      preadd_over_flag1 = 1'b1;
    end
    else begin
      preadd_over_flag1 = 1'b0;
    end
  end
  else if(preaddsub_in[1]==1'b1 && PREADD_EN==1)begin
    if((bsign_in==1'b1 && b1_in[BSIZE-1]==1'b1 && csign_in==1'b0 && prad_sum1[BSIZE]==1'b0) || (bsign_in==1'b0 && csign_in==1'b1 && c1_in[BSIZE-1]==1'b1 && prad_sum1[BSIZE]==1'b1) ||
      (bsign_in ==1'b0 && csign_in==1'b0 && (b1_in<c1_in)))begin
      preadd_over_flag1 = 1'b1;
    end
    else begin
      preadd_over_flag1 = 1'b0;
    end
  end
end

always @(preadd_over_flag0 or preadd_over_flag1) begin
    if ((preadd_over_flag0==1 || preadd_over_flag1==1) && PREADD_EN==1)
    $display("Error: PREADD result is overflow!");
end

assign b0_inmux    = PREADD_EN ? prad_sum0 : {1'b0, b0_in};
assign b1_inmux    = PREADD_EN ? prad_sum1 : {1'b0, b1_in};
assign bsign_inmux = PREADD_EN ? prad_sign : bsign_in;
always @(posedge CLK or posedge rst_asyncomb)
    if (rst_asyncomb || RST_sync) begin
        {asign_pareg, a1_pareg, a0_pareg} <= 'b0;
        {bsign_pareg, b1_pareg, b0_pareg} <= 'b0;
    end
    else if (CE) begin
        {asign_pareg, a1_pareg, a0_pareg} <= {asign_in, a1_in, a0_in};
        {bsign_pareg, b1_pareg, b0_pareg} <= {bsign_inmux, b1_inmux, b0_inmux};
    end

assign {mult_asign, mult_a1, mult_a0} = (PREREG_EN == "TRUE") ? {asign_pareg, a1_pareg, a0_pareg} : {asign_in, a1_in, a0_in};
assign {mult_bsign, mult_b1, mult_b0} = (PREREG_EN == "TRUE") ? {bsign_pareg, b1_pareg, b0_pareg} : {bsign_inmux, b1_inmux, b0_inmux};

assign mult_a0ext = {{(PSIZE-ASIZE){mult_asign & mult_a0[ASIZE-1]}}, mult_a0};
assign mult_a1ext = {{(PSIZE-ASIZE){mult_asign & mult_a1[ASIZE-1]}}, mult_a1};
assign mult_b0ext = {{(PSIZE-BSIZE-PREADD_EN){mult_bsign & mult_b0[BSIZE+PREADD_EN-1]}}, mult_b0[BSIZE+PREADD_EN-1:0]};
assign mult_b1ext = {{(PSIZE-BSIZE-PREADD_EN){mult_bsign & mult_b1[BSIZE+PREADD_EN-1]}}, mult_b1[BSIZE+PREADD_EN-1:0]};

assign PRODUCT0 = mult_a0ext * mult_b0ext;
assign PRODUCT1 = mult_a1ext * mult_b1ext;

always @(posedge CLK or posedge rst_asyncomb)
   if (rst_asyncomb || RST_sync) begin
         P2_reg_PRODUCT_0 <= 0;
         P2_reg_PRODUCT_1 <= 0;
         P2_reg_ADDSUB   <= 0;
         P2_reg_ACCUMADDSUB  <= 0;
         P2_reg_RELOAD <= 0;
   end
         else if (CE) begin
            P2_reg_PRODUCT_0 <= PRODUCT0;
            P2_reg_PRODUCT_1 <= PRODUCT1;
            P2_reg_ADDSUB   <= addsub_in;
            P2_reg_ACCUMADDSUB  <= P1_reg_ACCUMADDSUB_comb;
            P2_reg_RELOAD <= P1_reg_RELOAD_comb;
   end


assign P2_reg_PRODUCT_0_comb = (PIPEREG_EN == "TRUE") ? P2_reg_PRODUCT_0 : PRODUCT0;
assign P2_reg_PRODUCT_1_comb = (PIPEREG_EN == "TRUE") ? P2_reg_PRODUCT_1 : PRODUCT1;
assign P2_reg_ADDSUB_comb   = (PIPEREG_EN == "TRUE") ? P2_reg_ADDSUB : addsub_in;
assign P2_reg_ACCUMADDSUB_comb  = (PIPEREG_EN == "TRUE") ? P2_reg_ACCUMADDSUB : P1_reg_ACCUMADDSUB_comb;
assign P2_reg_RELOAD_comb   = (PIPEREG_EN == "TRUE") ? P2_reg_RELOAD : P1_reg_RELOAD_comb; 

assign sum = (P2_reg_ADDSUB_comb ^ P2_reg_ACCUMADDSUB_comb == 0) ? (P2_reg_PRODUCT_0_comb + P2_reg_PRODUCT_1_comb) : 
                                   (P2_reg_PRODUCT_0_comb - P2_reg_PRODUCT_1_comb);

assign R = P2_reg_RELOAD_comb ? P1_reg_ACCUM_INIT_comb
                              : (P2_reg_ACCUMADDSUB_comb? DPO_reg - sum : DPO_reg + sum);


always @(posedge CLK or posedge rst_asyncomb)
    if (rst_asyncomb || RST_sync) begin
        DPO_reg <= 'b0;
    end
    else if (CE) begin
        DPO_reg <= R;
    end

assign P =  DPO_reg;

wire eqzero;
wire eqone;
reg eqzero_d;
reg eqone_d;
wire eqzero_one;
wire over;
wire under;

assign eqzero = &(~R | MASK);
assign eqone  = &( R | MASK);
assign eqzero_one = ~(eqzero|eqone);

always @ (posedge CLK or posedge rst_asyncomb)
    if (rst_asyncomb || RST_sync) begin
        eqzero_d  <= 0;
        eqone_d   <= 0;
        OVER      <= 0;
        UNDER     <= 0;
    end
    else if (CE) begin
        eqzero_d  <= eqzero;
        eqone_d   <= eqone;
        OVER      <= over;
        UNDER     <= under;
    end

assign over = eqzero_d & eqzero_one;
assign under = eqone_d & eqzero_one;

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2016 PANGO MICROSYSTEMS, INC
// ALL RIGHTS REVERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
//Library:
//FileName:
//
//Functional description:
//GTP for HSSTLP_PLL of PGL2 HSSTLP.
//Parameter description:
//
//Port description:
//
//Author:Gan Linghao
//Revision:
//  2019/08/26: Initial Version.
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1ns/1ps 
module GTP_HSSTLP_PLL
#(
    //parameter    integer    TX_SYNCK_SEL = 0,//select clk of PLL0 to tx_syncp[0], select clk of PLL1 to tx_syncp[1] 
    parameter    integer    TX_SYNCK_PD = 0,
    parameter               PMA_PLL_REG_REFCLK_TERM_IMP_CTRL = "TRUE",

    parameter    integer    PMA_PLL_REG_BG_TRIM = 2,
    parameter    integer    PMA_PLL_REG_IBUP_A1 = 262143,
    parameter    integer    PMA_PLL_REG_IBUP_A2 = 0,
    parameter    integer    PMA_PLL_REG_IBUP_PD = 0,
    parameter               PMA_PLL_REG_V2I_BIAS_SEL = "FALSE",
    parameter               PMA_PLL_REG_V2I_EN = "TRUE",
    parameter    integer    PMA_PLL_REG_V2I_TB_SEL = 0,
    parameter               PMA_PLL_REG_V2I_RCALTEST_PD = "FALSE",
    parameter    integer    PMA_PLL_REG_RES_CAL_TEST = 0,
    parameter    integer    PMA_RES_CAL_DIV = 0,//Added in 2019/9/27
    parameter               PMA_RES_CAL_CLK_SEL = "FALSE",//Added in 2019/9/27

    parameter               PMA_PLL_REG_PLL_PFDDELAY_EN = "TRUE",
    parameter    integer    PMA_PLL_REG_PFDDELAYSEL = 1,
    parameter    integer    PMA_PLL_REG_PLL_VCTRL_SET = 0,
    parameter               PMA_PLL_REG_READY_OR_LOCK = "FALSE",
    parameter    integer    PMA_PLL_REG_PLL_CP = 31,
    parameter    integer    PMA_PLL_REG_PLL_REFDIV = 16,
    parameter               PMA_PLL_REG_PLL_LOCKDET_EN = "FALSE",
    parameter               PMA_PLL_REG_PLL_READY = "FALSE",
    parameter               PMA_PLL_REG_PLL_READY_OW = "FALSE",
    parameter    integer    PMA_PLL_REG_PLL_FBDIV = 36,
    parameter    integer    PMA_PLL_REG_LPF_RES = 1,
    parameter               PMA_PLL_REG_JTAG_OE = "FALSE",
    parameter    integer    PMA_PLL_REG_JTAG_VHYSTSEL = 0,
    parameter               PMA_PLL_REG_PLL_LOCKDET_EN_OW = "FALSE",
    parameter    integer    PMA_PLL_REG_PLL_LOCKDET_FBCT = 7,
    parameter    integer    PMA_PLL_REG_PLL_LOCKDET_ITER = 3,
    parameter               PMA_PLL_REG_PLL_LOCKDET_MODE = "FALSE",
    parameter    integer    PMA_PLL_REG_PLL_LOCKDET_LOCKCT = 4,
    parameter    integer    PMA_PLL_REG_PLL_LOCKDET_REFCT = 7,
    parameter               PMA_PLL_REG_PLL_LOCKDET_RESET_N = "TRUE",
    parameter               PMA_PLL_REG_PLL_LOCKDET_RESET_N_OW = "FALSE",
    parameter               PMA_PLL_REG_PLL_LOCKED = "FALSE",
    parameter               PMA_PLL_REG_PLL_LOCKED_OW = "FALSE",
    parameter               PMA_PLL_REG_PLL_LOCKED_STICKY_CLEAR = "FALSE",
    parameter               PMA_PLL_REG_PLL_UNLOCKED = "FALSE",
    parameter    integer    PMA_PLL_REG_PLL_UNLOCKDET_ITER = 2,
    parameter               PMA_PLL_REG_PLL_UNLOCKED_OW = "FALSE",
    parameter               PMA_PLL_REG_PLL_UNLOCKED_STICKY_CLEAR = "FALSE",
    parameter    integer    PMA_PLL_REG_I_CTRL_MAX = 63,
    parameter               PMA_PLL_REG_REFCLK_TEST_EN = "FALSE",
    parameter               PMA_PLL_REG_RESCAL_EN = "FALSE",
    parameter    integer    PMA_PLL_REG_I_CTRL_MIN = 0,
    parameter               PMA_PLL_REG_RESCAL_DONE_OW = "FALSE",
    parameter               PMA_PLL_REG_RESCAL_DONE_VAL = "FALSE",
    parameter    integer    PMA_PLL_REG_RESCAL_I_CODE = 46,
    parameter               PMA_PLL_REG_RESCAL_I_CODE_OW = "FALSE",
    parameter               PMA_PLL_REG_RESCAL_I_CODE_PMA = "FALSE",
    parameter    integer    PMA_PLL_REG_RESCAL_I_CODE_VAL = 46,
    parameter               PMA_PLL_REG_RESCAL_INT_R_SMALL_OW = "FALSE",
    parameter               PMA_PLL_REG_RESCAL_INT_R_SMALL_VAL = "FALSE",
    parameter    integer    PMA_PLL_REG_RESCAL_ITER_VALID_SEL = 0,
    parameter               PMA_PLL_REG_RESCAL_RESET_N_OW = "FALSE",
    parameter               PMA_PLL_REG_RESCAL_RST_N_VAL = "FALSE",
    parameter               PMA_PLL_REG_RESCAL_WAIT_SEL = "TRUE",
    parameter               PMA_PLL_REFCLK2LANE_PD_L = "FALSE",
    parameter               PMA_PLL_REFCLK2LANE_PD_R = "FALSE",
    parameter               PMA_PLL_REG_LOCKDET_REPEAT = "FALSE",
    parameter               PMA_PLL_REG_NOFBCLK_STICKY_CLEAR = "FALSE",
    parameter               PMA_PLL_REG_NOREFCLK_STICKY_CLEAR = "FALSE",
    parameter    integer    PMA_PLL_REG_TEST_SEL = 0,
    parameter               PMA_PLL_REG_TEST_V_EN = "FALSE",
    parameter               PMA_PLL_REG_TEST_SIG_HALF_EN = "FALSE",
    parameter               PMA_PLL_REG_REFCLK_PAD_SEL = "FALSE",
    //parameter               PARM_CFG_HSST_RSTN = "TRUE",      //Only one pll could make CP_PARM_CFG_HSST_RSTN valid.
    parameter               PARM_PLL_POWERUP = "OFF"
    //parameter               PARM_PLL_RSTN = "TRUE"

)(
//////////Output/////////////////////////////////////////////////////////
    //SRB related
    output                  P_CFG_READY_PLL,
    output [7:0]            P_CFG_RDATA_PLL,
    output                  P_CFG_INT_PLL,
    output [5:0]            P_RESCAL_I_CODE_O,
    output                  P_REFCK2CORE,
    output                  P_PLL_READY,

    //CLK
    output                  PLL_CLK0,
    output                  PLL_CLK90,
    output                  PLL_CLK180,
    output                  PLL_CLK270,

    //New added
    output                  SYNC_PLL,
    output                  RATE_CHANGE_PLL,
    output                  PLL_PD_O,
    output                  PLL_RST_O,
    output                  PMA_PLL_READY_O,

    //Used
    output                  PLL_REFCLK_LANE_L,

//////////Input/////////////////////////////////////////////////////////
    //SRB related
    input                   P_CFG_RST_PLL,
    input                   P_CFG_CLK_PLL,
    input                   P_CFG_PSEL_PLL,
    input                   P_CFG_ENABLE_PLL,
    input                   P_CFG_WRITE_PLL,
    input [11:0]            P_CFG_ADDR_PLL,
    input [7:0]             P_CFG_WDATA_PLL,
    input                   P_RESCAL_RST_I,
    input [5:0]             P_RESCAL_I_CODE_I,
    input                   P_PLL_LOCKDET_RST_I,
    input                   P_PLL_REF_CLK,
    input                   P_PLL_RST, 
    input                   P_PLLPOWERDOWN,
    input                   P_LANE_SYNC,
    input                   P_RATE_CHANGE_TCLK_ON,

    //PAD related
    input                   REFCLK_CML_N,
    input                   REFCLK_CML_P,

    //New Added
    input                   TXPCLK_PLL_SELECTED

);

HSSTLP_PLL
#(
    .CP_TX_SYNCK_SEL                                      (0),
    .CP_TX_SYNCK_PD                                       (TX_SYNCK_PD),
    .CP_PMA_PLL_REG_REFCLK_TERM_IMP_CTRL                  (PMA_PLL_REG_REFCLK_TERM_IMP_CTRL),

    .CP_PMA_PLL_REG_BG_TRIM                               (PMA_PLL_REG_BG_TRIM),
    .CP_PMA_PLL_REG_IBUP_A1                               (PMA_PLL_REG_IBUP_A1),
    .CP_PMA_PLL_REG_IBUP_A2                               (PMA_PLL_REG_IBUP_A2),
    .CP_PMA_PLL_REG_IBUP_PD                               (PMA_PLL_REG_IBUP_PD),
    .CP_PMA_PLL_REG_V2I_BIAS_SEL                          (PMA_PLL_REG_V2I_BIAS_SEL),
    .CP_PMA_PLL_REG_V2I_EN                                (PMA_PLL_REG_V2I_EN),
    .CP_PMA_PLL_REG_V2I_TB_SEL                            (PMA_PLL_REG_V2I_TB_SEL),
    .CP_PMA_PLL_REG_V2I_RCALTEST_PD                       (PMA_PLL_REG_V2I_RCALTEST_PD),
    .CP_PMA_PLL_REG_RES_CAL_TEST                          (PMA_PLL_REG_RES_CAL_TEST),
    .CP_PMA_RES_CAL_DIV                                   (PMA_RES_CAL_DIV),
    .CP_PMA_RES_CAL_CLK_SEL                               (PMA_RES_CAL_CLK_SEL), 

    .CP_PMA_PLL_REG_PLL_PFDDELAY_EN                       (PMA_PLL_REG_PLL_PFDDELAY_EN),
    .CP_PMA_PLL_REG_PFDDELAYSEL                           (PMA_PLL_REG_PFDDELAYSEL),
    .CP_PMA_PLL_REG_PLL_VCTRL_SET                         (PMA_PLL_REG_PLL_VCTRL_SET),
    .CP_PMA_PLL_REG_READY_OR_LOCK                         (PMA_PLL_REG_READY_OR_LOCK),
    .CP_PMA_PLL_REG_PLL_CP                                (PMA_PLL_REG_PLL_CP),
    .CP_PMA_PLL_REG_PLL_REFDIV                            (PMA_PLL_REG_PLL_REFDIV),
    .CP_PMA_PLL_REG_PLL_LOCKDET_EN                        (PMA_PLL_REG_PLL_LOCKDET_EN),
    .CP_PMA_PLL_REG_PLL_READY                             (PMA_PLL_REG_PLL_READY),
    .CP_PMA_PLL_REG_PLL_READY_OW                          (PMA_PLL_REG_PLL_READY_OW),
    .CP_PMA_PLL_REG_PLL_FBDIV                             (PMA_PLL_REG_PLL_FBDIV),
    .CP_PMA_PLL_REG_LPF_RES                               (PMA_PLL_REG_LPF_RES),
    .CP_PMA_PLL_REG_JTAG_OE                               (PMA_PLL_REG_JTAG_OE),
    .CP_PMA_PLL_REG_JTAG_VHYSTSEL                         (PMA_PLL_REG_JTAG_VHYSTSEL),
    .CP_PMA_PLL_REG_PLL_LOCKDET_EN_OW                     (PMA_PLL_REG_PLL_LOCKDET_EN_OW),
    .CP_PMA_PLL_REG_PLL_LOCKDET_FBCT                      (PMA_PLL_REG_PLL_LOCKDET_FBCT),
    .CP_PMA_PLL_REG_PLL_LOCKDET_ITER                      (PMA_PLL_REG_PLL_LOCKDET_ITER),
    .CP_PMA_PLL_REG_PLL_LOCKDET_MODE                      (PMA_PLL_REG_PLL_LOCKDET_MODE),
    .CP_PMA_PLL_REG_PLL_LOCKDET_LOCKCT                    (PMA_PLL_REG_PLL_LOCKDET_LOCKCT),
    .CP_PMA_PLL_REG_PLL_LOCKDET_REFCT                     (PMA_PLL_REG_PLL_LOCKDET_REFCT),
    .CP_PMA_PLL_REG_PLL_LOCKDET_RESET_N                   (PMA_PLL_REG_PLL_LOCKDET_RESET_N),
    .CP_PMA_PLL_REG_PLL_LOCKDET_RESET_N_OW                (PMA_PLL_REG_PLL_LOCKDET_RESET_N_OW),
    .CP_PMA_PLL_REG_PLL_LOCKED                            (PMA_PLL_REG_PLL_LOCKED),
    .CP_PMA_PLL_REG_PLL_LOCKED_OW                         (PMA_PLL_REG_PLL_LOCKED_OW),
    .CP_PMA_PLL_REG_PLL_LOCKED_STICKY_CLEAR               (PMA_PLL_REG_PLL_LOCKED_STICKY_CLEAR),
    .CP_PMA_PLL_REG_PLL_UNLOCKED                          (PMA_PLL_REG_PLL_UNLOCKED),
    .CP_PMA_PLL_REG_PLL_UNLOCKDET_ITER                    (PMA_PLL_REG_PLL_UNLOCKDET_ITER),
    .CP_PMA_PLL_REG_PLL_UNLOCKED_OW                       (PMA_PLL_REG_PLL_UNLOCKED_OW),
    .CP_PMA_PLL_REG_PLL_UNLOCKED_STICKY_CLEAR             (PMA_PLL_REG_PLL_UNLOCKED_STICKY_CLEAR),
    .CP_PMA_PLL_REG_I_CTRL_MAX                            (PMA_PLL_REG_I_CTRL_MAX),
    .CP_PMA_PLL_REG_REFCLK_TEST_EN                        (PMA_PLL_REG_REFCLK_TEST_EN),
    .CP_PMA_PLL_REG_RESCAL_EN                             (PMA_PLL_REG_RESCAL_EN),
    .CP_PMA_PLL_REG_I_CTRL_MIN                            (PMA_PLL_REG_I_CTRL_MIN),
    .CP_PMA_PLL_REG_RESCAL_DONE_OW                        (PMA_PLL_REG_RESCAL_DONE_OW),
    .CP_PMA_PLL_REG_RESCAL_DONE_VAL                       (PMA_PLL_REG_RESCAL_DONE_VAL),
    .CP_PMA_PLL_REG_RESCAL_I_CODE                         (PMA_PLL_REG_RESCAL_I_CODE),
    .CP_PMA_PLL_REG_RESCAL_I_CODE_OW                      (PMA_PLL_REG_RESCAL_I_CODE_OW),
    .CP_PMA_PLL_REG_RESCAL_I_CODE_PMA                     (PMA_PLL_REG_RESCAL_I_CODE_PMA),
    .CP_PMA_PLL_REG_RESCAL_I_CODE_VAL                     (PMA_PLL_REG_RESCAL_I_CODE_VAL),
    .CP_PMA_PLL_REG_RESCAL_INT_R_SMALL_OW                 (PMA_PLL_REG_RESCAL_INT_R_SMALL_OW),
    .CP_PMA_PLL_REG_RESCAL_INT_R_SMALL_VAL                (PMA_PLL_REG_RESCAL_INT_R_SMALL_VAL),
    .CP_PMA_PLL_REG_RESCAL_ITER_VALID_SEL                 (PMA_PLL_REG_RESCAL_ITER_VALID_SEL),
    .CP_PMA_PLL_REG_RESCAL_RESET_N_OW                     (PMA_PLL_REG_RESCAL_RESET_N_OW),
    .CP_PMA_PLL_REG_RESCAL_RST_N_VAL                      (PMA_PLL_REG_RESCAL_RST_N_VAL),
    .CP_PMA_PLL_REG_RESCAL_WAIT_SEL                       (PMA_PLL_REG_RESCAL_WAIT_SEL),
    .CP_PMA_PLL_REFCLK2LANE_PD_L                          (PMA_PLL_REFCLK2LANE_PD_L),
    .CP_PMA_PLL_REFCLK2LANE_PD_R                          (PMA_PLL_REFCLK2LANE_PD_R),
    .CP_PMA_PLL_REG_LOCKDET_REPEAT                        (PMA_PLL_REG_LOCKDET_REPEAT),
    .CP_PMA_PLL_REG_NOFBCLK_STICKY_CLEAR                  (PMA_PLL_REG_NOFBCLK_STICKY_CLEAR),
    .CP_PMA_PLL_REG_NOREFCLK_STICKY_CLEAR                 (PMA_PLL_REG_NOREFCLK_STICKY_CLEAR),

    .CP_PMA_PLL_REG_TEST_SEL                              (PMA_PLL_REG_TEST_SEL),
    .CP_PMA_PLL_REG_TEST_V_EN                             (PMA_PLL_REG_TEST_V_EN),
    .CP_PMA_PLL_REG_TEST_SIG_HALF_EN                      (PMA_PLL_REG_TEST_SIG_HALF_EN),
    .CP_PMA_PLL_REG_REFCLK_PAD_SEL                        (PMA_PLL_REG_REFCLK_PAD_SEL),
    .CP_PARM_CFG_HSST_RSTN                                ("TRUE"), //Only one pll could make CP_PARM_CFG_HSST_RSTN valid.
    .CP_PARM_PLL_POWERUP                                  (PARM_PLL_POWERUP),
    .CP_PARM_PLL_RSTN                                     ("TRUE"),

    .CP_CFG_RSTN                                          ("TRUE"),
    .CP_GRSN_DIS                                          ("FALSE"),
    .CP_HSST_EN                                           ("TRUE")

) U0_HSSTLP_PLL (

//////////PAD/////////////////////////////////////////////////////////
    .REFCLK_CML_N                                         (REFCLK_CML_N),
    .REFCLK_CML_P                                         (REFCLK_CML_P),

//////////SRB related/////////////////////////////////////////////////////////
    //Output
    .CFG_READY_PLL                                        (P_CFG_READY_PLL),
    .CFG_RDATA_PLL                                        (P_CFG_RDATA_PLL),
    .CFG_INT_PLL                                          (P_CFG_INT_PLL),
    .RESCAL_I_CODE_O                                      (P_RESCAL_I_CODE_O),
    .REFCK2CORE                                           (P_REFCK2CORE),
    .PLL_READY                                            (P_PLL_READY),

    //Input
    .CFG_RST_PLL                                          (P_CFG_RST_PLL),
    .CFG_CLK_PLL                                          (P_CFG_CLK_PLL),
    .CFG_PSEL_PLL                                         (P_CFG_PSEL_PLL),
    .CFG_ENABLE_PLL                                       (P_CFG_ENABLE_PLL),
    .CFG_WRITE_PLL                                        (P_CFG_WRITE_PLL),
    .CFG_ADDR_PLL                                         (P_CFG_ADDR_PLL),
    .CFG_WDATA_PLL                                        (P_CFG_WDATA_PLL),
    .RESCAL_RST_I                                         (P_RESCAL_RST_I),
    .RESCAL_I_CODE_I                                      (P_RESCAL_I_CODE_I),
    .PLL_LOCKDET_RST_I                                    (P_PLL_LOCKDET_RST_I),
    .PLL_REF_CLK                                          (P_PLL_REF_CLK),
    .PLL_RST                                              (P_PLL_RST), 
    .PLLPOWERDOWN                                         (P_PLLPOWERDOWN),
    .LANE_SYNC                                            (P_LANE_SYNC),
    .RATE_CHANGE_TCLK_ON                                  (P_RATE_CHANGE_TCLK_ON),

//////////clk/////////////////////////////////////////////////////////
    .PLL_CLK0                                             (PLL_CLK0),
    .PLL_CLK90                                            (PLL_CLK90),
    .PLL_CLK180                                           (PLL_CLK180),
    .PLL_CLK270                                           (PLL_CLK270),

//////////New Added/////////////////////////////////////////////////////////
    .SYNC_PLL                                             (SYNC_PLL),//SELF-ADDED
    .TXPCLK_PLL_SELECTED                                  (TXPCLK_PLL_SELECTED),//SELF-ADDED
    .RATE_CHANGE_PLL                                      (RATE_CHANGE_PLL),//SELF-ADDED
    .PLL_PD_O                                             (PLL_PD_O),
    .PLL_RST_O                                            (PLL_RST_O),
    .PMA_PLL_READY_O                                      (PMA_PLL_READY_O),

//////////Used/////////////////////////////////////////////////////////
    .PLL_REFCLK_LANE_L                                    (PLL_REFCLK_LANE_L),

//////////DFT/////////////////////////////////////////////////////////
    .TEST_SE_N                                            (1'b1),
    .TEST_MODE_N                                          (1'b1),
    .TEST_RSTN                                            (),
    .TEST_SI                                              (),
    .TEST_SO                                              (),
    .FOR_PMA_TEST_MODE_N                                  (1'b1),
    .FOR_PMA_TEST_SE_N                                    (1'b1),
    .FOR_PMA_TEST_CLK                                     (),
    .FOR_PMA_TEST_RSTN                                    (),
    .FOR_PMA_TEST_SI                                      (),
    .FOR_PMA_TEST_SO                                      ()

);

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2015 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_FIFO9K.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//      2018/06/28: timescale defined
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps
 
module  GTP_FIFO9K
#(
    parameter GRS_EN = "TRUE",
    parameter integer DATA_WIDTH = 9,
    parameter integer DO_REG = 0,
    parameter [12:0]  ALMOST_FULL_OFFSET = 13'h0000,
    parameter [12:0]  ALMOST_EMPTY_OFFSET = 13'h0000,
    parameter integer USE_EMPTY = 0,
    parameter integer USE_FULL = 0,
    parameter SYNC_FIFO = "FALSE"
)(
    output        ALMOST_EMPTY,
    output        ALMOST_FULL,
    output        EMPTY,
    output        FULL,
    output [12:0] WCNT,
    output [12:0] RCNT,
    output [17:0] DO,
    input  [17:0] DI,
    input         WCLK,
    input         RCLK,
    input         WCE,
    input         RCE,
    input         ORCE,
    input         RST
);
    reg  [13:0]   rd_binary;
    reg  [13:0]   wr_binary;
    reg  [12:0]   wcnt;
    reg  [12:0]   rcnt;
    reg  [13:0]   wr_binary_next;
    reg  [13:0]   rd_binary_next;
    reg           empty_reg;
    reg           full_reg;
    reg            full_val;
    reg           almost_full_reg;
    reg           almost_empty_reg;
    reg           flagempty_en;
    reg           flagfull_en;
    reg           dout_reg_en;
    reg           sync_fifo;
    reg           grs_en;
    reg  [17:0]   dout;
    reg  [17:0]   dout_reg;

    wire [13:0]   wptr_next;
    wire [13:0]   rptr_next;
    reg  [13:0]   wptr_rclk;
    reg  [13:0]   rptr_wclk;
    wire [13:0]   wptr_next_gray;
    reg  [13:0]   wdata_buf;
    reg  [13:0]   wdata_buf_d1;
    reg  [13:0]   wdata_buf_d2;
    wire [13:0]   rptr_next_gray;
    reg  [13:0]   rdata_buf;
    reg  [13:0]   rdata_buf_d1;
    reg  [13:0]   rdata_buf_d2;
    wire          wclk,rclk;
    wire          wr_en,rd_en;
    wire          rstw,rstr;
    wire          full,empty;
    wire [17:0]   di_in;
    wire          almost_empty,almost_full;
    wire          global_rstn;

    reg  [(DATA_WIDTH-1):0] mem [(1<<13)-1 : 0];

initial   
begin
    case(SYNC_FIFO)
        "FALSE" : sync_fifo = 0;
        "TRUE"  : sync_fifo = 1;
        default : begin
            $display ("ERROR: GTP_FIFO9K instance %m parameter SYNC_FIFO:%s, The legal values are FALSE or TRUE.",SYNC_FIFO);
            $finish;
        end
    endcase
    
    case(USE_EMPTY)
        1'b0 : flagempty_en = 0;
        1'b1 : flagempty_en = 1;
        default : begin
            $display ("ERROR: GTP_FIFO9K instance %m parameter USE_EMPTY:%d, The legal values are 0 or 1.",USE_EMPTY);
            $finish;
        end
    endcase
    
    case(USE_FULL)
        1'b0 : flagfull_en = 0;
        1'b1 : flagfull_en = 1;
        default : begin
            $display ("ERROR: GTP_FIFO9K instance %m parameter USE_FULL:%d, The legal values are 0 or 1.",USE_FULL);
            $finish;
        end
    endcase
    
    case(DO_REG)
        1'b0 : dout_reg_en = 0;
        1'b1 : dout_reg_en = 1;
        default : begin
            $display ("ERROR: GTP_FIFO9K instance %m parameter DO_REG:%d, The legal values are 0 or 1.",DO_REG);
            $finish;
        end
    endcase

    case(GRS_EN)
        "FALSE" : grs_en = 0;
        "TRUE"  : grs_en = 1;
        default : begin
            $display ("ERROR: GTP_FIFO9K instance %m parameter GRS_EN:%s, The legal values are FALSE or TRUE.",GRS_EN);
            $finish;
        end
    endcase
    dout_reg ='b0;
end

assign orce_in = ORCE;
assign di_in = DI;
assign wclk = WCLK;
assign rclk = RCLK;
assign wr_en = WCE;
assign rd_en = RCE;
assign rstw = ~RST & global_rstn;
assign rstr = ~RST & global_rstn;
assign EMPTY = empty;
assign FULL  = full;
assign ALMOST_EMPTY = almost_empty;
assign ALMOST_FULL = almost_full;
assign WCNT = wcnt;
assign RCNT = rcnt;

always @(posedge rclk or negedge rstr )
begin
    if(rstr == 1'b0)
        dout_reg <= 'b0;
    else if(orce_in)
        dout_reg <= dout;
end    

assign DO = dout_reg_en ? dout_reg : dout;

assign global_rstn = grs_en ? GRS_INST.GRSNET : 1'b1;
//////////////////////////////////////////////////////
always @ (posedge wclk or negedge rstw )      //wr binary addr
begin
    if (rstw == 1'b0)
         wr_binary <= 0;
    else
         wr_binary <= wr_binary_next;
end

always @ (*)
begin
    if (full == 1'b0)
         wr_binary_next = wr_binary + wr_en;
    else
         wr_binary_next = wr_binary;
end

assign wptr_next = wr_binary_next;
//////////////////////////////////////////////////////////////////////////////////
always @ (*) begin
    case(DATA_WIDTH)
    1: begin
         full_val = (wr_binary_next[13:0] == {~rptr_wclk[13],rptr_wclk[12:0]});
    end
    2: begin
         full_val = (wr_binary_next[12:0] == {~rptr_wclk[12],rptr_wclk[11:0]});
    end
    4: begin
         full_val = (wr_binary_next[11:0] == {~rptr_wclk[11],rptr_wclk[10:0]});
    end
    8: begin
         full_val = (wr_binary_next[10:0] == {~rptr_wclk[10],rptr_wclk[9:0]});
    end
    9: begin
         full_val = (wr_binary_next[10:0] == {~rptr_wclk[10],rptr_wclk[9:0]});
    end
    16: begin
         full_val = (wr_binary_next[9:0] == {~rptr_wclk[9],rptr_wclk[8:0]});
    end
    18: begin
         full_val = (wr_binary_next[9:0] == {~rptr_wclk[9],rptr_wclk[8:0]});
    end
    default: begin  //default x9
         full_val = (wr_binary_next[10:0] == {~rptr_wclk[10],rptr_wclk[9:0]});
    end
    endcase
end

always @ (posedge wclk or negedge rstw) begin     //write full flag
    if (rstw == 1'b0)
         full_reg <= 1'b0;
    else
         full_reg <= full_val;
end

assign full=~flagfull_en |full_reg;

always @ (posedge wclk or negedge rstw) begin     //write almost_full flag
    if (rstw == 1'b0)
         almost_full_reg <= 1'b0;
    else
         almost_full_reg <= (wr_binary_next- rptr_wclk) >= ALMOST_FULL_OFFSET;
end

assign almost_full=~flagfull_en |almost_full_reg;
//////////////////////////////////////////////////////////////////////////////////
always @ (posedge rclk or negedge rstr) begin
    if(rstr == 1'b0)
         rd_binary <= 0;
    else
         rd_binary <= rd_binary_next;
end

always @ (*) begin
      if ((~empty) & rd_en)
         rd_binary_next = rd_binary + 1;
      else
         rd_binary_next = rd_binary;
end

assign rptr_next = rd_binary_next;

always @ (posedge rclk or negedge rstr) begin
      if (rstr == 1'b0) begin
          empty_reg <= 1'b1;
      end
      else begin
          empty_reg <= wptr_rclk == rd_binary_next;
      end
end

assign empty=~flagempty_en |empty_reg;

always @ (posedge rclk or negedge rstr) begin
      if (rstr == 1'b0) begin
          almost_empty_reg <= 1'b1;
      end
      else begin
          almost_empty_reg <= (wptr_rclk - rd_binary_next) <= ALMOST_EMPTY_OFFSET;
      end
end

assign almost_empty=~flagempty_en |almost_empty_reg;
//////////////////////////////////////////////////////////////////////////////////
always @ (wr_binary) begin
    case(DATA_WIDTH)
         1:     wcnt <= wr_binary[12:0];
         2:     wcnt <= {wr_binary[11:0],1'b1};
         4:     wcnt <= {wr_binary[10:0],2'b11};
         8:     wcnt <= {wr_binary[9:0],3'b111};
         9:     wcnt <= {wr_binary[9:0],3'b111};
         16:    wcnt <= {wr_binary[8:0],4'b1111};
         18:    wcnt <= {wr_binary[8:0],4'b1111};
         default:
                wcnt <= 13'b0;
    endcase
end

always @ (rd_binary) begin
    case(DATA_WIDTH)
         1:     rcnt <=  rd_binary[12:0];
         2:     rcnt <= {rd_binary[11:0],1'b1};
         4:     rcnt <= {rd_binary[10:0],2'b11};
         8:     rcnt <= {rd_binary[9:0],3'b111};
         9:     rcnt <= {rd_binary[9:0],3'b111};
         16:    rcnt <= {rd_binary[8:0],4'b1111};
         18:    rcnt <= {rd_binary[8:0],4'b1111};
         default:
                rcnt <= 13'b0;
    endcase
end
//////////////////////////////////////////////////////////////////////////////////
assign wptr_next_gray = (wptr_next>>1)^wptr_next;
assign rptr_next_gray = (rptr_next>>1)^rptr_next;

always @(posedge wclk or negedge rstw)
begin
    if(rstw == 1'b0)
    begin 
        wdata_buf <= 0;
        rdata_buf_d1 <= 0;
        rdata_buf_d2 <= 0;
    end else begin
        wdata_buf <= wptr_next_gray;
        rdata_buf_d1 <= rdata_buf;
        if(sync_fifo)
            rdata_buf_d2 <= rptr_next_gray;
        else
            rdata_buf_d2 <= rdata_buf_d1;
    end
end

always @(posedge rclk or negedge rstr)
begin
    if(rstr == 1'b0)
    begin
        wdata_buf_d1 <= 0;
        wdata_buf_d2 <= 0;
        rdata_buf <= 0;
    end else begin
        wdata_buf_d1 <= wdata_buf;
        rdata_buf <= rptr_next_gray;
        if(sync_fifo)
            wdata_buf_d2 <= wptr_next_gray;
        else
            wdata_buf_d2 <= wdata_buf_d1;
    end
end

integer i,j,k;

always @(wdata_buf_d2) begin
   for (i=0; i< 14;i=i+1)
       wptr_rclk[i] = ^(wdata_buf_d2>>i);
end

always @(rdata_buf_d2) begin
   for (j=0; j< 14;j=j+1)
       rptr_wclk[j] = ^(rdata_buf_d2>>j);
end
//////////////////////////////////////////////////////////////////////////////////
initial
begin
    for(k=0;k<(1<<13);k=k+1)
        mem[k] <= {DATA_WIDTH{1'b0}};
end

always @(posedge rclk or negedge rstr)
begin
    if(rstr == 1'b0)
        dout <= 'b0;
    else if(rd_en)
        dout <= mem[rcnt];
end
always @(posedge wclk)
begin
    if(wr_en && !full)
        mem[wcnt] <= di_in;
end
//////////////////////////////////////////////////////////////////////////////////
endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_POWERCTL.v
//
// Functional description: Power Control Circuit
//
// Parameter description:
//      
//
// Port description:
//      
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps
module GTP_POWERCTL
(
input         CLK,
input         STDBY_EN_N,
input         TIMER_EN_N,
input         CLR_N,
output        STOP,
output        STDBY,
output        STDBY_FLG
);


powerctl_gtp_wrap powerctl_gtp_wrap (
.clk(CLK),
.stdby_en_n(STDBY_EN_N),
.timer_en_n(TIMER_EN_N),
.clr_n(CLR_N),
.stdby_flg(STDBY_FLG),
.stop(STOP),
.stdby(STDBY)
);

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_IOBUFDS.v
//
// Functional description: Differential Signaling Input/Output Buffer
//
// Parameter description:
//
// Port description:
//
// Revision:
//    06/18/14 - Initial version.
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_IOBUFDS #(
    parameter IOSTANDARD = "DEFAULT",
    parameter TERM_DIFF = "ON"
)(
    output reg O,
    inout IO,
    inout IOB,
    input I,
    input T
) /* synthesis syn_black_box */ ;
  
  initial begin
    case (IOSTANDARD)
    "LVDS", "MINI-LVDS", "SUB-LVDS", "TMDS", "DEFAULT" :;
    default : begin
           $display("Attribute Syntax Error : The attribute IOSTANDARD on GTP_IOBUFDS instance %m is set to %s.", IOSTANDARD);
           $finish;
              end
    endcase

    case (TERM_DIFF)
    "ON", "OFF" :;
    default : begin
           $display("Attribute Syntax Error : The attribute TERM_DIFF on GTP_IOBUFDS instance %m is set to %s.", TERM_DIFF);
           $finish;
              end
    endcase
    end


    bufif0 (IO, I, T);
    notif0 (IOB, I, T);

    always @(*)
    begin
        if (IO == 1'b1 && IOB == 1'b0)
            O = IO;
        else if (IO == 1'b0 && IOB == 1'b1)
            O = IO;
        else
            O = 1'bx;
    end

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_UDID.v
//
// Functional description: udid Logic Control Circuit
//
// Parameter description:
//      
//
// Port description:
//      
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////


`timescale 1 ns / 1 ps
module GTP_UDID 
#(
parameter               UDID_WIDTH = 64,
parameter   [95 : 0]    UDID_CODE = 96'd0
)
(
//input         RST_N,
input         DI,
output  reg   DO,
input         LOAD,
input         SE,
input         CLK
);
reg  [UDID_WIDTH - 1 : 0]    shiftr;

always @(posedge CLK )
    begin
        if(LOAD)begin
            shiftr <= UDID_CODE[UDID_WIDTH - 1 : 0];
            DO <= 1'b1;
        end
        else if(SE)begin
            DO  <= shiftr[UDID_WIDTH - 1];
            shiftr <= {shiftr[UDID_WIDTH - 2 : 0], DI};
        end
    end


endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2016 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Filename: GTP_PCIE_E1
// Date:  2019-08-08
// Author: ccmi
// Revision: v1.0
//////////////////////////////////////////////////////////////////////////////
`timescale 1ns/10ps                                                                           
                                                                                               
module GTP_PCIEGEN2                                                                             
#(                                                                                             
// PARAMETER  PART BEGINS //////////////////////////////////////////////////////////////////// 
// PARAMETER  PART BEGINS //////////////////////////////////////////////////////////////////// 
// PARAMETER  PART BEGINS //////////////////////////////////////////////////////////////////// 
                                                                                               
                                                                                               
parameter                   GRS_EN               = "TRUE",      // FALSE, TRUE
parameter                   PIN_MUX_INT_FORCE_EN = "FALSE",      // FALSE, TRUE
parameter                   PIN_MUX_INT_DISABLE  = "FALSE",      // FALSE, TURE
parameter                   DIAG_CTRL_BUS_B2     = "NORMAL",     // "NORMAL" "FAST_LINK_MODE"
parameter                   DYN_DEBUG_SEL_EN     = "FALSE",      // FALSE, TRUE
parameter    integer        DEBUG_INFO_SEL       = 0,            // set debug_info_mux, 0-15
parameter    integer        BAR_RESIZABLE        = 21,           // 0: no resizable bar, 1: bar0 resizable, 2: bar1 resizable, 3: bar0-1 resizable, ... 56: bar3-bar5 resizable;  Please do not set more than 3 resizable bars at the same   time  Default value is 21 which is 6'b010101
parameter    integer        NUM_OF_RBARS         = 3,            // 0: no resizable bar, 1: one resizable bar, 2: two resizable bars, 3: three resizable bars  Default value is 3
parameter    integer        BAR_INDEX_0          = 0,            // set bar index0 in resizable bar control register,   0: bar0 resizable 1: bar1 resizable 2: bar2 resizable ... 5: bar5 resizable  Default value is 0
parameter    integer        BAR_INDEX_1          = 2,            // set bar index1 in resizable bar control register,   0: bar0 resizable 1: bar1 resizable 2: bar2 resizable ... 5: bar5 resizable  Default value is 2
parameter    integer        BAR_INDEX_2          = 4,            // set bar index2 in resizable bar control register,   0: bar0 resizable 1: bar1 resizable 2: bar2 resizable ... 5: bar5 resizable  Default value is 4
parameter                   TPH_DISABLE          = "FALSE",      // FALSE, TRUE
parameter                   MSIX_CAP_DISABLE     = "FALSE",      // FALSE, TRUE
parameter                   MSI_CAP_DISABLE      = "FALSE",      // FALSE, TRUE
parameter                   MSI_PVM_DISABLE      = "FALSE",      // FALSE, TRUE
parameter    integer        BAR_MASK_WRITABLE    = 32,           // 0: no writable bar, 1: bar0 writable, 2: bar1 writable, 3: bar3 writable, ... 63: bar0-5 writable
parameter    integer        APP_DEV_NUM          = 0,            // set device_number
parameter    integer        APP_BUS_NUM          = 0,            // set bus_number
parameter                   RAM_MUX_EN           = "FALSE",      // FALSE, TRUE
parameter                   ATOMIC_DISABLE       = "FALSE"       // FALSE, TRUE

)(
///////////////////////////
/////PORT DECLARATIONS/////
///////////////////////////
//clk & rst
input               MEM_CLK,
input               PCLK,  
input               PCLK_DIV2, 
//output              MUXD_AUX_CLK_OUT,              
input               BUTTON_RST,
input               POWER_UP_RST,
input               PERST,
//input               GLOGEN,
//input               GRS_N,
output              CORE_RST_N,
output              TRAINING_RST_N,
input               APP_INIT_RST,
output              PHY_RST_N,
//system control
input   [2:0]       DEVICE_TYPE,
input               RX_LANE_FLIP_EN,
input               TX_LANE_FLIP_EN,
input               APP_LTSSM_EN,
output              SMLH_LINK_UP,
output              RDLH_LINK_UP,
input               APP_REQ_RETRY_EN,
output  [4:0]       SMLH_LTSSM_STATE,

//**********************************************************************
//AXIS master interface
output              AXIS_MASTER_TVALID,
input               AXIS_MASTER_TREADY,
output  [127:0]     AXIS_MASTER_TDATA,
output  [3:0]       AXIS_MASTER_TKEEP,
output              AXIS_MASTER_TLAST,
output  [7:0]       AXIS_MASTER_TUSER,
input   [2:0]       TRGT1_RADM_PKT_HALT,
output  [5:0]       RADM_GRANT_TLP_TYPE,
//**********************************************************************
//axis slave 0 interface
output              AXIS_SLAVE0_TREADY,
input               AXIS_SLAVE0_TVALID,
input   [127:0]     AXIS_SLAVE0_TDATA,
input               AXIS_SLAVE0_TLAST,
input               AXIS_SLAVE0_TUSER,

//axis slave 1 interface
output              AXIS_SLAVE1_TREADY,
input               AXIS_SLAVE1_TVALID,
input   [127:0]     AXIS_SLAVE1_TDATA,
input               AXIS_SLAVE1_TLAST,
input               AXIS_SLAVE1_TUSER,

//axis slave 2 interface
output              AXIS_SLAVE2_TREADY,
input               AXIS_SLAVE2_TVALID,
input   [127:0]     AXIS_SLAVE2_TDATA,
input               AXIS_SLAVE2_TLAST,
input               AXIS_SLAVE2_TUSER,
output              PM_XTLH_BLOCK_TLP,      
//**********************************************************************
// DBI interface
input   [31:0]      DBI_ADDR,        
input   [31:0]      DBI_DIN,
input               DBI_CS,
input               DBI_CS2,
input   [3:0]       DBI_WR,
input               APP_DBI_RO_WR_DISABLE,
output              LBC_DBI_ACK,
output  [31:0]      LBC_DBI_DOUT,
// ELBI to SEIO interface
output              SEDO,
output              SEDO_EN,
input               SEDI,
input               SEDI_ACK,
//**********************************************************************
//legacy interrupt
output              CFG_INT_DISABLE, 
input               SYS_INT,
output              INTA_GRT_MUX,
output              INTB_GRT_MUX,
output              INTC_GRT_MUX,
output              INTD_GRT_MUX,

//msi
input               VEN_MSI_REQ,
input   [2:0]       VEN_MSI_TC,
input   [4:0]       VEN_MSI_VECTOR,
output              VEN_MSI_GRANT,
input   [31:0]      CFG_MSI_PENDING,
output              CFG_MSI_EN,

// MSI-X interface
input   [63:0]      MSIX_ADDR,
input   [31:0]      MSIX_DATA,
output              CFG_MSIX_EN,
output              CFG_MSIX_FUNC_MASK,
//**********************************************************************   
//power management
output              RADM_PM_TURNOFF,
output              RADM_MSG_UNLOCK,
input               OUTBAND_PWRUP_CMD,
output              PM_STATUS,
output  [2:0]       PM_DSTATE,
output              AUX_PM_EN,
output              PM_PME_EN,
output              PM_LINKST_IN_L0S,
output              PM_LINKST_IN_L1,
output              PM_LINKST_IN_L2,
output              PM_LINKST_L2_EXIT,
input               APP_REQ_ENTR_L1,
input               APP_READY_ENTR_L23,
input               APP_REQ_EXIT_L1,
input               APP_XFER_PENDING,
output              WAKE,
output              RADM_PM_PME,
output              RADM_PM_TO_ACK,
input               APPS_PM_XMT_TURNOFF,
input               APP_UNLOCK_MSG,
input               APPS_PM_XMT_PME,
input               APP_CLK_PM_EN,
output  [4:0]       PM_MASTER_STATE,
output  [4:0]       PM_SLAVE_STATE,
input               SYS_AUX_PWR_DET,
//**********************************************************************
//error handling
input               APP_HDR_VALID,
input   [127:0]     APP_HDR_LOG,
input   [12:0]      APP_ERR_BUS,
input               APP_ERR_ADVISORY,
output              CFG_SEND_COR_ERR_MUX,
output              CFG_SEND_NF_ERR_MUX, 
output              CFG_SEND_F_ERR_MUX,  
output              CFG_SYS_ERR_RC,
output              CFG_AER_RC_ERR_MUX,

//radm timeout
output              RADM_CPL_TIMEOUT,
output  [2:0]       RADM_TIMEOUT_CPL_TC,
output  [7:0]       RADM_TIMEOUT_CPL_TAG,
output  [1:0]       RADM_TIMEOUT_CPL_ATTR,
output  [10:0]      RADM_TIMEOUT_CPL_LEN,

//**********************************************************************
//configuration signals
output  [2:0]       CFG_MAX_RD_REQ_SIZE,
output              CFG_BUS_MASTER_EN,
output  [2:0]       CFG_MAX_PAYLOAD_SIZE,
output              CFG_RCB,
output              CFG_MEM_SPACE_EN,
output              CFG_PM_NO_SOFT_RST,
output              CFG_CRS_SW_VIS_EN,
output              CFG_NO_SNOOP_EN,
output              CFG_RELAX_ORDER_EN,
output  [1:0]       CFG_TPH_REQ_EN,
output  [2:0]       CFG_PF_TPH_ST_MODE,
output  [7:0]       CFG_PBUS_NUM,
output  [4:0]       CFG_PBUS_DEV_NUM,
output              RBAR_CTRL_UPDATE,
output              CFG_ATOMIC_REQ_EN,
output              CFG_ATOMIC_EGRESS_BLOCK,
output              CFG_EXT_TAG_EN,
//**********************************************************************
//debug signals
output              RADM_IDLE,
output              RADM_Q_NOT_EMPTY,
output              RADM_QOVERFLOW,
input   [1:0]       DIAG_CTRL_BUS,
input   [3:0]       DYN_DEBUG_INFO_SEL,
output              CFG_LINK_AUTO_BW_MUX,  
output              CFG_BW_MGT_MUX,        
output              CFG_PME_MUX,           
//output              CFG_HP_MUX,
output  [132:0]     DEBUG_INFO_MUX,
input               APP_RAS_DES_SD_HOLD_LTSSM,
input   [1:0]       APP_RAS_DES_TBA_CTRL,
//**********************************************************************
//misc
output              CFG_IDO_REQ_EN,
output              CFG_IDO_CPL_EN,
output  [7:0]       XADM_PH_CDTS,
output  [11:0]      XADM_PD_CDTS,
output  [7:0]       XADM_NPH_CDTS,
output  [11:0]      XADM_NPD_CDTS,
output  [7:0]       XADM_CPLH_CDTS,
output  [11:0]      XADM_CPLD_CDTS,
//**********************************************************************
// PIPE interface
output  [1:0]       MAC_PHY_POWERDOWN,
input   [3:0]       PHY_MAC_RXELECIDLE,
input   [3:0]       PHY_MAC_PHYSTATUS,
input   [127:0]     PHY_MAC_RXDATA,
input   [15:0]      PHY_MAC_RXDATAK,
input   [3:0]       PHY_MAC_RXVALID,
input   [11:0]      PHY_MAC_RXSTATUS,
output  [127:0]     MAC_PHY_TXDATA,
output  [15:0]      MAC_PHY_TXDATAK,
output  [3:0]       MAC_PHY_TXDETECTRX_LOOPBACK,
output  [3:0]       MAC_PHY_TXELECIDLE_L,
output  [3:0]       MAC_PHY_TXELECIDLE_H,
output  [3:0]       MAC_PHY_TXCOMPLIANCE,
output  [3:0]       MAC_PHY_RXPOLARITY,
output              MAC_PHY_RATE,
output  [1:0]       MAC_PHY_TXDEEMPH,
output  [2:0]       MAC_PHY_TXMARGIN,
output              MAC_PHY_TXSWING,
output              CFG_HW_AUTO_SP_DIS, 


input   [65:0]      P_DATAQ_DATAOUT,
output  [9:0]       P_DATAQ_ADDRA,
output  [9:0]       P_DATAQ_ADDRB,
output  [65:0]      P_DATAQ_DATAIN,
output              P_DATAQ_ENA,
output              P_DATAQ_ENB,
output              P_DATAQ_WEA,

output  [10:0]      XDLH_RETRYRAM_ADDR,
output  [67:0]      XDLH_RETRYRAM_DATA,
output              XDLH_RETRYRAM_WE,
output              XDLH_RETRYRAM_EN,
input   [67:0]      RETRYRAM_XDLH_DATA,

output  [8:0]       P_HDRQ_ADDRA,
output  [8:0]       P_HDRQ_ADDRB,
output  [137:0]     P_HDRQ_DATAIN,
output              P_HDRQ_ENA,
output              P_HDRQ_ENB,
output              P_HDRQ_WEA,
input   [137:0]     P_HDRQ_DATAOUT,

input               RAM_TEST_EN,
input               RAM_TEST_ADDRH,
input               RETRY_TEST_DATA_EN,
input               RAM_TEST_MODE_N
);

//wire grs;
//assign grs = (GRS_EN == "TRUE") ? !GRS_INST.GRSNET : 1'b0;
//assign grs = 1'b1;

PCIE
#(
   .CP_PCIE_HARD_EN                          ("TRUE"      ),                                         
   .CP_GRS_EN                                (GRS_EN      ),                                          
   .CP_PIN_MUX_INT_FORCE_EN                  (PIN_MUX_INT_FORCE_EN),                                          
   .CP_PIN_MUX_INT_DISABLE                   (PIN_MUX_INT_DISABLE),                                          
   .CP_DIAG_CTRL_BUS_B2                      (DIAG_CTRL_BUS_B2),                                          
   .CP_DYN_DEBUG_SEL_EN                      (DYN_DEBUG_SEL_EN),                                          
   .CP_DEBUG_INFO_SEL                        (DEBUG_INFO_SEL),                                          
   .CP_BAR_RESIZABLE                         (BAR_RESIZABLE),                                          
   .CP_NUM_OF_RBARS                          (NUM_OF_RBARS),                                          
   .CP_BAR_INDEX_0                           (BAR_INDEX_0),                                          
   .CP_BAR_INDEX_1                           (BAR_INDEX_1),                                          
   .CP_BAR_INDEX_2                           (BAR_INDEX_2),                                          
   .CP_TPH_DISABLE                           (TPH_DISABLE),                                          
   .CP_MSIX_CAP_DISABLE                      (MSIX_CAP_DISABLE),                                          
   .CP_MSI_CAP_DISABLE                       (MSI_CAP_DISABLE),                                          
   .CP_MSI_PVM_DISABLE                       (MSI_PVM_DISABLE),                                          
   .CP_BAR_MASK_WRITABLE                     (BAR_MASK_WRITABLE),                                          
   .CP_APP_DEV_NUM                           (APP_DEV_NUM),                                          
   .CP_APP_BUS_NUM                           (APP_BUS_NUM),                                          
   .CP_RAM_MUX_EN                            (RAM_MUX_EN),
   .CP_ATOMIC_DISABLE                        (ATOMIC_DISABLE)
)
gtp_pcie_wrap
(                                                                                                                                                                          
   .MEM_CLK                                  (MEM_CLK),
   .PCLK                                     (PCLK),
   .PCLK_DIV2                                (PCLK_DIV2),             
// .MUXD_AUX_CLK_OUT                         (MUXD_AUX_CLK_OUT),                                          
   .BUTTON_RST                               (BUTTON_RST),                                          
   .POWER_UP_RST                             (POWER_UP_RST),                                          
   .PERST                                    (PERST), 
   .CORE_RST_N                               (CORE_RST_N),                                          
   .TRAINING_RST_N                           (TRAINING_RST_N),                                          
   .APP_INIT_RST                             (APP_INIT_RST),                                          
   .PHY_RST_N                                (PHY_RST_N),                                          
                                                                                      
   .DEVICE_TYPE                              (DEVICE_TYPE),                                          
   .RX_LANE_FLIP_EN                          (RX_LANE_FLIP_EN),                                          
   .TX_LANE_FLIP_EN                          (TX_LANE_FLIP_EN),                                          
   .APP_LTSSM_EN                             (APP_LTSSM_EN),                                          
   .SMLH_LINK_UP                             (SMLH_LINK_UP),                                          
   .RDLH_LINK_UP                             (RDLH_LINK_UP),                                          
   .APP_REQ_RETRY_EN                         (APP_REQ_RETRY_EN),                                          
   .SMLH_LTSSM_STATE                         (SMLH_LTSSM_STATE),                                          
                                                                                       
                                   
                                                                                    
   .AXIS_MASTER_TVALID                       (AXIS_MASTER_TVALID),                                          
   .AXIS_MASTER_TREADY                       (AXIS_MASTER_TREADY),                                          
   .AXIS_MASTER_TDATA                        (AXIS_MASTER_TDATA),                                          
   .AXIS_MASTER_TKEEP                        (AXIS_MASTER_TKEEP),                                          
   .AXIS_MASTER_TLAST                        (AXIS_MASTER_TLAST),                                          
   .AXIS_MASTER_TUSER                        (AXIS_MASTER_TUSER),                                                                                                                                 
   .TRGT1_RADM_PKT_HALT                      (TRGT1_RADM_PKT_HALT),                                          
   .RADM_GRANT_TLP_TYPE                      (RADM_GRANT_TLP_TYPE),                                          
                                   
                                                                                   
   .AXIS_SLAVE0_TREADY                       (AXIS_SLAVE0_TREADY),                                          
   .AXIS_SLAVE0_TVALID                       (AXIS_SLAVE0_TVALID),                                          
   .AXIS_SLAVE0_TDATA                        (AXIS_SLAVE0_TDATA),                                          
   .AXIS_SLAVE0_TLAST                        (AXIS_SLAVE0_TLAST),                                          
   .AXIS_SLAVE0_TUSER                        (AXIS_SLAVE0_TUSER),                                          
                                                                                       
                                                                                   
   .AXIS_SLAVE1_TREADY                       (AXIS_SLAVE1_TREADY),                                          
   .AXIS_SLAVE1_TVALID                       (AXIS_SLAVE1_TVALID),                                          
   .AXIS_SLAVE1_TDATA                        (AXIS_SLAVE1_TDATA),                                          
   .AXIS_SLAVE1_TLAST                        (AXIS_SLAVE1_TLAST),                                          
   .AXIS_SLAVE1_TUSER                        (AXIS_SLAVE1_TUSER),                                          
                                                                                       
                                                                                   
   .AXIS_SLAVE2_TREADY                       (AXIS_SLAVE2_TREADY),                                          
   .AXIS_SLAVE2_TVALID                       (AXIS_SLAVE2_TVALID),                                          
   .AXIS_SLAVE2_TDATA                        (AXIS_SLAVE2_TDATA),                                          
   .AXIS_SLAVE2_TLAST                        (AXIS_SLAVE2_TLAST),                                          
   .AXIS_SLAVE2_TUSER                        (AXIS_SLAVE2_TUSER),                                                                                                                                 
   .PM_XTLH_BLOCK_TLP                        (PM_XTLH_BLOCK_TLP),        
                                   
                                                                                       
   .DBI_ADDR                                 (DBI_ADDR),                           
   .DBI_DIN                                  (DBI_DIN),                                          
   .DBI_CS                                   (DBI_CS),                                          
   .DBI_CS2                                  (DBI_CS2),                                          
   .DBI_WR                                   (DBI_WR),                                          
   .APP_DBI_RO_WR_DISABLE                    (APP_DBI_RO_WR_DISABLE),                                          
   .LBC_DBI_ACK                              (LBC_DBI_ACK),                                          
   .LBC_DBI_DOUT                             (LBC_DBI_DOUT),                                          
                                                                                 
   .SEDO                                     (SEDO),                                          
   .SEDO_EN                                  (SEDO_EN),                                          
   .SEDI                                     (SEDI),                                          
   .SEDI_ACK                                 (SEDI_ACK),                                          
                                   
                                                                                       
   .CFG_INT_DISABLE                          (CFG_INT_DISABLE),                                          
   .SYS_INT                                  (SYS_INT),                                          
   .INTA_GRT_MUX                             (INTA_GRT_MUX),                                          
   .INTB_GRT_MUX                             (INTB_GRT_MUX),                                          
   .INTC_GRT_MUX                             (INTC_GRT_MUX),                                          
   .INTD_GRT_MUX                             (INTD_GRT_MUX),                                          
                                                                                       
                                                                                       
   .VEN_MSI_REQ                              (VEN_MSI_REQ),                                      
   .VEN_MSI_TC                               (VEN_MSI_TC),                                      
   .VEN_MSI_VECTOR                           (VEN_MSI_VECTOR),                                      
   .VEN_MSI_GRANT                            (VEN_MSI_GRANT),                                      
   .CFG_MSI_PENDING                          (CFG_MSI_PENDING),                                      
   .CFG_MSI_EN                               (CFG_MSI_EN),                                      
                                                                                       
                                                                                       
   .MSIX_ADDR                                (MSIX_ADDR),                                          
   .MSIX_DATA                                (MSIX_DATA),                                          
   .CFG_MSIX_EN                              (CFG_MSIX_EN),                                          
   .CFG_MSIX_FUNC_MASK                       (CFG_MSIX_FUNC_MASK),                                          
                                  
                                                                                       
   .RADM_PM_TURNOFF                          (RADM_PM_TURNOFF),                                          
   .RADM_MSG_UNLOCK                          (RADM_MSG_UNLOCK),                                          
   .OUTBAND_PWRUP_CMD                        (OUTBAND_PWRUP_CMD),                                          
   .PM_STATUS                                (PM_STATUS),                                          
   .PM_DSTATE                                (PM_DSTATE),                                          
   .AUX_PM_EN                                (AUX_PM_EN),                                          
   .PM_PME_EN                                (PM_PME_EN),                                          
   .PM_LINKST_IN_L0S                         (PM_LINKST_IN_L0S),                                          
   .PM_LINKST_IN_L1                          (PM_LINKST_IN_L1),                                          
   .PM_LINKST_IN_L2                          (PM_LINKST_IN_L2),                                          
   .PM_LINKST_L2_EXIT                        (PM_LINKST_L2_EXIT),                                          
   .APP_REQ_ENTR_L1                          (APP_REQ_ENTR_L1),                                          
   .APP_READY_ENTR_L23                       (APP_READY_ENTR_L23),                                          
   .APP_REQ_EXIT_L1                          (APP_REQ_EXIT_L1),                                          
   .APP_XFER_PENDING                         (APP_XFER_PENDING),                                          
   .WAKE                                     (WAKE),                                          
   .RADM_PM_PME                              (RADM_PM_PME),                                          
   .RADM_PM_TO_ACK                           (RADM_PM_TO_ACK),                                          
   .APPS_PM_XMT_TURNOFF                      (APPS_PM_XMT_TURNOFF),                                          
   .APP_UNLOCK_MSG                           (APP_UNLOCK_MSG),                                          
   .APPS_PM_XMT_PME                          (APPS_PM_XMT_PME),                                          
   .APP_CLK_PM_EN                            (APP_CLK_PM_EN),                                          
   .PM_MASTER_STATE                          (PM_MASTER_STATE),                                          
   .PM_SLAVE_STATE                           (PM_SLAVE_STATE),                                          
   .SYS_AUX_PWR_DET                          (SYS_AUX_PWR_DET),                                          
                                  
                                                                                       
   .APP_HDR_VALID                            (APP_HDR_VALID),                                          
   .APP_HDR_LOG                              (APP_HDR_LOG),                                          
   .APP_ERR_BUS                              (APP_ERR_BUS),                                          
   .APP_ERR_ADVISORY                         (APP_ERR_ADVISORY),                                          
   .CFG_SEND_COR_ERR_MUX                     (CFG_SEND_COR_ERR_MUX),                                          
   .CFG_SEND_NF_ERR_MUX                      (CFG_SEND_NF_ERR_MUX),                                          
   .CFG_SEND_F_ERR_MUX                       (CFG_SEND_F_ERR_MUX),                                          
   .CFG_SYS_ERR_RC                           (CFG_SYS_ERR_RC),                                          
   .CFG_AER_RC_ERR_MUX                       (CFG_AER_RC_ERR_MUX),                                          
                                                                                       
                                                                                       
   .RADM_CPL_TIMEOUT                         (RADM_CPL_TIMEOUT),                                          
   .RADM_TIMEOUT_CPL_TC                      (RADM_TIMEOUT_CPL_TC),                                          
   .RADM_TIMEOUT_CPL_TAG                     (RADM_TIMEOUT_CPL_TAG),                                          
   .RADM_TIMEOUT_CPL_ATTR                    (RADM_TIMEOUT_CPL_ATTR),                                          
   .RADM_TIMEOUT_CPL_LEN                     (RADM_TIMEOUT_CPL_LEN),                                          
                                                                                     
                                  
                                                                                    
   .CFG_MAX_RD_REQ_SIZE                      (CFG_MAX_RD_REQ_SIZE),                                          
   .CFG_BUS_MASTER_EN                        (CFG_BUS_MASTER_EN),                                          
   .CFG_MAX_PAYLOAD_SIZE                     (CFG_MAX_PAYLOAD_SIZE),                                          
   .CFG_RCB                                  (CFG_RCB),                                          
   .CFG_MEM_SPACE_EN                         (CFG_MEM_SPACE_EN),                                          
   .CFG_PM_NO_SOFT_RST                       (CFG_PM_NO_SOFT_RST),                                          
   .CFG_CRS_SW_VIS_EN                        (CFG_CRS_SW_VIS_EN),                                          
   .CFG_NO_SNOOP_EN                          (CFG_NO_SNOOP_EN),                                         
   .CFG_RELAX_ORDER_EN                       (CFG_RELAX_ORDER_EN),                                          
   .CFG_TPH_REQ_EN                           (CFG_TPH_REQ_EN),                                          
   .CFG_PF_TPH_ST_MODE                       (CFG_PF_TPH_ST_MODE),                                          
   .CFG_PBUS_NUM                             (CFG_PBUS_NUM),                                          
   .CFG_PBUS_DEV_NUM                         (CFG_PBUS_DEV_NUM),                                          
   .RBAR_CTRL_UPDATE                         (RBAR_CTRL_UPDATE),                                          
   .CFG_ATOMIC_REQ_EN                        (CFG_ATOMIC_REQ_EN),                                          
   .CFG_ATOMIC_EGRESS_BLOCK                  (CFG_ATOMIC_EGRESS_BLOCK),                                          
   .CFG_EXT_TAG_EN                           (CFG_EXT_TAG_EN),                                
                                                                                       
   .RADM_IDLE                                (RADM_IDLE),                                  
   .RADM_Q_NOT_EMPTY                         (RADM_Q_NOT_EMPTY),                                  
   .RADM_QOVERFLOW                           (RADM_QOVERFLOW),                                  
   .DIAG_CTRL_BUS                            (DIAG_CTRL_BUS),                                  
   .DYN_DEBUG_INFO_SEL                       (DYN_DEBUG_INFO_SEL),                                  
   .CFG_LINK_AUTO_BW_MUX                     (CFG_LINK_AUTO_BW_MUX),
   .CFG_BW_MGT_MUX                           (CFG_BW_MGT_MUX),
   .CFG_PME_MUX                              (CFG_PME_MUX),
// .CFG_HP_MUX                               (CFG_HP_MUX),                                  
   .DEBUG_INFO_MUX                           (DEBUG_INFO_MUX),                                  
   .APP_RAS_DES_SD_HOLD_LTSSM                (APP_RAS_DES_SD_HOLD_LTSSM),
   .APP_RAS_DES_TBA_CTRL                     (APP_RAS_DES_TBA_CTRL),                               
                                                                                       
   .CFG_IDO_REQ_EN                           (CFG_IDO_REQ_EN),                                          
   .CFG_IDO_CPL_EN                           (CFG_IDO_CPL_EN),                                          
   .XADM_PH_CDTS                             (XADM_PH_CDTS),                                          
   .XADM_PD_CDTS                             (XADM_PD_CDTS),                                          
   .XADM_NPH_CDTS                            (XADM_NPH_CDTS),                                          
   .XADM_NPD_CDTS                            (XADM_NPD_CDTS),                                          
   .XADM_CPLH_CDTS                           (XADM_CPLH_CDTS),                                          
   .XADM_CPLD_CDTS                           (XADM_CPLD_CDTS),                                          
                                   
                                                                                       
   .MAC_PHY_POWERDOWN                        (MAC_PHY_POWERDOWN),                                          
   .PHY_MAC_RXELECIDLE                       (PHY_MAC_RXELECIDLE),                                          
   .PHY_MAC_PHYSTATUS                        (PHY_MAC_PHYSTATUS),                                          
   .PHY_MAC_RXDATA                           (PHY_MAC_RXDATA),                                          
   .PHY_MAC_RXDATAK                          (PHY_MAC_RXDATAK),                                          
   .PHY_MAC_RXVALID                          (PHY_MAC_RXVALID),                                          
   .PHY_MAC_RXSTATUS                         (PHY_MAC_RXSTATUS),                                          
   .MAC_PHY_TXDATA                           (MAC_PHY_TXDATA),                                          
   .MAC_PHY_TXDATAK                          (MAC_PHY_TXDATAK),                                          
   .MAC_PHY_TXDETECTRX_LOOPBACK              (MAC_PHY_TXDETECTRX_LOOPBACK),                                          
   .MAC_PHY_TXELECIDLE_L                     (MAC_PHY_TXELECIDLE_L),                                          
   .MAC_PHY_TXELECIDLE_H                     (MAC_PHY_TXELECIDLE_H),                                          
   .MAC_PHY_TXCOMPLIANCE                     (MAC_PHY_TXCOMPLIANCE),                                          
   .MAC_PHY_RXPOLARITY                       (MAC_PHY_RXPOLARITY),                                          
   .MAC_PHY_RATE                             (MAC_PHY_RATE),                                          
   .MAC_PHY_TXDEEMPH                         (MAC_PHY_TXDEEMPH),                                          
   .MAC_PHY_TXMARGIN                         (MAC_PHY_TXMARGIN),                                          
   .MAC_PHY_TXSWING                          (MAC_PHY_TXSWING),                                          
   .CFG_HW_AUTO_SP_DIS                       (CFG_HW_AUTO_SP_DIS),                                          
                                                                                       
                                                                                       
   .P_DATAQ_DATAOUT                          (P_DATAQ_DATAOUT),                                          
   .P_DATAQ_ADDRA                            (P_DATAQ_ADDRA),                                          
   .P_DATAQ_ADDRB                            (P_DATAQ_ADDRB),                                          
   .P_DATAQ_DATAIN                           (P_DATAQ_DATAIN),                                          
   .P_DATAQ_ENA                              (P_DATAQ_ENA),                                          
   .P_DATAQ_ENB                              (P_DATAQ_ENB),                                          
   .P_DATAQ_WEA                              (P_DATAQ_WEA),                                          
                                                                                       
   .XDLH_RETRYRAM_ADDR                       (XDLH_RETRYRAM_ADDR),                                          
   .XDLH_RETRYRAM_DATA                       (XDLH_RETRYRAM_DATA),                                          
   .XDLH_RETRYRAM_WE                         (XDLH_RETRYRAM_WE),                                          
   .XDLH_RETRYRAM_EN                         (XDLH_RETRYRAM_EN),                                          
   .RETRYRAM_XDLH_DATA                       (RETRYRAM_XDLH_DATA),                                          
                                                                                       
   .P_HDRQ_ADDRA                             (P_HDRQ_ADDRA),                                          
   .P_HDRQ_ADDRB                             (P_HDRQ_ADDRB),                                          
   .P_HDRQ_DATAIN                            (P_HDRQ_DATAIN),                                          
   .P_HDRQ_ENA                               (P_HDRQ_ENA),                                          
   .P_HDRQ_ENB                               (P_HDRQ_ENB),                                          
   .P_HDRQ_WEA                               (P_HDRQ_WEA),                                          
   .P_HDRQ_DATAOUT                           (P_HDRQ_DATAOUT),                                          
                                                                                       
                                                                         
   .RAM_TEST_EN                              (RAM_TEST_EN),                                          
   .RAM_TEST_ADDRH                           (RAM_TEST_ADDRH),                                          
   .RETRY_TEST_DATA_EN                       (RETRY_TEST_DATA_EN),                                          
   .RAM_TEST_MODE_N                          (RAM_TEST_MODE_N),                                          
                                                                                       
   .TEST_SE_N                                (1'b1),                          
   .TEST_RST_N                               (1'b1),                           
   .TEST_MODE_N                              (1'b1)
);

endmodule    




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_RAM144KSDP.v
//
// Functional description: Simple-Dual-Port 144K-bit RAM block
//
// Parameter description:
//
// Port description:
//
// Revision:
//      2018/01/09: Update display informations.
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_RAM144KSDP
#(
    parameter GRS_EN = "TRUE",
    parameter integer DATA_WIDTH_W = 36,
    parameter integer DATA_WIDTH_R = 36,
    parameter integer DO_REG = 0,
    parameter RST_TYPE = "SYNC",
    parameter integer DRM18K_NUMBER = 8,
    parameter INIT_000 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_001 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_002 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_003 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_004 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_005 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_006 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_007 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_008 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_009 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_00A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_00B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_00C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_00D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_00E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_00F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_010 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_011 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_012 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_013 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_014 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_015 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_016 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_017 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_018 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_019 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_01A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_01B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_01C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_01D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_01E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_01F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_020 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_021 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_022 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_023 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_024 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_025 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_026 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_027 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_028 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_029 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_02A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_02B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_02C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_02D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_02E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_02F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_030 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_031 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_032 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_033 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_034 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_035 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_036 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_037 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_038 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_039 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_03A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_03B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_03C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_03D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_03E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_03F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_040 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_041 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_042 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_043 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_044 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_045 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_046 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_047 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_048 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_049 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_04A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_04B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_04C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_04D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_04E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_04F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_050 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_051 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_052 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_053 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_054 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_055 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_056 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_057 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_058 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_059 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_05A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_05B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_05C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_05D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_05E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_05F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_060 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_061 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_062 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_063 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_064 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_065 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_066 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_067 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_068 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_069 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_06A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_06B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_06C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_06D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_06E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_06F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_070 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_071 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_072 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_073 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_074 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_075 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_076 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_077 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_078 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_079 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_07A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_07B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_07C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_07D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_07E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_07F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_080 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_081 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_082 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_083 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_084 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_085 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_086 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_087 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_088 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_089 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_08A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_08B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_08C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_08D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_08E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_08F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_090 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_091 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_092 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_093 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_094 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_095 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_096 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_097 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_098 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_099 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_09A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_09B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_09C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_09D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_09E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_09F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0A0 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0A1 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0A2 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0A3 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0A4 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0A5 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0A6 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0A7 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0A8 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0A9 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0AA = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0AB = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0AC = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0AD = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0AE = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0AF = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0B0 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0B1 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0B2 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0B3 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0B4 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0B5 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0B6 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0B7 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0B8 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0B9 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0BA = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0BB = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0BC = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0BD = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0BE = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0BF = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0C0 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0C1 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0C2 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0C3 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0C4 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0C5 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0C6 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0C7 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0C8 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0C9 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0CA = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0CB = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0CC = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0CD = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0CE = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0CF = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0D0 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0D1 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0D2 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0D3 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0D4 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0D5 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0D6 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0D7 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0D8 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0D9 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0DA = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0DB = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0DC = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0DD = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0DE = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0DF = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0E0 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0E1 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0E2 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0E3 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0E4 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0E5 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0E6 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0E7 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0E8 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0E9 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0EA = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0EB = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0EC = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0ED = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0EE = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0EF = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0F0 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0F1 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0F2 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0F3 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0F4 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0F5 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0F6 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0F7 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0F8 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0F9 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0FA = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0FB = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0FC = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0FD = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0FE = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_0FF = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_100 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_101 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_102 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_103 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_104 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_105 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_106 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_107 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_108 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_109 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_10A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_10B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_10C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_10D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_10E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_10F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_110 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_111 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_112 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_113 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_114 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_115 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_116 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_117 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_118 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_119 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_11A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_11B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_11C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_11D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_11E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_11F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_120 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_121 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_122 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_123 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_124 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_125 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_126 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_127 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_128 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_129 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_12A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_12B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_12C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_12D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_12E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_12F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_130 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_131 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_132 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_133 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_134 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_135 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_136 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_137 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_138 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_139 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_13A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_13B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_13C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_13D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_13E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_13F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_140 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_141 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_142 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_143 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_144 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_145 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_146 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_147 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_148 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_149 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_14A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_14B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_14C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_14D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_14E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_14F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_150 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_151 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_152 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_153 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_154 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_155 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_156 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_157 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_158 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_159 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_15A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_15B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_15C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_15D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_15E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_15F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_160 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_161 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_162 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_163 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_164 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_165 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_166 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_167 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_168 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_169 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_16A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_16B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_16C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_16D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_16E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_16F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_170 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_171 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_172 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_173 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_174 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_175 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_176 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_177 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_178 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_179 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_17A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_17B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_17C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_17D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_17E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_17F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_180 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_181 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_182 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_183 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_184 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_185 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_186 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_187 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_188 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_189 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_18A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_18B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_18C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_18D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_18E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_18F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_190 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_191 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_192 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_193 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_194 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_195 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_196 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_197 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_198 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_199 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_19A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_19B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_19C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_19D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_19E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_19F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1A0 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1A1 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1A2 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1A3 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1A4 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1A5 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1A6 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1A7 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1A8 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1A9 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1AA = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1AB = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1AC = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1AD = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1AE = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1AF = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1B0 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1B1 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1B2 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1B3 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1B4 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1B5 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1B6 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1B7 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1B8 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1B9 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1BA = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1BB = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1BC = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1BD = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1BE = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1BF = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1C0 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1C1 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1C2 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1C3 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1C4 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1C5 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1C6 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1C7 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1C8 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1C9 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1CA = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1CB = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1CC = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1CD = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1CE = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1CF = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1D0 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1D1 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1D2 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1D3 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1D4 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1D5 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1D6 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1D7 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1D8 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1D9 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1DA = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1DB = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1DC = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1DD = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1DE = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1DF = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1E0 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1E1 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1E2 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1E3 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1E4 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1E5 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1E6 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1E7 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1E8 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1E9 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1EA = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1EB = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1EC = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1ED = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1EE = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1EF = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1F0 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1F1 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1F2 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1F3 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1F4 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1F5 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1F6 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1F7 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1F8 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1F9 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1FA = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1FB = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1FC = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1FD = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1FE = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1FF = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_FILE = "NONE"
) (
    output [35:0] DO,
    input [35:0] DI,
    input [16:0] WADDR,
    input WCLK,
    input WCE,
    input WE,
    input [3:0] BE,
    input [16:0] RADDR,
    input RCLK,
    input RCE,
    input ORCE,
    input RST
);

    wire [35:0] dangle_a36;
    supply0 Gnd;

    //
    // parameter check
    //

    initial begin
        case (DATA_WIDTH_W)
            1, 2, 4, 8, 16, 32, 9, 18, 36: begin
                case (DATA_WIDTH_R)
                    1, 2, 4, 8, 16, 32, 9, 18, 36:    ;  // null 
                    default: begin
                        $display("ERROR: GTP_RAM144KSDP instance %m parameter DATA_WIDTH_R:%d is illegal. The legal values are 1,2,4,8,16,9,18 or 36.",DATA_WIDTH_R);
                        $finish;
                    end
                endcase
            end
            default: begin
                $display("ERROR: GTP_RAM144KSDP instance %m parameter DATA_WIDTH_W:%d is illegal. The legal values are 1,2,4,8,16,9,18 or 36.",DATA_WIDTH_W);
                $finish;
            end
        endcase

        if (DATA_WIDTH_W <= 18 && DATA_WIDTH_W <= 18) begin
            $display("Warning: GTP_RAM144KSDP instance %m suggest map to GTP_RAM144K");
        end

        if (RST_TYPE != "ASYNC" && RST_TYPE != "SYNC") begin
            $display("ERROR: GTP_RAM144KSDP instance %m parameter:%s is illegal. The legal values are ASYNC or SYNC.",RST_TYPE);
            $finish;
        end

        if (DO_REG != 0 && DO_REG != 1) begin
            $display("ERROR: GTP_RAM144KSDP instance %m parameter: DO_REG:%d is illegal. The legal values are 0 or 1 .",DO_REG);
            $finish;
        end
    end

    // port A for write
    // port B for read

    INT_RAM144K
    #(
        .GRS_EN(GRS_EN),
        .DATA_WIDTH_A(DATA_WIDTH_W),
        .DATA_WIDTH_B(DATA_WIDTH_R),
        .CLEAR_TYPE(RST_TYPE),
        .OUTPUT_REG_B(DO_REG),
        .INIT_FILE(INIT_FILE),
        .INIT_000(INIT_000),
        .INIT_001(INIT_001),
        .INIT_002(INIT_002),
        .INIT_003(INIT_003),
        .INIT_004(INIT_004),
        .INIT_005(INIT_005),
        .INIT_006(INIT_006),
        .INIT_007(INIT_007),
        .INIT_008(INIT_008),
        .INIT_009(INIT_009),
        .INIT_00A(INIT_00A),
        .INIT_00B(INIT_00B),
        .INIT_00C(INIT_00C),
        .INIT_00D(INIT_00D),
        .INIT_00E(INIT_00E),
        .INIT_00F(INIT_00F),
        .INIT_010(INIT_010),
        .INIT_011(INIT_011),
        .INIT_012(INIT_012),
        .INIT_013(INIT_013),
        .INIT_014(INIT_014),
        .INIT_015(INIT_015),
        .INIT_016(INIT_016),
        .INIT_017(INIT_017),
        .INIT_018(INIT_018),
        .INIT_019(INIT_019),
        .INIT_01A(INIT_01A),
        .INIT_01B(INIT_01B),
        .INIT_01C(INIT_01C),
        .INIT_01D(INIT_01D),
        .INIT_01E(INIT_01E),
        .INIT_01F(INIT_01F),
        .INIT_020(INIT_020),
        .INIT_021(INIT_021),
        .INIT_022(INIT_022),
        .INIT_023(INIT_023),
        .INIT_024(INIT_024),
        .INIT_025(INIT_025),
        .INIT_026(INIT_026),
        .INIT_027(INIT_027),
        .INIT_028(INIT_028),
        .INIT_029(INIT_029),
        .INIT_02A(INIT_02A),
        .INIT_02B(INIT_02B),
        .INIT_02C(INIT_02C),
        .INIT_02D(INIT_02D),
        .INIT_02E(INIT_02E),
        .INIT_02F(INIT_02F),
        .INIT_030(INIT_030),
        .INIT_031(INIT_031),
        .INIT_032(INIT_032),
        .INIT_033(INIT_033),
        .INIT_034(INIT_034),
        .INIT_035(INIT_035),
        .INIT_036(INIT_036),
        .INIT_037(INIT_037),
        .INIT_038(INIT_038),
        .INIT_039(INIT_039),
        .INIT_03A(INIT_03A),
        .INIT_03B(INIT_03B),
        .INIT_03C(INIT_03C),
        .INIT_03D(INIT_03D),
        .INIT_03E(INIT_03E),
        .INIT_03F(INIT_03F),
        .INIT_040(INIT_040),
        .INIT_041(INIT_041),
        .INIT_042(INIT_042),
        .INIT_043(INIT_043),
        .INIT_044(INIT_044),
        .INIT_045(INIT_045),
        .INIT_046(INIT_046),
        .INIT_047(INIT_047),
        .INIT_048(INIT_048),
        .INIT_049(INIT_049),
        .INIT_04A(INIT_04A),
        .INIT_04B(INIT_04B),
        .INIT_04C(INIT_04C),
        .INIT_04D(INIT_04D),
        .INIT_04E(INIT_04E),
        .INIT_04F(INIT_04F),
        .INIT_050(INIT_050),
        .INIT_051(INIT_051),
        .INIT_052(INIT_052),
        .INIT_053(INIT_053),
        .INIT_054(INIT_054),
        .INIT_055(INIT_055),
        .INIT_056(INIT_056),
        .INIT_057(INIT_057),
        .INIT_058(INIT_058),
        .INIT_059(INIT_059),
        .INIT_05A(INIT_05A),
        .INIT_05B(INIT_05B),
        .INIT_05C(INIT_05C),
        .INIT_05D(INIT_05D),
        .INIT_05E(INIT_05E),
        .INIT_05F(INIT_05F),
        .INIT_060(INIT_060),
        .INIT_061(INIT_061),
        .INIT_062(INIT_062),
        .INIT_063(INIT_063),
        .INIT_064(INIT_064),
        .INIT_065(INIT_065),
        .INIT_066(INIT_066),
        .INIT_067(INIT_067),
        .INIT_068(INIT_068),
        .INIT_069(INIT_069),
        .INIT_06A(INIT_06A),
        .INIT_06B(INIT_06B),
        .INIT_06C(INIT_06C),
        .INIT_06D(INIT_06D),
        .INIT_06E(INIT_06E),
        .INIT_06F(INIT_06F),
        .INIT_070(INIT_070),
        .INIT_071(INIT_071),
        .INIT_072(INIT_072),
        .INIT_073(INIT_073),
        .INIT_074(INIT_074),
        .INIT_075(INIT_075),
        .INIT_076(INIT_076),
        .INIT_077(INIT_077),
        .INIT_078(INIT_078),
        .INIT_079(INIT_079),
        .INIT_07A(INIT_07A),
        .INIT_07B(INIT_07B),
        .INIT_07C(INIT_07C),
        .INIT_07D(INIT_07D),
        .INIT_07E(INIT_07E),
        .INIT_07F(INIT_07F),
        .INIT_080(INIT_080),
        .INIT_081(INIT_081),
        .INIT_082(INIT_082),
        .INIT_083(INIT_083),
        .INIT_084(INIT_084),
        .INIT_085(INIT_085),
        .INIT_086(INIT_086),
        .INIT_087(INIT_087),
        .INIT_088(INIT_088),
        .INIT_089(INIT_089),
        .INIT_08A(INIT_08A),
        .INIT_08B(INIT_08B),
        .INIT_08C(INIT_08C),
        .INIT_08D(INIT_08D),
        .INIT_08E(INIT_08E),
        .INIT_08F(INIT_08F),
        .INIT_090(INIT_090),
        .INIT_091(INIT_091),
        .INIT_092(INIT_092),
        .INIT_093(INIT_093),
        .INIT_094(INIT_094),
        .INIT_095(INIT_095),
        .INIT_096(INIT_096),
        .INIT_097(INIT_097),
        .INIT_098(INIT_098),
        .INIT_099(INIT_099),
        .INIT_09A(INIT_09A),
        .INIT_09B(INIT_09B),
        .INIT_09C(INIT_09C),
        .INIT_09D(INIT_09D),
        .INIT_09E(INIT_09E),
        .INIT_09F(INIT_09F),
        .INIT_0A0(INIT_0A0),
        .INIT_0A1(INIT_0A1),
        .INIT_0A2(INIT_0A2),
        .INIT_0A3(INIT_0A3),
        .INIT_0A4(INIT_0A4),
        .INIT_0A5(INIT_0A5),
        .INIT_0A6(INIT_0A6),
        .INIT_0A7(INIT_0A7),
        .INIT_0A8(INIT_0A8),
        .INIT_0A9(INIT_0A9),
        .INIT_0AA(INIT_0AA),
        .INIT_0AB(INIT_0AB),
        .INIT_0AC(INIT_0AC),
        .INIT_0AD(INIT_0AD),
        .INIT_0AE(INIT_0AE),
        .INIT_0AF(INIT_0AF),
        .INIT_0B0(INIT_0B0),
        .INIT_0B1(INIT_0B1),
        .INIT_0B2(INIT_0B2),
        .INIT_0B3(INIT_0B3),
        .INIT_0B4(INIT_0B4),
        .INIT_0B5(INIT_0B5),
        .INIT_0B6(INIT_0B6),
        .INIT_0B7(INIT_0B7),
        .INIT_0B8(INIT_0B8),
        .INIT_0B9(INIT_0B9),
        .INIT_0BA(INIT_0BA),
        .INIT_0BB(INIT_0BB),
        .INIT_0BC(INIT_0BC),
        .INIT_0BD(INIT_0BD),
        .INIT_0BE(INIT_0BE),
        .INIT_0BF(INIT_0BF),
        .INIT_0C0(INIT_0C0),
        .INIT_0C1(INIT_0C1),
        .INIT_0C2(INIT_0C2),
        .INIT_0C3(INIT_0C3),
        .INIT_0C4(INIT_0C4),
        .INIT_0C5(INIT_0C5),
        .INIT_0C6(INIT_0C6),
        .INIT_0C7(INIT_0C7),
        .INIT_0C8(INIT_0C8),
        .INIT_0C9(INIT_0C9),
        .INIT_0CA(INIT_0CA),
        .INIT_0CB(INIT_0CB),
        .INIT_0CC(INIT_0CC),
        .INIT_0CD(INIT_0CD),
        .INIT_0CE(INIT_0CE),
        .INIT_0CF(INIT_0CF),
        .INIT_0D0(INIT_0D0),
        .INIT_0D1(INIT_0D1),
        .INIT_0D2(INIT_0D2),
        .INIT_0D3(INIT_0D3),
        .INIT_0D4(INIT_0D4),
        .INIT_0D5(INIT_0D5),
        .INIT_0D6(INIT_0D6),
        .INIT_0D7(INIT_0D7),
        .INIT_0D8(INIT_0D8),
        .INIT_0D9(INIT_0D9),
        .INIT_0DA(INIT_0DA),
        .INIT_0DB(INIT_0DB),
        .INIT_0DC(INIT_0DC),
        .INIT_0DD(INIT_0DD),
        .INIT_0DE(INIT_0DE),
        .INIT_0DF(INIT_0DF),
        .INIT_0E0(INIT_0E0),
        .INIT_0E1(INIT_0E1),
        .INIT_0E2(INIT_0E2),
        .INIT_0E3(INIT_0E3),
        .INIT_0E4(INIT_0E4),
        .INIT_0E5(INIT_0E5),
        .INIT_0E6(INIT_0E6),
        .INIT_0E7(INIT_0E7),
        .INIT_0E8(INIT_0E8),
        .INIT_0E9(INIT_0E9),
        .INIT_0EA(INIT_0EA),
        .INIT_0EB(INIT_0EB),
        .INIT_0EC(INIT_0EC),
        .INIT_0ED(INIT_0ED),
        .INIT_0EE(INIT_0EE),
        .INIT_0EF(INIT_0EF),
        .INIT_0F0(INIT_0F0),
        .INIT_0F1(INIT_0F1),
        .INIT_0F2(INIT_0F2),
        .INIT_0F3(INIT_0F3),
        .INIT_0F4(INIT_0F4),
        .INIT_0F5(INIT_0F5),
        .INIT_0F6(INIT_0F6),
        .INIT_0F7(INIT_0F7),
        .INIT_0F8(INIT_0F8),
        .INIT_0F9(INIT_0F9),
        .INIT_0FA(INIT_0FA),
        .INIT_0FB(INIT_0FB),
        .INIT_0FC(INIT_0FC),
        .INIT_0FD(INIT_0FD),
        .INIT_0FE(INIT_0FE),
        .INIT_0FF(INIT_0FF),
        .INIT_100(INIT_100),
        .INIT_101(INIT_101),
        .INIT_102(INIT_102),
        .INIT_103(INIT_103),
        .INIT_104(INIT_104),
        .INIT_105(INIT_105),
        .INIT_106(INIT_106),
        .INIT_107(INIT_107),
        .INIT_108(INIT_108),
        .INIT_109(INIT_109),
        .INIT_10A(INIT_10A),
        .INIT_10B(INIT_10B),
        .INIT_10C(INIT_10C),
        .INIT_10D(INIT_10D),
        .INIT_10E(INIT_10E),
        .INIT_10F(INIT_10F),
        .INIT_110(INIT_110),
        .INIT_111(INIT_111),
        .INIT_112(INIT_112),
        .INIT_113(INIT_113),
        .INIT_114(INIT_114),
        .INIT_115(INIT_115),
        .INIT_116(INIT_116),
        .INIT_117(INIT_117),
        .INIT_118(INIT_118),
        .INIT_119(INIT_119),
        .INIT_11A(INIT_11A),
        .INIT_11B(INIT_11B),
        .INIT_11C(INIT_11C),
        .INIT_11D(INIT_11D),
        .INIT_11E(INIT_11E),
        .INIT_11F(INIT_11F),
        .INIT_120(INIT_120),
        .INIT_121(INIT_121),
        .INIT_122(INIT_122),
        .INIT_123(INIT_123),
        .INIT_124(INIT_124),
        .INIT_125(INIT_125),
        .INIT_126(INIT_126),
        .INIT_127(INIT_127),
        .INIT_128(INIT_128),
        .INIT_129(INIT_129),
        .INIT_12A(INIT_12A),
        .INIT_12B(INIT_12B),
        .INIT_12C(INIT_12C),
        .INIT_12D(INIT_12D),
        .INIT_12E(INIT_12E),
        .INIT_12F(INIT_12F),
        .INIT_130(INIT_130),
        .INIT_131(INIT_131),
        .INIT_132(INIT_132),
        .INIT_133(INIT_133),
        .INIT_134(INIT_134),
        .INIT_135(INIT_135),
        .INIT_136(INIT_136),
        .INIT_137(INIT_137),
        .INIT_138(INIT_138),
        .INIT_139(INIT_139),
        .INIT_13A(INIT_13A),
        .INIT_13B(INIT_13B),
        .INIT_13C(INIT_13C),
        .INIT_13D(INIT_13D),
        .INIT_13E(INIT_13E),
        .INIT_13F(INIT_13F),
        .INIT_140(INIT_140),
        .INIT_141(INIT_141),
        .INIT_142(INIT_142),
        .INIT_143(INIT_143),
        .INIT_144(INIT_144),
        .INIT_145(INIT_145),
        .INIT_146(INIT_146),
        .INIT_147(INIT_147),
        .INIT_148(INIT_148),
        .INIT_149(INIT_149),
        .INIT_14A(INIT_14A),
        .INIT_14B(INIT_14B),
        .INIT_14C(INIT_14C),
        .INIT_14D(INIT_14D),
        .INIT_14E(INIT_14E),
        .INIT_14F(INIT_14F),
        .INIT_150(INIT_150),
        .INIT_151(INIT_151),
        .INIT_152(INIT_152),
        .INIT_153(INIT_153),
        .INIT_154(INIT_154),
        .INIT_155(INIT_155),
        .INIT_156(INIT_156),
        .INIT_157(INIT_157),
        .INIT_158(INIT_158),
        .INIT_159(INIT_159),
        .INIT_15A(INIT_15A),
        .INIT_15B(INIT_15B),
        .INIT_15C(INIT_15C),
        .INIT_15D(INIT_15D),
        .INIT_15E(INIT_15E),
        .INIT_15F(INIT_15F),
        .INIT_160(INIT_160),
        .INIT_161(INIT_161),
        .INIT_162(INIT_162),
        .INIT_163(INIT_163),
        .INIT_164(INIT_164),
        .INIT_165(INIT_165),
        .INIT_166(INIT_166),
        .INIT_167(INIT_167),
        .INIT_168(INIT_168),
        .INIT_169(INIT_169),
        .INIT_16A(INIT_16A),
        .INIT_16B(INIT_16B),
        .INIT_16C(INIT_16C),
        .INIT_16D(INIT_16D),
        .INIT_16E(INIT_16E),
        .INIT_16F(INIT_16F),
        .INIT_170(INIT_170),
        .INIT_171(INIT_171),
        .INIT_172(INIT_172),
        .INIT_173(INIT_173),
        .INIT_174(INIT_174),
        .INIT_175(INIT_175),
        .INIT_176(INIT_176),
        .INIT_177(INIT_177),
        .INIT_178(INIT_178),
        .INIT_179(INIT_179),
        .INIT_17A(INIT_17A),
        .INIT_17B(INIT_17B),
        .INIT_17C(INIT_17C),
        .INIT_17D(INIT_17D),
        .INIT_17E(INIT_17E),
        .INIT_17F(INIT_17F),
        .INIT_180(INIT_180),
        .INIT_181(INIT_181),
        .INIT_182(INIT_182),
        .INIT_183(INIT_183),
        .INIT_184(INIT_184),
        .INIT_185(INIT_185),
        .INIT_186(INIT_186),
        .INIT_187(INIT_187),
        .INIT_188(INIT_188),
        .INIT_189(INIT_189),
        .INIT_18A(INIT_18A),
        .INIT_18B(INIT_18B),
        .INIT_18C(INIT_18C),
        .INIT_18D(INIT_18D),
        .INIT_18E(INIT_18E),
        .INIT_18F(INIT_18F),
        .INIT_190(INIT_190),
        .INIT_191(INIT_191),
        .INIT_192(INIT_192),
        .INIT_193(INIT_193),
        .INIT_194(INIT_194),
        .INIT_195(INIT_195),
        .INIT_196(INIT_196),
        .INIT_197(INIT_197),
        .INIT_198(INIT_198),
        .INIT_199(INIT_199),
        .INIT_19A(INIT_19A),
        .INIT_19B(INIT_19B),
        .INIT_19C(INIT_19C),
        .INIT_19D(INIT_19D),
        .INIT_19E(INIT_19E),
        .INIT_19F(INIT_19F),
        .INIT_1A0(INIT_1A0),
        .INIT_1A1(INIT_1A1),
        .INIT_1A2(INIT_1A2),
        .INIT_1A3(INIT_1A3),
        .INIT_1A4(INIT_1A4),
        .INIT_1A5(INIT_1A5),
        .INIT_1A6(INIT_1A6),
        .INIT_1A7(INIT_1A7),
        .INIT_1A8(INIT_1A8),
        .INIT_1A9(INIT_1A9),
        .INIT_1AA(INIT_1AA),
        .INIT_1AB(INIT_1AB),
        .INIT_1AC(INIT_1AC),
        .INIT_1AD(INIT_1AD),
        .INIT_1AE(INIT_1AE),
        .INIT_1AF(INIT_1AF),
        .INIT_1B0(INIT_1B0),
        .INIT_1B1(INIT_1B1),
        .INIT_1B2(INIT_1B2),
        .INIT_1B3(INIT_1B3),
        .INIT_1B4(INIT_1B4),
        .INIT_1B5(INIT_1B5),
        .INIT_1B6(INIT_1B6),
        .INIT_1B7(INIT_1B7),
        .INIT_1B8(INIT_1B8),
        .INIT_1B9(INIT_1B9),
        .INIT_1BA(INIT_1BA),
        .INIT_1BB(INIT_1BB),
        .INIT_1BC(INIT_1BC),
        .INIT_1BD(INIT_1BD),
        .INIT_1BE(INIT_1BE),
        .INIT_1BF(INIT_1BF),
        .INIT_1C0(INIT_1C0),
        .INIT_1C1(INIT_1C1),
        .INIT_1C2(INIT_1C2),
        .INIT_1C3(INIT_1C3),
        .INIT_1C4(INIT_1C4),
        .INIT_1C5(INIT_1C5),
        .INIT_1C6(INIT_1C6),
        .INIT_1C7(INIT_1C7),
        .INIT_1C8(INIT_1C8),
        .INIT_1C9(INIT_1C9),
        .INIT_1CA(INIT_1CA),
        .INIT_1CB(INIT_1CB),
        .INIT_1CC(INIT_1CC),
        .INIT_1CD(INIT_1CD),
        .INIT_1CE(INIT_1CE),
        .INIT_1CF(INIT_1CF),
        .INIT_1D0(INIT_1D0),
        .INIT_1D1(INIT_1D1),
        .INIT_1D2(INIT_1D2),
        .INIT_1D3(INIT_1D3),
        .INIT_1D4(INIT_1D4),
        .INIT_1D5(INIT_1D5),
        .INIT_1D6(INIT_1D6),
        .INIT_1D7(INIT_1D7),
        .INIT_1D8(INIT_1D8),
        .INIT_1D9(INIT_1D9),
        .INIT_1DA(INIT_1DA),
        .INIT_1DB(INIT_1DB),
        .INIT_1DC(INIT_1DC),
        .INIT_1DD(INIT_1DD),
        .INIT_1DE(INIT_1DE),
        .INIT_1DF(INIT_1DF),
        .INIT_1E0(INIT_1E0),
        .INIT_1E1(INIT_1E1),
        .INIT_1E2(INIT_1E2),
        .INIT_1E3(INIT_1E3),
        .INIT_1E4(INIT_1E4),
        .INIT_1E5(INIT_1E5),
        .INIT_1E6(INIT_1E6),
        .INIT_1E7(INIT_1E7),
        .INIT_1E8(INIT_1E8),
        .INIT_1E9(INIT_1E9),
        .INIT_1EA(INIT_1EA),
        .INIT_1EB(INIT_1EB),
        .INIT_1EC(INIT_1EC),
        .INIT_1ED(INIT_1ED),
        .INIT_1EE(INIT_1EE),
        .INIT_1EF(INIT_1EF),
        .INIT_1F0(INIT_1F0),
        .INIT_1F1(INIT_1F1),
        .INIT_1F2(INIT_1F2),
        .INIT_1F3(INIT_1F3),
        .INIT_1F4(INIT_1F4),
        .INIT_1F5(INIT_1F5),
        .INIT_1F6(INIT_1F6),
        .INIT_1F7(INIT_1F7),
        .INIT_1F8(INIT_1F8),
        .INIT_1F9(INIT_1F9),
        .INIT_1FA(INIT_1FA),
        .INIT_1FB(INIT_1FB),
        .INIT_1FC(INIT_1FC),
        .INIT_1FD(INIT_1FD),
        .INIT_1FE(INIT_1FE),
        .INIT_1FF(INIT_1FF),
        .RAM_MODE("SIMPLE_DUAL_PORT")
    ) bram (
        .CLKA(WCLK), .CEA(WCE), .WEA(WE), .BEA(BE),
        .ADDRA(WADDR), .DIA(DI),
        .ORCEA(Gnd), .CLRA(Gnd), .DOA(dangle_a36),
        .CLKB(RCLK), .CEB(RCE), .WEB(Gnd), .BEB({4{Gnd}}),
        .ADDRB(RADDR), .DIB({36{Gnd}}),
        .ORCEB(ORCE), .CLRB(RST), .DOB(DO)
    );

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_PREADD_MULTADD27.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

//P = A0*(B0+-C0) +/- A1*(B1+-C1)
`timescale 1 ns / 1 ps

module GTP_PREADD_MULTADD27 #(
    parameter GRS_EN            = "TRUE", //"TRUE"; "FALSE"
    parameter SYNC_RST          = "FALSE", //"TRUE"; "FALSE"  
    parameter INREG_EN          = "FALSE", //"TRUE"; "FALSE"
    parameter PREREG_EN         = "FALSE", //"TRUE"; "FALSE"
    parameter PIPEREG_EN        = "FALSE", //"TRUE"; "FALSE"
    parameter OUTREG_EN         = "FALSE", //"TRUE"; "FALSE"
    parameter ADDSUB_OP         = 0 ,
    parameter DYN_ADDSUB_OP     = 1
)(
    output  [55-1:0] P,
    input   CE,
    input   RST,
    input   CLK,
    input   [27-1:0] A0,
    input   [27-1:0] A1,
    input   [26-1:0] B0,
    input   [26-1:0] B1,
    input   [26-1:0] C0,
    input   [26-1:0] C1,
    input   A_SIGNED,
    input   B_SIGNED,
    input   C_SIGNED,
    input   [1:0] PREADDSUB,
    input   ADDSUB
);


    INT_PREADD_MULTADD #(
        . GRS_EN(GRS_EN),    
        . SYNC_RST(SYNC_RST),  
        . INREG_EN(INREG_EN), 
        . PREREG_EN(PREREG_EN), 
        . PIPEREG_EN(PIPEREG_EN),
        . OUTREG_EN(OUTREG_EN), 
        . ADDSUB_OP(ADDSUB_OP),   
        . DYN_OP_ADDSUB(DYN_ADDSUB_OP),
        . ASIZE(27), 
        . BSIZE(26)
    ) U_INT_PREADD_MULTADD(
        . CE(CE),
        . RST(RST),
        . CLK(CLK),
        . A0(A0),
        . A1(A1),
        . B0(B0),
        . B1(B1),
        . C0(C0),
        . C1(C1),
        . A_SIGNED(A_SIGNED),
        . B_SIGNED(B_SIGNED),
        . C_SIGNED(C_SIGNED),
        . PREADDSUB(PREADDSUB),
        . ADDSUB(ADDSUB),
        . P(P)
    );   


endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2016 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_RAM256X1SP.v
//
// Functional description: single-port 256x1 distributed ram
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_RAM256X1SP
#(
    parameter [255:0] INIT = 256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000
) (
    output  DO,
    input   DI,
    input [7:0] ADDR,
    input WCLK,
    input WE
);
//synthesis translate_off
    reg [255:0] mem ;

    initial begin
        mem = INIT;
    end

    always @(posedge WCLK) begin
        if (WE == 1'b1) begin
            mem[ADDR] <= DI;
        end
    end

    assign DO = mem[ADDR];
//synthesis translate_on
endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_IGDES7.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_IGDES7 #(
parameter GRS_EN = "TRUE", //"TRUE"; "FALSE"
parameter LRS_EN = "TRUE",  //"TRUE"; "FALSE"
parameter DPI_EN = "FALSE"  //"TRUE"; "FALSE"
)(
output [6:0] Q,
output [1:0] DPI_STS,
input [1:0] DPI_CTRL,
input DPI_STS_CLR_N,
input PADI,
input DESCLK,
input RCLK,
input RST
);

//synthesis translate_off
wire [7:0] PADI_D;
reg DPI_P;
reg [1:0] DPI_STS_R;
wire COMP_BEFORE;
wire COMP_AFTER;
wire COMP_BEFORE_D;
wire COMP_AFTER_D;
wire PD_BEFORE;
wire PD_AFTER;
wire DPI_BEFORE_POS_REG_T;
wire DPI_AFTER_POS_REG_T;
wire DPI_BEFORE_NEG_REG_T;
wire DPI_AFTER_NEG_REG_T;
wire AFTER_POS;
wire BEFORE_POS;
wire AFTER_NEG;
wire BEFORE_NEG;
reg DPI_N_reg;
reg DPI_BEFORE;
reg DPI_AFTER;
reg DPI_BEFORE_POS_REG;
reg DPI_BEFORE_NEG_REG;
reg DPI_AFTER_POS_REG;
reg DPI_AFTER_NEG_REG;
reg [7:0] shift_reg;
reg [6:0] capture_reg;
reg [2:0] cnt;
reg rstn_dly;
reg [6:0] Q_reg;

initial begin
DPI_P              = 0;
DPI_STS_R          = 0;
DPI_N_reg          = 0;
DPI_BEFORE         = 0;
DPI_AFTER          = 0;
DPI_BEFORE_POS_REG = 0;
DPI_BEFORE_NEG_REG = 0;
DPI_AFTER_POS_REG  = 0;
DPI_AFTER_NEG_REG  = 0;

shift_reg    = 0;
capture_reg  = 0;
cnt          = 0;
rstn_dly     = 0;
Q_reg        = 0;
end

assign global_rstn = (GRS_EN == "TRUE") ? GRS_INST.GRSNET : 1'b1;
assign lsr_rstn = LRS_EN == "TRUE" ? (~RST) : 1'b1;


assign  #0.05 PADI_D[0] =  PADI;
assign  #0.05 PADI_D[1] =  PADI_D[0];
assign  #0.05 PADI_D[2] =  PADI_D[1];
assign  #0.05 PADI_D[3] =  PADI_D[2];
assign  #0.05 PADI_D[4] =  PADI_D[3];
assign  #0.05 PADI_D[5] =  PADI_D[4];
assign  #0.05 PADI_D[6] =  PADI_D[5];
assign  #0.05 PADI_D[7] =  PADI_D[6];

assign PADI_SAMPLE = (DPI_EN == "TRUE") ? PADI_D[3] : PADI;

always @(posedge DESCLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_P <= 0;
   else if (!lsr_rstn)
      DPI_P <= 0;
   else
      DPI_P <= PADI_SAMPLE;
end

always @(negedge DESCLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_N_reg <= 0;
   else if (!lsr_rstn)
      DPI_N_reg <= 0;
   else 
      DPI_N_reg <= PADI_SAMPLE;
end

always @(*) begin
   case (DPI_CTRL[1:0])
      2'd0:    begin DPI_BEFORE = PADI_D[2];  DPI_AFTER = PADI_D[4]; end
      2'd1:    begin DPI_BEFORE = PADI_D[1];  DPI_AFTER = PADI_D[5]; end
      2'd2:    begin DPI_BEFORE = PADI_D[0];  DPI_AFTER = PADI_D[6]; end
      default: begin DPI_BEFORE = PADI;       DPI_AFTER = PADI_D[7]; end
   endcase
end

always @(posedge DESCLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_BEFORE_POS_REG <= 0;
   else if (!lsr_rstn)
      DPI_BEFORE_POS_REG <= 0;
   else   
      DPI_BEFORE_POS_REG <= DPI_BEFORE;
end

always @(negedge DESCLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_BEFORE_NEG_REG <= 0;
   else if (!lsr_rstn)
      DPI_BEFORE_NEG_REG <= 0;
   else     
      DPI_BEFORE_NEG_REG <= DPI_BEFORE;
end


always @(posedge DESCLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_AFTER_POS_REG <= 0;
   else if (!lsr_rstn)
      DPI_AFTER_POS_REG <= 0;
   else   
      DPI_AFTER_POS_REG <= DPI_AFTER;
end


always @(negedge DESCLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_AFTER_NEG_REG <= 0;
   else if (!lsr_rstn)
      DPI_AFTER_NEG_REG <= 0;
   else     
      DPI_AFTER_NEG_REG <= DPI_AFTER;
end

assign BEFORE_POS = DPI_BEFORE_POS_REG_T ^ DPI_P;
assign DPI_BEFORE_POS_REG_T = (DPI_EN == "TRUE") ? DPI_BEFORE_POS_REG : 0;

assign AFTER_POS = DPI_AFTER_POS_REG_T ^ DPI_P;
assign DPI_AFTER_POS_REG_T = (DPI_EN == "TRUE") ? DPI_AFTER_POS_REG : 0;

assign BEFORE_NEG = DPI_BEFORE_NEG_REG_T ^ DPI_N_reg;
assign DPI_BEFORE_NEG_REG_T = (DPI_EN == "TRUE") ? DPI_BEFORE_NEG_REG : 0;

assign AFTER_NEG = DPI_AFTER_NEG_REG_T ^ DPI_N_reg;
assign DPI_AFTER_NEG_REG_T = (DPI_EN == "TRUE") ? DPI_AFTER_NEG_REG : 0;


assign COMP_BEFORE = BEFORE_POS || BEFORE_NEG;
assign COMP_AFTER = AFTER_POS || AFTER_NEG;

assign #0.1 COMP_BEFORE_D = COMP_BEFORE;
assign #0.1 COMP_AFTER_D = COMP_AFTER;

assign PD_BEFORE = COMP_BEFORE && COMP_BEFORE_D;
assign PD_AFTER = COMP_AFTER && COMP_AFTER_D;


always @(posedge DPI_STS_CLR_N or negedge global_rstn or negedge lsr_rstn or posedge  PD_BEFORE) begin
   if (!global_rstn)
      DPI_STS_R[0] <= 0;
   else if (!lsr_rstn)
      DPI_STS_R[0] <= 0;
   else if (PD_BEFORE)
      DPI_STS_R[0] <= 1;
   else
      DPI_STS_R[0] <= 1'b0;
end

always @(posedge DPI_STS_CLR_N or negedge global_rstn or negedge lsr_rstn or posedge PD_AFTER) begin
   if (!global_rstn)
      DPI_STS_R[1] <= 0;
   else if (!lsr_rstn)
      DPI_STS_R[1] <= 0;
   else if (PD_AFTER)
      DPI_STS_R[1] <= 1;
   else
      DPI_STS_R[1] <= 1'b0;
end

assign DPI_STS[0] = DPI_STS_R[0];
assign DPI_STS[1] = DPI_STS_R[1];

always @(posedge DESCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      shift_reg <= 0;
   else if (!lsr_rstn)
      shift_reg <= 0;
   else
      shift_reg <= {DPI_N_reg, DPI_P, shift_reg[7:2]};

always @(posedge DESCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      rstn_dly <= 0;
   else if (!lsr_rstn)
      rstn_dly <= 0;
   else      
      rstn_dly <= 1'b1;

assign SLIP_d_rising_p = 1'b0;

always @(posedge DESCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      cnt <= 0;
   else if (!lsr_rstn)
      cnt <= 0;      
   else begin
      if (~SLIP_d_rising_p) begin
         if (cnt == 6)
            cnt <= 0;
         else
            cnt <= cnt + 1;
      end
   end

assign capture_en_0 = cnt == 3;
assign capture_en_1 = cnt == 6;

always @(posedge DESCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      capture_reg <= 0;
   else if (!lsr_rstn)
      capture_reg <= 0;
   else if (capture_en_0)
      capture_reg <= shift_reg[7:1];
   else if (capture_en_1)
      capture_reg <= {DPI_P, shift_reg[7:2]};
      
always @(posedge RCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      Q_reg <= 0;
   else if (!lsr_rstn)
      Q_reg <= 0;
   else
      Q_reg <= capture_reg;      

assign Q = Q_reg;
//synthesis translate_on

endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_LUT6.v
//
// Functional description: 6-input Look-Up-Table
//
// Parameter description:
//      INIT: init value
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_LUT6
#(
    parameter [63:0] INIT = 64'h0000_0000_0000_0000
) (
    output wire Z,
    input wire I0, I1, I2, I3, I4, I5
);

    wire z5a, z5b;

    GTP_LUT5 #(.INIT(INIT[31:0]))
        l5a (.I0(I0), .I1(I1), .I2(I2), .I3(I3), .I4(I4), .Z(z5a));

    GTP_LUT5 #(.INIT(INIT[63:32]))
        l5b (.I0(I0), .I1(I1), .I2(I2), .I3(I3), .I4(I4), .Z(z5b));

    GTP_MUX2LUT6 mxl6 (.I0(z5a), .I1(z5b), .S(I5), .Z(Z));

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_GRS.v
//
// Functional description: Global reset/set
//
// Parameter description:
//
// Port description:
//
// Revision:
//    06/18/14 - Initial version.
//    03/23/19 - add global signal
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_GRS
(
    input wire GRS_N
);
////////////////GTP_I2C/////////////////
    wire            i2c0_scl_i      ;
    wire            i2c0_scl_o      ;
    wire            i2c0_sda_i      ;
    wire            i2c0_sda_o      ;
    wire            irq_i2c0        ;
    wire            i2c1_scl_i      ;
    wire            i2c1_scl_o      ;
    wire            i2c1_sda_i      ;
    wire            i2c1_sda_o      ;
    wire            irq_i2c1        ;

////////////////GTP_POWERCTL//////////////
    wire            clk_pctl;
    wire            rstn_pctl;
    wire            spi_wakeup_pctl;
    wire            i2c0_wakeup_pctl;
    wire            i2c1_wakeup_pctl;

////////////////GTP_SPI/////////////////
    wire            spi_ss_i_n      ;
    wire    [7:0]   spi_ss_o_n      ;
    wire            spi_sck_oe_n    ;
    wire            spi_sck_i       ;
    wire            spi_sck_o       ;
    wire            spi_mosi_oe_n   ;
    wire            spi_mosi_i      ;
    wire            spi_mosi_o      ;
    wire            spi_miso_oe_n   ;
    wire            spi_miso_i      ;
    wire            spi_miso_o      ;
    wire            irq_spi         ;

////////////////GTP_TIMER/////////////////
    wire            timer_rstn      ;
    wire            timer_clk       ;
    wire            timer_stamp     ;
    wire            timer_pwm       ;
    wire            irq_timer       ;

///////////////////PLL////////////////////
    wire    [7:0]   pll0_prdata     ;
    wire            pll0_pready     ;
    wire    [7:0]   pll1_prdata     ;
    wire            pll1_pready     ;

    wire GRSNET;

    assign GRSNET = GRS_N;

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2016 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Date(08/02/2019) Author:dfpu
//
// GTP model of APML device
//
// History:
//      initial version 
//
//////////////////////////////////////////////////////////////////////////////
`timescale 1ns/1ps

`define assert(condition, message) \
        if (!(condition)) begin \
            $display($realtime, "ERROR: ASSERTION FAILED in %s, line %d: %s", `__FILE__, `__LINE__, message); \
            $finish; \
        end
// module declaration
module GTP_APM_E2 #(

    parameter GRS_EN = "TRUE",  //"TRUE","FALSE",enable global reset
    parameter USE_POSTADD = 0, //enable postadder 0/1
    parameter USE_PREADD = 0,  //enable preadder 0/1
    parameter PREADD_REG = 0,  //preadder reg 0/1

    parameter X_REG = 0,  //X input reg 0/1/2/3
    parameter CXO_REG = 0, //X cascade out reg latency, 0/1/2/3
    parameter XB_REG = 0,  //XB input reg 0/1
    parameter Y_REG = 0,  //Y input reg 0/1/2/3
    parameter Z_REG = 0,  //Z input reg 0/1
    parameter MULT_REG = 0,  //multiplier reg 0/1
    parameter P_REG = 0,  //post adder reg 0/1
    parameter MODEY_REG = 0,  //MODEY reg
    parameter MODEZ_REG = 0,  //MODEZ reg
    parameter MODEIN_REG = 0,  //MODEZ reg

    parameter X_SEL = 0,  // mult X input select X/CXI
    parameter XB_SEL = 0, //X back propagate mux select. 0/1/2/3
    parameter ASYNC_RST = 0,  // RST is sync/async
    parameter USE_SIMD = 0,   // single addsub25_mult25_add48 / dual addsub12_mult12_add24
    parameter [47:0] P_INIT0 = {48{1'b0}},  //P constant input0 (RTI parameter in APM of PG family)
    parameter [47:0] P_INIT1 = {48{1'b0}},  //P constant input1 (RTI parameter in APM of PG family)
    parameter ROUNDMODE_SEL = 0,  //round mode selection

    parameter CPO_REG = 0, // CPO,COUT use register output
    parameter USE_ACCLOW = 0, // accumulator use lower 18-bit feedback only
    parameter CIN_SEL = 0 // select CIN for postadder carry in

)(
    output [47:0] P,
    output [47:0] CPO, //p cascade output
    output COUT,
    output [29:0] CXO, //x cascade output
    output [24:0] CXBO, //x backward cascade output

    input [29:0] X,
    input [29:0] CXI, //x cascade input
    input [24:0] CXBI, //x backward cascade input
    input [24:0] XB, //x backward cascade input
    input [17:0] Y,
    input [47:0] Z,
    input [47:0] CPI, //p cascade input
    input CIN,
    input [2:0] MODEY,
    input [3:0] MODEZ,
    input [4:0] MODEIN,

    input CLK,

    input  CEX1,  //X1 enable signals 
    input  CEX2,  //X2 enable signals 
    input  CEX3,  //X3 enable signals 
    input  CEXB,  //XB enable signals 
    input  CEY1,  //Y1 enable signals 
    input  CEY2,  //Y2 enable signals 
    input  CEZ,  //Z enable signals 
    input  CEPRE,  //PRE enable signals 
    input  CEM,  //M enable signals 
    input  CEP,  //P enable signals 
    input  CEMODEY,  //MODEY enable signals 
    input  CEMODEZ,  //MODEZ enable signals 
    input  CEMODEIN,  //MODEIN enable signals 

    input  RSTX, //X reset signals 
    input  RSTXB, //XB reset signals 
    input  RSTY, //Y reset signals 
    input  RSTZ, //Z reset signals 
    input  RSTPRE, //PRE reset signals 
    input  RSTM, //M reset signals 
    input  RSTP, //P reset signals 
    input  RSTMODEY, //MODEY reset signals 
    input  RSTMODEZ, //MODEZ reset signals 
    input  RSTMODEIN //MODEIN reset signals 

);

    wire grs;
    assign grs = (GRS_EN == "TRUE") ? !GRS_INST.GRSNET : 1'b0;

//rst selection

    assign arst_x = (ASYNC_RST == 1'b1) ? (RSTX | grs) : grs;
    assign arst_xb = (ASYNC_RST == 1'b1) ? (RSTXB | grs) : grs;
    assign arst_y = (ASYNC_RST == 1'b1) ? (RSTY | grs) : grs;
    assign arst_z = (ASYNC_RST == 1'b1) ? (RSTZ | grs) : grs;
    assign arst_pre = (ASYNC_RST == 1'b1) ? (RSTPRE | grs) : grs;
    assign arst_m = (ASYNC_RST == 1'b1) ? (RSTM | grs) : grs;
    assign arst_p = (ASYNC_RST == 1'b1) ? (RSTP | grs) : grs;
    assign arst_modey = (ASYNC_RST == 1'b1) ? (RSTMODEY | grs) : grs;
    assign arst_modez = (ASYNC_RST == 1'b1) ? (RSTMODEZ | grs) : grs;
    assign arst_modein = (ASYNC_RST == 1'b1) ? (RSTMODEIN | grs) : grs;

    assign srst_x = (ASYNC_RST == 1'b1) ? 1'b0 : RSTX;
    assign srst_xb = (ASYNC_RST == 1'b1) ? 1'b0 : RSTXB;
    assign srst_y = (ASYNC_RST == 1'b1) ? 1'b0 : RSTY;
    assign srst_z = (ASYNC_RST == 1'b1) ? 1'b0 : RSTZ;
    assign srst_pre = (ASYNC_RST == 1'b1) ? 1'b0 : RSTPRE;
    assign srst_m = (ASYNC_RST == 1'b1) ? 1'b0 : RSTM;
    assign srst_p = (ASYNC_RST == 1'b1) ? 1'b0 : RSTP;
    assign srst_modey = (ASYNC_RST == 1'b1) ? 1'b0 : RSTMODEY;
    assign srst_modez = (ASYNC_RST == 1'b1) ? 1'b0 : RSTMODEZ;
    assign srst_modein = (ASYNC_RST == 1'b1) ? 1'b0 : RSTMODEIN;
    // input registers

    wire [29:0] xsel_out;
    reg [29:0] x1,x2,x3; // x register latency 
    reg [29:0] sh_xo;
    //x cascade output bus
    assign xsel_out = X_SEL ? CXI[29:0] : X[29:0];
    always @(posedge CLK or posedge arst_x) 
    begin
        if (arst_x) begin
            x1 <= 30'b0;
        end else if (srst_x) begin
            x1 <= 30'b0;
        end else if (CEX1) begin
            x1 <= xsel_out;
            end
    end

    always @(posedge CLK or posedge arst_x) 
    begin
        if (arst_x ) begin
            x2 <= 30'b0;
        end else if (srst_x) begin
            x2 <= 30'b0;
        end else if (CEX2) begin
            x2 <= x1;
            end
    end

    always @(posedge CLK or posedge arst_x) 
    begin
        if (arst_x ) begin
            x3 <= 30'b0;
        end else if (srst_x) begin
            x3 <= 30'b0;
        end else if (CEX3) begin
            x3 <= x2;
            end
    end

    always @ (*) begin
        case(CXO_REG[1:0])
            2'b00 : sh_xo = xsel_out;
            2'b01 : sh_xo = x1;
            2'b10 : sh_xo = x2;
            2'b11 : sh_xo = x3;
        endcase
    end

    assign CXO = sh_xo;

    wire [29:0] xir_out0,xir_out1; //registered (optional) x internal bus
    wire [29:0] x_post;
    wire [24:0] xir_out2,xir_out3;
    wire [4:0] modeini; //registered (optional) INMODE internal
    assign xir_out0 = X_REG[0] ? x1 : xsel_out; 
    assign xir_out1 = X_REG[1] ? x2 : xir_out0; 
    assign x_post = xir_out1;
    assign xir_out2 = modeini[0] ? x1[24:0] : xir_out1[24:0];
    assign xir_out3 = modeini[1] ? xir_out2 : 25'b0; 

    wire [24:0] xbi; //registered (optional) xb internal
    reg [24:0] xbr;
    wire [24:0] xb_in;
    assign xb_in = XB_SEL[0] ? CXBI[24:0] : XB[24:0];
    always @(posedge CLK or posedge arst_xb)
    begin
        if (arst_xb) begin
            xbr[24:0] <= 25'b0;
        end else if (srst_xb) begin
            xbr[24:0] <= 25'b0;
        end else if (CEXB) begin
            xbr[24:0] <= xb_in;
            end
    end

    assign xbi[24:0] = (XB_REG == 1) ? xbr : xb_in;


    reg [17:0] yi; //registered (optional) y internal
    reg [17:0] yr1,yr2;
    always @(posedge CLK or posedge arst_y)
    begin
        if (arst_y) begin
            yr1[17:0] <= 18'b0;
        end else if (srst_y) begin
            yr1[17:0] <= 18'b0;
        end else if (CEY1) begin
            yr1[17:0] <= Y;
            end
    end

    always @(posedge CLK or posedge arst_y)
    begin
        if (arst_y) begin
            yr2[17:0] <= 18'b0;
        end else if (srst_y) begin
            yr2[17:0] <= 18'b0;
        end else if (CEY2) begin
            yr2[17:0] <= yr1;
            end
    end

    always @ (*) begin
        case(Y_REG[1:0])
            2'b00 : yi = Y;
            2'b01 : yi = yr1;
            2'b10 : yi = yr1;
            2'b11 : yi = yr2;
        endcase
    end

    wire [17:0] y_post;
    assign y_post = yi;
    wire [17:0] yi_out;
    assign yi_out = modeini[4] ? yr1 : yi; 

    wire [47:0] zi; //registered (optional) z internal
    reg [47:0] zr;
    always @(posedge CLK or posedge arst_z)
    begin
        if (arst_z) begin
            zr[47:0] <= 48'b0;
        end else if (srst_z) begin
            zr[47:0] <= 48'b0;
        end else if (CEZ) begin
            zr[47:0] <= Z;
            end
    end
    
    assign zi = (Z_REG == 1'b1) ? zr : Z;

    wire [2:0] modeyi; //registered (optional) MODEY internal
    wire [3:0] modezi; //registered (optional) MODEZ internal
    reg [2:0] modeyr; //registered (optional) MODEY internal
    reg [3:0] modezr; //registered (optional) MODEZ internal
    
    always @(posedge CLK or posedge arst_modey)
    begin
        if (arst_modey) begin
            modeyr[2:0] <= 3'b0;
        end else if (srst_modey) begin
            modeyr[2:0] <= 3'b0;
        end else if (CEMODEY) begin
            modeyr[2:0] <= MODEY;
            end
    end
    
    assign modeyi = (MODEY_REG == 1'b1) ? modeyr : MODEY;

    always @(posedge CLK or posedge arst_modez)
    begin
        if (arst_modez) begin
            modezr[3:0] <= 4'b0;
        end else if (srst_modez) begin
            modezr[3:0] <= 4'b0;
        end else if (CEMODEZ) begin
            modezr[3:0] <= MODEZ;
            end
    end
    
    assign modezi = (MODEZ_REG == 1'b1) ? modezr : MODEZ;

    reg [4:0] modeinr;
    always @(posedge CLK or posedge arst_modein)
    begin
        if (arst_modein) begin
            modeinr[4:0] <= 5'b0;
        end else if (srst_modein) begin
            modeinr[4:0] <= 5'b0;
        end else if (CEMODEIN) begin
            modeinr[4:0] <= MODEIN;
            end
    end

    assign modeini = (MODEIN_REG == 1'b1) ? modeinr : MODEIN;

    //preadder

    reg [24:0] xbv;
    always @ (*) begin
        case(XB_SEL[1])
            1'b0 : xbv = xbi;
            1'b1 : xbv = sh_xo[24:0];
        endcase
    end

    assign CXBO = xbv;

    wire [24:0] prec; //cominational preadder output
    wire [24:0] pre_a,pre_b;
    wire preadd_sub;
    wire [24:0] preadd_s;
    wire [11:0] preadd_s_h,preadd_s_l;

    assign pre_a = xir_out3;
    assign pre_b = modeini[2] ? xbv: 25'b0;
    assign preadd_sub = modeini[3];
    assign preadd_s = preadd_sub ? pre_a - pre_b : pre_a + pre_b;
    assign preadd_s_l = preadd_sub ? pre_a[11:0] - pre_b[11:0] : pre_a[11:0] + pre_b[11:0];
    assign preadd_s_h = preadd_sub ? pre_a[23:12] - pre_b[23:12] : pre_a[23:12] + pre_b[23:12];
    assign prec = (USE_SIMD == 1'b1) ? {preadd_s_h[11],preadd_s_h,preadd_s_l} : preadd_s;
    
    reg [24:0] prer;
    always @(posedge CLK or posedge arst_pre)
    begin
        if (arst_pre) begin
            prer[24:0] <= 25'b0;
        end else if (srst_pre) begin
            prer[24:0] <= 25'b0;
        end else if (CEPRE) begin
            prer[24:0] <= prec;
            end
    end

    wire [24:0] prei; //registered (optional) preadder output
    assign prei = (PREADD_REG == 1'b1) ? prer : prec;

    // multiplier
    wire [47:0] mc; //mult combinational output
    wire [24:0] mult_ina;
    wire [17:0] mult_inb;
    wire [47:0] mult_out_s;
    wire [23:0] mult_out_h, mult_out_l;
    assign mult_ina[24:0] = USE_PREADD ? prei[24:0] : xir_out3[24:0];
    assign mult_inb[17:0] = yi_out[17:0];
    assign mult_out_s = {{23{mult_ina[24]}},mult_ina} * {{30{mult_inb[17]}},mult_inb};
    assign mult_out_l = {{12{mult_ina[11]}},mult_ina[11:0]} * {{15{mult_inb[8]}},mult_inb[8:0]};
    assign mult_out_h = {{12{mult_ina[23]}},mult_ina[23:12]} * {{15{mult_inb[17]}},mult_inb[17:9]};

    assign mc = (USE_SIMD == 1'b1) ? {mult_out_h,mult_out_l}: mult_out_s;

    wire [47:0] mi; //registered (optional) mult internal output
    reg [47:0] mr;
    always @(posedge CLK or posedge arst_m)
    begin
        if (arst_m) begin
            mr[47:0] <= 48'b0;
        end else if (srst_m) begin
            mr[47:0] <= 48'b0;
        end else if (CEM) begin
            mr[47:0] <= mc;
            end
    end

    assign mi = (MULT_REG == 1'b1) ? mr : mc;

    //post adder
    reg  [47:0] pyi; // post adder input a before inverter
    wire [47:0] py = modeyi[2] ? ~pyi : pyi; // post adder input a after inverter
    reg  [47:0] pzi; // post adder input b before inverter
    wire [47:0] pz = modezi[3] ? ~pzi : pzi; // post adder input b after inverter

    reg [48:0] pr; // post adder regstered feedback
    wire [47:0] pri =  USE_ACCLOW ? { {31{1'b0}}, pr[16:0] } : pr[47:0];//post adder lower portion feedback

    always @ (*) begin
        case(modeyi[1:0])
            2'b00 : pyi = 48'b0;
            2'b01 : pyi = mi;
            2'b10 : pyi = pri;
            2'b11 : pyi = {x_post[29:0],y_post[17:0]};
        endcase
    end

    always @(*) begin
        case(modezi[2:0])
            3'b000 : pzi = 48'b0;
            3'b001 : pzi = pri;
            3'b010 : pzi = zi;
            3'b011 : pzi = $signed(CPI); //both branch need $signed
            3'b100 : pzi = $signed(CPI) >>> 17; //both branch need $signed
            3'b101 : pzi = $signed(CPI) >>> 24; //both branch need $signed
            3'b110 : pzi = $signed(CPI) >>> 16; //both branch need $signed
            3'b111 : pzi = $signed(CPI) >>> 8; //both branch need $signed
        endcase
    end

    wire cinv;
    assign cinv = CIN_SEL ? CIN : modeyi[2] | modezi[3];

    wire [48:0] pc;
    wire [47:0] alu_out;
    wire cout_inter0;
    wire cout_inter1;
    wire cin_inter;
    wire [47:0] c_inter;
    wire post_select;

    assign post_select = ((modeyi[1:0] == 2'b00) && (modezi[2:0] == 3'b000));
    assign {cout_inter0,alu_out[23:0]} = py[23:0] + pz[23:0] + cinv;
    assign cin_inter = USE_SIMD ? cinv : cout_inter0;
    assign {cout_inter1,alu_out[47:24]} = py[47:24] + pz[47:24] + cin_inter;
    assign c_inter = (ROUNDMODE_SEL ? alu_out[47] : (post_select ? 1'b1 : 1'b0)) ? P_INIT1 : P_INIT0;
    assign pc = {cout_inter1,alu_out[47:0]} + c_inter[47:0] ;



    wire [47:0] pi;
    always @(posedge CLK or posedge arst_p)
    begin
        if (arst_p) begin
            pr[48:0] <= 49'b0;
        end else if (srst_p) begin
            pr[48:0] <= 49'b0;
        end else if (CEP) begin
            pr[48:0] <= pc[48:0];
            end
    end

    assign pi = (P_REG == 1'b1) ? pr[47:0] : pc[47:0];

    assign P = USE_POSTADD ? pi : mi;
    assign CPO = USE_POSTADD ? (CPO_REG ? pr[47:0] : pc[47:0]) : mi;

    assign COUT = CPO_REG ? pr[48] : pc[48];
// DRC check
// pragma translate_off
    initial begin
        `assert(X_REG <= 3, "X_REG <= 3")
        `assert(CXO_REG <= 3, "CXO_REG <= 3")
        `assert(XB_REG <= 1, "XB_REG <= 1")
        `assert(Y_REG <= 3, "Y_REG <= 3")
        `assert(Z_REG <= 1, "Z_REG <= 1")
        `assert(MULT_REG <= 1, "MULT_REG <= 1")
        `assert(P_REG <= 1, "P_REG <= 1")
        `assert(PREADD_REG <= 1, "PREADD_REG <= 1")
        `assert(MODEY_REG <= 1, "MODEY_REG <= 1")
        `assert(MODEZ_REG <= 1, "MODEZ_REG <= 1")
        `assert(MODEIN_REG <= 1, "MODEIN_REG <= 1")
    end
// pragma translate_on
    

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2016 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_RAM128X1SP.v
//
// Functional description: single-port 128x1 distributed ram
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_RAM128X1SP
#(
    parameter [127:0] INIT = 128'h0000_0000_0000_0000_0000_0000_0000_0000
) (
    output  DO,
    input   DI,
    input [6:0] ADDR,
    input WCLK,
    input WE
);
//synthesis translate_off
    reg [127:0] mem ;

    initial begin
        mem = INIT;
    end

    always @(posedge WCLK) begin
        if (WE == 1'b1) begin
            mem[ADDR] <= DI;
        end
    end

    assign DO = mem[ADDR];
//synthesis translate_on
endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_DRM18K_E1.v
//
// Functional description:
// Fake module
//
// Parameter  description:
//
// Port description:
//
// Revision history:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_DRM18K_E1
#(
    parameter GRS_EN = "TRUE",
    parameter integer DATA_WIDTH_A = 18,
    parameter integer DATA_WIDTH_B = 18,
    parameter WRITE_MODE_A = "NORMAL_WRITE",
    parameter WRITE_MODE_B = "NORMAL_WRITE",
    parameter integer DOA_REG = 0,
    parameter integer DOB_REG = 0,
    parameter integer DOA_REG_CLKINV = 0,
    parameter integer DOB_REG_CLKINV = 0,
    parameter [17:0] RSTA_VAL = 18'b0,
    parameter [17:0] RSTB_VAL = 18'b0,
    parameter RST_TYPE = "SYNC",
    parameter RAM_MODE = "TRUE_DUAL_PORT",
    parameter [287:0] INIT_00 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_01 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_02 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_03 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_04 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_05 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_06 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_07 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_08 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_09 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_10 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_11 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_12 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_13 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_14 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_15 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_16 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_17 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_18 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_19 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_20 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_21 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_22 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_23 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_24 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_25 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_26 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_27 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_28 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_29 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_2A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_2B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_2C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_2D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_2E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_2F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_30 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_31 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_32 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_33 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_34 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_35 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_36 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_37 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_38 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_39 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_3A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_3B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_3C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_3D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_3E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_3F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_FILE = "NONE",
    parameter integer BLOCK_X = 0,
    parameter integer BLOCK_Y = 0,
    parameter integer RAM_DATA_WIDTH = 9,
    parameter integer RAM_ADDR_WIDTH = 11,
    parameter INIT_FORMAT = "BIN"
) (
    output [17:0] DOA,
    output [17:0] DOB,
    input  [17:0] DIA,
    input  [17:0] DIB,
    input  [13:0] ADDRA,
    input  [13:0] ADDRB,
    input  ADDRA_HOLD,
    input  ADDRB_HOLD,
    input  [3:0] BWEA,
    input  [1:0] BWEB,
    input  CLKA,
    input  CLKB,
    input  CEA,
    input  CEB,
    input  WEA,
    input  WEB,
    input  ORCEA,
    input  ORCEB,
    input  RSTA,
    input  RSTB
);

    localparam  BLOCK_DEPTH = 2**(DATA_WIDTH_A == 1 ? 14 :
                                  DATA_WIDTH_A == 2 ? 13 :
                                  DATA_WIDTH_A == 4 ? 12 :
                                  DATA_WIDTH_A <= 9 ? 11 :
                                  DATA_WIDTH_A <= 18 ? 10 : 9);

    localparam  BLOCK_WIDTH =   DATA_WIDTH_A;             //block memory data width

    localparam MEM_SIZE = 18432;
    localparam width_a = (DATA_WIDTH_A == 32) ? 16 : (DATA_WIDTH_A == 36) ? 18 : DATA_WIDTH_A;
    localparam width_b = (DATA_WIDTH_B == 32) ? 16 : (DATA_WIDTH_B == 36) ? 18 : DATA_WIDTH_B;

    integer  cnt;
    reg [9-1:0] mem [MEM_SIZE/9-1:0];

    reg [13:0] ada_reg = 14'b0, adb_reg = 14'b0;
    reg [17:0] da_reg = 9'b0, db_reg = 9'b0;
    reg wea_reg = 1'b0, web_reg = 1'b0;
    reg [3:0] bea_reg;
    reg [1:0] beb_reg;
    wire write_en_a, write_en_b, read_en_a, read_en_b;

    reg [17:0] a_out;
    reg [17:0] a_out_reg;
    reg [17:0] b_out;
    reg [17:0] b_out_reg;

    wire grs, rsta_grs, rstb_grs;
    wire rsta_grs_sync;
    wire rstb_grs_sync;
    wire rsta_grs_async;
    wire rstb_grs_async;
    
    reg [17:0] doa,doa_reg,doa_mux;
    reg [17:0] dob,dob_reg,dob_mux;


    wire CLKA_for_or,CLKB_for_or;
    wire rsta_int,rstb_int;

    wire [17:0] rsta_val_int;
    wire [17:0] rstb_val_int;

    assign rsta_val_int = (DATA_WIDTH_A==16 | DATA_WIDTH_B == 32)? {2'b00,RSTA_VAL[16:9],RSTA_VAL[7:0]}:RSTA_VAL;
    assign rstb_val_int = (DATA_WIDTH_B==16 | DATA_WIDTH_B == 32)? {2'b00,RSTB_VAL[16:9],RSTB_VAL[7:0]}:RSTB_VAL;

    initial begin
        #1;
        doa = RSTA_VAL;
        dob = RSTB_VAL;
        doa_reg = RSTA_VAL;
        dob_reg = RSTB_VAL;
        doa_mux = RSTA_VAL;
        dob_mux = RSTB_VAL;
        a_out = rsta_val_int;
        a_out_reg = rsta_val_int;
        b_out = rstb_val_int;
        b_out_reg = rstb_val_int;
    end

// synthesis translate_off

   reg [RAM_DATA_WIDTH-1:0] ini_mem [2**RAM_ADDR_WIDTH-1:0];
   integer p;
   initial
   begin
      if(INIT_FILE != "NONE")
      begin
          if(INIT_FORMAT == "BIN")
              $readmemb(INIT_FILE,ini_mem);
          else
              $readmemh(INIT_FILE,ini_mem);
          for(p=0;p<20;p=p+1)
              $display("ini_mem[%d] = %b",p,ini_mem[p]);
      end
   end
///////////////////
// parameter check
///////////////////
    initial begin
        case (DATA_WIDTH_A)
            1, 2, 4, 8, 16, 32: begin
                case (DATA_WIDTH_B)
                    1, 2, 4, 8, 16, 32:  ; //null
                    default: begin
                        $display("ERROR: GTP_DRM18K_E1 instance %m parameter DATA_WIDTH_B:%d is illegal. The legal values are 1,2,4,8,16 or 32.",DATA_WIDTH_B);
                        $finish;
                    end
                endcase
            end
            9, 18, 36: begin
                case (DATA_WIDTH_B)
                    9, 18, 36:    ; //null
                    default: begin
                        $display("ERROR: GTP_DRM18K_E1 instance %m parameter DATA_WIDTH_B:%d is illegal. The legal values are 9, 18 or 36.",DATA_WIDTH_B);
                        $finish;
                    end
                endcase
            end
            default: begin
                $display("ERROR: GTP_DRM18K_E1 instance %m parameter DATA_WIDTH_A:%d is illegal. The legal values are 1,2,4,8,9,16,18,32 or 36.",DATA_WIDTH_A);
                $finish;
            end
        endcase

        case (WRITE_MODE_A)
            "NORMAL_WRITE",
            "TRANSPARENT_WRITE",
            "READ_BEFORE_WRITE":    ; //null 
            default: begin
                $display("ERROR: GTP_DRM18K_E1 instance %m parameter WRITE_MODE_A: %s is illegal. The legal values are NORMAL_WRITE,TRANSPARENT_WRITE or READ_BEFORE_WRITE.", WRITE_MODE_A);
                $finish;
            end
        endcase

        case (WRITE_MODE_B)
            "NORMAL_WRITE",
            "TRANSPARENT_WRITE",
            "READ_BEFORE_WRITE":    ; //null  
            default: begin
                $display("ERROR: GTP_DRM18K_E1 instance %m parameter WRITE_MODE_B: %s is illegal. The legal values are NORMAL_WRITE,TRANSPARENT_WRITE or READ_BEFORE_WRITE.", WRITE_MODE_B);
                $finish;
            end
        endcase

        case (DOA_REG)
            0,1:     ;//null
            default: begin
                $display("ERROR: GTP_DRM18K_E1 instance %m parameter DOA_REG: %s is illegal. The legal values are 0 or 1.", DOA_REG);
                $finish;
            end
        endcase

        case (DOB_REG)
            0,1:     ;//null
            default: begin
                $display("ERROR: GTP_DRM18K_E1 instance %m parameter DOB_REG: %s is illegal. The legal values are 0 or 1.", DOB_REG);
                $finish;
            end
        endcase

        case (DOA_REG_CLKINV)
            0,1:     ;//null
            default: begin
                $display("ERROR: GTP_DRM18K_E1 instance %m parameter DOA_REG_CLKINV: %s is illegal. The legal values are 0 or 1.", DOA_REG_CLKINV);
                $finish;
            end
        endcase

        case (DOB_REG_CLKINV)
            0,1:     ;//null
            default: begin
                $display("ERROR: GTP_DRM18K_E1 instance %m parameter DOB_REG_CLKINV: %s is illegal. The legal values are 0 or 1.", DOB_REG_CLKINV);
                $finish;
            end
        endcase

        case (RST_TYPE)
            "ASYNC",
            "SYNC":     ;//null
            default: begin
                $display("ERROR: GTP_DRM18K_E1 instance %m parameter RST_TYPE: %s is illegal. The legal values are ASYNC or SYNC.", RST_TYPE);
                $finish;
            end
        endcase

        case (RAM_MODE)
            "ROM",
            "SINGLE_PORT":      ;//null
            "SIMPLE_DUAL_PORT": begin
                if (DATA_WIDTH_A < 32 && WRITE_MODE_A != "NORMAL_WRITE") begin
                    $display("Warrning: GTP_DRM18K_E1 instance %m suggest to use TRUE_DUAL_PORT RAM_MODE if DATA_WIDTH_A and WRITE_MODE_A: %d,%s.",DATA_WIDTH_A,WRITE_MODE_A);
                end
            end
            "TRUE_DUAL_PORT": begin
                if (DATA_WIDTH_A > 18 || DATA_WIDTH_B > 18) begin
                    $display("ERROR: GTP_DRM18K_E1 instance %m parameter DATA_WIDTH_A and DATA_WIDTH_B in TRUE_DUAL_PORT MODE:%d,%d is illegal. The legal values are 1,2,4,8,9,16 or 18.",DATA_WIDTH_A,DATA_WIDTH_B);
                    $finish;
                end
            end
            default: begin
                $display("ERROR: GTP_DRM18K_E1 instance %m parameter RAM_MODE value: %s is illegal. The legal values are ROM or SINGLE_PORT, SIMPLE_DUAL_PORT or TRUE_DUAL_PORT.", RAM_MODE);
                $finish;
            end
        endcase
        
    end

/////////////////
// initialization
/////////////////

    initial begin
        if (INIT_FILE == "NONE") begin
            for (cnt = 0; cnt < 32; cnt = cnt + 1) begin
                mem[32*0 + cnt] = INIT_00[cnt*9 +: 9];
                mem[32*1 + cnt] = INIT_01[cnt*9 +: 9];
                mem[32*2 + cnt] = INIT_02[cnt*9 +: 9];
                mem[32*3 + cnt] = INIT_03[cnt*9 +: 9];
                mem[32*4 + cnt] = INIT_04[cnt*9 +: 9];
                mem[32*5 + cnt] = INIT_05[cnt*9 +: 9];
                mem[32*6 + cnt] = INIT_06[cnt*9 +: 9];
                mem[32*7 + cnt] = INIT_07[cnt*9 +: 9];
                mem[32*8 + cnt] = INIT_08[cnt*9 +: 9];
                mem[32*9 + cnt] = INIT_09[cnt*9 +: 9];
                mem[32*10 + cnt] = INIT_0A[cnt*9 +: 9];
                mem[32*11 + cnt] = INIT_0B[cnt*9 +: 9];
                mem[32*12 + cnt] = INIT_0C[cnt*9 +: 9];
                mem[32*13 + cnt] = INIT_0D[cnt*9 +: 9];
                mem[32*14 + cnt] = INIT_0E[cnt*9 +: 9];
                mem[32*15 + cnt] = INIT_0F[cnt*9 +: 9];
                mem[32*16 + cnt] = INIT_10[cnt*9 +: 9];
                mem[32*17 + cnt] = INIT_11[cnt*9 +: 9];
                mem[32*18 + cnt] = INIT_12[cnt*9 +: 9];
                mem[32*19 + cnt] = INIT_13[cnt*9 +: 9];
                mem[32*20 + cnt] = INIT_14[cnt*9 +: 9];
                mem[32*21 + cnt] = INIT_15[cnt*9 +: 9];
                mem[32*22 + cnt] = INIT_16[cnt*9 +: 9];
                mem[32*23 + cnt] = INIT_17[cnt*9 +: 9];
                mem[32*24 + cnt] = INIT_18[cnt*9 +: 9];
                mem[32*25 + cnt] = INIT_19[cnt*9 +: 9];
                mem[32*26 + cnt] = INIT_1A[cnt*9 +: 9];
                mem[32*27 + cnt] = INIT_1B[cnt*9 +: 9];
                mem[32*28 + cnt] = INIT_1C[cnt*9 +: 9];
                mem[32*29 + cnt] = INIT_1D[cnt*9 +: 9];
                mem[32*30 + cnt] = INIT_1E[cnt*9 +: 9];
                mem[32*31 + cnt] = INIT_1F[cnt*9 +: 9];
                mem[32*32 + cnt] = INIT_20[cnt*9 +: 9];
                mem[32*33 + cnt] = INIT_21[cnt*9 +: 9];
                mem[32*34 + cnt] = INIT_22[cnt*9 +: 9];
                mem[32*35 + cnt] = INIT_23[cnt*9 +: 9];
                mem[32*36 + cnt] = INIT_24[cnt*9 +: 9];
                mem[32*37 + cnt] = INIT_25[cnt*9 +: 9];
                mem[32*38 + cnt] = INIT_26[cnt*9 +: 9];
                mem[32*39 + cnt] = INIT_27[cnt*9 +: 9];
                mem[32*40 + cnt] = INIT_28[cnt*9 +: 9];
                mem[32*41 + cnt] = INIT_29[cnt*9 +: 9];
                mem[32*42 + cnt] = INIT_2A[cnt*9 +: 9];
                mem[32*43 + cnt] = INIT_2B[cnt*9 +: 9];
                mem[32*44 + cnt] = INIT_2C[cnt*9 +: 9];
                mem[32*45 + cnt] = INIT_2D[cnt*9 +: 9];
                mem[32*46 + cnt] = INIT_2E[cnt*9 +: 9];
                mem[32*47 + cnt] = INIT_2F[cnt*9 +: 9];
                mem[32*48 + cnt] = INIT_30[cnt*9 +: 9];
                mem[32*49 + cnt] = INIT_31[cnt*9 +: 9];
                mem[32*50 + cnt] = INIT_32[cnt*9 +: 9];
                mem[32*51 + cnt] = INIT_33[cnt*9 +: 9];
                mem[32*52 + cnt] = INIT_34[cnt*9 +: 9];
                mem[32*53 + cnt] = INIT_35[cnt*9 +: 9];
                mem[32*54 + cnt] = INIT_36[cnt*9 +: 9];
                mem[32*55 + cnt] = INIT_37[cnt*9 +: 9];
                mem[32*56 + cnt] = INIT_38[cnt*9 +: 9];
                mem[32*57 + cnt] = INIT_39[cnt*9 +: 9];
                mem[32*58 + cnt] = INIT_3A[cnt*9 +: 9];
                mem[32*59 + cnt] = INIT_3B[cnt*9 +: 9];
                mem[32*60 + cnt] = INIT_3C[cnt*9 +: 9];
                mem[32*61 + cnt] = INIT_3D[cnt*9 +: 9];
                mem[32*62 + cnt] = INIT_3E[cnt*9 +: 9];
                mem[32*63 + cnt] = INIT_3F[cnt*9 +: 9];
            end
        end
        else  begin      // INIT_FILE 
            case(DATA_WIDTH_A)
                1: begin  //DRM TYPE 16K*1
                   for(cnt=0; cnt<2*1024;cnt = cnt+1)
                       mem[cnt][7:0] = {ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*8+7][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*8+6][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*8+5][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*8+4][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*8+3][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*8+2][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*8+1][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*8][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH]};
                end
                2: begin //DRM TYPE 8K*2
                   for(cnt=0; cnt<2*1024;cnt = cnt+1)
                       mem[cnt][7:0] = {ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*4+3][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*4+2][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*4+1][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                        ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*4][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH]};
                end
                4: begin //DRM TYPE 4K*4
                   for(cnt=0; cnt<2*1024;cnt = cnt+1)
                       {mem[cnt][7:0]} = {ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*2+1][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH],
                                          ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt*2][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH]};
                end
                8: begin //DRM TYPE 2K*8
                   for(cnt=0; cnt<2*1024;cnt = cnt+1)
                       mem[cnt][7:0] = ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH];
                end
                9: begin //DRM TYPE 2K*9
                   for(cnt=0; cnt<2*1024;cnt = cnt+1)
                       mem[cnt] = ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH];
                end
                16:begin //DRM TYPE 1K*16
                   for(cnt=0; cnt<1024;cnt = cnt+1)
                       {mem[cnt*2+1][7:0], mem[cnt*2][7:0]} = ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH];
                end
                18:begin //DRM TYPE 1K*18
                   for(cnt=0; cnt<1024;cnt = cnt+1)
                       {mem[cnt*2+1], mem[cnt*2]} = ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH];
                end
                32:begin //DRM TYPE 512*32
                   for(cnt=0; cnt<512;cnt = cnt+1)
                       {mem[cnt*4+3][7:0],mem[cnt*4+2][7:0],mem[cnt*4+1][7:0],mem[cnt*4][7:0]} = ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH];
                end
                36:begin //DRM TYPE 512*36
                   for(cnt=0; cnt<512;cnt = cnt+1)
                       {mem[cnt*4+3],mem[cnt*4+2],mem[cnt*4+1],mem[cnt*4]} = ini_mem[BLOCK_Y*BLOCK_DEPTH + cnt][BLOCK_X*BLOCK_WIDTH +:BLOCK_WIDTH];
                end
            endcase
        end
    end

    always @(posedge CLKA) begin
        if (CEA) begin
            // high to hold the address
            if (ADDRA_HOLD == 1'b0) begin
                ada_reg <= ADDRA;
            end
            da_reg <= DIA;
            wea_reg <= WEA;
            bea_reg <= BWEA;
        end
    end

    always @(posedge CLKB) begin
        if (CEB) begin
            // high to hold the address
            if (ADDRB_HOLD == 1'b0) begin
                adb_reg <= ADDRB;
            end
            web_reg <= WEB;
            beb_reg <= BWEB;
        end
    end

    ///////////////////
    // task & function
    ///////////////////

    function [DATA_WIDTH_A-1:0] mem_read_a;
        input [13:0]  addr;
    begin
        case (DATA_WIDTH_A)
            1: mem_read_a = mem[addr[13:3]][addr[2:0]];
            2: mem_read_a = mem[addr[13:3]][addr[2:1]*2 +: 2];
            4: mem_read_a = mem[addr[13:3]][addr[2]*4 +: 4];
            8: mem_read_a = mem[addr[13:3]][7:0];
            9: mem_read_a = mem[addr[13:3]];
            16: mem_read_a = {mem[addr[13:4]*2+1][7:0], mem[addr[13:4]*2][7:0]};
            18: mem_read_a = {mem[addr[13:4]*2+1],      mem[addr[13:4]*2]};
            32: mem_read_a = {mem[addr[13:5]*4+3][7:0], mem[addr[13:5]*4+2][7:0],
                              mem[addr[13:5]*4+1][7:0], mem[addr[13:5]*4][7:0]};
            36: mem_read_a = {mem[addr[13:5]*4+3],      mem[addr[13:5]*4+2],
                              mem[addr[13:5]*4+1],      mem[addr[13:5]*4]};
            default:      ;//null 
        endcase
    end
    endfunction

    function [DATA_WIDTH_B-1:0] mem_read_b;
        input [13:0] addr;
    begin
        case (DATA_WIDTH_B)
            1: mem_read_b = mem[addr[13:3]][addr[2:0]];
            2: mem_read_b = mem[addr[13:3]][addr[2:1]*2 +: 2];
            4: mem_read_b = mem[addr[13:3]][addr[2]*4 +: 4];
            8: mem_read_b = mem[addr[13:3]][7:0];
            9: mem_read_b = mem[addr[13:3]];
            16: mem_read_b = {mem[addr[13:4]*2+1][7:0], mem[addr[13:4]*2][7:0]};
            18: mem_read_b = {mem[addr[13:4]*2+1],      mem[addr[13:4]*2]};
            32: mem_read_b = {mem[addr[13:5]*4+3][7:0], mem[addr[13:5]*4+2][7:0],
                              mem[addr[13:5]*4+1][7:0], mem[addr[13:5]*4][7:0]};
            36: mem_read_b = {mem[addr[13:5]*4+3],      mem[addr[13:5]*4+2],
                              mem[addr[13:5]*4+1],      mem[addr[13:5]*4]};
            default:      ;//null
        endcase
    end
    endfunction

    task mem_write_a;
        input [13:0] addr;
        input [35:0] data;
        input [3:0]  byte_en;
    begin
        case (DATA_WIDTH_A)
            1: mem[addr[13:3]][addr[2:0]] = data[0];
            2: mem[addr[13:3]][addr[2:1]*2 +: 2] = data[1:0];
            4: mem[addr[13:3]][addr[2]*4 +: 4] = data[3:0];
            8: mem[addr[13:3]][7:0] = data[7:0];
            9: mem[addr[13:3]] = data[8:0];
            16: begin
                if (byte_en[1])
                    mem[addr[13:4]*2+1][7:0] = data[16:9];
                if (byte_en[0])
                    mem[addr[13:4]*2][7:0]   = data[7:0];
            end
            18: begin
                if (byte_en[1])
                    mem[addr[13:4]*2+1] = data[17:9];
                if (byte_en[0])
                    mem[addr[13:4]*2]   = data[8:0];
            end
            32: begin
                if (byte_en[3])
                    mem[addr[13:5]*4+3][7:0] = data[34:27];
                if (byte_en[2])
                    mem[addr[13:5]*4+2][7:0] = data[25:18];
                if (byte_en[1])
                    mem[addr[13:5]*4+1][7:0] = data[16:9];
                if (byte_en[0])
                    mem[addr[13:5]*4][7:0]   = data[7:0];
            end
            36: begin
                if (byte_en[3])
                    mem[addr[13:5]*4+3] = data[35:27];
                if (byte_en[2])
                    mem[addr[13:5]*4+2] = data[26:18];
                if (byte_en[1])
                    mem[addr[13:5]*4+1] = data[17:9];
                if (byte_en[0])
                    mem[addr[13:5]*4]   = data[8:0];
            end
            default:     ;//null
        endcase
    end
    endtask

    task mem_write_b;
        input [13:0] addr;
        input [17:0] data;
        input [1:0]  byte_en;
    begin
        case (DATA_WIDTH_B)
            1: mem[addr[13:3]][addr[2:0]] = data[0];
            2: mem[addr[13:3]][addr[2:1]*2 +: 2] = data[1:0];
            4: mem[addr[13:3]][addr[2]*4 +: 4] = data[3:0];
            8: mem[addr[13:3]][7:0] = data[7:0];
            9: mem[addr[13:3]] = data[8:0];
            16: begin
                if (byte_en[1])
                    mem[addr[13:4]*2+1][7:0] = data[16:9];
                if (byte_en[0])
                    mem[addr[13:4]*2][7:0]   = data[7:0];
            end
            18: begin
                if (byte_en[1])
                    mem[addr[13:4]*2+1] = data[17:9];
                if (byte_en[0])
                    mem[addr[13:4]*2]   = data[8:0];
            end
            default:     ;//null
        endcase
    end
    endtask

    ///////////////
    // memory core
    ///////////////
reg CLKA_active;
reg CLKB_active;
initial begin
  CLKA_active = 1'b0;
  CLKB_active = 1'b0;
end
always @(posedge CLKA) begin
   if (CEA) begin
      CLKA_active <= 1'b1;
      #0.2 CLKA_active = 1'b0;
   end
   else
      CLKA_active <= 1'b0;
end
always @(posedge CLKB) begin
   if (CEB) begin
      CLKB_active <= 1'b1;
      #0.2 CLKB_active = 1'b0;
   end
   else
      CLKB_active <= 1'b0;
end

generate
////////////////////////////////////////////////////////////////////////////////////////////
// ROM or SINGLE_PORT 
////////////////////////////////////////////////////////////////////////////////////////////
if(RAM_MODE == "ROM" || RAM_MODE == "SINGLE_PORT") begin:ROMorSP_MODE

    always @(posedge CLKA) begin
        if (CEA)
            db_reg[17:0] <= DIB[17:0];
    end
    if (DATA_WIDTH_A > 18 || DATA_WIDTH_B > 18) begin

        assign write_en_a = (wea_reg == 1'b1);
        assign read_en_b  = (web_reg == 1'b0);
        // Port A operations
        always @(negedge CLKA_active)
        begin
            if (write_en_a) begin  // write
                mem_write_a(ada_reg[13:0], {db_reg[17:0], da_reg[17:0]}, bea_reg);
            end
        end
        // Port B operations
        always @(negedge CLKB_active or posedge rstb_int)
        begin
            if (rstb_int)
               {b_out,a_out} = {rstb_val_int,rsta_val_int};
            else if(read_en_b)
               {b_out[width_b-1:0], a_out[width_b-1:0]} = mem_read_b(adb_reg[13:0]);
        end

    end
    else  begin   //x1 x2 x4 x8 x9 x16 x18

        assign write_en_a = (wea_reg == 1'b1);
        assign read_en_a  = (wea_reg == 1'b0);
        // Port A operations
        always @(negedge CLKA_active)
        begin
            if (write_en_a)  begin  // write
               // read during write
               if (WRITE_MODE_A == "TRANSPARENT_WRITE") begin
                   a_out[width_a-1:0] = mem_read_a(ada_reg);

                   if(DATA_WIDTH_A == 16) begin
                       if(bea_reg[0])
                           a_out[7:0] = da_reg[7:0];
                       else
                           a_out[7:0] = a_out[7:0];

                       if(bea_reg[1])
                           a_out[15:8] = da_reg[16:9];
                       else
                           a_out[15:8] = a_out[15:8];
                   end
                   else if(DATA_WIDTH_A == 18) begin
                        if(bea_reg[0])
                            a_out[8:0] = da_reg[8:0];
                        else
                            a_out[8:0] = a_out[8:0];

                        if(bea_reg[1])
                            a_out[17:9] = da_reg[17:9];
                        else
                            a_out[17:9] = a_out[17:9];
                   end
                   else begin
                      a_out[width_a-1:0] = da_reg[width_a-1:0];
                   end
               end
               else if (WRITE_MODE_A == "READ_BEFORE_WRITE")
                   a_out[width_a-1:0] = mem_read_a(ada_reg[13:0]);

               mem_write_a(ada_reg[13:0], {18'b0, da_reg}, bea_reg);
            end
        end

        always @(negedge CLKA_active or posedge rsta_int)
        begin
            if (rsta_int)
               a_out = rsta_val_int;
            else if (read_en_a)          // read 
               a_out[width_a-1:0] = mem_read_a(ada_reg[13:0]);
        end
    end
end
////////////////////////////////////////////////////////////////////////////////////////////
//SIMPLE_DUAL_PORT
////////////////////////////////////////////////////////////////////////////////////////////
else if(RAM_MODE == "SIMPLE_DUAL_PORT")begin:SDP_MODE
    //port_A operation: only write in SDP MODE
    if (DATA_WIDTH_A > 18) begin:PORTA

        assign write_en_a = (wea_reg == 1'b1);

        always @(posedge CLKA) begin
           if (CEA)
              db_reg[17:0]  <= DIB[17:0];
        end
        always @(negedge CLKA_active) begin
           if (write_en_a)    // write 
              mem_write_a(ada_reg[13:0], {db_reg, da_reg},bea_reg);
        end
    end
    else  begin:PORTA    //  x1 x2 x4 x8 x9 x16 x18

        assign write_en_a = (wea_reg == 1'b1);
        assign read_en_a  = (wea_reg == 1'b0) ;

        always @(negedge CLKA_active) begin
           if (write_en_a)     // write
           begin
              if (WRITE_MODE_A == "TRANSPARENT_WRITE")
              begin
                 a_out[width_a-1:0] = mem_read_a(ada_reg);

                 if(DATA_WIDTH_A == 16) begin
                     if(bea_reg[0])
                         a_out[7:0] = da_reg[7:0];
                     else
                         a_out[7:0] = a_out[7:0];

                     if(bea_reg[1])
                         a_out[15:8] = da_reg[16:9];
                     else
                         a_out[15:8] = a_out[15:8];
                 end
                 else if(DATA_WIDTH_A == 18) begin
                      if(bea_reg[0])
                          a_out[8:0] = da_reg[8:0];
                      else
                          a_out[8:0] = a_out[8:0];

                      if(bea_reg[1])
                          a_out[17:9] = da_reg[17:9];
                      else
                          a_out[17:9] = a_out[17:9];
                 end
                 else begin
                    a_out[width_a-1:0] = da_reg[width_a-1:0];
                 end
              end
              else if (WRITE_MODE_A == "READ_BEFORE_WRITE")
                 a_out[width_a-1 : 0] = mem_read_a(ada_reg[13:0]);

              mem_write_a(ada_reg[13:0], {18'b0,da_reg}, bea_reg);
           end
        end
        if(DATA_WIDTH_B <= 16) begin
           always @(negedge CLKA_active or posedge rsta_int)
           begin
               if (rsta_int)
                  a_out = rsta_val_int;
               else if (read_en_a)
                  a_out[width_a-1 : 0] = mem_read_a(ada_reg[13:0]);
           end
        end
    end
    //port_B operation:only read in SDP MODE
    if (DATA_WIDTH_B > 18) begin:PORTB
    // SIMPLE_DUAL_PORT 
        assign read_en_b  = (web_reg == 1'b0);

        always @(negedge CLKB_active or posedge rstb_int)
        begin
           if (rstb_int)
              {b_out, a_out} = {rstb_val_int,rsta_val_int};
           else if (read_en_b)       // read 
              {b_out[width_b-1 : 0], a_out[width_b-1 : 0]} = mem_read_b(adb_reg[13:0]);
        end
    end
    else  begin:PORTB  //  x1 x2 x4 x8 x9 x16 x18

        assign read_en_b  = (web_reg == 1'b0);

        always @(negedge CLKB_active or posedge rstb_int)
        begin
           if (rstb_int)
              b_out = rstb_val_int;
           else if (read_en_b)   //  read 
              b_out[width_b-1 : 0] = mem_read_b(adb_reg[13:0]);
        end
    end
end
////////////////////////////////////////////////////////////////////////////////////////////
//DP_MODE
////////////////////////////////////////////////////////////////////////////////////////////
else   begin:DP_MODE   //  --x1 x2 x4 x8 x9 x16 x18
    assign write_en_a = (wea_reg == 1'b1) ;
    assign read_en_a  = (wea_reg == 1'b0) ;
    assign write_en_b = (web_reg == 1'b1) ;
    assign read_en_b  = (web_reg == 1'b0) ;
    // Port A operations
    always @(negedge CLKA_active)
    begin
        if (write_en_a)  begin  // write
            // read during write
            if (WRITE_MODE_A == "TRANSPARENT_WRITE")
            begin
               a_out[width_a-1:0] = mem_read_a(ada_reg);

               if(DATA_WIDTH_A == 16) begin
                   if(bea_reg[0])
                       a_out[7:0] = da_reg[7:0];
                   else
                       a_out[7:0] = a_out[7:0];

                   if(bea_reg[1])
                       a_out[15:8] = da_reg[16:9];
                   else
                       a_out[15:8] = a_out[15:8];
               end
               else if(DATA_WIDTH_A == 18) begin
                    if(bea_reg[0])
                        a_out[8:0] = da_reg[8:0];
                    else
                        a_out[8:0] = a_out[8:0];

                    if(bea_reg[1])
                        a_out[17:9] = da_reg[17:9];
                    else
                        a_out[17:9] = a_out[17:9];
               end
               else begin
                  a_out[width_a-1:0] = da_reg[width_a-1:0];
               end
            end
            else if (WRITE_MODE_A == "READ_BEFORE_WRITE")
               a_out[width_a-1 : 0] = mem_read_a(ada_reg[13:0]);

            mem_write_a(ada_reg[13:0], da_reg[17:0], bea_reg);
        end
    end

    always @(negedge CLKA_active or posedge rsta_int)
    begin
        if (rsta_int)
           a_out = rsta_val_int;
        else if (read_en_a)
           a_out[width_a-1 : 0] = mem_read_a(ada_reg[13:0]);
    end
    // Port B operations
    always @(posedge CLKB) begin
         if (CEB)
            db_reg[17:0] <= DIB[17:0];
    end

    always @(negedge CLKB_active)
    begin
        if (write_en_b)  begin  // write
            // read during write
            if (WRITE_MODE_B == "TRANSPARENT_WRITE")
            begin
                b_out[width_b-1:0] = mem_read_b(adb_reg);

                if(DATA_WIDTH_B == 16) begin
                    if(beb_reg[0])
                        b_out[7:0] = db_reg[7:0];
                    else
                        b_out[7:0] = b_out[7:0];

                    if(beb_reg[1])
                        b_out[15:8] = db_reg[16:9];
                    else
                        b_out[15:8] = b_out[15:8];
                end
                else if(DATA_WIDTH_B == 18) begin
                    if(beb_reg[0])
                        b_out[8:0] = db_reg[8:0];
                    else
                        b_out[8:0] = b_out[8:0];

                    if(beb_reg[1])
                        b_out[17:9] = db_reg[17:9];
                    else
                        b_out[17:9] = b_out[17:9];
                end
                else begin
                   b_out[width_b-1:0] = db_reg[width_b-1:0];
                end
            end
            else if (WRITE_MODE_B == "READ_BEFORE_WRITE")
                b_out[width_b-1 : 0] = mem_read_b(adb_reg[13:0]);

            mem_write_b(adb_reg[13:0], db_reg[17:0], beb_reg);
        end
    end

    always @(negedge CLKB_active or posedge rstb_int)
    begin
        if (rstb_int)
           b_out = rstb_val_int;
        else if (read_en_b)
           b_out[width_b-1 : 0] = mem_read_b(adb_reg[13:0]);
    end
end

endgenerate

//////////////
// core latch
//////////////
assign grsn = (GRS_EN == "TRUE") ? GRS_INST.GRSNET : 1'b1;
assign grs =  ~grsn;
or (rsta_grs, grs, RSTA);
or (rstb_grs, grs, RSTB);

reg rsta_grsn_d;

    always @(posedge CLKA_for_or) begin
        if (RSTA) begin
            rsta_grsn_d   <= 1'b1;
        end
        else begin
            rsta_grsn_d   <= 1'b0;
        end
    end

reg rstb_grsn_d;
    
    always @(posedge CLKB_for_or) begin
        if (RSTB) begin
            rstb_grsn_d   <= 1'b1;
        end
        else begin
            rstb_grsn_d   <= 1'b0;
        end
    end

initial begin
    rsta_grsn_d = 1'b1;
    rstb_grsn_d = 1'b1;
end

assign rsta_grs_sync  = (RST_TYPE == "SYNC") ? rsta_grsn_d : 1'b0;
assign rstb_grs_sync  = (RST_TYPE == "SYNC") ? rstb_grsn_d : 1'b0;
assign rsta_grs_async = (RST_TYPE == "ASYNC") ? rsta_grs : grs;
assign rstb_grs_async = (RST_TYPE == "ASYNC") ? rstb_grs : grs;

assign rsta_int = rsta_grs_sync | rsta_grs_async;
assign rstb_int = rstb_grs_sync | rstb_grs_async;
/////////////////////////////////////////////////////////////////////
//port out
assign CLKA_for_or = (DOA_REG_CLKINV == 1) ? ~CLKA : CLKA;
assign CLKB_for_or = (DOB_REG_CLKINV == 1) ? ~CLKB : CLKB;

generate
if (DATA_WIDTH_B >= 32)
begin:FAKE_DP_OUT
    //port_A output
    always @(posedge CLKB_for_or or posedge rstb_int)
    begin
        if (rstb_int)
            doa_reg <= RSTA_VAL;
        else if (ORCEB)
            doa_reg <= doa;
    end

    //doa combination logic
    always @(a_out)
    begin
        case(DATA_WIDTH_B)
            32: {doa[16:9],doa[7:0]} = a_out[width_b-1:0];
            36:  doa[width_b-1:0] = a_out[width_b-1:0];
        endcase
    end

    always @(doa or doa_reg)
    begin
        if (DOB_REG == 0)
            doa_mux = doa;
        else
            doa_mux = doa_reg;
    end

    //port_B output
    always @(posedge CLKB_for_or or posedge rstb_int)
    begin
        if (rstb_int)
            dob_reg <= RSTB_VAL;
        else if (ORCEB)
            dob_reg <= dob;
    end

    //dob combination logic
    always @(b_out)
    begin
        case(DATA_WIDTH_B)
            32:{dob[16:9],dob[7:0]} = b_out[width_b-1 : 0];
            36: dob[width_b-1:0] = b_out[width_b-1 : 0];
        endcase
    end

    always @(dob or dob_reg)
    begin
        if (DOB_REG == 0)
            dob_mux = dob;
        else
            dob_mux = dob_reg;
    end
end
else
begin:TRUE_DP_OUT
    //port_A output

    always @(posedge CLKA_for_or or posedge rsta_int)
    begin
        if (rsta_int)
            doa_reg <= RSTA_VAL;
        else if (ORCEA)
            doa_reg <= doa;
    end

    //doa combination logic
    always @(a_out)
    begin
        case(DATA_WIDTH_A)  
           1: {doa[16:9],doa[7:0]} = {16{a_out[width_a-1:0]}};
           2: {doa[16:9],doa[7:0]} = { 8{a_out[width_a-1:0]}};
           4: {doa[16:9],doa[7:0]} = { 4{a_out[width_a-1:0]}};
           8: {doa[16:9],doa[7:0]} = { 2{a_out[width_a-1:0]}};
           9: {doa[17:9],doa[8:0]} = { 2{a_out[width_a-1:0]}};
           16:{doa[16:9],doa[7:0]} =     a_out[width_a-1:0]  ;
           18: doa[17:0]           =     a_out[width_a-1:0]  ; 
        endcase
    end

    always @(doa or doa_reg)
    begin
        if (DOA_REG == 0)
            doa_mux = doa;
        else
            doa_mux = doa_reg;
    end
    //port_B output

    always @(posedge CLKB_for_or or posedge rstb_int)
    begin
        if (rstb_int)
            dob_reg <= RSTB_VAL;
        else if (ORCEB)
            dob_reg <= dob;
    end

    //dob combination logic
    always @(b_out)
    begin
        case(DATA_WIDTH_B) 
           1: {dob[16:9],dob[7:0]} = {16{b_out[width_b-1:0]}};
           2: {dob[16:9],dob[7:0]} = { 8{b_out[width_b-1:0]}};
           4: {dob[16:9],dob[7:0]} = { 4{b_out[width_b-1:0]}};
           8: {dob[16:9],dob[7:0]} = { 2{b_out[width_b-1:0]}};
           9: {dob[17:9],dob[8:0]} = { 2{b_out[width_b-1:0]}};
           16:{dob[16:9],dob[7:0]} =     b_out[width_b-1:0]  ;
           18: dob[17:0]           =     b_out[width_b-1:0] ; 
        endcase
    end

    always @(dob or dob_reg)
    begin
        if (DOB_REG == 0)
            dob_mux = dob;
        else
            dob_mux = dob_reg;
    end
end
endgenerate

assign DOA = doa_mux;
assign DOB = dob_mux;

// synthesis translate_on
endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_MULTACC9.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

//P = MAC + A*B
module GTP_MULTACC9 #(
    parameter GRS_EN             = "TRUE", //"TRUE"; "FALSE"
    parameter SYNC_RST           = "FALSE", //"TRUE"; "FALSE"
    parameter INREG_EN           = "FALSE",  //"TRUE"; "FALSE"
    parameter PIPEREG_EN         = "FALSE",   //"TRUE"; "FALSE"
    parameter ACC_ADDSUB_OP      = 0,
    parameter DYN_ACC_ADDSUB_OP  = 1,     //Select parameter ADDSUB or input ADDSUB
    parameter OVERFLOW_MASK      = 32'h0, //PSIZE = 32 OVERflow setting =  'h1_0000_00XX , bit width = PSIZE
    parameter PATTERN            = 32'h0, //compare pattern
    parameter MASKPAT            = 32'h0, //pattern mask
    parameter DYN_ACC_INIT       = 0,     //acc init value dynamic input
    parameter ACC_INIT_VALUE     = 32'h0  //acc init value parameter 
) (
    output  [31:0] P,
    output  OVER,
    output  UNDER,
    output  EQZ,
    output  EQZM,
    output  EQOM,
    output  EQPAT,
    output  EQPATN,

    input   CE,
    input   RST,
    input   CLK,
    input   [8:0] A,
    input   [8:0] B,
    input   A_SIGNED,
    input   B_SIGNED,
    input   [31:0] ACC_INIT,
    input   ACC_ADDSUB,
    input   RELOAD
);

    wire [31:0] R;

    INT_PREADD_MULTACC #(
        . GRS_EN(GRS_EN),     
        . SYNC_RST(SYNC_RST),   
        . INREG_EN(INREG_EN),   
        . PIPEREG_EN(PIPEREG_EN), 
        . ACCUMADDSUB_OP(ACC_ADDSUB_OP), 
        . DYN_OP_SEL(DYN_ACC_ADDSUB_OP),     
        . ASIZE(9),    
        . BSIZE(9),    
        . PSIZE(32),    
        . PREADD_EN(0),
        . MASK(OVERFLOW_MASK),      
        . DYN_ACC_INIT(DYN_ACC_INIT),     
        . ACC_INIT_VALUE(ACC_INIT_VALUE)
    ) U_MACC (
        .CE(CE),
        .RST(RST),
        .CLK(CLK),
        .A(A),
        .B(B),
        .A_SIGNED(A_SIGNED),
        .B_SIGNED(B_SIGNED),
        .C_SIGNED(B_SIGNED),
        .C(9'b0),
        .PREADDSUB(1'b0),
        .ACCUM_INIT(ACC_INIT),
        .ACCUMADDSUB(ACC_ADDSUB),
        .RELOAD(RELOAD),
        .P(P),
        .OVER(OVER),
        .UNDER(UNDER),
        .R(R)     
    );

    INT_FLAG #(
        . GRS_EN(GRS_EN),
        . SYNC_RST(SYNC_RST),
        . PSIZE(32),
        . PATSIZE(32),
        . MASKPATSIZE(32),
        . OUTREG_EN("TRUE")
    ) U_FLAG (
        . CE(CE),
        . RST(RST),
        . CLK(CLK),
        . P(P),
        . PATTERN(PATTERN),
        . MASKPAT(MASKPAT),
        . OVERFLOW_MASK(OVERFLOW_MASK),
        . R(R),
        . eqz(EQZ),
        . eqzm(EQZM),
        . eqom(EQOM),
        . eqpat(EQPAT),
        . eqpatn(EQPATN)
    );

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_DFF_PE.v
//
// Functional description: D-type flip-flop with async set and enable
//
// Parameter description:
//      INIT: init value
//
// Port description:
//      P: asynchronous set
//      CE  : enable
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_DFF_PE
#(
    parameter GRS_EN = "TRUE",
    parameter INIT = 1'b1
) (
    output reg Q,
    input wire D,
    input wire CLK, P, CE
);

    wire grs_n;
    wire grs, RS;

    tri1 grsnet = GRS_INST.GRSNET;
    assign grs_n=(GRS_EN=="TRUE")?grsnet:1'b1;

    not (grs, grs_n);
    or (RS, grs, P);

    initial Q = 1'bx;

    always @(posedge CLK or posedge RS) begin
        if (RS)
            Q <= 1'b1;
        else if (CE)
            Q <= D;
    end

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: Internal simulation model
// Filename: GTP_INBUF.v
//
// Functional description: Input Buffer
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_INBUF #(
    parameter IOSTANDARD = "DEFAULT",
    parameter TERM_DDR = "ON"
)(
    output O,
    input I
) /* synthesis syn_black_box */ ;
  
  initial begin
    case (IOSTANDARD)
    "LVTTL33", "PCI33", "LVCMOS33", "LVCMOS25", "LVCMOS18", "LVCMOS15", "LVCMOS12", "SSTL25_I", "SSTL25_II", "SSTL18_I", "SSTL18_II", "SSTL15_I", "SSTL15_II", "HSTL18_I", "HSTL18_II", "HSTL15_I", "SSTL15_I_CAL", "SSTL15_II_CAL", "HSTL15_I_CAL", "DEFAULT" :;
    default : begin
           $display("Attribute Syntax Error : The attribute IOSTANDARD on GTP_INBUF instance %m is set to %s.", IOSTANDARD);
           $finish;
              end
    endcase

    case (TERM_DDR)
    "ON", "OFF" :;
    default : begin
           $display("Attribute Syntax Error : The attribute TERM_DDR on GTP_INBUF instance %m is set to %s.", TERM_DDR);
           $finish;
              end
    endcase
    end

    buf (O, I);

endmodule





//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_PLL.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1ns/10fs
module GTP_PLL #(
    parameter CLKIN_FREQ = "50MHZ",
    parameter DYNAMIC_CLKIN_EN  = "FALSE", //"TRUE"; "FALSE"
    parameter CLKIN_SSEL        = 1'b0,    //0~1
    parameter DYNAMIC_RATIOI_EN = "FALSE", //"TRUE"; "FALSE"
    parameter integer STATIC_RATIOI = 1,   //1~64
    parameter DYNAMIC_RATIOF_EN = "FALSE", //"TRUE"; "FALSE"
    parameter integer STATIC_RATIOF = 1,   //1~64
    parameter DYNAMIC_RATIO_EN  = "FALSE", //"TRUE"; "FALSE"
    parameter integer STATIC_RATIO  = 2,   //2,4,~128
    parameter integer CLKOUT2_SEL   = 2,   //0~3
    parameter DYNAMIC_RATIO2_EN = "FALSE", //"TRUE"; "FALSE"
    parameter integer STATIC_RATIO2 = 2,   //2,4,6,8~128
    parameter integer CLKOUT3_SEL   = 2,   //0~3
    parameter DYNAMIC_RATIO3_EN = "FALSE", //"TRUE"; "FALSE"
    parameter integer STATIC_RATIO3 = 2,   //2,4,6,8~128
    parameter integer CLKOUT4_SEL   = 2,   //0~3
    parameter DYNAMIC_RATIO4_EN = "FALSE", //"TRUE"; "FALSE"
    parameter integer STATIC_RATIO4 = 2,   //2,4,6,8~128
    parameter INTERNAL_FB = "CLKOUT0",     //"CLKOUT0"; "CLKOUT1"; "CLKOUT2"; "DISABLE"
    parameter EXTERNAL_FB = "DISABLE",     //"CLKOUT0"; "CLKOUT1"; "CLKOUT2"; "CLKOUT3"; "CLKOUT4"; "DISABLE"
    parameter BANDWIDTH   = "OPTIMIZED",   //"LOW"; "OPTIMIZED"; "HIGH"
    parameter DYNAMIC_DUPS1_EN  = "FALSE", //"TRUE"; "FALSE"
    parameter integer STATIC_DUTY1  = 8,
    parameter integer STATIC_PHASE1 = 0,
    parameter DYNAMIC_DUPS2_EN  = "FALSE", //"TRUE"; "FALSE"
    parameter integer STATIC_DUTY2  = 8,
    parameter integer STATIC_PHASE2 = 0,
    parameter DYNAMIC_DUPS3_EN  = "FALSE", //"TRUE"; "FALSE"
    parameter integer STATIC_DUTY3  = 8,
    parameter integer STATIC_PHASE3 = 0,
    parameter DYNAMIC_DUPS4_EN  = "FALSE", //"TRUE"; "FALSE"
    parameter integer STATIC_DUTY4  = 8,
    parameter integer STATIC_PHASE4 = 0,
    parameter CLKOUT0_SYN_EN = "TRUE",  //"TRUE"; "FALSE"
    parameter CLKOUT1_SYN_EN = "FALSE", //"TRUE"; "FALSE"
    parameter CLKOUT2_SYN_EN = "FALSE", //"TRUE"; "FALSE"
    parameter CLKOUT3_SYN_EN = "FALSE", //"TRUE"; "FALSE"
    parameter CLKOUT4_SYN_EN = "FALSE", //"TRUE"; "FALSE"
    parameter RST_INNER_EN   = "TRUE",  //"TRUE"; "FALSE"
    parameter RSTIDIV_EN     = "TRUE",  //"TRUE"; "FALSE"
    parameter RSTODIV_EN     = "TRUE",  //"TRUE"; "FALSE"
    parameter integer CLKOUT3_DIV125_M = 1,
    parameter integer CLKOUT3_DIV125_N = 1,
    parameter CLKOUT4_DIV32BIT_K = 1000
    )(
    output CLKOUT0,
    output CLKOUT1,
    output CLKOUT2,
    output CLKOUT3,
    output CLKOUT4,
    output LOCK,
    input CLKIN1,
    input CLKIN2,
    input CLKIN_DSEL,
    input CLKFB,
    input CLKOUT0_SYN,
    input CLKOUT1_SYN,
    input CLKOUT2_SYN,
    input CLKOUT3_SYN,
    input CLKOUT4_SYN,
    input [5:0] RATIOI,
    input [5:0] RATIOF,
    input [5:0] RATIO,
    input [5:0] RATIO2,
    input [5:0] RATIO3,
    input [5:0] RATIO4,
    input [3:0] DUTY1,
    input [3:0] DUTY2,
    input [3:0] DUTY3,
    input [3:0] DUTY4,
    input [3:0] PHASE1,
    input [3:0] PHASE2,
    input [3:0] PHASE3,
    input [3:0] PHASE4,
    input PLL_PWD,
    input RST,
    input RSTIDIV,
    input RSTODIV
    )/* synthesis syn_black_box */;

    wire rst_inner_en_set;
    wire rstidiv_en_set;
    wire rstodiv_en_set;
    reg  inner_rst;
    wire pll_rstn;
    wire idiv_rstn;
    wire odiv_rstn;
    wire clkin_set;

    reg clk_in_first_time;
    reg clk_fb_first_time;
    realtime clk_in_first_edge;
    realtime clk_fb_first_edge;

    real clkin_cj;

    reg adjust;
    realtime fb_route_delay;
    realtime virtual_delay1;
    integer tmp_ratio;
    realtime tmp_delay;
    realtime real_delay;

    wire [6:0] ratioi_set_int;
    wire [6:0] ratiof_set_int;
    wire [7:0] ratio_set_int;
    wire [7:0] ratio2_set_int;
    wire [7:0] ratio3_set_int;
    wire [7:0] ratio4_set_int;
    wire [7:0] total_ratio_int;

    reg clkin_reg;
    realtime clkin_rtime_last;
    realtime clkin_rtime_next;
    realtime clkin_time;
    realtime clkin_time_d1;
    realtime clkin_time_d2;
    realtime clkin_time_d3;
    reg clkout_lock;
    realtime clkout_time;
    realtime clkout_time_half;
    integer clkout_time_amp;
    realtime clkout_time_real;
    realtime clkout_time_dev;
    wire clk_valid;
    real cnt_fdiv;
    reg clk_gate;
    reg inner_clk;

    reg vcoclk;

    wire clk_lock;
    reg [2:0] cnt_clkfb;
    reg start_clk;
    reg [10:0] cnt_lock;
    reg lock_reg;

    wire [3:0] phase1_sel;
    wire [3:0] phase2_sel;
    wire [3:0] phase3_sel;
    wire [3:0] phase4_sel;
    wire [3:0] duty1_sel;
    wire [3:0] duty2_sel;
    wire [3:0] duty3_sel;
    wire [3:0] duty4_sel;
    realtime phase_adjut_1_time;
    realtime phase_adjut_2_time;
    realtime phase_adjut_3_time;
    realtime phase_adjut_4_time;
    reg inv1;
    reg inv2;
    reg inv3;
    reg inv4;
    reg clkout_reg;
    reg clkout_1_reg;
    reg clkout_2_reg;
    reg clkout_3_reg;
    reg clkout_4_reg;
    wire clkout_0_reg_n;
    wire clkout_1_reg_n;
    wire clkout_2_reg_n;
    wire clkout_3_reg_n;
    wire clkout_4_reg_n;
    integer count_o2;
    integer count_o3;
    integer count_o4;
    reg clkout_div_reg1;
    reg clkout_div_reg2;
    reg clkout_div_reg3;
    reg clkout_div_reg4;
    realtime clk_vco_time;
    realtime div125_time_div2;
    realtime div32bit_time;
    reg div125_valid;
    reg div125;
    reg div125_reg;
    wire div32bit_reg;

    initial
    begin
        if((DYNAMIC_CLKIN_EN == "TRUE") || (DYNAMIC_CLKIN_EN == "FALSE"))
        begin
        end
        else
            $display (" GTP_PLL error: illegal setting for DYNAMIC_CLKIN_EN");

        if((DYNAMIC_RATIOI_EN == "TRUE") || (DYNAMIC_RATIOI_EN == "FALSE"))
        begin
        end
        else
            $display (" GTP_PLL error: illegal setting for DYNAMIC_RATIOI_EN");

        if((DYNAMIC_RATIOF_EN == "TRUE") || (DYNAMIC_RATIOF_EN == "FALSE"))
        begin
        end
        else
            $display (" GTP_PLL error: illegal setting for DYNAMIC_RATIOF_EN");

        if((DYNAMIC_RATIO_EN == "TRUE") || (DYNAMIC_RATIO_EN == "FALSE"))
        begin
        end
        else
            $display (" GTP_PLL error: illegal setting for DYNAMIC_RATIO_EN");

        if((CLKOUT2_SEL == 0) || (CLKOUT2_SEL == 1) || (CLKOUT2_SEL == 2 ))
        begin
        end
        else
            begin
                $display (" GTP_PLL error: illegal setting for CLKOUT2_SEL");
                $stop;
            end

        if((DYNAMIC_RATIO2_EN == "TRUE") || (DYNAMIC_RATIO2_EN == "FALSE"))
        begin
        end
        else
            $display (" GTP_PLL error: illegal setting for DYNAMIC_RATIO2_EN");

        if((DYNAMIC_RATIO3_EN == "TRUE") || (DYNAMIC_RATIO3_EN == "FALSE"))
        begin
        end
        else
            $display (" GTP_PLL error: illegal setting for DYNAMIC_RATIO3_EN");

        if((DYNAMIC_RATIO4_EN == "TRUE") || (DYNAMIC_RATIO4_EN == "FALSE"))
        begin
        end
        else
            $display (" GTP_PLL error: illegal setting for DYNAMIC_RATIO4_EN");

        if((INTERNAL_FB == "CLKOUT0") || (INTERNAL_FB == "CLKOUT1") || (INTERNAL_FB == "CLKOUT2") || (INTERNAL_FB == "DISABLE"))
        begin
        end
        else
            $display (" GTP_PLL error: illegal setting for INTERNAL_FB");

        if((EXTERNAL_FB == "CLKOUT0") || (EXTERNAL_FB == "CLKOUT1") || (EXTERNAL_FB == "CLKOUT2") || (EXTERNAL_FB == "CLKOUT3") || (EXTERNAL_FB == "CLKOUT4") || (EXTERNAL_FB == "DISABLE"))
        begin
        end
        else
            $display (" GTP_PLL error: illegal setting for EXTERNAL_FB");

        if((BANDWIDTH == "OPTIMIZED") || (BANDWIDTH == "LOW") || (BANDWIDTH == "HIGH"))
        begin
        end
        else
            $display (" GTP_PLL error: illegal setting for BANDWIDTH");

        if((DYNAMIC_DUPS1_EN == "TRUE") || (DYNAMIC_DUPS1_EN == "FALSE"))
        begin
        end
        else
            $display (" GTP_PLL error: illegal setting for DYNAMIC_DUPS1_EN");

        if((DYNAMIC_DUPS2_EN == "TRUE") || (DYNAMIC_DUPS2_EN == "FALSE"))
        begin
        end
        else
            $display (" GTP_PLL error: illegal setting for DYNAMIC_DUPS2_EN");

        if ((DYNAMIC_DUPS3_EN == "TRUE") || (DYNAMIC_DUPS3_EN == "FALSE"))
        begin
        end
        else
            $display (" GTP_PLL error: illegal setting for DYNAMIC_DUPS3_EN");

        if((DYNAMIC_DUPS4_EN == "TRUE") || (DYNAMIC_DUPS4_EN == "FALSE"))
        begin
        end
        else
            $display (" GTP_PLL error: illegal setting for DYNAMIC_DUPS4_EN");

        if((CLKOUT0_SYN_EN == "TRUE") || (CLKOUT0_SYN_EN == "FALSE"))
        begin
        end
        else
            $display (" GTP_PLL error: illegal setting for CLKOUT0_SYN_EN");

        if((CLKOUT1_SYN_EN == "TRUE") || (CLKOUT1_SYN_EN == "FALSE"))
        begin
        end
        else
            $display (" GTP_PLL error: illegal setting for CLKOUT1_SYN_EN");

        if((CLKOUT2_SYN_EN == "TRUE") || (CLKOUT2_SYN_EN == "FALSE"))
        begin
        end
        else
            $display (" GTP_PLL error: illegal setting for CLKOUT2_SYN_EN");

        if ((CLKOUT3_SYN_EN == "TRUE") || (CLKOUT3_SYN_EN == "FALSE"))
        begin
        end
        else
            $display (" GTP_PLL error: illegal setting for CLKOUT3_SYN_EN");

        if((CLKOUT4_SYN_EN == "TRUE") || (CLKOUT4_SYN_EN == "FALSE"))
        begin
        end
        else
        $display (" GTP_PLL error: illegal setting for CLKOUT4_SYN_EN");

        if((RST_INNER_EN == "TRUE") || (RST_INNER_EN == "FALSE"))
        begin
        end
        else
            $display (" GTP_PLL error: illegal setting for RST_INNER_EN");

        if((RSTIDIV_EN == "TRUE") || (RSTIDIV_EN == "FALSE"))
        begin
        end
        else
            $display (" GTP_PLL error: illegal setting for RSTIDIV_EN");

        if((RSTODIV_EN == "TRUE") || (RSTODIV_EN == "FALSE"))
        begin
        end
        else
            $display (" GTP_PLL error: illegal setting for RSTODIV_EN");
    end

    initial
    begin
        inner_rst      = 1;
        clkin_reg      = 0;
        clk_in_first_time = 1'b0;
        clk_fb_first_time = 1'b0;
        clk_in_first_edge = 0.0;
        clk_fb_first_edge = 0.0;
        fb_route_delay = 0.0;
        tmp_ratio = 0;
        tmp_delay = 0.0;
        real_delay = 0.0;
        clkin_rtime_last = 0;
        clkin_rtime_next = 0;
        clkin_time       = 0;
        clkin_time_d1    = 0;
        clkin_time_d2    = 0;
        clkin_time_d3    = 0;
        clkout_lock      = 0;
        clkout_time      = 0;
        clkout_time_half = 0;
        clkout_time_amp  = 0;
        clkout_time_real = 0;
        clkout_time_dev  = 0;
        cnt_fdiv   = 0;
        clk_gate   = 1;
        inner_clk  = 1'b0;
        vcoclk    = 1'b0;
        phase_adjut_1_time = 0;
        phase_adjut_2_time = 0;
        phase_adjut_3_time = 0;
        phase_adjut_4_time = 0;
        inv1 = 0;
        inv2 = 0;
        inv3 = 0;
        inv4 = 0;
        clkout_reg   = 0;
        clkout_1_reg = 0;
        clkout_2_reg = 0;
        clkout_3_reg = 0;
        clkout_4_reg = 0;
        count_o2 = 0;
        count_o3 = 0;
        count_o4 = 0;
        clkout_div_reg1 = 0;
        clkout_div_reg2 = 0;
        clkout_div_reg3 = 0;
        clkout_div_reg4 = 0;
        clk_vco_time     = 1;
        div125_time_div2 = 1;
        div125_valid     = 0;
        div125     = 0;
        div125_reg = 0;
        #1.01;
        inner_rst  = 0;
        clk_in_first_time = 1'b1;
        clk_fb_first_time = 1'b1;
    end

    assign rst_inner_en_set = (RST_INNER_EN == "TRUE") ? 1'b1 : 1'b0;
    assign rstodiv_en_set   = (RSTODIV_EN == "TRUE") ? 1'b1 : 1'b0;
    assign rstidiv_en_set   = (RSTIDIV_EN == "TRUE") ? 1'b1 : 1'b0; 
    assign pll_rstn  = ~ (PLL_PWD | RST | (RSTODIV && rstodiv_en_set) | (RSTIDIV && rstidiv_en_set) | (inner_rst && rst_inner_en_set));
    assign idiv_rstn = ~ ((RSTIDIV && rstidiv_en_set) | (inner_rst && rst_inner_en_set) | RST | PLL_PWD);
    assign odiv_rstn = ~ ((RSTODIV && rstodiv_en_set) | (inner_rst && rst_inner_en_set) | RST | PLL_PWD);
    assign clkin_set = (DYNAMIC_CLKIN_EN == "TRUE") ? CLKIN_DSEL : CLKIN_SSEL;

    assign ratioi_set_int  = (DYNAMIC_RATIOI_EN == "TRUE") ? 64-RATIOI : STATIC_RATIOI;
    assign ratiof_set_int  = (DYNAMIC_RATIOF_EN == "TRUE") ? 64-RATIOF : STATIC_RATIOF;
    assign ratio_set_int   = (DYNAMIC_RATIO_EN  == "TRUE") ? 2*(63-RATIO)+2  : STATIC_RATIO;
    assign ratio2_set_int  = (DYNAMIC_RATIO2_EN == "TRUE") ? 2*(63-RATIO2)+2 : STATIC_RATIO2;
    assign ratio3_set_int  = (DYNAMIC_RATIO3_EN == "TRUE") ? 2*(63-RATIO3)+2 : STATIC_RATIO3;
    assign ratio4_set_int  = (DYNAMIC_RATIO4_EN == "TRUE") ? 2*(63-RATIO4)+2 : STATIC_RATIO4;
    assign total_ratio_int = (INTERNAL_FB == "CLKOUT0" || EXTERNAL_FB == "CLKOUT0") ? 1 :
                             (INTERNAL_FB == "CLKOUT1" || EXTERNAL_FB == "CLKOUT1") ? 1 :
                             ((INTERNAL_FB == "CLKOUT2" || EXTERNAL_FB == "CLKOUT2") && (CLKOUT2_SEL == 1)) ? ratio2_set_int :
                             ((INTERNAL_FB == "CLKOUT2" || EXTERNAL_FB == "CLKOUT2") && (CLKOUT2_SEL == 2)) ? 1 :
                             (EXTERNAL_FB == "CLKOUT3" && CLKOUT3_SEL == 1) ? ratio3_set_int :
                             (EXTERNAL_FB == "CLKOUT3" && CLKOUT3_SEL == 2) ? 1 :
                             (EXTERNAL_FB == "CLKOUT4" && CLKOUT4_SEL == 1) ? ratio4_set_int :
                             (EXTERNAL_FB == "CLKOUT4" && CLKOUT4_SEL == 2) ? 1 : 1;

    always @(clkin_set or CLKIN1 or CLKIN2)
    begin
        case(clkin_set)
            0: clkin_reg = CLKIN1;
            1: clkin_reg = CLKIN2;
        endcase
    end

////FBCK_DELAY/////////////////////////////////////////
    always @(posedge clkin_reg or negedge pll_rstn)
    begin
        if(!pll_rstn)
        begin
            clk_in_first_time = 1'b1;
            clk_in_first_edge = 0.0;
        end
        else
        begin
            if(clk_in_first_time == 1'b1)
                clk_in_first_edge = $realtime;
            clk_in_first_time = 1'b0;
        end
    end

    always @(posedge CLKFB or negedge pll_rstn)
    begin
        if(!pll_rstn)
        begin
            clk_fb_first_time = 1'b1;
            clk_fb_first_edge = 0.0;
        end
        else
        begin
            if(clk_fb_first_time == 1'b1)
                clk_fb_first_edge = $realtime;
            clk_fb_first_time = 1'b0;
        end
    end
///////////////////////////////////////////////////////
    always @(*)
    begin
        if(BANDWIDTH == "LOW" || BANDWIDTH == "OPTIMIZED")
            if(CLKIN_FREQ/ratioi_set_int <= 100)
                clkin_cj = 0.45/ratioi_set_int;
            else
                clkin_cj = 0.45/CLKIN_FREQ;
        else if(BANDWIDTH == "HIGH")
            if(CLKIN_FREQ/ratioi_set_int <= 100)
                clkin_cj = 0.25/ratioi_set_int;
            else
                clkin_cj = 0.25/CLKIN_FREQ;
    end
///////////////////////////////////////////////////////
    always @(posedge clkin_reg or negedge pll_rstn)
    begin
        if(!pll_rstn)
        begin
            clkin_rtime_last = 0;
            clkin_rtime_next = 0;
            clkin_time    <= 0;
            clkin_time_d1 <= 0;
            clkin_time_d2 <= 0;
            clkin_time_d3 <= 0;
            clkout_lock   <= 0;
            clkout_time   <= 0;
            clkout_time_half <= 0;
            clkout_time_amp   = 0;
            clkout_time_real  = 0;
            clkout_time_dev   = 0;
        end
        else
        begin
            clkin_rtime_last = clkin_rtime_next;
            clkin_rtime_next = $realtime;
            if(clkin_rtime_last > 0)
            begin
                clkin_time    <= clkin_rtime_next - clkin_rtime_last;
                clkin_time_d1 <= clkin_time;
                clkin_time_d2 <= clkin_time_d1;
                clkin_time_d3 <= clkin_time_d2;
            end
            if(clkin_time > 0) begin
                clkout_lock <= (clkin_time > 0) &&
                               (clkin_time_d1 > 0) &&
                               (clkin_time_d2 > 0) &&
                               (clkin_time_d3 > 0) &&
                               ((clkin_time - clkin_time_d1) < clkin_cj) && 
                               ((clkin_time_d1 - clkin_time) < clkin_cj) && 
                               ((clkin_time_d1 - clkin_time_d2) < clkin_cj) && 
                               ((clkin_time_d2 - clkin_time_d1) < clkin_cj) && 
                               ((clkin_time_d2 - clkin_time_d3) < clkin_cj) && 
                               ((clkin_time_d3 - clkin_time_d2) < clkin_cj);
            end
            if(clkin_time > 0)
            begin
                clkout_time       = (clkin_time * ratioi_set_int/ratiof_set_int)/total_ratio_int;
                clkout_time_half  = clkout_time / 2;
                clkout_time_amp   = clkout_time_half * 100000;
                clkout_time_real  = clkout_time_amp / 1;
                clkout_time_dev   = (clkin_time - (clkout_time_real * 2 * ratiof_set_int * total_ratio_int) / (100000 * ratioi_set_int))/2;
            end
        end
    end

    assign #(clkout_time/2) clk_valid = clkout_lock;

    reg done;
    integer idiv_set;
    integer fdiv_set;
    integer swap_set;
    integer fdiv_int;
    realtime offset;

    initial begin
        done = 1'b0;
        idiv_set = 0;
        fdiv_set = 0;
        swap_set = 0;
        fdiv_int = 0;
        offset = 0;
    end

    always @(*)
    begin
        done = 1'b0;
        idiv_set = ratioi_set_int;
        fdiv_set = ratiof_set_int;
        while(!done)
        begin
            if(idiv_set < fdiv_set)
            begin
                swap_set = idiv_set;
                idiv_set = fdiv_set;
                fdiv_set = swap_set;
            end
            else
                if(fdiv_set != 0)
                    idiv_set = idiv_set - fdiv_set;
                else
                    done = 1;
        end
        fdiv_int = idiv_set;
        offset = clkout_time_dev * ratioi_set_int/fdiv_int;
    end

    //vco frequencyOA
    always @(inner_clk or clkout_lock)
    begin
        if(clkout_lock == 1'b0)
        begin
            inner_clk <= 1'b0;
            clk_gate <= 1'b1;
            cnt_fdiv = 0;
        end
        else
        begin
            if(clk_gate == 1'b1)
            begin
                inner_clk <= 1'b1;
                clk_gate <= 1'b0;
                cnt_fdiv = 0;
            end
            else
            begin
                cnt_fdiv = cnt_fdiv + 1;
                if(cnt_fdiv == ratiof_set_int/fdiv_int)
                begin
                    inner_clk <= #(clkout_time_half+offset) ~inner_clk;
                    cnt_fdiv = 0;
                end
                else
                    inner_clk <= #clkout_time_half ~inner_clk;
            end
        end
    end

    always @(clkin_reg or CLKFB or negedge pll_rstn)
    begin
        if(!pll_rstn)
        begin
            adjust <= 1'b1;
            fb_route_delay = 0.0;
            tmp_ratio  = 0;
            tmp_delay  = 0.0;
            real_delay = 0.0;
        end
        else
            if(adjust == 1'b1)
            begin
                fb_route_delay = clk_fb_first_edge - clk_in_first_edge;
                if((clkin_time > 0) && (fb_route_delay > 0))
                begin
                    tmp_ratio  = fb_route_delay / clkin_time;
                    tmp_delay  = fb_route_delay - (clkin_time * tmp_ratio);
                    real_delay = clkin_time - tmp_delay;
                    adjust <= 1'b0;
                end
            end
    end

    always @(inner_clk)
    begin
        if(EXTERNAL_FB == "CLKOUT0" || EXTERNAL_FB == "CLKOUT1" || EXTERNAL_FB == "CLKOUT2" || EXTERNAL_FB == "CLKOUT3" || EXTERNAL_FB == "CLKOUT4")
            vcoclk <= #real_delay inner_clk;
        else
            vcoclk <= inner_clk;
    end
//************************************************************************
    assign clk_lock = (INTERNAL_FB == "DISABLE") ? CLKFB : clkin_reg;
    
    always @(posedge clk_lock or negedge pll_rstn)
    begin
        if(!pll_rstn)
        begin
            start_clk <= 1'b0;
            cnt_clkfb <= 2'b00;
        end
        else
            if(cnt_clkfb == 3)
                start_clk = 1'b1;
            else
                cnt_clkfb = cnt_clkfb + 1;
    end

    always @(posedge clkin_reg or negedge pll_rstn)
    begin
        if(!pll_rstn)
        begin
            cnt_lock <= 11'b000_0000_0001;
            lock_reg <= 1'b0;
        end
        else
            if(clkout_lock && start_clk)
                if(cnt_lock == ratioi_set_int*3)
                    lock_reg <= 1'b1;
                else
                    cnt_lock <= cnt_lock+1;
            else
            begin
                cnt_lock <= 11'b000_0000_0001;
                lock_reg <= 1'b0;
            end
    end

    assign LOCK = lock_reg;
//************************************************************************
    //for clkout0
    always @(*)
    begin 
        if(!pll_rstn)
            clkout_reg <= 1'b0;
        else
            clkout_reg <= vcoclk;
    end

    assign clkout_0_reg_n = ~clkout_reg;

    reg CLKOUT0_SYN_n_d1;
    reg CLKOUT0_SYN_n_d2;
    reg CLKOUT0_SYN_n_d3;
    initial
    begin
        CLKOUT0_SYN_n_d1 = 1'b0;
        CLKOUT0_SYN_n_d2 = 1'b0;
        CLKOUT0_SYN_n_d3 = 1'b0;
    end

    always @(negedge clkout_0_reg_n)
    begin
        CLKOUT0_SYN_n_d1 <= ~CLKOUT0_SYN;
        CLKOUT0_SYN_n_d2 <= CLKOUT0_SYN_n_d1;
        CLKOUT0_SYN_n_d3 <= CLKOUT0_SYN_n_d2;
    end

    assign clkout_en = (CLKOUT0_SYN_EN == "TRUE") ? CLKOUT0_SYN_n_d3 : 1'b1;
    assign CLKOUT0   = clkout_en & clkout_0_reg_n;

    //for clkout1
    assign phase1_sel = (DYNAMIC_DUPS1_EN == "TRUE") ? PHASE1 : STATIC_PHASE1;
    assign duty1_sel  = (DYNAMIC_DUPS1_EN == "TRUE") ? DUTY1  : STATIC_DUTY1;

    always @(*)
    begin
        case({phase1_sel,duty1_sel})
            8:   begin
                     phase_adjut_1_time = (clkout_time * 0)/16;
                     inv1 = 0;
                 end
            25:  begin
                     phase_adjut_1_time = (clkout_time * 1)/16;
                     inv1 = 0;
                 end
            42:  begin
                     phase_adjut_1_time = (clkout_time * 2)/16;
                     inv1 = 0;
                 end
            59:  begin
                     phase_adjut_1_time = (clkout_time * 3)/16;
                     inv1 = 0;
                 end
            76:  begin
                     phase_adjut_1_time = (clkout_time * 4)/16;
                     inv1 = 0;
                 end
            93:  begin
                     phase_adjut_1_time = (clkout_time * 5)/16;
                     inv1 = 0;
                 end
            110: begin
                     phase_adjut_1_time = (clkout_time * 6)/16;
                     inv1 = 0;
                 end
            127: begin
                     phase_adjut_1_time = (clkout_time * 7)/16;
                     inv1 = 0;
                 end
            128: begin
                     phase_adjut_1_time = (clkout_time * 8)/16;
                     inv1 = 0;
                 end
            145: begin
                     phase_adjut_1_time = (clkout_time * 1)/16;
                     inv1 = 1;
                 end
            162: begin
                     phase_adjut_1_time = (clkout_time * 2)/16;
                     inv1 = 1;
                 end
            179: begin
                     phase_adjut_1_time = (clkout_time * 3)/16;
                     inv1 = 1;
                 end
            196: begin
                     phase_adjut_1_time = (clkout_time * 4)/16;
                     inv1 = 1;
                 end
            213: begin
                     phase_adjut_1_time = (clkout_time * 5)/16;
                     inv1 = 1;
                 end
            230: begin
                     phase_adjut_1_time = (clkout_time * 6)/16;
                     inv1 = 1;
                 end
            247: begin
                     phase_adjut_1_time = (clkout_time * 7)/16;
                     inv1 = 1;
                 end  
            default: $display ("GTP_PLL error: illegal setting for phase shift");
        endcase
    end

    always @(*)
    begin 
        if(!pll_rstn)
            clkout_1_reg <= 1'b0;
        else
            if(inv1)
                clkout_1_reg <= #phase_adjut_1_time (~clkout_reg)&clk_valid;
            else
                clkout_1_reg <= #phase_adjut_1_time clkout_reg;
    end

    assign clkout_1_reg_n = ~clkout_1_reg;

    reg CLKOUT1_SYN_n_d1;
    reg CLKOUT1_SYN_n_d2;
    reg CLKOUT1_SYN_n_d3;
    initial
    begin
        CLKOUT1_SYN_n_d1 = 1'b0;
        CLKOUT1_SYN_n_d2 = 1'b0;
        CLKOUT1_SYN_n_d3 = 1'b0;
    end

    always @(negedge clkout_1_reg_n)
    begin
        CLKOUT1_SYN_n_d1 <= ~CLKOUT1_SYN;
        CLKOUT1_SYN_n_d2 <= CLKOUT1_SYN_n_d1;
        CLKOUT1_SYN_n_d3 <= CLKOUT1_SYN_n_d2;
    end

    assign clkout1_en = (CLKOUT1_SYN_EN == "TRUE") ? CLKOUT1_SYN_n_d3 : 1'b1;
    assign CLKOUT1    = clkout1_en & clkout_1_reg_n;

    //for clkout2
    assign phase2_sel = (DYNAMIC_DUPS2_EN == "TRUE") ? PHASE2 : STATIC_PHASE2;
    assign duty2_sel  = (DYNAMIC_DUPS2_EN == "TRUE") ? DUTY2  : STATIC_DUTY2;

    always @(*)
    begin
        case({phase2_sel,duty2_sel})
            8:   begin
                     phase_adjut_2_time = (clkout_time * 0)/16;
                     inv2 = 0;
                 end
            25:  begin
                     phase_adjut_2_time = (clkout_time * 1)/16;
                     inv2 = 0;
                 end
            42:  begin
                     phase_adjut_2_time = (clkout_time * 2)/16;
                     inv2 = 0;
                 end
            59:  begin
                     phase_adjut_2_time = (clkout_time * 3)/16;
                     inv2 = 0;
                 end
            76:  begin
                     phase_adjut_2_time = (clkout_time * 4)/16;
                     inv2 = 0;
                 end
            93:  begin
                     phase_adjut_2_time = (clkout_time * 5)/16;
                     inv2 = 0;
                 end
            110: begin
                     phase_adjut_2_time = (clkout_time * 6)/16;
                     inv2 = 0;
                 end
            127: begin
                     phase_adjut_2_time = (clkout_time * 7)/16;
                     inv2 = 0;
                 end
            128: begin
                     phase_adjut_2_time = (clkout_time * 8)/16;
                     inv2 = 0;
                 end
            145: begin
                     phase_adjut_2_time = (clkout_time * 1)/16;
                     inv2 = 1;
                 end
            162: begin
                     phase_adjut_2_time = (clkout_time * 2)/16;
                     inv2 = 1;
                 end
            179: begin
                     phase_adjut_2_time = (clkout_time * 3)/16;
                     inv2 = 1;
                 end
            196: begin
                     phase_adjut_2_time = (clkout_time * 4)/16;
                     inv2 = 1;
                 end
            213: begin
                     phase_adjut_2_time = (clkout_time * 5)/16;
                     inv2 = 1;
                 end
            230: begin
                     phase_adjut_2_time = (clkout_time * 6)/16;
                     inv2 = 1;
                 end
            247: begin
                     phase_adjut_2_time = (clkout_time * 7)/16;
                     inv2 = 1;
                 end
            default: $display ("GTP_PLL error: illegal setting for phase shift");
        endcase
    end

    always @(*)
    begin 
        if(!odiv_rstn)
            clkout_2_reg <= 1'b0;
        else
            if(inv2)
                clkout_2_reg <= #phase_adjut_2_time (~clkout_reg)&clk_valid;
            else
                clkout_2_reg <= #phase_adjut_2_time clkout_reg;
    end

    always @(posedge clkout_reg or negedge odiv_rstn)
    begin
        if(!odiv_rstn)
            count_o2 <= 1;
        else
            if(count_o2 == ratio2_set_int)
                count_o2 <= 1;
            else
                count_o2 <= count_o2+1;
    end

    always @(posedge clkout_reg or negedge odiv_rstn)
    begin
        if(!odiv_rstn)
            clkout_div_reg2 <= 1'b0;
        else
            if(count_o2 <= ratio2_set_int/2)
                clkout_div_reg2 <= 1'b1;
            else
                clkout_div_reg2 <= 1'b0;
    end

    assign CLKOUT2_sel = (CLKOUT2_SEL == 0) ? ~clkin_reg :
                         (CLKOUT2_SEL == 1) ? ~clkout_div_reg2 :
                         (CLKOUT2_SEL == 2) ? clkout_2_reg : 1'b1;

    assign clkout_2_reg_n = ~CLKOUT2_sel;

    reg CLKOUT2_SYN_n_d1;
    reg CLKOUT2_SYN_n_d2;
    reg CLKOUT2_SYN_n_d3;
    initial
    begin
        CLKOUT2_SYN_n_d1 = 1'b0;
        CLKOUT2_SYN_n_d2 = 1'b0;
        CLKOUT2_SYN_n_d3 = 1'b0;
    end

    always @(negedge clkout_2_reg_n)
    begin
        CLKOUT2_SYN_n_d1 <= ~CLKOUT2_SYN;
        CLKOUT2_SYN_n_d2 <= CLKOUT2_SYN_n_d1;
        CLKOUT2_SYN_n_d3 <= CLKOUT2_SYN_n_d2;
    end

    assign clkout2_en = (CLKOUT2_SYN_EN == "TRUE") ? CLKOUT2_SYN_n_d3 : 1'b1;
    assign CLKOUT2    = clkout2_en & clkout_2_reg_n;

    //for clkout3
    assign phase3_sel = (DYNAMIC_DUPS3_EN == "TRUE") ? PHASE3 : STATIC_PHASE3;
    assign duty3_sel  = (DYNAMIC_DUPS3_EN == "TRUE") ? DUTY3  : STATIC_DUTY3;

    always @(*)
    begin
        case({phase3_sel,duty3_sel})
            8:   begin
                     phase_adjut_3_time = (clkout_time * 0)/16;
                     inv3 = 0;
                 end
            25:  begin
                     phase_adjut_3_time = (clkout_time * 1)/16;
                     inv3 = 0;
                 end
            42:  begin
                     phase_adjut_3_time = (clkout_time * 2)/16;
                     inv3 = 0;
                 end
            59:  begin
                     phase_adjut_3_time = (clkout_time * 3)/16;
                     inv3 = 0;
                 end
            76:  begin
                     phase_adjut_3_time = (clkout_time * 4)/16;
                     inv3 = 0;
                 end
            93:  begin
                     phase_adjut_3_time = (clkout_time * 5)/16;
                     inv3 = 0;
                 end
            110: begin
                     phase_adjut_3_time = (clkout_time * 6)/16;
                     inv3 = 0;
                 end
            127: begin
                     phase_adjut_3_time = (clkout_time * 7)/16;
                     inv3 = 0;
                 end
            128: begin
                     phase_adjut_3_time = (clkout_time * 8)/16;
                     inv3 = 0;
                 end
            145: begin
                     phase_adjut_3_time = (clkout_time * 1)/16;
                     inv3 = 1;
                 end
            162: begin
                     phase_adjut_3_time = (clkout_time * 2)/16;
                     inv3 = 1;
                 end
            179: begin
                     phase_adjut_3_time = (clkout_time * 3)/16;
                     inv3 = 1;
                 end
            196: begin
                     phase_adjut_3_time = (clkout_time * 4)/16;
                     inv3 = 1;
                 end
            213: begin
                     phase_adjut_3_time = (clkout_time * 5)/16;
                     inv3 = 1;
                 end
            230: begin
                     phase_adjut_3_time = (clkout_time * 6)/16;
                     inv3 = 1;
                 end
            247: begin
                     phase_adjut_3_time = (clkout_time * 7)/16;
                     inv3 = 1;
                 end
            default: $display ("GTP_PLL error: illegal setting for phase shift");
        endcase
    end

    always @(*)
    begin
        if(!pll_rstn)
            clkout_3_reg <= 1'b0;
        else
            if(inv3)
                clkout_3_reg <= #phase_adjut_3_time (~clkout_reg)&clk_valid;
            else
                clkout_3_reg <= #phase_adjut_3_time clkout_reg;
    end

    always @(posedge clkout_reg or negedge odiv_rstn)
    begin
        if(!odiv_rstn)
            count_o3 <= 1;
        else
            if(count_o3 == ratio3_set_int)
                count_o3 <= 1;
            else
                count_o3 <= count_o3+1;
    end

    always @(posedge clkout_reg or negedge odiv_rstn)
    begin     
        if(!odiv_rstn)
            clkout_div_reg3 <= 1'b0;
        else
            if(count_o3 <= ratio3_set_int/2)
                clkout_div_reg3 <= 1'b1;
            else
                clkout_div_reg3 <= 1'b0;
    end

    always @(posedge inner_clk or negedge pll_rstn)
    begin
        if(!pll_rstn)
        begin
            clk_vco_time = 0;
            div125_time_div2 = 0;
            div125_valid <= 0;
        end
        else
            if(clkout_lock && (CLKOUT3_DIV125_M >= 1))
            begin
                clk_vco_time = ((clkin_time * ratioi_set_int)/ratiof_set_int)/total_ratio_int/ratio_set_int ;
                div125_time_div2 = clk_vco_time*(CLKOUT3_DIV125_M + CLKOUT3_DIV125_N*0.125);
                div125_valid <= clkout_lock;
            end
    end

    always @(div125 or div125_valid or odiv_rstn)
    begin
        if(!odiv_rstn)
            div125 <= 1'b1;
        else
            if(clkout_lock)
                div125 <= #div125_time_div2 ~div125;
    end

    always @(*)
    begin   
        if(!odiv_rstn)
            div125_reg = 1'b0;
        else
            div125_reg = div125&div125_valid;
    end

    assign CLKOUT3_sel = (CLKOUT3_SEL == 0) ? ~clkin_reg :
                         (CLKOUT3_SEL == 1) ? ~clkout_div_reg3 :
                         (CLKOUT3_SEL == 2) ? clkout_3_reg : div125_reg;

    assign clkout_3_reg_n = ~CLKOUT3_sel;

    reg CLKOUT3_SYN_n_d1;
    reg CLKOUT3_SYN_n_d2;
    reg CLKOUT3_SYN_n_d3;
    initial
    begin
        CLKOUT3_SYN_n_d1 = 1'b0;
        CLKOUT3_SYN_n_d2 = 1'b0;
        CLKOUT3_SYN_n_d3 = 1'b0;
    end

    always @(negedge clkout_3_reg_n)
    begin
        CLKOUT3_SYN_n_d1 <= ~CLKOUT3_SYN;
        CLKOUT3_SYN_n_d2 <= CLKOUT3_SYN_n_d1;
        CLKOUT3_SYN_n_d3 <= CLKOUT3_SYN_n_d2;
    end

    assign clkout3_en = (CLKOUT3_SYN_EN == "TRUE") ? CLKOUT3_SYN_n_d3 : 1'b1;
    assign CLKOUT3    = clkout3_en & clkout_3_reg_n;

    //for clkout4
    assign phase4_sel = (DYNAMIC_DUPS4_EN == "TRUE") ? PHASE4 : STATIC_PHASE4;
    assign duty4_sel  = (DYNAMIC_DUPS4_EN == "TRUE") ? DUTY4  : STATIC_DUTY4;

    always @(*)
    begin
        case({phase4_sel,duty4_sel})
            8:   begin
                     phase_adjut_4_time = (clkout_time * 0)/16;
                     inv4 = 0;
                 end
            25:  begin
                     phase_adjut_4_time = (clkout_time * 1)/16;
                     inv4 = 0;
                 end
            42:  begin
                     phase_adjut_4_time = (clkout_time * 2)/16;
                     inv4 = 0;
                 end
            59:  begin
                     phase_adjut_4_time = (clkout_time * 3)/16;
                     inv4 = 0;
                 end
            76:  begin
                     phase_adjut_4_time = (clkout_time * 4)/16;
                     inv4 = 0;
                 end
            93:  begin
                     phase_adjut_4_time = (clkout_time * 5)/16;
                     inv4 = 0;
                 end
            110: begin
                     phase_adjut_4_time = (clkout_time * 6)/16;
                     inv4 = 0;
                 end
            127: begin
                     phase_adjut_4_time = (clkout_time * 7)/16;
                     inv4 = 0;
                 end
            128: begin
                     phase_adjut_4_time = (clkout_time * 8)/16;
                     inv4 = 0;
                 end
            145: begin
                     phase_adjut_4_time = (clkout_time * 1)/16;
                     inv4 = 1;
                 end
            162: begin
                     phase_adjut_4_time = (clkout_time * 2)/16;
                     inv4 = 1;
                 end
            179: begin
                     phase_adjut_4_time = (clkout_time * 3)/16;
                     inv4 = 1;
                 end
            196: begin
                     phase_adjut_4_time = (clkout_time * 4)/16;
                     inv4 = 1;
                 end
            213: begin
                     phase_adjut_4_time = (clkout_time * 5)/16;
                     inv4 = 1;
                 end
            230: begin
                     phase_adjut_4_time = (clkout_time * 6)/16;
                     inv4 = 1;
                 end
            247: begin
                     phase_adjut_4_time = (clkout_time * 7)/16;
                     inv4 = 1;
                 end
            default: $display ("GTP_PLL error: illegal setting for phase shift");
        endcase
    end

    always @(*)
    begin 
        if(!pll_rstn)
            clkout_4_reg <= 1'b0;
        else
            if(inv4)
                clkout_4_reg <= #phase_adjut_4_time (~clkout_reg)&clk_valid;
            else
                clkout_4_reg <= #phase_adjut_4_time clkout_reg;
    end

    always @(posedge clkout_reg or negedge odiv_rstn)
    begin
        if(!odiv_rstn)
            count_o4 <= 1;
        else
            if(count_o4 == ratio4_set_int)
                count_o4 <= 1;
            else
                count_o4 <= count_o4+1;
    end

    always @(posedge clkout_reg or negedge odiv_rstn)
    begin
        if(!odiv_rstn)
            clkout_div_reg4 <= 1'b0;
        else
            if(count_o4 <= ratio4_set_int/2)
                clkout_div_reg4 <= 1'b1;
            else
                clkout_div_reg4 <= 1'b0;
    end

    reg [32:0] cnt_33;

    always @(negedge clkout_div_reg4 or negedge odiv_rstn)
    begin
        if(!odiv_rstn)
            cnt_33 <= 0;
        else
            cnt_33 <= cnt_33 + CLKOUT4_DIV32BIT_K;
    end

    assign div32bit_reg = cnt_33[32];

    assign CLKOUT4_sel = (CLKOUT4_SEL == 0) ? ~clkin_reg :
                         (CLKOUT4_SEL == 1) ? ~clkout_div_reg4 :
                         (CLKOUT4_SEL == 2) ? clkout_4_reg : div32bit_reg;

    assign clkout_4_reg_n = ~CLKOUT4_sel;

    reg CLKOUT4_SYN_n_d1;
    reg CLKOUT4_SYN_n_d2;
    reg CLKOUT4_SYN_n_d3;
    initial
    begin
        CLKOUT4_SYN_n_d1 = 1'b0;
        CLKOUT4_SYN_n_d2 = 1'b0;
        CLKOUT4_SYN_n_d3 = 1'b0;
    end

    always @(negedge clkout_4_reg_n)
    begin
        CLKOUT4_SYN_n_d1 <= ~CLKOUT4_SYN;
        CLKOUT4_SYN_n_d2 <= CLKOUT4_SYN_n_d1;
        CLKOUT4_SYN_n_d3 <= CLKOUT4_SYN_n_d2;
    end

    assign clkout4_en = (CLKOUT4_SYN_EN == "TRUE") ? CLKOUT4_SYN_n_d3 : 1'b1;
    assign CLKOUT4    = clkout4_en & clkout_4_reg_n;
endmodule




//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library: General technology primitive
// Filename: GTP_IMDES8.v
//
// Functional description:
//
// Parameter description:
//
// Port description:
//
// Revision:
//
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps

module GTP_IMDES8 #(
parameter GRS_EN = "TRUE", //"TRUE"; "FALSE"
parameter LRS_EN = "TRUE",  //"TRUE"; "FALSE"
parameter DPI_EN = "FALSE"  //"TRUE"; "FALSE"
)(
output  [7:0] Q,
output [1:0] DPI_STS,
input [1:0] DPI_CTRL,
input DPI_STS_CLR_N, 
input PADI,
input ICLK,
input DESCLK,
input RCLK,
input [2:0] IFIFO_WADDR,
input [2:0] IFIFO_RADDR,
input RST
);

//synthesis translate_off

wire [7:0] PADI_D;
reg DPI_P;
reg [1:0] DPI_STS_R;
reg DPI_N_reg;
wire COMP_BEFORE;
wire COMP_AFTER;
wire COMP_BEFORE_D;
wire COMP_AFTER_D;
wire PD_BEFORE;
wire PD_AFTER;
wire DPI_BEFORE_POS_REG_T;
wire DPI_AFTER_POS_REG_T;
wire DPI_BEFORE_NEG_REG_T;
wire DPI_AFTER_NEG_REG_T;
wire AFTER_POS;
wire BEFORE_POS;
wire AFTER_NEG;
wire BEFORE_NEG;
reg DPI_BEFORE;
reg DPI_AFTER;
reg DPI_BEFORE_POS_REG;
reg DPI_BEFORE_NEG_REG;
reg DPI_AFTER_POS_REG;
reg DPI_AFTER_NEG_REG;
reg [7:0] PADI_POS_fifo;
reg [7:0] PADI_NEG_fifo;
reg [7:0] Q_reg;
reg [7:0] shift_reg;
wire capture_en;
reg [7:0] capture_reg;
reg [1:0] cnt;

assign global_rstn = (GRS_EN == "TRUE") ? GRS_INST.GRSNET : 1'b1;
assign lsr_rstn = LRS_EN == "TRUE" ? (~RST) : 1'b1;


assign  #0.05 PADI_D[0] =  PADI;
assign  #0.05 PADI_D[1] =  PADI_D[0];
assign  #0.05 PADI_D[2] =  PADI_D[1];
assign  #0.05 PADI_D[3] =  PADI_D[2];
assign  #0.05 PADI_D[4] =  PADI_D[3];
assign  #0.05 PADI_D[5] =  PADI_D[4];
assign  #0.05 PADI_D[6] =  PADI_D[5];
assign  #0.05 PADI_D[7] =  PADI_D[6];

assign PADI_SAMPLE = (DPI_EN == "TRUE") ? PADI_D[3] : PADI;

always @(posedge ICLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_P <= 0;
   else if (!lsr_rstn)
      DPI_P <= 0;
   else
      DPI_P <= PADI_SAMPLE;
end

always @(negedge ICLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_N_reg <= 0;
   else if (!lsr_rstn)
      DPI_N_reg <= 0;
   else 
      DPI_N_reg <= PADI_SAMPLE;
end

always @(*) begin
   case (DPI_CTRL[1:0])
      2'd0:    begin DPI_BEFORE = PADI_D[2];  DPI_AFTER = PADI_D[4]; end
      2'd1:    begin DPI_BEFORE = PADI_D[1];  DPI_AFTER = PADI_D[5]; end
      2'd2:    begin DPI_BEFORE = PADI_D[0];  DPI_AFTER = PADI_D[6]; end
      default: begin DPI_BEFORE = PADI;       DPI_AFTER = PADI_D[7]; end
   endcase
end

always @(posedge ICLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_BEFORE_POS_REG <= 0;
   else if (!lsr_rstn)
      DPI_BEFORE_POS_REG <= 0;
   else   
      DPI_BEFORE_POS_REG <= DPI_BEFORE;
end

always @(negedge ICLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_BEFORE_NEG_REG <= 0;
   else if (!lsr_rstn)
      DPI_BEFORE_NEG_REG <= 0;
   else     
      DPI_BEFORE_NEG_REG <= DPI_BEFORE;
end


always @(posedge ICLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_AFTER_POS_REG <= 0;
   else if (!lsr_rstn)
      DPI_AFTER_POS_REG <= 0;
   else   
      DPI_AFTER_POS_REG <= DPI_AFTER;
end


always @(negedge ICLK or negedge global_rstn or negedge lsr_rstn) begin
   if (!global_rstn)
      DPI_AFTER_NEG_REG <= 0;
   else if (!lsr_rstn)
      DPI_AFTER_NEG_REG <= 0;
   else     
      DPI_AFTER_NEG_REG <= DPI_AFTER;
end

assign BEFORE_POS = DPI_BEFORE_POS_REG_T ^ DPI_P;
assign DPI_BEFORE_POS_REG_T = (DPI_EN == "TRUE") ? DPI_BEFORE_POS_REG : 0;

assign AFTER_POS = DPI_AFTER_POS_REG_T ^ DPI_P;
assign DPI_AFTER_POS_REG_T = (DPI_EN == "TRUE") ? DPI_AFTER_POS_REG : 0;

assign BEFORE_NEG = DPI_BEFORE_NEG_REG_T ^ DPI_N_reg;
assign DPI_BEFORE_NEG_REG_T = (DPI_EN == "TRUE") ? DPI_BEFORE_NEG_REG : 0;

assign AFTER_NEG = DPI_AFTER_NEG_REG_T ^ DPI_N_reg;
assign DPI_AFTER_NEG_REG_T = (DPI_EN == "TRUE") ? DPI_AFTER_NEG_REG : 0;


assign COMP_BEFORE = BEFORE_POS || BEFORE_NEG;
assign COMP_AFTER = AFTER_POS || AFTER_NEG;

assign #0.1 COMP_BEFORE_D = COMP_BEFORE;
assign #0.1 COMP_AFTER_D = COMP_AFTER;

assign PD_BEFORE = COMP_BEFORE && COMP_BEFORE_D;
assign PD_AFTER = COMP_AFTER && COMP_AFTER_D;

always @(posedge DPI_STS_CLR_N or negedge global_rstn or negedge lsr_rstn or posedge PD_BEFORE) begin
   if (!global_rstn)
      DPI_STS_R[0] <= 0;
   else if (!lsr_rstn)
      DPI_STS_R[0] <= 0;
   else if (PD_BEFORE)     
      DPI_STS_R[0] <= 1'b1;
   else
      DPI_STS_R[0] <= 1'b0;
end

always @(posedge DPI_STS_CLR_N or negedge global_rstn or negedge lsr_rstn or posedge PD_AFTER) begin
   if (!global_rstn)
      DPI_STS_R[1] <= 0;
   else if (!lsr_rstn)
      DPI_STS_R[1] <= 0;
   else if (PD_AFTER)     
      DPI_STS_R[1] <= 1'b1;
   else
      DPI_STS_R[1] <= 1'b0;
end

assign DPI_STS[0] = DPI_STS_R[0];
assign DPI_STS[1] = DPI_STS_R[1];

always @(negedge ICLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      PADI_POS_fifo <= 0;
   else if (!lsr_rstn)
      PADI_POS_fifo <= 0;
   else
      PADI_POS_fifo[IFIFO_WADDR] <= DPI_P;

always @(negedge ICLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      PADI_NEG_fifo <= 0;
   else if (!lsr_rstn)
      PADI_NEG_fifo <= 0;
   else
      PADI_NEG_fifo[IFIFO_WADDR] <= PADI_SAMPLE;   
         
always @(posedge DESCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      shift_reg <= 0;
   else if (!lsr_rstn)
      shift_reg <= 0;
   else
      shift_reg <= {PADI_NEG_fifo[IFIFO_RADDR], PADI_POS_fifo[IFIFO_RADDR], shift_reg[7:2]};

always @(posedge DESCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn) begin
      cnt       <= 0;
   end
   else if (!lsr_rstn) begin
      cnt       <= 0;
   end
   else begin
      cnt       <= cnt + 1;
   end
   
assign capture_en = cnt == 3;

always @(posedge DESCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      capture_reg <= 0;
   else if (!lsr_rstn)
      capture_reg <= 0;
   else if (capture_en)
      capture_reg <= shift_reg;
      
always @(posedge RCLK or negedge global_rstn or negedge lsr_rstn)
   if (!global_rstn)
      Q_reg <= 0;
   else if (!lsr_rstn)
      Q_reg <= 0;
   else
      Q_reg <= capture_reg;      

assign Q = Q_reg;  

//synthesis translate_on

endmodule




