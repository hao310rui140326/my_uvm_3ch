`protected128
P]NN[O>W#][=% >;S+\0;[N7#N@OWFX"R$YTZ8^W=D-MQIDQR\:B<L*@_O- +*<J^
PB[1)7/T-+Q:'T21;^8=\/U80J?)=_&?+'Y<PK+YXJLEW?Z&Q/<),;7EAUQ3?S GK
P:M,WM#6'ME@% )[*58;0^>ECK9V=SL%RWQ[Q;[LKKH&ODF-F$59G'_(SSH9>7=^V
PNG8PJYJUFS*533<WZ3Y>F0[@:KD>VR'S/Y+:(,!+M3\&YU#M3\J@1S6'^^\&W*5C
P+-@>ZS&,J:$ 0@DM@L'R,6[T_,Z8:7Z8XV%;A%S''%J_#N-KW@C2I&X0*R!QRJYR
P]5!5<EHS[S(;^.OW_21]"FXLX^O48I,?DQ32*UV8='WS)'H3*2<67#X&D")H?6 C
P$O<-B<A5BF4G!FW16FYTW\B*&@V(O9?]]L$Q!07_URV=<SJV_@Y%;&_$J+1F">AL
PFO4O82AY=JG9?:VOMR7G<!/535/LBJSH8?GDKSN[ZZ6V)7G28#"\'\RM&G.16<F8
PY&V[,M/.)G=91%FIH;(36?]>IX +],SU;J1H@S?P)6AZ"O:1!X\R+#,OZ24WTR&=
P7Q$OX/AK.6&#B+I3E6@/NJ[$^F#*Z,0V0CDC#L>^D*U>Y0A?>C'18JYJ !I*B-5"
PQ!@NI+J?^\F)**.2/#B+6V$\K0I)H&LX6&=/(C3PVZ"+1H$^2^)TCA,@G7T)>;SI
P8G"?!QZ%99Q]L(3YC-9=.L]B!OQ/<5^\Z-Z[DM8M/G3L(XH.'"1;@,CSMZXWB 0C
PJZ!/+.C./78N8IQJ\CRL(1^WD:^.&6,Q"C>0AS1K?Y7&I-%]2Q+/=CP-D,&U'RRU
PC"\(ZJ(C?D2F\/FHNXN^5!;9Z_D(J0W;DF?0JX(VTL6W:S=%_;S,_AAB(-?O59BK
P:*?Q&OPHO\P (N*X.OUA%$0"^L B50:/:=DKZ?5.,@-EP)J %.DG K>S#GGNN4>6
P;Z"/IVYMSR?4'K,US/9#]\D]:$6]2,E.5_%A6=M'V&>X$FL @8$BXZ.A"!!BXHEW
PH[PK!L_T5MA3-4Q?.C-3R#A3J$.: E^)P&^+==AV5?0P^GC4+_"XK4<2(-CJY;,;
P%_HS25*KXYTA-TM@.B"^_X-9V.?>8&CAH9$,@GTPNZO=NKX3.T(7#;( /!@,.^<D
P$B'($)SL2/2 =YA9,M'1'[Z0!_;KL=C51LO828']* I)X.E"X0\LTWO._: A2FWV
PHM#__SP"]P]XE.H.,<Z8EO#4O$3%BM.S7;-\^FO?\TWEW>Z9K.=2.UD9"1;4;R)Z
PIN6;J;\BIE#(UB=0Y=:6K$X..B7[*/[!+C([VV5'6/GB96B#V<#(/"M9"^%<+GY+
P085MZ*ES9/RU5 "'-Y^AT'9JV3\J^2(9T_B#<I>.5BYOX1:8!0H NX0UIIM\@P'T
PN*>E*1+* F;,?5,C*?V3EX?+2N9VHP V]J[#R_!08]()^M?C=J*'V.WGN=2E51[@
PF=I&XVLN0P/REM%I5I)N TRF8'^>JN4Y+3RZ'L9G.>)<&.%YJ5;W75[;F3M='6:Q
PCG=2?&QL^AABJ]3H*Z 2G007E#-+&P><F=KT(]$*[70L*X;J>O*.@7C:W&["R5Q2
P#F8!D,;LUD=Y !3@8J=#'5\4N(WW5@<IR!18/0A89H$D%3^9+AT!K3SBL^T=N$9R
PV03],H'PI=++D0WS;AU!C?;1S]'G@%S<<7)*JH,%+])HPPQ)DP>J4ZG"+5/FV""/
PK'XV7V%YBZB*N>%FIF;%!%]>YRB60@; +^L:9H&]UN[=8$OZSWL^5R21>M\EB5()
P',6^F,2/OUL 66+^I2IKP(R"[]X@PZ(;N9'IZH!@2!P!3%#$ZJF )4/( G$AHN-K
PK%_-LV/%EE _1PXH5&*?0D>N9)'%,*M/*"@F5;T"NRJ50)YB_B9O]I&$>58R)0'1
PU!._26G>TJOUIV&.O(60XZ)7NVA?:B=.ZB?8K]]>2B'-U F[U=L73<(BBQ!D0!*D
PLAC9P I,/S>Z[<GK!A3I"@U52I%<D<(C]E.ZYZ%(7D?=G%.B Z2"']@FO])>>=J"
P\WDYV7TN.-H0R5IK E@F72,LV:,*H.Y1" X"NG3GV1BS7)/YO9S22.+X* ]L=P+-
P4D)PQ@\\]U&CR0+H=N*U+@= SJ0ASCA^^]R[1/J<.G\DX8VX=UN/#MANRMB<=S(/
P4]SBC.14>=)ER;L354?&";9YIA*>&J'E^GE9B\B-)I779WJ:^K=J\X+2Q\7R=0$"
PL"IZ G.*!COU$S+F ,9S/'$\,#4W]D6;LBPNI/<3Q5.<9WRN/M]+3ZSUT4%B4IA6
PV $<@"^=?8,FN&T"5!2]T<C^D#]9(^Q/!ZX,:Q5O&85;;>PI:HO1 P;+#P((][]U
P%+DD:?KH#F'VQU4W5='.7HK7YL\%,[A[0)C^)QP\10!S1PQ@EI] ^0JZ7$J#"A_2
P&\%FS>*.9H4EU*@GL;KC48P,O\MH+WH+*E<1.,5MYL$0UD,0!8H^7E,'71O0[,&;
P+9$S[\1OU[B*U,J*8Q*/NM@KTG%F'+\"O:NKLE'.\??_GH%CN(>0OP>SA,M?H2"%
P"D-,[L"?7*#67F^%]2""S0P_GBYLFME=YIC:0?M$J$^]19H[5XH]"9X>C*#Q'>: 
P36.>9/H]!B:<X:#6#T);H<_:_>AT6FSYQBO$?E[[@D P!/X0[X%4]K3"!7"!E4SW
PIW_?&ED,K0],BC]ZF'6ODN.&R)&X<^6#^/>DM\:61:]U;G/D:,38X&9;1(R=Q2B<
PXJG44+;I?XEI2>F[3OAJ#LTMES0H'0_><5FN66CF^4@S1(?9)@(IVW!;4ZX[TG![
P=;=096U5UM].>>4Q4/W$2QQ/?3J:_)J#+C2\H)?(,-#=JT^&SNZ7'BZNX>'Q?GY2
PU-9"3ZDA#U/PI&&(C\ZFR6%P^@@>U9&]]I."U6JV1:).P@%A86Q%X'&LW7C.1-]3
PQB/MAG[:V.9X(U*,VG8_U35\8A^U<<08^? =^*2B%)^*UC5@X^QWF>48)'-A^058
P*ZX'JB[C/"GH!5B@S<JVSE[VAO934?&X_)QV#8+MA%\;#<UTZK>"#,_^CU"'V%8!
PA*SJV_W"NLYM5*3#&]VZV# R<V)>+3F; >=R!C*E*[SC-50M3JX3+ JMR%K/C'Y:
PZ!^%.E];_?06K,Y \O2?6E!2X_L46$2W:['U.1CM%^&ML_355>"%_3Q4B^*"4DL^
P5_ &R,10FI^+:&(]V1K\-<XP9]I6@8*7I5/#BLY/1.-#CZ/([F2HOHS<2)<2HJV1
P::JUE%9#>VJ5#$A#1.8+1Y1U319V&$;^L3"QZNX]=:'Z#]Z]N-W#A02((-?M/$#5
P>A\:'LZ\&+"8IYI:R SW:@X_L-)2^/AAE"H'!]W$OVK6?: ? PJPZ$<*Y1!B[T:5
P>MO'):V*AT6+W8U"B/S#IYD/-$I*Y59YM;# GD\^25<^"FZ+1IB%'<$D@IGJ#5"(
PZ=I%R+/2 4""=I-V3R#X_;9GHI:-9%'Y$F+B51U>N ?#:=287>?5$JD:UEJ:^-0T
P/.](6BVX>WQH8<T4$R-:5B8:963(908!61=;N,>6)E%28(P<= UL?YX E2E9/F<I
PVUY[\F;E:SUR4.7?L8EHNYO-YX3/^O@WT<T;()?0 K1,4F6A6+^G[7>3>_;TJ/)/
P4IO]Z8*WXZ>MC>:P3N8I4G37&^>#]MJCG&!JWU8IZ/LR-FX&"229ED2:$%^:>*YM
P9@3,A1K+V EL_1-L^257M.V&9?O'N5!_EQ9BU_HQQIU..P3?8@LJ!A5H/?43D3/G
P(UM>Y6 3EJ 4/#-2D?KA8C&.<P*\3P-M.Z2Y]4XW%4]@&Y@C)1T7SQ$U3">K].-3
P#]Y"#LY0Y(UJ0@/2*OOD\O="AS//G!8_>YLL@4$'M-+ J,3]/U2=$TL'Z:U26TJ,
P9OG5%;6S)=)R!@VK!MB-U=4Y5;] B>WN_R G]'$\&71D8(;JYCH85/QBYIN #2^8
PIH,5(/B!UFP[N1?K+#?6&VXAJ!X*$[%8=MN.Y;$L^MI88 0"L!?-%:ZR/^INH\ =
PC:![H>]<_ 7.*=^.S[1#.6<KPMWYB'GUWDM)(K:KB6>$]"[TV.'7]:LW +5'9M6,
PV)N/:O,'_+!>-\+?"*=L' G0U60[=\5:WDAQ:W"$")O@@CT(X2Q27<P"FKME8Y;$
P#"?/6[TWTP,<N)AE?5A^$GD%U"39-/^9BB1X(IG;$-$64ZP_L#AS'$3O;%8ILK N
P)HZ]G!)"'/SP?VS$9E(%X_HD(,1^A SG=K0KP;6&E":Z>47)$)\*"BR;N8&#W+?#
PX 2.=@['<R3MFIE"BK#7+6;J&G)Z?(33J9VBR"QO5!+-OW$S:>!'+KKZZ$4K^,[G
P/KI75CE>)[$N+DR0NO*\YD%FQH,;!=M%*?\M[=)%9P2F?D"XW&IXX:Y@4<6S:_.%
P+@"=Y08ZNG^;F=X"H$EI/B#CK"::B#9#4MFZ1O'_<PU6X=LTCVKU!5F.@(_(KHG'
PZ(83-<AF<\4"X5VIT :C;AT,2Z++'X:ZIVQMW;@-SGJ,,X;AI-?79VW!M.W07[A#
PP-Q*M!PWC)P&!A\50][W_-+K!';U/',-)D?:V/CWXQ-^5_ATMV:91-3J%T7SV-4-
P.QQW+11]< /4)%]E.O<8&E7R(O<V7)#7:XSTI\.G/-&N#,!3 SPBXFZ\J9.D-%-X
PFFJ#G;J3/?),S:88?3/6'E1DPF<9UBY?W\_"8G5&)^5M2#SLOBC&?LWPM@M3Y),M
PX*[#X=?5BWY27?O.[]>27\+D%_A-5'R7K="?;*P$Z4[PMHQ'U#+QFI%"YC?5I[AW
PZ'G,G.8D]/0YNK5L7SVX9I PO2&U87[;&SV0,;T&6V:O+"?7\!+#&%C6*LP^_"C@
P>B?K S=U>]76B+H%"(';2 %H-@UN*UVXL"&/@#AT15S6#9RU,$IA4'W&)?'$DEZM
PTE0-2TX>$AQBR3?C$+*J$J#];"*0W/X18U4,G8JFKA6L]H5GI)62=:_NQA@A01/P
P$K=G"?)UT+1U^HD@B^.7;H@G&O5\ ;2$D(9#(XT&-3=,J70C]OM$V1<*&TT3\H,9
P]RQ_*,:)]BH;;>OL38H9O)EP'RZ723EY_[--.WAM,A$=#?!S6 \T&1L",.?X_T9T
PE3@&1CN*N^C;%F7-/.0B(RH,_F-$WNMI08B\JI%]Z3EO^OH$[ -)"]'6@DR3ZF-\
P;C8;HWC^WJX HK6H[V?]([U(IX=#M"CL%']P<:8@D6MPXZC'G%&F6U,E^P^"A,<D
P-(C)8Q__;T3Z%/6'QYQ#\]D=W]QX80X\#L=^_KDCJ)+T"2N?=JXWB6^(!G$=*Y?_
P]**[AG?B!CSV9E"9]@ !MR:4+T.9]]]X$N%A?IPCF^S\GBD^DG]7DYENA[+G/D<[
P%=]&T+E!F6X$ "W1>W^+'##Q'&F6_85%>[,= Z^,X43I\:0<P6G&<HN154[$S?HE
PF5\92"ZKJ@JG]Z&\K:2S]FFR3E_Z71)"VMY[',6G*^[<IC+.2SRJ(J1&\LU4G<4(
PV;<@ HY]8!)[9SC\Q6'%9O9 94]-EZ9YQZ$T9GIR^N.JPZU+Z E)ZD=-&#M&O2_L
P#F(/8UL6 ":K^V&0#J?-U6NKRXLTS?>ZC7^,Q;)AL52=OTELJ*R<V?CW%=M3FCM'
P1E7)/.+-\!3)V;3./^ZEIAT:$GSE]F,8"Q)P[_JGC% T3/J0/2Y&;I"+=4+P4FC'
P_G16W=+$":=Q5U'-A$;_2@5Z)!?" W^9*>E_MDRP;MH$[IXR1!3J1..-SE,/ V9D
PN[]-2)G?+Q/<78,0'FQ?45<1^#5Q?HUOR\.QI^MF=6J7:O?FU]%&::$MC:&<ZLQZ
PGUJSB9\L[N>Q>@JD=J* \++(/.(-9$L 2KQ\K>]QQBB_I4#W%1&WR"\>G,@X/_J$
P!K+!4CR2$O[E3FTOI];S ]S!ARN0!K0B=";<;.5]U[/)?NO'D2X ,=?'XE*RBEIQ
P$>OP"(OJ),YE2R^?AK#B^[]/BB1#IBKC:TB1@ZS?-ME@>(S;USG,T-A6[#8"L!<0
PBY'*S"U7:XK_1SWE9MR1P;ZJ09/?-2P.K42"037A#=S;E'(QWR$NJX_(!!FE,4CZ
P:"#7[8W"*EY!P=:*:*W+D'>Y7-4P8LZ?N(%[K%+8DU&4)_2BSOM/8B?;WS0 0HJ6
PL7Z"3,%&OH[L4/UU;0&C&/A&=VWXS,6K7R6(N8*\#J+CNJ%JK-Q07+\Q]W#43CHI
P/3C-C'?(S6*QTE(AKOR$494(KNMY[ Y:UYA1C"X?KON1L4W\;;?INB8*NZ=5+\;Y
PBX5)-RWU\IKSTT26X!4L*JD7;&-YW!#7TGA:N>T]6.-=IAU=71.CDV>5P=TRAD];
P*6ST+FWQ+$Y;CQF65_XJ[8O661>JX")]Y+@Y,=>/5WY??FQ^O.1<P-@[R)2JKV+<
P)T8<U==466+MDOOI1AMZ$,EHJSU;-'1+P0I5;<I1&),,8@?=2-/<;MV]YST@O8<+
PM;NS/\:28:G/9NG _#Q=D47BI+6F(X*XP _4EB1Z#:(*N0\N.;K"Y:O90MK"V!$&
PJ.SV0Y@_V?(NB.E_JDJRB:#K7H6E&$D0+D4\IZFO^KO+6OUZ(DC%S<O!YKGAA[Q=
P:F.N-+$_CW"2 '6&D5J76+M9O(%R:!@XL1[0&,=;]8@,#Q^6YX* S\&%JV"$LB_B
PL-1J=E;@]!\JA''KV ;BI,_+*YF)DJ[_EIJ;@9\06U7XG8^5W5,<7L7D#Q) IEOM
P,  D+-Y.J5CS*<UZ,A[0&#=3=;@D>CFEO03,1\OICKT]NCDSD0B5$A0\,F)$^1E1
PC+)O!Y+@9;F-!-(AY(T $?&=,Q=8V?%8_@20UYWU=_3$F.PZM5<P-,!S\(K;Y'@ 
PQSP N='788]3X9NV"KY/73Y33VVRQ^ Y!"0GE/[/; 8%.T.<6JXB;_T6B=R811=1
PZ\*Z+/J--7N'"=;L/PU5/!M+<?SVFI24B*);PW9VKMB&[A.-[XEI0963>+JHQ02Y
P\-X;KL$@SI)+N,/I,@$7&MWV9&;%OB]EE(*/=0*/G^8U@F7I5O<HQYP?J1SWSZ 9
P1OBXO3!=4XT0>0HP%R3I4O2()JW83HMN\A4T3?3U8%$B=/?5&P+=;^>)C==OHF2$
P%CYL((F@_BDU$3#]FJ*VZC4YC*@(>OV"=;(PY).8&Z3 \9NUQ\DRN1TE%9E\+EU5
PO[MUF>^;K8]CJ[^Q^!#17[<?9!8AS(FEB^5+]N#;B(?7>&RUGC_Z8)Z1.O^K1TN#
P0PT9-5YEQS.K 5$/%  F-G!S[F;GQL,EYM[*/E?;0IV=49D[)?I6+67 <IC=%;RM
P1%^FPS5%<1OF\?%\#3GYK?WU \7W!F%@/6SM"F6_$76)= *N!&:^\I ^("H3;O*?
P.'+6_#A4^NX-,QF=RA6SU</"WF:]"9U$48O$$\[R1P ,% R$1.]UXW!XCM][E/L5
P[]XA^AE*:&^S-W<#G $(/9@8V7W%O+5R!\A;K(N#PHK2?Q897.JQO>%2.541:NN\
PGM6AEJ^1%!B?(A<)GL]%G-!)RAP?@K>*3TRCTVYI,%10R%Z9GN$#"3\6Z6O(5RF.
P>00#,&5TH!04;A!Z:BS#Y$ ^%V':J=D 6FRT;[$M:K[]Q&?L]!A!/BC7QT2RCB[+
PVCFNG_%Y/IUTD8,K2=Q,@9W ?\N4?5DR8FHPQ_ \TC@_3G"26*0HG@N>FH.:?'*#
PP#A21[UP?6<8PHJN0:;5R>)VQQ0XK?=>H9A9%_I3;''ZW>&*-#^ 5P;GU8<*K7P\
PB!O&&:6:V.-=T\,EM' R_+;4430S:6A5STI#,%-GP^(O?#V_LXAET4DUW5D?/I:6
P8&AN!MURD7'[AQ-![36,3;-:JJ.%XV$W=@1A ;-"SI6(_ZDJ4;[Y@2D.;^'"2HD]
PT*[%[W>]_#$R,\LJ]#A/RMB_, 6 "_YAK9.$A999-!"3BCZSLT^,IYUJ"%UU9&$N
PP*D[R?6%86S(BT:YX]#,$7I+&G%\<$41DO5@&06N,BFKN+IQ'MMH4-J&&[2)W=F+
PL<1,JWO(RR9[ST>N"&A-LW$1P89RB?.4-R@, ?1@O9+6X!ME5.XEM-_SB%FAE)S_
PHN!U>*#\:GSH.H<\^*#\#!UNYT8D>BS*[ [G-2KJPDD22FX6JL^'CXZ$7,<;;[6A
P5)$#-%(.)S5^!;+S)(*ZBB2$B[\9$*)8G:NE09*X /(I*(C(!13=2$!+AL.#3O%J
P:R%@>DDMG\K5?B?@%V%" HZS;4>6'RXV>-$:>RZ57AL5-&)"(10;[LL@22H%&M$;
POM;,-3N;=QE:.@\8G*;L<,Y@  820PK,]SVP:E=_7U7:-2N+2YR/KC9^8.1)&V,V
P/>1T(W)UK%R#I&--I'W3\[5:0(6I++U!1P<+#UB^%Z8"?9:&00B_4B)M<O>OQ/7*
P*G1,0I!M-3*0U2V2B)&8N0F\NGD %%@O+( _I*3%"7#'__A4:DV"7#/KOWC*E8H.
P8P@D2>(6OBN:_<ZQ5H1'JUQU8"A?/\*4%+M1U-YH)A0PH=;1I\3T<8*/:XT98@<V
P#ZKT*-6VWWRCL;:W&$\[HN:QIB&4Q=&SF@WH.B+?592P4T@OP8XP4?LWJZL9?-L#
P)_6\]H'"&.WGF)C.N"X/:JV!L2205P?!S8E008XEWG<%E4NW^^R?#->F)0:#H%*$
PA1.K/\;\$1F'1?^H05>]#Q""[V0>_$"Y%7VWT8;=(6?AVFUT0F:6KOZ#V0=5"RLU
PP6GE!$T>NZZ/2V,EL&='--(_>X#'C7%8PR?)"846(55<,,5USMA3B<XE5P:)0"$>
PS5TY M#A9_QFE6U&A!S(S6^G+%!6S?1!ULM"B\\W-IQ:4L .M.":IB5;JO*5/G*1
P*;WZ,*E.@CA_^1Q+W+OUEXY+50814B3/?$5.9KIC]@.9'#[PD-;D/]3\)DL'3Y#'
P@84=&=6T^F=&39\2C0J>QT<O\0G1*1J%RM)XU3KNFS]Y+.V7 :I*_A;8;]IR+_ZY
PYW,8[?I/KYFD_'&(9/$'^VN 7LH9:P(^@%2X#?$-J?:RH[;A/22JKDGKG&N/>XP<
P^>&A1K/[F6CW'*2&[$&D:MAVVAJ*^^,97>D^R(E\UP^  M=-I/]:*^I@\;ZL0D W
PFA(_B.(*J"C_;ZK"X-2*5;)I%CTLGC)H!T37UR[V;H"T?>VDRM;\/[C,&+70/(O%
PY^U;3^8[YLS^@DKP6X!8?^,F>L>$11T@3V+A,PEH+Q?#\]E72-QGD;*1Z^KI32%8
PQ\%]BEU6VB4+X7X0<IK#(&R#QI"G'_G3WVX+P!7Y*_*!)SCFLSR*W_^H%T84F4)B
PL\)&<TYC$FJD[9?N[WM^N?O(@IJ+;/BUUPN_"W=%@LC Z90^_,)F4?,4-0H]TC@)
P(IMT'1U:)FE[47=R<%C=\># (YNY+OJJ!_&[/*.0=POL&8D41,+$U $5NWRRP:>H
PYV&!2//V<::,^W?%F Y=[J.@?Z^UV4E<W,K]+2L@W( LKQ"\P"X)+9#7859R->UX
P&T0+;$L'[[9P&#(HB0R"XSRPUQ+GS8U,#S9AB@DHZ1@B#K/\1! .+9S[25PJ'*(Y
PK.W^+^1B^Z-S^&/5-TJTS)!TBY6EN>8A>_-%H:M;4^XYX,L$5W($*1.9M.;EN4T6
PNW5V'M*%.6I4AV"$\<^5U+_#L6Z@#KWD[OW#Z['"*(>0L##D&FOPR.RI4&\U4]'_
P JXE1UKQ0H'++R-IYJV!%J2L7!*Y[^[!?2[TC&B)L71->=CFHN=M@\F$72U!XPR0
P4-CJ@I*!X*O5MD&C4V-?BCNJ_O2Y.7YA%L=R*$5H0W% 5JY7#Y"HNS!U_V&*P_BF
PE8E!BEW);*+_W1BC08["D9C"FC1*>/BNU1%KDGZ5M:LB-MS(+O9(^C=3YC )BK T
PZ"5')-WI89GA$@P4@(G%N/%@+'GV4F3'F<J%%^S<-MV]NF9_PL\W//P@$&MR38^%
P4-B&'1,JC4A.C1)KS]]RJXI+JC^/^U9<VDE^=!'62B!'TT#900E*Y:^9J4U"08*+
PR7VB.[F$N<+ON6-)P\[SN*V]T67R9-3T"YRNGJ=\T'?2J7YL-GKXMQ2WUJG.@ 7=
POH3&M38XD;D$UE3M3]DU"=%J^9NX"X]RI9)M>P\J+3$K.*AAM=359X N*GMT_SSL
PL$R*-N4T4Z@9 ./>?O#_U3--G #/H#IX@LS0'S^9L,ZJOMW7LVK8*;'FG_VFG[R$
PV/O]DF>=T>"QLV-" 7-T3W6N2+C@QO#XJP8>TBX()$TL*I^74W:%I8OZ5#RT\-CR
P1O0)C:4:50ROJ;[XA5CX8Q:.]95P+I=QXM]&^]["RS$37TG)<IZI<[!\^#!-,W:U
P68ZZ_DQN:+IC&J(GW3F*'_5A;P^QQ)Z$S4+=J!?7R@)'//$FU,&9JI<7/"^PC$@4
P<C;).;%@9A2J*7],#N@ICGQG+6[F*?/<<16S0_I1*K]X$#*S99-#F;LLFIE9;EXZ
P]<@1GG'(2%[ =7'$ZO+ K;DSG2+*7TC,Q&T"$T]*HM4647Q;2W?V<X5&@+\<6!S*
P4]H7BH8M6G\V4YV$ !JAICL/C($60:XS DGAX--!(387J* K:R>D2^WG8VTTEQ+9
PC-,_Z,V$FZ<62X:ID[846$Y&<;1\16$:!U0G'[5>T5@H?S:KOZ.$4D.^W?@:A@A3
PY2\6O?#3.GU)ZO<::C,/.D*DRGQZ87A0*'D+/=I_)&NM18B<#W6C(XFV=@+0;9^5
P*E)![D)9QE1@.%Q(>6M03"-BMXR\[\A.MT.*,"E<1OQ@I9:QLE?, )>I!VMXL-^8
PT_SMR= HBP0=\GI]0>[A)(9HPK8N>DF\?GN=_!-[EG:VY@9O?<-P(E,-ZC[@D&EO
PU,GP TY4DRY/$ON*]?F?D1H_L@M[K@<I)5 FF_[@GK-2LZ8?)7* B\"HZ%XHI@U9
P(V' <M"18"*$9*>HQL0(,:,$9,>%-*23KI6Q@+%D(#7U:0S'41Y62!%$P:"KI8!D
P6<6J;L*G@)IJHU-';+1*/?NJ8N>6R&PF-:=B2$QXDU_D88E;[6B[L>A/VQ&JXSRB
PA1QTISY* V1YGLP9>C$V:Z[-;3!)T84BKD]9O;F5?<RQ@Y&M3"H$Q>"Y:_+UL#F&
PF!VDY_2^R;'2=RUJS9Q-<CCKA<%FA+7+ F5J4_4=-]YT"AEJ>Q50:W$4]_4"4'C<
PY#T/1VW431N*0X!= 8N>ACZ@_D G\M4&_?'#*SL=N9@1[6/ \XV2[8 N<W2.<21+
PD>3/[S7P(7;=-6YS9AQ"1- ">(R,,ZIQ5&AU;QQGO!3TR/@^Z:89D!FC\:"7137[
P/A@/C'%9C,C]8<S.$E!IWB,H>4"XCE]E1S3O^DTDB*/]FZ00('N4>:J)<TM+JK%I
PFX2^2.\J$]M4%1Y>T+A?]5P6;/82!S&5:(?5BM,Z2DJWX"O>YS?WUA^=H1%-6NZY
P?,]5!!*-T?8I2\.<8==WX5%A;UJ^))JNELAW"'7]3CVF$:BJO<+U!XA1"U @]M"!
P[NF>[1<[00^IH_#(NX5G@#^9 )\;-N6<Q&(@B6WC:L.Q,C08Q2^^;N.%Q)H-/828
P.N0"^(8I.J9)]AH2!:7] Y#2.1Y&ZR'K13^GTO1#4 "K6\6]T;EH\<.)?1]4^9 B
P,"%?+CDJUIM]RB6UC/H/\>R&UR?KHNZHD6GI;[9YL4EP].RX)]  +J5U4$L&#KF7
PBP/?B8M6L]]6MOB@)%/[MF;66"![._<>M%8X#[_3<%K:@N%IMM"3YBP_E0OT<BT/
P0&L%!_KNVE+)E%A[Q7EW@'-L4'LV"XIU[W_3$H8\A[EL7[E6#?%-7BED>7O/99VJ
PM<&T0*,"A[;#T,1** HUW==#$FV#OR"ENZ !5\E>5-S[P(C=X7.OGCQX4"4,!N52
P1IUQ)59XZ @Y!H,-G.U_I4SO>XJR>&7F0E7**VXT-=OJZ/>]=.(3>D DR4^#-X6:
P5T^/VY!\Z"!>)/Y^L[TGQA7O(VQ"DI +Z*^YK1]081>7?X>;+SJ%&1 !3=.\_06Y
P9-AA_"NJ&[2*GQ?]#Y3F  \6\"(>]C&3*DQ:D%2#&MGN]W6 H.K%N 7,^]PD45=P
PRZTHIGCS+H6IJ:"="<^KN[V/ZM@HA.=^J*:$GD+*Q3#I40X\+NY\[QX#&D?L D =
PE0KQ?).<^6B:;*=$H&+%15_":@<@%68O03%(;<_E1_/52RM1Y;H_4J+T9?$1M=? 
P1#TQ70P3:CE 02(^;')K"W$5%7<J/=(:"&+;[DEVN;1#6/(_P@XIN3;HD^5<$54%
P= ;-/U50 RMPH8I[;JC0: X(@0-*QI>TJ5@^W%M:#!^ H3PC TR#>?1WEPSMFH\F
PS C 3T>88!,+1-F1WK(;\@3#%_+U5;IN*V!5HK)1[Z:P4:#$9LP."SQW"YHPZR@O
P3I<E%.W51-0C3&D4QR+.Q5VH[B7:(G62=0I1?8K835220*=F^$':EP[D'V9?AT%I
PNG"7?J7&<!?Z-UH;-+>:U7^(:6J:)8*SN?_#_B <:4=X=YNPE^%313US3M7[KS/<
P+3L[OG[W#_F9F; :3(6JU38]LZ<S7C0*&%\O2ZC S9C5%L<A[HBX80H ;I;S.DS@
P#N]S>X594G@ UZ&]7A_5@#&)!"<_-:92;N\S&?O#S;?;8?/\_K\?'L5OK:YSU+0T
PD87[;6XG..62(\IS+J_+$(.[!.#\Z7 'K7%IXTYWS')1>8RN "\!I=QOMYDYS?">
PQ'.?D\B?2..WD<1?7S^/>VVC0U=LZSA"."N &!_%^'&)^N\UT0.'Z_O8C=(#3UE+
P'X(R"K2K\J% ;.@Z5B[P1U\%5?O"<I/1G'X[7D(9D)!P#2/<&+)-6:KVK,F';^SL
P!))5CH?;7;VC(_9B"$:EZLMCD6H?899YCGV!UW<HY7Q;]:#A6VN4H+*,@Y$/1^"\
P0UI\98A'MS?!%/()T0_&:.S+,K'@3AOD#!*!F0."9/]R>FTW('?? QU?4C>_K^+1
P83<\_SPPV;V_MDGR-9HX(UFWOF[A<9&"@["A-'UX0]ZWJ6>(<%<-;\GN?7\]NJII
P0ME@7!_VYF7W/\ 0"L.ORF\AQCBCT8CSWT1"-8P-8=YMF%IK8'[EAEQG'["31)'A
P8^<<=%YQ;0E'6W\&>-9_EOIB'E"-GL(H&O0J^DCH-ZK.+]8(K%!# 8=F8^2,-*N;
PB<ACO\<!/_#QZ&I+UXP)F".Z 3H6T:&,=8OIX/%SDN,K%H)0K>'*TD*/U9<"'0.W
P2.,T_\0EE.'!C$]C=J/F9*E1Y6K=OEJ%]7D2$>7K<2BVE7]B:=_0B:A)&8TXR(VK
P?"X L_BD.[ ]GH'88W?>4%-=A^5;2&^/UOVGHC!5:5',%- :;BX@0=.'E>W#(6]J
P!:5"H3_!3X 5QM3ZLY;?<)@S?3$&=9+/=&'.(B<XN+24]C/6YT1B/-704S17EWVR
PBO<LE1Y W-U]<<8"*DKFMLXJ3$>21;>"F:0?5.^DY]C>F$T["5J"1Q1<FU5)H];7
P8Y0VHF)A#&3Z7.BZ)0.2](\VS4\F/_/TN[,#53, J)AB]36Y#_5T360,RGP6 5;,
P(IX[""Y-B^[8#F;/-AZ&=':7BU$JP(H%M+OFGN@PI,;;FEZA<@GK($U]_=-480^.
PB<.W9BS>?6,Z00U&SL)A"T4"-Y8QB\I_,J7G"/5_I"Q6>K(EP:Q.M+VH:=W%3AK3
PZS>/I]?O=$D,I%K4DY?-C0@0.$>%H*>H-"I%.P'$)LO:PO2Q;$RKDA^FV[V<UE4U
PEYYLD21;W4S$.C\=VLZ=*^UU6Z!\9MR #-3F(9 \O(>[\>81L)D/HUL0YUUYEC/F
P#00206:^Z4+C:MJ4<OH_S4V1CO3LZQZ4W11 YXT/QD.(Y6&97*C(4O:5#^/3YU+]
PLV+OG<!QMU4S%S:=%ZT^70"WQ<2_7]/BUK5<D1:BW5>4/CQ"BO-<YW).$8_4_SC,
P86Z(JP>:HP*C:GKE5ERH7!J%:HK%+@PS-FTK]TZOBZEPNR9HH!$_ T<P[9#7==B&
P;]071G>"4$!I'>$@1#Q??M<(I_P?4S >+A>>;XVQ=ZXJ22!T[6!N)5;-3D/S.^?U
P)VT,]O]4R62N""\L7P;*# RU0M[,*[#UA-SS)H(PJ+J2E/]U%SLF''&JI"/.QRT9
P3B#)@'5QIT<>B50UT^+QPM1O5B<]6B70;Y,5A$Z7/:U5= T$((41FFC>N4#,[ G$
PJ-4:)+TB"AD1O-2^4#+J QR$V1IDH_>2/-4F-#GNG"YI*X&4I_MURCO9ANBA"I3!
P62:LBHJX'0P(\AG7,0*)7.Y);.9V2SNK]P4PUT7*E1SAMEGG;@4V0'D.H9_2@/>H
PGJ. 9W2VQY 8[Y3U" V/1U(XL^L#3YYHDL,PZQ@;]3[=PFKYW EUZ@PG.LN]?[?$
PHL^H4@ 5I)@4'-ZWBIZ_]\<1/Q'K[]_D?MJL=\ D7J]*[?_N;3\XJXXSL='?5/#'
PWM2IW?]+3@&QEU6HPX4.(T $UC,(?G)%KZ@A_!"O(=T/=9Q;9PR!T#I-#EZKKB3?
PM!(9'*<^7Z)*L490WP(*#J7KB+5U@*2"> 8*GU7KO>U?I:9W1TU,MPN:H0E.YE[_
PJ.P)&F#[!#HABU=!?I=.:32]E\#D#/2(6#[%O$=5C O5SL_.<6[2+;TZTZ[ V6/*
PVBO()A-?DMN'SP:@#[^_8&L&C:7$G]N$C[998NR,,=CHG@;:!M;W[FKQUE ^+\X>
P?-9B%OSR^ EZ*7X 9?B]5.CC-79R2.UH("$.P;+#8VIA.4-8C]FVQ "'Q4C8E>+T
P^T%2P*;P'#FF:^&?F;'O.6LKT";4O.W58NP-[L"@ZRF82&:$0B9Q8%*LO#!9(!W4
PYA17T+#ES'#8Z8UK['H^K.D7,15LB%\O-67EG/65'0:M?*%#%00U='U(8#>;>'#"
P4G6>0)NE)WV/"@ $!@\-H%DZ*UBY&-"TV[481MWSL:W+CRQ L9\(PSCH!LPX\K7G
P+ 9J%@-UHA\[MF@)C:>R@-,>#MP.9C^PK/6;.DGY&#:0XF^,Q2MY8*G<-&,W;I3D
PXBD"N +@_,_J5Q;GPO'RXDFG$ F(07'AIECHP'\+_N[R/KQ0:9KI>=.XH&/#2*KT
P-'TPY&SKW5*>H:H+/1^ZE0\'9<6?P5B] X^$8K+:*8@Q[VO14T0D]).<<49!U"U+
P,+)0]XWT*P[A<O*YF 6^9@/9ED_NVG*P@#(?Y:IJ"KQ;%X"R<V\&1(Z,V2$?RQ9F
P)]0&_!>G[?W6$LBHW>73,:H10T;<<O7[..7] L7ZLHP<($7 R-PBFY<2@2/V -N?
P_OD=8:,>^P5R/;=R=H-4$(^)G:58[R'D#%Q"BXG]A$NO6(V-C92+-2ON6$0>R%.P
PQW1\C5C'Y_);?F^[CO#V  FNP-K0A=SJC:9IZB1X"B)4?O>6PVRQQ6X@M3CDT:.N
PX"_3]]=:H/0XI5?DJF?G]5I":#)X4(HQ MBD8KNZ\AA$RZV*-J$#E B\0NB1I6D2
P> 9*?@4Y1P.'J/?6\N)];.X* FBU87?Z)@C[,*'"=>YF+C;DQU,63LQ:E'$LW0KE
P[*-/2:+X>>N/<Q)-C+X[7JDYCERK4SJ=A4ND[WJT:-F_$\Q2I(3&(QCKRG.UW%+ 
P!',X_)@&DT%L@BA9KY$A88L^K0_TP"9-IWZ0G_9?/WM_1HH[R9  5FY*%!)B0!AL
P,M2C%V;$02[5(;8'$PP7GDT4&0M*_-%]IM,%SV-D;*.4N#UDBV_]4MN1BC2CK#N-
P($MO__ZK,LR20GQ#HQPOOLGU&<>+>8_2)6E:&1TUR1."EDIKJ<$\ 9,,E#GR9_O>
P"P[F%6S'OKKD8L-OP6*K=ES?(-,W.QMVDBF[FT?_UX_A-/<W&Q7SB( 0[6?(QJ(<
PR++\8YTE:6^@$Z["W!#KJR'K_"4V2U%&1Y-0S<) 4!V[,JIN I"3QAX&Q!(&&D.8
P$]+WWJJQ/_Q0Z]ROW-JIS]4J.+F_BN]@<BX!*\*-[V.G*UB[V(U2]Z'DY06@?<&P
PZ'&!=>16>:M_T)Q$YNP)AWD>0^ L#C6+R;D>FECA+L7<3LO[4V?I*%7?)P\TW3PK
P.6,&HO92BG6>5"P ?4*>#.7F<[1G<R=@7ZD,:[0?H&)=1=J;0)C-O-,B0 %<9N-M
P^0ITL6)N(0VLT*N:Y%Z)Y(EUM_XH$?SHS<37FHWP*+W_9T!3O3)?;55SW>S4(4]6
PYF=8S.2 1I.'N"A9'40K9XE"LIJH>./I+6WH(L--I42VWDW(QZL'M!V)%E F)-O<
P9U7[@%7*)_ADY@K!C1@OO0[SRDPPBKQ)HWV%U%8@=)I'++OC.\<R967+80;??(MX
P!5GH\0A *V>= G]YF8Y,W\+Q"!2CCZ* )1G#"5-_9WFP4-$@9,:NSO3'=_BUH' M
P]47$R65CF\P[ELI[,)"#HY!.R9[C85;B63Z*TBP.JXB\<C4*^M3T1AGD>YV+(\SF
P3 @68"3,;B5]-DF0K?UMVPA_"+@P?@F]*?87AO\G0'CZV*G9R7*_:PATZ(W+ '4@
P=:%Q"]3*S8FWG17V_(T 6!7:]=]G:\SNG-[?#!FCLJ,"_?UM-<!#K=%AVOYEG812
PU&=;J)YU7 9UM]8!&/55V3">]P9S%6LM %_:2#6-W<&Z+5/5#"^TH<:6R0M&["I 
P96KPN7FOJG?@3)=XYM  ;9!8^)L.^.SFSO#ALQ!*A$^ WNLC(H9O/15(R-WXL822
P#P_(2H"X-"1CL%2:MGHVV^U[EG6IOS;7*MSF<EU\Y>?%1/B$[XH":,^ZB7%,9&>[
P);S2<$O:+!WY)3.WN?=.CU#.M]4*J(#JNB?(#<- &:=*7U=(XS'E]"],5N%&IA'&
P<7OU%F=?TGPE3&(_F.Y%2HKZZ?_4@HXS[[H-3H\K)@D<F6/2P PTHN\#WN3<:9.A
P+5)^EP#E#2.)2 :+"T1\8#9> (JN<@A9<F-OX35/NCOT[A0U9JOV9]*$V[J1(SYC
P?8:8]HF/%U5];S!3X.E#6!9H54MJ2I38N8_L55G0*(2.K@0A#EJJ@V&)>F,K(U=1
PG.LB'7UF7&%X+4CU[%Y#;IFB!,!3*A)L*[[QOPQ>Q" "(!6[ZDP>^D]S*(4<8UU+
PW\>>&&2!K@M&M]X/VGNN;[K7U'SIYI+^/(Z:4K)]#76QJ+$N0IK"O3F\3-X4MT<6
P:44&QP<1_'%S3%>252#".E2*ZD;&-5ZF^T))'0U=$/98:T\_"+WL*@?0O82W,GT.
POR$>$QIK8EB$O!^P5/ !.0\DP@(%4(Z\%1745P9K.I(JU(^21=%\I$C\(43>A+]>
P?3W:\&R/DZ_.]"[V%J\V$*4&(W$;B#/ <J";D/ J\"&]4DJK 4X,Y[<DP8>G6.^G
P'OGI!-*/WBN$T%,($^\'E0_E =>%UAL8U]S;RGR9:KG3,!'_UVPCH0.2AM-EO7SN
PC!KZ*HM9*<5X)\5#?K)4*!MFYB?,E*F2$KWQO;>,6/?VFU3)A"5G.@;S"R%"2+YA
PI!/6Y1KD?YM.F52@P-O.56[9@C!5XJS^K1*BM$()Q<?V":"UI(C]J8\VUMQ/+&*D
PE\ DU- ]MABAYQ"@XZN7Q/&CBSF1')DNX/CP=>C=FY@EI-7(\'E/@73EB$DW0]JS
PYL.9UX'A8S^?X9X-07CQZ*W H T3R3.2+6IN1U6.^N.K>5S.E'D2:&_@Z@1U,(NO
PRP)7W;+>VR0M;7"[Z7T$XT"%$GZYA.&*5\=-63D,6U/M%]5NKQ>1&@/Y:HA*Q]X8
PQB-QP^*C,:U*N840N2P05&ZAK4:W,"9\<-]]/=TFTX5Y6U'V^GH@>UG2E$Z!SK^_
P*?0TM+@<%L[MC1#9I02\RV9:=GIZN!IOG\%ZG^-:-=P2(%3K$RASQ:SH3,"20U%*
P98ZOZ00%G#^"QO-E;3T]L;HOA 8/ RG7$5AH7.$!"E6%Z(LN/7835-_)"79'7$[;
PKSC$ZZL!*%6(:H$<V0_;$<N=<%2!-)PV?)TS@")9%X+P^W=R0Q$DRKQ:%!M<7!;Z
PMHV_&$/#M$8C80X$WZOL>^D?I%1!G&?S&AZ2<%I8Z3+;<+ZV7JPI#A=SIA.8>F-!
P@?-L*PBB6P.+-4_K"\R0VJ?6[>IG7>KU7+OZ1ZY7DQ_=\E8?;6B] OGPZVUC,88S
P[:=DF_34D0I!:2?'O6N)*%MA15:Z%%\HE&QV*-$!-V3F6?%:K.59#FMEOMV(U2GJ
PQ[75<>$5E"BWM*M/+.6S#,7O>\<M,5%,=,<)$6.\05@.=S@S%:H6_5#"'!DNIK@W
P/X+QI$EJ5O3RH/D/6.C?'&C=@72+B8<, DR2QT[H#0&P1^EKZQVV:!JN\3QAD=7V
PPB[>I,$M28LP'N:4;U'^<GS4^A)HC6NOG9<15,*#')6/V![P+2U4OI1VEWAO7/R^
P2WXO&HO;9FD\[):??4I[-& F""C9#J3IQ5BN>K%,D8@*,,_,:)<+"Y 6]@]Y,9RN
P*^H;H)@MH5:-]C7C!<I*&]6]+&\F5@1J;,K"1_5T1A=V]T?:/* ?FYLF<[QU)4&7
P6=NOB@V^"0IH3>=5TFX"/ZD)>$15;(KW.!VG-IE&'C_@"(3 '(4NPE(_1@\.LWMN
PS:<B#T9<]<V813QG(ILRZV%Z:O9QXT"VP&\,3W(NMUF_!29M,:Z*EJY;[IR')B\+
P][)R+D/ T:TG_<_?J00=/W0JT[>.U!+$5QKJ9W\T* &ES[1ME.SS@T]YV,A 40\F
P0G-K\T@\X<Z*N8$N:/W(51;(\K64F;CEH!YU_E2_=Y6PC>?8KDVAIH)3=)A;WE_^
PQ#O]8-,D14%%<5<@[0X,($DFM[\U S#V,KJ N>=E_=VWI-,3X/IGC'W(2*M(&/]E
P/@L$Q*&"PM#Y]/:?=;72"[OLD6>FU=2I!BA.MT(3 ,4\H<0^#% -/%+X!XLPP_: 
P[ XXY,6]Y8^1%NW6!WO$,68)K]X7*3[/EG%STT!RAXE?065:AF(1>R;/>.SWY+:0
P3\@TBB_69@BOREB]H72+I"$%M[LA NTLNB2\S"T^-U$2N' W&0/&<KL@MX7:L/)!
PI=X*E7%XYCPMZUDDR=L%SQI>OUM3Y-3^:G%>$.2N$;F4P1! ?L-5Y-P;'(,XD>T'
P6 _4.%X,#:X#;F?:MN.;#NY:Y;Z:=68&B@\XMS_<T2W<)X$/\ZKDEPS0@136"3LV
P5-!-Q<0A7SZ"6XB2T35J1_1&E.T)"!!5&,I;Q Q0M "]8=2)AHYFZ!:92A15E)K:
PRJFBC6^9ZH$DD#GV\B&?6GA7I==JWV>H>=&$[DN(>4DS..&+Y&"?NB8B'O+(U[C'
P04+3A#9]2H%7[UM>/<<9-*2[8]6*(VC#!1*:(!H,:-OFXUJVB_&-MD@P&7CZ$*4P
PO;O4Z?^E)UG+M4-S+TW6LFJ)%>TR#3EUEDU439G)]S+# [[I+X'&-^?WS(7JBJ(C
PE\+>^BZI/!N/@8LL'L;#'2R\+"?)-'P3^XC.5VVS<") 1":E91M_N9M:DL"6I? U
PN1W;*029='U&(U!ODHQRV[J_J:F(@6SB'WKI.XU8C.H=K$1W6DVPJ->Y@FYOX"R0
P!_6U"Y7I,(.I<ESWF](<XTN<#G'E<)5L41-NMTFY;)^7?IQH@+$DP!5(ATAV)J@F
P4_%:Q4\K>.%X^?HBJ41,9TBD><K"'*Y%OL];B!5]+-U!HH:HTI\L$/B2=O'NZ,>]
P=(>H&!H8 LN'1!H+F+<0?Y8FU7D]O_O7<'R8GK.NE!SGEX. W@%X;N#K&<">P5'0
P2(M%N=HQ^%-=ST\$'CU3Y:$?)L/E[6:B5>(=D8@Y;N$579RS=J".)2-S++;[?,^B
PF8U$N2.H7&81G.?^-- /%9!),'O^2UZ-XFU[Z6A]Z29Z!A=J#3!&8Z<M#&?YR&;W
P@_G@K7_?;"\TV"TNQJNG(?0+B^^FNOSRC<<TD:!2@W5R8XL@\+T48@R:RT?0Y+_?
P$V(1A "1U4YLD) 5D8L+="G6<+'7RM'/DR[-B->"X028O@?&-3SX+F\''+OY2C]C
PQVMW#H9(UN.2V06"UTFXDYL:M9(K<F>Y+;4PYU17EY#U*4_B]"<XS[D$N-1GY#0L
PI"+JT"Q,Z84;*/(IOW9K]Q&2B*-@H.%WJ0<@[!G:#%+@"[.'[_TL/<U&+'JJI3F4
PW"_I;AYBXQ0$+'ZS]@CA5QB!FG$C=;J!?$(6$WO*&/[K\A< *<AIJ.'^TM2L0(;\
P1O4&QT!9617X.D7'$ '$WAQRQD+/HND4\D\;TDLL<O2RR?RP&[:IVQPZNP"71!@X
P_4[&<[H?WQ[>X6"@]JT)4?XK":<V*>V-<39TY>:9WH@UUED@L24ZY@]2*<E8)-_@
P11LJ)2S(L0$%AD8FP5RVW#=S57%%V4Y-+0/'I[N<NJU]BC@%:>#MYC"9J.\;T":]
P]R0"R%M'RNS+W)!26PUW;5'*$3<W:+7UZ-#JSF^)Z:@%-"VT6:] :25CJA7I_M_S
P2!4XXJ5-%3+/>6>6MK=84;@_#[MP,"2L>M+5$;JSRP(-'UE0!,]O#]D>U+ 4R?63
P_%NK!2&;XNXL*.D"-_(T88Q^^AL*GY&.C%[$S,ZR@0<L!WH*,7[M-^A1]SZ-Y+C(
P,M3#'&>"-2/RC&LG"#'+S$84*[G& L;>1BXN$LK.GS34$&;L4,$F%DT8\Q7M:GJB
P!BS\G=&P^VX\9!,]=M6.L6\I$.8G6M]56WKA=,,5I)6;6/>VKLN16:MN&.179KS7
P@9Q<+S$=I%V]/J.1%"'#_RNM#U"3\2$\D=;RK+3"%:;(-5>=?1XYN]Y&/_754L0,
PXLQ!W&_TY6;C^AF$VJ8 -UL]QVFF\CX$:CX%%]JP09CJR>B9+:&X]U0'G->Q9JD:
PKI35S'68U&B>*%G4K-3$LY\#OJ5R^'U$H?:D5$-/^O6RW>#KI)HHK]P-O_4D6\4<
P&?[=>U<A.A"P4XV@TL?1P, I.TR" :EI?429S^%S'3;A,_(^A0\PL$: L+_U."HU
POYFS%N5V;QA#PQ:= !<8'1B>R3=I07BK:]U+Z\=^,Q>="Z6:, A;!_0N.=L%8ST[
P/.Q80;Z,-R^OCV$?2]B:[L)XF+\J./M;#P8'^M#UF10=U9W\7Z)NIJ@8X4_/24I(
P.6*JT4/$INZ8K#KL?+1J$"Q=7PUB*WKB[M<$^7F;R/0=-G<AZN[?>:$+IQZ@V)4W
P10&8[2'#9\>00C.5<FZ_^(**RX8<QCDW?!=961#->G<UN_%7;!(DTYNA'7PAM4Z]
P\!;4C%&)>Q""42N9JIYZO6U/$-,/2Z*J2OU]:Z$,-NH>58XQ.E!GI.SE;A?04?OG
PT=3<! FLDM+\]5R4QR;L8#Y+28%'FBH6AWQV_RDM^&U?^>W_^OP-SYKVQ(D4O=L,
P;??@V2[R+QO8EDGT&VGH(I"/O!JMQ\6G T]5H+-JIT<6/1-DY*\MG'J/I%6);?#3
PA@T%X#G:Q?9:BMIY0 YF,M_T%KLG%P6R"6)]Z^L,D9*X75U_&8NJF3#WI9-0!V-"
PCO4K^PNH^3EFD?L-N#N Z#M,>KS=Z-OEYGANX#\HLUFT1>^OY329EKLU"4O;LICQ
PZ;>=^5K 15VQ>H(T2^UJ.5*FDE1A) #9ZB+E22>T3D76?\V4;>6N6]9DP1$EJI<U
P(]YA+3T:MZ."-<'[4.**AGJ5$-$> ?> GRJ;CFL7WBOI[Y;1G#7A,H/('+^#ZP*>
P^'E@)BLW'N_CYAB2<%%+0Q'P8][&+O^P7U5??&D8ZD7(%9*V[@.DFAS"<#N 7GHI
P^NDQO8-:H)L%U1+[N6UVF@"D3UA :ACY_'(DZ9JR<<U@'; AHT,.&4@8S"ZD#Y84
P9$YPBS9_4?^6POY"#FX2@_U<W&"WN$G:!_XJ="D\.&=7-5/,^/PN8!Y<LU*X9:1 
PVLRO36Q3R2&8>!/1?8&+^\EWCMUE8*XX!H=!Q8/7VQ [,EAMZN/I]NC<5?$^QCB[
P<5'R3,LKXKDCWNQ-4WQ_VDQ$OA1X/4=*::2K#D]BY,J<0FQU/%DPA4D+(75EYZ[0
PH!F",-?>9+LDO6@O7-8L5S-"^&*\<LPC,IHUB7A"\&NTE#$.O'> 4X#(Z8)/%B'P
P)LR1>" >8CV^"7D& 7FTV>3X$<(%895>]S3YOZSB+^/5+M]2>WF\U261IKXMWH+8
P-OK?OUD?AS3N3])<BB?N%2G!_"<(MI[461ERI38BL%'S38PDE:S1F9F5AE/N!Y6^
P(T"4.\J:YEX53V4(1];2-+>\#$DX:?S$I+?-WWMK,!C52S6Q@JKR=9O"]RJ9/&R^
PC9WX6E"-;5T1-([,K%@$XE[WH?-?:8*9Z &/*CVR6H@D(8J/C_F0/M=[' @U9E5A
PFN4."$5&N2)4U'"$9[DFU=Y6$?P:P2'Z9_<%/7J1-QSB82.I"0Z5_K5VK*IO1*EW
PZ?$1!7:,D]GC-SJ%+BC9F\2_3A5V\=!X,_<^O/'S_68)AZ)$G+07I-\_66&G$R-%
P%IJF]".]&./>K;"XUUG9-M8$W4"I59?(@%-LS.IS)>#<8( ;[A(>_/K^6S<>?T@Q
P&]&E(N>:Y7U;/%[Y3B!YM6_N@_P.VF/H?A>I/\#E5@JH]Q\L0.Y03+%"W>1Y.]$S
P",JLW(_+S^J1NTK)W%UGW#_DO#O"'[D:'87=JO<E?S#V1@J2>GMU*(RREDKQ^O*+
P+O V\>.G_"9CV:5#6=5<RFVAC5[Y7<9+-T4PY-@LO]3&-'.[-:;*W(RWW!]2?5C:
P(B/"U5"FHW1 G2'[)7Y=]R^?>7=\]C.:"CEA+&FJKH+7Q!K7PB.5OHWQ>I!&3QI"
P.+AN(5M 91VW.&>N?P(PN QX/0\2<;(!0= E&1MVS[*#RP_'_BYI<^RF&@IL(O+\
PX1S_+3=[!DPA0)&NV^RZL(_L:(I7E>C+OJ(6G.DJIJ4KC34S7>,:0)P:;D"2AAT_
PFJ14T($AMCQ]=)KZ;L)/$S^]X5$-']D.[80OUMGO9M^?QI?/3?FWUFX.8E3X1^51
P>R X$JWX<[SQPSPECW F^^OOM>#4F4Z&(&HC-K.=<O=V;87M-O=U[!DED<:I!;Z>
P3$O[T.&<K^-L(DNI*B5O%EZ,766<"@'($+O,HX!O"!OJRZ$^DX]Y/ I(8E??:GWO
PAPI!YM^J<JG/^MLCDYGB*< DYG&1=GTCAA$[?WELV':[-%5V$9D@.W,+4.XLK,.:
P87.FJK(;%XSH86]F&:DLX]1'.;+:T..5J&I_B-:H?V 39*X3[UG*5G?=6G'\U.<Z
P5=IY3-VM0LI8NAK2H0C0:]P_%?9I6=L+!6T_/1Y%]/U+/X$/)VXUO#^- @6A1-R\
P=74$S,I,?!\(&])@.BC]5(X%AO3;+T<;LD8$272K%2Z 4[NG),))9QC2>N*C,W)/
PG]OTQV-&?'$\.'VJX=X'S?9R &'-$VE2'2,LZ,#EEM[FI?I'.-=[1&.X ^&@WP+"
P ZHO>L^28CZAVV&[<A3<B]N"?B'F_3IGS"M!JJ&*4_?ED;/DE\=B;W965;C)2_'U
P)5S B_G1&3\I->Y#VHU."!]R1WV'_<%O,:% ]*U7YS% Z"-$T?QWRD)8* CXO6G+
PK;A;T3#O<#-V#A#()IW+RM&,8U13*=Z^+F3@FN^8_F0MPA%/<,=[4!%.Q!)F\T6O
P(77,H;%GR$+:E<9#/W$;_164N# W%V9D0^;VAU/P2#C'.D0+Y"8F\1)FCX/*$*6;
P<]P#'7U]B-<OF==K5,\J:BO=Y$.:,T'K'L#Q/F0SMT5 **J6AA<#>5RW_"LM+\8M
PFZJ[V[>A7JW'3B5-.S.0:';(LO^4-4X4=5Y/3_D_P1GU&!L3(.GLF=YYZ69PTG'$
P@Q%2P&F]Z:R>I6[*$+D"5_5BVK%*X$8A>@7_W/"6$1S*]#P=>3L%+I6#Z(8A?>EZ
PSG)5+ZGE=ZAYV7G'&HPY$L^LX&5JS.17':2%:4F^"'>O,7E5\9?W9$_B-V  522E
PKWL5)_<^Z?.FN\D>/?E#F$[*8JZ$B*V3TZV"ZTAD[$0((*U&0AMU8RS9)/ $;'5(
PFKG[&!J0X8O9YB3[9OFIL/-LZ/4I,GJ-)FK\>"K[P PBQU[+2  .)0_27.2P]E-T
PD@.T^51>>++4,P:0(67Z<M^A3$)TAAY\UZS=1."-H RBYCBX7BYNL[6!ZF]FR=;)
P+D+ AHKT&?LX S4UK9?)=2VP4[G;?3)&?G377!9.[1,_)ZK#L@P3"G\*V&#S#)N 
P9$BO/N9%Y6MJ!$L?3]_'FY[CIU]F:YF9RK>;[,5D4X4*L(*=$U#<CW8H]Z^8"O<.
P8-R*&VV( %&I!P<\C@KJ(!&+CM&BX@5FJS=(.24V9P+9DVA(%K2LU#&.KD7//S+.
P4Z[<!0&R>OF!<]H]B("#&P*C%F_CX%GM?)+* .7+@NRJ+\S$E%2IMB;E<0*V&66G
PC8V(3L*V>4 "*6;$/+9T'JI:Q<>]XTM@[DZUYAY#E;IVJT0,E3(2:5C*PN13D)@"
P/48&^>3Z&<-4$U3]X:L9RB<%'AP>PE.T#Z7=!<,A*N+89]"*;7,R&J.D6VU8[%5H
PZ\%CN-8T3 ZP:I8;>LQ(,@*>1%BA)AF\V!,/THXH"I;N\&YRRM=Q#$->0KH204;+
P!W%7(#;I!O'*O :8Y.FJF@87:T#7(5]&V,*B9 Q>+/K;"^(J&$F>IV"E&:-<R@TG
P2."TI0I9@>'BM'X? 0HLQ$=2;!L%R>X73/\7ND9RXW/KQ![.:_QYG=&V0+R-+!73
P[T6&"IEO?(%51TQRK<XXA&*.:F($7HC1(%7+*IYFW[/'SN.F#M61-&=:9',WUAGP
PL^M^H]Z-*,\Z&,-^Y2.B#+QL5[TE9]!/^L>-+[6R/Z@XH*#K<QS"T]0CB)^M[8W3
P1V#4'>7?_6Y,J[XE<JIT-?4&(UJWX/9)$'P^&*]Y@BRKK+]!]XES(->%Z9WAZ>%'
P VNB^?R:7UN]%: AZWPW?#)N/$=0T4T1MJ[6.6LR8>%!DOJ9<FV"OOW+-^6!6U\$
P,+#,.<STP9M1[\5TY@:'.!7OVNK1/_1:GM1__%T>=C%/U?:_1I=>>O6@(]_<*;B<
P;@_$5I"_S%;G3W3ZLZ!RI"J+8ZZP&')[ V;M@Q2("'6:_=9^YM=.!J/JU_\QL*<5
P,Y]7%O-_H2'*U@,3)^7V!E71@O8.MG6/.SAJWP37,X=0"&!'\E*362VO]#RXZ8/P
P,C"5.S/"X;0@W[+8YPIUL)Y()A2=F-3"R>1%D-3JVO- =VXF_;+7TG#'N<!XZ?<)
PU>O3/=71L@>W05_<&<VQ=-#K<:*Y% &^N6[D!XT!TN2<3EN:E[BAL%OI#U9%(G+W
P.)V=_$J# /81N":-C%BV)?&\W:S[ )6T;_%Q^R03YW5 3;> KQD_6$-D3VS(=:<S
P+XER*ZCUTG:""=#3[VQ/"D/EA<O<))26^N#A&7S;698Q:[/GC1-@Z<^(N(S5*H67
P>7/!$WLPB\S4(;QHHK=+20VPR%$!KLS!//OKCA37L8W@XT@^1^PU6=.3D4@W(-;F
P#(M6^[TA*"Z%]!S$CRT3U459$Q"KTS/*;,[N[JLKYO0S>@9,5\$V@7$V6<2E32X\
PW-O>U704QV=5QK.5WQB\;YAO+ I:J&3^J/@ZT]#:H?A\8E]*LCNMZE*:Q\T=\O>G
P!+C4A;A;CK"-)3O_KJV#>$IFP8P($Y>_"^)E&$)/-(!@!,.*]6SHK0ZNJVR82LYE
P. C8V.$.0,P)MMP1*.%B%<$!S0T[A[S"^(H1_80"("PQ!;2Z)\(R"T:UE=O\@M5H
P5G[BL*+VI6CLH^F;%%5JM6'IEM]"Q9QG4__.IW&=RO#SG_4EWR:@6DZUCVU?,QT+
P:)(1D@,/69VD57QGTI?B X[YI^)' Q0V.L+:EHQ @?LFSB_CF=,T^>@<-%8Y1AZT
P4>3U]B#-S$WZWS8]ET& ^ CV^*U@1B3IQN^ ZT+>1OV1?81E$"TX/O):>:VT4-<9
PO]FF@1%0.V^^P9I,>II&4_91 1;OD"IR 6<_I $NX\'7Q_M@:A\)9,9S+K6-^T[B
PP^9BGBI$#3LO(I%%Q9G>U&@ G2U$:)_IHTV,*]Y,=3'0##LA%Y5=)1-WG&IC_MX&
P)*E@1S&&N++!HB@KR;UT\7B?-7=4L$VEYF,'VLX%)R?A-Z."FXI#?=3Y%*F0[XTD
P?!VD2]1:<&!ZY(YP['A,0_A3+J61/J/=IS-BO\"T8^040X0"J]CC6D 8@(R5LN D
P1U\7^9*Q<B--)44J[U$:$J,7&@;%I^X"L]!0!%WR4DI]'M8\QS!.54-* [<1N]/4
P"?[,:R#WOGW_/3Y_@B]L+Y1J)0\#K5<\32K?>>*\1@1J6F]]H^QX+]BFDJG)3;%.
PVE"--CSF<XX(*SW?7 4$<I'U&W1_Z%[=[W?![:8G?(%V553RG2U?_[@U@-4!]';D
PBU(SR0[E\4%1G+>L&>%=Q"IA!@I[G&[A3!Z*:<3\>:LL7OSP;RD8O9H3Q)1<_,<,
P^BL==RH(\D$I/:=K*.?9E])8'E"P!VI"L4.6$D4J.T<X@N'2&]Q"V=+Z&SE,<Q,W
PED:^OY5=Y]69IK(AU1M<DR[<PFT;A\\TOR=[ 4/LSXBU7E+L% O%R"6,V!("&S./
P?ESES+LB83:C)5<8;N5_=_':.>KQE)_::5@H\)S$<W=I :35D%%M9'2'XX;1?*"6
P(>UO<SU]]B$'LN@%^0[):C"LC;^][,%NIJHX_N=X3/8V,CUB, /:1:1;R459,6HL
PF^>!,F9>_OZ7[Z>2PU',4P15(/,?8!^55_%# [76[TX<S08R@KDRZ_K5"5"DX*X7
P>C'J8N(,_GJ552]A25K*,%UCG^:C&7=XK/Z/5/K(?:_N7L",\NU, .HV<@$9=?WN
PT0!''Q19LQVCL\ZG\UJ6(]4"APFJ>U?CD_N&(M[R: =OB58![MR,O*@VBLLJ.)'&
PE5#E'G8CZX-T'L%E)@/QQB1XJKAQ'Z0B$M74)Q*#SRF,6_2!'^J5%6?M,-6S@D'=
P@D?] Y&NY"K 7Q*APNGCKXJ)(U>Y>-)7XT7^4@O;H:RM7-[PQ..K#[!D<<D\:J\ 
PL LNNNS?F2'6-II@S/*&O<<Y[YT^@V-IVZ'7\(MT$^*64H1Y>QE&3>0QCK4/8B;E
P!37N60OS&J<G>+*PZZ?X$M&R+:6J.P"$Y(4@G;>C4W;[A.@L% ]-- ;Z6N_2Y9^=
PY.FG;*X>;&FOIN.K :5^AN_G'.R ;UNP(],PDC>SJRGT/\5/+RP,24&&:)<@W9EA
P8Z6/V[]%E-@-$N=5LFG&R)R#<&+8IG/*0ER'\U.JKTJQP9QIM<^R>^0_M^*SE!)]
P@9#X!,Y(D>0U[*]4M[6U_2VT7YP"NWZ)G1:HC6@80N$TM?JY&6<P^93&?E^!=!H$
P8U,QR+@-'.A]7&( &7FC_&OVV$/&=)#(' _W LW>?!O:JFOWN^$1F*)9TSACOB"H
PO!U_A>QO+RO:E'!OB/FZA+NCE\G+Y40P]?$J/5*'2S/_,0SZ"IV\;[!!4^Z6D_RD
P4GE;]I+OPJJEJ@\J\'+VTZ$]BQB"4MO+S5P.OB.N2=ZM-UE:1C05V/''FL:=@78)
P*IXX"WH?W]'=]U(>I1@F$EKT'Y45#H,6G):D\C7U'3+/[("V-+>?7=._SP7-F,<.
P'?@3B'3O42:BD%PX#:7=!B%&,-TM;.3CO#6_<BEMQ#.CT'P3:C[SVF%L^U&QZ3F1
PZ/5*%OY#U;$;/&%3VOUYI$ZMH1";&?)?L3.8EF8IF>/L$'R_HY?!]S24;2Y%VCOR
PW=^W#00M]58:X>:;Q9_4AF<<ES=K?3-L?V2W+KB3+75^:HQ9I$^O6K9K%^/"C:0W
P4)2HS=8>)#!M@%R<FJ]BW2WX/*LQJV[<Z)E<91FRZ4XEVE=7[25Z$ .G/HE=C[S@
PV(WVI-E9,+\PE^08TCJF1I--@&G;OU[UR5AC&;X[J)6$OP?1(+ST)@W*0WXKVKI]
PW\&)!0,J4V:S.;K\#FXATF.B6H@$?^MB,N,>N%>L&1HTFCB6;5UC"OP/"M$,"37R
P =V$JDEP5(_7%V5Z\PSV35P9>?OCOEN!S3OCR%DL309)Y'?93SKJ@W1\7K3CC+Z&
P0/L!/>P6J4G[2>2\A+C!2+;QS]1*;C>H__I@07 \FGSE4C@)Z#)K\N"I,4Y#NT -
PJQP0I;%7/5W Q@X&ZFZ0EVS=PHWE3\$M/D<X(%AOHLQ1)O"<U&^9ICEF6!&I\=(>
P4K;6(N,>]$_@GWR^;*G?Z'7S<2UD5FU...\E%-+XO1,N]/E=L?E)WO(SV4+'9N8?
PM.(NQ+WX=YW7;$D9K"F\A73"YV:T6.+9QGM266&(<K/Y*44ADRV&>%KGZM-F]E_:
P]^#_32.'!E* P-=12CI&S4?R,7_@C#&SHV#GDH;'DS$9#!"Z0_C-0AS@_U5)38S4
PF=?M:!T1$!M3-RV\)DYU/1]T&;D*]KG#P[UV:"<"!]X 2RA+%*)VC[I^1V!Q.D#)
P^&"-RPDW\83>[S8/?:_DFT&??"JN.*3F4JS]FRN@4]O^J^^LYVA^\[<6N%LX3%MP
P"X62^GQT7R"*!P/KUI(:G$YCC^I#M6815\FO:6J2)ZB;05&7!2DQLQ0AMX86XMDF
PH<:I1A/H!;^DQ\G1PCVW#"!G5@?M?+=1^^/GDDQN1%QLBE19D26;G[VF4,5\M1'W
PO\"#6EFT<T%\P,'-D/I+Y#25,*O\CW L)@U$HQP1$ E,?AO.CJ1$6.&895Z/X=\$
PLCD -3Q4H![?/$FK/3ICHODN+?%7J"AZ?,Z"9UOK;S3?A'$D?3Y^M9*-1=HK1RV?
P11URG?,)]_]$(S7E,3=ZE+Y@(59T3I\W4G (%WRX)7CBDOJ"XA>C1<_T.);!C6%X
P*AM-M8>!S#J\D8J^W/E%,HS):M8)VN%>UOB\@4GRD,/=C+*MY48KO HLI%KYUA;%
P>!E\\H+OF<F<[:24>'A,"J194BBW]24>QYQ8%G>.O",F\NGMY??E/V<]\ZC0R*+4
P)&#2'O<3.Y6XX".386A61*$,K)"R%:",3Z9F9JV$GGE(\AUJ_HR@1%<=>P3REN\K
P?-RF"D52C(UXTWQ2G%S?>UREFGR3R8<#5'M4 L81^N$I&3!&['*E5\FCZA;+0S9Z
PU;H;R)B6_3TGZ<XG9<5C<9*L/WLFX>76%K""9.7MJ<,CS:98T6.1!1P<,5&I:_ID
P."X0CT0VS*NBPFE.M_R<W%:WAB<V5I9@A2Q)@;S2#P)'Q_QVES&40J8YKQ^,[,@_
PPW/U:?DCN+!][?$+-J!BIG)?$@0#ZJMG[(685)L?A<VRT0Q<%">L4KVT=N6#P\7Q
PIRG 3\UFL9N<-I7+TEU9H/SR:A"Q1NOXOU<=6;9MAX8/HW_WO^ZIVED'W6C>6_Y<
PS)K!S^!-N=WW#XXHV(FTY4XLDGDN"K&JAV3&[-07P-Z,AEQ+NS4&OG-W7(N1P'Z0
P7>E3.2$YN\J7S+P-.HB"H]%"B7VMQ::ZV$JOK*_=F];":S:NLTGV7YD$#O[?#"HT
PAYVW& ]DMF2MCTZ,<,"8HDL_6/][Z(=W?TY_<'M:#0HYV@PMG19Q9LWC0751NI-^
P5C8)?B8\B^^YME5M(2$M86 %_ E^-1-QU-@AJ5YKDL$NI/O3?L^-9F)\"PB%N L$
PQH_BH Y#U0ME4JK+GL B 1HH%[U3$_[=4@\!H.?003<F=^,3!# C8XKFH+2=UPA 
P$0,AA!'6B%39#4L #L']$Z46WZ\[)A"[,>9;H5V0M$@<XQT%X$VGY; %MWL%EK[<
P@[<ZA8$Z(-6I8DQLR5E5,[5T[RH3(&[X)V:] ")K+^=XG4!7S4T*8IY+AL/K@S&?
PXBFKT2CX8/)JJ7,1\U&#0^%?(DY2Y/_BU!-+XR!DP8Y TOQA-S^8;KN@*\@=!(I*
P&]-#E"2X(V3,>A RM!YC>*=P*3TM8N?>"H ZU!Y>-)",A[JVO%_;C.(^=54-L)GJ
P\SL3[4M7[AI 0%I0TMX=YEWTTT*HS&!%7\['7=D ,[^73=Q/:.ZR8K?I=O.0RJO1
PZE;W]JH(W3RE2/:!<OKSR(YYZ=$ 'MFQHGU(:=$C#?F$L%''Y=_],[:K_KH1[2P=
PT-\O&;)8M[D--#S YDS&6*XG)JB/!PW/B)N:*YNX=TE%BD=^;)G6[WVJP5H@7K#A
PBF1)3,LXD&),A3KLVA6/PW2)M>G"3XKU*=#E\?M)=3G%:R0NV:W6=+*W6=WPB,E4
P]U+>FA#Q7?V,96*NST83A8-NXJ$N"FF%$B_.-2$>'B//_]F];I-[G 3&?''&L='Y
PMP^))MVW[8GLON-27JHW4OM E>;;6)P(0'@W%57<!&L+'8)$XEU$H%5\\N(?1[1>
PTB;6%.X(*"R^-O:_S&F,UVH=1T'8_RRQ',]R3[O:-#D'O-7I=PXM*-[[E(LRP/<:
P%NN'8<AU_O:6[Z\'%['%M'9D*TM;.BM'8EE8Q-\:IMNR/3;>@6ACTWY['1(42:_@
P>W$AS=Q@#'L+0[$,;D]IQ!9Y6[,DS<J,0#5^9Z%/+8_]A]V/>PHEM32?(W>DZOWR
P%NS=E:GZ9,T3PF>7%YP%=K?<+EK6H&%#6$1_%G/S4+E9N6:]T(8E,_6D?8/V_.,Y
P&7"2I5]4&W0+E2\QRGSTNE<\(S'!KRK?[Q>#-J  (6F!O!V9CB>)_V.H:%&9ZY]%
P+DRYRLE/<E7/38/YF(D8[#'-E=&3^=2GG.08.&D&M_>'<"E?L<-1IG:4>>CB(VP+
P_I?='>[<#7[:8'Q<D'ZKCL]M,^[U%33XRD4<Y[@K &'?4+9EI--'SY=I,*@G&@1,
PYFB:-5*JTUV__P\M1XAS%X@\_E]A!.2"96)&ZO.H/8GJ^#'%T/&=H33D)LM3?<_2
P\YHRQ0G10*'RWKS6E 9H$:>=PT^:\_LS8 K&RBD,)2P37,$)5)R@V5*PX,P*@$)1
P5XVH8-O8LG*W/<;EN.@@7M@71CX-DYPR84M5YE$ 0Z.<V JI]:&[=L(RG,((Z%/C
P&SX5X"]<4UXJR#4R]RW+/,A">/_07O'V+X,UZ(^"8"4#P$-;KLFYI\T%\P,!8BG2
PC2_'\B-*@;#@HQ-]7QX>]2C4K.5IKU%$AJ07 X\#TUUZR'YD/$+04"&2HC2##85=
P=@N6KCC90Y?-KD-\MD KQOA6TO)&TG#"\CR%9[V2E)=16O0W ]U1*]BV.4)8LA2@
PXR/!5_4<?QR%MSI3,PML!RG>V^7U%_PXR-:<;<CWG&P'4]4CAVP2C>@!_C=J68E,
PXHE^>RI/#>RWV78;6X>_1;[:?\ZNK4<P4*M_S.6YAF#CV65&:4EQ"M93'7"F<3$9
P!PLG62%.[NFOA5<62O$<3;I."Z<A,&VPV3MCB]C/**6R@!R'R;/_#K[\G(\'L +L
P8+TDFV*[OL-Y6?V=C;" C J"0_G!H7JNADK 5QD-%YE&=3I@6O%8-CE6=3O;5V' 
PIXC8FVY/(^ZYE!.7KJXO>B5&="9C7R&H3<X(L%CR!\XV#(2[,!JS&$/2_SA?\"&R
PW;T\YAG*]+H'>&HS0=HL%B16\$JV1P_M2^5#<(+*H+P@5N90Y*?ZON!*6SR^UBPE
P/>S0/0Y?,.=\*#/GIF*'Y&M:4Q:YJXZ+:X"C&IC$_"["'F\P"-[V&!!A0W[L<;_Z
PW:1@DC="#OU,L=P U0V[S08U3JPC9?#?#>"B4#"KI2VLI^,:O-TPU$+\4VMY'_FN
PEW2D=2!W(NY\R7M1,?,+)DH,@]3%B:0AZQF5 16IGQNL_3//EQ]S>1GFYH+@=NFM
PSD?\6F%6SW4J3N*,GIHE:A9B0F;>G"L:RWPUG.&*5[KZ^508S%81-'_8W(1W.%M(
PZY#0:$JXM$';ZU!7R33EROB)A#UWP.!1X*<OM>7EP6)OGKT-)$D2X4Y\?ZDSX,5U
PVE;L/]05;\#2</^\IO1G**&*%Y5C3 59(_FU+OS1]D7ZY?OT0U2!8@G,[I+DB:83
P0[H(XX>B)PI%4^!_6?:"">UT[1Y[B8+?+N;'>WT&FT^N.E@$#!-=U?T_'?KG<KN,
P'LYH0N]?CG7._@ QV(,,!*]RW/M9N<\L"LTWJ%E;=1X2TJ&EUS;CXN9UQG<M.'07
P,J#1&A9AS4^3]K'+]!,1N/N@UMH" J,'Z_TO48D'O3FE8*^8L/1!M,JPAQ&LZ+Q6
P4%#MT/C]D!7,^INFZG0((?&L+:L$-X.8UE2>.A:-P,@]0?^_].VJP%2D>I""#*_5
P,A "P()ENW4&PEQW;#MC8GG&V+%+TKCN1BR*0)K.1!7#4&\[F\-F'BYKX?M=+OJD
P<E(?X)OAE<=WR]MG 83?!1[W3[2R',B,=W3.==S'^)7'U8A4YX@&+>* 7L]B+S+)
PFC&38#B6@KJ>M,--$+7J@18U(,\["/O*US#!O.8'>H.[U/^[088)2D7&6><>[]K>
P[C5>/;TZ"^9;KE(OBF @T\@T$HM0MR<BTOMI7(,M83]O31HC+1#*/BZ2F\WGW@UK
PB10D=DV$THND?[]="?RX/N=N(CRBVS182V3%H:@FFL%0[#9.:^8GU#@<(J"GYIO;
PT!WN^MV@'0>('BA+(,CPD]=9#C P[/>HXN ? W .5:-:#]4CB)76D],G2?TOH;[;
PSDO+\&@CVIB.P6NE-[T$ .DY*F*%,9^+ATT=4.'XTW0X;V0C0J,XDNY+Y/XH[=F=
P"1Y V5^FC-3(2*L&4"]6M6UA]ZI&76-_'K7C!61)M^KOS7X*05:P QS_5]/9U4@J
P)2GO13S!.NG13E7"#1/34MD.5MI ?Q87%F&!P\X2;:3NGX7[#MGD.F7<(.9*M9&;
P6&X-\I"<^@FH%&U/A>F>I'$JA6H+W(;7 DNFP7>,T^(&6G0;0P=.Z7[5?EP11Z'N
P"R;A,:52ML XRX_TI&YLMK:P"P4QMGA-4&",(YU[#,MO$3_X/FJTO_4*CB!^?=1#
PN> TG"D^"UAXD.$U<4/[->7/%67=V9\P[K]EIFT7\M28*1'VK2]5TE5B@YRA9 N/
POT(P5PU(<2&D^(#L1;)Z=7_*>MXCEQDN$IYXL7>LGJPJ=_ITRR][9SHW+=L<^9ZP
PB;@T6FSCV12/O@+VK/H2H=KP>6%*O5^(T'[IJZ0(9]PGI1'_4R&J46@5$3#@>/P 
P]<U 5"'"M>3\H%4&0S*6HH1PR)?Q:58C;:HJ9G\-(/TS, YX>_EU:E,:TU1]F6@V
PNA!I!*4E]B(4%E W;L?C[[#X42O'B>K AK;PJ8ZR/^S]4LCLR;RL-WHE; @YA1*0
PKER SP>YTHWDOR)[N+9;)*G++.,:R\L1JJ6;6W;^V*)V9!<XF; X3@N4<0[7/I?%
P<D0.Q34^QBK*^N?60N!^.546F!^5,*XNVR*K&+F5E-[%<+L1M:XB<FK=#A[]H!1?
P5K5@,R^BKO8FB5VRE;PJC$J*-THL8AC*O-,C2X'OZ'J.^BBN#9^T'V+O:DZ#31,4
P CO_!#_S8;(53*2GFD@__>A8V[OMKN@_L)3AN;>Q8\/E,82+;($AU?%!J]&:EE>T
P\9W5Y"Q$7;_EFM:D1<>!\<YU8 XXKT?)8CI-)"S/=\(F8*M>BAR>) 6BX/O7WSS?
P\(DD"@>0#[J.VX$NT<':-E3':3?-7A9]&I]S6AECA\5%UA0K]C@K5+FI60$ACJ27
P"'&1HK#9L,BY]U?GK_W >;GED^;%B$_R6&R$[_LF*JJB%*(OP?3,'S,3V=Q.BWC\
P6@VV2Z<!G@A,IR!6M "L7M?CQ)!1?3@+V\E$W  6IJJJ<I*GX_HPUC_!?:UX1=:E
P6U P'@TAH@2%@#^*-,_P@DU)5"B48!MX?"UR/ZR\?U]47(RNBGU#)UBUU^C/3_Z:
P"K6"Z?LKL<X3?;.KT@T",6A)JA2'N2O#KDK8F&J<TF:2D\W<R!D]:1C%]FO9^'F2
PDP^B;\072&;<N:S1,[4?A%#J3S[A<OF4VK9;'I0"32*K#)+SC%"YOI48&9@9VM)H
P1#<N#1H\UC#ZK;D<3_82I#B ZC7FL 7G8";93-!Q1(O18;6VT%*PM+%!)H(HL"1^
PUBT -/<QO9&7CCQ@>$Z$(L0*0P3*+UJ#'N+JU26 $@=;2C;@T9F;=5,4?JB,.Q/'
P1J\[.&)K6TH+W]&W>[^?)@YLR&O:&M E!2(O4G<?RB>[+<\41^7_W4XK<#"3E(W+
PSQ#3^E&N%Q S$_ *DTD3LP *.'(D "TGR0?/),)@)*^)/($QD05T>N2G=@N'F8?>
P:08.2 [@Z_2B?VP9_T@-S5 A:Y)2/_\B_S+L/]A2,6 .6U3B%D0\=X4$*)#YO-KF
P1-*\ G5^<F,$Z/)E ;$73#*[:HY6';?<SC,SB^D:NS2,&Y;-(\EU-S$YJ.>Z:(1)
PBQS.R1T3E8!Y^JR<);\#XC.4879^Y*Q>;:EI_BSSF>'%$7UQ SFI82B2.?-N<:KW
P-*;]8^5M"VEG XZ-#@"_D%(-^U,P 9XLA^8H?;LOVYP+-O.SR?6N64H1[(P1FD<=
P!UT44*BXC-PFY:I!-%FN]2*$XD0RB+-/4B=T3 GV:K=@*ITXL&[0[+&J N*/5]\B
PXG,289Y@Z_[WI,VV"!,GC":*\91L=)2)D6Y1!@EG\'LPP7B-L,&0IE&DQ-99V!NL
PW]?<J,,3)*-);;G#A6F2]EPA)X.A2'G=(^C]^6[47+(O%,>@L!P4X.867-37PDMY
PW&-BZL FLBBJ6Z^_MW^IT9 B6H\*>3(2TY-?T9;UILDT\L$8E#GT!7#(F?=!:0!"
P)R4K5/2Q;@@T*H^R#1()%7GIZ_%=5FM(,$($[3=+*E9X;#D$'^@]6RM%EB8RUC0D
P+$S@U@BS+M./&]8<58XA>" V?TIHBK\[16<HZ0N360T,40'DH1VN=3HF!3]@XSMB
P!7P).<@2I#:/ [300ZF>)3\?+8:X:5 QO$=;)FVH.P]8=*%9VSOHT2@7D3F3:-_Z
PGX0,'2+0T%&1B&O8#5#.Q.%6?/I,_[ZD.( '\9I0X$GUKJ!+O<"F41FS&H)?G> M
P0.?;\C'I0ZCE04U^&@X@6]9,K74$,$1PPVD>2R9.D>^109O7D.:R=B,V,HG\O?Y^
PSZ9+[<K2)IAT@_2?DJEP8K=ZOA12"[\1R$B6MG'@5M0"WRR6I-N'4/ XP]2CIK8J
P@%LK@WL0-/GT?)]4-A.4AX1/F7/A\-4W*R;%RL0TR<I2B.[^,B3N )<%TB>0BD0,
P":;;(:L*(E%1I>*]Z'@0C@595.R)GKY)5=->5GXJ$SP-W8,VL[AK_OSO8E*- E7;
P0K.V!<8X<B@*KA#A0+K"&:J$8I41;!\RQQSYT%OP#-A*M(E<RR#U&P'O^?!R*/#2
PW(EL7)H+.PGWI\0X^RM:WP:<9A?*NE^<W#R3#X\?@+NM'6?74('FW.R!9Q=;H?QB
P;CKHAD+.L-.C.XO%>CQ&<'-N;QIXT LX]6\]II/>)EBMK3A+ADA/*_X5S$W9 NZI
PC^&N%HMR:#B-MLH'Z:" ?,;X,G@$%[8;G[%Q.DE; &=/^R&BZCT8*T'0K(W@0RVR
P2O% 'R+G%D YTAI14-CM2F4MAXJ55#-E4+>#NX,=)G;92DG?4Y75SUM_2D."0#(@
PU)OU'X9+\PIQCX8?:*:4JXVYTJGFO-#B_^%IT9ILM :8[^LB<^45<1YTCAX@%3K3
P+,%MJ6J8?J@H<T[V$B-@S^*PJMB$@:25/?+6[D=YV; "_(B:,V0P>Q#8LJ[@7=!<
PA]>A=11#I*_$,A*G+JD='CKA=1Z"$K$_N38G3+"D1W[]GAN\H8[V9Z83JM8J&21>
PJY]80:Z6SL.?K@F1)PE]3#A<%W[8L#4[&<)J$'SAF- S'$[&Q0'$ W)P!A8XKRU 
P2G!]]-=BL7.>PS4NHFI\I0C)P:"Z1F&Y(''7[7^@@%ZMI<O+%PZUA>DZR*<MBD)A
PP;JRI+\P*+8X^^)8!JW8NWKO8W4=;YIN6H5L=$RLO-S9!@@9\!/Y#C3S4VP<*)_]
P_1F-?!KD6:IWN(*FME9PTB5PB$BEMQX 9HZO#&9TK("CKJ%;9[.*1R9@?G$?J]XH
P)*2< ?L #9J@L:TTYS%F&NM,!>G+X<_,LY=Y+@2R:C>$E1%SDZ86E)<GDG!=7 9W
P] DY_SS;56G@YSKOF))J6H'W_YL=.D?BUD#MW@FP\^,XD-G0OO(^JW5-\E!GZ;S[
PYSE*E4L3.#=;[,0?ZK\O<4Z$VE7?D\;*P?K@J3(:;KYA&R5(B2%IH-,!G,P:A74R
P#ZL+D8PV7EF;,*PC-"$"Y&*ZXY.U'97-(-<%IG?WC0EXVY=;<<KSO_-P;D:'KQ%.
PQDMWE%K#_IYED*NVWQXB=6'2D;E5!QE<PUDUY7(6G=0$792I'/\HK$&# =K INGW
PS!4%9.J',I1;=$8RB&D<US==E]ZI116"%@FNH?0?Z1GB:*KZ%!ZY8\&2R ONY!I_
P_*-'*9(JO1]K82OM3,1B*'=(]P&@27@6,6>@W4W0B]^P9#GD)-59):PIU >^>Y(L
P9F@'B#/$>F@$'?]+G,D0)<O&^SGI5"KJ-?]'5+XP.O3GZG-UHEF0_(2[@L)0[&=_
P]KX'SYS>1T>G8>\AG,*",WA3\$G-Q.,O^X$2_N3VV\A V>YPB;6ZR! 7K&UP<'O8
PS7[Y1\](/#?'NKFQ.AIT:U5GA"3Q47(B(&<M7CQO*RQJ-@X*ZD#-Q!T65OJ*Y^UA
PY<**9G0X6:*<(#G2&9<MKL_[;JO3.B:T,_\;JR,9HJ.,PE?;HP*L#/N$R7U$2!/X
P7/%S1>],N;(W=F5[JC?P]ZD'M-+6C8N-#$%@X<TAO$7ZUO4QF8VD)[>H3;GJ.E.$
P_"WF$EX/GL8KE+R<0TB6DTPA]MH-\24GO%<3;OQV]@O2=7P5E%PD Q77,85//IL@
PH('-O&P J$TVB X1,.24S_1,X+U(Q H4Q(QR+.0<0KC9E3A2WD"$XAA9N0805DAE
PT_$/29/[H)><>;_-;8&:O+G1&(:/MCME&K#=]_O?B'SP0:;N_DW#[ Q,,0!8RHP"
P%E#6C;Q#(D85#&W8>-K*WA\<M9%%@"'MEAAVH9=BO8XYR0P?[R.Q*'QJO&3?D$5N
PZR;!^F1_;]Y"UT>+)H"94J:7DNU69NVJBH"BC-W<(47VUOD!QD@NX>TL'@_BL)9I
PY%(+2 J,$62B+]W[A/!%":"9U<&]5Q91U4ZB8&0/6E$XB( !26KI"#XQ-,';_C/[
P-.G86IYR"6+E%S?K=&A<,S?6@7:#&0_C,)(@6$#&Q49#C#IETX(2BT>,-)#VU<A.
PW>2($W#5QX]NT9;?V.%)1)F^8'>NNZ'-*8WDFE'0"$B[G,5:P^7]*UX_04"Z7)H<
P MJ%;PD&KC&>.1QUI?U0^:OR=&J5/"'2'?";7R,=\G,^#/LPMSN')5G5(\\WDRLS
P+FOGQ<=CUEEZ>B'F,F*]HXKD-#\!CD [AZ9Y*&^Y9*=NBC4J13S+!S=&4="BU*D5
P(^OTM;;VCM262HLMB$*J4MAE5-:B&ATB@VO1W$Z8#M1N3YA\K3R*PKJOV6;A4 )X
P_\RYU  ?L[XA.6E$^C[=)Z9V#J6M@>/=B^89+DW0%\B('.8J<-QF-D6OVOO<ZQ /
PU[?&U1:TG*P=,=U:>\98HUC^GSTREDG7Y,GI!A:*;-(.>W@Q#GA"#D7*"L-C#& &
P>=3V6O.18B<<-?!:$5O]&A[YXE_M8'U[1#W.IY2V 7IG0K-\N5V+C0+GM9(=DR+H
PB()9P$Z6Z8IW*Y";JN>[G'^('U;KJ.[I#K1_(\Y,&82D26COR!>V$ZJ&ZUSC[=I;
P;YL0]ZVD,9YC4G/'[$H_2^CHE<!GB2Q7VH^$^TREA, !;JC&?QU43=4-F7IH^*(%
PZJ640K8N"+JU\A7J1MW,G4:S)\YQ5>%W/97]^5$O-%U9,.H6)N'+F'12:#C:8V3;
P;)S '29S('Z(OUK9Q]TNY[9IGB@Z?FH>XZE.Q,I ^/)=[(;9Z"4NA[)TKG$CG$#)
PV6@;'3JH>DD'RGQCY$*MC$R57<KS,@-C2$WL,4Y/7@?>RH*#>&P:%?(YM%P->QI#
PS08^.Z'2^R=UPT7G7M7PWUHN IR8G-ML$<7$O)X2]F T_J-4"'Z8:>6]IV]@Z;90
P[R?B9L3JT4FZID.%U=XA+Y"+5]:Z,LB;V7MT%C'XAK(#*CA%/D/=7MML9(]#+KAX
P_'Y[3'%C-G#QQD6.0%4?1?;KU E&8J^DM?%7ZV5\1%\:9O.ZT\O\)HG/L.;ZY+<(
P7AS0*@M,_3P^V\VC2>,G2T(FFDO_Y"P=IW!%FC&"+:TK.V/;\$GR5P<=]HG)M@"'
P:?2MSQ,K%[])[@^V;VC\UU8H4D7MALI9(VA 2@2>8BL5&D:!01GD['FE@;R";FP$
P[RWBOWA)R!Q86R@M0%X05?AYS&HL6WC7M.E?/C/E-Y;: 3Y&P'RF[&]K[;4I!X8Q
PM=""^_"#\?F%TA6:*=:K_)# _!SC(^"N4<.PNYK7H0TLKAM2WE1SJ&B=6)^'Q':>
PC%R&8QM$#B"7N:-);JNG,.(6^[*FY.;V3M=X&[14,IX3R[[?S8.W 1,W'T^+CAG5
P\XON,*2R>HDH\@.7&8)@<<**?E4ZB@",\?6U07*;RHC?+CMIEH]),Q:D8%%.\M^#
P_U&H &NVKRY60L.)@J\)4HC_%.!\4\;T%#.[MZ#RINN-FNH=Q%R)_J\V](LPL:-Y
PL^?)$#Q7-FQF5.GAEY$-4!"AX $ $\#=+P3-YP0B=T(\;@)Y0DCKA1]J;@>(C+S 
PA/G2)?&Y(H_*C^-SLL7=E53<E"D"J0$>C-UBXF"V=8R!-'0W\J&T YIL5?J,3!]_
P7O%+,;O:,'BGI**<3RSL_+9H'PX.'52 B4(LX?N9#)H3L%208>"$TCVG=R8HO'7$
PS"/-OG,S7S0 ZR$B=UA4I^[0T":>FQ+X9SONI+],:O55&MCTE",U8SSSS"A&_I1>
P,.'/TSI,BS/,?2]2R)5*LRA#BNJG\>CU>>^>:-1PA#:M37"=0P09Y"JRYB[QY3^0
P*U>5\?GERL]_]EL^76H,R0M^Z;@[7)$9Y).[LS-.(TEH2%FI\T4@7\'EO#1,H,[:
P9'72F#O<[1"\4D51?&B%;D^:%0/?6O'<T_*)4*T[$MXR\#"T9-I-ZE=W^(=_OSH+
P(/HNB_>/%/A. L_30$8!TS1LLL8D% T%>@+[CG!%1#A;#IU3=Z8A%%N+'"TX=HP9
PEOYRDP5 7&@@^;MNGF@&&D%/(:&@*2(<D@!NKT+@6Y<[3.1.G5LT'J_BF?Q1J(+=
P99J @C429<=E8]PT<4["Z-V2F /W?(0-\<R2*J68<U)(Q<<%?:PWQA[+D56T$*,9
PA]WH_5+!4PEB2#]^Z?^+[/7#D'(77->'2Y WIBE'X<CX= %Y[K'8;Y.963II3VHX
P2Y]0]BGC*>@#$$_N4?4>HTHZ@:/>..*D/!C>U"*N['UPW!X1OKMX#F7^784F2H46
P@TM$0,ZW+EX)SL0SG'C3<D6R97+@!7U<,&\FETJD41G!L9G:XQA'>*0,Y903"J0;
P[,X)^@"GIECIYRBCA414+K3=.X?'I)8BY)*_D2&0D\LQU]+Y52S-GY<WEDYS7H=>
P,3\4H_I:.7L_*<4X+44*OA9FNWH6UO:T$YN^T#>O_3;&JD@+B-R?-"9JY)Q:_>,Y
PP[KB!UUF)+.QZ60*#9^:1Z+%N%(K!O6+</K79N94ATG,PB;?*D8_[SG$;/A2KVS$
P8L1!%O>$7KEGT#A91JGG)O^Y)$<"JZ/_[DQT1[K9%@F=^?="1UNKO%[<.,H\C+ L
PAI5XGNYVK@P63,_>8U_W*X]I1G'3VT&0G(!N W1O&/PKQ_+5J,;=;4'H7.3"><>$
P>DM(GO/A@ 4C),JJ+BFK$?UAM'1.\VSB:_GLM2/FL:C/F%9Q(?8/ZP%.Y%!9_2;<
P@WZ:<'.HP;/;Z^P#DD -HF0.'@6-JOU*9?O< RA"+:R!MV+54,-XBS5Y\[S#E_8)
PWXLD\-B^!+1^5_/P#XZN4?K\0)32;,#X7H1VRFK.+=)Y&J6UTY.J<VX_VVU^S_8V
P7%:_%.5-=\9F8/:N$ C%,A'A=]Q30\<5#S!.B7'_Z VB)H0/DU: >Y==,DX:F23C
PDG+' IMWI+]GH0:EFD3VD%FX6PVP0:;]!3.4"\TC=7D;ZM5[H)%/Q)71NK L5P>%
P^UAM('5\6DS3'%I-P5-8,_L*2#G?N V3_,.+ON27M"X)PM917"ST#>8!M<=[/OQ4
P@;?(6M4!-[ ;9'$_Y5.,UV>,Y! Y%_@V%>S.!M8[U]D8F8L<UMR5:*@#B11N:_^S
P^5\:IIVJZ&2 >A9Q,75XOT^]KC=14X!+ 4R5[U=4(@I$X4G N )(\?_G:%RQ+ZP8
P(E1 -1ZRD&[!NSNO3K+V)H]*N%16H@51'P1B]?0')K!Z)Y!FI.&T]](V>]AZ"[/@
PW3#WY9B 58UI>HLSRT8,X8."IA2VMVP[+J*]5<PM!AX^HG!P!]\,ZGXL>:&%_K)@
P]'>&("%=";4:-> GVT1O>8%YP50#=9@A_V1;!$40,7+6+4S)E#UYK$!@FI)\.J13
PBK->XP-Y44>UWU!#VS7Q_JU[>"NIR4@>N^$26F$>-W 6YU6:5F)<%OL5ES/(4@H7
P8+#BC:V(V(:B4R4PT1%DD[3RT;QBXKCF.OY@O4_S$JK>Y"[86=L#-FAX$I2M@7CY
P5VBQ3H0%DITH;.4RUKYL775 &^]86HHN52PU/(R8Q@S.T)95#W[2?"S2_?G:*-&.
P?;,1;(6PN96TJ62&#'WT8D;TUUE%U2)_D[.X_Q4&^1&S5$CO>6VR)S!N5@:%&P#3
PY)Z-OUKGDM&AZ;]V8X2^J7 .E1E-0!@$M].UE-OLKQ69@=XH57^6#=Q8)=PE-6V[
PK]1$]"Z6!$Y0DVW'B@(SY=KH5XKJ+#72>8&[]P*,9--!LB6MVS6H&2U(0LW6H,W]
P&S1)1DAF++IZ'5IH)TC'*X@\,3C)I>W0\!6Z\K>)! &APJ@A:_BE%W+W5PQ"D:,C
P[&/RYYM7U_?HPE_!MBEXVBJM.C+".\HNW2K)9?3'V; TH$YR9AH]:B"1EE@,44=9
PAVC;O$'9AXD/V<"+IYO<,48I$P5\0&-D2?'$FGC]TTC=^")*R18YJZ%YP!]>#9!!
PJWZY\8T!KMOWK">W*JI80:8C6RV360HX#2$GZ+Y40"<P< 7197@/Y-N%.:AB<SWU
PX]$8FVX?EZ0D94 :E+*C8J?:A@7AZU;["-@KP!GF_$*02(/._-.P+)J!2*(FC\KN
P(=.@,L^/WF7H?Y<9F.X*"/4@3,(#AB(T:>;.1N9O+U M5#*^)K. &9JQ?VL2 ,B>
PR6\[@]AG[^*C81*M'4OP00^]V2*ALA7CC<R%93;R(2?K</LV".\)77BW^;5IDR=_
PRO'+3J!_2T,1D:^QF8)J1IOMHN-MX\9UHA#&*B]!W8@R1MKKVPG<[Q*JO(+@\11W
PF4<H1%4Z.Q8>AE1P"0OK='XZMET=4P*Z^BS*30Z$=JP5_'A7)<7N0\G,@-$F]'H)
P7%0/G=+JTJ#O<X&:@#1??G4Z#.;B99>"]Q@;8R/4G3E,?#H1YMV^=N/%#5#]HCH#
P5[H3%$_C;;GL$\D#EH5WWJW%AE?-B1Y6F*$P 2@5T@E'O5L0173 [J?-]S\P#3Q@
P$#_SVXXA"WVU(U[8^[A_"('U-?,Z4Q-\\:#I2KM?F$$$B<HY>Z PUB26BJ!.^,_O
PZ]W].C )L6!-(??UG]7Z52Z-E7L</ =M;)$:X(*;8>I3GI;+\67P,J1[5GBB[=9B
P=ETD,H7_'G10?,X09FDE_Q-G%O?RQMQ=X+L.]Z&+0_H.V4;2=[TRA/O2>C?J$Z@3
P?D2Y"MRF3R)&0TEB?-:4U4YBJQ'G+,&: SB:N'/[Y]D\)=*9 !-'Y4*6Q22Y>01H
PBCK9@KX".J\<0_$_BV3_^TUV9FV3*]2K?'CAX'DL[U*4"VD*@L( :>M_JR]7!^(<
P%Q+%)]\RQY%G75+4$(X%+\M&@$HHCM@M/Q7'OM)89C$(4P!@=Z&@2;5!!)H0<NJ+
P/SOSDLA% O"R%76F_)=PC+2P!>7UN[&@/SZ1!&L*CI]'"ZZ-@2>NZXM!J5@9_86#
P]GN]K(\!(S$8;X032]R$H@81[3E)0*7-3;7Z8Q[T_)8N@([.MK^4&F]OA(F^RWRP
PBH7]1"90$%KDB,95#VK_M9WF06G%<%GP"?LM#%SA]ZX[WL-3&OD6P(J4*!U>L@_N
P9JN6]#!T-0W7Y-#R:LM\ '\A.4)9R^V[ZP<FC%6U%QU[.1*%H$\1++3$RHLA-.6$
PUU.'*X.5A%.2"U_H<3C[I!GT-N2AJLMC!2M7<RV&^@Z:\P>C?&_QP^Y%QU/!2(I(
PN>T4%<".AOA!0!<4D1S9A'!YV1@Z\$X>R? FK;.Z7JWS8:U]^%J,%3*\0ZL; QJI
PK_8\K[ARQJK\%H.<U+$3J< K-SV[&K<L*=6D"MPG25V(V^34H) 3YO"92?RUM979
P1XB8IMZ[?0"O"0""6GTD!"@XAEXX<65A41]&N?V03]J4I<GKHPX1E;W18,[P%H-C
PCIC!L<ZR"?![C"BSN8P WQ.&S>9^-M<_0SM'+P<JM"OTEDT:0 !*>LX'1B&JX:ZH
PZY_0B0C)'&_6]++A'%?O@X-P_()IN'\U4F6D%V6GCV,M>VA^0'KL6E2IJRF^FHTY
PHB6MA."QHG(*=#<AU'*TCC-VHD^UGIS9_P6)<60)6-^;S 2@,&XW_#@=E,O@;07(
P0_E'+\;+4A'T]@!%O;(2H-B)17BVX&'^E(HOB%(=-$^FM;>);]OL-?F "\B>/4PQ
P3WTS_8/)PIB;>A&1&58U1(/_=!BJ*'WCAP1:,&,7GJTV/0JJ3)R(0;1'WFR@&WO<
P0BDRL_+@Y.- Y;@;VZE=IOY&=^]HY1\Z=08J0Z__9<M5"44"/=4R3.J\]+K+KO9]
PF,74SU:O2)22%3(Z?F57@ PH0<W9>D1C5M0K2'@Z\9HUF<3HD)Z08/2.J^W7+)<,
PBI]ZZ5.>Y-_I4V#!^8$V%:;)\?IP^#0K7C9HOU3%5"][TNMOL*$JC(A2\)MX&?/V
P\-$P$@Y YL*4ZD6EK3[CJ_;D@WB(W7-#!+9^A37,)OUF9YZAJ>D^R377)T"X[.#,
PZ=A5!'CN^7[Y][A]I*,$0X;SO_&X %Y'*.0R6'"B;\KIFYJ&W$I4V 7PW)>8;6EQ
P _6*>S@0^-+ /7^Q9FZJ4K$M%=M%H//3=G6P'?%FW7%?O)#Z@72%('3C>3=_JJ^U
PCI;YCTJG]UU8Z:8N":RXN+=NK/01K[%W*Z'/#>WI T/CK4P>?,B/U.CS\1IKR22?
PM_Z6G,1"H6"F(@H -F_X.T-/*=3)O=,2ER>S4R&N>6M /?26P>VM=KD1\EBEMT_1
PR:&UBSZIP$;7=QD0! (OBV^*P/U3@0(3(D:?AZL.>B*6&IPF2R7M$WG@L:P;< 8I
P_ECYLVS"6PJ,UEJ#+=B_?)*Y7J%6 \S,+2]KPX@0)K6OKJKYI_/G(!%YA)F3+QTM
PUY?5)W'L,3[KO<0(JIE-!U;HW3+Q,\I7<V2SIFO>!3BA7[^$>]!\(.W6C%DN9; V
PCR$G,?76K'::A)C6BL.#;7W*_>&L,[9WL9*T?M,=@80BK%IO3 0K*0[;)1G7^WRT
P$TMJHSJGVO"XM"SZ.04S.Y$I#02ZA!%?C.\TH4#..@*)$L%$K\Q8?8Y;Z<#:-J5?
P@Y,%R2,OV^K/W3!_1M0:U#@#_E/['DMW33 @E)JW00M,S!>UI8S:.^;OIE:!'\LT
PO_O(HR#6+&D6-B*'> QZLK+[Q4T0X#,,<:IA?:A8M0, 1B!SNJQ&N'6-GB3B@(]I
P8F*!'G]/47,CU!^719-^HMBEG0= LM8C\2G<#2!L3PC$ZAB6%XR#=OACH,CY9:\R
P=B7P;O0-P-+:8Z#1+;VC"'3NHZ4^9.VCG77VG/2N'5+#WGTBR[GRCY,_X_1NP]A$
P<..0@W(^/N'53("*<$K^ZJ4>*"<$B0!$W31?A#,)-P[*CJ]VRAJ+QZE1V]C!7N$.
PC3^UKCF:+42D5S9'UTHKU+;3%AC.2]"P%HV=%&_Y1/Z+K6UNWVD;Y)KDK0I +2']
P'^2"_NB8TDL^-@LF@2,#,=$0.F<#2_4GGKI";[2L_=D_ <BA%>MR<YL;16UU2G> 
P!N#W$E;SY^HDM5./,=]MP>ED3*TJ663_+/X#5<5"7QU%M7H>]1#M>CL7ZV/^FDTZ
P _FQ,1-8GAK=5/C :37(J5B(A2=&+)K&0$CQ%QJMPO+A7*;B\F>8'_Z'_9B<_"Q*
PNI6FA -Z]P8@A.E:9:>#82#4@*L^640;WO[2#?#>L(ANMDBF3Q:.Z6(L7.^>Q6@U
PA4+B9<A8)-;)ARN&#1W7K&3X.M6^XUJ2_PN?>;AWU+80M"685<K'.RR+[T7$5\4-
PV+;]!,:#9&G<F.S>G_=V<3W)V$(_\IM Z<T3:L^SQ!8#SCDKZY8$.<0#78(O'(N.
PL7'@C)HHBM\.M ._S .!F5(_]."(JAGXJ8"?60-G-B:-:KM_/N?U0RB#M5.EIFX@
PA/IY!W*H PA>E64Q@2S.1^MIU HAZ,C *%2L5M7" 7-$$1A(_0H$58H7>RE. -N3
P*72/)6<P#^."3==R<EIXA)[R/)9SD[AO0$KG99B6GS?G\[0T!Q.]AUQ4HMO-17.+
P=,_HLW5Y0.WCUS!+7C"$X:IDEZ4)!$&*D-LO@%05^!9XGT7:*&<T8SUBM)K:^,-.
PPWQUR@$SBZ@&U?PN;*+NN?_4]$>L1IN,S[E:<FI7\>*XTQ'Q,N @U85\MTHB>TB"
P<?XCFQ'%TUYLV9FY@:AA.4%(DDKJ*K>+'_%[24CTE/*K,,HH7EMJ$;_)1CQ?3B,@
P_"5Z;4ZB9/9]M,]BZ4 >8M#8)QB#"Z=<KTL&MH& NEE<HI/,HE,H1<[7NH3AGW>2
P@@"96FZEML6J\5Q[(LT71MY+@>-P5X&+D"VXNYP!T;/@(8<K^;U^@-1H\@[5(CJN
P<5-PN]@HT%!J\'7PM+&5O[A]=ATK".>(7@4@FOA,O_&2Z"\Z[978V0'AG[O1Q*4(
P69C"V&[E97DU[Z6HD?"F8A.Z4B_[MH2X8@]PQ&H.'(W>%F1A@I<J/<IPEQ7[+1W+
P#3FV5?L<%/<P*#7.HYJ"U\UICYI*9Z?.)53*CBU1C<Q3=1<>MNP6*==_VK]\R?/@
P1Z4]TG#ZQ@P*2IG-[E[%OPR56&<[HRH@T5)QB+(>WDM+C@][L"D H>-&:W/QRR+3
PS\%;,(39S*F@)]/O5&L8L!7XBY=/M#$?BU0S/#L/K*#4/-9S)"JFIU PM#A%094^
PCGT7Q:?ZU=Y3MY@-N*H>]&B9EC7DC4&@_)*B*<**?K6+QG+GE+XJDJHKYNZ_UK8]
PT![)'MW7?YRP#$'2)E\4?QE!/LY$?3(1=M=L':]4H2#:$213-CGV'M(MX-:,:1A'
PE&;<S+0VNIA;.*M5U\3LN2GWD\..GL(&[5GV48HM/I$$)QS@@R-,PBWN$"<4<A8N
PT'H))V'!KY85SH4JT+H14&@-1?XN3,X=UFN;1B&>!5Z=G<>U3L:L:GL82+OM>(8G
PHX.!?:U=KU-L,F31W1H.VSF=OX\JII/<@RP]KOGY;9  R?\[AH?'ZS8W2"_V*:R&
P+L*-.L<DCWJTA">T;[\=7@];MCARN5;(%9/R<)\V#@&!65Y:E3*R8P,5A;X,[5-A
PP"ID%15=0\8LH9N3RWVBKU*!UEL8W6#T/;3#L2=,@2KUJ-6>'JI=V\:S.%D)E.V\
PO!9ZS4T?PWVGX*<++\H P@X?J^MO9!HB^K)YBW3"F)>=F0['H&]1NE)K#(W$H;A<
PH7E?_&)9!=-AQQ6XVB&K&:0-PM2'2QE1BYX_S 9X IH2@27M>2J^U#<%;D_P%M8N
P4<%KW3F%+I>X!2C^X,!J&>S NTHG7M<I7Q\5(061XB%F5J 9ZPC\J2\*.6> _(+M
PWF,0C*,"Q-]M&G[>V8!==K'O.]OH-TI,?0,/_8;>VR=J7(U<W[]'?V0;;,2"BA$H
P$A3.M!%\R1$:<^T4KSOBNHUA31%0F:L0U#*Y1\*0,EB*0^7)I2;<\1K#JBQ@N=H]
P#:VM=)E:/P!Y<2=,$6,Y\?IWZ>_P;L^9CU\ONU!AV=%Z_MPUQ."((#NS>''3- SJ
P0A=3,-B5?+P<;#E^+26NI-VD,RQT126!!>G /JF8Q"@W&@C%H/:K@CQ*%WZ_TN^O
P%G>JJ@3/#"?[REY/+P*-@:T+:/C$\JOU\<N+J VPH^+$_]WSA%E<X]) B28VW<N,
P:Q<5>".??LG>%Y/S+PZITSO_*&#I<G(H"'^'B::J4JDR@""WWBAC>D<?"FAVA:42
P<N^B?D*K &_>J,GUJ-6U%<COL)!RS"E"6KX<UX#JY\I*F^)?K$L(^9Z-D&C9KM,;
P0<32RYJ5_PBG3%X'LCF5,DJMOE#36T*P5)#GE\8\2L!GA$'1$BCHT>P8I1EA*&6\
P\AI332_%C GN^*(7V9[Y?VL=]H!0J8,V.(68\39&%&HG7V>4DO%R .4]2_UX1?\A
P(^TWSMR'7^,7Y3V,)Q,#(I<2G<]F$[4YE\M]('&M->L#<]'4'Q7(9=NG-BPTU[A=
P(W<8(P7M_9'*=7[%/&-+6D>5S1?D$:EE#,=W"AF1)OIT?$)0&[[T7UA,K&;V3> 2
P96,>\U ,MHCX\5J&.Q(])A4K&DQ!7) HMGCV0 EG5 ;8)OSS ^%?E&H'QY%!J_)D
P_FGPH;BLWZ)X;LCG%/A^$M2A.K1M\+474Z>%9C> 8<Y=\P/ZF U5ZNW*=+KK;@@Q
P\X(9_P%_235YO\KA-(BR^/GY\R+]P O);_6)8G1MQU;#X 2:VVC86N[/)[1XMCAO
PT"^BOXTUFP=K,]B+D5.9$<\25C%P(+<:G<F<F(]C4]$V/]_%N.[6UBXY-HGY1T'Q
P6^J#\:(.#C)]NM'/'&-/J) TY'(> [M;7Q3#C#4+]R/"D8$R1=],3<_G-FS3*Z-Q
PP_S8S8[ 4-4I^+7/Z@&J!._!C(9")E.;H,6K1VZVZS+NM3FK-'R->.?R&SI('Z[^
PI%V(:QHS/=4)H]/:?0D_QWNI+AT5PWMFIVC+RY*5[!B0L?R5")CPDC76&'R4G8GR
P _7AD%/YQUMN?+.HLC.T LZ,#ZA0>.!*?)X2,.A!T?-# E+>=>DH!61TA+R"D=PB
P811S#A+^N+S'^STLZU8Y&.VT]:B#_%JSD4F>=$XNN@R6]T22Q-?C*GXZ5OGAA P4
PH;PB'"&XV$"RR6+**T:WOKI:!J<4<M'P@G"UZ=%G0[:G/#STK5%#KS)@M3?(S(BB
PA<L99=PDL*][?W9^+8CPZ7QQ0 #6MP=QPP4WFZ@6'$%OV!6ROG\L-Z@)%SA0T9JQ
PRP!"?*%WZXY>-#/))Q7%6. 08B@O_-KYK_G7''F3@H.742!7J[WFOC?O7,JK "!)
P?,U_Y9V9V-*NO2@7<;S+[-$'E5ACW>78MBLD(4M[C39C-2&EF&6RF!MU!JZ0S>P]
P:PX+R,>5,YM/9J)3U5,_/6\_'@DE3+RBC/UJG?D?M_34(,!L2 J954--Z[F9ZWO 
PDN'L_)M(>EB7)S-F=I^+M0K)P64L9T'[%XPOS^YV$%Q,L"X-CRX4+DH4@P;]3$<!
PP509-_%ZG#F8,UD5C*PY\Q_G,"D9U5?1+J]8K9WF[!.^7$N9/#E4@J3M)>@Y.KOY
PC8R<F?!55%.7+C?GPO*4VBT@W42Z1F-.O+OKWS?8K5@LOI.RRS-;.-FPGLMTQPBH
PUM_:^4=7]<L\[2"#&U;^>/5KKDVP25FD6@,BLFNRK#?'P!UAI'3ZZ%?5"SJH&A*"
PYZ /H',5+/$W=;;"RBJL:IK@O[1Z=@D?>=9_\G$1N[:8@!3D32 W4]WJF>UT)T4J
P)5'A%8'G=./Y*?%,L&L!:%Q[4N0N/9+,,F5D8=.9CD\^'.A#JI8U1BH(_(_9][=>
P+!"/O@U_X/4UJQO//ZJR_J;B4.Z\\PJ R9]?1VE[X2NGHQVL_F7&MLQGIZB_E;6#
PYY<VUM,X+3"<I<?D$E4 A:<5]DFXFJ[&6*/6,&$L-,]9W$#/10SI>/-'P>-G;A_,
P-UEK L(C*6U:)Y@!S9)B0&*QD[URW6OR(I(#Z TZ@I],EV?ZF=2_LX!F>IZ1",%N
P !>@K";8*GEZPMDACR,H-3>AI-@3_)5LBBK2P(%CNW@<;DSM@C2?'RBCJ21R<\@2
P"BDJ0/%0CZER %0<^3]&\&\W=Y 8CP2M'HNB'76F'_#=+($30S9(38FHD]>)H2>=
P9BG$U77#[.X%:\-RU_@J72F81BO4RQ]@ND/Z;XK,)WTGR[L04YQCJ_,KM"G,W6#>
P[Q#\I51D%R>\W2."^Z1=D6L)XV<#^I!J&AN@K:?N)DE_N0',U= AKC\)X*^IAM*6
PQ67(8=CM)>%OH7V9=<\1YWW;!0IL98W6\X>Q'V[T+?NLPA<,^CB/Z/PS%#'G9FM]
PZG>S>3:G<-MC/A[A%_LJ;8SM)=34@%Z/0+Y5[01:,3&*AV>EA[[Y1M)JSIR1^9-2
PD9UC8F+V:UOU;W?_7F>-M8GMJ227C&O3%]MAZ&(**Q,\F?ZNS^B>P$E+GJ2O$[//
P4J>0UM J;U$CO+Y'A2#<AQ^Y;IY+$DV<<A]W$; 0$.%,7W:HMBJJ:1&.^[FH]W<9
PX_M7[/V8[1#S+9X'-E9,/(*R8)0@"K#@H@] 0CC/E41@=(#U6@(.E#S7]:/,$0>@
P=ZS7A03BL_^6^PO_$(3E]\?%)3T^8@X ?J?:@I6NE/&8RTY F_)])+/4R_ORC_KZ
P[KA3(L=K<_$XS4K79AS9"H;; R,ZD_AOGR8W&DZ(O?T6519.*RTIMWG2/Q*E[<C6
P(_:GF(X%H\?'L['W6J$_5MD0.U:UU+S$)@.;W(9%SK]/PK:>.YEN]X/=ED UI_NT
PWTSO?9@O,6U.\JT<YC(Q >'^VQQN?H*R+?UH?[GB5*3MXM6B)9M^CF.#!M>,-=),
P>M$5$5<&&#2ZQK22HB$ZA+HTC/["9&WH]9[UB^?QYYY#'"+UA6S,GMA"[ FV+!L*
P+)4I@UYQP6[>:%!93W:)U0LVOJV']3*)W\WOBA<=]]V]M>!8C]%JZ5I6DHC71PR>
P,96=P>:>RIK8%2C=DMOH+GPFD^\-2D%=X#:Z=A[#LP2E[0DS)1 .%XL\2QEV"^ V
P#>JOA0+/5R/W.5K5+;E/=D]=?U%A3_AHH^13XN=:(/PL4SX_!X-K)K:C2R)NX,$\
PW%8J*KR"S!HB=?OU[.;T['C^J85S?E>[4#@ -[&<(,,B*7F&:68L,2RE15^W[I.9
P&U#W>7&9V&A.[TL4]2L-!]1Y3;Z9B1Q0(K&"I;;YL-U8FK@+82ZI]R/\CP'#9^I3
PDP@/MPF473ELC1BEX6Z_ZBF$'"3ZSWF4TX. R%FB16W:GCZE;/[SF\5$V^D(F$?.
P0=8ZCOLT<*5R0'EKRI&>;=:ZWQ&=X?&IGE05-UY6J"HS$.3TC+>6 \S<F/"@[G?F
P(Z%G?B_YD4.&,F.![G<2G6C"A23'(QB8$A"L;^TP:87VJ,S"*@(>%2V:G;\YV9":
P)W-2S8/>MYB<%@G)#W:&W2B[$L'0JE^/-3*N6A^9DI?@BV2OS2PT&_,[%^#TH<-J
P BKYS_LP$2&$A^_$'P0B:<$8PW[P4] 9PK@%]ZQ#6+NN4RX*@+(J_.;S =#-RQ%S
PR)*XSE7AM.$? ?,(]A?^7Z%;!G.M0+X=[V&._'"]WB24C<F6-+4?"7QJ!C>K1-"[
P/GI2D=:OS,+A\B18^5CTB<+#!.X4:KV4^8Y@>&*U)3TCV7N@[(\,3\N.CDCP_32T
PTW@ ;C'TA<U@G$[E"U+O0"K7VO(B336Q$>$MI&Z_YJ,KT>ESS!> A)ACB-("VF@T
P +MF#H@=F"_--(DMVPM;/.ZC(K\B[0\7UC7?S<1]1FIV&0=B.%#XRVWN177^9C$.
PZ;.,\&;3[%W2^H>LW$@WM>K516\7 .,<$U2K12'5,G[<5M@&;DHXV,M"T+2R0,0L
P$]RT2H7_>I:1H2[-)64IY>L8%'+80Y<=UQI'";N\WKK\!OP,7R]58GRP=XF8B%SB
P,D-)Y\XY1&7$W=*]7>4BG]\4Y8]1$[-R#<+N#FT)3&AY<X.U998:W%]JCM9HH7[^
P]@Y;>EY"T_MD4<+$>/AR'R\K1\/2<^<Y)-?I9WS1"X6 5P5!SFC'\S&P6]?58?_F
P]U956+0CNWJZ$E7.FEHXJ<:./"?4L1U*LSDQ##7QE!YCH^+1N'DB5<$&5[QN,05$
P,4VSF(J:\MT*B]^_R1Q$#;!:^1LQYMZ8IOMX=0M5U&^N)T*#;,8#\!<H^SD41IA7
PI_W,H8>E89,\$^@J]0K!>@#E806"HVM1VX1? <5]WQNSU!T32QTB(H,=@6?J/>DZ
P%7D5FQ.C#7\I# OZ U@7?\#0'S'Z-UM3T4=E#U"X_5IVNXYFG.V9Y-@;Y1@\07#9
PM7C1<Y>0]HX5UG$VHMB_Z8ZWV!/R(#$P2AGY&/AM\R+47%3C1:9QP6O_MYCU'/XA
PZ3OH+W=HV_XA1_JQU2BB]1 2^R7H*D*N?E/9:W@ UX!H1R7M:ZJ*L.^"9UK(4HVK
P,,A[)L(/9CZ"I5Y^$?8O30&_GQ4Z&KL-[.!G7E@)!IQ6I=)80JV9+*MEW.8+;3U,
P(@Y>3<><NZ8FV4(W4>EW'$-.4Z=K_IU;!-&;(WP?+R91%^GHGDS%.0[&$/Z<E%*V
P[V?.;S]M$?[_9(O:R(=\B_<6XG>719ZIS_45XQ?M,E4]<1A:]JA1%W$(O1%IJYPW
PF.Z&*SUZ K;WPZ@Y#QJS<]?H"+'O3ON?_0 AB B4VB.TK#5&-S@BZ$;X*AM]P&3]
P1I)6&P04GL"VT\_;J(]EH51OG#U\V!T#]9E%D%J6F:A\GOPJC-D3L1NYRI\*14#)
PVZDD#@'Q8L#-K>=8&,<W3A/=^FY:$/ MK6A&PPRJR37J46,;#6ZULY9\C+PLP+*P
PZ?Q0>&FRJMVL57XSS1\$6.(B^N]RW_7L47N_ 2S9A:/A6P[O+R>W&SX4*DC\23"/
P+ 78S^],E_'IY^'B;[_P,!%UZS/5_M(9$?68C.LJXC,NI9Y;,!J#!E60("\19NZ,
PLPF'[NDT/KB*U9SVKF,+NWHF3 X!]&)"YU@8-#Y;31YLV1]F>E.&CD#"\BJ=F .T
PBE'B\"'*?D7)L/5&#9F[6%5S_$8><$\NU7<.=>E'@I)JG!JH]+B:W+B-3-HMT\87
PF>=E]*'ML*!J1M0#:0;7T-8CK:8[QJ3>=T!SUH0.+3>3R\4]<<M1SM;IZLR<1+)6
P!U'?_[HHO"[]ZLSB<MXCMZ3 ?7_H4AXQ=DNB4GYQKBCS=CM?E$&;#J"68$CD09S"
PI(*AJ!X/=Y1JLN.2@X'( EF5KA,,P_-XW*9 0@7>O&: (>S*_.'7SQ;KUOUZPS2N
PY[H8C-=VKVG_S(P)Y^,[I372_MJ'Z@[6>7&[GAO:!X7@VB% D]C.LSR>+CUO0P%2
P !F#UA=V4=)='/+YV!X@/=][#JPBJ9/(WKP7MFB14SWXZAUECCQ'0U#NX!A=</[S
P3DXU[NO"6TGK-(?$:<V&)D^#!,3JDM9@/!29H@^FC+6IB8^_104;!I2XW?;60L7#
P7P??7TA\1_1,1?&[&6X0R)9Z0E?5S&)"YRCT$=1LF5?\--\>=26C\?O<G\A"<TR'
PS!%J5204[P2Q79T/N!"?H)X,L?D$7QT-RI!;NA+#,TTW6S);@3U3E[;TA;/LX>+!
PA\TJJK$5?$HH\U<K^]H1AX>>Y!I[PG\,"]W?V**80S7(]R_Y.9SW,/+5SUG3A+"*
PW @\3PT:#N8\S$&G.X*4DDT\;I%"KLSF=/UYQ[#(8@Y S])Y-MA&.LP(>JJ^G FT
PB-D"Z6/1B='3%ZVX5*%<V$9/O33-JM L ;B9G)?UKW:"\TR-XVG5[RY= Q=>3 0:
P4"+@Q.%>>OZA&95;-(F2CYZK"P*=[S=Z.&+++NI.T\A#E3MRQY">9'-P"98G_XF;
PO6\L"='@\6;;>:!4+!?ERTF7A-@Z7>@>9/=N_Q+7&$O,4%#0]I2$A^OM^J-:U:"=
PO3?TA(AJ-S\J\O4YTHI>@LC7P-Y3>"H-+*-Y(8CK?8LZ#\SPE,4$=]OINKI75\YP
P\[ -@SW&H]" IL+V#WE$TK;L+V/'Q)T%%U\%P-UYHUYZH'+@K<1U/5)=/E'Y^(S^
PI,D^$TBTX73VC45_8'Y:A/W/QAQ_F<-FNWGFN,>.50_^K>AB8=R^.K(XUSV-F)B:
P)[(>P$)$)=+H^)*[/:Q E*RAKF#T#+2'&J=#=4VFE3X(8@IOT5?^D?'&AHU'K!)\
PY+TS[1JM 2WSW7 &1"H?:/57N<(VLM 8G(1I_UT,[(R=C#Z$++M/M68EJ]\(HL>N
P7O"R(QOG,6BZ9WBVR5_ %5"X;T?,QOJN3 O6Q<8"8-F+H%= =G-9ADZM>VSE061M
P[[859C^2;[5/E&C1>G_ <B]95Q3B4$],4E8X6%)>'9>%21G4E  20!E%.DQ3E%=+
PSJOJ E2DXO#/OXH!LB!H>CN+_<]<U+Y9I%-"/$[^O84K)L6C01=+MZC0<+!J[\FJ
PD)FB4IUV__H['KXQJ.?]3AN<]FXPI,TS%ORN[K,-L:=ZEVC(5FOY,B]P!%_)6*5_
P:9Y%QLFK<V\%&()0:%)(_.R[DGKA-0\5C%7 +7K%(TY&?_S71Q]L$G="7&C9_,*4
PE*UPT-MN35/* [SX9S5525*RNO@W6@4"L .GH8 >F$#Y)DOW1[=.=O-!PUQJ.B0%
P^'U^.YA]LZ3$5QC>412/YDF^+R?PM'GU+[]9^U:I%RE6ASD@L>=R-$XP@R9'KYZG
PG[S93V>U0@XO#BMB];CZ84R:*%FP%ZRP,4TYA78_C_)CAPQ\G0DVI YQ)&]?)YT'
PUH8ST)J[0+ZOVJ4(JBYX& %CU;C!=0JPO=W.M<.PDP)_=I9JOXOU &+YZJK#C.4S
P,&R<.G=1GU9;<V1RM!@6?M6L<D3'#00/[T8AGI*!]@>QYUK.A_2^[E-/$K95'ELK
PM_I,!^]@T[0A ]:E>E0Y'-U*:KE4_@IWF6&L?QFB.'OT%$K\HQ+L V=\RKPOON2'
PXW@)%2V]0]WH2HP<?S:B\=_-PXIX*70DM2/[U77IK15U#S-[R@BF[/<A\9'T#:,3
P-C60&C7X2FG[K'&&W6WG#]=%5>Y]V>AC_;$M.WV4NU[?L[C*-6K74DQWC RM(?J2
PHPP. N&9X).O&:"O4+;;PPW9LY@4%U*ES&N%41Q\%LZ!K H(*C-Y%:CF"HK0ES7K
P+70!(FTX>-ZE+\LVY'3X:O+CIEYSC-)2P>-0PI\BVE>(%E\=JES>.DT;(QUD^VL!
P0,,)NL%[O#M"@'/92G5>'KL"^_#X89T<_9[LIPV9HW)\#SE0.53L>KRAX#5NF<TT
P(?2XT^.<WYIF$2O80A9+*68(MVA-Y17U7$"UFMP$[W;\R$WC4D9A<@X[=VU)EL;'
PA$E9&H*5M/P[V):,#, 7Z8IS''N;UR@NHL;C+"$3>\[\$5\Z))J)+_D+![2S0<+#
PU+U00F/+0H%5%B),JM")%&8?$X8>,QC/49UF3$SYX; #H"GOO 7$$07)AUK=D&4>
P^#/IK\^]^"@Y)W%I-)%VH[O#P,H6%_MUD\0=<C[H4*HO?F&)D/BC]#;;6/Q> R<9
PCD0J?+5>&NP8]@>4OL&; ](+SAU:%S7PNK!%#Z-YIY(@29]UN$%C#9108SLW^$4^
PE<PZ"RC5S>H?&FNKQ4N#!B=90%NOHIO8\V4KXZ5N.D=H?-2+J%98RNAG1:X*9400
PNKP>O9WC[%=]J<B"0;6N3C>^<_I;5LG'%*0XJQD)F\M-LCN+N6<P^,<BZ^#8BLGU
PB/(D0FE!A:M++0$IO'7_2 &0_D3$K=#.>M8M-!!.*"(FLEX^>$&S6 0*Q*Z+N\Q[
PG\,0XJ_$_M0^;%"-V8LSH8R"DIH[:GLP<'F K+1>=$(>I.2S(#6*_#P[OH^V/VZ'
PA()I;K%"?BVK29B#$5BP:M4!XVUKD+B[5.EF-C9^-($>\LC-3Z/],VK>9+G)]JO&
P6@,0088<[?5S%V39?8FMFC=2PR.(82Y>DXWJ][!&EN40(G\:E?N1VVW=441?*P1H
P59<RADT?>7I_/Y@8:Q>1JUZ*N"W8P,/4 \N3ODY;I XFN16=XF<XPK>Q JLKJ7"@
PB4XRG./'\DPA.*S8O!8@*]-N=!A $\Q+VH8(R?9W$5 '"K8EGM=P9/^FAA<.!<[%
P3FJ&_PA[$<%RP;(B747,ICZ>^J&+7)'!7EQP0;(5@TB%[ ?Q74"?2E$X(OWM6<(6
P[<Y^=_NLA'>LDPT:MEA>*J8!?03N,Z-O$FAM;'3E,BC7S4D9FW_->,7C4%X[->;F
PLP9*1V84[^9U*0Z'Y\/73Q"@@7VL1Q;;Q7Z&HK:;,P;#&^I]"*:4@" +B4H->8UA
PR/7%6DBA-"(U&Z)]4D<A]J^V^(_Y)S>YAJ_0>+ZJ-Q ?B.V=/ AOM/,#,@?C_P<[
PUE,_G[4"19E,G)G!9_?3:F?MA6.PH1EEU+4Q=NM(SB_MEFW6.V>KM7FJR"T_LZDB
PN"_38*/^,"TK\C^LJ*E.20]/35@1MSI"Y@]RGGWS8"P]R1_X GEJTIFX=UGQ3XOC
PM64V6F\EE4[--'Z:#5[!,(:SOQ5T+?]GM3:]=P]W:$[<H]JC9$?3J;DI99&'**D.
PIE)N?5'?*KC_N =#294W-?$$QPHI6M<BWQW"P"I%U6P6JE5QM; )]X0DU[NM:O^=
PDCL94":SX.-CFFNR^@?*GG%>P82J]ZHD(Q<&3]X,17LN9+QIM( 2M-  ZDQ(_D?T
P63D12&-9)'WZ&)I'YU89[_P:+HA6AW!]?D@$B@##_8PE8'G R0RJRE:O00(D:/7]
PLX23)T^ '"&O5N3_+1RXR*  \1OMM1+:E_*J:#L_X=0.D:[<,-O4Q1+TU9)8"*X>
P!1@?/&@UG^R:_2<E[-R2_N6#<)QHH"#(AS^9RJ. LVDS!T/X?4\F(>D,") [B5BH
PI0\;C^<](M+#EB.U]AH_SI9M^Z-\[YRRUP- +IB5Y]H+3'=U!C%D^#TXS,:45XH[
PQ:#,QY8]=R\#R'9]9I0%O=4^Y0=C3?GL8.E=X_-.R-!LIC%"Q,\#&R0F6H1_:5>@
PY]V4!2'^.U1[++N4;^2FY(,7OFR;*DSL9;Q  P5@,)LS4UB:V$I1N/H^=XJ2A%P<
P*4QAD# $#RJ"4PZNIVCGK[6 G)*(K>DT!C^+'E/S.@9V#Y#\1_:+%GC#(,M8B>93
PQT7.Q*K!&23YVMGD'[F;)P-TDR?^6:_TD86J4'YR '@JN3=C;_GMJ<7T;T^1-X^-
P0=.:[8K3Q5-RL[:6):D&5X2HCI:,U->85MF^Q-2_80LA^"<_P).JJH2$@*ITWLH/
P=@21-X8%K>)\K7!9@@$QDQF;,QR[>92:!8,/[L#%)OJV;OU \]-^+R7A+5T3W_CB
P>^37JI/6G4\J]B'UF,+_(H+5/@1LV@^< O*&RNL5ED!0<_$KI_[ %RO7=?;/HVK[
P!1=JK-Z=+K>!%KQ,2S3=$[64F"#16X[,2[/O\)'-R8!X)W&1XZF4(FT-*AZ)0(?_
P]A$TP0T>4'2LY]VF?CFOV$+Q#CU&DGJZ_Y1'!O%E/VWXWKX7(H9?WGO_BFP,D*F:
PH9'=#'6WS4WS?1,<F4/7EO]0INPXY.TJG@6=8PD7,%)Y=@6L'>K)C='%]=AEC)67
P%ADNT,Y^W=:#K2C $"_;K^O,]#ET+<*7=H0BP_;%EUG5983DT@," I4%6Q#>HXA9
PA_><A&E3-PY%;(>Y$ES:3_YX4*EE]<#HN]"^P&>VTS 5\X<\5B*>EE)DJCHY>_H"
P3(%^AZ!4?ERFOPKUH?C4E0.YX NXSZ+FX^-Q0HIYQMH=*64Z?2*\/GK1U[PD'Y+&
P2AF5MO;MH(,0-%5"CLEP]U[3[;'B=!&N_4"\7:('D?M?DU,)#Z)H<ZEP/W8>N\L)
P?:M:[#I#* #%A'/RC17-X8CD-0,U\6VOH- '@1/W6+%;E(4ZNC+R+F1Q'X,C"1?<
P9SW\+D#\AP075&2"Z82]5;F_D_;/C LV$+RZ(* "4!D_D8O8Q@LV(VZ P(X+$M/E
P?C;HW]ZHK+Z\)E^8)4@7$\DHN\NHOJ$=NF?J%.V:#YZ[^,C(IW;J2(QTYU#UL;%<
P<G*5ABQMN]F8J5[/I8#? [1+0,-(:[6/-*WJH8] 4#>&$0KB(SB9_ROS@L%_+2,>
PL4Y?S(]4R9SHTM)6>=-(WV8LG0^OI)]\QA(8J-U'*S53#L<+@#]*7I1$Y/D6;GW^
P]S/(=Q?/87R#_D- 8.\MYB\#I,(O!\Z<-$Y4]-GGC!88HJ@&J _ENH.,*7IK^\P<
P%67J3N];QN;2UPWY>+QK4Z OW(ZF- ^U_70%D.-5C6APVN6'.='Z>@E)Y)FS5$(V
PU!U!15Z31PVP[:O1T\,>X6'00U\'9@+3-5[\>W;!'I>?^!!&8T=:[XFL.H%1N5NF
POQ4^3'5(H]3[Q9"I#B16S+T'BKV'D[4=1[=?[JXTEP*]SJ+-M$D,)GX T>J-PV3F
P;_.^N-I5IJBL5B%U@[^.$RQEV9<7XWFC0X3&MN_N:@88V!=B<KB46/#*$X:><B<7
P\';+_312F<.VB>M>C08"A>NR89V1$URNO?TJ-BE=8$$NO66+FKN9E<.Y1Q/"Y=.;
P;+8?6=R3_:7QC5@?3F4*T9 EA%C7YONB3J#[(OMD8.U3;WF&#1.W/XA9R93DYHV?
P%)0F/1.E+@?GI&MF??1 VP=1A9 &\TDB&\(]UQMV=K;#+8\\M,,02[)F #=3_W!S
P^U]_6&-Z9,$D[=;PHB@S&40)%W!;.*=+ Q[0UA$EST#4)0U#OT$]-&BZGKU$GC#!
PA_[QB8L0FG=NT4@7G=>-56)]RO3A'8WS.K"!P8%06_J=!K;5?>NBP,,^^&EX5+UG
PCPK+?-%JRSBJEY:DDQAS'B"2I[:&]NYFGE38(A0U*F&*\B,V<$D&)H33BOV6B'ZS
PKD\I]LM>=-S5!IEMJ02%FRT#J+[XV>:*(;R&N%H1+-/NT1WSGQ.,,%M%:=)JZU$B
P"/IE>RW8]=/PDC7TMXY!BSD"A39]V*$ZH[=TXW4]Y-R<512=-9ENHC_QB-(SUCD"
PY&UK']#%@#0,'6.+#6/OMP&4YVDA)9J&!.+Z[L@&(6F?^,0Q.5%&CTB/>6(OA%'X
P_F*.3#N%BILIN,F8!FGEH+U98Y,$LEK#5I668*7J="X?U+@9Z59@0,HA8'JH2,A7
PW6=NG0])?2K_Z_W2&,= ]A>)4_-*@L8ZE\+5[Q[H7":!KYJ=B5BYP/OE8\&>DMW1
PK.UGFGJ-,\2C^,38^Q[0W2B1] X*$WD9?I=?/X7]6U 37XC"C_N9LS,%6E ?F"? 
PQ^U\V=TT%] C/WEU"MTBB%^A$"" 4[[4@L809EUY@;OF=<" \?>TS6[%O%>42@^5
PPM LFU$2Q][M*F\"%)<[2W)7)7W$"[&$TI<?",+6%(D?3^.W^Y]CD!KCGY]_,8JO
PB3MQV(U,2NO0A*IQQHZC2[3L-0$KTSC IGQ'[8;K9860>M9V6=R@G[U,.,5@17U9
PEX')?(8KSFG;5<\$01>120N$K&W7Z9IAQ"W)G@['MXF!:;WA.1M9F):9]-VCU@:.
P:G=\61DE('5(W= ^$T?&H6/!_D+CH2X-I2#&&RM"^:&G2W09,@ORKS3"9M&:^"Q,
PRX)O\'WR"9\$S#H,O!)P;978MUZ?0OFA7\RKO2XN99,;.[F=@^&?XUAP2M 3">#(
PRKEIIA.X/>ZW2B(A6N^$UQ@).NR)\L41SBFS$:C31KP,0[;TU*XN84=CQ7IF-(_B
PD_KKR2"7TX.('%G'UP7I 19)GSN(,I _\,E3!,&#CE"Z#:HK7^)(Q?OV.7F,0.&S
PV/;V\$C=6F1]G\G_@S4@$"_F 7'&#!9+9< CEI^*ZUVA&RJ+=+V\_07M3DS88LS$
PXIN-Q2F>!PG;#:+Q:O71/F6(M'2B!,9#2^P6#N=I>J\X5V,3VG]B%S7MDJ.?U1?7
P2I/E^ "52PH6)?KG5[<4'A;^Q?T7!(KJ0BS11_#3"'':!D8WBG6W<G;(%TW W[0$
P-R036=L!Y%NHU'Q]@0#@Y^V'IIS]- DNJP4%TU32.QT$66R6J[F6([$O>V&[<R<^
POH<ATE.T!.220,E)>R'J6N5K3"H'D01&S;'Z:Y10(A!#T]30GVHR[Z"!VSO!/HY0
P%_G?&VK?42EOHWNU"[.RGE$G6_W?C=V:'7K:AZ%PO",/]CL[HW&,><6X\$1/-\'1
P>"0,\(_$%9PNLS$)X?[654KG$)4$PH!TN&>MR+(W#_9LLC;R.AE-W3VS?G9MWV,N
P$1#3JH%6Q'GGC$@YY7*G?:Q[,8:&UQF6$*)0YJWM3'PJ+E>V;K=>YQ_%\!_DAX'1
P.0IC.NRX4]XXA]@7AENP:.Z$I+6L\V1OUW<\4_]J36N0N4"%FA=\0%F=B'4_@US$
P6YLYZQ46(OL$])(> OQ+T39[7,0Q7[^H8*IGYQ9 DW]S7)C4]=WP_]ASOF'ECM,:
P2_)L"G_="UXAT7=,8U=6H>?,4;S7\+'Q.4@YPU&&BVTY#(XLMZ_7(/G)F)YKL:.N
P=\G$VO2ANEU/#7CVXP!U\;2YK69A9 -Z@LOKU'/H["+=L&'7/^FN).'/.]!61[-E
P]IKSCX>[Z#5ZM4.B@X8-S3)(W[/_C[,N,-%+LSNC (T &Y]-]=9LQ\'_D\7[ZDAJ
PF!%&6;<ASN<-?1Z+&'BU_B^@=])O-\CG)G#TWG]^]]_N%Y#);<B.Q]1C:L9VRLE[
P.AFW2S:TF5 23#Y=WWF&KA+[UTJ29?Q[!T&& 8R4YBIW0>%XR(%/A &-53<)9EE@
P_B#5IWQH)CDB79,W"1C,[5Z*V,O%4P5^]R$)]UA72"H8E*<^-*#6 $0KIMGLDQ+Z
P,9ME)K2'J4I(D2XO1JDT$9MHN)NT&?$N//D4C2E$B\&RM"X$YR@U)5B 8?*/HCKB
PF!U,DNF@"[$&=ALLB"W+O)#$&'81'[3GZJ>YORT:=- 6J0:NV"RE8.MP;)-73'L6
P9-%!=N>$"A%2=UZE]C/F!,CW*"V2CO=0L)^?8;WI=V#BS9[GS[5NH_E!\WYN<[W,
P#0,2\Y<HI":3@1W"'J*[\ZB?[\VJ"1R:\ -HYS5<F:NX14N%)*_\J&9HJ)\-5\Q8
PG'/%AO$[EKQ+W>W( QX/YXK'UA9"4JGA$S>LXX^QK0_4.YDIM*W\'!U:S))[2[7Y
P\+RJJ88:E+5XA:U!5T\$\WPZRM70HZ>'TEV[;/PNK&W[QBGI8^/V=+-5-50RF\S?
P='%Y2Y]RL6;+D.'L!:K@&>OAJ+V=6CB%-BN9#SI.TSY4_YB"NF_V?Z5H(-_?$%JT
P1-Y%R1<J8N3:3>0D7U6LT<!CZR2.78]BFJA.*1LWRXZX\+Z%"A[+/%!KS[;<-NK^
P%6 +'Q369\<<@4_H.5C?2<1>4(/*\/:7ZJ[J^=LX=+OX 6[K=X2+5A^]@/Y?=N*T
P7!\KLJKFVSP*IQ&HNY H=/7+!8/\VS LZYVBLI'MI)D0&Y6WI$ ^A<8JI^D,2]R9
PFXYN7NE7!?COPJUJXH)@(^TH%B/4>IBLHUKLOIW\XZ_RDREE&D9R.]HA1B:KA)3R
PLAL_>'T]WW]6$/"8'/^6GH0=C6*Q+9#(I[1%QXHZ6/QUDJFKQBT\ER59?3IA/-,=
P?AQ0X_,!/7V88M<3X^F*J-VKF/L'FKL[4+W=(G;[6FBZF4DHN7PH5]3XUA[07I:G
P)S,W#?=_']MVI#I%*US(+$*:!F5P73&=Q42%=X%>ZB>E_U%]'M@_]*: (K'./@9.
P6KFZ.'4 \BJ&G&8!/W%A#F?D"%0-KQ-*EE>"J5:==*SAX>>>LO"S#,I _)A,8T(D
PZ1/I""H%F,[M,&3_.JTS+"BW1.>QN!-[.*J@;1 2NK^G6K/][KNV/'>F]1CWCDTO
P./8MCN\-#WAYO39']_!_= CC9!22.3*>ULW5 OD2?)Q#QG#J7\[^;4A[6TM%I4>/
P(!]!L\N^NJ25KR-:RWZ"BY'R+]_M=3XNE>GS@^CZF0%,G;K)3G.Y3\>0#_C%5"H?
PJTC\)T_/$,&Q+]?E%60@*A+!Z"G=I&EY:B_GU394FLEG1[%-?MZ%V>@]T^UME)WQ
P'H6T9RB":L=4ODM_0%^$4)]G?<>:\TKPWJ'YM#"DM7309SX;'=/%D0J(7Z8=?OR"
P/Z"BM''@>S#?$ BL0E_'C7<BIA'D\P)60>@X;1_TQGEVM:M9DS.T!L+FA'O@#1=H
PM=&%'PO5*9JZ,>N8/U9JR4+&7ILN%==J2D*F9=F-A$X ]1\E9GPQOVDP:@"SJL7>
P;>P3V[B_K0>VFF$1(/W.=VV'WM=/28")G#A*=/B$VMK5WAE_3B.\,.":S/*GOINR
P*Y^>-8P9$$[L;.O'59]@+]B%&Y&P-N".G;2)UI5$Z]0]:#&E\PLQ+Q"9/( J^C_]
P7_3+9RYKX4C[0FJ%D'>'U/B17K-L J(O;T^G\134-9XTWG39[T]#F";G/J7_T7M-
PKE6O/;V/?=W]/_E3.+>44\4@%TS2*[-03,!#*FT#:K'6H>$L[MN0(6Q)$D=WGY6.
PQCFJ!14U,E5U"AI.TEQ(RTZGV<V)!?(\05SV#SF_8?N_3V'^&-82><_V J HIS1\
P():;(RWL]5[G,$[+!WS!5W7Z!1K4>(1"_YK-?TN3>KF2'G 1#8",;7S$,X+Y+EXA
P5C@GN, 2!PSZ]_N4)2\ 3FK_XS.RW%.8L*:'\UL\+43#TJFZO$P.YL@'7 BP.DI#
P'<6.J*@+TI*3Y2XQ)LW.83%I"6W"I^RFESB2"G7U8GV?7F[RM[0)Q2K4V!;T;A^J
P.K!P@7:MZ:55,,ZH* L\"C SE6X/2F,IQ/_O6\ /?&1U3!^,IM',%?1$9JV0OH>A
P=/65;(/BQ--NUS)*FL-A:^:?M,1'C6.$[#.+KX42M%V.KXI>)=)]>*7A!_$Y<;\_
PMRO(I&<;,3EQX?K3 \6[U?E1C=/50IO<F,Q* 1ICQ2)[V!KA(?B"IL4JF,RM#<33
P13-;Y#P)]:7\_BI8H9\HA!44#)$]=^Q"1 D]1<AG5QVO%\@+].->\XS$+XZ57-7J
P$VV13V#K8Q$9)?/V6/:CM1;!%LR(4) LKV1H5RQW_%!:1(--OL"HF@2=M5V=2P0F
P)_R'-O6DS?)UH,9NI]'"0BF6U]7))E_WY^[W7?J+LP[\)'** W"'#P8?@,Y@!JU 
P4^$B:$ 0!URIV\I"/,YT(5 Q'+]FT? R]2W1[GF&%18FHN3-H-=4'_4<C5T\2X_"
PGM7H</!?DCP;]$J1EO,? 'A S;*.5[EGGG%M<TA/0SNA'X>C/7@\=<]E,>F<?M1&
PHJ@KUJD@<!L\*CM?=$ B0NJ,$Y1YZL347>+$YB*?NM:3<X;=B\\;5(N[EFY"7B]4
PT(\.$BGUJ@_O@1;^689Y-4M$QPN-N=*[0_/R>5R(94?_;[1_N!0S2!/]*M1<, S/
PZVC/MD;T<B*;$)6>@OBC<5W] F9I@Q[I@3C2X66*ZY)LXRR=-<L[1-MN##/!NT]$
P>=1\8\'I#ZOA+?FN2SP[FL+\+7T+.V2&F+I&# :V9OL\_V.F_+<23-AH3/@6NE\8
P>-:)JE0]R9K/[@'/@2SD'\X#94=&;&OK&.F6-ZC%"TC8I#]T*:PY,>JGI5=T^NN]
PD 4.<+IB0#$5="\&XD4#0OI</,#A\[#@SH90L6@[^?XZ"?B D)X=D#[=A^+$55]H
PPIH;MF$%?TB[A4QZA;-AR\-\<]Y!IQEG;9.Q4<T2*1Z$@+)0$TV\VRAZ1$3#78QL
PT[T"ZMX1!XINI[6/-U!2^/G\'^S;U*;OTO*70]=N3BLUBA/D[0H*$['P+Y"Q%PNR
P@Q1T_M%Y><XO ;4_5._V62OZJQYH?4G!Y*K?,\W+[:R)4<>_S+OO<43E-:+$]9.W
PEN#,\GV"KUB.G5'Q1)N[]L<&]#GY+Y%/@<E%J$?W^]WPQTEZ.K\T+:FVM?9!>,])
P@!<B$&*W0K N(XV1BXVD/5KVCEM<2^K5/T11!LO@_$%#ZD>;MD_&.SY[I;2&=Q*Y
PAD9XL#&%.7C+[0IAP>"-+:Z3)9F*^3O5H5>)VZ7H>D)BT0_PD/'XO!GM9W5>G:-=
P.4(5 U#UTK-BJ.>TGG.3T[MR:N-]ZOY%@:+Y'<R?-4<]W?V#E)2-XFMG^?-%XOU_
P8JZ"'WA+8?EZ8DI7PY,R>5>-0[ 6IJ7V^(N)$KP$S!&$CZF:JRS["7=\7JSN2?G[
P4C0LVFB_F/JWEQMCE1V/-& (_Y>A*'^PH0+KWIQ4[3/;L3_62)-5I]\SZ:?78K-?
PCB6;RIN9NEEYD[.XG<NX"KXB""D.@SKD0"Q1 2;FPS*.*Q((ZV\ _"E!)V%E<_]%
P^+^Y)IN^;R>;D*O]*.<6?<J_]'_&S.8 @)]@F;%Y8R("?U5#!!U-A 32^-5AB7>(
P?I2)2H9S+!Q+(C\O(43-364_2JI1;W?$\(I]1SWL[?P5%'0*AUU=85'8>"1H=O,G
P(V2O J:)K&DUKZV]&HZ=@UYB,G/UBU4QH*GXG&[:SH0?QFLL-2VI D,7N83$/R?W
PKFHT]:W B6#_X3&WL7I,B0'<#P]#8=(U- V6X6>>Z3-O>6Q@['#6F\/WBS6%W1_+
P34= 3$?559/ /H,"5?2[/W6@''(LB@PG:YRD[*(/&U-RK[/#2[58WR[@"3K(P]93
P.$^9L5JRZ@;;HAHSM,80PF0;/A802HD,GRN\.H_L37SO@-"4E#4%R?6_?P&0WS\$
P'A\=1/&9#6R]K)\,70PNFS)1FWY[T=31/8^EI.P.IN^V\&%B+N 6Q(86H0!*+R1I
PL\MJ/"#01+:]ZQ[-:E58+3/8Q!!%,B(M3M8M>.Y[T]>S(5=%UN^!CCS6B@6?[W]Y
PANF+,^U$E_!*GCBY6=,&>5?2J-?2!HJHF6Q'R')J^F^K^D[)_*,4F\,4\&"7=B&(
PJQH'M.K/,H$WO50086^,7?"K$,BWRPN>%> #B"TY.*SA:[M&D3/DC!I\0 W*@U+<
P> SXM36 3D-Q;$):0H_ J4)Q>C(1F=/-,V%=W1[T'?=(1DG#,,<.:=6X2]Q<_[L]
PRQ$, W(8HL(,% /A"O*].X(X\(6:8DA240X<%?=D%%.Y8.*U,>X*6RG5FLC:J-,:
P/Y*DABD:-@GS\XF^1_R3RH*@DB_]O!<!IOP6V866F+B$_)FU=9K3\,)S1LI<^U1(
PE-"X-F+OJ[,.!ENP/#63'7['/=XZ4A'_2.5!249ZRL]2O O/(6K6AR8U4Y#T>2U#
P%+?=TR,O^;Z8'(=+JO#>1 OCJ&.B$-MX^O<_=PYW,'E"-:%YI5[QR^.'<22X5O<]
PZ_\Z)2N;0?XUBU/S-F//[/T6,U_033)B8U#6*;]"GF/VQ'_'30JF?#8#<JCVQ%XX
PTH7@I88=^$V]B? "9T*\L9HY;D<X6G4W9*8T3])-4K?0O+'?>X',%&Y]G40$(0FA
P.^>T*J[X#%6W31$<GF(>)PWT6YD>[K5?QA ,9AI4#:_^^(IJ'TF=XT*A>6Z)X-/;
P:E]-J<>Y^" HT/AF1'((@"G@17.SZ*O+OA6)2T:&)02^%9>H<'GLOXED^"!&_%W,
PPXZNJ$$@T!)4+2A1-I-(K0\J]N/@5R) ZA]5@45*,FN>,A P_>WX#/P[ ,)9QZK\
PCL]5;R*;'7=S7-W$R%*GRD^$]SER%_O:^R<J581GZ0( ELJ8"[#%/___YQJ?CVGN
P@(H:8 K(DO3?]/S/OX%G ZBS4"W[F6::G*W'&&I^?T3>@OPEN3/JP/0"BLV+ 5F#
PSMIV8.LE_LV+I^\>HZ% 9^_"W^AD LA5 " NT3U1W"]OX-\H5"\RYA**_,]V9HY>
P!Q07[,ID9[5'U.6?+7'O^&2]6R1%(']@X=R6U5R&-;OS%+]]@T-+U2J;ZAY[<=+3
P&G,%:JW12B5"LW?9RF#^:0(F1WH%:WYGD_ BN9*5J9'J_),('O/5/+R1KC'6^S"C
P4_O]-'&.,[1P_QCQW3EL(--SN,&"U<.ZM@T!V=^%3LYU:,"/YK1W_:7$GUCZ#S%2
P<,MMS\II_WWZQ+T 59)^]/":9J[YW235-5/R9E*E,,4/=MK_/TSZP/4)^(@];O=#
P/OC@@S1#%"*FX+DFN%G).DM=MPQ39Y(]^ "1@YHD\S98%?F-5BOW[64P":/, [(\
P4LVM>I=IBJ"Q#WF@EF(MZ*9T_+F8*CK?-IJ%$A3A?^C!$CG>#B3HFB0!%Z$^?SC-
PBD2XG_C<T;Q9*TDIEG[6B#9X>@TXIQ/RQ,T4J<T-QF<W#LO!= Q8'CYDX)#KT-_O
PXJ&)BPM&GI?/'K6)T)SUK3]EX2YY<G0Z7L=6O#'.7!*@(7,>_L"F+U3-IZS6HFVM
PA*$6X(,2?[)(Q-7KCW7(@/;(LK@VRRJ$XX3@[F'B<*X<EDXTX?:O$_CN8%_"\LEC
PMGIA;90P2W)I2_PN6Y07JP>7\S#-5(@5-&2C0!1<2%H@#U9(W*VM)BC LIM9F62)
P6T>4)@+)2>>PD2$5I)9C %=W+!ILF6-V^B""<OZ7OQ5 8.,1!Y=S$P/V%$A19:N1
PFP#>I4T75<^E\5+0B/"TZ+^(\[*TWKG8=<W+:W2V[T2]16(&\-F/#TOFO/J=1)/7
P6<^7E:*2)&*ZIG'/O(B,SIUK])NBD.@+".V4%>T@L%M>F(CB%^"<>1-"M#CXFD))
P0P!(B"7._VPS^_\3+3AAW5;$:K(#4>FG?%I6:JA*G$Y(121#?9]XW6M</O)58\/W
P[=9HE8?9!VU$$WDXP*/>=(N\Z&HH<K&_N^"TPBTA7W#-*J3B20.)+;^!BCY#H%S+
PO7>,[Q?/!14,R@.,191$OBFA:6 . 0\V91S%TO07NMV^KQC"J5(F"5\/$E&-")[*
P'_>.46#I]W1DK&=B( ^PV>(#'XYKMYJN\X3O LF4\\H0QQN"YW;C\^*BZ:>L/GA]
PE5K6#Z#<IF807EP5Q#XFS'Y=DTU #FF4$84..2U=*CE_W;L*>3ZV/+98D-P_M/*:
PD7YU1M$/GB.G70KC@%AH&,^/[1&I()IM.;?1UZ_VYA]89;) F*6F<7;S,9K "MRN
P):<13D _D;WM9,,^2J.1B@Z51D(:(TFDJJ#PYK5_M<-6'3_-MR![;YQSIW=-'<-D
PB;TNCH3L(T-_(DF]'@1+9V'G/@N&)?1SE)3HYEN_"B'Q$NYW&IO=G5&BM1:E)8HA
P>OPO18J!/^#-K1[I>&?5043Y+=HSBQ9F\WB,86B,DN%Q+8;72_;[$]BE>,R9GRFF
P\RC4<:;L'CF()9Q.8)=*84%;@FS8.W2U*>?#+]NQ*P&RAM!,:$;M$[9'6,P%?/FU
PX2'5U=E8J]DYTI'(+Z[0?<[AP$0(= _>S47%U5G-HK,#O89%;7F.;!#3B\$LO$*S
P.^>1L6::!SUG&Y>=%EI5-PA3I7UD_1@9:)IFMHBFGNWL==[4E%2ZX919)$AS5LCH
PT++$_Z,3/2@N+\) E95Q915I3_ ,J^J*^9_8Z8PU/5^X*MUZ2B!*8-F3L5@8BT*-
P]-G0TQHD&0@=(E"MMG%*F^/ KXN:+TQ7\69*K*QI4_@HXOZ3=J8BJ_.:5%46YR34
PH955"FS]/;]LBU1#)/_W&;[=7W3%I+D,.V!:^DZI.$CU8;1BW'OACJ]3?"B2EP]=
P LD)Y6["R=7>V_TQ*=C 2AT6&FHM%E(:K90V,#.MDL*6*2;(0,]"]-'7>-FN5:CK
P'12:4Z()/9@WLGYXF$@YQS!V4GI:VJ1>O?X[9*^1PC+.WQT2R=P"/U&6KH?;3$V"
P8,V.'%9QR(#L\]>,,JIG")GT%L<EP6!WG!T=T>78].-F\2?4ILUD>K54ZZ_4(2I=
P#5#<\L[ED13BHQ\KC4,Y-EK/7[B*(MX/D':'6;!\^%H5FNQTXCKD^W(#L*PC!WAX
P()#X8)[C,#.8E6& 4F17H^](-,*<&&@?""<3"'FO8U[.E;B53R'T_:']/7.>GOXZ
P13I3Q=SA*F*<79RZ>-@3U72][+@[GKE0&R15H&SSO1DC* B#(3N:*( QG^Z2PP;H
PY'EU7$![03W471O80PE)+!EC8*NDC&/?.83I$.:=\LPK=>EBM5HVA]RC@[M#C\H[
P<I,=9/< G9<)TZ<AJY,'3;?-1!PT1$6BBC"D?GC^J?KH:V83O/#B'7R<?,M-\*++
P\3OL MNJ4>>NZJ%5:X0MGCSK\(X\3@_T%%$S%\O',-[\=-%218&G"_,T[V*"1L-\
P( ]79<"*$&6XZ<2 L&F#;#9!O$=\GJK%IT&M@:OE?[F#KN87H=H/Y_IPQ@<&7V3C
P\<R7OWSS 0(FF>_:SMX$<7N%#SFU@68&7@0IC4^'PC\_"R:L:/4(H4L..=OQ?%([
PXOH';;)6"0_6>,$-].->M\$>.=)?G[TBRG>HKITQ#$63220K1ZQ936=U +SU24E:
PMV#&Q3[O<]+B,NJQ3B9J,]_WC:RS^L(]DZ1.:Z3+Y!:\$S"GM 7?OY<+ XV- HT$
P$DT(EX<VPC'Y((H@O(_CYGP%YCR!^I!JN4^,5U3#5JC2C54HA6Y(1<2UQ=2HO8\B
PA+UQ3'$B.5G< U7%R@<*J!@/J'+9A@:[$&L\%;A)@_N?!+?LFD$3[?9WH\>B%W37
P@B;/ H(A]>3YX'7MH57VA%+I2\LL$CO=[*/=*NH.,\0[LIIF=^8+(1,QN)^3J/+S
PXT=WG2GPB\F$8 *3ODH#3[(9'0(P7C2WQ<U/Z4=24^+MX:H\U/MW[5<(:@&U;6(Y
P745O4@BU;-ISSE8G*K^FR 2D H13\MV!:<+:8"(0+]S'A>!?CQ?]M<#J5ZHX2D2D
P!QZJ% _SW-ZA?0O6^TT&RFA+\VA<.[]KT)&4V"@;"G'G(*B8:P+U?*5N'7_EZ\[E
P8R-:08E 8Q5 @(#)#&EA]*9@6'S@]+%*1.WK1*EY?U^&UQ)<L1S'8)KZ*VQ\-&O%
PY[J/-GQ4_%CRXVCWV6X)FK[&[D3ARMIP6WPD@>;,#Y&> G7+?[26 FK6A!RH'T[5
P&;Q^%73]V[2$DH&*PH33D7:4=ZJ3]N@Z9+5 JPRQ/[(>R$]>EV*$&(/"S+Q5NAP'
P"5JM:-R?H_5ZT)N<JV<= ^/VBM11X%2O<#.",HEAA(GA#T4L0X)R[V,8A2*8[ )_
PTK%185K?/I_O'WUS5C'-D8J^UOE,##KY <77+%.Y:>U(C/M<9Z/RZD5_DN>+H5? 
PAOKO>],+W588W;6)VSB7(HQMAR%@.,3]W<#N3MLD/.9%BX0X8BR:51N=I_D)]%I,
P7_UM/" Z@C&1!\4#+7&N&9?/?1<@6[4*\ LEY $<\/R/$EB1Q<.MPT?1$BI1[6[S
P$9NFR([0S9O_7$ZYK#!F5,7ZC]X=N1]EDO[==L\XY H2W+7#7^$]UET#( W>MY^&
P39N8$=QS 7@=UT8_@3K,N[ I ??SIFHS-([1V@N=(VP(:E]3,]TB([>P@_B7R;C4
P=GI=F5_&G6M8U=54CL9"NR"5\US>"']QE5NE E@*IX.$/4\CX8= <!&J>N)ZF=@5
P+JXP7:T<#SSHEBBX4M4KG(D'K5N%*4NMJM\MRQ>O<C?1>"9@A4Q/ABWDQDP13[C1
PHOG.),(2E;+7H:Z]<ELYC#*?*CP&X=PF#_4@(J=5S+L+OK&AZ"!4K+<HVE-\97]O
PV]T>?)OT=J0XBI/X_O;Z2MQD&%?R(TRE%::'H*0PFE(1Y-9/:X?G#]JT']' F6=^
P9[FZFP_7"_-*P?C8!ZL;+FV=]W6W.\ZPYTG29CD_UXPGP:\72C&.@XU5;UV((G:5
P:]1'<$N,$;/K\[=>VK2SAM<J6W&$50>B-%D;.(2-VOB@4^RE4\=DY'=@((:J@ >#
P_NIAG>'P^9^X6*<Q67T0>"5,^ FF_*+;BI!U??EOY347MNM34?>_-^R=A*8W\*VA
P7%9R5%P9J:-W.4R5P'G/_=]>VB2(#5Y.)S30S &2]&B!7QJHNO"=&J/;I+5J2%%.
P4)=7@#.YEQ(@Q+"BU "8( .Q&SUD8#JH;[:_:=4>TA6%/*"5Z)JVH_"*-!$\@5;$
P*YC&$8S8QT*BEB-N@\W,%/=+-2XFIE2!,OCX@<-VN"(@/=$C+;&U[DX  BJ(OLBJ
PI_AZ+UD>5O':JKATV=' ;&$U.J>EWM:Y) Y[ P#,9SF1AM5,;9%+"@" D^"'PD-!
P6!R:@$N5WG9V4$SE%F.,2Z[O=<@6V!D9Z\3Z#Z6^%=]J*4?$:B-F<MZD3>2-)$B0
P9NO,$FW^ AU.EA3WD;)2FZ.H^#$5NS<#1.X&T!CL=/__!M-PJ%>Z\*5+,!NNP0"1
PE9MSK*FRAE2L/3MV%QPB%MU\J!V-794#59VXE)B$(U'_.P;9G9VFG:]*S$0;!AR3
PF)8H!<A4:9&(JQ)]>T)'$)W9R/1=)2*[ NY_-IPQ*0L1!5%7\A \^"UV#:14!F:V
PJDZLM4@A,8[HA#D_#LQXWOB&D<!'C%+JDR,ANYQ&K#ZZ'U*Y'PU/MXQ^2F!<^(B]
P?J-R,2403=PR05I;T5)KHG6BW!E&8?9'LKCL%X[.(ZV93&[LD9Z'QRC\?@*2!DY3
P,##F>%0!P+KK[_4DI/L&.,3M$"*XTQB:I$T8;T:7.7OE@WU)AAV/[OWHX#K*]JW^
PZ6[S\6'/^.)2#*#]TI[FP9$,##3%#WX43*;_@CG0KVO*=%+ @K]]RH71UOP]=J6G
P6M\QTWD7/5&.;FPIIU2;Q*?.@K>#J!GEBTS<[-L)1<R:L(/K1OM1H@Q_(3(9$OY$
P FSLVQ.:V(B?<\'3V9U#=>(Y/C!L7%2Z:-FJ*RP3PJX-P&6SQ^\E:#"1<$W.;Z;D
PL(Z^_E W*6H5TUV3[?_U? E!Q?./6K>3L=+HJT<FTD+^ Y?DZRE(> ^/)<4TC7ST
P5(7'.RA"JGR[9E<UAM&^E&^,IJL&YJ'Z;,Y1U?:V<-Q2A$&&BR*.#>_[1 _I9?CB
P.^S:B8K_559(7;/-NVPNRJ6:X\'U:N'$E#/]GSL''G5)/) +\$S"M#&RQ#!8KW?+
P\X0=8DC!MIKXCTJ\9OT1$8FSG@>1H"5!\R)CTS^@FG(F(8473G 3P:T8,R7$'PV\
PW>8]<ZV1V2O9:>5GBQ23FN=O!QWXX/6CGVB++\WO2?C#ZL;.O%'D+7K>7")PKW_4
P5O_,J2](P!MQ&\56UJPP]&C"Y\L<WQ; %J]SY(PW&0P I @3O1<EH<C-^PONE8VP
P&-)?IF-(DTU55U%WWG;.'#5EB[4>^*+2C8_^CM,)13%8WJP03HBQ?T4!+U%"*<AH
P;=(>\@7CU,6@85MU']#^I_F@46>S7\>"C,Z*0POY74^3T)9YTF7@K5X@<RQ]6!4G
PR&%85#WNJO02A_IQB2[*M'__:(G>,,02@C'FP %SCC?\:RW7H6VNLN-J*?2U1EI'
PK5+*N(_ AUTMB"@+VXM/&4M"&RP<>\%YB22"H^3M@P.'"7_]VNH>.F7LZ+N64P$6
PG8)@)RQ$\AN]6R1;Q'S 40#"I8*5<D0+,ZC)V2L]41_ULIN,#2RI,QH51A7$=UZ_
P-Q'[V!S(ZFCLF1$WT$)$;-V51WQ$:G[VBCDASI+'/&%LSTU[$[/WS&B9C)T@#8EM
PBY0/W(L+4I9'Q=6#X%CP CAO2ZO5/P )"2G9 HT7B*VZ-FT<TLI>E%%'<7:H@#'(
PT\4H-1,"/MGEO W4> I5CK=6!N#L=BDH*&1PP_'9)@!@^#*#J^8E 9"2ACJ-I=/Q
P1-*!,)>\T0 7GCJD/;3?)=1&]-G&6KC>O463%I<D.E0Q%/+*RIB'+0?],Y)XK"J5
PPV&PE74; (=3AN6FFU:0I?@<K\&]&6G8WO3EM,]%S@@051"-"<48+&(*W].@/VHK
P:5Y/QUK+WI+O1TZ/8ADK>42K2I[O%X^F"BD[A&!S@_LNQE0'V@S":&NA "C) ,\2
PDH1"6<&E^]&#2#6T3OKT]4.]7N0;7SZ6X&J1-8N6XF-H *_5:PD/GH'\5OB0Y: =
P8Z+86Y85?\L<8R$4AR)AU.RY;0_HS#27*^]!A@O-.HSKM!H#]J91]5!15#,?$G0J
PL@2Q1!_*R#=5Q&_Z!:".BB!&O;-&*G^(;IQ7*#*^&V SK *>0$7$9D VO*>EH\3E
PH<E&O9R-<#0515/(;?CJ\_.0%:D7:J<4F_^2#\7;.!% T%E;*YS09U1=IUE!.=J=
PL3<R5'\P%7N#'D'6=3/;,KR58!)Y>,Z@YBPLKOI1:FQ""HZ &*87EH?UX"G$SX7"
P@98?P]^:QP)#M^PTNO[X>/7?3M+6?G-7LH#Y<-&Z7KLY*-#=FMMKE:@;=^.9VC;E
P #PS542-8Z$1$TPE02X%9)3R(9Q@N43_*?PSW<8='*]DPT,I\XWM/ITYEFQ'WYG]
P!=W(/OLK5X<<9?HB(F.$8;DN6T;YI>ZN?0$6BT6@3I1RNH=)7*H7%F)P>&SG]Y[I
P%D%QW-?L31 G#.78[S^TB4D:M)>44##8O05O@WW(E4;$V"'LK  (51M*$,N26_4W
P,D[R"1BM;I("@OL%EGNWYA+1+Q=?K"2_3$FX*DH?Y<G.?T13Y%K0(MUJ1BYRAQ+*
P$XJHA7)=D$,OKLF#F0IL#%&6[Y;O[Z.-5=%QL#:)9/E- TPN!H\-;">(^O!-9UJR
P@VCRP+@_2=8_E_I#IA(ZS6SE=,7 G>4UJ$TPQS\/Z/[6%\I?]_ 2*O=-.N_@R(N/
P1D?%Y@NF_=5*.#^29.E;B8;0(+3K]%5N_2&3UAB(>S.6Y6-JS3TS*PN/+NUIQY!X
P<#H1]-Y2>EVM-#"QL,S1Q0K$W%@( =HRKKEYG62]?82%L_74@]_%L84E@U00Q 9:
P<I$NL!\C74':XB?.3!&'(+&F<RZVU??G=6RSW)%2$D]!4C-/RZ'K&XT$7.G'7XR,
P.MMSY"2VZK:IS*&GW+DG?\;RP!>D7J&C6OWJ)BD,WUX*M(VY:Y=H=PE:80(8G-0\
PWFK$GGC2N@$U]QU^>O"G0+]HD^K5*@R41RMKKWC9F<QJ-U<'%BXJUGKHYQ($E6E$
PU$.J&#?-X-50:UV0;5*/Q8)17N^LJ&LZ6#.NE^#''#X*,H*DSIS]2=T3WA#5<MY]
P^4#D1JLD25->=C/NNUJH;%+P87J)WKW&#.,!-X$,0W-!!"FXX1E2[0.++_"(Q^5;
P#WA;03R*4#'9/=86\RN(@1P<:MD;+-.)W5TO+ _34+V$*6K>*<%F[59E7'R84P=G
PD2M(4WALZH4MB,NZU^3<#6K&@-Z:L%5^H#YZ.EFI/W\S^,C P8];'_IR1XU0NSDC
PXKMS41"DJ 7K-L>3BZC)HI99L(!*\2=[#D]_,,H&)XV[#@[<N,@KZ2*4=0^X/'P7
P%%CC9EX8-G(9]-BCY62T&"F'$,BA?1$OLQ1#+35%9R^^U2D=1G#$*3GJM&3$KS#G
P2+)D"XC[U/H6#%/R )D2[_B+8QP_L0B.)TWMR2>YB5]:F[DP2X#F&@\6M;'+I4RR
PHWDG&#MI.LG#@HI5F! II7HUC1OZ?0US'RVYXM\O-&;1?NS ^'N48>XP"VV#!= [
PJCN#?E H2$3#]C,^C--0C)\5N.-SY73CV(RGJ-/??UDM/,V,Z0>:7!>?@7;AY+>4
PX)"(UYU]X#F@,$=X:,#:=)F3UP%.&W&9%Y_%*P&I*2'J>P470-!H4,_\)'? X>(O
P]DQ>USA0Z<-D$:_J4UQ-!E7EO[DY7K&O51!!@GL[/CE'XAS)DV(?T$FA#Y ^)V!K
PS:MJ5&CT<>!KN$P6JRP))B%&\0S73K63*@Z]59-PVQI-PC"<_JS++073C1$=00QL
P0$U.G/71SC<<7S_;""31.I2:R,TC!8G8M\Q5O< .]Z%F&BQ<XD\MBFD=C\GWTD1$
P<'W+EOEW!1G 6H\ *IY])4! .%4"SJ@AG77IZ#GH/R 9WP]55P2@EXNYU"SPI)!P
PL+/!S(DF8$<P[93-U/54HQ6/GDR4#]I4QN(V0)W6<-Q.M!8&$[ M+TVV?HI-HBW#
P^J!$*+4@J:8WM$.:$;8(C<D6-0Q+0(=;)Y-&*8B.12[/GP:/N)%"&U@$NEQVZD#2
PD4N5-6)6I^1$#*%-$XI9J6(%*\TB9RYXF$/)-:J8#(7PF]4 )?.5!'[AR_J';F1P
P:= &@7@:O;75PN^XA9.3BSBMSH[B"D^JV)."]#1K;PC%"U9EK :1L4A;;A@219D>
P5/X3I&&BJ-# [\[QQ ?5N>!E[H+*;S'>;4*0)=8>='YL8'T-6?!;,/">B9OI46<G
PKN45D,Q G\^01<1V TKU%S_#Q^OM H'W?[2!6_? H-CA?..L*D6N?LQ:%5!"KD)T
PL^:.63Y\*I(P7D8[2_;25Z' 'QKW#GE>1]4!TLYKG@<4=*>@.$2V.*B(;:]&6?%T
P+';! I*D,B$G?CA*L464_- <Y%8NVNT7]QN3[=8.J2Y>ZC6QW);=D#EV3^C$FH&?
P_ M+C5E:.T 51^L/.:E4FE,4>K4*?OT871_@L&$=>-V.[ Z [XPSQY,:Q.KZT:N5
P0G3ZN?YVC5Y-:CW#VIJ+?*4]B?H24*,R*T@<O5P '-C1\J2E1TO]:^+4RY+E:-GC
PWWDXY,1+#N=-&XB!59;N]:T_D3C&CI$U)#^*5J]1RKU1I$MT_)M I66F<2@ 7@, 
PI6K,#^<ZT"(&O>Z4/$GVG_B=;5\%.MT;H 5L !N@A"B")(LNU<_VI\H%Y!B@#4^L
P:IRN#M<;LU&?F<W1OGDRTE=:TRE';CM#[L#^$Y0!(!><D<7?$3X 0@&=JC!Y:1_T
PY60[QK#&_!QLEB4..VG7<1_;.JPW,C?,?RR%&B[@",L1W2! C6*UG* DE^QYZ]6O
P<"LS-CI-4';.+$']?%Y\%O1O1G:',=F:K]W^J"KC#P,%CO=7<(:&"T'/Z;+K-N/*
PGZ")0LXKB<&H46.5*WL/!)7H0>O=*= [[U?1Y%O70FU71'=22=6;8>'5&L=\IIYM
P6#16'*W<]QC4C N<(T[+1^6/9P4HHA]83UBE]WG0#X11= B3#P"T3H^1W/YG4B82
P[%$I?&#'W9^INP,/I*:^3$9HCJ-<K.U,];_=A1/UU_,U<0<:3\*1F+EIS'9\5<YI
PYY=KZP-GC"*,Z1;SV'&[>@T?/#.2K=8K"3'01\E"G4U(^V/Q!Y@0Y!<EQ/VI!U:5
P[."$0)#8-AHZV5?/^]O,EB&\A= "ZH3*4HXQ< P6?K%<K[TR)%B(T#"J-'0D[V&2
P#?5]C$!PG$*KGO#P:)K %)YQAR'6T!.?]"3QFN(A%%RE.TND3X8;<]^M!K*YZ$QX
PXJ;LS-X\LNS9I-5TL^@T<TIWN' +7U/YWMQ<I\=XPM0A5@CQBP_6^OG4Q FM232]
PLP(]8 #I'V#[PJ@VK*NQ/0=6$8@^92?E:46-S5?GCA@(:PPIM?+(HHB-OWO,IY_>
PU(/_6>0H$RJQN%J,PK5.Q.=!0@&#BP7S1/S#,*;-/:4*1UA&JUFUL0#6A!TV*PH\
P1DS[H!8W6T,:1)P!=I600C-2B?86RNI]&@<9DE:N"1?R)RNH8"^F(_V* HA2P"0G
P0Q+H,J6$U\SO4)AH*\H[-=J?:"=M-KC?@V0<9(CK 2+2E=.86N\43L;(95-+C.]W
PO)RS6:X4KPU%W()7#)[ANMRY4$Q.(<^W=H<OZ))F*'U1<4'':*%,/#K6!9]1*?1"
PLSD:[>\A?Y)JDMEV[T)HUE@?_8>)KFU"KA!>@KDO#*B&AN98)S,W'1NJBO<!+-ND
P$BHZYM.-'RH./(8!EE<Y/_*SSC^J@RE^OZ/.%!KYE\=74S;P=U[AW'@8APCAW.[G
PQ>#<8Y6LQ=F$^%".+^"#F/CX#^=<86T($GNF96:S)RGMW?3IO.H^7M1_;3H;+X>'
P61CO!62*GL?!<FII?C$"W.M+W^N@EI)8 \KYS\(V2&=%2@RX$^)9:\TMPJU' MB 
P>TC%F5?_ I2=S-WT!">Q_=0$5XI;K]:CZ,.BR<HCM[2GRVF:;6S8UG+94Z$J:$ B
PC.IA=;C[%$?4CR52[Z'EF.L\\Q%5$67548D%IZ-V0N]B(>#_FA%J!QFPD+]%JLGG
P2L53&O'=7G\EM>X2#DAO;2*4B2._'/&:58;M[]/?%-LX:.B:?VN>ZJD^9&@IUD9B
P<9M>^=A@;K$7AI-FVQ*H3OC3[#Z(7D1J!-=.]0P6,[]WYE'_2)U"56'B[X]*1HAC
P,2[>$-B*(W$49F?BO9B!NQ7A1I;),O0X5MEONBB4/3L4:\2(1BJP[X1@SM>EAF-S
P2IVN.Y.2>=@G]B7QK]78%SWEH1/WL(Y)T(:6K'+?),-(]<4$&>':0*&>_SPO?M8W
P,-;_]C<3PECW<+8N6#NZ*2 <C1E"<-&G&)X=OG.D:(5[H/^H8+>;J2'EJK2Q+=0$
P64T.V+ V-NB'.$M(,[#X$DR)VN 7'(]>P\BM6L'AWC%N+(8'6=12NDCDI!/,P^W!
PRR-=I4UQ/5SC;0]GMY\>:])N[6&N\G<LIND2DCRLR@0*%SR8V;S-_HL+M!$L"J*?
P=@?/<6($LX:B.QFSS,8)N#&.C@4NR(F %KQEN$XYWU)8G<]SR.>Z&\Q\.&E(%G?H
PJA[5E-?XB ="$%H<31O,2C>74[-:J:M(;212*6 5$558+SAW!AC07 Y=K"'T2PF/
PI\##H/_ %TLAB$RE9^IGW1(O^:-PVU/.-$H]+9.\.K>I,'?#4"IA[PHI@P-W\D>%
P\%;6I+&HWIXQ7G'\%C6'U%@##=V]XZC"*6=/3V/WK^[YL&RL(+\-U)4HW[ _8].N
P4\/;K1 G"+5PC<FA #01!.S2<3(RN0%-]*6+'AHN3<Z&@/DJ\PG]LVM*\S*JR7JH
P9';EXSZ[@O@BOX"WP<FG!:QN2'4]?OB62T@MI._M.IN$6SX&TN!VBK__12ME.5P$
P0Y+@%SFL@@M^C]-MU"C;EKT,*E+;,>6(A[$E:F6:5 4QOO&R>#/Q0A7"SK8[Z!]N
P&F[/V6MTNCZWI,M6UXQEYLQ8\OC)L\[\5\:"]+:FJ!06: /Y_<FE00TGJ<G3:_>V
PG6DKF*%>8OJKXB<_S>+-(L<5QZ0WH9M>SW!H^$$G+6=D*H(ZB8Q[_/58Y>_N!5M;
P 420EW?+L%YN?@/PG1='?1_QU+9<;H [%"]^W-Q7:.;3R7L+']Q0M[51HKDX4C")
P&>^"%#'%> N?&<U=""0^DOP9UT!S>PXK6OMB):BZ-JQ+U8U<;"05$;H6>J='2R0[
PGZ+2%_%'])XF=S=,43I2OX@&[0X(NRCZ):62!?5W0Q1Z9S3#;NG! T(A<=BLW!FR
PY:*(N5I=M11/Q2CL(->.^FQ\Z2A9JL'7 #H]:"^>X^PFFUK7#Z&N_+N*U"O+NXYS
P7 8GC*X/M23S*S[!#BS*.9@BSE\F.;A"!SD]N$#:K[X 6_,#Y6+,L"<1*_^]5)YP
P;@JXN8T'=5;B4U4[L< @ID]PO+#'36B\:]]G2DB>N"$X8#PQ-*SHH+@>DDK457$?
P$:F:%K5,P<[]1CBU]M8\9*53_>A*P1=5%6^\\H7+JMT6-B56IC.YTZN578S6!@E@
PJ@5AQZ="'D*5@7B;D<)RT5"0*.-"K1?DH"']AY\ ;470/V/O+U! H[)SAG@GI+IU
P2<RAPD>962*8:C^)8(M@6'(_VYVYC\3XVQ[T!8/#@X8/S3W2^?%.U:S$O37 Z_A^
PQU2\E]BW9UYIKFQ'^U*M9M22+9>-"6UX:@_ GZYRR#1CUETW:ODNR/[ Y?5--:AO
PLM:%/7<^ET@.J1E9 KFA"N1'.])#PAR_E[L(Y(5GTO56NAIQ O-NMLC]%BS>H,6+
P"]/#A;I;@9>1NR4"YMW.],07TM:V^<?\O+3NP%%+AQ:G"!YCQ:'K"2%AN13%*AL 
P-A<T79!QL-+"<T+;^AN%]R^8.=N%"I7<#@9C,LNJB^0<R>KS5RT3)2#1T%'=PMRS
P8/FCA& 0W$9SF:;J^;HJ9NI)DW64^T5!$0DR4@KK:JX2%GFUG /=QY"J*1XU32,A
P\V+I\!I3X>)#1A_-@=/)?EIG>>  R"AAJPN6 5\]*)VJC/C8LNU% 4 /]GHB?Q]5
PTYY/;W2'@0K">#K*0;_'YKRZ-8&E)!2\QHIO\SF8+*N]T[4ZW_QB2<X7T\"*(/'N
P U I/WJ5JB'+?K\F:-C;.!RVC1@P\]G/'/\U_A.Z#E$W,$,AHRB=+4Y@.)"3653&
PADFAP@[^;OS@J@G?M/;D-A*@VZO(6$?,= 373H,4=W]92_K%Q$+W^N:$I+72/<8F
P_.U?T2K1%0X8(<VY408++Z2AJP9\'FQP?VT-7GWKF?,R&\\=9*!/W]%3?QF9+0D)
PF)_S<[:U?\NTF7^9B@+*BR>1!,+)+&JRO.M?WU(E#,8=86/#^8%W 8%.[RT??!=-
P1I%\2N>0X<0!3+6RGB)&%!'ZX3G2+F>''! W"X$-6M_3];$P5# P>8Y:,)3%Z$*<
P=(HK;T\@$2BJ :[S&_EX\X<TS$ST I]7CEG1I; *./G.3[B<@MMI)6R"O9Z%WH"<
PB#$,W=6!^M?;_1 /YT\+R[$\/BH6?@:0%Y'!UVV7+VXVRB<9:BDE)Y]J_X>8E%;]
P0,K<UKL<!(\3+AT*?.\/@V._8Y&%OUBA#-%2B9X\;ZIB+D6TFL/2L\#"DC,'F81<
PHY\BG67E$5OA@;>MT1U\?=(KH"1R]PA_Q,O;.G. 4AUY\O=DZ%(3."Q)+<@>"Y/7
PVT] O.QP0!X ][IP6!Q5)Q6'=ZT(#1UB=6GXPWWCG>IS*:O1YU7"(P#%S1?%8!(#
P1X,8[ [Z_I%+83V?W\OU>7#')%B>\ !-DT F$L&Q0,/DU7)O"\ $Y\_&),*'9>[+
P1^P&BDO! *RQQDQ2'D@2GD!"3..1>_:\!!^U29V7, !<1NE\^M9Z4P&C1_B/RUZP
P?KWD RZ(>Z>5)!]I^AX\M,O0P64SKQT$H-*EB*+:1Y#7Z4#P?!0%3%L2,O/^1QV"
P%D800FSW!?BC8.E<.7X.:\C^W9J*]>:&BO7-D.;R<28FD;L%WH&(-"&S0_?<:_YZ
PQ(TP=D@6'YS_P?[O4P5+Y4F BSB3]@'4W^L\R_*NAA+D"<,.*J'AX5NN(6C!+XP1
P,U^H9(_5 :(2*>Q.P4()L<&!OINPSWIEB<HL3^[_!1PP>[E[&.XH_PPV_ Q(T>,&
P&RP8AK'2%I9G-?XVJ%FMW^>JYG:D[ GGRL"^I=G13+J[T=,LY_ [C*4+Q[F+OY(=
P0;\^:?&X4YJDB5L$,@>4_W9$^D6>$ZY+&+LN%Y\,;58/X'HN2>T;,<E@&4 0>+$@
PY:FB\.@AK' JXL1>H=69/X:I93+8L_%;\')7I2.#!VV EIG(P&Y95V-,M$#;#K)6
P9FWOQP]\7J6=?]<B*OVT_#.420F:[@=FU^E@1$0Y+&+EJLS1R"2_K^A$N6M'"938
P%A5BM=9Q#3RSDMW748">>Z=&VU1!2&QLC*+I-99HXIYB$2?C[UV7E;2Y]/G?1>M8
PWA0';NX#G!2A S,FD)0V*514PO251Y4 JO^0O9O8/_:JJ0>UY($6RU/HAC-H>9:T
P)+NOB[AY>$QND TV)+D F *LU!+\. <)V;^3^B>\< <CD%D@A^=4EJ/'#)3@0FW7
P=IX876X$$)T= _S,PC?;Z](?_$$?#1);WXTIE<0')*PT2V")R\B!BT8GMZ&A/_] 
P,S223,^I!;]SE&$QR6MR^5[.>Q#Z:!GZ-LX.;K)E4#/8]7F)'-^=DK++9M:GF"@,
PZ-J;V*QW7)H_$MDOXV&WD/N2EE\/T,,?;0<"C S.X'7/J_Z7=:6C!='@C$78O..J
P2^O![DXOIFAJ,C5_6O25JVLMV[%NZ!M]3FKD^27UJ35P25>AW6?MK=C!GT0\MK9K
P*V=H"*[V1_;G&0A_TIDVY:A<*^0!^J-:!39<10"&])T41;!?S9/[^DE[87+)3F,T
PZ<""_]S1 +GKI/P%7*+P/DN0+4K5QG.X210#N6TG !.SW)#\&8PVP+2N51W8+CV6
P)=](LAC,NQQ#EFJKZ0=)*[D<S&^.[!AF''A"Z>9D6*E'=0M7[C-C/T?9KYNZ1F'5
PALNLW\A82=S9&^UM+'[-K*R>W'?N=1%ZLQ_ECT5P:NV4ALUCMG]B&+%ZD'/)K*D'
P,_-LT$>)X1=L3N<-<]\>-F\-F'CJU.JGHC)KW^?31O&0M<\5.?IT;E]X0793?80W
PE.OU6KG7U'K!UX(Y>L!%,W"XBQ2H5DS8HE(#3VUPU#(/$BU18-\O7TBO1ME2/T^O
P=Q_U+;RTQ&)G^;\4XCC7-/VX\9;\:C'.E;HZ*/" 4!))^G(+!%FIK6<Z-?H?L A$
PQP["!Q40FOMQH$[BTU8_7\IL;H<WZH0V.,^6(E1+QV4&N;*T'X+I9ZE?&3);KKS*
P3IJ AM ,#WU$<B$]&\Z[_GZ>)RFG81J+89C:NX&,Z])G52:K%,QX*97Z8>-3?&2>
PR[V%"?&)XS&'-@O-QW?:$;0QT0C:;!Q3(  +F[N<:Y#;81[2S*&);R8Q+0T;."IR
P"T%W:;^=PFD*=)]O0< ;4643>'G;(UC\*;#1O+9=<#4.INU&\FTEW8+>N^E'^19T
PY8GT8(11ZU$>KJG(+K9"X%<QDNI6/4LCG\!0O.@GGL,5%+45"'@6FJNK8M$.\DV@
P]\,O/.+A6 B:5"BOUM)MX_-)R9'QVF5T[\_!>/H72>3EM63O:!V<6W"T<S!D;-M0
P8RAK9T: XQ<U?7HK:4S9.NZR35N0U.V6)@E]S:#13H_L;:,7+E&Q<7I)A,RF_XN.
P#^:;>T%-KN>X.@T.R,$E_TV,_)X/Y^>!0[+!1H=:3G^!!38=DO+=4%I,(X1-E;Q%
P&@& -;;?FQ#[I+[OTQW'5 \$FP*RQOM-$#\",F)EHBIK%CNX$8)DP:X-/ZY4"0^/
P3N )^W"6.[Z!]$4KJ,3JE:C"4EZ4/0Q0Q) "0XQ3VV[V,?S7B18V5X((Y;WT;[B 
PQ++G/@7BD4@;=:O==(>\#4E@-2;^AYQ"_*,OP4^"Q@@C2?%XE*SEABSU-.I=K@&)
PIY<742V*T.P?6'&CJUAI5\[5&+PTF126T9U@:O4Y);(X3'BMIR_XXFO+-]D6L67Y
P6>T65M#^CB^T=IZ9XU7PN ,"XVFFT;XF,\0GF_ D_B'SIS M3KWC/0XW^K2\A<+S
P.V;7-'S(##PJ]3L90#H1"<W$A5 1R.?1<:WZM "W,FP_3B#;&B>M= (.Q;4**,>:
PRQELQ%-D8V3NG!L#;5+\@/]')O*X0P?-6(>80 Y?$O#-!0+\_R.WM3N@ +.MX2C>
P>6 4+M7K."[T0V=0?HRVTM1%BBDD7Y\E01@X0ICA22Q(E[^;UN@\SH)E[A&=<*:7
P.K&9=)^JM,+ORK0Z0,%1N>]'Y6=G1]'%E[)_HEV!T8=&^LCX(D69SCC!>3=^X[JQ
PK;,=1@RPT;HPI"U&+%)?1K'ZS!F%0#:V$DN#^T2C1)BI@LE=).]5%[^-3_GY;H?"
P60"-1.MRN-;LN'0NQS(RC?28[/_[U,%Q]>=4@@>BYML=?Q)E5#:,>WE9T,V,R54K
P2;UVTYCRU._@IZ>M=]^>A)']SKO04.Y[M6:RB,(*)BCMHO\7N?KD->W37G)Y"L=!
PB[6G>-'E@\*Z-%K>'@[T1ON1N]^/!YEU91EI:3DS%/7IU'> R"T@7G'DC6?<H30K
P[DN1P%BX4U[?.R]?/&R:-@Z=SPIV:!D.7C*S*??5.?@6E?HX]@@?>\G7%<_X+#:8
PD%9(3JQ(N'"/(JBJ"3;>*>)L)L!.[7PB<=*=4-XO4K;H\.BJECHKD[!ZT#YGQXR+
P=NBCY=W?L,)(N!D7'5UB"%-J@GP\C I7>?RK51KCXX/'XGAXP- >5H'C]1A<@^7;
PS(+.H2&.(.H^94 ["PY/790!Z/7#Y)C;B]-D&[MR,HPSV,;+BH[IE&W$R>_C)"(N
P(T'(@M@*WA(.&OO[AS.+!/DMJ$0 C(#34-M9\]X:< I"2?5_1_=0Q">L/\_\&YE@
P)Z7@W_>SW["_T,V3[)GT(W$MC-TNV7"TO'?O"/&^IHEE'.03UP">V2==?55[;U;.
P?VJ/C5]:7-[F\G28[XXY_&^$%O19U\@9W[DZ$TP/,:1$;M2$&8XS.ZROB--O.F<7
P!4]X:KV9!>-]V-H(XR:[T3!5$QNMOGV<K$&2XF\269CMK6EKQ2CO79;;JP9Y7_22
PCZJF9VY ':A:4#=2QI08S:K0/,^X)L#>XQW[KEP.8J>J1-@F,Z[4;=@U9[1RU,T-
PQJYD8X"B'ZQ3AV"M]7?L9+22FN&-; @:>C[NN-60S +J(?0=SD37MP76F.(&AG[X
P''9OUALKT  O@V309)N"\)T_DCDOY.+(7SG+<$D#7AO"32U$]2>OH;^)9<FG-Q68
P&E[5LR ']A$?G!9'OWRR;Q*NFEL#\+"J6740L=8\@H2:8RZTI"TQT@4 ''^=B"E1
P&A0,9#<,8O(PD71%SYV@9AL)_0OQ C48T[:U>?T2!Z2':1)]E$,0^E7'=BUG'W4]
PY+<BAID.!709VS)7_BT!U2NJS4@KBTOK=YEXJZ\J"6B@=ARZ#*H'H&%?$B-3\#C=
PS.1&2:::ST$'/&JCJ-ZC"^$BGS_ZC^#=&[8%L7"RMY@UME]8DE>)Y8$T96W3%"K8
P^]%MR<#P3*USFFZLFUV2@WKH=@?QU"L'NH<$3;0MA]\]/FB0\JHNH,1>]EQ\XL-J
PL0EZ-=*EF+X,5?S$\:T$9M<>31D9(V'@7V'57ZTBHGM+D-?833GIK%R@ZT;5I:E9
P=E1?D^Q@*&B%S2Z>+"[*B,Y/=7TXU_O<4A]F05>36"I$+Z#LZC->[>S?[?-B7>D*
P&O[Q'VCU8HYT2"&"8L RJJ\&E:%VO;_@H=EE:)B2&<A7D';24+_X%!K <RFOC81Y
P5#2+?7,%#1@3C4[:UZ:3NVER9P W)4=\!":]-C:43VTVFE-M;;0=;3Y15IQU^C(B
P16()".$-,S1#>:L H\(I2O"S\^:+IIJ$D:3MZQ(;-) XOC)0O+;5*H:2)[8'HKH;
P[K_U=;E6[#M_/3!#2-$6#9.) 0DK$+!1K05T98'_#/LB>(#,_Q=9F'_,&*W.@K#_
PL4N"PA[+2'N8ODD4+DL0)<R2NAZ/*MEI!KE.U[BO?J&@NNJAA1?-P\$)@S5X![SJ
PU'TK,$ZY!&G8++%Z"+<$&340]:^4Q[+I:K__:IR^H4\1%[XD-WKY4U7\F .]5'U<
P]=(M_T9H!+$-J'T60+']=4Q>C$@05K7X3ALHT0R=P<PBM<N ZL3[A2V;25(9@T#J
P.<=5$E++F?,RT:CZ/U>,EBNTL[;GO_C7.LB%2]P,&D6!PK28+FM6[I8KWIW22LA5
P NYA^G3/M-3ITNIC8-U@.C;CIR&#)HM%JSA-B*220E&F(^">IBE;M]L\/V*>8KFJ
P@806S%&7?(F<1Z[\P?KE2/)WK[ONRB_9/$(9Q\M_#;[#B%B6&DOLI*#$)+";6RN/
PM%R&-=JN0&?O"SY\+W%:NL;-$S'4 =^WN XR>''V>P<NR '2[*^&_W62#BL;\4JM
PO_K?4EWJT6"MII,T*G;G[M*!<[OO3-Q5"Y&F8-/8ST0/6TEP%':8!Y)_1BH62LO+
P,0;S72;QDR=7JS1/W=S=H@5' ,E["X1A7,BOWPDA[:+$C..#3C./<Q>H0^UWS7=*
P#Q)WL?8)%#L,LXM@)$X5"HF["PYB:7O?$0H!G<SI+<'=1%Y<XK2IXR[C!6WZCJ:V
P2F[S/>%=Y!3=6& H4D!CCM.CIO^@3EWSWNKE6EHQ50FB?F2-]D^!Y[\(+4:6%_C:
PY6D]-NYVUGXDAM(?%H,BW<3%,Z>=$)TFHL=]K-$/N@CFU*_G_>["'SIK'%N?!Z-E
P,$]52?F704CYVI[('[8*F28U)=>T5J$G*J/#:U<V2I<OH*("FX/Y2QF5SL$"J!+$
PQ3YRBEEV2/G57+GY+D]2'Y&98N0J@G"OPMR6RM-4PSVB*/ 2-'(-QF<T:=!N*U?O
P$W*%E'*BQ&,=KHU%_-]G$Q#^@#?5? C"A]J#%^XOKNH^Q.":PYG=BB(]9*8Z!A9_
P80*&DOWZV']MC*.&GQY+>W7*MK2Q(!@$Y/?N>8QAGECM6U'7Q3L*@RJIWA%X%C7S
PMII0W?])_H)V_HUV!'P35+IF$;/XE9>#POH+\Q8&H1/@*+YEGU5^OU[GKAN-N9[4
PD+Y'/[+Z6A99$_AR)CX-E0$*-PL6J5<,.03B$E*OZ%XO5U$>IMHVYT" /"). U7/
P,\B1B2 &4YMC7[^E/L,\$\Z[/EUVU0D "8GZAL.0><V,]$TF",ZO6[V@*F@H-V,_
PTTI2%M'[<*IZ$9SY7*S00-MXZNJ\"#!"&BRYDL)SFBJ($;:$GJB$-I*[7ABE+.1N
PHT8*?8=R(S-7XAO2;&!Q7_),9;JY-,$-";>&=Y^Y^<*1Q[?"$))Y=?NXQJM6.I%]
PL<DG^)N+];_7.\H\9IU+X@_-M"'&NN$/$X<:2Q[^%21QU][W10D5J(D'[W%*&Z_+
P7A>KKK=**/!UD2NV*4ES^[LK+RD,4]5D2PPH;.R X'E5KZ9,'41U_*0D@M,1$'JP
P,_R/>)CXAEH/1E>%O:D8KF YEP."R/D8_\)<'Y-1IFT'+X46B?]*SY@L.,MO^(AE
P):.PZ;^2B#^Z]_P%%,;8=52V?$H"A.C9^E$THD/?]L&,O99>9,?@H0IDB+[NS;2K
P"@2!-KJ@&P''*H7:?;UJP@8T0/46<@Q"K%\H%)N2Y)EXW'!PN#-1M[L2Q7/+Y-1H
PF5#D\B@9C+[7QC":AOZ@]IL\+6]Y-7W^\@]8/YT_V8QX#\$I!!#2"<BS=:R?^"]K
PQ_CBB&H3PE6KT;69+K[L(5B9@0?'@/LV:/ ;FI+'_FGX74:0HD7K<\''BGX%PI2'
P?[X+<1$TTZ"$8[.;CJ:L3Y11@7Y E$RT4<+\VQ;%9\K'3)&N, NE,EAPYFYMX::)
PZ-ZO'D1?&;]U)T<<![X' UBBCD-818RY72,LU.*,:LD0#@1>>&"M_^ LRH 3M\.Z
P?7IG=S I0#@'/#&AYM)C*JG(S]\0#AF9R#NM?MXI&6B(Z ,J&9R#MGH/C"FB)'E0
P&3JI9$B,)LN8')OW+O673X/96*<D=Q58^" ACRL;:T_@O\[U",V'-^9!U#O/SD42
PRY$"-@?MBNJ(@^O.6,AA# W3:R9_*M*P?WLW>0+IFI.J9FQ_15>8A8;8'[KA_OLY
P)RAYH8@+7?0ZE2^M7Q8A=# CPTX)7LVV7R93U)'1)IE"TZ%F!:3X*"4AX,^9**4/
P#B0$@U ;XT6Z%J*(1W@%>6[)KP;4M*#Y1>O#W*G<JBZ6/D]S^M+*>[C&T>%;K,.7
P*T/)8Q*(!YWPV;]AX*$V(Q%2'+@5!?"./9*.(T-JB%5WM):AZE]A0G'8*=(&M&(D
PN$J.;H?OM!\#2%@TR$1???BVMZ<S>H5^LV5G<RL]D4[:?0*[<!!'BL_*\,!(JM<O
PN!['PP2"@U?6YC6@R!Y6Q9RZ\#4<E_OLOV&QFQTMXDVON07<)LH.+1NHZXDE:F6&
PT?UZ\O7L<ZF)$P&UNM\DZ8A06V1^1VFTQ:IQ92%!$@G:)N@VIOZH[;1>GK^)ZXRT
PPLAS<^?_[L@>9+2S3-12'PCDZ3*5:NDD+'8?-*'%1FXQU&\2M:>B7K7U2?H6SA"#
P>QMT8YU+M/7-:OV#/A@V(5_N?*\5T@WX:_RZ7?(/,[(P_&S!$\U0HD957&YUJWO"
P?>JI[?O1KK4?Q=/R]1,PZ=(D@QQ)G:MBPY/6#%/HW2N_6;2#WN) !%$>MXK+@O=*
P#5+D!K[29()U1\Q4B_IN76VCS=S?;.DR:LE&4;[%)\B="ZM7,B"H\A^_AYICR9^*
P'-/$A5@!)9U.0.>+5#W5HWH32&[NYC0!7P[K+-.S[37_=F.GC^H>+%W2F$BQ5PWE
PMVMXWV1<82/IRAJU-P&4FYG<#_\[[LK75V.HFOJLH9 ;)2(IHCI)C5$Q1#H9^-T<
P3HG)E UJ(">.&:?Q*706V(PH M)GKWA+ZT'Y*'2.:?N/X2S\(.-CL%B\.F>U4-9-
PU,BB"K#R:&%EJCPIY.9\1TBH11/,P8?9_9B?8._B1K.9O9.,=9FS05M?CY\OZ-@-
PCX1Q'L,142HS,P9NH/B27TKY9K5H!'B&0M$T>BGQMZ$,RP 8A9IY2E;SIOT/"SN1
P)$L$\.K.Q5WWR?!&WJ*LRK/:T=M.F".(4YB"8O;GO$$>Z )I%)]]9E[#;O)J,Q=A
P-=.$%+6]RD?8X"##'PA*!1$Q;@TA-=&TRY7(2^:S<,E?VX^6.$Q%0Y-4^QHIY&HK
PAT$'_Z"CZN=@YX$'^Q(_N/-:P@EL_5?6,-RT?8RI=<4-6]<82,;J&S;24XX6NWV5
P.!Y8?M][Z* !9T<!J*&-C$IUK>$ETG!5OFL<*%-)#] ]B%I##[+Z# I*CTP-N 0&
PI"";*[_L'@N4=T"NJL"5(:F B?-@] ;K11A7;3/,9BLQI!2K??&XHX+7)#:%?@6<
P%7[1*0MO7@LOZL@JC*, T ]24ML]7#95BKF#3NB.U\8;T53KI<'1>'WH@Y60A!7*
PP<D%V)M+<?6QJ$+-4>.>PK&N\NRZ>%C-F(::_S>VB0^< GF"_5#ZDX-?^ .17-/0
P@%I8((:<\FY",-E8'["R$_"X@:].L6]0L?@.BV9,*/W=3F=&WL 0^0?5T0XD\$RF
PIECP2*76L@"O=+X(G6TZNC = !7&I4P17?/]A) P9-QP:!$JG&. *5A3(TW8?%%7
PW(J#$^C0%$9C0G0[7L#'(S[HJ/L5_^:2,>!914.LUX,?AM,*(ICN<6*X(8Q\<^]-
P7I!7#>3,>Q(.ESJK-3$_'<;]%P(R =2\0R1RAH+(.!H1_A1Z8HSMIE**U-C#UO#\
P"%)+1>JGQ)-I[2+Z*?FMM^U?*_T/\"=M\)1V<JQ!T=@%C1'&>ED[%B!4.Z]K_VG=
PD7^KC9!IK#/(-'O@6W4\Z+'Q1XS, :!$!*D8E<EN=.#+3UL'6H+@#3V '0.]ZM]-
P[J(TG&4%V[Q!N"7R_G) V(YU<0L40P^SJ FG,GKHC(88M^P-O$T 0.<16_AD.R:.
PQ%%D?!\YPW1#>= (=I"91537C.DV,95AG! > M)9=BT&_BWLD!N_]\ ',#FS(#4^
PPZSH=B]4#J)K5E(9Q#O+*TRB$(WJIWW!?]R(BP8C')MZ.JX2FG,*V)!.;LY!,H8;
P&ILR/"PV/>X'<79%2H!D[UF::U&M0A<T<PD@$__;N>X'&E5+SBMBQ1\(M+6*:^ S
P6M*ZBX \A.9NW++NW#?'D)*"395C#*:[-!5\O:V2Z_&(P$;%N#6D,'GC73,R2XW2
P"A&/UPSW!3<*Z0'%^LQJ(+:2]U^>V&]:TZK5F:&/S1J"?5VZ,N/7F1I3D6+@)R8I
PP<VF;"T$]ZVY$SH9G) NCC<J8BA-6&#J9N#-YZ()XK0>L'(@E44W;Z(K=.B2<-,G
PVM%G9NU>]+'N:1/8TH4/%,?*AK@X3#.UHF#=(*]R8*<\OC]<4YU/U%PZSSG19;7*
P!?9@BH9"44*+0ZHG4AYU\(UW>9:1_0S*:MJB+ UYG2M/50WWG*_.AITU;@:FE]'!
PD-1(?TX:.QZ!I1Q/%;ZP434W/+^5(WKQ-T##*.CN)4?*[[H2.S7J.X6N66)'G*A\
P20?=V.N\DA,RM;@E390<&M-C8'8^P5P1,*K,L/;4&XQ5<RQ1 ZB=A(.H:>.]-XN2
P[-35=>1$YLAXRHT2/)1Q9/OTN^,H9+%BHC1$B8+ #):1CO?9[&'5,O+]TOZ/P0><
P7O'$6N:C=VU.Y.;NPQ[;EJUV%H/XL0]<J,>DH=TNFK'.TYOF#RJ[?X XP)BR* I&
P:%Z;U $:C2@D&+:-UFYI+V:]IB& 0N0&2MY".>8UKR*Q;IY:RQV=FB+=;*S*=,YI
P3$*.!=?;U3(>MXV =IFZX=KU&_6"S3KJ$6U&,*Z']?WV"!@E"?LN$"4SY'21.82G
PS&0381K&G?2VY*K,"@AW(MU*'3OA'E.Y++F(I.[;E.PH2=8M;KC9FB8V!#SNRF]X
P)#GI]OMX&LG(N!WJC:-' ]F.Z!5 $^)VE%M@I,#[?,VI2SPJ^-O=VBM>@;U<69!=
PHZ2;646Y"=.%CC,Y3F +-)XP_FSE:(-KS9MM9UT^F\KE_'#7)>E/I<CB/_#CLGT'
P*\ 2@KF,8O1*9KS+PJG7F5,$[VH8*W9,4,)#%Z:YE; #;?]73-NU+OS/XRHGH[QF
P)&!4TC3,, @6G2KKK?3@E9Y"(WTG730V5D0@1-$5"!"71JQ*(Z9.KP$S9+UXS6TT
PQ2J@ M*:,X  LJ,'I6Q4PNRAT@*X-!H*EU2TI*'A.=-_(>*NSJ18X!KHER#3\#-Y
P9""X>/'Y@PC"L4ZTW.\^=T]HG-ZX$+D,WWJ]Y-APS<4KQ!"86&)"@@,7E)XY#(OL
PV.(-R]<3$NP>;GZ+HK\\Z>]47V@'3V6Z 9*^718"&(+W;X&[:O\9&UG9338@Q7B,
PV_9]!]](3'*BKR+7G !S'&YCBSEVH?+*(9\P"J[\"7#4:GUV%/&D)"XU+QGY0O$*
PT?6YIAT[.+,Y/D3&?]8)D%+T;GH F4)ATPI>W"/X9<9<YT@L8ZDSY>W)$>:>%$TQ
P='.<#E9(QP.H\&-YB-K4Y=45AP:UR^DP?$Y(T&KW@_4]T!GT)\F#$%4P]1FF'RM<
P'071X0R'J&4,&"DBD%*8J6RJ'S8AW@,\JBI"-.XD@V7[0:6LE<)+*JP<*X5LJQMK
PM!N&@5E7[?+[0DLR^L+66S3MCEZL5$%'29BXM6< ]82%.8ZB(=C$87NW]*S)JO<R
P3GWOM"WX9K$'OI\(]D282QMQ,+_TD. /A\":;WF!8H,DB<,3&K F;\/F*K^K2>.Q
PM]"IF:EK2:TI*?KP(SIRM ?>V.^##0](OIEZ5XV:(_\KK)OF%N@B1='JS5]#.+Q"
PA;XNOC=TXJ@0<W.DD)5T1_2GO@&/C?;._T3P[#QA#EZC_2*<8 $E( V)CHVU28<D
P9+M$E9[O+D_C7%^Y,^714W+/I&J!9I**.]?$9'@[!0>79$=C:BW*UG*$TX^&J0).
PXJX 9#_XLWH=.P7\/K7LWSQ]GNGH6=.@+,=W0)%D7F4WO*]B)/%$CK\*_]/\B]2X
P!3E)X7D;OQZF\L*7RWL%B:W+AZ9GZJ65ZA O@S1*D[Y>G-O$FB_"I"13K2MDF<>F
P8;LSUY/#\0ZEC7CQJ,,BMOO2<C469 +4-.^&]$SP3WL'<(G;CUG"GL2>&_5<=IA1
PP55-3(8!HH0\O<#@<Z(-;:9WA9TW55EQ:L&J\Y6 =\IC.'\*$4/B[W#S,T'8<U*%
P7"*<P\7R3R'0:O/]XJS.$&<XK]Y:]9Z8K[Z<L7C9UNUQS4_A.Q4@%VD3S'R!H!84
P,S-K&T=SG_XV'XB:Y^.3W^ 7<\EL1BA-\2T_/ +JF@,7Q?6S6)'!A.I%#)*2]8DS
PE0G2WSP-E0.&^]D[ XUN=3R9L4G-G^#&9TE;R'C 1@W+\)FT$FUV'^KI]SJPPYZ*
P:X,HT8F)N9DMO,RM86ZVB 9?2"7OL@P,\22Q7.SE]#-F,,.D/ST80:SO"Q'ALN-#
P)*B3%C( GF2.5@=(:1R@P/!:G?*+4A/[$F?^4M[VC?G92'0S<#IO@Y8Y&\\UO8#Z
PD0\'$FM(4)#HP]@>HSZHD9U#_[ V/R,/V/;#J#(D)P9_? &?^SP ,^>$;BS,,2W=
P-;7GPV3C?)4G,73$Y=;0)Y#>U0>?@9?3E20^A(;4P2V-J"[B4X*VDP,E,1REVF8S
PWQM%PMLE2(7.JAE%I$XUB.U:BI#<)CP9V!3N<.5;8%S@"HFZO#._1B&2W%&' V3W
P$XVI,9MFT*DNQ")"G:#E^Y2?0QQ2*C$B  ",\OTL83:1.V8V:7" Z32[8 JN7;AN
P8J0KF!C^I;08_6VY^EE83<9/Y5@ZPK?7B_&K]E(*ZE22GCM>-Q[2OAABO#"[U)M)
P]"DF,9HAD3^[),*%I,0J&!A$6:+:\>FE[^V1F6EW']JU2]H+\EXU6*..-R#%$3)W
PL-_/1QXXH/%#2G:MEIQ5A,J<MW6C&D+N\>*X_!W5#"R*9P4JFG.BR'-K!0#3L3M-
PZEK6)G &S&_W,1#V?H?=I2$Q]%7*L5<ABDZ5,.=:<J4(/0EBJ^D*!N)/PPD=(<!N
P:1+1;64N\GYE2WX1^[CNM"$$@3/RPRW!JW"N@1N[#C;A,T9"9#\\_WUY'*V$ ! W
P5T@STYR! R6MZ4WHSYL$*+-K('\)TAH5#Z%X)U&,I:=PC63WL!%H*L6$&6'/Q+-6
P=A9Z=I9G(B"(M?K9;2H08&U;6C&VT@_#WH!1SB"<R7&/G-]T5'@6AQ7)RZ]3=3L,
PAA<T.S0>EWT!W1XYKZR-0EL9XS4H;Q>4]XZNSW%S\JHWED3/2*S,00;/<#-^G_@D
PZWBN]_B5V<HIDMB]' E&L73)!L=$#4N>#6@EJ&YXU]H2X"M9)EJ; X#U2-,5OJRI
P7:+.L-O^]\RN=,>".#X=@*N44:E&2R2>K(=X &-?I5!ZH0O:1@;3='2P>W3.I*C3
P4A+\EJ KY!;9P*>P1YB: Q&)10K.3C;NLL'T7_VD49(&\+DV3/6XL 7FSZIW>OX]
PMCXG#"7$02/P6".=>!E*7*OJ_H(V RU9H\ICW%8[I6VGP_Y+"\GY]H!X\B#K#1F;
PLBV%M'L8K&IHY&EU.&)J'K5$3_O?E^/7M1!T_;_.<7S^);25^<88(7(L,16^>8[-
PLN"BR; _1$$Y:W&--!$BG%A0=+PJQX^$[=>(8IE6$!M'4H<28*=@C8!&1-B<-2J8
P, X.8LZ[$OZWP$&Q<(5N[;8^#.KT'(4E5@C>=0KMX'[T@S5EFB0QQB(?9/V^<!QS
P+U5I5,Q4=$VI&V2,/+]W<7KY]YZ<O.(^182)QH4CLJE(&\CW? (V CQX=Y8DW_Q[
P,.6G.Q0]KP*>/L1_4<55VY4C-*1N@;W7O=9]KZV->@P[E:M1J;?'C+&^Z^1]CA'+
P.\.N $WW=]G"*U<S= <'#?E:2W] '^FE!=ZG':DUX!\.8@X/YO0HFB)'K^"6WU-B
PO_L3I*NQVM2^O'R_M@A*;6$P=E2[*.;K)#WPCXK"Q]#!C@*%+[5HE^+7V+<_GHU)
PCR>[Y#8(<A$)?@,QL4&IMBL,IRCF'S2=B?41S3IU"?-U7ZDHUOWV^?*=2,H>'GU.
PN.; Q/5;##LU@3.TV1?_Y[JZ&M64DB"9KQ-%],W[DZ$H"@AQ-^4+T[YMQ<^GXHXT
P'(?.Z=)"6&REAU,=&?N82,;&L^]S*>(CJTO0:26X9O6>O$+ ?F@K. SJAQMW*GN1
PS67RCFV[I;+;G3231BUHQ@L9IK*'R_E2"C!,P/LY[U  *JC,AI)R0C3ACQ9:Y!>P
PM]]/-9S1P9N[RN+") -C*L+1=)QQO^RL+5W:B"J>7*,/>FD92*@,3I9.UX<KC"%Q
PY8L1!OYXH/,%%% :*M3=%]Z2#'PBQJPG5;].45M K4!=6&7TMP,K=5AB<3Y&0YAU
PA3L]F%D<ZU1H9[\X=_?OL#8#2\QUXFE1?_DJL+N1)AIB !#KWR+\>(>40X57?<,$
P0Q@A$PKOS1)WA\>SXVI^/@Q#T1QY/WGG$/@ACXG2'W((_6"Q<,TWNP/BUIOA <=H
P.#KA^G!3!T_6(5#0Y8\- ;O(IS+DP7D5-#9YJC/)@F#&"-/>U$A5+[F'^_E7AIYD
P>N$(70]##D,1C&-R1F<F++(<9%G)SR)T&U2!_PNE)^1.&/14NP<10?X(9@X9WLKF
PXEX1=R7B9-W*(P0O3I7@4'KR+NBBFP;.._V.^F)S'R&GD&?U2N>5T$^_W0RDY*D[
P2%R6.2YE30_?E"2I*E&PUF52G!5/J)?87VT+84D+YIN"^4E0J^36+T 1QR@ K<^(
PGT6E*+:;PGZ6>(I &R%  XSEIOCWLZ#DA:S;V2X-4Y'0['/N%FC:A."O<-.(<79]
PNS?CG^.+0O5%,=Y,03I&VKGI#1UDM4D=?)\6DFMD,Q!TX7<E\7Z"TBPC4-;CG@P(
P1EK!**[RO/#QCZ""@9MO#ET8E4M,U^?D-F5[XS]'-/::,X-J-.N9%I X!CNJ(=7*
P/7%/N_O!Y*\ZUBJZ)3G-]%C%'LZK>5H:Q>]GDMP1,QDWC88C[!!$V\AVH,0W>U!<
PIR[UW5T=MIF590X.7#^?RA_@9DZ7O3B$(0MIR5;7KD';WH2#F\EO.%* ;;6-BLG>
PE=CDB'HR\.ZPRX>O44G?=CU<*S+W^=3%E (-R>RA:V^P66:O>WQD_WL4^1Q@7,6E
P/51*@S/$!T/P:> \DOV0T:99:"1A.0"DU#**,]?[]@.:;SZ6!P1"2ZK97WI77%MD
P5T I/H'1& 94@B/L:]ZU;C# UJ8 ;4/6>:X"_6JUC(F-BR.58%&#.K]\3HJO]C< 
PQZ$1F]9@84_0[+WC)E]P&!J<I^\Z+_]7/D]^7PU(B7;+;C_ BA'YC+R@7B$8Q6E9
P6WPZ;0G6'AE "T[SM\TV+W>W6_Q7J5S F.?3UZM<\J=CX- =E[#;*UE;ZS B[&\)
P -GM*^PK=OZRR,NAAZT)XU:6L-.P*#L:S+W4N<(G'ZY+ZV >&L_"CG:TCJ,F$"Z.
PS!M!-S-9R;C6]FW1B0D_ZZ_=OW51R0@[OB,(RXEP4R?/""Z %P]\RCD7?I=,M.'B
P(.[+ULEM60E?*++0(BC5;4<96RHIB[%O)%JQ+!\2HQF*KF*+.$,%2:-YJ1?QSWT,
P=(B;U>!C2E>PKH01_NKGG\@VB*)5)J?'_Z)?>CSP&RXD0.EA%M=_?/IM&T;CQW8]
P .]]4Y2.*?S&%?18FOA+X>XT-CJ-HJ&7RJ%S"@^MFO:=HV[>/[91_JE&$$!\9#)V
P-"C0)!;M\M9>D$!AD4Z2(\S5>&*N?Q%;V$(C8%.ATEK\9,_CT;)55M"WD;'>N^#\
PXK?8O*I:BS+K]7NU\4%;C>=P'-=5::)NU";CP-D0"4*U*2]Y8/JA< 1/]MC#C!@H
P?H4[7%/Z9?GOD+F Q,41T@YG\1!&+RYLD6B U+2*F ;8K;:4BJ+PHZ#]M,5[UX'=
PL2M,/SUY67IK&TO9S<D*D,RQM-^R<R3Y <5 0_%U-KHIB,V:_E:XU^E'H$+0X308
PE (MHRG-/(=6#"XKOXTK4H\1J*)8QDVH=F]@F%FM.0HG@6L<\>RL]20+.3[6Z&0I
POYOK:81"CI->TPNI$G'&N_5_\- )]T;8G'^5/B-!"*_0ZI01E;1+A$^\[O<Q6R U
P7$'4R=WR:!2W]RSKMM0']82A;U;N>>^55O[]1/D3AC8JCO+1F*EWS;[2F3Q\_!MT
PCS-[^M7W0S!A=7MJ0Q=JM\QT&A*"* MKN+_CT[G(M-$R<FW:,@R4X907:EC)^<1%
P1?2-7(Q@,EHMA@C$>(-#><DWTV=;@[*O0ZX7C;]\DF<J]3UD<"EM[0'Q OJH6<"D
PEQ*+,U^/)L!L?G8W0G6!WK@NA7_P(]IB6=P&/H"8@JXHC->55O)L<FMM/=9&G_$0
PLO@]&-6=WJS0E1(Z:;_*[L=IK!2/V+7,28:K!$&Q$E4.5:_;"^R<<:B'__[MOR$?
PQ^CNGGQ\>65,)*8#)P+-N B[$<18+X<[G7J:#X4/C2BM1O"\1UOX:^U.;:LR]5'Z
P_CU2U-K6;N\?_.N!:F4RC6,L;7J^]$P9MKB2-_N$TCR<SV;+RQ9@^:/YN?28V8(#
PX&+:DC>3L=2/&-?WDM-'7M["KWXHFZ,1L)X*T1:8X.-772G!"'Q5]\R--!W5X#BA
PW=5^R;R8 H6D=<[2 :HK=ZZ_1 &D:3E,2$F2HZZ"8+,(+_9\0>D7E8?' J 9;Q(A
PRE4C&LD->#A2?<D1_*;4A55"15+.*F6Z&DQ)D4$QL2NJ\H+]]%3L_&SS\1,#7G@>
P( 5"ST90!Y,ER+'V9!$-F?7?P>A<YH*>(,;="?WZ%U+7XF]7C4AY2$RH+3">=7OZ
PA)YMY@]:^B,H7[I",UE0J%]!%8SOE+,2K=H-T('#MTVI,:@[X R(]G)0T.+.I*S1
P;9MJK%,<0V(^\OMJ)YAHT'P&A/"5RC-XC@?;'7X?R50B5'3&]C)FO'9]@ 8V5+ "
P!M.*R.H43PI]T\=;@DNI+;U'N-/_ IH2,FQ$C1&$*S465Q%:<9?SJ[6]#!4^ 51A
P>[($R*ZTK2QZ4:S_-]X4.E0(T\A]7VC/MGAED."7_G\ZJ-)S=DX3BS?+6B$1S8#,
P9T0*9\U5:[L!/9#RS1_?%18L7YYCAINI:>$%*HL++MF0-RQ[:[J,;1W$RB-%:6C+
PFN7I5/$34:W+REX)KNW69";<VI+ E,IA]^A5L!8V6/MH%>B[^"H$#^$]12ZDWOO1
P"PXJ!!<$4B=-J*)1U1%&P7C'"/C8@T[>Z<1.<-H([9T1;^^"KC9 _">V4B)5KG6N
PH%G3.V,H*L:U 2H+<9)F$+I$.OR2 ;N?A^+Y]AI4OFTQQQ1,JQF#.?$H-#T>L*)5
P*I<1PH&7!UHS=JKXN!9P5D5NM->%(X]+%$ES/!$@0 HUW"?RRRS1#17K8;./82C>
P?@0RPX*96A1W<T,O%3&<+WGEOYC8CV=QB._6-M*:Z4L2]5 ,5-5MLV.'HN@25HLY
PC-A^1:?*-@TFP3M_H87'@B!2DRCXG, 3QX6<)&@TY-N_^;\I7EWO (Q4[4Q+RX?C
PV^E3U8U=]IF=MS;\!!3=TN;M9;FRZ(%W)N6F<_>','HX.BWLKK"3SBH5[ND^DM(S
P^@!N85A\RPQX+>S !ANU8[D$OZCMYD6MM3TP('!WF047?U6&6>K$/ V_,W^TALY2
P7ZF^T"F%Z$WS6S=F=4AP$SJ_1ILV)0F?9)@D",A2B TG'^?YYXBYZB"<I$VOFAH4
PKKZX8)]+T+LLP8.'[5)H'Z=28@.^>RI2V"[.J\!0[='4G")-U(.45WF1 AU9"X8O
P#(TG=6BKZ7:Q!];\4 H?'FRB.H6!R#4SG!C_<89R%J$[/V#IW5)=@N6%?)LT<,G0
P;"H;Z&ID9#.N')OTZ+1LLD:<\) _ /,Q>CB&<5Q6C2:*EU<3UIA&'@_(R+6U3#9<
P-B7.EGLD[01O4'GQ7LY@YU/P&_E&3H.%W3BNK9/0O>7"LUH%61QC]#O='\MC&P18
PVD[^)4'@ZPMVA4)*!< 8!^\S)E#(O&&QFSBJ#B+@4JB1\E*^,4_9(MJRJ <JXE6&
P"K^NSBP6<9C1=SE69L>^9N%V\PP%W&IEL:)EA!;RT4B\[XV4TWY/WD!FQ%G/Q"9_
PMN6ZW4-808]^,&LEN@-_')P_F)I1DORD(HZ%J_P%^+_69VI=9P0WPI0?<4-NW9'7
P"_4H4KNB*R?R--)HU9+QIM+JT$Q6F-)_9/&!T;X(?8Z$S*?.V,&,!70FS/EDQ_$S
PS@V1N9PA51$7$<:2++XR../ ,(<]B*Z_M,!(CO6A)W\-&>67BHXL@O2YR&?4,/PG
P6ZGU&7RNHY!7E.VO"46!S8-UL6#<FNG5;.D* KZ2HH='EXK)MC()LPI@-8OM]1:(
P2QC\8>1*FY1;S>%/,OG=V[NC!A A%#V_NT)LC>D:O.=BYUE;7V):>OI20L5L7(Q/
P<##<TE"\.,-&P@8["8<7G?AYR7<_+U\;91W'NJ2)X)HCNR\@9*I-D-YI8P<\O\@'
P;!NR*6-V4T26\M:SR84FWK0DUXL.!QV-96QX#!-[1\G$PIC=+UU)A;RG T6EW!U;
P%V=(W3)FB'L@P:*IWQ6'-D6BIN$J?^"20P<9-6FJ;\RIU2CR8OF[K6ZGH**IC==1
P18;0-PCBQX2;JZBC9'L(/!P^>RN1$%(,W;\9[3#@N_J1L<52R._+=,-X 9G0W3X#
P(?5%8=,\NN0A,DT\+,US9*=J; WF+"U)A.5LA@H!)OV.FK2'KF)=G6D)\FG=E+U$
P3F.)2?E]0DLH(RD"/F'80-&L<A3I];L=5CVDR,9I ,K.R7;3'Y <4,19A&5D,C/3
P5+N1IJ]U9N@EL8NT<>0\-OGVCV?>WR2"YI ND,4OQ@0,UEK GKQ&H>#?5)R VY'\
PK1TF*#\IW7(SIXN[B;46/G]]*V_>'=QK8[!. L<%]$-NN:-B *?^&!U?H5I:;CD9
PX9C"+:"TU7D=8XG1R'SKYT*/*L MN>C8]ZD#WT3:PWMY?'S+V;*Z[KO_Y=E(QK$I
P]X@OP 75,)-)5"&] =MQU8>+/R>1,U$4R"T%&"ZDA;=3((N$ST,QQN9VN@Z@=<^Y
P3/<9&W%3V<(Y@&=%.<%*X8E ,Z:]5RA+;,G)5=I$6?+'RM,/A.C]G;J8ZAB%K-;$
P+U7^LI2=:Y%B7!M"8+4,RG@4WYOG4C.7'.M(/CO'R?"RQVB$W"E&"XJ7RXP% <?(
P)%1/*T _\%X[0&6%JM;>3VK0*[/(FFC 1-?=K29C9^U@]W(4&@U+<E9N)E]F CD"
P!*'4<6?.@""TD^3U!Z<&<I-6-FN*Y:2K/1J /YP(Q3"TY?TG/4@91M#U;*%-)M$ 
P*%GT7<;<9!9$PBPXH/L@VN$*\( VX>%*BGM'%:?+@>?Y7@*)6BYK(CY/'+5)2&7=
P^G0BVL"USE0\)8OTK#7#?.)(L7I/K6O<_/W5JPVSG0^$XP.!V4LW,+=%"=9^LZ-V
PCJLCA0:M$9TVN@5,-]8JEU:X59?7Y(6)D3JI86O1,T]WKL22WP=+'\'*E9&X0G%:
P*+H?\E8]F$$:5J-'8-DA!I9;TGC9/S>"BLT%NV*7&[X0U-AAA+6ZXR8I7Y3%JIJ"
P?Z8W56Y9F,K6 I4C+.!A-)R3K0V"44GW00H%C6@?G;5"9Z:WGO.3$=%&912A&?"D
P7UW,FT$X%RE,"Q1@7O$%/;,3VVE=%I7CAM :860*#%$K2Y@/S- IB1-U%B!<;"O@
PJ?@^L&N8&2\5U:1>8^9/_/')D_3N[^Y0Y?<'UB#F#!ILT0#!:T[=!</M87<M'8;3
P1U<+9*J8+I^M<3ZJL?L$BQYX<<_:97X;\+&5:"6=(JU^LN /,RLMZKI&9+VNU10?
PCXT5J'Z73>NO[;]:U@LZ%(BRF$K[0]]Y@1!VQR#=>-:1'_<L\&34O&[MI?[8JA;O
P"_*6ILF'@;.DJ1Z#T@C?"G:(N"-U8.]D#N&4OJH%*.@X5PVK]8/'D=HZ2Y\2KI;P
P\SK$G@R1;0!: J"OU,R\S\]'DA#_N+$JUE!K]H*8I>1T3X);^O _O8;8[?#;<ZA$
P#O$NGDF_-S+2/O\R!+F*_L=W?#RFNG 8(E=5?+(T][/Y6AM#[/:_WA0;'%T_Z%FH
P:<9OF6_5-,$<@4K<Z1%E+RJZJJA&;Q=6D]G<(1L)H1!UBE,?HDT[H\=*3:ZJF/34
P+_8DUCXHG.I*=7!0MYT3IE,3U,W.*W9.\>:,ICU9$-G2F;]9.5&=FN;W')H.451U
P7!UC2B.'DK::93DGK<8)MI:[<P[FP3AZ>0RX5'_QJRHM4"-]"_17\QTHG#YJ&?W 
P:<(.^0*]-6]CVMV&,RYPEBB/,VYB'NKQL!F!J9CXBG8Z9C=L*:,>#CS.<^/:ZU91
P[8E9OQ(9?BA[F385,',K+TKD[D%!"%N&MZ[%^I[Q\1')U)MTA7G6V$$]M\.05=]Y
PE+Q9I.\WX7)%B$P,>4A^W?>=HR%=,_*_:5;9T@VU7^SW["A_SFP"+"8E1=[@&0 $
PG-\JUQV]I"RO,YS<[-_.QA:[R@0$P=#XF\(SDY&B8"1R_NQKUE$X')]BXW!)O+<F
P_9:2^' ^"529Y#_EZZ]A;XKZ_*FN2A8H%X@*XKIH1(XSKZD8\#$#Y5F'C+*CU(NR
PU$"8)#Y>LPB%U8]BFM*]/?F:BS.+*FXY)9%*V^2"40#-?9(AL3"_4KDA#_X38X9V
P&]SQ-! KD;:@.B;+-U26MOSB*2N=#S8J%G,IV[],Z;Y;VK/@R 3OO*+3PI_2)I]P
P8(1Z74$H)'_2_$<IABF+"V!4 5%L5W;MPEP'@/D27L7$<GMIN2-/W3/SK"?.QC/0
PC]KW?&Y*H']JZ77@+;B0H$1,E\\,26C)_HRZG1(662WDG1XNY'ON2#*@958M&U(L
PJR/3Z !T/<K[$N/#=RIJ3I '<<*O-ASU(0[)H"1#F'?NQG;/<A<3%63A2)1BN'M@
PJ#HKL_1O?UHO<@V:R 3G-!V]%]/[.LMU 88\;\$.-RH!5 R%3U=G"U51_WAG_/)F
P3#-PO-CGE&G\@_+ $2J%3;!^:J0".(!+R+P]:'%:">> 3$'#.$CS</4(&QT@^KI^
P9I/=-NL3\6NVP<V-R8!M(->9]K JK0,H+01UJC8$'?+>!\Q9$6YB%Q=773L_?F\E
PYR \YL2DA9A>Q?_OOG5.G1_!OYUMZT\O6C/>D9<([^FV-5GLK&/%0S)R89!-)@4>
P;>EL%*9>.*:3&6T 0J]<W3F0]D^T%6BA#(\R-4E(?L2?61^/>P-W^5&+1ND=32G=
P1V@-P9*TH<\DJ+=QA:Q&=O;FQ]+*6_8#M ?LF*9RX[*UF(WYTF4STD_<04(+(HWZ
P24&_>Z/!?1OT!%$3/F!YZ8?M"9\06:M BTZ+Z* ['^#1]E*#-HOR(#W(A5]F36;'
PE%9G89^W5%37#AM&:TKM_6ZANPO0&89,%+DZ2S@?".\MXGGS_$MYC\8P00<Y5%,*
P":J>R-DR!EQ'X3JZKTTEHP:X=UMX;$XGUS>&A#-)TH\B=RU7HA46GEIGXU4_?_TL
P)"V]@(Z>EUJ>#]$?S%.(PZEM>'A0<]73HD HPS]!T2"GC$795):@6< Y54Z[D,M:
P',L=1=7.U;$]M<--!4D@@[/=N>',OWT:E5<^@[+P& ^8>7:Z7?MK2ZG25D,?>D:&
P5WR]8.>&MM$VP<D2\GFYOR5UWLKA^C7[ %'(&IO%+#BGKD!/__Z0H(F'2"!V43:"
P2F--JO.8TU"#>+[5Y6=],Q"L<Y?(/>(3-@0OA0Y)MYG<7"^45$'$SBR$[Q%KCO_S
PY!N-!QN-V6[KH:)-)@IUD'71BG!9AO'9VB/]'PSXS<+0QYC#-KP?PY9@.0JF4#>7
PYT"?LU1AJO02)\>46NI6:XU3>2YP@VD!)\6Q#)W]0!QZAR/7WK'WJQ,?=&2"B4_N
P__US38/86')YU++ K>RG-XJNF;N/)%17D>EHK: J)/*0LA%5K_-0QX4!?%:H%8$$
P=KQF?[%@J7,K?D<JA\VH('VJ#$SPSRKYS2BX<T;>*"1?.)SC^X+^U^V*E'3DR>F\
P8T6YTHSI==E-D"+?OR-/]#']FK]X,'LY7PEL@W"Q895-P_5L4X-8['X>[QAT_,7P
PCQ01<YU30Y5YGXAQ26+YEN+(/EL[<CX,1SG#)4C)7MNQ;;,W>ZV^:4*L3UFT5DB_
PBPS\PZKQ5=C11RIPJ'U04$5(N;*O."$U\AZ"_N:M$][9&]E*D(HN^ .B!Q^2"U.4
P&\LHA31>%USNTFJ^+KM9_E;O+O4WXN\ZC BD#3RE.*E.3&@([:4[,:;3T\PCACAQ
P/LA+*G,.6(DEG<[ &[SC?+PA?L;[EUK4!7B*:5D 1,5<RXJ9WN4;9V(=-2?L^=^<
P^#54;K'.CKUGF/4%HE1_V/!%I0O ^D6JB'Z:L5TQY@GD ,0C<U=.^]^W8S=UXE;2
P2,NQ;S'IP4WB8"-[V.!^B[AK6A@,.)?V8@7.'!:I$74.7CNUD/.9\'=M$<?X+?%N
P?UP>,G2-T +G^+'ZZ'E(S%&^LL4%LB4G9&A5JHY,WR?.,@BA3O^=QHB+J8(_P40P
PZ'KT0J=9A27(=H'UD=40:R!GX%PNH>G &FUH!RXKK4]'6?7XT,Y6!QJ&>N*1ZLJ#
PE#OHX?IZ3DD1 HCJD^8L>Y<%>VK_F6NL'>"MM#!@2002;Q&2]:3'G*;N;82#3W]J
PGTVN+.&[EQ[4/@#!&AEB]P;@_%['<PR!]U2 5]/'.1<Z3;F-$J[B*$CH&C3:PBE1
PUH'A8!5-DA%_F!(SL.CC+:ZG+J%1])?5 LE:>SHJ).Z:O,(65G37X\$9$D2W[9;+
PPK^H;[;,J'RZ++;8-;C_@SMCG/<YI-('TH.T_-005WQS'G*F@;7S,+OH4> 'D_P]
PR', ]+.-8"&!0;CNITMX[+U;Q1A1.V0;9.3"! AO<TFL*]Y&"<%I$/,53;:CCV6=
P#E(538?XP)&V'S?N$L=7T.Z>R/G)@TBW(<4KP!@0EW[9%/J^)\"-U4^X+PJ^;7[?
P;<++H*^+IKE91KFRB21JKP5RY<[29*/S])0CDL)+)9-Y\V1+;VY^OTBH=+L,GQ80
P0A<]JE4G,8.=S<#\.OI.26>8ZL19H\AMB6GPM;F)ARK%T(2N;$X@JT-5EKPSDO-8
P*>0H<*M]0G4_AC $&;$HP?GI@>%,2@>/K<]@+$P_VNYZ<9,KTZF_AHP?D@]:2 (I
P53W>)V878NS^/#(+^5< ]IT74^Y9KP^'KJ'%#%>]XVC]QA*7GJ_J@; Y6/,H:66H
P.]>G=:"Y!%TXWMZFW?(,A-Y;E_P=([XL<Q50 '6J[(QIF39NO-W<&FZ7+KU),9A<
P:W\NV,V:Y$VGQ?E61,L)>A4<8QTH#&VV9-TSL+0Q:9,Q/?E6VW\)()["8D7''#&J
P38Y82%R%VS@]58!D%FH<B;63.P&'1@Y43(]+]7NYF7)J5Q42[.T<3F%&:-),2+!I
P*_@"2ER_\:G-BSM[E+H%9Z7S,H.VA=8:P&M3MT8.50NL$E:CYT$$WD:-WS:(F$F?
P\IR+U'WU[<PFF+NOMQ%38]I26X(B=ECH'PAJKL$#,C&DH!W9$I'N U2FH:9Y$N3M
P-!]=Y5XI<>\^^=<8,6X^;\CA,V"LDX(>?S#]MI1)I:O9/GW.1Z<)5L2$W966+>K(
P9TP3X/#WO6KC*5CY<S!?JP7 CB&7;7+1^]4J>"#O%H+BM7/8N(RH2DYE#)P?[T=A
PV2O4E(B0;9@+W> 3S.[&G^J5V14NH$P#*$92[I\K*3TW=FZQ>\+I6]C,Z1&#MR^A
P%.?6 W2VYZD#[7V4CVC@''=+>HS%()SL_H@*7N=3J(S*]&46Z'L_1@I9BKCI,TG4
PKTUB'4XZKS"P.J<H$6Q\W^D+_T];"WI8L%HDFUT)^(F%/6T^>=$JIW:SQ;9F7&<]
P(JWAPE3.?:BO&5A@:L#7_$Z)W)=<-Y?4WZYVU=T@7L8+\IF:4U.9RMO4?IR<C6EY
P:(3.-AN["0@$SJDIJ]8&!NU0%;"N&E24ERLP8[I'05R@G5'N$NKP.<F+W/M&L!CP
P:095=15>0W;A#=15XB;&04NIYRCK7^"O7 1*7Y)Y][8SG)'G>*)VGY;LCW$]J&2^
PV\?-''LD; 3G\>!$;"% 1VEBE,JLBR9B"FV6"OV4S7B\>XG_BO5SI.)R);;,*:V6
PQDUOUO(3XD&)7?[GA2VY<IC' $-L?T:!CJP;9^0%J!,<*(&3S9<B=IN4<0RP \^@
P>(!X-Z:35?#;1LF=8R'-"2[X]RD#)D$\(S0@['_UI0//\>!98$YJQ$&[:4DBV27/
P1IY)[(6OFT:H8"HJZC2801S,Z*#O'@*@2<72(3><D^N^40<T[4CZ*.G0G)#0R>;4
PRD]'5_0QD;EH5.TDZ.!$.]$D"-CR,BV2R(F#@%P5ZJ>C5^RC>KJ.^L+?0P7-UN3Z
PG'BY$@&:[&4-=0A$.QL>6GLU64OD&K-!+QK *V>9-Q)6Y:^ZG?,ZO&NIYVM"TCW)
PR#N@$RTP8I*OI15K+!H* (?AOYN-!A2&;6YO B:1$=#(]YH$%:=J!H[V^B5_IA'.
PQ+EM2I8 91.+X'U-.R$*UW+",L]'^R9U5PLEN:)$5D<@X.KK' 6T1,?1(6B; PT&
PSO(T6_4U\.GBE8RXQ7OXK..EM=ZG\]: )IA#J5'X'7G)OG4 _?#8>]KBPRJ!P+T:
PYT7+ 5>&P_\FQKLDT) (T5?9/77LMIR(S3D(0[>$*X3=*DXR;S7V@=<ZW:%L:#7L
P(G?98)"AZ;,$_3$50AGSI-=U.>8M9P5;I]*8#1U<@6:*SNYG @5:7SA5'")$6+3Y
PRP(F(:7&BRA18^9?C\=R;;/WR4%>7,-_"W%<8"U[-^*.T0IRM>G0):I$<?JOKE0"
P_HJA6X9R]=6VRN'IN+BU$/1(Y]7HC6\6!O(<7^%2Y)SH2D&]Q7'?:B 2J&1OIR%1
P3X#H9]NTZ)7:KLI1N@EL#J-DVN[ZXZYNOD5&"@3/706N8AE=O-2N=\Z12&0Z2VGH
P%Q. O9NR3=OE:K0T^!>M?W!X#1#,%XS"LK_X81HKDL\I8L-4)>B2GU/-FXOP-0/J
P*Z3I\]?8'%ESK3&CC;P/,P]-1IX&I93^4&FU.LN&.QJ X:PKJ5&(CXH$'U6BP.(_
P5;^R7AF\9-4@9?."MMIG$ AN"U"Q%?N:>$YJ=ORZ)/;MK2LF(G7R4(Y!XLC OG\&
P:P+G.P$'+B^)/-9ZKIE+]&"'E2; )F_W5,]B@J_0XT:.@E<-#<B$(;AB_1V'DYRL
PL;RX!)IQIUN9E<:33#)&C0Z018:M/E$'T0 $T)#+)NT!V?7/8#N0M>IJTV8"&G['
PL#'5YQ$K06+IZ];7'"*F0-OIP$9.YQTGB;,CM[ZQ0/>Q9F%&0>A\7"_[8V,81;'+
P;-YPO> &<A..T6E\36M7<%T3ESG#JSS:5LP YPN*1AP-:616W=E)#RDIX+FL]92G
P*@L"AK4+JD_2Y,7>-J&<!> RI*5VF-U?<HH\ I5K](^WS2)QU;'7[%'%-A9:BO>Y
P(M4.TF%\&-J.A&1#81.,5V;,G .9VJ,/WB! 4VF=8SO30-7(4$%TO$K%CM$"G5%3
P]KDKBNLN7FS@8//^D"II92WL(O<\SG^U+5WGWPP$4O7NT<=]=U"9M_EISTP8\<-R
PV!>!X6V5)\7P:+2!D=A.X:R%H'\$RW1#<H@=)IJ'B4N 1CFG=FXR)W-.FXN(%7#(
P4]NA NE6D8A:3>JIQU(6B"+X?#H)APJQRRI$8\&QA7B .$BI^/(+$WU3]*9WOS:N
PZM+4_8]W.;#)[0/+R9: GDPN? 2=+NL!&L^^A9=\B@8[Q^L$]>!#S@!/*V2W?+_4
PR)<$(Z3N%;D<M)?=GV()6_@VX3ML.]4T!^<S4)K-"X;<<0QT%PB_Y#0%T9M6ZF'1
P:-@A6)R@%ND:2O)C_TOP]/]R@!_VSC-A5S$'6N%\N23=5#+L0@'11+ ^I8B: EM^
P@>>GZX$<R(GN34T".^U4/X'B3N35%4T\UZ91L'SW76N)KEY?R'V5Q?!IN7C]<YG^
PVP/O"#)J>A+!V2!9% WHQ:1][ T'W%-DH4>(<#4&EN<4,_K_6P$O]^,CTFJW CG>
P$!X'Q;BHOM?@MW/KRWDM4?4-D395 >:I%/+W%>3.UK 4LVNH3#1OQ:-$= =MD_F9
P;1L>?T:'!X0\JNP0NKG)3"6#7.-F[K+0^8]8<-UNTZ4\?8<0<WPC>*5_=^,B9<-*
P%)4[O?Y^)_'!8;F2!B6CW0TW2C& J/YO,)ZE;S]L"!O//1LKAX )?9S9\@CFRI,.
PMO;DR2(J:HB;[+)%UGI2Z&'/(V=?V\\N^R\0<SD8K]B,W?RZY.78VT!*;@+#-S82
PP33P'^-5.WF9RR]L,DO"D>H^8L)^;-FL\Q0<,08V1DWZVY Z;H=6K/#>-&EC!+4V
P389C@<DGV.9_]+L*OH;4/1DI#IZ%<O&-3'%!_QH+PKO X]1,VCY[A^11A^$ #&#!
PX2^FY.(S9U8S%6,C)TL,PSR[']K'GCS1Q@?,)A7EF++)A>2 >:^HC.W#KP$77=0J
PAGQFJJX]4J!O,;4EN+Q&266'WDK=-J(/R>RP0D6N4 TXM9_Y:GJ[+6N_P)3F,\.<
P$K@Z\PT4YE]QCIY%W6[#J:;9_1U=6YMV^)>XKEV\#\.V/7!X"ED9 GYQ<Z6%Z=AU
P>R22 @521+S^\5K-JS(?@*4/%C!?JLFRVL)V@8DE"+]'.ET3%Q$X,T%[1_Y(Q#LW
P8M=:Y[6Z_2A?%N\6+X8\P+>.<I4VB+;[FQ+,"6I P;M?/NUE0]+EBH(M=PT_LI!P
P=)BM+K8OBW*CE^%D!^@O2G5W"J]:V/(42ZC]=U)+>[:D6AA^_$H.%\8Y9QKU)(S*
P]6T,USST#BK*&KFY+=E.GOQ3;;0.7:Y7]6%]!G!D1?MZH6Z.<*CI#^'/%$T!1[OA
PUX(9)3P!*;7'0>1_!GAXFECUO?44W-%A29@C#V"!ZWY\KM3"+WRZTLW'OZ3J3-S_
PL*_3[/X7#,]:%<L[!D=[^:NX@01!.M8#AU:2'@8T%S=DT?.@ PTN5RHF.L<7)@9&
PS?.F@B>*"\Q((G",%4.?P,!'62$6-.ARNDX["E*,Y:P?NQM@S\8@AK;NRI(2>?]7
P/Y*[1"_7A,C)*,7>5S_;6%>613+WX8N+7*39N^CD%CM$XJN9(]D&NWW-3'-G%>FU
PA>W2HL:8Q+3+A"'\+/"FI*FXG2"_O:XA[)! O<_:V&&G)FN .!2=?J#R@/ M5,@!
PH1G2PK;*<4<?EZU^F# _9 _WO73K]I+]P*]K,Z:MG_?H2 M3K9?R<U#5%H)'F.$7
PS")3R1J:30/1(;-&]SJPL"TM\UM4JH.V<V;JK5N'.S>$<B@?4^I39G\CP?^OY'?9
P/>VV4O&B4 O%)2#;^%018>^'59%$@&V3%+^25#N@<GR3[>B 9(#;2=$M[RQ<98'V
PV36Q?'3O+@(,1EE @%7"IF%F.-6'YE8?5L07%L&CW1(N09LB2]/;E!DG$1<HW[BF
PY&C]_ !E]]O4_7W!R=#ZX)CAH#SEE:K6GK4%9&&G@.Q 0I,\3;.8'"B_/ +[U:@^
P5I'"#7GS]ERON_<-=F#:HM.S!9"T8+Z4F'QC1: OV^D7@!VM1CJ$%L9  N6W^9=P
P9 ;TQW/HMN'AK1TALVGMDI//%OH=(UZB=;Y))['PS"QO4>YP)J[Z7<0BF_:6]@I2
PL3W'"=E68U@,,[7'1#8P*H@K(^\[^TY^#-01OQS\<TU\IDJE^I[7]5>JE=:=@8NE
P%JO?*D@@L&2-GM,TZ[\N>OQC1(X:/S5B1^S)C_"?F-S(N__E8_Z:ZLZ1T"2F)C"0
PO [1WXE]A):T?9XS7E:P4HXIRIQ7J7&ZIN6DE9,HMPF&7B +R;]SI!MD]CBN(*/H
PJ.)%B'];Z"S&>=RL! DU2$U/'WB=.0PZE<)A&><+.H4%>V!-PLU02@KJ$K*)77X,
P/,T94_:B.J(0>7$%:5AA#O.$6437U_ML84V;0&C9'FL"="H2J%/=AH_PS\)_3!DD
P+#B.<T]DY&RZX: \R:PZ.;-?#NWQMQ8C$G]K5U0Q,]S;#4/AK#XT/-.K=QK$XL%.
P#3WHR[=3=0QD4'4+YRES&5N_;:1;*$D)W0MG+(7D6%?ZDV?#K1 XDHE;SD8JY>8%
PNY\3BE8NBJ6(\C%!G2<J++8-OR-=[72<Y]C%ZE[KOK3(!7!?K;23/H*QS,.6N_WS
P^/8?M:YN6K33)"(U.!_+"'^<>':R*K2;9B133J8[0H.9DI<W6EY.8UP<.=Z;B&]A
P8>ECN<UR^K2: DY!G1[BU34XGN/5(@_9>3E)<K#_)./=?]Q',0VXPZ!-WIN04S>N
PC5+@.8Z-$U/#73#B0XQDA7K"64;K'A#(0N^[:)RV[M,W -85[WP4>4ZB'AL *&]?
P?OG2T35<3X6_V52Q=]RFW*HIKU:IM?4E.97EW_F=B5ZH'F!>Q&HX]+V%-S>(S.\"
P%-%P<+2%J00,\_K6M?(3(,#&O-SV7#Z%00=+<6B?4_(-7N>XF3]%?.""[=@3'@Q@
P&+?/\ITY)^#*%D[D?/Q&*:23/3#D)B1LFT9#X"-8/C:WB FS8?A5"H =<W=VGY"-
P/5@V4JM81:/_2O8=VA-(>O;^V9<&X9E03SF\WS)K&!A,-+M[64W"C2@9 8.P<G5U
P\EQ0#0MI #R0%,=X5&1892^CXOM?D6((0\UZITP+6*EQMXD,6AF<^RC?R:=\47T^
PMWHX]3!'X1L+;(5G'I;S"Z5M]::S)XL:81K3)#3MW['RYH-ZW5FBP *TT0$DL3Q8
P=?X\@XF=*B3J+=J./5R1$XP0:0*6[^/0(#"%_OG57^_&ABT'QY.U]&UL$L3M[7]$
P/9D/++?MZ PCBZ$QUXB32XO71Q2B:$SQL26*.==E !^DN]H0]44TK\G)VBD\MV&W
P4LT+4_0RG-%D;PN4:&PTOKXK++A5Q),:I5_*YOJ9N#M(NTV?T7O"X^A$Q!:;CN2,
P>R_!)DI:P/M%K"DB;,3]>V/K%F<S1BSUZD(JQWG_L';$MZ3!Y!2ZP:60DSSBU&MT
P*X&RE7MC3FC-2T?YV\Z/63)%/1:<+LZ-;T0:G$%>=5%37!#:*#GIUK7G$EXY74C&
P7J?\]QC_T2&L:I6L-;OL.#V;6VU\?_8Y77N%CT4*3P5Y.P/28#0_'9)0L*K8\$@<
PW2><HK$+.VRX83F3W1XIJP.*I&8,P5A[F(F4[' E,]P)&HV,^'.MBG3H:GM7\X#C
P7V;VY!^HJR&#45+0'P0F(FV\D4\6E]01Y?6)WO.>_LV)E-3Q!6L] .*GL3B0S_@H
P]&H7IM'\]/SAY2>;#/^$R"WW*?<:K$9@)G5)LCMC89C@B58=37B;5O(/2I5>\+;G
P4GTM_(70J4^9H23[JC9B3LX]2LC%D V8R0>,R%$'9\(IYJN_W2ST=R[6^(MCW<59
PZJ@R:0]/J[J/.D4Z0Z.TRE%A^:\ OO387K*@D5HXP@G^WE$C6M ]H6(O):+GP$SJ
P&')'>!ZUG8K &XXYB Z@(U-*UBU'(Z95I\1AM7@HXNKY[K\<>\IO;>O5309'%%<K
PG7;E,6XK3ZXX3<T]]J/SB_$]3QS[F2$5+#4+!==)R0)8JJQI*C4N?#\KV,C4%CCE
P?!)R?=#R')GW)A'\(EYS"LJL>)1$3W,)&;&D1)L9F79?;[:^R'!(@RL@*17*R3!,
PU@".X1H/%_<6<BDEJ49:Z].$E8IV+O^6G@KC.1>5SP=^UO'HGN7XN^TE,;/<(59R
P/<[GHIR(B2@?1HX-]THP,ET-=RP^7$.[F<^WB:C- 0;(B%-SD)?"%+]>N*KXHO5D
PF+J4(YA9!>)2NH#F,J3##)J*25GPDO?0S(_8=CFZNC1A&!^* D0;Q,AH8S:#X"]I
PV7)&M_$WG#&\"[;QY8#&,WG>+(>MI#",-3CZ(P/$5[RCGU:A1-U818&V!*_EH_-E
PT70"<SO2*H,(I9[E@&W.S6&;V^>"++G:_,NR_5!^_4YX8"0SS=':D&\7!!F\+$L+
P$80RBMP9,%PBB=USB8%-J8YH7<>Y%)#)(6'1C)S5(_;%).L'LL"*KQH@SK_8:*JD
PIPC>BHJ]#)^5CXY_B2/-R&4'GMY.HE.H[K"<S3,'?$X:GV&;":YHKLD?*_!X@E*F
P@X?^XOXJE'YEPN%9+[I51!->YA\IS>>FE;^/7+$U5M MT&F^"R.8SKA])6\H(2(Y
PYH 7/.<;#C%T:1EOIM5)K;::K::1[0"=?P7@\4TWP\YTWHQ%!Q'P40LSC_#ICS[V
P%^=M-0^Q24P*7?51YR"M%\.PM'_A!,UI$M%GK@%%"E@R+*3-VF'IPS,/=&@S6V>]
P9U-[-U6PQ0,[:\&.$1,MCK>6<ISR0"5A<5^]>X<M=4JT^7.F;//9[WB">L %NV ;
PG(BR^]' OHYHPFG=*-V0+YYP:^:& ?6!LX$#[](SU1_$S=U]2%:1+_,G ZF6CFJJ
PO&A(18CF:V$T?R 1I5I#/=8^#^(KAZ)",'( OU)9H[ )[6\8E3Y O;K@DPJ, ,"I
P1)3K)QN_\!BK_>AQ<Q%4X:5\017K.U(IJPD0]25-*]68=A&WR.88=.9XFN9-PR +
PFZQ$;?/GR@*L0;U-[Y B4A;MX3N0OA3J^)Q36MR#WJ4&6F%[AUB@W'0\E Y@D S?
P^6$?9+E=OYU4H+CD@OP?NGP<D 7U%?FAK7Q$PJ&,S ]6&OU?:P!" VK&!.H'O3O$
PI@%]FUX\]R,./00VEG_%*4[9FS4TY#BMPZ02&7RI$4UD$@B# %6RJG^*DI4W45)M
PFFY5<K2J$J=#9_@_>]OB-CZ[DP[<,LAY^"AC( %<C""7<#(LJ+>0-^F*,#GW%KTN
P!#1,S>A1>J!&G8IY^F=!>Y[J?%/U3 %?VL!)#*E/\FO')G:0FP<M_*%'7DH^_@2X
P*DOYEQ.?\<K7)([O3KT/^/C4928ZY[/BG:6$'.MCG_=S6A62*^#='09,3>SU(1O_
P@@I=ZF#U[ H/+/A1[#5[%:;K>ZJZ/RI<IW_Z5<#5P6M@4+YH5DNBP. M,"<^\1!:
P<F24KX8>$<EF87(ZG!F;_=<3"\#(W!5?+)YBZ+'D/0",8B6(]#"OVS 3-^A#:^/J
P=0\T 5]^I+X,75$$C%<4FL81>@BWR,;<SY&C"1>':[1C0/)G#NC;-S;UFNK6EG!:
PC%3.77 E<"T2*.BY?!0^-=K2@]B_QO.-80G$*SG("1I#*6^!"IE\!9WDU0( 2\Z6
PCD(!S5V\B1#AX3XUKH;BJKTTSPY8'5VU+=>%N?4$-/HOS26[!">S,P0X_TM"3'9V
P&E)$ =%%(\9&*7L )CP.<N/.7B+-MIZ"SAWO)S%_B.J!UGQ_*VY_&0FK-A_Z)=R,
PSOLDW&_#9(2B L!MQ\24(08)%A9F-ZBVE[(<E&A( [-\@]F"+Y4DN$5!9A1^ORFF
PV-15"+^ Q&UN54$V "W30E\#SXYH!UHK>@FS/6B\K<;F/#^<Y$#4W0\7TES0!&"8
PTB4Z.<C;=5*XO6($1K_M M>=$T_B>2!%KJGXC3/2 B)O/S;,EML?WEQ60XD%6MZT
P6>(:RJ<T3A7*H:AVUCJ'^;S['.Y\+PKLRM&BJ?$0",[\0$) FYG+B:%;W838)E2"
P-0?J' 9%3'JX <25J5,9\!,)I!6B$\9'!YR1BEP]9Y\A6"]#51+;TH4*B=*X7)T^
P%I=_AQ8+@2'7Z_:IFG]FX+/NOIHN1OWCNF4/,!NQGX)#5D!F<7K[!S)3ZF]' C!Y
PWO3;+@F,\+<2@+G8//2 IE?0>1-NQ31@U!$21S44:L+#3U;K<O06:W"+Z(Y-D1RF
P:'&"I7YU/@6L5YG18_(_UM"4G4!D9"D7!=F&_4IY E3U[\T\G( &_.B6_-!L;-]$
P_X CYGH4'@9W4XY[#)(F'5J&?[QP&*%81(@(_OZI*^\(;SQ@-3<(78M9FN6J@EVN
PZ4&F*:5L7\3I\;C$(:KS]Z*YI>Y(RND.6[5@^S[ ^<OY\F2L0';>Q:NUW5MM9-S<
P5[SRTZ4"E1E*1.4$H+V/A>;D'*3Q[/PX$3^,#FDA(A@XG1MNSF=!YJO,4I_;4%)N
P4BRZ:7;02CA>UH/']W,:DQ'L&K#NAAE H<,0$O'TRZRWO+_GR<NV/)'O*42_8.[\
PQC J*09O_! 3EBON4*8(#6S/T3QWU5@3_R-ZN=9)44)77.KN3^M&"[@F,]^"Y8&K
P;[MX^HPA^\GA=/2$)W]0GQ.AV::,)O ^SR&_)%TRR5#BFV&.]> <W(%TG7@5>X!L
P#!7)3M5>>(#9RM^K5/*-B!NP]'DY^KP)_D#O-E"7"J#9YNB"-IM)=<FH).N7+]UA
P93[HS#LL %#^,X?J#AJ%LZ$*XNUXXH1)SRB[#H"TT[BG5P;(.C"^'7[O*K(L7$#9
PY/R*XOWZO) X>_-2P+4?/HNJJ5+&K*&S_O09#S%D\%Q=CS'X>7-0=/K0Q*VV"8?O
PE:_#^/+C0/:Q6?S9OP,!XZF(.K6%X5HJ1R0G\3,=\F%U):F[M"!R[2[8[*B#"#H$
P"H^0<N_M%,L>?9)&Y76ZBD!*&- -HQMG&_OFI8D=ND3]X:BM;A%MS\Z0'\T&"H2-
PAL7;E=+=V]&XY_ ]<K(E;>.\A#LM3?4B2ZGT:;L8&#>$W;24RQ8B5/O6,:7>I/,D
P7OD=?E.:.=S=O8ZE+U5S0_.T.>L$\%O0Y6P'NF /C?$"A14F2>V**WG"F]_*@[P#
PB/9,%C?*H8,W,B-E[&O360]S'Q(+0#5S)/YM,6U==NI<Q"^*YWP=ACCOGM<1]2U"
PF:[R#,?"!?VOAJ'>C/KJ";W2@5"%) ].BM)['.64PB]!WR0D[I26+D@C[1K7?H90
P'!(PS;&L/6DC<A6U!037?&R-] )/E9@:Y]B9>>O YFB/S2 ."V,!9<)8@#K9_A1_
P*3$82L.CD/9]<I\">\>H(NYQ?7PGP?\@\A^Q3$4J!A6"?+R!\>LHDEN#Q[8:;5'?
P#(@';>21O_LI-8E1"ZDP,JKG,%$1@A>&SJB&'A9?_V>N"Y/FB2ST3ZO;J=)0&RK[
PSQOCRP(@?JQGG5'VVJ,.J65FYZMC"GA"93UPSLENRQC:95C71M!Q7J5-&++DL+2!
P%_GQ$AHH7U^4B@[(06>(+VTYVRZ?MK/P#Z]=Z_%>2$!U2R>E6BGEGR[[%212G$7#
PG;+ARRL!U(Q3MQWP<57-*$ .6T;%XUF?#OKQSA+C:(*\^O\GL7I'H(/PQ5#$?S#6
PMW<TXVP]96??!AP=VNGDDL5GNIXU_]_:=*:FZ,865=_')H5'23Q'9-O<M L]]3Q3
P SLL%"A]_G>M_47-3&QEI!B_>R,/C;6U<^]*?\J%&<(+:0V5$_O?("CSR-.U7="1
P$P^MW[JSBYFX(4":A0E*\<>95]989EYH2:NT1GY^VXBA>&?S4QZ:+/"2Q^\H(3"\
P@X@UI/1,\(,-<KA-@7H+HXM'6X.OO01[9]?I>"\;8><I/2HA*5*,!P9DB-QS5W 0
P89YKA9L>F#^-+MQ36A^-H>/"'RL3=('6.2[3P6B2U5%[H7RU.MH1BO#SB/&0%VJM
PO5U;6*1IT^\5-KI?J6L2@!>+!D/H$_DTY)<B6^Z<D:76<5M)XD7@8:Y@W-';"F_(
PQU=_5(6&.XY#__=(>W7^ F&W:C+)!2_(,4CU'\H&TPJ+_&K%5FCK+VDY<<^S*?Z4
PM&8R0)/8=V_33'Y1G?K@A#%+'V<YVU6#V5M)?'H LPD"E[H!"T^)O3\K3@A"[_S/
P%6Q^L%%O0_BQ(*8'M9;JE^5W8)F38E .:C8!7"S#NM97HX9S;5A,21U+,JXZ?T>Q
P4/P9BZ6&HW6B'9V-_ )K@Q+92@MMQ;BBD9D%:Y2"PC"6NWL)'TZ-Y@VH-=CK553:
P?RU&);)53TU27%^ZP=(Q'AC[TQ0'D('H^;,V,H,O>F!@3C7 1*V]9A?>EITUM&<"
P9R?[P8[[DGJ5_=/132,TC%+N*WBA7%2?%BZX!1);#(F />!NQF5V_@(]%S"GHAG%
PP"_>Y[)$3K;)9"G10CTM:+LZN1U']R7@PS<5O%4# G-8J5_MA2*$DYVQR99,FJZ7
PMV,2$X=*6.YPR]8I03N5]LJ=/\==2D]+4-!C?!\(OU!W%?(D*MR8=2 _GNQSR#Q#
P&?EB><:87H(>&GHOZ1V(='ZH3)'+_[OB=6B>;/XL]&UP"@-^@]SRX7>%NR-(?['T
PPF6B6S\U9(N<P!'-N6.7S/"U5(=$,R\!NN0H$5GZ2$EV= JN88@4:):%H@!B%#=K
PK,#^OW/+8[T$\>A/M).[=O=/<*YG@#=H[OL,>[TI&>ZNQGE02X\?K*2*W_;#?'35
P)+=X$ZK*S2 8UM @3Q88M7WD/W2Z5UPXS#N^76?;MB(])!NEG4K,D=='K">YKD48
P2. <D0)E=X1\6R"M7B<BRO8A 9\?F4$EDX(S%V1[5&FS+NHM%+__]9YR\G=T35 O
P1A_Y%(3Z0CGNY-90)KCH10"A)#*;#0EO]/2&NX"A=8Y8R1G88%/$PJRDZCA1\=^>
P7<$32WLIA.C]DC!@>HW7/=3#G_<Y03+,3"B\:E4CI6A)=A/>5,V,Y;VP"?;:0SJL
PW\=!Q&?FPD%W^.H0 \DK*\#A1RF(G-R/4<\#C-2;+7<49KH/AH=A.IA\L7_.0$@+
PRN++!\CATE@:$O+H'?Q#R8Q*-PA3Q+@-,3ICE,*R3=1:])Q1Y^69KA!\@2C!T!>N
PNIA92[N6B"FI!^\\^2LAHR-S$-^!PX8!F^29(FMYHP(0Z4U,8>0E2A0@4WI+N$X$
P:6^L[X3 R2QZM?]>IG>K)]-_'PGRSY^,&$K\T^,-.]#LA@( #.1KXL-<ER]O5-BP
P+Q&[&G]AH*O:]&2R-LB=H@/M"74D#V*R>^(F^NMHVX,8D)%@KT?:]V32V+\9?7VP
PR!1RT)&7UFH,P\=)Z/0 AA[PM(":S)% L:2&6/^CI$Q!+"+*XO^.Y5A8_[VV8=EW
P4'E3)1I07]1N=Q=.M1P%N"O.<QWCG *DGV]>VEW<PA\%?1Q4>-95=;9SL1;ZG?#K
P&L]WI]3QO.EZA-]0C_M)58VW#_X?X!0H9K[)50ME-K3G=RZGS84:)MKEN(Y#^EA"
PK;D[5U3R>C M6?U5VJJ<[&-]E]@/\X5%")TFLV98O&0K, JJ9>*M"KWFCTKV/]$.
P]2989.A%9"S"5I0INX_VM NW%, U_V7N=<K4.0! &]B,K'_L\J$"H=97.'M85\T^
P[%FQW%?L=EFJ@4IR:C?MST$%+H"8K)P!I=2E,[I3"?>9KC(I$QT;?*VC&1B?I5#T
PBCGHCJX[E$N3I)&GU2S@ H7UE\0=+TV],S'<8CG2X]4*LN^?_0,U"9B=7&UT>#Q(
P1[FB@ ]V\)IGIPO0_IM+ZR4?>* K[]#>O:&%T7<;BB"[IL=A!H/]BEX\I@Z@I<?I
P*F#8W7+*]34!=\?) R5UL+J6>($ \9N<>E88BG85SC/R#/E;4/Y!9!+-P_$P0T[C
PXN;>\^N>+[W!1T'8M$.8W'?D]NQWR*(>[B]..-#B.?8O+A'?M=3 )Z-U"R)6%G\$
PMBNE_XWL-N:_Z"VA[!;WZ\>QG7:F,=W^ZX?,D%YVXC"<=<@,[]@K ?N9]-$4%+LX
PL\9M#K2Q2"&?S'>LQ\#$?Q SGK;FAT^DQ;2)>\F)>1 3Q2)S!PR!B%F; 'G.291X
PF5:-<Z,2VMTF$K\NBTI+$:&\YINZWPMU[1[%CV8//RU*JJAXR!9H\$\8*3*2:CQM
PTA0:Q&<DX#/ FC/*6]F7"-KCI8^E*PDZ.E3IB@*=H6[>,_/06XS8C+57]XCT9A4V
P\Z"6FL$*"D'.%&\C1D7F$YD%W(^\:W$>6)%&B/!W<)S%Q[AZ9<+4.-#&\:!*)I:C
P=B8#2*VJB@X#&G-(=9MX0'M#W-G\&^X6>A$3W^F+Q._L!;R/*(]\[<J?F3TQ') [
P2Q9AZB\63(2M*@UUHA%TFD^O&(9^QSVFV*FD^%16RG^Y3#9=\R>M>X?H:82QG(]_
PE0O+PZ1 MAAL3=H%F9BL4/MTV:@T%_#S/D2![]9L5SJ$;T^ %DFE+JD^Q@JBR9JT
PC9H!ND/[3MY.F\JUH4D6$B5_%Y[QH*D15_H1QYZ12:W:)OA/?4,74_T,OAHC*._A
P)CM@B%I5D/(N*''3-;1N_'3][!^.LG5Q2"'\"_@G@7T ^269(\7$N3)(V-0&J"=Z
P^MEW<1]YN#NLQ]ZP$S7#J*TQP*K9MKHF\Z8_@%1I6N6CM1RD.GIK^:@=K$AD45?D
P#C#@Y[A6]'6'OI"_!9[A#,HU*^C4<NSGQD4Y'"UJDRM@,B^>&LCG\(;J ]-V^!_H
P<4K<"$0P\:]ZRFQ]NBE8_6HD>UGEWOX?LO%U;Q'D]V,I^U:?,9/JQ96?OF*+7M<-
PF*0*>>M<>W)(@51W]4D=G601DZ<M6L&SD)/6DO[,87J 3V3\$)+R&B%.Z\VP\&(6
P33\ P/96A8H6UUSB5F#(@:<82.+K.>&^'ST5<71K2)Q_^-I]Q."FVM@VN(+:]MK 
P9_4[J).+6TN+9X*6,28?T"0U3T3RR^PE#S4)I3;@*$PHP4&>'WSL#9B%&E,0Q*_?
P:T1244.,,?*1VO<_WK?E@Z,8L5,C.OD=P,IO@^3@L(XNO BEK8*E24X(NZ6PWC)3
P:A=&>=Y8+SW^AZZ\C 1DN$=&?\3TP:1RR(U-\J0TX3'I.FL5*;P+;&"-3RRGKIRY
PP[H=41<Y*$$AY8_46"V2%62H9CL5#"F*4'G2(**^MT!&!SZ^Q$"O(],'0R\)S9V1
PQ%L2(<C_H^"S9S@VG<?Z@"$2H&QR!/I.A5<\/XB)%3*3#B6*M^ZG+$6SCMJ\>MZ*
PS$2&B91Z*N4P5.09?V!E\Q XJ]?1O/->&0VU.@?9WQ)!I$"^%5W4^--$XHY26A&+
P$?M^+.MI2C),Y0<?*4*=6DI9K#=7J$]CJ4FGG>.\9>#\$&>BZED3KMDAI(ER19!@
PJ@Y!%[=&PYE>Q_83RY9T]F\@]A<# Y(=OO7JM"CAK+D54*>X=1A&,O7J]R4Z6>O(
PYX>70$G6XQB&0YW'?'DTOD99?6<$^S) 7: EEO%0O1_<=<J+#GH E#4HM!^22$9Q
POHO4C2G_S*PXDH+8_&AB_(3(8GC$@ D"M??:*/$+ '- 80%7H3'6](L46F2--? S
PL9WW[*E-273.%VX"K^M)^-1;I_P&@.49C=*XRFSKQ (%M/@1'V"SZH5&0QA=+96)
P7(SAG'KC"4C-J)3?G!5WN%>]FGD\R=%9K1SM-DLRS;/Y+._0TK)O2[CWC4B*#@D^
P >LL%\!L (XQ8X,%WF S*D>O[,@SPMB'1W]R]#*:)3CHG.CI; 8&SEMB5NZ!)Y[.
PPQ.R [80__JBH$UB@A22:&ZZKRW%AR6!T+JU"'.[@NV'GK<\"ATLSOQC56@Y=.(J
PEV^\5@/7%:N4WTH\%:S[L6$HV12RT.S%>DX^Q?"-M0A+;)1B;8Z/_\6<VO;R+M""
P9KQL5X=4H=TS"@8DF-:4PR AX)$^SZ!8&GFB!QG5E@WV9'5=)%B7'5;]ESMK_D.@
P?7CA,S:F7UD\8&29#07CK_+W3#(_ [)CF$%B;15CSK=-LH-X%"S^'M99.05$+7,@
P[;!7:?1Z#KESE*L^3NTHQ+H%Q@!L(CGCZ5^V%?&0PGEU&*9PEY:RMSI)O0'YFZ ;
PJ0=G(%?^6+&(E=+[60'JG9\NS/_N:W89+'YY\--+9<4YZ'!75IT2#M(K16.*[;4'
P)O)?] ,M^O^8I[Q0U\<IQ9CBOA\MK5*2+RQ_7?%6;YZ2JX%4!40^JPDVA*&8U^['
PHN"1O\@*D2=@'<H=WO/Q*PP0 LIT?_6JV7DY @YX'A^M;#[][J#&)*6N:2H'3G\^
PM(;!RQOPM&JY,^? R#YQFH(!Q&["*#$,O994*&?#[=V^S!&$XV!+ \"-J6W2LE.Z
PK^IBW_2<7I^P.\>N#:767N8+5IOJG.PU/7 #U#FAMQAJ9.Y-R^%=14U-Q4RX9#_-
PMMJP0P%*"A)NR4R#W9X7+A07PO[B D5RK(C<0.GG1Y87DC;6:EWE3?CZPEC[(*?_
PD\W8VX/,51**<ZM:2J>3XT94]!<#Z^9F+AZRZ/7@A\PPCJTOR'%$UZX,KU[FLP"[
P%PQGJ,2**&VRN5#9_M8Q($E+# 'P$7LLM%^;'1O6[]+C:QKZ1^.>$45&<9P'^9X1
P.;),_B.Y@DSP%K@Q:4UV[3( A?+H!ITGQZ_=9.L=N\1-(82C!*Q-6$\UA-I*/U)&
P8JO#R7.7UH(ZD#-EI.QVC57C:.S0LB]H"NOE_%VJK*"I7DK )Y#F)@"#(^"CM^S@
P=E WD(7@JNVUCQ,1:FN[ONU:R[?J8*X,848RKK5EAAN /TXF9EFL?5TEXAC4[)R2
P]^;Z"-I59KCDN79AZ3"9#Y=^?(&(@7Y^@+9Q@TAW]F?2OL4LE6#+OE4ZV)AT0-*Y
P-]A"!2(G,S12"<O3US2AT79? %O?;N.?="6&8C('\V6HCQ\'!F=%\:L[IQEDPUE0
P[&N_&I?2X;[-\'P_?.NS*_I^>93 R(NN<";2QFG[<:3@/T[#&0 470UF34QPR;5%
PD9PA48Z+-"UU&.8@YITBMT4AMMOVK>45]OD&@MCL3L&AT&#=$;?30A1+(:+K@X"R
PA _-M4KG\GRO.@68*![@8%[:Y@8=-QW^W@+["!AE'K,1P7&*F@4 /K"*;6F)TUO7
P]3Y8*^8CH>+7C=7KT#T4;7I"T][ANTF>E%#]^[3F2**781<W(U[\ )^M#.95)&50
P]V1EZMZ,(^7OJ68XODBS$33NL9.N[J78PTB^MP<K@H?R'N >2AU,;K<H@L]8@6G<
P5_S5*!0;/(OB[>;QVM7EX%;4D _)_(8-8'Z>VR\?N2YJG0FD%@@LJ?X2!#Y5('9#
P/1W[*RVZH_I6W+Z.4P&7'A93_X04Q4H1]7DE'A^9ZZGC==KYS5JC^)9 F<.@<V6-
PJAL/=9+;\FH(6A5EX&;BSER!A<R\CD2>6'Z5'19+F>7)! [)J3I;03#P!:A@2LKB
PTMAI!J7.M4B@=E90S1*6R].W04_+W,M)!=6/B_@6_V3,LVS'P>!%#(>3JBTV73-$
PS3$B1!\S\;L) TAQ5M+7&37>$Q[;[BJ[VW-_M,2K2<S#GO?V:7-21#.^_(0GOR4J
P,!] V;%QUR$Y(V 4!P&W@(2I'1J8<03.5A?/_32!IFW2>J8@/Y$>QKETRAL$S ^P
PU(TZ[!"C<!RJQ]O7>;U:8)\CWB*E6@@$UF95U!"DLPEFL*Q#HO=  4$]2T/4,GOX
P9A'W LZ4[=V#8J8FO 3IA9W';[7O"N'LI-Z$[& +C)RI/5JH6ZF2MAFR76 FL'SK
P E%M;@WJL,[D$<Z 3IR$D\(46$>;H]0!T_H69/IJDE8[H0I^+9J/%;=23%BRQWM$
PR014]6!-J:TU4'[86&D#P=<HM;^%C>1@+MRC7M8@_3<Q&ZXCSZ'0BM<>2?&WA8\;
P Y@A;8JO,0/.Y-8S_2_:+/!35)V0?</(#V.2 -EE@]\-J7FO9H(6Y"Y;1^F6U5/^
P&MA$O%&%*U7^^E)=T&X:T4/R1NFI($T#3HP KIBJ%5L2"\0+PCG6=<IO.@XX?UFJ
P$P3-@+H7>51]Y_<<W[.P/0,^4.ES0WTRSL9&F+^6&)E3XLW7(3)$5- J1<.[@(;U
P)1+!1!L:4@*3<"WB89_W+::)P?3BCJ3*+7NV<\U#).-9W=^["X+AQ@PZ:WFOZ]K2
P=L5;_HG%%)X4Q$63^5T!UA'J7UZ59!7.S$& 50Q;WH!A;+##U75 ;/G$U<*%2>:F
P-$"?@>OKX:NQ$@,1X1V5+DF?=,XP4<U?:NBV_K!&)8EJ.]-/$?9.67:ZPJ_6S86>
P/T$C4GY>E8TT-I^= (O6!($%/!OED#TG08Y>_]A?B!&@SQ<5PQ6D@R<BX')OG?YS
P/7<S.&I;Z6:J![O2<0(CNP[L])(R?@[NG;;%)LKJ1/$Y*65]25HYI BQN&52Z*.F
P<56"\STZBS/8SZE+TP/]YM%O)X>ZD(^HGMENEF?1;<*;X0*Y/E>F![E] 2R7]*]\
P_MK<'O\ZC=T@Z9J.?(6NO4%AIO,,:^7*[H(N6RF8:DLN+GF@5%U;,,%Z4TO?LQ-)
PU*6;-])64!23LC7%[)C%>A_6!:W;;5*G<DJSPRH2/R</7^K\JM""3^OZD^:: M-X
PL.*PENN5 ?%EC$8)S78"^E=!2-3L"?)_UA&[2K]>.6@@%WIQG7;ZR)B#0@4Y.22$
P_E7I;)JT,FT6X59>LL\JP98KQ5#V?.%%SRCB7P=@GG>:J44U?$9Q]<WG2?2J5LPM
P':;YZ[T-I>0W3)';),'K>Y[,T\,=)P'#R5W0*6ON:93]1,(OV_NN=-'T[]?9DX]6
PJ3LX.Z&8HZE4DGP5#OG+\(A!M];]F9I:FYG%68VS_HANS)I"4U5BJ)C9_Q9!OST'
P!A1JR7@)S] 1Y&I9\643).HDFQ=V<8ML"T&MM0[0)/C3'&XM_&53T1!'MPVY#HZ:
P23O]@Y(V$B62FBD!.TEG,B,,F> !:8D[?D*\89=A_ODGJ)HK+1$5J>"6Y1C=Y2<Z
P+:H^GE':&@""S9!<KW,%^R-<4^8*G,S &$<]33Q7##M2TSDK1D]GR@ZOF[5M@1[P
PW.$'&@IYP'XU()1K<?*O_IJ"08 (S:=\%#$93C8LHOOBZ-8,OR].52IX'U$3IC 5
P];0NR)L$:F[1WR^4%@E%BP=:K]+,Z=,]_2B1H%A2I"CK$V> 53E-KL2)$\Y9.UF]
P1,JP4@!HW9S ."'+&^N+7SNM5<)UL"IQR4KOO0GB5_>6%V4D?+PT<)0#V4H FKBZ
PIQ,.&*&P.#+I* ^.!2E,Q"%-PLGSKR3LZZFL7#G\K5^J9":EB>3QN-Z>#J><E&GC
PD9VK"S]HI#H:3F6H/O<T9ERD^6UU.=.&[&.\UFB=+1K0#5A2X"GU5S#?<8 (PSWV
P0.W7Q#UXQ"Z9P1Z?Q;>GSRT3EA8"._)WQXW:8)61%Y/C.01"IH?]Z"#OD^Y%S\G;
P)D7Y8XI&J$"U@PZXHF2AS\X '<3<!'Z:8Q1)<XC9-S40);.N+X2",_ B0$NPET/I
P.'$1_AIN4S81?QM/96#)Q&S%OU.G5#15=;9O0$XZ=)66U0=^IGJ4H>FLK2G3YJW'
PL_81O3!D,@E[^1&0/F5RC,/9K(BBJXY<5[IP#XMARU#IYT0]QYJOTP^VIIHI;#;L
P[D2;(5@;\A4FPWDM&P&F=JA+[<HLZ)6XE[R]\!5Z@\.@3C40+FA][\'PY!]$(F8@
P /[:+DF@CJ:0=RF(1"<GW5L29<%)'L&<>,!*TEF17S#;<$?VAP*=19M'2:7^ACFS
P%D@*&1E[, 4??45U+ZTXSVM%XM-_WHB+^XVO0^.2*W[&JG;6FOQ2L*8(S;W+G#U7
P=>[57T,J97ZRJ=1G9I2B+*8GGY:O_,4 7 7H6X/"?U$D.-]/EK,70Z\_$A=<P7ME
P:.#8IBS^;/B^\I+VB#$YFOB4;98=@)_F?^+Q%[.LO;7LJ8'%#IQ(TO^IA8DXTU1F
PC@Z78UV1 B/KXM!8$(*$DEKC\N@7:GS.15M7 L=B]:RBVC8T)T&$7@GUB8E?^*W,
P9T'CBB2^( /X@THO7[JU$F3[>Z862?5';'#W)J\VRV,RZ]KPY1/)$G%E\X,WWL24
PU- Z_O:7L/>VL,C) D\%'!*H*JZU;49WZVSLY8*@972R?.[GC8WEL:G_\T-70-//
PW% J4[<R7$R:3L6F$C4%V]OYALO+6M6*,RJ_ 4M?FH&_JU#*:D".0O5'/\F=,=$+
PNJ^3-Y- WKB(QMIK2,6/TS"0,+=>SJ("J#OM[BC]A\JS=@A9;D[]CDX.Z3;>NI+'
PMMN9!+8G3NU&WULLW[WE_"7?7UEC.;;[WXIFL LY2<%S7SD9TRGN\9S_;@,:U)0;
P96T=R0W$1HJ+5QD;^DE2PQ82E [7<YOROA/MG3AYV %WS#07OG;&'K-,X$^\D<4#
P)PE#B6O7<*V\,WOAN#NO+]D& B>QWAXE7F$5Y[W^"N0)+ +<@6"H2;'A8!<O-X?I
P.['..K^/<="(V1_,@VU-@32"\<(!H[1:^%D<(EP8.$SA/*QRG\ AY=5>>7?$R5;-
P$RHBXH\2_ZWHO1E+*9EI)3<&@>JX3722Q?*/CS.:P^T5VAA9F^N?T^V$XF9!ET[\
PF(Z/[ #<&58O!Z*B[(1+*3J/3QF3Y\STL(G-5/TVBK4%3GVE9KE7@!TKCM:*G?\E
PB"OKIL6,/<-N.Y\PE:LN/[=_"?"N<O]"+'A1?%T%%0Y[LV1DFKZ99 2L6(^>".FU
P?GKVU0',-M&[WX<&=NNZ+Y-F"+DEH#+I.:EI62OSCR4]SA._67LVZ;Y0HD 20&.6
PK^;PV[/"58WWKHG,>:?>W6+:S-7'MIQRP;[Q5;A>G8$IR!I)XE-XSU[ WC(2!3(1
P.<(]^L+\20[)D7AV.< RD-OF^Y-L-Y-L54MC"[O V10=!JY_3F))7FZQ[W(-\$4@
PC-*O) !M*A0,B#/R*Q?O90L+2&N:\KA:I#1PK=)2#9*@,IIPFI55+T&.I+N$Q/+4
PW&TW*")T<C_Z^'"J7U96SD]'"!JMCBYA5I ??#+9-I>_"$@P;<,5@5M; 6@!PRPR
PS%&=:=$:9/"15+YT7W#UU=LRZF\Z6^<9[UHAB]D#QBTTLO"-F/'W1)$AR7.5QZ8E
PUL_5KI_(&$7@X!YDSA3#?6 RDJZ@+V#P_K%[)%8QG:QF9',G.W2M*YIGS/5\B_=X
PL:)$PO[(D, O8EAT7 //:=.K,"T^&S"XR:+@_5 #@5?)L*ZKT)Z>F3EVVX!)*U:"
PG>!V2\R1\;*_&=B;U3/%)[%A=3U>]]0KF#]H6B"20V&\?.NL9VOD]!DX8X%Z7J5S
PS_*L"#"MJM<"V(,RDE]YS)9S>@J/XC_#;FJ2A4;R5X%^",_KW+=2<UO\*S27'R'F
P7L[D"'OJCF-H@UH[6"HRY6TW ./TCIYW@*B391Q=_7TS^>:ZN"/(;T)>@NB0/W.S
P +VM/L4MRVVBM4?I[RD8<U 9I,9YACV"/\$6-B!]$04<&ED9S$8QJMON0$@&<>/X
P]I0(%FLUS*S+2DG2['B)Z\D7;[5C0P;AB#D^1L'H/>>W6;:/X%IKG-Q ,T>,-"P;
PX =>IQ1/Y1)#*$[S!D2+7,+\Q.V47]O.8[9T%(K_)P]#PX;3AZ&*8&!;KPKU[^*7
P;-H>#^2P_BYBB][N.MWR/QI,OXA^[[VN0)#,<M8=/.\MEJU>),&NE"H^EGV2$_LV
PA-Z,E@'M');\,9)WD5"$ 4;VQ[.F!7XD&&O(CX-5FURC] I0H4T3LPM=.)\DRPO!
PM"..CE57FA!\:]NIO-SN3>!9_$QV0@)E-4[1@D:<C2(+U%4'FWHFS*0V5C-XAI5F
P-5GB;$VCK;R,LM,1NGA=G\T]QJ=U>CRLID^ET;I'#2ET+I[BN"I1P';UTZ'#0Y*%
PFF<P@]OIX6W"%"O819F-W*.>I&\;])$FL(4RH>)G1_DR1<#D/MN(]M$6HL54DZG&
P2R1Z3G9C\/A[Q%B*%IU48-B/UOQ\7?%<5 B%4)*!V<#H0.I"*"J^O-#<VQ]Y]E8"
P:F^0C2*&U]8']/5I9,UPU)"@Y.H 21VIQEN;#/8E:@";WPO-,!MCRQ;ZQR90W@Y>
P;RW&@KBGD>-KM(^I-"-<!]H6,@PHNDW(LHI2KQQ36S#&%).+_UYN1?!'#0V +9,[
PZ5-_# R'G$=1,MP,7TII5!$0#H1BSG1S '!WSC\1' 2N/)/]5YYANR4Z\?;!@^I)
P',PP"TMH38Z$-!+B6*$*N3W,LXXSX-PTW,Z4:6:436FELQ%/0TUD%,*5[[,2'=EE
PXZ3Z*)TPM*FAY4WD=I(U2$CC.,);E'9&S58?,'Z.^URLA44Q, TLA S?X2;WA[KY
P%FV3\[4WM2I(JWA4(!3EV&ERMN@O&KL =7^DP+!.)[8?S':(:!:\[9NL%R0U\>4S
PI(I18[O$IL-@YB):@$OJ>@=A.>SK87T6MSND9 R].>XM &X##>F% G&-&DXJ#M3&
P%NLG^]J&38TN72B^$E4[Z#;]]S-!?.SDWE0C9\D1>V/^O91F:<X^SO! +R9S5+=X
PC=DBE;PJ1&NU:KC]4%?F9D'K87QL_J>2:[2KX&]2Q&P  ESR-)AI^RRWSJRMOIQN
POMU!3ZE3QP;PM1#I 9PU@<D0PN77^^ M="-W[ZR'0.LY$ZSL_[\1.I73O?:PGSM]
PDE'&E$'TA&>VJ:9K1ST'6$"+7!16"VA\$W[QB%,J<>LI6HF\CKCB6X2!N+F8:8_I
POE1_-=?3'/[5/5]<DB>=4?Z3>'@Y9."#I \!T=01SI$C6O]S1@:M:)P>0AK:[<EK
P/+WA-Q">\"](,SS&.ZY=@G,L<H*:P$^(LPQ7O:"N"V+-T[$][$>OTE\_@B) "%:S
P:5]^X7@65?$=D,L,F,D3%?[FW6+YH]PP5X(J8IN8D)0YO(&XZL"/4-V,-L&4>']E
PVZ6TEEDULA1,RD'8K%>XML/#KD6ZZ>(#E;X^(6/+$0(3@[L"<H-%_(L/?$MAMD;F
P#M34WCBG[-PNQ48.^*IQAAJL\"G<P6_:6%>+Z'Y5M>D/:\K]R[Q%H#JS_%4.??-S
P+Q*JM#D 'ZN"N-C*Y8_(Y)E>_68T7V^*2=PV@O+;;,>%Y$2E&;UX!1_0R%?#3Y8:
P!D7!!M#,0RH.+H>%[V1PM_= >@'A$1;?;6+1;OY[[JAXERS!E5/"2 _6!Q0#IYD^
P$ 0-$X5,TB[#^"^!)U^,4)7TZFW]F8Y!_/R$0G8OOBKK+1N0I%ZHE0?56]8Y"EWD
P7%6UF+N])WKH7U"SYV8[_='1LVX#=:B?=X1>S15'D-Z:DN8O\VB&;;JJZB$ <6S6
PQ47&$+X-[+V$>H:N+J!J068*$17(:M)D[*U9;WED/+"\LQTZ4O:2 ?9F?>)RQW:K
P]9"_2C6'7A?+NU;D/Z8T$$4*\_PQK!%Z!%_\N?E+FXP\L,O3J5Q5E2,1(U6+>&53
P)#)R](*70_Y8XYZ;%<M# (-H8>V5S;SRYBO=/%%4?G]=@3YO!N'V;L=HG(>)7#?Z
PJCI%38W/,&-*"G5F213;18Z\W]!%':44T1;TDVRIG3M^%Z.-9;Q@W@;X">*[#HY>
P"(Y27)>L'.*\_LT-;TXPSP[%BA='??(V^CQ=>]J_75%8"=071!RVN<N()PFLWA0V
P3-!$AS^/[;Y0V>PT=6E)%UY09%A!\TRE(!6@EODDP;]X<3[Q)VA4"#M!TW02OX*#
P5UO)=[-%NIS PSKW([(WUC:+<$Z+4H&(J814.?*$*;O[H@E1,P2C!/9!88B@Q78$
PYDO*#F(DH9PV#7G@$H]FI9^2XIP3S/.9,$VS.3.(0GEC@@+/BYXT0/_M!YM>M\\.
PRJP'[>"\!C*/%L.PR^EWL)#-Z8<!^I;+TSJFM2*J5[C:?#'\VT0RM2ZHE*'4L0I'
P8$F.=)D3=TET[6>[KT#H][)9/]GC\ .0/V*OM\GBVJ9]?5#*-Z"2&/ +UT]P(%67
PCLY9!T::/->8OUK86D+4EC3K%W,BT [Q. NG?6--BAL^0"1% [*3,U%N!MM^OK62
P4]>M)_J,7^"90 K!2 ?ZEYY1&A O22F"*FR5IHUJT/*A#-D;UV:]\C2Z\N:_@?F.
PG ?(?W@<IF0S8/VN5G_EZ0?\&\YJ##1DDKX-<L6$?CXM!;+2S7&B5'\C:%!^TBTT
P3-BT?K@EG*9,>EC:=Z39*P/5&*Y84WXW1&B;J=J?%#J&G4759WF\/%J&FWMO>Q99
PA-L;GJ%J#<^M1F?T2;@LH/B-9TV(MW[>[C>2/U?R53[U T>\+K0L03/PT>5_R&5Z
PJ%Q$>/<M671Y/E\@N8R:? 2FI8J,5*6!Z.6W>J2K5]\I>V1 -2/1UT;!DMDWS"W3
P][$7O:HJ&H_9_P31H-?%P>W.,2,PC3<P+8I)+4,HK*N^C.V."E=S20JE3&4AE%*S
P/[!#W[$O-E\8W+#R2TG3]P+5^\O?S-;%]/"E^HW'K[1'9RAF "TJ=6NIZRP)+=.R
P^YLN\]I_;( >0/\TZ4X>@KVP+523PND4MOTK5CB'(<E:%3G=OJE$%[9-\3#U"B$L
PJ8IAWOEN)^)TVUQP8.Z8ZL8R*,CJFT2M\-&#"1D9G%PK@^\AFT'&$[92XF?G+'>S
PQS[OI-R+QL=@([%YZ9<][]B]RZCKC!ZYVBPI/.ETX8PROQ"+-[PE+IM30V\ AM1[
P!(!2Q+Y2 *Y 6=>S]1:=C0C@95LN5%R8@=(H;?]I-[DOT/^OJ_7\]2]=I#PLL.+-
P"[6CJ YRI!Z((L>-4P8CV%%=4*8]WMK&M[CW!F)K%"[&6*ORRMNE<9:N4?0"6-J)
P ?7IB%O8D<R>4X*Y-<C^ VWA!4!6ED6YH!$V[W[C#9WYF>%; KF\KU(PHOA1YA3+
PNZ6:0;OZ8&!O>H/KE"LZGZG'MW2KFGW(B&N(D;CP2A#DVMB1W_=?ZG')B%)2_2>I
PV+"ZB(+)<$;Q3R8X[505C#8,/V;] VZ[)V"MSXJ=)2.J/N-<\/<_C*R.5T9BV+,[
PG]'*W.M1\'.7\U;XX^.AGL;YQ#7HB+[Y@"*>Z8='W>7A@SO$AF:?>=/7_9^N;/6E
P]1ZF>E;"OX_ZF_R=T5'9]!M[Z\YD0HD2A*/ +0-7G6H:V/;.ZMGFLRF= <-'_KRR
P&^UM*T=J8(Z;.0R2S$EPI4YL4>)Y!"_4$:>%"P,SUWH-%(0N63Z+F&%3_8OXJ+&H
P>^5-QIQ]53",CMK"?E!@]#8S1Y7'3@*#J[WP* SVQ>:EU2NUP@[#L!EX)QO(_ .2
PV".PO#L7<O5Z&SW5IXV56N@A,H82PYG"+7E8#P1;_"&'B87&+\70?]S;(DQS8/0V
PS].6.IS$G?[A%E2 N:%65XS9UXRE"T3Q[4C&=?)NE]0'S!@K=X 9KI1@/CN&&@85
P)TL=\=C[4<D($H&ZU,.FK]7&_2&5T4XP9M8-[IX,9C+]87Z,^($K-<3&0&CT\=9#
P]&&!A^1V+(UV9&VI26-V$TR=E.9WKZ2#C%8"YYA-1KA)E@'^NS:/V.0X>?Y(\Z9B
P>SC1V]:@VHT)!'KK.ERA/+M_B5T&!(G]MS"?E84B0PQX)?A?@0PP9T:+F["HI!8*
P)Y=Y-'^<F MZ7-_D(.8;22^=7/!*V/L9C6"CPA:GWDK" LD*H/G%#5B:FY74T6V[
P 20RBO:S6E?Q+JPN/@EA3/>1U><MT<]Q6-%[/,X;[N\_+D;QRTL-;$WJ$;$U6AO[
P_3YEYB2QBV:XH )+8'EQ&>KD78[A+)8'[,Q9XE)1B"H-%ASZ_8<%PMGMCRT%R897
P!R5]5P*-'Y]"2:/T'9Z ]67]_?M?I\T\K2LB1_B$@Y@2#O8!QF(1._/NS]ZJN-UH
P2M2!K6]_L91,I*G1[HFKL7[H2+-8 <C;C0G<O#IX(/,65I>!N..D#.(^WZD]2#K]
P1EI H_HE4*Y; E'S,774R:K6]$BT>2:MM2@YWAY&9G?E,;M(]Q<W0*- C<=,5P_F
PF>!^Q:%C#"#=E8:"P PZ9SFB8K"4\5(O+;%[4A=9,0?9O^F11<Y]A?.M4H=1EF5I
PY-[HG&51 7"(DMYC&8"BY=O",2*6S,W%KV^]D1P?TTMB.TSZES,$HX-H-$2C?I+E
P>E9,Y1E.CZ4_":*=7KJ;!<V1E.$L7CR?)F77.BH^TE.!M--FD.2;H9DQ_43;Y#:X
PFX!6'I;[,F?N^E*8FR@74"*Z>NO-3/5\)/IE;U*<39H?"V,QRZ*6?,&#+.:-1D"/
PR2#G?4(684=KP)/C*O96F./#ZOO1==(>=92E?_M("$P85-H"CAB>TP )E>32Q51>
PE-R.&:E8*TO+^$PB/@,MFPX&X3:?D;W4TA38B%)RR!,)8)/H+&CS>*/0@\BWM\WC
P/[#Q=P"+XV&Q-EJ0<JJND=PM=N[,16YM<@$<IQW?#?1'U%=S3(>Q71F[G!?EK[)I
PZ)'5P%8!^*IRPY<5)8!&\EE7KXFN79=4+$V!:'CPW+J+E%W2DSH#X*E'%U?!H(LV
P8GHQQSLPB0\9FMOH5KJFYT7<VX8-S6H/?G?:.K%'RP8RO;AAH99=<O"<:L0GP<HG
PF&&;!I6_S4+1]##I@CI%82,>-S5DMP[2_9U0[?X[JHLBDZA=*4(N*$SO]RN4".1I
P*'EXXL$66>;K,Z&1[24.CN#E;W;)9?D5I>I'3_9B%3+]V9X=#PUA-I9'*8LIP.VM
P7Q6YT_$@2K,WT[NBD<B6O4@R[&>YZ[/G6E$\.:E ]O;&A''Y@2\1@:<4OQD<#.> 
P,E,KN7N\A0O >A<WNIRSLG+MZ%Y> Z!>"<WU 3FI@O>$4;*:H=7URI+#;X#II*O?
P8HR!6-S55>B<T*HAB-?-0PKK0MJ5A5$A3H!_3.;_@>'.5OW? KX(H,MW,(2R-]' 
P3T2RT 0=P,EC91JW['3/G*L>M4J]96-^N,A("PSH.([4^()PCF*]8$B#*YX2S#AT
P1PR;4$X0)&^ZCVI4G$<S=AN1;"&=K-NN_99A>G]T(3QX&UD]?(\HXPG1S(ANA],0
P[M(B!,(P #V0T+]"ZC([_7,Q3K4:G=NK33G%1:]:M0-N(RYVV''!P2^99GBT0BQ7
P[0'E*.G#67A^,J%<VGW#4BTY54Y"?@^^P[W4,#N$*_34M@IWIIGW^?<701QU5#17
P)K?-6<"T L Z<Z#%<0OYFG;XRAJ@_%<@.^1-E:_",%BETH<JZE95Q8D:3HIJ#2]O
PV:J84VZ0Y?++8"U$047FEEZP:_V'A"@%RP7(K3"&HP$<[(9W?=C0R?$%W*FS9WNP
P:5K*4Q6-T@1>!6; EA)_JK-VCIBSX,E>YP^!;>8BE1==I7WFPS5K#]F_.[O'I44^
P1=Q#%.K,EPY#/'#\NL1FAX<JMO^$3J(M[XRQ>%:K)F!L FEGI6,+'TSPGL7:0KC[
PWY\MB]I5M=R][\L_)HKU")L8OY)9F-R\W/M?_B^7$,Z3;8MK4CH/>!/^XF6H2?UX
P$D>6(W2M9?T&FGQAX5YU@=UG41XSGI9(5Y.0]4W -O;:)*AS^W318QRY-E(W( DJ
PVQ'/1*J0OKZ82]/#RB*+74K+-C^6BTQI:#2P['_+YI2$9[@4"JIGF%IXJC; P,(8
PZ*6@Q:OE9*%,Q:EU20Z-ZVJNJG<<[7V>-H7=SP%ZL5%@2V8&FA@X4C-N64[+HHJ]
PQ6J[I7AP:Z'IV\@^^=R_6%S^$(FQ8<O#PO,E+/=&"H'+!H%^<W&BZ\ SG2DQFT<H
PS>M:T<.[<Q9XS_(=EN<I:#2&W7E,%KRHT,$I=697WB8PXW(;39]E/Z7^60DTI7*I
PNA4AEY54C$8HK[TK?(-^!AF]1@EE\GEP^2P;.*&XW8I#7LC]R]W,'TX<+U5Q8 *Z
PX8SNE><%8]BD[=KU# !Q=#/-[8S).)]:*1<V/2T_+1SC5-WY*)#(7HU))&0M%!]E
PQ#%DH1.TROK\Q&&CHD4(WYA0 .B+]<XB2)!0_+1<'NQY@-D</W7E"F$J[!\5'F2U
PE($!4F(\'GUP+G*&RKWD:! 3&P&.?(ML^/!XG86A4::4QK5YR=]< _S[VQ[&*/L#
P[#(G>;:SDYVK&)1"?K$2="33D7INH4]+\R\1@$<WM1QED*MT*[(PHR2PUBNC7=#-
P3:/(/>!U_MM*R8W#I#S.F8@$V7XB+%R6<<7?Z(*KKJOZ\3]3[V/]LHTPKLBXTSGB
P_Q>SW!ICUFSZ5X!O0Z+:R:6.E7OFQOUM=XU95/(5<XN2K_W[ 6TN9LG6$B>E/8X 
P2:[?MT(*.$ I>:ZUBO3 *=8Y8ASO*KP),LO,ASO3$%W7B$" ^L62PWK/XM%A2[["
PB1?5?+]YQ6+2!AO#<A\?EI%1QFI?NMAJ<+6QQR320#"*$O&M&+G/!$5$K([B@8N7
P*J"VUM. ,7#G,;5T+3KYS7:*(%^\R^G?:*TK0 VQ'35Y%^>5A%%1HM"K1/#;303W
PGMV'O<0"DEL<X6_"&A81]'EJT N]4+,M"QPMI!Z75?"I$EV9R[75R*%H+-156N+6
P'<"*R:#=+F[G)*\* (K]N?,1!UR6T7%AID,$LI\^47Y81ZQ-!+LA2>X" ^,JZ$;=
PR-TE+_3UB#*WYK88$V%X-A$U8M00=GJJ5,U )W!^;>G_Q4;P533;)?'2X3=ZJ]=Q
P7X#W_KTSA(S-E!N?4ZN2%3GXAE_X<=-Y.)_[ALAVQT4G24?L)]D^@<H#W8QC&K)H
PC2Q4UZZU/3^7&RFIPQM\:V!ZC87.$%4[P]-=:OQF3&@DPA7--]MI>TU':S+>P0R5
P6T=FOTZ,4:M^2-+FF&]D' I.,['L"TMT!XH8).F<W FUZ/#'O"9_"^OS*_1.5LTN
P@$_;:W@]>-E.+"Q3691^>),X%H=+GROC=><YN],HZV!$<G> >$)MF7?]/ 9$*\;L
P>3KY]&Z6/N#D%.A:D=XH'*MR[H)/7#U^/A%2YW0>>$LL+7J:MLB"5C&@"WUDYG1D
P[L6?UV$=+*&]NO!#G1+LUU 6;AO3^)17 1.>;HLQOVJ,S8>,U)R0:Q\IFUA-?( 2
PQWH7[ALA)IJEJ^7RVJY0;',]'-Y3!35H2;:_IIO*1&M<  E?K>^CX>L(PT@7@W.8
P\&JQF+W"=/I-BNX$5K[[X%>5W80FRTYUA[\Z*-9T=<(/K=>1J8V:S!+8(&KY_Q)&
PI%%L?'7<X@UR@?;^ M9:O71NE\*'-W%DJIXH:,ZC%8B9@ /JHBP2I) !5^7-D^S!
P.#FEL]+5<_<C=/CV.>A?)=-P'#92WE3)NI%X@)'9B%XUPOWOX5J]^DX_^E5%<3R'
P5C]A;E,\NA6SG_BTC40;?K;DH:)M@-[3A^F#IR_*2$V0^$3Z#H Z=;".30IU/$)N
PIY:\JR8D.H"6P.<L\&-7(^7,C.>-'A+-@>$94LUVOL(ON?6Y7 $(\E+8FBW5^9Z[
PM\=7FJHA2[<VHN0-/C96("Q7N6<IWVZNF'0/X\9<G7+C;, A<9U"AE#DR8X\AO_0
PF6GI#<6UD:-[Q7CGMM#:IT"R3)@>E,-(E2-*$Z)#'Q I>S[=37WR\,9,/]AU*3VX
P=XC5,OS<E6=#&)3F6.5[Q=2!J-_73_)DXO^O##Q3<U:\I1<12)F>&"^(7*SN_M!$
P&!AJ>>0%&W*%Q7RL&[%V-P!G,R#*04/D@$H_%_Q\0>6MDLII6]^WAHOD[<XOO6NV
P5JO1S SRRO\/J?,U>9L-/F0U,,8'YY/1C]9SUP"68?FD5'JELAC94-"*J9V]<&JC
PD<O27;"(HQLNX])X\"=E%X%H5IQ85]6),>":Z<N(1$I-00E*9QNIC ]QM$I9!\T!
PDM;PW)&\@OX<V<JQ!VI &_)/.*GP)7C%7F4?6(,-5(S0SFJ7TRYK( )[-K.1,&Q>
PHR<F^O!G\JFG7 $;QH6^FJ8ZD]'M<<17IQ1T5?.]A7.7S)-<VI24JY45E0Z"_]:!
PUS1K[H3BSSAVOLMNB;[+)N-G&G6K\BP=P'':5A?0>[JVN7UZ:()5)<.N/X:P535)
P9.-_Q@G&U'T3&8=F4;*S8+&4O,Z\)47:5Q0Q>WS->.";&PUE6Z/[H[M"\E-2T.T$
PVN0(B*S;DV7B:'* (4:MZG$8XS<2/E1,+B[%I:"=QRTY&OWY]9R1'/S)HF"T/B+-
P&HIT8H[FXX3YMS10+W(E@C?&<@4 ?N@X3VHAQK6Q**>\LK[R!.[+T'IC&^)BBES,
P ]$&9D:1K(@99*'-A#47(AL"+;KJ#RT^=Q6GW[Q2HI,Q;&DKAT88+#8@_S%(Q;5:
P'O 94 JIH<\:B+JY&VIABZFG?QC#I=JA^'B6\+$P-S("&V9_.390E:E#3],-G!GC
P:C>VAK;-CL!!3L#T&2=U)7'9M;UY[9O#I#,U6B*! W6;-%F@]Z2_]KP#FKRBH@!"
PEF=$@I51$@8OPEC<?(RH:8K_>XSB8'KVV"(4_;U6?)840LO8G:&BUPMM$B32EOUW
PWFLD-X>].-^]C+YW_UK8SPX@K6#PE1^-T3 "#GWF'(*W,O%Z^?3Z$RWAH?G+IC'M
PHPLDTP[Z^)%U<C@[:<Z;I(N?$ 9S*U9<GGPI9 )F,8K&^0>,9^>D9?CBO$'L1W88
P;$F;-4@*GN#(;\SMF7+L4PQYM+&G&'*"%Z%$HL<UR%M&Z#-AFG@D;V1G^F1+9Q=Z
P1.6/O\3E*&@B!C3>D8)SXQ]_AQMB55XRWO=='!YUF\3O]ZT!WI 9C5OI+-!7[$Q8
PI-5\EDRWRR7M36;O+&*BO%;1?809V:KFM:=3C=!=@1/]PK*G\P%>! K!42C64%!G
PBOWRLMEZG*:S0SX:^$UJM$E1Y .!77=;OGC5T. YR\V9:1RAI32,!R=_MDF%',,3
PK$9]/M(+^-@S AM'30Y1N?Q+]!3?GJ;GRKDI7!V)"$&R:??!J> @VI".S7DZGDF 
PD'<2%YCIW.=TM-$5IGOU>>]83I6C#S #9R[G.6JA2D:TS^5E(.P8\G9JGB,-29U5
P2?%6O.#NHJ"Z87,_2D>CMW,16_["PE$<RHYN@[]-T8-T^QXRN+E-Z%4]'95&=WBP
PA:+@)[EK+6L1:+Y125BZL_@B&Q!=#^'@>41/ZN73,#&H7Z2:]$K5&K&AN*V\)&9+
P95#L3I+;E"%3Q"*<!& 0"N&,!+$$.SW6B<@2S.KR9B^/H6[^8,+W2]-:HTY3FV*0
P%H(I7<IJKY0>AHH=N0)U C$D;]''=V+3&!?^VYY6:^%ISY0G7(V%68P%:44:_071
PT8>8]E?P182HXV%)#IB-O>0\OC2,\+4NC_13RE,$N:F=&('W#50_3';<.<\P2LMK
PQ(D5IKY'4$]MZ)Z!?[*"<MV:0)32#'%TP-B#+%4J4FRGMX4#R#J!?( ;#'![7V/G
P]DSA_X=$W4+D>PESMDK/DF;QYD\+!63M<Y,KB@VQU@ZDA$;:0# +<Z8B=5J<C'D5
PS-&)7Q VC^,K6)&_L3H4I*X0>.T:_0$X-ED/(1K_9D5RI2(<@2[82B:SCZ\XPKZ4
P\@REM^[YH<J,RW6QMAA@I84^6RF?/&I.1SSP3M*I7!K60C+'LMJB(B\F!176.@\O
P/SS 4[9!X>X)[JAN?%M'<M2PR'0E[_O?(C2L6)Y*V?H;G6P$VX S5QZ+5XPI9:<4
PWQJTNDZ2M1;[<!227 MO[=/>YZ.$J[3:U$TT8U0_!8SZU$17/_I3![=E7;:7K2W!
POJZD$%G56$;$$#5CIDV@W] 6D/ 9AX!B$R_<+_MA,;Y9?)&*.@.P50;%!3EK"<QV
P;P<([U1YJ'IJ_8\#:#[BIFT-FBM$\RIGF7===YOZ$:GY>DZO&Y:UT.:$I4UEK);1
PJ*=^I5\/=/4H07K35L= #)V)R/MT3]8ELC,"J:B4DP-+@VJU7>$,:_8PHPBG+A=]
P$@]Y 1N#7=30AS;S!=>/Y7C?HCCS0@^N& 6?^WM"BD.Z2W)0TMW+09BN(6*K:.G0
P-16,.?ZBU74RAGTJ&XQ#V66%:UZL3Y812_-1QNQC-6CC;&OV3[DZ%<<BPI3.1]P;
P*M2+@E?>F^ZKS3&_*D9.XR.1:;[S@=[#E;A9.@R!:R.'OT\P/)MIX/M!(;_\GMI<
P*)MUB=LRHWQ@:T$;D7U.%A5.H?JI^RS7 "YPLYBHYB*)H:*,=QPH-QJA#WWLLSI7
P "/I5]2MG^.F"GX-ITCP4F=\/VQ",KG$X#[Y0T\[/VUY"YS5LZN:JZ3>[)Y+#E"$
PF5A:XF3 &YH\WVC:/U:QSNG]9/AP@#&&7ML)2QU:<1$HYD,Z8E;6_[4"L,FBS?Q_
P4<L*<Q+@]-'X#^*4:(Z9%7UW /SQ.>._7U!T57R<AJ]0^K<V<+G'+F>#Q7]GS9L8
PXG!Y/8PJSX.%?8.0W4Q5#QHE]!&_;5&4>9!L<:U).;B$0;EHD>#)QJM /"[())&S
P9Z4S^/T9DTBB.9M+ZWH"D-I5\C!W/<)2@/S(=9B5NL25@3-F5(H\<TLLEH:'F[<)
PPS;=Q2 /.]":#+?"O$[67PAOR#M/,6OK:4N*S,V^ 5/L!& 4H;BGNJJ7S=EI.,;Q
P6-"V=$= .#BHDD9:-FH;'T'&+<-'Y3]R]J[BY95YT4(&'][P8NE[(*"LG"(Z,@$+
P"5<"2]ND>7@[LS5XD@F#@,\<JA5)CK)=QW]E&Z;D^/;X44(NE"%TP-).N.96S@ W
P*2&9"-W*UE'[YT[01]ENH\(F 9+97+]+E3>-W[H8SXYW^5J>DQ2L@#4F?AC2$L1[
PE71^:9V30:8?0O+S%N8]%ZZFHE3%R@8'-Z,2FG&ES8#XYC.W<XM2@=ZR^$K2U'E@
P!J%_;,3*IBF\%[:N%N*'%:A?SH5!=+&3'YD -3NU^37L0=H 6(+ZD#%F.%>:]92)
PM1.9!0J^Y&H]I83;%< ,=-_J\LK4W%>+#BJ&#*>K&V #SSAR[J;:C]/)\][I0&F[
P\V_QN#=&%%.!J>DG9]6*P-2SUV#0D->[8ZE;^*)D8,$960EKW'2?FP7\;?82],&F
P5'K PXZV1J]9!QU)N\<,7 MA?UU*:'>CZX$KE).&N7N8LQAL8Q<3]?0>_C4 $POX
P"D-2N&SN$BPAA80XQ>Y%D^IP\B#@;L$I5V)@WFZK'O*85HYQ5H0>,)FZ7%S\9(/_
PTBB5XG"55T'IMX<>%@^!%VHNJ6^J)/6DR3C4D^EIOWZBAV(2 78"<\TMA/LOU.CP
PS&S=?LM1UPU9IW<R*F/:):!G*>+9'(=4M(6Q=N=V%%7'X)96D&_S#MK'2:EP(0>R
P/YW8$1EWS%Z&E"XD="L(WF<K;7/>4WOJJM)!ICH=F^6>;NR%P//?JB>EGH0S>^=U
P ,18I4*19H_^9+C3O$6IU"7F7:I#LP%E\FQV0>" U%2>*/3J[K[C_+3B.-K  _/5
PK8.W4-!^UY_&VM<7GIVEI M#I  XR[FVAHN1[JU8+K%S6!>7)%'P'Z04BZ#0),30
PHLO.TL@8 9R#-L#!F15)K_HU7$6. 0DTCA]..>DKM4FD<Z6<) N&"'$U_R-C'\U!
P3PH?UWAMO7N'J\-L!)/@6G\\"KW,$O&/J+QFB+W .'; B;[VTV8OC"1G>7D"A#?(
P'U:<X04U?\Y:J@\IC3&RRZ+C7^NY#+V?#0:O<EVMY].DVI'?MY-#FLKO1/WB-3 ^
PM2-Y\[A_O@'I%FWM%.V0:P7GB:+X$FLBZH,A&:VWF9(ZU3/&"+'E$$])\"[(V3^?
P -[L$=#&"97Y6G##S,/)6#!W[RJQKWXV.WQW:+MAA5(BJJ4PM9QOA66KH27N:KY.
PL6K^;*(?7 -ATNE[T(@FN O,LUNM\+R*?K1>TOHP!8L+4YH_[5 O>>;>W)F9]O*>
P\Y.8Y\]6Y8\A8<3 J2I3)7J!;59:#17>*KT5,3!/+Q9I5[FTQ!*^L(ETF\?GV*:J
PV Z7PV7*\6%+C([</7PZH^*#T+R*5^/"HX7!8Z\%2';O7S:)O5A1WI2 6#7\?,OG
P#'#2IJP83LR7Z3)$5\>8P9L#*?^,3EAJ?X2U.J1NRPD[;-(Z/^AA>'#&#E4LAD#'
P&X&>PS8 1/D&A[*K5XGKP2+UUL]C&!# 1?!0R'B8(5HE+\(&A4FQ>%I^X!?"LG'R
P7?_UZ;W5@'L\^M=ELMFMCFQS[P=:7EIN=+**#E9^4Q2EA(\!L"/&OS._"M?(YTL;
PA;VM!JX.E(^""4,<*:=BO=8)EL_ %BJV3]O^?4&0_M&\.(3"Q9N'>U4K[P&56KA@
P+$TX10/F?G<B _)XQ='5V(/A,.ZIK%FUSX"!/[0PGE&7@(C2'!X%+WF,#!O2F90&
PT!X/JLTB:/GHFD4#BZPD1&U()T?5U7RB1\\_9_G]+4 >/'#O#UR2@ "M887]E?:V
P>'4!;^AEU \"JJFP5R-:23(T8$@<W3T&'$(C[7\$ME*S%MA9@0YM+%NB&A2N8W&G
PQA..$I_2CW!YA'<;9"^7O5%L^WC33]N,S I7,VT%!8LD[$,$FTKVXCROT=760)SL
P2 4X%TN,WE(3LI.%!E]WRLL\JL'$RK9TI:!3XD>.>U[_T#X&8(65$NE>S4#W!6I'
P1P>ZA/V!X*_9=X!U)][.F@B2B*'-6M/A BDP2;*%.U#]9V_)@-A_9M[Y.HET6,B3
PBN @#FKE>0$*$<OGP /HM82/@", P&10T^,ASWEX2$%C?F\+U,ZR!9\D8LTF4.,W
PP*"2=[RZK'^C*QM%"*/\>Q!\2)5^,K!T -]%FAG# E%>0].J9>"XR8$\%FR&#:A,
P<43O-R$^3.!<]6*1;(+J0'T*,"0<NJ>;"#<\;UNA0>3H9US\6>-2"8\$2&5"A_/P
P%^*9511<CN&^@7^QM-8&&,6G"ZV4OB@KMXE9G(@;XQC1BYDDR5CMWI;&XF[LXJQS
PSQ]0SD0&#W>94>"K<[*0..4OJ%</H_-?(F]8O)&9A0B4W9%ZOQSX<>-$QS4A#&JJ
P/L@NC% SZD- G5IC_U8%9B<=J&9RH$>/+<?$-^TS#D?RQC'@[:PL68/#O#)+<C"=
P=Q."BEP%D)G1]B" NB*',(AF6!>9]7W1^CG25@RV-HR\;[V6/O/,9"H9M^VATVOR
P[$7([+#U)O>"\&37Q]]'0(TP;9W@[TB-O,HX@XXR.LD8>_'4N9WJ!&.-Q;]\S3 G
PO/PT!./?3!@+3DPQO('XT9CP['*Q\\5R5$HVL-DR/$NZ(:=A@W8P<8Y.63'GBMFV
P*Z!^]MGA1\"'?S<,34) HZHH"K5\@_\"7'<3]A;XQNDZ5F--^Q_JD.6)]_'.5W6*
P:7'G\S:<#QZ[S>W FF?C[N+C=K\G9+HN-SI N*HU/["?B*Z57Z-"X9E>K$3IHG9(
PD=[9TA!:-H*+_MJ.\'.63;#S$N/K=/VMB)K>X9('PSO61 E6-:PD]R>$<G(L9J]U
P+*K+I>#V#VSV@4ZVO I>4E$6[7BUVTJR.O,ZW2%G!\B21Y2:F=%'S9[L,?FQR\^L
P$2X72E]^ILY1A3O8VR=FYWIG+NCLNBI"9NFG4Q@R3A>A1>V9I@N('Z;P)K,P.DR4
P7I$N**>\!ZUN*H35Y:C(D[P/<D^= ']$![9Z O7R=(A0@B Y\:9MH]A#[H&IV)70
PSS',DZ1T"%4&;+Q?O_H.\#<0>(G*70P$LQ781N,8]=!1>PTAT;<(F+90W'OC3*)Z
P4K SH\<+O7VC^%;-4L7O<?C3]S:$_(0M*:M /"X0IN ]F=L5O,W@F<8*$24^P4X]
P:A 4:HK(^PAETY1J3LJ,7FACWTD1%F-U)*=!0W6<TK,N+R'[#BY5[^T 41PF+0K 
PK;2;!/,!/?V2D&>,5:$\/7I-P78YE*30AK5^5A:0OYZ!"CYDSQWN..3?4R\)!R/V
PV1J/P%-F*QNN>YE*C4YJTR-#>$]WYDB:>DXZ!) TIT4(%H\=A'Y)!<DM2.NO@-8_
P<\7@U^>C"V!-8<EN1..6M[[T(>A/?[+,7P+BP_/9J5E[O[R_C:U]]?G49F#M9!R"
P?*,RPD_G8Q,_&:)+LT&EV*(,%#&M5_JO@,ZB/($-![WV-E47WX!/)6C89V88E2,0
PC^2BZ,6E*\O(MU?-TV$-U2]V/,DR-W@:PO!C+[[%8'A"XX9OGGIO#1B\'@OM8GA=
P-W_#=O@6L'_%?T22/8WW5X#05I![ZLI>L]W/6V0F$ZCQ_$N4CZGADD5DL.]^.(5#
P%#U"\? *!/QWME8?5UYEA 4H5EO$2SOH TD3([>@Z!RFT5MPRY.<MB^ 0C=>R!<X
PMBSI[0 #I![L>EQ2<>X#@9)1@EL480MYB&9TU*)[Z$S@> 5M_I(NH!':T[\H2A,]
PQEKI$_H\2#S64=GRY [%C4I :#'D)XE>QI^GB<&IS;0\+.G#:5S,_A+%\'K.K[?-
P^ CK<J1\TT96+H(F DR9\#']L4_"3/$+AQM?E^QV(M:.QM4O?2'<1:J7=N:L9(8#
P&U:TF3?K1UM4."=0:H$;&W5@JS!+R5YEI@QFVNV%W*<PND*W(3H_Q"",DS-'M,8A
P=CIDQFL1V)H6:#N5Q+X\<W?\*:U<!L)10?SS^<PJ$J!'Y#AZ3L,V\D?[V8:ZCOGW
PCI]TI\Z1GNZ<LHAS'^\R0#5)0] * 8 KS:@D^0;N@SZ2>GB'7EY!G6TJ]#@0A5Y'
P<Y(![<I3P+RB$5,:-\,D@'UV%IW:3H^]I&(58(W1"E^L<]^O4D$II-5(VF3763C.
PBRE6G;R46)CJ99EJ-2693>_6<P="'XP>XZ?EMGO#[3N4F12&W?C$<^%F1UGE*W42
P])"]UQIJ#UB[:.L<W??M\C8]+E1C:0J89"!YL6VW*22(^Z4H160L5D;=OPYQ0]:B
P/EGKZNE4-D<A8)^IU*MM)6\Q/<.",RDJL\AMJ -HV1TKVRG&+^KG('(ET!OD(,5I
P&E'3TU&M5Y6.C9Q&X?=MSH7YAWA^I1A4:@P/Y19ZJFDP_N$3WIXZ7O-#A,8[6^DI
P$4KQ0P0'6.07 Z UML24']7=%_5/E7,I)UKK$'@*]'3]SK/3*"OZ\G!?!.[7QN]O
P#DS9<J43+[<_4$"QEZMYD[OD; 0>R56(S..H#].=B6+#>Y@]DSW]'+\$U;*:JM^4
P;$WZZ^QXETQR%@#>#^WRC.:&29NXHI]F.U<9/,Z%^XL<0%(H[IWBGEK@L.U!R(IC
P7W8SZ@UXYD)EH[WQ)6+#I@SQ/P$?ET#WMGB3TNG:B?O\:M)Q<;$OK6(W/$: [;?F
PYMLU6DI8RA^K<4324)H_J5WG8+<@!LW$#K;O0 60W&<M;>#>Q0VE)>G&7?R^Q^U#
PS?SJJ_83%]#'7 @QQ4N\YB&6!"E,'_\BDZA5$G>M*-9<SS- @X/M1C/2;=$\R6]C
P07BJ/K^+;MU4G_#;5_O[3ZTCN#+_9+6:A&:C@"#\M"&/=+<#4+RR,<-)":]T7 4)
P6D249MD?10$+YD?]<H\[[E(HM[(_2&OJ-E#10ZM6>)R;TXU1V%R3,!S71Z7,C C(
P4L?-22U^?Z ;/W*<SE)U$!J8*N OTSGBF:>;/D_WP\E@WWTQP-QE:&GMKD6&.][U
P'?7]F1IW?3G'ZUM,5OP1'%_-;GXGDD?IO-\CH0>PN14D G8JI%39EH93VNE-B74;
P6]SWBB#WY<_&LA>$L8G0WDKJ\OMXM(VFRA/UA'&X( YM"@6PI[NZYWUK.:HHNYFP
P#[T?;&) :($1G8.[!N/?ZZ+*?7_--#:W[*OW:Y-B1.&A@R]JQ9_*VGA,[3N6C<L(
P5_4DRY&2-?_[!KX]3="OG&HY*+W^.<-BQDO^U3.6/DD[AW?-W@T0]3/H&(=ZL-'A
P)KJ=TT+3!QPA FN%Y"@;1_]P=U@!%NGP 5L@J() G>E\U?QK/#PPH6DQSQ:PTK##
P)]_'HAU!4&"B]'B6VHP&8B))C%]^Z]UC9JBP;$2WB85/_YM@=@F@L=4VRKOAPW^D
P+$^[&ZY7><?YI>YNU#%\6?9);1%ASR@80" \<,\VI(C7!OE79N7-)NT("%8:6%]+
P 7-$56ZKJY,-E^8V-]1[Q%C9])KZ*U%9ADSR0=TTZ"0)X,_V8=4OG&#B+C[J4:Y6
PW9E>4$X-(TRP5+SN,A.ILPB)&@2".M9$@R PC 0[,"O%(]1XCG]XWXI:J:[\-:I:
P0_3K:N0^-MVUZ_=F!B/ D?](&MP,FAS-+4+K"XA8N3FQY4L^F3,3X#W#;^ZZ9\LI
P.#:@6%2E+3(<DQM+#0UFP1B1O\)L/-<]O9Z,#]^4[ZRT48WSPIA&0E;J<MFG."BD
P3 [ U!-57\64C&6TR^[W;!F.;6]='#+1:#LM\O*,."0Z"="V*U!)!,G($?7YHEEX
P1^,0$FX1+ZREWUB P)*MY)3LSMTTH"$^:$/)!?*55^F7^YJO),$P-CZ+.<Q35"XN
P5.^>M;U8_BU 3:J3&N?GXQQ=$F)6<\JB0[89]#F^CUOY]C29Q CFW[". GP)4W*;
P"GRK.)\:IY.08S4JB4"'<J<8FQ_7DQEWJI8?=<_O$*&<BWW"?CIXQ1,W5Q"&9C>C
P='[@&KXL_KPS8N#0AIFUI(J=\Z=B$\&TJ&@[83R(!R.;84@"7%3HBL\2,K>'C=V#
P3 'JLFYM@@HF!"F=CW=&U40TK-YD@>13PB@!Y$CR)K0=@4ZI[N^<9UNT3#0T@D/#
P*OF*B3/?A?Y34,XT+0Q?Y*C*E#I(6HW?8< C'G,<63",_5E2FHX :R4G';$^JLG]
P"G?3D<J1;:M#'P2+$HX#5^>=94.+\)F6S+4QI6_+]1XG,#/F7E[A93,@ZBTX6KM1
PAYSP?$!=,H9)C=Y%(#$YBP[0PA@"'.*)T1OYF! !G]7T/L!O0(,8^DJ;:;KVSP)L
PDDE@8/([;2"2MCQTRI@]J-'P=*<#C""K#J!BEULMB,[(YDR9D0]5%/WSU!I,^'K?
P+Q(OC.($!O)R?P@_0H8&_!'#[SG-O/2^,R04%#;B26;J&_OW%Y_REP:KO^C@6#%%
P,];>"#\0"KQA_)-<&*Y(5D;)0.8Z3Z,I*<TC58A<6FZ!M4<*SG8_]3V\5C)R2/VW
P-\B&E[12FT:F@R*AXQK+W>C); 8-?HJ"]IYF!B<7;*3R*M=,QW1>JRWQ9>_/>T%:
P0&C@%6'7*LW.0H$%KIIV1989%A:1:T(ANK4V,"B1-ZAQ_EL]R":KK%94G:@?^['<
PY$+[DI*%GSXH: .4NMN:"3Y9&[69! M*98PP5\E)G']2(+DJZ&-/7WUCI& N;-&S
P9318'=<?9Q*58.)*FA U0_\/YI7UTI@2;)7%?R#[^ET/(?F#Z6YQKJ8YY\_Z<]/?
P 6=O@E?RF3^_@1]&9?!)<G#9,K#@N57.ZU _"=>!"@J04AI;0QXMK;LPD*0:V9E.
PY*$;H^XRQ\?9-/^QH\&$+O(>2F378ZJ9.(;4UAMU@M<K<_5F7LWAL'U))K>]-3SM
P;IH91SHD2;O,^Z$.-?AQ&"ZH? [O:.V,!U&V6AXJH_"GB4H1SX24%/D=X]"J'3:%
P98Q[%\?>$1Q2^9EPME2[T\C)W+Z,N^(-ULN[FQ#@\_N>@:K:\$^L5:*CZF3,G+S&
PF=+]1$%B7Z<@G4;O+2N@%_>VY2C$46:Z=97! [?R<=!E _ !QH&'2'7C@H@ZZK[;
PM1LHHZ_K_I1=VR/&1;TE*:%" J: ,O=J\18F3RKY(7'\2 K&+64P^J0-;PQ,!8Z/
P2\$M'>>U@H:'[H<"ZW[YHQ4P<4@C"YY0.GG)-%F1# J-O>F?CH@DIE2(F#14RVE2
PF2/1SLSB_,9S^\F1"2L$T_"#!B^3WZ%E)C=ZG/M4AEG V>BOMN(?L[ZK0=A]2G_#
P#&G-_#?H*XE1G?LUW]M#._ZF.N)7(A@*&PA-DA9\,K&4JQ8P2:93H&9KRL%-LI!,
P)/?=O_4TDK5XHH:+.8*$U]>,]Y''[$6WNP5%M&3A;-551WJ2$PXQ=\8DE R>WL _
PST/A/IC[P*Q*/RG1WPE*53/,[2^X^1B>GI:1/3 #<Z'L'P);(14V^Y#NN,/RG7."
PC72T*6O[&%7IFCSF3Z\M>?L9))U24-1<57VNE*'!#7,%$OFIW< #L[IV)&"35J^0
PE);3<D7TH1@:1%H=II!/=V,7 =,-KS0^(INZ J1E37N)*ZB%E,Y;6-J=DM 64X2[
P.+809=CID61INMSI9&[LB]'XEJ(G41XW*8_H=&9LC19:KWE^C T=_U3!JDBR-\=N
PS8?G :WR.@MPY5S6QIF0\FQ?F[5 2D8R#9?S [ZN"+SZ@N E "1OI?+*-CT>D>8^
P[&.CCJWZT(2U^]<O*F3K,1F.C2>I\_+R%SU.I<E_@V*Y:"Z'?%H*/,3W_K9W[V:.
PD0C3D+!V_]PPFBXYY_WF=.#;D\4F@8I)<;-#^;JU"EW%N.SU=H\L1V5>(38WS,D&
P.@';\@8"N.^#30Z-_^^-=DZO<A,D=MEG.W0GP.'J(57[5\/^ZL7J\/E-T$("Q^FV
P:RE6XP;I7A98!_"^T.[I2 3[?6J=!"C1KH/N2>S$FAT.U=J.Y<1R!]-V1S'=$N;R
PI@%OD"G5B(J^ 7Y3?!6P-@,XFRB@;"SY/"](DCQY[1&?YPW7S(28U^G);C[#F>&B
P[M*2M\85^&13871T6Y!%D,=Z2#A$'"=XT2I"L6^![9,DN"*AH[Y] XK1[I?K#:7;
P*;VG;<0X@K3X#&NB;ES:.&UK C)N67[U2G=$;L[#NMJ\$Y%K==E\[;PZXQVI_'.G
PL9!R RUCJ6E_:I(F8MP$8JKKS0<@+-6I LM*LIOWTZR5S86 E"4&6J0(';O>*"E+
P*V)K.F%_:Z3%+3TX6$A0B4<:1O? S]>SE3KM!'BWQ]BH( %#^G*EV(D0LN.)GH%?
P(A" ISF<3^]E#DF\(623B&*O6?4$[GMNVG1>_3G64'WA"/LW%H=P?:>\#0'(#30+
PO]ME_]LSP63^$EY4F3&BG--3/#UJU76$X-(H<D%01X9ENK*LT[[-9:X7;J]VSG87
PJ87"W"F0LI ZE5!J>WR;4\6<_P!PH7_/T*>$"'N33G#%:F'^.BN99X/@Q1B[+<C*
P!3"$_ ; OT<C(4)A\3;V.V2]0S'CF8W6. A^[A#5F8WDZ'#)&?R2^NQQ$Z.:J;P:
P1+ZW"=%V:,ZEJQL1S8BW;=PC<?L\4^&E_B_'=/$[5QT,[&.6SI+5,O<YS:$B@*.L
PVGT[%&;J*K*/"WV\-=>'TNB>W5#>HF\/^=^:!1Y\QNGFNQ)TP>Q=)QDI F'7B8&#
PK).;-XN7D=C=YWRY[B>1;Z G[25GP+<QCVO-BJ/FU3J2=;4P:C ''8P?&><JE:]*
P.=#@;-W %9T\$N%RO?-=^@383B3ANGM$11!M5)QJZYMHGW$)N,*A(5NB3A6D="!^
P.BO&*B9X#D_>3XTU:89)\:&*64FKXSY(9;:,@=^%3>HX7.8,F)J,^1%:A5D7U<&]
P*0]P^MQ)T]NBC8J@/$Q!UZ97%/I)K3](<Z!C@G3PW^#^EQA<RCK&XXO6QMR]7!(#
PKP3"P6B0& NF#;&%'VVC'DIMNS\YP9IRQ!:##*:>P_IQYP58B6L&..5QK) RK*9J
PN'V$$]1MQQ#G1HJ28G \N/$_RC<PN%6,+1YXBVLN532&FA.=]#T]:FD0,,T+I+Q>
P@2YJP2]&YB5N^/7C5L14IK+4&K/LRJQO0EL\ZG)SZG*9NA&\<QF500X)H/4?C?H9
P]3A>:V4)4%@)H-E1BWWC8B(PY4+[&._^+QD]-^RY&US [ CU3)/-F2E\-3B/L4],
PV1T[%C3R/D36;&MO$E'6 JDZ!/X-TADSVOMN*F<DFZZ<:*/@'/_XA@/G(E.[L[ F
P!"C!\@"B?3("S(YNK)F:(O^MWBP$Z P_59CJWSA.,ZAM5A3 R)#K'W/81PL'E%T:
P<K&;6D99N =J9L7XIXP'TWY+9C3=ST]=JJ%BE&AA%ML-JNH%'1V\Z20(W![!2S8&
PE8,]*J1NS46#PC!%&Q?R.=;>X+?RF2Z>D^*0G'B)*TO=KC5A4]B^^<,I#@,X,H$\
PRU?TGJE=SL2Y=@3_@\QK-*>33C)8UFNA-;V< DTKDIA!MI1C<H.$<\VHJ,LC>Y:<
PE8M;\C+#!FF".[+^LDDYLDP 3<BCL.@HHN3@0&97>A;D-\>L+KQPM)D2N.A%.5#R
P0K!;>@0AS8M4&.&B.F!6'>DA'XV^O8OK&@0%V9%B,-3&,<>N1^,&(==80#)DLH$V
PC/*F1F+,?0?*0+;Q[%]_Q@G[CCYFI VZ<C*#QYUK/*& !I92TP^O4L *;'<F]56\
PX[*E5"Q0QP.I?#D;#PUA#&B0MN;?E9%]WSRJ@XZ4'/4#D)MGA&.WRI&+N*KE _QA
P74O*5_;W7'>">_M%G>>MD$A:\@,:^;*Z_\:E?PZ(C'QK<(9-)"(>YO(*B/X8ZS/D
P=)BM+=:Y53QCGVI@61$KM6>H_;_]D3 :][!/^9GH [MW$/?T1M?'@J/Z?*[L*/$^
PRS["O6%[MMFOT0X3Y8?ZXYNV/^<$W_C]>_?40U\P-'?O*ME57D((5="B#3O'\M$A
P#ZUKAMPR:,"?&N=;XR*Q#\GF1Z<_)NYXNN#*:A,= JLKX?*Y8,*%W\U#4(BK76.D
P-JQXQ]R,D0QKFNE#7Y>\>U&LXMG9K,MDG0SZ&.5J>X\4-O 5/)O2J%;5T#3,>XCR
P+BK[[W .E_A'>#(C;'5Y#=11RPHV=^-#4QZ/[T.F1,J>U00X,N@%@,<P^E/B!_OW
PV.5DFF0E+6,E>**:@K+(+BLR_<V(1\]_LW##(XX94NA/<+P#(<+<%"RVGJ"(X3XY
P_.=E;JXI;<1>67$KB#0IZ1I;J<(2G/XZ+P?=S/[KMBG+%X26ZEH9:E'7/UY 'CWD
P4+5N[S@>GZ\]:Y@(8!:Y$CF]0R#?7'SN,DSQ50;L\-OKZC4CKVS(+R (O11D[KV+
P=!XC/"RT2\SE9!EA<-DC4RJZ^J&/3=.SI:YIC_',L"&<0HM-&F5;7C1I.$^?E)GJ
P/?:40YX7:%X.&[5L5('X5MN41<7=FC5:& 4^F)C;*,RDE6)U;X<YVCYSQM42A5"3
PU:Z0SG;8,JZ=)KF6:BX5P%\Y:EN_:5X*61Z%O@R\:S5K'!]8![>+2?MJ:["^;]%9
PKWA?*Q_)V;:)V):R5"S*=2R8!OWN''>%K4*&Z?,=B"A.R./3]JK(J8>R\G@;1U38
P?CA>$4IZZB.NU"E&);=)1+!:("4\)H]TP)U^0"XS#9/+J!HY]F.?1+44W@*GT81A
PS)T_2=@KX41S^Z5N1>Y"G2$R\ QAI->MR-U R5O),\F$)%VCP&Y_#Y5T'9 ^H:'S
P2',!JZ1<%6?M9%<G$-CWM97KW.3E!%Q$=/L[<IH] '@0NHM;8\_T:G))_D1VS^UJ
PB-2$G2;(ZFNX.$;,O^VWS=$P9O6=0-74%$TD')J<VJ\TJ2)<#FP%MRM)'"AO?QZ0
P[DT9X&A\AP'F$BA@).O9=)5*E6+S73":G].XU90BF02C)3-FF<L?(TE8'$-@5HJ7
P8D_98K[6?PM9(1W-(0?$W.8/05;/>S:ET496T9NCXXQ&]Z#N=N1$#H;QIQDC3'%(
PMG8&@>1G)BV&$QSEN?$W@#H==@IU6F>WM,=#AMV!>CHH&ESY@L1M,$=M54GEWT*X
P<]KB.]=%.O9KA%96P73/>5MLU<P6CH2Q]'?[1+RUR61GE)LQ"P,X(X]HK$ ?VHNB
PNTB77V^&8='Z.]4I74E#/0J'T ;V//O^AC_U6/[S<ON'Y5D"I5;X5RC)7"P6S;,Y
P)#,7/4AJ7[#+>?:3FRKY&H\H?V;Y)ZP-\;SIT8UDAF923>_-K"#WP>0$\[VW1H#G
P67A! ?> (^@!>6]5R1WW67<6?R7X_G@UK@Z P/C)QB%9@&ZP]3+TY?T?=BI6WEYD
PNV\06CR?_YK1K\'*1X8W'4#4GS6/UT5)9<,R:4T3OR\@'-/8Z[95&*'!V!@JBP'S
P-(8K69-\#-W)HNA3)R K KLV@K"CC^?VIM01<&_LMC2>;1L[5@1)['I#%-%)-/"Z
PDN:60&5^^\M6\7Q;+2Y!;3P$3K<Q\4")JEET?KT*-9,^B(=.Y>A#CO5SYI4O+N)[
PBTD4LB?[I%[8Q9Q7?@CZ=%]WTNRKL:Z&\XG;]V(*9OD<>P)R!1;LB@SH3I8Z41%,
PJP.K8>H\9WO\0D"=#.1JY<\Q*EG@V'AAP@!^^\5D0-$^?/#']]0:%4KU2?=@2M*S
P2]S]+8EX9?%V= ]7VC%!V7+MCI:SUD)0>3EN0+!W&Q6]''8K[LR.GBN'A:;O-%;:
P)=F5SD'KT!_8_Y)FM1N%^J-K)"@Q1"(@JP&2Z-ES_*?7AT9%GP1=5M$)V4P)S")L
P87=-%DGD%7_#T7#Y(%#&6*1Y99?ZJ>5L5'6R\X7K)JW)P0FBVV.*('!XH475 $*Y
PY"TH1:V^:2E&)Z5!)QF)M'UH&%O< TD_UUT=)7=2@_"@D6Q?*8VE75;HVKT_M* B
PHJY+O0PHEC7+WN9PF\QCZ2P4I]C(,ARMK&%_W_:LT:?1(I.^_XLU^RJM*^48F;C^
P4J03A3MW<!*@3Z0M"A/)&4;<0W(&8L,2+LT.9G)X@;DU2&M9JFE,OXM].YT;K$S@
POG0R%H4Q;C0!</A>K6 2C6#K>2UKJ<.:)>)@"4-3_0FU8+>IWRIM?B'M_]F7ABM&
P&FC;T Y:HTXD1GQ3MBTF4G[176;\-9^2V.W>';DF7%^,W):=V! HD"BR[(E+2<2E
P,J_N1Z5N_OBV.MSZ)5B)9R0\1(%^ 96P^B_L5PI!*Z=H# SWY.YO#1RVOL %-."&
P,F@*M;D#U*_&I7H)==T/DW%)Q9K5W#^4V&SMZ$GF_''99(#XK"E=;.=1#304W?:#
P_7*P@NYL9E= M<B5OV8N$KT;(M&^3PJC]0_>SSAAF<C!D)OE]:H)4V ]8'"=;X/#
PU.W TMWG,F=@Y/JHICBPP#)7"/YSM^);R)\9_=[8],V3DM;(AOW0XK&3&V/=3++7
PW(];Y$(7>":_"H@_7W022ZT6=N,M_)7AU1!;UV@'+E-> MU$\/MC,B?L?FI=NBK.
P"(?JQ2'RWQ[UA$\9';GYO]0C+@H-Y4CR0G:R1!\/N3RNC9!)TVUZECJ(30MB&\-!
PJZU54K[ZWY SJ)2>3>$ #Q(?9N=KSE>:L(VX\&L!GAI[Z%K@?+DU*$$V+O8B8>NI
P&-,A0C0^A&;X@$JYG#H,^OAJ5XR])3#RGP,@TF0.86\WZIQTA3BKC*FU3(;=R6I1
P+BF8U09WAUARF(Z*I^:WW3<QN6B-(_SI4?*_;H%]VEMI+\_[=GD6%YY![,'4>.2U
PZX*8S^9@GMG*+/V/P^>AG#FLU ?@ZG\%>$SBU2;^<DO6D6#ZFL8#/;*XE!/#N\"<
PE;G- '_:P879<NOHN/W##/EBVZ.7.+5_X3JPC9UUA]92.(_'LR)*H#3_<:1LA>"J
P$RAK.S$QS H3\0&0=UM9VLI!O.&PST47-A#57+V-Y4(<I+IK7 ZW=+9MEJ]HKZ;I
P+?(Z1?!KAJ8QI<-_JX\8!D0!F2*#["T+D.%9WN!HB\$@S=OL_@"X?,)%HRD\ PB!
P(\I(.NMI*+Y'3._&*\N\,2>\*N'Y1L4@"AXN,22QAW)6Z7\[)!H Q;P@4QU_N;ON
P:GIV%KWZOQ,%]8^C=9F.^._:3.-1M+9->"=3\EKDAK3N?&7L52S1I^KO CJ"ZGCH
P:2-US'M!$CA<?/A[3#9KJ!,2*EUJ%_5\*N\M*\;M)1_2@P44@0@V#LG+E%IV')-;
P"_M[1!G?(4^WEW#/+A$H$$[+;6"O\B\N-I;-?^4:8ISI,F2-(5@XU_GK-GX+W@61
P)/,#N $\*UY5 /U67/L@>Q$<FWRGP4!)MG=+IX[:P83!GH^\NME388=FZ!;2$@YV
PAR;7_+O*C78NLM,1 H7@-HGV!G?1(JW9Y0L:5#73,(!S%'7"BQGH6%;W=KIQ[JS'
P7:1P 'E$!FL7'MFJ@F_Y@OT77O?] :"86D>'+Z)X%,J<*DS2/'RP=1OD#')6"SR/
PA%3WSN+/H/"@ !W_Y9YNS*Q70IN'"5[LW'90+ =<0?85Z7\*KD*$NM!X(GBM@$8I
P10B7>+@S(AB^-(C[0LA:2%)(T2W$]EE>'[.U$':J=-!-6F7P4"0B=BGV>'EQUT(T
PO!/F/$T@S"D(DU%"O9B?VF^?BYKN?K?<+\0Z35;>O>$S4?P\CN3W;G:O*6&)O ,Y
P\@#E%:ECJ+93X/6U*WV(%<2BM73K\/(7J]I??BJ@W#RTP/!:#$7]$ #^-QD7QS70
P&_"C!APQ#WXX>GX^\6B\2]F@83Y?&"$CVU!63B5M,3,+&[^0;++".<+0\38VI@E!
P]&+ W7G$:SR^PX"'-'+D>*67^.N@!'V9E1B=_^?M/SDKU?XY9^0?V-/486$)TF5%
P-@A?.\,_9?Y;6?Q+LO//BZ%4@P\B/\\;D0+61$ODGO@:&ZOA58>0CO^S1075VE8W
P7VK-ZV%C&#5)(-,7$-D/[B'/8%.;5)4FU=ZY/YU)#C-B<$XUM$LOS)3M+F7P"  #
PR.(C&U4Q(.">FW=;!01/ S,'9C.A>J]3K);6<#LL$7PH64YV$N?O'O-0W7GGT !3
P.'QQJC1SW&;9DD*73D#@.T3 Z_LABJWUA"DSS<TU$Q^P]_GT93!U9E"D\[^EXY_1
P15'HWG:PCGU#U2-4%BM^$+"A14/87RP2E^59E<=R@H?:T6]Q)"K=7=U;98&BI.%L
PP4X;<U47F[3H"C;ZV?MRYS6$3&^$[9ADX!']4GM#B+R(DOQ)-3DU#M0>>W3?VI2>
P495J(&&8?$XB<RZ6^7+Y(*#AYO':AG\5CLT)5M5/B.@#K:;+ERJOX= &15%Z?$\;
P<<HPMJ>%K%_5S*"'H-[V03FNXV1R49:O;Z1+]'+JOB27T>Q6ZQM]7]$ @"NW>4>C
P(TM2+RF*0< !J$^#'D172(M@'NLG\#[- _NS"MYC*GN/E#0]_S$%N.B]^?(&K.U<
PMP&QL!Y-W&IX=#)2E4+H %V%F(EQ7)Q-?>(=B)U 10TW66$=T/19*H\Q@71#:M^K
P#)?1]^[A-G-BUB#%>$'$_CN24TB)G<4>/2\><0UOV%+%> ^$%<!MH$VP*P^0ZY$*
P2(@@6K@\FXJL245DG+0VLR,5Z&U7'VA('.HJ@ZFF^BSZ_ ?O]@K.(Y5AU8A#J2+-
PS&DI#*T>[_A(<@,6)4;X7F7SJD+:$D",GL)">0)-6AHN#K.+TU&%;4T2QFDZW;*"
PSF0)9\#I./$*4*+>CS*]B34L_BT9GRBZ2+T9'^7IXI9-MG,^)*8-?X#7[S$0%P[5
P79Q<;*&!2@L<$GCAIXDF-5P"[R)4@LYK>>*BQ&EVCV",AM>:@.]\1[S:%(XM7MWL
P]X>NPJ6KFL@B1.U=]9,R\V82E@&^K'KGVO[\BCP4 KK*X.GI2P6NJ#QQB?N/D8M_
PC#A-M6+$?U]#R6OCG-T."(4P'NHJ5(MX1HZ--P2A&1UMGN&&Y62'XNUE[)P'NA8H
PDKB4K' 7Y<Q38%@C_-,*E(?E30/K"G-^CMH$R.QI-F-Y-*,(K"#X$%2A)4H58&G(
P-$.V7SB2GPEC?C2R&LFO81RCJK='3VL\0JJR6G?;G/D[D-N<V)0]J2Q5<1\:Z@5%
P'@*Z#),^"P4GH??'V=&HP\RL]6I1%S;ZCPG4W5-HWQ(S'XFGR^YAKZ4<8)R&!KD8
PXO]E2F;=.*R=,AN4>!0_V'WAK';,/Z^N!4=!3MDPA--$_@?<;\46?F[A<'YQ8Z$D
P@@3^WYXL>8940-JUTD33\>"BY?N@TER8_'I77("0-X?LNBLK+;?@I4]C%VPH0/8B
PU>F@3ZI)$($IQBS#X8P?[2O"ICPP51$W (WD?CA-78$U]XX7'??/MH7#E)1-ZP.S
P5QZ*UH1TKY0#=SFD^DNV^,B K.-80H)7S'A]84X'VLI''L(C+JSV*@1[_!HZ]K*T
P*_O!H[Z)!HJHW&&[^X*CF.?IJ6SP,<LQSKNJ&\=R_?KKU0#X<&IS@_6[R%_6W4L%
P![:#>YBM;TKV:K#WB$5H@]?9[]=XSAN<-&<I&^HLO0K[@!D\GB"]GPA;5+(49)WK
PHO451'.\J._ &)Q6<4?_$&_BC^SE]48^SJODST5XW3NFVIZ)NG;31AAJ(Q"[571P
P6? 3^QVP3B5R27L56KUU]"3WQ@#8TXFH^[8%2R&*<N?PK<[/5DI@12Z/)DA] (HT
P-%W)T<@G\>$"Z[7ON>BZC5[BTN:K0__*72!T748<"& HACNE!CH\1)&7LRP)_[]>
P'V%9]7,>>+CD-DT]&UMEZ7B@)IQ=UVY_N6+1G.VZ:14S'5"/V_@"J56(G<&;F_UR
P)N(##GY8Q\8TG:X8H,R?9J9N'\46U %QMB4WARNE_/%]/*O\& S92KT%B12C4G,'
P\L6VBM$40>Q">PPV) \G,+ML 8F)3#$N/89.6/^$[*?DBT-IGYDX5,,TG[E<LK@ 
PRCRFI2"AX@CP.8Q2M9K].JX%:]90+FZP>&/B;E@1)>64K-<I-U^2Q4YW"UDS72J\
P8O2W>)ZFI=Y)+J:5)N43:4&CP.KJ4,GV.ZX#@C:ATZD 3^.M27A>W)=9I]EM57%?
P"AMT_-MYA;3A&%"1]E6!WC]Y59.>52[OZE][6A])*6KKP M[*H8;#6;B0->6F"2H
P3[>>"F+NI"^PG5\.[G?1,"VFU/VO"AY 99H]J:*1#>,U:17+Q<+YQTW W\?:MMK2
P:"G-8]%6'O)>$C(NI Y:]C8>5B!>,BN-N:<L80DC,'*I,WE9NI=_?\19"#[E!%6J
PV?VT.J/=BZQQ?ESDMV>#7EYJF>60@B%W#X-16.']BV_I6WBE@)D0=0OVFMU?*?*N
P;!X6R%S" *ICQ"T@Q$%Q9.6B.P 680ALW/YK/2,Z(^L<$U*^HEO\F:H.;S+K%U6M
P.135I4_L(ZM61\8-]I<P R@ G[DS6 ^TZ]FI)6 *C(9W=+ N\\>U+22YN.>?1^XP
PJF5K,%"9*(!N*Z\Y:>C ?=UJR#K?C'+W!2<S'_O\WK&#1SWMW.TV)+2_24L&<>_1
PX$/M_)/8!]U-W)A#J3W4B6N^J[\#=L#H@N3ADH.\"])+SGKB2N/%G)\6F!QO&A% 
PC<?D5P<.3#[5,BK]M4:!;<@\^+DA%QP3(?1,VUPP"HL3I09/DICX$:3#M7P)HTVW
P25 CS JB=<YQ@MI!C_:_"H*J5P[1B7>PV!I$[YSBHT8PQLHC:O.34@3DE+L&)1W>
P#;YN)-48!8&VL8Q*8:ON\!_TJU3F<=+3TW$=9,.O4-X3/8PMIB'2.=8'B,)('A*L
PBRV:]N9BG7$JXC:;?LCI[<*S#':QF],K"LO$P'K@HD$[*='4L+'E=:#=LUB(K16L
P'XL@FPP_@MHLT>H<.%AC@W7QB'^D11,3IK^&TJYN+^A(2N?TV,I0+$1A\\3A]\_#
P[UKU.7#B'K(RJ!=Q@!2- QYG+) &U)NV3C/7/.%2XOF=- V8F%LO^Z=L3*FZ*"M$
P.'FU_,,!(,2D\0\:H['T"%UHX 1G("#+]Y/+@Z[RU+);1L7?U.P?H0)XERO\E.Z_
P</\$ZYBHXYB Q7+K'!<,%_0#XY4D"4[M)CD/Z.,'K>" />X[P8LE>*F'555G+9$M
PFE-G>WGJD*Y9*W[&ZTQK<W5S""1%9$&X/?"%+E>>5QU;[Q&O41D6BA?D"STR-T]K
P6U,<WD4HNH1.\S!TC#S)S6N]]VQSJ-]#P'O%2ZW3#D9GMQ.\T!MU%X<^60+D3("/
PMH*ND';2Y*NO^OQYQRCP_)+#1!L.)0K1L)\\.*GO.K!BB.2'IJ/PW_5A^3?Q38^5
PW2Y.<1[XJ#F_U:JO6'BZ[V8GOD1%#\69IPFC&_QX#*X?^^2M 256C3I%Q$P#$R(]
P<ZI\#N[A>:5W<\I$R*]S)R,'&FP\-MI]#Y:M5^M35+[>,4AA,8K',68 "DW1=.D[
P9=2)<'TUT)(]!5'$:=<O3/"+7SFYRSN0-3.A!1NQFNI/Z,FKWO4M6+O64RW[W%Q1
P0Y%,ZR9A8^Y4&,[S7@X"%C@5=O%Z?&A1^&,]H_#M[I Z'Y84]^6F^W];&N9=D1GL
PJC*5@BI><C6JPEQM,:J"($"-2HG<P%XKG#>]%5_?@YG5R5FJ:?%D\M@Z^R]K ?N-
P/ODI!^4]2":(R,T#BW8)QNVZ=:(OI,3%L\51]+.-GI+?;C;QTN;=V--^8"F'(HUJ
P)?W@QL<O&,()PP(PU$%K3K'Q!E4U2X\&_9+0O$HWU0XDD7WM?1ML48LWA!'D &H5
P%2[ZN"W#.K:*++.L9,05HJQLOH/W!F+[2D4A9BRB/4<EPK G)'T@.O26?"@D,4"M
P 2+RV I3I2W[$$1$;9A;R?4LCJG$2T\)ENMXR"!G[R_#IE&2RYJ"(1"$1H(W4I3Q
P8%EP"*:2#F*K.]X\BDL+[G!\WC!,"FUM7LYK)(KNG9LEBR4:\_#65@A8V'-%[K]-
P[@$ZF+_[O]U.3$#CF[GGK_BKK;,__W\ N\SBX3%6([I UA!$+B6]\$+NY2<8/VI?
P $XF86& L\O0#JQ)=(\6%>8UV"8)U:;:8JB>1M8+ #W"AZ]$>[E+DT@A?<5X"_1P
P)+%KY.N5N5S28-U031=,9=ZA2Y@,#_1T#Y^D3CP64X9"X5_6X9=NV+I$<O&^I(OD
PM57V\--R^PTPRWIS]Q*^ IO^RM.ARG2\L)BVT 0ZICFC:%!*'Y'H*GJYW9<7!_XJ
P6!V6A>Q5"%2\;<6DI(AK4?!)]4^Z(XT^_$&.:,JCZ0-P=QV=6;\J>#G]XF_FTY[O
PLWOJ,2L$J4BZVX)JG.&H4C&P.EQ6JSK@$BEW6((S<HM[)"["$&%UTI08=@502OVA
PF'<RZ=P!X&&9*GN ^B@D)BK>\H$F,SC/5[<3@J? GX8/@'3Y1*,HA%][@2'(D?^Z
P0071#PZTF(%2P_+!.#MP O/D<%\NEFU=>_K->RM@=%5X?J*^.Q$Q@:(=@8LMK&9F
P0UK1;IZ0\B5W^\0]:A'N[*?VDV47&%4R&1NZE?NOLG%(V26K4#VLBZ%W<-JA@R6M
P;C;%BP\L*INB7\]^GS(A$# N@G].EG#%[U)37'1EL @I5U5T5=M78S'^)8_"66!G
P! ]W:4TOA^AQQA%>V$C<O3#EPFHAR)6F*&,NE<,9$]WAIFLM1VF37U=(R3V_S9*>
P@[8ID7$O]X]#A6LHFY O&"1VC0WWY];S@W]UN/TK=>Q;#H]Q*( +7;,4"<WK0=XL
P0:P:-/D555YT83M_?/N.IT^?J?;2PZV(L;HT0I0%4EU8=\%*$-VWIJJA.VCG&X)R
P85W2#MB=$G#\ 4ZLX?-@_"NY"?0]":3 K/WUQQJ4\:"1\5#^*<!0%KO,<0<#$*@Y
P;0!P"]=AC21QW$VC8/Z8(N01^7:WIE5$.TXFQN\4=94\65@LT $D7%,Y<(JJ2VIC
P5@9:62L0T&8O9,EU%UW]Z86M:"=$H#?URJG69^!5T<;H&W8@?O4H7._1;!0)75^I
PB<%A3%RJ\6@>QSX?K,[:LNX,26_/]17G/F;D^ 0E9 /R62P3]B;6W&=>(Q$=E\,2
PDQIZ?P?1^Q!-0[?)C+JF[^42QDSS,.YN^A,-49P*K@L/VM[RZZ,>4"70X(K7";+!
PZH#DM97H+I.W\=&QJJM,FA=%8F_8U/W)[PD@.G/44!=$MI5J2AN,* 9GUL8:K346
P I(+K#F!L,\=/H\HOQ)]X>]J^GMP4?5VY85?FI\ET60!4Y!]K"'I6GU@#O'S"A03
P]5\]H ]_ ;L6^.LA'-=%&/OBT&2!OD+:57$^<X,>(Z \Z*M!\Z0N(VWHE;AM'E9F
P?$GW]9Y6Z\K;@3=C11D4GWPOMP[57S@+/#R,GZ*N_\ZM[69,M1JT;U59.H4DY5=%
POUX'M9%@;.+^$.T?%@$JN0W&_=D?VJDPE.\G7LNZ5BXQ#?T@TACO4BIZ+5K@+!> 
PRX3A0MICG_)Z1$48'H\;,:^.([:!E/_]:6"-@Z]2R(Z,LGZ7&(9=]7QRR53L1=QH
PD_GZAG[6%/0;&XYLS-29NO*,R];(>*> Z%!=WU#2QT$'J"KMI!Q-'MFL5.6&@+J:
P=.FDQ*,M:\+)"1B&DCF 0,&\.*708=A/;*IQMIV7[AA;"%,#J'3:U3P$OLG4*"H7
P(V)(FY[YME2*#F_N$F1.JZQ]8ZS*9]]_18CTPBQW-#:7 D'X_-6#]!A%C92QM%C#
P64B>*-H>BJ)FS-N-&6.IQO#%6:P77_<"\G0$IVJROT.V(U%M"")71! $,"YBUE*@
P?!CSYX]-^<*\'Q)Z_*E1Z\Z 8;R@#C,,\1LU9OTZ5I_TNP(D9%9'./HW75R!<<>:
PS> *M?'HMR* ;\S[P%4ZI.%*)'Z+--40LA4IX:U<JSB4=N"Q34XX%PQ_%H QUBWZ
P5VVJDC02WF,QD#PH[_)*&J8A!T+G4J8&; /WQSIY1]-,AM0&<WU D>FB^\T"3!_1
P9GE3CVU_V:2Y;;Z%$K\?O;E^W\D[;/T/JO-^>WO$^XJKO"PHFK "(KUJ-3;2%%2/
PZ)<+2\R-_<Y@F6F6NWXV]:N2USS^$4@*;M?(Z(VM9:N/F"<[XQ0UK+>@G\U<V@F%
PSE&XQ9GT^VD+^7&.%(KV*_0S?YE.@O?("V3,%(DTT!3"6W>'5QF^U;!!U7T"5-_4
P>'=W1\S U-$]]7,F<LG81S(TYO;7:D;YIJV'P$/J6(J+PV@81;G;;H#TTB.*,^7P
PU0##W#^BB=+^D#*/BGUWK9(83N<<I5!QT:.3^<QG2OK26ZGKDPG''9)&IKV,V^:\
PJ.^#;Q<]3Z0N;9?U4[S8&L02=2=F(B@.4Z)1T&!.W!C$M3_J6> Z4;7%E*N9-6(L
P:-)P24;@^=4T,KF8\]P$S- , *+KS$Q9B=Y>P8+LY"O4ES*VJB++!]%$/+D5);W5
P5?"G'=I8CZV3606] *\.G"Q8L8VF,VF5UGM>O!PT?C3[=(L]:H,WM$0PU0[;TIW[
PI[HRMW1:M%2)_8==% :@.7[OX9>F3A3QR?KAB>G%-&:?Y;-5@/ 7F]+JDWR$RUU\
P3\ZG[>J-&&75Q5OMI0Y0#&T885'X^DVNI. 67_Y[@]ZX*L\KW'%#7-^<:!2Q9.XO
PK2G$/P9Q$C/S&:*CU75)S'[, <')\"5^!H()FOO\B<$A*_B$D(FDN+.^8AZ^7[*2
P,"M9L)1"3B+?25U!2(= (9\1;F9%^Q447G./8;F!3'O0C=@9+&^2F #(A2[P9&L)
P68>GL.6XXAV6_VNY>8OT;<+0!3OCC0/IJ-S["<H ]$QWDIR!WD&:?;N-F*C=IFH"
PW>$8EFHI@T!@FH25M?2BHYY8"5I<K5>YB5T2_^<&D3]+G.+IKK^3$%A/<J6 \_<&
P)R"EHXAV8Z,[=!#RA).W:O.!NLA2CQ!Z/5:G;%O3W:2+?XIA431)(>Q$0]J$]_>^
P1_OI#A>K+KQ%.W1^?Z;ACI2[AZ0-5R2&KM\:*DDI_J1:^+N0\-?YA02D[K3K58#@
P$D 1!/= @_OPZ)_B1TW,3#,6M_V Z3@9RGZK%1;^Q5%8:20>++98G/7VZ^'3V$]+
PPMW.7AV9PEY@!16[7IGUVDH2B!;6DCG\V6%$:(0NZJ&8+V^J-D8 >[BLV#XSY/ J
P1<U/5&UX)JFB:HDVJ;>< MT.HRT2,HQ%R0,!B-"0\\XC$]^71X@U.T?8_/GTV%YM
PBDTKI *Z#1>%_^P^=0(6\SOQ+ ]QMJZ$S<J1@*V0A5F8%&-8C[+.Y@.IXSA\&J?<
PDV+/N@WS3: #V/1 AU']4\Z_A7O_$.'FU[J&IEI^9?2&^$F$$BTD.&!4B"4^JQE^
P_I^J$*4?M571CD+\-)K':+=#.E%H0A]CB)8E5Q4!Y.O.A%U;G1BUU-QV_I(L;G8G
P_87=3&F&+." #G@40K#=+YYI$4VV&QM#ZFFE4IK,;I%&5)J#L*JEMDEZEG%]%(\&
P@]#(EV^;IFRV7PV8JRJA8JJT3$\[:2O>^=D3G'3U;#R1QHN)@!(V]Q.E4D'_DV9I
P[C=<90YD'NPA <G Y)$O^2WJFC^:7CVH&F[5"G\QP[:N2G54T4?5%^062O.JT,V]
PSB9%TRK=C;L:#[C$V4F!<(#4U[>GEP"A.N:.WE-X/2V" X;AL9U>Q9H4ZU.JVL8*
PI295>V9G.J^6%CC!;O$W9;H=0'I;92X57M,F(_>-3N_":3=Z;R@FSF<HLO1RXMKC
P8CP4Y'1K<)8 2[#[XXY</^;+2,#?Y2QOT0$4^MO1;JT@\D=]*;2TXN]&/G)]9&XN
P5!J(L=JL<.,/=0^K9 9Z9%__X7QL);^NZLK5/\(1PJ@I\QR5>7LO5<[J%4AU#H96
P+68;Z9<7X!:>AC1O6</!TT[%H:ZK]07S?'AC;CLA>]NH>S08SV^?H" X774U7(W+
P.$*C=.:H0#*:V!=8BXXEJ4VQTWHQJ,<U5$Y<^PO*TB.(5A(SC ;J3%E**AH*#D'M
PN3@(X?&'/%4/*'V)M?!>Q@(#L8DP+D*ZEU")^18%^DF;!S4<$_[E<NMAC;MI,$\N
P1J*0GKHSQ]PH#<A%JT;!^Z!ZL\CIGJTFN')]*$[VC#P+A93AM)1K45:=N :?C8K<
P_=BY(S#C[8\L9XQA;HCZLSF4W7QIJ"#6I(Z)?,^G_D%A*:7*KH,AD._NQ.GB#7?I
PR<N5 "\$7;\'XM?)>H1?8(\&L]S?-V./O@ME/H6"XR-J622Q AA&6^J=BT"OUQ K
PCH<68(90GFI!'F_T%EYIPK;OCJBI/5]*1EWPQ87\A?BT;]L735TK:"X)",7NQS5^
PZ'T\\S[?]VP[GKCD;&CWKLQ&^7YG2M 1E1?":<.2N%Z8,.FW_"&P>):<E'G)5SY?
P1!AB86W>&^&:BE.C2M^UYP@3Q!\$[N/G.%3_P>\M35#''>*+H&*2%[S24II8Y&9G
PU1N/R[_MP33G#E0":IZI5&DA53GL/46Z^9F28YW,XNY*FW=?M6N$F*'D]O#CC3,[
P)7$03_?C)#3F#R3(JOMA^;)>$>4,8K,P_EK >3@[(T)B* __L;L(SV_(D=).6+00
PP&/J%D7280V^">I -VLV$JJ9@-8O.F#!\.4 5N$M\U"W<9A(!(&!ZE7\";[2?7\!
P_/31U62G\D'0[[.WZ^L\R4;;F(WW$XSLA7<IZ^C_?I91,[SJ-/R_"P>'W9620LS2
PT:\TD"MD["R.^N;'A.I7]8)T(%O'+-.GB=*H-1/$&1,P\+%(+V&.;<3$_]T[QA.'
P/N-B9*??RM<[L!,I/@!@W07R&N!8;72?GH1/?(2]EJB*CQ5%+LN(PNK)@5>%.\9J
P7&A9H;0;BP>>WR.*^<L-NT++?+-[J'P$:U<*E9N+O>_P4@)_KAZ '!3;-6_&P[Z:
PB!T9L)CR#';')DPS)"$7LU.4.E.%?(+H,3*4)B=!$^\*&'7!^0>! [P()^;7,,4*
P@^V*S>["*^,574G&WR4[-!P@/TNB03[34PT]%B;)Q_=;N;T+"JJB$0K//GL#9*/U
P^:T/$R(SI4[^L)EFF'0D<U?S"32T@VJ>)^EDZT%^7HCJ+6HEC/"*ZZPF*X]P,#@)
P^W90@-Q?=4&LZ!K=^$J*99>^/U@(:;!.+BL,-E8)7M<^,]QCD?NG1JI;>N(T)OE<
PCA_&N@XCT<!OS9;#X%\Z- Y;_#!+H_7][A&G:J1_*DW;%VVL<E9>[?DN*KX3OWCM
PDP5GHU-<NI0N/X1I]2&YB"_UX+<_:<JE]DESCNQ+U?RZ"] /XP'@\:3)2Y#HNOEM
P!U=R?H.*O?:P*XRS<!)X ?%._ZJR4G>"39*$2>Q46J CHP4J?@ %]5J8Y=UW+S4&
PF8Y2Y%]MR>H"LUL%U^9?8(G@NS+HFUU:H>+;;@NF!,<*7JJ9H$%KSU/=\CM?0^T.
P7E9,W!>:'IXN'-;YI7K3]H[26@W1E9Z%.@:SG1B9%M$8B)/5G1TT"X;<B/&6_Z1J
PVE0 VGO#)XJ3BB;>W#A?6SJ^Z3Y?U2".#=CS1O-TTSVF;%UY@P#1C##@ :AWP9@2
P(JR1!<3\1^3X;=B)I]EY<G-@R"YWM$PWF_CFQ9CYEJX$Q0Z![EDTJ]=4ZX53FU3#
PYMD==02<#D..J:[4-K][:?.128D^?00 AG\8PXXH2Y!['HN+A>F%'./4\2!SS%DT
PIEJUA#)1;E?6-9'_*MXTC<WDKJ[;VLUC($/ V ?$454'$(@03=/AOK\4 J*9OMPJ
P:EJU!*)XB6P?&1?E['8B<1DF4I0YJK]YAU]=1 :>?S,J++!!.;CV"]-"E;UU$)5T
PLM-!6=293!R!UT\,I'3%WEXRAB?^XCR<2R(B:4&_U>#XYW<Y3#X$B\$*YC+]J-\$
PN;$T4\B(&&9!WTU&ZVV0<;V<D76)JSEDW?W5YL%' U0 4*5F;<CE]/+H9O)9O/L.
P3C3>U:=COI%>/;AAOC0>=74=$^-4A"%O^\5#NDPNO[50,F#6Z.V3%M6X+ L2$ N*
PW'![L866VG$QTI]3NE0<_H8XK] LKI /A),7_Y&1_GC/ V2!#O$% ?.@%J'EYIP@
PDD#P_K!4\WT!EMN<'249=/M\^QU!D($73?IS0N;EYY3J_)9(MD<H@3^@0)#WB/0/
P7S<4]@G#?W-D[]0+X1F$L:U$Y-ES0 < LEC6/7:/6PI?8D0G^XM(,95E\\W7TF(5
P:DANR'Q+]DN82Z<5EN<#+OUQ$:H:HIT?(.'%1$QE F>L=]N$7-<B^])#Q67?M2RU
P/'RM-HJQIN;_0<K6N^D_%6>8*,\.@]J/UBDGO[E:T^NPB]=YI4DU@;98>AG.X!8&
P09S2.+!T<6[P'L>4QJ_/2$;Z]I3.41MNE&;$(L(2&3VLR,,0YWLU-8(':$4;DU?G
PLS :?1B1)H7<'US.&5V9^U#4S*6*0<";Y9N2_FOBPW2FP>9>2,E<-6PV.L;+'X^!
P=7'4 IMQ2H!/U(U.I $>;Q,$5AE$+VQ<IZ>&#_AYIXSUV9!:4I%0$/_)!P' LS*P
P.?*"AF6+Y'K,HQC:,=4@\]%:P3WG((6O*,CLAJ7"C%-PE.V\7LQ/K,D2N!-80K]?
P-T@F2BL8"6VW2-E :KS#O<P^F+(YNALZ#)5VDK&W, G+B0FO_E;_>HZ_K?H+ 9!'
P(M]T28V*-"%GQZ&AF\;>W:3"A?\^46"O-JUC XV5=Y W)U:IM2\<9<$#D"<>71&8
P#%O8_-'#QO+(Y5&9;(U'V@P"LI:K5,_L/H@$(8E8*6@8Y/.M*G;0?G.6<!N?L&K 
PN7/7 9%>;:("*N[RZ9&'GY"$$%L1Q'FJWY$=X?CWI29OM"7+KD%49R-H.HXBXE53
P%;=EGK(5 =\KK.AL'VX]#\,97[M-RHG1#E!!0-XX;:LW#O;X0+5O1\#IS :RC!"-
PH>_$*8&V'CY1O4\<5YL.4,=*<0O[3,[GI'K3A%UX\G>YW?A]Y7B*$AGX/-&2K_0H
PJS-HLWNVBHG$C>06Q'6^]OK=OV8+BL$N?-*I5NI2VZ$WDA/DR8#YH8L#CN;]G+2T
PLBHO=?N*)!E6/ *>^F/L86)9&Y*+=(SB#3<<.9^=+84!!_!U!BRJ*$HLV-WW[*0Y
POY#2'"$/YGI;"'KEJ."$"C\:_-W'-&+VO]&-?#AHW(;&8/S-3^LW?:$^@]S!Y.9@
P"]U%CK^??/*V&M3*+7US)]7]M?6( _N\K+-9WO8?(< *ZAC+)GM_4KM/@<8FQ/TA
P&0_LP6;7;--DBSGGFJU,U,,\8BN/ %V&-#BQ4&JLX:'5W$5=Q+)^6\M?WF%+1OJD
P=0I'R^9/%RG4;5U]7:T.7^(YJ<Q>1)4<[F1_D?Q2@=64L3J-^*HT3U_ <;0LLJ3*
P,SIV/=3"2V7K[CXMXQ\Z&Q1=2I+S 7MW,_(Y2=*R&D#[KZI=(@\;OB*]!SYX<KJW
PE4A.&)GQD[5&Y86=3\[GU790K"_^:J/$<C%T;]&%45,NJ0UJ7G,OE].+<3%<Y3;=
P]1GT_=C/7$%/$.[N 3[[_D.(6R3@9@Y%O)0<*J_^L W7]?B+#+-=NTFM.MZ///&^
P-AEWW!:)J\X#'B \_O=IC19/RPBKB+:OT_R"C--D\.(6BM!((OK1IVBKA =@V:8/
PI1HU^23)TO?7(LKHLXH]X;#@Q3$]B#3[[FN]N:QK[*D\OF8ICW_=KWTB:3)F2!G2
PVG9-NB88<7S"V@=_4Q$&)8 9Q :M"/EA-!,+!S8.',)B-E3$&.!!R$7#J1M RY"1
PT$4W!N $]LQ_KH:C6R:JG#-TL6)906JJ9$_Z4.88M/7T@36\?SZ@_</'$SFN@?[Z
PK=]-/_"G]"@1RG M=_5\M;NN??5\]ZG_8C;LIOCTNLQQ^F4:9,@8(LRTU^-#J59%
POQ20 6/4?5$Z%>M0N3B0L:H$"3K%J-?21>GF\3QPQ/\)BN-["V=G[O^">Q=V)2TK
PP/Y R<1BM#_\@L#>@?-@\?*1Q2X.N3CZ=>HY(,%6H</J_./X<)D<B6O+A@UU9?UH
P2'2:_5G^]"-!>+/N@UW@F(FH&L6MB-E9L">1!6Z+'#J2CN%I:#: V S]2#=Q?$-C
P3VLXY6X54G*G&>EK*; '[.W8D>_=3!<Z6A[5B8KB'_'HQ4H7?Y/M/#+SLCBK]M+V
P.- Z*+$=/?FK(G(-P16K'W ZGA^:RJU2;UY36I3N4>F]">7HPF7(2*F!7VD# 8#.
P#D$HP(\WF&2[3@I@NO@0.O*0RM85A6(H J"D3JU^EP8F@:/S)ES1C5JFE0.H8WO[
P& :3C!A'"AT:E_2O@$Q:3A#MSY*8RDW- 8<M\7GF5E'2;FHFR"8"YEQQ8>TYIO>K
PK/UJ_6R@*M;Y>2&\/_.P TU2-'&&U3)RD9J&#)HZ:G+"TJ5)1E[X+UTF4$IO-4',
PSWG7<&I;QAB&JPE0#4O-X!RA)L.V ?^Y"BF$3;QUNI[S6[<]C_2?CH>G:9M_5<VG
PQ^F$NNA5=RY_48?HM#R>V4&8T_^W%*. 3@*LB=KVN]&W<YSV,FW-$KSP9,Z]#_?6
PJ(TH;Q/ZX7/\H.=/*U*D3F%W?\%R!?FP+,GL).+(1.R*,'+IM*GAUOC&WE(.&2SE
PQ!EZ,*15VC=A*8?-ZK&_] ,5!\*I'YX]P*(FW>!/X13#2 #H?0;2@W9;4O74V*_1
PS&I U_UA,#JT<-XAK[MF("$NLP38*S3>ND*R)9UY\W.L ;GSJ 72"1N_E4/Y*,3(
PI,*-,QW<6WCYO'/A B=Y=D]FN"N  IZCYI]*^^&4!O 9.-Z1^\#4A=RUBM&6%'VB
PP2;2AM7X%U?Z \MC4LY;O+G0/[+#]P'4W9HB?_W)SA$N8 WB>PY2R=&=NP1)BX'J
PS$ONLW"&$-43PZ'ZW7&BCG=0&3]"\<TA5NQ.=C; 1W[+O(M5>/OX5#3<815^"IP0
P^CC<+V)HG ;5ZLZ)LIA2BX6-.XN*27H"V3@A#H7OR($F69#N\<92;0[@S<S-B4%T
PWMYU7/->92/#BNFP*?96@(#[ [Q.RVD@(ACUH0H]X4#GOY?AL1U^B*^1^BA!/'$\
P _7DRX,@BH]6H1N"7;9)6N47\%J1TZ@T)\ V%8FN"I4Y"_.9' _+V8ZTLEQ&;FS+
PU^N^595;LFZ&277XX;^V6GK)>5](I>+ARHS 8"JBE-]U:^X1&[HZ]5#!L0RPFM*&
PDWN=(="..2H)A&63G<0NT@5-?!=PFGGEOP*Q@*E#;C]E58RL6&HG0*#]EV)"R!\=
P2HOM]!SA*# A J"<'4X(W_-56[^R&R)G,>*:5PKBAQSC+T*AW(T9(73 %/&NJ\I-
PCQ[?"<'O;RQU9H[9E&D":)5GGB?_IT=P[N- 5/1&:7DZMH<@MVQ'"=H"Y_A; $A>
P;X%8Z4+X/GV_!^TJIW$ Q?!1J-#_>,T-RQ(U\Y(#E?O,=MCWGG5C"]F/XIJ9!P"^
P=+,<J=05D[1]HC7[+I42D(1.@+D2[#)LB\O>,O/\MMUD&X<D.BLRLQ37-\CO>5R2
P?G,Q&#;-JG"G0C1P8;T5#^EN__Q#V0W9?=Y6ZJ<@W667D#F]N^[' TSW7SCD1=,U
PZ_FQ1LAE\-8G\:6JRK R+5>)!/0@CA!O5J#2GUB"!8'#J/;M_7GI+5PZ%'(]WQEC
P+_(TEC#O+PAS"5D5NF<V_C0RUV!JF]QYF'L 8I,9@^E5@SS[* QVTJ.6G-K@\O.%
P'RG6?7M:;X>UA8/M^8X:YWPUPA0'VP+L(FXX8%PX<:OZ )A+%"A1C#@189DOMBD,
PD6]%BN"Y_$PQ)+3SOAD2ZQQMH7!G0&43N#!L=39&H.[.9W"36G=F?/Z%'7=%\&>+
PUVFU![^M01J=$>B6;_0BK#R*J]R3*&(0Y$C<(FB:=D24TP>0[B8V6KZ><MV#IX/?
P3^GE6UQN&?,ZD]"A,//=U1N,T^Y?T_EGBW]3\%3GT+CZFU,"\;X@&U>&C3%\O$L^
P$0MW&D-DTBF!'FW@!B R__Q(]=.CG%G1N@+.)*IPZ?1C&9V'X1MI$"T=T-HX2PJ/
P6Z["T:0/--MQ\2A"5YPJR@.AXW['3>^B!=?2B,_R"C=&.,1YLZ&M]:)&$-?W"#IY
P(G(6)$J,PEW.],^,S+MS!Q.3U"\[ZZJEIH+P3R_N]7#QA/?M06U@OM,]%>F="N;?
PZ>(L3\L;@MVQZ")3E6%'I!"*?G7"6:(#01L!AW]2Z7:6.MFH#S.HD[" 3X\9_9WX
P%MPH_!,4@[(JN$Q\Y"27&"94LT)8.'"0%A>@J;Z9-19@@)M]5^[[5^ZO3)QR)'^8
P'+XJZBVB_ '.CJL<[Z'ZQR3J0>J2";-*?J^#U[*(2U;,UB@AL\&7N"746!_*=05X
P^ UN64I4<2G/J/"\X.'8O\Y8 =O]PX+!YG4ASF^7_K-U;;;EK .MKGF.?7"P]'R5
P\%=ICYG[84M=/I:%8C%UFX&K#*MT7=M3YMF'$.9M39VY7M4QME"D]6,5'ZNK?S;D
P6849DU2S?AF]D%C,9 CFT2G4'A<*V5*-9C8LO9R9VY,L3\"*(OT3>%:'_IX %2"*
P),B%]WM^9*X=6"!+TYT>>8QM1,3\,61 +[[)GUV=)S3-IW7)+I8>_#(NH!%[.V+ 
PT+\\PZ,X!'.:=K3F9^>>CV$;&ZWH5/7UZ%HPV^RL82E&WJ &1@^N'SU%N[+H(!<E
PF\(IE4RYZ:<__/4=GX$<?5 7TU#GY$38?]+&OM([&KU[!(//7?+HYG*UIPW4;(R\
P9OT?19K W*\:."!?":VK/9]]_05($$Y!()[$])!OG=_F1'QR7"F_AZDM";<R&^-<
PMYY_X$R#Y7/M#*FIC&_8FS'3L2B?#[].>.)!]8P1Y-9V3_JFK! DBT^"\0^M>YFB
PGPUPY1&C8\LCSA^L%ZR^5N>3[#8]\$=6U%\)3CCE_PL\$^'G4V#)]DO:/J5;ZHCE
PZ(("PUWSMP/EYS"C^5YMI*[CYP[J@I+T;&&NOQ)NU;B-<Q1I383%!<VU:.$U4++0
P@^G[T .C\W>V!K+4 +$2;"LR",^M'>P$-[W>HA(!?+UF*0R4H<GEC-<1'*U4/J-Z
P#S5X-!J]GL+4?-KMHFJY.7+NQED+ JD!/GJF[+?_P@<V&]1:+-WRS8,D^JW1BE@-
P&:AYW3TF!4ZRWE[:CX=A- H T1MQT\<YEF1V[5+;GEJ.1R*29K*4O^8@X'PT MJK
PO\B_*J[A0K/HY;/<!L*P19.^W3X3+?HE0Z_E*S(I:L0>^F_: 402"3#!9["7P@^2
P1Q S=R;[&H8<0&*)>/A)%+6R)J2+96<1;#4M(J%_B8\QKI#S%$?;,)$-?-A)"MY!
P+2GE 8 *;>)8>/YNNXFS]);GZZ6%HG^KH'5FF8X-/%FWKD_L/%\@[-?X)S.:GLZ>
PW/YL;3G(^#3_P0&I[WDJZP&&EP7]PAX;/4".JAV!A7>.MFZ:P#[5:@UJ%ACTPL^Y
P)H/@V$\7K:3U:I&&A15+#!@.1&?>,%%-]O2,D1SB>8G.OMV"?JC%"'')G]Y7<8B_
P'I!/3R8;@7?C(/P05>*,1%=5I:XVDF;G!DUBQ5$A8]Z)II/*( B6*H,Y<&=A</6>
P:=W#C^#.:[;\)&P>5F3B9'AU5%Y#EU)N@^N 9 ?MB'5OQ^]>)F/C]:=\^7NQ;"N^
P/VH'E7R-.A<EQ1T)>C6(9@X=$.KYE[GSE]Y.?=R[&($130/'M7 G2J^W!*-)EE%0
PW4&&VL,VW/FTX*ZN9I<,ZFN%-742X>IN$[&L'+K,4DF@-R-.[F S*G ]JN?WV.+#
P#$-:7)CT<('Q.0-/+[:8(SGT7S"#RH;_6:_^&' LH,2M.;NT8Z*O&DN#";CY\M\2
P/3=3MQN?60HI'^$PS?6.'/>15 -W!K!<3C57+,VIE@V61L,TUJ6:4<4]46D5]'$^
P4D=V_L%-4)W3QC3M(P&]P>C&!C;^-0RC@+3X6LBYEW^+R D>].3 L_$C7LFN-()B
PGQG+U0P!E01'[.EBOE&X0C@J!>S.O(B4U&R$]C/@H->5VMY?$$:37LN>!PZ ZN(8
P?5QKY?X7J*PKZ1_JD'BB R,YJ[W:[J<B7DX'.ZMCEF\MS"HXC/!SE#5I7+[IGG1"
PG5T+\5&L[9PGMY(%;(;'R2A'7^'G(O V'@1GM'_ ^,1$9(?<9CQW65NK,]\ /N[-
PJ&'RA6V']II)VY&,+*YLS!RE]$1F(&%8^QFZ4)O\G3&>8)YN"_IC"W3_8&UCN,+7
P;\;ZW).^$=O1.]Z.Y][30'S/YU<ZU'F>+]XZ&8[.';PYPC$>3RA$@*-B_2I7G0[D
P_<9Z\?8QH:J6',(O,U*67*6!Q?,Z04QKW)^;.*9\PK)[_F.B7[GV@ HY<F9Y73?]
PM*OH$%E'0BS1(T.UI], 2GV\V%V,#>'*(5#X%A*<$J+<Z6CWE7C3',(LE%,4DA*R
P49W'X/$V(D47@6>#R+Z1/6#>FFRCTQXKP%E[$?N#BR(0P_Q$Z/AK ;W3I:_$LWYD
P<)(;&ZGK<T0@)&9Q(.CD@>/O\TQ5N?4L>]Z"711^-_9ORY$X[S0#]*/DW8.6J=N>
PF0CNK/:U7CI'.?K&,X5E$]X].V'&BV%$TW)X-U("'\H7@P([:/TAWY8MJ'5B_HG'
P'IL( ">>-E]DD@5K$/U#ER#/.<O!F,8I*W*55EWN(TW9XK$*UB"\M<0\JD,_X;U*
P1O97J$!25'M[%>X')6$ BKIAD++8<NH6FE(G[Q<A4BXV:UHFY;#T-LR+3\W$(Y+@
PV-:$OEB&Y?K/&N][;'WMLAW0C$-YK;0OKVQG%$V-->YR8-!+$A==6;(O%^MF9"JW
PLY'4:^<^N4)N\BZ]^/?E;=<Y@MQ*J/Z"#X JQLG/8XRSI15A?:'/6?%(\<H<05.@
P'EZ_68AT_O:-0E\V%BAG4'WL*F1;F2/!.!1641%:! ]<:[RLHL,;@OCH.:5,7\KP
PS(9%\# T.=# .:?MC<A8O<@E,+2\=+WB;D+Z<<:UT?DF-]]?O$;9U"@]E"AQCR.<
PC?529/N#V^JB6.;*2#GX8MSS677SQ/_;"8R$!KM)$Q4Y$.:<],H&M3OW#'4,71X.
P*@Z(F,2P]F+[3V),L821X:Q!%:"I(#B@</Z0^3=RMQY-DZS^#@<_Q^MC0\&02:+V
P)>F)&\,YI?0>U21!@9%J7&\UOZN3XNEUE*S?[U39=\>.G(&=<$&(SDH-R0/@6M]'
P*5_S@C7#5+$GN'KC7N(FAH_XXXA?TM,JGAG]SSJ"+$*SN6TT(7XCI/CZVH(6 :K5
PP)^2YHVJ/7)G"P</C>VBIFZKRI8U+4#00%8OU\OS^.46=M2>$D&0N]R<!CZK!?V#
P+RVBGS\:ST__   M45WM,J2(UIJ-%#N'FNU\#+!<^VXNM$4N3J9<,PA\0SFJAE=T
P=K\T7S1/V1I&!(5=D%']HDX8<>2&W9'Q9K1AX(.G<[=2$A79Q^5E5ZQZ^\,!'-V&
P@0->@TS#L[S3K=UD'@1@:4N%S;CDL3UF70<]*O6_'7_?)_W1M+BAB0G0C5'4;:M6
PDXAS;(LIOOCF*K*>D\9V@0<1#MO?Z/K)KR(]#,0W DZ R)G*XOZ Q"+V@8TBO*WH
P&08"><36U'?A.O6BE\QV7WJA&1 >=9:*4MUW+X76\@GMN=^'*#S0=$-$\,"8UG\E
PTT=,Y(=HDR=A4U=V[HOS1FQ:K2_U\_>]WWVSS_(!J >%9$^E&H18$Q9-'\0AKA8(
P.B6M,@MBV/VOK$3,L0) XQ\2"[9)'OD#N"6#4$T8L8)\FK[- 3X H&^"UG_;M&PZ
P0N;A,,537.MR?^0H-GL:.1& Z"D)G @%E@4S6MIJ^8=Q+>E-[*O#R\U0F[ QCF'N
P8[%4' TFEE"E"NR+N]X<':-*+"JAZFD*VBZF/EY"->=,Q)$5W3(/U6B [&*"8/L)
PW#N]]@SFLQ-KCO!J<,B&E@160O%B+LV1&$7IY7N8HW]HT377+72\CYA2 ;>SC&OP
PSF]P@,9SJH](5.GJ3K;R0XJJ8KRH^^U=:0O?0_+X1EB'\';]1WAAX#[5T>!L=* D
P9RJ+>#%96J<0.EY-E@?_F[^2FGD[_TDKLU%3_B:1NN#.UDUE5Y[#]ZXR*\/&2/^=
P5!O(A&69%\O*W6;)P>["GI[>KL><[Z,+\M*A6 _UR =O-^_&,KX <$4!*!1A '&>
P!QY2XK^WL..6F;.6;X-"D+=:@'1^ 8PEA3?MT/V!-0UVRSP>6TY*B83;\@+?*IG0
P4U$1501P?]'5-A;[L8!<K>AX/OCN31Z[ LLBY,(J:^*\*(B74ZH3XQ77%KC4>*X+
P-9SV<!H-.!RE"+X1NL]9[)YA4 %"+-]5W34)8 N\<:4<7P07JG9?GF\@(&ZFN6B5
P/#5^98'M4/&63)=55='C#% :N #A^M^UQRS_.RO6';!T19%_;\8%?62*6T@U(R1 
PV2;;RD&WJ(]"RT '%>R #V(>#=>) F.HC!3S[4^O2Y,P?D\[B(./W=OC/Q$-\/V*
P$U\/_(.8CA\G0P22RW+05P)KQZN+.@$0VP!A,KF0Q3RUR3ET$9>L;]X]>2O.F=T-
P>6])4:N94L[^XIGR1B3>^TQU=1UMN8,5[-, +'^J,B^^'1'BH1##!2X\L'96=(_A
P(B:F0"DJQGQN3C@BTD\EH/-K?NEGNDB8Q6;AG0AD" /(.18K47I#FO.MWW8@YWNP
P+GA'XXM;X=\P09P&L#'6.E"9++&FOO58< GM>>N\:Z(I^^+*)*HOPS&2+NI&H8<!
P+ZE<N7X3I]VU0S86^=%4X3C_V"UE  ^Q2E-I^WY16(-@&SY$)+[2G,!:K*DSL"72
P!P=1D.:1*.J_6*;SS-J@.(3PZ?HK]F/_WN 73D?"DRMR.(,F1:SP!_BBHYLV_$J[
PI[KZ_/[BTO74ZGV8=3S><U<M<@.=LXN K/K)11F99(JXPB0\Q9&Q?7L"=TI)X#J'
PR([[)MF>!1M<OI*/9Z+S 8&-?&O$]'C#_B\WQ(C$-2@CT[V5GA_+80I6G>+?^"]F
PRHN4#X^+2+M9Z-W4GFMZF^:[H:4-@+T1E^L,Z*F\MZ6E.V2[M#3L 9^@Q#'@3\TJ
PKZ":6X\7PE50PL\7GN'O-!/_E0 +6X1]&E]L(SQ)KQHV%5M/_39( >UJ =9I"/5R
P)P%EQZ>M/.<$$OSDGW8P888C4XQ%$XD]J3^KNAUF$]2% R4W<0[]"?'SW*IPCXIY
P1FRLL9*">&4?&];\0'&W$A+9GP/GIRD*YV0'62'E1&L+W=NZ;-A&;4;'=:)$+&'Y
P7L_5N^9>C[Y7M$"+<4&,( 443(A5QEUR,'62"T97>#I\5+P>_ [DQ(-.^0NI_,OS
P(#=..<^;PG@]LWI4HSJ7%:R>!_L/HI83$2-T#L#H_'!B9Z1"1(/\B)MS,B.V,>E8
P=H(*.HG+4F/VZ5"$.*.=#@04L])66'6XG-66_=^N=D+ +X]0\=50G@/=I:<!Y6L(
P$*###)*#H(87ZHM"-TI6MW]S4-+J&2C:JY7NQ>)I'J)DAD_H?EO9ISNK<GZO^RM$
PM*L [S>DN)=J)B8Z.=2^43RCM<8QIS6&TIE?>-^MJ64N[+KJGQ(9UV>%WAS7*T;1
P_VM'!;9<4]>*8:MQCK(*+$)(N_@'Z[Y8C0D=F;J]E,ZG3WJR#JV+<H^N!W_2C+F1
PTX:3M16R&M*SA.'RYCJ3W4XI*8VM0GN0]>E1]<\/($?<A"82738(\R>O9*W)]A\,
PEV4]:D).$X<A(,B3F!.X?2C.S+MKQ[B%*"<C5YD/4L_;R>]F8O1488-I+B3?G, 6
P8T^O1LWO4ZJ\-[#0Q<#:K0\+IC'3FB>(@"U;^V06SC]Y'X( 5,6&/;3L^6SFR>[$
PFKPE?2>^NFPK52?II2R3-F>9RIK^+M=FIP.#E&<_=5.5QT)3*RC1'5^)ZEV:<U+T
P2;_X,96N0EV:8W5;,K 3LS$H8,29&]B=%L8=[YP(O%KTODJG1(POHU. ="F_=?!F
P!:FH:'H-][DM38LU%90 <%"I11SLO\)F2EV$YT 1(P10PA? E(.(K0:F+5==>NY9
P?.*)L5\S#@9X\H0B!@B>0"7),,PJ0O<A.E:=J'#]#>&N/&FC0G'@ U%!V)*=-1M2
PSX"%Y!,QUL5> O! XNCAW)N^\H[7B8-EUA*17BV?4TN<O33']57#G%">\T0UUB%X
PRJ2[#72N<=TO?S;6;"FYXVIC/!?!5=6X/JX^]*0(  Z[47P#?FXE=APY:PA]$,@0
PJ9/PRV5/OTB\/*5.;Z[(YOE[;N\[[8QQ$4)T KMXVHE+O*)T_*02A&E4*N1H*AZ9
PS$R'<;>DFU7_M$)M\<8(*ITF#IPDRL1!?[>\GP8C L,%7#X)9<]T0LTO<B"47LN 
P;<O4^:@Q'$^ #?4&CE6-K@$]J F#1"LS:-GK/,M*8F\).8%&SM&F?)IYBQ^C/]NE
P-POTCONNX*("T+)!N>W-AFMO$4)'/Y<CE+:J+79T(OI&GO.X<J6Q4#A4F!H0RYL(
P"B4_R9_+((N\TEWJ^&$;V)<KE5#]; NDMX,GWX[YL6%K W8J4QZ&#CLRNUXVHRES
PA6ZO)K)6RB;-1SSWH8W=P*>)JC8T%4"/11_-Q&6$^I!A7AXJ7SF3)+IL'!5-C'=?
PH"@<A].'NZ.V4&3TU-Z9KM.FF$.5WM_KUB"Q;*]+\E\J1$2UJ0U)OE:8XD4*CZ@>
PZU8>[Y1Q#!]&_=RR@L2:YH+F[.L!83MK3-OM*=A0Y#'%@+#ON+IWN2W]_0.]%?+^
P5T^,L9_5",^!_(ZX=*945:)I+NNFZ(MI TP@%^WF=0)$05_LO"H&7YAII MA2G'(
P>6T(J=:P^A(\47O/\V2#\QZ7<BWZI\R8=2SE91@4<Q+RZ G[9B_("#0 $?Q@*P0>
P00?J_-X6VV,-O)\],-(B3A/OZ@%YQQA4(CJ%J.:5Y5W*RFCG+XF*7@6KLDPUX;^K
PL(W]XG,\CS@6R.*"3:QQ>2WSU0![53!=BR6H6"GYL.2<PM1=08F].;E+)HUJUHD6
PKWO(0X8RJ#UAG95,)/M?N(SX;*8?:!84%MNS](!*#C"'<%GK[RX&P/ 2Q*&*ZA&Z
PJ 5RVT]Y]RB,L.[6?RBRTDG H,+%; 87"PO,9EZ\SC=SU7\&'"/7J22A@SBH,;[V
P%+:/,*R+L=+L<3A7D<D+1N4'HY@D[8L NU)202YQ[R7B?>IF5\N1[;1ZV;$$5=C$
PE@F+[0@1)FH0[STX2?/D42%2YF_#<E,^WER!L[P66U=?1?2CJ/C0@>?79Q,=_%^(
PD!S[/:ZJ2[/%Y#._(FGW;>JN37YZFUQF1EXFH$E"1H3K X<^0E2%;$??5!1>&C/V
P39TYR .OPKL/%".=<Q_*0PO]I>[AQ---3?[BS!?0F+];"8@-3J;)!Q:LL(O6OML>
PT6_&T^LK-9:>2I^[[TAR2NS>^<Z6QHMFW?^W(_</EXB*96>_K#;3Z]3ZU [J^4[]
P7H-&'96,R^H-$H.^N$(4OC(X_DMX6+#5!<#^1#A(XH8C1AWO6GLG.NHJ,4@_X8#,
P^7$29,>(BHD>9GV)])G-Q/Z$;?].X302SX'IC%'94I"C&WCH=^%=UI.,*X'?%TIX
PZ>3]AYF?QHPLJ\U6\V0#W?-TN[ZX[/J)SZF@>1[+<=!6<*<Y:'_V&7C]@4(XL1A\
PQ.^NNR\:MU'1()ITQ1=SGPL5D8#&N>DPL?=1P/+(%-6"Y/<YA8P.9<@+T*D%O\\X
POBRA#RF!N@'J*I9ICM9:X6.'OQ,:IUBZU8W3/(7Y"'2W0=+SZMTA$M(GIVM6F[_G
PLB S-=CJP$;A8&<]D)HA(RI5S33A>:)'?,YXAYUV;?VN+D\+?S/ ;/PP&#X&)OBU
PDIZ+E/37Z%96G"AM0Q,J]MZ0_$I=127) 9Z&-\=YE$'A^N;45IAK-@C<" F1'OZ<
PNWMX&*X@K2]9RTAL<Y/<*@#$N^7-;JL3:\^F-K1&<U& /[]#3'YLEC^54AKK"#^:
PN<"')8D[7PDS%,6C9)D>Y0T'&&:)HCZ6O6!15?(GHYI>-GX67XK?3T"-3*Q@H"J/
PL$:-&FMD\RIE45L\.@1;T;@=)4>->WI9]>9/848(UO2>+*I:D7T57BA))C/I>U"3
PNKAYW__]W<55^^4I9:C!<X/J&/T"COFY40I8;XJ%]P$?/C6'J3RA%@<LZ\_MI(?U
PQ*SA%&:= <MEKZ1[@@*HCJNPF+&XS@H[8@"[HQ"]GF)>I%3!;#T*@</5XB^7Q1%P
P(WN8BI#D&0JUN$?=!T?K>';D3IYV\_,.K'XNVW9:6!?T]9BX1SS<P$1LE2,4+Z'U
P"?RPKR4=4> Y2+K#>8E+I"!;TH=\P4TW-Q< (:0@>FH/=WF(V&JCY#!>LQ+),S(M
PX7=6D@0 .)//85D;>#5WDEM$\RP3(T:=5.LT9QYT_IS.I521;&R=&RU+HEZ77RN8
PQ\BU7B2G8V-S\4\I?1,">'-B)_&;S ZGB5X#UB%S']!*M^!^FS>+7-@?9-'FQX0X
P4?>#R]9PDR.*?)K<FC0G+9L,I/XT=/]"B,+.9"$Q"51I4/M6_^(OB@"Y0E*$;.ZS
P-Y\ZW=J):EGI7\+VN(%S6$YL1(\(5@#X/YU._!K<1C449P+QI[WKFK%[_+X6;@7S
P4 5ZIYPUB25=_M>Q*\NQS"=YZ72<>8%$Z$CA5T;J_$@(C+CF))B+B<:=Z%N'%]N_
PM_'&?IMZFOR[#,'SKFY[XBU96XC()C7UYR:TCJB?E^W/A%!1[Q'8Q,V$$UGY51GM
P050._@(A?' 6&!E@E)N,W-43R,0Q.G7[E,[;BOC7U. 2GL'<5H93<UNH03B<6]1Z
PVK8"<\H&%E"214,?BMI/O60IH@=.V^;9CF!G245Z+QGM=P?TJ$-2 @S;@4'*3<:!
PA-T>0==@.@3J/P8,$1ILJ &!==V.T0@;$[N:RN =?T^"M)+4<(U*C"TR-[ ;/CS.
PJA:(I[)1)$29"3>X?RSHOE60B7OK^N\XBH*&@3R.8."#6HV'K[-E5VO710-%%_D#
PP74NM(Y!)"S=2V/WHU>9M!%EC*!?F2)Q1?)(RIYV*,>C).7*],\HE[<&6#/W/(A>
P48BM/"AJBPR9X@AP2R>_<7"@5NZY%3G&9Y!:"YF_7HLZ2,QKYM)_T@R0BS/:.$!-
P@OGE3?D?/Z,_&ELJ#>3 ]Z7@/_FPV;ZJC%[J;*$NZ=N^*K,:E31)OBK6U.K+/!U:
PI#O=$_=P*[T]CAYI,4=J @?3K$H)QAL+]&Z*>%U%?L&UUU@C':FC6)0+F0)BZ4G%
P:?<13[EYV.;"] *\J8.V]F+70 35(;:.0MR.YYPH^ES:?F7V%SM)5DD1'CHD'+ Q
P, >%8ZA)-)=TC>VA3%F\R <8T,U:,5&>,1X"$)/(R1R!-RUNV[Y.*]T-P-ZZ(#PC
P(6A6K\?J'NQ[BY9:H2*-5FH&30M1@TSCMG(C)(8%XW>DV,ZYFA";V!N7!:4X&%'5
P3;'L&^%?S4%540']=L]26[E]V7(DWF\9AL[)WZA-4."2A>E>\UNOK2YX6?GKLESR
PEOU&IH;I80D1-_S$'5= H!"833<4X=T[@F>(*N;).UCDUC<1'.];PP8"H<1A*,AX
P&@L'UZKL/R]/(3PSU&!DNIV"MT12$A5G =O\YH:])21<V,32!]36!7-.WH-S^+:A
PVW$S.LIB.8%#]<.)E+  IT#O(V#,SHJ5)UJ.!-P!=Q&#]S1'7\P), D([5TCC X/
P)A2H]*6OW(B?'-4_9(WT&V?.S&XH+DM,FROD]E&S%?1D;J\K*7'MI:5*E] ;_VXK
P%@-F<)5E-::!';C7!"69BV2!4-$'5"WQ24"AUHE*W\/6\MT!;J47?28XO@<QS\N9
PEO"PSB+7&>HD'*.22PB=QV;#I ><:2WU]^\(L 4VPC-Z2M"]ZD IR)R20!N7U#V 
P^J -[-'6)-I,"U'L0@[&/(<01QBY&I?Z$7"K&+4]FRKD$1-0A"PVH5#I_^/F0 #A
PKI@V<'@M6X;?A",ZD'ZDKAQ-@!_,/ROOOC8\BNVS\G$^@I>N@%W=VKIF#.J;3EFD
P,O]N1,_]BB<"!H%ZM\V7KBU'9$_ZH]4;IY89E?$)0C8--MW_Y>5J9=W\M-:O3@])
PFN6K!N?!H_6+O<FOP'B$=5\NV9\C&OD5?QQ<!$IP&B;J*7R0]SW#Q6G%\0]2<O\O
PO&:"S:BM'7P=4^;DD0&_3P4IL;KH>C]LB4L/3#IX81)\/_N0,QD4@?NTB/Q%Q?+:
P8T7+C0O=7VW=MIGFKPUI$[F=L(F@+(XS>9\OHP?4>5--I3;RY2E"?%X!<F@P]_>]
P+37(51VJAT.OZ)Q:Q 9J#0<>+P>%S98A?E@ATW+^*)/C\GJ'LYJ[HIM!EX/<94?R
P)QLPJWG8_5K=A>2Y,1!2U5"/.U@<"5/UY&L"5S.Y[XF5EK!P"=IR/(1'5:!\/W"P
P T"LV>[MEW5@PN&PIZ#KR\9M[!7)7_2=3PH9PM69\"T$\PP4.*H]R%K]I1M<7QA.
P)'-GWFI%5\*O-V'!UANGLQEU0VE!#RAI>K3L4->-]FJ0$0N%B)[,9<R@VM>\]I.^
PN1:]>9]9J^E4H\!D=T+1.+Q=C6981E%RL5+M)-^9V:Z2+(\LO.*9P=H:YNU&,N7S
PS([E<ST;P"'4KP%Q0BQ\Q(U72UW,3I)YHJBLC_S QN%$BTI!/R2BK3Y;=KR7PCST
PG1GS]6Y11W^X*VI7#"Z](R69]>-Z-)(TVID:!1=]O^VAIN%<$'E?[^=-":SJG!?"
PXX"0)37FVNQP((_<-"#+8+\_^ASX9?7J2^!<OO(T=3'I'4 /85^,'#6UO]XG\JXZ
PR]FG"6QGF"\H*@,Y3?!4OFHYH +5 LA)U\:RO:H".2+.I!2DJ\K7=AY#D;"DVH_&
PWCG"?-78"!UPEF/[X*5+C]OR VG6T!ZN-X0K*O+B=OQ;0^7:\S/%IH&R!,Y10U ?
PH6J!0_^!ER0U;E/<GATI_37#$GF@\Z$71M^M6!& /0_SA*WKD"U$FVGZTL.L,]0R
P-EB'07ZB.^^VQ-'9TQW^>.FW"^6V=Z^(@-E6 Y7.>2%Z4#8ON.Q6$N-G/1X(B#<S
P4B1,4_@:^*XU'+B/?Z$81<QJO0'SM<T](34M'W-8D"7GW8?&_'T$3:JJ:#;CT.G]
P0?(9( =RW)PP=FM:BVA6=%=:/!>5AVR9XQ8\'I*7 ?G:);%%3Y=AB%_O1YVB_@@W
P[+UTE'/]E8@."VV$"0B:HP<3OJ) YH-%C'155X)X >H+$_FY(ICT.(QTINNG+F@U
PJS0O9 'D>+@A!MX[D)BFNRE8N)I=2QGT?T&0A<)EGL'&K10+3;4;VHTJ5YORG>+V
P(<\[&(PWW]<+DM:CM#77@9X3LP,2 7U5Z9SE;"2[N40;'.N\MK\)Q5LWLU=)!0C?
PK^FSVY=?UR-B9+U^ ,KL9GK9:(,7>5$)!D&EDJD=E)<UNOJOL4[27B!XF7PF\R!1
P?=XMI>;<"O4LY0<D\3]EJ$NX=(K8_<$<+0&<'<115!L']WH-P\5\"371IV=R[!U?
P%1)1-X*EH.V&23CW!2B4 %E!1N9[8!)4@!9"H:2Y\>P@(YYM[@.91FTGD_0X$/Z"
P@^J_-R>^%B'19$\8Z+E9Z_N4.4KF\-]J[58N%80?931-9F5756K8HK) G' .+,#%
P8<[ *;T0?J;W,[5OU8B[IOE/0=.EPNJ9_IW7,2_V .ZM*I(/D[^8YUCA<Q"P"0\ 
PU\V$6@/?^Q;U=9FG2%+G'VK\ 4/1J22@T+;^N@X7*V\3HO5Z'$ 8?O.8C=I^]>W+
P^7))CLD[0XE&[-JQB-O*1# !?H(ZFUDYFW_U HQ%,2_P2XC NB)/U7F7UTKGY=>Q
P;$3U$N$/HON]A.\1G<WB[>"'>7D-6_-P%&7L'Y]>\)^N/5BG'4[T91)]_V*:+:*$
PGHH_.&!>>L"0S#R6,99K8#E7M4! -$X/GGO^MIG(=S$*;S6CS_-X<@70.M4CZWU 
P6E&+Z:4GM*Z.5<\PT4>9Y];B#V@$MV0>A_/#UR2)J*4.5P+KP/!:%AY%7 E%9R1E
PLS@-5A-9XW3*J#UVY/!W:%GNP43](7 J0(.M:TM>(! (+!P,;R\7:)CL4?X),<7&
P\4-(7&V-LAH=E3/_#Q.7S$Q(DH^R^T,1T*1R"#"F*CTT+GE(4M$KP$=.,+XS]?JL
PPR*,[@.O$Y%"I&U<V:$LO(J!PXV]A@I_[EK8DA#2?-_JV _0V@OAK(_1<>$9\3#X
PY<3T:!$6+%?PGX$5DC&F/O8V+-*X?\H(^RNL W72'G(.2;)KI+P4DH==;Z$@^W1 
PH]SU6;!RDJG73B!R:A]6,E;06/8G 9F9=0EVS1GY !Y!+)(?3 GIIH4UIJYPS(ME
P7YR/1G!BT[J;:B"OO]F&%Q6)J9;W][LNGL4H<<>"OR1B+G2P9O&2K4?UR#]7KA.Q
P!>$?%F *K_HI,57@H2AZDUHO?MF'SSX85#<._3*4KY68KDTNM;\'B 3&>3(DOW N
PE!8$,9Q)S7[%7S^(,XY)=!6[?YT<"(8]6Q\+7B<K7I7PF2L671-[.H_^^6L[ R*V
P!49?*4@[H%(F-HM$6CPBUB]A,M:D"YGL3ZT),G?2A,[#W;_LN6))4,H3EEN:$*/4
P%?JC1!+'M'@0CVRT090(;=BT?YE"4A9*SXW>6T2*@X2)9?(&<CMT]L#5C3))W*;,
PA'NRYYMSO7L2&CG)MU-Y,\-E2OEE;%I>A_WU7<)III9J.RCU;1^C2%R>$QI=&X,"
PZ!HX&/!RC8![TU(W^@.Z* X6*[XH>M-V6/)C+T _M-G/WSULW+W=P0<-$"W(WUKD
P/'.)_UUT^(B:.3?TI]FQ9PC%6B6A(\+\!V.A !_;7@FUK0]'/8#0&S39IEN6]#@6
PF Y:)0$7SHS@+$:#_U C;!SQ4LC#XXQ05 BVV2:G@=5K?/<Z62]1/A^#WF+X)-I,
P8]>#K,8X%/UIPU;S,ND7BD#W54UI3B/EI^3VAA"S/H8SN[,IF8 ]YKF(P^-=:]"K
PYC$Q"X ]7&18<#T).K="? \[<F+(822L4.">["BWCP]S"!_>Z"#/!8Q1MFAI4/N*
P\3#& D?B#_WB-#E+T/OHZ#1["C/1,#TP0S]R'Z*!W\VL^0.R[\[XPB)_%5I=8P!$
P+ZG\T_+I/U"*,7TT0LT(7O1?%KIVSG+N#S_S)-,5N4+F'39_ '7=!!30C'?92]BP
PN+0%+.E?"D"7<DO8YNU0;E$4\9+Z&HI"A9.8ULV'I3/LK3:HTOGMNO4;*U7Z@LM3
PML([KX/5^(MWEC$J0.J^3C]&!?0I_R>3.9,KQG)"UG18&C=ENMNF<-1O:J(>C[&%
P=6%S+<Z0[46 "U\ZFD]ZXBRAJ1T#]UC,%0:KG.GNKF?:STMW3VJR*&-17#*BNXD:
P8"NADBB67J\4(&!9"?-6OE,X\9<]4N\HV> [[9NS;FFP41)]@Z@5E;S\_(71$=8J
P_?]S?W9&=WALM^M7P0@X(8WKJZ0;JKM@#U'B&3=QT"@T8_!XC*B;DR 6Y:EBH$PS
P^;_7XE5FBG#<\;,@ZW(4C=R8SF*OC^9B7IUDREZ%*K(M)D'6$!J'R9.@A[\=N#;A
P5Y5$(%'T J9FN 1W),F4Z">- <P5YH"L*W[Z2DD("^K2"-W#+[VHNF:02& 4>NQ&
P&#FU*%!%]^<!;.;I_5'I,X62UB6Z<+= 5VKU\?XN#F'CX"2DH=<Z99GC._<S1!^E
P>)C;CDO"DVK=^H-<F+M3+6302PCOZ\Q=VF&7,^H3&HOTVLF<@GY)V-FDO0GGC0;*
POT@S?G-ZU^6M!S&U&=./D!NSEO.:*G2P9[ :X9L/&\8@J@S(V%TY1QW.[# Q)Q51
PS%(4+LLI1*&*?K)R:,\UQ,<$$4B&&U;QD'29HA.KWP-=.KT2L?WGCL'!I+"UC)">
P^T>XP7 $<3/T[KZ,S^=3^N";5!_WKY:)E;7O&0@Z$_6KVW,IT,'K+9C"J5 R8L>S
P,=2(<=KJ80 %8]V%!V8)*^JO);%<$87N9M*FS Y(>!&-5]AD!O+7H-"QO.S 'W45
P?':BDY!N"*^D9&4;SWEW('(3-T+S-F350&#2+MGB1)DE+5=]BPD[E&Q=\$+FK(Q%
PIB49<;EZY#<F$DS"2SQ[6-QED-?'#S]N!P,([/GA&1">):$D?2QN!O/5$8YV6I3F
P]/+MJ<YUFVH-6_M-<"P+4 "\7#*_/@>$)+GP.IYN88Y]*4#*!H@()B?W.S]7]')8
P6+<H'SIW5+Q7TC<I]S#PJV9>/C\!2<1NZ9CJ+^8^3]2OM0+37_82^>"?FOYX%+[*
P\5P*V<3=:P(#E0'+L"<+UW$84-/:SU&VLCJEMSM<#7 'E!FF[X+?90=70A"M]9UH
PQ(5&$.+2WV4F57SG)$25BBY*?!PBF295J9I[K_^^M[0'@H=K <@2GGXM35I3Q97I
PD7_!_DZ!59<?C]Y:&M'N^E^D"8)X^I=NV._TCSOQRU'/GK0F#*D2DD3F>PW>@=![
PYRDY@L1K&Y=OO[D6P97+9*,0-"M'%WF6Z5DSU57:^*U*+.).FXJ1JADOLB@(?P1_
P6P.?7H+]]R)I0R=HQHP<4(0C*NV;[_L?F6@89[K8ZJR=,:;+H!Z>P+N(;1W1F#^3
P+CZ;X=6%__N ?T&EBD/C._?KRZ[93@ME\#]4BEF:$'PW;3<JU5O45_:Z)MVY# =X
PM5PTM*HK*K:\@* Z/32CD_]D;=G04DQ!W[.(*A7@9*>D*./JH:\0'_?U!%#LHMGP
P7GG2%5B(G%-I$4Z_:ZJ'>YIC)[.UORF)W"9;2 0T:4]H0WZ&%WDA:-PJ?F$HQ_:C
P$ P)'K"!QM1G@P^CU2RE:F]R^_P25CC/F.07;4\O)D9?Y/Y"=E4\]#T:( K$_(4<
PH>)'T-=0!."[,5SMJW*1VO YZ_4'IZ%I]$J=LYV"U"G]<EKRA46_\"XU9FWT]/CU
PJ *M=:&M[G)^R+\<"O*&QSX@Z@>N1@LI?2)O\J;$E2YH8:0Z;\0JQ/GE0>(K6((K
P#T5XF%STNL#4'RTY6FAWWV-<"T*N>R5/,OQ11,"8L8;E8=^8XGAFSBVK[8";$9F$
P%F(<&4<%.EB^*Y%E8W&-4U?:S"X,&K3+<R;,LW$J S!;I63(:W.RS'&"<>'0S\_'
P6&B^QK)/5O'&JIX_5Q1)3<63LVN#V\<;7(!CCQH_:4G+W2E#8^C=@"U%R9\;)?Y\
P;[E%+D?6AV'Y?V%+0M<K!F#R[WYK-(AJ$;HELL,0_7W(8$<X.ER_<"L#0Z=QM85S
P_Z*96$"(ZOO[\">3*&%V+D7<O[64\RY=BD@\8$:7<YP#8DMQU$M*^.)P#%XZB'>@
P;4RJAY3%I)J'&IF.5,%]<ONPFRT>^IW43B.TN1L^_V#FF^=0#!6T40$Z"D;%P\1B
PZ,_1!#TW,%L 2H&7DO  ,2/*97[<!I(J4JD,QF\Y^YF<^,-AQ+/+",R$ES_G:#?>
P$^CT"Y$1Q!8V^F]<*8O!EQH+3\D%1.5UJE%#%'5X-58S6>0!8R<C6$K:=ZQQI)Z*
P8;DNA\.;3M5JY337\FMR37CG W&KAEM>=I<,,RZN&Y4#H7?P WEO.XV[G*8$B&,,
PP&[/"N!.1Z40_<]V:@A#E4P3=K9E11IN[P,<NCU.T7LHS;*$ YY/NJS&=(*=SVR_
P/;2'O&V/9P6F#42R2>Q3=_QNG^S)GF>'3M%,%4M2[_W"(WX+7+QR#/C60 G4% X$
PA.@<WB546V<.79@]2\]]-O=5?GT/T--@U05(\.VEQN5';,7\TRK74>CT9Y=$M$$@
P O2">6_3 ;#U#Y4:(?Q;&Q^.#^PO<'6VO@NG?J77@&KY'/_$JES"QWXTTS;A(P$.
P-JHK^>J'(HS8-J=BGY4 8XI2(G3_6V6;*J NJI/LHV8,3;K##"FMH]:C0AX/NW[U
P^KG?D3:]J3T6:)GMX^86#W1?^^[I7U)(^7S".;Q'78U:%/#MI7@I,C41-/!;]>;U
P1X?<HF8N#M1 ;\U<[NG/[D3\5[@ [B6,$B>)<@C7],(MFI5(GVAI#S2-F>AN=A>O
PQ)Q9H96R[+,\"=H"[OZ-ZGSD8>XPF8WDS0 C1/3#]A[A W@5X1TGUT!1"1]Z$U#Q
P^.PC"QRB_XPA,1'6L$A%>NG_V>>U^NG':&Y[+0T"Q'J/I=#0A<=:H7J5I_1/0B+B
PQZ79U$3^4>L\6,]_$C\GC^((K,ZG$!:;;2]<6]\0A[NW'*9OY*]XX?MIY_"4^,'R
P9I(_OIZ$X7I.#F,)*[&%;@X;Q!Z]X_.V/#>/IK9_' &;GIIYE//_V4[_Q8U&R][U
P6"6%]!]6"UZ:HQ4DA&Z P.HXO&0-* Q/'-'P+?J_LDQFKQY.[ 6F&Z DBWU5 2EU
PCQ<?*0;HI4;N_??J F(\4.2 35K6+C,$Z::(OP-AFW(X-GR!H$YFW.!8',)V;Q9B
PT[NO8%<-W56SI]"CPD7W*2]X87_1MDPK,,NV@D%X.7RAF/>_:TI7"6%T5.[D?SYU
PSXBIGT_1@$.0EQC+;U@&.CR5P=I-+-[A&=T'IE=-0H#V<W@MW0<5"O.9THTK?@E6
P\7H&E&W$!, ,BWYX^S4[,Q))TU*!^,VV!Z041X77+ L_B"\YX%-'<D2<W7I^T8QJ
P_7I?SKW0'QQ>B, JY;'6T]&8R^Q0&WCA;2-^$>]W4#2US#5/94#(8*JJ3DCC4YC,
P30VF6<:^"]O-)O(1@S8#0^R'D6G@*:AF<&+W]].FR.&T3752.&G?,89//M8>Z\I<
P"Z*7Z7.2:P&P4O H6&.$FT;=A^]J2WJEV9_(OLL<8ZN?7,4G\EI9F<L_5)=MJ5:#
P8LAB6^.N3P0U8Q1DB=7VB"=X<J.F\:T[G>Q+,$SUB<&$3EHF+$ B&4^F;T4+91A.
PCKTWNM=8?4%U[ F(W'[QD0"E2>0A;Y)4X7SIUOMC( #+KG "@D)4H?9XMT#"E*IS
PMC5O2)0F=?_PNFA-M*!R?P3Q%CDY!<O:E%_"MIES469<%;=;8S$B+9-=$<^F!9!!
PH4\$+Q  7,*?TJ] +[BEO-V&@45$0MRA#K/3RU4($^E5CWVHH ?[-]J5DMA*'1]<
PBJ8R3O8*>*UT4EVK^4.Z;/$E<.5"\ZE\.840X2)-8'JOB87J@>9X-:9?"0!;IE4B
P>)@:H/1=8'@4V>A:_,Q<+@&C[,X\S%.% ,K,71R,N5D4RA^*4\.]58C/?'N>8+</
PU--X@"6S?N\E&WXH9[BR5[@E)6UTH8C56Q?-9;:(<5]'M'SK=-WJOBIK0*1A9=2I
P?)F^?G*UEHIQ![OT^<KC3D2T90&CG;ZH>7CP#.UL[X,#FBOCI]OKRVKE2E!D"5@U
PXF7.@BR02M/!:/HAE>SUL%-G/O_BGWBP$^SX'RUSJV]PL'SPB=UIYY:,M+PMH)%5
PHWU4IV+&97LL6^R<JV0BD2_<KU:2L^']"3?J90Q'MUCC%6'MW4[\&'>Y,V4W3MOQ
P>9!8]@!F9%%X/"JFMT#WZ[4KF4R_X;R(SKWM=^386]JD. ;]JZ":Y47L>L32JVU)
P>O$&7B>%7!"B!DHLB8C]#5=[ZB E:!9/6B5/R[O3S^'?2 '"NS))'X=]:H[84UO 
P]KPA("B :M'1[FN,S*T4DCFR<D3MCZ__*2, 3)]8]:/=3"M"_8;2M]+#R1EV].GL
P-<GI[F!),9XD:Z9P^;G=HFL## B334__ <S H]X<&_6-NKO,!,$9E_P(31*F-.P;
PC]1(I8Z=U[LO)2>U;L()E9^HDE#\RDBM6'QJU\3V=2ET:F''UFLTV&F+8@7;\T[4
P<>JRBO[K+-H_#5=$_C<4R!]RX9AT6!EPK]6^=7,,:0;R-B1:"9_2N]*ARZ=@4([(
P4]W)+H*FJ8NJVNZQ<9C'N,RQ80").BZE>!^7$^0[L(1O5;@#U1VH70N#]E>2F%BR
PX"B%"\G9FKDNR/F7A9$DB1Y="QT% +^!TDDG^7*;YE-^%Y5J)(X_E(6?LG*)N\'&
P*KRA;;*#<C-M8&CE=%*5M2D/L_[8?RZRBI%O:M\CL 9$?'H.Q5MQ]P,]_X8K.A/9
P;;A=.'X3CN9GT9]5124:*8+64;C\QQ.6,FP#:5#3G@6&CO=[+:.7?3D#.] QVI)4
PFJ'0P2R/@PF&#^1X(;<G[\'[^DP\MQ'<66G>47I=HLW)49]H9DX!-@F]+2-N(](-
P8U]8[&OJ?GFJGQT0DO)@7%?;T__)B">!U=6)D&'IB?#Z)3<OKA:;3Y+8W+R4W^N@
PW=0CEHQS7;-"S4'3OPU$)> OSSA[ML\ G0+RS19[W2^V:B[+\J3+]K+TSF65>B7V
PRZHS<%I]4"-^WM43](!U+,+_5D2M'(S0(1]N_TM@SWX: )6 66N.0A."J'M61NGD
P6SDWR#FY".E GH9[G0$'#@(*/R.-L:J/"M!MV9,!//H-[H!O;T^OFB,UQZQHKU"2
P<SBI!9B@,?B@!E#'!-@A>^6RA5N,J\C^$;EC7<C22^[ROB4R"R<R6[:QM[+F0[Q_
P@'/'\D-,$5[I$S$Y:_(1=A3@"Y!@>"\?@7WEX^ S+G"2H79'/BLB?GE9(5P?UOSR
P TSH/H%(C)F(CQX[75T*CN+._DI<45C:IU',I>5^D_33S!C7?]ZN\H5N(2HIS;\P
P-.1D5!4+\.UNJDX3>W0-F\],PC[R@]M,><Y+=?:6I[ K&  3D9;:+9D+T",SY_+&
PVZYZ1!$2QXK7<<6<952%JDH^@DV82--^O_;*LY3_ $%SJNR&Z"RWUK>L1[,!M\M:
P6J=!<EI(%#C*A#LXNP-RA1/$-RT!O<Y=NJEB*\1@N00506IKK;S1A!4F)8^8'XX7
PQ=8/=R=S99',\KG&P]J'="C#UOVH2Z"%^/L(GEKKP=(-STX+.-&)2J4LZE8S]JL"
P@IH+(JDG15M3<DPKV'P/QG@!CTT!-[K,BYJD8N1L[/(13^4WYYB$V-('*  \)^$\
P!Z& QHS<E$PX*O(2O J+%RIVWKF/XK5Y!EM[Z6F->+=5GD?'K]CIH.=MA8!44 G"
P(+(Q=<)6666C)LE97@9/D326KFV/!,67WGZU5LOE@GYVQ-/P]2"H9'--J8<Y7N" 
P<O-OI#&R2<?V4T9I9S:[_L=P-62\^=&[C'^,OD0A5E_J3G'] ?4\XFRXZ7 \N7-M
PGH10WIIV7/;U&@I_>LKDNVC.:#U1'U4E[;:%>J9\,#]48+*PWA(&9!5R!\:QJ6B9
P_YGP5[V^SF>/'S/KXOHX2_8"\.CV(&U*UC';V%)[I 8^9IG6*)BWVF2TE90V1S3F
P9'<U)\U"X8'%^;=1^]Y"%(GW__)+9$3LNCG62\@WG.01%/%F#E,9JX&.+?U:2E.L
PJ!\*O80./;"ZQ>X^>)>HZLZ+!!(;5N'L[CHA.8V*HSEA'1<E%!1=7O:9@'8/A;6T
PMQ"=H6#F19!5'I.'.6GB 52'&3+Q66^PD10>2O]NF2T+:VO!MN7_J:)%.W0>&L%$
P4%EEU(/YK:D9H!3KD$SN8&8)P<,Y_!687E^7'4HGO31@U)2C9%_16QD!:DD[0BIF
PD9&.IP-'J6"YV#1(+:&RCQ;H<&I&JNOU9=EE$6NP^*)2_C ZO@#V\GKEA\UCJ'C\
P[B;XR5.M=FQ?WB>=MU6?,RW:5OA0*P><WSR',1T%&B=V1=X+S0-B1^0B2LQE%Z$<
P%CK>KA.T3?]1+8"8(%*G'!4V$+=BE(/"A8S45EUH_Y7V) W'T#% V#F2?504[V+^
PCJO.6[/MA\$_]V+79,"_1I^@]JN%[D.Y2L:AFI1@(*3-TU(XDSQA>L0EA'_^&L]V
PF[CIT;2 !Y%[%$5JOKR<GC!]\\2]=08]'A45;N3EF-Y,I2-$4%)N7#OZ7$2%WQ5^
PZ+_QF HRD"N+IZGD47*#0,]_KPL^_<O<,F*,E@R(DO.BS):HGUR4(B/[<NX]CV^H
P[+8V>:[!L/-8SZ]I,ZL8DK?\3A@BN?$9#QR3K<0Z_^N7KV[+R^;2O'0^\GP0IDCR
P*R>[?-L8?NMUSXL=TSM).*!.#/^-#3,U2 2@UB=/AT6:>^<3A<*^>%_0!4+(:EM&
P0*^/B<V!UU)T/.35,C2^D?=2]8@D'(,;#1% .*^G43(<*QWT@.+JSM!T!'(&2=ID
P7F(D/##S#_1&P']JZ6T*P%5;P_\&HYS7<-=5^<@25U;AN)PBT"==I17";C1QQL:-
P5!0>A</M#!"Q5Z]L/D3SRJB3H7KN0Q'1]]P'?Y3UN:5$U";8U88A'CVFT*'G=N:8
P-,T2#VRE=L(QWE=+A;:-NJ5 6"60*%Q]F1;Q#7W?HP^I@J,Z+@!;,+S2H';;:$I%
PCCE)V<WG3P$KVUX&*#=GV*T5WU30#9%FQ"R]TZD;/?' A7W]>]1UT"0K&$@RZNM,
P;@"#!<<YFJ0KVIE,'!2.3098*6:T1PTM_W"E+-$&R_MYRT%JX+_24?:L*$.!-$%,
PSG>.A.S>S04HL=7(OTEVU!7%-JMMG<*V,"\& 0(RPZ \X!FFQ(6MFDMPK)Y_-R:C
P"0&&+_#5D9N))."+//C@\XQ\$-J.(G8B.+?T>>@ULICE(^\ZRNZR"*YFP/DRQ0JD
PE;VXT.Q,1!F8L5/V41=)FJ?R("QY\C!\%.+SI,M<A^XMF2/4+?@[E\*N'),&CTO5
PFG+'28TO5@#N]B379A427E+R#P4PI;,6J"^.JDS2/"*N0GM8QGT_7IM# '/L9V (
P$EUV"HPOB,>P#9O+Z2)OMTH;N-*[HST&@&#VCCF2%Y B "=%L>%V>/?O45!@P_OS
PX=R49?J&E-4SB\DCT&B:C^H?4Z#'0^B5*$M0>[V!#[T9#J(@I1)FI]A,\7:K40N[
PS-^'Z@$>YX1N6,I:DH3 9MZ$M.&,:/F7T5+L8QC/+_9;W0C@:M;,^[ J5!@'*1LD
PRQ^.)D7H'%F4!;W3/ID<;%>>BCH_YVN18O_;S0",E4!7BW-!IN4-)N:<:*>*8"L=
P(YBJ;=MCM)!,.#1<542PW6\1D(&5&QW,Y6W0ML+_9:B 8EESZ7=K%=%L9**:$.#E
PX)XJ#;]K#]B.)+6E=J86?""15Z;1IC!]')=B3:[H()@7,X# 8/'#P<88^\:5NF'0
P(N"8Q6]$\1+84LI.,2@!HA6O(7LP;S:G*4BQ@<NS9>7/G*WRXA?E=$$H@G%&GI8%
PBX<X"JZ1F=CTQIY<23N>'@W'C1# BLH!*1[C];H:UP(V_ZM1M0V=&9I7\4N0&;X9
P)*E%*\'Q_K[=!?F(?RLGPS)5!WI8.B") ,'#^,ER(DQ9?\]&U>2*&8!,%!"^&&LV
P$0/S0]@'X8'FGR$,7?2YPV]JO[YP?>V&D"N]CUV DT6# AX2BO5><U.2LHOY]Y_^
PA\U.CQI9X<S"7.O7_3+^\NQC'*/MCB*=;R*4T&<]C>J5002#$@X<1D['L#3,6?F8
PQM>&*UGO4?S.*J4HML8PU]($-AI&1Y_L6?.3+S!6?%$;U#$H710"Y@.8EN<*/2O\
P[38(DT#PA@S,]32L1;\!;916.K+V84@PVV70OL-=W<"I[*OQ_-)VA0G[5$.3Q9#M
P)5;U8T#G.4\;1$M-#6_=?OP+X>%3Q:VCY';M]8<BW6@/'9I&23']BZX7'^7L-+2K
P@);\[QW8@=!?1S.':6B?#>RP4^#P[^TS),$;FA[X<218/OIGF[Y"S8K(5B@# =:9
P39D^M)_UQ7ON'P)2U!8O4>E@^%-F/5A\L^MVB6684T?S0H';," $;N]$ZS7EI];Q
P<;7[1$R?;8;H??I!I2=L4+U(8W,E^/M7'RH\^\TRR'P_!RM\ U[4>6BH:]/E7$%T
P00D*^<P<.U3W<(,*7!'426'WJ;Q;N4-@6L"!EI/N$/U%D-11UU/LJ/:^36FR@GTW
PPJ#CA&4PMG0_X+.K=A93Q2*K'2=(N0C;<@5ZVJ 4"*-)+)+K@#.1[&B;L$F>RZ(X
PYN(=CQ7=!"7F5.6>4)B6^Z(9(T?$P;/@%MX-IW7CLT%J1S:QVN7'V;J_-/G*^GE=
P9*(F]'I1[$!YO*+O21_E8PD)#CA54/S8_G_M3Y#60: I[OJ<27#RS]XSX7L71P*.
P$.QU4-("VG&R;-1B!J26&XK7C[^ZU+@4G3>]MF!;OVM1\0$HYNAJ*+8%NI'GKLA;
PRU90"<S XJ@Q%DN$K&!+\WAH. 8\XK5N^*/I&RA54WUVCPFO%V)$FR?D+0 @[ZPJ
P#M_#JCBL562"WA@IM,ST>J)H=;#VK0&;B'+(7D#)99)>X[4OYG:*^G>4(W@#"OBH
PE*48$ (>8-M>MN%_7OS[@MAB6+'3Y]. <L+Z0<48530D<;V-D<LS662C14;X-E#9
P9N.(+!GX:Q:09/\+8ZK='+WB8X+W%JV?AD[3Y-. W97EGPH5A%UZK!M*9*:1PW8;
P'R/J "-F8+U< ZUD? 2EI:((Z7AIBJY#*,IK2JA=?M)8F)#$#_OLSXK6V:-A1QLB
PHR&&<]%Y!'1; J&I(M2_LYPHT:*&7;L2ZEE(U6IQA[BL3Z%#^7BL;'K79(SLW?Z@
PK@^V'1$ZZSBU^OQZ3-8@OD@A5K"]3,L# .P^]8S,U"ABS5_4/Q8>ZQ^[;^I\E7AX
P-7MI\+I4[7("5$B:H.$<LDTT*%6Q7/[V5IY;OX$34V?F0@5$;Y$A$8Q"TB_*I-/C
P*)F66[*XZ*T*LAT1^;F2Z%=*B %HA+TBF0(+8A(+;,T=PXT#U]: A&?A\ILK]442
PMC3:U;K@&H+R8F5&/Y%%P!]:V1\GHY)M) TE94,*(+:4\%W?6F;,R-'46^G"GRE,
P[RH8J*^:5:B15RNZJNWB3WHG_:8T %<>K.!*M8C F%-(L>V;U)O"*1[SG\MB'9LS
P::>TOS &@U=XZ)%L=!RN@[=1[F>8+?N%3@A??*R-$H<O(C*5?> 9&>0CO%3^$8"'
PT.;U,59H391%G#! (#>@K\1B$95I:DV#P3%/G6G&H*EX_KN,"G='>SRA*O]#):++
P9<@N>UJ@<ED6D_];_+@]KTB3H,Q<2JM:;_W@<KL*)S>%:*$[T>ZVMM*CYL'KT-OB
P,##3N8D]'W$GKJ$C66)X7BQ&[WL97LX[K9]7^&%N=]O.8_$^-+K3?HBUOM:=*?VV
P@+]\Z7NF<N.,F"Z599D=1JWB;<.;.1[O#3VFMV5!Y$GB?\7JSD*6W\8^Q@$+5 V]
P?D]2WV=N ]AW0Z\?JQ9MXSX"S:!L+IR!XUXA5N;6#[+PD"%U=<2K8:@O$+$3'.%;
PF&V)\S'_,0S::9VH?'\ *X+N#G"HR4C!Q"\I/39T4R_,N=0=J'IKDQ(Q)U0]?H0:
P@[[.E'U"CWUMH66IZ;S%FFN%L^F-&8@PWQ>W][[&;7)""J:Y@J69S*"<D(F.+.PH
P %K(PWSML&RMDYIH.V.1->>[ U0/J.(7;'+^R+RL]Q?>S>J'_N*VA:JOK>99!T"K
P+VED];/8/?!_#C=!DDS%9#C[Y"L)TK[V'"]",O//2\J'BAFL6MO&W?+DM%?.%'_)
P9;;4;\2/W[1,*YX6\Y&4IS>GA@%RWC!P3#N,\[4XS*O< (C&^?DG6,KU,W/RJ9_/
P[?5?-/H<S5G>@%Q*=/65?JVT^)6> M^K+]V9U78/AG)\,L'72:FKRKOM%[C 1-F$
P59(>SPZ#="[P2*:,0/^Y"D!+;G5ETS%=5?;OFC0)7XO+X9T0IQAZ.D4@\7:CZ>UU
P_ *]$@VSE_<!"$B_>$%7#+B H<'(F&"Y8:4[W<0-,9WX<VM(*WC/:;SXMDIBZXKF
PTR%&\B8&@P-C"8WMYU^M!$/<AX]EJ(/"0M99L%3!T09+5C'2/*R,.10K^OWK\$S3
P4GEQ2S9ML@>>Q@VK!'?4ZRH_":*)\N<XG +Q \R2#G1VRQC>$[D_'R (^) )5^HD
P<UO_F[W@2>P$NMW")\^1Y*"'N33_5 VU%XF?A +%O,Z6S7N1O:]('^<#582YJZ7U
P.0C\EIP^'4T$NJV?5?X(-?8VF%2Q=0R?.4O*H1>*^L7E.L3]K?WFJ]F@01H@I:+G
P)B,:[CL1KSZG.EN2[;)95 F%PTCHN:9/Y.AX71>6R+V][?N82L!]DN_G0[G(*U14
P/G4Y .] >9JU1WH16VAI99?3.K)U8JE)G'MMV?23GE"BL!>;0_6)<62VG1KR[U80
P(2L\T\39"V6O$HUPPL%NH*DR<@'EJ,"M5S;9^M.*R'"?Y/PH&)8%HONIQL=>4A5/
P.\D8#N70?%Z-F[2H[I((V$\V*[C>593&T,CR\" <_R'1)VLEG47[,S3Z(5&IC"]<
P3^849@N\TK[BX4&Z[(P9[R)K+EFK"C(R7MT*KZ-=++<!7G(S2#< .&4>MU:*H L 
P/8O]=^/)8J09@['X+MD:3('0#?93H=#]31/X*VBRJ/*:C&M=P@[#WR!# <?M<<LG
PWW/<L,.N"V=?&!?/BDS'%>':)\@6&JUD0K R]>$JG;K'+(##LG7:"M"B8VJ]L\M=
PIA8Z^*0%L1L?0>NN&'3M[N*G85?AEX04%/8/4OA+WPH#"C=!"_X?N5],/.+R#/QE
P9^0FK19:H+[-'[+I+13-)B7R0HZ>@+.&Q,+,YOBNP>:Y%PCX\)H#;4FC*F5Y/6L*
P$GJYT+%RN](U>)K0E97>)78:93FC)1N&E8[6_R:@]IF&J^D>L3D6 X 'Q;V8*^J)
P%;K)=189 ?R"/#A'_C#_,CXALT'D2CZ3(IL7I2VK)&V9&=GT,3WQ<E+JL"Y[F9P7
PJW$\O$C0U*$H4,G[,MKY(U-2X-=_* NY!?$W/I_%.GH<5</P+9@1=*]S"G#0O+-5
P7#.JMH",,4XZRAI+'*7-A1'OSG<B.T!([?EF!QW&HHN-(V,Q1XJ$]9Y$BFMX?L%$
P'HW?O-?&0=VWEL</]DK%QW6"&K[;$T8&$"#'9PUM.@ED.4/@%/-,_6HIR!-S9\*:
P'+]G;7G\',WF]M#@&%$!*99TLJA )N?F:4[MPB\>%_+F\,)^%JD1*UI<W)>;C[B^
PX;TZB,5<U#5K4:E-]#U[">2F\J7Z>>?78/?ILX)^6K*)%O_@93VFV*1:$(>5-=KV
P1U>=;V7DB<K+_URWKD0\]1A6I!L^8K.K968-/*HW8)E,+G_=RVGZ$L5](8O8:D@/
PUO()1S+5J?Z@O3XK"+@YU@&P<25;DLT%4UJJ*1L01\RB$TAXOB*I3/V'Y\QW2!BC
P0>\O PC(*$[FCJD:IGM"S<_KS4EEW%]2N1F\#+/I$# .^*RL"O35\;YOF4<-D8#O
P1W%/8V=P& ",=J;X 86@0B/DD@CYX(G/90+QS*TD[:I)BOJSYO^Y.*4!*+0C&(O^
P"&M/J9(J54%MEBLS84K I4@UA-X^1'H:Q%\B/D1M+(1_3\Y$K<^EHK/5G0'9KG&,
P5!-XS0C^G4X::>2*\-* 3Y4"_Y86L=1QBZ'J^R>9(W;=_4>@7&CZ"-)??9-1<!@5
P)F*ZJ,?=A.H+]VFLX+ZQ1<(<JF]*T,BU16UG= B297ZE::"Y=&DD=L5>!]C7UK'L
PH-#8(D ;[0R-="1NB*N=VEU,*+J$L6GN4T>6+P[!^HSX#BD#$EO)4(*,LM=2NQ\G
PB_2^-@6XKI(O7OP?)*E[V1 F\&9K5LC(IK]Y79UU$Z6.%[&*2QXV?C^(X,<EH8G\
P>^9WJ9/)!7^XR/8\/T51JWAHHF)L>=J64+ZCNC6WL2*MH IH@'MS2 - H,^M5YQN
PI275M$6!XY)/;X*1J;51*C6?>*F->3JPNRG?MX)_;[99++I\:AV&MJ[-L$1G7?S:
PI<B-4B@XK(LD7&#GL:%;7(]7/P6!(O0._Q\2"1W)'G48]-[:IHZ.7F6I_QB[R-OQ
PP-D738M,H710&7^07CO(?@SPNT'2-QXM&Q#A% -%7Q](8G\#1?FF8A?'B$Q4&CJ/
PR_/[^!]5D[V76M/2.A;BX##CXK%$%I%F:KP<]>?C\V5L D)D$EW[ZLUHYEYPS2VR
P%R-U)(_6%@X18D2D:*FPJ(T\I?V<^=!Z9'KD*"E?C=Y,XE=,$-8 RB[EF<S117MV
PSV"7)[M/J6F'(L-J=@@:;XVFV/B$(H=S@NG#D8'1_?L#R0[00P= 74J^,JA=!E[Z
P>2!:"+5F/_ZD*0)2SI CE<D28S=*<Z7CH(B_:5<%)Z2&_.T:H!B[KN,JU6RN*U>!
PSQ[+43+&23WDVST$3_TD%LS30  "U5,;02E.UOH=,[AQ6!&EY"+1QSSNF@(<HGV*
PD?<1KW7L$NF&@:2W5YJ7+)X5/,A<(A>2'M^>=6@5]CJ>G/:Z]LB?(DCFCQPLJ".!
P(4+V%9!M[ML4W@('JL-&WH06R(='O E9<+$#\;A&_^!5K,V#G\\AM12//_2V%9X9
P"W84-[Z[@6)+ZV/N6SY$E--6?9EX_W9=3R+8E,M[3D7\$B+>$H,3=P M-\!GYM>H
PA"&FONL&AVC+[5-2$2LG(?"AN@3L ?# G*:_[?<+T'HH[\_C?\-LD@(\6TS_]:>)
PE3FK7,_:6JWRT:.XL65Z6P^]L@(6^L6L[Z_BL?X1SD/^_\Y4BNMB'X\M]K<J+0=Z
P@33,R)WV=N&?:VHWS:%RTP^XX%F;]<*NM/V?[-OBO3#1"ED*;M8A-M-TO<%WHI7?
PR\A_FX88DFRKEV(*]A4RQ!E=!)*O5";\5:,;7E[ZB3E8U;J19H7.3"?MAHV3=RS^
P75?"IN!\<)N,WXHP63;*^82-CT=6^D!QR3C>07]N[H@6LUF,YE,3IQX/.A^";>NP
P:,=@!$L8,M)VO+*0UM7CAGVT:;S6O0 F*4Q!P;3.C=C=W<*6(:5(R0G*[,8B<P.L
P@6FP#DS3^4T(&L+P(Q_9KSTU+!DXF6NQ-(A021::W,$=(Q\X>CB$O##<H8ZX^9CV
P!P$?KVMS##3G$W)A7"ME%;?>:*@3AB&B>7\ZW/SY_@G!:NL[N58>W(4YIL6V"*K&
P&FQ!O5>>3NA72MAK%"RE -JY$";>,+<$[+?!NN_4U4)X\](]TVBECAR'CP+(I7 _
POU-G(FG)E:IVE.@5)2CTA<WYP(U,;7"K+JUC0ZCJ'?I2&>A5-;/D!Z65<D_-'>39
P+R9B?(&U))JRH4989<\($9](+X]H;=FY(87J#F@P_M'%ES]W2TY2[Y6$^.PDXB4D
P"Z68_NIUPE],N)(0871]*"_IP&G+L^X@3LB+&6_+5?,Q!0>W016PBVU"NM(1*1HR
P60Z\A A!T;8Y<Q6VSW<P1D7 =8)TIA5MB5UL?\Q@N2).3B733\ETN>C^M$@S"-ON
P0E*JV-&]5&[PS9DLO,_HKU7W-P>/>1R-R['7@DWK7LSMU#,]$&\#BRVU;Z$,E;K!
P%/J1]B(%8W:8&%F._-= +A:CQ^<F^ 7>S0B>P^B<KTX&TD+J(O[+R.  ]3?AVZ$:
P7T5<_^]-  78]#ZO:E>H,LBO<9YE::'-4(1LJ+:R>VCB[Y&TDK*!Y2$ ,F INFX<
PD=-380L+#1[/P.W0MD]G^AIF1)1S*_,@'(#I<"4#:=K^V2&F0.=#)6*K,\C3PI>-
P6+[!Y2_=:5E!M"">HW8$C0IZO\67XT=?MB?-8)F\O?OGHQ\[BZ#7.GNC'?T^W$OV
P/3S&X3]$)4$QE<9&<&8'/5?(]:6;49XHVYZ7G"7F.C3"HI3L@& IH*D9'K6,2?-4
POH5$1Z("QOK-V&*J\<)[(; T^<@:N;%3QD_@(P)P M3YF) .O<K)<Q"X6S,+,.%I
P%=<%6Y$0)^NS$O&[^2* U1]^N;C3VD'!OVPS$HZQ.O$C,C%&ARTYNA=$M?#9X,[*
P@BW0U9!Z#.Q0_)D+JN^;& EW^IU\-,_ 5_)O$LU)!A):N7>1QI:EZI/U4G7/"7,(
P_[#E#X1+8&@]\=FXEPV7)UE/A_*;[L+9+3T O\5R.A]DF>J&,DEV+?A;2N$CC>ZB
P)&0* H7/=KUA]6:Z_J07WX-W- 6=SLHG%X]WYSQ@%R#G)_IJ*23C%9OUQ_DA-4T$
PJ<6J%-$"BK'$T3W8:N[:_F_SW8!>X6^$O#XJ7+2@'G6OHR\'&<']O<4'2H"!6J6#
PV-,4D=2Y1I(O#>B&D1<&_3T9RGBSM#?+U11,\2*96&$ &(+3#?'87^4-18]?\=KK
P3=!45(5&]-S1WS3(5X>0Y87F!(!Y* 9"XC("V>ZAX?Y-DCZ_6S^R">N!1++,FE+K
P/<2U%AD.;_@TO8U\8Y]I2)1.9)E(S9.N6J6^F&^>( ;Y+L2VFI'=2V38XA'"B:K@
P5WVO1P=/WA%VF/XVA*9W,C-TC@)Q2 42T99?C+HX")X]6"[(V-AF%%60MR_>6V?"
P?LQH=CBW]W9.AY\%6K//=67)C[\"4Q<5C?=UI[5 %XS>,:+;'9/_Y2V;B^S7./9H
P(S+4I8-\X;1](Z@)<8:["W$;DAHCK/?I.H[RBP#MBB+"63H2LQ?!:H"'P]1)YJ=9
PHT[L75]I@!#7+156H@52X?-?K_S92<4]O&UX2_*S^9F'(<(@'OX$E0DP-#]83 K*
P/2#2)CN)ZIT]*:R]XA->3\)R<\]H^A)K801Z?[LK2HZ7ES]BNW+[;\?KR:>@]^7_
PQ.U:-:(-?9.JGCA&JC>]R(FA2AZLN$\A<5@+C 09/61S;LT2(:&P.$OMBMTZ3?F;
P!/O81H$YRG5#](7D&##ZU_3S?9K0>B=Y7NTG=Q\B-X43=1Z&\_6K9'P?F>[U8&@)
P@A[E#<]$W^@7E$YT0%!)7$=/J_7* ->58F!!Y_)\1:/PK"8*22J4/FAWO,@(+9@K
P=B+->^%28J_*+, $M<&TJ;_'L2 G0X]W;%Q\Q\U$)Z)>'(^,T,#QV57D/X*:YIN.
PU">V*R L_L^1TIIJD''&,S/7S#/"%TO6>GN-$+@=CMPP47=V=+B.C/%7<ES#G %Y
P$FUU%B&VV/OFP[^6'5919?,O\Q6;"%U6A=3Q,\R&41=W544W1,XO$BJCO/FL7RX:
P;$$C;A0&2R,C=E:*'O)XB!]JY6AO>5?_B]T4UZ#MP/S5W5OJH)N<G_.AYSOPV&M0
P%-8K9.F_> 15:SIW(X',-R#A%E<:K%)BO;>.Q!6.\#69K<8;^)WOD0>ZZ]%>/Q'5
P>K/C12Z.K:QO#A]"L'] L9;[47P]M_]^I7Y5\^'<0**'H+O:TIGLA]V'-]:ILU=E
P?:#C7Z!0'M#JS4RYY<E\8"2W+M2\P:3][^ 2GO5G?6'$%^3V=<ELX^: >Y .NKS(
PA6#%W=/C5^>7_DD6NAY<[]);7<Q<V9/"12\T^):PJ2O<@4-J],DS:B(SMS.AE3(R
P$,>8L8/\-DK3A72C88K%Q\%'TD#=6'RVZWRW[I56MVO8]0=[V+=5A(H/YV"A;\R.
PKR=/V;^6D, 6GF?I6JLLMFR[>78!,$D!;,::B[2&;"F0^^JF\0"]XR_L#;,<;O(W
P722C$SZ$\VI6GEVHQA%7*N!F@:G(1D2N[K$C1.ORQTJS7'*X-2=R>M6"U);RILZO
P%7<0U.T$CRD*&#I1#>  3T!2A G4)3QC4@R0NI?(+!^B,;%B-O1++5/FGA"7%5F@
P8INK\3FID?1WN^R7_3SLS$XWGHLA='DMQ7K>3P9F%5F/"'\D/BWWD)V_H%,&7]3 
PAX[PTE9%I<Y\&"-;M#TKTB=-PJ1R&T2GX\\:>'W:'.*<A&)KRT(<+@:1\D_\IR&T
PV"80_OUK%&_E&X_)RID?+-B2@:[1\;8"+9+'A$9<_XHYR"FJ[0V' 96M$AXT#$7R
P<&<;O>@>]Y_JA9H6?6Z/4HHOU3D\\C8[I-"6QLC]HY"I[KT$+M% O?_<E'UEBX=[
PH-9A=,>Q=:$QG_TAFPXZ+BTG-\V'%)B$!C7&JT6M 3<"HA\ZWY"Z<8*;(0<ZE[#!
PUQQD@_EU*5MM:'L*;1X/\3PY7-+'#YA FA*W(U/(X0J'FR'3>&UX'<Z;="M%M-R.
P,D;%6+#:;6$0[@Q=%-9NC&8+SB_'!8H&5&!YK-W"S#X1^/E<'(J[7%!RUM4*$H]S
P"+1F?8/"<+.X/&U7$7>CC*A!,]_$]^P1A[Z<<$;9IKJ%3<+"7!>PU5Q UWGWR<$!
P+"*UXF+?:A2521P(Z\Y\WAYH<9O.F1PU$I\&A1NWZ(>$Q]K"-+F[EI8Z$2'$W[L1
P%V6"$#Y7C2VC;C#W >DG>CWORVX>^D.@U7:"_@#@/LJ<464.[ 2CWU2IO-0Z?.@\
PO*@0.\$$PC4H>?/+H\UODUV?S!.[+M##G+4!(N^O\1,H2(09:,3 X'@ST'Q0E_Y4
P&2OR'2L5=)\-9&((U&88M1#LC_V9Z@T*N4ELN!H+_TJC2A%0$GE?GLX]5:S-JJY'
PQ$X #_O)SU41EJ*[S8'?MZ[6H/""9O'FP4VYZL!3_07OU-PL[4'V<FC,_+)M?J'E
P :,"-2D^S+[00,^+$?/N'-WE)1-95*'/W_A>YPO$>Q;A_>B'C'A(2#2 M'+KDX=;
P9V%?Z@>I&LW\T_?L([,Q!*$C#<I^).F*]QR_-]&#<3=N+27+$?W\:Y3ISCGL0/DE
PN$'GTGF6SKB"?U6O%7KED$E.WT< /&5/'DRAH"608+M':.O+$M4^ YO/&*&IMK,W
P;1CS+A<_[LDR-H/:K1@8X59643-ZLV6>)M,LJHT6'OHZ)T[U]C?X&S@D::1&]!12
P>BR@B0]*D)5A8:(.UZ@0$]*AB1?XR(J$'E"BNVJ 4.1:<KQ!CE0ZKS) +V_RE4SR
P3F?7(;3%9<7JU;/Y;\RW ^;*P;;MW X6+&Z"+[NL.;<OF$P\ M[";.PQXKYBTUBE
P2UO+.6.2&9WX$P J,PJG5(V@7*33K)QPXR)S^WM.BGHU=1,VQ<083"D!'+#,PDZG
PD+\0U^XM:1_JP)HCD!=.=[;/!BL"$S+EU#<+Q39BQ=AU_9%4"4,QD@C16^TW^SWJ
PO\D?VYNU8&JXW.&K].H].SK!2LM.7EW&*WM 00$==(,Y,/%<48ZO/_XP;WEQ<I;T
P(UNL/Y\:/I;A'2P\Q :HF@O-*SJ*K(HG<SDX[)NWW7E+N:V?F=<6&/(QZ,J\H>WH
PET1O9!6E=4NJ:K@3PL1?)IG>U<V.H,.T,M+EKAZDA<:[".^&7_<9_ZX\,TQN<@M]
P5<,;"O[K_1CXGMD.$ETFCGPRZ/9OE'382T,2I$DFO-]G'#5!T\NE'P/7;/SC:LW6
P0GN@^_(="6;U$-!0@(G6NX(XTB26%PQ:'(>3P?MG4, # C4M9N2P=13$37)+5Y/M
PA@?"6O<_,!)$E9X5,4_7O"U>XCM>I7(H:U4%E('#(4FNJ;<O['I78P*6(]M Q"?X
P5@8GF<$&% \A#C;%]N:*7KVFM)C=?46YQ_F0XQ%5WB>ES+#*\0#S,:,[A64.3$,Z
P+,YA1VYM:ARK0_@NU25*Z"0C$?%VK8]+N$-@;R))!Q>AX46^@SSWGG^[DQ+X2FL1
PI76XLV<TX?_.@ TXJ3FO3<N!Y3M2@!)59@&;'DO$R%[*,KZ315,94L9S7Y:IG=L?
PP@[];^J?'7\<%4#=3IDK@/;B_A6?W ^Y39^9@Y0SZR_S"P=PNU%/8(3@%=A\3[VE
PXNHDJ:J8_B_T"R:2->5><#VW1;?HC*%V%&J#+.:X*-MZ\O]<LQ=7CCNW2HRZ[;G!
P!' *RK4ULC&[>Q#:Z-UB&F3H [M4O=#$FA43#\Y;_E?3V@X_%>I]F1+N6 VR8"@Y
P4A;:O_S/I:30!,0-CW,DJP$WH5&BA6I-8:=F[#C&*8%%PHL"^W^-]S/W:2]"%!<O
P+Z&%B6CBEZRZ*=4 DPK>A7!U;V= AR.+#JR/:K] SKZ90MVCR5?^S^*^FMC(+Z8,
P/.P6E8 "$C S75+48I%&4YGKAOZ35W#@Z>DS?X*+S0^ ,$CWQQ835\EQ"#1]BAJ;
P11K)]:?%)[7:ZX& TM[S\ 'N0KC>X3*TL'#/9XLHMM;3EQE917ON=-Z_O4]:(S7?
P",3LCH_6M8EH.D+Q 2?"GLQFJI=9X+^RLSP!K%H73J=HG&5L[YSMM^S;I\L.LQQR
PXM# *\NV0/GPTN:0?L[4:"XN? ^-_EO0PF"F=@ )NV#%=9=1Y]:1!#T2^FZ^746:
P%""R77%#B4OK1&0F8N05W U7XS=8%.ZSJI9QX[9"%NM:F#%:F2C/8!ODAZ7CHQ+'
P>:XH3;M$X"_<S3X)DJ'H-=KE 9.8AW5^4EC=SO?O"1R?ESA:X^W>3V!O@R5L3CG:
P5&&;@;?#9N)PVOD<'R,\$B3T!ECT_XE8?!*[ADQB4AJU@^PE%KRWZ47N=").FV*/
PFUU,F6$Q<PP^X?9W5^-ILLM1INY0QXZ^G+C<*NJ+M.7@%JI'/]U90-"Y 33U:WEP
P5=9+XA4A_1<_;FML1HV#M0?2^(.GJVMZL!W(DUDCAOVU0#7TKJ!FKQ=^W&N+I>N:
PV>+6 \A+ $OZFC^&H5PM'S+?P]BZR"K,I<Q0F=;>@1L##)$<&7.C3<@[L4L>_1DU
P7:CG]6#(1JL]1+H/W4Y%& 8"[0/[!ABH#(]^Z$Q8OR5\VL>OX]>?VC11N S<U%1&
P)!XZL1_.0/BC_M_EB4[\#( DD:N34 -BHY3/FVJ!"K+:6,'H-/,K)[]NF@CO5AI,
PT%0=/IB:-!>1O0Q+#:+9/LC<1U&$N5,WT?2?6;>=$AAH^T]IG:.EEGJY@J]2&,;Z
P*ZIY@=Y^+%QF^\]?"O\-5O62'_546V#A?#O$'CZJ3-%C"@/I]G&5R_Y4L*K$>YH^
P1??VB3T46#X [D3WKY:'/VEZ!+5/NNA+U5^ZHB"KWY>8*6YZ_F#0J:"Z2O"R^+.P
P6]3R_+%)!%'U)3P0A[\QG]I W;_,5R$8L[_@M0I"'^[.[ 0S07VA[7'#,?+K=1<=
PJO L6.=[EFJ-8J+E^=WYS[$PHGER0M!T &= O$M*C].NSF."%F[6R9% R3N8:R3V
P0SFG<R6%DYY,!@7 WN;MV:$=M&UEWV3]>^)EG?&GK4ZV]O%Y9R@Y%+D#2$2NW"S:
PU$<$E7E-ZKO)J=GGP>NT<PXDD9^XDE0)#-F3\&IP4',/E="60F8A@;/$(#.3<KVA
PD9J^@&^0,=3%;2^\NLBX06+SUC%R:8-ZAE_4+W,-"$ +E6PM;$=LK-%X/<7@MU_D
P]F1=$7' 8^HL%&XHPX=MYF*I+5=P1\W!/.F[O%<TK8?-:Y[*J>:"0XR8GRT0P3?S
P#1I_QR1FOK+\1^;V1EPW$A.V//P(:YQ=?<[PF2TFL7\BB@CC3GSZ#X[I^2#\Z-\3
P8X.6-7=06I9\[?OQF&ZQX;O@R^0%-\2#-HT\ N*Q#CJL$#+B30CI!4E7*(L!Q>S[
P(%NG?;84'=H=S_UI6A6K5]@I&1@V=BT4^&(((_(FK>IM0]C#N$HNB\:!)-VE_*@Y
P16W5(]:K;LT!(46$U>3$1:+^4G^3,)2"^R&U2K)#$N-<J7$CX*II<(U2:EX<IIV?
P6.4&[B1CO9"HVKP!-+C-QQ..>>SPZFG;Y>B&/XN?_4;/[1L@-@GB%ZODK3]/_56$
P805-H:D<,')?,LQ+K;B2R)6L%OK7106*5'1QN4A]'"X$(%[)TD:M$%=5;5%)^C:]
P:^V$OA;J"'/Q*[E=(.I)U6O<E@-MR/.L"Q(5-=GS)]QBKSX"J\N;W3\N#)F@:\PY
P%+F0F:7>$]?%BQ%V3_GSV4VY0=0?US1K1#,^*]+_Q0/(56MH0VF%$7?%1 D+MP_M
P3GFB)#Q:G<1)%4J"(ML65?]OL71K"SB-6^P"HN129>,@F^%4^C*LK.BQEXR_U!,X
P>+9C.>-71?I(?@3;11LW"DKPPU<@O--Q=H00$87V[=J4*SH=$82>X"] ,TY/]J@Q
PI5+C&G84W>=SEPP[ZYUZ9\(E,3./69N28#+8S+>S!X/CGP$/NOHQ28#;[AY_#(0_
P;M1^2M/, %%@R#,,0RU_L<%([:NEE23E?R;IZ=$ZF Z&X.D CX)25A*-1D9G/0=M
PN,IR+R1*H#.7!7JJN<[W#]G#V/*8VI!XQG_9.9%#+ZH#OLV$70X)>UIFSP/.#*B2
P=MX&S7.3_P$09TF>]0_]K-RP]4O]4&^H]_; I7%K+/-]^,/A1) :(N/1(R,(@#G'
P%0KASY!J?J4FC8^C,W"0NX^?\OXA%YNF!=&F1>S' U+R)1Q^7MO KGO;)G-^X;#>
PAVU3)'8R]=X4>HQPKY$P^')!0"3T"[;1 !GO78?.6E40S,U^7B2ME6W**AQT8K9J
P15@=L;"AZ!H]B<1T\8VA-P&WOF8GFF02>I,C/#T@&OK56M53M5$'*=\1-YWY8Z*U
P//P.-+7HP)N.*TZF\&&%: %4!3Q&X0F-]F!V9[2 DC?21^=:<6G7@FZE0DW[$VQ%
P5CA*TI$][-B\/Z O<1]].(38>J[3X)P2X>IPBZ&S#[JJR)9"8^C613\8WR;"!TY:
P&A@U#,@;:88-0>XS:,%C/@L;$6>''\,P'Q.'R7G,GHL'=1R:X2Z;QB_2P5^2>V2_
PTIO[9HOH[;3:L^77'!]IN"9O,46)QI2UTIP72E2)E;3P<9!V2X/9E<"<Q/9BEQR'
PTO SA>W7]:BPR8;/&KW.)W*L2*0]EE3JJR7>YJ;\H9TUY;M0$X&4_5NXD@"Z*HYD
PYICJE/2-?G^/E+R_.5KK79@HNDR<.&BV[<Q.90L<ND*V-06*)0D&J?YKE^'RU=^8
P CH+\$UR#@BP(-H^^1YX54[720V%.83.%Z>24:7TZ<%C%38'_A&CXF1?3RLMQ#HE
P1[EVPEV@ASGR_7_,K(>(&EU'(NM:A1^U"YJX?XJL"C:1-?PP4J][)H7H!Y::)$ ?
PT:K#3BQ?W;Q+5=;=PTXYFF&JHM+05\QB&2I%<@X:_6&XO49*4-&V'"J9V-\U&FH,
P7.]J5G+&F%2_H]?S"HRO(M'.2:'*9::TRC(7T<U8'0I42?ZYVD7-$$6BY/Q!WOD%
P*G-:Q+FIV(N!Z&Q>'E)<$U;U2:@NFV*!Z8>!A-Z=:.._OYQD970[JV'"/DQNJ(AI
P7S1_9+\<7A2>/^Z>@3+HRJ/VP9])# !"FH2PW(L[!9CF0,7&P]-+,6R=TKDT5/8U
P]L]<1FD\477WY\<7.OURBJD9Q\JIPT0Q:^P@F5 1\'Q88_Q>6?]/$5K[H#G(]6F$
P@)F*Z8LL0[;5L'1@FZ#(H7]=E-7!+Q25+V,3518').$TK3E$"*= ?'L:SE+%E & 
P(KJ:3J>B'5O*$UQD:<)RH"%:K8CO,ZH1I'K,C3FNK 9+L*CD/YEE$D@#J1GZ9!IW
P'&.C-)[D)TH:.>OE58/$?WSAR,AZ.C89UF3O^@5YH($QLH5&FOB5_,//$X=X%T$8
PYM %*ME4M[D$=H74."FAC,156O(]<5/*J7]*500(2[%/H^L5@QX!0P&E=;$MUE,<
PQ(:>$/;@) X#_@"?1A$3^WY!_=%7DHNB0EU6I&(Q;9/ORDRI -P%N#CVX(0BY4F!
P+PID"]<710.+<;S5G0 %4S@I)!6LS=&W6.@>CB;M[[3W%_]X_WF +]DF2X=\.B$5
P$B] 1'9CW+-D'!)/J]OCLPDB75L)F /G=XX>^+V[ST6;H6FPXK'%H9PST= [M.U6
PB&>S;!M$!4_:1GM[FB4NLG40TAJ&!?9?K:<=R5BA'DD]CQQ__F&G8)V;.JK8'?B@
PEP1KB/\II]K\=CI:X[T;-O)E0"L!^Z;.-1IYRJ_)+V0I*2!5\]K7,D>@ /.^#CFD
P>P9<8%^N AUL^EWRM]C]&SDEWS-QSI ;EGC^Z^&X<R.M*.F<9Y!  A4Y=5R"2* Q
P7/5PK,[FFFWJ_M3':;9'LSR&.3*;8FR,I\\J_FGZ2Z2^F[PERS)>P*JRM)=8E*LU
P@0KMG2.8M$YY.2.SP^IDG 8(?M>HI^%3XT&\ZHX49;OHGNCC""+2FS)58/<6HBF[
PMHQ9+C0')0_<)X5_IW%1G/9O@ZTQQAGP:Y')JY8#0F8*JMP2RV*,$%VX&Z&<3L -
PW!JJ'(::("K'OFOV+$%PER:\!ZD (^S+"=Q,Z#DJ:S[>9U._=BOJ9#^ ]IK94N8!
PK>Z11<OAJ<A2V,'(!DW6#FJY3FR)J.LD/QT"W[-D!R0Z*4,$9:1L\GL63&(CV->H
PFTR$&W,.EH=&P@S0-CW/U$A_.\9I /0K]X:W-WDNOL):$. ^Y+Y#T5??E@&K5O:W
P0(?G[HC@<PAK3'*(H6L3YBU\'#C%MW*H\RFTJ_/6DV6;#D3:]$!Z+!4!)"EQVK=D
P;T/%G0"+?[ZG]KF1 :7ER?ND93##K9H\R3PYE0I,6:QX8GE[#$&V4CFUWA>@;Y2C
PNF@1+YYYRX_ %R!HQ#_OOR)ZV[MDGK:+FJUW%/G1<N,*&:XYWBJBAHF9VK<O76-+
P5/QBO1(/&((2N.DJ<*NI]/H%Y@PPE5&?T<R1T9TU"$??;MR@,<Y+#BI(1-4/8??+
P<&>?;F*68\A RF9"V!*KJA!NT[8A>N\RB5%0J R5.6_$M"S07<JR'GF_'$ :F2VX
P<*#Q\RO]=/- <=ES!#8?21)@ES@K<\X]>\AC6/BG_=7,FF%/54EJ2R@44C\&92BI
P#@"?%NKQ2.\ QI7$6 "/%?/-&9F&3Z6/&9YS^WBTA.BJ)_>T?)L@E"4M=2DGHS8R
PK!F">&(O'->8&A$4QK?T3]7*H]#4K5,0RNENG:@8U8V9I( ; O2_K;2^KBN5C;H"
PXM<H)F/GJ<@TL$3P+8:TZB?DN^1V&-"R?"^P@5\>=J!!16^F9]'7D)@\2_RI[W^Q
PJ@1+ZCZ;?QVHFPW;E,,"AASQ^LKD;JD07<WM!>K[7ZCT;TZH5'0'D([7&.UV]AM9
P7(#8':567SUKE>"NXRRR=!(<D>YS.=@-$<L4/UC/A/J+*&=*V# E3&M5+3TG9T,-
P3:4O&A'W+>\!M37>O^7<G+ZRA4RJ)*O3-)3U@6J/K6Y7VL!",@@K.!7('*&^,E?U
PE&,1>Z]O4:%(T4L#8,M,P<<6S8LD[@;N^:W]ICY7N5@M!"Y]4PU=J?X^SWBZ55"=
P\!6AO4UXNM!;&6W$8;'Z[L(NC+$#/&+_)L[>J,T@I6XM-!9XLLQ()VGK5S%MK)GD
P TJ\%:PEM*WA6FNQROS7Q6.:5+I%-7S@".WXFSI6K:Z^$WDLJJSB-NDL%/^C]0I!
PN&E]]Z+LZ"@5S.+?*B]Z.*ISWM=(Z8PL"GPG\B86_FOO&S>? >MJ1Y<@ &BBBV\Q
PL6L1\;=U^&[.4W*[<4Z4T<8KLR%E;EP-S=TS!367!:XN7ZBYFDS0N,X J^\-\C$ 
PO1IH-1=+#Q9YRRC4F2[JW#F"X'+-E3*'A'E."NMISV'>0,W,(CR,K_'&LU@Z*_1A
PLGWP ^L JR(M .H_5<>?U5;)J05(/K_TAP1TLRY7@2C]J>:*0DW<=YW9R[WX4H\[
P$P2IY.F BXHV?V@#%P7*"/7U37"G:.%)O'R4KU0WJWN,HN?@"<<=J0U ?'ZCC-Z\
PG@ (&; H CE,_RF6ZYW7*^+"F45))5)N!.2O]%R :6#UJ_%S&A%_LIG0U*NWQ?PU
P/&SY&&"[\&&!:@+0GT>WUX9:CY=+:[6[T#XHG;7E;_\% !$EEC^@1@:)E1P,Q4HW
P/4^617'6QIQ2?X+.I8(B+*LY93@_;T<W,U@4]-IK$BW;OQ#[@RK$;QAHPARV=,+[
P X."#?;<7SD4&S_1I:3]N8+F1+C%EF=U";N=E@1 A=W>*HLW;J^0=='N=5BS5;7W
P-? +2UM_,HV]:&7:DTP1ZF"K2I"P/7I9UW_HY2:O(AIO0.O4"#&K#!GCM%B8S*@:
P1I(Z:+D/H^@3MW)R0+D1U#M<V2=:]7=SHKTFG@58_]82+.C^S(1RIOMKLW],\0U.
P^]>%+#W["\Y:PVPXA-0T:,6FIQ%Q:,+QZ+\MR":F[^E@?((ZK4Z (7<25*DU6])S
P4\)2$U:GE60,#8@M57"B]!+.L74_VMS=S>9:B&L9R.Z6KX62Z!3*Z4A1$&R:-Q;+
P1)T*,OCZ5LLQH^4_!@!XQM7=U@C,8&!$W'Z_9T<$P3,P!OD4P:Q?#UV-OM6U \(=
P?M .AW/-.<]=$%S+EPM?LJW&^Q6HD^)@!L1RR95#YLEVHY]VT/5O3\07M4A0A%1V
P:R;CK&YCD$)@-I$LY2J'=N<];"CUHO1E?;3AZ$WIX"1W+TVY,S:U\!VV% 4R:;33
PAY$307V=BN5Y7LRF,"+)S#EJJ>C'WLO57#=:[6Z0C]F)WL7SM)59/JA_T,;R;%RG
PUE/GN\107PGFLL],Z8\P8$H4B>^CDDTQ7*L$\Z#8 @3L;%BQT8ISLV<(%R#_>-$@
P+#C1>HAC:^? A\FDY#-CK[S+R=G+M\C).6YI [[C *!8D>8M+^(?9]EM)G/>0NO"
PMIX)-XL,5U<GZ&-,[?\0%1C[UK-ZI^%088>KQ5^*C:E-]<\:V_+< 6>=C-4A?!&,
PF[&I:UOL7"9^."%S-]JT'K>;13'#*+$&>P^/V81M+<Z_^#.DO<\AXN!\/2E]!7WG
PYT_/S/BN2Z8K7/Q>$JZ37HD$6"ZC(&MD65NZ)+24-U%1ICM;\7F:<HV_1XXC_Q,+
P'8/TJD/45E?N#VP4ND1L[X\D+*C&TLL$ ,6:!.MP3'J@9;0!U[!T-P!1VY!P=+8S
P<C<T(VS&-/3#QQQ\B]'PSY.:_'I5RRZ[;6=LAW8I#X%0'JB7M@<2C.68*_:8GS*N
PZ7L"X6.@V/ >8H=RE+L]P,KS2C_]I-<E?'NYC4E=B5N+[N!] ZLR1YHDIHAGFJ=U
P21R[AXFCUZ[A42A%'J/=8;SD_1-.1&',7W =>@_8;?3V3@#0AVB;/$.F8,?@L'G[
PB,6"4;W,L*[^HD#'CA065EXW-KRUU!Y27_[4>A-:S8!.36D,09[K(G3,D !RR<B2
P)GD<^F+.IST8$X; ."5OOVA\ZQCGC9C6VLU?,(&TX)H(/3/O8]*'H<#["[K<<I1R
P8)+>V'C6)PYGP 25W45S\GR*FFF<$KJZ[B&%+1DW2];"_2LT &+,G+)VF[UN :H)
PG9E!%-<+_(L*(61-+JS_<W_JNXFA!\2,)GJTH0 5'DN 5=TN+ZPC3L;R,X8I\LEE
P/_@K%"<)4/1'[HW&0BB9;2-,0D<41OY*83W_ SM$R7)6C>OJ>W836;,FA:$C70+]
P[?'^FI/T)W&2(2##!FC_RB1=TE)A'##I/'& =;[6F,:?=_%:&5&O\B<V4DMOQ6[L
PG7LU+.YVA*Z?XC)?1*S&)(22QPL-J[U=-FSEO**XR';KZ/8\D]VN[3R!LC/+6G))
P\\>6I#P?";(/]M;?8D+%U81TED7JY*B_R5V)(0L4)\2]].AXN 1X'96X3P5\]L=Z
P0ZF-.M2;-QR^,LS_?%CD8;'SO@+83JL!4DSS$$2H+/CX[7.LBD7/(40J-QGS2ZSX
P">SDD0N $)ZP4C?E:Z/-O<*3PNA,A2$^EFFT)@83$*<6FNL;AWO4-]@2Q-/IG &.
P _ZSE7ADJT\.N$<&AH"1K,6CQ>5L,?P&.:2?2";%J;F^6%,2QENB9V7.R"7^.]LS
P:4 RN$RA_TACLRD.Y.+U)F4::AOX*&[#1KG9*6^5=87:JGU//#SH5V)SW3PRLQ[5
PRA6(IF$%5>KBMOKIJI[816VWAH5",_2T0I-?1KP.-:?2$CA172(ZI'C\P9QQ>&HW
P;TU% ^,UM?R!$-Q.=C1*/.1W>CA'FDDI'(8D\#.<:6;N#WHM(B#R&W/B02B&R)WM
PTA'E>1+@DI.H//K4!WJN4Q B+6VXQ"@[(5\@_/[&<:"-_B8.IA;JB%WE.#I@-TO-
P:[G6W)TD\::YWY"R])6TXW0!.1BX0=^2^F6&ZQ."JPT9H0X]XKZH4"&@5+,3M=+0
P0TDAQ*:X_\/YH>/:]3'Y8H72##RD1^-4;N">\RK+54["LW-C_'RY2ZB+N4SNZ![?
P_X]-V3M\6Q.YIA:XXR+*A8*H'_]'3 :3'1"\YCIT$<;?>O?-[6<_*N3"4B[0Y1=T
P03H7$^.DU%B-M&7^[CLCN=DE2#S6:VMT("))-DX&]<U3FI@%,O1/&W-54KN\41%I
PQI6&.ZA<5GL.APH$:I&C.NLZ<%2^X4C>,?0+40^G%#-'&E#Z.?E)64FWT[Z?#CS3
P!R<2V9'$5&[@QRIOD=(?MF4 EV19V4,Z^Z9DVG,E-CE*'B!T:20:,27TZ/S#.XH.
P@7PY6U) [TEL]C5^[VOTQ"4=Y<7>X#7K-AR)O6K_S$;^@#1G'_#4'^LT1F5N!YA?
PS2&0P9R+ W?>3,!%;UBE@R>QD$CX9"Q?G-(-&:&KS6C8^CJVV$JJ51#(*&_FYF!+
P<*"7]>B9S[ZVE2H 9=/4S2>K;=&,;*"G5]31(:$-^.ATXQD:=V:3FO%WI_J =N#,
P5! V[X'.LC^ #BE)(M+4-),#<IEE:.8"QO'-V7RN.\QTJ^._3/U"#"5^F< ]^KJJ
PMS'D' F0;:)0$VE#]UN51/8JK*8=#F($AB4FN@+U\OJ$$/1T@5B@LU(PUMEEL4(T
PXIKUZYS:D15#F?3*.R6^2(H8T'F@CDSEH9<#C$5%E$??YV&D8ZF!07@$MOHDW'4G
P'9>0R50+H<X_C;D#WU%6SE-)/G;E19'D$]<(@WV^*VRYA"CXBGVRPU _=M^X9]HN
PM7XG6!2,@-)'&6F9[RR&Z&/,/FD>E@<3*:L'PV+$T);*^]@/G&B+5]5']N2GM%2>
P]VL/6L:D^S/%*NZ-7HSC1K+4NQ;SHZ"2+"G+O&5'-7QW1NA6)'-F\9!R!<QZ'KC*
PK8;6IEV][)0N](WHCO$0&AY?0C0.:?ZR&>(T\HDRA$E$B--Y!8I4\:!SI>61C">7
P'OB0BZ2P@=IE[I=S;HF(Q]4>RGALM]Q!Z);(37&VOR2;U,58$W]?#P>M'7X+\I*1
P^>V0XB)C#I6YWKX,5)*.*WQ3F7OD89)>9 TJ_PO\BST\N,6U_F:8CQ!T08*BD3^X
PV(38G@"JY%N%^6SW$\TVAZ)[ZRXRD,#$[]2T')* U<-!HL1^8BC<4G:@ 94RN.]*
P!I#%6T6\SFM=6BBO0]<% [12IN-CZYR<TN<$@BD!EXD/DM83";<HR"Z'D,_K&"'-
PTI9C.E]Y+E2G1L'J7Q0B\_2HR+8:9F+-OA71C</.^:.S]#<X],? %BAC8^K%%@?U
P5&[0D:GC14X.+:'?(CFI0FZBJH1$25N3VBT=,R,>T2$3$XQE/?1MA<-UVM.>8FBR
P[5].V%1@4>3HJHZ[0@MEIUBH;;+Q L"TA3P9R?6&E7!AV/0WFLK&7;;_ BRW'B>9
P[XL03<D_XZ8_3/V^XO\I-/7KBX\NK4%40S!^\21^W1$XXLM)17N=IV),;9/KT,T^
PCSQ<&H\\ZS<H\-!*+!Y5QH49W%NL63D_6&LJ:LU=>LT-9#.'[CKZHIU,$-A>!*.%
PK"P=AI1JG*@:$WC"(M.*408AJSZ8PD5L3)M*1_+\8KJAK;;JOOY&!+9&[(@KCK(U
P+N/D@2/!+I@7,@  1*NW3#]ZD6G)C#6"E8;T76\9KW\H/GQ!8]G45C!ZT*^E?.<[
P(EIDOC^*#'"D?A*3ID842,I4(E#ELNS4\Y0]A*ZYN,#"D-E#OHXVX1XPSPBG+N<D
PQS3^1%  _H-S.B J;'[O-JRL+(M4W2@H368>ND;ZRS#9!,KM1_SU!(PMTFHV*V9@
P,YT"&%8<.(ZYAL1-.Q\_[/8NCPOZ?G/+$U V."DP_.@_,IQ;C#610./(*2OHH!J9
PS?>%#PY^D43-T-Z>ZR"3JRM%0T+YX<.UGUL*C6*T=_=:X-"L0&L Y+^\P,_.-@L_
PB;,<W5/;!B<U::-;3V='&Q)A/P(.;>2_SOY4>Q?MNZ?7CN#Z(X)A:6"!0@LK0R)7
P.(PV4(3J46=2EZ((VLA0M6L21SV:F1X\^"J&SBR?%B?_GG#E.3%NWDQ_D"N&-?TI
P4+O,P*1Z)!<E0E6V$1X%:TJJR_'..>$S;K/[GOO>J(UQ*>[UAU&OQN5J^GO6-JB(
PBOP:Z:1ASX_E%9$]VB^[ #((0&DR\Z2DP/:$6V,M$AC[/.+OJ$^ P+JFW\[VB+QZ
PU)"3)<,R35PM^HQ"K"6#JV(- /]C\R[A&H^#=#9QX'/U0[<Z!+5O1/OSQ%LNY#E+
PWOQ,=:ACNG".G9@&_@LZ[Q>30;_:?'9;4@M;#6WW$4JBN7@.6*7[P+?H]T4!>(OW
PGR]^Z;431_2"VN12\=WN1_J97+'WR T&"P=X/\S=C@\+K=_&9@"J;P7]Y7L6\V*"
PV/HT,#^@((D5XG3_P8 )U:UUG.=D+?=GK3:T1K,,J<P]G <@EX8P[?+8OXBF*;PL
P,OR647Y^K;Z7*Z'P-X[7"A@EC&*\!Z;PZW(P%$LVV?D=-.:TA>-9R*^GM@B?\R@,
PP?=GI VE!MEY_%_N6TA, [J+V=RRHGC"=94D 5:Y+,^%Y4\44;$_N7[WG(=FD9W8
P4]*$N4W(:5IA.'+IUSTD,!P:O><+("&DX'D* 6A=G18P1NK:??RMR/ZTS<$62<?$
PH%M^*^Q?%;OWP1)LCXM]TCE,6]$XFZ4+>O,WY4UT7=5(@(@*G/P )8?WW("+-;1P
P>=*JGSDTX*.C[:;6^C"DDY&\X,"U19/O>YTE[WGU_3W$06) 3D5$@B.T$%?J';-G
P91[CTK1E+S/X=[V EK#$HAQ$+J.Z(Z6NFU5W"_"<0-Q+8VD-70H*G,1(#^\CXG'3
P%OU!!1U!\<:"JLU[>29O7]+A*QO+4\CE'%'.FGCUTV7R"3>1 N^UUB,)>_-^X,+N
PYAI?"),L6$0US5Z_I$R=__&4L*'I.:&WG6&S)SA^TS)RJ1S:)D</TT,C^VI9!\B 
PT6[(0$[0%WW]HK%RW/2VE]I#G]5S-I=Y1(51$]2:;OJP\M.ZJ%=H%/W6#QKEKJJ 
P6MY;6 Z:]L,GV<S7>^MY7NP!<IH0_ MA4:0E'7Y(D5,7#3D/M%<#+9U,[/CS/.3/
P/MM7,6]&VF)->YF8$C*7'WTQ[Q%FJ1[02?6YTHZ'U6K6-U/;E3[;)+VB)DU!18$9
PE%[&5T);$4 WNRY(NXLJ-#8TS'\$W)6NB>:?-+\&=I6P'A--P##BK\) U]S4)X@5
PEORFTR/I">%:$5J*HS%"T.\"ZQ<$';H0@IJ%M!NF!UMX/]D[N%W%@K!(OXMP2C3B
P#2-SD$F#E]&9ZLW$G*;:L[XD,GAL^YM#5"(RE]GB0[+6)*> LL$+0P'\BJDT]FG4
P9;J05$L&-?C4;&EXLBOZ-\L%OP.DG'G$KD_V.^PLSWS6G@QCD^?K]!!%N_4X).W:
P_DD[43!I]V?4'@.?[#*+B#0OD4RLK[&-M&[%F9&4&8OSN)SRDR;P^>IPN&);(\$;
P.2Z,3'%$->/9 -<@7H0T%J+OI7RHP['$]XPZ>]B!>?<7C_/!25XUR$M7 (\8M* T
P(-B]4!\7#'[Y?U:EX%PC1/-DE)<!)Y+^S ;GV;8K"-.[4ZF2[WR9_2^@P27=V1P9
P]VO,R#E.L/TA]+X.:5_,]JSZ QBNF3%:I*OO(+M1':3ZEH#N$(;2E96]T<ZO;;:X
P\SUP=&^P"H&"-)&AIR7*24RZ#TEX:&BW@JUX(AWR(V162NH$<I5+; %;F\.(YVR;
P=FC:&K'AV\W?7K?3)%B?*7M&Q8PE4I8:WE;@Q>7:0D2U6>=3 +>E)LH&S>#Y'ZTC
P[Q$2D#6 VK(P7R9I^>8)F<>,X[/$Y6>_^DY?2'L;6R?O<A\;WFEB6@-,U,T-3(G8
P5_;SP0A 2B:X3:_^@*9LOTL6Y<NZ3FYHRV\;LY8+3P63W<Z;Z"*R;BH_ZE5ZSZ-.
PCJ-&PC4/6*PQV)09-CH>,M\@#PL)8F+3\M<UW,Z/K@@I_1!L#$[$*G<FZ8:#);0A
PI(#876@CX+M<1.E0"X50XXZK4[$FB3NE#TX-U?T_<?Y/3P2 Z<C^=T/J<DVS#8_@
P X@?=C+KQT2_KD33D!""W<SFUZ:"%X)(?/'G#7JA[#*+4G4+6DS;" D5][V8#6>Y
P1_=!A'!VGWC (9@,_U57FQOM)X^AMXE3@"53 QBQG64VEI?UP;X,_T).&E8EKEZ%
P+3-.N%E2EG(7P4[;VLHYLZ^>U)$O<CLVU[;8W,9I:B3/4?AD@!&28V*A\O2 #*Y?
P2<(:;D5E..<I.J9=QNJJ\#2%_?*WESVLJ:R5U8OE(]&0U9"++57/4&CGM"JK (R"
P.%FP:WO.J*$*W)O';V=U6_CSJ,(D&JJJ?)F,5= %?_L4OE5S@.IJBR-9&W[>5V(B
PWC]\!B(^-A  @##Z%.?)JE=EUK.$NRI&BY?.X'G2^!F'E,UZLV;>S5-$)&F_WU$/
PC< ;WUSI@A!TW;Q^96&)GDTHKF\.^=3G;G8A)N"7"3E[-K;S".NVO"2;=7MRZTPK
P7B^FJ51M$'I43C Z#=KK. [/_MU]Z WK1_*O(*9&HS,9QR,W+=X70UL >(HH-67@
P5. 4(<PS)S2JFNE4IJ2[B00M,(0!^"+QZ&#]*<G?:?SD]5="^2$3<_Q@V'\F??\5
P3DXH8TY_D%J'+87G6I[:JM;H6XSB8*L9)8$$2/TLHQ+'N5G="D!(L*H23M&TXLRE
P7V.;<C!!R_14H=VY+7B&F:CU\\Q@UIY'5JV*DU$U0>1>F1!EHKE8@+XCM?VAK,'V
PNU1=^I%Y7=Z3G+2%9W3*BUY_IS?,FS "I,%R>>9"QOK;05-7B.^*+>"L>X*-C+;0
P0RK5WB5_OTRIO2<9D@J]?T9T9IW""%.#?MTHL9V1HA903GUS/;!"(4YXZPY(]9\,
P$1W!Y</,+%W*QG(\,HCPF$B3T\J.>=]D@XS23?&60T3(<@0/8%,&_]J5(WLY\Z_H
P9J\*+Y1U69Z2.12"S>BEEG,_T,HWY%:I0M\NZDTRE**(,$WG=]&RY;>5<X.@R,!X
P8@;8368>_T@$U%'9%9:<G'@&*%$NCX4-078L[7FV1L8-E8:W0+4QP;.O0>4$I:Q!
P154G]U@H-^GSR(Y*G7S!Y6<*[WIVO%OO66JIHVU06-I2@.4*ABN)CNO0'^0]G^IX
P"1HH2;R\6N  8_4MRD["Q]4GNP(1M]*#%-)ZNE PR2(/]/8C)5 K8U2 B4J55ZL)
PBHW=6QZ72/]?")H;B833@<D@+[S7M[K.RN=4S-2+I=GT/$R,GGNQAKS)FDA2+,F:
P+6,JT-X2NGK/E3IK96!V-4&F:* ,!#T4)].41^5<EO&-,X:\P4DFOON3\ID?/-8B
PQ0T)U4^I3F\YD,C//J*S94P!VL2(ZA5MO*E($WHG6/8E Y2B$3=Y^6@!'])*2WE]
PN$P;QF*1M[/QK(R@OWK+3K&6X_N*6Z\.7$K=&'L$G&EA_%9P\ZO:BUTG/<)G(A;<
PA@NY;R9_ 3'3:$?+NP *B/6LJ5N^,UD/*K52-9"2%K],M:[Y;!?T6B#TONETE<<,
PY+T$&7%8%A#%#,;WDWZALABMH>D2!V;X^![[CFMP%,C<@$L!+,WN;)@CLX)F3>J;
PZ_*OZ\$BX;F=;QSE!H9<+=DY5_KO24G8ZA9X\();ME3EKB5QZ)OPB2/Z 0-&?]J+
P1+BF%@\MI^,#.[PI)QJ+^/Q,20_,P;5D ]O\$;9E0G):D9 +V3[&LU=>>2D1HY.C
P]@6,\]'?07Q/#%:9W5&RTA^F]HK)T)[ 0-#8NO$'HCD&=[$%5_C!]NPV>.VVA8X'
P53,+?3H3(6S1[!$[H/I!&-;&)A6J7<;IB2EL>R>_3U<"S2ZWYE4*8Z'AD!IDKVH.
PN"%/COU*)J3QHIDI2%%/85A<IP(35$,W$%?^Q4PWC=6WX>D6#F<*2X7H +;7ZCBK
P.:[_#8J7T@00;K^\?'R$.VAALVVOGB)-&:031G!L@7+ O,VC#HHA?%)<9_<IXZ*7
P-'R<?L1DH3<-LN9J ZY#>9 QV!,'01\+=-A)\@//S!#*/0/TRYD<TX 3+>,N"S@@
PS<7KY1*[F\%_'NZE.X5#.*9FY*?G)O:PRC.IN_M#>)KQVHLK1761G*0\#<KW--F+
P5O*R?O=JU28(?8D<NRZ0 =D,Y_ ]N]SQ*+;M:MS*^?IFZ[S0,D<7O!\B'DYOD,Y#
P$9@NEZ"W[O4H9,]KZH3X!<,Y+2)B7U4"?BN+':DKO=6B. J+J(]Z7) V9QMC4[JE
P\<AJ#L5!Y5HY#EL6V'P*AV_%M>]L!6[/A.P6@?9Y'6KNTFWG0DP<#M??B]HK] #_
PBK[ILG>%)S;=]H#R'_Y/%,=M1N7']V#QFZG+OZ ^/".TQB)#MO,NI!_GNJPE]M>>
P+#1#_<6E)<4QQ+,N@OOYT;E>46.BY:,2(\F>E/79SG'3(&LAS.L6Y[O[*_S9PW$L
PO#!B1 X40+CUR)AE.Z,V>Z3W)BS()"7C>)FV7#FB4Q$-%J<<1%0>&*^P(!5V# G9
P(;%U9M\:_]7W8S7GN@4+.P/U"WP"ZA%35")_PE,,G=T'O;:ZF5268+M3VUW^4%!]
P^H-PMU8_;V2$X9<FLBO6K;0);BM/6U'OQ2KV;?://G;2UZY2*_;> 4A>,CZ1R]"V
PY?Q%D^>T?QHYV:CBB9IQ7%:R\.4%[W/<DQS]^IL-?/^[_;7QHL$*")!G'FU2<2NX
P68QO_HLR>=CP:]PBAX$&CEZX$FV:22-BK)W;7DOW'Q!'@WF7,+>/$<PM4+@:FF@?
P+NR]1X,'+68I4<HZ(FX\#U_YP HHA&X1M2 O;%UAD_ANI59F3OOJXZLX!@:,1&GV
P@==I,C(FO7AIO% Z;47]SV%< JY%8!8^OZT9V@V+D&#V1])E?FL6(U/?5AET'F;%
P5U+X^%Q4NQT1 YD)[5UG'=FAV0H-?M5NMWNQ->J7R3QM:UC& @I/-#Y4V4F7TZJA
P&M:( ?!5@=*@ GRR6K6*B6F9@/8R$94ZU:."?G0.X",%F$X()K_RLG5L5-$P9N3'
P8-9-Y,\!>A0_44C6ZDGD(TB.)B5=PB8(<2E_7,U[Q1> E+)Y]4L[&PJ2^#M5 <[&
PFNV<;EN@^I<1=S!IROU.%(<.$+">'_05W$E13M'%WUI?4Y([>@.D'E-3$R:EQ ^M
P34G6'AH?M7!QR><>UJ[3_T)')X'>/SX;%[*AVD]%7?IS B PSN96H!)NXY]+(: ?
P'38<R?(]P3ZV D[7+*H($\*ON#(LH\.Q/$-(I"MY?^455RLY=OU=T"0)2YJWD.+U
PF\SX*-\B!F!<M?1-';5?MKBZ<KT@T2;?^G#M&_$IIW5V9),FNE6NO1O:-L+0L8:U
P(8^Y!O>S(SJU*$1&Y<L>5M5%U\Y![+[WNPYGIDD9':[J."HN+YRHER/Q&C _0IAK
PA++BZ%3OUE(#J[EU6\;91SY^_OJ1C=3^0^6'_+;"B% 8J=8.[R_7?7)+T+$ H)E3
PU?(*_.(OK1ZL_0B$A@G,>C7QTYN.%S'CT 6'-2L09Y1C4UP;I>Z9]I]: KA=#RLS
P+,:# RFY7@YB7.$G<4JE_AO C%?_7] /^8[Q0#%>W=! M&,3'#_>D0_.Q$> 3>DU
PO'ZZCCEK7N%D]18&O[FA$K JG63%JZ>^VD*/J]P%VT)+.T=Q%LE7Z^G,HJ5D8=B>
PVB P958*"8)"U9N=U?!)66U*1(6,!6!)G%YOR9*ES%0F@2$_FR;MD&D5L,5#-[ZO
P<Z1_"7/ 3P0B2*$-)6@9CK"N^%2OZRCY2'I!X.L_YF+#4_T\<"&7]5Z+\NE\-$$R
PU\=3" ^#HIX95<WQX)+@9/&AU/.Q3;=EX5K?*KRDOHK#M([;9@$R1#?7T$@ ^9AY
P,Z(1ZC&M<G(==8Q[O\V+MAH9ZWFX=:H6_\_.GM,2ZSDQ2 <[3%MOD,\I6$\T7V<=
P3 \DJ!P<ZU]T XKY\.R W[X%)2I\/3A0?/8JQ&(E$C[@!.-K? JF-9W'X1B$;N'A
P-J#:9V1)PA [,(K%&'I'I5J8E]#D27>AV2GR$2^*PQII=1)&8'^%^*2?44-'!PNA
PV#1)3.*3 )JM"X\,Q IX(AE/Y-Q?;2_Q*(98_.$[U&G?I8FE]8Q2H5X(N\^F@3.Y
PK1H<EXV_+C]JU4*]G,']Y4*#M4PH$CC=KT;48*/W_6&)95*MS21"RYTWUUG*\RTX
P%=2!6=UY;P!MI7F4V=ITM/)B&?\C=C:-J<BIX.X,0MAXVP6%,O&@DXNA@NK+2N.+
P!/,L%?,+-UH!)("!OJ90BTL)#H/D@*'SD6ZN/*R3!LT$10R#FR,,@0PX5D,)Y-W8
P>*&]$RD[M>3.BT]:^D<R]1-N,-01+622&&'8RINB[:I)Z ] I2KW#'KO+EOHF6+R
PP&]ZK_165EF7N!J3^>R:(BOBB?*1^&9/"#2C%HG:?_UBD,3HGNQ$\&L@0N.\EI3!
PO\O9@@PR4E'. FATD.TJ+%\MCC1)16EN=HV;K^?N"SY:VFJ6FS_LR>A2%,<A@N(#
P^16S.4I+%Z(7(06T/'2^8,A?Y8HYPX%"X98!<K[(!:E\6#*^N 06JWG9?4!I;-ID
P1>E7,3@U7 )A=5K'IF/U%*6H*PSAS"_FTJ;O0A,T!ZPJFO7'(]MZ*)+Q6U^GL13'
P:JZ7SYFW_#:BQ\)%,KI@E7\2_*\2X!2L&U&?>=(1A/1Z\D.[LW@?=#KA4)6^/ZHZ
PU7%G3H?5F!=5)^TM%Z+E&SP/C3N,969<.;NJ"C[F6)P%MSQA7]N $N=%R.^4H_#O
P=:EL)NI^.AA9<&2HW2MNH,!034ISHK0=!.WJTM$X^6A;<B6I:W%I/G96"BV:JXH%
P\5._P70ZW)^X26G1\C>6D0#U 42#M:[[Q <H@<C#AAF9OCYNLXOD2[P+QP_F&@:X
P(J\18/4BZ\R==^/\8\/B-(P!__.A+#BR_/6F! XF8M:YE-W,V@2+>.0OO%[*<?-E
P[![*[, GL_/,D6(S(0+3\\$'3V"A1^1/LU/4S)%+4: 8B_%X>5Z0Z[ZG\8 3X2NK
P/U-7<XU1B;9P17+&A7-K5+#@O$7*4Z++6[&!3M8X9R-H3 :!LPQ5,?SA&?BH8,0*
P_78I.JR(RY#L9;]4[AV<A2$U=*&L/TD0IVPY^^U#M#HW!*SSGAE%;BMN$"Y>Q,^6
PW/K'U<:2F%1R@;*@04Z7]'%OM5*^"(5*1\P2X6E<@-Y?(/9,\4KUA$N]B/'(7LF'
P6T&![V,IKZEY" VM[.JJS[UZM^B3%BVAS/;="J AEQ2ACU#._%H<#5X!2'X53=CT
PDO^@Q3L/.A(1&VZ2V)HU6NQ3A1,.S#]#SEH/%TRHR$+=#>*2GM@(*>R+R94NK/#X
P&@VE(2]:M:P(-KHW@G,G^F1PS[R1=5'6+*]+7W63G7K_A#>:Q)7.0Q8Y+%L35\JR
PL=ZPB1%]#FI<K5Y?E-<#<>4HA"&_XN<L3,M5*52-;M'K,5PS!;F\#+A&;\%)PJSK
P*8Z58AZV;#TO9IJ3&)<>U!!8F+/C&TB^<?!H$MI,D..9G]IEJPZM+[A%1$9VBF;[
PGIR)&;X'CGF;*G.P(K<A-K(W+_1 -@GV,-T1F(^_ZB\'07KM9R)S<?2'?6$K?PNC
P35-:X%RBNTXGO$LB* AM.U**012?='2$K8;()[PY!R@NZCWY"/,IW@^*;R/3K86\
P1.H.%7(HRPREM1UI=[URK&C*'IB<6T<]C8]?.,.F"[J)BHY)0D2:AN_.40)QC'0%
P/VYU9<$7_EX@U[T.^) L7XM-EX]B?U[2&D,9)1C K/^D"198XG-UT@WGS,U]8JU^
P[CP KHF>#Z?,E#++?T?U3.[[$MXH"WJ<SQ'[I_P(-/QC=)H!=AOTQ$ &0UZ_6-.,
P^2="TX:_TDMO] $UQ_S9E^<F:9^QFX7R7XV1M" IQ&V+P_RE33LUOS]$Y,TTXI#P
P1]5'\;=91"C&2F&5I-=D/[W7I)MC[N$D?DKSA%8%@RF1<=:8;N:"@@?-FC.69.,;
PMVKV4+L,.%5$((Z%,-5Z<OZG5\5 T63C3Y?A!VT^@<;("U7I=4[OEMX_TR+IUC&P
P^!'/ 1([9U^%-_MJ/F4>D56V%KAZG'->T7,<Q[:<A\K&56208[K6HE>C13)T$-"9
P8W/G8WF?_.?14G:2)0F2N8EA>%'CD85*A;*LI:_RA[-E5^VF,_2TIU8#PM_X?.)[
P6V#DM+N1DU&*%5="-$8,^(<KHJ]/=?EOXI(/$>4P9AV<VN#3!H:$V3=IN[B>*_7;
PH-6 9V%VW(I"AT9PA=2FZ:>?.N7W\F!5&N3[[N9L[99ZE)FZ+KD=7V;=U55LZP4T
P?TY^IQD93@Z)10O?CYI%A49,BB5E(%B2?WKA,8C=35M&@*O[WE-23I&O6=]8U',O
PF8C*T:]O#!XRK&$>,N%6&%,N1"]]RN'EG.*\"G^8-JB/A.:0QP/BYMT/'^V85.T'
P2W<;A)SO6(G)D.5CWEX[WFX>7CR@XT]71[I2L<=/E?>7Z@<C63*T\3:(NNS=,I9*
PE"%XZO>Q6C2!$!?29&0C0GUP_2@OB'EKE!)E3FCU5:Q_\*XA2=BWY=QKAO!4VA9T
P@UW& I5U#)_MBSE"F&CZ4&WS.LMP>1WREP"+!/=5E$(ZI?6'K0BUZ."ZR1-9\X$L
P\DH-&\G4<CH8;4]$KNB?A0YYT6SR'H ,F2\\[S=@)W04YT+%Q6,@P8:)+)(M$_=Z
PN<!0>V2@FED^E5:76!O(;,[\^U;DZ/H>'1"^*.!-39USS\Y'UG"VTUC%R0EL&EPM
PD);T5:,[2&4I;$"-9=5'T9Y*P9>V',KU]N\B"]^KG):7#A"\PYT;W?4IB#I7DHZW
P\B+]7^="JXO]^HC=B3Z**>"/%ZZ2MT>*?#VD=X52G:/Q%P4V7!-1LE2?K5]=D=NN
P_K_JP\N'R)646!/@#R*[&T_ 3UPPOR)M0MOP=9#?1?]RYY(A"QG[L0@NC$FW,@JC
P+E<(;R:?5D<:TDS2+EC1^:S'#9ORYI;B-QCQNQZ0D  \2\W?9A0:2:&60U_R>;DQ
P3@1[-Y-DN!),H\9%(8:(OA;_R!#0J01?:G6&G6XDIPP7:EPZG+'.NBX'%MP\94CZ
P O%QL3<I^S:GM>#IIM^>F%7;($@QB?H-3N"T/E$8W/Z8SC*RW1U+U0^K1,A#0+.>
P$Z#LP'=7!M#PI/48!Y3VPVD8FFX6JBJ)/A3=?J?TR'_.+5Q$LM?XN6ZDNR65ROWO
P[]/H3< 3XQ^/I!'\< 8#1O\#B"CJF!2D4#</Y_'K]UI.(J"C!L8]THAI/TQ\@/LR
PN,L_1L9>[SS<RQD%:.\7O*2]HY9I?$ SM3 :8HGR4%[*?S^-4UE87\8XQD5P;*H_
PWG. ^D)SYZ4J=/B;D7/G5/HV>F["*QD&J$ZHWU*B!P3]B/>,P],WL6Y<"D(.TX['
P12X6"\VIUHNT0I;[?\<"40IM0.7?]:+@BR#*/-D9+N>W>7G_P(CEL48 &!=A/(.E
P%50F^WKKE+?E<*G W V@KFY@"KB]@EJ?\$OF/R^U%"H<ZE2;C.Z+[*AD?F:G=&KQ
P85"O2NSXABMXAB9/"0XBDI\C<=G:Z11A3E=:WZGQ!M2FP<]0-*9W39GWT9SL8_=-
PAF!OXTO)D' X?O-* 'YAR3A><[N54!"K<M5=O4FR;&3R.H1.36_32J,48[P::0^)
PNV[>6T/'W%&'=; Q;.X@4C'BC#EQQB:5]H:(QHFVKOX&K,$]B^+N++O?09GR=*XY
P",]GGE+VWR9<Z#?*0M<F)EW^4VF"//?R&1485H%QHP(2[1W0WUH+CQ?\'J/%>[]U
P2&A]>:=$Y:O*O?8$?LBY)GU7B!2*E,QL;)8N&H.[GPD(BP;=/R&]P='&U( H:B\!
P;%N:>.6@:M U\A.'2 +8.4B_,"+[79?&L'V"O  +#[UA_]_V!!*UN&7G]:%Q:M>-
P\!T@2JV@&BT:ID(')Q_&:B5L4W*=):\9#!$T^ T!-\!K^=?05=DPS;?^+%&T<E6\
PO&:<3UOXSH'EWY@.#V^$2*.X3C>L[+-+XWDR>>NE1L?@=OE<\%U;V6/K@_W6<^R&
P&E$0AW6]DQ,45^L$T?6ZXYA679P7BIY_CHZ/CX4I:-9QRE^GRZS]0[PCK=;MR"DP
P0444]DB8K=J)4"N 5DN4*X_]/#*#HG](T=:H-^;:KKKKG*P]_"'ZOMZ3" 4.VJL3
P^5"<]*./VD23O!VX5+T!,1,K !+SLB=?9HPHIR[(>W5<&8Q+PGY[]@67]D,+5@+E
PI8D[++)\D->2"))6NZD@2 MLF?7?+2G"#NXS$WH!+;NUOIS_6BXX[,YTZ2 B GZ7
P=7Z[>S_;% 9#^V7]75W)8J>TR#V$[>%5K4H$R*O\Z[/U^192+"U&;W;,WNXT%*+B
PFT=XTS2M0A,.$SWI-]FY5 GXS;*1!J=F8CMI46U8'?YCV0P_R0SETGAI\%<V!EKB
PB>_1%79^/#&_HVU[.PRKYNR)GR<5LGY]Q#V)2/ 8--3AP_J9["#=7Z6?;O*;3:\L
P4#.<KZ1>]4#361*QMSHZ)>7=C,-MP4S^O%VZM-%&_LE#Q**"J3&S$:18="33M[A!
P*?BWG;R+K*$T0.?_[K6WE&#P6YR.R*Q3=KP5^8[NQZBM<%X,;I@<.IU'W:RX[H?5
PZV$"L,*'TK^PO=GL<)RE/J[KR!L$SC#(-3.X[NJW4\:'Q#B<R^W+&C'&"K$SL?F<
PS[IL+XJJ#9U=B[))<RNYJ\@W YUE2)I,;'&/^/1&3(*]T'S>L644;I8_*+<$77PG
P.E1FL+2-X?O1TQ'E.D1/17%T65U=LMG.Z#$E9"^5\XB6!S]E[T@L4N^J6^F$DUWW
P%S:WM@6M9WG=/:".B)TAGH*79F'&WUD;^?C90&I&K-HSIHCX4H+X<=+SUOS\U/*(
P@PRXU_JC#M6?()#8^3X-%0A9X&%T0"B0IH:ZU2X=/]H3W44/%Z#J$F-G!4QBA:"#
P+F,F9J_9QLCJ*L51I*A?+!@0JG@GPL=+ZI<743*/7Z&N%*DCM='(ZO#+E0B6L@('
PS"P+,D*ED&M38O:@!E3!KC1XC\!VK^H)'$&'<&B6+?[2@*(OII5G(;Z=Z[;\'/1T
P?1P@^YA,U!0$DWC0]IA\%M>8@J<00-[>6>-$8QNGTLRI9^DD_NKOPG%+R3!HT9H8
PM\?K?6H02]-$">LIF#/245O,\?G(G0]"O,%Z8BOIW,<'_GOP2!'VIO>5!@-ZS_L:
P\R74BCQ7;$L7%@UZ<++G+!>DZDNXZ2"HJKLF;$FRUGPB<' -F^L2-]2*Z]C>'JET
PW;__ZFEQXU4G@P:KE9P>,+YG;?CUGC,O#D%A3VY> (?,Z\>M1RD:6Y^C7.F D'_W
PV/'0@D].7R =!)S^#6HCT:[*-9%![,[BB"4X68 ]72IU5N6J/VY<VK!@:@(UU=.(
PD?#^SJ-,#YJ/&WZKOYLAQ/V<%O<5Y%H<-@J'*"99_ I=89V1I.071UV"U$PO2>"W
PDM5_ 5#\_QTV!@>,KM)TQ-N:T/9Y:;'_XZQ5,U/17B%_H9,V:KKE;[?E$-'<*VK]
P^IS'W2KIRIG!?$IBB_[:?S!'L7AY%J2+%.\A%'ZEC>:=K\V93#6XW-@].XD3\97_
P47A"NROASC@(0N_$+-+S,%XS\TI/+BK2?H53%EQ1U,F=PGAB7PO587TU$=BZA Y>
P-M!Z.@QM+F8U=)59 ZXU4Z#GK6I22 1%-Q+_U5-;9,OW<7D85KZ)7-7HFV,OOC;0
P'5AG[S1M6.& D'ZS*=7C^(\Z\4N$7 KU,<Q.3I#Y$L6I!#!&9G2ECOKMHL0)OT^:
P/E< ?!(&C91HP%!^9*P"] +5+Y*]&;0M,R=-2;U]]8&%C]Z![4/8F]CJ]8H3NC)M
PN7W&1-MD"E#>W22PZ3^:8R!RA[E?E.E0##*D-+Z+@_)"=$3=,!Q[\+%O3+=X(]AM
P"N(=6&WQ>^_ [G+AS-!2T--=!>VU O-ET3\+*?AX>./9HHKZTZ&\%)B< )C20OL]
PNT. '3 IE3<WJV"8UQ>!/W*.LCO 4-5BW_IL[WX)"A:@NNY,FAA#7 W)_)C569!B
P?M0'T#Y)*Q*X5PU?@H4D@I5ZTK@.*RGQBG-X]B&&:9?X6*Q3"\LEZP$Z'I4RY2K%
P&T5SM"I)!!6II)X5]:)O.%FO>12RCS[KU1@'"W.;+D)_P=#3_[G*XNCOMFV^+KN)
P)[26M5^ >RG,#;13$>-:S]J]TJJC>QW*.R0A*%MZDYB<(C !P*AQ?C\Y-KH,+&<N
P[/U!W_BS&;ZJ[_R0H(6:M>=XH'DDKF[2E\ EJ$P4Q* 1)YAQY8FV]GBA=MTON4G5
P JRATA  ^F"5BJJZ2'IJ[MR%@H85FYCK:W"D.2V8XOGI#L1CBB98LU\?O8-XJB2A
PH3(71H\'EZ'XNW-Z;-4X8PWQ5Y3'XD3]::_(#,'BN[!WZ*#YBE43G](QZCL>>-#[
PC[<*P&P7COQ5Z6.Q:TY2Q&P0@7?IE,P4C%(@;*=MRQRMZ4,+ /!O>R;@.[N)X,H!
P;@0MO4EN8[#@- =;+J53=*P::]['UN.5$&BT 8'';63_N=R%V!%%%VM<5^4K"WWY
P.,.BT -@3^21Y[;-E?/-3_)TUY@A'0/E[C3R=SF[%"^=68L=]@@>B. 8JYJ-RB9V
P!=3^R?>J3(@EH\*RB,L?# Q^DJ(W\?8FG%K<>#X*_*]]-;K<T37^=<--'V:,M_28
P93#F!<>%/$> V<YPU-$O[5[XQ82<\*44@<&S?(P!=JI30,VN?)1N5P8 YOQ>7;6U
P@)I=Q@A=BIH3X-"6>U+5*C38Z+^S6^[GNF>&Z&B>4BF/M/T#6I-!K<K(FM!38:TO
PXOX80=1\ E6O%NX5YBDHTSW&YVW? 5A)'9&(K)Q0^$W8"9[05)*A6CZ++*"W)]4%
P*=AG*AN8LCX%(N_1S^VF>47(V%I12F=(53  *ETK*W<+DT>!V-Q#"C>'S#L$4=O)
P!1"D/A4]1\I0@37\ K/YT]Y#_>6N].V.0:YX@Q!U41F#0%\9#&],ARU "^ Q,CSP
P&RIL42RG7K NHTU=^WI'7((WP'W93;F7)43BQ955M9PRN^#V7,Q@L'M1Q!Q XTPU
P3/]=XF\&RH;2YC6"]0.S]MV.Q<&HP48VGS!*T"P5F2*WLOLC[I#'P'![1N_J?$T/
P-/&*ZY2,4=RD7[4_&YPH(FHQ9U1$48WD]E\U$Z&)9+.A:,61?.#><WX^;%O/1(0*
PDB/R\D1(SX.O)+9!<'RNT 1&\)?-+_+9+.N2>,99L+58ZBY_ANF9*<CPI^GY*H1[
PS;8D>EZ.VAG,582"XGOI%\$$)Z.$K-J%[!XJZYH$>]&;J#%XVB-3V1!,^P\QG@'S
PWA<2:MW_O#3II"X&#1E:PW]9;A;.">O3W"L+*NMS]I?'N>B +?_$O17"B2;.05FU
P_7P%6ZPVPO93N'6XW@K5:8NL.YF!<U&&.JO8@M4;6NXSMY& G&>BO>;Y:2)>&]&'
P#_G\WH"@+@Y.%R@_B$P9,QCQ^-\)5O/ ;FM2>@6C#T!XQHULN"<_QM_R77RSY*'S
PWO,RGW(AT!%8U;SJ7X&\RE$HKT:72;*GD'C88&.L>,+'9P%H,JPCT?:Z)@?Q,?PZ
PC*#N]TJ0E[9B:>[ 22C+!N[HW60_]<G$&2S?%?JO8#&41=(MXG2T<ZT-G#%0 ,<?
P9B];%G3&S=DOJ5NF<CBMZ1%&%F:F3YGO_--:\.<V(**QSPPM2,]$9V,U*K/&>*0F
P*[H;^DUM]4L67 PDHHPGGHX,9[L6E9T6 XQ&WE'UGX/$_+*"#6;\X<A8W;;0G.63
P<Y__AUN3L'9S?3>',T67DZK/5O6T7(2P*A0,TX0"J/E)V)"H.'?Q9=3MAI;2DNQ,
P]=7=\BR7X&WO'Z:5H!&(YQ'.2<^(M]HU#!4 H]CQEBU K2!2<Y8)UQV8[54 YFA@
PO6")F!M$'D>UWS5]B4Q[#?+QZ&6&'+\KP,:+.Z YN9A4[0]HW5E\!;JT5 XB^ISM
P!EWON^$'OVF$==N$,XW< N2>)Q<ZW:%'&;87$'K1#6GG%GF3DFFZ?\W%_V*]-VDX
PK8T51F^XOPB_EC0P?V1IQOQG05IB"M#$D!I(TA\9^[GZU+/?^F)G-*"'.$T*M+E[
PN;KEC8J;8+Y_L VQ9%V#H'(T)=U.U@+A07?,RL& QZ&<M'/55E)UU6A#+Q!(F25R
P>XNNTIT!$O$^YHK0K&I=GU#!F?T$MQMR9\)T!!U70LM<#O97WC(9CJ80GO?'CDQ>
P1KXGV<S9P@XH3 $@:83JHHT6>,&MQS2(3(R!H![Q8^((:S:DOD^%)>N>]QE)B)5;
P=(J2S,'7?K5)37NF290!))!MDG[EFOD.#JFU17IIG6L]PEH"=UCWZJ#@O4^#"9B2
P1D6]V="H,#K73J;:HVZ?-T3$>U4-M'1/![*K6Q&H.:JP[Y[O!)229]]YA$L8FW6Q
PAP+ 8*U7$Y'(HTO2R;G_S'ZY/P5(2:,B//2[95E"6IBVH_R2=G&HG[[B'=M]_00,
P1L%]=,*/BSO-[%1U%DI7.-/[GA9%?=IP/S\4N^0:OFD1 AX6"N??X482.H=',BKC
PPJHAP(3YP8AIHZD@32MAH<E>4CE.,X+BFW4CR:8&"">#8*Z(H&J_P9M?;,,N7/++
P%%AJ!DIP(3O#',$LG<T5T?*F_-&H](O/3K>^9@=NJ4T6<5?3%]2+K#S-6/M?4#CQ
PN]L7<L Q1&VN<2^PG*+D0Q7U#UBUJFF!O\/.<?;[B/SH"YCJ2=$:>NXCPDK$Z83B
PJ$5+G^=<;C(ZC@)[G<DTEK^7+U<4#;BW$0VK9^@]V##NW81:6 @,TWO0ED%-\LK 
PKN="\OVGKZ[I]J3I[E@<+P-<5_N MSSR(>N,E+Z4A7/E<"M-AG31N^_)F+<IIXFL
PXCPJ,B 6M*%*#*)K1T;YK#'@J?CP;!U#_\3R>V;2 ]A?O_CLR)^E+Y[0?5E/]Q_O
PWW"_PU_BTS_O3'M9)8 G%5+63+H4P#A.2*FNCHPVM111/VNE"9+96G71O]Y3)7U7
P0<7&^^5-!O$]7&W0E%-*/W;!ZYP'K?#_@APUEC6CU#13MCU:+SJ<()&;.,P3O*U;
PW'%@@<'78IL8!;06_@*_E":LLZC14=!'MWEM[\^5DNO?1\GR:UAJ]ZG?W3:Z,G&_
P%FJ'_[5MKX.[ *(7VU0V0P+(VRH+3SPP3UD#KT$NE8X05KC=:-?.$A8^_@81OJ:H
PO40"M,QL54?##6*1\]=;YT>*[BP59Z<E=7E1_RHMS?2I=+>CK<2?$-M04:\W>[FM
PPC'5#.IV?G#[^WWCQ$I=AZL816XN&Q[@,R*,&Q(CD22LD?O3-IM?#$"20.8Z$W\[
PWHF.N+L9F7')S*#K.G=RJPBG_C-2$@#^$PDJ[#;/$UU3-;T6X>R(L'VK-XXU]C>)
PM)#QYU"T7GT(@9U "2$MX7']V<I0K!BUANC*P<0A@'.7X'A1BPN-S%&>IX:R,N?%
P?O_(AT19'T0-:6/<M[Y'%9)#I@VVJ:R*@1L/T$8+J2%4D0WE9^1KA>H#%V%#&MQX
P=W67U[G].?4_Y>W3,Q2)2&^OX"H(1TUB)RGZR-*V)O:?$ QAN?0"&]7G5058Y+1Y
PUN0!<ZD\#A9LP!BH8]V(3KQNE]L&G'5\L-9D8)#3!A71(/4EU<Q6+HVI"X5<(/7V
PCYFM.GF@M:CJH^QE?:2PZV9 P&K)QHVWM>^'?;'H_D/(I(LM[CA.+JY;1L]L"RUX
PIG02[5M<]YF-.5@#7< Q2TSNQY7_N92&QBH?[T6X'2_R$[Y3"\L.3O'JIHW@?_N:
P"7+SD"C!)D0KC54)'WT8<GAZ=1]&7)P.XT-'+0A(EXW4M=7P@/:&92U$2]2X;N:V
P23 L]J %M(BPL"H]"G!["ZMXIIYW!N] Z<#KS(1Q<Q'W(71'R6^C40NR^@V #AT4
P X<N"KNMT"&7P?,#T3%/4_I8X'"&9OCUAF&79$4]E""#SX$;HNW7#E7(A)-/Q=7A
P/36&7IJ=ASA%K&EF/1*+K\G^DT2)8C=@%5W\I2%]//Z4UI!WYP-\F+9)S^C!RKZ#
P_3^RHDD:YV=U@R_6PANC#YDS'3&F5P;2VP+>#M]4H< T*SRQ%P:[^887EL2L.%#;
P/EQ1PE!)?HU+2[@'')@8=O.9)@Z!4?LM:&!V][9KGM9J6F>&?3[:$)[>TEB1@VD)
P4:MGVE@:V2=2]MV.W;%DHSI\[]IG4!9<NA9NK_2X3N/%#A=M*UZ,F!!LIHBI_F"V
PA.BV;'7P45/^;(U;$OT3J#2I@BL.QW1D%Z,"*VPC1%82%@=-?H8G!D9NL=>CNAM$
PW+O2!1]5P"+YSTBC@DAPE)W?$Z"Y<(_TZADLZ3S %O;(5)3Y5]P0! 10>, WP+_V
P?LWRU:9!,)58EAN3]1M"2 IGQ>WH:<>IV8RD-WC4"ZK*QGF.H5WAW47I?&2&'JT9
P- ^N\ZQI/4S#MQ\50*\<%M& /2CSRX82"D%Q6_AULGFZ7S-5(26WUGDOG=?F;3#6
PV[[60J:T8M[N=E-%?Z$I?1(RHRZK(W.7Q#2(U%ZVW[KEXM$KH5?3AT=1+?+%0SJW
PBIC&4W. &ZJLJ"5\#BD09;\Q*7R NS46-PX92+48BT X8S)8\BU.1T#9%;D*!O@4
PHN>LW$RW4FA?RG# 8R0"=+\#E].Y:/*I+QW,TM=7#/*^5-Q'>K%F LK"7%<-S+9-
PWNJJQXT\RY;-7). EH272Z$U^3$]D^-ZJ\3C8DLY(Y8NTM$4_#K3:1<UPDA4_Z/U
PVNITG1;_&7Q2BP NJ(S!.0CG$C);HP=U?Y+:,M, T]B8$8".9DV3V =@@@X\ O*I
P'C]4K8P(9?[OVU7"GVAUI24^;)"3IMI6Y<(_HMK?\DS- U@NJ:-4UC&[C@Q;20Q0
PX(T=JX)]7?);.PKAD9E^>5")GW^;*R=KA :E8]]IT!WD%E)LE;Y.)Z?!!@4<RNP5
PR72ZCAM$O."$B?:T>>$AZY$+'7MA!QMT?7V'3E()=-[(Q9?F;/-E(J3V5F5SY 66
PY^[X70\T<IQ@L+E0W/W<DN]&8>_NN4X-K%+3E#%;([U-HV'&U4S!7BIC:]4?L"]?
PG?0*<'PLU1?C4DCLM6JXD89B/>?*.-@=EG'-D<,-C!]1>:9G1#5H?>@BG;!UP)&W
P$,VGB-9M4X3X(;,T4"X4HA*S_TX^H.LPJVL&Z1A?H69W =U&H,B-GVC)5 R ]UX:
P$F$:U?$S+/$P$@@KM_N]$1Z#F\!,C+2%G44K88]S?7,.C/Y\2>_J"3=8$W76)PDF
P%,-:4'7_Q63SY;U[6'O=%617J5/2)KNZ6LG#2[ 4HB/G;V!).&74GJ@.0V%=R4_;
P:OL(CA?=/JQYAU73HSFPSR P48/;X";6#:[54A'3AFTT?4ZE&TU56QY1G^38DW*(
P'9H@Q,?5X;UR5PE)IJ"+,I_!.CHK>9=EC)!VIZAH-*HLBMYB_)X@"I+2"(*SS.M:
PHK0MC&^-?XAO$65.7Q+L-#)Z(QK#MU$]25P\.5WHNF"XH>IADGX1T0)\_@L0T+R 
P+@/1A'ZH_QHNE"17M=X_,@UWIK'#ZY9_/5:=T68RQX-OQ+S)YHC$U"0:$Q]Y/XVS
PN=W$'NMO5S7<8>X?Y^7LPR"IZ6"FU\WLT7VQ@^AFR%4<GB#3#->\;;".?XPH-?'C
P4L!:;E)402@^[2][UEEH6HIR=:*N "2/QY*VVF@V+T<$"9C?9\)F!E"I4K(6&)X3
P_I8PW6@;T)K[8F2_>OOE^>GMIKRW"U@P T!'DX^MS_1"A=P#)*%<U^2APK6F- -L
PD-_TFNSILC<6)(I&Z)_[&;TWZG[M- I45R]IJL3@@?(;F."?EMS!:]M!?8W<1FQ"
PAD$7G9$-Y+;-U/A&R$%O6_VB;[5G[] R,I8\P)K2057 IY"04_54Y?!,:]G9C56/
P&R=IP')%'\&Y=NQ*G"$I,,KN-*U_+[G!@YD%X5TF:=;[I9'IY%5;RDQ#.+&*P'\F
P.R:V]YCB^_\86@93N.(9.G#I\BV=XK($5!C3B4$CD6\8F;9C0<):[TP.JF-WN\&?
PKC]*)\LH/Q"XD5C0B:=LM-+"/J<VQGLPE8VZ#2R!G040!,8+4Z GL[T #(SY)1F3
P>IXDE4*8W<M_5&9#EV*AD[^!=#5NOH\!" RA\KX1S6B>V_<AJ$TXZMKH?7CQ(^@X
P_6.-CA/55U8O52(-:LG,2  JGLL#00I\<)QGSPKQ3F<S<*V/UH7((,XKIY$Z?+.4
PH/&STK8NA<J2Z_\V(KL*4]VO%Q^Y<J\T:$FP.FC+[ZW/XAL'CBHXWTD;",Z]OZ-!
P8>JT"Y4" 3S;7*C%5'ZUU<2\DPF0/T9[ !IV^MK_IR9>5TDW85BZ*";2MSRLI_K;
P9/?/WU[0\@==K<'ILYMJC<!'.4+0&^&,19>V?()5$RN_4\*9]?ANBONE:K*:*AJ1
PQ\9W<#89"(>K,7[RF*D6:'.EC,MT5NS2VQ%XOY-"+7!5)H(X*SGE94Y9:"LR2$SX
PIOO5E(<L)F*4N,&)-)PZ:37$YSB4EO\0)$PI<JLAG!(5C^<VCY;)N )C4%KDZ0=6
PRNB>5T<TG\%F36[ W'U>*!MRXV7V:'SU374#!]J:U&[]..B=3*UU'A/NB[C>>&T$
PXML01*]VCOQNP^_37*"KNXW(H BPB*@3A=A5FE):Z0B9:_C='!L \,-1MLC5,*^Q
PT+RZ@Z4'Q2M*)P?;]7ZEPO<QN!G,1/QVRN[)10HLV-1RW^H=3:##]T<W]#*(33Q7
P%@A0QC0QDY54)%=@&9Y1F!7=6OC2+WOE(UX1,3Q2LDD7?>:5K3!4_]-BP9ULK1DK
P*=3X>^<M)"?#6!+QKJIHM6AW).O830*DE)ITK'*% CZZU"* +@E4/V#T8,RM?FR1
PE: MK!2VPEV"Q,BT478& WAEP4Q;%3V*"@3&4M$1EII1QI HJ]E>)9<UY"5D%4JE
PU(=,RS\@OV ^@E8EJR.IIU.4#2 @,-,@N[K!D'O6VW+0&A2CS?PB@.'3^1$9/P%T
P=(S/[#E-)&4=$[PDXRGI)7.T10LO(]4-\GQ"3--<_ES$MP2GS"FR1TI"[;%,ZKYB
P#+84>+89^8OJ.?20(0M>6?)BQTKY#LQN3\L@4S?/3 !0FND.6CY0ES4@\M>>M]\]
P>G>X>GP&!;%PP6E8<Z1$OJ83Z=7S@Z@'5)6UQ:Z9-V S77#-H)H![UZT\[F&*JH0
PP^4:?9YC]I;"_.9#B%7UF*8G34DD_[9!7*\4%=TPX:0]!FL\W-)D5G5PG9P GA++
P)(6F;'0A+"\XV02(M=G]M!=QL Y J7"93X;?L#7"I0+.-$\0$%LN7AF]$7Q/12@?
P[EM(H&]T[",-ZMT2ZE%PB56 I1\IEPE= J5%]@<#R*7V[*Y4N6"0-><9,J,G<?IS
PWG0[KY;@CJ!O='$(F;]OYB^^3R8-6:QO4"B2_4W<NL7?',&D]=,FV&WT<AA[D(T.
P'-*,)O>,>. 6X^-LH130Q9E%.TX=_B:A6SEA;DQM C*7=D,TT@JRL)I4F$K$QV1W
P:=(/.)-*U?-&NNTAJB91G?2F_'J,#LL'@*70<>;<'M1Y@<7A8"&'Q@B09[#P9D;0
P^<0G@H-JS1U@YQGU)8QJBF.9G-JJ$7IVG DB$5;\/V"$J?I;)EG0(T8#$;KD<DL8
PIT'^O4_@.]4\&JAH+_*5?Z>Z(C_24)&1\6S"M X'&,NM\[&Y?3C<)>'K>-AYU@-)
PGQ;E+H?QF)VH__TT]<K4N5_E1QJR.ZE\*H6."L*T[A)+6CS7XH.G2:\\FFT?O<,"
P&-"4SOF9&?(DPZ>PT>B688_Z+VH1,.(-E_\R@P/>[]&IQ&L7>X@G[D.E0X%$'MDZ
P@C!H.K!^C$#<0_W)@#U^J= M)"YTP^>$[\E-O-(%LY-EQRC^]=$T++QWVR#H=KA-
P\@?#+8.@TI&&O)P*W]V7TEQAZL<-Q&I*KA;#<?E65HHM=+!XL?V<28,EJ$>&41W(
PP &2().7KM'F7T4#.42]SSA,5BG:A/G)O84WD%=EMZ*28&Q3-C,(Q2J@=^D7Z-QI
P";6?=J-3M\F_\\#WN1>Y-6VR9?V8YT&B;STBVK3 X]2PX9N]C&G]\,.YI'V[^!!&
P"H]5B ]1W]-*QFL]Z'$#1V8$@LT_6:@>BOCLAF-0?SH0WY&28!X/\S#'0VB[+KC2
P@MJM30)MCZT"5=O;F#'CT[/$3D+X!G:BHA=M1R;M>G!X1CK87DJY2/H[Q^!P?F&5
PW2_"(J\_^9Y(\/<:7*W#9B_I$7BL8]IZS(FV2UG3R^Y?D=-Q&OGE'5?)"#6_XO+F
P5U,VG,-\'M0INA\^6@ H+%I0R6%SL#Z>YMH^AI<X5+:$AB:'SJQ.0FJH]&13Q2K<
P)YIYRKJ$7Q3Y%1/?Q,DL9\5.;N/' :N\5[N^@P*[3F+IW5B,IUJ2*Q ^8#/E0MK:
PS3XSTS$S!_QB_._^BKMH:PGO(ZCW%":B2L%;%UQ[2JH0 / =Q3/0;5"P+@$__9^+
P2)1B91(LS"U45R_^$$28=!+2VB<:>1 ]>M!9@QI1F&6(_.\;_8P)K?VV.8KLMGZD
P*(V<RSR5-YV=-3LY-3<H GZ"V4-7 \'J;N\Y1/0]2CR^-_BK*A'J^ (%P\X0*Q0H
P)*^([9/A-R*(CN;0)&B+^W7BY1_U8A]S+J5%-^<AA:X#-3%\7,]K,(MA(N?R+_63
PCVV+5:R_KJ">.82ACT1D&-NO;_QJS@?-R>AEWQ749UKO:ERWEQ+A)N609[P9;'=Y
P#;&I"(L_U]FWLI4QP!G^NI&3]U/J\3+8Y@S$\&CC;8]W7>= P__4!*>T7H)T6:P^
P%R^O*WK':834N(?UJ>#2'7><?VO_RUC:_:CJJFX((;S\L$#+ #S]E0CI0"S)DX+$
P<@Q=#_O)T_PWG"9.02_:T%(X= , :LUWFD^%&D#D)PO1**! ^+H!S& /QY$<PG8V
P."64AN1OHP8AE4^GFXT0;<@&I]PLHI\%!5+;2,2;U6#RM1 RW4X8@!-Z);-:\RDU
PLHT-8! B."R]B[2="^96*4FEF 9$,,+'['*13Y-TT8Q'+/2G[NW'VU6E,5B!\]'M
P)Z?Z.WH/"D#FAETDZE5]]-).IAK%/8:R5Q%.DX.]&.=L:2MUO8"'5R/:/(_D8\=Q
P5Y&!_FZD)5@'Z;73<SW!-E,]^!Q:=C/@3^6U,A)^!9T-[[[<.Y9=43+MK\P])X'K
P8\A/'*U-9C'K'^VVN?N-)E(JJLGS$P).N(R^5_U-8+!MV=PA6YBEB-GNN5EEH'?F
P"$!_H(@Q1U?U8\D%JDE[69H8L4B7^726'1A-T A:'*SB32.T\0](%$L6RA#'FXO.
P[@M35^:"Q65MD +:]J&C[RPT@(USC-\+8C(#$CC#;D.4YI,(TN_)%1HC[Y^7SA_Q
P VYBI11,KK1AZO=:4H+$IA(+'-_C/"K+R(SLCNMN(X@9WQ=@10^TQO.Y (-!.E5N
P'U!^[/4U/HA'(/A&<F#?68QE7!&2UR_2&?13>,P(59>I,T%U7X/G1,<3.#<,^478
P[FE0+@&//$/$DI9/IS7"*X8A-\71(6.RX%HE]^Y/+^6<<:GP7U?O[+-')@3U MD*
PM"Q[+R&6SD3DTJ0>(,6\:1)6OBK]Q SRL[8N4A];@T(IO$8J'PU0)>5%J@4N !P*
P.L\>T%=J:$JWEL?V:?"#BF.'?<NS-4Z;\7I.%V@$/P)';-_JZGLR?RG(AVE(69GS
P0#@U,"=L,B*D8=5K'#6:8/:NJ D8,)HJ840$I]+\1I1Z$2>E(>#4. .3G1X<9[:5
P):/+ICG6OQ#:=P*-M<* _*:@6&:I#>B>%]!V428M*4\6)[F,^XO&7JWCV,^Y6H.,
P/T(TU4R7$3\&$25,9JNJ5BO)PL#^ U=S\[*C&GT6)8>7$RUHUQGHI:PKAV'LF[3#
P!* =.STU<#5$] 3=Q+5:NGD(=11'M;.-SKK! YFZ$U-CW(T! ZS^B,7'9;*K_0B_
P4G[7"*MS"F#D_>U;%EHR$5;786%QXI7SCT3!-C5IGH+N7ZLXL]L>\RHWES(*9$56
PP\>K>3UP;1?Y*KQ<..VUI4<.7 9]B3S))S5M<-S7^2FUZN?3"^5;T1@G06?'57N%
PUOP!40L<$F^@ZFW)!!UN1G_N^H:&!1OL#AK<XI_'#AI$/]"4$F:?].QCWU <4_::
P_$V;.E&;'09"S%^N.R8%**,#1VKZ-L,$S>#S672CV5ZHP7VZI\7%$_5\&7]1>\2!
PSRQW*U@YSB_HO84C]%T-:)HG=7(3I0X:VLB\[*GM-P9OM:W=SBP$0P,(70KR FO6
P8FFACTD-(Y!/S/#D]K&.J/BY&Z[M5$P73^'NY,6"NYV4(#:A-):D(<J&D4>K3MG%
PL_60K&JG"VBJ-VPW)D/1+6I!M0>H*Y>)FM$['.K%': $FWAXH4K' 0/X_K0U1KLR
P)T^Y9%O7PGH5BSJCMN?>J.]EPUQPO U'[G6<D/TS3-4A[)@5QH CJR15G/NM]7Z@
POMBF2-FV/H:".7RI&\,U;EK5BO2D73"R%[M(7%Z'+;(H:!"FDJON\+*0A_L9@";B
PJL(SR6[-RY_4*');(GF?)ZSQXL\*6$Q27Z0$J2S*:'PQ$'T-Q>?:*@DZR@1 _L8:
P9<\ R@J"3 N%+G2&BC[PAG!W4JH$O.J))K"<W<=B@3664H3M!9(][,$*_A6P#DUD
P!R;IT,4U\[Z:M@#>9_O]?WN%146!WE5=5LFFP(SMB>&=[LMB)*G']&\)7][\SPG*
PN*0%/X]#^>B)I.VN4>?'0F3<F2B:!!<-->%%EUQU8M*8F@B1>/+O$T<$"!@JQDB>
P.!=2>X#S_S.0!HS]U3;81WXWM+WE.; 3+ +CBM==O?B0I4W>ZD.[K6=8&C1 TH46
P'6!9#$,G!W8A#V[-O8'2:M^@@/BB<Y/ZEJ7^ PF"45?8(9^@^=""$)UH"IV%G'E5
P- Q:!'W)ADFVZFM(.92W$CG[\C/D%?(2JO>0YT(.=V8/2:5J^&_T&; </7G^9TZ@
PA<]73G%#S7VE!4O*I5^U'0.5Z91#4@G;H5W=E,#ERYLQEGI$R'5Y\@_$&5#R8M2L
P6 J8U";PEL)W6#!&__71&=,=XZ:Z=D@,*]D5A'T@S(%6"-(?.>16(WMH,TE9,(9A
P[4QLX'0DFO#XBRP9DKKL=G&2_#7Z(5E\'-P R&[5LN%FD4G(&Q9[D*,R X;4#M%J
PR0ORD3C<'U<UKG9VN,!G=68OQ_FA1IS5*)L3R/WROP;N[?</=]$6KM.O<PD#3C2Y
P4@6/PD <9:\\<4WA1%QQ7A%Z;C,U)VX\LZ92ZRSH[+U5TO[6GE/$;\[I#=]T/[VB
P/O^]MJ4EYT1^M8<YH(+S&,R,VFL07;T,SLXMJ?V9:2"G-1L.UZ.E;JD194CYVPP?
P^<.A(PTMS?FL3*<U-N5]A37\?3D>E"POJB5"+?F9\<[%JR4*/_C?+D8-ZX43L$%_
P&CPM]CYA:::HW0!:HK[DI^\JT9AE@*S>?J;XV^V<GJ-8WNNRH@-1M^(#_=&BP0L&
P#+^%WBV)?H+<V%@C0DS'/<;XA#IMIW;Y7$_ Z3:P0BEM_S/]D.F3R\0G!"-XQQ,F
P#V A$0W28$B5::]8%+ 8?8CWZ;:XF'QNX^?:T7&BE[N&;!5<:NKBN$Z>_AK>EH+#
PE0;M -%!>9(-3JXLR(W@PWB%Z!Z:D<.7GU5VI21O?.%2!R8K%TEDXY==N_O1^D5?
PB=B=7Q**<ZT#F/AL:DM_2/QCAMI4D5UAJ!_8?KC.<%2*_R>9^"EZ_Q$JET?=OW$^
PEU@RS@I/@MU8!2%'U--69$ 8\@UT9*WF"##7 )&)S1];P3LQ='[CA9HZAF'BMWP-
P#XJ[4+B:*["'V%+U#.EI'2P+T"5:_>1!'PDP64=HCPRF%C[=M5?#.P;Y-;KNJV_!
PO':7SD)*N(VW"5;*$H EJX$D]%*SU->04-P$#B'FA<C7-XEMH)RLTZ'8C4UA,,#<
P[Y\,V/=G(&L?S&RN5L&HAW5&Z 4J0L7>)N+#>= $P]_I)J8D(M(9O>@%!UV_KNUT
POKJ)5#HM1 B\<Y$3B(>6V9CS91)IX(6OJ\=(**B\%13_'DV<_0(#GKAGKCAV!9 R
PK&EH&>YK$Y,:F^:&F#+[&DF6X[SJ[UBJB VXO5/;NIJUL"HAD5QXSMO\!2-?T$^"
P;@<COQZ2EO)R5DV<\LY9PH-LXM&^(-+ZE]3:Z&Y8-#/5_,EK[*Z4CN+J2NHA'=R4
P*Q>[Y9,RCX'@8X!?<:!ALTODD ^[]6T N3Y46N.<#*-MMOLV!Y1'%B'DB!2NI6;K
P+VM3,:)BI;E=J=K?:%-2BUH4O$P&6-Z&V%2KV+2&\.RG.P4K=.:O_] R07BX%JS,
P0V4@'C?/H,DV.YKT$=1S4.',R%+?VW"\PDMOVM/NU&J(C9Y&\V[7N 5XE:N.*YPV
P^_9@C1N^E"NJB!BXS5S0Y RJ0@,#'U8'9=$'RE2U3#/%#20EVY _>=C/T)E.:S.R
P_]!EW5:"0X^!S/G$2Q(LA\7 BSP!/W2QZW[E3B\)\/WN4T=4" ^KMXZXS>FC(:U=
PO<E+D,9VKNVW10:/UWAQ3>Z7+OQ'>!*C,R,U6OF&F >"%LED7RF^>W]CK*M!1E)O
P5!2.ER8@:^MH<#A5F&EV4@[H$4'HTS8"%IBEB5+XK4O]9I;M=":32]J_+"D#K8>>
PGQN.KLZ]4::>&-_(BWPI&V'A%71:27ZK9GQY7=Y0+!Z'U?3IF3/,#+??.@F!E%MZ
PLGU#F^H*A-_@F:ATR.9W9R)TU[%L(3>6.FE1S7POO@!?6A.@&"@V*LH*34 F-0J+
PT?IA@Q8.Y^JB<=?)QV^5)9?O@W[B@@#SHF\&=-W!7,)+59D\ U,8[;G5H"NOV,)<
P  _,WL$$ PD_-!+=NV$0W$\UD5EPN)D^-Z:5WO5T&=5QN:.-Q1E1%_\&.-^1E*40
P.!6;I; LQ1%9B_1YKWWX\4I]O#R7W@_+WDM9+]"RXRUHZ+P-5$:I/XUE*$S>+G]J
P46ZE HAAK\6BS^S-,%M&<10/$\ZF_<@NTDEN]4$QB.R/N?(9ZELU)?(,"7[V_C/(
PN\0P:F@<-#UMOEJUZ.KZW-+'7 +JC<>9H).[%Q[FN!-L&+=E;J6F7OB3L:\SA)F[
PBI>9$4#3RSSD2RWI"0<UJ?[B>=JAVY'GB1@CHY'LY=[5^ BT6%[GS;[(DDM,,/YT
PRF]A^L4X+FPE)B*:L!ZOC+!P3]_!>H%Q&K>&BQY":#EI^5#F\G^!&4*%WU$+Y )?
P8&(; F0IJJ1,*?%#?'"UKUXI6/F=-*&EJOX;*#V2ZV4ME^R N+XPNI0QL1"%6(U9
PDJ0=?,'FQ2BUV?\_F<=P\#)Q($3%V3/D??C$CS:H*:%3L0!2D49L9./##I+?)-.9
PZ.]'UI[:/V9[06[I%O#=FD^5><*FY4D"O!3<"-;2NA%E^C4M<#?E%L"9N5EB6N)Q
PZNS=)IT$*4 HW!\E&YC:*."C-84%AZ'C)'\6^F$@WL6B.'%YF\=PGTFW;VK\SX&Q
P]OILM/!7)E2\R!(@%'Q<D$R\$>_0-9:E.WK8W&K9O]BW!"\ 76Z9HLW',#%KOO>L
P>0*5;/>C^DA"+DPMI<^#-V<3:X5#1Q%F0';R3EM2\UMW(&*GSA_[U)P3EIX#LAR"
PV0;MX[G4RD?>2E7P%O<["\!+ACH>W7T4?<O2_N:3KB>?%X=>(C-Y1\%R<9I2?4[T
P18FKEQJ]6;=0]3/CW^N[_-"?U5-1=W"0\<@@/92;9M5YE1C.3/^CND &<DOE/7Q$
P;.=B3LC/HEW+QP-IA>Z2:NUB!'(S4FL@OEWWTTZZ;.3H783IN_)D*NI2P[S1NP3K
PD:O*J0ZPQL L!HJ=X6QSDNFS/QJSFI]3"V-W_%27Q);S$X2W]"Y[<2\*$Y8V37@;
PZ9 :K$AU/@.-</WZU:0I4E9XA@O.XFS%#MG-7#%P>\_>=QY;OW;3!>XQ?#<8);]D
P/>RO:DO$<+,7_]I7U,M!!D(LU$$__M2H:FRR7S^%B3++B$*".4K*F*;F)FB".&,,
P14T$?I1XC><ZWTP%ZB=*Y=Y/O^$C\..J [VZFDJW\CBH!:NH\1,4T;W3M:$<C,LS
P@RB N+;N3N)VH'X8)\\K-5R:U9)K$2LO^0.IS[)V]&EH&_2">$N4'("6B31UQW]0
P(T/(0[@4.B<$O.(T=BZQ<6EWR3>=32U(V7:J:48='L0"5/:@/N0#XND<VN*GMWRV
PU?XO(9 &@*M$<7NU +R%W-=(\D,] ]0UH:-'7#(Z3TE[UB01!.R\[0X51; P>J9Z
PNL):O%;)@6F&(\(KS8&QL&-B]@:T1;0E1\N_>$S:(4V\F^K':0G]E2 ])PXS^19^
P#0+H)@IH&7T@W,@ZO3HU1#DWFHV+*(&X>@!V02)A&$(7_>2@GO2H:/M04&-@V\%U
P#*E^Z\+S]\I5_IVE&SGK>2YJ?QW5J&*9HSS.LEQ>'K4H]R^YS+A+?XQY7]O_; V\
P$Q\^GZZ5R#(*03\06?4I,T$N?1G-@H$[1\1=4J/BU0SRS7P<1ZMQ[SDIQI>NP,]3
PWUU+09C1!.)4&B=<*]_A)A>1I=BABG.^J _6EEU1CSH4?7C'&\J[1L'T^WF;.EQL
P/.7T\W.(]4,0/!5JK?7PJAZ98K_BSJ$YEY?BG.X;=;5&O&2:R,UPR)D^0 VNUDEP
PXH6Y[F7L/9CB!DQ%$H2J^P79:F4:==5 #Z3'%6>HAL/%GRCIR,IY! RTZMP7!=PA
PTKWZ_NDJAP:![ZK]BS %6%.SX"P]TJ\!K >YJPB-A[PV+N?"E5[C60/3]8=2\@XD
P2>(X[%;(]<2HGH!:11O"-;G[7"$D5QP(1KP1DX ;[E*Y"AO@^:3"=%JK'[UC^^P(
P?ZQ;\3>3/H3L*/P8B@[K(M%B55JR'T%)D?I)M2+:.;S\QA(30IM]XFL^DOMK47VW
PS48X$'))^>3<Z!#MAK[]T=T/M&%Z1*>_,9V5(S3YN2!R C E$T3'9\2PL\*-"W< 
PF8]M@Q8%;'(EP&A0=M97W*=N3-!8U)Z4K[ [YB<Z17P&VQSXW. R;+8CFLE$$(._
PA&<;-TK:) Q[I>HO.6J<-IUR@) GW,$CULGI$D:[5:.;>NG']&B!1 7I%(NK>.)+
P"8__S1@,/9(KP#P?7(2;HS%<HPBV8O9\ 3WP?A]P!)=K(Z%_<*F4)N-02YX:M9->
PY>A:- WT*7:?!SN[&%[20+B\J>.?/_<0@(D6%B7^H3[HU+0P]K"?)NLDLW[6_R^'
PT8%^"&W8\TLRUSVN6N)FL?$;# Q;V8/I[DOEXD#?H'"K2-VA@-#!832"7.JH+\\8
PX?3]6+XODDM+V;>!5RMX07+KC>])9038IKU263MC]W_;;"8I#;5^&T;,>L@*_ \#
P(#ESL93#-A*5U1MN@%;#<DMY!,:,5IVI.OW=-M,5OY\HI&F9%/4GKZZV&O56)HM(
P3\ZV_OB "OUA$KZ-M0<9FB&'<$XP9#C.1K:T5SU^[R_NQ.(%2HR3,XSK9>IR0- S
PK-MH;#3<WDU=JC\5*ONE HN!K@U:C<?UH:>3*H2:^AT(2 WK>\1G/-U*QSEZ0%==
P#\5B=[H\.M_ 51.:Y<9H-*4'I"*)IE9JDC^7UJ]ACWR)98N*ZA]"?+L&'Q0H8VRA
PL96ED$#^DA-=)TL@<OH&Q4>( 4R:SK>\4PYERJ3E\%961_M\[.G5DO+-,$7 VT2S
PNZ3FA/TS3(^$N>JM#U1?LU_U*JV\[,@/]"WW$ ZOJC^,&RW+52^6@I2VJMD\;Y>E
P@M!9R"7GA4S05^+1.52UN6VRI@COV('7FEN.,NB6E+%>J=IM>RP&N9^IK08.JT,/
PFJ1N_8^63%(7+L<#A/Z!+3R&+;L%DVAG%+/PBF1^#YQ[C 7F%96/4WW"N0=OBK<>
P,K[.\+FSS!81;EE9M'5*3$ZHDGJE2Y[HJ:#E3C%*,J].2W[4@A9H!C=KWBYT#W*1
P*!GMI_HS+N/03=)JST.N,2EG3(S!U^0=W4Q:>G6;D: 64^5WP+AX(B;8-6I R$+6
P*=YBMG5\W7=RAIK/R<U>!M/FE!IY6#X$X[>OWYH>\<]W:FW6+@_2<A&L"A2J9: J
P<*8MV_9)HF&/=7.(0G]]V3QTS::%W\_E!TU!M.N!FUVSCIT<\*9T>'_?'%IB7U/^
P]>^G;>9P5>9CT]*M5^PRAA$0P^)MXEQ Z1I:(]B",5/0B;:F ;Z)AODUHI>1\/U>
P^2V]QO+H&DU5@T*ZV_)8K&[L)NTY:0+23)V8-/J;2D@9B)8/[89A_3I^D#/ )0:O
P,1HZF*@-_C7*0\FG?I]>LJ\[E-NQYMI\/T>Y,-14:Y99EK8O8X[2=Z:\,/0##'^@
PE\%M8-TQG=TJOHI;M@19.J>?KPMTXF2N.BZKHQ3CLOP:]JB0W9ZTIBHY9,N=W'""
PG6W6UI(IEJ'7P2N/_]_;G@*(<Y,]H!2RZN$:2T_@3)S/WKQ0)+C6I207W):YN_KQ
P!OK5D@N69_Y[]'M ^-JR9;+3O9N*%Z;:=8I&)5^1Z0S,V/W%O,[\0_90K$2L^$^U
P9";L0[I^#:<'>@3G%IAGSI51\E89H(;]N/*(H=@1%8(\_S;HHJIS+^)A.UN(-KFH
PXU9N>0EA4>LH^EGK+ZI>"X)^.RQ\4!B%A)K%J5.&L%IDN8#.Y*3X#L(=D0"JKE?E
PC]IYXWKI-C$Y/>BW>N A\FP&G1FX3/#'SA*TI/RIV88V)//P9!!JZK\EM0QGJY!S
PNRAA/.4.$"QGG-;0Y>M:8 U2G&(9E^26ILP D*LON(2#15*D'P,3FLR:7]OU>*I@
P-^)[L5\\CZ<MWX1#D@R)O>[5"G+RD1MTF5!"]1YK/9JX035?:9I&C]^UM1%[L&DG
P;?I#IC@/SD>=ZOAP!C%W(-ERD2V&?WPMSEIAP3\L+\YWG5O0<&,>"&O.Y)+H<7?H
P0(2"IK-RPE2%:5?MK4.P'P91^VYI"FJ5LI#%@DX[;%@&I3Y7MX\%BD*/A&,X"*L'
PMY367(Q <(-V6P[S1SHR>B,%I$?\)/''-A@H X&).\SGS2:Y+#YJ0#/^?P!F='QB
P-=M_Z_@*2N4;^OU"6Y>:M._VH5U0_PS,]\Y4*_43!J9C:<#N@RRU [;]U[4AB5>\
P )5JVL??;KL-"OC#0;S#C:R@8+85S7:&95U7;%5H5KK64-;M1O'3"%B8\2,YD_GU
PG,>O7I)V_Z0;@Y$\]% R8/*D@%)!S'V!6U 5[]A,28]BT.F5!\:R6B(D_&KJ"R!,
P7<?Y/_V74EN)42@2MD^:I4X<;*];"CG(PDR2HEDK#M0^VFB[<G$-_TDX" 1Y%BE6
PWC)+Y3ZC NOCG*C7!D05*]64>2* O=&%6U7$LS*I6Q>'81>%XD\(##-4=]-YRS82
P:^;FZ5-,'H7H$D4<IU1!1S]C[P>+JE/MG1I[,6J6Z0%ZJPK*U*WA/W>C9.R&F%R 
P^4\BUJ^,.>N=P,DT@%MV*10,C[7H^:<I9X5^?HU*?O@7;)0A"'M (>@.E\]\G\^:
PG &\,%UT=YX(WD65_X2\@UWJ[-MG;BOYR[U>Y-=]S9XB8HA?1E9("5[[59JA2?>@
P-L)BQF^X-118!V6^]O6DQ082&;W[H#0'BW*Q/S@1^^B0BQ+)6E M/+*Y=]H'$I!N
PNS >.C\RN!F9Z+\7\$A26D>/\4:G?ZS@]D,_9@(O!1?&8MC6RGRVHLY(#;F\NR=X
P<>W?QZ]>J,2#8%MR35_ELM"O;0:1,^/]%!2W>:\:"7YR] J%!5AYR JHB@-4$_@O
P+X.?:X\Z( RFT6]'T?AR;W=PA8"?R?1AW5"N+G&597LT)/.(D)OGP8>SPDASD[Q^
P4%>!2[O'E,H'BD]L=-@,AD!E@YZ3\V<X5#*%)KI<7->!WJ>4K<S\>&S/#Q;1>)43
POA0_2X0#_8$4F+***Y+%1)\ 9%249I7\_X@BQ;,:0CN[G3XN>%?X7?C'F"Q.A'BK
P/]F[STG'*(#D,GAJN%*%J7XJO':W5R@D%4_SA#;+[;Q_1.\;%J?*#(:95KF5$_O]
P3@"LE^&?!D3Y.H#BR14Y1QA/:/2B941(=&'D'7]DCK]%'^"!AH8[/=P$M\LH;)E%
P51VRJ>DK!1??T:_^4]<B(&A>PD.&>^\P&3)26=)Y+\0"N4TW[F2)NX@ZHXW<MF,P
P G>Z9EFT^R_#E8D]V(UG$-=3U=2H$Q@T; H>9>EYQ?&X#JOM6UE*@Y8.DU&!ILT:
P,JR;ZF+.]A-(;H+0X&H2XP]@!XA]+%/PYY,ZQ@-E+F&Z"D$ZICL%+9 V[RLKV[F>
PU4E\!4*2'0;J\RZ,\J-1I_1I'MVC_7S8FU,!PT;*TTGU:3NR7, O.I;F9'Y.Q8S&
P=6:24!0-T6ZLDJIT%%5W+;/^%#!?4QF\>(TVC%POU(Y%7/?B_.W;I#%*V;O"X5PF
PW_#.2@E2QE4@99;@"^K*LB62#R5MPP9TP%!"\RWU/6\!K**IFT!!]+$*2;EY8,:J
P(OB"ZHVW.2;$Z")4!BZ;KEP7(W4%V(]RS[5W_-$;1EN::\#$Z'W5/@W&#NV-^8@E
PH!F3!K=)L_V(^G%B53R;D<)'(OCX)M\E1_CCGFX^*;SV#AXI&\!N_?F6LBU+?%%Y
P&FJ)S)'$#.;A*FL,\]M@/R*B7MBLC $<0QE*ACU9H5]QQ/G9H$9#(PO:P4O5)-?:
P]R),65@9]^L8^AV,'SN +\]1%,F.&#/3/"\C/ &R/T(0/?L.,1>7Q'7*8-62O/Z=
P/_$S9M(F)A<)\"@1JZ/=^8==NIL@*J_?(@$REI,5=/7NN_:$U%8/<8T@2'0B(;3N
P*,Y?B.4:3<@$CX,+/J/2O@'B$35>ANEYXD@PS^H&SGPG%@OU8Y0B;A9N*!JV%53"
P\$U]D:S[B)M_I# DK!$K1$++AQ5LL Z3BUHEH*+4EM1D3",B;+IP>G57V V)32+Q
P&)ZQ7-BT,SA2^_0-*X,+(+#L2LCF"'WZ[J->QU+OM@G>B6+6]II"6G ZCIHD98(8
PI]JG#Y(%1[#:)/2D/O'^FY]0/N>.PZ[O-X(8;5M5G(N,LAV*S+;X_6!.\6EF0#Y]
PVRV>7H5S3WM,[[9HQ[-:,+0^$5I&H?T>O3I28IG%]J 5L:>"HE\'\'8V&R:^:?5 
PLW+.O-NCE=2N%6R.^X*B[+:K+A]:R:K%IW%C8'(UOU3#OMSF4<$#)Q -7.&9N9IA
PY^2MZ*$*G)2!)"L!.DK,9=PPJE:U->TLYU0C;4 OVG[.^^*V[U%!\&#.R;Y*E\1@
P413XV"#@4TB+S.3+VU'II,;J8\U1!W$^IB_%[&=L3-4/<_'_U\FPS@8\45ZI:_EX
P0@_2CI4Y_MHML73 U=]H%,(ZCJSOT>B4)1BQK?)_32QGY2LP4QA @ARMZA@Y]I%3
P*/>DBBY4'1W8]NXVRFC/M.'#_+2\Q+P!D_]QGK0E*HI H#*,M;7LSW_B#<?%EMF)
P@7&&7A**$#A4+NVY33&OHH'B/T#^9V<RR0R37G&U#]E*M=[Q+M!C30?!XE-@69)Z
PP^HBLAGP$P3+L[ZX._'CFYSJ!5_ F1>%-HF^8:RVQVNK1._W@$R68<P"-\^ $4;?
P_W1L3!IO1<VX.20<?FA$1DL-X46! #9NN^"Q%;(' NBUK8'-(M9N ;=+%I4SWLHZ
P5*@1M>/OKDMO[,T?X:)--T\>YI?6BS6YT6$^I(284LSYYUN15_]9;PY)_HDI(9S+
PMU=Y).S(E#R85C^=<"5]"]($R">5JYAN.A1"OD]E>06/.,88KD-#LD7;NYM_;U*X
P<7 VY8P%)_.[.8P#BA'J+UX_78T=+AOG+D?/&+FCE<T5XY8]_R@'FA(*UL"K6N3B
P#)!!,IX<D)<K$X?-I7[XQ1B&MAL\5CA <GI.8"+\7:2$0Y P1N5:Y[Q-=!\DH8!D
P?FS#\FNBP!3G7<;U453]9 &?@(!<+D/B&FX$QWA2J-TI642Y,4^#F*5H>5#;"'8D
PLVJ5>JC714NETYSC?>DWG&O\_9I](\-EL0O>UC90UIE:@"Y*(F>&X@5^OI3]#GAY
PX64PJBP2/QT:M>DE9ZIK\4B65<KRIXP%KU26+Y#8'[/#$X(J;CVR#WGC&%G\L?:^
P^TK@J2#5A.%E4F'+_^0C;[-W#)8(X<^;I\R/:T)S^F&1Z<AEB\0B^4_V;A/ *@23
P#U6M&V;M_/"P3)*O*F*NW$VZKY6E-H6< @!#+[#C<X[D3US_QN-S,S0(-SB$N@7.
P2RA#%6MG'0KHOSHC'/U/5TW!T2 Z#E"J+[J2DW'^6#(CY)"PK=3F_7J[@+\0'.,$
PBFQN2RF,X,JO6: )RD=#0\XXJX@04?HDJ*;0ZQRZQBZN;K_87NJLENUNZ,%7A@;\
P0")+0C&XY1E@COEYL<2+#8%T8V474)N!A-?RE+SKN2=%M79-W^ZGEN8L@QK3)T 4
P[4D^WXAYU-A,"V\*GVHP(<-G8'*9G26.%@KNN(W%6QXEP*TGSR&'=;'SXEFP#*%A
P!<GDYN+TI^<E]A$U*4\@.BE52^4RLHI([=I(JL429>0M-&CCV%Z>L2)0Q %/U^[>
P].WS!7U'W47>8$4'F<=X1*X85I32?IK4V7>B2Z@TWS+1/7GT7(/F[&V[932M0N$@
P]KNNA=L:CG:"=$;3]D-8AEGM I%,>D(_R_"A^=7OB\?"5U;YCT>F(ULP2IF"%0,&
P(8'/)G3>?]@_$]9K*_7^4#"+:*JEZ((NIMG7+\#]5 I<YDA>K/6(..MOX%@O-Y.Z
P6;:QZ.\2SVV(JT0$L&#7G0;.\'N%Q;&V21-=B&/=]2EAFSX!?1DJ5(#Z4M'C["IO
POF;) G6&Y*]8<']?8M]<MBN)7((3)ICM'F/+B6QJFC56<<]4PNY$V2D:B$O=<QZH
PUT1 4I!N>]3DGA!.KQ@_5O6+1NI;NDKZ7?Y.67RFJAZ[T!^D-1"YRZ[#\UUER8&7
P*5+9.G\[ZF^4U=$.OBE$P>\[LV!0X^;_KW>E3!9$2$%S;[ONJ%#@K?>= S%F84YC
PLX! 1*W?K O^:HYC?O]JI]A'!&J)S]:@Z9QL*Z""7=K@G%8=!T=8+L.$,M*;PBF 
P@S YR)6>*_Z8K]<7LP'^AHV$*( U([_&7>8RQBC?;G6.34AS$<\;G$_I5_0-86EE
P@$KIPGW!Z &I\>Y8>>NG6NS*!S.T@V8M08Z\*QFF!DWTI)JQ\,!CH?2%?=TS0\,R
PF^V88#_J,O;YFW>RN3YD96V4H5@[:6WA96Q/$PB'=U/EY<7CG\=.G6%[O&%?2U(]
PV6 2##D:8%1,5.C+2Q%E&^SX)!XD,]))\5H S1(BM^(GQGM0?874]/S<^ZGNE08 
P%/C5P%AZP5\!-MU[AEPD9+WL(I4P>[ERV>%9C,H*38X-_I6PXEHQ ,FLBS9AU2Y\
P=9?R]0YYD!ATD=S0YBDHW,N3U^1 81_'%;KK529T8X[IP?U-4K+DK3<2HVJ''531
P>\/Z)[6I1XVMB:Y<Q>^=0.A]&%[H?2A\Z7Q(@F69PSR>X7K(*.K#? TQD]L#&PT#
P;R[4Y ,WF;Q3/A7.8X563%_KDE8$/&/FQ,+K<-#=_6R<EPG(R 4UOHY YEB!Z^YG
P/1E#M"\F& FQKKH2FA[9@*FG M1Z*O 0[#:D=B%'.:-D$\SLX%ZW,-_)WNJP82%N
P "-/$'2BS:@(YW?8F-\I0.H?S4<E=$N#\NV%WCS/']Z1^47B3-MMV14[DO[/[W( 
PJK"*.6UO'*+PP9]L/:/[F>&]H36Y(IO?'5[G9-O C:41/9(?_"GL(?"*3CD+(UR%
P*,@!#X)\6-).9JZ*DR&Z)%BFN9 "CX3'+.BU10HP?&7.XTN$41T(!D4VK<4 MUS'
P,^WV$XEPJUM9]W1P_FUL55V@L"\_J NOAVV>#^]D8<$2CP%&A?&:-$8V2RYDLU@@
PN]O'7UYS#[M419]@+&#<7OLR%8(V9N335DQLYT5^,B#@PH2^:\N02B+Q%CMMA(B6
P#B,B4R>Q(1.VYNE9/U;B9IG!?0A66A7Z=(JU3(_'SA\8B[6=?H3E&2??4TBN0UEB
P,%6W_8P@9GC[1PZ3]Z[I.N[[B13RSGO6XF%:%ZZIY$B[)*P_>WL!VI2WQY0^.0G!
P=E,@3T'/$%4$F$W2A;6_RX(\]:G7_#/!\!7V\#6L&:4S@E(.5!L0U]C^ <H.K_F%
P,.G=KB()^9C@6!%TB27R&WK,B-^%YX_;YP!/T/+G/KK?JRPJ=BA _/_[*'+!T5GS
PUI?4A#SX$,:_XP  SYC<S>XQQ-Q(DB8A;NCM&3<A<XZ75\_5PF[B?)<_Y.I[6T4F
P*-3UQ* HQE&<$ZJ/67SQ/6(A2@14A(&0<A1"O(I7@\WH]1!A6^'%H>$D>A>]2@[1
P+T#Y0!6=Z.YNI";FD(K3;K_;?W'ZK+-85HM<!0T2Q8#OX+68Y1M>=+I+;Y1,7NW9
PDHR@;SIQ^ZSN5:0WTHQJW44T1?X:"/878[;3>V^GH(2GGE)6?L*@H.!(@_O_=*ZS
PB%^R7&DM:4[D84!5'@0L#?W\&393/\A_/!0IN"^OQ%[M=%MFIQQ,%69C+VT<:G@9
P<IX$ZC)IEUGJ<VC,=307>BH6GT#;-$L#X4^1CD[+=BBV@!P 5##\%3P9D)H+(7'2
PG$TN=5W:J5-)0XDE,QIUG<A=5=,D%L^ ;=XRH0[BS>+H2X',E48I4[9?E&O,[YW<
P%031!:"?QRA-A8AA[)938UI5Q[Z/E3#IYVA3((9JMBQ(U@SAHB3FP!%&J\(&&A0P
PO'P(5^)UZ4?,"!ZPL!EOUA!?D9&O!,,'Z.E03=KMUD2MJ:%*=SS1YV+DR$75()<4
P'[&;2 !SE^""5;G%LZ3#1,%PTKIA+*_GB'Z&'#LB6+;R0A^6QRFA>!YC345V^)]9
P%X[;:"E?OLH\7&&Z?XD];>@5&B*V_L][260T$N?CY85CKP([[5PYS3!AZRR;[=_Q
P=O#RA.>S&>+R/=#-RRT4<EZ$I9'K]=OZ;?),H2I:=ACT-$Y@7EB!TIV@78Y[0)\U
PM:E+B4OOWXNHD;H2NZ<[:G#A$?D#Y#@-+I,A)/F/_RVGQKPV/J-.0N76<J_*H@Z6
P&6M:T9^*U(LSLQ:SR#YTS"+,<J/OE03>-#-"JDEP)+)3ZVCFB@1\W>/NO*9O0CT$
PC/]XJ T8YL7M5=V"X,]5?O,Q5LB@_U2[SOW+AAR?%C1T\4\](' 26\DDPXEF!?"L
P/_#Y <3#UTGT*;YA9A<G\T)G"P(G[VV<\(C%NLC<)[.U6F-"T"TKG;]/,>/]YO]N
PI-?<RX:FW5PX.GC^Z_[?<=PGCFR6E2,L4J:&U]BH0DKKU0#MJHM%[Q?8OU-#.P"V
PY05B2F;5]I1:28Q],66C52:B@GSTL(V[0)O>]!)M!I:@F2L0/TD1'HA\8;%,U^U7
P 5K7<]@P\,&GQ-.+X;/+5')WZ$Z7F/%Y&$C'_PU>@Q[ZI8$=R0-P?^5S"LE04O98
P:,./TY,V3S>XH!:(JU<UD4X.2GD0).P.5P9D ./1D[3/E(B<'7;MR^) XVS8MQ[W
P^QC.-\O[)"#<S8NW_+>==F!DJY504M&0H0*\8_<T0.8%ITROH(AC\*^!#AAAIE:@
PKC/V7JXK'J&ASI0V0D$&_.RU3QNTP9GR2>!C::8NB1);$B.)84;X30=2F\:^4N%0
PAK +>29J/$"1^5'L1/Z4CC]7%N%1_A3<PZX0\W8&,!-; H<I9,&P05N9%K,!Y(')
PJ)KGG>*$PTQ_:3L[$-N@:RKE%%@$D5&2E3I[EV#:)D)/@+2S6I7K8Q8PA\K<&6-S
P\<;J#AN*@MWTF7!6QZ?;KE#C?A9(KN!2RLGV/P%.B[_]*5]>Z&B77M$0'984F^B]
PV6)RK(D0$%\6B^<W]$"&XFN3!CZ?.I2P%%MV@5_&'RU#R<0J$5&V'G.SZCT.G4D'
P!86NFQNM4]@S2MOIA , @C1-'?AGQ:527%EOP_A-]@E8^MD!1?EDPCHUZZ -^ 1"
PX*A/_P1L V3):L&>N'>.8BUE_Q ]E$^Y<X<;_V?TS&V,T[VMT +C8I).D%WDJQ6,
P2MOA^C@VL,&V9K@%AR>:*"59L2#IG^FIH/B8>.?-\8,V$1.-$!I_ CH.&:6V-7LB
PF0YX.V![B]07(HG#9C&&W=CW/B+APOD)(A#0Y!I"-1I-)<GJ)K@AGP9EH?:FY-?&
P/-_B:,J)0T_G;"D-]O]]<MR'!)<XLKK.ZDOM/-]5V6W\ZSI=@'@^S<[,0IEC4\11
PC54-_&R0_;29JC"=!04+F*IQYG8HQIEO@=U,F"IFA++<T'P4 CV'R7TK<U(KIK,7
P44 ZA<E]V;F>L:XI]E$4YN//EPQWAMIBL.[F>&XGMZAH^YJ"8PX_K"0>.?1$;)V]
PD3AQ 3U_ *6R'?1'?$&^K< IKI!Q(10("<(H0B$QAX//8P-7A//K-8SLYAP!ER.Z
PO^$_14F=]('B*Y5D&($&AO'Q)*"M4DMQ4_TB.N.HBFI-U^1S'*9L53 $\JV*L)/[
PL=1:$V=^L^QID;\##A+,M:PBI[EM4VKAW;VK? X1'\7J*'X1Y.96IQ!$W//V\Z#S
P\)9;*U- R71>P/Q/.'J\,R)86GK+L5]U;#&<SE)4E@VJOB L<:H[7DI+KO'Q"SY9
P;WXAI)MJ@'0O*$@P'L2S?=='H=VOO$V)[J]VA--S3&OK4<#&4\R(;LM%'_XMQT&\
PBOY>6D$*\I#;EM>B%$UL^3EE@&3S$0H--O"LMOQ]5\IO$^H+$0F?K;_H?D RHL&T
P94]; 5^D+A+L_:09K3KNC;DB@*GB;4J#KR?),2M>ZPA#]<-E3&F)MI\1@&$'&GHM
PPY6LX\KH< ++9_:0G1EY"WE7Q;(IN&RO>3(5[7W#G=:4[QS3IMMBYFNBK(!7UM/A
P>,RIIV=1"AS_N8JO+(OF]*)XXI+OZ'JM*"@O[G9YOKF7DH4[%5#81F+U,<JI$"GS
P9>/QS9UP5PIOW\4,$B'[/:Y%"!56.KC>A/1Z&OKCA<)BT)?C-JK#=,V;;F 5N?$G
PZB_#@:\)6(M%$[_)'?73!G R2F,Z,#')D8<I3,=8A#(4LGR&GH #\"XAPQ:47& %
P,>Y%L0[07W@JEE.4=1FM?3R3VU2M!.W/D\4M^[P+RE\(+GN2B>RDMNAM"EG^00>2
PW&U:$IHN?K:X\.XWU=&Y7+&(*WC#RDS$5;&:-G(3!]N01&,TGTD78(MJIOVU]9@R
P2F2J,U04BN7.:M-<>"^3I0&U;2?KT-8O!&%V;F$2U%V4Y26VL2#\1($)[MK]5'DL
P[&D@K;  2$&P][W!UN/.M24!+K_R/L:4D,S7S5DCN FC,OE,EN32V+5AX:N37@(?
PG%/^'N5NJTFV)Y!0*9<;21%F[ OR(YU$4T./>KH9];D\>Y0%-GHM<\A(1/EX_0[5
P(U>_$LZ;!85?B.M=+]9WT^)7 &)N<BU14T*5G$(V!R T0C^[D4O[G8INJZ:F)(_M
P5?_?S\P'17LC@E/XFW"9=]LQ[1J=Q,0(>M=]'O9Z%G9G^6L:[@N!282!(*&)2"5R
P[U"FU#!=!!_/DL,MKE(8;;AO<T,L#ZK/N>&RY@,$NZCNR4:(\ S9EV^Y%AUU;DE:
P4ZK.=#&_.IVX64VT]$I;B+](JI;N*\.64/V(-HRU9ZE9>8ZUS&/>K6?NH\/YYX=S
P--H0!@YI3/Z<&4^W)Y*<NMO^\X##G/T5IY"=BWQQM,]4UK^#&T4P,Q&*L1/[>O47
P5*.?*D!QM<&UYB-[]<X'2I(\:?DK8V5/,*YJ:0,@%DAPLX^:%BE,7X1,O ^!97, 
PF1^J((NGSNB@K3--<NW_;&.HA"AOK%@%JOV[X(8GL&2^[8T/ '"X&]Y@OD+3.D7F
PU=B6W\,M<E89>(&P6'7^I_7M)8K#@^;)Q"C0&'\RZB,[6][$D\A]/BD\TSJ8R^6V
PNMPNG?!&@FE]L2S-U$"9Q3F-U0;Y4RCAEU*1RR!WTX\=80>C8YHCZ>)K.P>_J7K6
P+%#-P!#0<\R,\(; $O4:D%;BNK6DV$YCYS; DP^R?&(]$+YL>*@XD"1369D&?F)5
P'=K-=FO/ME349W)CM49*52O(<;?V:+8IREI.S30)..5-=>V<9B$^^'481/FS=!##
P3C>Z6N0.:6>)2MQ\94N\P5!.M,A)I*(?O-34S(TS#CLT \FR/+;+\B/6\(C5,=P;
P2E0MX#QJY6YF:L]7WB-2!,,<-.0;R ]G3E+2A.M0*I'(VQP KI$"_TV"_#4!HBH]
P^J&."@_'P6DBD.J4D8;+[3,Z1);H(/R5/;HT!W7\@&KZ><-0SF-! J:Q-!2K?S%7
P@9L?1SQ>D,Q8EH"O.X#WL"C?'9+):/:]=W,>0M0 "0_NA_'%%RS&^V"KXB_N@(=*
P_6<.5***9,K!'DR_7+H2ZQ2EG%%]+W K8_E1'F1/A3'@\AG:ZRSWHCFNZ2KJ"E>\
P8C4BZ!108?_2LT_M=EZ$-!ZF%)@UW8BK6X FI+HD$9$BP QH(CX4S"EI!8GLQW,]
P6_Z=C?Z[+#NN3L5EJ)?WOJAL=E+-$"L2P[1]7\$Q.8-PU%0C<<FA_5+4:5A2I'9>
PA"F)3WT $+SPNCBDB:USNK4B2_F;KN8[^0LB=G#\K$ J']84?%FF4ZYO\;G ->$B
PO&9. DB59X-T!19_,A[G41PDY%J=]$+VCOQF]B9Y_KB'P9&>[_*=[AE-HM#^JW:E
P^E^'8Y:[ OTSXR5C(D+7-ZI ZJ"?*<V=,=QP<KUP2:OI_6+/W#."M!F9#G2CXC,0
P_B,E_257^ZJC&M\N/C@(M9A&)K'W%#:A&+2+6,+OBD-[ K/ 74(? ,SFMX[URH,H
P*FP\%GB#DB[M>:.00  ?>SCVM'=7^S1^X/I+(M(KOJY]?(&YK2X56I$FV;G ?SL\
P *E#>$/>'BE!$=6 )-A\>5[9LI&L>D^+^#8++K\KUJN%3JA3I.PK?9A?V:N36QTI
P>#/#$M/XO!4(!H1D;Z0/BU$CHSL[V%W!SXS/SJPQ"08RO#UJ??GUS'MN3=SYK43Y
PX\VVL-_E3#9<05T$>?1O[MT&4J' <_N_[AS;?^8+HW?P&]A >R;D4ZY5O]ZS HD'
PK86'@1.%F<:7>J6:REQ)YF[GJ\L.EKM,@:+HZJX.-VP<8*:AA,L=JO[2<<BK'Q@7
P;[IC_R(DG=2@U%)+5)S%+<N0Y],^5*);$;I8%!RL=1H5X-+Q;/3U B#%;F#3'LGN
P<A"+,9V&&47 /M>$F,2\T%4K'6,Q[\$@]4ZKX'PR6.'(PG.I/GMI(9N^?<@M<'M&
P/+07>)U:SM!Q#4O+,IMLU?<8 #A#-J0U#8:2U\VTX9IF#1#^59L/8=7M.DM$T,_E
P_@[+8-A)![40S4;&Y$0*#]++K4D.:!M]?T>1,<7CC1_<CQ<'1LL)Y#2FWU>Q-'%K
P6<N.F!I GF+(3=KJKBS_H=NR65PAD5,G"3<$ =Y:_M>HMSPB&K?8EQ&,"AU6KTHJ
P.U#>P@&E(#@WB]2KX1OAP6'\YL9XDJ33?+8\PLF& M+#*2+X?\4E^86+[OVTG-!M
PBA^2W1S%&:6NMXF]J*7R$5[F?>E&H.*;-2W+"JGA\!CB%W*TM9.TXO;^\![N<1F?
P%CXQN$RRXEK%>YW_5Q&H:1+\7BSBX%IK^H97B_\=[(#EV 77]>-F!&-6/9=Q4D9W
P2<5^P<B\AJZ>=_4XOV%"ONT+OJ#T_AIAXG\BM45@I'O&"-0 5] T[%$$'ABK[5J:
P>M.&!&+)#@2*[+1G^4ONMEKW8"[T9@[T-9MQ$YM<.]*>2!,)>F1MR,[9"-CZ-^T3
P#1>U06Y4)UEA:@H43H3WV_7?'/EQ58GX$]WG=_.873VCQQ+J5SH_OQ1ZT73RVA1[
PB/EIT]E$>P>#Z,8FU0[=.^]?7\18@N+YX=T87ERJ>'PM\[ :=!>KTG!*#4B+,RWJ
PK:BK#P9Q4(4$X\_1J3-HX4,C3V:*^3J/?T=:P$(S/?]4-'<?!?ORYX03X4HZHD?"
P5OG3$'\=X\.#1$#SMO:#>""1T]8Q.8IVLMCD8!^0!7?<L<QS3((./J"_T3XX-@/$
PSAH2P;I">H+WWJBS\[:WTS*0\'HO24@.M4VKS$"!#P59-1@6UAG91\$YY6#XG3,G
PP+J,WP'(CTFO]@L12E-SUG1+T"=3SLI!BD42=1O0&"CJ^M01'[JN_64=JK;5<&VQ
P5VTC<'X7_F-%DIDNY%-6Z4 RN?E 1T/3&03M"#+Z>'KDP6F?M0..<N@<@O39WR*:
P] /X <H=$Z3H(*77%W2>6.[T2; H<[]4#^>^.3PMF9B9)M]7+LK%TKT6K6.%AC^1
P]<ECK[I.G'1UGEV1@5#^^='ZJKUUF]YJJ.^P-8ED'P@8*UMS(_T %$BS+;WINTB:
P$A#\SNJ]%%GEHVZ .6&&*76+&$\(C1L4OS<,!IO,I8:L$-DB@AFX.?_ -<69R!'Y
PO3FXB/ZYG Y2'0ZW'B>@/] 3F7-]@<HK^%@Z_%9#T==K$ :ZZ/E?6 1@U5:(AX4P
P1%A>3&0#V8&%Y!V+<,?FKP96G02^DK*UGS)<#=\+-0\;X9R>5]6;'?]9$2,_0KI^
PK@,E1;_,FO?,.:+9YDSK..AQ>.Z;T"JT9U-ZYBA1]&5V2R8V7FJP_:>T*40D:)=H
P582/BAV+S-N5WA*U7XQ HVSI+9<AC;O;'L9*K#4)-@[=;2JH:L+@'KCF,RQ<,VXK
P!284FN6H5PM0Q\',NM9W;-X'4.T'/'S@A#'*4Y#5';WNR.8B:JHL3?O)P4B(9I!'
PE5-S"(C6^?S?+F>\"[\OE[IIEUU81GYQ>[=+-P4L!&*+.[+)%F> *4:GE:5RK.OI
PL,^*)"UID'=@C5 B)/C&K:07?[SZ,FW[LRL:H*UR.E6W_XXJQ&I\$O<J#/$(D.Z<
P??6: R?FPJSF-HU39V^[!F#\(2P6"_L1K4YY@@5L)WX!E:QCDQ&%#QFC"CLF1L,_
PN])\JI0^"Q_ER0IHN8K]$+2!AU6.,R0"(/#%2Q(("M=!6(?()>1&V<O-554DR??8
P4 3JL7 )# ?U$"2/VG-&9Q06:G'M_#(B:]G=&BL_($F5A->6<>-!(.ZJV6KETJJY
P_A8D*L]8E *O]%U@R+<(W5SC+6NW66U"'&%-]L:R :,\_J*:I,MRBPCRKDQ._'N&
P9"X7GC6!B)6CI6XK!E[QAA!OQZ%+U?(B<=T)-5$VX5MD]1Y!5HS>(B2B7%C"K+J_
PUEFLFW*PRR_X8VY9>MS\I#%T4RIA :SZ%HGG[JAN]35@?QUS$.E)L1PWI3?0?_@)
P@/' *8:;O?SL4[NHJJ)FP=Y)]_VW =J(56A.1LZ*QH;6W":Y T:9VY;S11KI-*DG
P_'L[]A9ENPF1%B#C>M$W7D*I"L -8("&*,1\;9J7I0O2=-T#2#U,\1@VH5.=1GXM
P'3R\/QLY,+EKF$#\/Y"5^PYF3*2@&*C]=CN6:#3@G1\E2Q$IJG.AI/-"-"D[0-':
P0(D7#M=9IH<^IM"G$&,(<D+$V>N>61EO9,>_MF.QSOX/GN])!TY)%&=11I#O[%ZI
P=-2B9%&DT3(X$[T3GCL*=(T&;DAJ5OA2V,1FM>G2<9:F<G9,FE?:K@%3_<_13C!(
PE'<3P  4'V8=;V1ZQ9.9U3LO9O>H/6\76#I;KHUH/9=O22H>D&K@3[R3_P6+;Z8B
P@.B]S7>K_R"MX5>[Y"#1'!X+S%-%X+\8O=WHY[,.[=.G'CM0O.U0ZO&7,*A*F^]<
P*TVU9<?%6&3)'5[::M\&2S)QIG4*I49R&',\$! K51+#!F7B#2B4F;UX)G]]-OZ(
P5X7.:Q7:@_V&-8(^_Z8*4K'G0<%.%*;!;E%S.'0B@]6)XTZ,L4[R,$)@YHSJ-D,J
P*&\!M-^"R!@$5#T'S)]98S?396SN#=?"NGQ#UI@H!-JJ7_V'/'H9^:CC1T<.N^5H
PB"-$5WBI:X&7V0M#J1BO$@&9L%Y38E6O%3"6R?)01S&QC*A%J.!T(3KE>7'LRI&X
P_7.YJ[B.^)G1W]+U_MUR<+'!H+^$SQP0.?$K)Q*C_(+EX@(-%98Y]6KZ:V=@'-8'
P?L*M(2JQM^M"Q+@R3VS+E+Y<^P1)(^7H!/G4.TWTB]7T1T%C=+W=Q[RKAK6U[']@
P/QN#*V72YF"1.5LD'M W*YD<K?"*3T8.:A./O@P[UV^R-)("E@U<=V0-_Y[< C%6
P])N03 4;#_LL'SRDN>P^-1B=(XB%YZ89%._\KAI!KWNG2! )N&)^P),7\X)H K#V
P"]K<4:AJ"!;OAH ;+B>GQVNJ3820?#ZI'1?%.V/?-%,'^IGP@CYV^E-M)X+W'9^[
POO=@?L(UQ#;- LC0J!'SK6J!%O4YL+A@7.2L$V8Q5PMWOQ0-J_161X1)?3V[0:Z1
P#27N?*F.#T1<4)7L#2Q5E"<<H 4W0!MK#T*K4LQ"DYRU_CY 84BP;##@/YI-KS>C
P_%]UF7/0\-$<:3*]EP0$NW-:20< <ON1N0!8._(<7CI3O/Q@QC"N)B8BR8:*\W]V
P"61!*239/#A@8/VH3H1SO2L?RH] 9IE"BYS@'+R5U1A^,,[E?/:I?TR'[(6I90P0
P/>R^%SI"O)A*(1G3V"?A*P(00_FQ&KAT+L?C!(C$BD-V,D@_:V9\VMG>7_80/7NH
P ;9VE*WPTHJ62V@VW(@9,Q>W OU">7PA2^D3P&AASM'0+.2+0/7?V0WD;\7X[O])
PT6N2_O4]"*&G&")(>_82,<!U'-@7]^E@<;X(;S:_^?)3W"K8'?K7TT[2W)DM*"9X
P94#(4W]F,:$&GMPE210>OPO> 104'AWIK@,^X"'!_<NV-/.L[4KSKI%T5(P2TL"H
P5%Y)L_-66@'C^?_8!OI#RQ\T1<!=Z'@U4EAR2W*H0^=2^8GFP7P&QMB]=C@YTZ$W
PI?64+FVG9RNW*4ZH*+8=-:3<873>@B3H+S- <&30_1*'HHD,XY39D$NS$5#V&HSS
P4ZP1PI>" \)/%DUW>2!W_(]@<AM^Q*->Z<,R!.7@3PFZ2(B[RUQ.MG%!%?698@#'
P-7K7+S!Y3_=<3=XRK7GK4.7YVI7T7Z?/ZBM<C;K!%@.>Q=IW%_@BJ$)TY5Y=U5X3
PX0;[WG<GD^K&#&/"X6".% &]'!X_*W4Y()^P0(OU#=K>W$7"7O7[*')W.=#SH^#C
P!%>J)&-2P=<KR0;'3M^KMZ&"Q;"GN?MA]=(V *1\"4Y<7?)_H5&VO\_*O"[$"L4R
P*+)C[GLQ?V/2=ETWAE/F*)B'LN@>A89Y*Z05MI=F>3U8-Z+)0AAMBBU.$H6D^Y H
P.9-)'DK=>NFO[P(^Y"XA L*??:?OG9C(UH-=Z4Y]%%>4'W-Y+:KO9TW]O@=\#-S5
PO_N?[ZBV8CZ!G\&W5HT2HZ_J;)".<WHYO>L^MR"L&CB-H\0+ !S7LU?DC;'3:]EB
PSD$*K*G>=9&P?ZDIFJ2.Q>)8M :!'2"\M%*!(IBL+4KSXJNNSL='3SJ9R5]A2?(4
PX$#$>G:1X8GH+O P,?Q37,%JM;+:QU[S#I^65VS%,L'W9_P5<)X27+6L^D7 AMF8
PX)P"/#(-3@,M;X1@*Q\)WH4UVXDXJG':IAVYTA4?:DQ(P[(91;UJ$7R1Y4_'0OH1
PM*O[4L:KKR@[P6% ZN26M9\2Z%[&6FBYR^[1<0<OGV#'A-118Q81 ?6GJRNFEJ\O
P5[N7@4)&5/3W;$?04C>I!-,<780NA_2[Z9X_6O8AXGRO4;%>SR]\?PZ"%O;\E:HY
PTC:DV\>C5@^Z"2\E-^_N)2"5'QN4@4JG@AY]#1MIM/$.J@F39 ;S]-!Z@R81T41R
P7!WL.@  O[MNV6YGJWBY5B]VW0D%J!YYT6@W_J'Q0)/0)D*XIQ7$_N^:QXK/@WGW
PNZ%?@9">\&[,1;QLV"[N BXQEV,=QJ4A#R.5G+?/?SBNY>4/" F+T$3M4H<1>"T3
P4DW@C%#*2YV-FM'(#D^UG:#%-ZB1Q3W D$HZZJ/9STQQ3(-L/],?Z&<XY3=D>F-4
P&8#:=,X#(\V@&)@>GIAV,V%CZ7822*!Y0_IX.JFGK1V)<WH-?O$T7",-5IPSL%<I
P%$,V,WPOKPA%(^ -Q.W1/6+7\E#:KVB=.1B =8D-2N!CEK08IT7D20@B)WU^H/PY
PI>(D4^3;>H=+21C=,*"4IF\'Y,R/&G05Q.\+/(>)0<56PF\+V0*4T:6.M(_IB8.M
PL$G%N5T@V^'8C72^HX_[-6'"HH W>^#-B-PP=^GKTB9I)5ZX6!\4=?CD^C8,>EXV
PU9E;3+"'BM9X0FDJ*7=,JXR?%1GI09$E\U'?#(A_VK06RR<\V5YDO<GR=V-*[/ED
P1VI+R'S+Q19)?\467RS,@"<:_KFK_)A9CU C RMNX#!B<<*<@#5M@JRAPL^9/4;W
PM-WAT,5&-"FJXR/QT/ \%KP# .0) [V@%Z"HNJI>YAJ'F!O!:K:N.1N23X78MGCQ
P?:OZ#.S?-T5_>ISL7#NDF[<Z'+3R"HO54E(B;XQ5!H/Q(B)GJ,0*>1*[!7$1'^[8
P"L*L$JFHQ268#%Q0IV)0Z%VA55;S*KPF*J/"\TW#1LJQF496GL[,/R8RYUO"@E:,
PM3*[C+E[#N@/4ZPJT)CG#7SV=443HS[CDHH<P\,VK O;3@7<#B:8-+-XD9V)$,PV
P0#F6KCL;LZ&-%V%GFF95U&CL]/*>3'-W,*&>_SJ6G8&':2HC=JR2&4/72:!(%[HM
PS0FA^P2#(?A?,"'N=]3_<B]Z<1VI0XR4+F+2>;.K4V.IAQ=Q#' .( ;!&1+WX=,Y
PEU/Z?YN2<6]Z6$[LB6?"V6=O4OD;5TP5=T&B?JRDOK*I)] M106%AOE9F:LD^(X%
P=+!<'S2E1[I[:#E7F!EM21XIQUBW&G88_2:U]D)82.I5^]NVSQZ3 Y.XN@I+P2?_
PCT.5=>A&4&70!<?I'@$^(JOB7CN6$[6P@BT$+1*D*GN/%;B(+=S!$5//R-P]U1Q@
P?5(=FJOA<1Q%'E.F\88>3F,($8&58#RJGQ'=9A5 FL-?B"Q]9IC'3Z9DU\FRN\K%
P49+@:>DT-&P7[-GEDF=C?=!6OEQG+UIBL4]D_,EWX97M):!$\,>BQBDE\S 56;!&
PX3;8BEUVKQH-I"^!=$(98(KZ#I 7.>;\J&:)^'5N)!VDT"[ >S\#LIUA+@/JX\("
PVO\WF6I(K-ZJ#]8K\8-\C& \$<2^$ +UF.@3)&%&"7T35E#6TQ*-N1>=JAR-+6T!
PO./>/5UF@?8@/XF#7ME\:0'P]_4Q\<A<0]5W/H]DL/"4QWINL"HU$;H[>]6\T'4%
PI)ZD=YZC"\DRB( EI.L6F3?F,9@[A(77=(7!<JB[5#%E<Q*\4K;F"IN8A^()P2 6
PQQK16[#;R,0ME/]2KPZGM9#SCA;\.-]Y@ZH#9K&WBS,0M32DG0FI^*^>:@+WJ!*4
P3=9?O5DU&S04"9R@98$IGYS);%Y&M]:S%G:\OUV1E7:.(A)=7/O3 +8$EP;6TWG;
PG##RS%/IGD,<'>?! 13YO&;5NM,7?1_WIWFNHJZ# M (<C'=YD0U51X32' :BC@T
PGU=JJVY&8V["_L3P+R ]9AR9,EL)%G-IUGPZ4%WF0QN],RT??&=YBDFW7)PVX26]
P^+#ZU_BCF"<E/\)W\_UO<H_-4N[Q5,C,CT I:OD;4FZTY(_FYS%I24,YA&%"H8"2
PU'1F]IUSQM*6?GUA VQ"T#EZ..$YD0*^A)+R:&=OQQ4'KM0T6^V>< @=G2P^+( 5
PI<#8I/XC9<_ .,A#LT566F^5D_9B[XVVJV:]JO"*7N+;N,A'62@/89(,F>ZC#<WT
P$F[Z$.I-SR3I,Y?-M<&V@\(^W>(ME*6LO;(OAPCQ>NEE[GL@ *#BJ7M'Q=<RV;5O
P[KU1DVGD&=.],'7DN,$:GU;#X;X,?G^JSS(6Z$(-J"(XVW*K^R?TPIE=B4/2$T6*
P%'1WX[4YB5S6G"\*@JMFPY_0A4:P)8K16R#OE86=^"L Z64!:&_@ $#,: D?I#K5
P9:D2V9 _%?9"(#;D6@$9P(60*ONU"/D0=VB=;$9(<?P1AI^9)6@5I(S8->K-0VPZ
PVW$DNNIL6/Y%9W!RS7LB=I3L*:=F4*R;(U*$YLRPO" 2*1A$Z@+(7.(F06D@5TC!
P$-J5Z@:T)5(Y*<CSN\\YC8[R#8T.]NN#1@9*_I$?&Y1ZGJ YCB\0.#Z<VUC4'AH-
P<R,F'TQ])4S[,;?Y_O8F ==BDL((] 9;A)1\%:+41?5GI*^=;G%$?O%?(OX?K@@T
P@14!(/4$ZJ@Z^U\PQ],*.1H=3/Q0\-JX.821;9MXY;]NEM:-E,>"K?+^+FC .L0/
PHI(J(J1*5P&'Z@,QL15EK&GJW HV3Z!D"N146M QS-\#43[74%2-V!^<;1T]W0$8
P'2QY\ 3L]"X90+/!HW^F-YJ$_EL;T!LDOS,37<W!AT7-$KSC\'.2K<@U3J5^\<&I
P'QJ]GXKU)"1@%<<Q+T551RIZ_XAN#@MFAWL\C[W[0 440,0ZM#6U4>(QK1"D]8<:
P$9M4XJLR2I+A!WQ).:LQ6"?%[QEC;@I/.!M+)M(**/KBD[/+$@@?4"YHU7!S]S4L
P@*AZ'KIAZCMRTG:F]".ZSLJ$6(/R^-\^>7'!1I]OW?^Y#BJ;RQC $$6P48;+Q<H&
PS*I"L7:-M9,E<FZ*D#*L\7:<WCP,KV$QQYWF%4K4QOVOYBOQ=LRIW$1[2TB: KN$
PBM3S1M*,_7:SEK;2<L<:.%K1]Q^0"Y]5IIE-J>8M5>F,[V\/D'UFYT[P@T%AN!/I
P]:G&^\UAG!_7S5I*/BE9Y:,F*\SJTX=5X4M2&+-&WR#/,X-:=-88VS>6KL&P)QT2
P2'L):7_BVK [!%$HD*Y4C@\Q<E#(3<!XY4[SM0O.E*90GW4<V\$W*)%=C($(\A[]
P9]+"X.SPUW1R4WZ@$53-1OG])YNA06K5)^D^+XD"$[\@ Z*D_&:I]Y+&$A?(5N&W
P^(3;7(+H"D8RI<AWX))"W\@-Y84Y_+H:&ZV^_^:NT>OY9$^$^2]<$%M:,4"/C_S.
P<>ILHF:=>>C]5, PW!,YH&=.XB@)).'[ED!\&3EC]5W[^_M9SO6M$";HNRCP-,93
P92:VT#0A>O'7"9J&%\KKJ,LB4G:^H=5PLDTS ;C$:\6)5P6M6SR6Q:_([WJ1E,!Z
PJPL0W]Q!"I]\.%6VB-SE.UHI:UH)>WAOY._HO" "MI0G03?O+=G+8=_'K_"(U^: 
P-W<_-?;:.#"VCM5BG1-&R1S&T-/%FD;+/:'6M81E#H(2]-]SRU%]G5AEV146S3'J
P-&NYXE3 [Z/PN<'+?(EE@@E-!NWY"Y_0N18;G);_"(0R; 4TY,[#P@YT >4!&RW0
P=FH']Q.%6RA9?Q ;#<1?'#SS#=22LW$QIE0BKA[WS=WM^S/W3I/;PA4]C/EB]%L0
P[Q-X9"T;#%\)]UR:EBF[C:%3QU;98:?+<RC$T=AOV&I\!OG0,1(]SYSI7<"ZB7 [
PP6)W(:B-=CD&O8Z'%S7EP:P%QMS\-S,%00L&!\(6 ZGGFW!1K,(0;VZP-;4.Y='B
P(]4^" 3IW;R,OH%'\#J132#0C6]_JJ%P%3Z0L3\5/,Z.B[IL9I=LMLD4E;O;)VXJ
P-*"S"M$5#-"%=P>+Q_T&!:Q+W!M"]S)74L!RJF@2DS62%%E!DQM$!<!8A6O>!?+/
P__!\LLSJ?,^PRB[EOBL"%R5@I5*!QQ]X0T&T?)0]\8XB=4HC"V )K*6BL56WI^UE
P/_MTD24NRVVKCHO(D22H@4_EDH0Q+KQ/Q%6F5DB&B=/-@6"^Z*8SZ2F8^:<LUT8K
P'A& LS>"1.62">P@)O!D=&00JRBS/#6LZE&\54=%38NY,>2DD.TI1?]GQG;[%@>C
P_'_+'W0W#%O1D-/?00\.CDG#)+@0W[7T37_!,-L<J,#%O[-.OZMEXKC63W:,4E7'
P DTT,<&R:M4GT9+OUHOMO 4B$NP1L)>NJ:6*T8R%O;E=IOX&-D_:BX20[B5?L#_O
PAE".[=\4V@8/Q0UJ*D"&7GN-!N:5W,LW=^+<"MG>FO?U#]4Y0O8 =<LYZGQ7QOJQ
P.--8R\6G8$9"5]2Z:J[V)])>TK#'Y^F%$M+RG4U+ 8NW%IE1\.Z"&O-Z!YQ=LKB;
P1DVNJ$Q'NVC>JQ4?5W "0C@O&"(6]0SZ>!KVKH)E7>0$4?:@91A5?7".8#5-I"RU
PJ6Q"ZA_O6D21/#'.0E7JN")FQ 012O#T)]H.B8S)8.?[!$(ZZ%HU!Y;C.EZ2@%L?
P"[ 3M.A)26P[NEB"FY1]U9(AFCG#,$ W?2N3[H+ITO6@^%S3UP4FCE>F:NLU0;+(
P'2[@VS#-92F9,@&SIHC!.XLY3&PZB/OO]922+L\'R+/VBOM\N\30GOM5=.)<:TQP
P%P/>&)(XTHTG2ISP@E1\;-FP"AQ7K(0=,3F,*(\WKXTPOQ,3U&/6/0%"@/V30WCA
PI%;EF?C(IR'#A?$]%>STM2XJ3<8.CKE6WO]6*"3XKWD0Z?W511:F1D&)>])6F]0X
P&AH+7&+0#\U^5JH)YU]DVD?ZVB( >+[7FFBAA=TLQ(0LGEB\6W8M(*@@ 9K5^Y[I
P2BO7 ]T4KGX2C-1H\A>7'R$X13>W"73J 'F9<A6?>[]=QXVET2T*#R.;I5JO,U&W
P%/0CT^PLVJA\"$/)_]"HXFKNW@\S\:W$.QW%<!2$VE^A8L$4/8+:'[MEGI1[-0YT
PCJ6[\&K&$.K"*?5&])#*X1J, >GG_!6K&GOE%K6F6YVPB]A+Q4[,G7-):,\6/Q-#
P#K_T;CFS9(0$D,E(:7^\7*,T6%\3CL;:^T8)(<5E;$ZG,;JI-I4N888D 660?LO4
PGI%#O&HX.6\4K8+A5:@B.?*C0[I!]*M5X0U_X*+G +X&W,3 (K!NRVP/E]K(HB.J
PO\MM6XCNQ>K=@EY'  J]$3*BGDQO8)>I@99@[--?<38KTD>Q_E_8R#$7LGS^6P%0
P+JSNVM[8_EDD#F770;9[(1!!\9*K#[<)HV@OX-F1%BN Z7,T3:YKT#_Y\["$X=C^
P>R.[Z,)P*XF.E;A2V!S--#3&,"D&+D)^:5YF'"83+'+(#ITY!^K?%T5Z3W>FVR:M
PM8Q:B<-BW+!@=F+:P$[3DIXE>ME"':G*?7_1YQ,]#N^T*>= 54"$FE9Q'#>"XF9G
PT;+4O7,:[FYO%;N6Q8-R7&K$2CK=GRSL4<*"Y9.C,O'5@_I'S,GY53ZP],H[JR1%
PDZZR*%;A.Z+<%[4!*%$<@<9.IPCUM="WWQ/J9&>[?46@&<GB\!67#>0A)92#V[E;
PDM1ZO&*>?T7+AB.5G-L^PNZ\TET_='2X>[AX^4#]O;Q"PR\W-6CDZ7J74ZZXH,</
P9 N:P>/3DD16)4%"10E('N>RU0@N,39CLQZ'1;>N*%Q%9[0*R8[$7E+Z@>QT33"L
PK8<M3*K*2"3F_]]XQ!PIT2IO0+X5R[)-YW.U29TFYR+73[,^_]RR+E0N/KFY$S:P
P!(5PFN"-Q\EV<WNJ8V*84'D#<,C%D4$ !F$NX=L,62P]KP_!.)UL6W(=LGGJVXT(
PP%0_+YWI#^2V?:!_%6'7YXS2B3?0V?)=!K#=N9XK;N:S]2H?E^'PP(7]F7AL=B]V
PW!OB4ZQ/GOBJ8;,PB_*_UWWHN^HS&M.U]XPFBSD_X%IYF8?SD5X@+#F.O14%OLO6
P.VNE]/V'Z,]><J+(_[O+,!@5L]*W.)=QCHO7 F8^>"JLY*?@9$*5KKWU"'\&"P 3
P2G>,*<7\Y-OQF%)L?-7;.Y9[PAHG]2*R#]@*)7C&-HG+B/L$.@&:DHB(!B#(W-B.
PB.$[=976P=9N[FA?/D$8B/#4@RR\H*[T0T7?1T?IN+0+SQC]P8Z=3T^U>.*[Y)'>
PUJH!@O*Q?/H$= I03PIC"4\2+T_AA*L1XO+QOTL]*;E&C4C98>AOW *WE0_O[4KZ
PN&*^_/,R*0DJX1##0_R?X+9\8QC%3W\Z&[(CHUN[8@(1@X%#\FT;,SY"9G@]QK>/
P[?U\>@59(,%\POECEML8MXLR ,<5^%BU=WHQI')>C@@\>4S'%F2R&9C,MVL\^H$^
PG(=-#<OGQ<'K"\T(=>A.:L<1?UQ88:8PS@EY85<.<*+E'8L,4<$<%W3 'L]1U<$E
PU-'L@ORHKOT_-U7,<%E;TB$0,[[ OQ@SX>]?)';Q9+Z\O[HE?T$NT(%]]&L2FU7_
PZOOCH!SEO+9HN"45\^0-@/7KD/I(=KS->V'/S"TQ@0#"4.)F26&EFMLK;X@KE556
PW3^C!-TN/("JYH(=7+]HCZVA?0LE*2P=Z\\*]+?0/NOZE*UMA93E+04/W?I4=L/N
PUDE_G=)?ZGKJXA<(;-))(G @HN"!::3<K11R VQ"75ME4XVD+\^Z4_[8BLI7?0:C
PK2#+?$:D-QEEF0B]_VH-/-BGZ?>(,XMV_B^9"E>,48LE:2@RJ-\=5+6U'Z>0\>SS
PA,AV%H@99,VBU5478V R*)ZW-_OVN3] Y_U8+0HI[LL6-H'-$U8I!V7KWVW/LH5#
PI65;G3_@<KLD4B*-'.N^$JX2<.V^,T$SSHT<,QNS]V(S,[4$H=-*A.(/I1>EE.M8
PN"69OS##TX:A)H3O)$MN(#-[TXW)0_&IX(H[949. Q'Y% :$^9I**=I=DP.'@LX-
PB7*M[FLY:%]TY->3TI/"X'N>Y.I+5VN&*5Q--L&IU&B>HY@\D PYS9IZ*#&_(<(9
PJT)\W':N<O(]NH\WVXVPQL8J9/.ZC?W5(4U2\6<,UE:AD=*9GK,5NHR9._^:USKY
P2,8;7PVO$H5>U/+]2ZG,E_8VKI7UNLN5]5@>CM1Y<G*B?@L6?AACX%FLE:IT<MEE
P(]8EM/9R>"-VJ* G5Z:,96FP=%.3\?YE]P&4KAJ(!+B#LHIPWUEK5MM?[1]LEEY^
P@"/DFE&M&A!8A3NOW>OS+^Q%<V]-@WA)\&TQ5F$L6S@NXF(*TT'^"]!.$L#4)4P=
P3 D+"+[&7,:J_RV#W";+B!;!4+AAS%F5J-2"-@BXX'=^JA/<30/$D"D^WHB\D-<M
P)ZFV[R,OH%?VMTO8H0.T^?1\4>LP@RNL-\K5/&S5MQF4GFV'8\G91CU*2UJ^V%73
P6()U^W$V ('XJJYMG.%*"OKA:0;VHOP/Y+;33<.7Q0.5E<D3 Q;KHU!M]RBOG($0
P@WOB+(,S&6 IM*2A("XXD$N"2F.=<N(%2?%F<GW#P05[V8QJQ%+1PM>5YZ#A'(5J
PMJC1I)>Z?I5.VV="LQA)?SF)Z*#WHG-<UQ3&T2BGL$*Y[P(<$A4CKUN-:9Y1[H-^
P[=9;H5 (I\L;EMD3@KC%=Q944AP,+1GWA'O$T/K?IF%JM3E]#7QD+)0CGE9B?CLU
P;=HVJH_#SE\T%S31D)[1\6:4WG'^KWJ]UQ1SBAQ^3"[ ]P37TJNHI.4HPE)@;H'W
P2'GT.ZA*/Q @U#\>)EE[DH*EMS/CN [S:&/TQ^\+$(^JZXM60V4X9WF%L!ZNHI=^
PC"',0^*"9V5+!B+A3D>)>>09 WY8(0<2"+-,%RFE,7WF_N3>^'::*]HD83TV$D6T
P9XR/'=&COC^\G/0-^X8?N6&G2JV9@V$!P&$#DI&$T"A<JV<-6PU*VC]@*'#!'9LB
PER4Q\(_7P2:_^&XQ!D^V_5]W\WR3T[AV$9@+9EWT98,_E"9#RQI4X-48("<* >^8
PT0N<<'&/GQJ8#T?/G]"G$_4&H'S/=JA$^J\$SLLXG/_IO)?L_XW@U>??-^HI:0.L
P5\($I%T#]@=7^2VI_.YT8+V.:ENW!BRWQT[%Z)"?']\V7.$]ZO?_@Z3X;)_:GF>R
P%GE5TBESB6J=T1=#<U 2Z!>O/0X@05U&9TH0M.;?8P^0$,6U!5XS"'\I"@SY,M?@
PV,=IG=J%D6Y0NOC@7I8(WJ/^^.0,,"5D(5#]/[$_^='EH(28&$R2RLB 9 KXM?72
P"#68MV,' #_7+0RQK#$X,)&B#Z3@_<Z<:>W&-VG!K8SQ-;/8EG.KVRZG-1.9JTL=
P<$(AG*1&* R)8]V446OSDO7JD'29+[$DH-9>:B/':L1?55_ .$;TQ3_<>7Q8I>>W
PE'UF01]?]S5::PD;2H)"CTPW%.PCN.88IGUQH>LB?8N!@E=3HLKT_JHDH<$ A[_B
PFT!_HZNW.][JSLOSG.H_CR&#-4<3;7HS11WPV,_CH@O1N'K%;4HYB: 9Q9>95?8I
P]-!#J?@(VAFVX4RZ/YNB 4]-4W'TX!\A^W$@DE* F)NOAC.)_HCF(J(+?W_1/G$L
PL-P(W,O8_NS:1VB0C(@VVLB0;MWN01/3/MH/'XD H9+%1QD5&B(\[%4=PH=,16VL
P=3*^&<$_;GJJW#R<;RK<UD(G@:<TG-/$8M_EX1!C9S0[!G&5HJPXC-:)AJ>*5X2(
P8[QE(#'M?9TDZ1#RW<;^FUZ(Z>[13%8^"=Y.9.2K8H3(G[?$K30=_!:S1CMKTDJ9
PHZ%_V:CPT33$):Z96+YCFE_]C+@C(0EWB((DKI^(>3WWOT\3F6PM+3D-6\B$!>YX
PH&^[*9F0:L-LE8L$&FW?SU?G=9-XT,@SE& @^V.I*?Y,]4SBO?U3BH?T>TNE^>MI
PAA:*^9Q@C5.\W.ZJ6Z ^WWWGN%:L_EPQ<\.-NIJNS;)W3]T4^032G:"+_&B,W(<+
P?W"K[E>S$MD_$_,ZB D 7>RGN)IARPVZIW=G,</^TM3C6G6A9#QJCQL%%<Y8V,WW
PW0P";5STH,"3JSLTTZB07]'\5A)K?6 I/_G]@?JL61ZN(7,A#'T>$_K,^J%+>M".
PM)]3@:IPAKK"]PZM(WQUQ=B\V6!YL.FOR@3'V=S%)=3 XE\N1A.JY5F[+!E#2!.=
P:KE\426)-AJ9\72XG<:[]@C8=VLN]W Z0[\7,? L<J;MR\LU*5 M95?ON0NTMD_!
PI-B?1A7]S7I_VSK86[V'_.PV6^XBGE L_T<K-!RBPN)7O08RXXJ(JJRFZ/50,.;/
PYSUVB"-!_U4J6$)&OB=<X@Z1 B]$KHRW'VZM(%1CD>IM2;U@#-HD@,_$ $0/+?$3
PVGN]$'5W&OE+U:#-7DMQCL@B*;,[<A #\[" Q/$5.>--LX%BR@(ZSC,IZ&>%:A0A
P/TCFF]],U0BUX6NJ.7P=XH31?Q"]#LK1&.V&N[K"?*Z6\=6*Z:%>A#^TI+X.ETAN
PIVM +*^/LJ B--$>24M-Q6CD.6T#%J;J6ZS; R0(+T^7G:H^FAY].]1H'5R[#@!.
P5>DL5B<G.)QPMRT0UG!=02>P3S'.IC=;6N0LJ99S;:;<V,.*!;MB&D@]0W9"G^U%
P/_2?S(MLRC7G^/'1)F&S>?N97^GX?6M9L00V3Q5:Y_?"]0]+?V?E3A-IZ/0'^ZN 
P'J&< ;JU6$<&N^8JMK&,?&*7S?=JV7W!T019^*_ 00P)1%'YNW[XQ#Z5VE KV4?-
P-R' LT30&U>"H=J$N" <A#BO;:I.C3(&8^*N7V09^?ZHMLV;8J!BKU(W)Z]?;6K>
P+;Y'O7E"=^RI3Z44G*6?2FUN1SP6L*.'?;V1DZ6:,HY/_$TD!4C__"*)(Q2A\3K.
P^O&=97%_!P:KQT%Z#Q&GG1 $L,TH-U4$PV8=.2XB858-0CH]FV\!7)8+B+8(E@.8
P@/>ROY'"'T1]/N'Y1VZX*C<3N'X5%A\7;#S4@0S/)CO!C8UKO\.?>X7^2_(C4&&9
P2'8H&H![_,B$,KNUGQ'E0JI !:>@>M@U\*W'5?-;3R%[3?)L,6+^6>-]D6B&J::2
P2(/$K/X^NG-5=<F!>K7S#US%<SU3@X!0U9\NHGQ3(5C6PB!;L7"3?.2Q!CM[,BY"
PI3Y:Q@0)Q](C_)&5;E\XT''ZB[UXF=W8)7K&:TDZ2$Z-^%?C X>S&ZF6>/W,BL@#
P,1?)F@'5\.TWZ.MHF_I:EWC0Q5FTUWU(>3<+Q[W:[XJPOZ;"]45RKFWBHBDF+DS*
PF.@A000N8?F;F;M_)TU9($&DIH0-O>19[BJNIPFBB??"P,<L"+9V=HN#F"4ZTN\R
PG$L/MD/ZE#,,HU$);&J*NJBF^G+4L_X5];'$QW+,/X)%_<7B=D]VZEJM =N#<6@R
PI;2/3P93D#-2+9_#69ZSA<:YK45R5\=.=Y]:<6:NNF@5=FJ=G*^BN5+B0R?28GWX
PYL=;3D]+ G=6>#1F[[&H!H"ZGS*KAJ6!J2="H]YA7'H9GH)]S2S\XP>#VTLLJJR)
P_K/VF^8A:Y^^-+*N $C6_,E3+A?1+-^N.*8VK-H ^*.YQ@W0G<40Y!F<@*W7MW[6
PN7!#,(]3-'B>T7K]"@$^+;)#?&5=:QY=0PA_E.EJPXE@!:4,$.K  SDT%TDUM61)
P8?^Y,-BRJM_/BM-;E2)ZI:S8ZY3.-F016M@P$TY^]UA":1CMS&!G!TB#QA^ I%)\
PRT=Z=4#W5:/9#]3P" 7ETH68V=T@M5=WL>!;INZ2Y<%]Z%@.1-/;I4=>2\PC"(FO
P_9!2YSA(KQV(^R-9$2&ZVMJN;=D[>8BNAW0(O@])D"2,KJ?&+ZZ.CB#? 4I3_.M.
PFWM6J!P&+*:EP,WR)*VK*E^'[HK\1<V2XC@'<81/7;Q[$NRBODW,IQ+%U$/UIB2@
P),EEK,@)@3K+EN:@' 8D #5!UK2/DRE=(D@FFTSR)*,^F_L7!$*6KR3-&++#Y?NX
PA?TX13ONV O65GQCB;/0PTB4WIK:!+ >HC&:L]5C=[_/$Q]/RQ??Z\O;ONO.RNYX
PR2+N)%X5IM\JQV=1>JI@2E!)#A'+)H[GSGJ8.[1"&2,]XH-4WCS2MP(E)KZ,^;=[
PM1]Y4=#L+/*6XS7";XLY06"HVV>X."0M\Y;7A5D3CT%CI!7$6YVU5;]"W!?0E&VS
PL#U--@M-GF\L \)<"';SJM\\.0/=;&I;<P("YG>VY0S,]$?'=#0)/SO=.9:<G)&\
P%6=P4)L)N%)8)8V<XZ[(2E<98-WU7U&SZWM<BUY/L\/5Z?_.&MW$W%HR<BUPY+6P
P&8NAN80,*?4!V!1UWF[%WB$-D5'3_GJ$QQKW>CY@GM&;BR&+Y!;XBR! OFM+8H"<
PCG%11$5UPH3+.T<"H)AQ;=,N6S8OTKP4FON6H38.GQQLT?\+GFXBS5>2]]/HS@LP
PAP +8% B-/HX_T!%0W/<+*%;!/\.V-&N?V9F+\E_M>NNT]J"X(YL7'&]F/!\O>?6
P;JX7N4Q.Q?C=_? RAEV2*.=7K#*@X <OR!+FU.A.YP#-F<;,!4\NNE"N0-EF<SCS
P&V"T@_!X4?Z)>48-6REQ1,J2!Z,VM69^_>J@RI==574<@PLXA21D/;,+?*D'TN.O
P80<LC^KX#6S9+2NLID'RHZ1A;A\^*C2X.(+:+O )\^J_9;VT6<&#U#PP7.(ZF*^7
P1HDQ])?4;P\-6I'24$G74EY1-L85_\^_]IH >[+^*^<"LIQ/>E-9W</Y=AP?2_VO
PO-N1[=?]F/ID;C=4#,:Z4F "@"(,?TQ+X8^H_?O.,M" ;'1\/'U'Q\M!RUQOQRQY
PCJ_B6081,OULF1WNQ6G3.3%D"T?LI/J!D3+>ZE1F3CBRG-11<9?CH '(=?SZIM9$
P(1];$Y1-R7RV(MRBI%!!'=>?QS2>NR1X@X<U!:D\RZY>9))F#)\81?%TS<V/QX&5
P6S044_R?5[2HG!-". D= \;;""HOJF6*<"[OSI)M1U3D2 EZ+:TY3SGC;4NCS51 
P=R74-)HU,N(L!C-:ZE,_A_'.:B._(:]KCNI%S;[=JU,WZCCG;P9&!@ ? U=?)YGU
P4H[OD(,X1$H("$_)8*]* J;BDF&$ >TT2R NIT@4ZFM4+@],/@ GUR;C,"+0'*3_
PZ8K7'M(]/MU;(RTM[Y=->F[Z/$=H;HU,13P!\0.F*OB\0:/G0Q!LI(AT3N^&OD*?
P0\X^012C>7:_#]U%YO!*>]^X4%F;[A>*U-<?$4I1_2PS#M;HM]-A7S_>Z]%8#CB=
P%<[$V#,8S)I.?RYQK[NS1F%CV2[H?$>_:QS=-5@>2%#AQ)^)]7_*V %_T_;BG#J:
PGM'O,NUO+,.0JL4>8]?3*<+&I$:/[I(?^)@D3C'9.6$+#XW% W+52UBM7;I+YHD!
P%VC27#T8IVHB72"[7D:=U!OZ02"S:%:QSF;NW@W(*J@C?\,(36I@R0!?=^3@_LDF
P@\^'/R*5D6P-#H33L!/D;I?5\K6)$%%IK[/->.2H*"2_B#[+U8E6"EDL^.6"(<5C
P=$7L#5>9:RD]OS:MUQC\5!AB;N.G)%TA_?3146FN!&6->#3^-Q#OY*16LYX@D"CN
P..[^X\'CV]!6J;-L]=>ER?PV<1+U<#-1IFI8C-J?4/1JKT<T!!\!,0RDN6Y7OG$W
P#(%UND*XOKE%KMJNWFRRVW!_O_(F<*'FQTRB\Y=W6R6:)8C03< LL?Z/!6G[*.LQ
P.X $ N! 2N?/)/"6*AE"8/WI.BY%=FO34T(D7XNVR<YX)N%(.I/YZ0J3;0"W;' E
PS $UDLQC320!ITQH/:2#$IEF7(643YDXP0@D4/[W08W(9+1H<::]Z8:"DLZU#A^>
P'9^/]OQ^V60=8&_A>X; C2<I(V>+\TN!?C<RE<L>JD(JHSYA%]Y6AX=]Z\XW17\Q
PKXIU]6[7)MZ9%L//6\KCO#W7Z2<?!T,?O9"R5?3@6_S+>QQ"XJ6BJCVV4Q08.%(>
P!;NTS#VI;-*S *]%;&-#?#YF9D^31](5^-#T&7-J1>(0:6G2R;M["<C!VPSO&9')
P!0'"!;&936?=Q\50=CF=,H^!Z!"'"[I<,+X4VI'13.=(QMU^3V?6G]BDCJ3D0MHK
PHC)[B8C+J0-P\Z(0PO.0+ %<D&&VGW,>]F(B"E+GA TUQ=-8A;:BD"LYG "0>,Y#
P?DV=LJ J_F-M"R1+%IL<E\<.\8-@WS]D)F?*<;_SBU?&#!4,41E_TCBLJ_D728(7
PB0HK_*]S2$?U.NS87H* <U4C,#'5A2HI9CS#)23Q\X, 8TYJ9ME+X?;LQXG,=*35
PE?J]T^3UK<ZMQ9WO9>]G0FS!"&:_$-AVEE&5=HPK0F?^.A"1ES,GN<WJ0NW'(A66
P(G5=6R(FB%H0Z!LTY'3M]U;U6<X?L.%</=+#GTZI@.HN2V>?B\8DUZ=S4F#SAN=]
PE:C;*>MB1Y[<?Y=(Q^GRX8QX$2Y/%EB^YA:YZF]. 9/WCUKX1=4#Q>E)QTK?/'5Y
POOT5_"4:MER;\CA-H:U=#V.3?1+*453.5542D,1$UDZ53G!<[_R]\.+\TOILKM6P
P-L"H 2JQ<OE\;V<G_;"%1GP"C5@ZR:[\<0/_E!#9K.[=?R&QSEPC\^PX6I\- \)^
PL#UU^:7?ZRZ+):.]@6\++O,7[//&ITIW?R-<%J$2] "*.%JCVQB\<EH_'\9I6R+$
P[57$XLM1NQY&^+0>Q?CNK50SSD/A,D:K>%EHP.O9:TNK:4M)CS(31!49D*7*=,'Z
P)4/@K9&,J\)E14GU"6A?M91^LG QI%:=<R[<8'(*H?'QK_&6&KS-\./K_?=_>VJ/
P3V14;,7U[\&X\*3.350D25/$!6BRF@0ARY[ZU+%N^Q"6K") ^5O1'UNQ;FL"F46U
P_=&XPTY:\HO1L:J35>J?_>R8??%&UX,B/*MI[6[PGA",#4A5HA&@&BAT>7"6?U3L
P 8TBX$IJ3I&(!8+;BF(S[]OF60=Z$VBN.W5#PKDJA9Q&]S/_,='09D:I3'^7'')G
P'AAN[>ZSI%]!YG+>L8Q'!V)0KD.+$H-FN2H!HEQCA9H^'ZU!<$,UYST-_5 RD_H#
PF-(U1%%DP="L*B9[=$Y@O.$XA..!^T53<H#ZRN?QN=VY\Y=5@+LTT)-U4 I'/": 
P@*Q DU&[N# M1(79CL&?(P6O&PQ>T;'(52+Z!L,YD[8/_MG@B1GCA& G0IE0TB;2
P_$B;!H\?(QK\[QQSV?;K*/T =(;NSJBTV3R7%UR!"W]LTP96<P0L)'W '7LBII0<
P*JTV,'TT#DY<HFZ>(\[D93]CZ])Q%%:)C/.E:?)Q]V?'Q >S/]'.\PJ_WX0:I:0%
P48EU[I//-EM=-W^(TZURHS7>SROALX&U=0\(&XD08KZBJE^S*>25>$MSHK!:BO!T
PX7(EC/&;]POS/<AQ,.4!I3T="-A./P,\WZA<AL"1S[/P\M%_9/5I'0L?>B%M3E"X
PW,P8 A_MG4_%CDC&[R4%S\5%?O=@>6GIK8Q0T?PE%7Y-\U"KKRG2 R'HIH&F8*UM
PK_ALO=_\L*DYI;/:2G7/99^KLJ,W++S)]Q?749H_$>WP>MS>-1)K5:D;#?ZROGK1
P2%@WV'D]K4H-0/NK36N"UYF?0 :9&L6/.GB;SYVC*3G3XJUM$9TXH-P"'E.N>,>5
P)"J?=/RA*J =I[P)ZT&8HE@YG9?E,@#_60^K'M6\3^;][2"ST L6^)>Y-_+-&QK!
P@"!B(7+5U-5X#&.M[261N\B^X>")^6H/<_*I P?]E@,Y(9!!X)_JV*FT\9V"13\3
P.4JPIDIT'J$H61NQS_.L@&SVIL<+B4,XBK6OLE>KE*F;_](V?8,&-9\%C?=X[8:_
P#G<,O+I/O8@<7\E+D_%E\W[B_!V+%\4 *YD31\[\$I;HFHZ108IW['H ,0B$("UX
PC5O@D[C6Z-P3OX@8%@WS:/$33]D-BT'?.R$*N!JMV92@2HW?0N$SJ<,V_/SXONY&
P,_@=X:M#Q J_5J%F"@SQJO+F5ZL^)\$V\D%'GH@>)#]Y(-/WQ,_D1'9D#W!$'BS6
PHV39AW+7?>T#(CBN"L\4[B6Z/GV=KH8DG\5_Q3V/$1Q3 7>G="ZJW)^M$,(OA>*W
P7S#W54[M1K'.0.S"<GN.*)! ,_.8[5.W)X7PS]0O)@4E?I^L_6JR"W@G4;F38&V 
P-348^2AD4^3.?<]O=7 K)<S"P%G@_K!M]L;7>'M5:%SBA>?V(Q=B&-H\<M;#:ME6
PJ00B=8U&1P+T5I'"_^MR>UC(KAR*A$JT12^CN/+>1<NGUX3Y@D>#9+_(9W@ NX,D
P1TN7D'[\Y?(ZP5+;H,L(R30&;K%CF3BN72(_RD19$,^EDHW77\^'OJF;,,6P.FF@
P>: _OI7 6AQ?$7T^-1CHST>GSKZO O/S'8YCGIMFI:0=V#'-E:XZ>PA3(XC*9.U"
PX+O+1_U>RC7%4S,'PCP\#W>;EZ(T'/5*H-V&#^@ID\Y+-?S>5'@&&177(TG'D5\U
PB\]N%=-#QSPW*O+M!'UBT+G9KG60@Z)Q]72+9I'G5RHD4LNU(E'K/-1![!C ]\E*
P\X%JL<D$4>,]W_[%+CH.7.$O0#GU>))+C&MPP*(-'6(DE#2M4'1YQX<?/M9A1MER
P=_X9.IMT#!^/U6#SAUL@)]NGUMA-7DZSXZ^:V0ZQLG(B$ '0I($3R\$0<Q=-#0;)
P.;8@M5TJX\S]RA'H\</' F4T?RE9CM[VV$606_QED4?:,2)WM-)A[@%E5V6O6IS3
P/)A! ___2P+V?7/L-H@_U.CZ+>+H^FL<M'R[3_0U-%V'GJYO 6LB17#P(<"GO\LM
PC8IR7LV^C0Z-P(>3"[#@7]2 '5OD[+\.D=W$AC$F!IWBB!4>5247G262@EI16=UI
P"^CB!8T;<^)4UHE$Z])SSH1  M.=-PE(ZYWV18R)C)Y.M*5\X;!9=KH*EU6\?:6J
P[[W.LM\_UUFC98ZQ8"XT_H!,8/:)R-=54)AS'@-88_,EY>\P'T:9W7;=5>,@5Q1.
PKOW^DE;M+4'3P?B5.%S-LWY.S;]$KX$.F;.,/)A*/F?RG)W38JI5()+Z:8\%XK,$
PQ9+**%$]<MW':PEVO\ZH$1=>]0@>[/"_!JV5>-ZX\L9&8_ HK0&?>0<2P4?Y9Q])
PR,KF:K%]APE++Q4NN$2XD1D#?J*X\1RL,PN-Q.7V$<3*#HSL.C-'PE _&YWK:>U@
PUMH1:@ Z4_<)=0R >\9_B,N!!^8;VXE#RJO6YN>W]_)6/^!U>C3[E1+=)!P%C"8S
PT;\=RS4<*S]=O[T4;_&5:+3C3&;WQJ%^*@UB(K:FE*\WZ)#@7HSS0O4?Z74;D^5V
P?4;]=*%8$)<7W#/I4 ;CJVSSUBV#6%^F&>9?)[U2$5-5&#?Z9@SU2SXYX3R1O M$
P:9(W- S,7$!2>=/Y2?-)36W&5%[!& 6[ALF[VJ>7G G/AH-.)B#[]>WM\9YM%04 
PA<_XU-((8R&@ ](<&DGE?0#"GR R*W[$T_^56BH;,=0(3CGCU]<$DRQ.^$9DLG:Y
P#$"&E%9BL*3BNY?P<MH"L9K*SS/7^5^E<6RFVS%N-9J#ARE+\NF)Z=[&4:!B.:;@
P9XKAO=?3XG^N:9YF*/^3)Z+FS ,"88)H=M/M+T=[\T;#[(Q[0_9N</[V#CEQ%FGP
PLF**VG2JP_N0=11EEY6=Y*UR)(_IBP#M29K;2&19A>04' D,A"FG*YZJQI,^>5=6
P) #V(JBH+MPP>IVDU(>I6'P6;\#7?2+T);CN+P^0,( W7!M8/.G^!+3@6&)9-\K*
PMWN+)!SANNQ4!*22T"Y$C'G4N[KKEC 8SSCF143O4,9DGKNK?-R\IZCNMPOW4KGW
PHF[RF+,F,-$0WY< C@0BBRY\%&Q(3V:#Z]MUC1D58*Z%>1D[GXRL]_F+GK/_PE1_
P7MKT JZYAWT!G6#8V D'18:9%K]A;H?EDAUQ0/6>6$QBGIZQEWE]KTBS:@C+,W5J
P60$:/\I#!]J/RC7J=YEEGN[EC QT(Z(:%O#(;/:%KLYW[ EBNR# )N35'G?*USF^
PV"^.4@D/UA[QWL2V]7M\(PJS5W3QH/1C>=FA7?<EL43:_9E^<+L=E(57KX6!9@!W
P2GV4-;(ETQ3WN72T?0AM!JEYQ &UAKW0KS ?B91ZU'4X+[)J??=Z0P$_,A[UAWR/
P^$60M\Q^2<V@1$NY!XPSJ/<9'$Q#(X!*97DZH9*_GH;*SR[Q,1X4.\;>ID,_*DB%
PN]424&%(RW8P3G(6J-A&B"1'D)K*$I./_I"N3WIYNJ'XC[T^/CY30>"#?@%>R)C0
PM>5&@^J18Y(*ZS1H22 XSO+0",&6(.LWBH%0UXP20*+T7O,G7IG1EX8<;[_9JD7.
P("/[RQ9J<H;4%!V#HUWYHR0T+2563/LU%Z61UT9L^Z$V3R&_(0'=F!M./(#;] 90
P'E\X#,C*P11"U%G'7\)XY>MT3SI ' QWX :$^4FE$,JU-+Y[<[=ZC[CV=."O;=,3
PBC[09QM$Q<J*G;27%!@ %7D[']&(.FF'A>PZO($9@=HC-.:/V^9)^FK0,\L +2.-
PZU&?+8P^(2NT3P'V!\<9]'2ALE(9<*T2%;3X28^#)[7XH TO!VXMT=_BE*1J0V!-
P$HI/O1WI/09HROIA\@!MDUB> 6HU"SL,6FG<3ZTHNLF!V*@$O:AP'8UM.:K=^"?0
P5%-,WQ^_]@1^RC'RF0..'I68#X6%)FWF:ZI(N6'RR"KEC>-+0S+,Y-2$,*2^7^MG
PCHQ9#_?H:"9E%[@*F/:^@PG2@O1F!,"GJ6]B!AA0G3@Z"DXL'AR?&4<SF0EP7JSF
P&<TA XQ$Q@GGDM#O4^_Q-.V94DVXGQ7_^(!6UP&%R->\/W;.D(:R2CD,PK&Q+CB#
PK50P4[;C+QZ&16#7N$]M&;*^O>!1Y0W+ IO,%%@QC!@?\TFK141O9QJ\*5B7UIJN
PUG$\PY!;E\F[XA"6 ^F_N]V^\+CJC'OP1)N8GH@TE'6CN)3WPZWAON5+%A20\AO!
P;0O\,EXWG/31PCD?:-F?MF.R1YPCE\KI5+_#H<\B4U'%Z\Y!B52?3>?Z%_?&YA/'
PM,P<\')[QADW2)#Q&F5U\*]BP7P.Z2];T8))V];C@13R?+VRMVU>?L2FU*UQ1 58
PZ!^2?N7$ZVI$UQXJ<89,S4.B<Z"SV1(#+0TP5YBE9!5%#63!L)+M 9UAFT)+ ^#-
PWRE. G>,'.=%ZLIU4/#B<!<?#-;)#1<[RAW73-A,AZU[^Y)H5BN.9S"E]4E$U"N)
P=<#?E6?^',#2.S)%H"F6A7TD@@ESAQ5E(1F(Y??GKQ>B?_&E/GVQ3L!Y?Z+*M-=:
PF=W>7?.M-^PQ9#'Q (=&81WATK O)O(84+G(9? K1KC"I5#0L ;.$MW@9_^Z+VA=
P. HA!\\E9%_(W>*Z=1H[:?Q6'S*'0OWL_M\RX!J<I%/&X3E:]J]M[?LB5^QF_Z"S
P^B\2FP+W9+9[W;)J? R*\IMA1!9*$E[8%98:C#/+S]Y'L+LKW-'8\9"=-QALM%EM
PJT3.GXEZMPPVP[+]'WBQ0,+>C(XWQM2GQDR7U%,:?4W;;ZC7^ID/'.YO6F'#8:=)
P$CN@.AU2I2U+123/O):LD,!?"\!2JYDCWJ9)O:VA(C:M_5!0UJ.1F;B,!ZRNK1=U
P5V>=.@\GA<*(A$7(KJ'^*&5;7DH(E-\\>EF?5.P63%1>ZP<O:\KIKVG/&+]-QET:
PW 7?NMPQ5$7K1GO8+"5TL0826 CNZ:/BKH&%N8HN08MJ'3["_O@',(6>F5'G!*@]
P),:$A<)=BJO*N5+9V/4P<!J7-K?%_^KJR9XF:XU&HZ;,_ZK+\-%T\0@2'C64ASV 
P'TT868QX[_J*]7S?N%X\K<;2"EXC2_$I=.R6<"Y1[X+<$D%+V.(PO=4R1(4?^7LT
PF$J^Z>8Y>LK3BZRV1_E2&Y\C+G1F>L_3/ M,O_T[229$X)H^L5P8X44STMT<'LVY
P& (D4%UQMXWA#,<K#Z1ND-;4J:.>-.,FQZZNS7-(1,,G97FK#5RXWZQ.]4E<0YRR
P?3G8,C$A'*!Z4ZA7/IL1A83997\M5];B.2"JC.>T9]4N',;'\.$:)';.D10T6N]-
P/M$P=^0+*5A T9 #8O)Y]^#6Y0\S.QM0E62A85CC#O;PF\=V9V,K'TPH+VS9*Y 0
P(T]H Y?=M8Q5UQHSH;H]5\9)#<CM:)^.,^>%0LC>AQ;G;X*!,GL<"3K#T5R&KJ''
P79N&!>"YNMV0<V[\QMN(TI^*53VVU"8E]"ITAX"7\VDN/>MX9YX39W%%6&)*.&]6
PV35^':S/A%H?NVY1S].7.GPB-0,52,9R9@AXP)/ .-K6$)Q&"1O&Z+:/@APM'YNX
P9=6W 5')XT/*E#VQH(=Y4BIR!R#C@ PL@KL/G("1S(2Z5=BA\0L,HB)HC62">MDQ
PTX'0'2H \W-PLE.&K>F'5HXE#E+5X06^6O%]P6XUGZ,UUR?[OY*,#!U[Q[Z;U<";
P6(-V7Z<*W'J>*XO(O%]8E<\,^76]9XD/ZFL\ \_:"$9>\$H@<$*JWF!E7#S:R>(;
P,!O.F3"6.196:&&Y13YJMAR*%FTT)D4\?8VB AT)CI-/0['#,E^ 19JGVX7 9I/W
PQMGTSO."LE7.2#C]0W"S:*L"&FS&=7]-&XR!=791 ,6B*^6AC!,^?Z?0$,[Z14_P
P^P]L9D6SO4Y?G]9!?Z?.\]8M[N@DVCW'J-XE*KGB,>-.7*T#%H8OIXEK&TYG50/%
PM,]>)SP]>NI!O4MX.DPA?L9J_?,-\>QD;(^MNZ$IA-\&M,A:224S<.%$R,<Q[/0A
PE<7[D>%RP6H^+:QV"CGZ/!6G5.&LU1Y1Y&5I!8GTF:Z?F*W9(11VGDPW9@2YEJ@3
P'(RV._63H]ZOBVD'[_ <R5&[(V03Q*WCUQLBK7["J& LU4P*2DQ;@FT&?'[="!"9
PPNIR&O3RIJ+.\[2T$[40[XI](QDS04X=@W8YBK#*9,N?IJK)%#)VKQM$) 1<&D^"
P^%VH7E]L=MS59'<L=B*7]VI73FP#'4Y_\%VH02ND2_G;;C;U<!=NA ,FAK>B,CVT
PE,9G]7 Q2Q@JE+B@!#,HG;%3R#]3DYLM74.@;Q](355S_,],F)PN&9B;F2P>_^(%
P'H,71T$#.MF&E/,PK2SB2U*&^(MD%SM+ ;3B0++I->J;]XV G?7.H/E -0$.;]P6
P7/JT O&I/3;D[HZ.(>.;3K#]S@VFORF-JFFW)L8W?V\D=P"EYF#[^Q\,=VG@+(&+
P4\ ,==@Z=K-P4UQ,$MH(P)%3&2?^!2:(LUJB@#[X<<<P*&G]4C6B>=TY\[9$[ @H
P 8.%<4MC/81.CS<2;2;UC&B-N;G8&C%C3P8TJ0T$' ?8G" 4Y<FTW]::=-W&SWMA
P$?/X> G'R0# +HW4YR<R67@B"01X:F@IHY*I%;.17\QW'B+-K_-<-S?#Y+!\+)[C
PZ4<$*3H>$RHT<+2;A4.^^=&X\] 68>GN0F'H-^8,1<2^?G"XP<&<A7"VA(BI=66<
P%Z5-V\KIF _H"+8Z(6T$2#NL,5 >YAVMX#I6I'R#?@P)D8+SE;;'=EIO7['PU9(V
P(A1W65A!*1DO!T)LHDO)U]9G5YG7W=FDF?4G+K_K($8#1V52&FPWI/%GX,0D"\NQ
P0_+4HXK_>1[JG(Q%#BO*<'89:L#P@G%MR,1E65^&A92$5[(@WZAS=M8:%6N/7:?R
PP<-VT3>\A%!M^#_>]\Q)<#H95 >7+=(9>%[2@>JK.#[(N&X ;@'0KL7"0?"=I?V6
P/HDU"2&3@/?,3[!S<9M18Q!'6M"!$V+J". _&$6UZ,KQP7A,85?W)O%\GP-GA+-K
PM/0S<+BQ]J5[8T2"L(/; JDL5]*^X:3MA\GZZM7_/NC&%U^ZN4^(R8+6RF>?-3#9
PL]1B.W5TDX)-L"?.^GRG&,-S%L^_S+/4<L;*_>6GYI;01@UJ![WJZ%8  ]=MKMP8
PLI3C^"(.(8Y>!6?^%A6@='NIHNU$%EES3GA"XN>&.2FI!/=6.IH,1C,Q@-D(G:'"
PG.7=(X;%YF.M+F+*;<)/NKM?7IF^23 6%TN>\81\DBQSM^GZC3_6L.\>819 I"[C
P,BFPCM>R&L:=;Y5;8\YS4H'3^D:Q%?Q YLZL-!+@NK<=RE!K5*&U))V)]1IM$+_$
PKOBXF@!N!H(3VCWG=I;U(4V$(]I*RX.:&N<)7]=ASB!MU>D.C-'>\LS?VDH9U$IS
P^US0-4K[VO&$_""X,.R>*9=,2;2!1Z5_%HJP:NYNGQ-4GN)2W*.$UX1+/KF3I<XO
P0(RZLK%>4)O#HX4?>G-+UG$(\WBX(J%W*D03JE?QR;AH?\)/S)^Q<T?!_RFY4XQW
PO)<[*YHE0MA)6>(7C>C7@L%^#3^_KTDIM3*CV \L*#E</X#2?8@"@&6WZJ_HW.:$
PS#>;R6UO>T<82%9 ^PAZI?QX@$+_1>WST#[=H[YD<;D#.T3Q9#;KQ'S,>#N%OFA_
PX482KQY05(\KH5(:4#Y^1?27LKP!"/EJ["M=+#:DZ ;>]F)KZP)*]L 9#%(?D/:!
P_0^B;X4MK>$0&V,OZ^:8[YJ7YR3]R_Q\*"6C&6^GN(Q6CQ7!C8:R4D 6W#;:@7X=
PIM15#5)TX"?BL\D$ME6^<=<7X0>K8]=7P48]OW;OG!]\6N_!CM^W7'QB"!)%1OGH
PUU;,M+#1WDI8Q'6%+H*0%E^WMZ1?F/*L]C^?>S6:1(YF $.^5,+S^=+Z)Q&Q _04
PHJ LWBLJ#9FG,>/^\SGT1L?*%NH;+S>'WV=1HZ(=8FS/)?>GB9>0LFN3\(R-$7ON
P;)!:0+V$3A7E/""=P):D&M;EN_!.QK!M7XP,(NZ:C&./#Z[Z_S^\4,DIVL';2OLU
PJ0GS<&Q=$YS"9E.=MP+A\&>>PFW:2L'1S,Y;%_!=(T+/E\+641TT"9M"IU<R=;ZV
P?<']5[PO<%V?<JB5/NTVY:;N[*%@)M[NL<TW=$8*?XVA_+FEL"( T\L^2OHMH.5^
P</P.2>7=T,Y5(#70(UW>3WGJ]"'/G;>&8A4;5_G:5$VOO=(^$U'>XISA)V-@RJ> 
P02;-XZ/_X=[H[@+_.%8JY: ?/EN8D@6,&0H[(J<FF=<TV'6&@4VK,\DF+BFV(*&L
P=Q)3&0ZX4PG@IG%B&IUK<'&"PQ((JR:M3TKMO?H_NV*B=I.)M^"3BQ(4B-+,#41'
P,*K FKLCRR].:,Q%&8DNW%\LRGU -)@DJHRN>1HA91,^8/IAC?]SA#_\X!X\[T+/
P+%$<USHPGRX1CZ5[Z-I8;8HVUL29*[)L&")I/G<CI#*501# %]RNJ(I'XK$ER:,Z
PV@-Z-KN23EVUM76+YC;=RN3D )MX3-&\]2PTR;<@() K?YS(M!,& ^4N$]FZ#ATN
PM9W0 ZQ&\]948G]VP#%MP92&D+WZH5B?+^>+9;^E#N05SA/IA(X8[U L1;BO7F=9
PF)VM&?7VS:JJ:G?IZ>3.+ST^YA50IH=180IU3=+\CU)K+@Q2O+:"91WN]*0BS]"#
P9K^X_*-N YG>7@]>^&>(/J%2GX4B$;7QC%:H<$: B;?TRS7@+?PXH^*6+&?=UQP,
PDK7?*&.84;$^%"_6L!" EENJHMG+F+V^Z#=F!@W9T9_S'DF[[RLU%7N?U(PG3:C-
P@NQ)$.<HY(7'5I_$RK!:5)XC:B50W)/1E'WV9=7?[P5&0+W 79O5A5W2/ )-K5U+
P+$+^\+:&EV^))9(W)X4X X)I7K9S3SB)Z3#*11B4:_?K!&!K&5>]":J>@\#:VO>L
PVT5?7<(_[?'6O0:S/K$TI8%FJO%GA(%ZC5R*_QYIVTT/%"B)N-V+)-*S-V'KMH,)
PH:.4<)I&X!-^:H3(87E3]>V'$/LF'#[_)KT58Y# KM;(;<TV,]$74$F.4'4Y_7P4
PAQ:=GIXW&\(88_TVN&K]EEZU8$Y%+.NI\.HIJ?B7XS0_)LUC$!).GIV2V8&48U64
P6ZPOVN\OZU2"T!?65BE9,@V*"_J/#U)"C)U(IR%"!P2FU8>WEO;YM;8^".C\75#U
PFQ:HVRN9<%/\ED&;&^T7K-Y_$7CM*]FK0C,^2?R,N2N?%J]2P2!QU@<1,U"M70HG
P6D-$5''<C?\"2C#^"GQO-BDZ2?E7&QKK -QD\IG$"#FXQZ32SKR*A?;OF1_!&TCK
P=&7_"AB.WJ]!1A,,#H>_R^5S%<#6;,095A<L)H)G/AQG3'HE?P48IH;[E^I=(ZD?
P>V0PVZS<LBZO!H:W@-B(T\H7Y:F+Q]QRB0P*BI,UR-.</WIY^"[IGNNGSY]TO0$G
PMB3DOKZH:!NS[K26D_8!X7LV'#[7,N0ZHZ6%?MUHB353"\**FG(-G;F#Y5'0KEE?
PTRK%4DJ/+C%S%-G1&3%U.#YVP#&M%"NHF1P''%)F\*UNIQ&/X)*.YA)P1Y_"'2=%
P$B6K4@!G*]6.TP#<32O8A;NT0N76U=&^%NVH8@@!6TT81R\GMSUYAHB;M(#)!N%L
PB*TE<0$?W2=NX[YK0D#LR,OWEEX2Y\CX?P>5;.]O*,K(RZJ=/+ZA_\W)N?.J*,AS
PB(DVT8!R-@D%O0*#1KHF$G0=7]#U[NW[<(\W0/6B_DZ#Z,/# 3PTW)!#$&G8=M-1
PBBJY.C/'>S5J0.,SMY+PY8T"7>E8PL>W0&\[R A8R.(_%-8S'*%G+8CGD(JDR>9"
P%8L78.BQVG'1E8_LJ=+C RW[-G53R@=N&==28GC-/1XZOT=9?WL\T673$U[>:$!C
P9BMU&!=;C,+-I=C(1<JG_CK)OOM01+1U6<DL!_!M9X@ 2C]KZ_8,SKT5WKW1V?5F
PZT0Z*(2F8!*"&DNHJ%SPF#K&0%>!=I%WR"638:LF]Y\XP*4J%<^JF=:V>#$HLE?A
P52>SNI@DQ9@RVW"[V;M>4*$%N-'-$MA'=J&U;4&_YS#5]+>YRQXWJL2  0?\Q==^
P<4*6FX4&SM\<VK&-#&P3F&%$N1E,*[FS(T)5^G[=7?(#)<2(4/&]?Q3P_\N?G=5V
PET$O$&=,QP!-[#QT,8R<BG-9R+"Q8PL$)T?IVL-K2DWW3'4RBY3UN,Q\P_SECJ!K
P_!ZO.TTDXY)6.5V&!I_?X5>EF3Z66_!..-4S*H-2@$;<"*7OU/P(0V:"+AB^3!EC
P"W8"W80'UL5U=T9T1G0+3B1VY9M.[*'8SSUJ+VR/2GDC['WN@];(II.R%X@2E9([
P_/5/_=0+7V(<(NP%^@/7E<%GW'!.".<5F60]3^8E[8!1</_3JRFDK[ZK>A/93;EZ
P+6NXV)WE/B &?>^.%!!M@H^^0_7.9,8Z1K*  2H_>/NQ)YDI\B[];QVB.SNFTNC3
P!MM1TUA1@]2N+L8E5_K2]@^NV0D]Q^.W0\. GX^E5*@<\D5?S8!20YC]MT^Z]^#&
P^)=SCFTAY12WY\_XHEP_@0*8CC3]*S)27B(FC&8CI*O?$Z-#P#(+:3FV&,/E*1U'
PWDW<ZDGT,4;3YA,[-PQ(OOO*8K:Q0]ZBLR*8&=GK#G95NI#XIX"[2P=->\Q#AW57
PSR$A+:_C"YAMZ)328KC,_<0P&M _I.CG9G)&XVB1T#V*,/#S] W !T))J!+)(MJB
PDB]+ @P)X\E%D!UN@8^,@<SV>SPLA&ECMMR@]1@\MTX?&Z Y":E4'L'<:;JHK)9W
P "![YKSH3]+I^8*=M]S92.M"PYT&?Q>\K392EPDZWWO2%(K_6"R;N4PO&L<[Q_TZ
PZOD-)*BQD*IR&S;UCXE'XRS &1 H!43"T>K'_A 7XJ6J5 6.9/^;"E\IT'AHPA9D
P" /[C:N92FEDDJ ;3XE?=LA4T!-53"=0.! LC+CSXX6:C(3F=E_<W"="9, FNV>\
PK6KXJ&U;RJA^NR=B)]V9O#0!LQ5> H#?>,AL/13]R3:-Y'LM0ILR?\X\#O8&HN&>
P7DH?O.U<#V,-N$?L(]OOU\Y.,%%Y-_WBX4W(4&QZ38D9>CF4 S'=4?8UY6+0>$-V
P>-%8%LVR&E/9FA^MU_<=9 R$$.',11""W(3-J-+3C]7G?O?D0&)V@0UVO1\H!SBI
PJQ!EO:+CP?J.L2\XT6X.ZTXECX^1BIC"26&Z%4CB^GQS*<+-?,)\DB723W[S3*;J
P7_)YDG_2-SBF6K?\J2^LUB9W%<18'8<UT-Y.@UN%99PP@:#P[JD/8V0JKQ B'^=%
P[NX00SD0<QZE<=*U*&9YE]^ _!>N[]>L1)0@%P'+SAB^0W>+),S5!]@"IR)+KN?8
P35Q0#\YE8;$W4_;)&@<J*!?-*[+R!T*' FK'EK)ES?*<CTC(P@KRT!(*%\E!92Q]
P=6G+!Y5XSKJF+A12"D#0M)A[*Y]Y+67+)XTE\5G'Z2<O?)K5L<^Z3UP68RE[-D@*
P*UIE=A;]JU.%^\LHJ3#QB&LHG(2^4!<0HE#^CC\J@ZF5]ACC;9*RX$#QWNAJT0N(
PB 6!TIV/??V4!"1)\\M0^JV.2I#8M063J'XVY48@;^$Q?'".87=TY#!N2X69*Y,L
P'Y&5I1[P-@T2SOOZ>^M.7J-P<C ^"9:33[F.:T4$BC>B1L?)J=*ZFDOF]*E/$8S?
PQW:/+V%Y56).Q6I'GYP![X^0U2EO]R,>:,\^3T9F<M5W+P/W7YH>UH-)&"TI*6D@
PFP.F) #K&$34^ LB_V#=JSLVV\4C^MI.TOQZNP (3K5@D"\DR)@Z$(Y#//XM%T@T
PI8AJ-T8K-=ZKG V@ =MY0= TM,*U4-<$*,SV!]V$:GV+;=9NM&M"XS12P<>(['U?
PT) MTEC!F3"/Y:D=9$T_NQTA]*#:4MVRS^Q_[@KP7:7-F#3CY5*#4$^84&+TRCH,
PKA&5#K43:HID@WNWJ5EI8_TAYO)RQI9)<+%WK+SS$CO3]1;B$4;Z&NI4;CD(MPUE
PT#);XO@@Q3 +N_LFHQL:[0 5-3N*2G)@_V:<IV#5'.LL%O=E\QIB5)GL%92H,-V*
PK=DUYP+W*FT(6:W$VB.&\2P&%!QS?N_9S81\+>\UB\,F/O/A EMN:B3A+.B A,X*
PS\-^I(-[>=@O-W_(,97XO5,8 B:RUL1:V (V?:7T^O=N0 AZX_!"?@1S0>WBUVMZ
P>+VA=/P 2\M+;=69/1?R3'P<IK=6_J*>Y=F!;J2S%?FB_0S:SAOR>ZOVB(N,%:R6
P3+VN[Y92!7$4=JIHE5-7[J6(,E+9)ZHX:^E[ECL0QT\G2G*EI0M7)NY95#R!)X'1
PW-KE!ZQV99I1(9< )^J?DAU+S<N4G1< MM^?ZZ1_1 G$:EX; @J#3WID9B92,E"G
P['0)4;XO@:N;K*=4? 24#^R;H((CV&R8>^3:IGPE 9!TX]YO)UO*<AKJO-26L>^[
P=[ 2&<'B@^+N)5]2Y<7Q&4UJGS7GYH>,7*".,JL0<F HIMJ(%72Z)(A#:A,RE^Z)
PUTJX3+4ZT*;%I1A!0?"UD1KMZJ.R,IAZ_!  H)O_]SV@I[:PH&XB5B&*8G@*%5[B
P'U_:59*V_%<4KXW@&H[>U*T'KI^,78IQ"36\<-\H.0E]=J9X4SG7+J'.*(K&6Y-+
P95/&GQF"%MENU,,$F95V1#PG:J,?S68%R&= %@_Q)@<"&@]W,^:@XQXC1VQ=AKRW
POF>U[,)5K9@;YN.)V0J4L(C2_C5"8I$8$-O:^FTGABI7[%$3N>NB\KK\B/.*C:2B
P^&HV%F1,-%H;'>??V.3CP&?*8>5A(L@[7?GP&E&=N,KBS-H!RX!'KS-1<_&TMOXP
PCE5.8W+,#$+*2&;PDKF._D$T 9M9A:4,9HCG'==>"O:?%+1"9T)L(+6)5@L2?[D,
P(W@MKS:!X9W)'P-N9:$LNG;M*ZU+;F<E*I!CT,)4LN(_9*[&-1M3VT=9(/#RVU;X
P(!:L@WNW9#JX&#H.X]!1/TLWHZ<X,@X?H'SX=1U&.=.+)S9%:^0CS)O/, 0$BP5J
P_T9!QBNCS:'5K^O#"VT\%8,S%T31)C5$R :X>=)=69HV/7#'\]:F[83<R1'J>/GC
PD)#;W504JQU3)!A%%VU"7C[]YX%-6/DW/1W]'_4\3/H']]?2RGO?$]=GR$J^)F72
P2+I$7!AQTP!3B+U(T3P%[!$*][)K8^"4299)*!@P'GHYF>:<EF/> P\LEUH ;W<C
PV">G'SMZ"%W1K65XBX>1F[0J1-#43[A4@=X,K41P2%HWYRWD>9@TPG[C'D.%\)RX
P^O35^W1*T!FN^^M$&#=VI%<,]G3".:4T2$S563<Z'O,L.2HJRDO"XD(ET\T,.0HP
PGR"@@<=H # -\QEAY1JY'8IX3<*+XP:2!\PLTV&1L@=+^P4]!I0R3,<4^J*GL,Y:
PQ7E?L6M"*Q.T+W=(U;()TID+R34JH<T[;/0L9MKUN;R\^Z;N<9H?\<V-:^?#"CNM
P.!];#RR8&\'[I(KN]C^ 7LZ<?<FI&,NQ%6S-$KOND-V3W";@+#!TV$1S&5Y4V8EY
P4R^FSK7I-R4O4>3#PZ&6H*(D@"^ _!^VJ(UV8 YTC?AQ*RTKDYNKV]-9[.AZY!C>
P=13JM,_/)^>$+I.4PND@>.^\S)^QL3.%WG?F-![G=DY'F!K[E4 YRR# T)]"R8A#
P&X^YEWIKO':VT.*?(\H4!'H2*NZ3,R6$L"ZBEMC3E.>;LVHC<GK^%:,<OTTIN6*K
P[J %M\F6\>3HS"7;H4-RQ,0MU%I+:MK-Q?A8_1UM@&^]W<Q:Z?;;NJ;6PA]E,%\D
P\8$4HS&N#:O#   )J\8_[TL)!4'B?H06?8WOQ4XOCQ7YA1!2N;FJJ)'PCO8?[I4/
P>OM*-+"- Y$J]/+:C.!/#T'4)4A[O"\G]C@ O'8B52+!#K!B,7RU4;_:GI^\I]C]
P-D(-P\(TEV%K<O*Q#27K<F\_''_$K5)3566;.M0D[,TE3%^[.$V&CFQZV\ .W7&H
P3LDET0+MBFA!KY3F*6>*[*"PWBRW=@5&Y6G6.7K:RQ!B-#7RW#F&.%;SKSM- -!S
P+O:3IOVGD6H?)_?=I.$@07#V.:W,4R\Y>+[EJ8K$V8L[YL=XTOXK5_AP\BV;M<,H
PLG<TFC+-\8DCD%+&5K%A'MC!Y!MY<I1.@@"JU&08-)X?VA@& ?"9OX]Z/L\7;GW5
P&=1A.V]0&:?N3;DV>0CM4'<AWNP,WB"&5 ZJ>EGBM ::SX-'4J<.&<'?1UFG1-<U
P\%/D[:<-+AID/#;I@(EI8BOYEI<Q);^ G^JR+P/Y=EVHNY$-ZER<?)/[8^HX%>AJ
P[1IQ'&2_"]T]?C7NK;V$S:NO!;=1]>P9@8&H\L$82F4?_$)Q>D$.N7I52FLHMR=M
P"4O__E!&H<6\(9ZM*V*5EV1NAE:!!X(@691=L$)*+!*9Q$*][5_!B5P@Z2\AHTZ<
P6IP3#64<*C$7US0QS]0%D1LB VVJ.Q<)BWUAU_@G7!A6R=ZJ*$>Z4@:J03FMY.HJ
P!&[&XX]F???W$3UO.N3"L;O\&?$*FX/6\4^"/QYV@9PO2!I'L^>SL7EPB1<2=ZZF
PGAMLD-2 +A%O_S?6G\ZS*_>)%$0I*20;)X7AZ:FI[SB;Z1<9"@J^190;%E"IQU.'
P:<S]I6=)[*] L@>PNL?;09(6SX$*6:WG;>@"]7K3:[='9]G<3#X$WBM %M#,*IXL
P_Q/VX3$ZL!+JMV==C;\$':9B.6(8[K4O$X#(3LWO^?WHXOC BE1^1&#9@BZF\U8(
P:=AHV=-K&J#:C^^"K5'Y*2.,I:GVS-/?L\2/5L7-V8)&S9-=D"I$5&K)N4<>*2F-
P-EVDLF:G\!GE-"\+THA8_K)MS-D=PUIB[#H-;G'JH'J]:5UAE&KGQ9N')7S9,<$I
P%WM_]CI0$PTEQSS&]IE]3CE"$0OE[_(['2*HKF=?)8\]96R[.".\]OV?<YOA8S"0
P/V9TB9:B<PD&]"'"2OG+4<MC9 .CD<LE]%K*"!5.SB)EW(^WGSJZH:Y2(!^>YN54
P%$"T/W+'27P/CK-PIVG:HF+?>>NJ4TR2QEW09*Y>)X.,']K$]?J=TN2=WUPO&U?3
P026X:L-U'R)@R00:I75%YQ %A#.7]#:.7;EJ("^;W/V6!F]*\F%)K)>WKZ;P=OD"
PMU7Z"25)U<VVX&0<=#58<5'A4X>'.=J-,"SP/%A%4ZM#X!#7QF>(0NMO^Y@O$6J=
PW_S8*_)R7-+S=\4=(3/R.']$!72BWDJ@@C1;."WTP8;,.EAW@UW=0##W'6^>0D ?
PTWEUGL7#N_E/UG\<PA"B(D0QN;K9YI6ZAM3 B6Y1;!U:E/ 0$NWY@K<B.WA&UCD(
P(H10M: \*5(=5\KONQ/G:[F\9D7G8BD-X,9HS@A_3,',['93*),P 3CRTMFF6;^6
PTGMP?+5((^-B?6)D4L:IS.78V5R#E;'$_MZ%E_&(8K!A"RO.UI?I7U8>8ZH/)U.(
P^;VO2.5XPHACTT-1\#H]$D*E7*))G'F5^'4C@/7K72V7'KMKM]12T=5Q.+'PHLL\
P[:/,R\F?WL&M_7S,F?:_5E1C0'=I%1^G]S"DXK)H'#<BD;\W S"<%8)07^*8?F"(
P:^N.7PF@X%*AJXGC,7:Y7J/&;X#KA)8V%;74_R.3FPU[N<&'Y()/NSLC<1R5H6C&
PKXJZ=/_C2'I8$0NY*#PT1&N<QYMSRC$ZY2'2'*W7-L]C >W;0V61W_=I=PY)KP*M
PV^=?2SE++=?7AZBY4%,YY\!;2R ;W=J:O1>46JW*B&CE6D!V8U4@5X5VEINT6YK-
PM:(7<FQP';YV#[BL2R3>MKYW)'#0Z'FR</UP)ADN,Z,HF9\L^1REAPUCLM6D1Q_=
PU%$5AI<)&/8F6$KK+]^/-F#;.NOKHXO6Y9CW>C$5F K/<GW?D2@(C,D*]1?HJK1Q
PN'M@1C&M]@Y-1I.<94HZWC@B_'?AIR[-2:?K3Q?(;^D8R5589LP[7K/)1(Q?[S3T
P\;'9,=[,+R_#JB-W]*_1I&6<5,N?4&HTCE1<"@'"^.N8 S?14T4TH1J2T+ KR>]\
PTALH'Y2XY;O].J#>=HAH9J%D8>S"C:'$B+2UMVY7\DN;;N2._<?U4M;1)JD#[.G/
P:=WY6]^55I392D3X4BZ'C&7,0G;6I 4B+G:F0'<G=C"Q):E?2Y4KGG&T4"O@&PEB
PN.J:2;D9$I=FTPI; (6\V;#VT[PB6;.SL1^A4\#D@D7VK@'3(%,IA:@GV2@FD1ZN
PN7@3%2]^H]"/>QB<1Y[-0" _!<13LOET3%'R B8!4L!Q<V/D[\^K:VD+B1#=\WY[
PAP]&B>3\9W'B'Y^]GJ"[I*_SMWN0+E2G\JSW5 Z?8:H0SK]&\J?$F'NJ'Y*8F"YC
PL#$[*\B#YA<SY<M/J-@9/KYNF":.@0U;G^!$A?U4XG1.D-0NG=*Q9Q&L\A=OO)&H
P.09[,"X*Q)Y-$^SP/CM)D;@W3'OIP'1RXF67.94" ^<]?S%1:^_$+EB.SU^MS%D#
P[BR2$6IXG D[CHFSRC[ N EHO'4#$D%[A2<JR3E6/J7-7KJF\D@AV1OM?&:'JQ(N
PF^FY>.')1\IAX'#[)*Z&)OY AFUL"N(C>(=&+>E^E^R61BW!1$NQD7H*%L<FU*F<
PZ<:>:9OS*RN8NM*18CYK/.6?*-Q5=/,WC9O=V*$8EP,U8H%-28'>']?=F-78J1N6
PQ3M<0S)G8]QPL* "<$FPP^ R=VR,$V=!MXNEH0'#S29JWWDM/W86N:)D+Z;--<L-
P)EJ0;;W:UH)&9$G"Y24;A8>/0CV"LWN5)$)IS3CZN GAHIP/( :N?_&+\!$C%/<\
PB_^SJ@*L)S8X8P7FK\( T*[S6UEZ&UZ7'79U*N-[](E,\+ACTZ!WFQAPK_?F8'OG
PO01!JKN,(:7A"U.LFT+ *\):K43\(>5IW(QNH1%5_0*L4-'>AHR9%4@,03K2JFF?
P,!WE\BAF++QR1F^$N"0CSUU0*:T=-X4<?WJA(XX1IUZ!=W@8@#'2Q&CFDF;U^.%:
P*O<*R$9?O)HI\'E:Z)&F2;]ER7U"T(A4 =6Y>3<8'J/%KN=V*S^1/0?':2J^.>Y+
P!9Z^L-Z9KB0M6C\5/;XJ2(HX;^SMUPE RT0YSEE^BH#B@ME>VVL)&D0ED+C'7;"=
PT&[ B7JJ0TL0M1-%JR*/H8R7OA\? [6ZDX3"&/Q^FR(R],A4QK/^D?MOW(\]YYF9
PB;8.T-BR@8%=LS%*U.Q[2%EFXD\*T>F0W(8Q-TLU<;:Y*MQT)FOJ S\LJ62=LHVE
P(?QU>,\3R4=ID* 6D YWKUMN^'S'I\*13-HAYOL4,Y>@U\V8<;Y1VXFGNE3W%E_6
P$\9HU4?+/4RK.A!6F 9KTHXF*@G:OJO0FI]4Z9Y!/5N$ ^W?Q6DCH@-4QK=@BB6C
P+!M'>?U(M&R&\1QR#,#+7G'^3RM(#)8#Z7$5P9DYW\*R=(W@U"9&:6>#H)X9SXGX
PZE7S9COX,X($=S07C:8_O@24%RP@,QI.XLTCL[4NV#@"Q*;'1K]I; I@B7JL/4Q&
P>B2)J2U54+X3]BJ%ZX*BNE[//K-*K//%6<REII5*%\AI,Z^L?'%[JL ZOHSM*UHU
P"/Y/;6"JLN@GQ9T:4&2)30W.>O@PL K:)YW\^ ]^S@^WI+.V!0%F,*&IL33;FBPD
PVZ?$0CH&P.9R^M4"]\5@6>26C+^?");QG&VXA3R7QVPYZTR_HAQ'84JNV7:L[V+F
P&YT^!0 $;VB#US&&G1;G2C)V+150F*ZNZ$&?Z:B9M"!PHS*9=#^WTEGT$;#O=XM5
PHQ6_/+^.&A!^AJI=FG [U!E;7YI=W\5HJHZ%-Q]0/$70@=]?+J1-CGW*]_3-#<H]
P%%C[_'=W-:U:3FLL9J'AW$M=\=HE:!IZCX6IVMCO5#E=?L!-1QNOEO<WJX3EKUQA
P?/W/ZO:9W@4H>%S"6LK#QU<<6XYQO+,&:Q6M?6)<1S#2%NIDNW^=:TM"[X4F4?T1
PEA$@YY2-1.TNCN/9]Z :9#N*\.*?A6*Z6ZUX)+!^_>/KGN',)H@S7.#@.$ES95B)
P7@^X@D 67\"H^:+7;E-S&_B<]BT:T62) -0#+(<@&^X%2,^?(1:OY!@V5+B\/1[Q
PU!J0CRDCLA<3;*=2!%[:RN<(=@M&^T[M13$5R3765Y3 'R,;;;Y6-KHPUW,9(!>4
PW/:?&7WP)"?L_QQ=#@NMZ&.4AZB2,WB60^&[I_G>TEVUQ6I6_(HX?-X+L,Y)!,^#
PEY0:<'Q8BY2M"#"DZJH[]^YV(:KM,E "QFL3QOM)U8?V,03T,9LPM1>=(X$)D@'L
P&(;R-%T0!HXIGK !MLMVRT1R:G,AM^C4U7;20W >6."BFO2R9@C11TIR\' CR99S
PQ\AHOLETE0AK%?=U53DT+&3E@)R175C88.<.CIY>Y$^\VDO<:D4MIK)"O&=;"IZ1
P5%7A_S _)SGU8F__91"8(G.T;9!(1.F?3_ L.V'@/;EZ6#:H"US[H&/ID[+L=OU6
PODE7)XUW@-FBRXG5N:P>GST*M22^+K'Q#([A:6([6TYN[Y_:G(LYUFG-HYL+D!Z1
P_G*G%R"(RB R+V@SU=^< MDU",4"OONWRI?,ZK#F]P%J1*B&5 H1"^DEAOBHI(GX
POB,8F,WMVR)D#N&K=1%XF6;E<>7F._;<W<0VO!GIV13"RF[R ;#-SB3"NQV3]<H-
PF\L4' AMO5A%F#8.V=(467*H>Y;[D5758=Y A@")5FD \:/46CIMH2ION-'3.P^^
P(!NR?<T%&;)$S]=W>\(?T!'MTT.)0&*<$RO+*Y)^5UF)!2M>H.=?;TP ?GV6PD/7
P9ZZ8AE;>A_Q1I0*A=Y,D8".?Y$@[3D1I2J"JO:_#=&BXBCQZTU_^I#G_=CR!$L_U
PD*9>(SPY[@#Z1KT7@-$7 Z'-8('E^09E+#C8VJB;N^Q3=5"B\Q'AXR4L0'P[>VH1
P'0_QB%SX)U3? 53$_5JUO./VV8XRX>T/K,Z OM2[V9\ZU@!U03?GF)C,VL^F22[#
P:V2TF<#(H.T"@PUXJ>SEP@7<-H4RE/')#M47T<@!; W0K<94O8^,2>F-+X@L&!CZ
PDQ IZ^ST09?')XMXO1/'<ZS)^^%48HZ:AM*4N9O$\9+LBJ'5J@\3_F*VMW0@_X%A
P2%28\M;70+W)6>$7V]5ESKCZ^RXFKU]4^/C8@'/_6VU29$;QI\@NK 1W#>$"KIZ:
P:)#HK?/S/EE.SNR%^;;]A]5L,Y_6%UG'J@)U5^6R8;>,?,#7&B5-V+YIR!9I\$[8
P>!O9P9CMG^:6"A:X$AOCP+4BY2"MB4S4S2$F&1&V+DZF)UMPD6WV,L(P90$.XS0_
P_.MPTM+/E@ (/'1<\_J);EETHF]S65^HW_KJO<5!M8Q#K%#ZN/; "1%.?P='CHLA
P7PO"W!?^J_""%Z[/]PV;1PIRAT\[[JZ<O2.4,I2C9<M[J6B:V]'RI,E0.SD+-RK<
PF7Y'X@46=J&("/<*,SHZ>*)GS$N+CKU_XBM*:365F?^%P#X!Q\E!PBN<$;WRM%@\
P(F#PZ]_7COXI"?(SS;RZ5-,!M_V&MHJ@C9B^@3L_#$[(%1B?=2YE5<7.##37H78\
P%BA@I?>I-4".+[23R^\@-<N[Y&:<KC[$'7[92Y2B(W.HZ*XK4-+^/..8X3ESA9J"
P*@U>%W?U7%JOH[=IS)>[VH<GDBD;#ME#U,MC)Q3[=00A+2**3/+;( [-C9ZF .W4
PP_%$P=6__*SYEFYFI>@@1U%U;7_O$2L/YB2O58[]W0I#>X[U;)#TD#-^1/W_@)FR
PL_&DCLU!^EMAR*V8 07$QOSO>5MW-E7S )BA$L0=ZRX8AB.4H+K:'KTL^7ATEC[4
PU?1<S9!^:OQ*QQX-[<\/X('NX"0V\YQ<TN6T8NASTXM3T\.JK/:!Q_,FYH-7O0E:
P^%$23#<W>.K-,*F_U-[-;(;I=.0%PY71W'J*][F#I@4M19 ?'T(D$=)'C<]=DV/(
P>VV^=$I4+<M-AGARP(\(J'+"BU*W 6K"*[O*"SNI"8E84SG]KO1=F";]PTOR9V40
P\\##@/F[*O$=8B]G/OE[1I"838>(05S."\2!LW[7&Q_2<64#S9;W,/HG@>H[:K,$
P]2W>?W,[X+OV,AMB=CO@]\0;7$IHA/-2^6+:8A-(4*=5]?K8>F1 2FXTOR1?M%$&
PG61\).AG<@G%E((^((D?1$6C!(DD&P1#T),":DZS^;!<+LQI!0U@ M#2V4&'P+M*
PX)M'9=I>L-PKEW=\M_I XN?3CJY'("<W]H3]N^%E'55":R!U6P*G92FR=\N0LYZ9
P0PVE*^YIY29XH( )5S^]"EVWQ^2M_!+Z\I&; )[?<0V>X([X_EUQS_/4;SQ4^K?A
PGQJP TFEQ7.+$E6H$1AKRA B*7<@:DX7)('_Z-W@@ J&_=*J-;D]"B!91:[XH-X2
PN5_.%"/.OS9XZP*G,'!]!G'/NO+I.7T >0IU?Z8+ONYZAGLA).P0K9,.T2E^O78&
P_R="Q1A(]2@BL,\^L!8\>OQ:(@;'UN^PKYG]5HU**=\SJ!DAIM8MS 53YP0-R3JG
PKN EUZS]M4MT@/E.AOO.$T"G,I$N %'2T2M4JO=Y0OO7"7 :K;BRDD.X%>3+@;W$
PRF"X^;^3-'\%IX[_]LLE94 UH!92!I(2*)'<A;:ZZ&+(Y&Y"V9IB9:8\!^<6  W*
P(<81W%5N9QRW5[GWV$I&XG2C5MY@]^Z)?)T]GZ-[C55TMM#'I!=T->0MC)?!S0 ^
PL<LVF1FT\1TR]RH!=4K#C<K?X\@?1L&<(PW_@US"B^3[ML)&NS3%O+?UTWS22/\Z
PTER\,=&V;B;14Q/BGH$*5+"CO$N;>U\MNCV45 1TAT6[*-*%&8Q&'\K%&!9I&G>?
P#GP9E70'Z;*JTC)Z ,-!-Y[Z$>.+:N^HEL,WB7-GZ5*/#.H#7N_O3"M36J#75[5H
PC4%+4#A3S5,ONJY0*+SRFJ,FPWLZS"+2@F:3L6*9! Q_J$K+9KT&XW32!/*H,RIK
PIC"1F K(':!6L(<Z6^ J*:&L.-2(5/*K%VVLLG@5 '/:3^/D*4$LMKF?=%\&ZP_"
PHMRC4&GK-)D(GTZ#?_OI?Q37+$WS[9#_/J2&%3UF%[M8_@\?! \1'%FM_-L:'%OZ
PCYU29[@(?F;G>QYBWE3_5.?*VAVM"'#+.3A.O-@H_2>E-*OKZW\Y ^EJ\YIH:,.!
P@"P<P>=$K>\^^(*#'9YB*C[C($YVR3YD'<'I/4P>9Y8;78+_/0GVJ ]8B.'E IPD
PIP:TKB L ;1[.3L5LRN)V/+<S2MGBJ6:>;&/F+?6\BJ(85Q5FGP>O_&H(,#=WH*9
P;8+?WO30SF8N=[$#<Q^ZBY.+U$$9N4(M?U\F\!=,/2=X43D($$3,#%6W29T^3X@)
PQDR]\]8%R, .I<_:)U\Z;13PY:NGA'Z7RE54T9/S<#$Y>IILS>VQ I7/FKYP32S=
P&];X=69W(9.2?N!.J%$X357_;\/B\>&GT(BU&0>+("ZAQ/-X..X/<\9G__ P<"^/
P<.PVWP"^=D9XFB9LW(VQC9W,H*EMM5 .1!"0JW6F>7F)9$4K(CTG@'(AANJR-*[(
PX$6#MVO-T:, ^"X#(WU&<J1"G:%"N++8P8POXUSAR??:SI"5$@*;896G-#-2'0K*
P2[%>9=T$Z=.E+; 5.<I"(&52*^4R1U0;$!2'NR1\-[+9YN.?;<!";6B"',:I+\K[
P/S=\M>ML7(SL9QR4RG*P(:S85Y>@5=6FB.64N2HI0'B;&)7<376.'BUZ=<Q,X[72
PY;"(CL3RJ252?[=<2W=TT=UI$_EAXT^Y)1-:QGV'VLC73<!BSMNAU%$,_"Q,R*'Y
P2GV5_^7N^6N5EZ-9SX'//?]>U>1C[5/:UC/?EL==L)%(Q9!.&^G3.NM/6OUV ?3$
P8!NZ#V1\I@D<K8@*I=; UC9:CKW74TN1>DGDM6V.[6DWR#5QRF[()BR9$3<2\7PD
PVP:0\<GK]3D=RBBB^HM&8%K*:;Y0[>*42CMHSH"4;*J=S.,PU,$^[=M!"_(^7660
P*^U9/_H<T(=%RG'UR4*0XVG4/*^:[,\!2&)\F %%%('^8B'#Z J5,O86Z <ES[Q0
POPS&D%,.%QK1X$3CY0J9XQBR5LK,(?)0B7#%QVX'8EFUK'61?547<>>5/[,\@6*+
PAN&$=(34G4FKX:&B)DT1Q>1J]J;+74^Y7V7@'.REJQ+;<9OH<657'AI'B[MI7]6&
P\*KIB$K_2?#>4VO$B<F%M3V$I7O;%)S$]XBR"C9+>7^'+YC2*H'CV=/7,APX?W+@
PN$EZ"I-LNF'YL4^MTC1%<5P' _?5)/5W";42:J=W <!L80UAYFZT;W1YC1E6;?*=
P5@;NX%J6W)T'!8$7+L+G%\ &DKYYH%-R  PO_I_]P'9-7T+1<.&']J@#M6T_J!1,
PE.X)4X XBB%[WZ^-"R&HA:D:?6 $JH1KYZ,("E1:+4#M-G V0<.2CY;/V#7]$.H,
P@+#.* 67X$=9 'ISD!&Y,S$8P_K\DOL+Q24B.XC=*WK\(Y0;1BS"0D)^L\A<64N(
P#^,97EE7W?4."V_+(]P9R]=F7PY! F+!XI=OLG#/*J("KD.?W[IO%"F^-X"I0T+<
PH3,R[LEG96^1*[(& (=L8BSF2)W@M*(D-5S;H;Y'?4R ,+7NMX_Z9Z8K&<6!VK:3
P&6309NZ]EDLTVU]/19%B1"^QUI&MYFX-(9E)SNU&Q,29:*0)W8&@.A*A# 4+ZO_&
P7ITJ7-6TK7[TN&&6@%QGJ;!_^>)!PO(7=ROPG&@D2TQ V%HQPMK*YWCTX>F4M\4;
POJ4?U#V+9S#X'Z^7/JF1&C Y.R[BL4$E#V&H.HW"N(.5:>W+.F8MJ,-HHVVLG;19
P5W$RD44-U0%A@<I?K71]JJ38$D5I A]P6DE_UH*/P4B0%[#_Q3JX%C<5LM0!(C4P
P%ZZ%WG[R/*#Y!/GH';P2XIE&M:D2F HA!>)H5*ZC,()\5-&2Z=I6$WP[VJ@_5'RL
PMM/LWH@S,KO>[*  *(0_3$QN2 L.4Z8HB'C"D97&B3WUAY*[P"+Z*,I9#$=K2*E-
PJ3#Z8MK3Y9=XEFK;N5(VCW_P^%;G.SX)"]6^C+7$P@5RA@217LF5*@\<I"H)53V(
P.%>T3D3\.Y$UD< R8%C]_K8#LFZ!7>FY\Y=@2>'I6KP+KA2R@FLXC74$WWEL_WWV
PL$9)QW'MB+-40?7\)E?PC&AZGME/("Z9^N*\"P(;,C:QZ<Z\Y7&0B;O5MY3" P[7
P01Y'O6H =F/);IM:AC7[P:@WY-3 #'#LR1 W^+OQI-PA*X#R:Y(CIJ&CD1M+VE;\
P>8^_XT#2M[9".LO,5=ZP,J$?=>YU#A/M+,1H>"K->8[2#FWU4^%O"=CD#'U F[VV
PLW+-83#)<U>;OOM[.R)"TGXZQ7J4&+RSUKQ-IE3H-0KVRV3B2+_'* CHKXLTUU7P
PG!#Y/\&)D_(RUU;S3BN]FY"2EI$BO_9$,)%'L(4_]R"2Q$JQ96;:LI6V1B6AN+$B
P#TR$)\E$E[2(P_R"#O,I)2F<^NW;YSO"&7<%-3PD5?&O+:%W%ZMM<OTN8S$YA0P3
PT(HS:-K D*UU6)W7]Y.202,?^.Y5X7U'9M);]-QLPSGM5^6#B(_.=D'F1CG686VI
P5SI6+3_*JT2,?@3AFU0MQI.XUK2D%,[ECS #&(<U;7J#!S\[ST>[W<T^S"L8JBO 
P&>?4(9!$5#F%UY>6/ M9PP4N-9[+P.ZHP3&FV_1?L+3T?(!&@_I9U^:&(EU<[:>U
P8QJH#G(R0542BM!M=\#G\KBGP@YNL-VFG+3\##V;74@8P:'&OM!5LNO>S+@IOZX@
P0+-\_>-O)ZO]6=HT"(WGIMI,Y2+J[]'*NQ^U%'E%K,#C=Z%JC/4B\[(2G*_W1=B(
P[-J8LY,DHVY)A4';8F*BB<U:N$&*<VQV.^)7@"+-SH,BH4<_*05G9U 98>C\RY:(
PBJK:*;12"QAR,A.0O^;@])%L+-_C*P-2N\V65X6ZR;I!9\_<O@"H5@R<;8G:S\X 
PAX00[*R.NZ"I:JCI#F_NR]H;/P-RBYF#1*IB@J8W(A.IF$BH9NN)1G1!M#A#W\4P
P_P_+=B(OP6UOH==^:I/-"Z'6"DS)$^M8;EY<X=KU1M*!S9JK)," (W$DWZMH(CY?
PCL_.5HM@>!$Z_/.8VG;78P0I;!Q"9\V[5%S,-W29H^&M.=U86OB&/TPM&CX?2WV'
PPK5#()31GR$'/VT_$5,Z7>H>EB C.D#H_TP6H@">&! !G1@MO,@LQSU*AZ4C-<<'
P03#.J&$&!C-="*D"_82C;]-&+)B2."UW#PMR!9L3%4B*4U*,]:ZG^Y6.*;NE/EM'
P*..V;B%@-LL#;4^*FT#$4]W05L$0'7S'PM+.7W6C8.-1]#*YS83>U0CAS^N$KP7M
PWVA=&T1WQ""D"\/;@=M<DJ6AVZMZ46]0Z]%T- H<D&S_/IS\7-C;*Z !4W7O7ZS*
P\U$-KUR3K8_8MV5]0YW??N[;Z.;7D+E6L8LK4R^4BYO47S:8W).^HJSEQG55&D9<
P<)+0A<04+-Q:F:.010EC<#5ACZT=[7.I*F[2"A!J3V>YO<AED9!&UV9WN8&',I5<
P=7F/H-.WH@E7-]TZH-992B<:F@4*P;/=VE\HCI&RP4 [[CC^R55G=4-4Y>]134<$
PE&NL1Q427/89C^*FTZS#*Q&^[.^:DBZ39\2L.NO1V<C@\%OTZH$:!ZTWY-_<SMUN
PW_7OM3MQH&E4S7%0 1$%.6;&3AN^*Q_!LGS^PG&)IU%Y[&)K[#JJ=YM.XQHYF19X
PA]!>Q3$GE^L>4J\.!N0X?';58T97:#;F)1[S.&*KYFZZ?:MKK>U;Q'6VG.HGMUF-
PCBLIA.UDJ2B)ON1KY_Z\ ?+8Z: ?,C\Q\D29M\=SC,C5[(+7C=^JGR1>(RBTG@:D
P>JH7]6-*G<PY2*8P ]?P/A% '9@%PJI&53@T?64QQ?H;:C]8;WO6)$;V>H'!EV*M
PSD932F()A<FS3K>KM3),B*DT3%2?(%-@$_J%3\LAYEV]&6M0V\3Q8XS\(^>,DRQ)
PG:M7+31O6'MK@S,]O[$A3D<\AS6*YT%?M#B^4_YA/@&6I>/O[AC/-*H>:J7%@\$\
PK['[>MI8OZ^&]5U.4.8['W7D-G_+R&QPJ>P>S)%"3EL*JZ%JE\HU&/6ED?(''61^
P-, !,I>0;"^77_44%@THOPT7?Q3"1-&JF9G9?D0.H:*>)NLP.BV.0;Y(&=ZC.Q,$
PE=8X5<3!2M?-2>H64-_U8-#X0#U)=R.Z&)AM!'&L[/O\O#X;:#?6/D*1/(QZY\F<
PZB?W2D<*RBJDE=W17!G!+/)5WW*P'IK\4CV8RXN@GR2'*EU)9./=*=EB2K@%,:NQ
P;A3EQY9 :/F$=I22=G\IJ-&\+EM@;/;+&>\-K8)IF+JHW'5@%A'KV6&\83%;\MF4
PS/ZM0P3EEK0'P(F2E0CZOZ!?,S07K]EB7@K<W,=/#H%3J!^/G^4U;K5116#M.,D!
P#?>FY^47:Z%=AY+AS\:^"OMQ(J.+\V2]GT,]5.J OY>GQ<G#H0RT:+_C+)73"=-%
PD;^P.9;]?32:]/V&76I$II@(YFK]>,W"C#G3@:>FZ27-!3#C$.:;*I9'37/ RRNP
P<T%4,6=K-0+;K+I63& W&:_OI),9_3ZG0_)8D90+$V6 GMX"%[C.B[\KP\M9[@!*
P0Y&R_TV5>B;7*>4954Q9[6\P" C(;<G\H%OR_E!PP]N&RON"R[N/ /Q&8@$[MXCU
P8T?R2E[#!&I0S%^9\IUTLT%7;QM66DX,N.!\<%D,&.3#'3V'*0!4*TC(0TB47SAF
P802@!?V=WFR78V!S>.S!ET1([)B(IY_<GVT-F#8,<?*\BJDN764"EI]S^=*_!?'&
PXR?A+NBL@*[=+VZ0S\WZS-3?@!P#(0V?G/J1,4H"U9OV;=?'=^BY?X\V!XS> J9I
POH^CBL8?^*+_!4EYG(R .#]_SG#XT,OP$$R'^(D3)+=)E>DFM]'P*@$[4P&,ZSG]
P'G&<#QB\CG=J,I7>%J(]-+S+:\,G^D3<[6HEY=/E=&K0$*DU@'\&@NI^<X7V5FOK
PM58J@&R$D(>%/>PB.FX0K'R5/RN^HWB=EZ:$,3I3B0X5)=#[7PB\M_$?>XFC881<
P_:O3[HR=N/TET'&#&DV, K(5D;JA$^"C=U-%,V1L+G5SVTG9%#HO:<T/P\KDZG*;
P?XA%S3BO:>.$(041.NSRT.XX]N@T,RF*>)C'4 FE\ )"G@RZ1IL(,.7?GB<>!AJ%
P?P6L1N3_OCI7#1ZCNF[E=&*M'&+E0I2!=.Y7FT=DNC#3'4%\7,0>"8/!6[D$2'0W
P]IQ^Y534W6K#_.;@72Z-6?W<-JA=(< Q<=!0'=OMV7 '\Q[C77)=&3"[S^::/6"7
P]NEM)Y:/?(0H)IR.@*$,8?E\R(ANY#]^HZ[8:OX7?M]\KC]5K,G85+&2J1Y@R0K8
P#Z>0K+,D08RWS%[?I- G>'CO%J_B_MFG5$]MDL#N?%I.-WE$#/ #CM-6#!C+$V*=
PJDF[XQLBI**@!;1H[._-"L^BG ;WH<#%]5)\ 0HF*Z_QQYIS\ BO82^Q)AU]\LLM
P_\>_0_*=0<&C'WQZTG<1<2^)M[U0^=UX_8&J"WRR(.BSART&^<+.<M1..W]G-&K_
P&=&O?YD? ?$6QOT@T92G?=OAB+S\H,/%KJJRSVEL@2Y4SH=MJ:OQ[_:MUH+%\9I.
PE)G%KYX@6LE:%PEPV*S9J;\#OBV5O5XT@3-)F#2<4W<2EI"5'5C]%,S;OQG<,-DL
PJ> P6TT-N](=FH[YFSYD1QSL^"PN!3&^HEO-)X_X'HQM]E>]_<DM<)!1VM10\[T;
PDIK>O2%H/SAY@%<-7A(A'06!@8U^;K=&2:W6H<OVHF XT.Q"!8C(8D>[>S5]=$"'
P*?Q(L&90JL<*3D["&[9A>:>,932[=E$NTRB$_K9<\EZW['R+\V=&!+>=9#DAPDY%
P.:DT$L$_OQ RDX][?G'%N9K[EWO41K>TOF( 63S#\*M-&>R<T'-]&T[S%77&ID'&
P(/T\88Z#^R-I<^\QM*-VPO*[5ZR)G?VSO/D$-'YZ9SY>Q5\SE4P+9PEI'/(^GYQW
P%?;%4MT*B[B%1S6S.8%T-HH!@!X6%^2;RA*J#*^V$WN@4#0G%2IZ? X*^?KGX/JS
P1K_P1U/SR@)I(JX&9!%8$OU.7V V,.7A+Y<4@+6M&#*_"+F($7A'L!@"QWR]="2O
PL[W.XLQ/5N%N&-^$[6VP4]6'QG[\().W&C?W'(^TGHW(H&LXG/[KQ5R]F/W\OR.:
P\PO?FV>5SAS.J1/\VDYM7L@)='X8@XR+A4GU]*2>!,&P0MU"R&:96&B"J/03R0W<
P"!OH0[HEX>K1K(@B).LNUL3 U=T:I3#BFW\3!-PHJF!;LAM;%K0]L @^>N\WHI0-
PR]-PP^$S^.>:T>O7P PYYM]D'ZS" 1D!L,"^\J9D@#1><2(D!;?6WN:9[-1]#[Y"
PK9TPH[I^+#YVC$?K27;!%S&Z\VM::<NS685=F,<S?G8C\URX,!S$(T%K3#-,7\ *
P^E[\1]0:!A'>J":BKA.+?5E0]IS-=(WIR+-/B%KY.N_!3D%GN:TD*A1FM$MQ,(G,
PHV3P$^HN?OU"0.5PZ\1;B.FH=B==ST!D$#(]IT$[6P%3#I-H_CM.=,3@Q[$WEJQ3
P=KJ2[&RG]-6WGZ!]VJ:@Z?!K<* + VZDNACU +OQ'H$0&E)#?.Y%"M2D U'\V !R
P+ZDTRG:S%9<TZH]\L,SVT"1B\]M%=7QQ4YA+$Q"1**()B265MN<X45?EFEE6HQ"^
P=VL)]W!,RJ)F6$TIQN5Y"+8N+U%^7NL&!.M0I /!BH FCC0?V#W,@W-?AKIMX,X^
PE2\[\IB:"5ZN:_3P*03#;?A<^LH?Q&N3JF&D6,^Q'N'?A$2O9QB-V>%TQ(<8<&P'
P4-N^#?YQPH:K=9=V6:H&,TX5WR[EI;G-.[\L9:7IRQL]!!UH[%(M7DN%3[:$U@. 
PB! T/T47&SRRDGY O_HPFQEL6TN\>AO@^I6M?I-BH4T?)N^?I%R?%MP@Z7"H>*\N
PW20\L))6W3>_7P]$AW4*4+$\I BC$]TDBH,QB(3>#V1?OAS<(J<L^1XQXK%<+Z:M
P\2K&AGQ?[$90:)BD5K-A7WX_29&OX_*^\&.6WTY 3?:N1I>">CR:*%#Q?B5#T@(D
P<M,)EL,I(J)<FVJ]A!8\!HTM^4\F[;GL9F7(P^5H!LRG5YI [&& 'ZL0N J%5D-(
PN <+9 N(FWS6@5\PD?Y!_H\=C>:$99"]P9Y,/J;:V2W^_@NZ[/Y82(0NL($>F,V/
P/*R?H?1=LK[0D%];#>\D-PV%!OV!=?M[C,RX7>[L8:(5UXC LRVQRD/JU%U\J8MJ
P&*)A-_3^ U,#85:PM@M7CD+0MEC+B4IN4:MU09<%B&',)QCHSOB@T,#0!:,Z]]<#
P! EIPSB_<D ]P^YY3U=1?'KA/7+*Y_SI^!KB5MTXLH3%INYR5G&2Z9R Z9M-> +Z
P@8K;>7 2F$9H3P+/WP)DBN6IEC.WUNO,E[/<#U/ _C1TDF7 %"$D@%-HN1N%'55W
P"69-$Y@8="NWCZ1%R25*F*ZG=Q:&[2Y;"=Q@S%MLG8U#D"L>\$-VAVQ1X@WA155Z
PWQ]HX+'#W7(:,0Q80*6S I3SV$WQ:TW61&'X.019Y7JHUE' 2OFXRK(),TU/6GIL
PE I'-3ZR*,X/)%XM$ VU0N<\4XY5F;LB19:\")_]D%*C1=JOF"9TKIL!81\].R#<
P(B#@218K^*:0!SQY.> %H$4%H9*7G<D\H61_3!LU?(:6LG00BDP4M5I^R5_%GGV<
PN_=O"QP%A.F[%P*F]^3BHBT6A<IAF$5@/?/@6?J!"\LAK;P$43VXC0S?A:]IR:=O
P<[U(E[R/0%Z_KT0KB#737_LEES*.//-YV;IB.3TJ61]. 1!?J=AEK-CK_@[.S0@6
P)-_@"8G <N+\T2<[%,\I:TQ:U5B&BB\5"%:9C=-GH#!!B2Z7JN=YJ0.RW'"MP^ !
PG30M4+F^%C &GS9O^RVW]%?#QF9RYW9[H'9Q"E+TRN&4&0ED#1QO_L#K25:1LCJ0
PX-QC;*?<"#WJ J2(LN<P3F/)I[C)4A1T5FZ7;ZL.684.3.^A0V]>,8 *:]@,YBIN
P4[;A)WNLV^=N[DLYXAUZ$H<;ZCA68D#/J:.LQUICCH0$/(;+GC[ZV]>*0ANYLI1C
P3@P;F'V+"'GJ$[+J(NDGDM'X)4"PFOZ9=5-Y0LP%)6&K>7&>;C44U%WS1\EDX$MQ
PD",I 6\N1< IGS/%@%R?FC@TD%:[J57JO 2\8TH8.-CG:I\0^5HPSW?5!'-= O4[
PG.H:=$ 'HO*84I81+,^^][6N#NJ!VLMM#U'FA.5(6VJDB6$H,V=?D2MGVWP[$OA;
PIV5NB;W-FV[-B6'HUD\YD3_61&\&@&]4N>.+KC_70C(9I[+R"T@':4ML#(+=3'IC
PP%LN&$-=H,@0J1%U@>6[S1_<;3MD*J_Z@_GA[I'VI(%FC6@V![^5!GG,7&W/SO%=
P_)V.7-QT@NR#4%9(\3=+ I[T1*J3PWEVCO:Z&O;63--0J#[JW/!LAZ/FIVH,3*XY
P7TE9%V>"38]6^V1J>4R98HC$L\>.(3?2:@EGG8BEN!XK3,)V*/JBU" EY$YZ&9-)
P99.GQ&WVOTZD;1D! F):FW'DX^,,(5<5V>C4OGZ,\R!VY^600K\V8]U29MH-P?<V
PLYB&%CIEN_(Y@W"(<: 6.^^_/!KO"TYN6+4X,_TKV$!Q,\TAICV6<[,]T%6_V!FK
P2CKN;N@1 >9G#RYXM(6CRPF FMT@XQXM0^A$XM4F#Q\>3/ 0FD&3KDZL3"&",U4]
PK9B;,>2M5'(M;0#WSS]"9"R]?]@GHC/]M$P!=3^C+Q";R GPPWF\:J%;?R\FP[J<
PE.$-LOMV  P/9630V-!1)E"^-_/MX7KCQ\OO (HWYFS1L!)=(:+[^]$9;&NN-*Q 
P7NH2,U! !9KH0*US"#<BE-2(9Q4:5=ACN?856&8S4^X2<+GUP\3A^-+T1B0>VCKF
P8BB+4,/&&NK<IO3XK1H\YD.0P>S.5F,F^3N&2P7D!]#@:A>3@I\%$]UEJ>J - "3
PY=^#03N$ I57:9*1CJ*LYT#J;T+8*@</6"  .Q56QCF$9D+6FSIK: 'K$2(ZOBWD
PC%/WDT;7+L8-3G^J 2)Q^4:93ZN=: QKQ"WA_Q]A9^A(5945_4OO*=IU+S:?@&U[
PU6R%TSQJVW]V-N=!W\R*"L?],T!IXP=;N:A:&LH(L F%+<-1<='*5G"V4%<N)L0N
PIC ,1'(@F4E4>>6$]ZGZ.J%=15WH=Y$Z[R- . QFL=GH5:IHKV\5&PSFA)U<.\O'
POGA[J !]O([=4P <J!B?3P &!SBFS!GQ]U?,;2=+RY!2>FZ4U(\+?6=X7$B^$:Z%
PNT6,#-2+WG6@TU'1F+59V^F%:V9=X0V)J!!5X6B3^)QX%E/AX.SI^/?/^$TGT.5A
P=Y6/TWA0:/A>__?U'S<)^BV*#3.*;ZI:SQ>3J=*G]']&1IP1QHOJ9M0P2RMX#]&G
P]8\:"?;AB6[K+N*"HAH-^B+M&],%2K%8L_/.%:=O_?AWA6CA_S.8 5%I\2+<YUX$
PO7,E88>Z5,\HRFU<A*&M-<WNULH.QX:>/Z9\:'+R)13I06[7\;9:;)K(YI@\<GD+
P;!5SOP; 41 :;=NQ/LWW+W@D0EEBYM APR$UJV/NH(2[=L!W:UV>I$@BOZ:$([U_
P3H?Z5DF]*;GT-CD"1QG5:CI+D"R<,6&H^;2O9B\<;/M6X+%GG(!$1ICL \D/$'<G
P:5*0!]J]7E>A(4$(=!GN@L$1#O=-EV/3.ROV\C[O@C;EM]!:'P<<+$Z)9<DM\FQZ
P-KJ/V![+&B2J.\B,HE*%M=#?1$J/-&[<+#R1_-#JH<#%=U+/Q 26C\1=ATJSPV64
PBR.JS6P>1#2* U\*@Y;+=V"6XLEU/N.(Q<1&@'+A7GQCZ,1"'/A (<>Q*LP&'9(;
PJI&,T/NN A44+6_&DK7O\,M2'V%!;Y/W\]Q25 +N1:&T%IYRMY-UF5-]Z]<VYB_A
P%5!#BT(GYQ-[9:6&KV"6TQ\7JQ/(B(A)"W:\[]6O3CY#]0H VTOT5FXA6'[ZN!J%
P\JYO-7R)3^/<0BN%1(1LXS#;?EH!6Z;R51#0^-G>O$9W$X,;N?^$10PJK+UPR>KF
PRFYTABP!-JT[&<V(;?T\]N>JHSOS:S?"L['[L@2J(YHSH=*5AJ'@M_0X@!&_XY@"
P[YI/SAXC+C!%;VG8_7V]Z([67"N6-.)QOPP/>@.P7QZ_-(72X8P[?0[=V"@T3*1%
PLX\K58A'Z<F:":,\RU;ML 8^5J9WR+GGMRZS;[V<E3@&MYZ,1Y@K/&)TXQS8+A69
P+YQP^"E%=[!87"7J),US=3.VPRU),>MEX81YU4FI_3T;;P/C79N']DC/YY#A5)')
PCBXU0WHA.E7L#)UZ_R@VF<C:@+JDV8X9-)$A<.4HUN77HD;6>LI(/JD[T$"NDP?N
P]J6D9Q=<%62PY8&DA>[YD4R&W-2G9<+ 6R*ZH[-(-L6$"KLF]?S_M,.@9+-O1!23
P=A+<%2,@,)Q IN/MFR_7BAF;,U3:NIB>G4A95('$A/]-,7 [\N-0:/*M->P\#C7S
P'#<OZG#V-@+5[=P/+K5TBW8BA2@#"^J'C4*92.(]N\*0.AHM 9K+/IYVBQ$>?#B6
PM9^98+#P1%XJL]F>837BX<N4L&TUA2]:\8OTN#>]IMY:VHD^)J&=5A915E.J05D$
PY1M" -ZH?.,0Y-SNF+BA?%/>=]X00RGE)?W)$CT*XOV<ZG(<F1*6(WEZ0E-?8_>"
PFF\C\/V'\8'7#,HI++<6\JX7]5I3FH%EMXB0= J[>T9VI0L'NA="*E6J'V-(T.Z7
P_+DPRP$R2)BTW]Q:"B'</>I\%'I%FF2-WP($(BS%#Q]YW@:-A"#]>N8DY90KOG*Q
P^K.PQ,^NP8O[.&X($B*?&^R9+Y)P:A\EDCXQ;[LD;/2^9&\,QZ_UO=IKG5)"H6]:
P?$53]$7ZF1TYV0G^U@.NVRL+)/Z9XGU@/G%LNI"1B1@XU5B[-T3_CUBW;.FBC+M!
P&"XV3)WHB9)-\X''G=0/*4(R-&;:>]1 (<4OE&69Z0-?I&I-?5N]L'&RYYWM(S(1
PF5D_O^UH2Y>>2-8@ V&*DXV ZB?L\?E,\V+5$MZ-<'8TYNZ2^(]T\-> :"'=D(HZ
P96J@<D7Y/?P[ZQE->\+\\A7;\!PM'@@RMTS^-#-8QP2,3(#^C39\N8XPHPTXGP:6
P!(=Q",6HL7O*JI2_W:0R^.\R[\Y6L>&L ;!;_JODVVH"Q[W@81F/95(H%Q^+5^_Q
PNF*D(M_ZY48/-XTKF2P2%RC2U*/G;MR8!>6#4 ^"YUMZ"I'HQZPP$W"S6ZP1I0QK
P] "G3P?^W!6-J7KO3WH#=(=_/"5^S#)G!.&=-OG-K-\BY\:LY,&QQH B$2_405@'
P(^R64J$--]!X/JLEJ;@7[L\@4(H";:&F1G)*^E_EC.U<E#HG;@^UK#,)\OH9=R ^
P;-GZP6*;@ZG?-/=YT@8]A /6VSO:(XBZ&N$P> '4E[1AC_.;)D*XSOGFRJVA$VP0
P\PZQTI9#HTJDQZN"('0E!<,F RRQ'P81W1$90R"J(B(S[<LY%*1Y*LD)"5YO"RD=
P$QSNLW%L\:0ELQ/CW9'->IH;']4:<KAG9J$O+_*9%]F2%7H@#0\/3R>FY(8[\>"4
P0R%\+.H%\6N,YNN2B@G\*QN>CB&I46""R<G22*5! H-+B3G;K++!7?/!NEON+T[4
P!GYD!)M8UDIO98M^&_UR&0F#DQ!$(8)XHE7-)FZ##FS+">5/Y@8;UN5H5-[J8BN0
P6N7D[,AB&<5?;:YVM5O5]E#":]-'&W&_(?\!9]/__63;G;P0G'<<];2H@S\F+'VK
PLI)K6]DCDSK";GP3_NW-+LX#@>$MACT?L10-;XV$D.9<S-JV6LBX'+$A3>XUM5\J
P.Z:@!@Y9(QZ@:ZX6E9%6B,I 2\1R"WQTZV'& R/'< +D;NDT1LZS$E!#;7_1 B*[
P]^0-^ZNSQ$E ;9TA.97Y3:1H)UEC 5^Z!;0==#F5A-KHX;^M"18012=)N6UL\:</
P/TC%I</S.F#HG1_U%"N.$]Y4DAIF4:T8EA3RQ%SPMTE[.(F&Z;JCPRYS,07*L?;A
PBDTZU?*9UO#RC<7I.UJ?3,Q=N7>Q5!! .0_F'>4"K50)AW,W[^8Q$&,/R9H]Q#RZ
P3,$JA<N;J>J*V$'89'.O%MC"95BKC75T6TO&ZG48UE&464>QE#MKVZK5"!XK+9F%
P\->,^,F/!!@)!D$")7KGRQ;+V()X#LYOX:EH[?;+.J^T8\5=+-N^Q[&0#$J47(-/
P9[2(PA@=*-",)I]*:'3:@ L;*@L!3,S+0:GPC]<&H7T3=JU+*<2H# EI3DKJ>O< 
P'4,YS?<-:UJ_U/!?L65O1[989<G!'_E'*%%TW&@.UD:#:FT@MRYC,";=L(D,KS X
PY(PX.'/%<'Z#" RAY(<VIO4OFM7)01FT;%M3:E-P[/+F+7U_P<^M0%M^^7,N[.88
P/L,HTVS7+8"&OLY28NS?6,\7X?P!$W?JC:.O\GM>;\#*K;YN%VCD[GHU\2),81"7
P("F FQCR00X5HLH%MV@%*9NV^?O=:I-Y!G)B7ZZPU8A<D$P;N)13O>NA)<L_,I';
P8\*&$_:LN&&*IL<^[%;J2Y=>L_?,&946Q3B.+BHSQ(A&RBB7EA:/L7.:_<0'C:UR
P#N$#!?(U^5<J:SO/H1]CMI84$.E+?,I%WN&13E6#9*D'4(T(D&.9KN0=3'- ;VUJ
PEP40[QS"R/46VYK;8 E+Q-L[(YP3 Q&:*I3=R9HOQ0V>$;B_<=,@PJ@DESMZR '3
P:&8;6+CS<UDS 4^BSIR6/H:6.PHUIP]RF9&.U,#K>_B6F[HC6;:-*</2JX\?/!B2
PDGL'S,K?0X!FT6$\O/0ZLS8FZ;'5C)415-;D2]HQ,6:=CNU/QSR,C1SS(/C-S#H,
P2AQ<3DOC_Z=)]S$<IB:ISL2K6I7[ )QQ3/"4^*/G]B=]B6MH[)8^=L1RXX*6:\;V
PO[$3?4:9:P[-N,?>2M,"-YA]_<3)U+W)K"TQS/8B1W)KYR+/>_: -YA0)Q[W+]8-
P/2-F;,&2PJ_PGWJ3Y'SEMOO <'RY*@R'%W]G@$?;.IZ9+_3,HK)1J0AD)S3]7M%B
PX3Z+*5&O ILH>>H+GR[?1D:31M2KDY$140M8YF&/1RF(/(5?*IJJ?[(ZBSPOZF?$
P%3K 8YPOT#2SRTK /LJO;[UCI;76%&",TNC0J&B\9=:JWP>O)UN1-C9CTN3U3\*C
PKB^G6ZY-Z^7U.RNH_-&Z*4'HKK0J_'Q2)8D/@!+E9QON,45U\>1"P+3)NRHI56TD
P(WE>B_L9;AUX0C.E46P)E@OG5&SS D'RYU)V'%"%YT=<61#ZR0\'C,<NJ'2>>H0^
PXQBIW_4?@HW\7>7B*D?Y&[5">?>NW4++K#$=(0'E(VP>:IL4V?S?ON45JD<F9:K_
P<\INJZ_=$SDNP N"\]>5')0*\ Z#75*%9K@N2";BH)C\F Y?'/#BB;ZR3P#HP^@:
P6WW7?M)O<: A7VD:@10!AG9;N 0D/UL-?@%2EE6^',^D6EO#RK2V](@F4=72E0,(
P!YK1JY])5(R.OK4G6H@P_NF0 $ ]"H[O[R#7XGLS>=M8</G()0D6ME.T1G"D7;%.
P'">+F%M;LQP?=%S\=$H N/IO+B]1ED/GLDHA)NQE^ZMKCU@&>9?=0M[VS7874/JU
P 31-DF8T '"U?'5Y[)M/">KLA&;<3F5+N)4WC._4IQO)(-1)_RBS[/H:+IN:'M83
PO,K,.RY>%^%Y<H;2)=PG9+WKOFA&2*#K^3P/A4P= Y.,K5#D37;MLH#<YV_OIP)[
PN:VY0AS7J)&!5HTG_'M#"XP24'R.Z\=0A9O.\1>?.:2Z+JKZF=Q\#1PG'^J<>GXV
PJP+-8]0O<JGUX3)9!0$W]W'<!0K*U?I&;BV=%]C\G!:A8'Y[;-+'9[:?TS#Q7J5I
P^U?]'N($N7L>$+H&^!A$[WB.TNUU?>V)(YDCV.FTY5PZ,J^>J?6L<1?M29.92S1/
P_GE""$GZ #4F]E"(P5+JP:L #=D6C/*RFUZ6U^2LPU%-&=V.1LAT1KB[!8$AIVG!
PDU!3/<" (1[W?O1_<XR$T*D=@0#*->5=WM4Y\;*@=JUMJ!N9_/?M"$-OI[^;PV8Q
P53)#25^R!)9/&]5L"DR9@?@R,4[33Z/T":PHH(S&WR*6-FZ%H[$P]2<[!R_T!RZ2
P952Q5D'-[#-TX9U?MGUN#^4V_6&[-.)W9#O M8"H 5=VK==D+<$46M4./1:0C6-9
P@L0"<(768WV$VQU>I35!,V_-DJ2LE83F@H*;X;M9,<PZO,;#LA6/CPMO7= )9G'(
P]+7A=I&F>-,VA7GSP;F'K:/EM^D2>@.+2# T8F94X_Q&]=M'=BX28?\G&./XXYJ3
PZ*U5K@N(HJO+KTEFZRZZMOH1=@0S*XKXQP\5"U,LBXI/EWM;SYD.Q5<=@CJTP$@;
P*G,:Z\>W2]FM3'?YB7N#+BE-"C!!<!511M- \LH^<XEO]8 S89L691+PY8RK;CZ$
PI]1=ETDQL%40/R4<%RD-&;0FN?XT^=]JI8(,Y>G9X+6UPTG Y@D$36+E21*Z\%PO
P)3 6FK:N-1]^?]WW06BC!5H&U846++<7)TY[KC!D1?_>]C"B&<]<%@^$T(8O)\)3
PN^U^TO2U?Q.RFK[7LJI>\*5^6D26#GX;K][JQ58KYN5\R+799C9.WD)!.R[D>!ZV
P5V5;<4@FXMT]=KELYRWB1#6=]S[FC?%W]:;,^SS=(@0T<;;*Y/YB?N'80EB1&7.3
PZ(3:J[:IH=T)B KC.@971(-9 +OD:6E#I^#D=%<HF41_=OE:/VD]K]$MYOB?&8G@
PBR3I4BHP?:7OX'C CDE!,KS#>A6=\0<%G:$"'$RM1W>*VQLP2[/*E-;82NAXS^&1
PHS!$2ZS2UB?;3S1?83M1"5BD4&3O_T/DZAO,TONN1:>MW+RY6@I&ECD$VY2:MU3B
PGX>93Z29M?.73PWF\<K#5FPM'6:A!G?)IN8Y2"NU2/%$)&04TZ"<3X3E?(D<@]=4
P),-C8%JBQS8G34S7938<!Q!@17-P'=K#E(!%=E,L_>@=55UW)@D#^ZH>I[\02T_1
P11!+U]N8:HFS8&]":S9J.0V<9J[[34F'K1AXI[UJK4TK\!"GYQ?E];_)<4C#/HE0
P'P4:6<44-J-) L.X\9EE)_R8=,DZMV"C($=Z-%JE<H_IAXZ+F##P2)U#&$CX49:+
PN?,B"@:*$#X,7U.5I'[#5+@N]U5\4\M\Q_7$\5\HWRD5-A-,M-L=7L/^HW']>@NF
P:*,*G)_!D4CT69"BWZ0>[P8-^VU"$:N#]=W$TW"^^D"'9Q$VX3_6Z=P OQEI^05.
PY_.H,(JX8:X;"(WR;15( T/)P^0'#C)!T;Y68R7')HP0:>2(0+<Z7S M/\GZ2CTH
P*X(*J_DL,U;1TL]*G")J);6%-RUB G /7[:>1ER:#,F'<;LL4/"[MCZ]BE)ZV./<
PQ>N*9?#2?(/E,K@KY 06&R>VC!NF1;.>Y&)=8LM1P9H ^_"[!#%CRK%?>*T_0:4X
PB.U$47-WT0^!-S@_[]3R<8'V \70H ;L&2NEG@,ENBN"O=X80R.';] W3/^]9&JL
P/A((QA*TO&.KHL0*5K;9H:Z*)!.AIK[<F5EQF%A&8Y-A"N*QD)UKO-_:80[1,@&-
PN_3^KL#XR!DV(:VW8/; _R/7@O?J]M_/>=11)[R.2%NC1R1I7^Y"'J6%][:!2<0K
PG9E=.\7R("2*$$XTQEA >EA<R(6FFK#F_@3I'91>ZAFE7U' H6:L'Y=.=V(6QW>O
P8]5":,,;&Z(:ET0567)*JW\J JX/KFHBF8",,0%U%0:.^5A%5<)S*G(@Q>?^L9[[
PW,Y+&UF#IL8N)&C3+01^ZH"Q.- XZX;CZ$9]PL)8H>W1'M UF 5RJ^7,'4^G==40
PR9\VZQ;MU$*['!>O7JHMB3^*3I"3=QH_/&!:N$H?I\C-\.V86TMPF!.JJD3;C-&<
PF(*-$'MO'CO>H@PTL6TBUJ'X0]Q ;;2H0K3L"H(ADS X_Y%'?Q/[.(P2TOB:*LY'
P"(V-)?[10@J8WC)"OB),&F 0YW6JS/2*)0:=?ED%X?*J)M8AT&;;\"Q+GGY:"Q2I
PLH.J?1,:A6Z2W,.%0K3\;F6@2/TK!$GX8JNS5!"5\(5!6BFM5\>P0$E=?OHW@\^D
P$1N*V&<O2!,IZU[MK\1*5QX%V$XA%L!/^K"A.T(=RUDF$CO:6V?Z!%\J)V^;\$?*
P]]&./QN;P$RY.-UE9"QD,DLIDCJ&=.I(!F8#[<+#'<Z5@$JL@.-+5XY)6;H^+DI%
P#+3\>)^2?B*M%@^_E&A0UR@_4^@'M*D7-]A#995@>- %$5 5;F(\70L+I^4"\T*3
P#RO0Y/3G^)#.S^&;$AKHU'W"7!Q[MY>\A@#, $L!B9<#GKHIC[1)Q><Z0Z)O$A,W
P>L>TW1(F:;)R.L9WEBNN56,Q: L-Y>CQ4/-4@*LST>IVX4Z4/&FHY<!&!>T30V/Y
P=Z!78L8T$@8\HJP##31WNLQ-<B('<I.5#(9;<%RXB'MI*@I.M7&S.K;?A!3C]\<Y
P9?#)9-WMC+6Z0&H[5=,SWWTU8=8@&WF2=*K=*9:/HXN8E5*!7EM#KV:9K+WI/;5W
PA">K^??6" ,( ^ )J_CL<:R[/CP4V]3-44,^R9DB;8Q\];\1AUQSV8KS4.Y\)>86
P!8RN:T&C4W@:A^ GQ=.K@/>:0,UBTE11_.3&44RH81#MO=-CNO7B%3>I2V 6FB:E
P:GB9IA\V]7OH9 %CJJYA;9S%8\L;QL-$<]8]A?Y(>Z3^4VB.6$I/7&@)X;$JZS@'
P2]-+>P>J]*:OG"Y>FV V[>P6M-4NK^\M[9^KP;W[6%_+BI*T,21QV1:(GJ^T_$/S
P@3EM7E9/&L)F7W\PG#"4P+N7@M1'\2APK]X(BTWHEU%QQ#_+5:8,9.7;#T/840."
P@+!UFI[)T_X1S/BB4,@*F;0?\5:S/GV-5=%3%.*-"Q[^WQ?W<1X!_A/UDI=P(D,5
PR M[XO']*ZU#:R3]/=PB5 *KSX;#'K1(R@2^5ML]6GF(GY](#'0IU4=#[E:>;-38
PWV[]M$1>8>[ HPU=*&-7($EB![E"ZI ;KBW&EYY>2GMOBZZHTD# [WAX@%+[W]$4
P)3Q04J! @/;@9'96#C5R#;Q>8A-N);BH3UW]9X"84^-^X.AY]-,,(0(48O.0\F(.
PZ=:EYAZM9.FM5&).@T-\'CLZDX[C9^E\8#!OH>M&(.(;O%>B!$4),A3JTUH.11)%
P-=@3' F+UADZO0MN#BEC'^!VR!;'/8T'F-TP=&=>1H.]^5/- @14*/"WM/M)/HCO
P%V>!@TRJE%")<6.^0NE:S9?F]&+BOWPQO"EP*UU%>U4A6LT#UK<AZ3SQ"5LK-_M_
PH4/SO1'L7X+T62^^4RF#]@<2VVMRJ Q-B^72YPT?OLVGGOJ+.PS4#UN;OS4CF8"S
P\M/+;0G)D[T&\I";L0Z3?UTNT<F2 =I54<I;P5FTX*D"IM;0W@MFPFT+"5-&+*V$
P^NOE*_"-YC:YI1JO=[[<PK2K5"'RMN6L*S^8M8)CIHT0I^:T'W*ZK!)9/YV WL8>
PB??Z[0T R\9="^,YW8A=>&I)J_4_'>NDY .QYW/KJ-PRI>M.:%2BR#X:)7DZC9EJ
PP<I&H>=P+A'5'9)UY+C ZR"<P_=:'7;<9.%QKV^L5C-%.2@?!\Z5T#-??M<6.($8
P4PX?=S6FV[+YQVT 6,;M*N/E@-P7)! GFYPQ0G[\D['<1_KLX$$N#UGCE_N=8H08
PS8V_EZ=*<1L+H+<0%?Q*(X ^!WSWN6DS:[,!^!SP'10F9IKSNHZ#)8)1[EJMKX__
P-C0AJOON<)R7H=GP=C5*$13<-.UO4EX'75132BEB8%Y""@AQPZ=Y#$LR8&+W]C4G
P,_2$;<4IZRH3.#-83LE4O=1T $)3\6HKM6W'T=M4U<D@#%M^N]#W?@*-8UU+^T U
P:Y-CI.;-C(W7#_2#[+Z\F.IR?!(P"@A86 AM7AZMV'8*N$?0@3!)?S+X,2X" [O'
P:MU7IZ-K26_#L'O#6];DN!U1PU*#PLE0TF\P+X8<JH^W_42^K&&0U3<%MC'2,=.E
P=T7B!&U,>G"%XZLE?N&X8B5BH)ROG\7PXP@V+UM>$!]OHC"?Q"G)3)#NYXNUFUX"
P[[6;F7)=83JI V@XZ"%"WR"CM#4)!GM8C;Q-A+3R;3/E#KS5'[[E 6$<PE\$1?R;
P =^K!Y5V]D#ZW7!94Z_D\VX4DUX#E-;F,-)#V$V[/)I5ZIX=#)R7"6O4G!:%)_S2
PIUL77"NCU=Y%B"4"&'*NLK7_GX5!<W)MM  G&Q03I5 1/C]T,3 #)X3D+@">1A&G
P&?#PQBFW9-H[WMGJ..9#6.@KEZ*##WYY1[<1AF7!.7OT1OF_&%E;#N>12^H1?''R
PW)ZSKW?E3  3*RU JC/7 DG Q:,T.%)6P;1."606-9WE_IF,8<6B O53AW@S]=SD
PW&#RGUX+*>U@L+6E?N5+VXC\34\ Y702T[&S7MKPF-A!%=L1<KTFD5.9)^2ZG"J+
PN2.UBQ^#WURMV=UT%N2^U!EGUIF/*]&A'^2U"LK!EZ2>SQ,,*0->5];2V-_;>!IV
P6]E0LINQ,Q&SE&NN)3\&I$6+U9:2R6Y+G_D@UWC)+L3L,X#"\$^ :LI=B#M)?LR[
P6(A_DD%:(EFD^>=B7LA#UESZ91[V%7D*[.NQMBTQN1XT>ZT?.3M-0FPHM<7TEZ$%
PAX.MO7B,_L$];H49#C_ I)/#VIE8%/S;<3I:A'T).H[A0B ^FK+"A5<U-'F8>795
P.0PJ9K<,N(;I,V+G#H2\,: 1,\P^VF/)&=$V!#8N?%<E7_@+J( \[Z% 3EAC:O#K
PQ(L>OP/YZNPX^*1K6]^%UUJ)'KGB5(^(_7>UF]GYC2U=K0%*F\$ZPCX9FD/'1$4I
P9'*G?9+..*P"UHX)(19_<N!9($^39)W8FZ8&ZH,%9Q:N*-;$]T6*-2 3JB3=@-D>
P-/DY<)V^RYI'SZ7D)5<$$ CH!1H73M?#XG""'<#C502>(T9JRO4T]GTRB]M&+EZY
P;$#7G0B?3LR/?6LO=FD%8>1L:^,5J#Q/"HSM(4$QQ1FHO?(#39ZU"V)>9VO: G;O
P(L4;$LR:*]E[SP,^G+K"=T B*,!.QB%3N%O_E8C4_##94 BL>&3-%G=>Y!R)D N#
PX930,_2?'R!G*W6<ZR:LDI[JCD\I8=QC191S#=U2U13_4(63IRYH>]+L]'PM"D)'
P,?!H/H!JO=_1Z'SWN</W9(T\R&U70/=DR;^"E@_2T+O;V<-K>EW3L24]X.LJ%H-X
PMBXEB>HX8GRCI2I?,N!D \6;=UD$O1W?[@96CN/LE+/H=_2;7%5J?JC9N0UQ.F3J
PD:G)&!J&Y+*?V[NBX@]O2W&I$&Q@&O/C**%2C_FY^ISKEA!@))K<T<G=O\ H*<H0
P.S? DYKQ8:)\70PWMFZ#>O]CK&MHS*--&N :RI/!UA]D2#@I$W"0N%B#N#??JM .
PT:Y6C6X:RR_MQ%!Z_==DRK%PT<;TQ=,?S<,WC$44KN#$Q[SU=-A<;)J/FSQ9P'[<
P!]^(02W^T<ZXGJQ)I)'.U6-_O\#C^L$P<0H<=HM F]_:I>_I-/)B[2(T&*<^VN>=
P']7NRH;G""99KJ7A90_D3.YW#\22;I40B[P!O:N:2YZRR03K?"5L+;S?&;T.,8[(
P2%(LB'^OIE9MAKP\*IL#;_).TBCEW6.@:<#'\,RYQR!-"?%4#2JR3W$,YAPC_@/S
PYC^WK?ZKN)45N8P99 3-"7$XL  RL\\XT.;(\TH383,]TLOMZNCC703JI()M3JC+
P/L,_$LFK^E%4ARUB?>?<-PR&LZ2'4B0>0T3OC7/@1/\>J'-Q -0R=D#?P[QA2"O?
P>NJZ@^+-;9QY3U=A:ZI3LY3*<WB;#FC"H=L_A3<;&*<9L,G?B"F T(:)WVXK7;_6
PE:;8&LKN@8VLS2D64.,8O@\4AE:J>9Q6P*R<Q$8Z>@IBNS$SDRY2")U3=M8*FM5Z
P"C>FI[WWN>[N0S@J^7)9?Q8!)D?19C0UR2>R)#@'9!,-_H%#[_UGWL"EC8IVB-6L
PT,)$63#^2X+5/75PSU20^V\9?P6")+:X7(.3J0>ZGC\=6_8>*8(G36)6G\7K7/"\
P_L9L;_3FO1:5&EI^);(PL.@K'Y7_0DR*2>6T8?O/[S..U=8E8]O[:R27OL,PMA$3
PG^2: A#Q-=++EEJZ.3R"CI6>3Q<VY<D MG@/=_A:IT=W*J+0^Q )CLPF6X66'ZG+
PZ0_\)@.>KF+8A@$*<Y36^Y1;#N'<@Q. 5*3F7GEW<[7Z(TY;93"?U8NA(4'JV253
P^%USZ3U6'4P0)0Y<L5G[NUGLJA'%!EW!I_Z1FG&R=!;)XM6"=W>7JG\DB.UH\5X^
PX82ZL4IY'CK$C0P/RFE@=6U<YGP%6)/8E9KND5T>Q!;;($&R0:2_J4"D9U[&:^Y<
PS!Y4]EDW("W/ZY_4.L#'V RP.(\I*9XG-*_F-+DH42ILV7$H!2\"P,=I#N]BB9,#
P'N\&$_"),SSA%3$T@P!^S*S0&QF"GCV[ZW%E^W$&!4X4]LS)@6AA$-9#>1H;,N^<
P0M^= O)I'53*\\%LA2-'H_3;G@]+*!.2T'?M,O\BS:@DG$08 OR?/,.\*$ LB*(0
PT(9D$-:(/%&I3Z;"FAY7W<2]RM1+H^Z?_.C$J*L1? Z7 55G'AQ4?;5<C]8/A:T#
PV2ID0Y:*Y9@VP&(.;^U:9<3)=DJ/F1Z+NA-P+?XN-%"7@IUT&=UL!Y'QQX@"!_="
PK55S0V.Z*@UW0]A(>?7P U\+-OZ@?!$L76<:))91J\6SL6U#E.472P))-]671_&>
P"NTH3IS=R\N,;LI24+T><E @@3,>5^]MZ>*>5H<-[JW*S@):?-SXP/OJ=WXY3K^8
P+ .NRJG$Z;&-PL?YB,;11=HNC\C(QJ/7*(,"LI2ETW&%Z)9*0S&(-IXY ;\:I(!N
PJ>OK+T%Q1-=:!MZLM?9-.W=E]]S<F4/1$$"=:^+S#&6?M!ZKF,11_NG<#"HJ4'_5
PQ<&5"GIGR=TTF1L[:C"3H*\EU%:%&Z"6QY*LXBF[\R=U=NADA6HB];F[1T8F#]8S
PEO9@L!>.D@/$[&81IFU'T#(>[RJU_CE!\OZEU;=8>-3 \TDL5^0E )[5^-]=V/C?
PM9[()"M11$]&-??1%!J(:#$%99-/4'E!,M/:I6],Y5331M5H:O:E+S10..KO_I:C
P]M+0[Z!VKT7^R3+5?0F1U3,2&?S<5SD'M#V8TP $+/;YF/G6!HJI6UKH(F2R5"YD
P!/6%NPGX>1>E:P1O7U,8WL<7<?); V3A,(J29 2,)C+<&:?>1%>9.6 P@O)-_;]=
P7*K?FN+BX'>ZXC:3! 71\ZDI!93W/50OJE\IQV>1DX3A&#E8T:H@!SATI)1!73%S
PNOO'A_!I%8PGFCJ8HR$MOF*J4+QA%@D;G"A!$LN 2I5J^WOA^I=(V!M;#JFQINRS
PR^=.JZ((+]*IA]&*RM0$FK)(^%9]K0 %33-?N/8-#G-6U8#YXQ9X0GSD?U9]&+:@
P+N15]#JI2C0\2%B&OG!163XI-N3I=E_1OB;WJ,F!Q)M=^!<#2 Z5H,(^KF0O<5J+
P5IHC<-ILY+Y;#5>DE< 69!]F'9*\4:3YMJ5L\3Z=C4@-<+%8M&007SDR<&\:FVJ%
P;B7;<_$4V='UD<F8.>#U35W><*P4]._C=>D)G*K-9D'7)!^@<9+PUJ:BEFV0<E;F
PC4:QI,]P3*"1:\9^3V)MCL]X>\=;Q8$9;5W21[]U^,$%]1]=-6@W@H!H>?W> F$,
PISZE='GH$*[2#6K<1Y( W2/@RL37P&FO;BTF)Z@VWI).MOC6A6>Q%!0I'1F'73NN
P).C)DF_X_MV;UF8<+52J3*O/ X46GUE:?3*5$D0-@!._&MO;"J<L4&((CZR(+\8<
PB19VCFYBQ.0WG>4SY1$>X?J(ID3M017J@[++K6;.P+ A3WT9'2G#(B[51%L($!5@
P2]N5=UH4,6 -!WUY+3Z7*W V0A/):8]4U?@^VAD06G#[R*I;TU*X0M/Q3D#JT4Y@
PW2#NO<QGNLAG!)8_=J]7VL;YTJ(_Q $+!F%JP!8!T0O3,Q8R*4Q>%/Z(UN*VR'K!
PUX@VO_JI./08Q-ILF'6C+TC+,=2M"8&!.6:K12>ASFL<!F1ZFOO3M?G06581!O=#
P!!<-M<,P450F"#PT=[BT=-WW,0PZ#1F?3)H$1B>?XU>[F]4[U>(!,P\#A8F,;9*H
P]*0O>2P;-8:+W]'J4+]@,?P9!BT-L=8ETYF<O,/16^AGS'>-I<GXVQ.]9)]8ZE?9
P"(_.)TT(3,Z"R8(H!@=@?QW(SP*GPTL?MAXOMHM4@]]+5I7_9LH'6HQ$!\9@9MA5
P0*:L@-5Y;L,@K'K8+9F+S*IH5?^/-*M(&60O&USJV?9$B$\ODH_P?, OZ8:FR?Z/
P4;>@F;5V5!;?6FTQ,D"[/V!\7?(RS[X12!X7ZPO]10BGSJNDY?BH0O&,)%U*N*?&
PQ^/C:A*;HEJ,#];?2B&QCEQ]9#6G;7?7%PP+)A[6^$*0=/2%(NP>H<2"G=?=\^UT
P^"C\_R9)R8"$5Z3.%[D[GFIE#Y]H.]<9])QYEO\:0)_DNA:I-'GG&SHD%,8<&1(R
PKW_#R(./W* &%R]QSOF)<V*^UE"[4%\.7J[L07SG_<W)(#LV#41M.9>J9 (\G#6<
PRL#AI"5()X>,X,<A-&O/:'C2J0*K/UV%.SA-0PQ,33O5*>WLTG5]WNX2<25O9,QZ
P?:(#GN*>.+Y2)=;'?MG )#'>4J;@DYJG!0IS+0"_A/ M4KRNWF'W-?1'?JR!,<H,
PU@1J#Y%F#50A)IQ0:4Z=".J*Y+\/[W+>Q5 \+/EEJJ@<Q3)"U8#O^'GW8'5Z\M46
PDM&FYJ_-&7U9XP=,QA6K!APRB96:BO)-IZ%@6H2;82MR@=WK(P%H)'X53;RJR,/^
P6M$LQ=."(F9MJWD(?TT=(W><:A)=WKHF8AYT_EKCLQ $>B+;_/G2&XUQ;)G>ZM=4
P)%"3JY\!AX):T=O_7%$4/VJ.]/TJ)*ERCT\Q5<.R>QN]_BEQ)ESMIA=].:$JJ,H/
PWGN<K6]](4[M]K&%+J&*XD:&6]-(D+@S!*Q204\N$@%_ #U$ZD_]+#9.?P10>98^
P14?*%5URUT:6HE5U+;UP6$>=68-_>9.]&F&&U(Z*FY+6+#FU3CW&05ZSBVDG=0GC
PAMC=79>@=JS3^.;T54%8)WI\%"6)"!LYI2TG/!F:.:]#HQE5A*EZRZR"C+YC+'T6
P,I!?JD,+;X31^J]DD1QH?T65.W6&):'\T/]S L/U!&W=G:R<J2.2D&1VKF4\S'Q,
PH9FC<(J!88-\/DLV=F-=UVK>*G2 ^AVM8 *&[5C+=4%A#:+>K%1APPT)>'?2S!:!
P24\Q[AN]O43/XS5<6%!O(Q5*.KR+FMBJY>R3&CV$.!M$O5/, R\\J+R^_UU"GB--
PVI!%I&'K-JZ'D(\3G2J+'C/=3T.7F&80U_E9:,O;;(YB"BJ#NXD\&+,N-6W*E$6\
PU=2?@%&G^K83)U;("H*CQ2DB@RA)M-N8TC%3@[(8@=DB*E2"/B+BL9S;Q-@@[.8$
PU/BE#T=G][Z'%[3\\LSGZ])AQ'USYO/,VS2$F=02[/TM2&"=F\C&%.6MD>=L]869
P1V*Y%8^VTQVG>:G'!F9) Y'D-(L;-M&Q_KF0;+Z09@DY#"ZMO29E %F80W8;G:XF
P8>.5^[.7EZ7$V]R.V5$)@?+Y5@%6\\FE_630F7%"M(#1R@=UMAKCJ1^6H%CB%SH:
PJV:6=QO^Q5(/#+7AF5N;>4R4]5P7!#>@U4,_$X)0R .%+N79"10?H-13D5L;4_$+
P]-4?;*<#0AFI6Y1 3\*R=MI+$]K:$5,U'WP' EEZ1!#8F:,_[[)+Z4)'$#=/#<=@
P'UT8$PGJ<G/MW0+;YM="!U(4XF2B6D:]D\6QS=E2&J+[RA3:PK5!VAP<%X(@K#S*
P\\E-%/APG/@E)U7_>C['"T:;LJ[J_XKUA\EZZ',GR19CF#G! (_=%:IF0^S W<: 
PX@:-_Y& A#&V^'VJ*C<T)Y@>,;:[.<50%S7P'U2*9@SQ03QQJ;B)\1]P#V&#@6!W
PT;&W-A9Q /F#]X Y9.5E#.8="]MY<'N)4LTCQEK&AG(UU'7$4'3H9%1I_A*F#YMP
P:'.PC:7FLLID1./@)P'>06C880?@+%6!DHR[CA&!QG_U>KM>+VCRPY655HLTN7TQ
PB'UTQ 7^FR$L;#?\EH<MV8+T31*$S@N +-^>=G3TT/0=Q>OLG0^G$IT6LR"3[G(B
PMTML5-)W2/ ZT\"'IM^#WWVA;!1!2CQ6A?VU<A0,?U/<A% ;PV0H9,3UZ&8' %T2
PR*_CUY3K&_5#"NR7Q9DVHZL.Q/H8/!4B3SI@!_\2;H;5LDV4"S+IO2=@UU>RAY:'
P%'#AE9*#R4?Y<LD7WF)\W/4+8?ABMDV\2FOPI(R0]<*UUSR4C?KP(%"E$AG_)WNY
P"Q0 ?8D2$7':\8U(:OU$S;J_3.CHRCT[-6\C1B1D6EQ.GOV+BCJ$;$VI<7/1TDF4
P!&(\#/. ("C-FO?N" _0IKB.8\]-<@ULV,$"@DN:P8Y4B+:YOWY)I[7:YT_$?(&/
PJV+!G08S3B7PX8MT'TFU9G!(FU 8#CK==Y0H6-.(H7C[M [8+XASKWA&<YH!<D\L
P0)%PPD%]OA"M 0-.2&NLNYWC[C@)MWJ##Q=7>;E;3\;DSY09&:%Q85EMZ2I7,L+@
PUA!A0X%Z'H\9 G.(>U8)@S5H+QJGBYGXVRJ-N\@GPG"?" QLM#@K@[9=5<?M80V]
P!IO:0X?)H7FM6DYP]_2;3&YI+**GM:A$!ZW@T<.JPPK6.HIIDB3UO;@??"NN4JD9
P.U;Z-URCK%T&(@QZ@!<'V5_O>@R\17"WAXBI[F@2%XG:IR9DV_GI=\S7*O<+310>
PB2ZR8:0._6EW:O?N+@Q9[SS[=,+*</:;U[ILH5^_"T\TGZ]#E RW BQ#U8B37HB2
P$ZF%LAUT@)/%J[P@P.8Z#)/U7;O5;:9Q%?_P1YPX/&'6A+G*;V+:,]##O!<P#3CP
P"3PA0&IQ"NT;$IT,E# #DPLN\@\XSJO4]#BRW7#7TIJ]$OA.^*!'8J![\$&RM'K3
P,L;93D8GT_M".9176!<T'3 C[TG+L0+<-/6JAOD_5TM2(6Y*T7X?NFO2 $V"[0P:
P"@Z XUIMJD&X2 ?XD94W8;). _#R&(I*-8["QDO(FRV0L-VC'"VOML?PO<[A V#Z
P9DKYGS:K2[<X1?>;B)[W%<=-RU/0SF[Q."VMZ%%.5"^I#CN=VQ;AP[%L> %IQ."Y
PK7IVY/>A,3U.&G0>/W'6^]:50X"9#_MLSEKY/ZY8U5'=AEPP;M\JS)^-_,U1BX1M
P0W628^41>6 )AKYS/_LI:7W^@IAFII#/;.'$V8]<J(;+]#L://0@>F-0H^2H#^^H
PM@D9BOQM$<W\ 9WU= ?4=*-AK.Y+E@T[Z!U#DV-W<WP\#?[@Y4??+NIYR%B\_H;:
PLR](NYX?9!G$BO3].4<9P.KEE*>$.PTTJ)T'Q*5[P+:W<,5S)>F\@*>YYRT_4^/.
P6.(M[42$$*BT=XB<3((@(E-A#V:A$[575MY"LCRPW4J%V587(#6A9^Z[7:K+U:Q-
P*4S+^LHTR)ZQT.LI,6I:C>M1)=8,^'2,H0LTY$[*AV_?@KLX+E[T)^_P+%004J5[
P))\?O:A-6&-OG<0^'#-0!N'+)MCR)P :$ED#=DFPRZUK:Q3!7PBC<ROGJ +*23&F
P!BG>784ZBF1&V=A+=)0T>KS%(IC$P*@QFW:+U!,>:7).K5:GR*SC[_C:0S#4AL=F
P9MPLX^YW<_0.?G,''K'TV((@OW#"?,,4YC_)6:>&N'3%)D;(K5?_ V9*1R/IW (=
P.XC0YE@ME>"@@!/32L-HR' =#C'HIBQY36V.O@LYF'W_OVU'^_%PMMFI.7X8%K&-
PH>H+V5:"/.*N&L8Q95&F0!-/)\I3BF1GN!H1,,\SV H-80I&L"?6L^O5["(I8Y7Q
PKEIJTE'+90J60"D%?*;<>SA,(/HU)=MJ$3S0?,5@!X4F*5(FY_OQ(PT[P5(G:<6:
PU+K</S[3;S*GY\+93AIK*QIENW?97$$R>XJ^N2[]TMN*#F22(_!P3P%_!3LC3CQ0
PNF'2\X1 .L$AM.*G"<%D*S$-5*>J@_#D++QPM?4#6 $<'&)_SN;G\Q6!K&KO[6WX
PR?@CVYC2!-J@< ?-K$8GH4,ZC^&7!8T' J-UG_HXICA4!93]=OG8PIJF[80_4:B&
P=<\5]/$R.[CQ90;",=Z^YVJ,+&,*^Q1N&=-E7;KOH"/$-[XA\>YNMU@9--*PM6/$
P-XW6(:.6S (X.G,W>>HW;HV>W3RG?UU&ON$#,^9<>&(?$?M9Q%1,O0/YZ8901PSC
PII3(MI\^8Q VHRE1& V?J([;>U#K(.[&W"MH*")S&+.4;.W_]/-0-M%4>SHZZH'!
P3[T$<IIJB.R(5JHB4LOTO:92:O @XXVJZ,2,:[5@X]^<Q,#"9WS3?K:64KN@LY%I
PLI" !"9?%L7O1UU:^((M=Z2XCJ8]-9(F1U0IHS+<UCC.W]=#3:3ZJE_"EL"Y><H(
PTMCNMUMS7%2@K?E1GA:U.L[JH^BTKGJ4-A39HC!= M4+R+PVN+IS>#^]X--NC:7.
PC>7I,]%>^C,^9E:?G-0<BZC*:^K4 4;SB23]Q:(KUH5Q4#<2^!_TP>$A3<<6L/X.
PB1&1F653)\5+FG^L7J>&GO1^I](8F%IGIR]@4RBRP6"[>X)S3I8TZ!G(4/MZ8ST<
P;V_4QNZHH:USH?/I@9#P-L:]*/I9[LB#'TDC$#&@Y%>IQ4S#LR9EKX<S4WYQ_ZWL
P+/;QTZ/)7+WKW<\2[Z]<PXI2 ;:*Y]4 AZTMFS%"-.SO1KBE@?K27: L@#R<1^4^
P0I5\ (QK;&H.D!-L5M!PL- *)9":<4?1US<O#I#]T7CT,)SG%Q-!%L%B^?C5"FG-
P L+D6 E9X]KY\4;]:=DJ^[G#15RX1 [;R+<)$&!M3S MKC) *.::_9[4TA)$.11'
P ^5OLR7<.[A!#8152\VC';!GO]/AV->JUKMO5)5KZH&-Y=M .>G5G]]@70@UAVU?
PZ/[)_. %1X'@$6+=P!B_398Q,!PX0  /;@RO02(G5*], &43B*<!P,%))KPW/[FT
PT%:FL&!,QSD*16R7IV.,(T^4_> @%YJX?/:G!^\1J]COF/ZGL<61X]$2$4697#LA
P:!D9:BF^"IKU^XQ4NQ0'Z-0&*[X<@>DP'UFTX\6G:@KP>Z/B"8Q$FGG5D/ZY;O7W
P_%^+66RJ-(LUA+!8^XY]6T#!=.C]6B-EBC292?.FWJ8(TH']0*&!)46,L]$MO8?!
PV\_<Z%,D?%D)<A02NZ3'<O%/PDI0:-7T3*>\GV@?]7!A0)[YY'[+L25W)I5Y/*ZK
P4C3YRC=3FSOSNY;U<+"Y="=DXAVEW62D1UUB!./F4,^H9]@C:R!^K=/WI*<>W7QK
PR37AD@=V<O*+2KGBA_M--M,M+!$4LZ7<WWIK%K!LOWZ6%A*?2FPW<>*8BJMX&A>6
PHUOI\Q.X;HO%W@OI<I_$YE#-\LU8IZ +LW(,;]/.QM>4&@KRV5.F12P_&$LBRFLM
P0E/!2&W4BJ\BD?S*#11/2A@K)EL8G:OK88\/_9*Y^*W8MR4=[8,?V+@)[GINF+4R
P6A4UQ*X_F'> 6G,\:357Y7T-!K\K(&5 "6WJ6U4K(TKK<UXJ/_:_]VL?P?_(TG*.
PU'KO_T5LX7:7C;S?0,4-$(>'VL"7('E/"%5=8(Y?4[4F=<%AYB256%VJG=4,A_%$
PBSX;%W+^J8G-*'BEUE9379U.]'N.<L&FN 4)&85(;;GC*8NL?0++NY/G6Q&O'CQ-
P,I/R>4TSM+R6).: Z]U")V(CY:[Z@:_ !=!KZ0.U%%4?DC(.A*L3Y+>!_:JO]BKN
P>D DAE;H$@O]J67==0^5+1WBR@JF*SV>(<ZLCXT'*1YYL]6<T.&JF_X^GU(70.4A
P[Q+0?[&K[6,1O [NB7-GR=B@^7:D-Q8D#Z,I(<F=/UVY/0YGP02$VNW8%/-!3\Y3
P]-<ROP3$W^/Q 'DN2<?/;1QE)(PGBS4(0$P\T*6PR1QU^ DQ#!4"U12>C%AXQ219
PZIA>&E8-I'UM[+2_I;SLN8PW\#.O2%7'9YD?%:C_\&9JM)DCNXRMP6:..: )HKD_
P/3[EDG+22)_-19VNM<M3A.,F-Q?5<Y=7F4-IQ(%U2VD=A;?")M)$T5K[>\0O>6;X
PG5%I^LS0H^=:ZK"KR1=)GI6O]$9MN/^'0=+VSO/Q%NA;+,!=Z>[ :ONDK?7F)V2W
P>< LX91"8.3\<SO=&]Q,+:DJG'*KUC/D[T2F1:9<G>$]PE30!W@3B'.P^(OG?N@K
P%">*F.K-J_2T.(0!O/G^_%7AP&'^KZXB  .4 /4QD4XY12ZUQ?D)O-[=-9E'B(DK
PRJA/I]?)QG;/TV%7Q<EQ#)$QF]_"^SI^;UR?+)L7>=G?R/SUN/?]U\0'A$U,3JQA
P9(YV&.D4X2"VUJ[H);LB\7;(_]*V6L=T<8SAR;]*3ELKE,X8S9RF-)3J6]?\R8:]
P2R!U,-)J-!7&% A[HX+,$SX#XB=E_!#)](61.P814DJ),%?'CT@GN236^>]=PN99
P8XHG;,>R1Z>WG2U8.GOVU%L@M2^"G@NJ98%&F<$6F5R@7E[,7XX(2A4?A)U'@$X/
P*@ YBCL#J/U7NNG3<DRH4>^[E6OAB50FNU( X2);ESTA=OU[O8$6MP\LY1"H #\&
P<?PX6'#KDAVBRG4:;H:;TK69-=+BFF^;Q_.;0EA)GR<5M]U$1KQ2G^@E<(':TW&6
PH\Z5/8"/ $-_OIWI;02D#H@Z!=@9>DE*@_\8 PSL.AI2*C*$+M7XU4&1-8J^1$0$
PHGB%RF:H:*1"^ R4]1!8JA&4"_I.K.F)LC)I%-F-*(^/]LKSJ*R9)A7XM79QW/&#
P)$--9DBFTOG =9;%'XLV;L2H8R!#< 4%!0B"L<G$<77O4*W ;(A5@&S\1X#IN);Y
PDKZ:#E*FNT"[,[,H.?AJ)\;YU[UEE>BCE=".F$12JTFFSWCJB^2]%8. ,IEUGYP[
PA3%7N9DW:E>7X)-+_M53WX/\T!?QVDQ4-S>\Y-_!O@'Q3'RV/\S<5)[EG,HZT%+T
P0\Y/XIJ0"^O9CH]VGLSF$#0%$$8)&W$,8,'Q%IPHN,;2FTB-5K/JRZAY/Y1P=A"M
PB;6F>G_)1-[/$- OBH8N50FD;C9/K?$*!,$#N@.G=:1LY,8,.?0K]-GV+- ;\5OZ
P@&\U%7'!6,?^B7:/>,<\=1= !T@ Z6UD7P/ [GE:A@&N+.?N9+H4TF&?2I!+VNOF
PCJWN3&&-+=CPKQH3+J>Y))J-"\+FDS"^L1*;F1*0@I$:.FYE?5KL6::Z&?X.DW=&
P0X-=+@+%A'(KZ<OC.N6B;#QJ^(FS"T91A/4NMM;@M _F<P@GKFR^4\-RUFZ>7"$^
P1NR5#Q5&WSW[Y%0E(6[ O)5S8!Z ^()KT>V6WEQ],*COB W1Q56&#.T:^XB6JMW&
PR?;4T#$%->55Q8LF'H>6BI_)$*^SN).=@1C"CZ!J25*>W'IT%<CAI*OG-NOB_[@N
P,!_&MVKF*.JJEJ*XL14.C\/QE,N>4N*W+";XZ8SD#J*0M$!B.-FZ$QQ$85Y'8/.I
P!@.@X6I6D&AS\:3 .49:F5\$T$#M[!7Q8CY Y\AA6M3,C:7-I:6%*81\ZF-+'+B=
PQ6?/]T,T5P3Z%()N2@O!K/7V<Z;R-[ZH[:G'%XQ895>*\TO^7^ :SL#M^RS;L_W8
PQJR(TD0SCPB3]';2[:;N7,PM[9 !3FUKR NZM9]GB#JEZ &3ZF7(D8ZKU!'=$D,I
P8I)"2!UYCNK#[S0INK>,0JE.$[@:1LP.Q=2T6;(A(Y3*W?V "1=#=,3GE9N!$H^<
PT+)YNK:KZ4M<F-%>D+'IV?PQO[S0="$Z50'Y?:6@>/@>QF@:8+'Z.[55I%4QXH'(
POP^7?Z<@7EVV\8?O$"ITSV^?XH\[O$C+Y63>O<@.(II#(^5+8C(5C4:KU7\\Q\-]
P =(T^AK2_I\UH^;N$\$GYE,%5[ :W)")U'L(]2GV])JN;1?ZCX5H!HIGH0PB3&#L
P%<] 2+;(6/GLVK'Z]^_XU;V_44*?<CA^B>43_61KZN#M+*H%E!.#16Y-'0!63MRR
P.Y3F84FLR;N;\IR*QO);II;X1UC_+39903U?E):2,_ )$O6B4"1DXWQ.,U2&9:6^
P9$5Y<9[?BO!LZM#]V479[#.<XP@Y-&M4%N\3CBZ%#MZ1/;'@M7W("5J3AXHJ[1*+
PKL*S*+I ^CX)N5;#HAR;_7_8-6B? A-0/*P -9EE('7S*Y.*9 ;\D%=@52M^QON%
PS0,.AF!N*($GX/?2#DV_[$("J% Q%%B5%_01)-C3(H/F<I$0J,\&Z5B7?2U E'65
PA]RP*-HP8'9;FFZ(XIY=Z^"O &[Z$K%'.&P@%%NSR$/H7[0$)56\!H]]L3/56'WS
P;HH/ +18R4GH)4$;-'V".].MHT^U:1\ZAK.?M'?G+C,.!X37'MU'Z#T74-!UH@2"
PX);O Y9V&QN/>_#,GV[-VECJ!+]E(#Q<JCJ]!^)Z0KW1#&DFB4B)(T>0\I"(1TA&
PQ+ZSZ.(?&9=EH5 %.]_EO%OTB,U4^^.$ZJ5M#=[Y^4@GSIKX2.T,*TON5Y*7WQO9
PQ3@6,( CGG1^]%!HA^K=_;27X!H- *^ [9;#$"P?@<,&O^DX%1&CTD:B$&U6[2%S
PVCM#B?(KC"C7>2SE>U+@U1&3Y1%$B".IJL^V;8TL?S5X(6IYP;T]-]0M_8W5*RN'
P.B^/)KL(*QHWZRJC3P'ZX2\1EE[RD"8&OE-VGMXV&*3X<7RQ5P;-.9[V5W'?M4'/
P_1L839*-'ERF"F;D%N/?2GB&;98&+-0LI59YMHLYUR:9,,PIX+KOWPS&LASW;S/?
P,$>,QWI6 _HDOC@U)9%26K&P5'[+')+6([V>(1Y1#.D<:54*Y^1\.M0()G8)_#E&
PT=JC'GQF%3:H4/6NVVC'?K0?7.)8.[919"!2W!&)&G*:)Z6DWX-OWE'T^L)O^-)Q
PTC@>[^8#4L8RB"\_,%<YL^==N TF4YIMB7!J+,;:K_D0QR$&RP.5G:R^,!GDFV9Q
PO):PCU"7S3LS"T2YXX'B)@&]&/:>A05BRG??26QS<=11%SY2WW-06>.?AQZYYD?I
PB8< :U/XA%7F0,F@%RT6T-Y,^&JQI&_!)$]7N4L"\&5-J.^.21ULY= SF]G"?,ZR
P\3 WX$TF!<<"KUHWO)HGKG>BL6=+X0_N#UVMU;LL\!BC,IES;S1RLWZ"B @>$B&O
P79<%$684*BW1H+$\'0$$I@_*,A=^>8:TK)=L\2:B&IE-$9QV^\GR *1X&$QX)9:6
P6=T!<]T\-+/5L@KE:]P^*&=\Y6:J\A<L,Q9!>NF H3-X!6E:>3<&&4J"D/S''C<+
PG-E:+'? S4QY_?F5LB_"(V_9*8!M<#,@T2 6J5(1^B3S=8"%&Z,L#S!SP($'\6*K
PD4_WQQ&AF%GW]3G_5$@?7F;8N6/_;UER@Z94I1K%]Z$UPP *.AJW$/067(J?X?Z)
PESL= 6_U Z4;"EK /78SL,PJV^U1,[CP$WXC9&K 7$Y*U9JU27]2-E]L$?51TA)H
PA[TO]@>.;*H(K RE3FLHXF*'&CR>YN58\PK_INN)!<R A!T)3B.6FP^CCE1]O H1
P^D)R<L0B9>%)$<S>E^V[RY2V[7GSA-%6XW'<<?3\Y@9:.I.YF+0>X=<0//+$M>.2
PJ4(VPJYDSGB%3=J9=[S5>BD0^N_;!_ U_CP&:/8(IE+=6*J>/,F)%L29?^9G)#./
P<>&;0]/C,#]D,7]]KFMQ.$B;SHC_08CEOH)V9WKE-66()HA%_3)AK,XL\(!O\J"D
PJ\+BS1WX6ZUK8B>S8#=<:!/7; YJT!D>CS6,&(1QMBN/RF4 ?$ /2^%#LWFTD^[,
PF%+U14-O\-U[EI\)4*Q:"^\=HV%VH;+9'6,Z)BJ LQNBU-BJ@\72N@J:PI%00+^C
P&J@L)\SR\:\KK;A('K6]-NHD==9;OD0C;_\FI/VD%9]X%F28;!' !'K2OM#^25VK
PX_PXZ@P\3VS[-G+&E0^TYC15NSRV"2<M-'_4AYG7.LGB ES9P<GVTDA^I2RQ'21?
P]9&'89F42_G\%76S<B>H\I;L2R7;FM((*'+?GA":1(&R"#9GE!;:0A_53G! 9[;[
P]J^1,BY:H.0"^-2I'-.WQ  W)C@2OD4K J 7&*0G)@+R\^L(KVLGRWR(U?T)M_+H
PTW:W?,2L2\C/1P'S(.6&5!.91C3%[!?8>E"#=I=(C6/]ER.G6'/ZBY^*],@O8PAJ
P=,Z=XJV]<G[PN:H@.SP\>?J'3-#</MK\/ZZP'A7Q<Z\<K&R6AUVG=O"1PFV$Y1 >
PT)GV_T^8!Z))?;BG&Z_U5Y-<NKO&18T/^*:O ,?Y+58WNK6%:[V]-+M\Q\20R!-<
PQBX?+JYG;.:NI/Q>S(%#-B]6Q[TQ$,XWAC1O"JS$-L60 FARB?)H'_,1Z$DR5QVS
P[Q>A*!\:P7V=BB?B6>1T<XI LB[4OHN*;E@R-'^ N^N]14M (G+Y,-P9RW2?'.E[
P#H(;T\L]9B>&Z@72JW"?NS7V9/2$J@62P_OZ%4I@& L?@2: 1\M;!5+]5QP -"6E
P7.SMQ)3Q,;%%\QCK^RSM^;3O2^8@J2H(74<<#*:WOI*^&AD%=G6D;+ PN&=S$IB!
PD#8A8I&V:N)3R'!,Q<[H+@[YZXWH<&S@WL[>'7.I3^I19+2J"GOTU4T_3B:%D\?3
P+2>RM;BZ-:A3%U11[X3%DP"-RU4T1H_L:^PILKAXX;Z?KANMJ[+LLZO,K;JE:G-K
P9SC(3]^*/Y?W'^$JB:\XD01M!1CFZ=1I4YQ;6</MH/L'U0/1XP-:)-V5MHTAY<+@
PP2"^G9>^S"^M?U- BMP.PUSC^C</NQA4\Z_MF[%\H6R#;XQ/*+#] T1N?(B5EP>@
P*I_2VC1P'P+L7?C3"U\;L; BNMZ'CG%37/>CP;!41A!C3$JY%0]R; G["5W1S+O,
P3W><N?"+3V>YTB]>$@HOS@8FC$QF*%JD% ,UEBBN?WL/($-0MDXP+UD/Q6Z8AN+V
PT>C $@%2[=71(ETWK_:=-Z@YY18-K)=1"Z2,%ACC5_#Y7@! TMOMG\;$.?+KCKZC
P,]@.40^V^C"$C<1K[IJF4J4&<8$7^AR7D% H4Q*$ /EL&U5VG7E(OK-VJQ_@$+18
P6N.=@1_#Y2^ N=6<,TG),VIJ ?P - [;D*7U+\ /NX,5C)C?5"HPM4*4Q7+ B80@
PJ%H0V=#<4Y6_^/=9#J!U'EY'GWB#%*^M(;E>GY08%=D6:80;F"?G U_!BL::;G0?
PIZ+WXQ!NXXJL"7>PKBOT #I W^0NZUA)/%:^CO*2H]I] +N-.JS,YY8Q'=3-"/O+
P%)^<V^BX!DQL6%-4PJ!A.Q3.AI.D B9C/@6&<IW8'CM=$<0(@[&E%UI1GHS.HX>D
P%KSK_/=)'9@LGQI[9#)FL1V.G X,5B:+;-WF)HE\6+QO,4/&PTQ=2-1B=OW.A7JR
PJTSMER5"52N$.H0 Z[RRJ]EH87U,AK%U8UB..VUBB"'81X#F?7CA4XO?=]]]6;Y&
PCXEUW'<JQ+%6-B8=FR3CYI#L]:)#ED'TCDA8"'#"-8K#FE< T$_=%EH,4Z"ZZ(BV
P.(#0)M-O2@::A=6/\D9OL%&K>RZ*B%.<YZ]#O% P0.$8J/5IH0.&;BX\\5F01$P_
PLS):P6:F>%X G6O@ H37R<%M-0[UQ#],GQ61.1*'[.7SG?U""-\J>I@_!Y:7I\^<
PJ'-1IJ1#2CQ%#UM\.D</=O+0)"XZU__9!D\)0VJVJ5BY\AQ]"?+>^;LL/(Q>#^"R
P%TYSHE_K\M4?$@$F*#@P:^Z*"E3D6JB7[IYH"]W,G,O#DD R]7]RBH;V%:C&1QP+
PN@\1QL.%IK/V$TM!+(3+T).OW?\^0)\;WI@-@2I(.D26&H!S,-R8UX46DMG_=1>J
PCUNJSC$"7AOBBI_ZA_L&RBGIN*G,[2-TKL^B(IHO#/A/[#C.G,:C]\_M@&-G)LYD
P/]WGVIC8)W96\BQAO,E6PIJ]8E\GDKH1XZSE:$G3N3C:V3(IVZ/7]D464/5Z*8JB
P6Z4^2O!I(6B/6J+&?6\!KQT<+GW+%DA+EK(.0PJM+Q$V0^.6SU<4#T:)]E:,=0X8
P%<^P\<[7FG^>I/'-@(-]K(&][GT#L@3+?3L?5R:7OG3+IC1Z;:JB87PU"A?<ZGU&
P!>9K 2+OVFPZ)J:?_4YWE7(;>I 2!70#""&J8;?%>9'%[CB>%-U+NP APL[N1(+&
P^9QR?K47AB4X">2=(J0S@^W,+ AS4UX@#> 5E>Y! L(USR_=^@/+(G[;'K4FXJ3+
PXYME=)9-WCBQ%(;(+5<F$A.$MJM&?X*M"7H!#4-&E]D1< &YM7I[HQ"<:(?':2Y?
P]XB=1OC.:,"6HH?_3W=*&/LRQ+"^=]*V<K %Q=P^WI0_O]&,_T7'YZV -? WZ%^3
P1O_4Y&G]&MD(@-9?-S?@AT"38Y,)6(..O9$"2TI=JG>F53AF:QZWI(%#8H<3/HHK
P^-K]%212GJC6T3PPAM:8E=>:V8E>.*]]<APQY='R*U;J2*DENMCF;NJ$KC%::K8Y
P#+@R>5P/AN\[P^JDT2]R]X[4:^/,4__<[D)L_*G&^H9W[PG&?%\88OM[1@=\903Y
P>5?B]&E? I3]**&RV6@W-8G/<"-56F0?/7NAX Q-M=WH(=[>3<'-G3T0V/4<LFX0
P>&KYD4@#)SYKS+#6MT;P(.:A20=#4SGYIPO3AJ@P/ P,'N8XGX!26+61RK5"G[9%
PJ4LSLB$.34DYN;MI&G;+%7A:Q31YJ*,P34LZ04HJBR73=L8;%K?3& ?^%5.+PMF-
PKX+8 ?,Z?C<.]?8Z6!^TN'Q#9U*7!8W8Y.'$;"=%"S>6,K(^K/EP_;'P0_GS^F*?
P<E<XM]3@B*M%BBH6L+<]^$#L8?B4$W7UA90^2(^=!=3T?<QU1#-!_G=W,9-\''6W
P%H&=FJ'O8TT0H[B#AH=B*>3_PWH!59Q-] D&2JV9?>:Z@X.6-]_/G8V_39T$-X^4
P5=%.QD_MZ7<<YXIS-OJ%A&Q+7U_0IH+\ .HFX1.WMMNF17 *1R9ZU[5X3I)>C\NH
P37PEX RB*6F(24Y4F"FMU<"P>E#$!'J56I37E^RZWXCC:.6AU?Y2[1K:-<KI/ZQ<
P8XSE=^3[/YP_?^O:$@&]OZZZR!OX#D_G.<Y.9RVVO#K(4@9I8YY".9_/6)>^X+R7
P,&W,\:FK9I8!&8J+8??[-7R:PT<MW8)WCY 997B*RK1OU=@:9%?<%ZXS.@ A'\#^
P(+<L.YZ,A^0%+I60X:LOI3\M4<8.5[4F*F#QWB[*N4CJ0*=%Y!#P]UO1;YRE#?)C
PBJ<]BA!".][Q-HHMQBVX[<J/$4*\$=[$M7@8*T$S2(IMG==U:I3Q^8]J !(W30NJ
P5L^ID#KWNR'3+R)0R(M'&4(H\N+SV<<\FYET>+Z@7CRO]%A]ED;BT1M EQW72'D!
P;E5OT]%SE=I+OSFZ\^S<]>,X:OF/1P4QAZ@^*^?FT#D)N!=00CRRJJ],S79V-73-
P>3W@!J[3MA7 RX^0D:HJM%P_0!"X/7&B@U6J&^7=DTOK+WC /2!GO,BC0ZUMK&WC
P?0O^I3Z76D]=D)N*SHH(*&:LH$6"71C=FKHEET,4E[D-FQ^Y^_+#, Z8.PPEW:BL
PQ2:J9MQ(R(#7&\Q@G:9.W3EJ2+4[, < PP^6"N^9:1$6/1V(L;TN0PC$$<M91+Y9
P*.!$BGALW#.[= =0=)%#"1L/F&*JS^U ;6Z!):3O,J#LJ]+[?+W&[T!:TC\E:., 
PI#,8AH: S3]V%JX@G$_<!1D_\HMA,_]?"*27\7XH^_:H"R3YB%N(9M4V4*EGPJ.!
PG&= 2*>3K^!NE+(PW;@G!?I3_6J:\3>0%'H_%\'< $\58QKL;WI6%YSHL_9,S-RK
PT]'NNIAVLS$%L=<X_T"!.3U/P*GGV(_LNC"GQ+;%2&79JDYA9&,)LH?.=3]/XE 7
P);#2 @]2'U#*R3VT-@%E]YAG]A=ONON(U<%,_3.6NE59Z<?LG>O9[?Q*!7,Q;D>)
P!8MRD:?FV.M5],A9@Z9Z CK*072:RH1FF)ETQ:$LD"?6!2Y:S5JU'0D(^K,RSE?!
P=DX=[==,9:-% #9<_^A6[;?;?%8&58TM]3KM$?"GX!-WML3E5 J8$7W[J5*D\[V 
P!I87/18BB^P(-#[?2^:WD6-QTB\0Z[1W;\((1C3>_:%/ ^!TD4P5AVK!6$#%?"M"
P'4\'&TJXB2=>*"+TVRP?LKUJ56AP#KK6%(GZJI@:K/OOH%JO *ZR$K,OCB,RT4N?
P_X^(AX9(BCA1*O_!%._1'?*HO#FI*X/SQ&-9<1YU4@:Q:DL50P@T-SJ4Q [IEK3-
P9S#>5OC]P7Z_UOUI58'+GV32O?9_^KE!XN4R4J)IUKU]$D[BCG'O@F96)L5<:!&%
PX6YJIJ-</MBR\PKVEUZ^U4P&V0U.K=5IL+D1DJH95LBS?%D9FI12-?R\:1PR_,;#
PI_^9@II\9)<#.E# O6^W\;5J/+N&E*<QY_!1$+)G*0 &6C@*\0@DWF&CZ+5+ Z$V
P3##@]4^2V5D" OB1=N_V2:U.J[I]5C^UJE5?;UE%L(<!WLQJVS^"$%=U[F]NNZ: 
PKE/LP[_JF SJV@L)?SP;$$&$H_4"&Q4&9U'B>K\;T_VHU,?8VHV1C6PP00._Y/?K
P.IG5R_<1YLIXYS:[MAL)WY< C=$#MVKOG'%Y! 3'%AQ%2?)%!O3=70]]E5"4L"W%
P.R.LS #H_M88MF.+N2Z-O/K=-)5_#\432EN\//NP+&+AVU2F[>\H3M$F3K:(V)/@
P_]I@K+'K<UQ/%$JPY1:\H/9L5&V@4@XL$0XH%:0@2@3B%S5_LBPI<6E&+0F6'K=+
P7L!.\K"/0H 7O'?? 5XHHB=O;YWGZ@ 8)4F3X=?(2-+Z#:1?+V&.4:GB] _1+8<1
PGREN21'[J",YL(WDBS*^084UT8=)A<I#^-=>;BS:%2X=-O5"F3(!U]X\]Q+$<J$B
PG>[7;#10?"LZ9H*L/2-$H!>Q>^X4E+5 //8T!9@RL.I VKIM*<OP0L[$U*.A'XVV
PRX*M$@8K$N ='JTY<3"D"85F,X,X%">!G?.$G)J'UPK M:2DK4S 2U*BXI<K6Z4[
PQ43KY-ROWY20F'IGA@6PAG WX@5T:\;JH[H'K,'$)'&LW-!"1X^) [*%L#"/?XJF
P$I\-^]9-S<FW9U7\&C:]6NC/44VLVH0*!R:ON[2S)KFL^7?M7+@PJ/G/S68]>M4&
PP3GSTS'@//X@I6V9BVMRT%*.=";HEUKPPC6TS5I5S!O@8;"1TM/N*RTL7J63'J6U
P\R&-%HSB&=#X;#V1>6WT5%"U[U, V53W_L]VRYX^I$%&')CX-3#) ;;@%T7F\'(;
PXVXN"S3\6.B@Z]/' _%Z>NY=:*GZLM<6=9XQR4<UF$WG4'I)$;[!2>0W6"8\&9:7
P2G*3"QC0U-I2]GNC"L'XF</63L8"DK$."V#@B$AG)-"*OD5$4A6,W+G_T\CY_SYN
P,U38J(SR8^&>-XXTQBIM*MNC+I9&4<9:00Y5C+[!\#P$U^NSM\K(1T,>J1;XM?Q"
PZ(':UQ@4A $]63$I\3R6O=Q:S_H\7;#3&#\S0:(!*!*B(FUJ-YV3S\OAZZ,J4%>O
P3)\&J,R><J;.\T8:8^ <TW/Q%!LJ=762*HV'R370[%ACXE%_3>-(V.LK[:51TZ^C
P<[AJ/SHOT,8R7\J?/H[,P_7Y"IYXO)]'N.KDJ_\U!#CHVA(\6-Z)X!.@E6&3,G'@
P>;^_/VR.ZRN#^[PA[_ZG#B RD@7BDZ#*+AQ"%U=E&4H5@<J.>:#ITFX_HVH7EDI$
PM@?^#JI_-FK)<8R>>.\*G3)6[F\R@=YGXWQL7RJ*9[&,95\ZT<.M62A+W =(Y,2>
P(==YNQEGM?2!V\;;%>(9P/[(J>EB$:=6_&NUB]68[(D[=K^V%3ZYO:=RA:CGJ3\9
PE'FB^#21G*9ACQU_$#D!+G/HTC8RDGL9'NF$Z7II^DW.'_L58S/BZ1-?"WID8/]D
PN-FTD6:)L'5 -:%'33F^7;G'_H.E1B;)&; H8=S'?ZZ7\5MXE;['6&IR'W6-%M/0
PHUK+;TJTTE#R&A^,3"IL\#2\RQC(='R47];&19:^6?8!PL*;39G;++S+J&#CT#Z6
P6R*&)L^6M44WWU[C[T1J?4W6#6B66G 1":P(>#4='_GP[>V [0W>67F6MVO;"\@N
P@-J(W0&;637AU1E-<B@X,QX/Q-F*]1ZC@-V1U  ,HVYZ#6QV=:]OTUT%I-$KHXPR
PL"H M,SGU %C),QKS([,"5]H#W2IXV2=JN 0$5SO$9Q[#\:N\/?9[C+S,GZ@TS.T
P"NG7SK0<;S!)O2_RI'FV@JGO+Q(3-U+VLS:@6DU"_U=^J71#,IF[D'[-$?J23L6)
P-03BA@"@!0]L@[=T^[><5SQ=Y><X=2M O-E(F/0-4Z<ZZ%(!),E/39 F>=F3DFV_
PK3%$:DD ,U%X](JJIXB7M^-$8?_?\/Y"G?^USHM[Z!XQTP]>4J>)USF3%PRQKFU7
P'!SJ7(,:J["<"SW3'*\II/FRI$WU"YBJ! 7,]I"SBM?S)V("!U5^>-U$<:?F,XHX
PD;H6.Q Q?R%A/9FK=$Z-*5B'Q^2'RA<9&VB*55W!GMPS:S\VS&U8<S"5PPO$,?BT
P99:TCM0-@QN#FX+GH^I*$Y4J]:&I4.UR8Q"_#UE@JC-IH/(;<VOWIRW9#;,W,"SA
P+K';/4)UKF.7DP#IU_ 3S.D[)L<_7B4FCP-;X(]7&HU0=(+CJB-Z:,X=66"RD?D9
P0C!0X.0O;EYEFW##KC#OE$)@?NS>;21"CQ[X5S@#"3E+2[S'B$D/&]&5A\81Q[KQ
PG0%#A4TT.R391J[JQ9PG%:CZCH.,PYEL7>//&RY9*3HI<DW\4HO&;N1&W6JLQ+"A
P.5> =IT<G1T,K@,&UQ)LUK=6,25YPZUH3& XW]WFC95R"3=@#RBI-?KSM0V3_>)A
P8X'H.R&#E,#P+O.$$#KGZ[@C0&=;L@A#[B2\^"G@ 3:L(9>>*M-WMMX![JY;.FE#
PJGE(W\CSJ$!'$IS#BS&KDY\*24&8I.Y8DV__-U.2@2KK2:\'DE),-5[I;"?@E[3'
P:3L=I]!_+RB&C50YJ3<]T?6I*Y 2[_RCCY!4!S5495#^P(#YDN9Y&@I[:8@EJ2ZD
P5@5#FU+.8V)^\!U1.LFV33QW1/#5L/C,)P\5GU,G4B_9]L"C15?:OS%[H=-1G"?&
P%>3<37HUS5 7=8SN6Z)%YFN(AY#=2DF#7;(X9J].3N^\4#]+?L%\P+2ZS7YCI1P=
P@ST!NI9.,)!:V,?JB5E<6U*=J\BY9\V9'0/54EJ.?/.\=1-_I?AQTS#FIE&_)2C]
PMG7.468GHHEN]+_Z'A07^7^'2F@D]$=<.,9V'R*RSL@N$]"4 <*9V@I [J\382!6
PZ;G H_E"7KF)YC==&7K AB".-U$+N:.;\A%IW3!$ROV@63N15'KQ!&;^ S1N]"8I
P!EF>'59TI4PQ/^M>&\GTD-I=YQD??;(8](\==QR@(#Z1]!TBX?$*]LIQN!:]_(7I
P4A!*;@*MGP:!["OI&9;U#&F=;&?:6SE'(46 JV\I/$.J?4=KES121*)%\-.G<USB
P[<3)97CF4Y.YS5;EF63]UY1C'[9/-W50)V<M^@S2EY&;%FG0ARA7.:E"YPM?VGF_
P]6)XV225*%]6/P_]WRV__F"0(Y-*#O#IQ$?_&U]G+123R3->?#1[I:2@[(X/I7(3
PDHO8[-AZ,/H1XAU,(2L.1"@D;W1\WZ<)ZE'W.];(<]AW(+LH)*[VB5DVX^NN/0NP
P\R<'Y8:(?_ZO "+D@RR ,!!>':?>X3J+>U[B'G%5B'I3#/L:N^FBE)N55)4U7"@E
PN'8,MG^B+Y>]MDJT#[?;!S-2]!9V=*6'$G%8;BO/-5\N&^\44#![5MX9\V!$ZXJH
P?(R"P$8'$^ROY]9,^+Z"4W/OYHHWH%#[X2)HMF!H_L@R=:[E8QB?7IK)YYG\"/6=
PD?S\1/HZV[OC.I,5D\5%*A5#$7]@!DXR[;,9\A<R:(Q=4"R!K7CU&FB0!FL)P>N[
P6X4N\R=2JA4B!EJ8(3"]%[K[=%QZM:$N%EZU+W[!MG9* XR[NV=C.O_;^ZCC_.:6
P*N] NM_IZ5CVS^&A\AJW--PTW'QZJZYP*XM*>M6"17M$,_YC;%%<0F37)9O_AR,0
PHOC5OJLV4N@?[IKUO>= ! 3BX--7,&/#MA9$4">9[(B=Y_)PBYK;GLW."U:DV=?G
P75I#KB&&WV'L^TY$8% H5,2_Z4>6LL@J/)^V.'P<P$RY14( -7,X,=X<WD1#NR,B
P;TB+$'VX1$UVU_C]B;NC ,:J&:PY870Q16GP*(7-HO/#E1(-Y(36170PTE&=53MB
P=$B*U39G34P"Z!8*+8@SG4\>GGSVR&F1(5\*TP_R"C;  S_/EM@JM]WT[[8G2=U(
P$?!9R<H@$+9Z-J@(J%7H9NK;C]%?.0 /VMCIM85\T5MG8)A\1OXO =%K7T)&T&F+
P;JQF0O;O5>%B0U>W@U8F&Q)>/2&[GK=]FKZ?0[0'!KRN-X.PO49[\T1'!,38"21#
P@Y#ZL[T2P1C%>7US?)\]EC14RP;R+JH18M ,=,+%=5T[MU34&@#\GS4JLSU R@IB
PUR^NL1ZL(0-)<TU:<J/E5Y*.#L<<?7Z0KMG#Y;7T5UOKK6Z:QT#:YN+OC[H'8XI0
P?%_O9=&G7.C:";2#'*5F"GYUYPL]V56=G9#;<>HC:[/R;R:WF+6U^4*IJZ/T(R8)
P!7[+AF^W@OI@/ ^9Q44H0L42AC.IK[AEL\!LH@U0L,@VAT3B$CISJB,JX&I%!!$Q
PWT/]MV)Q9$[5F_DM%+W[\$UI!80'[>[D@I2F%?"%1H";7BL7&%$D#>F.0\JN;'LA
P"A=@4&[C%5HS_OL+54^0-?BU6+=W#JK91>;#$AQ*0/@CCU<N;G0)'Q^W\>S5;@J[
P@A6Q^@RO )P@DD-];3VW1S_29@I89-70[<YD#L#8HW]ZWI[:KCAIN14I;;X&SK01
PI#EL@?(K9'L-.JT,D)A.6H3'W$D!J?$#P$[(?H8G#N0#3SDAI@D<$;)"27!#GTJ-
P*%J,X6&1[QC\G7WNMGCD;A<CSK6,T]XTPN>WF]2B_H'I ;5IP"WK/<LN2\R2A=!:
P'=\*^54_'[#4(,P!&BH\>W UMESYI?_#9##AH!#<*10!A0Z!=TBQG?AVBL2VK_>R
PF#8<3(2SE)?P##S,7Q7L]85BU98WN<&5,^1M(,>WX"#)D?LP8BZ0>.//^.LR*YJ4
PGVY#O3D7-J<"=_T[;9@SF9_^8\H1*ZYVMCZQL8PN[,LZ@YDUH\(7.D7:94ZCX75-
PIUAA#(PLLE\<)VWNP"GL%PX"R)$!0HP7.A:ZRT"CIFNPK;#[*]'/!"]]3I\@4<$)
P9KKQ*8H"4._1J_@0A=M$N4PF0;ZA6D!)D*&O%AR%@'DM1;\(/MA'XP-XFE=53_;]
P1Z2Q,)MW!FEJ5CE/DL0*1+0"R93(H%GMF>(:]TU0;[UI-E 7IE<, <6U16=W&X74
PQ38O9=]#(3@2)6D8/<BU)^'EI]3F]XWN/Z:!,A'T\-X.DK'RF=(_*+)7D!/$7X]3
PW"=\J2V^V(0Y&=Q])%C70K![DTW7C,"2O 0.2@SY=Y(]L*A-$'U:Q'D0U3O0PD.L
PPG6GM0;KL6V3"S6GD@V6OCJB3\W^,7);]->5>H7BC)NJY?.B"B-*4 BE/[\@E<]E
PT]1>.2W5H? 0W0J6TVT;A-A"KR2P6?J\_=9E>-H8=412(-<L^;HXH E.?(Q@10-V
P%['DPK8=QW1)H?LI4_!%:19UZ=(KU=X@^N1Z_G5.**)QMDG)Q3]M7,O0+[A_90E-
POR5F @H^<O6QU>'NOV*:.]E_4E1A>?#31TIP7QP*8"!&1Y7;?.Z1;#SG.VF\S[DD
PYEF<29N_D08V2U%T(;"@#:Q)*Y )RM=SKZI<--G[I[25X74+ITB6(HBYHI+%9:.F
PJ,P7JEX+<(H,7"I,;C:JKQ"%-\X5\[#'$))U4:+UN:RD7DH+K4$]W07(/C'*1^2J
P#,M]&N[BHA$\X[N64W[\@H%,%;J(4J!=KRGP7.0@126"Y;]L$FEC_]K.H-2)+PM(
P+=+Y_7N&U]]*W\9J636:&1N"L)+V&QK*A3Z4W]-ZO?^]A<;AL:I$%FE4C>#RG^I%
P:42$^DHM8Q]F/*MZ*+0\B\,?'PCPET6&19J4Q#QL^W"O\1N#['>EI9Y+'"[>2(R,
PYG.O(E<-A[I9T>KPEJV[P4= VLV)<2B=BG.^-GBK:!)R;:H9DM)G\&-PLRO."@KJ
PB"V4\/Z+B&>04LH!""NYE.O<?JZ;\>=_N8ZB:,\&N,F<DHC%/'#761KW&WHR^783
P98Y&J(XC8\*4E0P]L["3(F[:Y#YH,4F6K3I8R10:.?!8.@REXV:<E^_RH.%,$-Y*
P5+I9LNRWP_J;7E37ZZDC?OB9>BG0QP,D1;2X'&OUZB 1*&M+4G.L)B]/-OTO3T(]
P540C' L@GALX+W0$ TGZBYTO $=DV%GZ);$LW^$KCNV61:GF#D)%IDTGM/I//S9%
P!*\4,",3>Q[9KG0?X=<@-%&BN\>T]#TVV%I % D1BKS&=./-$41.3)BG7C.4:D(B
P6J ;J#FZ=M;K724-N^N! 7B<(QRPR-/AABT+,74"+O,_G!R?]NTD=,8L2IB;&DW"
PVIQ@"V!>( W8]"':W *"*/7F6^I+$SB@'\= Q7P;H8+U$S(2GL!D],9$[:DWS5-G
PMELGZ:%Z*QYO+21Y@R=^FE*/5)!?6YG.)-APRW*C#)/O.T3%62JBVFR0XZX:;HHR
P63V<HPRH+A,7D];-1YK25!,D<V^!Z@K#-14SG= )T8F/DD%_Y$/:FLV=[QZ"I_(N
P?+F0HLJ#F=W66X;I,,17=#YLD;EM@J\).$Z856X) 7BKH % RAE_3)UM&['OA=PR
P@%&G35VLC.>IL@&I$"8'H" '=%>L@=9)=,4@P_R\(OL1[AT/F4G][$O*GS 3@/#6
P*M$KA<^-\9*AQ[7XV[MC-^O-+N_.A!S:GMPVC]E&<^L^*1'OFBM\2!.UYWN-OXG\
P2"] 1T[BEY1YT5],3ELV>EXBY]J+WSK/*R_VF:@_9EA&>KH1H9V)NU>@Z\BKMSGR
PLEB&4]+]V[N%6H+L[,K@>H*D?D;)RR!+_!,[@P(/%8:;2!J:U&+X&%(BV'Q_"%+/
P5M' XP%(BCU18QSC9ZA/K$D]1-T#7!-_O8+F&CAKVF?C.<V2ZTI'%/O7'+Z\>)M]
PL3XMD3^-1>P^/E/#3R(S!'F2R3)<-^/E>+JIY^X7WM7TUF^$?VGS26&3MQP/R.I.
P9V\24F4F47E8&H GUTF*8CNVZ&UQCA:>Q+6=@EVF*</%406,B],%>2 ?0_6,%$6+
PJ/]@<]K5:>: 725NCBMVDAHXV);?W#FX&+?ZY+9C9_Z6+U^>K+G,(3JO6EY(>RV[
PF)3IO#_<^;YLF%T >]L5DIE(-HHCC,LAOCDG4U2\D&VS;CRD;!LMA%8N@@=L4=]V
PYCJRRQ7A;_\R?*L<S&LYUY@H*+:"VCO\)Z(74\?=^Z(_5:IE5"\;DN5*T2P$W-LH
PWOSQZ\L.HZYN^[17_.1)F4X1R!)B'5'ZR[NEWSD+1XAB'\"P8ZCB-XDJ7I4_=7CU
PEE [6,UF8S9,9;#VN[+UW:%?[TE5XU9A_QN7'.MG;__,G0FK74=P[U2"%S"-A) )
PI4SBWC"<-%,> JYX+D.D&7 _<4K&8/GN'TFZ9#L TQ6"2^(E^'GC @L&CY8R*U2:
PFLW6J-[?YQF!OL3@L&>&3F!R<S]OT;H 'O?FFO,!_^N/4[A3#0Q[>)E5@^B!,1&F
PJ]Q+YR?^F]M"KX%1!,;_3L(OS?V$B;MWL75,,Y-?Y*L>@QXCEZP8#PF3CY0P!^,R
P@:T',31JW?9 $ W!_CD =Q3RJDZ?; _?? +L2(1E:)_B_TMY8X?<63HC78^!O;*6
PK(Y%1X!1TJ.2-"T)8=^<^0 B<[9"A_OC!)XOI_-6JY=HZM KAWHZJ/HA>)_WBE=7
P]O6;IQHT[._?M@&N^S;@K=)>,!_[@:%Z 5RE(3<.#5B/*V<\[O?'+PO@4_W>\M=6
P[?&JH'P(%5Y:-P.@9]Y0<1B)R-1!<V NZ/L@BS#,.-=U86+L]A4'SV"BR0.[CYX'
P)J!)(MEL0@CZ.2U^AIF4T8@BA\*/>;-/=T*Z"AMZT1L]#A)HZ3];I:WOPCUFOTW&
P"D'%(<F&876;'MGMV6:<SQ@:O>8L(F+.S-_*A.J ,>F<R<7(S;VPU<@K^3GCC*<H
PF=3HU\;_S2G22TV$IP",B=G9)H@/UG9!PC>\"/^LMG\=NA6R7Y].\?WAM5PX&K'Q
POV[,?53@[D'!?5C*>CW[*7I,--1_GRYG&-[?O9 ZXC[5TAR]964KN?+AH29/E%3N
P_CZF ?+4,\"I&.?C#)ML^K%$>JV^_+T>\YLB:2$_A:K@4?KX;.70L+T9M/MFH/Z8
P<OJ%($$)>)?B@P*IT82A/=5,"NMR>I].+:.JZCN%._.3=8!#OX5$<E#$P[M41]DV
P7413VXF6G@T,=NW[-3$\%4@BJE$'\)<9+H2[=.AKE/I_)TMIB6LN#=VDL@I" CYW
P_F_ Z3KL?"DGLE7(A8J7<<VKIP,"T6=[B_+%9+,,,R9WV ; 11(J8Z"I=/$!)#4Y
PC<&91N.PACU)-7X<\_.D?)O1VRV0*B8%==48C:09"W%PG=V1,*L71Z!!R0. EHNZ
P5YQ._O(>SS:,O1ZCX60]EA3"FKGB?/(2W8 /Z,&]Y55TY%/#RYEQ-XZXF.,R,D,%
P/T?HZY(K_>I1?(*=JNV/ OPC3DJ3.;U2U^2%NJMA+V1_>-7@!9:GKA8@7Z0?@*C!
P1V&>V:0I:,'AQ-ZF__@LW#O!W>YQC_QF!?G! /93"7$A"AX2QJ66YNH"=#\,"VR"
P<))Y-JQ4% K5XM)2DH3A.A$OT*V%_S!.9MG[9ZI@*HO%47@.[!E# L(>)/!M!,24
P?]#T*GY$A_F)"(;:S7)J+DX=&G>N-S=:T"*RO^>45@!_PT__CZ+K&ETPSGH$_85D
PLT3K55&PJ,44FM/7C[DCB\&G#R5-&O7XA-$+ICJ-N.$4J(2T'.DD51THX8C%@3.M
P+AJU0?F'&VB'I'&\.'*T>X:79C-;B$:R5; (5$D6%\:$7X_KQK3-ICXQ(2;DP( E
P,!,%UO;[O/V 1I%W':YUL)UM:02UO+;V/_,IT313HS.PU'KG&26=D^MZO45B0LN6
P#?+4$UG"P$K C?F'A:7LG_[_@/.41ZY4DPE]T0Y"0H<#HL.*2D NF;\YYV,:J#_\
P8A*2,<WS\JY*F<J#!KF%>[QJH>>02X[3F<OZ :$"![9Y<8;/HI(F&78>+-W >B3D
P61YV*5;)V;B2QK7FH@_4$*Y^IG=?W'SI\=3E8,2D]?(-A5:TFX6?GK]?8GYZ\\=U
P4ZFT:.$4>V2)U((XS[1[1@R("':@!MR/5- ) 4!F>13U29-B*<HWP8L,T$3!5015
PE/E*5PG4!F_X55/DE@CZCXY"<DX-VIY$3Y8&+A<^]-_MA6A$:C\S/&SCA$\-%#L+
P>1O&Z+O\X<3:M.D!VM@G:S=D<<?M5$D8KH$()5 LW?H*/>*5ZL8=L%6KX9V-PH/4
P4RLH\^QEC#G3[4O>M/!WYB8'%;ZD'^Y[IN<443"5S7K#:\&0X6B"HA(R(%C?0FF]
PT6RJ=N*VN21D#OE)J\6+ARW$ESN+X _R_?.U00 (RIG423MT^;0FPWN$00"G:YU<
P6_:55>U>%2)8,FLY>_*8[S>C"S<^@9:X*ATGV+=N#S!_MSI@TQD%/&MJGZ["\ZD]
PIW^\S3A.7PM8&9@/4>_^K7L$_]RJ=2N@;(!W&T:#NV[=6;YC4)M%6 *]S>.-ZAA\
PYEE)$...&JOI69U@>XJ?1=PO7!JK,S[=(08,'U9_V;\S33$N-VDZ:7GRB(6%F5(A
P4VVV9*'K*XJM5*O9R>31S5<9&F+^,WHTR/0\$+_P#S0I^7;]C0#'_)'.3*@5@R'6
PN6Y%_D@>%/P%DL[S.0>@C"KIZI8RP#BD.8#9@3//*^6#Q0QV0$M>M3_R"1B<C:'8
P>F;C+41.)Y(>VW0C VT(3)XVK]<4N8C=\RK;!.$9,]W]NUZUP?3P\-+.&/9)IT2+
P#QH!RUC"@"A)6E/;XQ,7L&54\_X.5-WL39^G\]0@@(47,K]Q0X[]*D(Y.O.69F<)
P S_X:&&R^\AVZI3+#2E3X0P,ZX9O%7)ZG.;!8=^C]69$"<^%W;G/LE5CD2@HX&GZ
P/L+B9W*S<]^[=OP=EMB0< LW\4<?]V;G+FP-X(JG ^$XVFK#$*N 3((*I5)EO155
P9Q39MV,SU!]?WPB4')<:.S* /!BZSQ,^@4' \/J01M">9I9<BL#D;2&DIQ)JP"HX
P#0NT'#3.R#H_-"<?/[;!)CY#V-(GPR_ZK<GK35AI4 CN%,EVI_8)EH4/R#EM94GF
PK-A ]?#5@*W[5,4TDO9U@2/FG!;VM19LTR[JNVF!]!W,W/JZF:Z.X)#6W,KI$^1 
P%$8?24J/?ENB5'T9=*O3O?HHURH0X_[E#_E3HW^8GO5?PHCM7JV.EUZ&.\ZTZ3B^
P=I0N!\K])MVA";4<<'W"3I"JO/')/P0QA>(5!H/+&!C/AXDNYBV:0/XD\K_JJQ;T
PVRE 0"Z/]94O?+XF(EI8WBK*M,S&92?P=O;5DV%>8PD1R86P;VX9@^_(?W6W</^7
PWCJG=_GB4/T?J,7G"1M[_1>-WHNRG+'?4G2IA-C-Z>8.K-.[=(/-W*H(>&?RAC5N
P$=*B(]HY)/(M'\F7GEOPVNNTU\GH>HR[T9+@HK$VU#<&L3, +-)6T\F]>N.LS0CO
PX)[Y?AS!Z@@CYQA-\R9@!37<Z@?[0QQ4TPW'[_B[OCS?-[U-P1"<8&$/OT4DYQJ%
P3LKA49@/B6>,;-O"_&I=%$Q<)<WTR<V$I'A&%Q.W%\*#O>C&FLEM(:7=-7Y5OA92
PX36F-$6+9@9"'5&(& ON((!2<XWH54^&(V8$=F4;QBR]7[RP)5/EKY6@Q!,A5#H^
PA9_EL[Z9#?<A+''MR!BV$$8QK>(-+OA3O9__0>>Q+O?LR<3E/4JW&.7>L5/>F^ZX
PX.M%<G,@IO@P&YU5=AV?Y^A@F5Q4G!.]JB2T,-2?>*;[?DV8K2/G,@ZLO;EQ4R95
PY71O-K12V/.)/Z[*L7]XQ3^SG5)%02[MCRDY6Q0?:@/O2V[-.UU(9V;SM!0<?Y?K
P?F8D?>"XGQIDHB!8XRN_\TE67)!]!37/4:HR>?:<[,V^U)PY-4]8MG! ($XR'R&=
P&DG\,Y^ "C3M#X/\U(^R5RG,/]Y(1A_#IRKBAWX3J2PDX,X/6LKL3&^P<*YIYO@J
PXOZ^.[F'N2]-?+IMT79SJT[W_RJIGUU"Y%U:8UV27(:%N:?PL"J=0I?. F?*>9O]
PT27+NTHEI6Y@<=$.E0]W1AZPA#<<72L 2%-\WNX!D/85?DMG#/?X4$]<OZFRZ/Q[
P4=2@K 42OS3N'XWA)"]50 ]N6[,..7+(K: [B-1,IZ]FT:N,%%J:=9 $8K8SV,2 
P G\+]GWZG%\2L9.]B$H:YTK,VMAUY\X.Z25_*K%#_&+.Q%^/N-AB.T C556#12KH
P^=_H*YW[]#9&'885N-P($P]L7 K1._E6UZR\2Q0*/E"XR(4P&7M)-'4$[&#IIJXU
P*P<\*<(4(O,+&*VWY"@[O"0D"EUK#12%H62;!7_/;0_ZK,-"*#FQ>V>RS9;(0=HL
PK=?(,QQJ/2!$7P\C1GU@L$FM;@I1Y#\(&KXSN/-98#>5KJ73=:60T/T%NQF;LNNK
PE<]!&IO6C*IZS_XE9TI7FRE@OX/=)R*'>)J0)S5/F G>] NX,*P:A,.":$TM(^V"
P/C,IL54)SD'U'_M@X6[$[4BFVR!(J%V*3W$\Q;W+Z:*LAH_56\=F!D^3X^'JN)C.
P">H25>) .J308+N3^G2D'L7J3: ^JY\^Z$;A-FZRG8X<L"1==U#>Z#)]VB/C.WN9
PNX16(XV(WO#0F373I':+(2'EHS\JL:=N+[YR7*W*/NB_,*@2EA3<7@:X+?);V0S 
PT+=JY@,^DZ:9>)%(,"'N'U=3%TH8SV*WA*Y81 Y?3BH]UCV]*#"40I@RH$$=,*&=
PO>5^*AX6#;2UTC3!TKO&>^+")#&?.-G&%T&G:TO!W%DLW)3<3L(YB+;;WH<C08D]
P21#B0: Y@ PI1@7/VQ9U:N^H=-[N86#T[YPC#D@E[<6R+!O7SE4 9_K,:3NU L1J
PR;)9;;0V=N5'TY-'@7'5#7,\MC;+O=@]"]H:<X YM((=>\^P*'>K&M6)[Z_F]/-7
P*E7_I4CU<2'[R,P$%E7 I\;=6Y2YBB'(YD&2"U3H9_U0"@KC'B_ FT+[SMC!B2N4
PIO54+%3DO^P8;\7-Q[\'Q6\DE8M4I#2)V>>V*;FM>!?Y_EH@#^;>;X3=USJWV<)L
P=.G6G-A.03=QHY$5B=;!!LR-2M30$C!I86;+TH8)$L3PW#&1"<V\5HL1T=P4+66W
P]"_Y&ONB=4^6!LO<C?7]&K]\8TG!R9 !/FU:LD(6_,7MHQS<J0(MF-9KG"F#>RWC
P#LD\E%X18F_0KO&PG>D+F'*;H$Q!-1A$GRH4._7#M*#CM'5W,[9R<WRO&2DFOF(<
P[=]IP>0U')]:NE6$$R:OJ$N33_'*J+MWS5NM!YA4&!6?CHVF-*;<".28:D@J8I% 
P4 [[HQD%R"==4)).Y_Y"T>"784P8 V5.64A.F/YX/'@ (X<<O/[(P[=@JB^>^*UE
P]5)8"DT">O^RYTXU10'GW-T:UQ6V7>D;+MDU#C254#>F\P2%V&JQL5L9[WPX04%6
PFLE4(V35O03+)(_F-U6:N& >XB\"W_O/W):?_B8Y +TA:\.4)\%S>Z8$;7X0_">N
PYX^6@JNU\1-?8P38E4<B&A!)COYP?W0SVH],-D2$/!#3HTRE;XUJ0:_)_G&>HZ0B
PH<_'1'!0WKJ%-WQR;HBUA1=>\=#SCDJ\*8N30(R,E:](E@\2F]X.,9TWSB'<XG#G
P9P]]0XA:!.,!0$)/O=,Q!5P0(60C-6>$;3L]C21,7B#I#DV'F#LE52KV;STN8U6P
P/,^R\'I836H8_V&0E9 \Y?^Z079JC)F&<@/6J1RN'3;EB"(*C/CKPH__K UQVDG#
PT_\O1YP#MANM,IV9>DI(!E[AR=$A;;.TCW;WR;'_S064TG0.]I5/YVH?)M33:W^8
P%!1H_3T=JA,@N-1*6U$D)K%QIGS>B1546*QIK27SEBN-+1*1^E18*]$7>>0%&#J6
P=.7,>\:K&I"/)EZS24PF3O<FWT'(^NNO<VGR31[?HY*D/+'MCE-KU-N^#?00*%*E
P2X*6@PXY08)6T.:7DD?,ML]"PW0#Q%[:' (':H8-(C0]\[N*91?)O;"_?.Q@'VEZ
PSB"&"-Q/1_<(4ZQV%P'/68#2/0 V_PX_6>1K,X?#LRZ-]B.I)T81?MK X!B(/D7_
P# 'UK[2?E&$<V/5O6"^!G3H]$XTI$YUH0-+VNOL"<0@CH5X1@)&MZQ,VE$0UR[+_
P)\B/V+\KLK@0B6?B@75- 5RZTU('D8(V.8I\&&1?8F\1DQ-;ILP@BD_-,. L2JCX
PW5SZ8L^.0R%G!(%B2"=J^F?0F*6SS!&WW9AS/7QBOHN6=1C0(WUQ\4G7=SLP9ZF\
PL,J(Q-U$@U*]O4$2:](MF%Y U&\%AIK;D_%LH?#MCS95%VFS=!YI9]RV$>7U ],_
PC>Y81A/<9S4DWW+^2Q$13YC4.D*<3-=SK[2ZD\Q,GT[)I7DD+RT%N($Z$(G)=8T"
PQ^M2J3-,Z/QC@YJJH=IU>\G+R<^!K5B4K")CF^^&-(A?US$W.5@1,53=8PJ,[*S 
P6Q/?#3K>/$JM_]W+Q;>AGI_;1/&_*<?4,.2::@>>RQKFD-$1D2!46YL GE %_H.A
P#@HB4=B.%" 6E^_797LW4^]"XC8]TGA7+5TU/V7E!/I63]DJ86#"M@?L)PS" %Q2
PY^@U%55')06$?)J9/W(,'%ES!72H\*N6S3M"@(-.Y\3.[-G-Y9KW-YK/^YK/XZDR
P:NMYR4 /]!F5NC5QM6ONJ0Y J\LM)3[W/'UA\=1$:B(L4&$1Z4MC0,<:JY^4CHOS
P9%/M$K4N2/L#F_;N\T2)P3$!WV4:SW+IN?4?']%=\'3G+5:?]X+B+H))U_?BMBK?
P<RS:8 @6+''VD.9K.;--D30KZ\W!M'V#&#F?-*P<V\6#-S55^0K#7"(?-;7!A0,(
PM?U@J!Q/-[.'X$S!^,H*NPD-3%Q?$H4_N="VMVC2U653F1+H:O43H[$_TT36J"YT
P^NR%0E=('1-#[V0&K&P!D)J3BAE\#H_PL;HM)(YRZ$3KR>0;]  >),_P2'C<8/C,
P[4D/4X?5UVA2XMQ$(!?I3RU"V]U8717 <F_ IO)I9!VEY/%$Y= SJBPO'5H9YM;3
PV#HKX"UY>5T42S6[R54/_G0!V?/T.00DO3'E8B05T!WR,2;!<H1RZ0DD'V.J9HW^
P59G<6O(_#CN%CZ [J9&ZMSB/\8$UB7J(@NT1#L?ED8?_NF-P-;7O>UKF=--9; \C
P@?UEQV(TN#B^#L\30,_XX2M,$1]D&%TK9P*I>*K,XL5 9%PB(9 ZJ$/8+&/_1;_8
PF?G+$%<I3:?4&TY\XSIH+'N#<!NC*2"I!PWW%[:0[0RZ3XN=.-.$Z]45UE4?IB'S
P^1ZE]-U@#$.3E-:7J.BLX5U%04=\&[YGAC]A+O\"\0B^, ._"'S["8]39, E%8] 
PEKFT?C;DT])"G[PB/(7CFVS5A0G=7V)!D'.G45J/+5N"]=W0Y1-K3<<H=0QO:$R5
PB?<BDPE;EF-R2P$(< ^L E]]FB#WDD 1 ^P17E,CL4.+@?-EW=<RJP<L)O.,DI8X
P6*=_9B!DZ*#N1 A_S:?1/U,H_LIS1*N#7N7]#HHF%!C.Y \@,6],L?6F(#(ISXL,
P"4$8H*-YQFM>*K;4R"\W" *Y3!X]VSP88+R(5XJU'A@WM<HX!C5W!9(:8BO(!<"X
P;/:&< SFJ5*WJCB"5)QZBVF0%AL <M>;7+4 T4*4#IIW:#HY3L/?6!AVV'HF[(=,
P=Z]X=,27[0:C?.Q<2!M%AIZ*>0PF1W0DU)S6VB]X[_ D0)QUJ&6 FGR]#K; IY]1
PW<.-13I4A_:I!Z8)5HBK',-PDC,M1=C7FTDYU(8MR_5HT"?, 4-Q7#4TD_VD5GD/
P^U'])=-S.5V@A/?D)C8<X8HBINEQH!WS(A[NJ ?&$V>K[H8>J'V*6%8_A*FE.C).
P=U0+_LI8GH54IKM.YTYB=P\TD70:1((+K<^W,R'-OYH!ZW\@5OC%R@';L"XC'@(T
PS4?2:&R90M"C5N"6'AE&2=T_2(8S)9#4<*-E?-*ZB/)+6U"$:Q3+9J%QB+>:.7C\
P\BNF*1%",RL\ USE"7':;P =I#C\<)A#LG\4C.$])FN^)!@!G;3M3G.PTEUIQ- Q
P/0Q*T@<9=VDV""9&/SV])/$#=H@3ZG:O<>)O(?[YUG@<<[X%@<;H0>$6LX"#[<3V
P8HIHB&H6_L_O!AJ'2!+V0'*=VYG+JG9D8P[1*';!#[4WZR^;U'+X$#+32S\\!^6^
PTL=+:E ZG:N:IED CA-"FO]PQ.OIP/L2D[7DN]R'XH_S4\A<AC!KR!JB<AG4S/_W
PP,#!P@M./,W?62C+-*;0WZ]FRI$[7,YYUH7Z.,C.AG?2'Z]8)^)7IQ/$<YF%%RG8
P>P$BL4PJ&*;Q!"/,"Y[T>C#/EI/Y&'SMD"*$6SJM76@ MK?G62*RJ-\& 1?NR+!I
PNV*DDWK0 Q=!\,K.$LP3*^QC?91C2OGV+ QQ2NW$.!6<C'!T2=J&D$RXO\GBZYE/
POO?21.E2@Y$[3#K<O^CH[XFXD+R1V;+ M,)LN<&W8%]_ ,@O2<P5[.GJ-2L]^DU 
P)G%JR=6H1(O*^7DW),Y+Z"2$,\CB(1-;5[*83N]B,;!4U!.>)? )ZW+V$*)P&,QO
P-GE']?\N?!2-J($5 Y$1+V>F8VPO$54:M7SM'B+-#XYOQ", /"ZD^(#*^,]35Q07
P7U>],@XD47)[DDRF@M0LJ[.2WJMJ]D)*'4\]:<EYW86DBW0(4<V%=,7_D%PC.6*/
PY'W2!2O9FWOLH^9)I8H6#;3G5ICNU<",<'&-%6!F-UC NL('.XZ=N:B?XK'F/<29
P8OYJ.&!\2*ST=K\\MZ=$P)WL%,RQOD6)*C-/11]7ZE_6<7<3&-!;A(I(WQQ='U.Q
PJIV7F6B\2>BKLW*]I*)FGS.+@\$7 9"JST$W%+<_R;U![:<OT*0?67;89J=XX7GT
PHFG>[!3\*SIH#:9CZISF,9-;4@\9M,K3N+#8*0G7,Q$!V?G)-9V2"&?M7+3".#AE
PH^3UR^:?''K^?NJLWZD<-[+3TU?(DO2MA,MO3J')@-(Q'+".85T_P%B)R>^/"=5Y
P($US8/ G ;8:]2_JC[Z1C4X'.(+!;N\;QW_VEL1V!Y3K^P\P0&+X=4P)G%;2^JQ?
P+?2E0S>)QP@C+_J8';"7>)DRO5D"1'IOB3*ZAG*O-PF*5%^V9[]W+'T&U\JFX/]"
POLFW)=0ON'SG& $P-MYF7TC<QCVE_CJ?C4@4?.1\A(1SEQ/S+XHM(Y_FX,$I* :9
P<X;)ZR*8$$F#PZ?L!5PSZV*6 OL#H1W8=%_&WFX%X4XI<V/__%U7['!WJO52,VQL
PKXP6%0">BC553Y4UI/,47"]N<&NX'B=M-Q5QB!YF64FSVRG"156L"F7 [J\.(45@
P@![H?39:INW.1M]Y+_SHM!9=\3^7Q!_'.9O289GNP/]"^^>@'QH@K8/=2\BMJU6)
P;R/'^D9'XNG3,]H[<W^<QNQ%Y_[?B@/'GR<OW;ZS4-_2U]7WTX7E"#>TVT6DN6CY
P,6CW,-AODDJ+VS;K'+5373<*L4<<!';O& <A6"_$PE/-R-(Y4 ='XJ0US3/ 7Y<D
PJNAJ$,&.+^6?JX;S'Z&HQ5S';%<]A?2;E+;GCLV&62O%ZXT!F?"49TE.6'X>3&X/
PNG?M!GQ[+9=WNB4D'>'2'V](K(!T5-6QU%]4=>7]=3WWEYRU"H>,TY\L".J[F)OX
P99V8M=G[+7O:GIW]6_MRW[[/C-WWEH4'7P2X[D!C+O7W?1!^Y:TSZXON>?WV'+6X
P>?=D;*R HKC!".6")@<T':/HKPT+IIS3"&P3'8ZWOW74.W',6FBE@@5@"$@.N&&6
PE;AJQL&R9 ;=XM_HD6)^^9" -A.I$X:KZ8CO](NZ_A"8=@M=E_A+&/)+%9E)_#(9
P6&$W+M6JF?PXSR)![\TOKUDDY;@<L-SE&<C\H*-/R1U 9DB9"#_;(3X,LH;^F/MC
P.BEJ;[N$(ZR9'/Z; <'4O)LE$IRO#V&4$Y^[$)>^=H5Y- 34DQ='QN#OO'4=1&_J
PU>CVZBW;:0R/*3ZC?_^F*[]3TE9DDMRR-=1]=BB,ZGM%#KWA)V$TEKEN]@*G6"KQ
PJD#\V>Y&TL4)HH7'BZ$Y:L-)OZ;R+FWQ#V]_'3(7/!+<_0UK&T?D?<L[H<XZ#T;-
P?F6$R-46//@=R\0I,@_&:7[.APY4@Q24S 1DRNUXLBH\ZF%N"US@R/LZ<^@ H\3;
P_^H<Z[O-0.H?&CX"+S""ZJ(M_RJP*SF8L8I+B'U;PQ ,=X-_D7H_2Y9PNM$>0"6M
P%\@^>E;(7/C4)ED3-C,<LT7$34>B,9T_3DWA6-=YI9T%11_#KEG)+)@MSPM=H)EI
P:Z6F]P3>?;JK0/&L89TWB[C[RG1G Y=+G.<+)NY_MI[7C4 K_9(R,-*-67XC( ]R
PYL$_,_;1UBQ2!HM.-II8_:E'-A42_7E./%L>.+@GCWK K>5J]U[J8,QD;C-J@I][
P!(0S9])ZX(/?%TP5+S/4*\AX2]GL.YNQ\(8"=X^]0,_+P@E24)30$Y<4C1-S@9B_
P:=H%"7L6;F4<=(=+/_GW"]A<'E<Q)B[W7,X-U2("Q418#00F/2C)$'S':])D@@4A
P/;2*#6W6GICQW*+X]8U.TZ&8-T7!68D+MC$T!@%^L<%_.6U.X8N0086_?Z+CQ&%,
PU8>/#H?U.L,'O\?D@'L6IGZT,)FPA&LF M6'($#*=/:D3YDWN@(#UF'6SBYCHU^J
PU:':E92=NLP4)R@=#$,[P71#X/@C!4EY!?S[!?7]%>=2=GEU/G+58&7"EZ!T>9+/
PAEFAB@G(^3\41!RA@^Z#=MI#P+F CZXZQ90CL+>VA(DK%1Y&-.DX41.CC4DR$:==
PC&'T4LS%1VJD&I6U@,VD71["2H?9H="_^:^H X* ;A"XNH9;/20#D,MR\E62)7-\
P;?EO2-[K+=)8WQ<(&!C:O;S?>2BWH/J[?<+L?K;YHMFRZ*D(>%;BOY/$QD6)DB+2
PG&XN]6O",Q2-NQHR FX!MD2_P9<,FQ3*RT-+-@9%'+R1T3-XT!]L$N?P&K(Q8W+(
P2B4BX$O4M<Q$PX.R,)QN.\[0GQH#4:O(^JH3Z;<S3;QRCG&':Y;#A;"E_@0+1>%1
PE!MA,2=4$FR%^['YT&[YC\B)#<HF$7(TMXC1QJ#[^84N1? L<^RX3=4T-JE?A&.#
P(("B1$O!!=.L?)UMQP#R75?31RH?"ZZ\5#\58R#?0J45U!=3F1Y3U1>/E"=UOGWQ
PWL;IQI.,8:)'ZG1*0!/-==O-:BO>XUJK0J&NFD@=B(=@-(&S_S 8\ILZAF%.U@Q_
P8ZM$'*'8[5\8_W4X,KLG>SAOJ3H^A<147T1\0#"8@PVF7 +9=N_]^CCV?V4]>!B%
PF[],A1(Y,2^GUY3=2WQ/I^E98>[@H.NX6/E:'.8,\4Z@.O+X[,%%18#8=**%-89D
PEB*7);F+(GD-6UN,'G?NO\%5IN>&U8=J;>2QE]'MH-\Z5A#7<A^:__ 97N+X WOQ
P#Q\<,\Z*Q+:_."H"ZIJ@;(*Y>TV94_:3*GY+H07O$G5=A::6[U3ZKAQ>OB\QH2,,
P[D:Q:W*W'?YY6H?!KNX,3M=6!/2U_FQ*F&XPD&N=Z+I/]A\,.*&%73+-,MK$%R-7
P+/-:?W:4?Y_V ?6S#W-S[,F.?)1SC\+)B_.'C]O2\@&5KJ>L7<#PW?KZ]P8J+<M0
PRE#:W[D_"<DPP,6R 'X(56'?2*?_O1)U>$H0@]B@B+)MFVB_WHRM]0'A(RR0Z,$E
PWA6P,<]VZ$FR<(.=JB"[@V#W%/6)X%LZR*8+TYP^D7U([O IX8Y2(G2,[]-07\^0
P\H4I..M=$(QR58Y5PIC6UL:N9;A_A!J@I7#=/@"A:1M>(3$8F,0\%;ZI>W? 972G
PS1M2KV7_M1I)220<G_=O!)EX!B5SV>D*OEGF&N;T!9Z)N]W^:'EWZ:Z9RO06$;O+
PLM:7'^:YT^X6LY.Q5K7XP&'6R1H^ "\XX&75N^$;Q-3*HL &6*@*G2C4FM\/RIYI
P<<G4O(KQ>&2_7 4&0R&OON7PVD3PE$?W@X):4]"GP_NSZ*O2V+!G@L=H'KG<7,.Z
P2KJ64=U**@$E-%5P6JUF:3CZBSS-,EZ=#'M6SQH,M\,P&:2]VJ9FA$K^"GO:= ,%
PK57:KQ];8(/_6"FCX0AN),71_KKC3SCO</S;,7V=.PN@5]/%ZMI=;5MR:']-J/1=
PJ#"*M:B>>Q%MR&REQL=(*N, ND5Q(,;YDTQ%NP+RI5YXKME?*N&8)T=!_U&4* K 
PU-G)[]Z6X@?NH!CPQ'Y@UL@/*1;8NSW/-/&"VD$'!B+DE;HY 1)7(63GZJOU)_VK
PD$U)SG/D6]!SL@>?C%+T]4VQ2XM#:285JB*G0N#.X6TBM_!L^AQ4XY6COTC_,6DA
P=+)&*/L-.C7W)]_+OI.!7"&&ALG[ QI H(^47>;*=5Q@-_:D:"Q/$"Y\W?+JZ6J7
P*''O\V5874F*P3++4:@L=+C\<^O=2?_C%=T5X<7!07?%0#ZQUX[5#3.PQP8.5=%V
P(=2'YC>F$TO2QKE-_1"I(0?>[S2P\:74LIO5U N A?_, A:PLO]-()E9 >)H-8)>
PJ2=[$\O?L>_W$JX9^,/1V5:4BQ.]3U.K<F#6$1ES>54=77NH[IT*4:"\_6\%5=Z*
P)(&?Z\YO]4'C8SZ#7FN%^BB=T 8@MA-Q4F P(MV61C_[?G_$9:E!R&FOY(6"[[R^
PXN.WTTZC]&XB6RV2S+PF/#5R9;#Z)I?<30(>\GD2%OC3NA]=9RN-5U[?!TJ4X0&U
PGO?08CBJA@.I&CW.&NZ<G-?/G6_2)LTU5>C4.L "B<U=O #AD$\.%*U@797,8KH3
P NAJ[W\(^_>5S\2RFDU.5P=E"!8$H=X(+>RC8*^S*:9HK.6_3V;8WM0!*0GOZ8"\
PCL ,O/6?2B7)?KP=-%O:ZPTP C?%RQ&NEZWU[Q@VU]<HWO/<'.HR%61Z[6Z#UD5T
P&@J0K5 6945:3;R%N3G^V-EH'T7Z8/Z[RV1O[R#H'CJW.5BRRJ^,F%E"A5:OLWID
PS^G3)"RNL-W0E_12;ZPO;:N/7X Z\?\N< 9&<^*,T$XJ[)9+DD/EDMB1LH1?+*@!
P;]VIOJS (&XFGE<RS7T'6R=$43+E!1DTBEH&Q.0V:/L :[=]5+WF"WN/O1DK%>X6
POC%*B*K1< </:HN">*^,JC"PE/ AYAH2[4_U_[EM;A*V7;LJOVZ7BO>G0\JS-DSX
PI$ *7MQ"+81.[IEH_5SWVY"=!PF\EP6#)4D_#5:)XS2;=JEU#2KM2*BXMP[>Z@CK
P)<HL$\"GLWT1$G0UA]'Q-J3ZS2;?9(1<^6 AEOUN&S]+ 6NNQ$S9:/R"+#K\8CHU
PJ$9X80_[S6*>D9LA[(9 7^-RLX2<++"G63%SSC7#\KE5$]@_9F);H+ [%@I-MP^Z
PUY\ZW7<RP\!+5YN9*2)]55<27;.1IBM;58=/2J>B4^.]M<Y$X%?_O/WD8Q9H;@#S
PKGG<81?IXE=Z'B.EG-9)2Y*ZL1-_];UAP^G"W5_!76WQ;$Z>(^?E1'[5QI1RP#,8
P'E5.A'N&;<5=_/ .>ZVWZV2 <;-G3$L7"T"\@GO9:"\_3SR@6%DQ9:AE#</XIV)I
P7"B4<BT>QXP(%^AT?%;3=D[2F;FFVX.WKQZQ^E-[=P N90D_VAPM:4PJB#:(_9A;
P%)^;B.*S !]QIB8R^U]L=P.[&[3L#Z)IZ*TYE7^R2S1J0MOFH<P0S/I/[;F-=@63
P=.E(4^C+7WK ^.%<TK66@XG3 BI<7Z;83O*[DSX'R 76S6C:@AT?4(4_;FS?IG_O
P8#!NG&54&&P1S-RX&?M9 ADZO7&@]#XYV$/K$\?XF<X@G@$"LL-^PXBFDHRN,$'_
PZSS6X'M5-JWC)V7#<XH?X3]X\<]9*8:#$2.,_;W39 @>1X:QB[CXN 0)Y[Q.E2MU
P%I>G)+->XFF3$+P/H,5O1K@8AV76[)UVU^:9'&J)[C5X+]':P*,-O@>_KYD!+G3(
P?0]]U)%88)W;;9N6IK-?1V[5:;/T)P5H["LM);V_8M+PH%[1./HV; @!VS+B1\O%
P%P^'J5.P1G02#'*LE*[9A&*U34E-F-2^,)9W"NF27_SK-)VU;(@4R2GR?_E(W>1H
P&Y.HK2' O0Q_T<[-1OMWWGRKHJ.@)>X8RQYM!]'7Q_3]#0$8:7[&!0G;)9<B-#FS
P6YX!&8YV@YX>,$+^L+%Y_?TSXMI;;$>!:\]1P>55YPWRJ$^'> 3].#C\[^I6DJ"4
P1+\29'_UQD1H-&6%>_8,3@';AQ')2E)G@=U_KN0&[MD.C.(:&%9/)!/\RNH0S8>9
PV)Z_&+KAKSV'[/\S"7K=635K#'9<*94J_JE)43@\@L0*%F8I>G:LC7X)-?39Q:+;
P.\XK%AVI3$DX,V.EV!>N4LMJ)CQ.#L=)8J7Y41Q^='"==<_N0 ^B5^)EB2/^OH8T
P"HS@!%WBNP!>8+\A'#:OE"##(PKZ0C_L9 S*B((EX52GR!-AH"EO)%QIAI="QLC8
P^ZF*L1W(L]H!S%;$5$48PD.W;9/[2<6"=OE_SL(*EB3+[ E Y;\,T ;/BM$.)^4)
P72&&.CZI;5[4R=9!:RE<3*-&KFW[X11*(UPQ^-J89G^,EG/@,C%74A*$^+4/.Z]*
P>,-W%&0486/V8_Y'3FJLST"7V$P#5@8)KTM-OU #TFG;/>T1^[160-")A;T,3C(6
P9TC$5>$\A#$TK>0TDW.+:F;6D ?#P&C=A%RF5PLG6K3CQ-[@]5K0:TBMMC9]Y*I2
PH >[;L\Q]]!MDIMRI,3!$3Q/QIYWSL1H;5\ZQ078AR(0R(I,@OFBVM 3RT7T2UO&
PEA9"^&2V\I# 5"Z2N3P91>&C5";$,(;M-,>XB)@'J5,185B%>-XN1J5L?IJHL5JB
P:Z24DI>X"X!*OX4%IBT&Q6C?,P%(8KF<A/XN+VBSY33Y3?CEH_W5%T=M-;/M[LB!
P!Z1>Y*E9\,9O-*DG*5.\UL!<%L[Z)"@ON25 SFBMQ&J11L\^70ZJP'NS7C!GO]V?
P#S:T]U7_OC*?*/@E,1Y #;"9BUQ#.U[WH!N--(:6L%\ #0KIC_>SMT4'DM,L0= #
P1Z'D(3'.P>.^L#CG.ZM,6>&R0X4MRS3\X<<A>(+(*#@8EW$;O-W0@=TY-SE4Y0/^
PJX$1CO_3R#KLSN_L5&T;EHW'L-DC1>1:0CO$AZ?25JO&-L)/DPZ6..MB&_&;9QO-
P((M2[6 EPS^";5M:?A'MSD9='.4W6%!F_U</@&(KW<5![?-WI,ALK%0</J\NFTI1
PXE6 :-87[%-B!>'2EIBO=OJ4,^7_M>(J*0A"^3NN2PE=*A&>5C/]'YTT8,Y:R +.
PS?EISY"AG'B$+#N%F;,0>_4,L7Y'A,=/_O[V[F(;P3$Q0IPP.MCL*F>0W1%4"@-&
PFEI=-'AO:&(&!5&_U7)J"^;C6R'VT3%S?>M/@:!<;YJ6^?P6.:#RCF!3:D?]V,,I
PL_@$PN*JA\UFE=_7(S6D/R38)P%X':-SO6SATV.S-D#B:JMQCOOWP3[_FGSMJ\T/
PF*>D\9GIM+'K67I?;S0!/-N27/ >18<_O>.0L2K/7QF>F];LO#=H?<;*%Q;4GRF-
P:G\O0'YU$@-4'V($:/6U$E(A*(^G-XNHDG<@7GI*ZC.EM/_*<X'2SM#Z0N[F+SK.
P'"B7-![%*P#CN60&M^9H(VP[&$"%DCU0^@/B_H1:!+3KLPXKN7%D7*VN?8#=\CCK
P*\7R C._"'T,HNUN1R$(M2QF%ULF/&)V)1&6$Y?[&L(J=!R["_]G80#$?1#34\MV
PRR?X$,=-NZYT:VWAI$.XCWLJG8?'ROS!7>T=#74MUT:UGF4?T![4JK4\I5%3ZW#?
PQ].98,YKG6B8S4S6V4AES;3M38V>A_ME,QO<VAPTKS"6<RG)0PWB7HR+4>\\!.<C
P-W4&KQ82SI43-2"?Z;_$UF_$&HM8L;(_#3/J)44_5.0MCH>NML19#,-1<16[C3.U
P4>\-C@-%2DQY\%,^28TVYXAP#$D!CI6E6VZUC% "J6PLRS26&B-<%&#< 8IQJA*2
P>2CO>O?'C7)P,1Q6G'\JUTIS-FTUY4EM1M4@%Y_WR8(K?>Q6:8<4N1?PAOG7.ERH
P..@-E@VM[X9_::H1-V4C 1\6-! ^6+9PQIA=SMZGT'UJ+%Z8WNHVN4;+:[O2)/N<
PN,&<"Z-"\]HD\):3PPE9;/YKI:<-V,( D1I-HHR:'4[.NGB")>^\TPJ'7IUSD;XI
P^IK!82%S\QHB!J,D> 3&D\)>V$?Y"$WV;G]6BKM=*ROSWM'F8E"ZN8 )SS[LZ4!+
P>/RWJWQ)UQ+&8'OIXJP"V$0&JYKF!>N<_6MP5U8X2=)Y<:[B+V<YYA?;=A(9WR)_
PACD8"DAW'O $UDHEN7C5='YKTGW_T)HI(#LR]@+GK.C:N"K+D9R+8MN=0LQ[D.T[
P*?\7_7OG8J"=>CL<UZ#!_'4NW7C!*1S8-#,3ZME9R!)#EW&GT2._+F#4 H+@B?>T
P45<L=7?$M\K)TP[94Y?.EZ[MBI/ZT1T6),#EY**)S-Q9$4&DH/AIEV]WH(I=4YW)
PEX+=2$6?UV1<X#<@F)'H$4Y?77X<7ZV#L)'?R=_^TD 1I[MOJ22-OYFTJ3G$_1E^
P#W?4,_.><_$I))8XCH.6E)2P0U'=36V!/=4HTY<COZRKP1;J928M<"07)!4/ -*:
P0*NFP(ZQ)L.N=>\!!!1U&Y26D);SV75=C%4M *<.GH)R+R;%],*\^&XX@Q3-R1SW
PETX'W8^-3[L*1W0*W0VM^WMM3!"88M]AB>1V:8#.G -+A9X0@!/:!D[\'?0#V+GU
P9AC1YO0YA>A!*LFU<!02Q(PQ&19KL<0!W?K5*S[90V9&!SUV(I^DDP:X8$+.:Z.#
P._:BWXM,-)N6=HGSVO3Z8HHR"CHW:JA#14(D@#AB(12>?L3A)L?4.5LX\R!/=B!A
PCCCI@Y3]RMBG$7#43AOD!Q+U6>Q'.+I7-"TGIK_)<T0=T43>.D)4ZFS>D"T<U-3W
P^T2]#][A.]L%C#I'XJITO]3R#;'Y=G?1$ZUQ??$EJ"3/Z+O_W,!5A^#5%;/:^2,7
PO=^'EI&O>@_/O09,,#[C4BJ14DM-.:I1FYXM(QEBP+I[M_,-;CW\>\L4)59!/D@J
P /?&-\ZR_6!&Q?R(ES.%CKLS8PK".H:QEM0!W9RB?%D$LVOH,Q2.["K<'-'F3)2I
P!%BC'=(%W[Q6KA16=Z_Y08D=YY_70N6$1#?@_HO4RD4Q"U>?Z'I$7XTP^#=FB,SY
PS>6B6_>%9)9BFGT%_DH_[/CM-P#)WGQD$Z']<!RYIE5T68S]Q!?NU7;#9UZ@6/D<
PZ^5>L3[8$)FWA287@4$5O WLRJ-DV<^K] ^ZWP]ODCQEQ;<RTG!P6V<])P_5,I1 
P'RQITW7Z%X+VTK@SF";"/U,3[!)#UU\>X"BTKV,LS!YU5PNO9AKL< V^,[ZORZ&0
PR%DS90]K_PJN$WZ94$<JT8I\BG-<D'K2T3UFLV9^,25>(8O_J+A# ONQ"OE[TZ8-
PVA0O(^X1QP5-N7W^J2K\GH#0:Z=A9\G[I,0'+8_35-9PHR"H:;@@03ZX!5^TXKU\
PL*#</X5S_12?G(J>#(W8$IET.C1RZB<8?AZH@<I6*05TS#Y110UR[I&[N*I=J1Q;
P*KG@7X)$A5ZL9E7[,(AJ_/!9T*<K^^UD?ERI=R(>>G 3=KTP,73)]KQ ZTU2D6;%
PGRO.*_4<!1\W;RED_DGR2I6PZH1)6SQY^EWP[I94=PR1C.L?HYKVVGK*AYG3C6V'
P%.X>1=F8!ORYSJ-T%=]GVM #=R:;"M=S!])&$08VVK+_XS=8QY-GJU>(_Z.SVX[L
P%&GW;KY@SG2)&)4_-.[/HD25+7#='6UX+.>1$[#I@R9MGN91KI>>0VW-I'I@N\-]
P>OA[$%78I&IG?_3%=RU\C7.X-%>J'_YZ/(:WVSQ^T-.B!?XFAR*P&^4C'[H/:6P:
P7-EGY->=))/O'5:-9L/BU<$B+9/)"EU 0X:-/8JVW-%^AW7MXU:GRDM8UBH@%?P.
PY63?.U'X/-(K-+UV="[BB\_ ^D7Z"Q=C*F[NLK#]=1SKAKLJUZA3E?';2L?,A091
P-=@4I":R\ D=+[%?P>ZD0LW&3&'X^8X"OCF V')7VID,&C-V;5+RU0&+,3P2SH;S
P08;LWAN.O%4_D#M5L+*U-IV#!@,##]T2=9.WX:$:N&PKD.N4TJ4KA_=Z;!&XE4<[
POGF&2?*%7^@VYD 075196S5?[4PU+;8&+L+:%,XSM/[;4I0#=4G\1S+.+5\;F/B'
PRP*W+3:@*M)OS'K5,'V%WBV!5N;#<@,7;KOLIAP$GH&-61/86H)L)%A+IZIHN/%!
PON4--(QI7NT3OZN8JP44IF:O4"PEB;,/C,I2A(B49Z#[1?LQJ!5Q0/WK<8UZL.W*
P+!B+P60O,?I3[ N5=BJ>#_H,;D!\DF),:6U+G^4C;+6@HFQ6PT#;(3;^M3N.2?N"
P;5&'C6]#1;^B8F8_"5>@43M:.=M72D/UIT+5:3\XO+><0Y^*P-MN..TYFLV^!/I5
P+V]NW "WNG,(3Z7P0&3HRP@NU+6W4D*.71AAL^4V/?AR>1Q\D0DB)P?<F@ @!,4T
P%!V,02X;/(YN$193S*$BSC C^U1Z(U.] F^1OH]"(K_05-Y9,4+Y01S$Q[&[QQT_
PZO*/"E33;/W.=G[8$C L/&CG2ACW,K?IPB3_[QI0=C\*ETN-U$]2.)GAZ&7W23F=
P57L+WV*O(-86O,WO9/R*Q#D=%*H<@;EFL@/Q,=X"M,QJSVY<7'S<XAD*9MI=^YM"
P6?9H+QR9(H:C0D1RFR%L&VR1*_@H86,_(<UU<,&JX UQ[126'6)Y+:BCLSA%!)?7
PH<"X396[X,V0L]XZ$0EO1(\G$3(!BV])@JQ41;YI >"0A@(N)F#R^CWG5 H:QPN0
PF[9/7^5LFA.'ZI$7V^EEH)/PBY&?H&S@F2K39J'D@Z!V:N&FH3Z6_UL,Y +.2,<%
PB36U#1'^I.":2.UPK]M]5FOEA,@DOVJ4G=K(WKJSJ0Z=,:ZM3$D VX>-9XZ)"68P
P?&2\P[6!,/4P9*]^EP5"JRDVM,+60%@ J>JY?(&YVX0="WX/% ,4>MA"S/-AS][S
P<W.T]/4RIWTT  %DU&+%DKQPS'J)9VI[\\W ?V)WJE#+FU)1D5_ O8!C.\KS-6D>
PW(NLUFQOXM:&_SM4AAJ>',40'0,3WU:)N1#GCR"[C_"EEIK6!ODPFS0@<+/*'3P'
PCD@[I*I@8(H"+L+:YX;(UXVK_B^!.C!"1PID%B_WM9B;I;7-18E%[ICS&9BY_ KV
P\+5\QEUO33!U8W/5WAZ2R[?@^MH*G0NVJ/:&R'<&]AF:PTK6]1+R0_-+08B8H@'9
PVQ*["GI\B/XA'FQ@]2NX/X"/-<B.(Y>.@JX1KIP0@U:OBSH=$'U2<\CT&YIMUBNC
P3HP)B \&/C@_/@^-]JMB2Q+R)@.P[GJ_:IWVJZ56-F ,R A?6]03.] _)LF:HMN=
P\.8[]3/BT#R*,%0C:J,2+(-/NEQ/0/ GA;8I(WYRI=SB@?$KV_RU8,36NJ=>M*@I
P(-;L!.C"SIZV+XT7,+W5!6R*#(,4V:/E_XY_TU=:2C9038#OE PP.C;3?#.9C/YQ
PI3F1EN*ZNP??0M1;=K<W@XZ+?Q5;L\.:-[GQRJ9;D;DF3%6RR%>YG[XTB$N<EWZT
P-/S05:RAQCZPY$ =%6>/-$QJAY=X19AD6E:+[&C4]9U!VLRC7"I86MIZ$Z8U<[\.
PV:L0!H;9&3W53HASLO6$Z_AZ_X/,(UNJ[>T@YS$QX.>MO0XBFUFANBK3)1_X(=8D
P%;^#Q3._[7@ GK9:@Z7I[]>%!7;TS0MB@R<<$>,(-L,Q'98;R,*4'2HK*.[,#J4S
P2,6J)0-<?:[:2?*&Q-86L)G4OKV;Q$Z]9;,0FB@(#Z\@^)N+Y24R7<62DXK863(Y
P':#6Y]>=A@Z"XK2<O!P.8Y9\GX<]31F[PD8+:<9728\5G&M=&V C#^8<WL3VK1=\
P'DL<O$)5FI'"QY#13OH<:94=;N#$9WE)#/4R=R>267(+:V>"-L.5@H((J88G11&W
PH3R5I0C64?418%FR#=4+V5<$H]B5[.RU&[AHUYM#R@@FK:#CK>P8HU]1  %*^%3Z
PWQ,'Y)L2I#MH;_S$M]E<(^)RH2@/8M'B8UXJ8P4$*$Q5=B$$MA-<X9;Q<*O"L,5$
PGR@FLO1;C3[=Y*:^S&X2-GTG#7*4OFPQJS8/NQ+59.?>)DCM$\'][O/P&7.1K&Z;
P:EE''Q"'/X]I+Y U CR$K=33F;,8R5X@;"#J47S/P35KID,A]78#_6P@J631.'6^
PMF+:0HJKX"3WNY]^G?7RK%/$>+O0R@._;OW&1*HX%+/)8'U8YW(7X!3E2SEY+L$W
PS;0I0":^&G;BMZ'L!QKZC[_)NWP?R_B39%"NP.JV'N3Y9 ML6QO"G-EEHZU&/E#E
PPG[\'H)/.(9EOL2D6U[DT\O @8,K^LUQ/GK]Y+<\A06G7;X'^C,^7]^4;@.0?3(5
P<]?N-^0&+,@NJ3?X/DZ'WS('\.U\4WZ17_H+$!MO&FQ2TC=I,?>?U^3^7/?%%@>=
PS!M/'TE-1+:ZKDI.:_B=YARQSZ *G2XI+11P_.>_A&ZLXY(ZU]-NT@%&HDOP%CKC
P!%I,*,I^T*.VJ<\(YCS7!C6!;EH:W5V9+^D(/RN?;Z)!3:L85_+V2<5-YU/%2 4\
PPALU?P@*84"HC?%Z52S\P#CAP_XNCP7#8*X242^MYACIJ]&Z<N\?AQ?$2'$0Z.#&
P.Q+O]5$=W_) ,@%B(&2$XO03,)LL;#2]3$>D)HJT1MBW&AT8"AN2-P;6X!]F+UO.
P<#.,^ FEVN5 FXI-&1-AI^,%U*R"&YZ\!V-6RGN-J,E_=KK'ZFFT&WR^:P2^N2/A
PF NPYU!B22_:=2_IP$A"%("$K7NMWB33M^KA?NB]3VX;5@2%<'"+G>*]I<"6R]HD
P01 [V&"YS<A9EOALF*/2TU/1]8IA@)"1TCF$LCE);D,LUS^X"95>=G9I3@!E59*"
P&QAT/*<70:;\G2[U@A=^E?2).L8EA8A1:_I-^\>JA=;?U,'.WW21+47O%QC C<0H
PWZN!*G2JH=W_9OW?$B:%2*%!%:SJ!LS"".,SS;5>V*M$1K9 YI0]ES32",I;+&":
P+SW4^!?Z+$?K?ZW],)ZC1Z($^<+SM7PZFE4IPM^C7@B#JBWE6M,-EUTEXH^0N?.2
P43[D14*.UC8>)$_\$?9S:)K,%>PLV[+$X_%#7BA3^HX-*@> QK&$)9L(/_-*#"_#
P8L;_U=^GB\'6=,,*[+M7X:-LOY=54"6]@JA63 M^IL_"V]WF]T;'QQ=^+^N((+&L
P)RWR.X'R&=^PPC=0X@&XF7D(3!U>OJ!,?_Q7:I:68T?Q3)MJ5^6?\LNRX F%'!4B
P$=+-P# E/^/M&_752<N55=HZ*1*%EF1;VK^=+4C=WK&@)_+&GK*^:6JW'U^B.?W6
PGOU<0W;7WUCDAJOBNDQU,6$]]$=W&0#4BH_RCK+HQK\3X(K1V(* MM4C6*HS8;-3
P^Z^3FZ.XS11<%CP1V47F( AL%PU,<?*6,N-J(<""D;R"?PY&5C9Q2P<%/P6S<:)8
P]03JM@:==]>4URU6V<^-UH9H;/LM-$KN*B":3QV*7F\/X::66(%.RUB*AEU[C1'Y
P4*N&Z%/O;E9E^>*_"73,I%?6+=[CAW*,H^*=ZD:\@-G ,_@EZTNNSD48Y$;\9%1Z
P*&,7PM'1'T$E-@E1E9P*0JYXZ($@"97Y]<6F0@>9#.?-:#_(]>A.:HH-/D:R L^U
P9;UJ$6.K5VFQI>;].@I0W"F&#\6U7!.$_ ![3$-2H-3R+#D]F#4<$W2,V">;==]J
P)?2_"[B:4G162!7J'7B0M3RFS"4PR[#[_JBWCFL!@TS>=*W%###XJ/H(?)F6SU*$
P[KZ=>EDF^<1 &Q*I, H#.=0%Q'L"OUP5'=ED&.;.__1<XC?3!<$!=16C:(:VP%^\
PI_5I'7CTK$WH>ES&BLNL<1'/J>\MSAH#"T6U!RH,>"V9:'*\B7XT!1AF =8>E9;]
P^0YHHF&571#>8KH>31=O=#NM(LQ\-UXEBN7"8ZM$SN3<]MM'+1FQ@1GM!% $KJJZ
P7N+@[OM''EAT$!<OWX;W@''VBJWL6:Y:'B9,1> 8N^&O%O9BG)+FI-A[7>%:7];Z
P".DK&OGTAN+JS[CU[DW&A!_K"BH('C\:'*T6&B:J3FW*60WXMFD2DK#J_]G=HF99
P(^TRQR$NI@#>)Z-_G[]82#L?0;%QE>>4#1!=<%1R)C'>=?4YK!029URM18@WOV[A
PU5V1\(@,2JC%Q,<7?#"Y<3T0E&< V["ZB>Q)94,Z!P 7RR9&F9[V?Y?1WA68FB9B
P8[PGHTO#/C;&[ (G)C2E<@\X@=L)06 \"H:CUBWS)GS?!=4[FD0YA835V^#6AB8D
PT7"_F%>R4'@X 8NG&5>2BVE[4M(?:^D7\!W$FCM?)<W:85'[7)?-70M7M1T^X.Y0
P$>\2[IY+IU=<%%Z97!'>W>Y_47[^+@ PKV15F#L\#EB#H6_*AC!G+ID$Q<]3^?@O
PE&H*GNFUFAQ@;9R83%/H%TF[^9<@@P@U>_&,O;D.58=5 _6Y$G2V:=+@EI0IBG;Q
PJ$M5MQI%R#&/C0,C&./(!H-RQUQ]6=7(M?RZ\=-__GU)A\';9_,+<B)\KD\!">0T
P1K$8,<G@F&N('L8W2OY)Y)O:6<P%[H8U_\;?P/O2.MZ[97'9CX'U_Y(-5XKNP6@*
PPZ*?V$JMGMJ21LQ)^S\3B^@[D64>\*5[>TMMQ*=?;;6FC_"EBFW50(2O^?%#H_K&
PQ.O<!VBJFDD%V%,2H&O#PAA>09(33L!B<KWQ0D4L,*VBO>X#H[^V/0Q$/0D@4\ZR
P &GH/PX/Y):%1 Q*)"[I\.FB'%PS^,K;)PR>:=($+A5\AV]/;'NV66-2]^;:/L"Q
PK'%*<K_1U]@O/Q%'V)W75$_>T+?9;Z./=X45)[.:SJTF!(,W+^@W5*?WE%I="H&:
PD";8O@OUKV+683T/YTS_1H:87F=#=27N7G-ZONT>_T(HL[WVPIQ^)KPML"]=\2-Y
PIF%+3D1VP'%:IA<9;GR,W[N4D)%D8()V4BQ 9TMVJ9DVO"GO V^L#QX-=,/*Q)X5
P2:&,H06T1XU"R8!LJ-FLO%G&0"1QM'E-*>FD)V4)=A^B 6#G; .>057;*!_EA)MJ
P>OA'(G(<^:=C%TM/FI/9 3-9F5#CQ&8UD(KG=['YQ^D(J-#PJ>,S6/*KR;ZJ(73P
PX!7OEBVR$03=)?WS_Y\9]X1MR-X;11M9/@?4OR<W!7HAYD 71&43Q7*.:=_>J.P@
PU'AFHX7+>8C:]%B,0%RZAWOWFHM"%ZXU#-@CK6V #]_D4P(BPWK!KL7\EZ$7%URP
PD>E?F^CL\K 9_6].$4+8=AA&^4ZRL4ALTBZ7JICCUX'-&/@E+ NOT5KPY UH?.39
P=EI/5ZP1+M)'#ZD]O"KKGHL,%'QZ+I.K^_9%9K\T/CG3RAI8MXT41;@D1]CJC0[!
PI_,2</ZC<E!GW1>A0%GL>XR*E!/GAD/8XI-^G(+%1#8U7[DT>9+=IJP*PN]O+[>R
P-7#\I/P%X]*#1B0;%HM<J\6 UWA +7S#PYS1O>IFM-;S+_?]TW4T87]S3<%I7-!!
PGO#[7+&D"E\73YJB+0LG^*<UDWNV4P\<O)7'A(>>C.9>QV0FB;MR9\G(OI+7Q15V
P*KE]3C[IN]RQLH>KA@(V!#?6V*:W93GIC0NQP;^LP<<^980&3,@YPNRX6]:XJ$SC
P?X]-=VZ[/P6.\JXA)YQ$RA?1#8T;9J?(0GT2M,D_QT,3TE2'U3CDX#"=<\LE24MB
PGZ8W4\^=EARUR=8-G=_J9'4[HT$!B/LK57"8SRDA>V(:Q8I3ZKY(U_"5+H^&BY)9
P0=#W4;&D273(@RLC09:_3?ZVQ9=)2PZ.2K<TYA%]%>N@8#/Y)15OVA"=#1SX9UES
PJ&](+,9GQ"LL<[0HB9V>6/?>(QA!'XS2NZ"5M8B*U1&TMY_T; ]$NMJG(I<6]2$Q
PK*=HBB/I">V,"?BV5@O%^*8/D^*RQVZ/%F9I!;"Q.^N%:UX"YZBFS5]I+*?UTIOO
PBWC]Y.+PCG_=2G#>&0M!V+X7Q(H5M[B9/$D_&7J[*R0">)?" C(TR#LMR$S/*DAX
PG3;2(9DSB!0!*'V8%VLQ$4A**$#B4F0-W>2K?=KH!:T7%DXTNT2M9PAA[>\Z"ILO
PT$JS(2\_W)AQM4Z P_4EFC(B.MPBY=82S":*N2B:$]*^I;E]O?TSU@4:[3\\.),B
PZJ8F.%/\0XEM0]AG;+(W8S*LJZE.+9H-"1:]AH8SH6^YPR0+^4]LJ&GR/:BWO0CC
PV=TM4R9_A\A1UIB6@+FWS2P_WR7P/S8W.KV$L_0(U9".WG!,A10WB(4CWN2=^7$I
PG=5&3Y?.TLR!Y^HVP7'R#;\C5[#R _ I=:C\$_]9NF#$_*7;D?W-?/?9VI=\[6E4
P!+<<Q82:-XB"UZ'8SJXLY@Y+^N3K QCIB;:2M(U4HY^2_FH$JGIZL*4@.@31*1.R
PBL8F,>-B$5G.IZ^29GOZM2;RKX)8]BG3&&GC"R*9Q "@<#2*V.Q+SV7XT3(QW7OX
PQG[L27BZM1-J:$=5Q2*R^1N#-;#2" ZE6)BM1?NY\WA80DZH;O? [A.QJ68SWW+K
P4X8!>FA,>G8M6NZZ04AL4%;UMKY?C[6:BY^^FE3@3N$%ECW)W .PN48(P$J#<@NX
P+?I;MW;"P8CA\3&4G/$YD1^C23IBXR,S\B;_-:^8ZOP0]L?#27FA8V-BI?K"K^QA
P6AQE$R\L"9[U,K5$D:5B*,OG?.B%21):H_$T;T+9<9-"C_S\=* $K9:_H9%FCZ?]
P_I0]Y;.CM%PSS%N'+HIP%N-9;:HLZ_"MC8RQ !WJW.W.1^IYN(R8.QW1AYQ<\I&9
PVJ4]IE15_+8+QK:O0\F8:&3QG-K2Y&ZSAFK4KB-MBA-5CT6I+*+Q=C?\=E8Q T"0
PI;0L17E]_6?GA+0T;@C;*&,RX)9N4^Q%0@HQ[]]1.]KY*RJR>]5A9JS\R/^8=O#S
P&[IV-NC1XHS:A8N 0@%RE@MU7BCD<E3B)SRSC$;M)<86?:6A_K/T9PV(=8BQ84WD
PVVY,)O$(RRD8<YWC/TUMLIX7O*^RE&:Z>+ ;MQVA.;THXXO]C&4%D6JOQ?>>JFWG
P6J=K!2(V6)%FO;V94BHYH57ZIDM8E910?6NF"[NF=-\S+C,])ONP^QNIKT@&CGYY
P;F=7ZC(K8WSGD'$@A Z1TO/H@-<'HZK2@7BI^(."FYAV>FRD;!DP$S]HZ%Z3M[2Z
P]*&3=$00UVQRG/'?,!??^V@Q(>30;U\R.)2Z5;Z_!^/<HC_ZXKJ:Y6CIL.!U.1=Z
P[RI/VX"KQ?3"[[K1]P#K\2F&-2%57.%DV@E2E1+&6Q7T34(=^M+W)M$0>'&SP&K<
P!*LH>^!.H<H %$M<_[1*EZR;$W_I?BF&C3ZF%D:+WN>6HCBX#.22CJJX(7>=88'B
PRJ#8IJZ,RK@%:^!F]MAT/^>R@XLI>I(U*O6(G"+6ZS?UUHQP#88S;;TQUPY=A*#!
P$M"\0RY9AU8H")9L(@&U\OVT"Z:<$S BK&VRB^M4UF]'\ET.1E=FPA-5GPG::*Z1
P(YRB F689A;I0BKWRB*%+=17=R(M*9;8.Q$9$"@#C/W,;M]/H$\MAU_]*Z7OJ:]2
P,6AL[9$,C2^B6,;1QU&,\'@ZOZV7 >#&=(!JI+N:07UI#4"'ATE.OJW9ETHCO4VQ
P_0(1&+<)I?$AI;LA_377EV*R!NB"K^PLK^:K-N:E6Q[G#D18!8F$+)K.^R$BS6_0
P&SWL2R(73_91<>I%05P.=[S28/QI5K@CK9FKL:[;>E##G+9O\LPW<"$'_,FS.PBP
PUM&CD6U) ->++LJ_.U[L6)[$@>?^AIL':HTY&U-0]0DUK(:7\UQ:C6+%WV Z7?:3
P1[(=L2%>2\["PY9V=B7X/ V%9;=T9 MQ7;MURJ6 >;2BU"=Q9*[26E2*$J; E=BK
PLVTF?R0B!6&]!QO@Q2E(L ,MWGZFGV2B]G#3TZP3>8*>LP?"-(ASN)WI[7Q4FGK@
PL_QM-%Q";+!M\I3_QJF4>-[Y:Z:0=CQ)YZ("9]O&UR4[) R"I:4F4G4>.1L%@HW^
P9)CP1LV;2"][(UK48&*EKJU%<N:5R=NIHKS8'RJ-%+I<E /ARK@ M%KX], H=S[1
P9J(LBEP5#Q#2+:' QQ-(8TL8[;=[8065XM_J5/<G1/W!6$XUB!$#R02*W1 =+N0!
PV/ZEJC%QAQ]0HM6F&AS?5KW:IA]H I;8-_FC*A+&<?CE444.G$6(Q'W2H.)'38RX
P*93_OQK#<WW)TS> CNSBJT]E@]2O83<2_C= [!5??9";GYS] TR&3SHIB)'8F( %
P]EY):64@-X*$6C+8 3Y^/+9N9W*.8:N2K47' [63FU6I6QYNWZ+1@Q-@L?^QN31*
P+XBT6_.N.9R9)_8NE]_!QK8TW8P9RH-,+9DB96.0ECR%<BID4W9P'?O[7\:0LI"V
PQ^JN:^0D]0)KAW@MBWO+$5HY.ROXAWS3RS2""_"=R(=HI&<_M=8]?;XKK/XN<3@0
P>>Z]\1>L6+W_TH8C)"X\Z#O)?0:L!&Z_:B/ZZ+6?GM>$6-G^U:#(/Q _?^60JTQO
PV%K*:-;R5=WU*AN2B^?D"):D$ET9IL"(C]OK9_)0?VJ8-0/_[-I<!L$EZ[O!$+@?
P^4.^ &%8"N9;-1./V7KJQ7&6< VT6D'AUBB'PW;/LZE=J,VRY($L?%@!G;7Z A$4
P_S>UD65WOZ%%^ 8)?+&D>)T8UQ#[^\1B=*7I9OXW+IJF$7FJBRBP^!W^<HO%E#5.
P2'M.00L5H0+I@KD[_'5IC1+4:DWY;)C(6DZER!X>''M]VEOJ]W2'8<^PRV%IYH!L
P@DRH=Y25)+!URSZ-1>Z'-[VU';3A7"&JZTF8[J<G.YU^ 7JA9 A&"DEA)<KI)PFX
P]61. (3]FB,B@9.+W/25A A;#!8]?Z-YB"GC$25EZP%)@$93KG:>"-WC$XBUCPOX
P\JJ:CJE!OT&(,5=F@X'\'X-FW"KD; 2A$H?<][]ZJYC<&J(B!0>]7+K$DV.+QUXN
P*+!],IM6YFJ2^M4@_7JS7Q>R;?H<!1C_[EHFJ74=B[+-\:HH41P3:VB\E3N2IM9'
P"OEK>U2V'/02A@?F+&Z8BD#&]>[]2D52L)9<QB  !:K/Q"_=FOC6_X;?9&:AUW9K
P)V]'7L^18#]5DHT;-LFSINF=I92DN/L"<%Z@-ZHFR;K-NG<(@?/C20>I<;[TC;L#
PD5#.<D2NH7<!JPB&U$2."*#C^AJK5W&*;8=@E7OS$HVZ4@D9DI(/ 4";D:7<)B)P
P'03')M.Q&NOI&=R6870K68UBL-5UI1O!'F0\MJP4R-=H6#153##.A_7OQU0M! .!
P; W*.K?,\E>5 :M=J6W8E>JPAQU\NB>4=;"ERCQ& D$D^+'%,BIA04Z# ]$8#MS'
PB1Z86:0T%M7S:@VLP @F)@P];KE"_X.-[R&\WA?4G;TK\TXB*602J&:>6//P%<*J
P*NE=L]M<D+,.-;RBL\570.OU.-98>'RCNRE&U2@A!@KT+7DG.6I#";BVA K5),_C
P%P,Z>E.>5X(W$/F?]UH>)FY1<_R9\<WEU]<:E5D)W8X@"/MXCK]\D_ R@2@="GG1
P//+;M[-F2549GYHP6+&'7Z-"\NH7A(E=IX7K9F42V/7_J^^XI9]1AI>#2D8=?^5Z
P0$C.#[@_!_\FCY*<*14].Z5XCXIZ.>8C#-7BC<+S^ $SQV<3HF:L&;!$47+1RG=D
P4TSNT4 "X0WI4U/7B#/U.?Y>_V[BH#3KVC?(Y^<UYH0U1,CQNDQE6EE(8TKB@M<)
P@B$UM *^,?5G/-'T6SBLP_S0^TK%5I$+QX2+\#:F5^GX5+RR*&R-/R]CHITVR-BQ
PJ^L6AH?FF:[&>B ^HUH\?)=U]CM#BA74<,U4-4*T5_+;Y'C-'#,]ZUDVT0Z:/TGT
P^WB?*4N#ZH'3D2VTP4+:1$+7AA %>F-E&07 ;L?SK$I&HW<F#M/2-V$B;R(Q8R-(
PM"!4M+/2G0Y)N@"M<=3,J!UE/,'4LU0W3@0-$H*],B/BF+LE*5JZ<8C*JC>7*!*/
P2,64AJTG *$YNF+/K9!DK4KKQ J6T5I'U^>QZN5LXM&D&S$:&*G+L3?@@[)F+1DH
PW:4<* QCQW0%F;9K7N7AZEMF769XMY>+]Z+ 8S'JA^5EH%70<9J!^2V6M8#8EA2$
P><2&,R,+D2O;,(%5YT8F:GJOJ5#]7W]*WQQ;0/]\0 3TLLI*Q_<'>_%>=G#>T:QL
PNED:J_ \V=&N3\1NERSV M9?/&0<LBNPCL,1Y=#$N((!V9M-9AK,ZQWL!T\R7V1R
PFWB?"AO_7A#>1-&%!J. 9FLB9"V,X$=P&3_H<JRY\C&ROQIS 0JEJXJK>6&[H74]
P-E4^ZU]VR;T!8HS6,R>WF0%Q(.]UJRG9I?_?M?S6[77U^C<N<TIHT_6Q 5PF3X.<
PFJ0*/X"0V0H-A5?\-<,&33W%MSXE)3@JO #5:U3WL& MU]C80EP<_BZ&$TX)MUWW
PG3W7=6#I8?8KC2+[ +O*#S'5F?^M<06&G#KV8M5N_#ATQ]B8-FN"T U+/TJ@6]!R
PV& /K,N%ON#3MV_F@KIT_]!\36V2883(.IV^=]/]4S\!EK1__:GY@:G55=X?^ Z4
PE93D\D@S6UNFLN.Y!"8[BG@(1A<=F6O=:\EA4L]2I,++5GVW&8/9/W\0^"Y\X7.@
P*SD[$3VR[%*'#H1]U'-C5",U3S4%//:6UT<Q1X[5OG^CC/,$LT+X N22_<O,4@'X
PW$-L(U!<J84I4?EOPJM9IWQF#'+MRCRFKJ2G^R@H:S(?OE!*+9 NFDK#N7X&"K+D
P^)H_)^NE+3KG=L$)BML&#\ -;8,>NOMSG2#P?26\]BXP02$_--CD?:*(9&(%LUS8
PRM(<]G_ []M%B9)H+1-_$MI'_H<!DDK3/AX5*Q_F"NN+M?IMV8[E@5[SJK3P3[%O
P*JT;H* 5//E<2YUVM]!]2PG04:=)-5G[9),>N]B22HZ4DC<KRJL23V[X7(?[;^T7
PT%-1:_.#LZ_&*V4_V)K"#]7:M"X#A8J0NC00Z3Z80Q%F3O;A#2#)L[Z>E*=HUE7:
P".+-*8$LA+J=,@LIK"J*[66UUQ\%;09:5LAON.[B3J'YB#9U2FZ)UC%L($E;X T6
PK:#@C2L70H>^+J_+%JN-51=\\2^6MM\#NC] P$34T&>(^/$Y/%U !7FHZIMKAC<(
PEN==S4*\478#>-2.& &+0;''L*I^]'$8T6GF036BP!#O61G!-N[--@UJX,J_  8B
P7"R5CA-@5Y\,_(//-*_TC5]0)"L;(3DOZ@3(M?W'.ON%S$8&%,I?=8^#:<U^BPZY
P[8$@@OI= J_12=58%A^^ J% FY:<#J!J%Y5;[43&/SW:!8_)5^*C,4NZI^\WO)C"
PAIY:SD327L6WL5!6F>X,8[9=IZ[BJ47?^H&M\TE=A!&&SCEOI<S*3SEZ3N6'<8$N
P?L,)Z+W7YY^E$813;_K=RQ](LH_Y%O[S+%J=O=-.XG[],IFUH$DB)=*[=(T 8,WI
PM6"_$]G*IW-1H5L*,4+;9_?_]$.<K]-RZ9[UKHVNGZ!M0O8IV3H&@O6=<J+[5LX6
P(;NZ-TH#B$1JB#B*RN$(V'25U_YI5,'Z0 YO-"7-*9;K.+[& >UY<5?SWQOTXF72
PIP,7P4$L3W< 6.*DTB*83EA(O</:!T8_]8E:>Z<3)@H3R>8O[1'L\<0)'7NP>%'D
P;][?;M4%%8_/3GG.6]&L90]\?! [[>;M'749?W!2U:/:K>T\F[YN*Q](J'H=IV?M
P&L#T7Y;G[ARO&[5;>30]Q$WGZ(UE*0L5RD&!+1EJ3I3W9G2R_GW[.#1?Y&&5?0R_
PG"ITT\_?V#2D625K,EDU(I3?FT\1>,>W"#VYT7+C<7@_JR"4]7TNYA*J+B9 DYZ=
P+7N<&KK03"@Z(XNT%:!=YK=XME/1UW1G9 #)2=M8)TAK%]W6%H]%\(#]"QH-()&Y
PZET?#CR]3=D0]K*I%&J;5&*563FR$70-Z'<HU0+@EZ,_3N5=&T"%C\)F/3,/]@AW
P,";#8?%^C]HDNWAT_P)XH;VH,:?)TO^BOBK-3C:<0I%(3S9E7BT[JRF7>4&<)V3;
P\6S*@56DY<3/'B9G=S>/[_?\H\W&Z[LBQ/2RQ*U[+,H(^!5#=77.75WSQM(F;$OV
P^$;YJ;(#Q&L14ZI*$M0>SYIF:>Y:74*;RAD1M3]0-CMUA ZKW2JDC1I,_3:61$_/
P6_.2ZD0$1TPDOGJM!$*3F#VX;DHR5[B =KXCVG18E-Q>7+.O;KY/O)9:?3@>H5"T
PL]H I/[]5S5.P^8EM#ERN7PR[7GDY#:DKJS,IIM*"C'DZN_-&$%TO%%ZTV[_NC K
P*F3(6%"CP]K>58X;=7.&NJB][SF:0^(TZPQ5)(QS&I,$T5)Y*D:_MQPW0S,"DCQ?
P286/9!'V1"?(V.4LWT4>K(#G-!><[Y*:/=?9)?Q/_5V\(*HS]UC:@55Z4PU%*CW?
PNBT"1)$0+QO=I2>=[&?%4-S>UX,:I*)Q;?)(!&<19FB-NFM5FE$RU6N_+6WB\U< 
P5X1U@?_N2!HPTF25FG''>4J6/8;8GA 2Y<X>P\&UDG[ S*UMR<,HQ$=I^;(P)DD>
P>D-,HU<D*;_HQ/R*O'5 4UOY',YO&,N GN_:, 0[J2#N'/9S8+<4OEN-'K%?O'6;
PIJLC,T)@ R\B:U:7*PNO(.[GE'N*L%"^,7Z7T,C+;C^PYU1T^'!2EM'#TG.]Q5/]
P=O.Y^ ]@^KBS: 37BG@N?X=O?V"/>09H(1@C(\Z?(BX@?F=$M3G''=.!C7U0Z>Q-
P%G>KE":+G:.N3 A]Q5*PCS)ZJ%)3R]MLA,:;:]:RSNQ])?W2R)'=&@=]+10?:CZ$
P90MW],/J7,"?X1'CWT2LA\'J:I%5<<\KD2B0-&+QW%-);F HX+\_&F#S@2MZXW'&
P+5X1+8-\W][%).967,J.YY $W'V+EA[CA6>V*Y1.\%G:*>HGZ,;WG064,3S#ND2P
P7+N.K/Y7 5QZ,NK-%'BG6=^&6V+L.6VPF$TO'04+%,B/S/6JMV/7Z?X;; [/](^&
PXCA/++-)7EN3:8/L1])CLSM?"-:.]#Q;VT;OS%.E5 3P1I)VQ1C&GK'(N6)EF/BY
P26<4% )2UT0_@%NF5&2N'C!^W\M#;JK+%F#ZX"G*%-NMTIX.9#,C@;)8?N'MI%+1
PF:+OV#K*5AT"Q27T!!!EXP!>9F66>F]7P!FA6.//B<]NSWN41MK+;ZCA%RAZH;3\
P_^1P=,<81YT3>!*J-U:T5OO&[!O00'\]; -]:G+A6._E#D6>,4Z"-.R <-)_IA1I
P8O^^R"B<2#$8DZFMTB^&Q>W*'0Y0WUM"6SI;H]NOT&K7B;U\X-7Y-(FB2Z@L'6;I
PK5@A(L?$N*6H[C+#2Z9(Z@D[$G>^S<O3Y7,B//U*2RT1".)+1*(SQ/!AWE15"T>R
P9@SI8EU:P6$U#4TA@J%,-SZ;*?)N)D4X\?T9G:R-7;B(89X*[^C&F9OZIQ)N7#/V
PXT'M/U*VX08(2[1C@=58^:B6E8LPK9\H-Z-26*R3HRE0_V@DU59BZHA\2->438G$
PAREP,?0M,H 7(V .]CG]MVJ^>,E:\PO93,HP\6R7RT!(+?NKE:)YKDBWW')8MB/I
P.T<!=8BQL=^*+YN)QHC@)BQO2XB6'=X!D^X66 F8@'6(&Y%=HD-2>IJGJCTIE6@J
P@[079?;8NCC%-SZ/Y"23?(P?P/AN.G*W'%(=Q!>E^>8(7"T.18Z;NHV)H$,$OG2+
P%]#2HAIJQ4CDL%*=!."#U3SN#J&%_*.)&6W)O;[D%/1C' ;>GX=:V;P7.M_;.!VB
P/1J/,22-V4J NJ&I3\^OH BRC+](:Z#&ISJ90P/8@KDGLJ4VJUQ;"'KN!:<3N3QJ
P$7]Q1%G#?F=BA$E*2A>X<M[KCNL79U<RRRGA7I^-;<>\<*WM\;'8&BH,YXSG:[SO
POQ1P&:9H.\GT#BZ5QB@LPF0N6]U X>].A4C@@S/+ZDZV:@@'KGD9E,(W'N,F,_W'
PPW_E4T0Y-"&4Z7R*S#?,_ACLG(*60D<]"SPNG##</-",^#/+B^'QSHX&CRZY9,<$
PN44Y.S*Y="N/WN"(8(->CX\ K)?3]N3R8552:@S' EQ,-J."V:!N)PG$RCPM>R;\
P-\D:SSG7U#48=N6933D\9^&/"<W;FW3_5](S"40@KJ8P>R@9^;$%+3DUN?\56*[3
PN,/T+2=;5['D=I"^$7?UE(3;9(B1RFRK-H:E-M%P^+Q"7!$'.6-7CWG;W!1[3R2T
PYN %ML =>3T5W$DF0VN4C?/IPM3V&1@0@+L3V8)NX^Y_\D3_/.@ETZ_ZX_O&!LE<
P2C:XOBI>,&FL[^M+0#$(N%=1=)H5FWU <4A06@-2U6&BX"3\QS;+ZUW$&E;X:F&R
P'J1-'06-% 1#P\-=!$?,36CN3U(\GTL8)0W=*-PDYYIU*E>?0C9$S"+A:5/,FJ$E
PIR"!V4WMAPR()W<:_ ^4Q(X/-*!*W+!0B*O?+G).871AG_2O!VO'N#XD%*=!%H;R
P9PQ7F]">0Y2D@M&./4LFDH!-$4DD. +% +W3A.#0(Y1F++O?/]?Y>'^G+R1XB8]-
P@L</<@9%)PE/$35'7[P,^F(8[1BN29>,<S%@9>6GQL1Y ?*7V/0+.MX/3M$]2F.5
P$Q%74@A"V0^50)?S1B3YUB6[RC]Q^I]>H($*4G6F:TM8PFU1#%/#5IY*P9X4()'4
P4ZQF-L#Q:BL\OBT=9A+0CCOL+\9\F$AY\++*H :5U;=7S(N'9'9>N$9/R"L_DJ9B
PL&&1#?7_%P5*I^Y[O?O2UR[EXHAH1E[VK(2L\MX=$A!&1WGG "AU._$[@@K'2RWY
PG=W563"=8#SRG_8R1GCED0SPT'P LB<?N'-AO//C]S469+OKV4MFW^H3(]](F?#V
P,C5\^$L1*62#<\?"5@^NOX&;49PKX?R48?$7ID:Z"HDP=O1;OW[RDJ8Y)6C'4G:!
PS0-D#9&1^@RFSX8&!<4O1Y1+V[\4_0]+_.C!QO.[''(HUB_3<3@S8,O?]12=;,4U
PP]0L2'FO"+6%"<366H"P>YQO]R(UIC;Y%W(C9"J]91Z.'WQI!;C(^%: PKS (T$1
PP*>I8.N@XV$0D_&)ZHC"4$T'T4Z>7!0=7"B?/)FT?G5*"%-TB6BAZ-,B$WOIN_H!
PN%@Q0SO<X.@-EY3DJI%(% +W3'J:=VGQT=VA#A"A7Y+KYQ(?EO3O/ZWUP;P2=+>?
P%<=Y M7 .UQQ#H[71GQX$)3A+QW9\8! R)$=2X6X2HUO*F"?]BD8+Z\DWS$.XLA?
P(EHAII_]M]G$M_LW1#BM@I2];%;%K /#J5Z9R##T8815Y2K;8!5N$,=**'=3!Z7@
P@_P!<#$!9TB6/O3O_-QIE\W)ND +GUTMB08K^OT0W1/8I=5X"]O6"JV4S> "J#67
PK N3PRI_]T</P)NPJ@0TF,U7ZG,>G,555W#N4BHX0(EY0A7+U/F '_>A_96:1LO2
PJ!\&&5-^'??G^.B<P0/QNR$IY$;U60RW0A5HK.I,4X!#,\LTT L;M%40I[X''5 G
P.'@,BZSV+(.4E48+'<327E&6\NREB_&2\$#FJL(O5=:RJA+>PD%!U#@)=CX%:O;#
P?=:T_R<0HXG7/ :J0B0;0['+')6AJ ['Z7 7984?K>BN') 01B+>$,\:@_IH\L[Z
P 8!V@Y U!1@YTVS)(,Q0I;>X%,'!PL'+LC]=;O/:DT<F4]/C\-8[KL?%A\S4[)S\
PQ!R6.AZ(]WC$*FQP]Y97SNI*]R)G>+P/*5O0S"H5OP&I#%'_JISD+>4?.O_78(!+
P?8P#O7A_E$I9DK"&VLT.>?K2R:0/4\,U)':60R2+ISEEM*3_K#8C.)FPL$&'S,1K
PX(FKB>?&GBE*+O,@B/DU)UZ7*B'(I0&F>-#+779^T<"S0,E$Z<GJY*_-#WO'@-%D
PYW-]SMPV6J;\9U_65XDM-LFQ]2D:S#:6F[2F?<JP>HAL/H<_CK-5.1ZLLE?'JR55
PGH%QN]P^H U+N9F,*]C8NOV%6+_\##>E]?@ ;Q)93*EL#MWS)M(L@X![(_D!5Z/W
P3:.C.7_7P7R"V\:_CN&-\*[LNA(!YG?K!TC$8D%/3$40@:=L_,F9I,C)%3>T'; .
P3-BOGA90V85B>P!*0H"C1IEV!*G,"=6^*G>\FIW_J1731D]HO\G$9\U8"1.W9_"+
PO*6Y)XLXRM)F15!/Q6+,)-(7V.8MD_T!BJXO'E^JA0L)]-\."FOV(7O+[CP\>68)
P)EOJ\-51*O[>3^FOYZ-F5SE 9>Y#ZFP-1GAV<.G5ARC+=U$;WP;<BCZ((^XI.8E\
P/;YG'MP=?PG;H79[C8K1H4*J=VFBK"#);?DZ$FA$:B-5/T*A003]) TUJEEBVZ;3
P6/^Y 7.504I"15#RK5MR;DD]P41C,/$M+"M@308*?V[TW^0\C'4M0,%X#Z&KI/&#
PZ;&;#3TA"?QCBU>^ #JC+F=V$[1*^O9^Q?UW(+ 9L.% G\,6(B7_E'P19 4S[P 3
P,YG=CF/5BK2)4.RC2AH68)]<WJ=T$$!^4QUOR=)>P@;JF2 7";M.OC+XM*K=Y" Q
P2?V._]P@DD50*+(T6^)FDO#6*?HW-=*'I3QTFELZ@^GTO$,*8H!2BD[ W;%GAJF_
PU7L<S6Q1K[O&)<\<OD7<P5 EQ9'"U&4%J7*"26$W48827NFH;<*,FN'?JD\&=V4P
PK<UCK75LNF.-LQK-@&ACZGIK@N[G!-9VK)VY4P6L"M6\-LUNF?S)R!=3]!_V)#G 
PC78&[C22\7A&1C2Z9#>U(U?"N BO/3+Y^=19+]98 GR#[S'71.-:X9@K[_GUB<A^
PJW/@R28"MYIW,..<KL?+FD'WZN1!+X$-_KTH\/FP'&/9S% 1IHP%=>*=I+QSI\Z4
P3,5@8O\N&:++_'O["V(%8Z5<;#2.9I<XBXBVM'#B/27&^16RDS\=GV=:Q&D,ITCX
PX=S;=!?/22K^<C18L(^;E6(_XS=W ,CX I+1IT^/QH1\8UZKUW=U3]3GL#A"ER2(
PI7"I [VX3J.1GWOW<=VVA_P!YDT IA%NURE,W_&8@T9@5/VZ](&X(%M]Y=[?OS3C
P2XTAA[KKHH%%C!>EV23Z>5AL.?>)RJ2]&8:(GO.IH0?HW?AF/XEOF8*G5-";%+9/
PZZZ7H/\X)'!!L^=XP?T$:*HTS4/)?@2$"9NL&,0Q-)$^1^J"?41-F!V+UL8?W<XM
PZ[/<9?[0"IYF9<#;:\U^VD#/D5E>&LO9($L%T?ARM^"7;$37$2B(8T8RD&&*H%X5
P=4ZOYX.5<8<: [(%DWD,N,7Z"HO[?>[O6*IY\PY T)D-W RAW/;A_*0UCYPE@/\1
PV\ 9]G/(!SR696=R<O&&LIWW!;&L+)\.@PH8JC3E7\>'E',+2WB1?<W*GBE>)WIH
PG="Y=)3%3*W?V$D"*M.I@K.5^\2,4/T(;]-[-GF+-B-+A@'JXQZ[VASY-E(A:++L
P^ML==+N,H/;'KV(8P8-7-5^-4T;5DQ+$L=[%((+_-?M,H%V69W.*_P_J,"_!0)-U
P\^??@QMN DX!GVHZPM;-9"1_!MO-FV,*Q(1074=[*:_XKAKK/410*S<HY2LKT=9-
P51G%CA!O(0C./8_2II+;0 DN'607B/ QGXO;XG[:OB@Z8F+)Y  ,VE[+SB<]JUTX
P]DNRY,X+5FEEWA8@'_ .EL>BQS6!DZ2M2NK3F,+P^E24I]-+FLMO.2:NC]$MWTCF
P#>LP-B7M)(J"-,VAA*&NH5:3DEA + [LAANJSJ-Q!)T4.+8_OX01B[EE1K^)A-:,
PGP^1"/NFH^UV*5/05:0S O[VL%O%W?)9M9V$JIIW0'@+=H3-X#P7T2UT%+MZC_O3
P5_GJ,G(""V(VKUXS1V.R%07A[G8X7&B%,Q[)2D2JP= 7T'OV(D0WNYQ$AP(41VPX
PK7P;IECB28^#:D1[KRQQ#=G(:2</DI WX&:RU]? JT 6(5"@^KW'QZ?Z(-=^5@5=
P!W?1[GL/RU=LTM"G&?P5*VH%5P_9W4>)/V66D"@D>M4NC4"1$D0\G5]C?NZETX*O
P[H"'1Z6)>B5(_Q737?WV'%-'@F^Z@XH0'1.F('A;2G)UFKH-PG O\TVHYFU<$ AS
PS"[?_>N\#.K,E2B=86>1*$T3=UONT&;GCU4GS9S"21KK7'!88G  K2Y] T::+EL]
PI2QYPO!9S9L-."=,M@9F*:][+GBMC9'S"['\9>M$$-A_1A[<K6@"V9_=1K#'&93.
PJ*>/0X%.ZU#'P^E(SB?-NL\'D;!D.CXBB=E+R(%[?)A>Q58 W*_K%5E?3"9I=4M,
P71$*THBZFV&U >+RR63F"DKC8./:DL%I#/_GC-ZAOK-D"[A=!;F]IA"@OI_5*J;^
P01(68,D!B1>#&\I'2B@)5GCSX$\H;CLMWS+8".%!,*+6D<J]+FYX//5+5_E*@%E^
P:6063X]K!BICP!EAU$\6C@"".0A Z;IPJYZ9#<U[$^NA(EB)\#7O(>T/ZH?[+)@#
P(GC<5S3<3!(R+UY1W1E/=)S^.R'M;=.W%"8<[Z1IOD&\XO",BVR6W1) 323JX!QH
P 7DF&.+^J6KQ3^655XFR)+!>EF:+#&JT"N1CB#[HE?JLUCC[JF4.TLW9]J26FYMU
P6D8H"UBHPLI+2X+9JHJF54,(,W,VC )6B78BQCFM,UC]122KE"C*BMR9QT(*TG-(
P_Z6U>F0ZE8(V/F,/_5S5/G1D7[6+I7!%S\W!0%%?9O8L=/G$5\ NO4(1*>I7,PEQ
P#I)>=6T[AN!YN8R8K2;9['X=$UUBO OXH"AZ[+*\QFF4, EA>\J(YY]O&7DX9Y&)
P!W'9N(($[NB;2>D]#XB!46T44D?7_@:\V+UA9K*JXW]IX]/QJ#HFY)#<$+GOPD&C
P+- W9M).P/FTL,X1T4K;;(QV\0T>3*=D^\UL3-?X&R0F#T#WX]"77.Z&'JRTDBJ>
P9FZ8(A2OG 8L?MU?. *I;&3>&FH#3T#4]#HO,(6X]-,./DE70]=WM<F@WCD&^'_.
P&T3ES*2D,2& 16U+G.N64 N?]8I?;BUO/MA*=5Y7-5#<*,OSMC)'8?K?BT[U+S"T
P<1REIRDSWEG%4V/T)*WSCVJ(Y;9E>$HID66C)TC+<2EXW=AI1<@8O(=M/_=T;D0H
P8>=T14:;(47E]J'G_<=3?SMHYA@GKJ7G'@?H\EIEU-%GTM-OP)*\;JK=4P3F1+6%
PJ*8S547!;VN(OM$\LL6BWE#+H@*U&#T9?BPB;O+*4=+R13763_A@D>%YLG4TQW#K
P<0'WF!:7Q]:!UA"V[0JIVGDI9:^*8YTQ5>;B+,D*2/,#,NFM\*M4"+#7(EQW:^$1
PL."=YW10I4I<1DI1Z5R$2IA<>,42N[OL9O$L%*9UWUH[NHRZ9Z2L83&!D7YD<P"0
P R$ZFZOPCJ65I8&89&*UZ]-F'6IZ]#1KS1Y#5 GCVEEO"E2E<.R><7J^MTE:L#+/
P/BC[!V.Q\Z7=WTN52Y-_0AP*8D $]I*IOCL&0+GH6#D/QO@U8AT,]++M'(EM#=>1
P>+9^_9X:PXW'-:E[^,4?>IO!D <@7'SB:0),$3?4PKX#]U9(BPH/01#]A[G@:Q@8
PE^0= *R@-9/=A#VO.SH-ZJN<CYPG^?X[75?$0]QD'3_^M;0Y,"4TE&ST'X %,FY@
PH:M)6*R&82=;HJ]Y.-SD9+C#[:LY2*@G"?(T633G Q:"^F'J<85QG:M&B8X*]^Q9
PT:KEW*U0P_VNS0[E"Z@$) '.Y0(0O'S[@\@78!2&3E(8T@9O]60=KMHH5(YJHZ?>
P6OZ_Q,,A0RX2*]M=('D%BZ^[LA_=' 2G&+7XQIW!W)DSQ)-<(#=CL&_O8IGLJQ]@
PK6N?4P9%,Y9+MD7*8.CC(D!9,]>5QO:OM.JY7P X,SH[Z+?59EFUHFQ'COOCS(H.
PG,1G=E1FCRL[4 CNZ+AH!_#><&7:_T"M$"!,@Y<2U^9&:,($>'.&> \C*-G?;]-3
P&^.CGK 3VP.51&:/194N1L^VW=0J";@?E3G(?]X+79PO.9U_.=6T\]:BA)[DH0H-
P5%/3RS=(=8 FXXQBFZE@F5"/SQ' L,!_"3_RC4W1:D\B5^":!8\S_\.4#6'L,'TQ
P3B/ZE3D!3?-%6T; [5/$K7]B^),T0S[()]@^,HQ+5=^]*E4XUZ QJ@0BLPXQ.7:<
P4$F EXUB2?8O)E$$L_'=U0#9Q4&W\$**V)SJP@Y,D]M*<Y<%>^]XKCL6-TH!']$O
P:7<L<JUJO7_>:+Y:VJI$X#7:52\9N@/7)P=2BKJ?LE.G3D>(40*H]A8DA%*FHY_B
P\LJ__:/)HI0O@ ;XY-ZOC[R*12P 1&:^F91P>X29L""[$TG'SLY0@7O[MFKW?JQ)
P!#"V3L/BSI*_362F9.G*HH_-Z86:$O]Y174QET94&ET-;KBQ2]?[FK6GF^1.QMTY
PUW)\VCA[!M(5',183D97^)AH2:PFDW/3/##?/W)I%K#%PI\VBMD4^I[ JZVBA@S*
PEGU@$ X#ISQ*QMUA26R<>V286RTM",FDT!FK!W_.IPON(='BGI5/1$LVF PU1$*Q
PX)A9!C213FRRN '_ZX<D:[I*JIRA4 LM@ (%+2@5I%[C_"B>=( D4_D/^Q?P23;P
PXDWCE0=0[,0_W:#N!R]^)]WINO>@:L7E/4]N'$3K%,^RL7<,9L+ -/?^>(Z,J=&_
P2":H7]?^EC=D5N*J& ^Z^Y18KXQ*9"<57HO9J,0(VP\LUME,$$&L4OXNE"!N4 Z=
PZ!$P%34;159S;2%UZJ0R_1KI1]FN!_;S(2?C&3NM-_\P(ZYJZR/&]?L70ZXYH^S<
PRD3IKX?\R4V<)P@JF2GM9OXO19F#!5RAH(JLT!R?-@I@53J-.V0)\"C7@45;@XYG
PY"#:.]BTSO#)+\FK2;NCYUI:=@-WN$D]]OP_3E91M:%H [*Z&(*)X*;?.W$])T.?
P&%M$;,,Y>)]YC?X+90 NXXZ:(B Z.?8S,WGFVK=RJXMB1HOW5FYL^NAKD&<XN07%
PV/ <D,;^5C[M71_3Q=_3+\(J:KT,XS$4HA+V H\NI-4702W_PED)X<>ES1) @C7Y
PYHD8G<WR'5\^C116OP^REPGUBY=*)LD!>+&88O%AQU:ZG'C,FU8S,C)STM:%BD.F
PZ-P[Y<.D^N2YIX-ADG:(#$/E@"N'B)/Q*K3P2K,?T+D2!_Q=%^ T9(]2O[;"%W_=
PQ@3D:5?C&VS;"NAVS#UX/00ZA<A \. 6?8-@=H\#:,]8%[H,&$><V:6C+9X2.:-X
PMZHA$)"-7]S.\Z+9\?*E27!B0J*%1BK:I,A$,FS2WF<^0,6<()X'8E3C2@VW3MUF
P9%M]!'J$WRU+(-RA,1KH+<;5$0U2%W;1WURQ[Q;UJ/DS2^S*@#G84]O7K&=/_1H:
P(I)$=>,V0&9OK\Y+R7[[KFM]<S0P3+0>W+&ON3.88]_G62P#K: V@9Z*6H8.J6R\
PMO+SE9J07_+0;KIDOMM4,B >[*KN:D::^C!H\4]  4GY AN@=%K"XA(+ "UV6E>:
P?UG[/8KIR6L>#(<8!"3R7TY_^\3 M7D4"0>*)(NW4\^X"FR-E\]FZA36M7J3XM[$
P%"]U?B3C?;L:7]"<MD*M';!YH^_9,I$SG='_MAY(>+B6.%6#NF6 0@.33WE(3AN:
PKTNL)&&MZ)=,@D/#5JJT<)O[&/JFMXC#>AWOX[E9VJ\OKOPE/$@7U@MJ4-94TJ+.
P]OI2S;H:W*!MGBJ 5 !^0?(BA7MXB36X9E#R4:^TT]436$M<.H'&>;#'M8L/U+$K
PVN]PPQ2M8<Z4H<6DQ2)ZG]C-YI)!()20$E(4"D\4NHQ=VXP*@< TT\!M!WJZ"3A1
P9*W./+:H<.,7 _AP;LPQ!%7;JX[:I<K0NIJIHX-%43(]T1%I:*'?+T.?O]YKJ#&L
P]!P!38Q;29E#L:MT%EX?M]"$@1\QO0T43LV/K)T_<<Z(S%ELRY\X-3]VV/(#+R3<
PSF$1].'%)AG=H$?B+T*>HW*[%ECV!4D[*/4=N0W3AC"88PQM$A9Q]_R?_.KF_\E@
P!7]S/?J>V8SB%VD&H<H7O_'<D4\J#!?O&@J65L1Z[O46$FY>H0S PTVOCQT[?^@H
P;PV@:HMW__3RL\J?_T*^? )@<OH:N9<V'Q 5$P;DSARW%)$7"-OT&?&D21,(Q<FF
P)4 ]SG**Z]J]Z[RJKL4%#%L4X#N\D-@H>Z=Z2"2PS\401"AKO[+TQ^6G;_#TH0?U
PZ)UR@G9\5W=$,FM\U+9ZP?:B6,,MY#X/SG0\(^QI\_VX-XH]FF-8Y+M[61QQ$CJ?
PIJYH4-Q[2QU$037P2-\MEQW!#Y6FE(%/\A78G'DEO"4@6<W: 6=:KSD:I5KG=S&7
P, 4/+>C?$2E(GQF2!ZZO<,(8QW0;!\LJ-T$8IZ^>>;_:Q-Z:N$> (M%G>9.EGVSR
P*YD5R!^_P'(.Y"2TD1&A )6::YUK5W4'O9/N&3@BIS!X!6@LVEW9]YH!(P4; E"E
P*EOW,M).R=D-U(C]MSRBE:8?>S;$O*[3!FA9%92S $N!LA0Q&GVU?LAQU^8D\/EB
P-"- >+/ [AI)-&<U7=7?/($5!JL<-3N@6WX?:Y/ QX3TE/)^A3LS_</ ,*@\KE F
PR$J#4.G1D#T\NK(5!&F#P@#-GA OT>?D;';6I-Z80/&L#FE]0TS\KV"_>@>K,NG9
PE FYXL=FZ*K^CIT/LV+SE4MO&_)<]Q'Q!_1!Y9(IFI#"$]/(V=&IBMKPB&A;GT=V
P8+N)>=\.Q[<&-.X_RTVLS&10;K;7!!USWD_,P55.L/7T&WT[^&@VD_B?OB'7OI6.
PZ'B"SG5&NW&XW[9V/DU(JRE: V>%&*6 CM^@'_8,ZNN(:^=FIM9N,K4P$:JI#D7L
PUO!@PBUN@&M+6XT_4%;?N[S5Y?@1^[X8RNPG!!#7?:(*4VK#>L#<60WHMS4V%Y[N
PRJR:E7K=-.=HT'0MO!@/TZN7QQM6:,HH8XF:W"O^G9II3" LA"VC#1:W.%CJ<B\(
P%;ZMYW1/_\9%H#TTFZ7HQ:7+IN2$T.,V4: O%M4PL&A(,O7MVJ5Y]G*M+/M!).#E
P5P3<UN[4ORKN\2]#4I<#;F21WJ<8FV]+P16 8]HW52#KP<Q9R.[[]SIHQ"AB$;;L
PA6Q4G=)1)X-:?G8K]"L!K(58WG90DN[T![7X$D0C>%$4\DYPAM\VP3I>,+[)L:/>
POY![<,@<;-D,$.WOEV:AZ+J=.6'33-VYCIN3UDQ8,ZK*!FW?(1;5%=Z(AM;;. TV
PU=A]F]T%6@/Q<<?Q*OMP_H4EGX 0IQ!ZD#%!S2Y1]9X_V60^<.E6%0"K%Y+&#].%
P@+E/7 \<@F$2>[SD@*C"01^7GT,U%V%TM%)+K1V7PKF=5UKB4-/$!EN"I3&%:"Y)
P3$6'FVI0K]GMP<P@CXQ!/[U2O6;, X&#7MA[D[,ALX!9W2>,5S4@=L;21^!M+IF.
PC5OA*4:?N%N<FO/BLX0;[R6=J]6@L;[]P(!5<ARI#[)%HYP8[9*OQNU<A3:72?0&
P+5Y(7"G]RMH-:^ZVU;Y&X/":LTA%JX_]%;H6:'S,BV$)UC46X=)(NJ'&8:%TEIVH
P106M!?8U7TII8-2T),TY'"S@ N%MW66A\^Q@WME1\M0ZGT#S_Y'"[BGN'F\G%O,7
P+63: 7:./0JXG,?]O4O%2YV6H<0WFKVO!QCY<Z;T)[P>&&*G+'%&/=R2Q/,\^1I*
P 6Z.2$],869H C ]"26E$W6DU&,@P2 !-XO*WN,^LTPHVYATP6WAL[TJ;S;#@G_G
P71CQ;KC+T+$OUS=B5(8#AI=LT]Z V[T)+X^4TF_PRM3E\B]NVGR3)3F-J5'X-)*L
P[J!+D"5\F:5M8]TC2#N8\_'19PY*[L;,5H@_O_5R3%M:J?G IM)3:;%8.)5%<PYX
P"M@$ZRS<!!3*_)6,6+Q*7WAM4RR*H>YZJ,N)-,DO]BZ):K_ABZ7GY92-TTQ1%:1A
P:+R6=8_!5J7Y_JVE8%[FI@_PHS4>_0YW^V!8'2DRC<M$D.9>.;(?(APFT:/U%,.,
PU?$FO) ]'<LT(&IX*D6CAF3=>%(L1C,;S+ZZ@AL6 ^TZEY0/K2*^58D),Z^WW#^#
P< \F,K!>QN(LZT1281%_E'[2&9D8_'/F#JV$[ZUKC7G_%$7J5.*/Q#I+\6SQ(("I
P;Q47/D@94WU/"%W@L#IXD9_S2HBM:^1X:1O [.L+TN?P6VNCCA%C*XX1-V+*9S<?
PH*$]=BB3^.R'D]+%Y"ZP.4]9V.9$>1QZ0\KNSO!]63#$QAM>E0)3$;NU-=';7H5]
PQM6^D*!4A2NLH_L"Z=IG"5P3'\CAED4#U5*Y9I-FTJ(II1J#<^D[H"J9.CF:29%W
P&0V=Z/=VF8PZ?D5=5RP=_9,O/7[)U;C'+;S(Z[)_3H&8G5J;3QMT=^Y-&DVKFX1#
P*NBH*/%>_(;&R;#JRA?RS>34,_)RM<OY-3CA!O ^_I=3E2:*FHCZ>/X>*V'UFSQS
PF8P*6D_<>O B;9J&J,^*U(A*#6X.H%.T^)H1A:72 ^5 1D,5AA? /K:3%UUQ+ UE
PBK_]EYN&L?)U%$AIRLI"M91IC;8\B@U4"M,^J)U87ZAEGL[=.C(S$9)RK TAA]@M
PH>-TX7?;)R:BL!HCI)2.F--NEC_C7T@/>$=CPLEL!XT4RZB.^$LT&.\YD"YIW_=B
P:%;[$/H)90,;CLIWPJO$2WH5-V$EJ0?&7(#%9%@ZG+)W]*)0E?V'(Y.136G;TQ"%
PZXOW3VJ@#*'2@\P7!KU4HIV?I?M$E%@  '@<+HG-RROUSQET,T-JS5/I\J;(H@J?
PZ7P\52'LRY2\%_<4DI??Q3+=V\G/B+8R"@E(J3V+1ATC(]IVA!O]'N>QJBW"&,QW
P6T@6%E$@7*6%4G05MMO49I]S"Z0$9B" *"YC#__K)D2&6X%QY12*)N1/A\L_W0QR
P!]V*U53,5\V_JE:E3'F6 )!^0!/-*@:9>MAIB/SPBL9/@%WP&&,TOTQQD+$;PP'Q
PPNG/H7FJ5TVC*V;4#_VFG+6A8O&2 ^CV>YH=D"+")@0/3?KI/19U"/'5N.9N(1=9
P]$%_^T#KOQJ:#_;<M?1^$"_T[C2I'R^4DN_&*O*397"J#.&5QJP->PA+!9OT$I$Y
P(M9U6./!<E<D-.9&RVZP+4OEA\C+-DCV#PL<H>HG'ASI.H4\$U%'IM FTZZ><LY0
P*(@!7=O)UEW&6\*7SDQLY)8"ZK%VKO.V<1''L]_M0TU\WK5WJT.9^3>[:>->@QXJ
PTL_W58'^W2M]R&/]BYG6*/ ZNEZ!:A:%^=RO*H@,96369OZ1\0<V^I_7[J%IJ,;/
PK)Q/R4CM;KY<!<]MH+17FJ8.]J &B:-#<#=? 5=%2MTG,7FHBQLK&-%&JA!LP E8
PG=K.7)%E(/(@!M6_G25#\T[K[,Q"8Z'.0<_K"@U*[3!*J# !?EZG<O;PQL,_2L6I
PH%OM0[^Q@1W9;:W:T>@O=@&Y?_,U$+(?GJ.(%:[7_82^_5_Q=RM8J?G&SFDL,+)X
P&/NK= +!G^MBPSO6E^8TT4MBE=^5BP1 !-DL3/ITVV5XG#Q<IL 3T.JD$:"5O6Z4
P*96*;G%/T:N',-$F>3'H6BMF1JTSC6@ID#RK#[2<&P02\8Y,.[\__&?,#5Q[6"?E
P!#MJ)(>FZ.9D#3/OL,0EQ(L'E9P&ON/ES)0PO3K9PDO3TQ#Y)@.JCUZ"1/FPP9)9
PA4 UW?N[)^,SQ1BDV>:I.#BJ!9&6-A?H@B*]G&@#OIAH?(T8Y.3.6H>1I0:6Z5B"
PWB6J-\XO\F^Y$MVD61%8+[9FE"HG>L#F$RK7AIJ"&U&]+]?V!RJIB](N7L-C6=??
P,19?=ITSO!#;&R^_QZ_H+(P#A'[HPQ]) 1W#'2AF(L_6O?X*=M3[9*0=MD]=5HWI
PO?N]EN&5!?M-<;B01;3/^T5@:DE@T_9 E<T8?F[0X^&D)Y$%*K(E$2'O 6D;+35J
PFX!_LR'YYIP;=5'[-'E8R)_?DJN'GX JBPUJGA"A+CA@!@/K&96S(OF]&<A,48H,
P<1=F(22SM=0!ACTLA:IH T!73YB=SE,YWR9%P5:03*+T/?;=TB"+#7[TTZ)+B.W6
PBC/0\QMYMH^K4#\%]Y+8%N3#'&]U7PWI)OE%4?P2.=Z3WI-['@\W[&YU]LCSJ>" 
PE1DB(97N$=1XVA%2'[\SVB+*3!7D;.CTAA7-5X8,NH3>*=*[".\\:@>"-SF(GEJ<
P3JZIR$ <K$RO'+G(5G,A80KF XZ;!="&9ZT5/D'3/>7^X</9D*1-HHH:3&7\,_\]
PIXO#" 8^8#NP<7FB9$S;#C\K4%9=9OANRF7C4&VM"'6_\ T$1O!(\L;:=L]S;I'M
PS]Y0M\Y^/S(Z4VA]][BZ=AD!&AE]11-_*^GQ!5T-*-@$=EN>6N"O\*X0KNK/?Y(X
P!)Q=T0E#UO%6BQ_ZB32)CU"0R_P\C#A4^G1D30%Z:9$%,!HO8H!)@#%1C*YR19<>
P /R;@_*)%[:K>@*/@&>'I2J;^L0R$, ,TEDV5A;MR6<'D+&'"YEA$G:7;PZ)">[0
PX$&U4C'9918K(^H8$(7]811^TPM:FS0/P:FLT3?;RY1-O_]O4]T0\J\2/QPSYS4'
P%8VNM%R(\><&E7IO_@D'#0D7'+XM!EL=H<"T)3@\[,@74*Y.M\(.;V02J1)R@?3%
PD1L+(9D!TV$$P6O5UU.']CW1VJ[5H?UT*6IP?MN% 5?Q"D0*W_-?^L] I#K D3WQ
PB@[!<-!6-$U#7^F^J01*QGYJ/O8X-:9X6YKS?)!2,<[3B<GH*!&&?6=69'$R,+_X
P .X.U+Z=S43%Q'W-OZPB*"FX,SMSH!D%-A2'9L'&JDFAJY!9-5"Q+RFYVV[3"X8!
P,^];!!/_NG==%!DPE4@31MNZ&K^)@DI]</5IT27R6.V[,L-)5D)@%;:-GO1I:5/&
P)H(2@<O'7$5#<:X>EF7^?(]WA27Y@?1<R C4GMA9_;A^7:!8M>)1C0_M^4 @"#+#
PAUY?^,X(8_37&>)"X3@#H>&A^,OBEHHDG\^GT5=]ON2YBCUYNC#'T GHBC3!ZF9\
PV*O,=R='#DH[:.WHO$>V_JD(TW28T1O%?<=0?\<Y69'(A=.)*4JMVKU2/+R)HLHG
P;$J&>43N9*8"BB\!A+LL0S.FGTI$8K6 .3)'&/J.P@Q@L($8*/RCB,P2+8Y!XP($
P:;WM"WBQ:)JO;"Q(E)21.4"K(C#I]_ 86T<\F_B5G3&U3$RW,JZ!",OC9I- N4!L
P%)R5#A(QX:PCB4B=V:%O-C%XRF_V=U60)RYGA96\!E+M6@;9=(L(->+$MG75RDV;
PQ3S?_QZ97^;<[0/3I)5K0D\/6N*'Z9VDO,[\Y&5(,4UMXW0D0QO9\"EO4% #)LH:
P=0>R3U4$T0 YN%+?)Y2PGA@H($F!8+RVP3L8X$RL8^HWDU8._W)JB2-85R%6O%J2
P";$9K@83;Y(K>3HI)PK]I!JWY>U*;9HT,LKUR'=F)#H2#MC@.=)#%>1U3SEY<1B<
PD+CIU9&>C^&&R/54%,P_96T2<(75)^\47XJ%3"/>9O%5BX"=X40F(5YA''-+QU%V
PK/^R,I)JG'$_X;OC_Z!"$QVU#BD*FV;QT'N^.]?X)2*LE9_J:6/EW"3WJ)9A3M@)
PT]:Z4T8?,^9JVD 3>J[):]>M!#!B<I-\JT+;K@#,&2]LO?C*K\0[(:^E4A=9<GOJ
P;D0:HMQS.8>X?*R?%$VOZ J$IJXR )0]/% ^/OP6*KFI##26<U+AK^05O*J,E ?"
PPW)NOA' E\U"-9?XZDF3"$AS>X^5P*YKF?ZH&\\T2.MGF[%#GV.NN"FUGF:L!"3/
P_VG_L!Z/Q;^]J-YW""E/D^_,K<$[+E*\."D@>4(<^C60[0AY+MV I/R)*=!(Y+#@
P'LH9WL70[EC @OFUL=//?NT![B)]3%L<2=J1CQX:=NK'K\LA-YIW.B579#$-J%TF
P7N>(ZVK][IRHH-D>%3./3YRKUM=UKLZ$5")A9 ZW\1$.O@Y-)C4V0,[E<;J+XS2?
P=IJ\6]G5HZ=)FOF$2@PI1I'BN5>C]S3I#LR[X_-F_C]@G"^U'-V0X,/<'<.!D;K&
PS <HI:2T45[,AZ)F2+ICY)FWM\N44%%(NL("7JZE1()/?(/<"P'"8U@J%90C7B2U
PQ'$W0KF,^DJCR7-B6/CA<.W-DKV%LL[/I.(ML(/[DB6FTS8YL3NP!QO?G;/V*:+Y
PKB*+K&/'Z_X0BV]B+DA"!V+5:1)]M2+%?9%YCHW8.;6"!^^I1M6NXWU[2A^/@DA\
P>_!0I.@;,'<OZCBE0GR)AU&3M"W_R$0F/'@E-0J5*I(WRG375AY//EB E#AN\U+W
P^?EIR\*_O9?B<E:X%D>%\F$4_5>W&BM>USDLM8D(/X2^MKUL^*."8XFI!Z-Q&;I9
PM9<)+?NQ4^(7'(J23#GB,:CR)X!D;>2T&97)<<,Y20L>#"'(TKP^S"/6@B:Z/IGS
P-II0P1EN'7A=V-S.&%V7+[#L!D,>/=<+, '&PV5/Q<Z5)"@6:YWI9UR4U9(#SZ$U
PBL9_^<6RU$MT5W/-FQ]T?8<=&$YXH+]X+!<GP4G=YUG>&,EE#Q+/=)>U'[ _Z.0Y
PSXUG:PSE.579(3*7D2,EWGJ8#*_<CDO:YNN]F$Q=@+6"*S+U+<V,OL% P8P@>BB9
P@/*4$6NRVF/J1SUU3PNZQ@?C6?"-31H5W5P[W5>'949PI6^7^4BQ>/;1>'_7L=L]
P MXA143!/;L_ZW=^0<G::BF:)+-?[6X ).,Z,,MZ)>F)L7:9F8PJ'9=OU,!!2.\C
P_<5"Y*(<&EE$U_:QLWCC5A&HJ(9C.$S;CT%HR]<<$S_4$[8FZ5KV5 B;#5R%8\_?
PO&!A9L\,=:(^_(]?O=K)^2W?(Y6"N))3?TF]Z]ZP5>*Z_7+QZC7+-2Y8(DMGER(U
PDT! TW8"*R9 .'[9NH,=D1PA]&,"#[BKL7DY*6?HK?]NCTS4<=7A6):_MQD82.7+
P["AS6?3UV>##R=+[Z#ALBE6;KX8-2I+H=K$V2V40AV6C G];!S#,'>5I]/@PC 9(
P&<N1&?9U 4.6J^R@R>2XJSC%>]V H+7 +ZW8Y<S\9%&O"'S_NY.]I:1I8L[RGG'-
P?17!F7FZ1._3O=MC66%7MI"*)W3T MA#Z]&&)IB'W.5QONGZ>M-4<8Q(O%2G7U>?
PQ#QT[]35DFJ.!L$^0PB8-^]G,V;(-?1O?/$/=#65!,Y<;SQ%VAPX.$"5X=/!LF<C
P4'75N9O-N.KWEL-R+S!WB(/N="PY;M0S;LS&1)2+E$57+8>T@%";R :STG9S.6>Z
PJ(=;.9"0G280(:)PW)F)QRR 7H<^"@I9/%6%>UL=$9HU3?![W'+V>1"[43FZ=]\!
PE=RT_(:BH#2HTP1CY#\^VJJK4L:0_JYNL$E(>W_6J.D-\AP8VD@3G@*)87NW4)"F
PX,^XDFMN$-\0"\ 7N4"ISD]J]-!^V=-PG[$GM3O252,M$WXT/+H:VR=X.H"?'KRP
PE"OB,K1*UO!.1BHP[TW/&S0L7],P91@1Q 1S>9QMG/;MT"P,;9U@'$  J:&&S=#E
P-AC9'^Y66Z<=@6OO* T)7*"*!:Z8@2 F[-QS'*J0X@LA5++,2W^"%U_.,#ST?FO2
P?F(F?TP3Y.'=HMR4(Q23& ?NUYS5_S2I00GI%+07?I =\J0]'I4JOZ9.Q MM/%]X
PC4JNJ7\V@UBR17AY!]W?+SF-'K;';#NZL0%ZQ'OK(QI%8NE#^-&;DVM!PZ=P&5>%
PY1W\N>8P!8L2J)2<MD<5J>8J)&WK%T[ O:G08,+[UYAF5R6/;E^8EY_S&BC9:L$7
P>*JKN(%[=(MX! =-Y^EYL!(8(U)U^".JT,HT);+]45H1GE.PYD<6@J' (C>GVR:*
P6>4!BLC:3LS^)KXC(7M.!L1/:5&G.JKU4D5\Q",E-F2]M>W>2.4 37!^8[L]UAD7
P]08?J]"V_GE7](:5U /WI$1JUVNGDBP=L*XHDI'2'SKAPZ&:_N6GBUEK6*NXVI/I
P5"7GONSIZ\S9/$S]M4F9;6/.L=B$_%/=7;E?D[O=]FENU/0@>DXH]$O%OQ)-]])/
P3<$G"@O_ +5Q<R%MS3"55D ;^4$&_1OR :#^_*WWX+8SM1D;>2$P(FQ&D-9JLU1)
P3O)165R!B(6(Q@/_8C6.L^%Q"8#S@^I/]U;5DK<C2 V,_ZAE>"NEWL#F$OK#HS0O
P[I128/PX"60**!14$M_MW8&],<:6I]WU_3YG?6=Z-(2B&(]C"X0<0S,#G'J:Q_^4
P]<X6J'G]?P;?+\2OS/O-SR7@*VW_[0XH'S5/ZD^81".&+G4L--BH#C&9M/LK<2V"
P_$IJ?"_J36@M]6M!'Z:3:DQ.A"PJU]951_V$EWU.11<HBR<G0Z 04[9 <W&O 8YR
P\.VS=SZ@M+6VV8[9>HW P#F,2 !@[A32%'FOU3PQ5J<%;CVQ?@ECJB.;D%U2 31H
PC,94QRX;64_E:$&LUY 27CH-:O7+B8 /C!?:,$  G,YT$G98R=R=4!E#*TIXA!&[
P59KF[*Q\.?3-S@D;*E\ZZ$FBO):J5O79FHFB)SS#\E8+3=1ILOE*S.*KFT<=HB5/
P<,X8%UI-]/0@Q4A,,B[^?V&NJ<\3*\+&+ J'5C0B1<4X0G+YR9D7F"_<-B2^I&T>
PKVEWY1$UEO5D-M"^F:ND-'5Z&IC+ZE:&J2ME@/Q0ZUN&LC6"&'@:)@J,D;VE4,&/
P_&4TC57'Y!T@^Y_&X[^S'GV^;9[I',?&KY'@OL99R@< #73K)\A[C<=#N+1_OM_W
P_7_>3,U8 5"%Z ^E<PGO=]&&FS8)HU.[1V:\_G^5!D'8:3#UBI+]V#.5C\,K4@9[
P&3;1:G[Q\MKOTO7.!5^'A"<ED'<:/2G>9E$^Q[]#[V_TK%#4[ ;_>I#I^OJ<GE=M
PC"(5"C44ZP;5;3PKU/*%?1)4#R-D<\3ZT)S!1:#]K9[A\*Z@\DER;RBG<XFS/:G,
P,.T3EV1;#I73M-]@^'5$Y6.ZF64MZ6J+RW8L^\_ZODS+Z.O:+B6O8AM^Z+J'*&ZX
PA^*%C%R.4Q&"]9BBZH,MU,G7-0%VA:I.PY5[*H@%)9<:$X7A_V,CZLN%S_DO6/[!
P @K'7J4\9&R!.ZEMK!])+3ZR*WS-1 QJ9\KF]04O^*@EE/ X;/2A73$G2 )G4W>P
P6S \H2& B<N1"NJ#0K[ [/L#FG!1X@U4"58C[G0"8&3X10EH?DSDA948!(QP666!
P10DLKW^?Q<.A&CC)N$#]T]WG#D(D&STAG:([(H^7 <&AE" !%!Q"X\#UT?I0(Y.!
PEDF>P()@)[\C"YA<BX! "X%5/=AAM$_55>H^ORT>0WIV".?XM1WV_]*&TT<_I#_<
P>+.SE>R'?-=3X=<!^4\X>QZ9_FB#0J:E"" RB\'#@FQU:OQD,<%W(+YL^8+?)C=V
PK3X^5\L\ZLT Q4'K-[Z#1AT&!R4Q#B)*,ARU0U]FKQFLE]6%.22&9MKL[.TEMWVM
PN>MQ7G5VT-(Y% 2H>&:/9.7VZ9!:H"2B>9?Z@_-06[%QP 0V[TL._&JJ7!O)53:+
P,33)O 4@D_AQT5NF@=][_1[V]DC =!]E4GS;#M)2C=A3!81?\'7CTX("R$ 99>T(
PKU^,S,SRW4@"E <=TB%_*,#M= []X"#/CL@Q Q78K5788+8*1F-VP%]#AVGP#**+
P:Z=4-JF@(*\]O]PYS^'=21>A&\M4R?Z^W@="GPI@NAUVMPJ+QJ<6!GQE1X_?8LB 
P&W!4;THVI]=P=#[GND0.+F0_.M#9R>J?\XHFF-?G0C$NA$NI:9\R;[ / O5W=*=N
P]N[F7IF(%FY2?X)1@=Z'MV3@;2ZZ&]4X'*[*RU&$!]V'KJ9E"?"RP(:U%.6H;S.9
P8QO#QTJ:R?[+08 9\X+Z5A[V_BE]*67:ZS9@/67))SGM541&[]+.&H3B3V<S"&+'
PR6=F["7=61$PQ).B0/I8#%:HLK6+>ZA!L'\GOM7FF_*\+[6N%F[)0#W4+&  ?KPP
PQ?3M37L(W7\7B4O[51:/R]Q]K#L;HG:P?])@93+TA"ENQXB^%Q$T_2MGL&/N?"S+
P<5M[XIPC\KD?) 8A#;F:>]<&J!L0L36ADFK-I)^RN@(?YD\6S40J+Q4\7(ZYP>:(
P9D&$6KZ6#Q"1)FGT'#EV^Y1W<?:OGU\#72(76MVTRN!5==I"A(ZEL9TDXR'GW55.
PW9IP>[;KNQQ?@@"9\36?&EQ$HK9>CV+E]P*:#])15-=116KVHM'Z,]P:O7ZE*1\7
P91!/BPGA*S.S:%OC$"NG !_8_#/(!$#G:*+\/L^6!9O8^95^:7KD^=H&0D>2;*@-
P*R08)YC>-OEXU7/)9@\:=SGR_)P]=1;0CA?24!/>HBJY&B@>_+/KBWT_6NC4&7/'
P9/?;]SE[YZRL*4=+^ZJH#N 2NZR:1KI&9W GCSS-W9&9UPOQ$,+&9F:254^X;LR]
P673X.$_UYN%8@S;-8?T:T^EO_+FVBMCYFJI3UX4Z^BS+Z6X=_M10V9_V@ZIO4.?[
PX,R1-BXP6PX6_&8;<C%.R1T2 LIZ>MI"!C^/7D)P>V%HF_K!< [@<ZY],6;5X R]
PRJ\JH+^A1#T"F7WPP3A&?/CESF/30+\K'X)I;\@K&A)]SE(@C,* 4!#Q7*;'%]XV
P1H@I8C7A&D:&4\D9D;NMR0+&^7*HIH/]35"75&<*AHX9V^>>ZN(8^ WO<U;OUP&,
PTMC:>'N[EI"*!PP,"4S,)\.S]C;'F(8,42VA8E?+^*#*+N4"-"2LO0\8:JN7_%@K
P-.H!LD'YU1[&)[ )C@45@;B9 $$"M;<=2*E"R0_2)V$]#G;*,"N!+PN&)Q D"&_K
P6AU)&,U#:Z17MWN?+'"?GXY.N+3X0"'1Q-8ZQI?%8'HQQH4ZE_753>?VFIQ#W)V2
P;B+:8U7\9UM73F0&A.A>3U(4W+2'>_&P0PQ@<A9A)P2#(69X@*V)$C,PO8F30/#L
P7$&9&0H,CAE*IZ/X.^BA(C.V*Y?!2O;D[DUE/LBG?^1_X8%72_$^:XK'U>B'H-OD
P/RVDDN&\ V;0VRQ[8\9XF S?,&SIA8"R)[R*QFT+ZW04,]!3""\C)SW&Q)_Z\%6]
P:PHM)V]U[N_#[BMZ[BI%B--8E[S/_:WK,C"/]5NNP=,VHL);#GL1_C?6$LZ67; J
P%GP:$YFP^D_+P)=#0-5Z<5RHBR-Y!2!:[":"=YE]+H(]2)O7:,%M*ZW5H7,;Y:B#
PN_+4D#<^)TF<4C7_$)]#Y+M\I#!WTZ%24G5HM"KHSZ*AQ021SJ8T"#@5GQ;KWJ]1
P&5R]&V+D-]GD?$0IU80S'1+T,A#Z6R=^EAUS>61MOU>/%^H$;M6.0(,$2!4&6"RQ
P"L)XS.'TC0=3@% 7NI^KC'XE!\&L<F\)[\H_ N-6UV3SS\AV$[6#!#HW4*SB>_W0
P>,Y*[N:_X2U0V$M=T[:1OB*;5.-UBP Y+8HPRSWY&UG40Q1MV%+E6OH'CO_ JMUI
P4 8ZLX4AT3E^)0A6RO/VQ[EJB)>/,:;UG#'YQE..7/T/G,#RR)-'&KS9@:@ 4*#,
P86=:5X3^UL<3E?GT'ZDN&1X>K4K66J1J)D?KE13A\2V2^*+*-D<S/L>&8,S4P*FA
P;Z;P0519?Q:W*ZD^\*@!*O7H16^H0M8PO202X-%H/#N'1T.SB*Y;;7/?23<J?&HJ
P$K)_T-FRK2\^672B@2$@;V:_R)HXB?0^]ZLV<[Z Z5"1A<=<.ZXN"A\2U &_4-M[
P9-=EANXZHVNBQD&.>Y P=_9VH6 D\8;S$+X\+[T_@#K\6'[+%.K #[?9X0EG(R:/
PR*]8IJJHD+*",<V5;IBN$T5^<T6'>>SXK1O/'CWL-2N;/3S;=8'5^+4<N*4F/*K5
P]K(#U\- JEW!B)+W.;)K@;LNB<E(]Q-54S"T#RD^JGJY*7%@/Q4V%HJP(I*F[O0G
PFF;\6P%^#6*AU6%;ZB)Z5,S.:>W"+QN#<?N(=YU?1XR28\@M E1(N)W]R6_#,'89
P@"7-CG31!\-(PLL8 ,=:9X(06Z>-HNR_OU22D!X*OHZQO'!98>L@\]&85([3%DF@
P+H#@\24=/:(> 3P2B:YQTB21$E"*GXU&ZE;FYO#-[PS) VF=;]O2[S*K<20+/^!O
P0:(S::M$YLB$\,$IQ_KL(5"_X6-9 ?T"&S(WVH#>A;^0 M[ $'VMX4N3O-83LG82
PCCAPC*"?^#6;0(\A<]P0P=ZPB>C&?^"V/W\[I*N#_6!0ZRC9T&Z&YLC>E1,+6"<3
PH*1L? 5?PQ?>ZSE^O NJHE%&6 PR>X1:2AO==O^PX$_(WGQC'D$G22>SZ!_$"&X3
PVQS)'-W("QBR3XN$2>)QX,#[3ER!.X-  Y85&/\.C6(7@? ZL'01]\2H?(Z\V/MA
P?A&KN@Q*\1^5$&]"07DU.=BI- $AYDW$VA<C28*D.'R%4I?@WZ#MT#Z]*7^?NKY@
P3Q6CV%SJ@::,ZO.(*I_M:&Q'%:DX8 =F&%!AN$'ND6-&T=?WM%2.+$6(C#/DN86%
PU33&$XLX2(C5\,8(&VC]NTO^<&M>1EQDEA0PD;B.Q#"@;JI6E>&<8W#%N$!J>NAO
P)1NCWC7HOO2XL<[0M0JX:G6"^/)@L".Y!AU6#;0X7:7WLY\-O%S[\R7@_Y&B9=/*
P=><.*5$#W,*2VQ6EJ9'-DE4OX,Z,O2T6CCM!9R&)@PBT+$0Q.]N1):W); 1C(^F$
PIHM9U^/OR&9/ U.>J@;P).>6.87T"ZB8H)IA*2 E5HB-EI7H:1" B81_8$.FS.+I
P,/OH) / \@;/?N035"LCIP,WF/+JGT 2LA1N69$FX8ATNR>A$;I8H5#*A*7:20P'
P)LM"]ZOBRU\X6_R4#V@Y^H*/ZD<NUN0XP </*Q[Z#;=W(,;KZXDTGKM]Q#@G1$#\
PGK[08?%_5W4%3/0Z"5\F/QP/;/?H5A[JAL_.D#!10PZ_WHF;WJL[1H=+B\K[@1UI
PW5^=%-/F6+0;W)R$O??(/N-IGT%@SJ4%%006ZDTU>1[;%>@KOMY:XQ['9=J@TT81
P_S;,D6KH7W01LQ2-@!GBUX?53R)%WC]BBD[8\:,C8XDB#45'/M'[TGFUN32<'LMR
P&T3'M]$;;M62;&H"O6Z!PA'P%C594DYG;^%+>C. %%GXS@0J@E^O3/>)S>_F_%I1
P++#?]<HV:.0[;-P"ACUYD/5NQSN@0<"8520_.5Y! 8#9$#\*H%@:>^"$P2$8M6K 
P@^$OU36EC5>KGE.:>X/3^W^R/+&DT6%L7KZE"@"A![V/&"T"+@R=+L^?-9H:"7>R
P.>R"AKT:&A +V$=B^A/0"=S-Z<)V+47S:N2JGC"NKB@WVD 1G>>PE4N-YQC^P2PP
PR[-MA_Q,'U$5PGN+5*068V5]]V9:7=/JK6 34V_)V3FA12:U51E@/*0Q]4UX9CNN
P+6"TUJPO^7N8$S"#D9*3FG=>LRL7GCO&)5_D'F<@+3M6\8C/:#TU7!O?HV+FM04X
PU%A!]!VEGAKOT.P8A@-!];V(09+J-9C=B2GCX$WF+]B"]Y.HXPJ.*_ $2(<5S$P7
P%T*!^DT+#2(6.WSYJ8-<CG04H:*Y?HU\(!->#8'FKBW@-^BZ;GL3"[\WO+&@$7E?
P9OQ]K]<4U^)A#L0(M?HK+I]:<F7)K/I73]Y*>%T!I&^9[EJX!-<,_9L6+)^&:/0#
P0%QN8ZLCLF=&I$M<"WR[T  >"E]Q%LN]%1QP]3=:TDW&S/,SV.IH 49!WG?;Z*%8
PO;?46WG9'&>?19D?44'-=$6 /Q/JL:TV57"NO\!;ZD9 0)Z(CI2D,-URUKT(XOE5
P3B1CH]30G!=" 84')W@_($"A=;_/N[<-JG95#/[4VELP<UA1/]/S[M]06Z=(U8A@
P(?4G;%BJ?"'MFU 7,[ZI%=V,Q4K-Q4 W#(H4$+73KDH/1GQW26B'%H6I?(\#$NC.
PQ]%ZZYNC.;U9AR<]V=SVQG1K5CROX<ITS< H6F8++O@F!8Z295;1/\G\^F;;\G-G
PD\4\YC-IPN3K5LTYJ]Z$9V35QSG@7N8I&9%OASPQD*XVT:GZAR_92<-64OD>5DUY
PS_P!M>9$:6+N-;JA$ -B(H4?1P_'=XYXU(ZV/;$<5N(TOS(BLV IC$GB"GQQ\IUC
P^_%C5#G+0U1,->+BD>XX]CRCM&!EWS8GH04R%"[]PENV-/R6MN$S?^!L;%Z0@L/-
P"+XO0 H)>Z7ZG<XRB)K1A>((15=(+Q,FC[S@]RJ3BU>R[0=DI!_JNX-&W+0(JM+E
PPFO-NCGS9P6?)4K_\.R]"\IBBFD[4^U=3FY7;G!.6$'YZI510-/4C#Y-6DW]I9NF
P('9FYC3NL_\_&$)>_$?#;PHR9SDI/R9\](XG>+ ?J1I73&%Y>&.+8W0IV!W1K9]3
PS&'ME(XON+M) \M]=2#K+_T#^I -)HNDG;;_>NQZYSVV/$K;7' L[1.HV]V0$FZ\
P&<!@C)#COBMJI<YL5&%5FB'CX111(^0MQB7X8D7#3-\A-XJ9IJOKL(E_5$G"[9/0
P_=?*M%BX3RH_\X_Q.O$%(]6O^*QM%=N/-3K4/-G0;7'W\5N(E(>L*B?3&\U'CTWH
P?V:G1$Z;67>5GU&(MW?KG=A& D^#[+$\+S45I#"XN00UZV//]GHR]R=W-LK#BZ=M
P9WCR&GQM.AE#OL7NC2\<5D7R[A$>6#AOF3: :VQ2U-OE>.4E=4<V1+_\ P46-,8%
PC520)C7<IN4P;L7>6L4CI+HJ[P5+$[/CL-<?Q":Q+7OE7HCS(S10(:0%4K+K48DF
P+X75=-J(]9>*S/R<%;1($/&_(&L?- X8'VZO<P3C)Q6WFJ"&T-Q&J17*/J=764X*
P*>K_$_ANNVAE9"ZT+%LRG,2_=0C*@\:I]?R"%B[9XE@+V*>7&#@@M>G6AFJ%6/>[
P][-P'P&'$OB'CZMXQ2AJM-K35%24@.>4+WU'4!DRIFG%S)RB/].D\B-^]L6].NQ#
PLG]=+%-?RL\_83D5S/=,/ 7SW[$1;@X HY7$L4IF6!A3,-!LEV$F3?LIHO;_T1KF
PFB^PO@88_R5G#G?\,XUB9@=J'C4R<KVV\EMA1^&*0>LS#+-%=O/-@HC[QF%ZO$_4
P&_K@""Q57YB?ZG"XED92:@?\6C>?O6K)[D]<K(1/K93.Y#Z$)S3%5C5HC!3\Y <F
PI%8#5,O6O+@Z77%YG&I2XQ33H/WFA=FE*\]I5DRGFIXG#O*:S;+RM.F=0T1_D0Z5
PBBMX7U;$(\QI^%F,K+RB^'?XC K@+.6U8EZS3W*@@.N%0WD45MCKX*C;(*@U=-OP
P;1$E)<9BT_$"&<CWP-,@1\A.<\DMHRC@_<3&(II:=*0/5B=9VCR ^S2VGE4>8\!,
P==+KM@0-%^H3$88H"%6OO6T7(M2+O>F.#(U%=FLH8*;F>G%U\% GZB&B*"9=MY+ 
P@RO2LQF=:T#'(6]VB*SD=H5T7C_O@CR<%?C403$F!SK4=P,!/4)(H,9X="X:SY'K
PZ%<*.")I(>FD;ZS0QNE6LK5;@F8!I0('JT7CNSMBA6M;^2_R3CZ3VC)2X!<:;?,$
P3; KGXB&'F"@X(#11C@ZFN*&AQ9;$*J('X</4ZGY-)O>3<'+HPO80S-3"*@=EJ!]
P8BHF#+#X*+2<8+[R07>\+PES \\!KM(I-+9B9;#($QL;;5:H@3Q#2#MR:*-?N!;^
P$E%8@'W&K<PCE;RT-.\1N\M,I1Z70]KF/U/I%%[48BK<99RZ9BG6%@%]4:@_S#*/
P<1M@4BT\)+><V$PW(O$JR%=*,W*! FNF_$,)!)ATV;)@=$;BFB3'+/?-+"8A13NR
P3N9EEN>+'1LPOYVW#%/L.DN_FB6LA2I.-) GF;<8HEAU'5[AL0C.;JP&TH:]7\;$
P?*K9(JDNRKNV>3K30B5 ^G72ZGZN#+OQ(1@_3DR)]#5A ^KY[KP'MOK'OQX1>C?P
P"^"I-/$B3T:H>ZE,G-FUUR\V5K9(DS!4 $2Y]6<O=CD,FB.Y^\E?Y"])%@M&&V\X
P0]$-N*$PEMGI-.NCS-A<%=OKNT2@<6)5E]:1,NJ0SAG6.("X)IE\3]QJEKBOE8^$
PU&TKQ9)C!E8NDJJD5WIF-T/9&16JIVE\_$4N^LPFD.M% =N";1R - NHE3J2XYY7
P]^>2SS3/2Y(UL*S*6O4<.HN( [>?9G;[ !51[7DKLT,C8WX,)TX_]%> ^8<B"D,W
PO$O\XW10;:I=MBR_$LQD^@R'U:E';.K-^@" @-_Y[LP[+)UG5QZ@^R_[#&/N<TC&
P^D<#XSDEF5C*M8J:VK4A,4A,0+9KT!!SMA,:/9/M<,A-V5:Y02A#TA7V[=]*S30+
PC)H("6>2=*Q0IH@QLSJB%E@^D*L)9MFRT2O_3 OBD>JK5S_<6FY]'4-DIB,M3BSF
P=-/YD_5F. C8(UYT\*8<VX'E#IQ(@H ]=BWB0,)/2/F"&Z/IQ 06+!UXQ!-' 35 
PO$C*Y0."46.HYD&[6V# VU7'$5IBU_F(F8KW4G\7GGPQQ:X@M2"ZK?(O6 9[_Y?8
PW#^98QEE21K,N#!CXP>75P!HG] .XT46R.V&^<F4R?/:I-"2?0-;/LQU('>RF@N6
PL0A@MV\N4=*GT3B>='BE6"<<4+2H12M@23CL,?1R6MT*B-HAO^)U<>!]F&4!16Y"
PD64RK7F%CMZ?4'_$43"R"$&L08\E2M$:OGU7@LOS8L$Z"I4<AF3A0+N/'CUEH!0D
P-[$="R41&+KXC4E$&%%H8!'R!58B#<:@C6"<XUC M' ^DW\8:&[ Y4J8C\7$G<G&
PH=8]$=0Q4;HYWBM<KM'NI9)Q2-:WAV2>F#8/U\WS5\Z-VU#?*FC>1,L"1;87$?1!
P>QL<E'8SB?,65@L<]G:B64QKX$(@:?)=#(@H=V@5&H@@H@5:B=1#NF*5?627Y#_X
P<E49<,]=[/17YUF8Q+LPS5%#;O;<2$2[!;6^'DI$CQ/;O%GOD\;QA,7"9=4O:8I"
PEH#E&,_]P0=$M'4-E$MRMQ1!M)\8\C5A^WFK<]BP\XT(H(:2?52,)-@(#G%&]>4J
PWJ%<U.[J>BY<?G/R_.KW?<A$/*1"E -4K#BQEAGC/ +MAM+%7TTU1D\$(2V14[@9
PBHCM-?O95%$,F6/PYEHJ^4PLKOE6;U94 P%F.)E!+,=:\T0J"/GVC/TH.\35]!G%
PI2QE8.N1 DK$A7C6(=>H3Y=%J7U4W%N@%YDVLJ(] "AX%K7%U 78EYJH/&Y1$NQ&
PR@G-2.'UF5#':22QEM7X[&CO=.1T6,\F7$1H@;W-71*CA%IC(=O>&G"!!*8[S(40
POI!0U2&9/?#&*M S>/*<_(]4E]#7_VS]J^#CD9:21=I)"]^E(.U&%YW;LP<8IVTH
P%&7CXEUK95;. 1QQRF#EU8.=E-!A1L91#'M]SB$/GK]E[UCO3U>I[JT@M_K<."WS
P4*BRH036)+-L+PS-?4KGY(TIS77/SH[&S:E,K3P4[Y?9OY 8ZY>#NE("U+!N;*N?
P35K.5D_2%@J#%EXXW1@;DPBH6@[.[CZA*-0R(NF&*$BFI<3G*6! *T(\O'1&HI57
PI^.,QOI\K4TIFZ>T%.*"P) ,EU0_C'.%(N3-@'%3>:K<?[*W G5]U<?4.DD7IA\;
PKN%D@8$1,F#IW.<S(6M@1F?,5_E_T/+/=OB)M##["QHX<,#VN7XNNN<<A41O>]_5
P'%CQ3D=J, U$S!"IL9<8JG. V)X%GKX5BY79?I;AWER8;FZ)B>;A)$?%__LZ#DQC
P<Z^.V_-%/0!A'97/AJ_B:4\]^P88,YW%S4[HOL+L>::)"%RP/T+]3A"+^!_"*7;L
PB+HR!Y'YR2TAQ1I_K#?[;6H@^_&9!8X"!]#3 3JYU$K1O7"N"\8LGM6<FRL$$[&U
P""D7]&*TK&2M"=A>[]::=F4/H+O'UXDWI^Y!E9-]B3#61''K%[KB96"]K<^#&%T'
P:863 WVEGL83$^$EL]9VG6&?>8^]7R"PWFM9$#0QQI(>6QCR3+=:=*IS+PC%>OA'
PRO/=OIXX^EJNI(4I[&GY;!NNE&[V>X\<4YA0Q4='ZA(!XZ.BI;7 !I#<<V9;UD33
PR4.CD"A*;W"5KJ=@6Z8M9>""E3WL6:-TUFY,[0T\44 ^%Z&!IX,H;1,36FO/D_QK
P'^:V0J<7I&U:SNV%YR<:_,ID P*5#MF[H7$PL\S=PDH7J?"$.R8,O+DG5GZ'+-WH
P]$DRGN.UY/H:%>(R;>,(WR-4;=]ULZO=)D:@E^HG3^4R81;'-\>-2II!V'8"3?L0
P.CQX !TZ)+ E48CL,#E$M'V$P+D?<>-S(Z1[B! R<6.^>.(LV%1 [3^D5.WI+R_5
P@@)/ -QS*O&8#<B/M<EC?U[+LSIU?]UR)[Z+K&4OU88JXAH)L 2"U?YG>;V37!@8
PUN(8H#;];CH[Z.S!CWDQ14NX8^:UX&OT!Q[VP(%BS!BUOR#'-PT.'&Q:YH*O_4^[
P&\!"2MD*7R#^H!3T@TD98R[\:CBUE,WYT#_A8= 0L!1)0R%I#H5L?Z)X&IY;O[ZY
PJ#OF2#NW[,<<(_4+&$TSQA05N2*C"J=\UAD>HV[\#PL][&4&E6E$ZT,Z&HE1+G5T
P*L5[)VLT71CIYG5%7W6)-IWH$GQO-M"_UR<,]4IEUB9M&[9_P#NT0$Y9:6;Z@&TP
PIY]?.JSYPQ4ZD<5"<YY;H@F;D&<S"QO+VDP&PB"=69 @LL><_J;%'FM.SVO!PA@'
P*<1F$XR4S+OO=.UV<1ZFDG FF(*[<81KZXKB6^LM?]+[J[8&.X&F Q(R[88B@9GU
PO_L5U53B+](4R+Y\7Y1JIC6T<S&?+MV[#0N_J6@0*3K8!:K'+;':"* MQZ];PB'?
P3A#<K:P;ANEXJLU1&,86W9A%/67'6$@%=E>=7GP)6N<*EW[<G(4I@*H/5!1?T,_2
PF7@5=Y6=!QM4IY!8<;7=$<?IG/9VE93JEFF=?1'O-V'$2U@(D$T8=XC$7*0"9MK@
PW$-,R#G8,"O.L*DXRBR1A]NE7J(?B%?>ECX$L8I.)*7 5TB=X/VR:-_&A2=52?%V
P?!A'4$Q8+ZA,ABGV@#182R/RSS%-?H"K#;&C+<USZGV1G-RY'MJ QW<<#4BWT>R?
PV977T7['M4'$0>B=6\\\7A8$,=4#03)&@R'")4"*'>L.Y:FLF<*@'_KR.[H'!?Y^
PR,#K9UWVX:I+I_>'J%\'J2OI9@!CBZ_$J'7R5*5E;(S+3'7E\MY!^OF].E+05FJ>
P6^7ZT3BEL1D8A\J -5X-UP6SU;LYTW$['TU.D? %V7B#!.?SU2#O)RS^)B+K8)6O
PMC<)F$Y)EX6< /=0Z<<<M4Q7YHBY]_ML1U-Q!HPD\E)A\)-3];<]1W%UIPN0J_IU
P'VTKY99<WWC3GJAD,<U,1,;;?9%RMRF5H9.<PG.]WDUNB0^U'D2 '[67K'&=Q <#
P'$ 6;2K9/WWQ5ZYZVQ5^@]@(4&5Z=0R]-?FL&%L(7@%!^I&;%S=?2M1CR)*V^<SB
P#2;A?2,#RO@P8NJ$7!IONM5RZJG"%QL+U%A%&'35%)AFBRMA_D6KGL/O2)MY%N-D
PALPTE(A=X2#&_1OR@&1L#!/DTM.^"2O57WY@.2L&(W]WA>+8=4U8& Q"9P/46R'>
P"7XX=F ANF9*H?]>K-LLOJF?16<OO-/WS4.U 4PD))2,G6GN*W@M4HO,?V(J4TQ\
P7!-J@H00LQ<<CT1[:T_D2$7;E:CB+B3-U:'V-L#YL]J6H./D'RK>8C+PG8'HIF R
PCJ.("]748/MEDQ\(F7RD[C5M5MEI&JE.YG%3]M]G+86+*<4JACT353Y6X8@LY"SZ
PC]2)2!B*"WM<TN>+KD*C_=M+Z.6XLE;@MGB=#E.O!K]!]^ D6$^[R%Z>*9QXG7/%
PZ(NO8]KS^BW,T]T:V=W'))L(@#-]YCCOS-G )Q\>P'K $XY>E_'AG6>"7O8)W0 K
PT@: @04I]SO$U1[H1*<G>3 =$PZ)F$[XT#Z[YH$J3=C4SR8BXR8,6BND0!]'>IW!
P6CW*>&3CCG1[;YJ*%K13&WF!H8<+>TU]SM,@:G4[8$(-5<3TR0E?G#GR[\,R;H4@
PE8.[88:PD5+20A/+]@<]DF6OZVS \'KG>:>J>[,S39-=9IZST)9-2IS[?I#1\TH^
PL%Q2$ 7D[0[(PN3Q3:QSBE%#,>"U)FV]TIO#T(!"/T<UB_+8DJCFBDAZZ\."K[/4
PL+Y'M.?Y6)21/@Y;2<I1[X4?(,"=6#G/JP?^C9*U !X_+MU!%4H"TO-RO[;&9F7?
P.:5PQB&\;L('TKK4G#@%$R+=?BA5&3] >+Q4=H(CZ(M(S \E*XB17O13]W.F;'3*
P[]DV]E[M6>SR(\DVR05?!!L28O$S80F/.&JKMU+K$?J/4JOWW9CJU4:'YZ2:.7GI
P4?7VU32#D">%QB08;B2C:X+HA@)_O/FL-Z\HL 6L.YH.V=]'UP350$MW7R0-ZOA 
P0;+NUDQA&*Q"Y-[V6*SDTB:U% CYO"X/!$U&)P-6&C*[L7@O2ZMIG[J<GR.9%I#G
P=<)2I87\:_(@>7P]SZL>>GJ/.QT56'X]08+@"S36JX)WN%B?SG8];8*LXZP4:;M4
P"D JG"V;[:6'N=* MM0B'TO+K /7?G/8.A31/"-S.J172]V&X=!UVSCB8,_":Y5;
PDSZL1+.A.K],KV9&>UG#5I39LL4!)/^W;@DX:,RRL5POPZ$F(=I9YR45C7!@TBB:
P.NZS[2RZ>D Y_0@+8&/#H6?#%)2TU*#;"]UI^R:.21P6M?B44AJK*[EL9:8QC"^/
P0X--^4@^L[(S4P$7_W>M;CY4MI8-D0*CGY\X%!.@@;Z0E^--$*PN7C=77'#BO3D^
P(1.G(I]81$D,TOMZN,$Y=C@[3LGT;2,WDNSMJK^] O\=]^R[L\(%J#\%#1FQ(XT=
P3SJ5IE)@_^J \]-Z__]MCA&W-]Q+/3ZNZ(=K'IQL@2M(=^$AA* 8M@0"0ENP1&[Y
PK>EM6L$=%$[;]%D2<6%#SGMAXM>R$C'N<]N*=8K"&JDO<X)T$HDZP,# X1&UUFK:
P\ 5H1Z_2:60N['6IVA%M S./HOK#W<-2-#^[XM&$,+#0SNAU"NX@=XF8+E^:_GH1
PMB#-(D657;8W'/_L"1?L"]PE[0$46$W=[ZE4@/5)HC)P#Q0%-P2S<#>X@@$/NZ.*
PNMV:H4_6973H'==: J1<D.4VNNJW-GJ\J,<-KFOD1FE6#9JA#(ZU+#J@D74GSU**
P8S%UKCFO@P 2[EG'$2,<T#@BCLO0Z+P",Q\B$QIB-K))%0UYLB?^_AYL*YTH;O,M
PIOB@0B4])3 NZ#]<3!E\(I07IJATDR-[9$Y06KX#2+5::8OUHXGQ\[5KC7VE8FS:
PV@$G< ;S&*3EEF=$J.UIXQ'%)>HKP[Q/S'I^),.<&L.QU[#M<XY1;:9/LDKD$^Q/
P!9#2SPU-?6/"7W?&)*;?>DKIL!692PG\+(-F5:J82GJCV8:YB!2!L]=I\E/;1KY^
PE7.4K'$M0O6F@1ER/^7K0Z#?8%80BHJ2A7HA.+6Q>W,W=M&<S;A>.#I^%[TT6S(6
PEC9P:/8]I,FX&9]26D.Y*^Y,H"X!(V?U"<N(6AZZZF.WT]:.]\F]M$,VJ&3^K2K\
P%NNX4L.,(]/XT$RF0UQPD#1$ITVQ0[HOM.:1,^>LI)UMD,998XWJ=BN-&(^QBYC8
PZ@,E<Z53(H-"OMWOV;ST:F@U&91CBN=\74%'-B\\>/MU159LC1>79HXJV8.,.Z5C
PP@B@IDP##0X7.V=4?!)@0DP^"X^9.Z$J.R70]"?<,-Z2J?KNRF1/V':4O80)#DDK
PM$1GHQ+Y,#5XYG6O[F;#U7P^X*^<)U5;5YD%6O MT^7'+%*T&@B-W)_@&':A(=AG
P81R<T62Q(@1V%#VNJTOK?R+[9[^6'2NFU#++>6;F?5H57Y"J*D*,KXZ@]6I1 7^-
P*9# QZ0%=^:FMK#OBTSBUK)G95\'@$XWS8N^//QG#_#2+8<'T^4R+1ON2#N:X.+D
P(F_"3(WBE6_/XQ^FUY-]6U/?6I8<XEG;*4G("C/PFM-E!R^MA\!6*^I;)X7M'2!\
PTX"W<*=CA\*&E+'.4/S3AF!?D/9CQSAK=$I'^*8K.-W:F7)G%GOW\]FTRI=+)&3=
PC"U9EBZ\P#TBZ#?G!Z)=<>F<\_:_@[+22_#3"#;L^119PAY#_1)FT9(I93Z'% DY
PM)\>3W=,QYV'OLW></!WF=S+@C$P),X+6\=O>CYK>AI5[1AGRQ+VX!DZC)'Y\!<\
PJ[#H<^>PQ(SXR9X5FLDD!@,FQ'>0!@*2V[LV$@(A=*\DX4DR-6_D5TU@V80QQ5_>
P#0+0SP.5IBA"O7H9FAY1A9C.]%:^'8L%.7S)05FIVDYIA68)-Q!*PZ?L[O;BUDCF
P FL\]L&+A3C\]9B(6JW<!B5=>"\UB4JH#E!^5QQ@?&8!GQQ*!%1>K]C-Y2X!+!;1
P&WDE+QCP$Q%_Q+/"T1%I.3XYIU]PD5I*[9-<2!Y)7<L^K=+!=FF=FFD:M4CCX0.-
P'?%K*%1AR<X>]>=T\"4LI\ZW#\1W8G"HPTYK\$%KH[JK 0AH%";!-BF^K<'?=*!P
P>/Q+R9O=#?0X:V;/GW<Y]U6 O\*>MB*X6'\&.,O+*R;QE>W3+/YI8;4E U6(]TY(
PVG'2="C(ZK746OW2HE8WK\)Z@RI=%&L[F08T8EGWT'O[T4N(7IW_=)LT.D$$,TMW
PE@H; >]1\'QZ/K!OD_)>Z#QHA2P&V/UZ[9:X701M2^%7.QPV8E_&%-H.<9U.F#Z&
PQGW+'G/"W]2B-B2FG%/&<E'#4/GHL/QC)UQWJCWDLIC"2O.JT3KL&4)-=GFGAP!=
P+'0[*GN+5+! WC35CT;,+G/A!$8^WO*<\2J[V,8Y*EV\6Q"18%[62RMYC$90!2AP
P'MPHRX#2+[=<TJV1^/&FEAOF6Y'6B%$=]H_=M[CZ0RZU"TD^%K"X)?J,N 7#W)7H
P%A8K?$QK_5N),AODW F*"^'*[B6'94-A0P(YC$G.^*&>WNB2*IH5R[QS]_+8V QW
PPVO5AS37^4V<DGD9^1P$5FUSW-T++UI7&C""^"_M@+2OVQ[EE5XP1-9HKPE\PQZD
PN8QI]EZ_6GE<T(D)!XD=,\K@O)BS"'C_H=2/:%*+QD(^N)?/:[H"3ZV9>ZNN+)!V
P<SC+7+V%4A2L![K;W;.W\5W?3+Z9#0-PP/FH CE?;@'%VAT8[F ;QA_\9X"Q!L;*
P?;Z1L8$]K!8[FG=O(AZ@.G:;DO^=+7.[P.+K;=ZAC2610/.!V(NKF/Y9(V4QZZRG
P2<5>.#!L1@<*&9Y$$A50L@Q\;"Y3P2GV%+B$STS?=HL9/YL]_A)QT&9>(40OLC7T
P#JQ9! QR,]SA4K!F@Q+Y. 4@T^8VT['^?7ZJ@Y5&%VHF37!A>X;)T'BBA*<]UD7'
PP$Q6^=0J*#T/_Y0G=7,&'R%<'O8,L&IJ8@;/O*'$@,940F#/B^[L+LYRORZ!<ZOY
P(/NRZ]Z]%A%80PU^7A9<!=60/9X5SY1U#@[I1\8\ 144ZGT.SKY*@JO7<\[-/<4*
P;E)C"I$99$F?+?J->JH2GH0Q<RH45A3Y0WM!$J:7&VIC<ZD3/J2/N'ZKPQ-+5 -^
P;VC!2I57CJ8;IK>U;!ZK+*&JT]"[==;N-@+7'L%5L*,L7R[B(S;SUM:H4\4P<^^P
PJV^K,B;_7"'9=FD8'$127%)25U-=#ME@,<UN*!VZB3/D,!V"+&)_TE\@0.!?_"S%
P)#+/V$2C;DS_OK+.ETU6!9L:N"GT7[:EBRG=F8A-WQ#F-0][0UK@*:=*IXP11JW1
PSAV.FMV@,V/XY!1()=40@_(^$G-9&7LEV4HV9IO-+)]@E.('_6J5#ZPV4;*$P3\7
PM(@GZJH_3I56.@X"JL?MG(ZL,V3+11+ =)5@KB"R3_CG2%?$ N/S4!&7>M@QM7R[
P[4:*^]@&&G'+"0_&$","@JL3AL'J85O,@<D[X[5]CJW3JQ1E102+Y?7RP\J$K<C@
P>>Y0;F5UAV*/!-9/4 $ZPYO=(Y1S6)+[4Y(A:(5M<@\1'_^L%O\4-7Q79;7,(-N^
P_[0,^'/"4<G;G-22**<B%H^)<Z;IIPM,-WV,KUH7P!K<%)7[2MD+2]$Z<0N?DK]X
P;N5Y,8JJ!RQIPP5[W)5V?Z3S\%_-2+,X"";HJ<A*U'#8U=Q!7W_PC*0$/?>J"2H\
P+&8K[2J&[P:*^0X',6B)>1*O:OD@1<HO;6LW;WU&715%\C]"OAG/3UO_.A*H!V:@
P!FRXZ\9!4N%#94X.K\A#;0Y46&,NOF5"W !Q+J?M0-R^,"N(_-/(O,;,)<T+@.('
PI[4,.,,>E[YYOZ<):333VID8=V"21[MVM%$CT@Q4GDY3+-7,-QL.Z[I/FL_*\.;=
P5*T%+23H"\UZ1?)\:_V3<06W>6KQ$V<10, 5QE1&@]F\/ ?7+$WO\@/B#LP[O"<[
P=R9HNCL&2KL [+T.M#6I!@EC:W?TV*,SEF6.IB20NL09ZB8_E]N6$:=8IA0X4NC:
PT^?Y8*CCKX=*IWO4JQ\]:&K!9(6:4+S:GCUSV*- Z*L!Y/UU=02N+[ +"_2+Z X&
P-/*QYF(6< <Z,S'FI6 P.?X!O^LKM$IB=^^+(C+WZD\$*+66&F<K/-SSD]'P$-4A
P-G'A%F'OV.?'\-ZT"QB+)D&JX#R6\#=BVS7>+W:' <%'%O>)1C[246I&I..Y#04?
P[+@.;!D-EUV?(3?;9MKDQLR=YH*^"VIQ+M2.;6NHX1D$VF(0T)+>'?09-3<JB=NY
P#-8_2_$9F^Q(Y+-%.9=F .O,$F8?P%E72J;N4:)"/HM:\Y@\1Q9%-'!!A^/T>/.W
P%*WMV6U;C@?O13MP .=]?L=W)FD\1'YXTKTWL!J=!:&W$>V_XR6_2I2QMP+C"B9 
P W+=C[ VQ0_.:GA0>>:J@B%JJQ0F;#P8"N"@8M&'C\@=7(#X+K-4?54JE<$7,,M@
PHZ$8-,RR6%#+/UZ>.$ON8 X1Z![%A)JL0YX!BKI-R2C^W*-E&Y^II@ FZ"LWMCI^
P:M@NA<F4* 7D5_T]!(Q#D27B0X[+)!'U/((*O_Q=JYMM=-7^W-Q8_:WNB =# [,U
P]?K[ZF= -&D -=<84-7>KSXPI; G]OJ/=A2$RCI_9_C=:.0L'0-PY^H7']E;6G!>
P ;&P@,\L>GB5WTFH H@)2^4;\)VW/4K(,LRP.L8#.'_%+2 SB;"WA ^7NDV&IYR+
P828 ;MXOMG0A9^:*7X=O0:SUY[(;#7TM+R][ZB!_Q[QR]66/[_F+F3CR$@@#QJ^1
PFM3E7XH]4@M1'N<3P"O&!7)-<PGT]BS/S,&I+K\LB(0"LUYK 6,[-SM'C81J.WI\
P\W0((*V_ >A.A,PT)V\URH*]"%39K59Q4YL*-([7<21(THYKL:HXT0F 'PI#N\P^
P<!#Y\0 \B-[V#=,%^5*-TKV2Q2XR1QY_;;),C@ST$G4@WNP/ JZJVV7G%QPC*.([
P<,#*W:OB1Q :!!:;Y@[W6["5<]>[=P\#(P]6-61_6?Y.:1E/#'XJE_"7'-JDK;(&
PO6I6KH60*<TC)2B7KU7]>=3E^6. !=%C4328CED;ONS"O:8[P#A]H7H1!1[$YH(@
PBCK'IWJZXJ4=NR>W.4DS.PH\-X&W.4K*[#H@>!A20N+W939/S_,(A=:?155R*T6G
P;CN_5\M:/RB'E#GG="S:D<)0F0+6C[($X[1K"LJ0(VZF\V3-.#NH>>E/A[B(YTS!
P+#>^6U\,U ,29XC_@-MA'J$VO2IH2S,?^;?9P')9-]'K,@O .9_8DYRC3;FYZP"7
P\_]WN ]/P"@Q!]1P%+\N-EI"3Z2IW,<][]"<8B/HXK%0EKS,J!>8!1D+]:(0-?&X
P]DA?T)K U%659"G>!(,)(^;J;)CO6R3"CB(9K$,-E%.%A^$ISQ89EA.+=IW4R.%S
PU[1JT R<3HH3TS6G*HIQ\9*!@9#(NB@!*]Q6'IRO43RX5%GP]D$AX(W7TV%0@6Y$
PH\ZA73G8DG-4@M5[E1'MPSM%+A?G95R-/M1\L_#'FWR &2'WK]G5%8F.U%!H,\V0
P!%S8:B:^<Q=Q]O[-KHEI+9W!-%U^G!//[,](V+'&HYA@U*>7LGKU); 6=I]8CD(!
P@^[B.K_UK&#C:;B97S6*=6J+=[[OBEK("H/NBLT*2UZO^.D.99&H#C.(X?O0H>PM
PG#X3LO+[UHY7!;B_=JL%3YB[:RA17'XZ>"&N<Y*;\3VB="C]3M8-S;/H621ZEL84
PD= #,WNTP+FF++);%RMT:(*SN'70AY11P,8F/<X<_Y)-I*LM,QF>-&_>NMW1_X]T
P*$%FYE(G5D<_AM@)N;QVBE+3.US*U8[2^B: EU9TD\X+/.3X\348ZDZV2FA Q%X8
PKZ0XT!+<;>,OLWKMK1("_%+P#14-)VP"BHAM&]8;U2H%LYX!.[@UH>R*Y?G[,(>4
PS)>U)SL:,VX%LL_1'JM!,K3&@#&X>4@X9YX"JEE6>U7^GE3GEZAD*;D>:EI6F)Z 
PJYJC+AWHS9$\>C<AJY,1)?CPO\7E+1X[09XS#I@(;#D]L;=ACJ14B?!Q@PEC%]6&
PY5.%:IP'3Y^WP">$AZELXA<YXIU;B._J4D5Q1_@>)XSOZ/J)=D$F_JOQ0)NM0*LS
P[]^:"W8]'#B@][9=+WCH*T>0P7<^E8)-11S.;R 8RM&/!,0ID+ZAU.VJJ]GD3M1-
PT^872 P$/U^F:XZ[EW=LMQ#,,[>!\H(^T+X-JO?$/1V8AJ_7[] "(U+,D9X7([QJ
P#+E,)>TM#7(+]I,+I-RIMSI][A$<3'0;-W# PO-Y[K\Z.FK,T]LW)G IR<6>90U)
PZ0-J5-0Z',9.XY^GG8X$=OK'1GNRJN;-9B"9B>!#V5-I%?)\P-&XT$54$Y(-2\@&
PJP/+'B^B4]L7$UM1)<*"^N/1U[TM9YKRS;?)SL@Z_>Y![UKVCV=/I\P9G\6LE4B4
P)?$2A3L.=NTY$*D$;W'W!E9I%;&U=Q+'=..%&9O5&3S<55@JU&UY@_RN32=<=^9"
P8%_24YO(]N"S)%&A>(!(!!4*A9F'0WZHBWI@(2+,;1,^:1YC&ZGO+M'^#Z.=OP$'
PD7\*HC,PL@UV2E9'0I\XJ?9-H,<L^_AM]MY^;4:H##'V%"'MTV$+Z+\O(F^=TF>T
PV<1(8F!^+P)$:EAYC&QY.2 "K3<EQ,U;SK?3$@QQ4W5$6C)6B=HCH#)/6;5(V8+H
PAYR.56&%)(Z+]<I,;>/7_H /8])M&9/'07T16N*:UP( [_ DXN5O(2HTW()A\M,,
P-3WB"T1:"G=/AOQT/WIK&4\5!D'X'+_^5M+I.\,RZE%(N3" *N12[1GU&V\<A4LX
P*I,@&/K]XRO-<S.1BZ8]QS ,TQ=2]&]L)F,P67E#2,.,EC$'70IWID6K)6B8;:&"
PB;F*A1F8QE&Q8MZUA (%+Z\_G3T"37?;>:];A'H^GA#K@;9ST)QD6)<1K^9GU-%U
PU>*%TE1F.S&-9MUM(\#OE[ZP7JE)P0^LE!P;[C+@9#C-V(#AJ8"<)*I8MXV[W^X$
PZ>QC->YXQ3P$_,:U)+?V$"[>M3J\VS_HS[[87THS?MO1&[C)N#.2A_H4NF!KN*2^
P< LQ16('M//2JH'*@KB/V.6\GJ6.'!=0<" NY,L/P @?J1O>1'$-HDES&R1%<LR'
P<^H&UFTC'08-M"2??R0) A7JGZ5$\CVKIPU91$OE;7JJ(SNS'(Y9#M\24C4^OMFS
PJ:V&0(W'#J#JVS*=<E5]#ZF[*V^*0_,?2+GN)@)(<K(GM(A'1B:+]V[19UW-)N/_
P+Z9C"78!Y3-0-S+S)=WI8&A$W!^(?3/?5%R/I',05H4<'-,_B.K@ZDG6TA#-8_M:
P-3F_C9=YP6=R@*#;/_)(R'81RD<$TWW93_257KVO)<Y$1_GSH@[YU;\!&"B<\X1Y
P^IY W-*AT!#?X[WNQJ-VUY(V>G;K74ND5*#M:=IJX/BIP!.7>5/#U)ZM52?2] MH
PM/2VS>[@8YJQP!I[C:IC<6MW!D=)2=I>\E\9HE$7-:)D9X'A7B@8$T+K/I#^JKOZ
PY6+&O8UV%B2V480X0)2JO):0W'&%;FC*/JAP$;TJNNWQ3A9Q2!CM(;6?E^DDHE4V
P[93DH8PF'-TP\Q&_$0;6HL0(,<Y1"<\*'';Q0LF H;'F:O5V&TS9H\[3"4@%QZGM
P51C"?G,%" Y.DM^YX>[-<21UK<@MWYK*$OFW\C0B%<!8]C8X!2NV=<'9^232?W(?
P:S5MYZ2Q9DT%N0L-1O:K&'U:HR75.]ON515P.+;_'G M[QP96!/Z(W,XQ#9<1=EB
PN2#AG19-*_#>LQ3" *A: ./4B+E]"/O*_PXZBLHC*>P.3I.B1^%(?G]@T&5"PNGJ
PW F*6/W%0FRMN<7=O]; T:#?_['"OJ>G3UEX6[0<AT,JAM,K.BV7#T4:6_)#)(\B
P[!UCL21N\E=[O^NJ^"/ V@I5JP(JL]_)IH!J_3R,[$"Y*>YWHZ2 ^- \PJJJ&[OV
P,,,%L(C,3M5V/,UH/LC 56JA+D/SK7B(@LAWDF17)%MK[Y6<_RL3F]/@FI4+&Q0N
PKA+T&'.GO$C0R*5Z7R? LHTRF1%'<V'/$Y3W=(J0$6'QAH83O/9^,9NSL.HAC?[V
P#FDHMF7ZPUGW0]:MB<?OZ?:+%(M[YZFS9Y*R<L>SH2C.]@9TPV%(,S&HNM_!I^&>
PSU&8]05OBO]J_CJ\(U;PW:S(+YMU@3)TK4M-W0A^OTJV3!<9-\>Z_C$3^&N2ELC3
P&\N?<C[18,_KQL)/E0Z:XU>VO]: F*+E(_43V"9V?NAR<JVW+6L3PC:&M1GVXD7N
PJ1CZ;U/*-: HBQ/Y3M4RA"V2@_PY,"O/\%F13CRA"=(U\244!)4 *2#W \*$]ZS?
P2C$TOF_;J"Q"!L@BY#=#6;-F??W& -!W+M^OE").QM""A'87_PD><S(1I!2\LY31
P4=HF2[;":EE*:)12),YE=OU]&#17XF%AO;EF-=;3G/W!@:ET6"X32!X!>J(1 _OX
P;;08T]L5YP('FXZN^W/&.7OYDG2WG:ZFB<S,@Q\3X4F9F 5V=QADQGQ\AR$XJ[YK
P;M_5\;W'<8;W=X.X>@;ZG['LF?3;?9I(1-#]HQ>MZ(0^O-@ SC$J7M[%QSZ2B;^4
P0OY&U?M$4)PP+FZ^^@OZ9)Y4U@]-E'+O]O(6]0=1<WS?XH']UL@>&\OIEWL1O6^X
P_Q1+.D(WL,-42S90;26KXI<(Z.,9D.P G!UJGV@62_^TS\@0EQD/$;6TVG/PC7ZZ
PW*0Q<9C*=4VKD(<C?$P>JKFF2EMC8B+337I,R;N.#$GSY/JV#_E4TFWLYF2N1#"P
PXI).$.S5[T1W,FR9WD.?P.Q6*#UP</%I?IW8;W##38R6$#H7?C)0JFS:-9I0!1WY
PPSK!=2/RNHW6H>SR060RJQK:6M3'SG.\3T]NB/O<G -]!\/SQLBN5L;@]72PVL^S
P()^=?-J)5T^%3*OT ')O9G?<Y<-<FE%"A3@N3:4N3U01Z[T="$6EN]0[B802XMCU
P6P\,)D7V#FS]9AFY=3@\$$[J-2W.ATLL14)[67SD!_"XL8A=W2^0\:-R_S:O0[C"
PBT+ZI9Z\XV7*]:9,);]KO=.BUHHETJ\=Y^FXDPV*.*$XZ 8O^WOJ/]<$9*V(_0J\
P**;(5]0$)N !%:FI_RDDVJ:<Y*FF"R"$7$Q+X.3*=6Q^S:3.4)2!=$@H@@#<G60I
PAVY4,;258G7D$O]W$_V*/(\%.#I['=IGZ6+XHV'VC<,4DS__,TX:DGI]ACZ61%+0
P38C]/)BD57Z>%,F$Q+?W:4#E)3[I>@H17?6V=:<KC8#2,OV9]OC:0GD<<84E.&\H
PP-]!3.CLT$\"*]_4&*9["%$S&R#LZGOU6 H+"\Z6^U7^0%'_"F8]E:*;EK$)B"OG
PX(O;.BIU#QPLSQXD8X=JD"%D(O!U,QZ;#. 6D02\6,4\+BJ,"+1N7%P4U#/X?-53
P0[LR)#RG3I8U+ >.AKWUI7]A'3H5XIRN(X/O=>WDJX1AT#8SU59G4KZ4(*%3BXF@
P"LG;IW]Q>TQ\L6[3/8-:W,P43T7MOOMUN8\UG-B<XE8KC?,K?H#MFE"3]W;4C81O
PG! ^:F?<,NYN-GY^Q$]HD>)IDDC6=PO: QRX^04FD<V 5LZDK2W2L(6+]/A'!']+
PRM$K+GRM- :?E7J%5L4RF]CQ9SE&HVW-#"S_I43NGQ#)^POJUJ05E0&Y-T;*NX+%
PQXI?HYO1-.!DMX] )72G./L; "J+TA(<C+55:=;=W)ZUAD338ZTBA#1([B.1R.O!
P<KZ7TE5;UU)M$Y$?1C/YL?=0/SY(5"%8:8(E[K&&CDHW,!Q<9];+P6?]SO%:/Z6V
PM<Z\K'3"GHG=)/7WD@F;.":6Y8T:6,,D)?K B%%G;IWUR)6((ZE\5([^E9K&UI,)
P)T^7[(YZ](ASLR0TOQ(F6N"M;TU.G@<)FS3B;(NRA'33;Z!TF$?;$<6B[I@847]1
P$ [HKU-1VMA:#)L=>NI ;C82@H7'@<8#K.TRC1%"@49(9A@,FLV-Y30(W=@(VW!O
PLQP)Y$><,XK=/'MB4VCZ"+$E)F^0F*^CZDX[*=M3<9[GH,OK4CD5J!*93:(PSLWM
P8, /SP8[Y.F8^]+E=9E0$7>\(T/VF8VHN3CK3,-6&S,%\K_G2XM_>_EWU]'F7Y,Y
P9C5CNI8<V,')+C[0\E&_WW@;]AI^C[:DV" T1'WA?@F+.V^]ZW!52QGVV.Q)VD4*
P%6CK&LL.F5*9R!=_4B4/O@@K0G? 80BY:+T:7*1KZI'0:U>F7&NY"CPX8SUB).?$
P&7F%H6C*MCD"R:@SP"Q-42AM\\AEZ.8<>_0KT>_"#E-D825<G_,OK.)UJ*=>=R\V
PY1APYED4J*]F#*C6WKKME4Y8@CW]#E\5O3^&GXD;N85[%^MU:-Y^J*09;*A3GSIT
PPJ4[Q"<-V:Q=G8@%.$89N_M5\=&AC2NX+RY!&$_]O,2_PVHPK>;#@9T.L).C;'#M
P^6>F#:)B.UNX:?D@-.BCRSRHV$%N2E-.E('MOKMH-'1;FJM&0T!V9TQH,SH5[0SX
P35YV#:,4SF$/C;RL8Z'2$_"S;!LKJX:+GS[0 ]P"&8T4>3[DM]>]!$R?03B?M>T;
PA-KM)8OZ4-@43$&R2TICV%!0Y2$<_'W>TSB04'&1C3\#K6D,+^3W:<@269G$,M7F
P.>3%:XF"@<<6X43S_^<JU,U[J;9ND;A2]6JQ0\LXI"*L@ 13X]>P]YN_[T6@9Y6R
P.Z=]/HJX2N>),K.CPR>[B+0 EB,!#K2Y/IWC)BLAKKPI0!8 3N2M;9$X%"W7U36R
P[V4L8!?C\6\6I %8R8..I*<@$/#1K:ND8%H1R]T>-D.1;[@N\<8]MH1,HKWR3KRS
P%94]#&D]);0;!<)UI#0F*6@]^@@+2:E]\EO(MI?Y?L B;K G:K$H!<-I97[@^I&-
P8,(]@!(9TP(6'_% .::J%>0H?Y>QTE6.EPM5RTP'P4^.X>' \QS[@(E5E@UMBG*R
P3/,.][\Y3H>,?[K!PQ2J6>3\DD]62A!6\]M"$R)0]I!'/OPP'N4VTW'>'[6"Y!+G
PIA!X/9X^SR6J5($FRBL"U09-0?PSJE>W@I,O_UD$>4LMS7/.*@2KU"ZFVLM/[J7X
P=,Z#</<[]C#[W\=:*UX'ZD1^PJ9PV4M:#3T*3M%AV!)E?.&**MPGH+U3^[$Z()GS
PI0K!"U9%A,J,!H=SP\. _U?S+%*_5[#P0NJ1]VHK)"AD\HK1L_)J5X6/=LR2<64^
PM*-4=*_)Y NHM^A6=M\O?@(UL]:_6Z*EH@Y;&EDB[@?+V*NR(?K,I'0,AMT_G8!G
P3I6UEIM3P%D31NE\ ;KL+&QL6]')BB3]*B5+XNG.SE.D'F#P)6[S&]/=/8?PF#+2
PU[%.Q Q?$P[F : (04,,S-?#\YJ-)5:QOA9/TDCY>4$L%P8WFA,1VW\ZT[[UN#EW
PEUO!1:_5J@QZYQFZ^.P<8)NIE,^/I>?H?&:2R:BN2[/QWRJ";BNWMW@V8O4_8Z)[
P!N/LQD!*MN1F[AG?)*@.*J67D>SJP5KQ4:F%.KNZ]1C&BN?!\X+4+ U7TC&$V1'S
P>>6QA(*  =W-K$YKR-_JA3V'L3\B'JBT-Z5$S>:=:A%J1(%3CP*=@/IP2"%7LM'5
PB ]V).!4*Q(:Q2B I N[!P<W'#+_HM+?,/Q?(F)@5J;LZ2"C_#W6,QC8D*,6@KL9
P+ES\]0=J9ZF,9,+\>4*4:)/M1Z8K]>$9T&58/;+X,-X WK(""U7':LOI2#JJ?_;#
P& 0Y/>G]&,Y\^" SO/L)1(:4X\U%8P,/;N$&!J!O[JYL7Z=N6((<@'1'>33T_UT>
PFI-P%G*@0\<(B+.]:O!3,<D^+W72<E\AI6;7*KQL?PKTP7'VBW1SGB2KM4.P5)12
P6^,N+P@JVYX#7-Z,N05O.XW6?2A8TNA^0?P+UQ)I5?12Q$?A2'$PXFQ>27(4HL.T
PLY6/[DN4)(=@&Q'DX_4@Z0G@'X1:?]/[GNR""VH>NAV-0:)*69"K!:%S*>WC[ 8'
P05?V\'9CWSIRIHV8KM%PW%\4(_ 7T79O8]6,P'FRPJ#K"%.Q!X1%W@*U^Z_2H=14
PD&[X_LK+IP"A8T#K5CAMXXJ5TD? P,.H8?MQ+. UY<B#0PQ"/MBDM079W5U%HT)@
PJ&$XPE:<GCSL5"/3#I0VPQ2YNB1CKL?P6@U*8=@X%4#@57P-N"D)%ZZX%=SB+R?S
P'^8DE]EKPD#T1<X[S TV.*+IV"3C3Y$G 4)UINON#-1CKF6NL"2-$@#U_.LMT)K?
P@4' ";%[2?M=DB;+W/)'[$<Q[(CC>%+HK2@$5S!OOJZ!%-AGS,K9P5(.Q&-CQNQH
P[Y[0])I<HN[7C+JK4VC;I+FHN#-OI)V-D>U:MS7O>]&V)0!JI7CD+=LR=\$ 91BU
PD8ZOD<'<@9<\ 18@ Q=HKI'^[Y=!S50>>H!;LI<!9,80\&A++SD8MRJAMW2=Z!>&
PV)O!;SMZ2^?#UPBCLK51[D=_B>#<+JL#O+GO$&L=T%0+),ZZ1DU.9YTPTVYU8<&\
P;P\S!+)1YRQ[U/?.WK%G+WR<D!P;_,=<C=^$^>!H5OT$F  ;GGE(H8$*</VPJ(\C
P/=!@-'UCHM=)VZK8>E*ZE#;Q>6DI(@6QC44)[M;+J^@J-X_"]2[9)XI;(N<*?; A
PZF,/)^<+Y6TTC6P;@Q-KKI?VN 3XD?PTY;H6(=/^J^ 3!M.$4XVG%?W0$3>B[(.C
P.H"!4@C%HS^&*B+E/G5P[/]%:I]BL^,1I@^TC4PY4)#K/QF=>,MMB%W0;HK51 _(
PL%[T,C0\XE'.PB->II1[3J5G&RUD_?33&V ()6ZMU"U75"#<539GH8:Z,,RH^/]3
P3,W$7XEG[BO@G$V"_+%^!D2(2+[P@=;K1JB7;//'62[B^-]E%2!1X1YD0]PZ8E&&
P^J0&J5G8T+\?+^7&<S.'-ZTO!.PUIA7/ZKLI/9#M@R<HC8L#*[ %DRRJFYYB >KC
P%W>_UR=>"\YH\*Z2ZGLE)5H9IH-CO(XQ64 P#VPC'6E/BOKG !:RI8 \=ROH1Z1I
PE&AC% /7AJ9!D_H-'5V)T$U?SC4+L7FB8S-BKE:/D,4[HBW"Z7K"F!B^<TDW;!B.
P5KJU$0<AITT[;=F=)0; W$W:$1A'[L_FM+4K>@=OS5PYW7#9I1\4._\]4OI0%YAG
P>,^L1_25O+EEN1R!;OH?FN@X:^PMS<8<S?@>0PTOQI5NR9K@,MW?R^:Z.X!%UY'6
P^3DO(A[O_6*W19 Y-ATY9X^HE!A#JW?(^8G%'CV83Z[;8R[$JE-3TSR-:;@4]*$0
P*!4T+CG [RYI^E#-1AR -#;BOL+E\[ 8X7:;9C@%(&@CS(ZC=0[S-JY.9WS+JJ#W
P-L6& \'&@.4*FO*BE?B-GFS!L*T6-B1G@QO?II :7,X'<T5I$AFF9UQ^:/[L^#2?
P[A[S)7<CO])$C01DF-8;>9FZ$7.R/7LLLDA9#BG7 'E5_AN '^UG>T+ ZZ'<V%?"
PL6QDW[6JMLB5^$SS(QKPF31E%T[O0D00.N)B3I_V#LM"  %%%FK,?'F^'K@,]S,+
P0%D"O#$W,K1]#'E1;>"AV#/Z?/.@W+_5#ZG/>FWON&*_\/<?:0<@B;*HD\\)BXZ[
PN*=.*-"C?#%:Y$V'<:99^F.)1Y'6B6'^*Q[GH$ZOVBSA_.4G6F+KH\8*8IM"%..R
PVH*%R#L QG) S$!RL?GFN1;[76]!(!ST2Y84TZ8<3'6/KE!FI)"&>%^H "4,P;=:
P")A",6D->]^2C?;C:9?BI)0B/LZK:,D3=G>293U'W<0UV>J\$2]OZ!X)-L$+8VJ3
P?KJY-W"']OY#GI=ZE@*WA\QLQ>-X=QLF T-P +2<D=KCD?6?YL"5F(P:(H%XK+K'
P:N0DXHR%-^L)1>M@ETN%[843$AGP-O_N#C@/%$ '0HWFS@P2*&JXPG5G9.)5T/OZ
P\Z-!NI1Y@ EF9XU1O+AU,9-L1G5\!_NBX"&6'E-\PDL1@4%"3A*!1P43]=R9OS+#
P'NF'6=U3SQ?O%^#$W/2P' *Y,; $]!7&@H[H_>5R3=C^C^$\K+SK_0[9>^9"FBTM
PP[EPMKQ,W+=#&=AABJ?$*X+CWW81MC.D>"Z&:81A:5<I#Z ^.6_1MA^G0&0^YEHC
P &WR_^,@.=.;=[!U_!4\7TB$7/_0<NGIFEP_XG> 3\62KC[C(9J\MQBUD$"-@S/N
P\Z.T6U96M8ARZ4(+EX#=GV2+ )W.L -AR8DP.T*J0=Z*JI@UE@C+^&%@;+1K/Z?<
PX>I(;JY]EV9;)X,B>="""5[%T.AD:'JWZ A#[4.2Z#Y2;<9X&&?/"Z@OB61"%0G/
P>//#FQ' *ORXVRE#]:I%W0H.3*N;74)&HAN//!G-FYH#2&ON/^T<5P^2W]^6(&\ 
P"G<,O#120"/C#8'A'H!\7GGBR+YQ1=3$#'&>NH]IO*/K$F$6T:FW5((**DS D3M*
PN7:QMA5;%0!;?=B6[%H!F+CG58",7+[S-MU3A7P5HT?)QYR+T4"ES:,ME+"58ASR
PHPP!:CP,Z_FDG.6)?JD=#_$P-]G*T6I;^(C]7T2JB#QDD^(OF9#6)KS^U6( '\K;
PP#E:B@QK-_,G26JL!B_N) Y<'DZ"AT?FWDO[!?Q&U68G.$14!^]\-LXV;X A0GA+
PX!"X%VE<F85<DA3847N.OVP1^-J<AY;@Z8Y2:PC+6%<*/%!1^(HK"Z8T@-4E]!#C
P6-GV?+RC'G(0SXIWS^%"E[.Q'*[C+D15;'IK-!^O&S>M%7EDNYBU+CCE9*TY8/<)
PWCNUF4>5TIU6:?;;V/Q2&O"WOI:)+'Q%Y#Y"/_E_2?%A3 7YUA[TF2.H(]N&ZWLP
PRV7QA2R)5OFB(;?[ 3_MT0"F GU/%0D-(/=&1[!L<(%+MUZ!#'"05NZY+HO9D.IG
P8]X5S)*#N$&(F[5_6.^C>M -L20#/U:77TQP@<A5)J(4[[;+I@E2:<7DE-7VM2M[
P47-]"RD""KZ?6LC1<#V@J8D70XTY\M<PZTSK]1\ C#0KN#\YYY9P'S3,T4;$6J/6
P& +>7V&:&V/G&W"(CX6/KU?5-D^._,#U?K3<8Q4C'[;?-?Q-XO-9F"25\ 2.FB_\
P(RY3'8<5E=%.]H]IOQ9/SMPHW:KAHY)LSV6F-%F/T,]U7&8Z-T(<"PWZ\/H34Z&J
P4;E9YON@:+/+:="#_?%E2<JO2+LGSBY4[X]FE<O=C6F8H'-,"3X:[&+*=9)Y4F2]
P4%-V1$DIG5; DT9BE8.;4A$_C S1JCGW_^!*D7+AZ;5#+&X,L*DH1HGEV"]/L&VI
P>Z^P7OI4%<P*6**X5LY!EF7L-/>TA+&C2,<: \^3['6RGV IAV6+?+QOO)A)W(,8
P,*R,BDV\M/H,34["!CK_MOT+R7 -5"3W>FI71_\A.5X\7*+ULGJ9TO8XIS/(U"ED
PO7$'%9/GVS((3^[^%GAY?='B(*?)>[.%/*KK%/5![6?9%ZZNZZSK),?HEM;$M[L4
PO#&=2]A/M_?OLL^2>0E[^32+/0MCPR9%&Z0"<_[33[04UK[R'M(]D5\V&A('3"[C
PW^"KI^6Y1(GK<,_ECI'?IQ0FR4T5]NXI;H4 X58<NU6IZA1X(*=Z@"W?^3RRI9],
PW*57GNF"H\T]NU!=[FH^G5072G;AMDM7;2OU*LC<Q \Z)K5H2*EO!KQFPR)8+I?2
P1H"_KDN#I6,!NPQV495KE3_,OPS>4 /F+"OWCV"Z;&7)4^$'1L-?DE!N/+U;GK?,
PWO24\]>IIG6-XXI,UJPB+C)2K#<//) Z;\GR59'7!0NV8-'N'/%=B@0^.F)G)/9?
P@).(K$7<D4IJ$I?,(65U5$&6'U39\1CU+_F$1A&KAF%N'C'QV**U<-AH?=JQ5 9P
P$(W:P7 _L5P(GD41J JN#?R M#D==ATPJ^O4R#:;$]![;5' .D"W-U'%^I<8)YO\
PX33[CRCAZR[_Q&NP%EN=029^KU[\5@7I$IV*:2_^\:4>$%PW_7Z88XT:]2FJM'(+
P3&H*#Q!?,*#V60XL$K]EL-INCF"<T^MM;28!6+@ZOXOKW&:&:#ZH0<(+LU"Q,LB<
PNMC>'GW42*MMC/HBW5YW,R0S-O5<W+6B'ZQF9%2/89Q E/Z<THVB4VV067,!V#P"
PUYJ.IRB @G'U?M]P:R7&^\2#*>V-=H.'@89R%IILY"$#?S,/0M9Y[<!/D1'EVT=/
P2KZ*T0Z\]6V30_ED^E:4'/)72UTY+O5$#.P3 ;0-]G*)753?$G 2HY",AKD![1>2
P>>R_DX7H(S[2'0SAZ0YGT#,-^/E\?(=6?K$_$AW=]%T\J =H]?[>F^Z-.8B/]"X'
P!#Z'@'OSTHK."W-B%6.D'78\$N?_S;,!!BTT\,NU,[+VSPIXCA5D % L6CXS>3\3
P58NN '6Z3P83LGC_6M"=>&U;<6@KUSF=AC?TB.;$80>,8\BM-;ORLUP+YQJ/,UK6
P5TO0YO.5%H)P M$:;:-.<*DRJX]?:A)EY\EM,R'A>V@T;0PAA$YP.T]^6VJ>?P<<
PTCN(<A9O(=J%5[ADP.G?"_4'\^VW+)^0^R1^4K6Z5+VW>PAW0<991>->MS=.#_G8
P;&<AJV>J_KDSQ:XS[\X4!E4/8R)ES"[QB&&5\N9YJZI[3.?YW.RT_PK4,$;9-<4(
P"&.SJSCC6Q.+,]5Y(AZG_XMD1]759R2Q=H>+3VP.7M<_N+CF$6!$:TMGADBGBW,:
P:.9)B60^-HC5>X8":S92BXN4^\,2;2@^SBZ.G3%NPA,V)PNGP$M870=1#V1=+#(;
PZBPFJ_F7J2A#>[\Z7+G[2$:2"KB,D'@2E5 JS-!E);&-94'ZW%@I%^*A= [DI(]0
P+C[U;Q#U->-5W:N-ZE !=20 $,<#LV($Y_:QJ'ZUH#Q-F7RO7<"HBF+031Y;,L;\
PQ6N4-1Z"?LY>8*[5\L4CE4+^O\_=BZQ*?,UMB&+3WENY>WP9JO02LML-]C\#'4O=
P-PQ:(0)#5E/&%*F94Q^A7%1_/5?:Z[R(9E!>9IM)@Z#AGCW!+0;$/5[\;H)FP+Q,
PO!0]O-3[D/I4-IAV&MC&\8/PVKC&.E=DPO.4()PGWQ6!*X$HZU1^J?@=QCYE5W09
PZK;M> @D-[:*&!5[99'HE+&YUP>^H4]_1F%HL3]8$/4R.+2+YUQJF=5C>;Z/.(0S
PDXYYAL.S[\1&F5,O= [/R\'>K%<H?VMM50Q;76!0(I;%TNLP@+VQLN16@HZO_+EJ
PCAWQD1Q _,,BU;6#UPU#Y,/=5;3@L)DD,M0M![M%4:NS9WSY 17#[<P0OGKNY7]O
PXI]WN#!18L2*R+9P "_]C120*5EP)V F45$&EODS];WR[7$8B$ OC,Z3F"/]-Y D
P&BIIXJCANY$.G#V(Q1CG82"?$)X&V]OX\/$\7<ABW!*Y@)O.^9I,N7U>#Y$J1T9T
PZD"K2%%D\#'"N6YF?/?DKP3&]0G$F@6KI_QNEH=49"KG44W)CS.K@,D%Z2[4&-L%
PL]<Q"MR/2H6G?_6,)Y*P#\$F_&Y2_HTR#XA 8XO..9L\H;N6=_AL$L(T;##HDA<O
P@9@.8A%33V_JAC1*8<JFHR,7)[T<JL?OHRD@3K.M)M'68Y1'DP*PE 6W;_X,(BE:
PT?3Z12CXF&6QX$9/[]L9T/X)=!=79-2S^QF-:;LRE/OS:PW%;B04;%[#[TXMX6H_
P^9IR+\(YQ!P-2ONDBXD$_ E\_:^X:',WU23H7JXHM%/(9;U@')6?R]-J&$:E?^TT
PB9>]AHYB55DA"C$_=CV2SB AG9IK)O),K'4PM@8\[+!0LBSC3U=I ]YO/V!4KBV 
P<JK8/(2(FXC"7D[7,N'EB228<%/OK4B;ALS51$WEWM3;5NO0/NP'MT^#T4599>D0
PI@DCGES?6R*<NEG<HZKDO.0=6?,*)%3XV91VP3:[_P+29<1R FWL^U27:UCPEQ.1
P=>NUJ\H >$*SC!B.UW@)D)>U37UU[+NLYGAU>SQG^$ K/(VKL L 3?UIF'C]2FA4
PGF;!Z*#C$G3UM>E0[AV(=%D71?MH1\T=Y^L$M7V9)JUR.IHG%CKF1WPE]#%BIHF%
P$6#*NE"M:TR/8/WT-73-Y^)/VSN1?*Q;;T*JS/.!"6TGN"8Q?.M"UDDI,WAKW7.X
PYQO?6Z3KO E_D_:3[Q,K9.526-_[Y"MNSS>M XPC)H8&FG:%VWRX.L#FR\J;LLCJ
P_$+]OY.]1UM\UWYZ).WUXV%W3@Z]PBR/?5DQ2>_#1/S'=%'#4:FJ# =Z$OAL6[[@
P0U9.R/EFJRD6C3%\U 7M+.*'IFCR;6Y:3[T8\*N%64_1*W(N-8L54$!]_$IF5^*C
P+4D&O)VX0D6<O6G+<0R09NPH5PX7.TJ.SRAMZ'C7'2 \1SRG\]U#BL(Q4I8^."M4
P/:,_AX=&")D?.)?9?C4P&Y2H3191#_%BJ8;6O\<)=/A$+.ED$@^4RF\)&O>$I=]Q
P-AC;NL^F=("S60<_%X=NI3?PNR ]Z\J('!-="/I<)ZDL'KJP=L\&4!;-3[$W 12@
P%C"0. >R8:-S]D0%;YSTG WYC.LVT,)C=% X!N[&ON''0_4^7R<9F(V=#@-('$US
P"GJ+,#:ZK6G+/T1 >)7 J/^L%1H*\.I[XOWW8P&?0+=_*ZZ99;$S+1J?VJ73)JIC
P3;:96!V@$36 K4RGD#(C&0OL[.U/O0Q S>63R3RH7FT[;NJ^,''%G+<U2(WAJ( <
P3FH?H*E&^6?'<\E$G,+0_KX@KLV KQ!O$%L1A*O>[6I#O#I9X1?T@'< \^Y]!=UE
P=P_X/!DF&RB+;U)^+'MPJ;PN>#\?2XG?R.88N9MS^=!1-=(F_F]0%FI;'J*@<&$K
P#CU ,X@:P_7:CCAH7"KC35>S*NV8!?EX<>=^?F?2'VCS.8/ 3#,_Y&I<JS[(;7.\
P_,=JK-6'059;D;&K7T/^?5&]E=:*^HMU%'C#I\[*7.0)PY[")";-?233_<->=@&H
PEJ<AIAG]BJX]Y-5I">.&%)!V%S<Q,JZ!E>KHUIG5AT\Z0U."/>5>,D3YY(,Z70?Z
P"F8?'ZNX6"S(8(0WW$S&?I7C T<XY<E_Y&+D.$FTO49^<B5(WV[_<(MYRN4-F56N
P[I"M*;PO@(_GIJ6C((,I?U$<P;^I!F0I&]'9N$W*/%@$X2,UB5ZX).W>BLI3^'B.
PM$\C=W&AT!F%PO8?3RZZM_ZN?+(33Y/!%&NVTN@Z(W"NX%JB!1K!\R$>A-99>-VQ
P7MEP=7I^ECE$@KTX^ZS-CMP='MV"D.8G<0)9,R,J[>W."G3"B/?]7PK((3UZL\TH
P[Q,;])K_/'U21'^BLW(7 XE:26Z$.FEYQ8*Q#U4J)[=[M U4+J&X<A/(*M,S*W4'
P+]SF*T%5(+ SR\:T6W)T<%HCR]--^PFM&=ZBMU]Q>DC&+76P,7JWR8))9D.S&9!E
P'/@9E5*9U\6=BJD'SQAQMV9YI.TW&C_NA\]C--* 7EK%\?&.BS68'697K*7Q%VNS
P5D#F %%A_0W2B4OS0GEZH9<<DD&2UAI4&DF?2H]+"N+2@DF 3+8;4<12^HM>?KQQ
P@A86BG!M-X?KVN_;,-<:NE[-;,5;SA^3L9-A^CV\A:IH!P3>%CDYK$HFCW\.>+I:
P43.<!KF5Z:H%"DL ,"-,74D+_G=4;C+))'"Q1][IO&*U5LQ_^@MM__A*DE91R9#M
P4-\"1P6*08(6#$__#%$=3T=OH0*8_;QE_('E-T)&-M([I[<LR;XWB"T&Z1-2JTL#
P<"7-,<WTE\GA_-9*MM\@HG4VVZ>QG><MU-;Q18--YJQR,!>W4\5O8EO6@3UI#7&-
P<%*X^U)Z0QY;IS=1TR=J@FD &NJPQG"6%QS2%<D$TZ;.4MCT6*B8KDB9;F>!5-G.
PIS#!K \:$%E&R:XO!-O_.LF2J5A_K9#P=AH0JA@PVL;,49)&C(-&('T13!/*/K10
PSO[9Z'4:#D!/4-P0'A&[<E3G06M*HM0A[W%T5< ,X9 P @7TO"8%7*<[0OZ9TUV^
P94"=E7.J#$-3/^LA-M$F&UN AF5!3UZD%O5A-?^G $SPZK[\; KQ0+9.O\8;_O)0
P-6#L4:4>U[ZWK%S"XB.KLIL9$E;(_'A57T<X'2VCUDW/*U/D!(S$AA5L]VITGX2C
P_O.F%>E PRBQZ33=US7@G\&F_,.@G+AK3 X$KN5:.4SJ DN93.VK*43)56_JCRSF
PNN.\$I5B*)_&VM<L7@^RP#(;'#+A_E#01HO^,!>-9619Y&7#KN@5E\%8[Y?=5JI/
P,%L,(]IN.:%#)C#,- 0+R[@L9J6_+YSIVUBSO:'E._09][Y(H(UH2>FI%1*B0<BS
P('+%N$Z)_&R>F^K1V?D)G=0]-/UCX>H.H)S0RZM\\$;1H"/D:[7ABU\H!YO7^<X@
PM6U8)$:Q,USZ:N5W.22@DW_0<=X:FA<^*RK,U%Z(,\Y4]DS;50A1L:(?33;35Z3T
PA2EMYWSUXW+1!-WHXFE#:S/'-":93V9(\K 8,!I(7X=B><H41HSX"&D##_OB;PG3
P1Y:PSH=68O9D<XK@NZG1J),FA'+%;.>E$_.DY6KLR_8\C\IUZUB6:,6M9706-9<'
PP/*Y-._8WOU?XY*M1K'/]B45#9;>"!Y/'F,7JK(NVW5C*\5(V7\OCO6<UZ&JBGH5
P ?)J3ZZMJ=(^<A>X$:4/SN3S81D<=^.QT3NT<I5Z]###K8Z2 ;.XN*X,$@ L<24@
PNP=>ZI\IN!*S'>J8U0DM6CIQ+CU339%"V T$\3^EU!T;X7_EI>-?[4\)BTW+^<;D
P+H.D7PH'8)Z9PC)$"D#;EACW."'A]_[_1AU]2GIR@(F)>G.\\1E\JK\R67VK2#3+
PV(MF_[*(#>I83C$E_[,J+<DR?3T*I^5@.$L_9?V3/E!XR;.A7Z+8_@Y0.-NF._D(
P&2P/S6++4#W/HM?;@,J%1B.')G5Z/3P))>.,^/B2#^;TW0U,*KZ5TED;R7@Q0JHG
PF]B$C$-G+"M'I4F;>$RCX#\.8="VBG.<B^2"RR[P0#/>R6Z\A<*[H!4W.>(X-URE
PR%%DD4[5;;I+M>=N-.14ZD=I X[)O;*PSNER)]SXK=<KIN[.C$F^+ A[I\<8E-4*
P!^G86+;>"/JPANW,8*IFC.Q#-H-8QG)/'H&\T#G:^=T8 +L;6J]1RZ@]BWF2XHX$
P&$&5.W'E9/;H03#D9MB. Y!&()6BA)ZIB];][$6VMFLT"1P!3-9KGXZ;Z^8 W'<"
P@DSGMU YS9['V :"[7L&UH731%P=VZ!6- _<EUT>,LZZ]_V&AW_&*?1\&:D;[6C*
P1K&EAOW>1T41=Z,GA+Z&&PVF.A& ^2!4M,DG^;H4G)R.EK\M@%2YSJ2=J\7NOFX6
P5W]PTV:#R?FY[R%+L&X3 ("WNBEH=_ 6 QS(?V<& #W)!BQG)*-?J]]L_"3):%P"
P-)T_:*CP50I D!%G 'C#R;V&<%Y6/^4B06^*:2/G<N3%E<+& ME7<633W2A)>')7
PJZTE6O]-Z<VO")P:3[-@Y&U@6G> I*<12_U=;W,L_8%ZK3B@MY-]IYO+UXR5)<1U
P_I3(RY8N=<T>)\5<$?7VW$F>WG==7/2%@[4'N UXEJ&@V^)JYEW&.1HS]EOZ(K"6
P+7>!UJPSHBP-67U$BB+(S4.9ZA9NKX+]YOZ@Y7GC\(GA*=%RT<GGB[!3++%<1\P-
P1/WLA2C+6T8.D\GR'6^^V8*C,1[Y^C/!_Y5*7T<,\H-AZNXB$<>GH2;FYC[ZZ]W%
PT$C3D 7?XBC8H"H9V17#I]0=WFI<2J6V^U<&,.I@;N?73M\X?;-@C'3\)TRG%6YF
P^KO)$-IR)7%;C^=&13Q>G/%TY($,TKRAXC77,72EPRC@H9W+@WJ@G";I[IZTU'37
PB ,%-T@<G=.OJFMU46@(U?9@/=#$:D@ TSG"2H[E+>:CH<G>>0%:?K!S!8.ZHP?_
P7*B2^!STBAL?F"L!D!22S&H(B'4![SS&T;%^,]C7A60_2%M>DY[ZOB94F/ LBNR-
P,B7<9A"[C*5]I!U* <U1[=G*KYXPZP1P?_Y%%V,/%V(6BFE[%U$'A6T]N9O$1K<2
PV-=IY6C@>5G8BN+97OX;#_L4,Y U3 0B0@PF7\<K-7 >"5PF W[O^F7-O90*GW72
P2D(OSQ2?=S+U('EM*\7#^_Q0WBX@TVCV@LXH\\3'N )0&XY0/2 3^)O1TG72H2N>
P1#$;6Z-4<7",E'<IJ#;2&SWCOG]%WCI+\PE"[YA5J&;XW4IX_ @U[[\KI"O._S7!
P@77P6_"GZ=XME)]0/*4H4,3]2""I3G[GX!0U YXGM<@';T-5:RY;(' )O%-5Z45\
PD,[VX7@Y4>7WO5BYHX>$)GKW9@I:E2-11B3&)PA;G.IV4KTOGTN =*P=>7C'CV/@
PZOX,#@[G8@F>FD&])_6!6J7JYC:)([47 C*K3(K",#9@S]X,SP#!L;FOQ2%24D<5
P'RZJMY&X>C10ZOVH/E!BV-A_JF](H(F X_('OJ!\#.+>+5?G* 2:)R(D1>SC[?T=
P"$D?*(2%8U@M$X^Z7U_DX$PI7%#S;?[W212B!5F\EV)^MXL..V:7]L)-RYH;F7)-
P@5?M$ &]"RE!-:\HV01C Y$ J9'$B"KM]M6=^V =7+=4=R[)X._U>*OO2PIL(>>!
P[W1/')D,*!JL!86!^V'[,CY!BT(V?>:S9@\(^' 3G4\=$3L!R8F1&BX\3B6&,U0F
P)5T&#CAJ*3#'>(ZSA4]]C(!NK>YP)R<8F12M/$LH%&9"Y-AL\2Y \!;0VITK)'O\
PCXJ0\#:K&/?\X"*<+'5"HD,,<TK[+N$MC(4F4KE,+)T_]3GPS#JSQ-DC M#5NU>]
PR!;B;7-H[% W;-XC$EL%K41\H-RQ(,)D8!NE73.O4%J7\#R=+NWC+P44AE)2@#O>
P/" 0>O1_)!?&U?C33KKK7F. ?;\EY3UC0NYJ)!R>'OSBM)L53)/+@BNE45^EC@ZV
P2KHR,'V/9G"6:QT==[?U1XK2P1F\,U3&3X++UWMSIA1E\^X6CA'P]"84+Z:@+7%^
P?\\1I15>M^7!!R)$MLJ6!7&K;WK$%X;4<D1TN4'T-JI((49ZZRED:-MTQK'5SLI9
P:;Z3K57UFO#B+;/%(N?S=(4K],X$VWYE!YLMF9DE;N@NMAX"U1)"^LN+)S\#K6VT
P_*+LROH3TP'\<N@N@L.K&R&!ZG#_;>?'?IS##TU>:+82$67>\(@[.;"7WJ,BW)_-
PZK%VL1@?<SX7-R#X8E1!O<8ID))#U(=Z@;W3+3&V_]QQ/5C>CJL25HPV4*\),:T5
P&TN'*Q6N[$,>X]F!5%_IQ%M?R26A+V(V(%(12<J.?-!WHV+DC)7XTD*A\J3M/9FF
PKK*0OON9,^Z]%F/:'GY,27NKS JC'*VQ*/FF?T*G*QK5?77_^';L_'%-RT I)18*
P#%E"*P !!S.R(E"Q-,C>F\3<^S-6%)))R13_TM:7E61Z(<82UY%ISCB4BKG!J)#C
PZ=U@3GH =8*&XOETM(J3AVA>1B5-TGQCF &JK_I>N^3"^\N",H(%JT7K' T@YY"_
P[VUG%O=A:446*)G2E#@>'VP6\='LG5_'-\NQE)*7!GA@\+:#C*.BITWR^Y3FW>Y]
PGE?9N67D9Q@B30=O>=4LT7ZE>U)KII51E-V>6Y?487^29'!4+R_D#@L >/2GE=;#
P)VUMH(.C[@FEP9/Z9)05\#AG($P]V,NJ4UH7+J#:^\LZ.X(YC)D#LO=AED0%P[U7
PFQSE8A"<[7_W1+"*!8&;'@'@2! H=XV!XK@K-M"%L)O:<4?Y(R92=2 ^+U<L]P&3
PT%8?C#?=(X:&CK@EU13C[%D(&;3N""]B!^E #KHBX?5A%^@^.+D<UB]$M0Y^/TFK
PNJD\KF\(24LR%PQ^_RW*6*K]?WFM)8?D2GGOD+2-!4_2QCKH+ODY_>&HHA&4DJ[#
P,M5/7[Y5Z F+9PU97F]F/T&=\96^S%6\6Y2K&VPM=B_OK<]6XS2Z*VI98($8^L[/
P;M=._,@KYBJSX\^^=1-S&4IU&&7ZO??+.N.G\.W\3M?D6_*"3F="LP3Z_F$38Q3J
P#C,?XD,2B-"-.KSFD/$"O8\EFZ"0HPOO+74?TZ(&KE4L1-/]ZDW?K__9H&Y7NKV3
PD%B2HK%V;.FSDOD5!Y%W]?K@S&8%@"8"$!(BCR ^3Q#]EZ@J<]QNM>IK0H2YM2;Y
P\"&W5#P-0^//@IYKI[O8'Y4.']H\DM^G,U_:K/M]C8E?_IU5MNS)>ET"T&#_L2K7
PYV*$HY8S7O.<\UM>$Q_5UH-4@<&H\?&3*J]%H^IDT_UW(TTX8>[CD&LG]I0J"-9S
PHXP6I> ##_.ZTP8^.<I];BVZW]25C\"+!N4-<(>$\74>0O%7AS@@S5\-#6;"L(JC
PI9YZ7U'[B__-UYN6^5L$V'+]'FC[04?WK*ZK("WRC4]G6*N:2[LUQ.0@\KX?>R'^
P/"B/\)F[MP7?F9_)JL>B6!EFK'45M\][J&(.]*$D+?2 @J[-.>:8J 3YV V?]V[D
P)=*#/'01X@.#RO92A(ZF?&"8/QI9 G&U83T]6^$1Z4)28\N?%U(>D(F'ER^ZZ+G[
P2F'CZLKJCW.!Q_^0%[%UTK\'PBK8_Z@\WMF@D[M8?QB74N?X4)A/?:4CL(5N,W!0
PSN(-VDBV^3$P(2N3.V&>Y[&UZ3^.EIV#5;RM0<*[6;HJ%7H V6Y5V*V_RM!7U[%M
PI^(!<LO;]*>F#KY3-L_'5._O-^3E*/KKZ/L_49THN<6ZGT?Q4OCZ+ZLN*&0PC7%F
PI%$6F(\TR(9_TZLSU2GTV[@&Q_N'1S[X\#;$6W]N(DA1#9#2\VT9@8NL"]$-XS%F
P*DC/(I7)=VON?BWQTGJU'SF^G[41BD3)7_$YJL,O"B?7M!?0<5@N28%/+F7</8?T
PVYRL2&#U*_#'-H UMA%%FF)!OL;TAC1JU-#,$*6J!TC]&T^_[]R[_W.GJ@>PT'+7
P= <'?!)3AF)>L) 8B9V_A/1#9QH(E7@,-OO*JAO8M><$F[Q^%;E9W<".,X)2!(Y\
P!EB9>+:/HKA*F>2DW R7[!(@+?J$AZ\4)Y^" 2;VF,>Y%&V2MUY*F'YH -O@[ 76
P?8O5>TFH&92]6^=B)7C3-^6+5($QW!K#.@J>_]NSK@0EA?B,U=S4+0!989D!;^P0
P24EF&UY\,J[[EV92 GO=$J]HQN2UG@=SI2OU8.H0DJ,[KUJ05=/4Z6HL(19Y%.M4
P,Z/?C7@3"?:E<"&.\C2=]1<9$RJ+]%VO^-<>CEI",>\?_XR8S'X_7Z[#E+X$X_C,
P=VXUJR#+GR>Q[(/>7$9E\S=W5/3]Q"BYT['?^OTQ=*],*8],7F- /J."^8N**9J*
P'[ZER+ #V\L,]F,YF;^;ONMMPE]>.]O9 <41NK C@)_CMZ]SI@2>(J/YB4YJ'X1I
P=(23U.@0HY;)@Q^D55-O^=!K:/(2;;HO6O("IF3TTF3Q>[2=5IFVF5>M>6! N=^$
P;FH+=6ZB<L!9.RQGQ13(/:D3CMZ!*OB CY_-J3R#I0(._ (B,[5; <C#A#6L"2.%
P/G$/1.JBTJ?@!&0 N#0IC"! Y06M.AYA%4A=@K13TZB X+I-B%#PU"RZ @XD4["_
P+"8&3':\O&[V@I1_4D><LLS'[6MS;_ ^5#A,O5834:BWOIB7Y!/"*+V%F3%'5SQ7
P<<F^02BU?F_1?6) )5(\$5)I]N.]XV!F.\V/S8&YM\Z,C[4+/^;)J];<R^1;LG;P
P_G#G??7:++M7J')"B0UW8QN"E>,=>8'RV]ZKG"U/@3(/2E;%]:[,*+4"]%"07<FB
PK,;R8G"#L+ I<YA)9&@HY1C([D/O[<;.TUYFE2&Y!D(838KK31C%W$9=6-2<RW!C
PUD;PSQ-N3OQ20,%"VB(U3-XX*1HVC/F<\<YB2:7[U4R[XOM!(AL#X_WT'CAZW*VN
P7TDKXE\7#811)*ZJ"\T.98:OHN.@+=5.OX.Q6XR3T-;PK!UE;Z9M!" 77^94Z[4O
PWD]SQIH:$Y%50JR=5YK]G-$5P.FTU@S.ZI(EC@0(=CMUM00PV_^.Q@/1&W3GT7RF
P6X8PO0?_>S"7?&7J"S,IL=N$B[U;31<S^HJ58%PZ6EJS-<J^ZI5WMW<7(RH/?,\X
PJ4)FTA;([TM(YZB7PP&D)RXSVQQ2.:(:&*OX%=><+I]NQR!"S\Q9-98N S%E0ATC
P?'C@:C&WNPOT2AGO0YO4NOOD,F-WIO:7DO@%\#YU8^L)>G2,P37!]!0PEZ58O62%
PK-CPY33O&<>N(>RMQU1/.OG:PT3%0\GQ8RPDK4,='>O]X3?Z=1()ED(&;^-53\'+
P()IWH+905I)$\*(UZR&!9VO,V1"R<@W(%;%?]!4IL-32OH%/=Q81M@O5M\6$19DC
P_R/'6T1!\I(M4:RH2IS8C%C-+SD?^R$!4Y;5E -BA/N"B&5X((JR1\D?YM9HI(#\
PI8;$#/HB7$7TDP//LW_)CI#6N2G+F&#%'%:YTOK6"PJ-L7+ABE_3]CF,'E@";UL>
PL#LK%$=FSEBQ<<V<5]MMA[)*P.U.6\G0[A<-.A&HFY""N2SPW3&J"#T TF)W')]Q
P5%=+EPA=9<1A%5:FC (QIK)(W&K,)2KO!06#H(#&E]Y1#%&RL*=,4DT5;CDY.M/:
P0A)GLSMKEY/1+E'U7;;_RM"4!S(&MY@*DZ7$?&(2;;!K*D5)HSU#Q+Q^ !J$%.LZ
PW-9G=VCA3@6C;:XY$!4@<A31$U="WI4V?T9JW6ZWW;XG;E!548['@/^XE'P[YT$\
PXK)&>H8M.N^?\KGDUZ&%K^;F #%,P[N.<[TS6C_<C$?0,%6BPKSV*@^( G_+#BJ]
PDBVNMAMFD=#A\57!+<!1U%:O+5]E;;N3QSTYYV<VA9P%K$;&E#C(/0NTU\'HM&J\
PRE8@2%28=[D55*.VS#CGAXDLTX"ZF,!G!$BR8(Z0%,BYMTCDC!1,Q8Q<J$N?H!B0
PF@D,*L15H$?P6VA@FH#[#7-7G-E-ZT-FO8!@D 'F2QQQH0F>74C*ZL6F,Y^)@JQ_
PO-N!W/&IZM:)15'/N\GTGA-9+B*WXXB0[HYR%"8B=]PW,C0=AW1?U(VC\U*:I-E\
P0S"C?=H5L="JT?-0XNV)+A\@'/ 2Y-83S7(U@>G@ )8 @8#@4\L:?U1&W?PR]<S(
PX]M7V _2 -=][5;,!FR<L?&^? X[462.&@,+^<B>K8[,SIH'*=N;0S?N_"\FV1^N
PD=)SII3VYXLT)*=6FIY I 8JY'?Z.X,0Z](&Z?0KWH0 [_IA]@8LS6<'%O^:#B5P
PZZ0QA5]0[/5U$Z;54;T5"DW0:I<\I3-@*C70^" /&@J.)*3&U[V?"2@?Q;H<Y9>D
PSJW?0$!>UQ]9]]8?6A$9C84_'V$K,-Q\%9LQ]/K;,9S9$S&O<XWG^J'^>15W[X__
PH,J1[YY?]?9%R.@STI:Q>;9^ZM_UPI&.:=XCL'3(6C*"EVU#-J< .)I@V<]3(2\>
PP>$ *W92Q4%,N:\;$_8PGUC>$0.7"<'2^[&@IP\G%)L4("H5IQ[ZB+X<K#_K_/0L
PMT1#Q=(1;J?)CUHGA@_[\N@6)XK7AZU$(-[=ENQU+Z]S'02$GXQ>3,M!E;:KSS?X
PL)6STS\>W1'QY"8YT69>2N7L9I.(:"8VA7='>NV,( 'RJB1I@+H@5(GO,)CE]4*+
P/V=ZP-)72DK2O'8N'4;1$TY&\$/;FG=46' B2!\U=*:*&.<ITB[SW\@!N%B:[@Q5
PB+@W-7T]S#GTPA$?_79SPW!Z&(3@M_N?+X".?GN3G_@2I'"H/DD=[+VID310-OOC
P-'KTJ(TI7./N76V:.%Y&U3MC>QIZG8_$J4#L6O>E[[0$FO:-TV(K?;7PIYVY,1F.
PV![%KVQ7(W-/ QN>O3A39M(+*G8&:R 700'8CL'UF9WAK.OI[7'CU<OSH6<9JJ?L
P[S1-/+P!B"?(\N\_*@&3E8,14<!ANU>%QC)NI-V_]MEYRSW;8D#0^C:]P8\2^L&6
P1Z[=YJ"\=G:3+R"G\XHU3=FI!BQCY,P0^=,5BPDIM%QL\\$(SEF\HC;%_VX-^$ T
PJR6EQD(FM(QHR)@J-L&"8A13\UNM'72!@0976FL2G"5R)%X2J%D+_"7IT'R8/ YX
P ;N_TQ]6$?>]M'+ 6>W6,\U/SQ:BTFWBXRI0'7E%8\3=]U!3R8P-<@@GX0JE*U)B
PS+X0 (SI+B_>H2 H5^:EITXC%HSS)^@V^'[U,Q-2$P4#OLF+P-C MH-AI]T ^["7
P95SN6,Z%&K(A46S7^(R3X-=^;:\=?'BBO%)&L1^$5_4G<]X>;E#GQ0H%JP"/0(FQ
PKCI;[73NDH$2V(7#XOX,S:MJRJD#AY.,8-<)K\%6.Q0@4Q,?Q11-0<N3> \S>U/T
P)./F0#3#R%U"0RT&NY^2&)1TNC3>VG[/ )>P\N^U:?_=A,<GFGMLYP_,L)S*;>#B
P67XK &\AO )F$F>?$#T-JI?81C )%&K/7%SG6%;HJX#7UNX;21)X(=E4L)'$'2RI
PZ]C1U\N.><F\VG)YGQV<R"H_EDY8(A<RM#KE&,I&N .:VCF%#-5/&?>W-GD*W/[+
P#J4[Y4Y19;91V48#H%R+*"^:$&P#&)Z*Q\^0B #%AAE-AN&SJSD]U'1E4199;)$G
PB0MD76.._-R)WD*P%*)S:KFS)D]@J*$+I>0=8/M;?^79:7+MR*MZSGXJ]*5YU-!T
PB"W*] ), >\ZHUNR;?7=*B$6 SH/VT#Q24\!0$.?5.'Q;O%Q)5LV'-,;M;9KB!)_
P'_1$GD1\1KJP#+2XU3''=TJ&QVD-"5QPW/W*R7M<[5=:M5P+2<.DLNGPZR1;.*W]
P5BK7OCH7] I4_2)G!NM[A#D*3MWZ;N@Z0-X3S$<A;F)/0F_YECF?/AID:OF-"Z*W
PZM.>HP9C^<2]Y4P\R-E3((!-G_/3#23N^09OWI8?CC2$?YCA H=\LU3*UWLO3D?S
P6)F^?@.9KH2S_$L[M=:KTP@_:O\>?/L1\/:C(3;A=+^8X22_"):X;?"9R;;&C(/M
PBIWPZ.PW_5=*0HA!&:;7!37+)]=?HX*D?!8=$PP2L?U[0?E4X\9,Z:7L=K2&"F#H
P<"<"M_)@*C!,U.AHQ/""DCB#G_HR%9/JA=3"G;OIPTB74E#E#?^"&M!OUV:G7QH-
P\G"9 #G(32!-OPCMMG]+L4*UX7-#(,F#*Y=)G[(J,M4KY_X%AJPYZ0$(2Y>J"1@Z
PV^ZC#0V%'9>]/\%TV%)QA=.74+4U(%+6-U4ADU0&U!EG3Y#::#X8D@M"V6Y11&X[
P$XK1MLW&N8@UY():T%O&-ZV3B2S''1FBHC9^!7B&1D*OD9@>7@8ZH>/N+\;>,I? 
P/_2@4,4?C+4?^_G^[TNOIZ61L_GAUEEEFCF[_;9F(&5".R+@S_<X!9=IBXU>G Z7
P_"?B^98-L.$<*$7+Z;%E:2U76=6)M7.A,H(T5MOA.V30A0#&A\URL=\+HR&ITYW7
P9$BAB3"ZK=O!&]BNISG,RL0P_8M9AMNQJ:P25.J('%OD68'6W=#%L/0%8Z..!2-M
P[U#O^ZVQ7LP!<=1 -@S,\Z"V5#&,=!N(FFJ!22/7-)AQNV#^#<T[&O!-T6C'U'@^
PS]F^Z$A&Z1F5:RVM1&Z^'\H!.7RLYNK@FW"#!A"-6L\SBVPL;/!*A'PS'B'YTEVP
P;"9HEEX=5<D4:/T._JX%AS0LA>^BZALL-QS@%O(@S6'I='Q:>EO@O["/NR 7^VW;
PE'9W<U@@S^OW8-.(T8/E_$QF$"!MQ407Q,^H.H*%/OM5=K9Q/7;,V+-J!/6=U4NX
PN?1Z'@I6MFE9^^:+:UZ9E=*9'']MD (4-'@(O%$/:_@@:BV66^[M!-N$T /*!&*0
P[GQ.-]'0-5^L*(MG\GPD\QD):X _"Q_Q]>FO2%C-R!84"X41@AADQ$),4!L%\AFS
P'#S=Q%M"JAG>L4%$3F_%2DF>'_!"@X*NPJG/G$2:<!W^ZV[ WEU]0J.U:-57]V)3
P8U"]+%US/9>UQ']S&?[ 3ND>*!O"3> _!0QJT+<KBJL!QG&G?T+5X04SAV!<!+Q!
P>_Z@RA-JSBVMD88/=^&U_36[YY"PZ#&5558B@W="@1)<L&O\ HGDFYQS"9MV=4?G
PQ#CN0O+A9E<H@I4&Q.PKT>P>CXTB&!TS;W(FH;>@=0C%7KW@XGL: &YH!YA^@?)_
P=";<0J;2K4/>M<EMT"5;+&R+B21^NQ(B1\*:8"9\9Y#V\:\OU1DKQ%MOGNRO)O#R
PAM:'&)178S8_VK4B:.:+N1W?4$UH Y?3Y\C./Z J@!.&3=EHR$R\_,?\"9>\(/,6
PV.V%UM*=51!4\]Y=<C!ON:OV%3 6AVYMH$&HAFD?1M")CYR%U&EVJDYZ9(E^<IWP
PK[[J_PW2;"AC)-UZ7WD?1.!TYRD.66A0.RHKJBD/KIL1!/O?]6]+;W8I>BCKI/'3
P[(D5?#4JW<T?B=>*&OJ;V1%4_$LTJ%5I+9Z%-CK*=:W:Y(/<GCV&IQ9!C2=RN160
P.%B:>=L*!ZPOD&")+"\4^D[.5F SIZ[;W8'MC\W)*Q!HY@WC&D@L_)%]GGNX1TA$
P\YOJ"Y2:CFU"% G:]R%7 F$N[BBKCR$O8?&VR!031A3KN>)GJ\'\B90,"%FHD>;%
P9*B*>H\$VK4;U7%R/;0#JX?I-_,0Q@"?VS^NTV+-K]J_BFNJ(L5S,#[-XD7!-Q][
POYP>6%9(*7TPHL7FC'UMA-D&PL_+^$F$NGIPOU13YG!*]FV+K2Z+Y$<H3U43'C<'
P4<!("615\!%V4WA;YP<VTIJ(*.*GR^DUC$.7EOL]K_49+)&7BVO>:+H-!L[5VAP_
P)6GN%';X:1.-'L$;##(7YWE>Z3\@A]%P=SE+B (DR38NI 7$B"(VNNX7$M3BQYG4
P&T#H%OUAF6_SRL3QYV^&IEBVQ)D71V&+@TP%*1C45YQFK.E;=LK9%]L6M6UXA><1
P)^T&<:@E=-RDQE^&]\==FB&=/;<RE3BW S/E,[!B Y$?0I*NYO$*M4J5,)9Q-O?)
P)#'?H1;M[@?"# (X,*1Y;;A78M:#?\\87T3\!8Q=HP]LBD5/;Z_>\;[84V8=]RSD
P5Z]4^YIFNO%:GZZ4SM!O<>3&G8_;_K?&1H6Z/P2)(F9*E0FW]U10/U3UVLL+=**5
P6\G!VC8M.PMO@H8687$6O'DV"(.(G#5IYSJ]^P[\$6LLZ&2CL;4Z_G4;Y98\/_'$
PD_KE<.1WN**9YYA&6HO\1VI5J^;Q\I)P2?9 )KC!+)3WRIS'O#5#QX&)=V_OB<]5
PN+,8''^54;U HCUOKR)LS.1=@1&_PQ);_?1Z[R.MGG5#O,MJJ4RR\G[%X8I9(T33
PRO<A-&03KSQM9UW=,D'I%AXJ1<O>D$TQ)A;#?&Y,Q $@:2_CS<#Y)<LMHK3-;S-<
P42]4M^@- ]Q,J*<7$/$X!$3;130D4PW6YG&&-_6 \A:;<Q/LOA2BYW2+4>X+;U*M
PI8NZEQ IV#TBHRG.HY]Y2?G'A! 01ZI?=BP+%$Q^UCD\(FJ@NVT9^[:-HE$H0'7R
PYC/E92!V@U5X$P2.',VUQ'H]U[G]_<Z-VOO)F[$'YGP]-\+ 77;3OC0;%PX:Q7Y9
PS%LI1%'I)V]3?H2^82]@YDZE% K<O3;S779@V6JKI,4KL\@04K=]O>0WO++FSK)\
PXKF-68###R[(*OPDV<&B+'N PP9.Q?U*LX7JD3+KKKD;AS_W^\A+X"N9TSON6X;X
P#N;D'.S\5O?7?R*^)+2H:5$MR4)2RW?;R\L)&%[XST72QB+8P-N>*[^O<NUC;WT 
P3]QUFP!H-\POS!@7] <[?#YDF_.N]MX]^\@ZU>790H4<I"D'"VV]L5 F0\?8D&/6
P\G4)$=:;>XCTEKJ+=K?AR(-W_NW(3C0<$=("FX?WM%[!E" M:U!"^"=7M7X62MM!
P"&%M.[7)O6%I$FU)&ZAO8C/((08[15P@P%Q;,(11F<:8;QHR&"9D=X#^@TI367/(
PZUZ@<2;6^AHRH4.YJ94(1N2PPFK@ .G P3X*XOZID=<V^:<2D%=F)Q:V!F6>#K'H
P:Q8Y"937ETAVERR 8G7[09G*/B^!])Y,J<%$*(1YS9F7HKZO=C3940TUB6/$-#;7
PO+"MXKJ5_((=8 CT-[TZ3P!R?0-OD_0 D3_ 2:&,(&X7M?R!ABQ])I3BL]^_EP+C
PZ=/!3-*GB8Y/>["Q#SE4*MW-@K-\EZP1IJP5S[6UW/^FLLG5T%N:.""&&5!X:XS5
PO5O0V?$S3^HF."?&R>J!@Q?4K 3+6:*[)\>C=(KC>+O4_A1[(.MKC+F3N=!0:!_@
P_CXT$OY+K@/Y/?DRBF7YM5AS"Y+)>!++V,R#]1)^&@P+I6D69^Z.H_A3+:U,4ZW^
P;\^P08]<OJ&L'LVW^G=T2XJ8^Z+SH"CBX:6KL"XYJR9G"O=DQ-L4@?(SN'CW@MJK
P,,5A>$O+((:O<*MGMPY.M+#T;:/?SL:(&#X4YP#.U^IHRS;%1"E/./C/Y.F[MXJ=
PWI]392+8/]FD,KCP'#9>^;R3;K_9F?%1^>LLXH>=QF-$K\=(J\!BUM"*'MG^5)!!
P(\0/'.UR?:*T27@Y^#^:V:OSE#ACJEOA:<1V_98R0C@\#UKLR62@)99Q3<A+5'/]
PX7'01:;S6L#03IH,'(B:8V),6RD<*8:<ML<4M RG(0O(0KYM:>7@'U7D!G8>7,WI
P5/+<,>U2F4VL2WPL;F+85!<&IN^I*.P_PCB3V/9_#-D-1M9V^?S68F*J&@A($GO>
P+8Y'+*0[.)B:Y:',T3DOA)VW+ @A"P<ALVTXG]_-*0GU5X\JL*$#W  M(=C#CR_/
PKQS6&N I^W.SPU83*#M4U(D,WSQ T6)?4Y-JG;-S'CIW_HA"1SKMN_8-RM0O,JO:
PYH:XZ)>WHV764/)SN@!KIZJ%%XI0EP)Y^U25GR["^X7:.<;IZQH%'>?W63.C$7B,
P3[FBHO"*+#Y;1PT5'B35KU#G[!@8MP]_*K7R$M:K"$YLNA%Y)^+/\ATX)>)_3S]\
P@1S7P@.1*#P=Q=AD.FQF?M O'D4PY4,*C#C+XFCH?X,[YE?15)R^E5=W\>C8X.\<
PBOM![>F)44 K0UDQ)].IZ1Z>>)]"JERAV.>!_*L]SW.95]AJ=(9$KJ6]300VN 8B
P"P$9Z.K:AS$RY1KI*M@<CS-0B_NU=15:4?R[W8A,;D":),MRR7>X<OS8Y$ZE<^Q!
P,%8SC>7-\\%'G?I4NU?'IBVYK)--5.7WX%2<,KH[_4QE!O$HOD DDP&17"T2+;/=
PMJFR7CTGDP$.(Q?RUPRLP\UBK%CEMS_*&_R$?APH!#$MU_$@+<#XCCQ8K#,:O^BG
P,16Y>#^/3CID3J\:&4M!V! /O'5@'Y,GG/\W,)D!H?+/8_9,"] ]5X>1\2" :0. 
P>16<)_[?+ Q\/\ U@K%%D)&/J6B/VM/4V;N _;:Y@%]&EN#S?D3A9B]YD@84O$F_
P ?P&-4@\:*U:FEDH$*3Q7%M[?2@PR@X"(''+MU.&<_1.W5)_M-C>J;A6AAM9LAAD
PV.1JP]\6>2;N%P]CJ8OK4]*"+IL)SF6+G5F]AR+AGI:2)^?,;)#?7*H3V\W6$4*6
P-J^W$F- ,"$%Q&$&FKO*-=L!$DLT-!N_J$<;2EU#6*4I2^[Z9,S5"C:U\!=OMGM8
P7)U'AR(K]TKRK*>A1OBJBG]K<EO\+'CY-4.#&Z_:*:2WPZ+-+]C#Q%*3\;&GF,.L
P^1+FV+3"$[6NM2]7.XQO<VBF31.\,W)7F859[MJ]IZ$=.>U:<L=0&)6&[E\5V:@8
P+'T^ZK-,=@"XS/%"0]>]XHUTC%@A?WF9:6Z/+=NC>=.D>YQJ:_G-08NQUMZ^.\+?
P#^")SWJ",S-O4/ZN!L&8M 9ZJDE?P>?F\%FSR 0O61-UOTW\:+4.CEY,;;9,Y^&7
PTX-FLKKJ- 8:F!3_(/@F%8L:&+YHH4OSV*LFZ=SF)E#'$Q$^@!DI^)$GP]K!'%CN
P;9G]7<?MU,:%LS@-@?6UR]R#%)O?0W4Y;\3IQ"%^#A;(!' 1%H3]_AM<$N@,<Y,^
PW>?[?/MB CP,*P[$O@:2$LZ@)@4RDG 41./3R_@U>]X.!YH+0ODYU67K"-J=,D;:
P 0XZ(G$$%/<,G0!KU1SNI/,A>TB&96& +DGLC$-J;M#6I=_C?W4!Y*Z8C(NR.BF#
P](LF--G4/?2MIB2_&@QZL!Y!0Z:5VC6#"?[:,RTI%![\1@0!IODJ5NV%NXJ6O10&
P<D %U'KE;>[SDD .HOV *8&(X2U,;B^57,H$"/Q++E6!!#XQ6CV.-R04+;9P9D5P
PZ)E!;P%V/FUDMGC-+>GT=I^&ECV@ZSHA.V6XC@+):\PR=8*H_>$"B,%#.;&EJ&65
P^$N4<W@:Z_WJ.; ?!\EMW/G(9%?@)3$''=O]"O!82?T(KH":M6+6 3%3K,#-:'=*
PAJKP"=G(D \3,Z3']BQKA*]_%>_:L=!@,4I3VD^"LAL=$:$5MG_O4$DP],?N (]]
PJ>[$)V%S\($KVFCB[,\AOL:UU?V/7?RWD(F:(<^TH=.<*,4V%%]0YSUN MS@%R@1
P=/Y_2='T9RO-(?(/\OMW:E6>Z&#AB1(>GG_W@]%8G<T]84[0]B+)26X1NE50I+]"
PPVQBAO=>#?SNBBK<D L@C%U3F?YKG XQ,<.0R\[*X JM[QD&0CU_DGTP"J<.<;TA
P(EDR-F0$\#R35ZZ--NMX@A-4!H/@V S/O2'MT4+@FTP81W1GS?#9];9.SGP? EJR
P44#*B?MXY^;1-C[_*LV.]#FM@&P@(Z"EZ,2D>>D*QAYB&>*G?38\)]GCJ^J]S%@;
PMM')7B(EN'R-XX7CI)E>;F!G,)_6X 34G1H"+#H?=;1#4P_0%-SO[)%P[9WR]LNR
P*.T>Q*Z,ZZVO\&7%(H'32Y4UWL1:DA7*[UI]6A65LF!.^I/Y!DQC^C'^VXVK:>S_
P$!)U>.FP8CJA;Z&80"YNG&&^&20YUD+4H;)B?7C"'U]"6MX!F5@$@JY5&;K-5FG:
P-GUJ9@VTS?U;Q%Q=(SY[0&2+8M2)XD'.MKQ1,W3EB'1$8V]:+'T^FO<[-^R&8!+0
PJ'Y\_4"Z(IE9F8)L!*-# 1=SIX<"[X7_H(/C,67@UT&_YEP;1+!7@C)V]?<U^N&0
P"5><;V3^##\^J3O&?2O#J-"O,6Q0/%8UCJ";G722!&?-&IXZJ\Y)_L-;&!5._M?R
P]@RL"L<PNXB^#B"WMJJ&"'IW,^ E<R!9PUUE6VYKR(G6:R^?EB2&<D8XER93ZQ)R
P:C$>126?=-Z5;1Q[41)"0;1FYMPJ'?)<#-*;W3[!SC=*=CQBM[T,7X_JT+.'@/AO
P>31> 5*+0P>F7,0V,(V-;E4B9U?9H*>DW)W8X# [K5"=^!<VA5YRM@ENOJ+++=?]
P*D())<&T[A7WJN5#_!C8352$6?_)_.PMU--9T-MA$+5U&*SFF"*U8@0%?!A)GB>3
P5A8-,%HLM!2A:O6"=X@3J247$LY2#6P0>08\,IK60\F 3#4\-8T@N:7*#0H>N)//
P!*@7=AY62IZ(X^<.)C^-@J>H/PW]E6L#I\Z;%IL%=+'8G(7(/KG\1E0N?U1S?"'S
P!)%UO,-&C:<X[2 F^4,4*3?"EX4)(PHE6?S6(3XRUG980=Z[\5T\,:P'[8<Z/EJ0
P@!Y/))O20.%='PQ51XM>*D55D M90^+:[-:%Y$F%M,NW)Z H;:@HDG;%&RY.=4&2
PO.1@R%_3(9STENEU]<HWT4O_9F28K8XLPILN)@@ ;C^FW8]0M#+^M<! (-W5I4>5
P9\E3I'<GZ:OGU:=)+O>&KU.G!,HU/BOC)Y?F1,ES/N*PCU<:V\-Z\\584^K[][7\
P3%)),3RK4Z7T)*:JBLA!#<_;KZ/%G+%18".1$O_Y?B3J8):$&+R IH<K9&O%EU'G
P&=PCF3=R=EM5T *&)HGF,6"QV[N$UW SD*W C,Z/-*/#+D0<X4U8#@:!C:JYE&ZW
PHX2:9EF#0Y_*Y64*OHVI.#/#<W0*>$!4Z!N94.9:I;PZ(IH<[?%-LDP+V3O$1&Q^
P-05&9V6[0?YI[(\/X7T&[A_W  0H4)Q0L,W FK/!M"]8M]^UG3)=NN"#?*32S=HZ
PJL,\C4R<B*[9RJ^5HUB?7OZE(',*MVFC8960NF!A.Y<W* GJIJH)20^U,S5DG%Z/
P^>6Q!*R#67'7SM[13S,O-#YH">'K #O()ZHH4=O GQ?+.NN3Q9(IF/>\-NM 0PT2
P B=]"* <D[]VN=/B3E&:/K'1ISEB#MN2\WX>,11_%5]RSDH_JU#777B*YN'5JEF1
PCQ)6(1:3CIXDU-$#0]M91?L,&>9%"2PW:S'AR<QL0^MJ,%N9AW+3A\G=:,K?9,W.
PDISEUFK;*!1HD7ZMI<[Q^E'N)=#ZT.\$PE:\T^ S7VP*#QQN<0M0AG.3O7/[\/]R
P]AX[#J<JSK3!KC#0'PWU-1<QO7?I-_M\.M'?_6!MZU89V: !5]=,:[:;H%M(W6U2
PPS(8KCFF$N':*I6$\8[<!]/3FFUNUQ("!1(EM0-ZEKG]L&\$?S<[!$_%6#;&ZZS.
PJRG>9]2[6R1HA16"P5I8'T)4=KG'67#"&G-BA4"#59$4@:=QJC64 CL3P_9A_!.B
PB6%NUX^*!QN?"]A>CRE+Y/G8$C3YP5 _A]>*<KY!>]@L?Q=#1ID"09JE[,&?+T_+
P&H^[+."\$1^R94 4I*<=!9RXZBN*;.E4_L4V =0[=K34Q76X^FN&7*0 $N&4[L'\
P+KP= 3\MI>JZW7:\(_*LDC"J6(4\OK0[-$.B+1;&(HI@AB567?<M7 #U[4083%Z#
P:Q8"TZ.1K8)VM^//B<#2_E@R)=AZZC'%1-?9VS?-VOM/Q^I;U_8__+%E/;I/)T'*
P%R=#_,<ISS"G2S3*Z#M.CK%EEE3P\ K*0->LUA1P^>.F=15(^0:Q=,S^00%=!L>:
PV*KQ*U&FTW="Y3R<Y-;6IQ^UKC<&#E9XG8#CDM4Q93KM)YHNP8:7 /6S9,O-]M75
PSKY7WZ0)S?CL%PPGR9=,L7DI+S1E/73!.*7.;("#+M'G=KA.0I289!QT$:(0A]6W
P^$ ->2Y!X;UYC>ED>RG'_YG2A2+3TB^X*+QT<NHW)Q42[Y_)]11\UP2K:^O!5XC]
P7-3#MYH#PZZGO()N#KHS1G88;??(L ].KX: XL:"3YPM=!8[B1TI2KA1H'WM5^5N
P8UV@HF<^E7),[,>6D#5'2&T#(@1"%<V1R>3EA,C8V]='T'67YS&D5^11DN%6OH*N
P"C7I:C$D,9/RR(O,L?NOARK>)UE1[$<A;(6 @]UH6"<4W*_G1<P@5'T9 98+  A-
P^J2?*)"ZT"%2O9D)))D/<(.M<T-P< S^0T5X\8'?WW/A#87:WIW48G#?I:+6()0E
PX%:)<U2-IY1UV?D,5X=G1*P3P*&8Y*[YJS=>2_""%SI@NL9RJIJJ?/GK^ 8Y'S]#
PHN2MG</GC3-9R<?%&PXSVVD'!OZ12(J,^>J![#<O%\9=?A5*RYA/DS%<+$#/&"M(
P+3%9S+AQ$0R_]="5AS6-IL>U[?<2).3 N$<-42V 5RM>:@MTO'_58)J>*87K*I&-
PVRN8H;>YF'S7LI%C7;$I]5JYBV"G9,?[LHU4E&$S-U]P-UD@;.)!>9Q%)A"0.MY^
P14:K/7DCA3JP&<(<2[FW X=9!SI/XQ6J45BS<&==Q2X6+X7[B+GOUMX876!M8[P0
PQ?LU0J$/53_9TNV3=I=$"Y&VD'XFE<1@,G9C."HF-F:'#2Y@*D#QI.>'7TX>'*V2
P/-)=D1KAMSD: N]@HY%$-:Q+E95=+!<B]A3;W,]:O8,43C5Q>]3&$0ERE%>UN\S"
PK5]=&M:'X",L UQ,S;@ATW-BYML#J) 2+HQ2P?&1%#Z]JH' 3B3((*S!V2[@,]F.
P*M8,NC*3"^YN@F"7I6"%\=P)RM<P,":,S\&7=<Y"8HL2M^K_Y>.KW!6:1B%"&?4.
P4Q.'H>_EX*A]!9MY.*?D3J,>@*=GTRPY=&2LVT';K:G"DS+[O5<'G15S9[7;% Z^
P:"%RH[*1["TJ&,[+T77V7A0NM!/=6/9LJY)])(3#HMI'A4YPK^"LI<IY1HEJR:_>
P57A>R=X<CE'4+GY3KLPP'N\\O=>_R,O+6'#+0W&-N$X71K,!?5!<)!S;N$S8;?9,
P&5^+CPY/ZRRFA>)UGV7#.HE/&JOQ$]M:BP]NNM[O# 64[G5^6E'J%5&JT)5S DYO
PH3)IYD3J&: _#AD\Y'G.:CVJ"9S5"_CQK3YU>.7+!/*@K@RZ4UJT!HM#R/:QO0,P
P(&[>S,/16LBMQTA%HIHZ\U'4HF^-TI2\H07L%NJ4K<TQWO?)^T7H^E6;9A/7W_FV
PS[NS3$51/B]!JSWY\EY-R$.54S<;*8:O<3:0<^.;B*+!<Z1O$GO) Y23!/PQ]UFV
P!CRY)S6<I[P__0A)*(WAJ32\,'[4FG>$HEX^T^R^03STS92!Y_//N2_5U2B%TC]5
P)QJ8^-41L"B1>E+=!9'7-M8O>>/*;MYRI$08)N'#1]]3;< 2>< ?EU@%RON)K1";
PYU.Z&1/Y&%K?(9PN8@M.W0T2SQ]^#YG:U>=/W03.E8\V-PTTY<0E$[Q7$(^*/V5)
PX#W-)#M(_8NC>%97E_V\R_GAX25ZTF0^S80)VHT4L2D^5#&8 F0\[A.M)]#XW&ML
P4N<F09_LD#S2;3N",R(]\>JKEYV\JKE(&-2[$7Q@@/P<+8C!2+@I^F@G8 "T\*?%
P4F,IG[14OMA>""R(S-@]]<K@!0(Q'_V$A?H;/WREW=#NWV8F;<P)L;8H<.B(L=UR
P[ZAK ?!#,WM*WN%^0-0&)?K^<D\%)TK$!CQ;1<*)Y*O;UO^TU6F(.8K!'L,]$Y\$
P-JJKT&':L[^HB_6S4;/H0 *\NB7 '7@9BH:7!:^V=<K0#F(?P.B2.5^+<0\3 '?*
PFM_3VS;[\7\%8LCV4"AUO _".-@=R,,H>EI&F/^CP_0T:3@\ ;;M]%'A>([S3*?]
P #]U2[@7GFH$JUL0K->U('/16C/X,N,B:M>D\ 3C%"36XLMF$?R'3R3;-.M&61?U
PR^GR!9(&N^<<[V_P/<(;$.'UH51B01ERV"5,SR<RU%+?SF^PE CD@0TY/3XP4;TX
PDXN3<OI&0)G@2^63>^':VZ^?&K\:\'K=7E*4LJ#& =B"2C%HVBGG76I6' +F339]
P^>D65F6E[26K]7+WWKR=?L$8:&#\6=?!A>)CX;_5UJKC'MH-N9@M%\'0QF6!=V5>
P ?9<U81*AZ7= I='S/SS7-]?P$@//$S $74>NC@KU+0#5P/:>LT+_::"?=Y^+'Z 
PUOSIE^+SU ;Z Z_ZTY_ML#7NJNL.4?K,HK%5_\"Q?6K[@R<>]4@H]F^3KRMI_*8L
PSL*U7(^FT[?+LL6"!Y;+ABQ1('UZ:.OCF'H#9YK68?96O!>;TAJ>6.N@' RI__SA
P#,(9AA:=WW H9/78;V8<]=T$V*@T)>. K+C2^B["R?8B5+N#89GM</.?J!9F$P&&
P!H!K4==@OX0_]CV4&U5,SW9YC,HA(<841,B+&I#(TC0L,Z\3;"?&F!)K2K"_MCTW
P9Z<>*)DY4GIL5!5ZG#V"6^2<9 KF^<9Y?TF>C>ZO7OU *B$;,WQ&L(E%>K%+Q^Y$
P0(CIY*AW!7>NK/]^Q(F_EN6UO9J4<(SS^OS!PI7)Q9K=)>QN=T/*04WE?XRH!W#O
PW<,$A2][Z5/H44I5(M 3\T,=OIOE&J/F1_^A%,TME-CW>/&/_Q,O9(>&G5L3J4VG
P$?6NI)%Y4/(?+G, 2X;\\ :'!*RF7V79)>:*->\;-! O6]K8KU;OS&#FQS,H5+WH
PWZQ(902T4\4CUZR(<%]'&XPDCBB5_*G40,5JP./8D,(9^VCNBG&R:^/TGJ_ZF5@?
PI/[D>2.I^:X?YP-/ENL\L!>#E4LXS('>&7[=VK.-P(ZPL3U]>G'AYN,C-\E8QWO*
PM^J^0OJFB3!MP#UR7%I&R%13CS0;TCU U-N;=MZ @Y!NGR!!X!KF$>[AE6+-FFU(
PJ&0$+N _]@W:24*5^%O,$MP\+56 C&SRBV*QLRI$$.I/W.-$M+CMN=8;&>P @^U?
PF1D3K.,C+1XQFZ8Q[WD4<4R[GN<6'[8_G=W4[K$U"QB]'/O]R<%68KIUEIM^",&!
P+2.FJO)(4:QB(_X-$GM5M7HW'QUKVT^OQQHV<Y0$/%(H#8S[H(.?'IE)E(VY'BB+
PY$[NBI,N1A3_@HN&OA>GW5=XW@)F.7=%5.^J")O<LY]/W25?<,6#*RE0P(*I=DO[
P<(J2*5BCCGET ;5#1%RI+(=':BW$9X6.%,6&]1I$<<MTI)QEGOO>++-=IT*MQMA0
P.KC3M_0)OOH[<A5!X>;.JY^S(_W)<E]1?%?2H'K'A/4PH%ME?3JMO]?/3LY&UHMC
PGT&IL17=3?V</!%2VUGZV&QF-%R0>U6'TG_Q#>M$]7=;(/-Y\=@2,'GV7@!C_R3M
P<N$,@\MHLLD8QM"1O;NM=:V.=Y5.O9IV)7?(%5W=@;T'=!P!,N $)8"0#L4&&J@B
PO)$0VAYCTF..WSL!F+K):H1>46!QP <M8"MT]7E1I%E\%]NWT/FN3%ZS-49(].)3
P1$LK<'80\5+UX?DXJ4<9J4W/*?$,0N:(Y;+]37O N<Y-[&RO ZA;V[N_,]6FK ,L
PH4HP!9B/T@PFESH$/[J<--_1YR?B&@\0F^94%@&%U;X3!T[I'=Y':*",J4E- 6:9
P]M:20;4FW>NY>)Q4&8#X.8LY]6PDI+*]2]CN. ;33,M^1%"%ZULPV[*BOI<?'IPY
PAU_Q25<[![IFIZ34(UCC7=[T;0T<<!7$:EYS>M/]TY>-#2E"(*5'NY^E6$^KML0/
PR4LUV=D_0>J8:[JX4SVFGROK76Y+MIV,:W5'1/LGFTG (M&Z-B2(1_>"8M^MR:4P
P D.MZLM8LYU?[5GRJT^^AV>YA6Q6,T@WY$P:_NHL.&!C#&RCGM.'7+5M(T>V;\TH
PMNY421GJ_+=IL,7B[ 0FKJ\W_8>G#@B;];,]F.H.%M[+51OON6H--IB/_PWFEOA5
PYY!VA5-C,,906"0HL)FF>N^"NA#O_85Q(X(&:5\N?:SX+20.#;#UYZ_0QB$8C/E8
P]"R6^TYJ),,%2U2T!^PW9$.&WKS'U*^!65%$@Q][E1CHQ*=ME^J/;@?LCY$FA)O3
PZ.2*TNZBO'6_V4,_5Z:H']35:UIL);!<>B9-_#1H4LI6!F!W)D?\3 L"TIH->K->
PFW\W?^L-7)/R-D7V;2E*2 ](PE0>66Z0Y $"I'O0!Y3Q1)5?$$3,MM=_F%?M(N$,
P""I2+_/A'K]ZN-E2O])\^DO0;0A=?0F$QCA?F;)\YJH@?(G<K5<77 BR_)V$8T@S
P >R=J[N;*E0!!E@RFUKH,_)O3!O(*-13OI $)BFH79];T0G]X%UM<B(/EEO7[@A&
PE* 0:T$?H6Q2Q[IQOX.1$[ VQ.1W=5[]C3/AJJ;HD<\7U)@X>C"DNSK18*B!!![+
PX6OR"<J2:*TV1U&)@>1@ -TPFYNJ?NUW#Z=^)RS5%YG2^(B02VJX]V.^R:SF@S?1
PM#R[D'8"\.GY5AXSWUH@$W]MRQ5&L_1^)4$3 VJ9AI(&>TC$O5ON2_ -%W]Y%+S^
P8%7'5:!YE-F7BS>!E?(DBW*9:RV[,*/!+!"_(NUGD'B043]M&,S(.DNFF[B,94 9
PDTP(#K+^FSPW=6W.&GW-SB<(E:V:22&*8QLP'(5)^[M*?<K\)[%@(!1ZO1"#_Q>&
PA;H@N"A]PFX[R^UYS58>B-"<> 3CLPZK5!.9YLDU^$ A,'HP4J3)7$DHLA,WRZK%
PB6<L[[;!:*9]=O&97Z051JL7,]B3[LYC#J=A:$'!*+A_S 7NE'I$( IYS>75_G3T
PO0HCC^$ MV2Z@8E@5&0[W\!R/!EFMW:'@3%O2F.])V/4P+<3\:,:BHWO#9C24#W<
PA]WQ1]4ZEI&1=*42<,-$-S"K4A2$PPZF)J^G#3A$%.N+-E=_[ =.=MZ1JKY )-<M
PKNX3./(-V<U?T^?[A6$+@L:I'RV5OPVQ=Y.7@^EQ!Q 3 >U6.G1G]*IWVOB"PQ$5
P0E6X+4>BNL#/56* 8;]2.TCUSQ\23K9Q*"S=MCO&?A!IY@Q*Y^->=Q</; Z1%/.I
PA9<7&I]?['/TH1X7,!?RN@/P8I]F^F=4+_IWPW\0.SY7/I^$]EXD>=EW9RD-%GH(
PZH[A%_'J$/IBK-(N:9JVQ@8TD'U9Z+K[.TE"!O_2&:BB+9 ]4_J-X%VP$Y^.'_*Z
P"-@S4=?:&^4C,=N?*'+2-?W-#?'T%('R/G;)69SY$A\B[MRT2RDNZC_U]*8SHX2(
P*$6SMD2;0OS]:T%W5;Z.2VYK@6>;4?2KT&3UORT_?;M9Y>#(^%-J1?(L:5S&!3?9
P223%$BB75A/Y";0:.6NL^WAQ,,-2:#?"5)LE\9R.5\I&Z#8!8]$ZM:ORGA-+U*[J
PGV-68$JP8V,N(AV<)MK-@S7TJ\*9W255BM)GYOI,PS@ $'L^B$Z@VL7^*4GQ,HEQ
P&U073P)D:M6FG/V;\)8G\18[@ 'NCOU@#'CXN!@C3<^7E;?UHW&VV8#+?;F3B.E.
PYT6]41X6 V]ZP?-\T70.3=:5O10742'-[E'DQV<!/#YAGN.V:]HR(R&1\S(+-IXU
P\7)F!;V8W2$JY.Y_"?\07GQ6@V75'%/YSO*Y]&RWJ(+YD!*!#%8RF8?7FLB']C =
P\QJY<4+$QPCI GVE:62=JV6_.Y>8.^1%_@2>(BB5-5R9C8C655>^4^W74W9=$1+J
PUR,TWSY0.B)6^%H5,^%1@ 5V)_;QVA&?F1GX'N13[@F!C"J<F8W?[S;89?G'*_L,
PZ:1)G<*:S,F&-W5[0[BLNS,BGGG^5%7DDR]!_!?V^DS(2MH.["L[.T-JL<IO@=LU
P2@]M3K!C[Y+/[LC\Q61NY! CL,(_;KP,APU^($R,=*3H9_*7/[Y7GGBAK:4/"8<&
P:=*OK&5C.!IU;@0E"$0$ H;D-JZ^0[FS@E)RV$R"ET)%6)TJ$RIAX,P9EB>ED840
P6XE#=;''Z(IR1R4(38QE<V)F+J/O/2/VO\YI-KF%-.:)I> '.B^C8O5&SSHV@*-^
PF.R4LI,78>M4M_*R20.\F7^<O^YK4!/VV<"660O+'*T?/ZM$3S_YNS0R_F'@:UTO
P-?[MTM6TGG655* @6N+EB1Y>^)=2J\N*_697(0KSS!XD,U5#I2.$C>\-ZZ%]Q] -
P_SW3(ZQ,HRPQGF],H-47[WB>/E%E,GKZ?OK[,4C>-\@VAK<UA^JAK^WTGZX^ 7ET
P?_J6]RTC'61:X%N$Y+M\1I-/TV3*!\T@<#VKDJB%ZH+Y29Q>&+_0 PU"J7 W\.N_
P[-6NO7(C\YO4,8(@,2GR$6IC!B<40I^4B"/R7GTAB[#9;Y:[ +:37@*JQO3#JWS,
P9(H1*F D[2^(X=J/YW-UT&5Z<#**1/"SUC_/#*C)6$)]F"4]V)<E+(&'Z8 Y\RNP
P-2,0HW73#WX._=KR<RKHLAJ^X"!4F,%L<[+NYF)C/SX;5DAMM1J]%[/KZ/G"/W#@
P8HL> !DEC;%Z)/1O75@".J'@KR:9ROS6?0V!%7%*2H6.6]Q'#M(-KF+GXUK=I6WI
P_L<WR2-_?00J#PX>J6^]_C\Y0DD@855.. ->H90LZXR$59#@F7<+MOC%[7RIM<+%
P4(!.[W=[?8\ 8;TB"6?S^L.WQ>OYZ.:J&@^L5NV1M(7%#!5R?9&1-8N2FRN>D;W(
PQO0OZF.*QTIJQ5,'RJY(#S-]KE\L 5,L6. 1:98)!8PY/SQPA(O71XOXBF]-V+M5
P0"<,^3&GTXQ$"K5H&2?['CB/%G1> 5=5 P<;3_GO+8#BS**..#)($:1M;?0&3Z8L
PM$5U Y8J%!?QW1?@Z!1R>[<_'%W\8@C^'R_5Y> YO@/.-7RWDZ()3"29A,@6/7O(
PD;WJ:4C;DTU@%"MKG2N%<R>S"%HL0++-H<Q<3QKP-RV'L-&K"!V+2T%4DC,Y6)JT
P,,!"_4[MC9+I-;9&$FI[C*[I2-T_TY'R%.1"9XT:$^;-8C29[XG9^R;Q1/4K'WDC
PHD*\<ELO+PQDV].2)H(3WP:#JHM+_OL'PC2SE*+06N04]"Y]EFN1@CD(\0YP'Z4)
P%@SDV)N.(9V&-4B<Z'D%S].Z^V+TS"P=>1LRL_VUK>);PH_W2E<Y@VX^J^\QV&6>
P 8!5C)_T'OLO(0'7AG*0,*NFU/WA=7P9 $]37D0O'16[.V!T-17B7>00F(VI(QH'
PYHY_*E%)C"E)[]X_?+3(%A2XAL4@P3%[]9Q-+KS;']U*B%3?UA2>WD>B5KQ%@.\S
P]H*-6+R24D\TOMS_BGOTDGNK)':BZF^9*_#)!6^9N_Q^;3"G^SLGZF*V&3+)Y+S_
P/$R[82AXB(#=F@A-XE[854-S,P[<O,W/#7;A"0\R3WUO&$:_6ZOM3E;=RLH84<0Z
P5*HL5WU/,9RC6? J;W55O:?U,#P_E+\3)UD/4P8;7P2 8;_[NR7!=!3A(^)B,.O9
P)X[H'F#SFE%1N$H/TL9NQF][,5.BJ9%.JN&J84H=6_>\\/(+U5$@_(&5!L_,)]TK
P&^HH1'Q/R*NZ#K)%]/0T>%1*;6U<W[4@ G&T=4 ;ACP!Q6NROA: WA3MS#I42HWM
PK6D5PP$YD87D^+9,LL29_@$(=QCVRK@O-2.O@-?/@<5?\W&;PJDFVIOSF>=6N[W.
PV(MAA[R2O-]%?MAE9S $L.7>./^]_W5-C&'=[;J]))]*34T^G 54@E^AHO,=4<#@
P1P-DIEHIO&C&$Z;%7O=5QT+U]3W1JUT*-@<6:T[#D1M,X"0N+:><K#^Q>.HLB1B?
P[?YDABHM#)W%*"4T@0;M5_WZXS6L,HO0DD[3O+YUQPEZY%8U$I/!! 4[&",(I#B>
PA\LZ[DB,9&\I+L=),'0:ZJQ12-8:2XP>5TVA;CWW8RH$#ILG?5] X;UX6<'B3ROT
P@"V <I-!;BC=/8\Q_\TN<^"F2QQ*FLX<)3_^.@*#T!X:&!,I5EQ>3UC?K.9C OO-
P.[4^KU<F-;246<98$48N.?!QU^ZUO9Y'R&[E6)%RZ;#$";E7.#3P::WJ06>UU,J_
PO/@2A;"E)]L[8T@92[R]DP32G.'J#+YY; '7];?NY8FR5@SB!HR+$)2?V"$A>+IW
P4R>V0 :#:O.QAR09VOD*"NXV_S$$11:SG\.\I)79*8")S,&+&"T R9VV/1A/WKZ3
PJ5--MP]R%5M5S.C8^7DZY,*_0S0XY3]!=]3:@<_6%C.E7PQYKMOAE>"Q6JW8%(+>
PB6G/I-_)L@2&<->0H1#.3U1+D8SL?[$;/(Q'O R]1C$__-3=@)_9!?D3"+6P;X'_
P?K%BZ^N 6P)6RA3/9'L@U/F6)!V<!;M8)%TU.&KHT4'DT#E\ Q>IE.HOD3^C1I1,
PLVLQ#V:?I:JPF9''ED\"[ />M"]@'0Y'?.!,-2_F5A"S]TVP'C9+OTFO69T!OBX 
P5'AG)2S$-Z2Q5O+ F&$J79).BP]C+*S 10"3<3Q1, (>C4F(G33=KC(T^:S+DP>*
PM$:$M"%BB2P^2:T]F4,L4,L4',7Q(Q+X9=^I6H^<(M\F*G$(BTK*S(CGOCROJR."
P<@C%^B_NYU8JR;T;T[?UY*AV2:SG);*7'+@62.F-#/0_%::Y)%5HO-_LJJH$C[Q+
P\.:+U?6"[>9?)::Q/S'>D#J9(CP=&,.+Q3ON&)FLL*Q(I&6C6?M#P>3C<$K:)^03
PJ$1-JM D=][3!$$E%#4J L<QL@YA<GUSV+?* "B/GJ9$#Z/]PT#I=Q9KO8L!0@\B
P[,-R5'I?_79A<\[ M<6\\RN'=?8+:+X64>8AYH/.QX,5])6-><G\J^N[0:A!3[N;
P@#L 8LH-P45&LJY-E=!TT]B,.CI7XCM+I_BL))S$=>E5&\\;HE7PY1+ID^L\YI_$
PDJ&N6]QHV=EO#P;E*M&1 '[8>OY*XL:?(5N$C?O:6U$L[APX.7\+JNPS&O1S]W![
PN=VK]Z],J0"<2SCR*(G>A##F%7OHH)UN\/2=BA'V'?+*:BSBBM; -/1S^H?W6*TB
PQU1('PD=R$NIEBGO;=WUZ3H.P 5_50:6'.]I>=2KPP;B>Z\* S(*_MT6.L:L!30^
PP>)29QVY_Q+W*;3X&YSVK,JHOMQ'^T*B)8EJ32R>T:@]2$C,D*YDP*F;":9"SY",
P#$%T*+IOS&R#XLJ807<\4/4*VHGI>(UN"J%PS"0?RVJ&WRI'H#EC#D1A4\ 0.[42
PY?PJJ2EOW[2$L9"]"T L;*40?!JRN7=+U*/^GG66("(&QN,D"!=,)U:7*N+4G88V
P026I-6O&N?O*G213^:13P3<M&G7,L$!<SLT:2H.D'XSB:&HP$_"<HKPHQ6U426J>
P5O4MAO;<'DN)S$(BS*-8/*UO.A8%/!R=TPJ188<P=\[<'@]\>;ZRCKDDZ@,GSP-(
PT\Z@^=;Q[T9KF1A%P[WE;NV $K^Z]/Y^!3;L[+*0QO/Z- ##N7!(@*I^$13 .A1$
P_PAPOL;N(0K#'C.?0-U;/ "47+<$S=H-*CKF=FLSY><U7GB_8Q"^&:R>ET\<>,S8
PZ7KI:#,<QOXCO!'IK6.BP2-R;"V A;)$'J-4Z3>/<@Z\\L'"S3"^GOBKF6/J^:+]
PMXXC)S&<L9C0/ZT0%-I'JI@.P#N66.,6]#;+:?X1O=#NN'FB+36- %9>\,G=I "/
P/ECPN&U_Q_N\6UR *>:UH<_WH@C0"0V9S:QD,04E*7H *IIX@V#1KP5P:=O&ZU8-
PIE'$QB! 4O7+FE1RSA=<S5U^)\YY+>$>]ZF=EQQ--MP<GNT9QQB.B4'QO7H'=^F(
PQ4]8RW7>1, +D7X[B6(A!Y&'7TX5I7!Y91.S</'=X1B'1RNY-FP*I3U_* 4UYV"[
PTG#X;K);'R)V1#O!F\BVU&-++'#JISZ\D.T)@'J(F(8_P/(S[7_@WM1D8^0%S(>6
P3X8*G*N\#ML1P'6_FYA'T ;U-?N72I9$0R1;8/.TKD3W<(AF=Z&_9A-@($+[:Q2D
P&+)3DR32>\ID]+G-"E3I$-]H1^ZY\N*]R4-'\$63EOC Y03/,M&<5-P-X@JKH@KT
P]_^#&FE<96];<.3IK20+U _$W\!/ <0YK:B2&940!!<J/?=/>)96MW9W(V?^NF4[
P<8+UA[W[!IXQR?D$\O4:'(<WFI+FFX32$3"<QH@PX4:FR,\@CK5LI=JT\6,E:1//
P@,O+XX)._/OR/^4=K<QN%#)G=O0B_"9/L01G@AJ&91!8B]XH"V*A2*JJ3Y-@]E<S
P )'"7/')!(%TR0G@&EN;74?/%YI53B[)R^ )UX)]=\*?&#&GXVW-KD!0_A_A=*%N
P!=<>U7PJL7.QK_JR/TK(03WV/@>[QQLI*9=>O9&DAJA9H^KQ2KR@PZ$47=R&AU(S
PN 6;7DO9FP%[U%Q2N*S/8BL*4HH$9Z^0"[RD RAA]O"*&C?8W@X=?#9ZD[N+#+UG
P[\=7*^!WWW,66HYF#8!+B@HI6[<,OMTJC9U86GZ??16HEMLJ:3S2^-+3H !T7'-4
P-'%!%@R+S,_'\1OA_""3^DNGTR1/F9[UL&*K1\%6P/*4;SNO&S5,$R<9D A).S&L
PZWF4?Q>^ZI)LD8.6SJCPS642PSM+,+0@*,7$B\;:Y:VN1T,'(S#@:5J>*076/##$
P:,B7/5.IY'G:^S^#Q1?!@AX1 C,0 5A@/0?Y-,V#% 'C0QHP:T\)^=6IM0#$#6U:
P69@.((N$.VTJOKL31#*PU8LR1]D9)YBK.EHCZV2WK=5,0B$H-*&KD@OT-:J Q</0
P&JKSDN3HNUDK+A'+IKNJX*I=J&EK%A_2J@*[:!Z5M8!&9Y3=MAIND^DK4;"00X8>
PK-,<#"G@QK1,OVJVOP8UK,IF2@CZUZ"R%GCFW*DD?*90''(!MQZDK@0J[[T G[LR
P<2%7J COQZ]+OV4"''G >RS.^4OWQK4"?*I0Q2!4U9:S)YW==MG-UN/O=%T/FE)K
P@X'+[Q,&.B#GQ!%:MKN$%,QH&F+Y($=NSNJ[JT/F"GT+(H -&BI13_@EW/S@5=@-
P,OPOLU4P-]@0CH1.?:(+$%5=CN3<V?:JURU9TA0'>T-M+TN]8_9JM9FZNO9+T5HM
PVYTM%BKT_<'="Z</0(< 3H5RKLGDPD96(FVN=2O->J+X*1&..'[H4$Y9'S'@_?_X
P*OTLOYZ2/NI\"29X*3#4]@%DI$TL.6I^*ZT\AK.OWA6R  #BS.F4LTVB*;<BL. B
P5([".J@'27-*=S>3DW_?,^3;/!UOR<Q^Q=(\GA0, %L_\#AVO'F.D5! LZM1KW2G
PM_GCHDR9$HT^TVX+C.J^!6AU#OR@&?Q64B G<EM)19<%TSJ)E2MXLA.V<(%B]3K5
P>,[]@<>O:AG%7#1&1^8G5(7'PM%CU&':W-^7]".R39$\\1O:X<'"6IPEDCQ&-K%K
PU+VN;\ZXYY16C\ZL\,B7A6TLF6&7%D@W)NN*G!U0,(5>:U45<O,*/8,&19[&XT3'
P$M#D5A0>20;;ZTCW/4@7* SU^A2;$OF/97ASYSVRO,@N'WZFHY.$940NBBGRXH4+
PX9@5)BAV^[0:785=FVV\Q&YDA 560Z.6J-@K50J)IS?._;/IV>NV11"6,D*;IY=S
P&S29\#78$2&@;[!,"#O!DQKD>I^V,[\6Q/&2D.CO1N/?0]@EC [2H4PBP]99M5$U
P4+EBQ\@O^3$[<AP^Q\R!POYWXYZ,VN8]67L>?V8/AGVQ9TBEHDY#UD(1R,\I=3DV
P^5,D#PD3@98L,"T5--ZRR+R ;]K+$F[X,=/SOX0O]X'X2_4C&MLO;JR3H_,M9JUB
P*&25;I$[M3<#6D5F9];")#I09C>XVBR'KC5A5B&9**K%+O]URDPF#/;$\#2D.2GH
PN]4>/8*%*&3@B/:?)#?Q8< #J+Q8'<//'%<K<; ],\JR>>Z'2_T98S423PQ0@>;H
P"3[T=?>-;2]F(!B9\Z1A_H:7N?MOF'Z?XYTF$;7[=1/-N&H0IJ#><'\>1XCNH_+.
PR-*2_&>E+E9AGQF$7H(?=*XZR_6_FQ7G!GG>_\.M9^]M949PN*^1+"9( R=[V'_L
P&[&GX"^!^$^KU5'8]=*@.79V'PJS)H4V!9O*6PFQ-TDJR/2H9\97Z%O0S&XX\\U$
P&U'.W1I4/L8?E REF*)$$8_PB9F^/=?":7UT5.E=R]Y"!6YR?8(:,$+F49.%I9^/
P<)6(D0,"*ZL,O6EJ.&0!IW<$7,1#6SII'^O/A^X:TP+V>^[TNNY:1Q,R%[?0IS*T
PAX2<-5$L5W/4%P,<\8.1=(_CE[,!)U.[>S#4,M\/@=(<8"JXU6]_K]?\*!)4=.T,
PZON+$/K9*KN;/M<K&2=+'XGP76ZP;;B@"T;\[^!7TE7_ JA2?,D9Q-@//^58K^$"
PPE>&?DE]^_5\C"8_<F)#LRY?.QU(0@">)C9BI^'I@DH'6@^U+$>7,>G)8?,Q7H9@
P#)9XIDHJLIRT#10GH5RREF;S6ECIF@.F=:2CWQM-E!2UPO\-R?TGDB4M[C7NT]<6
PK650L]B@Q.U%MY5\MM]P222DIZQ="4".X>P='GD9 9+QAA/\A',H#E3AZ6:!V.E/
PNK2QL%PX^LKVD#Z!6L^%*H =J(O+]7,DK?\KD+7(?)IQ=\(-A+WO9L?+K@\W="5#
P2KZ:%Z)W<N%]2UJS9#N.+6#?V<85+EI,0F$'IZ:,B#0</AJ ZQQ1*=90 55_R3&*
P!TSB(/FZI(UIVKA)ECZ<4-A('FVD-A"MR.7#S>FRP;<&NRKY!F8D!0Y)%$+)\"7!
P&>WDGP4X,^$R<5A0.;1CF<#T"^A_FR7)B;1$@\T)+V:.4E(HEF"[J!T8V^?E-,42
P N#T$JV#];$YCCN@-^-DN=#YKV9)O$]0_]W]<;[G57?:L@!A, -OS4Y5@L'P3 \A
P%3;B:8/M>DG@*8$& 6W.V*$(+XF%+E]W/ 66*ZGF7YW+>(%^2,;-QH"-47#?>Q"-
PP(!CFX8*/4Q38Q?V&5,?3DU/4R6)20Y2N+8HZ48?<H*;7AJ[H@(_?H'6ZK/ICO?S
P1!3N)\82>%,JGQ2_*#>6;W0 B:5%[2[6;";(:"<?8D>43IHO'E>OT<NT?AAM1QJG
P#&%/VB)ZNJ.%TCMA#MYA*T"Q3]S^2_AF.WY"X1QQ(;Y<9E&[=.FY1, -D+NH5)Q;
P-9)VQM/-<#P,06:@YH;JIT8,$-!@1%W1/1,!D,C.%%J"C50*:E0L2*E#W<R BDG9
P"^JWY!N *W*,#;6 .Z_KHP>&@;QI=Y_;Y]OK>X=>LNKFW%;#;![&K6.P,$UY'IXQ
P$7V\#8J$(DN%K>="DAUQU$-G$U/[1Z22.9SM5L\&T;HO%V_8?B. (] =/3WJD1SL
P5?JSOS"E1=F7/$GHA] KX@"%^]6\.H0C@PXXA"!+P(BE(DE2>8<I)Y0EI0C0+CK3
P'J*);["G)_Y&0<J?/!VH<ZPV<CX8!\) 8RFW]5P;I\-^\G..%$.3ZM-8PG*69=F(
PTF@+_=MF%[TA+[+35BDXMY8(H]X;H1F240,.E?$@VL1;]O4)75RRQ@Q(R--_@X#1
PK'FQOH2F_EF;_<G4@+)]X!J>AF,%[(VA =(K?+34[_N!GAM$T7IJ.:FP" (3TZCP
PW2WGR_^HV+TI7T&=J>[8(#Z4U%:,,OF(*DVT$YO7$38F+A:<,W'W6I<O)/P,)EC8
P#-\]:';<F/_?_PBCC_L-PRZ9-!;09S% <-PW*4C:D/&:P[U6]<OYO=ZROW$)FAMM
P<<BH\))VE-52V_T9LA6=W %:V]:"(N'C[P50#ZU0K<>)9;: _>&H&;8X=7/BAV"Y
P(4&\Z%=/TY\(STDPN^AJ+^W)H<P03#A04_YG+(8@*SAOR/Z=IT,(MF'3"!D<#LR5
PL@JCI.M,I0L3[IY,%G_0T.(OJ"MMN5$[K5$J6_;;F"R1<'&R,+;\P?E-;@.HM<KM
PP%9[D'VW=;+K1Y:4_GV9(J__>QW=#3JX&JWZ-2@9J)0"HL2XL$W7G/FG"C4;EMX>
PB4VS.I> AT7^TGV>+ 'C'U$GA_^31X".P/Q#JE:10)[B 7T#\)2<Q_5$-F:H8XK5
PXKW>.?$*4*XIP)4C/<ZG$?5W_OSEBYU X5)8%^G>8@24!LK<)OYR^PP_]"\HZ4Z;
PD&KZ87($.YZH8DK7HU(\P\#E;)8Z@>(ML?87BO3'>**G58F:21$-H3*+$\>X<U5=
PC!/MWI#3A&.QSV"3>N2C+B$9U,$7U'B'@CG<(3#N!+</0X4HI6ZA8O9#A=#O2C$7
PK&Y#J RV+$,)[F-@%.Z8+_HQFYI4%XA+L['XP5G4#!.JL4H)$8W8;1."-00S+A.Y
PT4NI]AQ"8B4^DJ3T*RNA':Y4?2XC1\%M9AL2HD,4B@8W+Z\FTP"X"QG2+,TT@*G'
P?\GF.0EY$IW?X6+- K(#"MF54KD([B*&$8!Q[U8X.(SU.9MF2W[XZ.L'E>1Z-A(@
PA#=-W/!66M7Y!;IG7)IUU>Q8P!$1@Z"TV#>I8VG[>A/.P+MRZ5(+VR&,!'+7HOU9
P/> 4W4I0C::4<<F%FR8RR6'F;W '"EYLK3TWOCU.)J!.6!PS^0JJT*Q%?AO TY)5
P\"."/E=]E073'\)4T#^EL1=5BH^2^K0\5\8W1QV.<9*3G%EY17E%U9SKLO5=@U:%
PR@$D Q( 5HM)X802C-;SS"OS-4ZELGGU;TNIA6*LO#HI8&[\%3#A]1(TM1^$VUT)
P]#AGJ!D2\2C(O?[<^3+^NOY\D2$=-4\G@C<H&B@#WN7/OW.U:T-A9>>2*_8.XC6:
P3'NI';NPY3CHM!)B"%WD/K5C'RO2^,5[@F0E6N_;5R7A0;-&WG]KVINW"MD_=BEW
PM5%S"B=Z;W%_H+!XD<4Z,G(=^%6NH*/:/A7.J^[G?[/\X"I6$"6DHNW-,PZ*+&'-
PL1<Y9RG@BT^3MJ$]X_;8#G3LIF8:NL?DM)@'7.PKO71RQI1Z 8K#%&)D!@&F.WGQ
PO3W2,0-)&44I$7M?E8)7+S&D,Q1THD/!9(4QXMO:16/I;'TGNOP5AZ6JB?+ I/$Z
PZ$2TI['L\H_AWT Q,QW+A:A+RV;3O64E7F^D\[^?,=5,O"RQSU<"QM:#6GJGX .$
P?D3N35QQ;(W%-A!;#$,C*^JE*VOW'3#R#&)A2_96P*6*&=V5X1LTX*G#*IJ$JW)3
P_I13S'[1#,:Z$F:&IW^.?$O7([W2$K-B)F=WKYY[=^OZNK7J= #T[0HI*V2P](L$
PP/4/N698AQC]AKP*>UUVO_QHX#&<5UG*/H [ZHS7"#DB."-8.3I#_&[15>-=VN'@
P=)FP>YR804F,KD?E7UIS9?C<=.#XU<G^HP_,])A>::=V: 39LE!I?J/#>ZTE-)[*
P'T4Y);4LJ)SDK'NMY;FM!R&]9_#BZUA>NV$/:K"X.0W6L'>9^? C&YB\HMP,3MX1
P6B [GR.-^%_,!DP$J.)FUVFYZDN=Y1^Y53NJV,0A>'J\M$69P2PF4)I;!"XV ]L+
PU@8Q.<+15OE7I3;<V,QJ\B]( K$ ^(%-^"A,W*/7#\9,0NLJ!0^F%07U& WI,$4;
P4JO1BX+HI4PY#P&#V,,U31O)1'M(?\89I ZML<Y:[M/]G>IWXI<K/ADZUJ,2=]KM
PN;FHAEB9SIV';"3K:%WG/W_L/?>]:.U(UAP."Z7N/Z^ZC$ECZYH?BPA2I/IVOF[2
P(G9>5#@_LE1S(^6S9C6BXJ3?V7/<.P6RMO\$4A1L,H,V$> L&ZVEK=*XCMJF1 -X
PR6T9X.NGQR->8'U(7J/(>5\(;C%U[2S5))-K7,S>3MH 7:Q!6C"[P8J$<.;Q_=#J
PHU#[W(F-2Y)A 3YKM<J)P*$UR^/ N\R+DS-7@&\M>'+86M2T[5[2DA.6U\"[]-1E
PG//H*OF0/C]<2ER2'Q7=-=?6D;\80.W32RT3RS;2/!X&B*O&=N<<W_@,2T71I=_7
P3-4L1KY;!,+HFU@31*_M-(*^QS49#M&=R[[FIR)@19N !K/Z 1*CY!%[!+R_7>RE
P$^FFGEFDU?Y&W:^3*A#'Z8R5V,AN(!1/LN<V9B>#JEB>A!>CCUTGV(V8HZ)U4"G(
PBB?PHF$!A8;#N-T=;6# XRK)C<5Y'4I(_'M,&+&$<<P.!Z+<B9<60%@_(4'RE[3]
PEF-,9 Z3]S\K,1;I,Q_[ L+1_9]AR)E^4:+,N[LVS(X^B&LIJ9_A\J&30!:ITZF.
P$T0<CO/>Q[YYXC-JAPA%'Q*D-E[P1M[>PH,)BZH;JCC1PC"AMRUDV5IYJ&Y''TP>
P\V:D.-9Q!&?E$C\<+FKN5OK$^SG<OH'AQ1M)]&[VHY%T5^:IH%UP"EM2"+=L,C/5
P=)$+!1)(\HFOS>P[G5A_"AVJ^YB'D887;W74,7-G/8<B^'M#^@+$@K5YZ\+6]A%&
PL3S>@A'3)^D(Q?_=E26]9HM$:QG04<))JY5\A2O,OG!B)M"RG$U&@+V+@C=8AEQL
P@B$6\CMA!=+0,_UF8K,E4\JQS3R-S)V=X1IJA-*+.D Z1O<<DD_FW!D-O3[&)^GS
P*Q5DI9'$[](VPB?*;;]C_I8J"PG@.^0U"0BT<1$]''J'SPX-=A<Z?/OO '6\NCCF
PS#G#-2B?^9RA^LXSISK_/GVA6;76PJR6..?)2I^SA997:<\]=2]!,PY$=O-SPD#$
P4WU_UCEN00O898[=W4[O?%"QYN!B8K_ *@\W;\OM1(LXB=<H:6 H=)_/$^W]<S&F
P2AJ&"SP)J=_%*U8.9<1PM.J*@!S/K&_]2A!CD'MY579]Q#NY O 6T8.W^F^<$R%Q
P![F="]'JV!.+7A2J* G@SK1,/LE3(2RP6N$X7/" 1ZNENR(0D(;W6Q^!^KU5X&32
PK&Q3^CN[.O06")>L%IY1T[#)42$L'-R0$C]L/9 *:2ARC^71KI8M]1<PLCTNI?6P
P,0.K/J@Y#E3YN)H8O:YGW19@ (6=]4+SN^']^K%D/C;YU%R$U^O']MM_BU4 AGKD
PU'<1'S%$)"&M)$]I#/FP]*C?9:+3 !?*#M"0,1:,0B2.5%IVS$6B8MU8)RIVY=)X
PR9,I+DF@"+B![516X*:O)-0X9ON(@G>Q&QI'PT+I=3QY_9LYBS?[IDX2HI9;JX/:
P(B_"646L,CNBRLDMR7H[G82HJ2O':'!Z@W\.Y=O8]<V034KS5=@^U@A&Y71KBUU+
PC?UL_FWIKT-2(&[^?H6=9DQYC;)&M5E=C[]6K-'HW0W;:%.=+XH[?CX-,54('Q+T
PEP3PO-SRH#M/97_VI$?%O&YCB.A91"QP.!\&U+9O5LR.U'=?V4%QAL0'Q"]>"5];
P\[8L&!]XO(X)\"FP9/GQ5/<;&A<P<]EM=2AZ3.,Q]]AXJ0,'']8+V@YVO'>#A<2@
PZXL\ >]HL@\O,ZDDW3HN:^ZR[:LNF\XG7\]./.-:(]X?:YRKTY;K7MRO;OD  "6K
P;#"&I3EG2YE'7WT7W6^7!^GQ77S:R;&R0[4V>>5;=!M $XHE8])_)GS\#MCMRA,@
P+76^@D#6O#F!Y-Q&P5?:D<T4[@A<'@V+!?E(I"83T?U^G3I0T\S(_SM-W2]H5,+C
P"% 7 G)%S?:EAAR+4O#"]9NVHS5%0A033D_+)DR2Y+RVU. $+.GO:9-O5%^7Q3<5
P3KPZR0OJDY@E0HMWX\45DSQ9MZ;$G7A_TXQ7W^JKEPK=T56U3PC(/7! ( 55U[L@
P^)4WP4]C?TEY$TOC*\NTD43$\9Q 6(P50"4-3[O^G.)_98!?:U1A6.'R53K[!9PN
PBP62*>XH+3<&$#%HT)=Y)&A&N-+DHZ/&:7M4 ZEUI-\YZ0BN7/H%G$0))@U_S_=H
PQ"<59'5"+#HFC0UXA-$0H-/*C[#*8ANZ72 1,_?J.]P(1;&)F^@I;R[GN$X+_HQ,
P+>=O*NY:P4=&2TBG4SS:;_+H"X//^0(\/_PQ%D#-7TY(]\QHT"70$7$NY".;_:@?
P"M!3^)FHP!WY)( _ZZ;2/OULNZQ36U$D4:MIW>QN!:;WNBX'XJ\F@6EXA7H5LF+9
PZJ<!$+W]0UNW:0KOD<)9(6M_!-9%;HCD/BJ V!_'CB:7@3<_5]*ZVO2PR^(SX'DI
P$@U73ZI>ZZ@-Q&F$"<BB4]+:K^)?8(-G'J.KU[.,ETI0XDPAQBY /NQ>'2]'<(I#
PB2<F9O,U#SF+0"X)# 4+V?JGQ(-JY(XKV#!5BM150C2D8*QFS]NF6$RNJV\'2S3_
P!* 8O5W_',B.#Q-;@?'A4(7T/?AVK#@5*T4];S1?>DH(QY^!8R;Z],U%\!$.DDH$
PB*?#Y<V@5WK+GVFQ^+PC=F4R+-$# N=14:R)Y>?N$Z>\7-H0@^\6,'^LNH1Z_T2:
P&Z/]@ M@>(^\^N=9RB\\1@3X"J*8YAP<0"5*6S&P2R)4F,^,2/6@FLA9J[54(XK?
PYNID3> _%'!HM'DX$DW"HN_16NX8(N< $Q;]/?];#IA',C (JV>E)4%2,>[VO<F;
P-MFL]KBH-C$WB]SL0$$8CNG<J+Q@7WMJ12+W7F38[Z(9-^O)O3SCKY3_<!+1D.FF
PFQ7\G1;V5=:@+G-<03Y&KLYL7?-6Y_G+8LZ!4,E;JI_ZO//X2Y2;T7Y_]WUAA+)W
PIGILMUY11!>W_[OPN:D[IJA<:W8CU#J1P*I7VEO=4].(L,"2Z5-9':=D?.1Y,Z5"
PT!<R.>Z(:..2($@5"AJVCK! .LA,LD*7)['4F/N6>?G[" EJ/80)K$2]CJL/<A?$
P:JPHD,U3=H%Z18S08T9 :Z\>G2EQO2H7K/HGJ@ZX:G<H3H]);A_ORR[HR[:WP_BH
P:@HD.%8'$+=<<+HSK:NEU3LZ^.V'X?3OO%!VB?S8CG4,#Q:4AZTL82^GP37U$MV?
PSL:;?M6K?A3F%D>].(6^Q4#-'O]0V5;IWY>H"H-N)JI"W$OE=55(G&-!O8C'^)8^
P@\34.70_GN 9E1(R/G'X#Y8SC<](7M@3)=>VNG-*H<@^HB(CF,R]9M.'=MM.CJ==
PKB,NTYNY++UBK2QHZIX8Y*$\_<CV*U60EI4XJJ:BX&4KS$Q=/F(OCX9QNQ4@@Y?\
P)>;6%S&H,+.-PC..D0 Z< OAB3K50U=<SBB_GH$\SCIJO"*_FSJR^R%(&\E!B).!
P-Q2/!-_IW3Q:S\&M5&(8-C0UD(6Z,O#\.G)I?S?K"<?[$@=&&89UWLCDK (7NN0?
P_A4F'7-"/^ET3PT,0$2U,?+EI EB;7Q?FNK"@S9R;SANR<P1CU!TQ'8H4S&M%>5'
P+RLHY[[]]DT(=TRK'>7E2Z@X6K.Q0'3"*UR51K;N4F"<^)-+0),/-02KD#+2 RVE
P9\QE&^5=11#F2&"E=%?0=/)U?+.P5\Y,E/R8^F)/]0V"=7Y?%<Q-T6?2\TS<"XQN
P ]7-R0>SRB];HKDOGB0!>R_XS9!<VLGE>9XG()AT;@0V_%4X64NW_:::T43(9,CR
PJO3<&#^0+^X=BBIH BB*)O9S;F&DC7S>_![%*(NO3B,+O>%^WB?9YF\:_-D"LQ3^
P[%?X<#9 G@D04&BLO;L#1'IXG]R'YQI/9U5+R[DN:E]YD=Y>4/#""O[4^OB'R20O
P5]>*Y/S,4&1FEHK3)Q;J<[,;8_$_4EAF&$]L9)$(T!\]GM&]^5H&F'6(8N"JGNDI
P):TA08TOY]2K350<@6ECW6N'7(T*BE(&4KS(%:\..9)F<4]LIGY?E1VW5-M?2Z^R
P9(\E!2-85(VCR':!?P]Z O,* W%G4L?'V3.21\?TUY3&@AS+5("W@'SC=T+@-U*N
P*K][*^0Q5>$ME.5^/X2=6"!@087)52=Y>ZZ-5E3G+\(\_U8&$1MUUA#]?L_@CKN;
P_LJ;CO-6QCB\3Z7M0(N'PXOHEH,PH^#/(N(JET](FFFTF\\I'T5"=CF*+@%5$DUZ
P;YKEH4JF@^YPNZ\ ,;"R;F; ;LS(*VO&&>V7##E0RP$MEFE;ZW;UILPD8,WG8<%U
P;/'G1FFYZ1\&7]6X\FU.U]M!T^67B5S',IW>1E@W+Z&-H37&+\U[@\2]!5*\"$<:
P$[UHL[\5<@7_O+$#OI5YN$I)?C]C4QK/5_.N ?GC*-?K)(8/NWLQ#J2'YG*Q=#$B
P?56J,K^@K:D?;R1*Q.9PEB'Q,AD@J1/SLNRQX%<$I]R/+Q8ZI=(G=@)>J4GMSV0:
P_)68AUN%V?NZ/#ZMQ&M1A,OBE07/PTN Q"',=%^ ;+<]GZBQ+US]16#1^<YR+N36
P@V+A)EYC2=8;T-2[..STFH97MM%V(U!$[0>\-+TZ&RP6K*U8J'&UD[95?W6.HA]T
PYP^1CF3@R=ZPB*.!1Z)ANR[U/:J/J2!XCGMC"+YI"0\M0 QHS5R*/3(>-OX\? *]
PR[]SJ.9C_-B>F=\DM348J2;81N3[O.Y9Y:7N^J$!?7]<\*891;QH+SK*\WI?[F#M
P_(E!_!SQEL7O50/D4#Y%J*^T8JJ[3JF<+1;W&W,2O:AAAJ)4'6.*\#HY^.?# M:T
P&)(GKF7G  HU#N,;_F%LZ^6=;S7NQ[5O<XEH2*!K= *VHYHH2E7AL%?1<A?R6]52
P^1V:7HW6FGU#YYS.L74827)&XT7/%8O\J3WZ61>,HMB#E6,=IV #_Y<9+E/I<#TZ
P_Q5!JL*? [HNZY;!M2N!%.YD\:5"GD2E,.D1T>[&!R4VY2LCZ*XL>+'Q_GG?3>::
P&DL[K@3F(7B4B ^;YK1%\0H NH7-F$6&7DK:JAQ:CU^_L5WX.J^A/C$.?C&&]7/I
PO<,AS.O,!ECS];I1^%<"(U%<\B:NY3(( G VXAI0:=1%_'14_I'=@1FY/O"K.0K6
P>!J/;JVJW,1"ER5$D\W\WI:&FV:Y8!\J'1,:^.RL  SWUV 4J=AC)6J&".R&^:3K
P$%U@.<&U+=2I1LF)E4?C5ND=%\G]/YJ,"A+M,>COKI'!!!U^YE,Z1_6QC[6CNMEP
PG<"YLQNJ0.[EB D-\W=J0YX:YA2BYD''=.4X@DE5I>;8X\S]"3[@F1_QNI$.J^?>
PL;_\ [>S=6>@#C_L5FW5/40H_4G9;(+;SD37U8J9+6IV#2&PT J;$BH#5HOF>0*3
PUE/E;[7-,07BJ10Z]7O#ELG?%W@31I^3$WRTU<8^QF[.&0,'COHIUZ#YC<:-O?-S
P JJ3*.[/+QMM'\MF.ASXU,HLX.!=@?8>F>CL*>TP2:G!?R)]4VK4^&R%,@22N8Y@
PI\2QO#1(5+=\_"-S.BPIAJVQIA0"ZLF$S7H!"W=U0WI+>Q/-&N)6[:<@!09"%Z&)
PADN0C&-/NYQ&!N,'K<C7L<J:#E6F*$GNY@N#CQ D23E 9-'M+K?#,?M/D*P6,E"'
P(0MU5'CM-\K!T.+ L[,6R6]/S3<D.@>_3/6U3?><9&DDUWOQIH(M=<$($C,?I \F
P6-VNTJA;-PP&;5CZ'3XOQW_)^U&9;B&T5%B>O0V99SF65JMM[EF><DL"QVEZS@\Q
P.GKGTNP [%.S:/)Q$M,Q5,>4@5Y3S2JH3K_.X=-.K>\XOE60"\OUZQ/7VL2[_,F<
P$ZG3DHF7!=82F$"OG=YHV<<C$$4668>4-3$#6IA1YI\UGCS2-#;]62?2^%/MYI9?
PSBBH9*??:Q9>==_@>FC7G\46B8*31<I 4[PC6EK FD13:@A.+7TH11$EPTWX@L_L
P8;[6+L:\BV3F]R8#-(F[39;=&."'0M@C<L<7*N<6"*1:1S&D?X8@ @8?21&%+4,L
P;6^]8.-],A4OX,Q0TYHK$.DCK !T[M%B)&@:!_CA*8I62+Y%E+HDV,9)=0-$'[#?
PYW /U1 0$U&P+I2]4Z9;++J/B=:C]Q'+,Q:]T$S>AJS ^\#B[LX\9C3 &(<)GLZB
P&9Z#H\/5EA<5W]1G(-\(.B1A1 B;2-*TBLBS8+SWO)6[+&8@[G)2[R:W'?^<EF9T
P/7@J-UI^VE!Q"*&7=A,2TNG<)#LCF<6M:+\RDA77D0]<;]Y0Y&L'HUO5FB#;)4W%
P-VR:5AW#?9M-#/'5EV3LZ8SHIL1^!5F0@<'/$4%F/M__@T-O\SR#+>&80Y@N(&$$
PG/'>\C-OFN<V6A)I!Q/ 3<"!/,9\9IG7])^' ?=\$D/L$160N5.Y(.NR##N$'],$
PV-[%4:GE8V(/HJ'JPZPL&VK4?/Y5AG8YPIJ]:CN)]?RN> N0//PUD1XE=QA'\K+R
P<OVG@_S>TB-8-],VKDC'@IUB>)40P>SA]OJOIWHGKV84=.EQO8'OQAE+R.AK5,+=
PWE)L(_%!/'J*!C*TURUFWC+$/R)L28NPH1,)/),7B]&8?B&\1Y+@XK+IQ(D_\OQJ
PT8YSY_2_:/GUV7*]7A<I*=P<J%+]80:H//@(%DMEE#SS+>+[C(@ /AGQ>6\>0Y@(
PK_PAT,^Z3\N7,[7G\G0D5;75/MHTM[W;QBEOJ+NJ8\IN<*]1*60OZ.*FY4GQL$E[
P;^W'TXHCF4NUW!<2NYR!K#6!=_F!VW+A_'*3Y=&RMHZ5@9X+>DZE9'X;_4$&Z8<7
P):M<;NI["BOG]^[[8'A@JT1;<ZE0_.'D;353GL'@$>J5!I0)=%Y-4#'CY?SB,O*1
P?%36K#CBZ"Y$]SN?MG7)4F@/&J">!-\F857 >*I'8J?36U$K6,34.,YBXP_/75>O
P=YHI5:\JA2]"G[HY/WKXY0J0_3>9E%0]-7B*WHU3M85@"2CEU'(JSVO=X?JU++!A
P\C;K1MYKCGA,F?9MKX44?EHH;"YF)2V/3B&^5WDY!W4H!_E!0&Y/YQ^ED*JLK.LY
P4T6%]%+ZYW.#&E4+#5"V,-M:E'^ '_\:U@TZ?""YIL!-I]16BGE*(PD:9E DPT"+
P<T KIK$54H2;,X@QMY1C1E,!<^YJJSEI)Z/?D[:8<L,-#M-;4-( =65W;(D?8[M#
P/0%AY&!SY+_VZG?&V6$8UL!ABZH;X@G_^(F&QR^P>7OV9PM7B>Q*EE@NU&ACC.9Y
P'D'_2."DQG0B=<G9R)):,,:<5/F7A>?FW".1AJ]$UYY8B[Y]<YPG/3E@<$>K?3>+
P?K&'VAX@'H$O"HTM Y:Q#^<?NGF6F/3YTMGX+PHKQE:^^)F9-UB"?H7!)KK7%@0M
PMPCT+>_=>;%<I%SCP#(VL[?39XAI67VZ_?QM>]39L(NH5O:AM&Y'R%/M)?%A-1/%
PILXAUF/8B*X:/K>O_M S1ME6+D&Z&"B=2]W-<F7H\. <#)-3L,(+;)?V<C!(J-4R
PEFJ8X^D/C$X_-J\_!>&8<\8:[^I<YS69\$Q/8SE4A)(T]>F)/_:;U38CIK]-,<YY
PZ=).]-/43?V!J7M#14!^[(1,9%67GW(=":R<8IE^+TB@4?YT![!PGR\[(=!@U5*B
PP F_G8I-3R=U"^FXGBBU,1&C.[A0]/,N.0#_/'5DJA<OV[YPZ"^27=3-ER1?4&]&
PI@SW2'C'A#MZJB4EW!HZ=/3G>D>!!X3.-"OADD[0IFDEFN'0KVT01?DCJ?B KEF.
P+*;-]OJ$]K=!) I>0O6X#E0"304L4/>,E47QS^U=&$/6\X,((_F'ESF&WH]Q+>W9
P&0MZN ?[OOS=UV/&BPJ?5G!>:M:??GW8,"<M8B<I]AB6;34',D NO_#C/23$J-$$
POH:TWG+J@3FOD!/A*FY8H_-JU\84DPQ@<^S>O[98$W+Z?R]/2_&K&,SP!;ZB6F?'
P)"8K)*^DB9,P53B\H3*N=RL!9R;HYUDKCE?Q4.%2#L"$+LY!$IY@8/AHN!<;5]CE
P=WI#@R!87#/CMBPC%L>Y!@D43S?^?[%9VFAXE!MG/K80)IEQB?](F*YIL2R#!%@@
P+@"H(+=RU)'/?$OOPP>,-'C#>UE9-#'!)=? WB#A6 K?Q>]% '[Y&6+&$JUHJU\&
PS]N*:! ?^:)1RVSB327HZ*"1F&^UJHT-6*WP[1SG)@\4H=(PTJ_D,TBTIT5@ QCF
P$*DJNQ)9W%>L_%1FWC9B^OGN_@,!2V;211*W16Z2G@))A9.QVDA]JR4S^HZP"XX5
P@\J_83%5QEMR]U1MTTI[TSN-_-HJ2+3S6#'713AW#9^4/I<04IMED%"BQ%4UI(X!
P>7=E':53Y)9;0GO9N84%#JG)^@RR4T.0_9:@(-GZ^ZJ"/8F(PLR$49O,J=,*1=^_
P&AD*_*$_,] &>+SGX./%39R,I -@M':IDZXW3/;9>^:Q65@E0%_]*1'V001;$A9T
PCI>HT8"([0=/@2-V*15^PGW0F> C#'(UL4BI-NSI4@'02U."O,BCK^1"+.:0:=-(
PE^;G=')> J\_PA -:&.$R-LQO#$5Q#7HJI0@FLKS*R<A)A^"[-E M]YT4;"NDZZT
P7 GONQK\:$:+(Z?D@\UVG +IZFLO=W^[,HF+39$]$$D:6C)OV@53_ 46!"_$1C/F
P7+SA$6=V[#D/5,-.5X#T;JJB:J5$!/>K#=K6\A1#'&^W%09:XQ*Q15"5'O[&6Y>=
PL&3S8C7*>)\R4N.PIKVDZ/ 6RB5#!XF%11SL*?/(Y=?+(IQ-3"_G^NWS!.6O ?\L
P'G**2'9ED#&Q.'<L[Z;61L49)<BZNT33Y<UMO!M&I\2(DK'LP^U9H+'#>L3QQ^-S
PG:=9<]D+':FNO.(4&F,L\][LG166I,)E%)S.E"J+8HUD-9'.#EC^%LD#^PT;/,S!
PTS<0F4CT:_WG,@6MJ1Q\4_=$R.&T#,QCL75XZ9[X5:Y'R#)JR2Z;#L-@J9DQ>A7J
P$4FC00QBIAS,Y-#RK%N@@*,5E.4D6:GH\P3(^_Y#%-?:(BQAVTKGS$LDKUZ\:=/Q
PR';I^*K>;*P5/(:-!T$;4UM'J)%&D>7Z]\C">H/NJQ*/HJH9M!(88^$-,L'03*]&
PN=2U%Q!)G\7S!,Y@MEOS X&8U<20@M!V@8R/DZ:IU9ZFIU;3'][,)M'H%'38NQZ$
P<.][W/,$;&)9)%B;6%(-1_4^)OD!2@8'L3AI(!AX61+9BU=MB->*HF)[#M_EF[.&
P.2W57['I7G]O+1_1TJ0"#<X%DH1)2I*4N9,Y^6FV NB XQ^?G4_WKD/%UQ?K]Y)A
P^[,M=/OCBYGHFRC(:'.^I61A@OZOHC^^$QQLJ#QI 4G;+X"VD:1,,P^T-WPRCC$I
PW2,Y.CJT[,6XQRSSB>)1YR@ 8-\7=+I$'[9;K<;%W@";-=C5;,1*>6ZX[S;4U H+
PGP-ULRS@WPI?8^Z<6F,W,L.EB7SW>LM)D2(BT]7SA!93WFAIG %G,T;#4241*G+6
P^_%2L]YUU$<.9[C=J+_.^1R68>*"$MK1=8MW +ZDLIFDR><;7)>/1)B@_/ .42[7
PUO';K&G>K:043IP=]59U"KUIJJBL ://<F7PI% 8&B0.%2D=*Y6)O_V@T*PFVIO>
P/P%"R;+@0DI9,CS7L&,)C+-U) 0<@P$(01WAY_>WSX<H%VPEC2#5^>Z+N=WZ&@B4
PDQ9ZG.H0CC5PNB\!08_H_O#?#^,(KFW?Z83T.4V9=LJ.@CTEQP#9$-&,R#T1BYU,
P6F Q'"K9<?2B(0B_!V+\1]53UHC=!5"O'H4GC$M0=+#?:%Y#?N6L_#<2L6'.PMI)
P=,OZL./!88E%FYF2>.B++5N"=JC">WPI]#Y'MY\^88G2)7^V"BQ3+2YJPV$C8GL\
PR2*4@)ZW?A;&X?SD3\RV)H.D=ML-=-E2%Y*86",W?UHR=!-@4D&O$C2U2.D<#&<*
P!'>=\0V-P:[*7+]MCT.]I!(NK+5GGHO7Z.RL@7:$@.OML/;/V-A6:E97S_$Y<AMN
P_\"-?;;N$,+=C ;[IXP@-R4F41ZBS@43^S<##M*P?/8WFUDY ]Z _: !+,E<%AH@
P&=TNW9AK&Z_T0E.FCBC9X$P(4ZTL+>ZSSL%'NMN_E2S/+=R%HUSFB/88<UDN2A48
P&^U4RVF6N0>Z#G 3JPPC(]HB3:EMFK_\F ;G"/DA)1<\1(M! L2EDKJ*?HD$GU80
PI? [9VLMF.$]T!,DU)=L(F(M J?2I6T)0.=Y]2%L?+DA?,G=X>/=<>%H9;*;,?JJ
PL*GOO?!5ZJ*QL%.AL&Y7ETJU-!^J==<8_T5VCZ!G%3\]8WV[[3>=?R+=D,5Z<&/8
P4C55@&+AEV>V]U%!-] 'EQ-=:[@]^&'S;3AUK=BARGWOV_8T+V>M+4EAM7/1&2P#
PPW_#=IKQD2_XQ.B_P5M\7JKDJ-SP/B@$O3I %N'V,1/X47;FJ%ZP.H_-^CLP\YD.
P>HXTQ>F 3/)Q=J(N.7&7XDRCM2#R-5B+L>'J&:##!KWQ;-$Y/?1'X/7U$MU$HV3K
PUT_7^31^--M#QJS2"#%K](6"\!,? >F12"Q'=B&:\JDF:.TVR!?,*0.Y*%6T];3@
P(0YT.Y3BG]\;%QE )<3>$<68IT^>^YH372X:EK5- W=@Q>10N:T#2'#?!B2>-V:'
P",3X!UH:NT!OWR2\,5J1OE+I.C+ON.PRD6#7(,6,JD7W(;!28&]Q?,2ZI>L$LD8[
P^9.;X>%;=_;U"7U?>_BO-0@]9T.N-BQ,Y##NL6IT>D9"2RV?D?*,4N/X:/J&D1*^
P.J6+VI:%3*7XPN0NEEOMJAF:16; $P*7%=4;[K-PI)!@:<.P)Y?>.<;^;8Q;=EG=
P5QC>O.X,_(/(.\EM#+W)4U0(38M#I9(\K1R0M#BU+6O:SQ5/66M+1^26PV/B03A5
P7UL9U+&:%ZP]UL/J,3=!Y\<5!8I_C [8,6'U.709?3U\>AA65ZFZ0#_3! SZC"V(
P!+#)$T&?G?V#VG']A Z[V/50+_,U:/3P2C3G:9Z*S5\QH$@G)4/U0\HE8<6WCK(M
P".["C7/:LC4&FK9A,,#D;7A:?FN.XB.<G\J)RJ?K#X7C]5R[V.D3N+Y>W3+.!C#P
P-RDH?[&^DRV+HJ[,B'+5AV@OP^P:>HRE)='G]5L#B_X/AD0!.??H((8'>.R0$T2W
PRR4%O-G0J#\[>01@,)$&N<L7[V@S1]M!P$9*I&]^]<$P4<,$#T1 H>LZ^B-&.+ZB
P <P:2WOL!7P,J^$B\!/G>34SBBU;OK)>+9,Y4;SXT @>LNJ_S]>+^]K31"ER-GS;
P>\\/"AAR5,P.EYTC40P:FB.%G.K+Q<N"3IR[PYWIO,B#K6^;5*W"LSY?27]*4]K&
P])3.W!1CMA]4V'JA;43-:.T7B!U(E!!:#%Y_1QT^A@CKMOCE1"+IZZD\+@XC$]DK
PY 6T74.P#LK'*TGQ#F%D@([-!EKF@UK1%3%KR-MU$4C+S [65/T[5#R_$Y0WB31'
P +!Q$K\6)NPWR[VYB$@/P8P9#?G)763G.NKF>@;K4@-R1A*H3OR>+7DAXU=O;<.'
P;5&T96UY!@HM3W&C7ZB$JP]D-G)8%'9Q^M,@$6-(^'9%=I,_5R, /8G&W'M:@$'"
PH_<" 417\#?";IG W5:.8+,,(+UF^V]# D]I+2@&@QBZBG9,!UI;9T.@3B5FFNHH
P!QJ*H"H7Y=5+L0/=#IM>RR^00TFL*;0-O3&M<3][*Y@?R,ULV:!L;N,#SP?DRD>H
P3E3#:B]R4<QA$Q(6E0#Y*3N/U,?,?QQL"G5;R'AXK</+DH"K\36X7-[M'4!0345W
P)WLK=EP[P%YJPU%6!Y#.$^Z>&&K68CZ.I: +<;R ,QZ+*TA'"S2/U)7^7(2D0X81
P?WS=NS'<$API'E26U::!9>V@7Y*F00@AZQZF&_E*U)_.DHGG2"-_>=S8A* G_NS#
P8BE$3-D1RR[1*OX<;+W6@I6MV:^6(#''$4:#>Y%BUNM7G-*,T[2>Z&GMZ+:X]^DW
PZ%\@Q8?TC6OS1W'?/\9HB8-W O4B57T-E]&M,&V8+?2F@/_Q  )@?UG3_I<7_J[&
PAZLMD:4#?Z,/M=.Q-TH;21A$95:LS[V>U%&.Y.:\BX8\VHR8$N6U5#]"'8-57,9;
P<?P&L;[Y/%VH%7)K$175+5[&)XWO/9I XH\CQ5K.@5'-B> :EVZ[RNIV!ZY7Z!W2
P127]__WZR/Y8N63*O%:099CI=?%_(N.':<*5L >%[J !-W3LM9/)Z'%).G?7K[=D
P4&="?%0 # I!VQ6PY&47!5@%A1T7PJ#3)U9'KWTSS-=WN6:/KNUHZUG1;&5'.>Y,
P6DLO<77^7W44*J2-9;>B#.VELPV]8B1<J^9="</<?E@'*GQ17_;Q<K'3$2XC5'F=
P5VL_J'<:WO/L!S+Z= 01_(IAP?7R>-PSRN 'P"EHCJ$R>AG-VQ= HBK+2H'P]#%[
P"MGJ'XEX?3L2[>AR^I:%5V0F5Q7$JF%QWRSY@H:(K%^*_@UOT*D<N-S]5W /;+9_
P9VN(<,@&O8-PMO>HK*C< VHF'OP%T%!=+DN)O/;Q;=&2"84E)GD8E6B68&2'VU/6
PQJ769CT PO0LGI&*DBE%@IS^7]?.OP 81N\3X6JC *6%.^DRBGAH@15P+[YNW?H<
P.AR<31,P#ZM/*%Q;'0_<ZR!,L%E]#2Y7?- P4?V>R\0/R(%RXO*GQ[I]O":>91\.
PJB$GB-_&NEH$<,QTK 3$I!,!G6T=61 >XWA9JY*6B4T;J-,#5&T0,'E&ZCZ,33?6
PB(<F3U]@EC8=JZ."F@87("292L\CD9TT6+ D]QWS>C+U--A<?'YKZSVSM^E@6><7
P@]&!XQ^IA>N\;P/#;7KJU3JVD8FRI2U6,XE'WP!KBG+'V8,T!]-7RQ105?"89-4*
P:/W2=!?.$8C5S),Y8*5ZA#SHG)]IRUV69Q^&C_PR8F,B^0'DXR<W),HM$_#K40P.
PC'<F(Y&QH;_>HM75KF_OF*SP#0&5-F-Y4LH#+PRXP&]_3Z<<3P'WS]EK,R9 2,Y$
PU"/Y).*V/*&QF)&=&O"8AYN/D_%KO_)"]ANZ7G":%KV'R$Y&+"#BK%5D?M\OB$D^
P7W7Y-23OSRMNTL<Y<5$5*1#: P1S%55)5>V=D7@L^SH37HV(2CVU*)IAURG'$@P7
P1$KE:\?*>(?1J65G\[/B-8$%WVWU327C?N =8E?O\RF8@42COT<4[)+73R\UM-ZG
P';64?HVEZ)PU1"XA-=-Z$JML!T5I8\E-=WQK$%I0T<J)Z9I$X@]>VRNZ+J>W@8=+
P[='#E%&:%-Q1F/%2:K;IVI.T?YHP_M-X==F?-*U^,RFOR:W>UC@^17@VR:\Q9 (O
PD8*)M'7SH(40^'139E]+W=>/"T="5I]55X)>X3?E+_ZN8'._38T]9[@DU]4Q]DM8
PB;THAJZ%FSB-_$P>W(PV%U09"66CB0M&Q(\'V*W?.?^O?.N\KFPS8TM>]&NAU&&8
P-ZXC)Q9\=<IR5)@3N  S><;>,>D&IP;N86SO<$,'(X40L:1=<6W8UW2K>!2#BP6Q
P+4]F?4D2,T.?RU65&*[M?9O/,DV>XC'*NUM=1W$D\XJU$T?[SISI)@J8Q0.;GW<<
PB)/-S^X,'?5%N KWVN'C?FUV]!K[O!P.;J8OE0^AF%\L_9KZU('JD'EH,ZW9%G#2
P:\(,3F:N<OVSK @I[;4 RDQOM0I,T-67B&7,+TS2:Z))E#U0GCB] %DB/O=AM--^
PX2#Z#Z!)!(=!SP^:KJB _.6LGH,NCY(]Q7T(I^!=;L[=+T$1_<CO@'J$I0SYL<_9
PJ_,.LZU4Z*4HUNZM])R^ASLD&QWWN'([+'HL/RYPU"EGK'C$T&_F?;G53R<&Z2";
PA]<('<H;?R$8M+/H$=-LXSP4H(_=7JEA (;5+E$C2V M_6"?V)_#]2-C"O%F[59Z
PU\_;^2VPFC:X#4"__?OA>LTJQU36^\YLV(+WS&@\4)QY1%/X&2-FU9)+D$<ET*8#
PJ/,Z)0]'P7CSX]48,=2$@C(<M.@#?NJL/V]:2_PI_^4;^3Z*J%K'C$JZ<2EE)1%$
P J&+=N(LYNYR?(\K#^H1BN@9$WZ01<.CH[D)Q%I%BZ:!8VRFUET&#*6'B'K//-4N
P9[I.E+GI($+?&J8,$^@L/"<3Y[NEP."?6&5PZ0#:@(\^')<W'9(:HDP1&6.&$MS/
P3!!=I71SR=//V%*H0L'X*L\,W1@0?I+5:[@Z; !;!Z?/!"0YMU[E A<R")7F>9L3
P&K^^[EZ.G@"PX<&*Q[[E.X((,1GQ78T@@S<=GS@%6$T7)]],3<D)S4&NX:+N(=]I
PG-ZNS3MNY!PH20E6Q[E .ULS0>BJ W#AT[MX4C$/?W:)85>#'1,5MRU-(M/1RNZ(
PGC6/M3.R(8%L_#^H%;\ 5E;;'SWZ)"A(@K\#6KDI^-9"FF*#YP)G3A20EUI$YA5/
P5FLOAML$E?/I7JWC3GN^#:VU%5VZR.4)8HQ+[0!=JK/VJ4J?E1WOZ7!VKL^0RL!\
P7Q9R95H[XQLGD;.Q/0.K[R=F1*_4+F^\^F3*]!TT322KL."9<"<8UW$4='#QI5+J
P5F)JJ6?"8ZLD@G_Y,!A81ES3[_"4,N,9NCL<*%A'R67B'3J=8@<6CLX6.Z:2A:ME
P68@*KP,W](:U()& ^,E'>FD 5.823KY3Z\L#;)]X"N&Z\PSD&3F8(K8\0FV"!@+]
PL7O'\Z<.>WXLE' 3N]F+@= 3#2\_!(_ 9U_XU[/.&\4_(Q>AMY0\Z0,3[%\B S6D
P*TN).85>#"Y^0,PRTK&EV5L.XBQ1R$)MHQ+CZ70+&UK"'?3)I,CMLML >^9-)0YD
P3@);Z@H+D,[M7T]+!7H($T[X309@<'5JI0!)HB+76-)#3F WJ%6C1%'2?QOM68HA
P/9RRBZA[_SLG-/].^2W K=0 :+L6\\HT0=63VC(#_AJHN8<S\F3&B29*:G[6\'XM
PKQ26KHS*G:Y8L'Y'FL:)CH9/9K5LRI]-&[9UX 7&G/;U2V,X[1'.E_+S[515KQ/6
P97?$U03,>55%XBIM<3I#;(N@2 *3;;X:5U9F1%26@ZA"]+V; @$E]$QEF^L'PB_%
P69;ASS.>NSPQ5@ DVP<:TS#7XBM8T[Q8X2B70P<H;:N1DALM8()7AWHUM"^.TG3_
P[9GH-P*KX<.Y_,<=\@V=O+0=L<\PN?RE'T $RJP$M7T%RE+V:P'"$O\?;SL$G<2%
P#/L78)J!JQ-^<_J&^YE!*^ZWI)CU9_H1/>9L^$"73!@%Q(_YVNQ9_5.B?Z\69J/C
P\FC'8E0$/#,!O=]!0C1)\S>S-1@[Z1J6^2"?&C0\S/L&:)H_/.&R&1N9/8TZ^O:Q
P5IB)1-W[MC1)8X&;F6#6;_02-MR&\<V1+#E/;-.M9E!+=[4GH"R]"3]DA$WHI<_8
PT-E^BQN(+<HM&3!J21G!DB9[G5/$NZ\4KY\QQ(1S[> ;JB@'LY^?$0DT39\.'^/<
PW%/UAH3RED/T.3[JQ:X!-DZ.?['#I!?M7"?RVCB7][9Z*1W0F_4'H[?79K^]*JK-
PLJ&;6HU; AQ&W<M)]_Z((1PM2_[N7"Y>I.EF; S^+ \#%P-:_3*HN=IC*Z#?XV6T
P?/8P^_Y(*.X6\U+4-ADOJJHTO= #K2O]V]1,%<@2N:=G]YF4C-H,(^G^:9Q3W4T]
P33C\UMS],:AN1F2OV,@8XS:=I][VJCMU3[TD@LQ\=<6/0;]%V<KTUT>XE>-;R58"
PT@G++"G(I"!QV^9&.TU=L%6B8?.FCU1NK7(5NZ)D%)P)X2RYR,![<"1266)+\R'B
PG%V#D0IB0V0?G.USL_\I$FURDT,,>7\LK Y'3TN93!F.,BA>P014H3R/LU=LGMLH
P7/]MI+IY,JB*C-B-5#\L4^+>D>3UG/C/J$G2>/6-_B;\(%9*ZMOP &%;#5?$N?IE
P3;2@)_H!#G0HTOU%WW2-YHQC"F0SF\7A4U\E#+5N#(C))BQ69PHD;Z%E[Z%, -0:
P4IOZM%*'P*5%@NF'4)- P/VDT\%.@>"Q%T<:DH+#U@8!>_5F:LD#)S(-\DE$'+ F
P%M1#+Z.&<X3A3YPC[?*5!UPV4'3:3598Y70#7Y+,KT(&M19Z1&V7ZI>*!6,T;L%N
PP^E5J@DLH'";DH\A,S:M-LS@M&MWG40ZJ>0Z(-RBYHA[P1D.A*@0^A>?XB*>LD$:
PD"39(]NY-NJ[L37+8U*KHMRP.YAWF) !M2*R-<0''@F];6F&AOX.^GVL_\PJ0:6D
P@38*$0+DW/D3T *CLUCL9!)3A]!:G8AAA$Q28VV;>/8FJ=E,_G2;2-':*BEH F2&
PIE0$+E2CQ%[=#WZ>0\Y/*.UP%AJ"3=;D!56-=Q:2M,R3N-"31ZR6[=TMUOGJ""G;
P8!TBAZ7==ZQ\%3E-(+FRCY;R4_\6W@?N<$^E/DF5JE:U9Q+6D9#?Y:Z=ANV"7N8I
PY)6Q*+5Y%5XVDMJK0_?JJ@CQ_NJ,/SRUZ3?GJE$4@BPOZ-$*@)E9^.R[":W71/Z1
P-[,JB?K.J$LUUF?H9:TB'\O80(4?)7ZH(F$QCK+";LCD)34#5_$Y4$;A4!@IJ)+0
P77[.;!D?LN$'BNEO$&/GE-IJY<3S.WJZ[.1SK!8HEV>-,J]7SB.0KH1;$GR';16M
PJ/P=@MG%U9"6D'(1JWK]XV^$JC)7V2=3?0_:<R M QA#Y7;^!-W')N-C\ 5RHUMH
P8:'5@2"WA]'*"A5B&8EOGB[SBM HD#C,Y_;?LQF\5"7UNF#J3NAPW=(<F"7+"68U
PQURUVS@H>BX'LEV5EOKX[\!7XU6B,T-@9+;82[29[;TA"3,_Y*BFGK79,!(;Y1.V
PK49O=\7PO@QJ[U[:^O1KBIT.)V1?S6W"U>%8UZVK<&R;HJ0]E^YT GE^(R*KITX]
P/H RV@5WJ?(/;M#140NX#\^2P<L<6VZ'.CT%?E 2D@K3Q]?8^ +\Z5*M*1E2:G5M
P#U$'3'KH3%5ET0\%U(E<!RN>#$DQ@+X"6\W/%]#/=>YF<]SG5@C>N5#L08N>":?=
PYBLA[RBP: W;GX/)MR<TXDQ%#R_4N-R(D!]D[\YJ:K>B;/Q#DX*X,3+ WR"U.=Z%
PG.:?Z]'@*1;(HM06XK.G77YGB.Z^\=>V%36($O1VE;"/4A_?E>"'_9SK<MS'J<+'
P!6U0X(LE?2+_=A\/NWE0\USF[U>@B!&&>5PW]7NC$7BM/PWV@<.QO[4[G H#K"NV
PS.'HS?P,P'BVBM@TNQSP"GD8C2WI>X@?IMA#"[]:^>+B=N/6)QD+H.5"A9UDI]*B
PB^\/#7Q/9/4HM.)94,80K*9QULA7AS2-:$<+BP\L/-H=#\:$AX,&AHV]5C8-*?*-
PL5IU;D>(&JL%GLM\\ID+,&O?-FO:4W"8FUV#%$0ZY3>)$#XJ5"A[[9/V0F=ZOSUG
PPVV7J/LKV_&2<?6@#">;.9K!OK<M^_O[,Y93NI>P3 DX[.R2NC-J**.*1"@1ZA 4
P^\8UV6B74$LG9LU@F&,^Q(, EVR4TB(@^7M/4PM6F(G+%C(;RC3SP"W)[$^JQ,#4
P?2>CC=U ,):6;<*7B[[0=@FQ3 Q+:SJFHGL9)PE6-S208A=-]->J#>@K+ Q]]4QI
P&KAO/5V+:G1C&.+$K8C[-%'E/PX/BFNLZ$UETLOH/]EED0'3*#?8*!K[M?'9MT3V
P3BXP],)H!ZA="^!0/T6[:Y;^<Y;Y?H[ 95U.""HO/VM^T[(%(D8I:'31<,W8=_@Y
P!'@!RG*JD'Q*PSBG)O[2WG]>9\7*DVDS&FD&A]O?8TTK5_+T=NSD2''XH??C!\2L
P6?QHS$43[#E@A-VRHTP2LWZVF#&2#\ DO,GSP6J<5<8[\0T H!!4%BX']9!6@/=/
PCA6 %:,.L,7/<6EGG?NS$9^68V80)!JO3V6G0K*=+ZDV'?N_()N W5@[)P9XKEGM
P>4B+,G"+TIYMR4Z0,80*0M"2T<">\RB]%UI!WQ0_\B..<R)IU4+HM#^"XTDYH_=$
P2"9>B$1*GW2C*69T"C^AMB$7/2R,AX?ZR<Y(,?0PZK2G5P[CF2%W_)K$F%9WDHQK
P0^O^GH$-'X8B]7'P=,*D#6#5S 0H-G/1G0DF=3YJA"PMF"C9Z'_XU3P3$M3IY>'8
P))#9<85J>R\.H80ZX[\]+XYD+RI^"0O5O>@B88"D$$"=6'X@>(!(JNY\#$#DKA7(
P;MU3D*O,$H=J7J%P08J21J$=/IM]N8*+"Z+LW#@6B#%?A!N7V;=6Q=3I:L]6Y1G1
PB=95!$[!?9PMDNN)]X&L+4,B.(5=S+P.ZQR!1\5^$M\EV^!>6ZK=Q"EJ-700QG$:
PV#X ][Z^0DM=B@ :<DOTG8UI5XBY,%VPQU_ 9K*<J.QH<RRH.#)Y$IOVIUYKS,XH
PO[6X!\/.>X(K.K_=LRB-JD9[,6%.X0-2AU#,+NZD*+>^C@_*";6'LE]:I]98E+^1
PD*#4T[T_NAI88E(WLU#SIPB0:XDR8_>]JHROI9E5?#%% U6>43TD#6&&_*-4]F+M
PPDD\(J+GI1B:P_[YI8@[_:E8 R_L,;O3\XHG I9ZAV7:XKZ%[ ]1PA_K/9TZ%Q6M
POW3_ HZ!T9GK/<A*Z_&UF^P#^\NH3NUAOU67A*-)> $G.J#TM82B^D9LV<MS*[8T
PC-QFR'8JN1!XX*_!_N1NZ&:NY_*68Y1[*LU</P=1?;$#F4 ^-?-,6&"Z.%AF4+#%
P,\#QXZ=B/ [J$KI^=UUO649CIXA1)8VWSN\>RCY#ZH0_@B4!#0RKQZ 0K$V<&20"
P3X@U%))K>3RGL1KA/%@;"N;2;E:F$+QEJ, 7VH:G]@AA"_,GDP_&BX"%NYU?E[V$
PVN&Y__O><6;RPT8,A:]WTZP@Y#DNML1>BLP;Y[[/CR7,#].+=^8+,-.@5Z4F0B6>
P+Y>*;4K&F8PX/]"BH7Z.HEL?5X7O(3?%HO<C&1IH8<Q3KIU.@5KHV)RO?K/N$,M]
P9!>.BOK5#%Z M!\]5 G]V<QA2_=PPS<OL!Z7S&6&_Q%*+>FM"2FB%LO.D4^/;3@H
PP6TQ^C'><R?HG2XS!CBVH7B96?Z]NM<^?KPHQ];_51JPJ9#"W,J<!VE/]./EB]Z3
P!O4\>RP!^# H*/*$?8B:Q^-")*?VC_L6>F286)0,S*IMXEE#NL@[B-,,VY&U$(6[
P<WBKGV0XJI/X;#**+ PE%T>O637[&!46*;WKI>0W<MQ*1LJN7;X#*7"'._CT"P$I
P@$W%26FC4>,B,($ZT$O>X,5+N# ^,3?=LP,+TZ&_PN"+-FG(X%,4VH;-B=J+W7_Z
P"AKJ#:!'2[_(5JR&L[H<^(E_F*#] KBTE-" 7SU64$J-DTS(@..HB(&E33)4_+D:
PF5WB1CURNRA%(& GH3U#-!4X'0WA1>A]B4GC":B,[%8UF_S>O;TWU=XH6#_+F88(
PEBN'55^X P*]"-'PQM02O(H($3-6A!\C0Z=*+Z5(_N4NGA#36#G&[MBO06MI7O\S
P,/ !:?7-K=1@M+,[PHBC!O=BLH$C%!YR9IU0%V:4L7X4^TF@1O MLRG]3F=(WW45
PDOL"U&LM)%_G6:40"_09C"?IER,)HOQ;HXN[O#A0:_/,,7+6+OC]#FK2=!NISE..
P7!SM9WXS736 )?*;ALE]B[6JE@Z7LUC#L+^G@"0\.9C>$E!&[1Y/LKSBKHG#WY9B
P7SS8<QRH@BSQD79PK-2C]3]6 J]"R-9H*C;J\U7"=DP_6%63/+I4G-<R%H$ /'R*
PA%1ZFODCM$_]36;*LC38E-N*8.0_M+KE)OC*&6NU.^(E[V3>)%.@VE081_E6AM_]
P.6@SD 4W87S-!..%;D&14!_'3/H:*[SBUE7/]LL4,W<P2]%8*)B+&M+B^2I;P[.'
P*4N[V5^;/_61TY]3"5#3FO,!7%O,M"H A$^X$V)/D<?$\CGY/;\(LWM+):>'&OR$
P^E"?E")>I6 ,S*3.QQ(X#MKV <B=N7"XKI4X6[^?@4X[I06V4CLM*B=7G9*-3>,.
P7]*GI:%/N\<USSY>&?J@/":^4(7.-K0*61P-##$T 6^]._4-G_@I&IUEN01J#8J]
PEX:A,&(D#2Y2 T=[1T&VA>7"5Z*I%ABZ"TCNJUP[4;#7>639[MWY4Z5SK:EBQEF#
P$CYF 4=SIN"9@*IZF?>,6&C83&[E:1T8>%C&;J@*^#E8RW^M'AD)$7U4]H@39?QB
P01^,CD#';#,_8+6Z8TW3DUF-"6^18J,'E_.F?WX;V8 T,D\GXM<K3 "F#]L+J.LW
P39/AI&B/KZM@#0VL";-*PLXT]!ZL<XB1>!B0BYXW)U<A8P]5T(JPTMPS0<Y%NW,9
PK&:DW5 F*."ES\+ OU^,5]%><FX(^!Z2?G^FH*>\&%[.VJAY__:&>6&H=[\G,-.-
PF22]N4#@Z A+CLJ7O&"K$GG0S2"<,K_-M"1O7B?D&LRWVE@L1?VZE#)M$@2WO^$E
P[Y!TD)Z%R:\.GZ%+/\R4W12]+O!&T(-H!-J 0H,V[R1-+,((D9/9460G+)M?<5X;
PHGPX ,>BQI!G_7' ^FAO4^P]G#*;M>[-ZQRJ$>1AIS8O3T<4?49ZA2[9*?CM]_O<
PN/24"'.7(L@'"5VIK-7W ,=;HVQ1U$NJN=-WZ,C=?W_1,2;2(?W/-;(R;2#%"^+5
PBTJ5);B&Q)GB/)';>1D.5;_)T+#,U']J",R- ;MXEN)P"V)%!9@YT@7.+%8^1'!U
P(%B1,T!'LOT4P/O1 Z0VD@ODK&L2BEH%M4.RKIWQ09W_?BD+?NHS%]P$J&1!.@\'
P7OC,[<#M=;*Y1G SE\C),S"004#'R(4:!^#U@<F?51DB) D9_"69/VX6XDF(R'.,
PO0Q+CSC(DS2\*RR'8YJ<9=TMW!&_C7\MB/(>>NE?8Q$VWU\M&YL\"@&VW?/S-N5Q
P"W"]C<&GT^?+](X-_C"YOLD^744&"W!D*>(D6%BEJWQ$8!XAM6T[>'ES?4,O,V@N
P#?2L>U,G/2?W$O_B=1T,^:A>Q?KL-#"95^!J<WLN$\:@C?C^W&H$K1^?'[9C5=7?
PZW%HR&CS@PL1A!0![AF+SUNZ70_IY.K(9N7 >Y@3?\H?DHX_7AM48^%\S(%? T>2
P\Z6@GG0(69FJ?FDD2A((":A@S\51G1558,C]\RI?'3X)B,'XA>GVT5*U]XI1H"Y2
P0,N$>8W"WLIM!::81)1QDK>6659'*".E/FTSER?"[9.#E2LR9<?\>!8S@Q0^AEK>
P!!*(U'3"X\EFIA.++UD_PTR9A_="X&$<[P52[AQ4-1&K^B<E> I?1"/8[>Q4Y3-L
PV*@UE5J:),;US($'D!%J4'3UYC4S,A967)'/\1'A@(\#D_969Q)[),RP#+6'-)+[
P?UJ7ZQ\B>&3$M#@VZ*?6DD33!S6^QDL3)Q '">Q(OA. =1'7H%4.Z9>HB7IQT8R+
P(TNSAC#^YN&P"!1,E2.B/2\/"<(;@A,8%KF;2<W&])P0RCT!D&ABV:\'R*WSA_?]
P7&4*Q0%TP>,=@(R)F',X:& #*17\9X_=>O70F7I98Y9DWJI?+35E=!42%73O%])R
P K?29*?8)V;4-#-M_TZH@A?G*I!MYBS9VW4=B+*Z.UM_:0I;<A'>I+(P,U"X68[W
PF^Z?,5MB-F\+9>55R>'5A\;=F'!Y6B$#W0T^LDT8I-X_6$S%O'8BJ5$9:8[PN3(2
PN;-7Q'+"9(F,HNQWJXSNZ\>=_SYTZ$Z<M]2\]G+?$P-45D.+_V3>L2], )I;LOV"
P[4#3%0Y>ZU^D-<-UUU?B-R$X;9BA(KFACB%@V0@D7%)'RM9C6AGI+?P1"!S;C<MB
PE7"YF4F)*9W^V>VI4)H16"B2OXK@HHWP/Y"4C28.%>NY9L]SCO J^X*BK'!@20V,
PNH8:G!_0?GMU4MAC/7(?.G0PFNAS!R@S'D7!=7=88 ,).Q*M&6((,'(17NC";6=0
PFW3XO!-$^9:?#LM?'!+K$09K1]/Y%IJJLKT$%(38) ;]8&7Z#4N<%3$%F[G\P>B%
PUE:B=E>\T]K9XVIB7HTU"WBU*:>FCP@,WE*L,L.;J(N;XZ6M2;^!D]I1]2WR&[?-
PB2BDSH$.]5CTLJOGZK,,HSQJL-G%Z\\1]/47#>;092UI_K;N_ZMGWQ[ E^I1VA],
P22VST_# UKA\VQP:F!D $VK4AY\8RY?2X $O<X!3UK074429 8YN399D0/_]YSCD
PS$^;%1=MO9;^AK7U\&C8<I%(FVW]W?;0%3#7$D^MI3 :F&ZS((PURP*-I[ Y4=Y)
PS-80VI Y'C.(LF#9N?<%O&+F$/9LJ1OZ_!$GV='J<(-/PB'HZ=/9L0WA@L JQ!6L
P&">*H'TNC5%=&/1)W;*1,/;4@['4P3DQ_H24^6+YF#;"Z8/U:F8C*ISA3!>Y4)+9
P2W-@44/-R\D9&>OED%\<G<LJ)S5<Q.&2[/!DRJ.-2*2M -LY,]Y*HD""Q54JZ=C.
PGJFD4['ZC3$OB)9>\@1C.063_"S!-5@%^B/+VI#J8:\-!P+R''\U<-VB1)#1MD=H
PI37?#0D QAOR]CP@%A,>;5G<#ZGOG[9_P5:9+3!V+/T"]3+\3*5RJLGWU"1&;>G&
P]3$EEV*;O-^UW\)7(?#5T;R?BN4KX-J01?(U+^<;\90'*YC1.YCC* ;TIA=1]85"
PH>%:RGH/1U8VRS5Y8$0FEK7$O#7L#I;]V_"0"Q'>8!!]XP(*+I4*?MB$A *G*X$V
P8CV[CN@>-:;_[" S7*Y U5"OO=/SPHVZ\L)%0U+*U?,9YY&B>]5\HJ=N9Y6.%B0X
PI/\9CE?!-BF^M:=Q[//#<(/YVT11-1<J[@-)C.W)8/FI"8L2<^;RE3)N24JQ*O=/
PP6R6'9:6OJ$_PG,NXDB6>[WNFT.UM$\4#W3F_40#79A2E%,/-+?=-F<C89V7:9V8
P=6<_D#HTR20,K=FI>.DTS[&VCC;;??GVJ,P.74 <$3$U9OGJA!$R&:FD X0\$U/%
P#+"H)J2<%]"H BXE2(H"26^'LVCX4%)2U<6CYPC80SM9JC/7;+6%= &XSFEQ/9/3
P#B%'Q,$:MH=?YIS6C L6FK@C8U3NR+I!$5K,T>U8/;%_>*)DN@ED]6<G7>2^)I 6
P.Z'H:,J*72ZE;/,.4'SC6OD%H891@EP!0\+%D23P=7(\ VGK5_*UD7+'.%^@3O7Y
PBGETK13(_8^:RFU6+OP)$Z$310E?RYCLU1$'T-_A5E!C994<."GS1T?BZ_#-RT@+
P.]841F.T$&XJ!]A6J^1*W)<_F8WVH0.232!Y.!\NX996R> $X5ES1;%UC\:=C)X^
P]#\L+OZP $[(D4X"+)[2BF.3XNUTC_B,5UFP#ZO)C\E. CO1P QGJ'%I& MAWA]4
PZ6!21E2<Z,BA1FY*,6T-)K+)+ZF2UH'4,*W#'*?L+F^S:[.B (V9,L\19$QU)M@*
PJT9#^L:6KUC;?S[#IN"YI3YTAYER@BS\6WP*9M0'Y:E?OV,:',<?;[T09)R&(OPP
P/I"?I$1PW:T\BOI'Z"N"Z#E&2%W J]4CWS9>DK-!7QX>.FN4'0H6^S$_C#A.;E 2
P.LYD;D2NWS/1'\#D28WP\X300"O#O,G1/[[XZ0"[NFKA5)=<WRTF&\W[,;J616DB
PO4;S_=JXM:V0.#76:IR8+2'AHD^Q7L(H-X=I7X;Z0]@O[R$=3?FW)VI;2W:E%VPS
P581(D_]&0>-+<$V[OT0,2W'_#54A-0;=VI?^PIK-7S7=[2WB#O8;=5BR+$*?XHRA
PTQZ@R_I$MNQ^2C\=<B81^4UVHV'/6R/.6>SY#GM/$NF1BM15:"[]GKG!X&._&.R=
P+Q-1Y(75'<]GZ&@-<@#6UA@D9Y20N'J[AU?_^&#C/(C8R1&1_@'&T0>Z(B[?@4K!
PGW<%GC5;]34?4C6XUI[8['D1EH-LJX";+5OED'EMBG2E(19=$BNP\T5NKT\EYF97
P:RF$EV GU' [# F;BI.HO)DRNT/7_]VUYKOAVD*CTM_4 PP\&TX=S'SGDA2JGG@#
P>P2=SP 2N OLI]QO7?)160=^4;PM\'\Q.Y[XZ?%-7//4;&7UX)D KEM'?M&AK[28
PD[$];)2KOS"TDQQ<^Z<=*V?0^L42JE8ZKUN&D$=6(R,8>^_;X2PX&8F20Z'&9O@F
P-J@^RY 7\!+<,F5.KQ28*6P,ETO-*D487!?VVE,LX!-DS7NJH)PID0B^*N>M<LQ 
PVQF+3+86Q5&<^[[2GAXI2858PLYH*T]TS80:6"."LYVT.N9P<:1>HWU&5* !LZ-E
P.Q_CDO.WH$0E.2]'FLP<(NOM?/WR!^AY_?T!<Z&PJ(290*UF;[BC@<)M;H"^Y J]
P>G&90$0!J)D]JODQM_<BL)'%^(9 W^:_0W?R&%TC%\1 ;:R_$H]+:A5I41]X1,-_
P.[>U;J+0VVTU6>#C>(&MN1C7^$8ZF;&CGL=ZDI:Z$&!K58B"6R%Q'TS>>C[2*[I=
PF>,]?3J5)/6A8-]&X]MLN*'K=B,0.C S</A(>[!@+JCK?K],!BA]WBM]>N7*1KF:
P%[T#2EL@Z&[B 2=^5O.$^B*P#LI6O@GYA*.G(5+7R'.<3BW1[PB,-P#-C ^3;RTO
P+R*P6VY8IP8OH%YD*'-ZM@V.RQ&B,S[-%2[;,4G_K5;187]9W DYH&]T->KIC:<6
P]3U.U!;R6LYY*]H(#TFOOZW[^U,<>%=MMVKL .Z2._,'U225(^T3O!J\YASKBQ25
P#0/*#NCD\B@!XWO(>E_*>>5%3O^4".,5'I2G!J"D71S1L%B.-\_'C,S ;P<F>=;_
PGQGWN\%MRV/2.CG_9L-/(QL]3P0GF"D\-ND(Q/@JOEP+ZRC&$64GR!A.Z._:D8[ 
P5=5A_\V@_0 (N%&='@7<U^!C.@-:5N[D0J .M3!.I"(K;F'%B>)GR_[1!,3C]EPX
P3MHE_F!^^AZM16D,_AW9VO:.^K;!-[H#W?-M^];;&M'4O#5F:8WB@VNR!AXLN&EZ
PZXM/K>3NB]0O'>&.%,5)+XFQ%C F5.WZ:\,2'JPQE\J?(213X*568=V*7#;-Q5OQ
P#3I+&Y;KN'SYFMC!F*,0HEK[K:,F48I-2*7.:Z-^8NQQ8Z\[GQSH7$O7PUY5"DWV
PZN\/7QSB55S;P4%'YKJR'.OG['TR(6:]\1%R;!3*DQ.56I)K9M<H[*[+79;LM'F 
P%*344Q=499$-_>+9;T:^P%N3_8K2 P1A(FZ5&V\G!@F#@OG<.7I3D+^)R'?MO$V_
P3A0K896O"X#D(V*9T&0GT66KK5+SC^3*5N/F QSP_!A*6SY@S\O6GT<V[WX3C<*L
P1.V=\),=(GFSU@9M6Y=H=40FH<H5=9]0(+1"O%BEYHZ^4^$G\48^>2&N7[X &?'J
P=W_O]?;I#DEO7R^;?P<96Q"Q)4%^??*F[W^$@+S6VCJBOSC(='2Y(QBN9GQ=\,1&
PRHR/1\*6#L17W\P-BQ\G#+0]3!.K!UYT179Q9];()EH+@M57H2NQWVR/BP^) 7/8
PN$R7Y3GJ70O"7R8K]O%]K:#FXP[-5,&A37>__5*#L_(8TYJI2Y(T\YJN$*[*GUH.
P^G+&</:O]UD8QV*/J&V0L$L)Y>?FI,0)V;KA<"&NS%\2+<XH5!+';H.*6O9&V9E$
P(K;Z>AIIE8);3&]!6B6F&SEG(Z7>/]^5^V2187G0!!=XU36EZ%O'+CVXMWF\ 5H>
P>&<3=MK$W1!K]>9LX_1><HJCH!65XZ(6<UZ>[A7 _WKB3C9U11%@OPME485D>+6A
PX],T%&G @)Y4@PP0=<)\.1%E0"\N%L'H9#[&USA MCW< &K7I C2<6)+Y@69MSZ9
PRFHM/%MXATW\BU,RI0*BK=Q63A83.=:+J22AG\1D$*$(*P_KH41S .HIN3B@\ "-
PUX5YKFIRX#Y -W;8'H0& (;599G,&AB)T$5C$]Z=/,X]Z$\<8!=S\$0!FLN>,452
P$-A-K[1T.32C-?XH1MG\N.B5<O!?Y02V[5NEBZ5O/A<@X"N5@87G+G%L+QL5J63G
PT 4WX-S=5D9L]$91WAQG1%NZC&6XG]6L)]GVG MZ1BZ0@718\&L'I42E^'&Q2<L*
PB$3PJ2*!T$. I@KJP!O&OB#WDRI;+M(V0;D38@X4O"1]1[ESN@3=\:YZ1O*%'!T1
PB5^]],TFH(^=HH=X&S?3[*"U29).>YI_M^XQ[P5TS)6>7MJ#NYJV3_8(/9SF3NY/
P\QE9R[*N;,"H1/B*.#6"RY,SB?J%LT::)F"#SP^IH:'48OO EC;P@;ZXF\L/>N0*
P;0T1JA^5.)LH*O,-!OP>H1,2>>CVS?M2D'<+3SQH+37SC R(/2% P5>>S2OWJF (
P,(?,DR2JEB,N3[174L^%;/))"BM>XQU\?!S;FYCI6CX71[W'5;'ANY7%(<"SRTZN
P+@R/ZWAK @M.C3^SW)P_N[?=0S&\0=U]4M<:,?]MM4\G>0+C;8>C[=R#'M2,^5+O
P?,+<$^9UT3W"*IZ+\JD6;C!]$6T)]+&! T(#UU,7(R+W0HB-QI1"7'N^RBR%G(U*
PN<IW4^5QIXO;IJ&H>,:1)EB"A>"BNA[^=]!YWR.(MAS(D'G#?XZCM%TGGL<[DHXP
P6JYJZ$5F#25^0TIC2RZQ!$-<M\ZS)LS3\W"2 CR- Y3W/9)7$(T&[0>G33JD??/G
P[3-QH*_B5I 981#%PE9^W N#M)Z4Y&/\UO<6*P-T4N[\U-?E#P.9Z8%A-'L,N.?1
PD?VU[+<^1Q*"^J-&ZJ6!6=/"LFWIA\P9/].&^MG\T.I78H R\OV\U'MJZH\2U9XV
PWHLF!VOD.1!OEN14O@=$=V8T_>L6)]6%RLD#+ZB$Q;P8Y''[HK2M4!S$<1A-X_8W
PMJ3>9?]XM90;@G!3<-E#V?I8,@7>30UBS#_J!R&>$NA?V71)RL%-ZCT5_:W80]8]
P5Z(MOU*)L)RDPY84>K#1CV2]QBAB0%0#2!7^BT3&+9<^JMEQNT-FEJP*\PR*.'6B
P8^:>%1#0_:HVG@-G5=7%,.GJIY[*W-G#2,52?+S=U.AY,O^?2U4^L"!8>UZL,_/M
P^X&4-J)$NPY+_/MQXR->10M#JZ +L4:L@FY6W0^3 D=Y"]I<-G60V>Y4Y+PN/"L+
P%&TPA.SE589ED3E@EH]PADF[$\G&>HA]#!F^@AYFM#"!;\L/S4,Q*\RK5([+H^NM
P2I_/H:(B"!V!#JZ[UOHD?N!4&!=T-X)I7Y[#:-&*#D GO"9L,)OS&J-_DF[,72']
PG8?V12D!'H+U$@%LW*-+%R;KVLG[-(Z!<_RH/83T)(44KTZ=P$WF0/^+NA*-VD^U
P_54Y06I[94Q7L=R4,BQF3KV%Y"UW.F#3.X9<>P^X)CX"^*Z^0K5-SQ>Q<FMT(8BI
P+1RN(B&]"[U8IZ<C5-^5L<]=$B"-=3'B<Q!,!HZY+3S#)5=N+R"Y7%]J_[D_U$0C
PB1HP_7=N[,%KNF/3BK$VN@_[GU:?:1") HOU/4@5K!/<',3AN)_P+="LPV/[."9 
P2PKQ]Z'T.!6^(.J>*F->80HH;)TU@2!91@@38E#%"DZ!XZ'"Z%#TIJ=J2^^"VRL$
PUMK=SQ0!0<TXQA9]K!8-$"N^7&.;&&+KC%=\;RK/]$@$.\36@(S'-:!Q$L.!5B4V
P-D):IE3AKP"'RJ*0NHXZ=[G.(ZP% B8%6UZVKE?9*L$/QL=WJU\! [2YI6O\'(@N
P8='6G1;CF@MZ>A&32OBL<PFU(9T7D?.+1";:Z#PKH3"\D4^6B^']<\206( [Q/Q0
PMJZ1-I9EH"D;KC]C!%M.=5/_^DL$;[G5SH\^$Y.5MH=3\ED=UEB[_^-^EG)KQ!\3
PWW2R9_: 0 N!@@^(X>!J:[M\1YH#UJD+A?;*.1JN^L,'+BCB:C$H#\H1\UZ;1NG"
PSQ,UD6Z3&J;EL&-DS'<TGI0-.8FMLN-MN,W)TR7*D;!\-5,"#HH!DR/M7VR>P#_$
P<\L:#.P+T76S-I'?@,0SI]LUZ?==Z%8!+%\!\MC*$!DU;C10MYB=[4:?Z#T$S VJ
P+"N5V:0QH200YM8_OVCE!ZYR[XD=:Z*:>'J/XEHDN$ RL]*'AQ)/2AHDHV83J:?*
P?R!9H-;^!&V#6,V:51+&:L1P'ZY6@1OIATHF_0* %_,!_-JA0?29)9?:'T<4U])M
PF%FC"#.3J6L"5@P(5;0W@=;I@G_>Z@^+FLL"B9J38DC>Q^;4\,N8 WR5=A5C>E@V
PM%G-;EI^#KZ*,:L?C6=T<\(:#NA]O?1/?H<P(K]8$8A9DBHQPGT=/K!#?4.N>F%'
P_Y*V8#3.(BQVT71^44N^R=+$@HX[1?K3H"Q^&%%8T[4])WO/E'$FVF^%K)P'1'2@
P6^L^<P'"E%V9""D-C*[Q5:MV9NHIS(73J;M0P*;.$U\;F3>SY%?E^_$#N[@#Y#DA
P["NPB?5&D+@_3N65GPU+LL:.443EVH=M-H>OY#\>9>NDRX"JRHKMOUC.W %8SE7O
P79(8A]%[&#+E$"C"9E,N;(^RLU=KX4)/V>$YNF?/Y*(8JV[FK'M]'QF56THUX$V%
P6,'H)U+N?R-(X:N[1IR97-'\^' %#<*1^T;_OI?'W[OP:GR^)Q*Q^$74B^[<G@I0
P%S41L6)PZ[)F21B?0\((<EI0<72+S*(*8<_(:%8&(C039YS3_PTV,QAR9:V [6 [
P6>=&-C&?X_H:8E#N>\1U2%[/CI-;_7O0_&U4XYDQQ/NS:+GFZ!+JFL.K4X*UFZ39
PCC0?DFC<>2.%G9[ 5G"IL^'\_YK9O2KSH5%^JQL#O(9L=8I'$@NAWQ7MWONN@>=(
PQHO?Z03V6_8!YR9+,=8!60P#%2J>NL+C?&=$91NPO W,XLTLI']GS)B7PFE<82:7
PS3AO['--16IO#-4YWL./\>0XI553T]R0[JFS 4D ?I]NC/8H'; VY@@O,D -.Z4Z
P\WLH-WIYVU$8P[<-:]S&='7\,,GMQOL@BV)'M4*ZK?8J/*\0@(Z =_"$L0#/#-\ 
P/('OA-?:4+^A,*202P)>6D6"953)I ^=MX'U)T$63Q-$=G=N!V@ROU]A!U"%MG6P
P"NQ:HRA8.AL(_=W L[8U#&JJIKJE>5!#AQQ>]W",S(NGFA_=P$?97LB=E"E^5]%F
PLAI//*/@QD0<+5/T[.,2!QBZC4I@3S3N)D@M5SDZ?APQAKSF_B"Z&)PP3OP^2\(0
P1X1J74<&>WJ3MY"FX+D6-\)L"\:8#-<Y6%'/OE5V,TK-$%%_'>#'AHTKBGSI=\$I
PRWSEX[=TH#=]W!%"SO\$EXE48=58*!Y>+2\MD.+C[_<ZI04S][[<_B9\Z'_@)_V$
P3X+S\!,E6DA$.]6EI5 ;:=,A$U-/+<NV9G ;]X=T&5F;H,%IYF?O%\Z9\E*,FC0F
PQCLXC]"L$>>"'0+?0^I;][VF[U>/,2?9;AY(A#G,:=@#=40^* "8BN-QZ7YW"__<
P$B,\;:J,SQ=_,!N>#[GEVM X))KJ\/<)EFK,16"'0:-.GP0!J,=JKI9'Z-EC+\5B
PP!]PM*&L0BK?$@<VQDC-.L]M&.VXN+BX"?+F'N$6_H)R^.B8563K0"+H[<B_76!"
P- UUS>1E*5)XS81U].46HL$"X](X1?%4U$!?Q#"C_JF'A@]9"ZC T\[WL+]5ZL%B
PW:*)IZWH^;6P2H' )MJ99$!#R-JR.D"Z7JM /Y&U?%_0P>[>)R(5_5BSG;F1JJIR
PP2G@ (=!-HTQE, <S;!F4P?Y#V>+8["!%3MH@_"P,)LG2PAIU#7EF.8:Q@;(_4"E
P.:F#%=.!VC0),#^!;>JHOALB$FU\0\\@BJU"!%[C_:PI&\Y$YQ?TDASZ71%=T,UG
PN*0L![IJ\>5066*KM0?!+ID^U&O#;]I.V61:D>' %&=TX(9JSM2:_Q@NB_7&E97>
P+&=QB"5EP\IXBJFDIN5Z- &D.=-@+/I:#RJCA&E!4X+WC@Z)CA5LH_6YA&@M^">0
PXHI^<N#D?O_A+6ID7B&XQP#D3P$ M '/NG6US4)+(Q,^A&E3#3[F!(4%?A7E(=&%
P+-A:QCB/L%Q(B''7)V)?IOR.TW%+4?()U$6#MKNC^=3_C1]#4)U(.BY*H/"HNZ19
POT_K'!BT5Z6Z#M^=^QB@8BU&=$[*Y2^Q0%4/MV*UG-@*5R6 T!"WWA71K()A/)!-
P?PZRY\KQ'O1UK6^QR0B%C=M6IV;OBY23E(W#<X9\LJ8HY'M2P?_2JI+$S'G+WBFC
P#4.XB)*0_^V68S3= 2MF]'G EB).X2RT9H]U1I^L))VO(-KW#FR3AX[4[)4=>.S.
P>@X# L.*/)KX]ZM-43>84'[9M] -.@XP_"6?<6&<4JX5PBF4K>8JT#S@@ 0%OC:)
PGV]%XTK>"]EJ77H.@3"Q69;_V=IJ=B7B-,$3;<5/O+,IWP+P6F'BO%CWU\]R$,"=
P7 P.%=OMB?<WCC/,5!\ANH8O9Y?Z'_$LL]Z6H71^G(KQP!/FOZG"?;.&"A(1W#CL
PE^,XQUN3"#SHW+Y=\EJ3MN@1-XNS5*\J&I]HZI7Y#7;=WUPB*"]-FJX)$E^\87RX
P9O=-]'KL)']6YU8(9I4.IZYL L3YPZT!I\^_RDTH0]7< 1@!CO:H*MGU8Q?1M"\Q
PBK/#O ._14E]X%FC4F4>NR-E6&^^E-ZR2?S/9]N+VTUQW'8)*;"Q)+=(_[4Z.3XF
P!">+0-M^-;\0;%\S%6QM[-C&0 (,3K!N8!Z^(4(O]+U<C;(U;@L\.M_TY^]Q P L
PB W&ZC%V_"O'U75UH*%C_A*AM"_==_+D(B?S#?+U0ZPHCE=0T0+J(.KI]S)FR 8/
P2BF]7ZF7U\YZDHLSWE&#=YK;H Q=CN%!!M.6=2\/.@H\?K-]0T4K;L7*Y2;[I4X>
P#JCKS6S/<O.*"%V%%> C]5T?GGT*-.];_,W,O@A!T8QU9F@R;:"!%--C08B:7+R2
P,YBT*QCK\WI?#%*@&K7D:ZJ_LM[TW2#PP8+_9Q]F^F1E@M27H(#ZXIRC^H+2$P!E
P.%\S#,:Q(1J<0*",N(PJ8X5S9><[W@E$#WN\=WIH]!A&&88%K6\G1ZUVR\<Z(FGC
P98Q:%+'XK*LA%669'J=_7Y4ZCK2C]*43V5H@G*9?VW]G/2IZY^C"IO#@:O# =_9B
P=3!ZF0.S5.:A])OD"]OC3 TC@9W#"P-[=BP_W5>_(%\QIOO"7VP89(@5YP=DD@3$
PX+-,HONS!E%#&R3GU:MKH6A,+;[&[OB2K+E 1\*DX9VI3;L%[_0^*E0M7;P99?:&
PK)LD-@AWJZ];''Z?EK?+9R,SSOKS\T-[I(B1SAYR__[DN(B2\(J_UFMTQ33TUDQ$
PRV2D%C:NG#? C@4+P2>M/8O GUV2.;6(]%WHATH52)0RET+0Y0O7GKTV8@1&];PI
P(KIT'JG$CQZE<+C^ XY&$?/&()5=L7&;CH5[X#K <Y?M&4'CH5- _6@*<*A5IW+\
P>?'7QBWI'2^DX(MAY;GWLCFJ^I_+7ZD=[9;"!R:[X#/%?BK_-1'=7J\<@4^1'3EO
PYEY-0C(=O!FFSIT"L*R[Y0)+'8Z(JA"37ZSDKWWIR8+T_ %NJVJJ?$HH.RR\[;"N
PDC@"];8.V/E*6>C%#DBA$VLHESL##PD\9EIL3WE.&*>>MR-S78 F5T&'#A*.6%,.
PJ*0>DO--W<HOHT3\$Z8H/K%/ =S%+7= Z%,$742R3U@H%:TM>SP%NSV"*&Z+]6\%
P'',/4X@S!ZDIG-L#BPEX[KS2P DE@^%1BN6(^C&SBP9B+8.D*7$0TNRQJOP /0\W
P$H6M-H$MN?F2C3$_24\M(-Y'G1.B(?4K:>(5-<_$-)F#7[7YR)??,ZDI8$<K]./9
PTPD0Q'Z*;>4/=M%&'S,QV&FVQSR;7T(-HV::)V"T Q1%-J5'G!VE<F]9V5L(:Q),
P1T"=B8+L";Y&D(V<[V?;?2G]Q;(GYG] C2O-"EH=^GQIJDV^F'*I;&XNM#+<ETP%
P2(IY'R4/WU]H1'Y<IAK529\$R3\18(J$B,S,8NWM_ <3A4DAPN^Q5EGRY^'Q8+Y<
P"<S+U%BI6^P:7'6"+#7V7??U+O6K) +"PTE#C;-*VIYG .T@6*B6)MS^$E)'+72]
P0>94(0@AT0<HKTU'FR7=)<[,])=0R. @Q[Z_SYI6F'@Q'S=FMVZMO-<-)Z7OG0G_
PS%8=^<3]]0C&=8V:V2O.BR(8[NRMH 5OS:KCPP%V>D@?9B!Z,2LAL[2J0W])'4?)
P3F8%W&>#_W6V[<RV#.F)@+Q1D@-[Q5;;UG6**;*_%DC!$V-@!B,D(@A"LIY/W65[
PGM)(! *W64%XV8Z1?ZF#YPIR?PXWZ9HFSL6HH)ZQ":GNDU.'9)6XKC ZR<94[D^3
PP%S]]+X?J:,L^$>4J7-[< BO78[L1'"E="'C"T]"DP=0S6(>ZNB?/XH,!V'^>RXC
P#?_5#2:/5BA@E"SR7$W33UVKZD 6B"0,";(X;7[ONK5K)]R2*<!<'PK6ZQ2335PM
PY68 DUI&NY6G[^(QRLG@<O?92YR=9A1&G^>U0_=<L@#+A.^<T"Q7ST\R@&7J8:W(
P],;(@C55\6#XMNLUD84,&89U;K(2/H>KRS,L#=)3,+]\C283LNF?!7HA%D9&7VOZ
P@)U>Q"7D*8!!^_9@'VX01NC!L%^IM_]E':GRXW//.?VN4SF,VY/XQOB@O7G^:B$U
P-S^Y8D48=ZG_?,TA7'5G(ET2[O\<6O21BMV2[3@[@&<A\>B12+X=+K-!;]J0#T!5
PIRAEW6/B^XSCT$&A<H%:FZ:1GM#8TBH%0'7U:OVQV/,$ +%1"[^1_:281O*E,"8W
P C!XX0RW\N'<[J\0*5/'/I@#F,<LD)I8O:(*%Y!>O@3++)#PY"/DZSA&K-"WG6HE
P B5VZS0LQ+7"-V>OA5@\$P.%(4*FSH/ 7EY\<Y]D,E3N:JN#SQ.S$M2]*">I%"?L
P*RA[)NH\/SKJ8_A0EVI/-7V2NHDD8,@*R3Y%N*4;X\SP'E*0G!@)8-,)&AV=8+RO
P!J[X+U1!XRF3Y57^PG5Q:#'%G'+/-E),TPJ,DJJ1+.FS- ;4A)_@&MWI_QCI1%^V
P[>+\W"+RDIR>PETTN3FH'K:"\G@+I?38!\<PM)K/ZJ T/WP1OQ)D4K53X3CA76.5
P@,S--^UM[9I8N#5NJ]V&$'LF>-+VVH*#M+ZM$%IRJ^Q;^4Q@E#>>N<J;@RZ='&7#
P;#7"DHNVJ-.IBO *)GJ^#9,__%*IAEZLF>(C$1'UN[<H0 PJ>I*VT=&GVS[/W60U
P6W6L?J SL1J[LBE!I6M)Z!@*YE]_"-9&*H76, *E@T#A_).F-:&=R*=EI 7V5@E6
P7]H77BKURMJ8/GF6(C\G)N7F%Z:Q#II')AW]Q0<6+@ /P^/G/QC&BF4Q(O/C413'
PP\+DZF8$B^C.=%ETM.E^,5FZ&9UF-9/Y-M_O'X&),7']FKTG#4Q$\D;?59'_)T#M
PU_424_K*-8 '47B#\%J0T2<B7$=&P7M7IU\.P+93.U6?I:SA4MVZO27F[D843'NT
PRYRUG@TS\6=PB:;MG^QH?03TULA7JT2DZVDAUBK)=S)QW4&WTTVYGSWL]HOSGK/8
PP6N:P6=>0"=R:V0;F'S"_?8P,@('9RUDGWT4;\W6-"O#\1J2ZOWQJ 4-41[9Z76!
P?38K!)-SGD2^3:7^S?_DQ(>-WK8&>;#YF2P63'W@KD5J-/PLO0J-8SG)VP3(Y82J
PW$CP]=1)7NB_E#J6Q'GY-2'EH9E\)&,PG*^=BC(T,M*KG@M72&55]!\=OR#&&Y>7
PRH(YE<YB9,][/H\[(\PM5=#^-<8HQP4/@.TB_%DG0156-#CFF3%9Y/RZ;3H]V!Q+
P8LXDJ6[1#(VP :L.=Q:I%2S&OC.Q3-XKP/%.^OUY%?[FR4LN-X6Z>A ;6%(F,@MC
P-2( MS]J^D)(J_>;0I>R!^ZPXA\\;5%W$U>F!]C-)*,/MR'!Y05%)GVA5!Y$6RO)
P[6"&3*T7/^C,#M&URYY?3GHZWZ@"HL3P;ACQ9!GS4]-Y8QT+3V2TMI@32M"@AW,Y
P%F*#6#IRL"8)9^F8KA23/EI>7?-Q^'5R\J^"+]Y^:@M7$9_6F@77FX+P+S,!7*#Y
P'FR/[J$?!UMPJPKPK;EI*97K8LHM:?;BK_3#RD2+-)78>D;5".X+*:4#JO8<_XB>
PV/R1!\HS@"'[KF3VS+MB>#*N7!D#P$$@[7T'?,74D=^AB.KMG=72F@6S46#68H<O
P*X$B^2-.2@46M("<A"Z\\0PH5X 581KWG^!^W\%7_JZ".]E" 6OZ7EGO]/35B,0H
PD>J#3^D93QGV:F7YL:@Z$,R(V01^E:E[)L;#IM/]+".'SNU*O,PCK'0 4022>(/W
P#+*\-YK(1_(IRLIVK./2.S8D:9(4V#LTNSI*"XI6]?@)6ETLT%&6?@Z*AX6J2H/8
P/F5;JZ7%'U<D*S>HG12Z>\[;]ASEY'J(F6L1:H@G"FFWA;[=0)HRO2H"81'?-YYJ
P!<4V55*^ BSR]WVOJ2JQTE/3<:"N']+7*^._D"A)9TPM<CV>YWYXN][[-%).<]BX
PA_8!O(!AY;,O:?:Z_F8JR %LTK1,#!I(X@;EIF6S0)L$>]#?B;Y_2>3;:G9+?WOK
PVE=VP<1(\[RI+BQEKZI O(%WKGT])WY*"'(2F.=VAKP*06:J.*"!Q<V:SDLDP<OP
PS2@"\*5="[8H2H%P*C,J:AYJ8)$_LFX^N!+049&S0L*T21F'N-8CUI$0Z<RL)-S8
PCS/1H@&])8!'L2(%0MVMB@"8"/3CO[B^25.:XDTDT HS\(*:+PC\8='-9 "A10FX
P?0X'5T[C'2?6CSQ.:D&/#O[P0Y#4?S'(3GH)^]<1[(RLM.5(O;B  %@<9R55AIUC
PU>HQ$X#T(-]'0,B&Y0X?(8H[EIG<;8VJCRT4CJ"XXT\8]UWE^N&[UU.C&T+H\)@L
P85,=WB$D*K@_P1S(RW;P%C8A2M?56K;YV.!3NVM5DT%IS/9$6W\JIE#F*'XX-M_0
P? 1Q]_HRET/SG(*<KYO'M^AC)YT&2XR*0QI U$<F:W6QTVFN47'*^^SOO99QJ;HV
P6#%BW"-V+9.YU0BG -9%2,871X?@_?6N*IX,>.+V@CC9:"IOZTA1?;));I-3[P,H
P2Y;LO[(U\_C0LP9</#VR"!S0 \_[-4W+UK=Z<6@L-_2#F .,&[Y03U#9)R=(*/ZC
P;+*SR:?X!(=3?C]+$<?:$:RY85^[7,_X.I%L%6EPKNFLJ6@]_77>AL?N:S/NU1FF
P&7I YU'5I$\3S/<;38W>N%MR9WHYQEO=GZ6!XAS@E '+SV(E&#XB?')D!V@H=?S#
PQ^UC(%8/T,*H<CGKD&#)%DU-VRR&SPW[M2A[['K\[!%1!4$G @=J +TK:H#2_06;
PMM(0Y=AG7*2E#8$E[LV&A 2O0,U>$3QJ/U)'&W_' P!"? Z<$L"RA(/?S:&<I9**
P;L%54_=!N/E?A#[>X^^PUQ,1'U4:MCKW!U?![K9K@_QH(C)-)V9;Y_P'><%A)+N!
POD1T4TD]M'NNZOF09<"(%90;% \RZY24,90ML)OPB.<BPN162RHM-C6-!FM$(L>[
PD7XZ#-]$=9:MJ4(H\K<7KZ[) /KLP+*T",OI3P8O<SS82C+N@S<J@]*O\_WIRQJ&
P\GPL)4\@)O!59RP()H@PKB*. 5-TV.I<MI$8/XOW?#ID ?+G]YS:1VF!5&4V1P'@
P!ZSZ6(>;&ICV?YO*NM6,0$1!5;-=0[NJ;#,QIQ7ZPP;@N*D!Q9! EV;NP(:B0.&^
P33X+1IX%"/B5,$[NY/:\6OR>!OU%C)ZJD(TE^?VV_5UQY1@,=F!I6:>WUV3 +1D]
P+SE[KB-21?E8[)\>A'+, A7CB/8=%Y >T>AZ=(@NYGUN&4+4(C3GM7<X_?L &'XA
P'%[6+I]%OZE2>IG+NC.6Q]#Q OYIMY$B ")67YQ07N>-QXS"YOT:PT]ZJ8=B;%^(
P2_0;Q)1]+1?)@YC$X.VH8?XRZ 892Y96.'!%R8!5F:MWVXZ]<X,:??V=QB[)(3OR
P^\*^J!!YW'GY;:^9(?D3PJS]?I4^=Q?3%;1/8"R.FV$=,#AFHJ^CF]O<[SQ5AMZ&
PZ;;DD.C&5X["XYA[#NXX/@A1^IW7[D5GDRI)8"J>'X=Q#!#H?:\!DXW=ZPA5Q=[K
P)YFI\L90WQ4G8(X8-.3#1X5N^9F8RJ1A1WL:A]!M6^(Z+C[XX4Z<ISIVC:,W#DX%
P=MT^BY@B --8PJ+%+7PJ"S\WTY<+@T["L_@JY9&]LO!5GOY^GK"B[M/+"S=SOH;Z
P5A7B>7:DZPZ 3R@U^2IZBVU(3#6VB:)C7T4F)0,^U_B@G#R\2LZ@Y(Q:_2)=W@;?
P26%$S8IMGG2E\TY=Q*+PF''<<_7)7)M!FD/=05?[I5NPL]]6N.8?2##'W@7=(\S.
P9[*/X%_4_V%S#HO&AP!YA\>K?WRM*RFC?*0X.%I(^\^=9QO]KS5G8/(L7EOAL@\B
PAG5'"*5?SSF1O#,51L6E@##V;R!W%^(99&[2/_&[:HYR#S&P&.?-7H5%==U'?!)X
P ^;X&Q#0JV78N*4[1^>QTQ>_<)D']B:<S >82$?N4RI,,8$"'6,@?ZHLZ3#UX6FB
P:4>P=B$,Y[_[NW>>J2=(=5F92N:FL8RHW697?I )U@5L\$(4XU9;9@ZBNJU-#0]Y
PV-9*A:_BKE10I_CJSW"9-$O-,4Z;!S0EY$C>7%0MM[U8_ET'6B=P@R1^+PC6J[> 
P5*V"=%C5!R!--C7=23 KG'4KA/D5QO62V:^[Q.CPN9U"?-F,."YWVO55V7L >8;A
P;J<_<)C5;5+X*-#<::!D53A]763B#0P";5>SVJ1UHC2 M"%_[F2M<970[M]S,4]?
P(6QFNG,F,'$*PVQ".GT@!]+G9TXH8VX_31C^=QV+*<_F6CX_9_&D DGG+I\_7SV%
P1 (/7J<R9PS,3'!BQ9H#9\VJ])H[4OK:>(-A%V+]Q&GFD*M(,H"G&GC3"R*('Y[&
P(8U N_SQJ:4:VC4QX]A4%M4Z)9G7D[%=+DFH>=+S#ZR/UE1"*)WB6+F>AACS><:_
P887]/"405%<QX[9]NKMNI&$B/?XFV:)IL%282_E(QWR$*< V_G=]-\F?6XV$<MR@
P%U].EK$WC[3N:B<EXGQ;2+$I?F'L1(>$(4]?TLTI*=T:^=O$E("PGT)N22?Y@DJ:
PSV/*8#%< U80B>523A,/L^=#Q"8\1]&*<L"8^<8*G%C"_H<MC[. J"=?@P/!%K]1
P;9&3.<XNS,]T$GH<T8@9)U80T_S8OKWX_L0$?!\S:4%_7/9 N33<)W-W-=I<7Z+!
P>-;#<]!WT-R[K0C\&O?!B=]:Y_J-&%$5:%JMWJK<,6KZ7A'SY!4$R[SIX"JP;<!,
PZ87!RW_L(SND.Q<0"UMO\ H]:!78^-V%3NE9F&.%JB:@OD/AY&C/VRT :UK*D'AH
P:%4$2.A;8D,O64"?X,(5?:=E %AKUR6'^9JK</P@&AISA6C]IMW"@<A@75GQD@^/
P&Y9ATELND3:TH:&::T!\&@6NZAOU2O)QIL90"Z#1I8-4 +245.U+@[- VK?C8@JZ
P D@4D%^V_ )59$34(#3)!_-LEZ=FF'0Y14HF%CK"4*/K)D?S_1YX+N0]ZK'Q4ADS
PPC,6/QT@/B,ZL&7$IQ_0QTOWB*0_X'& B$M@5"8U6'153QPY\6.M8X0:S*%MO#V7
P*ZNSQW(#'%%*&\$L&ZXWE(B*C\-?=<]&:31(S3%2/2;E2-FG0PCPA5U4PO?]8[L7
PTA;" >%EIH?&T1Z=I+PO7@EM/0M,HSAP<UH016=W=> ,8;L1=F8AR3+2*=AO:4P>
PE#UW97L[AEH.W.U,+UX1YA^8B\OW+Q4>@"&;<%":IJR-CM<6BV2QT\3)A+UQ]+>]
P5N:OMN#P;7&C[,T>(TQ:!>VG^!NRB" 49]"F:+S:75I6$PP-<4EX)(_8.KQC=95I
PE]$1A?>5Q N2G9@*6' _UY3P<)Z>VF=I$+32GIUME8D*5^$%3@*^6!(<H?94X4$6
P-3P?V$;?=+B_:SF%_'?U"J>@\B>LR^3@8&0_J*?VD&R/+/2?09_,T?0 AR)2IS7Z
PS-(N,FMNGPK@B]A590:<L%2*LNY:B+U='_J\G%"U)E;BP%LGQ,Y@[1HOJ'?[>/"G
PK/>"(IY<2,"I*K$H:E&&0#WV24HCB91R*:^5/_+7*>ET@358ZQ\V];;]7CQ4&\%;
P3W+6ER*'](RD\P_6(*%B]OQ_F@(,@9914-W<%E0 V*+&:Z6U7'\Y7T29TO&0\&@L
P(81\^S_<L$K"73-8!8=49'NE<P%-_&9WL\D[H'=,,V4X5;V,U0Y6>ZWB ?+3UORD
P^3HD3K> 2![B!GX58U+C.YHX<X%A1PIE=4>U6K4-GJ0Z;EI=<I2X*)7+A(;UGWBS
P3NV+M9JS(;'!VF&V=?GK$WY)(%?;] GAC=&$W/-C8BMGMS>W$0VTB'P/_.OC,F#:
P;$X2>O2HLS%M .W@)LYW'M0CT*/='27-9I[+)[T_!J9R6W;%%KO0? >D.Q/>:+;V
P]/ Z\5C^!,;;4=3=U0-+"6\HPF]+G*_5TU-?V%!V9P/NG44ED07O4>!0!XLKJ&P.
PV31[BW%]M:*(Z.C3B\=B"\_X^=2^GZ&7T$Q)[ZV:_\_JV'F4>@M?-NCR>=RJD7WS
P+1/^^^#B9'&++'NDQV=2XWL13^@!;=7#85<I2; -.D%6PT-GHS4]Q9_[KY/JYT.P
P+#FF$JV:%HV_.W0 IR3E_?:O__YBH#Y94_!2"DO;LAS<]D>6(Z0]@V\!Y6/*(ZBK
PF/=E0VA*:B)W"ZR$F':1\7KYSA"R@@+*PFFYT!WA5(I;X'N3R[.18?O(EL.9MS6A
P@H_FYGO;W&(E\IX6Y8%]_+?)84F-W<>]C1U,NG X U%HA8D6HGR=T?)\>ZCRA"C9
PE)?8S&'V.ZU^JQMW0+A=O+@@7<AW\4N@:G^UROVDE\6=5T 1)VG4S\!RAL?DIUN*
P*2093!19\216XX>64116XF^>)B(@TLM=VV61\DQ;OJIC Y. JWG9G5A+B?'!T.G2
PL(3!]QSXBWS$D8[$D*%^<(TB07YJV)BK9CMI# ZY[\S'I.X:-6 JE3"2G/GJ[!&A
P\M1*]4R8AD$[.JW>CM/\6EXY)\])Q*Q6'UT+52BZJD+]_@XV=A*=5=-6; .G5L)S
PTF9<$\ YHT1,4)1C(;LTOKF#KJ*1U/,P?U+_B7$=@29Y\V+/M.79</<"OH0[\*9;
P9DY](QK\(EQ_'#W>S#I/)JUY&D,J:06AD^ZQ#?WAC=-&'UPVJRC XFM5-+=]NJC.
P=$WV).P\@DSL/6\R#TFKJ"?_TXZK\[J6U\K8M3N!;L-).S2Q*^H(,T^Z]1M @VGV
P]&_400ZR,D5G9:J>AX31HAM/6Q$4E(:X H/?.$T*]>"VH).";^Y(VH\'3[U@(.F%
PQ0WW(@<W4IUL7[+F8X-U@ !."TSD5QD$\>JYBKY7N;A%W?<I^FCK=FQ*=!7YALAM
P39:].6M)5FCZ*,NL/?&!>=N+K#E:R-L:9IV"Y7[^;!UH83J[:60A#[WZ50@CR,F>
P#-773EG+GY-7O( EH5-NORH/ ,8BI%_7$MP%OL%-)LGQ(0.:'+#47&5<![  %12^
PB+S:?6QK7,PPOM'LR><3"\_:&8$HT6+!/$%Y=]_GV3.4ZU!02W?)QZ+Y(Z$:.F\ 
P.:%!SHCM<'9//5QQ^%JS?TTN J5B5P<,&B(EIR:^$+TT[*(B^ORT(SB9U>CKD#DU
PR4<@2UQ?^#CX=!<'(,!BO9$LJ.E>$Y)3BI!H?,D<A-5B)($<B'4_)2FV#?<3,8Z2
P1L:HCH*-7=/D!O%MP0TF<8[A6^NFQA2ZD$0C*LJ]#8V7;1N(74 $2P8E@9H%0 9(
PM(:+1=@+;!NU:7[]1IIH+Z"NW;C";/)S2JQ3"7!:[1]>RS8 ^_#+W;;-6G/E,J^^
PR97$C'6 XQHF%HM.6SF5J99H:T]+V6]T"AZ,,2P2\%CV,_QX4+'<0'/_G[[= SX!
PGC_;6"Q>+@"1\%<0[GQ)-:)C=R".(Q3ES:F"IL#G&(: P:N_J=K@)=*C#S=2)6#R
PM O^'J#3FA*H'$] *%L9T;E*>-)L.ROTJI:TGR6ZM,G[JNY/Z3G@1-J9Y_[9N6+.
P;;P]MDEAE%*[ SH!U^2 ?_:<J3X,342?8DK@E2J8<N];!+%?SP";#DJ5$:]Z&U$:
P'0!WA7;A#&[1KX "V]')Y!JY]B$W@*X ]AC+'9DI;(M;O1V$(H'S9Q4:IY@(@WS)
P0JCH\9(GMTBLBNL@&>L'K;^YBKO$4%M?NJ=XXE7QA3Y#9;DU#U93T-1B\8O>@1)'
P7+I75Q;$#P':,2S[Q64L#HP]Q7&4;S9,*#M8%37K)EHUQ'=&T'T=B$W1<J%34R]Z
PPZ43,$%<5H(]TT6;;F]E/[=;IE+.@++W'C_GG)]DP]^\XM1DTD*9U?#@A;3D3 KA
PM'MOP*04)MHDDZ^>;)%(6V-:X1GH,7/D)^]]W:\Q"@1BV**%<6[F4P2XT?<&\D2K
P,,ED%0MD3.VG5C^WS (F3GYRA^+G/DP# K<P1%QBU%&6R9?T7=B_"11US4\'(R&/
P_)5*_[)ZAOSA;6@7 CR>6_T/A""^O0KMK[1I)O]\4L^E=5O[T2']OC^P]-L45 #.
PC^4G0^Z<H^BS_>YN8*6DQ@-$=,1RD@IZ1PE=5VBIS?1(R':WL,3[4FM2TO)#0&E_
P>A#=R8IZ!9*+7!VEEX6EEZ9-?E)6_&YNZ+O.)[_/%)X/M?VZ"@K:F+9C"13NE3GB
P6C,Z28*(/[:W)-I'?S])&%IDR=M7]]@V4,T1:@#RMDO$%JCR,8Z^+G(YRR0OZ>W 
PFU/C@.HN)'I;9A7NEFE2#E9>X$!KND4HQ.X^ H>1YO<-T>XNE_5PA9W&+G_^.YSC
PWEI;PBL6\"*,$V<1:MM"8 _2NUB"/ W^G'C(D?%"@2.\3)WH'EQ4%X7SW.!O4.3H
PZ)MA96Z=:?!4PVI4O<Q>*[&DB(GIY%SZFJPR4]O'EM@FX3-'**YKV3.R&/D\\2^"
P<LMV]DK-=&,]1,Y2:?P<A^,OM J!IY<@9L: :9>2*"YEKR-CCR8X,N1*V%"4:^ @
PD0)GCSK2_'='2B T\(:CCD&L0I)*?1>N>M_CJWEMCZ_12S0O WA1%3Y'VM2_/_BG
PM%A! R7#(=L7E*0._2YH<+!(!$1\-7JDX<;@^_A4!L.T"-'_Q$G-,GP[_LOX'B?$
PQ$X&6;HM4.<&K:%HG'!>/AUO&>MB-3(<;-D[^#PK,KUQ0E%7W7YL.5>%[Z"V+H;K
P@8B%J5MELP.[=$_LP<G_TCZGE2*-'!6C^]71JY;*Y3L3##+0"2CH%5&P**=7:W:J
P9>>N=$606%,\;XE\JV9H\:^+ 8#WZ<W,E76[N/TSB-"M:P-<;\MJHX&6*@V!? AG
P4SU*Z5_-N9OO/4$!4:4,JE8*1+L-M(Q!K,\RAP08P+HTI#<\RMIBX^:Q$)BN&&6D
PI1"MR@88U[0L012+-BZL]  ^>N#6P"^24H_'BQ;]99J9&_8F(:F!,";O!R.VK*!V
P]?/CX]U)!^VHK!@/39YP*."BSQ+FJ-L< YUBF9N/L@K#5UKD&QA,:&?WM,$7%M/?
P]714RN1:_TMDT>Z^^F=&%$;PV\A-NT\7M)_7M6\0@>6B^^H8%Y%<.?=-+B-OC>R/
P,C@NV[")3'E.<J\CZ7!#$C#K,C/@HL#I1Z"ZXK/"_%[W11>(^)J:DDH61DQ60K;\
P "PB!W125D\IN503[P#4L=?X2H0%=]*C]8-6=3C1Q,@:L&1 CF_G0S[5"\(L;/#E
PM/44FHBDS-!5<;-'H@M8K$ *E@3,]&()A2V$P'34T@JH&K%AIS*X1)D 6X-0:\S%
PE7(!O%\)Q4WWROGUEDRIL;1$>\A1SROI#'OZTY%0 @OP%]5UY3W-!4>RDPOJ,U '
P;0=*CFK@\)2-%<9808]?FS__>9XCRX<;:.SY&Z&\R7+$_6*ITL@)K!CX4'MI4;]L
P?F,^P]=+C;MOHFR32L!J%+6*L-4Q+_D>& EOA(1W<^H%3A<EJ'@ N='0 SU#8RXS
P0'=JC=#@^U50"4:]C<C&0B5;!F\Q2S_4"3^R08/9UT#<HT]N3ZSMM#12" M/_2;E
P51QERG<QKXK2IDY%EK&MH9/\B2QY==S!KC",:9'S8,;F@ >T,SWF#QJ@(Y]A6\-*
P;D*UO\!S)L+72E"2T3(VF'!V8E':\R?NIV"%++RKUE)9;BV,@:0"1='_S?L2J<B&
PBMDWT4][+UGD<^)6H55'#B%,U57FT,%B+FHI2!GV-%$8WU8;&7L%6%R@/Y<(0QZB
P])SE1RY8Y#ZVQJWA^:!_2WZ1)TI(JD*%J?2_3=61S)P-$I'9"TIC8".A70]76D::
P^<O7MLAPS<( 08G0!Z_I=W2M?,Z^9(LY^][ME?7((H(% ]7;WF$*V#$V?9"@#(CE
P86GD";=;<2 +IWY"^OMD]_![:@*06YU8XG/X2&NJ(\!"Q1WV(5?VV#F>TD;>!H N
PAUZ:)I&SNNFDL+O$PRKBFPH\KQ=#@-@1:_(T#WP4+YX!U,OK-] 1"^M_K>L\JS:>
PAN.^3#9-!PP%/78SB9Z%6/?2'G'?PV)3'(4MG*X?U-N_MG,%2KY5L+AF%ZK3GA8U
P?,.&<>NME^:="@/"K_Y?(^>XXF/*,QLJ(73-]UQ  #Q;.Z(G/W E>,<E*7$@ I)S
P%O_L0.G<NIB3J5I)JZZ@:[5F8BGO4QX?%!V%[T=SW,;:4">UY>.?>8AJK,AQO933
PAA,-?NJCA2H:EM@(_E!OHFH.AJ'X8O1-5O7)1](?/BPEMIQI_U"+6\\>2*6*/J-V
PB=]4/%BO#CD723U93?A"(*177%U!)#%C3&S4INLM FC,0\_X^+U[=IG*@%AXU&%U
P%U,\D.P(Y+;3[V9R@:EBB2J,8KVU3G<*]OSFB8+F R?5"HMLSUTF?M1B?[UL"!L>
P:H.RFVHC"FA"6RS(>M+(1*^VZ@7Q=_.;T545\^\ ^U+9B5+/ (]IRB@:.FJ1\6,3
P*/0(,4,KX>%QC[4:4V9C8%14K)TB .6_X8J&T4#%XIM5/1Y5OD>BMX7&\:VA5):F
PZ03"$/"6?M\:CO\QI1$#7%T-$]L:*W<"Q4.BN*>9;O0TXH@E52H#NQQHF+/</1,4
P#<?WU.V6PS-6KN8]T0S.:2@XYURQ4=B*9!+,PW*F[SHIT-+-Y(E&EI5[H)/./RM'
P-#.A[?8(:**R8: T:0F^.B MLOY@:@MYW+@PT3MU\M^Q6]'D[,VX[GLKT[NV+HL?
PP=_W;>V$B=)9OK+_.,N+>,X6B\?E]ESX+=\-8ISO^[W.MS:FZ)U#8[-DC8>A+<;%
P4/1-KW$_0!LP>H^>BE*U(A412B:;HQ63QVJGVOV3S2(H^Y<-,[LYOWL %)--Z3EP
PC\=7GGD@#<':69Q?7+*0K-BMGCPP%K6?BAP(AW'#)IVA=-"9GY#8MW,SB#J6V=8$
PDQB7%U8?&([%X6]#UEC%T\Z]MZGEOZ:'<V >"'N]^LJ+6T2Q/.U7U4+N2MB&]Y9X
PGZJOF)TO"WP7=P\>)X#Z=>5JC ^84QS!61 UN-I)]'ZA.('/?*FP+[9',0'?[?$Q
P5N+D(-3ON'-"Z#LDMM%^8L13\,ID_^,5A9R$%S+)^-)SRQS3J S2: /'?"$2O&65
P5,?XDNQL05<=%G-I)1$:CHV);VT6JH%H,UV5]-C\P5Q>H;I=W5YRS2S^=K%ZMOH?
P"]OYE'VY(?'@8;#:.B0I23FB#G;"X2DMT9PQ>F&<Q7H:SBWI- Y$P13/45P"EL*6
P^%#4<7@+%<6OK>3O0ZDWZ=W0C:$)"0"?[^G,BR3AAWR3)H,27<K@D[A!NE+Q8@*F
PVT!EAMBMV31T#[=*;XB*=,M&D=ET7[%M;G8<]3F561N]&7PE:*T^UNY99.?8#S>&
PS_U,DR>)+%2%Y/M>SJ 5_]H9FGG=B2'&P\@"+Y\PX1B[0)H2>P:*4A9TQ=Y-Y9OO
P.XEB>II%TAX*.&U2^OOL@N4LU?TN_3C<AS/"(^A; )H-C>5I=3I5TE?&'P!^23\%
P$K,I>8'7^!#,YS7U!Y9$!= CY- ,'=V4FH^+V"\G]0Z%<K_6\1&,]#G#KDF$0D%#
PJ):+?&S7=<\:.=]EW'^W PJ2!@O3:A=+P$ \2(W&QOEG(%;^3*,2ZHH\HF+S\&\[
P0>\\3#?2)>1_HM;:JUO-+MD3!EY*LB"(" G[2<)]WVC_*FL^3,0>1,=-=GG9J0?;
PUYMV<HQI:5*< 9YN^V$Z.4(G 1%J+TOR+(2Q@!JO2Y.\U3ZWPG3:Z1<MW\I#GG<2
PGZ0!'(AGK^A@Z33_\GNT/[(W!,VW%M;.[$I)7P%T$:8O%M&Y3=XJ[;IU37:95LZF
P1[@YUDBZ;]R"=9F7:/NT0J^Z44@O%EFC\, /YMO+Y;8)(F3!MM9=(>X>VQM6J7P>
PD4U4=V@EW%D^#UJ*N?;YE'I2S!N7^F77Z?TI#Z9L7.:X]1T1UB+>&8-A8$L<0&BA
PJ:DO/6Y&+5PYRR=EKG2I+J,^T1=)L'&A.U>@5"7G!IY;][W00I]$/>M#+<A<E]O=
PM3#8W$2,$OK5K7LTIEP[=$L,ROQ][/S>@N+]:ZT)PM&=6PA-K2B[T@&]1T<XB;FP
P4=-/B@)RXX(^]WZS;X3<HG%T#."<&#0L4 AW;9BO5=)DM%#9UF=X,'<[C&+X(>(!
PC<@VG:C-FBY#97+VVR:TE^;#23SZXQQP27&>=+)O/YLS%&E!=Q3)J69J6PN:MD9+
P19.V"'J.N%X9"PFWLWR&\[,BG^.ZA-3CG\I+J(P))#^B_7DSZ=)?L,\UME[N8X.E
PEAD4_[%?,009T/;%V=22Y.HA DL4U+=$-R=$K/3UC; 9O]ADWR[WK1FFD9M= T.%
P#TG\R)X>4Z$-OE_J6L3Q/:6$4D[9%6KX+-E.B2XF(PA8Y3"V +]9Q+S:WJF9 7=\
P=[Z4RB&W!_O[DQQ>R+C ODCK1\A*LQ9$")PA&/+MF)YWBIQLK.<_YNX8006V%KPR
P%8BI,4X+MKLBQ\F!NPU(P2F8Q+VU\0EE^MN,X56YI[Q4F40YE<\D%SC07Y40D]RO
P19;U%YGR"&H^<=CVH\[9A$07@[R?D!=['V% (=(@1I#>6W3TXKAC97F1L7>U\86>
P.,&;P20$S^GA9884NOY4M>O?_^@IV2I="0:N0G["@&31=6;#HW<%$>MUTUS8^Q+R
PD/^OT07RS=08/F5'K$ 5M,A-Z:R9Y9DC/^8Z/#!> AU?X(?X^Y_C8<G"@ $,!I'3
PXG,F\.^6@CB0'(F[3NK:+F&G5( [V:]Y[H%/)"(GR8]5JVAT=5=.H3Z(WGK(+L#$
PW6*PAW#""I,PY!J_2:L*ZT#ZM,))AMK<7%,T2UZ7@T(4VGZ\R!EO3'1B4$4*,&A>
PCJ<"ME,LC 2V3,5S?RD>^QL90I;H96-^#:^6VJKO[_O?FRPU.%*.H<4F$6.2EIY:
P>?@,GW"H_X1"RV9K\YYF8*L[8,'NHLJ/QJ2@V/R(F&O#X=; T\P;B#,-AL1TCJ$.
P4P%>",R"#A0%?)ZFJP/^SR&46A],F;R'=N=[8C7GKPV4!(,..;"SV'/I_/YJ.O7K
P51Z[-#T!%B3-0S/0&^*$:SHX8Z_L]75F>:<08C6\T_P+90J2<E>9'W6UY=, (0S-
P[.]4M5TF;(5!M6R@QR<<T7PI;Q07GL8=&*;@F.>7%X+>E/L21USI/[K(US$ZB1!4
P"J^>:X<$#]E:\6W&/J'$Z9@[HC;9>3(BPT_ IT>[X_ZE)<+NY@HQ0 F$Q5OI6+/9
P#]T]1?5,8?Q_^1=;+XF>\CW<0>DCK%\B!9L<:F(E+ RG;?*K4T_<T,&6ZH>8&0EB
PX"EK/CH!G[/%5^Y@ZJERQ#:T=27.P?IK,%WG1PO@^U*9C[/8.F]!3.%BO#\5P00G
P QF7/[T]9FN/O"";OG2'X3&]U!ROM^0\!U'&WHSIBQQFY0+.018@4"O8/(E[Z"7-
PW&6YQ^T!$%7ORI5]'0\QLM)R>0<X;RMU@NL4W!V0V*]  28JL+J[T&(6ETJ&):=>
P;(JXW(J@_XDY7/0N<B-WLQ"9R032:>@_G.36XG73:0;<PR#']DK 07-D'0"HE!R?
P8A4>D$ITKD4D,O><=ZD8PBHE>=HY13CY*B9.PY(^]HM@*G"TBR&D*;JR!GA>0;*^
PLT<O;-)559I?F]H+U%,>)PD5N]1-W,7B7V-7E4ZNANF^4J;<TER30;!AR^1J&M0N
P9"C^%>DSZ;5W>C&B-B.?4%CJ15#@Y@)L/>@5/]3*[SUOJ "A6;RYW=N+F%9*QY\7
P 8Y%*F#GC+H__8&S9?QDN^BQB"L++\I%P+IX6"FRI6I!QRZGCFHM.J#(!YA(9,..
P+]G/@EIG(:XH:F@_0R<NL^<:M<OXOG\Q8I&, :V$0==8WNC]V?1EZA$PHT(<)['6
PX-=D,-X2Y_^U_?_NV->?AYM6V<*Z]YPD/P!\,?$]LBQ5-R=ILS_7WRMT6((0VW@2
PJ PSTV6'_J##\"G^[NWU09$^^(D*U>2+O)HA0SE' 3\($>XQOBS :X3Y^G;H$@=U
POLO(+\2WSD1+%\_%#,0Z4<EAF;!"4K&#W712[O(S0EZ:B0U(2@3Z042!VDO?_ML^
P0*@;YZ5('QC9G1V31R7PDBOWM.SJ_7)WO69D)((7#&7P%.](VJ;=[O5@RL%KWE=$
P[XY(%$??$+M)J:WESUK$YBRC$V'!=5^0([F.-(2@#W(TIO=-9#ACW#134&U;LPT&
PF9C)A#Y5FK\F='BD<+/!D1.95)RENK,8;1&%6GZ>Z%Z^G+U(AHL"0]A2J/ 0P2#6
P'WOXU8J)0.F6 ^MJ* ?_H#A*C1=IU9%E,<SM2SQE"4KG:,"=J:#\\H\JG'J_Q?7-
P36!F?%X\8L$G]U-_'D"<8PE#->E?FC"T*/H[=^;M::/"JL*+;J*VC-<V14GU;06$
P?_6T:"GX>].K,O,CD?F*O]44- L'6"'7,:,M5%35!K@[&R%S4E'P7GE0[4L+LLO+
PVRK0?49=:P8W]V_H3>8T5$-4DSAZ=^KUH8/E+*U9]91EOE]?>T?]66[LE$5;]C->
P\QX#,^-3R/'PE+_D%E R1C!&).18CM-#KSQ@8B/2Q\R[$K[>UQJ;NSP-C2G/]^T(
PEIX(6P/=5D>(+_&#R6V:AAG4\<0Y$A-O]* )Z4D1LOZ_-JA\;7^"+N@O,;':]%W/
P+,J1LL4:I\^R !1C&J[U-EH2$W$SX+L@396+/ERC5YB]%.' V5-320I/SFGK%,@P
PH4SSUVA@GS3D>=(]N!->QRSG)KU"RU1N^?[:%-9!*X'\3^7U[U>V0CVDL6=([B+:
PQ9'XTT'A0S/DC3C%BI6D-NJ"S)-W'\LJ0!)'3JK COFRG2&FHQH51O^OYASUL7+S
P%;].9L!RR$\O\7H]0=K$^=:FD"!U."!:Y*A/X8$%G"X$C7X30L99&BUS(X\>GA*X
PT9X]:J9GYJ1SNV31!7\2*QQSNNRW +,T<QOW- [M"<<N]77CP/ZD\%<5OR6^PFJ3
P%<S&)=OC'KE<3AFK=#(1 0* ]AK6O^WGRNN54!Q)%R'0#ZFM *R++T^V9H]HF6NQ
P@!IP'_[YF5-]QE>CB24#VH]K1OE,"W%F2?1D'E!8:+A[:<U>>*QWQ0MAW5'#='W(
PQ"_N9KV#?Y[S0L@GD"(*%^H/[5XL_<!DGO$V9^W+L)V=M;!Z$VDJDO8D_AC7L-6:
P]8J])/U@+3SS/8TA,Q&1LH(W8V8H?EK 1/!$E(4%(&%"#/2CQ-O86H#B5 VKG1W*
PTRK)A-465N-[MK*7]I?H/J!TQ](_+@N4ZQVN!=BLCAD!5;U.".R) 7J[;44648WB
P/.@?_)>QE@0,V6]4BX6 XF.DLK%C,N(_EX2$(8H^[KHN",+>A#W.&OZ^XA5U=5A&
PL;(>///N"0=DW;$7.+\K\'?V<BO+24H265#6]2QPO[9/]_M-65I<< 2MK:HDH6K]
P.@/@[W=.B&Z5T*:(:?$8NU"GBRAG,);45*C)O_WBXX@B\%7:$V,$]D%=:<D+IP('
P24)LH/Q*3NEG@AB6 TOJ!U4_8D#G1Q&O!!/_$RW#.NHPI5 [TXR2RT'NQ62??2GT
PPJVWJZ9])A<5VV)$R9L-'L2,JCVZY4NQJQ64<5'A/Y5]UJE^8AG=DH^ K:/$KPY8
P81,"C5V[!G4-6-DW=\3!<4O+V<^$N$AH&^UK_*X7@M1IHX9\45:\-,8TDA&!)^)?
PNMWCX(^_/,=S8.[ZZS%>-4:0=$+O?KYE5ZB6%R:<I/N2Z#!9+]D7IX.%M>225.!Z
PQY!#+K?!?VI4 \!B615]&I=MF0;P_@27^X?BV\J]B9[(IZM_W.K6U[6).H>M&<\G
P)%)#S']0,3@/*\2Y9Z(UY>:96QN=Q_5$PJS%#K,[UHI@AO7H*BK?'2%%G<*F0_%1
P97IM*[Z[)5X(S06)S J.'UX18#^8[H3+'K7S^-E@&M)TN^)V@<=#S,O@ ;DL.$/P
P]QG=:RF/O5'2A?>2>/H7<M'@'WTEL/SB$ IZ[CDR2GA5MLQAR0EJGIW7N 0Q4,'3
PG1\F2>5]-%@$.X=!^^4+([N&!E:6'#W%\@2M6"X/&D$:L+2?U;_I?')"-V2[W653
P]_D#;E],7$4C1Y!GFDB:LS3SN4AC-N\$Y5]O["SO._',.__H>.9K?8D(3!;M-O@*
P$9^M#;RZ*&I-@!VF:Q+(:K"C8XN7;@EX:@:Z,J8555(YLFE 4Z()/I(U%<I"TC!O
P*0D(V]PUY,'N[RRTBL>A,2'(FSD>WM02I$NSNM]IL0D!<ZK'?S(,H)FQNAE'$;;K
PT)[:/-X5D?POC3Z4!4SJ@SE!5NE<H+D: (GUR7B^#:6>1$72&0K<( 9O)C'-43V2
P%'U*'46K1R$9)=SNZYE<,Z]V89DUI$ZG,S6A=S2=O5B*@K8,'8>HW+;^+]<$>:ZO
PBJZ%4:^GZBF4;CB.SQLL1ZDAN?5#=)DR8%J5*^WG"M!@5P2#/&WBL,\3A%9O6([%
P6,CADJE5%IB6Q"(/3$5*FI&KK'(7>0:_M$_ "?ZI2%HHE5OR"E:;E\0CI'(1J7_O
P2E%L-:)$ V05@G,UH\T-^]J<_@0/6)8'PJF"5;LA-$+5/1VN*2[F(R]0)M,I#K\/
PGD8HH<?8!X[2$D_[(42XHB\&BO=O1-]@IKW<(2EL=,-1_]R5TR34EE[D?KE@%!O\
P9T_&]Y9/*'OZA^FB TXK!PS_AX5_2I<KT\3@P:\?A'RT>!GUDS^S?WO.MC9KSB"1
POF%%:/ZQJ*]R/E!S+Y"1E&PC+E'D7TX&S+U^T9W#?W9=5:SGCJEZ,!#X"-T)]6[&
P]>)1 6,24#\\_F('''QOJ?G"@2.+15TA#WI+HCIJPM0..!;X==GV"',[K_O_D]$$
P!%O$B// <'P\\U@";SH[ DFRN-003'3;K=(A5PE>FVNV]&2.F]=Y9<HPWE @& F-
PCR-?BR&N#Q/H^5*@V&9*X;W.$&92.49;DF_L!-@-EX_<H;B]W;0DW1HEHD.ATTS%
P F%17&MFE%*PF\M> 2G*!2GWAWU4.\L9G8P;V3M)"\'+S^CJ3>S.7OB<WI\3=9\ 
P,,:H:T5-S /J ?3Q[WGL429T6-V8(#2J#2%:BZ$YBH/J)F\S32?E^__\+<%GIBM$
P5M%% G_ 'YFD,PHW7><>85J(<L?B5HA_7IR<)(@GF/,+;I!I2Q-"VF;I/U\"IKK/
POWPZJ\OU"%SH\26<M\"Q]DXB5Z[D(/'1&@%Y?)&T%CF62V*I?9(8QA?O3/NPQ<5!
P:M\9W8-][G=VO&5+O</LW"Z<*X,_=,)%<#H '[<*Q6H [9QP:V!R;6L(#W001FJ1
P-P*W7[@M#A&Z"N(H?K_%1US>#3*MO+N5PKI0(^!83[-SYL$/],8N"C!(5]>L'+>D
PP:<:"C,UFP(4F;0T[,?A-- .\<CO^QV'@1.WF+7.^TA;O5/;C)<\?+=U[>4X]<_S
P+.?=Q1YO1E^G*8W,(@<R>*@P;NK=_R^+P6/<V3J0+E:*5.G+85AYEEG-FQE2W@_*
PBEU+/^*V" _FYN&^0FQ(OLN.Z8(!_^)M91.[2,]N711^6MI;_I=<VC&5<7U4/4IL
P4/(DG,=#KA]]TU;[SE12^;0JJ:$9-B6[6.2K,2'A,<'76=Z!-F8^KA]$C& TZ(K!
P:W7K?C,.BX?,@MMS#T[C<)?\.KNZTXNSW:(/M=]$,BI%>@R+-F-S46.6><A>C A.
PO,P$:K<?>[ZQGJCN E?('X,2!"@!20;XU'[]/0&Q+0]M>,BTO_#/KUO<_!0QF#+5
P#!%J [\2M",[6*06L-B!-@O:O1-1I>X"$PO2T1QN!'<QW5XM2#91Z&8LD.5+3-91
PB[5I FO6'1M?=U@:XNZ8S/DG]A_%7=9J.((E-B8_<17T_"[0Y@O&N3=7%"UC2 ^J
P!"U94T1/6$$;NXM?-X]96B*YC)N;TJ998SG$?1A.Z'Q(F"%?TDQ6^7<\-$=[0O2[
PK#\440/0]9 #;(LOQKQOC'UU>!7D1[/L?LA&PH/8\&I8 P&0=RXR(N&@]O'+N)H5
P9ZWP,>27BKF\=%WGC2XYD KE*A2C;0RE6N119!12=*;"! GP3OAI),K :[Q)##\Z
P5ES#,J5Z+J%Q&$#'*=PK-^,U)BT;@XT9RX_.RP)QW.!KW?]-2V!%EU=<Y34&S:L-
P@4O>A98#E;1VH0_R;K1PX$GNM[U;E+(FNA(GU]=:&8[],XR.YUY'3D17K8?-OXVD
PVRG0TK6H_I-R 7W@IX9_M D13D?XYV&LWJVI\D$%#_Y!N5\0RVO2\AO\%R;!GRO3
P&TV3F'D^@^6BI1Q_=#SXTGV1,=C]"VJ]=&S20<1?2L"J +B'(W#,XA$]Z=_,":\,
P4SZ#3O+&X3N3-WBKQE\_77("*F'W&40CB:B<Z!-,?U%SV^2A..[8S(=SKDW?XOJ9
PUM"9.C3P4:P=KI0N$]7DYB4R&)8Y3]^\AB"=N@P!Z.S$%2I&G<"'&(CYN$U)F5#\
P\J#65J&ER9W^)^A6=E,4P!1L20;VF2AKPC9\JYGL4&WX0-/_QJKD[E5-92UCLBNP
P2D "015"#L?A(OLO))<Q_]\V$?MIO(W,:/ZJ($(D2#0@<<T5.+(A8%+23EB6]R:4
P\5UMD^1^OIHNKDZ:7:8M&[I,*IP[NE4?;O-F9TXF!2J4MYG ?E%ZJ09@Z:OW<Y%3
P^2L=+&7 1'O>5:($7KJN+K;]5K@$<E%Q#YG,:#-"V]B5(41'C9!S#L\J1HBA!IR1
POWD'/WC6GPNRK@!L*$50C7;B=*$IAE9_*=-QQ3W_)JQSO,C^?/+\VEBK>@SSM.C=
P85!G#?HD#:=__>LD*0.:VM6\4%A-OU,-<Q2?_Z_^_Z8DF46= #&(J.9N\X<,_X?6
PI^ 7VPCKOY+LI9<)GLAW"OA\F.P<@]?"O7M_)C/N'=LWD<%E?B9EG\8C>5GJ1K&F
P\)I0I&S_^'I?CC%P /'.'$,AZN\&'&V+V]!NY'#LO8TO=(F$+Q 7UU^;ISP0HSQ)
P&0^^2Y2W4EB08X]J04'2[]=U-\/^V<IJO8H.<@@Q%\*5WHT;H;ILZDR7DB?YF?%D
PPR4T4YG%AX]R11MB99^LW9S=EAVY_6F%C%ZF$9%96E!4/\;1/=P9,-..^H ]="\G
P"VC)P[R73LPC[2)39*$4O<S9#0<^<&<#JR8960^IV- $E09EI@N3YH$ <S#N$7(&
PXBT"*+V&.J'EYAI!W0!$@,MT43$5J9\X4U51_AB'3W_N:I1L>DS6$HIN$)8]!8:Y
PUHK09]#'.Y-'XJ_5$V@&2@DBB8-G5;ID)X"K'_(Z0_^<_1I&S"3![5PYG-HY'D%8
P +'K@#@#2G<_3(A<O.SR\I48/.'W&_78U04_Y-(?@+1UFEO?!/I$Y$;S\T%6SKS$
PN*8KK.Z<I39228)SI'L*^H1 ;K34C)3-"[ZL5TYPL!"0M4+H48Q#_75=S];F#LK5
P"-ZYS4\#3/KW9BDDBL/-C(&H+4V]EFE2=UV]#\M/&"+</<]%)AU'-#,N%A=F%+YV
P;W(W"!R:/L10:GXFJA^E!6#5$G/V><[9TH)'<C>9X'=2/-59T2SOA_%XV!\V@/N+
PAN41E[&@]M4->B'4:90%I('K&<:TJ(B"L5J[>AJ$M')>Q,X$)A&0I@$X[[$4B'E;
PY?FM[2M6HF?^H(/Y<1=.U.H]^ZO0Q[;%HH3 !S\X,W#T;JK9ZS:[BWGI7;#NC5X*
P#[[]1&]*::[[6[HJ^4MU9(]4V&!! "*4T/\"GRBH-AL=!TT^8/<F(:DT5?VTQ.S:
PV9*YFNKKRVE\"+$Y=+9!D3W(8=,B$Q8>S"+XA[66,:MZYII ]5_^R4A?[4V:MJT'
P4:4J/@1BN+3<521W.JAP K#HW.*M[:-Y3:V>VQ*GEZZ\_J$7JIN@-K%%W'ZU5F=0
PA(3VGBX+Z/0^D1!F NZ;1_O>4]N,O \CNI_>0#H-8("&\VR"T8^7:VE !XFTD!ZB
P=FAWF4=R('U'4)J'ZV3NH8L5)9OO[]K4LA-"3' :H9C\V ?M\8/[;WT(S-YZ^L,*
PXM:)NS!\ZJG?;;>D08PI% 6J$!]QA:D0HV,RAABD")@Z1'"]NN4@F:H!W5:>16%U
PRICYZ"DAA2>. 9>L(X>NJ]L>Y7V9[<N^_3ZM&9O>WTA 1!)W+]7YC8;;# J%_,4Z
PH0U@S'8 I):B&] "4&\5 <]C+".R]L3VG2)(3)IK>]]L%V)D_GB>S%QJ#3=&!5'P
PLS'/%=IYGLI-*1-1+M44"FN5<Q#8<F0HC/W(9TFARL&MP?\<J+RLM26V#HL&2QH6
P,QJ@=:':($5H9G36$'J.<K:X53+F.'#/\S4RA@Q \>=]Y JD6UP7G/GI[#MY9B^P
P([[\"DI*43),5).4V#!GF2SD/%PQ&]D@4K,5P=->N4[,@22,)%*84%>KRS[KD]=-
PZQ#1ZRAY2B$3DJP\),5"S3EV_$<7-.ZG;)@,^N"Q[,T4@W\PTR*$60W]&K:AO@FR
PW<O,FE9GQE'7)GJF4I_[>X2>@S3'PI/#E]0E0!K#K8OZRRHOZCM+$1L/QG$N5Z8J
P&]2@)Z*#.UVHRQJ"U2HCAXVW2N2 XYNA'&@/./M:YQ:O;HYGZ*T6^\-1 3_DTA=@
P-I8/ORQ&Z0$U,5MU,^ ,7EXWZT!56YU$R%?WLQRQ<G%XA^2H+KYK8JH/3#(6)L/P
P 47);&-@MC=->+>\H[ 8"-1/-+3*%QM5_CA,/7/('LF(D>2P*<ZO.=0#&.9@V+B(
P-&(OW8D2$6U)"+/X3*FGVS 7\Y,R\.;Z, DO')/?"A(!)KNN."9-# F'9 <^<?HN
P2$;PBC[,C?Y;Y 5MO/N+8PF,'6S#(-UYI8Y'__P7[(9?J$[ZCLEWM$M/WZ"ID@;L
PK')+0@^7M"B"^C6H-U'E1I_HM I+D@\]?3'4P2R#-4ED9 ;&^3+>K%68X0B(R?)>
PN$5$#XZ9P7^_BMZ]3$YWD8Q2,8D,I8;?5LU?^MT_)ZH^<ZUT"OXB#Y Q#.P#9+&/
PQ+]9CHT]W\7.7!_]04<2O!"&9D\T$K>1:]WA=<JV<P%\S+60:PZKNU_86T')Y/YR
P' );W+=>DQL5X<D.,PT<-N*HIBO^MW!9>0N- C3,<=,R;6D"[V*_U#Y20SNT/(W'
PO48%%&W#Z$R0%HTKS=-Y>+9*#H4(#:TWL-\E6T %V;+S$?\P5]=<[\.#WYIM091Y
P!J= G\1[0%;)O(HF)8I*J5J*K;S=M!M_XWE-V^\ ZXSX8>'Q15PEX1\4Y,49<-U/
P2*]SI# Y<0L/901Q.<(\I!^Z!7^"OF 1@@/D]%-RV7OXS ,;O\[F>V."E#2&JXDC
P=?^=M,1U]JG'8T)@;^ \U3,W;YP7]'DX?H:+>E(8E0 @=]:0EF>F'EN\PWM9QZ=(
P4$AU%?VLX.!^WSXLO&07'XDD*?0",TFA*G^TO2P$U!O2NG;*+O[>77%V_IGA9*N%
P"O:NY8]!V[$&R@M=Z81%]6U @CF:V!N?8'FYUSTDLE2T<C.R8REDXB!M+I;&1O=!
P+!H])_(U$@CFP%4D6BG5MP"B^-K*4/7Y087_O _!L03ME-?"]UR3MDL[P1XAZ&@Q
P2<'BZ1FR;&A?I>LZ2<0@KUB!YSH=#%L?Z%Y\I($?^1I9R;[,T:O'W("TLM]EW\1$
PD7H6<A#\U6&-RP#MTW#2S> %/UR=:W!FH:\(/\'I]9;1)J.>_LT[:F<LV)V&MQPG
P!QQ0[]C(JO_/LI3KCAI5*;2(F\9\<XHA%]S]@%QK@75.U@#MB+(V7K-I6JBX^D'/
P.]ND.0DL_/YY"" 8,2&_AD&.(U>$1R_=+H='QHN2VJL1V_X)50#.3UNCI47NXHVN
P)"'#HPM%R/W@GDG<R#23QG$#JW@R;>I0YB_!1+B0F-G4LU"23HT9B%K7?QK<B<:H
P:3$#&6>YXT4UZ%\9%76<=9911@<C@_KX <SNT Q@$F5-1%>S)MU\\" GF$QIKHSB
P 74Q]^RBI;V3 W\6J^-$8BIWBVURF..$<S%8ZZISX4H_+ZQR0T+W!@!B^R45;E--
PLK#!F\ZC6O#W(U.FMND&(3&$NDA?1K?#(F!<1,5]C[HR-M^D5\R4X,@"6J'2&"CR
P_60O?Z' P=O459Y&--4P=E"<((,?J"9^D CA>KOT>7_FX8H;[C,[PW*[T<?;OS?:
P3?=1\V?GZ"UJ!D=W^[4LM^Y*+!G>[?9KF%:])<%;D.&^,$GE^E?-TSI,CDLWMU0X
PRQS*[VZ@\WP4' 6A'( *,BAV0U/Q%GCG$(\4:S-?*Y$__G[@7I$HI  ^5VPL/F3=
PW_GD>X5LH0':,3>8DG>3F0Y+DU+W@S@++0WK#HLA;=[O@T:BL-"^1(8!X'*<._CP
PSQ8I:4GH[\O!%C<M-;Z$1X^!;)8L'H&A-3<(F/XP_-3DV6^RK(.ZJW+*:@S%OZ,>
P']6;T-&0[]#1$,3$J.XN__?MOP'+WA7!V0@O-%@..DAC^@A6^6,3OJ3U);B'BGR"
P!1S6/RMZ6)=,(,/U-T06]V(UR55Z4K^R58.-$UE0F&FH>BGP#?0<V*N@KCR8)$J0
P#<#3CBW9D.U(!C6DP:ZLH0V+5%FZ^?(WDLV\$D[>Z1D*,[$)_W@U[DVOJ)LO2%B]
PZ:MX]B&I23[M%][5)H3"^M(.$D<T0B+6'9%SZ'R+4INB70"1,Z+IF&%<:^+R8AID
P3C1.)R191!>=OH:&:FYJEI?Z#(0&G#YU""F[K,$VCZ%-8LA%8.)P$)J-C/',/U.R
P61<#NLE9,"T&'\ OQ/;PW"C#J"JIU9GU/P/C%8\6L^U@)2* NG.P%]*IZJ,X\DH_
PD=S->BUC\E7/84N/<OC^Y(+I*%UD,6'+8U9%8"/VDB/$&+Y807)QER\C**E@T_L6
PS7G0_2Z&L!'\#@IR/5ORW;PEFGQB+#QUQU.O<CE442/N"CW[>^8U43],[9CLC>1A
PL]Y8)IR0.H?1)9$=:12D$2Q[(!9 K68ZF0:1M.FM=4G$$S']MTF5:LNBT)$0A,U 
P<[!1/KS"K"H4W/+S^3PK3NSW1F$5F0T=X+99@_W=%\\E;&I68X)+@==#J?'/>(5B
PT[UD0F^D!3Q J4- 7^,M<88XN$M*>CNUM\"= 8UF-%I 0,/A:T+G]AM%FY-]X^8+
P9N3Q.L.[#!9I54#Z;^XR%2L*E>!8[U'0;EORL//-%VM,+!.Q%JQ=M?J\ -N8S&1U
P5[X>R8V?"=HKUVJI"6*'<-T9%]<J_E)]4D;XC8.NCN%V87JI+VJAB@6F.2R(L&EQ
P%I_P12F]M>&W1^9G V"\DYX*WA:_;-U@%0IN0Z#)8ZZ@(_2=[<SG:7D&(!QVUF'&
P!9ZQFRK_/TM7\ V127<!E=,SFGS599>'>+#C'N0#?F_5@<JM"V&^^_I0_TY70C;-
PC9HI5^X:D*>]]ZC^."(TVMFT 58(Q-O$8H<6H9G1#'>@VJ+H!EC7)K.Y,WFJP3Q5
P0Z)UW(OL,^C-3 Q73I$-HX;=0A&/W/(^ID)RAT5/P9:K'&N6;>BNFP&,).G&@*0+
P=B;/Q# 4,IC<0N@#32T;#8/Y(5D9Z_YU_:=THXSF[;UC+0?JO:_@8J-%#MZ=(I>C
PAI802]MM)R9S1SL\'3-IMCF$A7T+$<#Z\Z, 3A6A.-_2NZ(]U#G#Y#B.&2;*ECP_
P_#P0+G%>_I<3*^5+PL?,NLN!8RMH]B9@O231.%DM0KD'WTLTU']/LS:CL16PX9H7
P)48=@PI3850O<T9>6SEP+1P*2W0([697NBXCOE &LA*B[6;[>$[M!24/H5H4&0V9
P]3<'^JWWGT4/E=$R@P9B-JR#V1M@!]V4$,;KFTY"UF%6GJ*UG=UUDOY9Q#TUVX5M
P^FHBH(FLGTZXVU[?(;CT9I#BFC_H)B3IZ\9A#,O-0IC^)I4&9]L.O3S"IW]"HVCC
P+7.06Z<LC*X.F?SERX#DSB])0'6I3CV8[ED'V6_Q@;,EL330C"[B177.BD".U*NJ
P[8KII,5D6N=CF1W,P YS ]>6!1!^]7 6S:YV =;XI._!*'M5XI)C>X[WS!FD!5  
P41"+AIS!7'_YS?<BZ#7M4@J/*0RL/GZ;BH!:<^PE"#= B"1IK.K_6-&6+X+P).%R
P%-OIJEN]'(Q' E:<3.,K(VL][1RKTYGBE2J/%IQV@WJ*KT?KD_ADPOO62/\=\XU'
P::$K>_L3IE! KE]/?-+_+W_KD"G%'TPYRK)LFJAE-Z'.@C%LS+U#'>J<"-9O*YOE
P7.\,::J2>Q=1*:8!J$0^3 .Z3;*1Q"("VI3FAO"EY<A[5A\E+[%Q@9)VD3C4,RC2
PJH\:Q#"],;<%B501IF$0AAS80[)G]910.8..7+?@>IF-LV(ZV,0&6==+G-3]GU[]
PZ(]GDUQ.T%%FXOIY#OQUH5)$!AW%8M=>1^L:8VF2[COAL3$*GUP4*JNLZI_C$G"W
P.W0'\EJ9NN2/R2"L5]E?*)4@*2?B17$[&A8VZ*",4^^(@1'7 7XQA(YI/6]8Y3>C
P$12Q)YU K9Y(MMG*#EL;07&*,G1?-B-.FK;MF$QDL8FULI\.MP1NXM9Q^](<$A8!
PL8XSLQB18'?WSN$LA-+7SD.5N+&F$C8XXEAL98A*:;(QG],+Q6OWAZ+"$H\;6E/>
P<T+N$# 9_5*Y(*USR6%2-\-RKPPL2\R!8?\^Q<;A^!3-P8,=-H-XI'X89ULT'Y_R
PX1]^OE+#\:>BRG>I>8$O)\,K@0)/)3LR)0,OD1]B'D$.16RP?0L=E>"(ACO-XICZ
PSM RDH77&&V?CA?K$U/%PVQ>1M!;F=#Q["QHTEZO8_;Y)]=T 4X#:7;+C[;UPBU6
P9X#^*1 Y8AA+L7S PG5_5OVB=LV9;%X=F[13=DYW$ZU-XPVVD"ZPT@0NNG<^I&!6
PV 6:0JQ1J.*A-(Y[C5*\$2$6;FYD0LIK/*4L&-CL&ER4B3(AHQ]^S,R,*3K]B:0=
P"[5Y8>1]XDL=NP$;1&>,+!%D6_+!V'2[#G$/9?)9A8.G@Q9VAZ9B<1M<]Y:\VE@E
PF6\";49AM$HY@VO:=^][F;;_D91?;;/%D@DT 'M0OXE)2S./(*]9K_MS4O<>GXC/
PNK+BACE@_^LV".D?>_3=&J0/6^7?Q&P9$7_"!JVSC'=@Z @?U2Z?:>2M P:"'Y!C
PPVVO  REOVBZ9<Y)$5J\P>*($65S$R3+"KX0N4_/&-DF/N+[P1L:22#1G:.5^10<
PPA&$0J62I_#'P9Y04#TAT+*8 V7KI1<+(_5?"^9H+M6J$>^&\X/@JB'-^6<W7VOV
PBDWL48'%J9/)."%Q41&H2(^5F ,VX/;9=03'-JT*EF?Y5K+0&E\TXQ:64H0L4SG:
P&@KY]\RF@0\_M DA"9'#RM6=[EP'Y5D^K_\"@<%NM&=Q$&Z8]XNO#LL,0 Q$LQO-
PG]:<KM/KY>0AMD%@Z5;.7FX$T/72T(!7D!W)1WASO+Q^-Y:I0WY["?X3'KFQ(ER,
P[WE0 J;2J?4+ELJ3FW6'1=HN%6)9DE(\Z_+?_,/?:;ZG-<7X3PR4 X 1)H*LZH-^
PB+HY$&.S"F--8[(%U4=@S&9["\+]?[S\Q+=BMEZR4UZ?MMU\Y-M8N79O@:BV,*/$
PIC%9X==*:J;344/AQY4(XO(\#^-&/W33ET>JL -YPMG^UWR1"6&A"3QDS#1T_/$!
PS%!IL3],Y^/F^\<B&66< #3(5R?S8J<$ /[3Y88=OPBO8[RI-\/V)]TQQ3)2L",9
PY,Z?N&L2M<,C@'7$7E+,4>Z<>V<80^PCO5B"[T<0? H6:MA"](_<:H'5$S?[>U*3
P?"O'J-:5DX\YF^)>D<"I/X@V$)69M.W,.!<+<%-S?M*Q<EV08&G]BLC=#)J*V$XB
PUPEU7AQ;*RT&=.6B.*I+4CP=1[G0$ 7,F;QVM3H<["Z'Z/&4,0 WIG[+G:+$\,'H
P_02L:<Z7+_L+PHTR;BQ<\N$"O4(GUB;(Z(9WER^)N7'&SPCF0-X>E33_J,T5W&3.
P\MH#T1.).L)\N<MH$*,LJ]$$2V5-! P?FL(1,,?6]]*[T/TGT)>X"K(& >##>>1_
P(FT>HS,5?KTQ;/5(>EZ30R0,-:@\$Z2KH'Z]H:YW H:7O2N-S1.,6.XNS6\G;]@J
PS'!0 ?0#5+8$J?E95OJ)F#?A'XV*1HH>>Q1L!3\#,Z U^ZS V'@.^5@12_1D"CUQ
P-MX% T5'_(@>.*SSOK0P70!+92923\YK<&+&!V>3T!SR31!+/K3GK)DQ,@1[61?[
PZJ_QHL1X10Y](3UC]=%*ODO@>^V%O>QQ'EIX246 ;!*:YWF- +29=8D@T.E(S[SL
PEKCG!Y*\L6P406'U%UL],GON1 7?M%G,$/- 4'4[B77P #LH/HW$3&N<<YVW 06@
P<8@Q$#,@Y%2I\+,]UH_Y[HD1QGR[:8H',>3^Z#='R!8:]Y:S!*SEPS(>!E$TM$3=
P!/O3UC6WT.QG6M@_:1"L7.T .3[:M7$CUE0J3NBQK.=?;HD(\3M-9DL+%W?D\K'6
PV0,:35WZ'T KHM(9CX&'(F(8._1DEM"<9J$ X\WV$FY;^KCI7H5V#*-SL"NXH%M_
P'L.(1)S5X(WP@'[-9>LY[0<NA/XFI)&LB*=YF]U%F(+:CCU!HL+C=PU>1]*#[+_#
P*Z'UPNOGK@/K7" >AMT8=\CL!/(VZ\^G5<]],DUE,EB)B</,ZB*B>A1,1+!X7-\Y
PHFEVX]&X D EW4C0#[IC.TJ<CU,+J5 \1%\XQT>N"H(>/7A278/BX<P?>4+L.Z@+
P^+G+?R2\]W:(L@48*/-6US3H;,6G+%1.DFA=LB=I"69M9$R$%?4N 0V55FC<3.LW
P6_ZL3>K^VDLO<D4QO<!XAEP_]BND+?\T9Q'JG1[71Y36%?,G3'#[R-34UQVJ%$2E
P!@0C,JE5R\_19K',0;QFJE7K HA%IX8R#$ !BT%M..\W7]SUV@7V8;WOW*\TBG [
PI#V,A1/?I/01A<-PB^, 8%IO+VBOJY?B#Z8JR/X6MGI%Z>4*\3M@KY(,(0W'#-29
PHB(O#SB(NO\##Y:GK7QGBH7 @_M4",[,65M)(K^])AW#LS%(FI>KB 5%?Y.; U L
P1NVGH.B0K"[4G3*A&\]R(\U3-1;C#>N.$,"2!:WC+GMB/@603B;@;:O\^!6:@<PF
P(>56<V'9N9>=6+$V)]/5=?G$;ZW=*$%FLB$8($C"^]71UTZ'O&!4";N<)Q+V.D>8
P:W5U(CD>"A3.&$[LHOXZ4.*(JWYB0(2'>0R=V1YE>O@!WSD+^5N*Q5^NZ8JI(HE_
P;J5S4\J6. A;FNQ^IB0 9!(G]-O8Z;314'W[D04BQCDAEYLFJ5.0@+Q4TZ5;5RA5
PIA$U?3_S4^WY>1[:/M3$50FT+ON1((VL>:ZRJA%YK7@PYA:3T(M,EUKYDZ(06^B9
P4W*=Q9:L&2HH5\9UCQU#5OZ#Y!6ZIF^][FS80@[@/(32H4D):Y3G,CBIA,>M G0U
P"BKNENG]32]J"E\_G!43Q[HS]VZ8\LPX@O'")+I[AL&A7,5D/EP]MM-[)2B2X, F
P&Y;4)Z3RD,7-T$+PM?T FD<6,0]+UO95/-Q LHZ[.J+%-LU)#Y81M-S;2?""CC\S
P'P"2YF-9,D'ML_.FQ#_\C8KM?TUZ IS! 6C)9.M#*BQPYH0IPJ0%S=VZT+!TZF9.
P<X/#O>XNZ46R%^%5Q"A]S<S6PAFM0Q6]:_MY\>[R- $$.R_M5X2GBV&:73%GH" O
P%2[8RO/)=..?K)> &Z+0VDBF$I/[&^7/^4-X9? ZQ>P#?>6@I5 <G.WSF5'>:72#
PG!&PCAM5]3YL.=^%E0&"P+6:%V==YQ]'<>H !.@/XAUH>M0-N$(*;[$P]_='GS9X
PLG'!!Y@NS@3GE2_)T[' @]?;DN]L!91A (> F,S)R9*6/&/NG?[9B(5H]>2!329+
P]1XE+NH,8731VI;,/C'GK<,PG-!LFSIP]GO7,/N%/I)PLJ.E>X_FBYI80?=HC8%X
PZ4I2!!V"-)A<=276TTG':(_@HPG:2:5$9&+TL6, I,N+:05">&$/"X<;,191+:5#
PG6J W?G;?>BM;=VMBWX0R@8(_+8EZY WJ27:8D(]"T^[2X2VY5_M*G3141%[JC.\
PG\NWVUY]T%Y87TE.TD3%W02R[V/7]3RY)YHIJ/RI;.#0/%\C+@G E(/T>KFQC+*!
PY)D0Q:?XM0=S14[M3+]QL-,@@IJ-J/V6=^'KCX7VYPGD.S:+&&_/ENL&*,4 <D\ 
P7 LO&J+S[DJ::3NG+FE,G]?TCM(M1<+UXH;68S^ID_)Q[.!DVR:CT7/%[</DW?1X
P]6D1XW-2*4H#['TQ@T +K_2-]R[^>D:R+SQH3C+C%HYKM=NJ\LAZM7J1[S(3W.6:
P\^,.GP_E*-L7YI;LXG/==?" E[M'^_T##P+P#7J48L??7D;/OXG0XS".6X*.MH7A
P2XA-(K2NP"YG,KU1G[-!JW&Z)%J@ML6F3AND *I^+K]JN8%DB_-_\042(O=ZRH.T
PE@_S9$!<T7>-'?RFFPE)^'ILX&*WG!8KM:ZNA2MXP;FQV6_,@8!1B>81":++CF^,
PYHD[DZJSU<O5J4'5G(2];#H3FP(3C1PY<EO%512H;<Z%[X%1771]K"F*M=_/JMU7
PB@?&T)7,#8,"V_WJ8U#^X.@PTE38@+Y#G3W(;A_Q4KG1718;OUB]UG./'8Y)YO5Q
P A@H+"F;@':6(Y/!^(J#<. K8U1UH$(6Z0,2605MK$<,SNK/H*(@GQ.]A)3?XQ\O
P2L8HWJ)%L J<M7XQZBI8RRPTM?J^Q:KIULBRG+%FB_>_=:/%R*P0 K68Z!S32+LM
PW:*[K5SZNH!+GQX>9M(S<XP-!DB(2\V[(2*EB#6QZD\U'!RP;J[!D$YA#I\C9M0+
P85'1E+6NK+S0\T&0RJ@B1\Z9YK9G\;KKPIC'7)47#/BA\NP4 =7"! +,51_\5,+5
P1,M+DR! /C$ +VDLV+@A*KJZUNH-W\_KE"2?0Z4/=V25=,;]7?\ZG'KP9Y.T!6UD
PTR\SP'K=TP/&C_Q4$]1K3ZTXXN_L8!XGYN1XP$VT$NT(X[3\!"59X[W#8X.+#/P6
P./863E@;E9E4(&2>2YMY/Y17PVQB2 NR=9X!O(]D%6[O?.& ZLZ1+FW(P>B)E11I
P%@YZG@CRHXR_=9(3ETVKEJ<FUG<3!ZH#;?BX<%'K^V?I7[=+\KCSFJK?U,M^(CY@
P?\JVY]K!8 C7%-T(A$]SFV)^];!4*R?D*E/-#$" UI>.J6Z8Z#E6&S8JL[F(?.B^
P4F%P]+NT?UR*:A:BDV)V8X>533N7=WJ\7;R@;M.)5 920@"GIAX7:\U.#;*=6JEW
P\%&G7AYX<8-6=9X$3O+.K$\_EL]L]4L!)=CFXXFQ?:".-Y0#&P54S5M1%^A;!X 4
P'C_P>5&UEPQ;B1(Y?_U-M5.1;O4X :BS4!=34(3 \; ;H#>;TNH4WI7UDS8BLS=@
P;1)D2G*:SM[:4^ZP@X<X38>H2@3J>,3-9HN1M1H4P!?PG$S, K<9ZR,45GI\]7(0
P1O7%[1XH1U!P%;R01S/S8LSC+2!OWM(FG[C!B)VEG2DRSI\/@,WM%Z1LU<S[W,^R
PV:499EJ!Z =4?<00VS+WW6)$UX"16[C_SMGSQ1: =&@]*DXN8[$YLU8C.(-,4)XG
PWJ@JGL!R&N)4MQ#R4?AH+M\9:_;P*.O5A!9S:D^?AG"C<."]+RB'R#0+7J\7;T;L
P2S05AY-OS5Y![\E2P\X:JXF430^0BV]3\<9KA?^<Y@M U_T6K.:G0W@^%W;&?J-)
P>Y$%4;1^MKWRXD/FE!9U#9.R39^<?(\0QDQ1P$8NJ- O95,RBUNSA&%_@HJ^+7D6
PU7V_\6R6'&_Q4PJJ7?_/L?7H;?'.9JFR!<M-_1 :I''G?G;84KH@#O,/HHP#_CRR
PMFZ2(Y%9*F.M;^5;XR)!9\IU<SIT@W@*\R?5IL1 +N^/$M-YP_:TB+@_);C+]M4C
PV%_] V%1GNNM=E-@O1?&86L0D<P(<CL\^6HEOHXZ#PFN-@ODG\1D'V=%-+%(E_45
P>2/I6:]1 >4N8 E*$PNX1,O%RO(N.NB7?RFGA&1.&YA7S(0V8;-N".!D98J 7@L!
P4VH)FB\CI-59HM7ZT.?Q$Y/>6KG!-B6#9]9$D]!7[Y2O=)-^?VVN; 0EHY1:J+P4
P]2)/,ZEH3-G.&\G+'"NB,YB1-+KWQ7@%ZJ=R:VTCK(>]78\\5.@)QF?8V@,]EAL3
PPN8,K,=\;$5.Z<XR,6 (QGKHZJ@UJ^G">4DOZ.WK0:#TFT[-XR[@PU-X*HT1-+V>
PBJ^D%E6'D21#1Z@X%;NF10K*[O9<@6>3Z*XIA?-<_^0?G@QTEBMDQUW"TL2C[I6Z
PX(C-!K8:4>^$@0"#H N"G+5'I,@I)HU+6QB"A>M='/M%1_#.>[XP6TD7\Q<$>8Q3
PLUL#?2QX%YD%1X)0#ZK)WG$Y 0=U&7Z;H6*6\W21F3]/^<KMAZ4KWCM-E4?[V?IR
P#V>FBUPYMR<:4;*'#%FIS*J$KUAR]1@CJU/S50/+YX#=P=37%;%O']75J=;;[[GG
PJ<8-E&(1^.-2EV(#F$^5 &\/'/[/CUFHGO6N*C[";0"B@THQ++_?%*2,*.4*4%G@
P#+=F7I1'*,DDC A&)1U<$CE?S+728P2^(8=UF:.51-P2D.M(?W+9(ZF)[;^7Q]]B
P6*WC^\+R4^-&+*.&K_(FB8%9T_0#7 62Q)KUADSK#Z]1N:+DR6KX("R+L-7B1M1N
PE1@#\"0X;H34N**WP[CQ;CRF-BT3!#L.9DG &'.\@]D"<)FNZOP!K:3O5\2DK%I(
P9 /;GIQD!C5Z?UIL>WFE)2J!*@ S^L,8WSBN@?\:O,"WO"'7HSTM]Z3RN5=\GM0F
PV$@<(89/%^_C__>>YWK0 L+H?V\H9]6M$A"RAC>@!#R(0'&<W%E/-@=*O!6L7 D+
PFI9A,[4="O_R&',LNBC:&(8AJIUK)2=@>5PL#%>Y:O+1N-JZ#A0$PNQMG0-F'A!T
PK(N^4II*BN$Z*6<DFC'EHZ%DCPG7U^3-GS< UHY:SHIJ4JN:F>;XWQ(/ RTY%Y$:
PM[ TY@=YJNM@(<P?STS;-T^#"^C+DXN0=XYJ3BP0)B?XIM2J!: RND%WF9C!1/0S
P(>DM&N.I6LMM0B\U/'C$?9-"$6S71JH/WG>&44V(L=T!'#8Q9AQW^K_O!E7;A@-L
PI8)2_CXFFXJ.0L.@8-IJ;97AFN_*S>*%H&C$!%G[,0;#9^>@1W6B/'PP=+L.'JP+
PPIFLN@?'BI1!LJ[@W Y*J_R34:?6):N,^>H+/& C3P!O1:<GUUS[,O.%"?CC]?F?
P/\V%J/4<R>SUGS^ZWM$/@T]53?$@7C-K="72^@66+QMX5DD# YI82?=<IDIG[:U9
PD<2RF]DLDN+U, 1N9BE\1Z-#/8!BT!_SK),/!]6\LO6K091J1*RZE'4<D@HRLUC3
P ]2GY ^$06]1X;).OZKX2[!L%^0:P#S&\TEB_&&&;%R%0H;>GWF98"K.R^@5H7I[
P+RC9RFZU4'C!UX03Z_U259FEF&MRZAC4JY3T[)V57W!>XGJ7GG]>JP!7$"O2&8U%
P(K K:W0[7N5MC?7KV#T[2D4,^A0P?M!(,EQ,"#](Z'$]QLT/>/NIJ &&=9>IH/F?
P*U";+/HJ&N<X *)YZ\E3[G'TT!&1(%8NY)?0I=3-!L"0H#]5 5R%-JZZ6"Q-6P#K
PCL?$ \VCIO_703"#T(,'F@7+LV-! NSC5A(F:&$P-GCF?5'Y?2@+4'#XTZ<$WUS0
PK$,"+P-CF HGSRUS9QPY=C77U'B?\84,)-AJZ+[OL-%-U>26/A(&D,+8%,#OC?84
PX54.=VR3ITST[ KR7FT-"P4/,LZ<=,;BO;?FG;(ORN0%A?^F7(LH)A4GC<?-?N/-
P_NI>!(VKH=W?2C 0!$2]4(ATF3ZIVH1M[+1%JEQJ<WU.C$1WGV>4$]^$3G4_Q,-B
P_^Z2B9 ;]X6ZE&;^W/_.YF*1OZ 2F4%!T\M-.#YB350D"> A0X3QN[9:NZ.&XL=)
P+EIK*L&T-G:K>G1D5(\-5<N9W)M3?4!>?;WI9Y WRHAOK\-%_;4K *2&Z64F9V%]
PA6K39G7X1'1S<.D_23N;F>(ISGU$AG&Z\SLL>M+"GB'78X%G_!=Z0[L!ANPG&V!:
P%!/"9[[>I/PSZ>XX07'BA#W;%<Z Q9YZB@XL(V=(XB@CK7*-EF><%77H=]IKV#.[
P#:P6<=6DVD 79RM.<H1+*+$J0P/:MP:MR&'UN/'V>?@V+JKL7,O*P_)LJ<),RD#.
P\['AAH\7?3!4X2-5HLE#H.A J']<; 'N3!K8CF!)/C3P>E:2&&PPRCFVPQOD?]7F
P#7A.P7D6^ZBLL.@I!>4^Y;(M+*R! T;X6Z!J]I30J>(XKND;X/]4I(<"7NR,Y*D#
P4=U5&4*?QE0Y:$6Y9%K]_.GK;8488566P0[77,*@E%1&$&)+8%F3GB-W"FCS,&CA
PHAOSJ^%DF!0ZC H'MO1]DZWA'V7TT?6&7M''/Y8\K2,8S>^?/HP, C#!?7:U$N,%
P!4=M6H9U<UBJ7OL)?YT<&P$FY*">.?;$<A!MP\QNTDC;$.%I*T_9_YTK?5MW:LP[
PC7>U_Z/:1*$<(Y:,*M\D*;<G^&9O'?$NW,P!UG&&*\8:ZH\OQ3_M'Z)GL3<J<=! 
P-:8'B5X*H;M)F&C3B7E 6N(WN:[AZ\&IZF2E9P]?("1UNG<KM*'@QT;SRBN,((>,
PM54:M+>C!H-L%9_*Z:D6<1^D^:!"[(4#B1P"L+'2[%X?7RJ]4*U)T(T)5(,;GK$\
P8&GGV.X3DXDQM\R(4%!(2D))'ED!]B[<]G$:S02PR,K5Q5G05[EN12]P-6Z.6/[.
PJ!HE/J9%X';S>5#YQGF((9!8L.=5V+G:H9N]C_P&5SIGRZ5F!2,N?/=7(?*1RC:*
P>//-;C6ZI2]WH[*>H^\WX@$VK8Q.51G3YY^C#WFEVX_J*F2H7QQRMCMW1G,X;<SP
P,4S/B5Q-E9E<U#(#J6_$%R-[>C<(4K ,VA.KR*.,#Z3Q03A[VQ["@?R!'B##M(MV
P:"9>L$?SCR*<+\2.!"M5@EBRR(^%<?QUM;WT2TV/2O,56$,&^X4>P%!//_0GHBF^
PMMZ"\NBJV[!@1$%S!OAR$#:\(L?&OR.J4'O<M E7_P^O;\M$@64+\88\D#6+WS=#
P19.YG@VJ&":) MZ:',78S,?V@IY.GVS6?$.8+"/+:]91\Z06N%G3=T@N3:69K>L+
P'5;H5KHCC:>Y>AI:I2P<Q<";PV8S?,$,O6H^X08=S3QI1.3#,OL=V+YRKX6_./^Z
P;H%3\VK0YR*U8;ZNL10E,@Z_[DR[@.]L-H\SYT6ZV;<HFVG7*\(AU*T);W2LH'AU
PF@=)UAS)*-R%WE2W(=1\#I[7]73EX)C9& L5>L$@.-O>Z0U*$1(B2+!K,\L07[&<
P+T7[>38V[OOI48^=]K9W4=6:7O)E V-)=ATFTT'$3P_7*.K?;&$T(6P0@[GABN!1
P"KVB6[5/-?-VS+0BZ7.FG.!'(]X%RYO+\Y<>=GZO2SE"]S;<"N EL7230(WQIT@V
P!J7' Y,GT2#'D-&!O'W(@14L>5_6I_0]WW>9E^R#.P,L&+\?^Z$]'CUB/U]^BXL?
PP6#N.2:J]R8A0W@ /M5@XD.HS\8T@/DWVR%/^B5;D\Q>Z0=_-2F/28?<WWXEO3[>
P5E\IC;^$0$M0)J-]#;.0QT$2@_>+T.(90(8G8[\IK!S6')X9M,9\\-5AWZ)RBZ7#
P6"/^?&=QI5$)MZ3<NJHC5IN1,;&M2#""  D.P/$#3RP<;QZ1$RO-\;U8JH$&UX:B
P8[!1D5)S%?-JJ;/+,"=YGX-(9. 5T7<IF#W0G(T^45-.(OQM"F3C1>9[L8\XHG3>
PQR,$3@PX2,I*"$[C9 27_7H_H%F6%G2G9->"A%7%YD1U&(O^<)3N[]=%8;5U9RY[
P@7I.?X__]7 $/Y?.A^D9$ ]Q,1P)(._%OPM"8P(OZV>>T#1U[H9,UD8@6[1WK/<^
P#P&=[4:2SR\]UL8AMVKTMJ+3R'*(OP5J=H5<>8G'V?2(5)%+.NACJ[Y-,RM9MFGX
P : F2^N]*./ 9^/YCA2@\;,@PL[K3G3,YC__%A_P00OO^MVI99SFE0_-X,U/J4/<
P+*59N,*]+JP_"+VI-L?+98L95O^LRANX+K?7[RW$$GK.!/4DH2)#,Q-8BQSX9I"H
P%O#R0=CO#^3!G!&((M4J[2.IBAX&Z'&_ZH_@)4X T"K.H#'ZOX7]?/0X?/T';@\+
PH.#=+LX/$JCA.X1#:.'_$F(O7V:U_H\ATC(HT6DTM GIA&K"UD1?:%<0M'P5P:0?
PZ37O,"$2MP,^P;MT")U<[TES_^!%LI&]+J&W?]Q.S7,:8B="8'ENV7:#Y.<97'6@
PX2L10.4J_(B_'X15OSBN]68U6F)<A(SGH@[ZZWU96#.(9O!!Z(MH[OKV>J0Y?5@D
P^YQ<ESZQTY<1#P;\S"QPJ_PKI-\BA]S2*\CGU;JOSDPFX'9+K#37CD6U!RF;D%Q1
P)R_2O,Y6<:Z'R<*U[)4O#ZL3P!D/.Y6X'9G8&SE-4\L>8BTFDA479B674IMTI)F@
P_RSI3\_,;\"+TW/CTI&LS1 ""]IE87,/>@V3^N^=".?2&<EDN5\\5@$K!45V 6([
P4&;:*AS+X$W5*R!JO,?"Q;+A($E-Q4>B($?KT/'\B'UPP+7T#6SJ(J,/2S35C[YA
PV04M'//36)]7I(6P#!*8[],:S>MIS?<FH(W%1)#RE)@T1E,#W1Q;I>R#Z=.9$3U_
P9X #K07;FZ6K(_X&_N)]C!O,@#>$]\#X%Y'#-", \/0)CQ?>AL38"-MO@(3Z]H4I
PY;::P8Z$)):YM-<-\/,.>/@%-XVPU)XN7R8I!(C^HD0Z7&DR;>E.*'9"'AMFW-C+
PV)B,3&Q%^@IS-W:TBZ)1#"3^'L=JG]!Y!QGP]S-WU4HYIL3U]F--B4I,)O-BUY*7
PS-X4L8/R5_3((KU%0\5'\)043JC#1<JY,&2?^3Z\T(I<.MD :$G5X"C ;4S.5%W3
P "^'?BK^7OYZ0::?'ON%_1R1=*.9U9PSF;,F)9-$)<<?2)5?Y9AS6A%% ^8AHEEW
P)R,*F2C*; E-6&5IZZJ-O<:6G 8;Y"4\;O#A=0WK(*,J6L6* ZF-_W'0I7CG]V_8
P+?H;>MI_GJ03;-V!350,:UW_:J3O]-#&8I$8V=U_34<N4-T6ZBR"]/>0*NO#[33A
PR,KF$@U'1\!I$U2[&#B%XO@KQ_^VZ#_" ,KTR3XU,-O<FSV ^.W&HC41,!X PP;B
PT&N!3KB&YLU,T\&[]B9(#.%W5 DR*'!!KN'25M9Q(H1'<,3@!LSF) ^(]4BQ2D'B
PVRJNA &:DEKXQRY9;"87YV8 F,YUTRXW\P,PLF5NT?K$E2QD !YTT"83I_Y4G[H?
PP)^T&&>*\" VU#/-NG2 /8<9W&M!G)I#]WA5F.:E*5(D?=J@RX:5G-A(FQI*2W.-
PG86JVQN!/^X5TDWX#XS8Z(L7?KP@8+-%5497.\%O2(J4\]/'ZP%E(=U$IBB&''5 
PA<@R%NZ:[DED'-( ($(33-,3S4*:3<H^8>(C%JVZAA6V2NVX2X1&UEG.-5@&KCV[
P(F6H$/Y1U5/5IU.\_,IK/0.M3GA S)W24&M7I!:?26#WMX4;*2PAM+"C3I[H[!,"
PJ[JKH0;\)IV!HV..4\/NYF6;2$Q7N!L=C8[E]<AX"31,M,8EE98-E*'=0JO-9U=0
P:A'Y7/9U#\,[BJ$<XEG?CY#3GZ1KH-L&S!<22UX7'5"31>(##S]Z\ZV0KU-6:QWN
P=]QX][O(J\R:5^Z8A^'P99C;T:Z1,X^]Y$93V.^^3I&B$-7*@ZK3W?L&KZ8IPJ@)
PEM)1M:.HP7ST_^ZMG::>^%PO,6)B"K\F5[03S7(Q1A^*S7@?[6!\6I_(?>5L^Q+/
P"+-3T5$""[V\4<W5);Y\,@-^%$U-G[$R-\&]#!"<!K88;&JWXI\W^.="H++Q?%Z"
PW"M.I*&%2/$7R:7@TE=PL%9>M)Q_;P/@#W[_T&4O9W 8[%=^=S+<R9VF(L<1_<;,
PTPTTW+N"OLNBBITKD9^VHH7$<N]WAJ1/@^<T6'%<:; =^S##NW\3P<J; T=18,DN
P4Z4ZQ[0CMGQ-)*R'W[;P-;GLTPI\36KIPQ\_X!N5V)Q39B<J[U16B$N#N^?H#W9S
P,!S)<?R ;(>EPWEV#KK*6?M4<#TH21RGZPJ;_ZT7W7<SB1WS<S?7U5SSY>?X*4LP
P:+X-7-"_SY")>(MI1_J^<H)T]"%* = ^<O<&_Q7W+6<XZ:%KE%H]&6WY3H[J=7<X
P6$7TTGJ=0(G/!+)%'*G/$ MA 8NBV1MEEP;:%B]1SZQ@I?<%E[TV"\FXNMLDGQO=
P3^426T!@DR(;<TUT\Z=E1!DIM"%7BUITMV>]S.US?.K#H\G$4CP=@ACE[6CUWF$^
PF2A8)\+F*J=I^)95,N9 ?GBY5IM@IE0*5.;;YX\8#6-24:#8#4[J4F4<O])DS7!0
POWIB,EVN)*&1Y(S>IEW02V/EHD&5]'0._%GOG$Y \S&_>)LI](Z\*A.HU*L[0(^E
PV^>=+1BD:J6RE8564/'\VT$Q5X@[D.\6990^A67Z9B:Z@'!6 ;TPA=UH;RR0B:O9
PLW3'&CI'OM1I$Y@DDYZ %$-)]55V\YJD9\2#HD:KZZDWZG'@F; VV62:J99I="MF
P$@*JYV%C=-!_7%[, !$X!)_QLJ6PLJ2>O1??GJC<-1\H1>6.0*4B\:R%"0CPA#:$
P+!;<E<A<PA3XP<#>>9/[KO-.47!)-QIE.H!*TT^K[W!:1\5(?EZ=%(R&"-R7J7\M
P1\-)ZLLSGOL(Z'=U9S9'Q_2)[)AG):*_!9NN-1V.=;7M"%7N/#^FG9BPPLZ++ %R
P8Z#7&GQAWC@4GH=JH?4>V*$T4^KJ?+\11A8<1^,)U:9@#8#O_[6F6OQMIJP#)4/)
POUS,4T>*-K6"Q92Z"@J4*]RT7#@%5Z@6_7A?]X6R&G?XXC+('NRWAB5$K0B?ALVD
P03X$!@3Y7UR^4./C]LI5>J<9ABJ<.$RI'U7;F0X3V'F7(NX3J3Y O'4I[>+%E'L&
P0L(%P39-@M\B):0WDHX0&WFJQ2.M;W6#0:+T_G3Z!_"R1RE[>:Q!R$3;WE1I@%9:
PI88*\&>%:?4A# 6"$:%6E7G,2&EI@P/!928D9(FGWO4M_'E_#36&JLC".NBPJ"[^
PJFNK1X+=EC^8SI:S^[RQ!D2(<2DZ$_;M!>^*[KR&G!UG#?2Z $ D<R!=MM83FZP9
P1W9],:S;*P/HB5,&EPMR^V E]@OA6PZ.DXL$S%:1*&]3W_YAUSG5C3%VE4>YKU30
P4:S_);R>% .BW9<(EQGMR9-8E_QVB-]8508'O-WD]*V3QK??3EK:I(5L1S;T)Z'Z
P$];".]3S= XPN;2J$8J,=_DO\,?%5OPCPL+W#.9U'NP#18CK[K2C0AN*58%S"8:*
P[N'1%V5=J,4+>5HTG\<RT.;+.TIWO2U\;BFSD]*H"?5^9>\NL_Y!5X\*0M!AU&G-
P$D9:+2P_8(4?9W*?(+P>XS T4(1P05HP^OL@D<$&"Q'<8X^(#%D;R*@F0TK5UV:T
P6TRN[--HB@GAN?A&U<8J>,T%Z$?,9;B0@V=S*0+X+^,C:O#>,U:(UE[I!%'\AO[_
PV1*"54+!  ^GI$;/\[,:VSU1JP=JG:&63\,LE769=CJLE.<]+NY8MO$!O1%/X<%D
P.AUQI3.F&$E5 ZS)8YFANW#']Q*J0.##@MGTA?_UQ6[KO481O+5NU6@?59H>"D-_
PQ5=&Z-8@L\!D]]<T2X^&EB*4N6I9K3(-*,RXP)"$<[2S;44W1J)5(EY%WHT^K;>W
PH(3%>;RF)!(Q1*'%.SUR)R.V+6DA.M'S5&#IWS?3'<H@;_()#RYQCO6P\!\?GA,K
PIF8E*S"-/[+J<ZW4F*A$<[4.9K3CV"=KQ@GDD1D5PJ7*;NRS (Q\@+?0Q HO-K)]
P32.+PZ4.,V[T$\)?HW"K+)7!&DH&N_$2/H_"IU9Y=$I<6TK,"2BXI\ )?&X(JJ:-
PB7.QG?> JD77^T2LS TFV*#YN6YRW 7P=(+1_1HP/8IF($O5&O\@TU_>+*GNE76P
P=<2CJ$MTT<TH=V&5D]EWZHF-<*BN>D&5_S!M4F8QEV)N!$NKB  IO17&L[&>I&Z3
PWO.XL0-CR#2Y[23\O: 4 B<,M7K7DMFVP\7-?B7><(NM7GKO2)$(ZGX^ Z!-9('I
P;A$Z@60[[W3D?L082#AYYY*GOO%ZU/RO3[^.CP$Z2:BN+X_'POH ]70O<16^R[?1
P_R@X9?3 =X+:G'VA]Q?6W]Y<+2)EL>G58 -YENV\5Z)Q!%/G30"M;$TS)4R9)DJ)
P9!AH0#OZURW[I4OVC'=7<\RI\IG"('P,' SB_US*F]=$CWU#5SZLYIY!+5_Y-C4<
PJQ5B0;&[#JJXH2.^$SYD&L=HZD.PFY3UNR2"M;PO3I9=-SZ*K5Y[993@+Y*C>\]F
P_)RT();7S>;#M[OFN'V+/P'"T4YD9TFV* K--IJD2'&137Y ?(P0'S]<\<<IDCED
PA0@ORXCD,LBI6>&%!A9R+>_H)0',"'\I4F/%DD\@-F4!,P5B<+.3K-5Z(J,@^&P7
PLY8Q <=N/K58$*1W:<MMWI5;EE6=2:7'XP.E_Q@3HM+D?A1/.[2V="AU$JX[Z<I/
PK1!3_]'DE' (6PUC]MOO\K-JZ:JT;)(V_[?]%9+!-K/5B(6NZN9/IHOFQ0,;!) (
PNB2YC^=O]3WXY+WUS8)0'^.>V@%G*B7DVJDF(<79J<UM&P%R\?^JR''A.'TJ0]-1
PH'A>RI2S:$7V4"A'\G]=2$</&)HF!Z;*8^)T_&BCS'B.C&'?)B]FY["V+O/M(?+O
PDY*O&S6E^1,BB[#"31ZJ9$$W%CE9H=3K"YV/WIXFC^]4F#J(#^!)ZU1-,/W)^:^3
P,A:R'6%$U4 2KEPX=;V/@J,'.GK) >(%&SAC@)E/)^P2@;&1SJU*B]A.V6^'JP[$
PC=D@CSW1B N=/W?=7Z/+ C/6+>Z/=9OZ,14HGP?3W5@X:C!;N0IH^[TAII]^6OY2
P#^_GY$H\[,6)(F'$65H3X59;CNRL49<8)M*G*]O=Q&GU:*K@PO"]<.D&OD!NV(J)
P+/2LZE#5H ^T>LPS:,(F'MSMRK'$)?VZ/FFAYTY7WS0)F@;#FPHEF;=*&JN8^U3*
P-_SQ#W#:$7I/'<W0J_@ PS!G]GM'N]=/.2JH0U0X'7B<M8>'V1"MT_ZY6(2L9;VR
P:SZ5YSZY,$!_R[NHY >@#P\?+LZ9?BC*R<EMX!ETX5\\^R$1+GXL/P4%KMW/_7(!
P<QAO7/5998"*IGR<93H8TE55.\ZE6-33A$88YI0FZY7^6N1:(-5:JB&D8:WXBT$9
P7]4ZPU3<@UJ#!5OSRQ!A/[V]P).$'U>Y#%>3R37;+WS__$.SX-_'2XUVNM$NK!;C
PE\(2#5/<\Y?U73N:L[\^[6L#/@< -'&K=F'HF>BI%RPB=.#,SLK5!8ZEW-)%$$!+
P)B+!$UGEURDD0QJ1$OYN3D+3?;#F1B^BB7V QZ>*MY8RJ$9K/&\F[0;N3>4N"DY;
PLP.2)=7;UW6'1+^&D@:G@*G%$V0*GPD0<0\1PMQ]676YC8#.O%PZOV8/D_^F%$]<
PK0,"O*!Z--Y(%3]DF5Z2))1##SAI@,6SQ!+CF>:*I00IR1BZ]^.:T"'-XT;QT% 8
PIP)9WKKVG,TK+D0/"+GH:4IE/DV8+@7[<MI0^PX#[MR+^$U-$Y(N="-6PE#+283*
P,P[^%&$VR2CK&);+@456_E@DHAHFMV<3<(YK0?DLKSV>4!-@**:Y21L:*FPDSJO:
P+&C2PFHG.,O'.#YNFW^XRD]HC]:5<N%GAKKO7VTYWQVV;#O/:61&E4^[,S%R]4*9
P41GE,]7]#;ZS^\C??W1!T\&<"8"(D5DH"E^$^RVH6E_'$ 65,&#3R%P[8X/#D1E\
P[1D,\$=AYP;MAF<.=;KY!:?P:95H>+")BA8&&PT/ACO6'G06*7C5W&E(:+=X7"SD
PUQ*LUX6N;)X)&9^$,Y=MS*?[@]G%NS<N P8'@]]E6WN=8W J6B&@ 1T$Z71"E.2C
P9\*\];[:'E&39@_+7$S_33,C,YY0228E*^.J2UMN;8,SV[ &G7RC%QN2]\]?D$-A
PG3*V0X$;^>+&L$ID1;90#@^I$%F^""KQA.)P7*M01B9:I!Z]J_OF3K?JMY%Y;2ZN
P76GZML1N6P*HCF8!2XC]=P=KW'O]IKM)MCCYB-8B&ET<_N'EUR?A(\*6!'P"IEF#
PT=4D9>N4:.#(?R=]UED5=*$4RPKN53[V<$_^<%XQ"Y$C*!(%NEZE[4I?<$J@&Q>C
P_K:B476IO27S!Z!>T:T4+V_F7T%_A_7X637E#/\_[WZY$ 9$SH6L;<03S-Z0O(-6
PF>8<O_@I42YMSO+]?O6T'5PJU)Q8ONAK-&_^0+E>^T/W2IP@O+S)AH'/A-ZKF<QT
PY"\;J@),:J_L@@Z"M'OCK114JG*IL\>"'@M##0/^IWM.?J;UI,(O4Y<!A_L1F_FZ
PYPBJ9KX>M]/IJ%1*Z,KW3'LDRN=5N)XV%U!0>PFH0L;N.>@?U%%^=Q.$8W/FE1<%
PWYGH;UOD1EH<[L D7VNWQ!!B\C+_#]D2&6K6S;&FNU+NVGS\TXMCAGI>*SZW7O]K
P)T+UH MK*DW_/LMR?T=&*R-^SD>';%+UP#7&V\P6'9N02XU$B!(R4V+U84(99!O>
P/=]N1?R",')4J8[6Q#5F%_9$W+7L,7DX)(+YP=H%^L[3HTX:'K'V../<"1+2%E5A
P#3"6%XY-GJ3H7PFY)PJGV=LKFYDVWV#E-Z"L+WSD/J#Y;&-5#+?^,EQ+Z0/V(Q):
P.%EU)FZ^/8UT:)W !:?>![Z+]Q]FF#]7TSFH?/#UUPJI:+Y-V>07/NT\-9&<=ZB8
P,)Z2<XD_:'4)\:V6Q76/KT-Q7O_@HKB8O2.,=R)K4X3:4,=@>-<45_N%$UEE1/!E
PEKE8V$#H$'G?-H&V#IE^_4?I:$"P?T"7+I9/I1#CJ('MUJ>.U&N3CO#T>+<%X9;Y
P"'FVUWK0@6(!^6+L<F61=!S7RT3.IH]Q=&])(0'9;*@* -:*P-55^V-M87BZ_5&9
PBU*P"#*FW\)NC'%!E=4I8E%Y"O/47F_:MR:<D#P4=X<>O:D!8I8:+*CC?Y*'BM#;
PM$6TV:,I8CNR8M*'9F%'<04.^*+]ON9D\VH]O;)8J- 7+BA[6;(ES)B/OC[QW"6*
P1%_PYVR=FLD^O>/HB ^"7Z 82'I!H-",Z48>22U$DZ1L$!DO7C;SJT]FBN:KK594
PWORH?Q\UE81W\K@N93&(7*G$_(F+<)V1'Q@!4N6HBQI-V.-)4L5?R>7&V!]-Z!#,
PWEA,A:P-W]_2P<ZJKV>J  JXT^XK4$VN3N[S_S/W#:0&W2Z$\3":4OD 2(X(.IW.
P(G 0_&2Q@'6L(/RHYI'<]Z-P[>'6\TTS_>3Y#(,A#<;LQCN;U#J#J0A 3P_R%^O5
P%>((S;M1#EQ4\HS02TKHV\8H@W]67?FFW$]-^8GU4ME!M4SP^0/##A/\Q["J<COI
P)#GB85'44W9F_H2:S"=I,C\HQF 2V,><!B+["G0,;2^Y9E]T5.$,'VM19[;V1M%[
P5",*FTA\+A#C=F5$ -I;9S:;GO0.2-#"[KUW+6B7'?H7X<AV'B=R_Z.<]R(F*3W@
P=84M=/L1GP#S-ZW! _J419&X[\H$T]0O]B -AH^U93]59[P1(T> ;><5-D8]HYH.
P4"^I6&BL/_^@AM,N+N(#*2JO31:N_%TZTC8V,7VU4SDO\28RG:-NH>V_4 Q45LK*
P1FVOI\D<N?-0Z9NZ74#LN<B0J641U^I7DO_/LLXT6/F';;8UH#'@P,C!#3+LSTW 
PJ_B%CF>BY<E%5(@E1<+P:!*Y_?W*H7,ZEI<I!1:T]ZKC$"8&8(7VG9EW?]".\4-&
P1S%5"8 6+LN]:S$.B$XS"UTU%1_/:9=$]+HDUF#,5JG$R'8RR1=VB'E$6R_HG#_"
P'F4M+ O8R]\OSZVROXLA&+<"GHYF@$_*J.VC"3:CHX0A&S44/LJSQK/4A6CLD5GU
P^\VH91^GK=K06,>JR<+9^5QU$HD5M/ZF+(3T'_CQ#TH0IW!F\8H6=Q"VYN.G.SAI
PM0(KO$0Y1$2])% W@V@Y$E$F=G;FI3^US&7BE6A-4V)JYA6[5"O(FH=5FK  =@?,
P[4WV9(JMLI,=D-COFKE3E;$6%]*$,1743?7V:'08Q>RL19N?1?)7U]BRA:@93B%B
P,8]96@%55U]BKCP!>\+&"/J+>NX[]8=MUB):#(T[2"Z%"[Y7S!O(_EBQ&"=?DP$!
P@]R;M)SNTL("28V?V4"F.C8\OP6_1:5RTVZ+4/0]FVY$9@U.+L7'>:F&V2'WN<D.
PY,)YQ ZJ@KZT\_N3-A-9C,(A6',Y6 _=<_>Z<1OB9?:(<:6VC\  EV.,0&1;Y:-[
P99D[#_:<_SHKG*V7:"&FM>7J"K8\,I.#3J*44.?3P/JJ>0H"N?ZDP3<Z?!!%LZ1\
P:4KN0Y9/::LO>)EM(5=O.1\AN%_94-UJ[7!>3,-,H5=)*%5]K#_-?/6C^4>_/T[,
PPO@@*@KX B";EA2GW9^G98O&>#/&2E2'<%=%J\<%)7H6&](0E/\;TBP.JLH?,$XP
P\E5_!%",S8?U+=Y0C['#IH8Q\=>XQ4][5P[[5RM$ ,TP8VX9,ME*SDK]88H6*?WL
P$(J?,D(VGYW_6@7NM+>A[&/PO:KTPU,(;-O^1K;MI?5PM"-#SDW ? !/FZ_T;!*D
PBYPV,]@ =AL,.Y!#T[OE.;E5_>%27M?5E(.GTLPI7NO6\#<R1W%AO*OAZJJ144QD
PV!\&LL,$V,F_Y%L7$RW;3!!5-OFO"*/7EC'UTF+P.,;QT_3PSZ#M/*VO9UA%HB_X
PU1GB3OG"$7>UEHT%>P\9W%0@2%,HE,L;%+-2H&]\_#JWOOY% %0Q?1??"2G7EH)U
PU20R4]>1;T*-:F [E)N!6G/_N?#Q!URW1, [S)+NZ>B(3)J$S5"Q$DR?DQM1=+P;
P\$6"HH6I%K:[H"\ZQE+\X&\7XG>?*R!+V=NX=F;2^!-VQK- HFC06C84W1[R<0I]
P*P2?>AJ0:(KN\' 1RQ<;-K8Q<^UFG_!2_I_D,T-<\ ,/@D>]QC8^Q_U;90<R$01$
P=8"M*4W+DZ[_7N@W-&>N<3U&M$;;*("1EX]=?'^=IMW'POP(>PQ%XZD^YW*/U+CL
PT//<GX#UT90=UT3T4EQR4<B_Z/XZ) AO-LD*$V[(. F86^8J"QDOKN3E!7?]_&HF
P"ZQ\[3)JP',M^T11DBU7V=Y>R-\&'\#^2AV^E%  @R+'EF'^=UF?AZ=6%8EZC5KX
P%F Z*S(H-G9.,A;Y'=SG:X:_Q%L4O=-4+4_%<-72*1./\6RE6.]3%0TA$>H,9HX+
P[J+1"L!2XE4*0 +77"KZ*8MB#O%A[]).%T@;X>/87+20JJK<I/6"_'5#'TZ?9.Z;
PQG"@ZFFJ$_6]D*.,%!Q32RBWNU2/:=HE!Q0G$:CU;!WQ+ IG@+:LG2H$2SFYX,-6
P/66Y<_C:C?D]6L.;"Q>5@@>KI>!ZPTF=#OX<X]4Z"#66(/^X_EZQV#^_W$8*;UF,
P:""4M3//PQF_#?Z>'T_D<*4%)<FI'[\WL7Q:#;"3R^\1'FN;ZQ<-R%QO,.3&TW\Y
PRD?=%R]<6LVC8-;=0/D&HH2C>*G"'J^H^-8F7R+%0X";NQ_T"9G/3ES%$;D$I5P 
P7G+^<IR7% \K0K]@"1H/MT1,(0-2_D?!C@Y,++[\FKTU"C96D3X.!$%)#WA 8%5"
P_6PB"&6IM@;VS8*:0;3N].CD+^6.<*=H/-Y[RI?(Z30-'W>'5GVL-!@-$NZ1I-#^
P_Z$$B^?I2L_!S<C\NW9,J^(1T/A%S5E@F$D39 %"Q:6A4:A%C=R_5YK.A2Q!?DZD
PC0L@EJ1X1IL%U "28MS]>!7!DH,:"XC@NA/)/FX%+Q)PCS.AU5W6R0/H](>TCX?<
P8W]:.=-J0N'<Y3JN%R!EB0YC04.0^^WY3P+$MXKW8+^[<ZVWHE&O[([4Y]3-X[QE
P5&IM='^!U;$(:T'LP5P>5ED P]-^@2<B+=E)-XT-?AW.IA+95<40J/OF:Y+.CL[#
P_^E\I(.LLN1=:771'^U*6!.2:UA4'=>'V$2@JIDE>=,B%9AZZ[Z@ ;C&GF&H+V>%
P7G^238H_%SLZQ10#@=O7XC\\-#>H0UKF.8!MYBW@=@(Z;I7K%;Q2'N)PL-E(:LI^
PV<VZV-BL_BO7Y%$!S0!@UPG=>G6D?=(T\^-[R>Z"(L5_NZ)(5]7=.[R.J*\P'S(C
P8U$"Q#9@N 9^E72 U[5G)W)@((T<3OQTZ>P((.^)7!:@ *$)8W58YHF'("!,]=,@
PM$5I#YIW"A$G2\\:E^?J?X0"IF"S5 G!:'M=(&'62<027!27!@G=8#V@N@T2D'_8
P9P9)G  !]X.A[-BP7GQMG+EW7U14_1INEC8!T.,HC&CV6:]X5MO4=LE3YI*BMNY6
P*ZP*(BZS[3:E$%-PY"'LM32DLDG-$/"TE.9=Z]6;FL9SW;ALT_E*P\<%DB_:=71_
PBBX\LZD7+*-9F+]GJ5,_L?V>_8PPY>D*13J;_K%L;"5ZD\S/L/$^!3-6_[I]IT+N
PP]P6VK U<R\5/.B0E;B^T'D$J'WDEZ0BRO@'GBT[6K%PYV*/L"B@XKL+&DJKW6/4
PQ//I#_QL4Y8NH[[(N04+A4^8X<38:?6ZLKXPG-335:2<2CTV7SCF#1WW=HVC68O=
PY^N$X7%..]4_*QZZ]T,>W-N\'1,#F'N&<"?4]BJ,=)$YI.6NBRH _%L0%>$%R!\&
POYB-1&VO_JU.O^5E9>J=897P6:#DG/'^Y0.0_M6,Y=V/6KX+:U^QFJ:)66!$_*Z%
P%G-]4C$FS-\]@X2IDX"L[I>6(-G#D3CNV>(,*'*^+(?8&0/-/O)SA\C5@\UKW6=1
P_37-4OCMX2.IJ4<=O>)9@56'_3W[ YN3M ]4&:ZJAUODG)D<@?[]J;6T;&@\QT]@
P*.*;%$EW#CK26?W\%.-"Z/P:QU5.=F62\$&33Q?!=:9(!?NBB !!@F(K-J88-^%J
P# [N4GK)^!?/IU\$O+#LW>%8=AM,?,^P(!7CAT-FF;JSCU,OCO_?93N#IN2Y.S.%
PCDN#J^>NY0,_W%?8D6%!8SC"=5DTR&&M9:- =B&VD(:AG*%3&S+N76\4X&BFVJZ<
PKOO5U+]"'3 T]TR*-T0$(@]HQLH%EP0O)?ZAWE\.&Q"&\7/*4(!*.%G[NZQ ,IAM
P+Q)+A<\$Y%Q)=5?QR7*1>] K?&2=<GHV8FG4ZV)BB[S[;SNR/IX54)9\M*LL>Z(A
PR8CC$Y)BI4!^DHD!B]5-RM%LXQH.@NR,S#TF??@QK4[A41.OP+:+H.9N Z>Q:-C"
P=50QO]3QB0?4:-)];'CIQL%_X'E5J.FR$&M]_@Y[RR3/41X!A9+)5U>6Y'ZEXAZ-
PWS^CZ1RNTWL!^E'N9M[R44QE3@N#IA_DD18J&&AJ7*E4O$WW6##P.$,#C5["=8?U
P_?R*'J=]([B*\TM?8?#%F!CTW)JUI?@$CA+KT;MQ3^X:G8?G.?4K\!F2UE2"S*"E
PII@+ NGK PQO,C.'URI*=U/Z@2DBD%2 2WE;G_IYA3UA_T,F#PY:MD2CQ(F64+*Y
P-946G'Q!W=U#/(JJ:F"8T&2['4/G;*9ELOI+%K]M2FE_T3^_T<DL<R_Q- +#\.$Z
P=F;0&^Z9)E1E6=L@M6@>U9U(K; Z_&-&>I> _!N3U/'!:,5)+\(=Z;JGC>XZU9R+
POFI;05=EZQ+ Z>DC<;JF2GK7\=V<,M"%KF"A531$68.5QOPW$<7& F[BB*FBWQ4"
POZF"_@!_VM@[W6VA78\1$'-2V_<:?_9+]XZJ,CS$;S2:'S+L1W![%MW*,*+XJ1P1
P+1"$Q*6AH6^./R'<QLJJ8#<HRK%G/):-0#Q@,*[:W*R5M9<:O]5Q\_K1Y:)YZG49
P;5!A!I'GF.\D868.!3M!4QPL$6^F$B.T=/,VO+(ZD6ZXKMOC,6WP-D27(I:F/DE2
PBJVE^Q*"K^1Q' >5"I V+&C*6/+P;+.,#68+-N"&^$(,-]O:G5A'SQ%W!&S!Y<BS
PIHE-DT3N\L&!LV^%_U]HG4>S?,X*)MV@-%8-/B"J?<^A0XZBX-#(LXXKJYK)=9X=
PZF !>W6HK*]8?;/J@NYMIMJZ90S&FQ(X/40:S"H[ WSQ5/^-8B@'>M1*S:+'U!H7
P'](F%A) SJO=^&PRU*)V>'JXJ0NNH'F#4F>KG<X&%UMZ"GF207U_:BXT6%&7F/GF
P!"*M/HSQS(E*"IV$D<_V9^T3\Y3\A0SF-51,1.=,O>[*/M$7=UOC>)U/N6@+-KL4
P03CN.+\-$MH]1.WKU^/BS4UN'I4/6^6G,PE=@:*?(PM=O7$GE"50NV>6B$!+VW;I
P>5.\P(D)9B9I.<SZZ[6BLJA#5+,<6O]@"V:J3P8_)Y-NC=WFS3,)T!3(RUN#55X]
PX*;Z-7L\O2I7'4],B.:W+XS._JQ-\IF"7O&(!85 E%4C"U@##<)0",^7_3Y1Z(8P
P$@B^R@XY0MRE$6I2*0T_P<2;J&C9F$Y[-&/JXZ_E8S=QG&<:EJK<1[/O5US#,N99
PN)AU#SPT]7.UOM&A)"TAWA [4W5CK\\C9AC@ ^O26R8+N:<=6!D'I/1^Y8QH( :$
P#JK:12&W\]W_H=^3Q8-@<'[]\? V=H;N,$J,<&ORAX^E23*.ZI]/M9"T]1KD;09 
PM\0Q]N#V@FR^I'M *P> 3&6DC9[?1*45\Z/#+-"W#!W%?]>IWV>("W$<E1,.L8W1
P0\*^?GQT93I-XZ2MZ*Q#<A8'_-\@@'>>T#]L\:ZQX/<>#DMYW>;4M-;1<;^<CV^&
P[G^]_CG<Z3ZW5I['KXM+_TE:16B.) 1P]FH"[I8J-_!^XG>O^8KS8&]7",0H1CS%
P[C(_NRY2D,,H9Y9;4U_J=YU)[:B0>69[,D1NE_;H+ UD;)O:[@YCU:Y,>R%RJD6(
P%O- IEZDFR[V8:;V< E2-8K=[L81!VY)#\<P?N#F3#C,<UZMQ= :DZ@\/AV4!JF1
PW^,-!/RJZ._UREV,M7C2]V6'Z]T<+N'X WUPN2L?7IK5>+!!N(YOT^0(]9(5*DH$
P.YMJSG9A_L2[5%ZK+N^X0 HX'7]MJ.\6K/1Z*V6* _\]F>>%_.27+8+;67NN)+$K
P$J6$ > %.ZXS=T8XUZVS@5EG.8I@-$25:?D6,./SJ#LADH(J0J2C"5'@<K-\-T?U
P W"_$)GS),M=*F^G[?JRXURNWW[SGIYWCM 5FOGW0K#;M]!-WO#N1@7 "S+$- 3A
P26F+W\-(2 0$JCVQUP"P5ODDK_Q+S(P^_M"I2X4UMT@.8#7+*=%U9R<#H=>?E%=F
P6KWI5%M@\+N?;\W@?W279E^1M'I3]'V0 IV (V)H%TGH9--ZMGPP93FH0../:E^_
PF>TB9#Y<9>#AI<L+V$^T!8V3S[2,ZVYQ9*;W@A?D?5<>0S_EZ#=>'^D&'>.5C!=1
PQQ_BL@BWZ\4Y1R(X"OTKS;A8L-#GEJ;;V^C&:V] :HF%_-V9>Z7EMY04FONV]I 4
PA_X_6:*' 8,LG:V;:OLO"R5P2<X!3OYQ\$$+@%+",?P2(.2A<S))M?X=T$^.2G7T
P ."$)%D ;)7==$D\0U#7)^[RGP-B:#KFH3TTG?8L(+\_R HT><7^DIZ%/NJF."D+
P!A),(F"8,'5O:/Q^$U&RLJN^IOI' /R*[:6WMV(92C;V-4"5_1K5ZH%,/*>=>:Q=
P[\$M$1$,K>M  SAQ6S,/@B=#:B:O^;Z/K>>W%B::0;]_[LIO)<,N +>8=M)7/9!]
P1<CD-'T81FOFB#MKZ[7F%YD>?#Q-E+5IV$]G^<'/>[SY:HT4(P35Y2*F*=NHA!27
P*F#+$@GY+K[L;_<-V/Z_W]H DMIX(/JA!F\(9GO'XXNJ$"W_Y:MC6,@4^$0B5 )"
PJPK0(MZ0%^CD\;<EB>#R8Z$:P3T<?0G]"+.6C ?$.ZZ<E9),OQMOU<\?^)7U98A'
PD70?D=:UJ,-#(COA:N!?&S -M))Q$D.")^<B[J^7"W'&U]%6O  #1-,8<\ 2+2'$
PHXN.9#H.CIKN<HD(QUZ3)2Y4-).K-=NLED.G)[%(.??0WSG\R39INOIR4UQ,VSG(
P#0BPQ[9)JPJ'-0OVV'=BEQ V,E0Z8V$II#=C-!^=EP7S'%QQEJWV=2)N$\RB3FU2
PUD+OF&YDP"9=%A9HV;%0&$+649]P,NX6AF)7.G76+*YC@%YIK]KU&;>3#/AO1XRV
P.Q:  7U"MRFL />P\8<%UG0;+#1QPG8VN:D''FW]5KS[K1B-00%&E[=30/S23V6K
PC]O7EHV-8Q,GO4#\@3IC9P=;'!\;HE/-D=<5<PRP"JR\G\&!G0WH[ U/J2!J'56>
P5M47<=ZPEWDW&\^7AR@;I6]$3'*FC23DR;C"<(0.^&$>)O=7LRE.7#<GDX/AL[0K
PO+Q80/^D>UF*YBH1#(WS$%H ')Y<@2K% J,6.449#C5R"Y;2*#7L46(J1':5>>A*
PH=2@\&.G;CFK"Y#YX?J8MR_C&G@TV,J\J9136= 6R[PLKUSI%<+9_9T+1-GIPLXU
P,AL#O#/N'0"UY&>?GFAT=->TJE+?V<FOB*A.M65'!FO8MGVJYWY!G.?%[$K24RE[
P5CHZZ9TDQBTD$MO$Y O'03*<@#"Z>97BW"8L#H[UIZ&2KNK"?T>"O<.F,$M6"]YW
PR).U@MR<5_Q>DL+WDLPT"!5BQP[N>95\TCNEAJU?1)G&-T+764?BLB]M"X80X21P
P6#-O"U>EVB3FQ,Z3VMAV5[ J(6X<2@]L<M<*ES-;KJQ"]LTM77[MT:;$W&;7<X+3
P,1V'&R>@3WQ1JL.89]L20D_]7YWGKDO@O'KYO^T"G"ZFH=_<^FET^2IG\L]"B)B[
PRFO+$AM@%3C6:^P$R_<RI*N\7UY& 2#+6L2>[D&VF1>_LK1B"205YU+N?2>P+A7 
P$^F#/3M/UX8,3C9\H8#!TJ$5QOQBRE$WD(T]UEMFO,=N)9J#EHW]/*=0(:ZYTQ1.
PE;PR*[[\].-F'%,"0<B_Z*H3ZR7R:6;OYXF(=@#%Q..Z'.IZT07@FZ_P8-65XS%V
P<J?@8>.T$U;O^0J6\\!L?^^_(GQ(^!36)X\NS](64J%/LV3G='FF0BZ;NG0GRJE9
P4.VZ+&G3?!>WI, @7MY]_OQ_HU'0@?9Q3.C,8#PV9K3EJ5-W^"?=H>B2_98B0#*A
P<!@5SP@$/6/CS]7'^^&2RE2P9[]@X"QX5</X^%5W)&N70.)"D5)2:$\E3]N!?)[E
P_:W)?[Y_5<9=B-)J0:*6^M^V(\#/6*JWSK.#QO+#7X%S-<PYL+'9FJ(;/D(GI<\@
P+7XM6YH:TY##>36A9D!::3F05E4SX<LS%L^%-=1SVV5: $!D]^=!4!PEN>Q]*"05
PDLY(7])2 G@JD'4\K2Q3E9<<TYL"C<\!%6G$6PT'3Y#IXC',(VZ-I:N::$T8S-&R
PAXSI;)O<X<0=%]3;G[B&GHM$O<<9>^EM46$B]Q5[F[_I1[TT1?W/) !HP+4Z^[O,
PQ7D<8/PHP?*>JAS9PWS6*XP2FEW1P(IEQ&CUMIQ(,@4TDB #]H[CH3,1]7"&^CN@
PM,BZ\6H67R?)STUQC!=P).>W;"XBUG;O.R7G09)GGPJ@@T&/=/:N #L3_Z@,4<AO
PEZHS4AK*96>SCQE;K!SB @KXLBY<;5MAZ>U_6BL,D"&Z)S&%LBF^*O,RE&PK?W_A
P?0:!P^1W>(F>-K8[A'[89&INL$T.@H3'42XC=EX:50D59?''L]Y@7,4"T]&QU%FE
P?YVB&L-X+&!]0FA(0D*F4'%,00QZ;2J=7V&+U1"OMI79FJ6U!#4>K1K_C5_WAB]9
P3 ))ST3?#PKIF-KT,I3LUT]SF_S: 652(PI0K6VX'"Q\&(<,Z_7%996'T1$ZZT ?
PN/EU4?(<8!RV9D%90S=CC9=[&-B\I;6=]>RHH)N\%=B@'4]M6TH@';(W_K #;/<F
PJTKJP ]Q.GY)-^.[GBT?J'*XD-21PBZ-(095OKE^;8AEZ2R"-?@TU$L\O-G63Q(8
PGK03]OCQLU^BEQ,F+DS6JZ9?)YEK^CW^)?E$?00?X$ECV?39H(Z0<Z^R)RR)Y\_"
P^$ IZ.2S_K"S803.;A-W7K GD0_B#3,5V,@RE39 B".HJL(0!G0FZ*ANX+L$F0R#
P#RW&_$/M>PH=\JS^@D7+S^ZU0(2'V>-N*_&P8?MOO6;#_9S";LX%'&:SP"OM1UZW
PU)NB>4^@&M-%=@A,>.7/"K]$N7-RP=3;_"V'S7S6PJ]+XZ[Z8O <TY3PX0-,2EK_
P;RO@91V(<AG*:YBSB5'T.9 1NP$7DFV45)%HGIL*C-$A5<[:WMB;>&-682(4>CVT
P:%P6=NE32,K%/JV&;1XO<T6:\_D:D )"(899FS@#3[N88/6!--G1PG2TS]O9G?#%
PKZY=,4_[+I"4RO:A#R>H:)$@B=NC9 >F>O6C$;QG780(G!VO+H"6UGAL6+H?:H1$
P/ *W,<\2,=]?,1WINM86W1MNM+CZE6Z;X>;2W,:S39Y\#(V)M'V5]A2^^I$<^UBB
PYL@QP8HM%Y/,H%1RM%UY1CIAK+J&++_F7@^R9*CZ*LH &B:A(Z4'97A=F?#,FG4+
PE&3F/&5WBG=9'0]14G('/BRO0GZSL\V5GWX$UR=$PA+DC7 7F<PS):4)QC9=[BI9
PR+DM, GC6775WJ#E>O,#2G<&IS7E;/L4U'D9&RY$PR3]+J]P*V'$D8>+)EA%Q@KF
PZ\20@>M93RTD^FLT"/M@;0?UO#'!PP1!T559=*!,BI$]W=A D6/D\0<^/4,/AI6!
PR9=XRJ^ ]M*:_M\*1R>*//;N\7U),U(US8'+?6)=]?"QXUOY$EEN5>K'^B[Z&+*0
PT.O?BO;L6SWQ&THH5JK/"L @_J<4]-];EC'"/F)Q'OH=Z0&/QI4@X/>(U)3@>.1O
P0MZ<X]BUV*$MFB]R%7<>$8 %X__%@NS7P[Y6*:'"N'M(%9GKU'[(;9&H3WJC+#M%
PH:>9+(Y5&J8?"44C:KR,O4M!IPT>= $PK0TZ4JZ@6( [)^Q78(MA";KI[A)F$\-/
P1K^V2$ 'ZJ_<HYQ8M?-3*F 4Z.2\F"%K5>@&5C\WYVV'$,PN&,0(1S,3>.>6S.DF
P^(T1Y*"WOX6NR$,O";@CB1C97H+Z(G4E',N\N?,4^(KKZ?)PXN7#Q87VLCR'U6F+
P9\P K\>\JFEPR.?]KV)XLVGV=[CN)^"N(E I'KG3X5J=(^DE-NPDN%K.IBWL9?-2
PL*I?\NKV)!JL-'XK'U\217*>"3TT/ N<(P_PA*EV\*A8. $8I2)4BN<Y.[\;"2W.
PO+MPWZTO##>6%8S*AZ)9A:/)ZL2C3([=<341*?)GJ#//_GE8H^EJ5@2M_)1=@(W]
PV*S'=I5Q_8J7'20L2(< ]S61W1;S[9M&X-<])DT\\+:X'MO>@-@"G&C06"?1?F%3
P/;K7@L2,Q/M-=$;V6C]C4:VM!YA?5$U>W+36DI*5\52]+Z,Z%\JJ%W9YQ=*%%H^&
P0M//&FU[48[7N^OTZLPF]3'\[@WEZWQL;:PX69C;PD+P'MA-,UX;_?\5R@6OY;Q]
PNQ1'?F6(]^<C7(HV@N[(BT=43N7!KS0G937IND.JID)$A!^(P[Z$59*"1C$D*NHX
P5& 8K*MCY.LK\M(+8 >>TSF5,]?A"A X/LIG 2:NXY5II44&<+^(^N?[]I3$OOK#
PJU"SFO%/:[1T;__-KU<N3B0;NGA]_R'_@<7ASZ"KVP#H#QS2+WL]IRN;!B[.WFK)
P;&I'"$A-/>,GO5SW>/9@G6#'WK=G ,ZN\%VM93,MD-:'@8'"P.2F!/84GL!ACP,W
P;R4./G3G+ZDBQ+Z?JRRL]F9/NNN*GW_F%51&Y:&=5('T!>5KVN1U&!=!3G\8$R@\
PLPU*$%;-I\ OM];XL&3DZA^,:_VQ'E)P2&Y/>*%4M'Y I>CI,;KG\(?_6>JMEIP@
PC)=KPJ(YPF30_( +N*C:O<6TI$)Y#<:/S1>X1ZO'RVU12TWM\1Z],)I(<68&LBWC
P>G<WDV%>GE=CFL?2!M3'$(N( _6CHVM2O??QX M,S\'ZH.%0_FJ E"QFHZNX>2>@
P=UV%F]C6Q;5^UR#Y!(A51?'^PK5YY.EM?1 <=*&_P!V" 7[?5X0G>!?6&RIPAC#4
PFCGOZ[&?-954T5%:&@G&<.=N $:MNRX>"%S?!4'&Y6X(_7A0$KK5A!J*C^V$#6;J
P#\V4FGGX:Q8REUI=C$H;V.9*3H(;_^9\;. ]*CH\]^?%=X[>"T_^$HK\?0XW:&8%
P2Y[S,:^_Y=F[ (;53I+]PH\FQ=,K6*?XO:!Z(4#Y0#ZEG 30ZO9/->M0]JI?_>V:
PL</E'Q%>0+0O ]R^O=T;M9[64QY[#;PT-.X1C-X).K1D:8.A7[0 RW7,4KI5Y1U.
P;K'=0@ V</MT7TJ1T?TQ&.]1D76H1XHW(P,N-$6T8X"?8ZY1S%*647 R+"]XU%C4
PL@W'K?V?=A5^09[OMZJ%ZEW6R7_Q"V>#JL/QBZ%W[S.;'#H.K2VYN+A\/>$@^EK'
P<(3^=$)*\#)"E06HT@^PX?X2UGBL?[-2A8QBXG>'&_Z!G@<:DK*F#=N9<0"2V;FY
PO_61FCEJHSQ*P#M!QQ9-01@,6,[A7,/%-2=QO. X=P(@*0K+.-)^R90J5-C3)*XK
P>W*8ONU@&"\L 7NR?T2FM+SS9/_=JG'">D\^ZS4JO,9JT..I_M:<$7;@\]DM6H?L
P9M0T+;J\T,=W(8B%,W!B_,K\%NV.L Y)PF_T1#Z$2.WH'B.LTQMP_Q" 4"8W642A
P.F).HKC)AQ:DS357FQFK+)GL\U8N3:83;F)7HTPZ0)??ED4FVXBNZD6#5:-P!N[T
PWUJ8>V'\A GXWIV]-:%]_&^I/][)"E3$D:#Z@L"FVS;)K =":DO75&Z*CP_J)/I%
P4RK3Z-?SU\6;XS;NMPS)FC)%$4[)FWB<.2J$GMHTR&'!E3FD.W?-H UW0 ES%F$S
PP_8T^W]R1/,.R3_#*0K?LGR(Q,&&<]'$G 26ODM%!^)8H)9[;0213PO<H14'^/5M
P^3YM9!C=O,_RP[T!8'\HZ?;H S!!@FWIE)>T"M=KD*+H.3,@"XK2GDS*!:&%0%3S
PQ>_CPV+MF#=-?"3++4U@B,E]2XA2;TS<87K+J"H[I.]HFL:)U<?9M@'M 4_K>YN0
P2=[G) 508JDK)&+!T!$'<1?6OX"BQ:68Q>8GZETF?7M!BR[ VG.A\6CFWQ^1Q(T;
P;[=D/KS'8#P\OTV&[#*K42*OCW^NQ^PR%-V9]&,YF8IP\-;>7.B4I'@E6=H)*P:-
P9OF@S5;B1J%Q!H4O]M/ITHP;+QAX4VTM,ZY*S2L+$49,KO,9P85$O':>$QL,%XPI
PSPHA&YU61W>Y#L?_127&@F?A4:RVQ2RU]QY6ZR%.$4EFJE'0H^ZE45(")$0O"._!
P+W-,/N0*5->B19)92A1/UGA=\L'70^ 7:(\4%VV &X OI@QD\'MZM :3"W88IH_7
P27>MPR-VMY<C?]/K_&:9UW6DQ51H.4+[:8&VW2ARM**/DD-ITAX62J9#2G?9>XO7
P]GM<(_9J YP'W\RLYSY[92$T&>B>FPTO'=ZG>BD@E[($)<-_;O]4,8X@)-?H[,BW
POJI+"DC^:43Y40 <>^5P@<V''N>7HN]R0O4,^0;=Z2*N@Z5%Q[B=],IJ'C[+!LNB
P/TY >.9,=EN,K:V"K_QO\9#=+?$A;_\>8^Q?Z"K@]V3HU_>F_001)%% G)6EZ^K@
PC,7RRI1.0/6<MDFSA4:Q6)!=5OD+8O86D3Y\*^=*!/G UG$J76HYIB=P:3O&U/S?
P5A/+"MPT.=N$C Q&@H7J&-A=%S7@$.42F\EABKI'IPCB_?RSIC@U %^]U>:FN]%B
P,'C.1BC#2ZRDNINA!KA%;VBSWAG5#C;G8\ +=M0/V7"Z805B/7QU]1 ^FG-/*B"[
PHJ$MA;166Y?W73>+W@PXU!S*EG[P)Q,%@K[=U8<0*'9%0LM4 5[,Q\;O@O>"(\[<
P37!8[-51!#.:[,Q9F1362M;#C7)NDI%!.>3]QV3Y^HT4V?\&((D%1J@JW4W71 -X
P,,&THZ5&')8PLZQ7"!N,Y\KM:$?NJD/CV,<IE1O#A6F#$DG<JZ\QOE^$6R_@Q 8T
PROS^^B1 5JB7PR GY,%G79AEZ^P1S_B\-:'[KA? :&NSR) ZDOO,+H._D?RXR90Q
P"RS74S;(@,MH5ZA'\Z7++TW46.:QKJ$JKJ)H\>P)IM"V0$\EI&8U7J'3=*LD(^M]
P6OMLM=ES)A#ALD5/K^/YMJ/TP=^)HW1JL)@B232=8#44GH7=YN%^I:@/4:"/NX\7
P8F\SMQ%NO^N=(\8ZJ(A-8YY63N'M,>Q#[N?,=$_U 9[UXLBQW !(S9;,!_LH^?6Q
P9.*HRU"5_U["7@@#T"EKHA1-2&/_[%'-]G!EB[<A%K-4V(Q;LO0E$8LP$Y46',R!
PJ!YY/"J? ?Q>&E;NH2)%P";G8WLM(BJX2;#'8?:Q8=*/9:55: BF\=9LYB^VIHVV
P6GPD9OYJ'O:X/L 5L I6(MU-;<S)RLGE_=IHHF4SU)^ZVS7;W9?2<&V-20I2T?6\
P*2E< #:/$LHW^@M5K-CZ#<+-<' [JW/R-GXM9U3*8VV2:DJ[E'FEDO?.O5MQ\O:D
P'NWJ89M=.76PZ8;."O:984PP87CA-5[@OT^\,7CQ@MP,0J35UG)Y1;%+\SL6G)@K
P&&C:)>O%\6:U^/I?LOX:SSR*NX0F^_LG/6>*54-\+GI@=R\?>E6XA9D0+(_H:SYX
P#^'4S<0#:I)A9=X?9DS4Z4G3L%YG;)Z.KJ7IY4HHJYZ%@@'I_:'Y!>R)=]!'/[,-
PT J/%7.9.?U1]")O-,YN/L:\[M09?TR5&XJ7S;,_(:GM5#.A3#,^\/,AK90/>QNM
PW(S(QM%!V3TD]W+T6_%Q3WW[<)5@T593_G2M!8R<+PK^I(*@GO,W<?PB9_;QD\JZ
P4HB/:SCSO,.&^ZDA98+O%QA#.!:RX_2_N3[K5IN+CB@LR\NT<]O)'G$K39 &E$!>
P-#$$8/=H4:A!305H$;1V97(0#%C.4C<)ZX'D:VE!39K#50E'47AH>V3AN82,\8IN
P(0*O -74AGN@+E1P@Y\O2E9"6-6/6<;/9G"SW0I8TX[X@_B4=1YWR>Q,UR"AG!C-
PZZ+U&#EW[L'Z'].-\2+C6Y]7 #V7;)'1=N3O1CA&*84.O=I]5SR.L%*+('!RHZAM
P3.7@O%,&\N#UE,!,@?*79I!J/?"[(%4)D\R8U=;,A+ZQ-(I# E*1[<$O9HL J>[W
PQ'I3(&M[!".;BD"&5V>3%<;K B4ZXF!6&JGT+FK???+90>/G6-("MM&=J S,I\VQ
PGL2<R"H.1"<VQ;&L]<*?N@TSH;T-5+W&0 53(O>-X+C':U\($T9/1J"IN# *I48+
P"$PFV-H [V;-*CA=<,*D\P;+28;.AEFVU#JR7EN O8F2*N%F-?*+61I$S1;PRQDL
P\$:O1DA^U=N6+HN07[E?A4*LPW#_;XR!\V/4C Q\1O^C_U^QAZ9%J*.=4\[':> W
P)CE5@E\"C"O2:0LZ9$RPFZAN#6A=A$SC0/,#EI)'@YY*Z=G<\S)L*//2@8F=T@1K
P3VC#OBEP%M2B&);(F<\(W9T42^;'J!*IJJA$TN24FCM/0NGCL=HO^/B./ :M^%X%
PG8HU?Z-4DXMD_W?A_BT=WBO6I4T' =Q'4AR*26^#&_&*I51S< +KR;<E3$AJ3!0"
P46 (2%B>J?1*8[WO+-T+'_.Z*-9HOA[S/K3CT]@]+HJ(Z"*H#)A5SU3I0[4]YGJ&
PII97UU?B/H4^7,-F=Y@?]Y".-C">%<.:[HZM*7DN-$%K0%=*.7TEZ+#8KW(,<V;E
PJ?/0R.4*H*2TFM..NDO0M\",")5LL?QK].HW,_.Q%IZ$W^.1,'*0"#X&R%USO0VQ
P/D#]G1QQ<6-E[ /69$Q-AYD0V6^-UBLW>W;$67PBY>KGSZ;:DZ(T4_MM6WJ'V;P.
P_38E0+!,</$*-(XX9R-'7.%1X)@*V1N< 4;@@///$Z_\69).9LP8':W(X!A,:6VA
P[_TRJ2@&65%B=[$V\> K^VM#Y%\HC[_;%;%<#T*+2$R1^?>YM%0P*@/I_]O9%EP5
P^#H.OZ%5,%D2/ $^UD^<F#QSH^K!E TTLI3OD*8=]B\II<WA2&">+L^PQ1]MQ ?,
PH&^Y8HG$<8V_ B0V5)*ZZ&68[P# B3%!O?FI5 [&-7SRAK)>!\-<G.NX>4MYUL8\
P[/E2.T-.@E@9'+XP9@S%'P20U-[@<^2BN<^ (%U'/11VF*B7WA EM'IQP-DQRF-8
P8KEE\N#X5. D>R5U#_"B%LY7*]FFFY&#+.Y665 T CNBQ].)F[Y7W3XLQY@'SP4*
PLHC8;$WI%Q9&H74<#0A_[ "SYB%3B_Y9+4<#[(!&Y'N#)$!<4F@1)<]5KCA-KL6X
P%!YS^6;:T2A%,Z&HF]MZWATWM ,)X55#YYQM/!_HQ5"H@8\T)3N/6K@P/V/E%R0/
PD ^8YTNG *.)$&XOT;0BNT4<T%.M5"7WJC(V#$"K;TG)'I:Q*U:OM9.227[\W4'(
P7_OU +OZM.];[V(^0="7_$*N#?9B2">?0PTKL:JK! ,,0/+:Y%?/^2"3E^,+ZX9E
PJV4.MX_G$ "KV^^:<2XIR.+NX_K=CJV!X =^#,?,#R3?A:;@ZX%'9ZZ>(:.4E(D=
PM&^T*'P^9,B,<\RU,^GU9WWV#OK@QO8++2#F5$DM2AF1LE)X<T2=ZCS2\J2CYS*T
PACVX,6;QR4%CF$GANM$R'!3%7M8Q<UC76J]EJT+Y?+6UU!5S<AZ:7V!L] ?8MU#9
PTXDZ6:G"TO@0-QFRS0!#F;])3*T96A9Q="U'M0"V^"(=Y<K'1B-'/RU.?0!=OB\(
P7U;,4-A#!0,P+A!7I@U%Y)1GV);G33(_ #[]_R=3Q5S4:DYK;I2N"H$%A!072>H0
P8VDDF/V?S-*1OA+/'H1@LQ^KTZ6@"L?-A%G 6\5R561I,9O2W"EL@#[2P$[K/K@A
P'%9G>3Z:\3< A+4#V.E.^C>.Y?< B[[X\Y.@Q" _B0*7DG<XR)UW[C%9(31BW',F
PW/,N.#Z.J@Y?(JB,\[?GJ+?C=WJL\OJV3]AZP,Z?-J4&^9RE<DM<^O_%3I%WLQ 5
PB_=RQXPX4^3R&R09*]==M.9)BOU"1:6[A&VETG[,O!^"#N.L^\7A];6@!ZJ4(]%!
PF_.C/Y.J .(_?(97KR@9V 6$2\D*4UQOA?NWS;F=8U3,AFU[\JVAVM7Z39^H&(F;
PM".54W09J\DIV1CPQWZOZHHPRM,_<'Q&;L*)>6L@Z"7+]!*#M-I59AV_J;I52,=\
P\HU>U(_D </*2Z3V9"41_?)BB+/DS14/\IH#S\==U &X>N/UKALECAD:=.:VM_]E
P9$L[42E?_KY9DHAFU-&?.:>#2(3[T;?.M%9I^49B:!^6\%\RQUU%V",36KU+*(E'
P"-4=A*S>H[&J'ZETKI^!*RRCDUI&)[=KF=;N,^52T,ZV+U:-%1N8YDD27?HD0=6]
PJ'6;2"Z4)-'WU:'4NUCX,ILIY+2BJ:@(?0JY$=DT@-+EA&A!81)QI(ALOM*CP>=%
PB14.%2MV/@FVA%MP=L<:WB*1NU<13.\THFG\_5+[3#:<_>=+-=(^0V5[*G%KE\X.
P"CK>0Y[G1GVE-5=;D9X>&S_.GSMY=(JRZYU\QS6^R%"%I3'2O)_Y7"3W"?X&T<\#
P<!$!_>YNS2S##]273.D6B1';9VZZ K223B-^G\'P::PIZN><\:J=!L@(_PY8[U(.
PR+3,O;:RSCC9 [<"=DN_3>973%IV5'+ O!$,O;:TA8"^1$P+,=;A=_/EA?:%MMLJ
P/AE8Z7'1 +Z<) 2VI2:&[&QK7<T^(@&*]KX>B79"\@I1+H#^TDRTY^B?3J]/!0XX
PZ7(EY=EK1!\XH5=/JO;L?<'OY)&"QGD,LJ(_2#0S2I3( NM+W&FS9.P;E>C*OF.,
P8E@KAY\MYS+,Z$XR[>#N@60442QI.UL^N945AQ88$E=-?<5>%@B^QY\;UHHI'(:R
P$;I XH(VV'0,]7.1MS*Y%TT@V(=0==3:V>?$BSPP#D76_GO_16+Q;<F;_''7W)8+
PL?OD2I4Y7$!CL?)3PHU%U$.O('O!!9CF!5(*/8*"BV]QE'>BQ?QRGSERW2<<I1F6
PB\>X+9^-\N//WTZ?.3=*WZ0I:3O@BSU=LJ0V&^&V%:=1>9$YM+SQ4DP9A7B!5^('
P+*MA*^A0_X^ A*6]"""VR.Q""+/=G>3;K=4MB4=!SHEX;(%^8X3ZB@=PY,P&FEE]
PIP*VF'P]HG4O:N#+U^VO2I_SPH*9&'(%JS2;*3AA'*2N.([V/ V'D\1AA6791M"Y
P*H4MW[X$?DEM#-CKNWB(5O>V?-)9BO(?FTCZR2K!SDG_^6\6T0+?^4%AZ@35:5&0
P2F!Z,Q=3+560C8Q+]K?LXHNW;U.,UM%&$O- , L95@^9U6+BBNDQ<D9EQT+70A#S
PG;I?8.<U-#W:6!!0[,$&&IKT)=MW=C\@TEAN/NA/WZNG :87#8)J>?! /+!^L%$[
PBZR\MS%?*C/:]=OO5KVW8D^<&?=#9R\O3]E^$WGPD@ _SW<'H?M!75*QJA1;XGG,
PO Q7=CO$Z=QA/"U'EI)O]4_7-Q@IK4Y;&N',7K3Z\=NO,D3QYD;PJN@PN)$2,9,K
P0K&'^Q+H$H]=_Y+2CUSK?JV.A@3\N/[TMB7QGALAY[5GMB+1A3+;PVZ!]5#MGXA/
P+3%,2CCU)'=70VIACA+L6)UI_H/0::]4148:*EPPANL4@TEWO[P1MR9;0.S*$S;>
P"&US'8->:EE>Y;NM)R]&B)S(.&6QG)DPQ!S<%WF:&>KE7NL#WB2!(E6P!.2L&BGQ
P%3TUS0G+@JYH\Z$U%]Q?X^$J";"#K&#1>T>P 0>SHDFT5Y<<Y8.$ETJ;^6._-#1U
P#V518)$ILKB,:?1UB:33=]X>8H6*5Z:D?@Y3]CN(S<0LF/LO]>#S<3D,/&)=OB6_
PK1)9@C!65.8TT!G;/R\(GY.=A*]=RA,#"XX(&$-Y" ZJL/MGFS\#S1IA7ZUL2L#'
PIPD,?TV"#=*>=@G"*43E"R]B03EG50BX35N06<6%T%9-*963)@H0Z,^[O'WX&[]A
P;919H1W+Y<2?"B!RFLD(O#+P_XVYT[@&%CS1")2(;C^T70#.NF+.Z!@)34R1P%5F
P!?EH-U*K(>'1=*37&5DB=Z'_!..#O;S!<U!UC2MA>4<^J"WQQ.;DLC$O=XLDH<>1
PE8]*CJW(-ZB7KBG:N>&X),RB#/7+^6^2+GSP82= 7DE/&.)X33T0-/IZ)1+#-8C'
PNA,$Q"H$B\BBJJWO\4:]&1-(RTD1G)JDQ;5#,2\32J0/LZ347$[;AC,=13Z$M69*
P$>*(;(R+U[V)IU7T2 60"?X+. <WY(MU@@ZZ(1K>K*>]Y[4N"<!2!9@8.69BC0ZC
P))*@'R[[OK^V]GQ"DA]=8!V3'^:47ZWP(#?E)EEC<CJ(9Z5U'$=&-[O(V_A<(_?E
PC3:AGT?&6O2W"[< Z!M[9*>17W>Q'JM==&@:DG$&NJ<*M:V+EQ[ +#JP@:O[I,X]
PA@PD57-KIRFO-X^5QP8_PL$1N*^<>8-]WR8,T%#T+C=, ]FF($/B;7$D+.D;X,'G
PL'5 1\7-P)!%JJKPA?4JS8*)AAKZFZ$IAS1J8&M'YL4,JA@]LELT2]G(O.G^$9BG
P-"4'%L8PLNT9%R!"1@,X601_"T2\_1@^S-%Z3HKV;"<E;@3^[*J$W!G7ZY6I/X<<
P5C6-)[;R_'VK/D)O0C$=%H0_\)J@-^$.Q/+ZFYN#]X7SX@F<]E1:UTQC[P]YG@B3
PH?)\'V[CLR0'&/@]Y*ZF)>[Q4#ZZAM@^1SPUZ%+7U17DH#KT9S2V*PT='^HQ(ULI
P3PF$0CHI@@$2([@TWB)%<6!7F"":7V9OY_@*@K#ZD-:D\50?E>5.>C]#JWEUC6U*
P(E,9X*M_H4P'_Z "O'[J, 6WE=B DGZNC4*MHHS')U!ENT/]\O5[,K<FU+7!(F1[
P'>^*RFW#]67[^#,VQEXS$DV,5BEFQ?AGDG^872W+4USH@TGH*Z(0JR\M\*/&0)X&
PE>J-(\$+@9_R]%3V#:7=IO>9CF4!KXU,IZA 3O5M!=_)H]0GA1?"80UFQ8K T\_5
P_]JLH%S2;W,W,G7A9QKXZHHCYZ"[._Q (&KBR\TA+K6\A0>[_9P;D&#A44X07/N4
PBW^:LTPX_TU74TG_3= '(ZPCU*H#E53")-"O^5R2.J0@I H#\R47%"NU?@'9NN*G
PX9BS,VQ[X4F9O[6(ZKV.:!>JV;&#,Z9!"X!7V.;F8-,0"?G/PD*:\OLME%3-4NCI
PB0$=L2V=6G0D?.YM&I2.)&8\]S(##9"0JG$O= ?$)W.L_1 )T.M]Q=DX DRR,@TI
P,&4F,?6UKWP?J%_=NNOGSK77J;%LX'HJG;S[4M=%DN3IH'ZC/B> +%IF*C@H1/K?
P"IC+X_QD#713D H9-/$8ZN(SZ[$=:+8%>Q09Z^6H:#B2//G]8-KO81+>83ZK=Z.S
PI Z&UL;>B%!_0^I?3+ H68,0G!J@95\S,WEPZG>4/Q;198)XX/&Y6<. D! T"CMB
PT?WI]$-PP^KZV2>[^G"WP)J]9@^9<]R*6OF_ ? :FX([M$IV+;NF*QL0PY_96N)C
PSMXF1K>?&PRBB$]Y(I%<GSYI7N@'X^NR@%FL?=9Z]PUA5^BX1R!,F3XG*6Z5>Z5P
P[ N?H\O_:BWZ',75X3H*4W_S),XQC["Q 51.!\HK7\A_UH- 0#@$N#';/S/J^*3J
P]C;L))L]SBKNH&[>-7Q!\B[T<:J4>Q*JM\)+0H?N:Q,W-,%:JO3I6GP&X-V\[/<N
P1#%IJKS&WWL,M +=@:LA:.;/OJ+?G&-2S(>6+W,T@0VMY4I?GS\CP*N@$-);OWVD
PD3V*S92=DIB_'YLZR@[3'4%,_YNDV(&DX.6<F&8R%N$G9%ETYJPTJJZ2:;TK6-LM
P5.Q.50M2A[02$NP!PGH5GY+ ZKK,*U5"2O8QPJI]U_,8X<^HG4W]Y3IL"+8'1E:\
P0CKC4@3\2_:V"Y;,Y5*M+!B&<]-O8GSVH 8R!P@5,WT-1W!Q^0J]9'4L5QMDU6I+
P#CFS %O\ O"!6AN)5SQM_; 0=4Z#<DBM3,Y=,&18A:@_%605OEFIFIP>5AH78.JX
PW,R]#YNMMUO543Q758;E36QL:*.-GK"M%!#<G!>V>KQM*,\?FRW>_S7(&?L &VF\
P->L8MH/%9777+F-7D)L;O<$\;V<G"2B$C?/"BR,=MXGLU 6":#^,K&FV'E@5!>00
P_.Y(L43 8Z!P'@)QRN>EX)M8$[2?W2D^A,2ZO1%FC&=>.,GB"S*G@ONG)5C!9HOP
P:46D!IP6CC>B7X32$9O\*6VHT=J2*9BH!S^I*I2-L0#,<P1"LCCM6P(9*N_G*\*.
PZ?@_A!C[_!:(@(NUZCBGDE?QDI?KX@>V_DKD\2X!C> 240&Z*FW82N#HRG&W9<^4
PUQL5W#RSR!N(YO?-M%0<Z\FLQ/81DX;&XE3*J\9]'O>/S1I(5@9L6]V*W;%$XT($
PFO;+-UYTCIMC#^45B-=$R;F#N5[1"\:FET],1LT+B2)D.]ZQ6#C4*[:/^.K.!+,]
PZ285VXR9B6PA>WXF:<\30FY"(,I#Z:%[6[H**;/B[:@4,/F3^0[*" @9J*@(5YV[
P;N@KSB.<>:B<]T[L,5S/>Q+0/(/D+3CI2V'_:-9>NC5IX&BBUI&UOS /<]5=3_G!
P+=@P_QD0-0A_'HYM".2Y6OK5U.I/_;#*<7S56LY7#/DFX3X$;+!WP!/)7WS7(MS(
P;9(GRJZKP,]>F'#L<@FH!+PBW:-+SS(@-DVI1CU@-#T;610G5E$4N>SYC=F'&-/3
P<'PT7(Z<^T\_TDRX\-)$2.+17SWTZ3< 6=9Z<,N7ZKK[&(2I%1$>":@4YG 6AR+J
P-P#R2#'D<3C%:[CS>]4:5=E8@CM9A XO6PAX&5%#2T]H!&R88V!/>WT%U1JM.M3C
PKDV&G2UB#P>4N;\S3#6OYX'$US/[[AMW1DD!!;92X-8>%E#L9A)@8%&J_8$!C5V+
PP]_.AD.YY4SJ%59),7O[,&23H=KE#2A35,I$=_8>(XU(&!N[=V5W)Q0H2??P)AWR
PV2O3>;WKJDQ00ND4O^+,&E(9>:(-MEV>V,04]JZ33\]=I83_/S/Z'.HFLSXB4N-?
PKX_Z9 ZE=@HY\*,V 6->&^UC\C1/A%-22XZ@X#Q-^5'UB-]TD&_''N1?36@)3ICG
PX+'YM1(.K-IG0;W7$(<&>]V3!\,-'$8$ ]M'7@'2C!'EM']^R+HLOLXM0P^X@-6Q
P>B.H@H,4_D+,CC+.ZIFK@!>R% @MP(+E@'/:#KA*OP%#0HU1M34$GL>@1(*>O=66
P,2S1T_DLCH!.O+++1^S^S-ZJR5<F7@"(@V"='F3-N[L),AT]L-><SI.&/.;^1<<!
PS7'C;\'O!(+:?H<'0VGHY?6N2N*I4!]5YAV>-5^[SL; D[.!UU>QEW,[W+1L(2>G
PULBCN(2C;@2>@/SU@C $58PGL\+T(P:KN*]H BCFHH5J50[XT63"#NKAGD9( _K8
PL#[\"I(7U>#_]\)K!7W\])T]W[5OCH7>%I6; D$)7M2^_/+R3!!QQE[7EG%SBN:F
P25$6M"7,J5+X$;"S^0=%EX7*HI997OM\L_[E*<K93H,_O$=H^N4%-#)I]:^W,86J
PK'TJ0TOP@J-7X5KXS ]K--T)^"MV523#J;.;W)G[7!"=YP7'\8FW^B%.*6H?TOVX
PY&>5_0B-ZK<283*D"HX5W,R*R6(K6NZU5;'QA-WG*88YQG\"M>.B<>];^O0\!46,
P&!E<>T,%"(,:RAC9V/I5Y"W.?:3QC;3L:'9$EY]"91S"O$)=_ME0RQBG>1-2S> $
P^N*S_XH\\:3"<8>@),E%B*8\?[5B@)W8G>_4D=UW[B?/(>G>\6&A-[P;R'R9IN+D
P5Z6 A[9W1&DRF\D]05ZN-SOISR!-R:>2+BM9\F'%ZOHP<H!%UIN1B4]I].!N(H*V
P!LF/M3PL57 Z)Z&4W%*%,>I:_0-'G8;;7_#,PXAWO'57DG,=WOY6U6.2!XS2JL2;
P595(Z=7>0\1Y=>>C+F<EUU#6Z%=-#/F'21=BF ?IW7I^P[CDCBA[+ZT/VH2$.B!]
P*L $6/SVJ#=% XOG]VQ93I)^F;CAI$ZIGWYUGPD *47_]8C"Q;CBT"ID<3#FPC3;
PBP44QR') HE$^WQ8*3'W6]>"N\R!@A>TDVS-/$8U_S!%_V,'%VKW,CAG]VV@^,<)
P+L6KQ4FHJ<,I1 Y[*>;5"/)6OAB'GHP\8LC7]!8W)(CP;QHH9W.RU#]V*0 WT(9+
P(8G]^?[D_?95/,H-@L%6B-7;LAJDK!!;Z]01'<)X3KJ3R@!R4KA,,8P>,Q.J[O_N
P !?\5627Z[ _[K,Y1?S"$:[K!!@?$Q2TA&_*$18,[>E$>^@7,SN0?@,$IF*=#5Z>
PKA& :5;U L%*[^#CQP^,O5+[X/HDR;/T/VCY!_ECK6-+&^TH(=$?M"28;R&>=?1[
P%)(9R#L4=S6_(PX!4N/31!I[[LV(Y,&@96<K!5"W(+-R#7FZCC3/_+Z""Z)9U*#3
PIV5KVU28@=_,BT-8>OU#HBL7Q\V*4K8E%8$^RF"=;!A?-@*7#]9"IQ;3$XN00!,W
P6<S(WKU<C@QK:@#?O6P5C02#*3;+*1-FZCH/51R2W(4<8N"AY?BJ>H @0Q7"=H["
PW^@,JO4 [/!'$_O6@;J/LKW+W<8I4[!HN75RCMM#2R^N5=\C6Q313V.!9(NOXEH$
P)4;<C&5#N?>0MB-6.;U+U7S\BF.DD)_ 7W2>S ;+@ZUB"[7CQX>W*L]'?JN410?Z
P%UR0+VV= J9^JA141?!F0#TD_^H6_U04QB"#V+81]48!>Q4PB\BE2&U>ZI(K^KJR
P,#-_+H8LAA@$56A*G\D^#<1+\$, 5/%&M7TCM-,>),"WB8PT1@+EVR8N,KQZ97/S
P[Z:5@/PYN]H]F1NT]#"?%KI2/E[4?-C+XD!\!3&_"E(11UXD8[("8PJ41<--A$23
PF R<]+<7?QR+ :I7UCDFF;M6^U])"W;1O_S-@"?@Y6\)$ZRZ"-8>!X*QM[W,'" L
P2OC]?KH<U'8INZ_Y5\JXH\N_#,'Z"4(K5YE.5X!WKZ@!+,IW=C4M*K11 C);22A^
P?%<D>B@&E+(7LR@\+ RJ?)PJ0=KCL'Z)RA; =+7T'^V8$H-(B5H?Q@]#RLM4J,/J
P/8\YD$>MC:>3M]LLMY"_8!2<RF"S7?&L4K8B>Y_7F2!B[9 WI:.'7QH '[WS4V)'
P:R7L:<>.&P\G[%?V'\PUL: A8*?ZZA$T_)]2CX"1ABMV6Q0X>(L_FGO/(O0YSY,R
P:<[$U,#5OWP%C9)[J6NOZZ3H:+VA[-ULG*-L??JKHN$H/"PA$,]8+#H.2]U8 0WM
PZN5+XY#)"R4[PH*0YV(3RTHA9+0%E9PZ&/];1.MEB1%0=2^^42),=+W)<],0IAUT
P D=</65<!F3YKO1UFWK+NM9VB RB'OD9RX>'0A9A(-MC^*ZS*SF&8+;U.@B-J[_B
PP'C@S >7L;NS4TVD*I%<91$!#>* F9!IW9CK9%8ZAAU!T:[/2D9QW@(4T!'F-B%%
P829LN_0NR2'$S^G C,>B4GJ=:E;](5;X3\\^G+]?78ZDZ>*A[G;Y3X1K*H>I+G1J
P8LIDG<N?0R_:.>$G(0.6UP0Z+]@T3O8"L[T 60P(";<T=N#HHTBA1"C@)0V@ZOG'
P!SI^IP;-2(88R3@D>%UWI'/:5:>!MLI9[UP6&B.2F*%MJQ_=]M6/^IHPW>Y8M#7@
P5V0P6GA9<D48"'G.6,_.*Z$:N"KZYBQ:2P80Z87 S#'HHNX^0NDWA%V#W=#/9 WZ
P $>[<+YN#[V1NFO/7D<Q\.58H5#^[&^0\[C'J(67:UV-STE(5T]ZTX+X7)9-8WU"
P=.27894\_M)E,^D/0AJ.$C)'J,2O >#'.9^8!JZ]6Y_<8O:PR?8"!:'0M)><%LPU
P4TOHTYQ"2229])+%YS<NW)*RN\/IO3:C.$QR-V.;;<69AF:7]G"P$F1[6"2"5G?J
P--SN,"7;;4V$,9S+%I4$J;5?*O>ECJ#)3,0;,W#9IYNE:7_UIU-D@$-&(8>_4 (R
PXV[<\L?W$824&Z@Q4@Q?$0: X=?V,HYZ^[I=6RD2'--E?7]AH-S9!T]Z,ML84R57
P6"W;/7 (0LG.EX+4$B?[G^:65C^_OVM"0$H-<$TWM&X$GY4^L.&E"@J_8?:K8]QE
PRH6XG(/MGM1"8X0YUF#LC_1%N"EKRYF HK[ U((Q^4_/#(*3X^*7,_\4]7'>%DZ(
P_,1-$3L\I0\-@0$'WU/0ZDI:_L0^ Q'P^"84&0T%3**A$$E?(TDCNVF:>$FAE#QU
PI%<\?BC-=Q+'J8\K$5JAB5]+ZPS=QI;.JI.D-933!I?L!?2>'U7N=T 5EV+]G\\O
PWD9O9ST$;<,UVM5>&!_Q[HJI]?8EMFLKI(6Q$KPGN]!Z3"+M*\FBSV[=L7B@+$&K
PG5OE4KDJQ+5!:P-P !KH_=Z8[+8#(_,CON<B6Y$265'R&]\CEXRM2],V2'\Y_!S5
P)V^C%70:Y*V1QO67H0G]0-*B&2.X/#"7F( RA"X BA4-Z/@HOE5@*:/E',^3[V0'
PXY<)O[C*2B8Q*YV]\G\A"^8KL!B_WY4^[UE4[;C:2+[, ((=_8MV^O+F9\]6E25'
PY#RQ2[,#&.]A/'9W)M4WM=&DGLY3O7TUA5&3TR/XQFI(37N!L9L)"'X;4<!0KEFN
PUKU"S)>N44\A]8:>%&\7WG4$[(/VS*(R^4:RQJEV85\6L6=_02OKHXD\.@M[/Z^>
P/T D7JEI8E :YD>6T$1$?Q$6R[[\ ?1@.\.78+I;Q\=(P_,+N.XUV'O0-1D*B?U5
PW?D.++\M9+LKB"3TAW!9T#.&?$+ E$#R,^JV?X7XCU?*ZL10WIU!NNBM,>T.6PFF
PN4BU9EUX71]DTIR3S0A"5B4]B]6H*O4JVND.Q\FI"AI%Q)>L[@* 9/JL>*(W:*Y0
P1JT<M[>W(?K.H-[)/X^?H5QN!+A1Y?RFW@(H ,:@8@N*1MPIC_CQ]:^#*L=HSN_3
P)CY\FA]7J>#\3&_6:P<OOQI4RTI'A:.&1P,(8J61%24=,JTG7\[@7I?1TQTR*=S0
P8[COX0XD8QF[9S:4$GYB3AVZ ME9-: '?D6J=$F?!V7>*1:F)#\I%OM2>]:V+%<M
P'EY;U4\!N1D&R$)87(9R[BXB'-54JJJ3WZ28D UEAYUE%J<U78>7"1JI[U5310$]
P0R WO,3-$M:TASRXE#$"*GC?W' P(R"\>?ET5_\<&U#NCNQKS7V[I6&T:T@"1=A#
P;NTHH/VD"<2ET7;P,H[5'MBKU]]M =^/\7(M]S=!7IA +T&"*,E?\DPTSK&6@*H5
P9EJU4YNZH"^W"&YI2Q%N&#2?-I>J8(!)R9OK<OB*+<.B+G\AK 93-STD(ZB\KY4+
P>B'<"/D.B%N$?<F^8*#YK ;EI0I1XS$7W)"\-/ !Y$"T4^.,1] *Y+[3+(HLWE2R
PWA;0N0+M/&&-%+BU'3^WJ+[6V*_EY8KVD29"J^508(1,YQ[! M=)Q7-YHA2?BI4?
P,:+\=SA#EDI]XP>07=J04C99KLO"CC.C_I< 'H%X'V5^R\P9NP)FSO,7D<%%Y8V7
P^%PKR($6(82;[021L?#Q$X7TT3AX8Y*=9PK4;)4<\[S<&(ASA7^;T^1!43-X[LN%
P<[ER%T2F9% 2ZMXL'B@;:A425+1^LG?+;A!$]38L=*)LU;U#;*:(R8]'9A:=J1IL
P R':A$7N$D']*OIQJ[_SR]TE5NC^@^L72QH16(%G@Y@T(]Q[8*D(5K&#/+AKW^$=
P#!#8]PEM!>6319J6TW=I]^Q8HW2L7Z9;[5(IJE]&?;$:..N9^+&LYE\P&1+-(\Z5
P$VO(\8(&3D#M5^!NK$/AO%*-1KI?BCFV9-E&XO028S'=C\]V]$]_%1E3$'0G$^?;
PG_*O)O45%V\I0 2\J K>ZYY<3'65N&KE_GYA90R9"RGVN#K*E:G<QFWM3,JZI7#Z
PC;KUD[ZJHQ7<""\]#;!P& 56^)MW^=[I?JA 0Q+)VZ:#X]8!G?YL*I&E3.'+'79(
PB_M\4FS1:_"4;DL6 N-< A'#)!<8CPC+!X\:6N(/3X9Y5PUKF><@<="Z#) 7-*BZ
PKV@MI/N?"XNKE'YA"0GU?A:?66JTJJP&'>#7+UH&+:Z0*O_5&X(,&D:?URZ1/N=-
PF@;ZFHYYZ=2?[ZD7@$T\[<[C&\YVHE66)5*\RW9EXF_\V#2"@OP@3?:HWU.58$4*
P-J-/I=QUQN2]!9 'G0,1#1;<<%)^>RY/GO\)&UIX*U!S%$<O],'1@1+JA8 +9>J+
PL*-3_72"CHQF :M:D'6L]\.4CKK%*WG[%K]=0"G:_0!C!$Y6;2-!TM876\;_@YZZ
P6ZRL!&K0+8ED /A$I)J79)JILK5"REGYISA*.B&5EHR_[?)XD+UQN8UON+0MF%6_
P'BSH_E3.+7+'>=KQ8"#1WZQQZ=L-3D/V G5T-W",E8RD<B;TN\.?/@&3AHI)=^=7
PBEW6H5MJ8#BRPL]P%P.[%L>;"I '5*+WR0;AJG+K<_M9%D,(?#E\LGL?!0^;;_VZ
PNBFQ)1H->4E6N1$NZ9+PDGHQ.Y_Y/)75;GW]V>/F9!Y![U_<)H;TB/M79I[+@8)U
P%Z@&FM&:6P13ARJD3QO.HZI<\"<A? EJ!UOB!2U(@SQNY+.WT@6Z!NF!GP=1?BM7
P;&ZF'JC,8)+E.98X-),1*9-.<<I*ZK>UX*NVPWP%^@&*7>=LAPDRD@4<5.VE'>S/
PJUW=.=[,/QHTZNJIBS/=(ZDF1E+T ,7LI"1,/ :0EWOT&YC%E5'MO+_F=C3:I>Y^
P%#]W7<5M87V/]F%T^ Q/: L$H ;7T 9,/O5G073!V"W%X>II[ -'3A#ZU#PC'ATM
P>TYQ68$:O'T3-<<G[T9U$4I?;BBC@V!10/N2/FZ3$]^#&GX?6SRBI;]BB=/QP2[Y
P!_68^''KJ0!J?[]@4N>MEXL/B7#B+!)C8ZB(.>\5*#[HY^%/_#P0<VV.!X2\Q3V+
PXL\TW,CIQ<DH&Y,W(19HSUG)OA2YFO?2L'&R!=1DV9?VEK_"NFH)G-(&G)L>2/?V
PJ<](,Q-OD%<ALU7&O&>9Q&)WVN;$[E3,]/G]\HT<?2+\*SN#A61Q=CW[.HM!UW.I
P>=KO:8XHWNBJ]#GRV\16Y#Z33MW34]BUM8*PG@@Y4W=4.4XW+I&;6W!BJ)Y+9H)E
P-;9\/&/=^?V>W1A6N[<8NG>DB\E#AH->'BKG07F]._53;%5MC"%6414V[?K^N6T4
P1'XWZ]M$";[KMY62YQ)7':'=E7SIN8&KEFIE]-1LJ9509E$.61UQ(O%M+-7!OL<R
PN'(FLJG0)['2Z/;1I?H?"*U!)Z-Y1=H&Y1M!*FF! E\<!O/Y@=6U6+A&J;!NCURE
P*NJ_F&=<!$U3((>^_KA)JZ&1N9AOP8Y:?:].O+$>-Q%2.&C6&ZXCCW8-3BX@E,&7
P"ZW5CS/2*-V*)\WHJ%&.^D%012P/BB'SX;BEEXR18C@9(LD;!&),ZFST-DN,&9P#
PY98"+9GK&;Y>X[SA=V\%2>"IM$G%$82@0U4R C-9DK!:0OIQ#R]P6O%NP^LI1.+$
PPE,:ZF@3KIG'K E^[IB":6C:L3Y/+3[DBXXO=T3!V6<(ES;K:[0.E4X*BKV]=W6R
PG$(F,2='0YC/?Q7_G:TQCIV$P'1^QB#ZCN564K.$P_RMS&/49_\0;\0OH%OXU$16
P//X(%-I-CW%+&>-B!I%$-+6[S%G> MH7$:4=G0!?8P4,=G2'HHCO ==ABR5A4.(=
PZ[<RN[K^F&9C1L\_>O#QP&# X[37FUAZJOQ9^J)EWF(_-03Y*I<AWU/:08"HPZ)/
PC$?@5_>@]PUV0@W]D)GCKE:N-,8P/NOD_5^2SV,OF$"KY@><@+07P=.)+V\Y.W-B
PM^Z:20G]0D)XM\HCW0Q*U,F_->DWU/:2FP4,6,Q:B>S(Z-,,.0LR,\2^[IL0C;:4
PD0HH9F0I\]#=D\\R;AEN$?N_>(<Y-;T<AVF:5\2G$'HJ*7>U==\/CF-$<=*-BUG8
P%)1XFX/O1=WY0RZ,%D5("('F4H$6$'JDJ&)H?FO4/KF6 (;2SU/,$OAY#O@&157&
P.P);[P@!7%Y&N@WE)*V75Y^? OD92_R,9MLG;E'N;H)4(P+PO=60=)>>CL4 L'EK
P@]I5$WE&=%0^DIWX<I=4&MTL3 .B20T""G/NYXS70X%B D2%"D7ZZ7W5K6O?ISNU
PE=HM(NSL<BX&W?C>1PP"@B/ULE@$\11GIO77MVA,:Z78@+.<E-?+8/LL/Q8!W=6>
P!-_Q4'W5UE;XG.1-Z;,XS@MMZ/P3LEP7_!:D+X*1:OZK(K+UZ3A2$V2#MS1.9+WE
PE6D0=NCP103$AI+'SFZ_;D#4D>@$-SLWRPB,5NTY8\DS1)%N*,\V:+YL&']C0EJ)
PSBK 0F58W\IGN)-8:&X<OQ]<-6/ KUX%2_'IG!14GP[:H3R:GES+47,0_+RV]2O4
P',+'J3*^LC2RW0Q;2O2S&8;E:CP3DV,S12X5B32U/6=AV/&0E^T=AB<E0 V0S%J\
P3KR:__&+P4VZ <$B(YPKW),':.]JL.B>KL+8Z)O/]^,W)^ 4SIH3GB#88! GVQ$B
P>H21P_F012I<H%0'24UEQA,5"1S.,DZ2=<3615JSI22MF]LVR)ULL;LI/@(T=HR]
PVA\J3JX'XHUXD0 #JAN,O3,39#LO]?XT'LV7]C,4PH %X&F5G5S+>:%%2C5_&#6U
P4*)2G;&W?@\[KRA0P?/Q)*%?!>*K':E[?E0="@]F"6_=W 9]C0#\V0/[:0 82U8N
PX7$WV.#,BSFS^LD]RA[ZWC<1U!4\(":723*,H-0IVH4;\X$KSP/KHMZOQ&>>-41,
PYR6.%R^ZAXY\,8'.['7OA9E<+ST5,;&4SZ<.M=/HK6;+Z1F,D4?&TA",94X-#,E)
P8R?9\_3]'\L]3U&$V+NVPW0LH?F.!'VS43Y-(9CID''R$F4ZZ?+X5?K60U21KG#_
PC:?R3@B]%0( =Y2BAU:76I^PQ=_[\XS^0\E^0*@$B6^0C0+XY-?JV9G05%CYG^!3
PV2*IXXM@#:6;3[G<F&2Q,S3DOY..+;UR],O, Y%*DXODG/#M>@M-%UGS=0P^4AW7
P_R+>_ S)\2H*.Z.C)\KX^XPA:W8!QUJB(DECB1Z(9CW7G[E68Z4.+#<9FN -+SZN
P]GZEB*FP6%!O@=GKLQ;!3:YC9HJW,[R_J"B0U.7KO'K>>R2WD%'"R5ITV;L283$\
P7FS^?//A('3U9R^GKC/?[1#YZUC2,*UC\G.!H[+5B9!IGVSKB,,$PB8P&T].#C)J
P_=/2*M+J;LLW'7_6D+G!D>AV":60YYKB$=<X\2/_H E*MLO_"' &G/PH__S-26FB
P6%L/%"\C):@9V?+:HF\LK_X%ND#CZ>O,@:HH0N&T&&TSK(^T\9"#%^3$ZHI(%,,@
PCNS]_(#I]0<&=0 !3#KVR"XN38/O#?1G[?\EE\783'NK5T\XX9 ]'ZU*JE#H+$[L
P(K/0PH>+VQ/Z#>D98,XE$1O707PLDW#^BXEZ4]3!1EI1=PE)]VBR<H=]-OW?<O)A
P()/>&TI=!'6#8&$V$KKY=6\YC-T,&RQC3LPV$0SVT=C WQ!E]/%K,3GOIGL+S*Y5
P/TRO.DOR&@R?VS9G,>^-A;:G+#TZ*(SZ=S(:KQSJ=@HTZ6GX5F6J'U,1!RDF91FZ
PU-QI%^4UV$:UT,&R[Q?;;'+%G5!:QRU%O74,A EG:/6,W0G<!G]37<+M!"%GN+JC
P7O%K;*[ZI:N<"OMZ8\L T@\&C5I!?VYJB5629JIRE?T2D2R]ZGC=TQ9T&P$;BWW2
PO#HHYT65<SM!(6;^H87\1R?R^7<.#5\KP;&17J\<)*^5VV=!C^ITO+$+6])Q(B S
P^+.9MIU:,MSK*$ =YAES.%B6.[VFTSSA=D4\>)T%:(8&N++M@;AW%B5:FW^UH)[]
P@DYX):7L&VY239+!<PT%7;6\$@Q49L"9D1_\ELM/9/^H'R22T"D65A1EZ,;90(G5
P(J;)Z[?8F5LG,\S2'MU+#Q*9/EEUL6\X0P<S94%*!$DEAU:7$C9.6B(!M6G+II6C
P&=CB'@4WS;00O!G'"T;',:3Q9)\6>/RJTQAF%FTVO"!S@I1X7K<Y"'ZOD%_)91R<
PBCAO_.;L%^7KNO+(Y:B05IR)OKK<R***0>*SR!U>X^B4)39O*%<X@D/UC)9VEL;>
PLK4#$(Z/:^JKFW7NAOSFA)A_FI1M"QKO[U_@V-J5HL=0_.ZY7IE3^#CCW79QL6%S
P,SOR(A3.*FY>PT!\<]7#/%<GR9X+VLIF^=U\ZMVJUW1O/KVTD8.%Y8%:>/F[<%M_
P*-B IU5P(AHG ,X]?71V1?EC'^G.Q\G?Q<;D(]3%<M25ZM$*A5R&VR!=]JKRJK<=
P V>3]3Z61,YD<&*0(#KEF7K),=6_<=I"2X!!?D)MYP[L5I1+\</8C>Y^U)<0Q5N!
P!.WQF(%R1_=G,K\P:,1*>P0FE'WNQJ/L: =1 .LQ!S';=VT7-Y([(0]5&Q6!C7UK
PP\DA4UP#,R,ZQHNU$QD&$6\354Z"MR1:S:[B.^V52<ZF&GI3DT,!CH$&5$N*^]YF
P65"\SG#"<T/MNP>*6_$?I%7 B,C4*919IE4?YHB#>-^4XL3,\RUE*T*6::4:\#-P
PCR-KWT/.1ZT2+&^-D81<(#Z+@\G?R/]2$RHQT+72W[$,IK*@9#U-.%A&%?B@"5)8
P=KQMTCKG!L^OYJ^Y%'-8A&*/!+">E\D.YP7<16+S66ZQ)<,F=X9S9JKY(Z$>'3(.
PZTWFK9?'8DA0FVKHC^TE=6Z$G]D E 1F:BM%0U5^6P]09OY[1V>#BH#]-[$L"P[&
PT,#'(D0=+HR.#Z<PJQ4L?R</DVM1Q?>H"M27<?&:/A.SA\,M8B]SE< GJD)1[&++
PJT9]3?:6!?].PF64CE.IQF.?I&UU@W'&%"S= 1PBIN;I]-V6:P-G?BR.*&TN+_!U
P@0C(?O3K#WA/A4.NWSB;3((*Z"?85W1_?P3O2(/?/RG(IPR@<@AEW"]0$14#/]GO
PH:9=\0H:/87Z[C2,1S3V4A[-J=RBZR:/N9!!C(WD:(#QN3!Q(OW6G\XQ47TH=MCE
P,V2 8!^T=Q@/7R#3PI#UKHH-IJU554%@)EA+0OF4<74?]3['/>Q$:&*XT[OK,P3O
P5=)9+Y>YC;_$$_-X0A];)OI/2J#:V[6D&JA:8_I=NXC6VA&&-$=BEJD12(Z*^ :O
PUOL,!5Q=;?N_UKU]3@(:<IQ_\PO&3 32RFR(J^B'2FE>O*)9>[([M3*P7*L3@=)W
P9;UKA+W&L8GIG,?K,IDM-\">.T10-1#G!):R02N;DBM@V%1:=OW"8)6-JT];L"";
P*,O;I>[^%FCMS5)*G#61 G.'S/:/->75)F'''$FUVKPGD?YOQ4=38R*OL'^-Z;.3
P:J U3C#98[^([##'J+4'@G(D$5V+#W/'4'^DD'+2S"IA$UP<5%O_XW7,M&ZPKZ*Z
P03$;M37?2 _OHX/_DSUY_?29E,D=,BJ%B,%90<B%ERBS@UMSB]8$)7*75KJ5DLX=
P-<*,+X 8B*JAWFV4,4?)>S)@&(,9UE^S1>Y&$RO/R6];S-(G[Y%A3DX5)$C&)N*D
P2K^M0Z)\C]S(5B^?>+BW#I?.V.3?VK32S;9*P@C]QZ0F$!4=!/;07T\1;13>[G#:
PH=D*9KG;(!];>41-:-;%LF0^*@=]-08TZ(RHVS@#V4GDHLG9W>I8[2),EYBX@?X7
P'F1:NQWX?6:'E] K5-NNWEZ4@O0/;9.N/L&._3YHX<Y?Y_LIB84-PGPZC 0D5IR%
PP7.,6/2H'DD78?Q01&[2W?.Q"JFB@72&C6355'*$S=7V&J)"9KZE!G?U#<G:%S4]
P.D)\RZ=K4QT_I)1[IUS^G:V&O 92 ,Q097;2)HT4!M.XL^""5"Z-]EV3XAD!\.]*
PJ# 9S <-2Q$E7EBKCZJ"JL.+) ^E"3_3_H+B+*()(VC4'9,'92(C ^8NYQ9TT+#O
P 48M^!EU<$X 2M3"IRI;&Y?.!RZMH>SV3L>%B?4KPQD"O1UR:)VJ:E ^, GX2!_/
P7@Z7T<#1M/PAPAZUQV2):ILQ"#_@5\C#CK1AR%)^)(LMY1[C9:_N]6D9976-RQ3V
PYXE;'0[8?^KZV<^ZV==*98M:GOL+#K3[0M#3U2B(1H!-GN, X^^C(WI1.MY@L'Z&
P\[YE4_>_#7RLZ._Q'N3KNB^2D>=N4RN^D+<B],*UJN)NGW6YC8-:0PO\0)Q$[4[!
P\7I$)F]438M7/+JOKOP+QTRW<%SB(B'015%(A2CGU>/(GG,^F^8*^WU'E'Q/< OQ
P 6A7:P<B1[XK< 8)YQ.7-HW;EJQB!2?_FF!-,HY+A? G)%<=9 XNR "G02HM!ZB0
P-OAZ05) 4_/4@$E0.T-(VT$G'RT/G_#7]Z&1B72 QP@UQ.K;:Y/CLW)@E857?N/I
P-R1YK@2@?C+5RLP!XFB5FU3*]P++-NWK(2CW5E4D- I9>..^I<\WO3Y2R9O'"$ND
PLY[^1PA%0!4J-71ZZV1H2U=>XZE$YZY>I+'\"B=(D!/@A<]NV>/GSR]6LS-2Q2F\
PHY](B4HB(P%[]=/%Z9F64T[J98"98!U)4<Q?T6FMQP[FV;!HQG6;4$*L=5E@ZU>2
PG8+BF4ZT,\>2 <N^JPO;P)F X9<XOLRJ2;'(L;,_[P$FF+S&M"&'0SPE ?&S$/3#
P2Y19P^MA&V5XMR<::Z:F=6T,NB+&";G$MM)F6%Y6#A_S2W!KDL]< G)]7J3CU@G7
P@GWIYPEI5J6Y/K#+Y#K3]R=<$/8BV^!1MWK7>EE%@4T=3>M1"[<-\IXU(9#\WR21
PVDU0>FV\16TCM_B$SV]=6#,*_1&B$UKXU8:-@3Y+)IPIL=1'\KE[=%#D@HAWS;?4
PL[R[1K+(U!\A241"E,<5Z/726TGUM'3;S/6>,Q"Q##\0'G>8//U,$.@9;DR/-S.Y
P7K9&8?//H7\47R&GGIK9)JU1S;^J^=X%H2K),%IW-)?)6>6X+?B6R!!,O&1Z'7A]
P9K6+,0F,K6]E['?!4>7'>J 77**72%A+60;CBS6U3KH/.DIMJ[G2!8)APKZP>#@H
PL@QBY84"OB^ NM$&?9+B5V?<U<^DH*Q%NBZ!*4$TW"AU"13>EOJ5B_ST$K.)+)A1
P&\T.2&P >##ULY9;=KGYA\OFX1.D=A-,8A(6@T(N8J;+";?V<_:_8A@\0STU90DE
P$PU)14A5JIZ"-KE[IX:6#J8?$*4#W)?%QB.+ZWBE\Y%C'D[[S-:99AI?L4+I3AWV
PX&2\_5QHG#&"C&0!',INZQ*Q#YY-E70P]Q&-SXC 4P=W. <Z^EIX/$LXE9MNS$L5
P3'D%F?NJ(W#;"@[-%T6ZO)Q+$%LJB@6T! NP2Q,%Q?[-Q"%!LXQF=LUUZ<&"0%OB
P:XB@/9+!4[3A4:A^$\:<C< S5EQM^3N=FBCQ=C%8H/5]Z;""L+_P#OB_BBM1$M?0
PS7\">#/^9W(,KZ9205AW6+J5HT8@+-OQ'=FI3]?#\V2MS)6W+-+,2ZHQP*_?P-I&
PCTH;L(.U]-&GY8U#_?!+T!" D&#-LZR!.50@#(5;??JLSYC5V\G!:9=;^2YGE(U!
P?%<X-P9""N6\$>D2160HR)E$P(;H"?> ?85_,Q>I2DCCJ@O-12'FH(A2:V1I-G44
P'&S:$9!.JF$EFSVM!'EM$4%DE6C:R.&7X"^V;GDJMDVF;6NA,]5PV]61JA(QAJXH
P;,3.UES0=DX]\1C%Q@PX$3UWOBN.DC-33C\'X'4W&QZFQ,L0$WA<G^LR>:RM$2.J
P!W'+9E^&W TD=%Z_6  3#X1G&RZ.AFF>0K+8F-S"ZVFB@')C"[ZA^ (W0;>;K)I]
P2@I/7R3!+XV +M)TF@=O3YG8/X+$V[/TC7YX+&82<JZVB\J)9D.Q6YDOG-E<,;Y(
P(NI6<63[A)CGRDU_9?3%LE7988 LDKU&VH8 D/>EY\N^81H4^+'75:3JG7"K9T-Q
PQ\@*.J#ZS^T>1]_!*F.DU<2JQ]KUBVY*L3+>RZ2+AJ$I3>WLWC\_"6HWZ;X<]4]J
PV'B\Y5%&B3'K;KQ"&.>FS<0XXO9OB&24QF*LQ2=8%<ADM5K.PY^::L^'>,@'B&)V
P-1)(3']EMGE]%6[\UT[)=<:"-:=:CU%6)2T>!=SH&G&G:%I.#N:U9-:GS<G4KN"S
PX#7!8,'+MD>NOJ5]_"=&X17QT,DTLV')3YJGRV&^,Q=@O-N+212L7+,ZGJ"($"]H
PCB)3_!8! %V3&I(^0G3N*U^;F*,!T_"EZ<ND( #MC9AD)JT0.DA^3W#Y/>YL G('
P/WW$(1AG/>D8=C1F[$K9=HAUQ2H-B>J7T-@?@_HB7XS%0%*V]MI0QXS43.-ZVR;K
PCJ28_1K+3YGB#KQ!SC4XBAOE=PU1;'MAML.M1,G@,"]646!:+A6!YFUTU&3 !7IB
P*32-JPK>U2=KU;@#.37TK53\,=2>$TK0*N7'4#M^IY]./HQL_UGI_D!Z7E2>.[QR
P,T.T7!3*!;,Q^0^>\4;5M/Y9#>+WH\XUIL6,Y-"UV'ZHH0K\4"H0.QX-"9X$MCL?
P:8]1VV5$>:RB3(=C*'@(OT(JL*<M^W"#?Z"74+C]A]RN%AYBUJQDI(A3'I1H AXD
P^"ZT <%EY=+$4;EMZ#O^6:>,: O1$JP-?,4LGSKA)-W7%$I/"D&;1;P'>LX&26]?
P[6_]_"'K]00ZH.<HJB*X6S,%*SMY(#OTV:=E=&E8V-PS[[RZ[+R ^'0\.,9*O/*Z
P'[8J NVH$-O>0K68I34%X<MXUM%#P]6/II_6('3UR@0LTO7 \7AG\CTE$J+.^FH\
P0P(M3%]3Z6.I,MA$T>S!@4&RCZK:YF@D$2TLHA %<"'QF,\U:SW#EPTJX_->^X, 
PY%I286,**Q!>/:)R#8FK3,]/RIY'%!#"HL5"Z7K=[)2QP@-)?L+60N",4$'V6C.X
PD]_HPG=!D U+.*P,WW(<[7S"DM*E/L36^55B(8-NG=CL B:OH%0<$JNF<\-$V267
P>C<'9Y4L]E@@,97B_ 0%^RFIT&ZQ)B$M-4/-S;/W' :EZ5'/N?[3:H15![3>9T"K
PF1ELK54DV76QM2BZ*%NC:M231)!B3_W1/@DEZ6OCJM _0,2RH>$,P7QCHL97CZ6O
P3&%TR!F\SN.RG0R+$ZK 8X'NO8ZHZ?T7=Q,-GJJ/!P%7\5!RQ$@2,-"9)^Y)O3G?
P>KSW,^>JBXO00=THYN-_"MOK"@KJ) /7FFB)B<#NT<C65>9M^&T62G5PPA(!W9Q:
PRC?+!(?)GJ&]( !TX.!)*'?+K6W^BXP'K]D]Q?0[#1V&>J(M3Q3 9/PC\CIO"F\B
P1ZG>ME9KA?@1)Z+=F8 #_3"IWG4%A.':_;!"SXRTG@&3\@=)BG7=4N)7B)U,N646
P:B_8X@7+<*.L(DK*CT7[DX-AV:TDG=8>G5IB8FDE0O6T/Z>_!QJX^,'.A$9.NWV"
P/56@L9667'2BW3T@EZ<@[Z'X=M6VW HA^*I1#<Z.>3GH^A7?,0-%,.'4R3W\VC?R
P^XTJR5;BO"F;$'7P,+$Z&/1_L6GSH+^) YOI7=,SB 7NI7WJ@-V6:I@:F8*(C2$K
PK EV'KG_1S;C/_MCZ_A<&J7@MGI+.H+2Y&!-*N(ONI4DP,IK3&\JWZM\M80IM#O_
PG$,P\?OF--AR+/34[U\7X/HP/>\7@,MJ? KNP<X5[^Z'6-SJL&.OX:/IG]EL):G'
P*F$B-8!#DR'.T*N;'+9ZT_=A:)K%JB, "T21RYSCAPB\%BL1GB7EG3\K=<W_VB'-
PO*(E[G-&6&!(0BM:;+Y1S#NT204'9X?7,J@7T]<Z!LVDU< >B]P,_VJ]9.7^1Y[[
P?-"/,AKR*@%O%WJPHGZ/+_!;\'W7KD+<?9:8ZL;%IF):Z%=+94QI[787Y(?B(<;J
P^E5<35Y6J-RI9G6%<0! @%BT$ ]WG-1,-_GDUXJF<.,8/^/0IORP9+:POZVP,[I>
P=)^[057@U4*ENI$%D_3P_ IW>"%]Y3Y@2*+QU8ED:@A+.9K37'OEW/ZD1CA*=+G;
P81=99L*27"5&^/.?1@H7)6)MC*F%:$Q!:1R(T1V(:0 4Q_?0&Q&:Q02"1GF>G!D0
P[T1E.81B3G T'SZ_C;EFH7.,\SRQ18$]DLG<A>$[/-5T8J?X#EY3BY"SC7&4.AW6
P%/Z[?M+W$G2+22H_A1B4VLWKV0^4Q'34B'/*KO'*[).$'CSA]9 A53)E)<'K2@0J
P"P01YP^$^GNY*%.P3GHW2V;5[G'(A 'FRGMC.)\*WN*!NUF<#"A>JS>7>V"^1 6 
PS4 Y-'B[7L ZU,#6RNSPW='4"2G(-TV@GL)WW@\@Y"-%AEZEU'$7[7K[,.\HH3F(
P'%X?;\[O1Y5QY)1?([SFBWL*WC>*[ONQGS"Q<+>1:-#Y('QT%5PZ'*'&F-KS# )]
PF9O[IS:0G3>X!Z8SZ_*NP1?:"1#.]_]3[Q!!5)PD$(;Q#/W#RUW-!EG!-EUT]D;E
P0,AH4S0N0A5F)!?;5!JS\F*?)\&YT@.F!#3H?5;F9I=95O1, [%$%1?3D+%#&[?A
P6>E]!Q(*!\UF2*2AJ^ BP6&'\8(%5X>7GQ[5JRO^_?GC6HM'@CYBYO8IZ>GB)9,=
P^/6'2;\FA'IK>:%+$4B3G_GW]]DM^G&?/SXD1KT,%?P[L'M?Y+=6/I.>BOA@#!;L
P?N%3S.O7OYM^8:IYY0F>$E$;:@123-*FB6![]=/.7DM^;+97/UA%(N\:B^HD;;0[
P0/UHBN6Z&_2O_J$'KS385U$/$%>^0#K:$=D6;8(I)V;"*#8T#[>*&<T$)98+AD$&
P3&NZB/A>NGZ.V>@D(#7AQ\(#W ^U_$6]KAT,R9ZLT8X]:7)9RKFWJ5V:3.<JHTSI
PX0E"'SW*UK4-MO/40I[#$DW83$^=)R1YJ#.6@YA;BL^RM;:6\(F-LK^?X6U2.BC7
P4 TR+"#M6E"E,Q[P.NR+\5-Q'OY! VFKUM3)^-/^XL'<I;3MV,Q*6R0871BF*OWJ
P^U"#"$@NGSY,G&'.R4E$B)2PY9)M!>93_[<:T1E;"I)E!#/ON>WV_C0CD9+X0\R^
PSI\T0"/B;Z+'$X#@[+D&",L/T/&Q38-TS1O%OCOK&B,63<, 5U7C_-V4H12GGZ%\
P<>#A#O!9RK5(HR#R4*"A"MTIW-X.S(*R<NZH&7\8!7["2QMH5!T3/N3'C273,-?>
P/ATIC$PMG2H#-5"7YY,[!TT2Z);)* U3E%'AVT4#U1]LETQUW'390"/><WW&W)T%
P)IWD-55@E""+KY*>F?EL$F(*MJ[:+W+[\ ZZVBY7CZ1$U_*0*5]204DI>^B:E _\
PGDE5GZW>P^<_-:SY:^)7%[M]^*EL]?8 ASIM5S7.._L&T%1A("0'B.R%OV.-]:S,
PIEV&VL:SX1MHSO#O97\.=A4NK<IT#\PD3'D<;0P<J5FP!)L+#,R%,^7I<":22P?+
PC]4Q>G@WF1!=60U5.1O%\4T:(,.RO53O_I*"_Q<Q(%8%TH%?^@0DO0TL<$R$G=:[
P)\TK@)_P95<<Y 4$ZV,)._V9X$]*D$09?NCG+P2JTT CL9V<WA-LB/$@FM*SM0*1
P;?%XQ24*3/\RIT&949WPA3>L%Y QT+-?A_BD!(3WHLNVJ(@TNP.,!6:A=F:DX1,:
PWBG72<E$:U",[JG[["_"$)8AWJ/(>9N)2O)2>5V4FH!K6B)"NUCV#=6F)=W<_PC(
P5E6?( H&Y_\.551%>%H)V5Q:^ -8^6Y-0)4*S8CG=Q[]K=0OU4)]IM)4W--&D>*E
PTT>6=A\K3V*Y^TL^ZE5/"92"&OX2N 15!9TI!#WCQ<+?.N6$5Q?+=:&A=$8%L>U0
P% &R4Z)/-7-$V1'1RP16K3"J7WH#4BP6$$;9"MM4T@NJ#R,;-E>8>*_/OY'QL8\9
P\;_/S-K:OIR5/&.0K=(W"[1V.,:=!SM.@,D.:,FLP?/1//^TW6O1JRT%Y-^JP3TZ
P7=E.EB.1'4^L1OISPQKA[W;,GO2\=#0C"HF1%PK!DKKN)7_4@^&>C=X8CCZC(NP-
P6^JU>R-++>>7G\X7N;]0=;F$S0%D\8-/*L,+_!4M=<PVOX4'00>ZY.^V)R]8H)Z^
PLOR*W-C\B*#AI @?B=?*U>'0V8YWB\;6_"PYO@^V(C&EJD[ A=J&]D)=,V"(RI5'
P:7;]4VBA'A*63-2BTFOY*.I7?[JDD6M8GQ%W^^PD>] /E-_ V7,H57JQ<^Y%+]4B
P)B0NCZ0QE9J$Y,E)<5D008)MT%:,?2GD&=.%8FZ.J\A[0FK)('@@%XK,H5K:BM8(
PU&85F.<= %_P%D(H__9&3A!="M6_"UF."&8AZ)DJN[1:1-*5UZ^LPNPPGF>^+J%3
P?4D]X'9";7,@-4T"KWZ43'9)=RIU1.:8+.Y0LF)W9\K51SXUJ8@N59ZHW,A8XV]V
P(T1/N&\O^..GZ^0B;]$\C%+0MYNF4+97<-]RI&W5K";.Y\$^-"'6=&TM*DC#.T=U
P<4]+@K2;^T9T,[0I8_"P>7[7#!-"03%;7/D!UI0 PW7('2(Z/()MYM#3_AA*$F+L
P!L]\VYR9C^Q2\!2Z\95I\U;9\."UEQ@!5JRP/]$>%5CF7JX 3V8/5!^HOK;Y=AX?
PW-, 7!7_B=)V#=DL3+ET9=KW +V'L$EYJZ"(G07N"#+Z9^T65&[L?C'YU#>Y/1IZ
P6FE6<OF:QGCAL2\-W%-@E =X",8]&]D +J(?\YB]#B6D3DK/_^F/ >9&1Z=TUBQ)
P/$5 U=208M,6N\6/I$,YO6O:SK/'[70+(16K_>,;D=33Y&>W"YZP)SN@+>YI"97A
P\7UU?GP4[K%@BYJ9&AI'YM4ZH>-8+*1LAWPZ9,G<9Q^D[&0;?L5&Q4Q/GIRDR4_.
PDU(\I,0!PU[NV_F(.V%B,+SNZX3[.&7]3-4W!E=/0_-Y-9W:V>"N@O?,8K@0S$%O
P&V!%'D;+H9&K?<5'0X];0;W373):!D:8/2K$\21BA<-R0KW3L7Z)<VR5U\05'-IS
P1#AI78%8UNLDMZ-C$3HXCGHI"^P^!5&,F=Q?9.KILNSK>NIR4*?0S%?!"22 <CBB
PR2:ZP^#94ES#H5UW,EYU(SI(5AN+L@%I:6A),Q-VQD#RX7NDOV4*3= *D]\ZOSA9
P*]N7@*GW^GD=BW^6E>_=7/6U][YO$7<9M\EX%TUTI/T@EI[)C.#UL,JK L&</GI5
PZ==FF0$]+I'.\<<LNPUS93AJ5R (EE%/ Y&Q=8/WXA;NP?XE9CR."BX#*-Q!Q)F2
P!*S\2;>XS,XYIZGP-$;,CMK'IX;_^-/Y2KSR.GH(3Q@4Z!YXNV2&W5_W,^;Y^?72
PTV]/PDOECZ9V<W&QXUT!P)WU0P-,D[/X_J-Q&9/ET.5VS]Q&6EHPB1KG9B;&<_-M
P>FJXS^IW3*@LV?L16&C5WPR@K+-NG^*WJ,8M%;N5'TJZ_V82NS2&FP=O@W0OL"F7
P^H<T;02QKW/FA<P]MEI8A#03E)O?[8#B%]3QI^M(D[PK]"DE'!W!"^3W?2DP+1")
P$\=G@\E.I8%Y");&H#2C$R$9L(L<PHA0*I?-*"_"+[SC7MX4RX%LHTI"VY;%6H&C
P2VQ2ZR]@)Y+RIAYV4<E@#&N*3A?#< \*S&3ZPEN8I5#_9TB\[H_-X2A]/M1".+DD
P/T9" GJG/V3DFRP2XD<M](^\M/U[T$)GS+L.\7Q'+7Y\.$L9%$-Z>9'P4?=+X'K<
P[;#/L71R5O'R"M@:I&CN07##BA#0DC;<&E609#V^ZTK\+=O^=KD9&&/ZC*@F+60%
P_%-WXI9^>]L1,OXL\VA2-PH/E&:$$E8B.BGI0%EK. &V/UUG_N#IKO X4^P=6T$=
PN(@6*8"F"XG;48MWA59SRQ8QS<7%P;3(S3@;(=CO7VN^//6+^__A C7.+RI:PD!M
PYHXT(ZKT-6Q#._B >&M&!/W0B +NH=\7@?=)V$L@9"W'I=,-;AP![)5WM=S!$V$<
P&.:2Z*3Y*%RAAG)_70IEJ]MLK28GB<DE=5F56S]^KR)=K.:I#[X%3TK\CN>['[(;
PQ*<Y)A <.AZOC7_*G,']6Z]8V&S(;0_&/?\-'&M9ZQ(OT<R5Z8R&#6?)8L7["_F;
P%2=1)F(QQOK<><9-G#@R)V^%;TUEF/U%LM@EPC3P7T9]"#Z34@[OT<:GRMX2<@.F
P.(O:EP''@<S9OEU*!1TO_,E]R,-,.U1@FO19"R*7Z3,IM6O?A2)>1ZZHI4?Q_&SH
P>&[D<E".'>?C4^ Q>Y2 0-LDV8C&:%D3W9L0($@5,0A_UEC'D&"L9:JT9?FM_DJ]
P7WCAS#80H'PS?[T_$QORPI/T!/AP@S0K/D!#'/JM$L:%6ZMYTL;H+DIP,VR7JH"Q
P=925K.#;Q:Y]^:F L=]'9=U.=T)8<0@B%K3N?R>NP30)*\B%X2*\':$Z%$8,5:C;
P":/6C)9Q5J;9>.TD'8_OE/,DOW1_]ZD?T'B(CCW.%]OW7O2FT7]1I[BN+M0T4CQ(
PYPNF!EHP5"9@<,QM&\%'O$S2?#*@0=]%F2>D]/) 5#VI*X6':#JS8"QG;[6W-G.U
P/\%B"3Q?>HI; UUF@D$J6&/@K)]R>CJ2B'-__U.4Z"6NP\82-3QZ<2BAW2F&*O#O
P1M0RAL&N\^2"Y\L(/OAID6<SUE%"+!";6;R0.WBI[Y$I+.]ZF;C3N*,5_1H<C1O_
PT2-6T;%ZV8_&ZK3GZJ/+F1][)<&K8JO4J @8IT3G/Z9[N6(,M@B52!Z6H?6_O!'1
PHP*9\$#<641- 1$X!.?NB?:!.J7,FTS4>*4 6 A,-\*0%8EKV]9\(GF&GY,6VJ+L
P]SHKERCW+/1+(MERC!)3>3UXQ6%UPRR/R[9C*AQK'+BT#GT%JRVPW\F1DR+1FU9V
PSNI. H$>4%G6FEZS[B;D(W0@5\5C5Q=J-17L4I@!FWYF-/Q]G$H$'\]5F#%KF7K?
P5K7*ED6D\<=_)5VI3M)J@[15(UN;ORWB"4'[U=F.EW'"5L9XP9!6>^['LB-?(C$#
P"I4J&RDYUC[19K6]"F=PKMI54[EZR!A5A;RK9%K7IJJDXE3OTX S3O!LA7/+IU-Y
P1!7*R9@_Q(E[.-IQ0:?GV+\APU9G!EJ>PR^W+U!2#</B.FYB"PB]496,:VGDW7\?
P1P35=>*-R/-[*_30-(BFS];[C/52NQ3P46]/'G>4LF,_>.TXZ D^ACTD05B)VLRT
P')D^56P(LNL^+?M+_$<QJ[._E*QUC$&^A3BOKAL5*E06CI].<SB:9 \'H6E+!W@_
P08IF2#]NLT [>_ULD!=SL400W@4%+J1 ]K@#\@H!U1E[EHXY$(YRYNGAJ]S114S'
P!9QKL))_7,_B^_C=O/3JYL!&Y>D(_ 4!A+8;BQ7TZ@$$A]J+LND<(8M0MN\@L(I\
P&VUO\8>_EI$+O5D&]P.4+2.RN*/3DR3\05F9KL!%R IHB/GW"RCY25(%_=>6$O<1
PA)FQHXW/L0!/90UN43I?Q!742.DR\XPZJ8Y+DHYNX40L'+K5'9 <:;I6$3J;-T)>
PY^S ,($Q"M=R'K XNTZ_QO3[!RZNN1DQVQKC,K:0,"S$5 6+1SSA%>3Z2?(M5UF,
P7J["K"&)$\4[X<QTH0')N03B'2ZN9TC+UR<\IU;DU],:*V)Z(,Z'(/SSC--^/>\@
P7')/3SJRZ6N?KFJ8AC_H+S:9@QTC$_YX&HPTZGUY4O*\Q&=-8060HDW-F-8^/20D
PK+%.W%-C74L)>!&Z'>&D<_';$3LN.ORJ4]"J0]9=/SS\V]]!NE^" [Y<V/-2TL&+
PNP(,H3/M,4+)T\QJ'C!#UZFEM<W=S35]6OV#Y''ECXE3C+$T6* C.8MI D66[L/?
P9!\XGL(FM4>'EDXL5>[%7')0:>HH9O>07U<'XSE,2Y;5\!MO]V,QF"N2$XS?@9A^
PLL+L="7('&P-QLM]>Y&IFPG&=1C_WX>$'W8_4J5 D='"[@L&;6W=KR=+ W. U%0"
P^*,33,7=)\'!'<]V.2!QT!H9FW)E9L=*647>OD+F!P^8TW3E,OL=WA&-&W<'F_%V
PO#I$5&^BEYN*RVJ<!,.WN$M^CK)R4=TP/J/4CH%_BUJ&S 5U^IHW@UP8]..7#]; 
P%;VR2X5AI[7<:X8AM+K4X'#M//'BY\)H3*D=8.0+756-5[S5,''%=1%TG[@?D+GQ
P 8.>@EIDMS;8O%YR;P;]-##\WJ'_ZV$4\T\,(8HV@Q=/&'<#+B>=AA7M[ S"<J91
P^-EZLJIBOXU%EF-9TZPD)<)\"A$G.2O+$4</O+H&7"KR3FP:#@5:XS#Y%\GIHG(H
PR0F+[C4B&[ _<J_.B-Y]QMD9PC2;9VCL[ZCF^94@%V=B%T81"^^KJ>V'3(^!KSND
PP&L6IF5GQ&JTQ$-LY;*%M7H"GUFIVQO0Q3%=)=W/!58;Y0K/Q8$G.7J;"ZM!AV%?
P"CZP\8-]W+/,YWFMARV"](\MM@V[CEW,?H#92*]M\?/'448[QV0SZQ70"YTP9C',
PC,RCY!I$2J&!"+;K2J/Q,(%8U;J@J +!T>!:1?1YZ;0/>7MV23^_S<0\IW%7G :M
P\TP.U/[D79/Y*!-R!@!R:1(PPQ[YC6,M1Y* _/KS^)8?)^LT_Q(UB9>&*>U[4\C7
PB+R6]\:"EJ.)N??='D/2MP_71I<))@,>_IC?W1Z+K1<J#0&ETFO1& ;\&QUP(GLI
PF03,P3_&I,PPWF+NL%HRM.^[PJ]VE>+8\G6NGGKC/D7[ U</SY(!#=>"A526]A%V
PSADSP-!+-^%#JJ9%"5^S[VL=NMFP MTDU : 0,F[V<T+/L6XQ5S8H$5<)/NB#CT<
PP1?$H<QJJ^IR%YZX2#R*WZC.G[9DF95;[,(DJZ@*S\SP7K.$'A_Q5-@,>JA<&GP:
PU;'S$4%.X"LJABVPEX567$O!H$&]AF[?)V.N1\#R=,'=!Z&'$I6MC'$Y(WQ6]+L?
PR:00_;)%^>(U'-SGE9R#22"2_#'?5?'XLB,?PT+#E<F_RP]3LM#YN047]YG^7''J
PNHF&DR,%N08/;-G7+MP(,'_ V<[K4^N+0P=^QLQQU,U!UBLR'VL^RW[D"16I$\+&
PC$;N?6,=GA.\HGEUV^\U-%0].2PR"O6;V]T'2LR1R;1BZI# '>'JIO""?@34V5!Y
P9E5$J01:?=L+V'45DYQ6X,(9ES/C!Y111R0Q!T<!<J(AQ]X()*:<E2Y^&$$'MO5V
PN=2=QPZJ7H7#:FD\ P?"?:96/^AV1ZWU:_'G&!%_A= 3CRF@?VGO<HO/A?C(U63O
P[-2,_XQH9EA!,%?,VG\G=3-%!>&87OP_'S+/4,XS7&4MEK'H2)M\&QBI56#(=? A
PD:M4XU_EF<:_I!2B=1O;98IZEH2EB/:Y***+I PI3%M^/7)#!]RZ; K*RO@_/#A\
P/,KQM<)-!9>*@<!&'_]F>F4;FWDGG0#\B>H3K<48<=2=79]]+6L91,*"XACIN-6[
PT^>)%88^R)Z/7ZR$'(7"UP\$AX,(2LW6R\9<@Z)H2EH+R06\^'SF-ESWS('0YJ/4
P%0?ZOIO5P'_>:]LB09PM%!./;TRE_B"1*\%R^T!>%C:1#H,@MIJ1H;*67LTM]K;C
P:W]61B=/?L3?H$/61;)(\RH_;BSHV5O4WQY$ H8!F2.141W$.-E!6&D%&+$K7KB_
PS,HH,U.%<QA)YG!++5M,NKV:H^$&.-5,_U+;\FLKI2HV.P7./.Q8?+#M= P^U?:O
PH,YOX^ZVT$*Q)N #M+'3ER8]B,S/&IF,I*16-#^8JH)L]$M4HS K)I 4"9YP9 I>
P/WAGWF=55'US64VBR?/1 '"L Q0XP:F_SLVP0N7=J+:8(;\:A*+]68(&Q9ZQ&5CI
PMJ&?%7S]CIBTS;>,;1D/67+SS 6($$(\ BT1<H8[?XM6=:,M,^/+DZ>SMR+8UJK*
P<9Q5 U^R+/+^]PHI"5[GWHC5@_L!+ECL^0NBLX-E7]0U-_74T>((6@=PW)=O>.<X
P*6O,DP@5I8?L_5@(4HD0[4\80@8!S?"?)XX:-!?&/KZ0@YBZS$0K<\6K!E8%HI(+
PM)Y/NE;_PN *7JH(1HEE"U^"EDH')1;\_.)[Z.D4618)J6\Z QC+UK_BB0JC$)J7
P^?-P"E@*/%Q*$9=[JWX'H^U:JFN&DT;GSERP%8E$UUOT3!3;F_+^-!:V:EFT NN_
P+$=1'3=/:CG3X2@&7B .SZ[%S@9\:3&50')U-''+4V'!A/M<5!%L4F\#M@5E7T6X
P(,=1\J%QJ\<N[=\5SULR@9,65J.E4IH3W4\2AYB'GQBR*83;@G=_W9=))O=N>K\V
PB@-UU8=HD2.VSE77->JI/3Z[!&$Y! [XZ>*F8SHM.K<VI*OKH8YV<W:JBM#SH$[C
P #"FVY2#JP=#'_]#=IW2?G,N] I,A?>F[P7TS![=Z[TT"F=P'EZM?2=521S3X'QZ
PA*QZ2]B0'[_-Y4-&@,=5H%M^'VUN@V>S0('SX_46]R*C9+!FW34KM! /@J+OC,W)
PG(8%C;K()!%$^;>-.7N]W %JZJ*KLI%ON>OXFYG?'J5[G D_V>UQBE& AE[$2=S0
P;]SL85ANW"Y)8U>KY=$TY-ZS=XM!Y2>(F#N.!#*B#W%<EP-D70T[CG<N*NDWPWEO
P;(,5Q#*%!U*R4(S\]M64QHWH:]WY) 3J=JC/8=#R?H .@F%%\Z95,^;/!W&>(-7(
PO!:KM;&3ZYA3CWAZ!NI\M1TA!3-P*9+P$)"=,DV"-3$*0A8MBO?$.2^8< )%7XO:
P3XD;[D)22_;OQ'?%W7>E!HRZ!"9*8!V2X/8_R^+E3=TEPR4V='/5=C^_G^/*0"E_
P]T@=V*<O81F*;3B6. \&1=8#J1.I(07U0F&JQ+)5CIU?"+%,>%'RFD*42E*PYS7+
PG$=A=#2GM/K-1C?G&>)](Z)&2NR#[!%]W//D"T(E/"44J/M?0 4ND+A>&"E-CMAM
P;&(,F1KV9'\WFK!X-U]IE>HGN-'D(?5J]Q^GCO2),":L7R/1('VN=<(HKVI<M3,_
P 7X:QQ^3_Z2>NTBA-.M^#/ENW$^IL+K-T"IFEE/TC:7]0S,0S"9$/RR^TU'K.UU*
P9._'"_I7O+$9\@.T"<1P/Z9?W5_5ID@T]55OF([L+B]?\@E7&!3H$CS[V]REO /:
P@CICTC.5<C>G=FLY?&%<Q#T#_?BJ8N'*!\:#01"%>R+9KZE2>2G"EMJ_1:T(GS7Z
PQ&]F8_R/=M3'3P(@S=0%!_P)MJB'ODU<M J RH$]Z"CQY*DG2C<1^0/F66D4;E07
PU!8-F 'GK'':J:RW791*.[VG;NS!4,DTI R*^[849,]5O[)X>K>X2W*$*$T"=:ET
P;>-$8S,@(WKL_X@1PQ!1=@R")99FT1V>A9)>?@]VT^\ .RKRW(:]Y4-$)$? [1&.
P4*^+2NZ$^2CW=PQ-<-@A09$-KGLK!Q$L]C= CM@J%3<9C</^45WX49N^2SX\G#KJ
P%,^ES7VG?'S=Q">J(!J"G-TWA^^8'Y[_]]!YRNZO.((.$>C/,]7Z>$>\W?&>QT^M
PQK!3D=8EB>6?1%-PQ$V=2QW4NTZQC*(O@M77W53(+ICC^P7&4/E$4T0R@Y9 )+ST
P3-.3LRX>CJ$+<4H#&),83TA!)Q;+ND/)*E_R-MNQI"$,_<>94LI9>5 X)#(J:JU-
P;(G0'^^ 0:5B<F=XM3=%!K[@+*@71+ZMW^.P68A"GTWW6RB5SHK6@!V71*B]P5X=
PUU,9)ZD-C;)#;7[C)_9JG%) /TXY0H#@V--GLO6ZEC4J>2>7<PY#;'B[1$)&^T= 
P,IQGR]V 'O?R(^>IL-Y0?I=WM/EL8KPHP$.": _S;^,#@@O#B>^AF4=1#*\RJR?+
P,'ASS8$<Q?;%QI>FJ8^,7?5 *P*\E(H*.-[[QB\W_P_E:@Q">Y;ILXR(6"3)=.SQ
P4AS(F2(06073-OC#E+G(1M,S4<0GX'%Z%_EM:.AB?")WG1F0YY=#P$H.N8BL6*0U
P+. AP)(-]9YEJ4J="?ZF*3M53\-[P[//_ QP'YR.7HKQ!3V-@?+D/KJH3(K_3=@5
P_,F5M1 @Y[JUO!%?1.K)'"N03G-LYFS.+Z.)?S-W'ER6XKL^.8-IF*RQRXPXB0AM
P:'<28UR=($T-0IA4.@GMN0C#]<-$SKFSJO<#^Y!HDWSG,;A1H!F-L_<)+''2,HD$
P0'\J9U/0< 8 6>582Q?P\UH.([DB-29602KP:Q!:HS[[K*3K)748T&YE7&@*#0SW
P88W",#?M3AQ(YQ-XA;)::GT*S1S*C]4<NSA49G;III_W$J2,ZQ6HRG)$%L:,LE@>
PI5Z40X\RB&V?]*"Q(!'STB<JW<R (D>5? [OB[V7LMYO1<LL_53^0Y Q-./T:0KY
PITQ=8X>5^;"6U#0SWXL&2'DZ(J&^!B[Y/<[1%?8QH_=>G8,ZD\C).UAYS41KRO80
PVAR(UD% "P"0$Q UNS]M+D:_(^9BY*I18KE5==NJ4]^UPLB?$TS&WV@:#_ ]7Y24
P]N7M+QLF3F 8I%O0DKPQ#_N5$ ?5=R4[EAE@4M$ (<$\V-V$(BFF_RE!"HKVTIV$
P=5)D<MB&IGE1?P9@/C++5W8#=-R[//!1;CAH ]5B'DA1:\>K *R._-A9:@T*69O&
P&?-UT8H]%K[L0U=K'O:J30@63'"!8DMW=Q[JV.K4NLAI N^PU0RT5;<MGF+T,X.Q
PFG_\UT!FB0.35UH18S,E<>+8DX)KL=']TTE*SC&W#VDV8ULB] A^.ASLV'B]1 =3
PWG&@Z2$U3VA'6IGZFR\F%BZ9*SU95)',1%8 [4M3831=?[Y>L@QSB3&?RQFO@Q&,
P(+KEB^!\*CSXM5ZMY5Q2)$PG'?=_NH"ZG-0O;$("FP%@@?\2.IST^Z7,6__(9S%^
PGI2/#'.#13([JSP%7$W8FPFQHGF3XOXU JG[2CR'BW=!?,4TB.*?1A0Y8?44O5;\
P%%;,VZ>P1<CGK?JQM^;'RK30:AA\C^YVA)C&=K2N3YD?I#%_#]K9YIE>;,3IO21Q
P7PN!S]KJ'#K]?+-$,WB5/0 &HZ:$:\6 J7#G1-VGX-I)G\&5D($*^XY1,E9FQ+#4
PTX1K<V#W:H1]';<]'S)5]6?<35D?YL7I^%J=1T\JKQ#YF^^)G(24G+E=BKY%?&5%
PR<=&IH"TE&U$KNM>J?TG9:(Y.25#OP,"^8&G&2MR;TB;]8Q6-8(I17HN!(D6IQ<F
P63QO$,J8F):1H%#0%JXDPNA/J+*=LD9P.XC%U]XE>!%W^7HLU0LW/AW4PO@/ZO0G
P*<=.QC_9T'[%B;*$52BA3$X!MY#Q^15_$MN0\BR'T!X8P0W8(E )O9'TZ!:LU.L&
PIYQ:F86N@63=@KJ+!*P<S<^['P%&+'C ^=F;UL4:-RR84^MP((G?%4+<QIS*OKI9
PC9WC\"-Q=YR=,0K*Q4-UV9CE1[RZN*;3I-F+<#0-%-&='\U-K+\%B@F++=%.>-5G
PM*\<>%<>VN+ZFM&3%O6!$&^XK3R)LW6EOIA=7^1;,\N]G9[.P#8-\1(L_/Y<A3V2
P?Q[ %FF*%U)FS>"D9Q9OP%Q<C=*#^?\6R< ;DQN-FNR;*6N96AGMT27EP1J<$;)@
P@I7$.Z]T76GD[,; ILU;]>D<[K4U*\JSK"&X D"+&>'BF)'^@@2G.BX':#D5498.
P%AXB\2?DAX.5].A!L:L<03#R50O[QA ],K$%;Q]_$5;;9SBW'7 2WSDTQ^_:#Q=9
P^W?^67;B-N2U6&)F,,"P#'G^B,MCR8Q$GT1W4O_I:.U\&OSJA,M![(3CJ>MOD(>:
P",\R5@Y[7,UJZPT1YBRLB.NH1X9 0B.7GHD7=7ZW;YC9>[6=<;("B-0^J) 9'WPY
PY9N M9J*O']1FHY"TUP53?$EIS:J\_4BRW) )*)64>N#AKKT0?6[4E:$=='\O@=B
PT?P!WMEW]E44]VSFA>+&9KL]X=!/P4]F_:DKQE4\9BNYGV@&>3VVF*\MEN0Z02+I
PPSR!^2LV;WG+G% ><J 8"F]F(J7&)YQ0_5RJT>-//7V?A4I>DH)TR<.2]C&E-/Q6
P\W+,9TW8^;WC00!I.X+96R2"RJ$[<@FQ9^L0O1[L<N0V0 E%O,+?V<A4=\24_:*T
PS^DXTA_6[$\T8V0RT2J*CR0IFD61IZV.B.5TT^#;8N;2@SX.M"QS )26T$8<'!1.
PVOI'%4VY>Z38?+!$B$.)ES[D1B6&7#EP@>(SKCVO\J 8+%R%I"&PJRN CLTY5)>R
PV519?1B %+F@&I;^VS$%'^X_[S?&<*;'[/HG<3BN]X)%^]E//N$?4Q;.47;,WA'/
PS&48HI5VWS8MAV[=+2'B.AW0(XD=^:0&:_-F54SL[K+^!RED3(Y4^)?[ZO?M:6K/
P+7F3Z4"(P82T+ +$95-I'!9OE _!28%D&U@PY=WV?:7*B@T H @E-$@\(8H\"BM8
P]V%6K- 7@GS3YDNJU0HW ^^K=/3NU'I!9"AM<HU4!X6U3IN.3704KKOI9FA2;V+'
PS:W& N&FEX65^S[>?5M_]\':]@+>*D$O&+:2;(+,V@5Q,B,6Y?3R4E3/) +4@,@S
PF+'WXP(1] E-Q)6$2^E LO'QU0&.+^ZR(HI0T"AS9M$A4YH92FYK+>H%.]+,Y)8O
P%R?E-HO46XT9 (V0GS_CB%D/^./9O V1^[%Y/"WZ"WX0!?5;81&4P<X> ;+:X>FH
POPIN3Z^[OJJ3^4SE)B8=PY.[M?JP-_T>Y!;'W?A-&HK]F[D2-/90>^X?[V:RMD%%
PM.*I-@D-?75;*R#PLR/DXN&:=J8NVZ]L*ZWT*,110$7;TFCU^Z<8/!BU349Z@M"A
PY9!Z,<"'7LOR@)N=F69XGP\0&9KEDT?U*=@BH'^&H5QXYV98T6Z-?!.[-ZV*3#RM
PB?&I?AQG\EO&,KO:BP2"[]B*3_171NW(!-[%W49#XJD,^@6/&%O]%F+;J3H^*;SR
P^0_18E.(WP[V9H$?,P3X]<$:CD,#_%1AO/''I&96@+WPHY5ZVY2C_94?:%Z08[.W
PO#NP")4COC3S:<)%FI<YR8-.F,@RUNOTK?MJOJ&G9UH3(%S[C!9C8#N?K%QC\A60
PVJ68/>W>U*J6HTC&.V!B(1B )(LQ:E6@KO@/X]MJ(N^!R_KB,&><B.&&P@I3G9M"
PP:J JA_<FMZANH>;8=HC(FH;DPD<.,L[V$L&H83#^,K\/AY#]LGE5K'3]!Y$BS\V
P@Q"(UCG4:GU\(X9H+@LJPU.DUQ;&F%><;@JV[(5X)<3U_"U9#1<>=-J2@K-%<:?9
P_ 77"CDB7L4FJ!.,N8S>^O+T5PD*I%U,=&+=V:1/Y+--N^M,8D"->=LS@28(;5VO
PBL>@?N<4.7_6<]E*7AQ5X&?Q&/,2_8;6"M3$OU/M^%V$0S8KP/*_)F'W&H@)XB01
P!DCP+ =V!\!'5F,;.H+5OKVDB1-N&HOWNTR!FD6WK$)#YBQ^\-SGV89I?4UKDD:>
P;+Q\'[?$8  5?:=^)E6ZD*AW&UVO_)G#CI8I-URK-*B07G57DG,ZW&3-<^[NXF5R
P.W&:F/0NZI;1UC<FA=4V:,(MAT'Q,GHC /K&=$EU0Y*!'SC=M&1W4NYN%8*<NZ_K
PLYH@^;AH#YY[G^MS\.<,4[G88""8[N4R U2=A43(8O+J%Q) 7%B"+99^_5S$\5#L
PH#=QIOA-4E?V4W4?_3X5%W(465I-D--;#1E^29JT8!<^.![I 1\6\L']_::!]BR^
P>P2$E>!RJ55&GT-_"\7 4MHWB?L3ZEQ1.53_;/#',(DQY)LF49V6O$(S>V"N^.O#
PL7KM9.4<L<.V)K4U(JR0_-')(\'4+TBJNI6.*NZ3?IMB.+G&"?M_4^5$@K9@86\X
P&(9<H$^"]-2U;+O)O_3ZZD/F)Y*TS:O0 0T;.B2CX2K/#TE/IQ&NL=<3Z!A284)4
PRJMKU.'TX5_ZWC<QJ&[WW5_01*&V7*5V[#^WH'IY?DI839I-(O$F< >"X3@ * .(
P%2-I\.8C'G*,6M+_?<L__S9L@>AYD<5>Q&8(&1O!S6FW[9HU5_2E>5E("K@L -JU
POA TU"_6):/9-\H<:L522)8[29C:R@+8/%>G<@;^S(;F_$-81?H=J0BALIM_L_U%
P-Z".Q23!<//MENRO<\N[I"3V*VW"%C" ;^ ]L"5P'"FER,YK&H9W/)W\J@I]<9MV
P7:7:KG-9=E9QJD44^VY9P+925Y"A*;ZMNPAB?=5C;@XPDI]L53P4TZE3 )8KB!(Z
PFH;$B]M1Q%B]Z4<"1_0/'?Z!I<JW?SD"WR'$0:S0QY'"/)!4O0MN^2TSU[JX P(#
P.AR3D][=J-DKJ)KW'[#^UHWZN.I$$3=@^9 IK#P>+!I6]JQV.!V24"RO4F+@;$+,
P!&4T3@ "F15SR,MP12.[_3R^DSD_)1KI48:UM =[>?!0;_4 HVV,;T*6MSH<K_L&
P%%^B-#I';-2V!I)LRV?#?<!$$+PE]QC@&[L,H'HZXH6H.$FD]BWMT,]^NA&';^Y7
PV<WN?2_XTC'OMC8-A-B-PN?+#*E- 06/8=A?=;UA-H:HVC[3@<*UA1=4TM4CDRR]
PQS4<F^"+%V&U9[#MG#*T\":!?WD$%<C&LX]0G1* XXY!A:"R)3PW.?ANP2Y5/ 9;
PLERE_L7T0A52WCF8E+2&0QM_!N%C3OITA5C16=5*V!2'($C.[KJ$1(B,!CF8YA<@
P=+%E\FA#Z[W9?YB:[$5SJ(Y8(;-OV;-=#A6=.LLOUR-V$Y1@T.%\:#/PZB!JSGL@
PE/[<LA_$Q]L9R4^&$?IPM@'\_RWCJJ"50/I"HSN"<)]&M.[W13T#O=>!7SY1'7/2
PXHE'C*@Y?%5%QRUSA )5H.LP2;B#^ORI%:=H@F4\\V,! ZM81N38&NF?]I]48+$%
PA@91]O+;]KXI36F2!5GOAA>R1_%O+NM0*<JP\G#'4)&1*MSVR]S^H$8"@F1E:KO3
P!]P D7YY'7SDOMQ1X)K DYN9>.S#>3XEH'E<1Q2&D C??#;;]!:/!Q<FF-_SG9/%
P["20@A:L('U?.Z-@I:(3&L7IK9#AP(+2&58ZA_].JS2*5@.W4N1[9 $)8VY3*H\J
PF5 >;\)_1/$2#K5$Y9B? C&>.08;]1ZQM F-E^Q*&8Z&27C?@YV,W.MRS@25=W]E
P,?6\[8+Q"A\$SO>'R%O&449"XE:FG& -Z[H48M=)_!8ZFWCI<_\ZF7FXN$#]BYSX
P9 Y!%2 /R9+JRC4.K@BH/';*I(R_*UM)OQ/25QL$5<S6I\:Q9%,O^:@Y#@!)G.J6
PA8?J=AJ.;*#7)RC\5 F@JQ9$F4I ;*^1UCA*65CUD+FO<FZWCU@F"! V(1X=QYD/
P<V'7<Q/VXIJZS3U[49A*(;H,1.XHV"XE-*8G^2Z/RC4+YP"6]E4P K7_&Y48X",^
P/19#GTB%BG&%-:=.39SG.^>+!B^UPRA2R K5T(OZMT1"V;F)2"Y!ZF-",W<_4@<G
PC'U>$T>>."+K/I^$IE@MZU&)1E?YUIRBQFS-9?\_U9VJ*_RK*%WM_L]6Q*2LE(>H
PS5(L7!-&V 6"7^4N7O;.!5;.95FBHN<AZT?"8YGJ'!ZV7)487'+(%#$B3''!Y6VJ
P^JJ-WT3>V8Y((N-X#!S^C/#0+N!LV:B)/_$AK+,V'GG0&'UE+C_[^Y]U9G'XC=IX
PNMT_W\V>H06,&A-H.!+((6&4%&M\AL[I/-YO%R75%*9C288WB/CA:$GIL68*3Z]Z
PI/6S!K8'J1',;#G(N)>'91U#9=3)#&H;C2XKECM'&$BLW0TD%S#P_TIF,<,A[4V.
P$Q]]XG&<#3.:Z=/I=L\@I86 ^%D0S5=:B5,(UN=M!QDU;;V1V*]AB8/23P=+@SLK
P#JJ3=YL&4PJ;.443L$Q#&.%Y'O"*$JC-=D+Z2V93#A"KG?U(4%)&Q^X'H4'6UTH&
PRY/*\ +;W%K(-C'&I+N=E3>]*-4]F;. #&&)L,03@=.0:5-J/Y\NO8HK+>A[IIZ7
PX6(G*A:NY0-:S>@R">H22,27'+T<@F!=Z(H%4$%LH&X-8 4T8C^>^BIQM3-*]?M?
P-3JW_P3L1F.BLPHG]QM>#@$_3X7DRRCNON>EW)S5A&,:)/\(<&\1G6V!F+;YF3!^
PK"2].CVC"8Z1?W"Y[4,SSJ#;,(!E5U)V@/V,753.R<RL9O+K,4 UI,#4B8#U#A$A
P#N!"]@:O#;S K+%[Y>J3FK!?%@2G#^W!GYO;%_'.?S?OIJ+1NS:$*]I$@_$FB?!J
P2M#]$"7ZTJ9F?6*U6[WCLQ&*N'?7V=Q4:%5"6Q,>U)76A8AMEQCD=3;?S,?A^_LV
PRUV-OOL)(<G5+DQ)!($<-BW6M]7])7V"BZBJ0&PAIOX7[Z,@A=I4M+R;9#+;'X(Z
PK87>DA6!WBQ6$4;KQ:2XZK[#;S4"[&$O==*O !'A3O0+W-,D#6<NOK]_@'0CF1Z>
PE:Z<C-O.3[3&)Q*0H;!$@'6+2I:"U4%;77V<;D]6"+.3*\CVD+Y',A"LA$1.GN0*
PG6G =_MV'@\2(&QZ)(+_%V5&33L#$B51? A,]VW"L[T ;GX>/G.26%\$#.^U0-=_
PM]ZWO1L.S0=:376&8?VI[#.PH[\!"D^MC]O)\-WQ\@/BH3O#>^4+W\$9A;/&?_;,
P]^UJ[?L8TD<42&<FI(+F"Y7RIYEEJLN\*YG7\,;E&KU#,VQ_R@CN?AB]T45:UL5 
P:P;9]=O]SG4?I98<.=V KM!B5$ 91:^<9(X7@C)HC.!$IBV%A/>(HK68BQ<FF&)\
PS 21?$!I<PS!NWI-*+NTGO@E4*^&! =8J;9GUE#N_3L2V;*HW/H'+*Q?.!.-L>UT
P0:+X:^<H?JOH@$N56^U7WQVYO(/K?\U7HK?C-_X/#9#^7TEO4;*^G\XF5"$- O+$
P=TM'4;LYT,PI5'$OE;,L45!9VC$I_KMB@P!>+5 U%IVQ+1)YGG,S1"T^ [<\(?"?
P(N.6H1,2G]3Y?TVN2*17+)F_4+NAX<FX< NV JG!4Z@A/[>J,*8;XU94KM=5GF=!
P_4?F*4@,CD+KE_)LT^B4YPTCVDXX*LA?W6[MWBL!3ND(0$^W9^%K:(7H&; 2+-)T
P(LD;]7QKEZ+0:':QB[%U!,+MPBL__+0!;1EG3?RGDA<W P .Q?ZH0[A+3T0B]=H9
P\V"6* G7 FFGC/<&GNY>DZF37E^]>^HE_,DH@UU1$:0D ;]"/NP\91L><".2 S;3
P\U 155!O12,?JK8B T6G?8EG*N6%H7VC"8R_JP;U7I6O\GK$U9)YZRV;6V+X0$Q)
PF-$AKP$Q(ZN1MA?!$@L2TSF[A-<<OI&GV&UG7C?=.NXZT2=+WS/#]X(5BS$1_UA!
PM3SV[VU_E19N]DFBD8P9#H.2J&VHER+D RM=*;^]N=9_VWD#!3U34"ME75L%E'C6
PCQ3E5.E+9BSDG%UILOX-$QKRJG,I1<:YM ]PRQ;<Y4OSVJ'HL**=G@@]/0;O]W"@
P_@]$K])$!]R39C9\GC3";1J%^VL,J@#/SIT4RLI%KB\3BJ&L4;%\@SWA/[MM$F2B
PLX7SRY4DW.YNI;<NLF,8AP8%&^GC (9H9TBU1!P=_,8MB0A!5;UJS#]*TFU WQDK
PO!XB4R5TM'^)V IDFL=.];A@!VA0L617A*FOP3$)[Y>#R<?^[^)VI1E^H7",0^P^
PX3N;CEVR$=_VBH7><W.6&I$+%,LE:\?' 1]U05Q/_PRZUB<QO$F-KP^__I4B8&SS
P2>3TUM2:#9E_&$VN"8 G3$1/X<H$297(^1"O=U29Q=\L3!:4O.P7R^ [%JJELM+-
PV;[$;GJGG*U)PELA24BX(''*HORL1^Q S;6+='Y4YQ.)V= [9\,JW]%!UE#Z70_R
P,DFVDRJE_!E[E&\4]!9[5.#6'VPNA%9HS0<==YO1!1E!>.P=T; 'S%:;0<?0J#]$
P#_*6L6AE&TO1S<6^54/[%P[^:*83%F*HGYY>-8FDLLAT?O^>@2PA'*1F+3/U9[ S
PKP4ID9+AD ]Y+&BKC1">?9N:$PB:]BQ\E? 5_+-!^<OL"J\"'ZJ9AFM!B?;F&E]M
P5/P24F,\;]^70ZB$T4]JJSE=8)IVUQO O(6>5Z7V,Z$@'<A$?^@9A=?@LF<N_\#>
P$GEH $PD4_F6A4;,UU;$)970L_5 "HC!9#X(>@5L:/-(6$2 UTR1^&Q'_+F8:, "
PP%[\<DBCU.U:1#+:?")2H];-N_S->5=B6M2]=!0'H?^@)11=:!#WVZK,W]7?*_L;
P^M"$_O(>:-\]016>!X1YH^-6Y8H/&UM\(2L6F5PM>%4-0<VK?*BS6JKZ?WJI*NVD
PW7Z6-':)&ZJGKFQ^&>>W=%Z5.EJCFQW,!0N=<EW&@-]M>JHJ_'@XRM@P[!3K=@JR
PH+$#*PO4HG6^HDI@,M1I[AZ^'[?_U8U([)Q&C#ZD+%AP+FI>YGTL+D!KQR0R)0P?
P>-L98JI</L).6@GEW<(_T"53:7Y5E@N9@.PEG-1?L@#'VN(]$"[:"GQ!LS^"CITP
PKL4FV>\N,IIY]_;L:R(I N(>!Y)P]-2@8<!DXX]-D-?LS*9&J67?!: &9:K>[J_+
PC;0BRE/9I+MJFS?Y9$@8JBNX(#'(M[N/+T@^'[-N=%(55N^:M2 @U:AXRZS^R%;)
PQBH=Z5G!#WS^O*-=-/9X)(N>#6 1;05MT@0A;4-TH",H:^P:/3%L??(MB/_"Q$]\
PJ+ ?";5%@#!_0DH(ZHNC?NUHI'Z^#OG%-/7=DIE QL^?:"\K\&9\%5;"C37KU+N_
PD8\?%[; (ZKFAQD@O3/<R+P<9=B3&'GQ%!$\0CY7N"?Q/5J,T8^M3]_4_HCI3ST\
PRB$.,A7A<JVV#7=(<U789P]@G,3*#;?HY,KS7D;X$"ERU0CJI$:20%T.1(+E0WV0
PI^.ZGQXP8%%7^"<U:@UM"8RK3T#MKA(2+PI3X401@WN]3)S0[&*LYWMEF4^5JPPR
P)^B*(,F1D7HA(4JPJ+8W LGU2";]I/']GO<ZO<"VK[VG&"RKEQ#JWHM&.0_-.=K3
P?1,.'*7AIQ]=A60085.M1>RR8*$G_HQ]WDSX]E)?&#>^%OQII-K<#AV*BI,@K>VM
PR86K16FC*$UP#N#2&</^7C+09PZ,VQX,I%L 4'PB,DB,18H-_C$.37;N20L>F4>G
PT#( /)HHN/L:\@,659[']S:L--W&[I\(&N%;NQD=CA ;F"HP'>B*:+,K(5)M*24B
P.)NF[CR6?;')W>"+=551YS^'FKKR5!>V+,[%:.#@J9/NM@!>&Z@(V;/@_7GAC]8,
P._[5XT[%@W6"J7I /NS;D"[=&A.6UVI3"\,5(+ _*ES5%$4;UPCJ\E^Q!X66LX6;
P5(%@ .S-N&I&G$\W!F[,]*SBS#*8R';H0;PSV#1M]8O]NV!W;A8FO[.A\WVX1B<;
PDIL.F4U2T%HM1*QLY]0(+GD'<<H1)6_Z@G!.K6A-W2",U ]&"!.+=Q3B* 19L$C3
P2M=LJ>][+&B7HCG50>#X6D&!)=><=Q9QS(B)6$/U?8%7"(=>[D/A9=>N[I6.Q8;]
POM1)QJ4Q-9Z*K*NS3'/'7>A8D>4!G0I. .T;]HS?L=:$@&#+"9DD97&V*-KRGJ;Y
P"F)]S(TW'Y5"DY<X]9I9/2I70R?"N$((9R!,NO)%>Z79 ,/T*-\)ROMEE4_Q7G4Z
P$A[UH1NA3U(G2H<5[,G]Y^U^1J3,[1FV#LN9"LH);W>9&,ID&SK,")@(XVGYJ2=+
PQ<&LBV".2ZE24Y/29:'@N!.C.3E,VMB@E_COD5ZHNF>4.Y\00GKZ:54)E3P- UV_
P##S: OW/X!G,+..?D?:DX,QAHT\T4^D]W0%"),BE%-:Y<L%VN>F2(M",S&E ?Y(D
P(6 =)/_J*C8D6S*<<%[+3<]+0V[O.S]$*DEJO$%G K95JFU5'CX.QKU+.OW'E_AR
P\_> &^_7)W/K3DK&B 8]'9WW^&U'":0 CMC1BP;M56A$#(V5[R8.]A1C3/#^EMSR
P- /XQ@I_].=W.E1!W+WA-+:.$^2#F'I>GN6N8\@8:H5ZAP\TL?EC4W/)BCHWF=&5
PY@$3"*(]^T.*I&D=%7F.HWIKP)K:/*\YW6M+@>WJ+9G#P$_P7Q0H\.0P*/H(A5RF
P8QA25Y:7PG?-4[R O+P=A>V2;D&(%7L(% %HW,Q"$LJ![B>^7H3TGRO8R'%DC5B9
P/+]M]!V--(-*P?>\7@IYR!/N\C@3EO3"<@@GMHC)!A0$;#"(6>D3;B0:33(QG@DT
PJNKS*#HN32D7! =C0915\L:!D2X&9'T$)#]9R,,YPEJ.EK8)=3J30Y]!7]W;+ B$
P\13LIZX)+YNOME->';USW>KS:AAB-EXD)OUC<W!*S/G/$[MLIY^H:VZZ;$C6'6Q8
P3JA4D"T'M?0HNBN?ES]06'^7_( 8[%.AA:*V67FM\+\9YO#XWAFHG2Y3;7;EF;;^
PK9CVNM/8)J6/\T(&T8<D]14+S8X6>*GW!L(P;G]Q\<FP$# ),RP!X="1X;DT?)#\
PN<0E-Z_!TBC[W&-GUYSTF0Z[%D++">A7#HW*JN[<8'M?T2Y94.U)N&B0BN-<6!3Y
P+UW((.U=#U-(0/9LC> 1C<#D!,L7$. \,BHJ[US6G$ *4C^?)NJHC5Z]AF")OBII
PO7!8$P)M:\W"0<>"?8?4ON7%/_R)@6G.ZH%"[/*0'A9)5/<8OG:2''L%L&E+LJTW
P[3&N+<L#41RL:O' EK 9&9@^HRNK9K<CW\KJS<&=IL@0$QD=B*B%]$B6.VW_&# \
PQ#]<_E\X_G]K4(5Z HH%N.(O@U!N$8<6QN']Q44-"U?Z6$G9)W9\B!K4\."I/.;A
P3='>#EJI[KI4TV$YW&('H^A:@I/8K]WJ&]$J5%N)_>D]TS,7TF[!V[6@Y2L\*<_7
P]F>-\/BL,W0<N#(0X[%$4_A?&")Y\^0#KFB8-\;<ZG?YQ\P8[>^J2!ND<U",MRXO
PI\Q8&BEP#5)E=-P*8S0'KI3))YTG,4S$5(C?3-'E@IWN#BU[[XHZI44M!$(G]-V@
P6LOF]Q9WT]A _PA,,-#Y4:S2-AX2B_2W':A/<'@SE%7&S5S2B59,MI9/[UQKGXNK
P;Y[IAY9FPDL]E!>!%Z10D\&QH"Q <,Z@>Q!5+3[ "I=WAM(=E$<C R)_"9)32 Q,
PZA))3F1!''I14;^>9IH\NZ4N#(N& D0R7F_DB:B9- H9NM-/*\_ZN]LF+&3X;4[Z
PW<>+&Y+ 8(E8=^WZK\(NS=2 ]]$D'?9"N <<?T]AIBE)QF5>*?#RZ=[1Y+*$*"_C
P(L>Y/Y$_#KZYI1N0VK^Q*07_=YY<29W,;^$MNRV!^59$L\@.TZ;2@];.>'0LMN(,
P!=1" E(F(T[- '$;$4NCE]@QE096>X$!+0B&?4=!>8%O);99,!!$WC/0KER!M'>&
PTO;+<=WPF/E"3>>[J3E[=P8J+!$&PQZR?+?UF@V"UTO:BHK3D[3S/)G9P@X=>=>P
PKRGAJE8JO",VJQ5\7.+&"30H-9X3"_$5"D! <LED;""L@%3VST)] G2#[YLJ(!2H
P)2$X'9GG$UVJ@YQ:V0J)(&.8-/DL:X:BBH0;Y*:4?I$#+@A-6)+*0P>=0V=1X03'
P:M=X(6ZGOY[WVO([Z05Z$M%LN5]=-,>?CBB#W7-.H*,V1+[Y#B#":,W8N^1X;H>,
PLL7Z=OC^7=MGM0[KL]G&EWVD5H)2\(5HX]+LE=M+?_)Q.+E8$V1* 6 5[QYNF'.3
PS+SONZ%*U!+U^3'<ZCOH[%5Q>/!J->-E5347CAJC VV\5I?K]* 05YU$0B'*2E""
PRM37P_KP+%\VPP.VM8SOE!NKVY$I]^<K>>@(FN6U]G\]'"(/2>:'L$%5*AJN7;%9
P@[W89XSXU J_:B!V?H%6;#+SL"/Y939GXQ$&WQ^6PE5&YD+N=NQ?2*\K3!12V\7Z
P(RV,61*9A'PK!ZL^:_9'(,+E: \+M><F4^YZ-6^><ZO(?L/F9T291NI'<*%]^99[
P@!D>+ZU)B*\Q(_<! Y<_T@ZJ1>+'^\&Y?_38OK;#*3W*Z[93NSPWL,'^(&8Y"M #
P#OFARJP=<%X#:J(-YP.YE&5Q:_"R8,P[L2R !?/+.-"DRU7M3?KR 6##3]136=ZK
PM#R(W*,T\C575&F0ZR7:$$)S+S*_/M1.H^5UD3JX\4,4\D\1725L"D:Z80VK?JF6
P[1B8_P%-4:5L^960D3.)R:%( ZC9IY3R'$#Z.]D:L*^;GVJ7H.((MA;U73LQ<K=N
P;%.:BXN/*,4TT"H98BR!%K,C\GU@)@;>(Z1Z(\KI.]]_0#QK]-@#$%R0$>*<(I"B
P01^*RSP-J#F8,P@.V)1*/"ZHFD'F3993S[ JV._'K3W\M*S?@*-PI(158S<\Z.1%
P_3J(KO(QD)[_9JX(^K1&T4NBT48U<8UPO]+M'(B73&UQ;C8OMTC>>#T8CZXO,/X>
P""3J\=X]WO>'_4Q(C.Y0=JN@=>BU>2JR%=%0*ID-Q/C]P73.8TA1/.8"8/K2_7 7
P@.AU/5<5.SR@">X@;$:JL2SN(+80NLEVFS7#9HDZ-J[3+N]80$&^0"RQ8@7M_/C/
P[ZHLTH&%!HQB^; QO)3L(7U:0V)\&,'N?^$IVAXLHYO:M!P8=S0.G!?_%%15HJAH
PBAREZ5E];G3^=/KG..G#K=-9]AIT-J)*G]C8F )!WJ3C0B_-F$;T-YGQ%_0<O41W
PL(1#2V\8:F)Q6.HHO&'8^B(1OM0DE7=O8M+CI?JT>U&P4@P=I=^(:@)@:>9W(LTF
P]PQDPC]<V?TZOZRF6DY:MBN1A<",6UQW? ?M#10BFKJ7Z7FS[Z[SJ_.63A#DF>[X
P*SR%UU7(+Z>Z";D&\S"P>>J0A@I7#(22[Y8AR"@[HKN5$T<F//?$GKFD </&LXN]
P[1,O[+4E)&_/JXK\F4VM"X=R57%:MJI,7NP0NA>-!RT2ZSB \(9E>O"M1Q(),:X_
PQO77Z8$>1<7#VO5&L. VQG=\I )/HWLCL_TJJ?(KOW^6)_0%_HQP$9J@?DC@E#2I
P4(9@XFVI2Z:FF+BD13(,1URJS)CCK =0Y@N&4C@Y04471K>:$/-$E[%=6QGIL0,>
P1B8O5@LW<6X&2^U:CG'!KTC,KXI63H:J0-X6;,BT;QZM5[9^''D:X_ULF^6$*4M!
P$BTW"+!1"H_A4N#V>\='A_0C6UTZV>'#7UW\_%8;IM8]5,LOKF+EV'Q21H93\<RY
PG' W.OHDV5VO=$92U=B5!P@A#;PYB*A+A1<I0TL2UXXV;@;-V/>XU]+J!RR=HQQ'
PB24$4XRJI-0 ;)M:I_$>*;=]L-^?A2AN_.4;72!T&/[3(= 7K^YYY7!L4G._8;78
PXCCE-ODCC[8@KNOC2AX89!3YRO5WU"@:[9T[G&V:6%Y6YS[MIO.)8]KF-2(WH5E"
P64[Z[MUE9 ?-9K?]N5:YYN0X\>1X&B:?U/\7HDG&[*_;SZ>0=*HAY*/1FI>-H+QO
P)I/-@7;D:2"2^>;_,=MMS0(#I"<425_^N99.HM^&P785<[#96U2+-N.4-DYI EC>
P@^U?RQ%RL)@OM9F 6Z=GAD?7_@GRSY1_"0'L5?*A_?_B7X&*H/]:0J($F,?O.<G3
PTWUL7"'#0#\,E QR!%$%57DT(6(O'9FXD=@-][3FU"0^(M%$*8Z0P?DP;![Y:FK/
P_ZK%,>A)[K+U$_V-I9QOKL. I10?>'W1]VHL,S,51$N.UHG3Y*F13&_D;QPJ(^E#
P11S72[W4O'^#4<(R#5^[?,M\*TY@DEFGP77*$5BNKB+4_IOG\>RE[G_3K:X#KD,,
P.XH$A+@1L45%.1PN+E%H8)Y\P_-\+]$<]S^QA7QKNCX5642Q@AOQK.Y\;3;&NTB/
P"S_<3KN5^$T6$W*FYJ\(?&!4VG:2,%0]L80**LPW@=Z\'#6W[E2OA9*1<MO[2ABE
P@3Q UD=C5#SC-R*W\7'FVK25A<>8'''@B#15KPP&&P(IC^2!:NP1 Y>)V/'$&/(P
PL?V61 ?E ?,?,YX#+@L&2&&N,V4^]BB#KWT5AFC< [#I/,4%CYPR9*[A?3384BU6
P#P^ZROZ1"E_W9V4 &7X<]8S-K?P"6@-#)%^"7[QQ2TJ]]3?&#_H0V\:4G!7:KQ.O
P8$[7[:&XW."QM'<AY27C9&M'@>"UY\JEA,1=/Y5ECNN &T&;.7$ET?"B;%7F?[2P
P(T>*GM6-L++K@./Y<X_DNS2N<Q#F),YM<GU3Z=PU#&-?%DYIEC*$Y-Q<OLWM=^YG
PK???@&US,.4P<#<)M4Z.[LJ[ZDAV(B^"O4X8':*NK&'>9AF)LT@$\L^@2M\?)*QY
P(-(WME,0;&AE*U'!SW\CWP"981N#D@9L0)C6$E>QQ_-KUG-^0<L$)25@@:[$/F^A
P*^GO1D>%P%4U-_XEFXG/K,=V&U)]K3E&Q_@-("ED/NJKP%9EJ]:5K" H7>Z8Z-R%
P:(3,5RO88;)Z#H?SW[XA04'GPJ<HD$)YW:W<TVUCO\BDKH<QX>L7?ZG43SYOW WR
PI2H*ZGFV_GD)SL5>;\UD%Y=T)]AD[HF8F135T'D1CA< PU&<2IIBVQHH&L,EE2<5
PP"_#SOX\43F*2/Y2U3KAQS3M'(/E]6X5)"-"(Q+[B&SNY66=B/^TL9BN_"S)C58@
P2F;LJC0Z-<\$2"#LETH*M5*.:&NI**10!ZRQ.HP\@[7=+CDO:2H*:NMU]$GJ'X'A
P* ^X,>SB?L'J/AU(D4X8E5L4S%%FYZ*)J8>#32RH<",WN!*)<W[\W3;<A@$+LB %
P!21F>>:WD]V<@++JSZ?#E'%VQ<RYX/L77P23%"G" BD=](;#UZX)9E-!/38:!NDC
P0+ETO\U$FR!FG9Z=MQ3\?7.&)4AEZ #I+]=Y=3FMA^U^BES1J4-[AE_TQ[UD0')=
P 8SWDDY)L;QRR_YK<0D=%"0: D(49 F"S&85NQ)BI3V^ZZ./!B.D/8$[I#E@ZLA'
P-I7<M#6%1"U=@!3R"@Q3M[&I!4M/*TIUPZ-'DZ,NA_Q)"ZG/ "6N;)]1B%;GJ!B\
P8+*&A(<Z.J?4I4X(_YM=APKU>! P.&NQ)=?DL]=BGS*JH;ST'/(#I"1GNSI?0RT^
PW.>._7S+[R59%!!I@2Q0$+<6XB58E&B^F)O+02:'8S750.9IPL_588SB?AQ5G ,#
P3"74F$*YWZOFBSPG9:B2;/ U*@].-&5<DT'Q4.Q&<,PV'WK'TL>]AZK!>.2AN^L+
P(SY'DQZ+=5#_A*J:[?QZL \K(6C=8R"A9!O7-9S?]XUC"LHD_EX[XB,%H@/O1K?0
P9@T"0V6?3LZ2<[XSMB+Q^U$X*4:)6:WJH6V1H.F&(G'G\Q\:,8IVO6S^S\C5B^=/
PIE?<E?U8A.2))!4RKU:Y_@0<-M#Q[\H>0),(#RVDIV:*TJM,>GXAN'1NF(O=1,(X
P&U%-Y',S$J;JJ]^6AVS(Y[C?S[%*\BEL&WMO%_3W!)48%](N".0PC>SKHF P6L_%
P^ BXB!W[#[52$UL_VYUXG/.;B14:Z-Z;SVEC]]."3J:%*P*Y5?,'P,PY_5P8)D*B
P'88'JW\!XM<552%5\-;IH@N'$04W%&5\Q36E\G5PU-P4U GYQ%N\*&%R9GX[OU)9
P*7@%.'S[Q<C(A@<@IB+Q&I\?)C9.S2@IR/\<!#($>)]A:#&<1_K$ 4)L;<6S>X\2
P>&C7G]45M(G.4&IT<?[(XT.?R+I &3PXWZ< T$6T;L07L]0SO8%0F]1(GAZK>2E(
PCB>KT4NC0F,E7H<.YE?RMM<L7C0G/8RGL6 .? GH!UQ9,@!7NRI?.'ZXW?I;B5H1
P]6GUQ[ 'VA"&_'(N\1%Q:8)E!1E' D $L2*V\ 9#E]DA[8\9T$,6]I2*[K)[_GV]
PR$YO7'7I1:WGP9C+M!JISQ<W?^*/5;WP#&=F%3L3QX5<W+ TK9KA3I _(_GSYAA&
PZX.I,V?ZLAQ<N%^V%A-\Q%W;?AM]Z+7&C>Y13T"3^&@7K35J(N@_&C%X;.EWTY8>
P3PQ)L/1[<S/J%%N6#[AT::\;CST"J$(.%8[[FV"!(E92&BO"[23U*'<]D<;<(6)?
P7<(]WJC 6C)99=F&$YK&$(*'K,^<_F>AJ-&I^![*]&=6DS95TTY@V3J.BI]1*Y(-
PZ1YK%GB3"-YU,[UZFC(^7[W&AO@!,LE? =1J$<M!</,WK[P5G:?WR_,&M  Q:7@9
P;&2E@\P'P=:YQP/R.)Q_*[,UL+*GR]/[ P&*B@4-JQ>>3276&&M6Z-72WDDQP7^4
P%KBTF26[(5*#A30B?0=I35,=A7C,JW&-? ;="7U_H9AXT='()+Q_?F%00.\NG</J
PBTF_8VY+AO:$5HR]E.X3 Z,^RX@Q,,00&2(]:KD&?Z^;0BEZBCC@F^WD[2(5['Z$
P8TU[^.9KY%2D&2%(I_D1.>H'0[YV5(9:17CAG'GGT:'17?QSLJLX:M"6KO:<F@GR
P40^]\0JB5&^M[P)C&>^COG@O2#GF!>U_.?9G#N??5]/\;1O9X+N3JT;*%ALNF87I
P)17\2D<4?H-K678ZUOU=HM:TJ'R_V)3NY#@NN)R!R)Q/HFS\ T >T5JM=;)\\48)
P@Y*!IPS3I6]"'(2F.6\X $A6UD^J@Y@@%ZDBZKVP6P1'2L4,'+D#AY-^B Y_VA^$
P_U,-]H4VB^MU$;.0>_R;D]690#>MB=>:' !&N,[AR\2_(/O_KP._\E>95]_&C#E3
P*XK5ER]4[R$0DF]K;S K8<]8]5*T-3P/U>8",8Q+X!O9IJ@]?/Q,N &G90;"M354
P^*OS)C7-9EG=A9=1Z" ^P)#Q"4>=-"K7GLU?IO?/<53=V\R_&&R7XY_;R)ONI8L8
PI?>:]*9GKB9OW6VX4$=R,6;*>J[NVA7NYP\,KB'\C&U.-^@S0W.[ PN)I+=UJ:#'
P70Q("/^$J0<5+LH^8S1'<76&\5L7;@-W+EE2I8Q&IF]C')V9(9Z+E18['R:]U.C<
PO4#N-=(S=*??;VR'GFS-5LKO-&-LBU'"TLF)9'PLZ<Q0-'F!#P,5-?$L1W(,4HNU
P%+1SV@3_<EI(7%.3B;XB:QUY6<CO_!(U@0^<:$X>/N7K7X[@-FKA_VB:UL*-5J89
P^FB%+@:^3*:0D/!!P@C8S#;]0IYD%) B5\N2EJ2A,L&E7@XM\8WWL[_2'Z<:IVW_
P,J]4O="[4'+L:&&U\K/:S\_DD'&>LP>$PF,&VM.72IS"SA>4P,7^>E#$#^OSL$(9
P]%\ B=(26(]CFU*>$F_O+(;?#.?@\9A(7IOJI@7@N/8PAP47\;7^V64N\]$;<[H>
P"X1F:-ZH9*)P)40:=2WJD0-3KFW ZVY#>?&RW4,"#(B1U2E'8WI-*6/F<0A\.<1$
P0VQ:4H\$)'B+0=76%(6.%]J% 7RV2J><(&T><@GEO^)W  H\%-5[KI6ZO/5/QCH]
PF9K'#C%#[]3D7')@G[8:32H'D;TG/=,EDPVC,(,IR$N,O1^?+HY%0<H-D&:C/Q#D
P3!T!86T!R&UM]7OH#69*CL7%<NHW0]UV?%Q+MI?(Q&,ZT@K\BQOGQ0,^^F-MT%D:
P8XN50AMYAA;L8F'K2#I++E$5$%VD:-6I&^6S&4:[*66*DQDNYST9;LVMM($N.L7C
PDGWJ(9E":I[I/C?*^$_,?^-,F<M]?8\NOZ:^03,DQ_('73=;B*ZBF0H]$9QPJE"O
PKLDY8,>4+2@S1:S#\-DP"%\9?4-OJ' :WA4L=UX=R5=Z092'N_G!P?X?$@FWZ^\!
PAV!FI K..O+BT:M 6R-G&S,QP4PD6"$M=!'9\3C5TSC:1>PO&VFY)<5V_N8$-0CL
PQS8[6&]%64:5'()T88U3?3C[8RI.U!O\2UJFW'V;6D.CO>$HW9Z>'F/O5X\ASGV3
P=+^1K:)=J@-/6"?=BIV7$--FL-C?:OQ=L_/%<XDXTRF(J+&#A;3U71?0TOQ Y#!"
PI6:;;CP7(C/5O3921@AA'+FD4?C7NWN]]DZ8L'P=Y(K%<R=EI_6H#D)N6Y=C4[\O
PB9K-+/"YP,OFS,"#&ZA!P3[D!_=/F!Y!&H6FT;+ 7H%_NLL>'??(:"[/W3[VE,Z6
P;#YJA (U >(!Q=0-)D;B@_6E#=3YU542R?B>"])M$[B(,*E![ RWBIG/;?.:.5:.
PJG@O35S,O?KV[J>.73Z>4FH0Z1JC0S #XP&'O= 8BWX)A#_<#8 '<.&T/( M/:X9
PTC77VWK0HF\7U.2$>YY:NQ/3J;M,$6Q^@.G?6_&J<QR3*' P4V8?Y\MD?CP\QPGF
PE/SE:+8]%3AULA>TO 80\\_:,U9)I*9+0\]99#29CUM3D]B1G#P6NU'.1Y;%$;:]
P#SC+5+2=9+]DLO=L-[$/O=HT#E[)6%3-?$1Q :V>'32%"$%[X?9P2^YRNR9_"_Y!
P$-5-V#C30E#2L:(_(;ZU\^Q"/8.T\>N+LF2T?:,V[RU<37I^#URYG(I1%5K>=R^<
P_K-$#?Z%5L6L"3*256-*&!!AS60!W9]]63JOH )I>9]\DPVPNCTST3R_@BI)AZ?I
P(>ENK^3VX>"OLS<FF> =/62*?UG4&-6K=/*J0Z#?IR=V8QT*7*[QW4X="-B'1"$C
P\P1[S/FW'=7BU$G^."-V!++MS[4T^@BEU#GQ?;:!K?ST**%_=EURWPM83^X.AO )
P55N?!EUC)?:1Z.'4OXD%(LJ+':C'(JS3LT:=T"<?&XK:Y$N [/5Y,%#GA+!@3DX^
P0[:(*J 6!2H&:9@.%X]VG.UNO!YT;.P<!7 "JN'(1'H5ECUQKD\C9B<=7NI-'@OT
P*1O9(V(4#<B&HM/7#^#'W2I$.*,-0IB^ *\V_.Y(-E)3DQ"K \0N3?XSO.@,,0[K
P#I=_^X\%9_[+DA3W42&/BKR,98$F ;4C6GD87I#@0RZ* 65]4EFQQ9\)YT4FQ =#
P>]PR\54?&1+8#L\<M>%I44LE4 #U/3#;*Q<M7XD#9%G!V+=!]^@>6M![=Y7K</1"
PQH=7>TREDH9!*)S.E#_%#C1RY^UO=7.=66=S^FQC^+WK!!RD5%_4YW5UW%B+$T$Z
P34]]E^+^!-)D2UZYV?J(L_] 1V-LRU.C7H+"J;(2U&.#ATPA_>G$GQBE'GO9GDA-
PM^&<_64J+]NKR@3Q2-[D+<T"Z]#.>*-Z0P_F-_=#0X7A5=]U$8.1N('CGG]+^2)A
P$$2._LO"/%FG#MZ?G*,3H&(^C8>W&ND!:G#/.F1Z6GIEON_3$&/NE@4B9V2WJ@/B
PK<D!#LU[X+_2_=39-D#S*.]6B 2!?A [L6[[FBF2%8E"<4T4?IE1W@:L+ P*%_\7
PH[.M,=^?N$S Q54%TOQO(O,"K^ 5M+!R8$1H'V_UDK Q(E!"5X$F5Y4VD!FC#2C>
P]1!;J(4OCC]2N]OFFU!1%.S$FJE"F6Q)V_SD2[$$&\#;0MOU66N+N_D-17Q<Z!R1
P(+8%H?8C80)SB$'%2E;?QT)ML340PY\)7]+5 K+I4M=RM!--"PC$0B65WW!\PMZ!
P#9P.DEQ V)[$0\)_:%<2F:B52!<@W*W3X1*ZU=0 6D= Y=R9B!"KK=:A](\R" AH
PU%A$"!$U#,;+8:Y/\:G7:!06!:> QJD!49O [O7IT=!C3'_4 2K7 K7X66_,-9@X
PT:EJ@W37^^T;@.MZ34<XL#%32QEQZ-,0@".RS"]RVYRG;\1$&75,LT3/<'F-/"I6
P.6TS,9 EH1NT?/AMH!;>?HIBYD_FUQ'7VG$)6-:N2T.OR<TLBHN]FM\B5H+;(/:?
P>OTC[F90H99,X/?:?6Z#1<^-/A91A>B%Q=BP-^A ZG4D^N,T)C;*$-/89R>'1="4
P/?&I]*>#T]8A5W?JRXYP2[24;^<WAH+&T[@HVBWA2=8;R*Y&*CY\O>2(PK-<.\C3
P@%@IRJ5 -;&:OR]&#_5A4-X@L)2@:0@6K:O!0]''@>)D&^KSP 3^^$-968^##+EY
P#=[N'FP&QH7:^4)H\L+=1*.E/)&>+!(H@4^E$J#-PE_=3N7@14L5^ )<<*3O,/A2
P(#I ]ZWY']_?NZ@G@XX8L/$0P-*VU'_/5H_U&>F+9>UZ_<S /.S2(_+VY'EFBOI]
P4MZ,_!-D6C\TI \G@NI7IF4 #TQR;BAG4+P,"DN!:.TLN$)D$Y_M/2:EG:-EZI"!
PFNM?1JRE=$Q'>S!;M(%")TP+@D*,;6'_ARLSV:Q2.V9O:PG6=K(L'F# @(2HS$D)
PM):&M7K[ZVM?^UK,=:1/^""S,3L[@/*8N-8D"(LH5_&J+ZX\UZG@;Y(1VA0B518B
P%,4UCG:R/N"< '0TQT7-]@TJ%E-G$$2&!I%1L!:R+J*8*MQFCX]JFIIS^-/)'606
P)&3G2;;]1K<R"%7!]>#D9&G68:/0G;O%"4%O1)(15]Y8,/>S/=]L*& E(3\L+YXD
P#"^BVBM*AT:0U.\_^70_)  )X7&2(P;/E].#"M&]]<YP*"B5L0I!+*G]?B'-[B&X
PRON.I>HX[E0H5F_DB*]:3(-6+'O]!>/PF;FDB, 5>;>-II$3D5,WHN<@)[SPI0ZN
P_6'/7!1,S5Q+0\QO&,1!^=(('#A^A)D9HVV4<WF.OIF4*LHHM\:/"PN2:FLCP>[9
PD?M.['[&!%)!"]N5*GD.4)U0"*M**'B)<1^/*F_9353T/^3DZ<I5 -:NQ-S [<C=
P3'-I4;0W8XT!I:(:I;<%@$U(4EU@KD4H\!Y&1S?0RV?YY'CN@<^I!14[RWT/'HN(
P<M9SZ5RA+-1'HIJ0W $MM^ERSXC,AUG(%L L'Q"IN26@^P]N"/>JC3-*.P*F2>2K
PPG^G+GT.;Z$$[U%K1QF<8"018CUACZ-+2+52R(&B[_%WU7:K6GA8'/:V6LVGP#B2
P+/UE**+,R-NFI+HBO(.1O* 8&%E4$PD';C[$;/*@A+*"DWQK-L#>8V$+6 JJ3F.5
PDW!O?AT@?J/#O*?(.VIV5KV0\P-+& 2[\1)OS\ZE9>K^0*^E0<]:# <098_R:2?@
PTSWJ2BU41"\CAM) !1?6 I\)13W]>6*0_BN:S=HXB8MB?I"NBCXJVX^#5EH%G<Y^
P&,!_]"TCF^9R_<LUN54-N=AT)E[5P,BV$U7K, T)WUHRI^!)JZLH7 H+E\Y<.EO:
PH7;Z6EIS("R,*'UM2*,,1(@_4R@--S\N4;]PC&"M8=-L*G;4$,U\1A*Z%A$<2[?:
PS+JB2BVN@HZ7HF*K01-OIX]KW?W\OUI1F=W4/6W__*(U=1%?$ ;'^1HK)^9'.&E<
P;($R&I@DGF,MZ*TQI%-( 62A34'?IVXX\,<HL,PNN'$;SM0DVE;#KO^"(S]&8J"/
PV7YJ.IHY'!RF 6]C5O6ENA;0<Y$PZJRBD3.$P?HFH:%VG3D[&/HE/(2 @03(;!VH
P^MZ5F&PAYWC:!-O5L-]7^<_LOV]K4+\;RVP#M6)Y!?AEO_1$M.<6\M5KPM]C8Z""
PX71(HF7@EUWOK9ZW\)/ZO0*A?2BAPP\[HXG(B4^GP(QD&/EH?4,O57? ;_&@6%E0
P095(?[9(=?!OG#:DB1-@\J-CWL@^<-!TK3"[%^:A7(<-<_D6XGZ)+*,^VJ;DLA!5
P<=E50Z8GTK#:3DX T=]RQ&)R]K!W->!EC\M;5NBL_"M%N5[[OL:^<0/M[C5EQ_?F
PYRLCJR.'GEM[?D"+F0M!@\*$BN-SQDOI1C'AN$]U;SZM'Q<%_R> !7:,C92K3.&X
PD/2QIMRPQS<4;LP;4&^-^F!Q@QI:1!^+*#)<P 0A3ZE);-\*NY2]IWWD2=L5E?V-
P,#!,/A\*>Y4#M2?ZJY*XJD]]B.FA"1_[CD0K4(]7A>79?&5&='^.6UU<7N==Y9%K
PR-50#@7@$-.ODNRI5I:_2^<R2M?FR^7[,!PR:(ADPS](/_2-6C8HN%E<Y0-$OP@C
P%>:EW>0-Z'E38//#BDU0PG(\B34"1\-OA&*.=*KX>0%8*F0Z'7/R;!Z8SHKS8-W*
P9^MTE9Q*>&-8YFGYUY_90.'+IE0+5(=B->:J-$QCH(U*G.!_@(^JL29V+=(3+F0A
P$,SE;L1GZ>.7#/#,GK.\1R,>]6,;* ?LT%ZI+FI@;1G"<:+L_>KN5()C(#,W ^J@
P >Y+5)QR+,B ,P@.LR'X0=/9S?]%L!L0*ZIA3)E4QU0SVJ&Q3Z_>KC5=V09WLE@#
P__4<VGN*>BTS?'G+/W\ES7@,6C@9[U/L98-/L2\+;FHVD4XSZ&\._T6A<^A0%U@#
PU*;*9-8M755(0K<UU=SL*BBMZ)6\M!M0;L6.$B*FA2UGZFGO0:FJ8 #?P6U>'P0'
P;_$Y+[ABGUW"TL9S3 N1G$+&38#_^S8)&U#C>(YX4B<D/ :XZ]?/..FL=Y1J59B]
P[5:N:E/S?=M=3^M:0@EJ3*8!%H#?1@P,V)K$2Y76PE;WK@_O>:0S)RA\"4VRUHIB
P<#WBZ<0%8W3\%0VRIGJ)8'E"N2#RU&A7.&G*WFDOH. 1XVX<D)NM .OY@;V\Y%I_
P^E:*%D\J<;.@5@QJ"O(JX:]_>#A28D] 4MB\D>:P#QSY  *\U1WE,7$F\MI0&4D"
P:1Z9D[@E C"Z"O&8QY<=[2T8Q/FK6;CE-(/N$_#C_1TY1[=FPN<&\=)P=W9QH@;'
PE6(QA37SOOHE4B[)NJ5U->\(4BT89YP8<086TEYG;*4<!%0]$Y1;>0'Z^.I06CK%
P%#%D0N;2#T=:DG*KKX)Q:TO6CA+\-?[^_'I<->&L,,](!>=>TK@];4.'9XJ^?)<A
P^FB7&_HXL^A+M7U=?G$^'EW9(5(+,8XA>GY.(D7HOJ31X( R3&6[NS.5%E>S79)B
P0C*OP.CVKI-BTXI*(-32;O#T#\'<3L3VNO'=W"+*NXT<%!_#Q)[AV^!@:3;2=H#K
P9*[NE[.&;3V4<1PYMN[KS@>/GD).O%K;Y&&#F[K9*TG<8WA*Z;%V>P0S*VAK="?8
PNGVT $/M64ES^%MUG<ILDU^]U@3A38$F@F_SRESJ0#5Q9%<=,HDJFE,+:V?8?S4\
PIQ('_@:A@NJZNT;4FFZ3?P(D%<.<OQ%[51G,G@70+/7W+N26)GEC+34,E:GD_T92
P&51F(FDH[Z4T_#M&ZU@1@5,]M?VME<>"I=Q".V] #ZHR\^FM4E]]WH7CL7L@!#T'
P0USH7_HVO8B>+ UY.<+2'8_B!U<)7?#E!#USUH0NQJ@%[M.!B'(RL,6O:Y/[TEP8
POB,V\BW%(4#S!&L7QG0=?@Z_,-V0:R]MXW<$)TP\50UD1H>]6^9^D5D^>*4 (A$=
PEPORN<ZO))AMY$F8=K1G'PH.E9K,M+)?Z@> #-B?>!WUO_*?^ 78-":Z$M*B%76%
P@@+6[<78+%&SKEH-ZUTCB..Z!_4.V>G*1IKK<YO?T7(%+#N!>6D!KTF_8ROE;G"Q
PVPCLU"5G9E,6\ZD8PT(Z%4@>'ZY*6;%OW.]V _^]6F44\9\VXSRKBA2WAU8[UH0T
P?C-ZMR?01LU?",J;WJZ$VCS?4]@G=&G6[!EX:>V9D&K!18NLF1)Q/#V.^^A,'G)*
P -OU/L&3-63AS80F<ZG='*/$F;S+-D:#88D92#Z*>J?/'>:R Y;"!@.Q!S9$2E@V
PF(%0R 5SCFKB4!&B/P^(2^MUHJE1?$#^G!?<[* ,))R1L*7KCOS\E*-Z=[Y??RW#
P*S]./P75@P.\(HQP<K^CN@VGXX,026FU$G?0\]$+:5-\W""[;6PQ<-;P (A'Y$-H
P5(->;+"'',!R>!HKQ!I53J[/*CQ;!GB,VN/,LSDV\A(V#B'T+C$E.R$/\@TO<#AC
P5HD2LBO'-'.D;$.)J#'HC#F2I"X"@UQ:HN@H957PTBVM#HP-%O8_":@44*]Q#V/M
P+K";'B8@28,_V*S(:FE(*YZUE9CTSBN;&F N!*=H#JR.MT7X+1,_L&=5-8[1B8#I
P,!FD_=85..> R-I>/)Y_?253Z]>Q^B;9!Z/IUDK4E^]S*38G1(Z:.=[12EZGI&$0
P@VW)NF1[WU1:A/MO!6S1\9G86KP7LHQK!-K1QSWZ.UZPRA*Y%@7-;OG+:Z,B",5.
P7 A+UQ1\M'**ZEG(PIA7L4N$.=.J5VV+DEOY\ Z<)H6C/W3:\=7E:FW,\\V:&Z#X
PB_QPGJ/T(E5$$_9 &_!-92!4S9ZN3<'_[DA[4;+XF"NH^@G][YSK&EI5;HY1\5( 
P2>(%-'/RS>TD.$4D:F*N?:K*F K@'NI/^\39,D62:W_]>T2/Q#3XU&$:U#5V#N'X
P![8@\@!F>-A<)PAF]&3%886VA-I!GZ/J-3J7D6'88=?]*$06QI7F0YO)),S[6$:S
PU$! 4XU9 5UNC#"(K]MXN87T)6]7QQX=TPKZ?\F:TH"':%J'U0799'F6"PR"GB/I
PLYA(D-!]K*VDEPU<DUM0!PDU"+4N3:M'HPXRF*&)5.X> ><)"H2HL,%OZ%2J5X1%
PG169%;'EPC^D&'XC7@DH$1ZR]<8"CL!E9+NF0;D7B/#__&UWY0A#8/5&H+P-T\9F
PA?=>#[_EA[V\YAI$[K_\Z)%E%*$$X74!?."]_T$B ::07;GWD1=:#/JT')=B,F"M
P+11Z5YG:)<6O?S]40%[SYUT:R@1LLK#+0VHS-B8(!9E2W-CE'+4%WK OB!FOIA"5
PR9*R^2Z)U ,6YBL]O;8=6/=<K,&U2>#-!V^/&00S+<!02*->(1QQEPL10G3/=N_3
P41<VK8C_X-=]-DGR3Z-U-TT-=F+L8UF#C\QJ!@.+>.51I#[]=#T14KQG3J<?B2V4
P[]R.BY_P)3)ZN7?!233L6JEB9J9[Z)O0+IMM9G4E[!O>#W9))V8/YC>^<ZA8OV]U
P53T+FGS,\P>89O;DL SAEUCV'F2$<3<]*[;D0Q(@5YBY153B?=E1&8_/668/I^3]
PBB$N=)=_/OV]2;D8[TBJ,R8D\M#S[%M(*@"^3=/S86]ADWZ2&,AU61-!4]&KSLU"
PI?X[7M856?,($;WALS%I/>#>..J%\@=RP1>X$'F,44#H=RH?HG<B>0+\M?G_6>&]
P-<FMQ%,?XE(C[7DX>O%AZ3O<N\$JA7.,]9/Y&T<0=8^M^V.?;31527V1ZHOKA1CM
PN%/-.:6F6%TJLE\G=F869\S9ED149W)DEF;10C>"R%@0%%I<QX228./1<)6>]\N\
P;#QVR"H7I"5Q%7Q>O^BFN* :Q2GZ<H)[^U5D90H&IVWKL]#BU@,*.+VH=*0S5BWF
P<29[ZO\:6.QD,V#DI+[P YE.7NW**+CGUPI]A'*17VR[Q:['^#<V.WT:L^LY-M?<
P4TE75 (;*EG@[Y@.I2+KP8?\KZHR5];8&W/>U41V1VBK[+PGV\H92_4%H7<M-NI"
P#!A>FQ09*70N%0+Y#JU/R164B:C[Y!S:5TF:-,,:)XU5[73;?:6DSR&Y$H=4$@9@
PP6:J0?GPYH@89\HZ,JQ=16JE^89L*H3K]P["MF,!\(1S- TQ##K\FWP'[@&_7.6D
P5",_52#OZW<,AQ*7'> +IZ]Q"=.0'ZCT'+^/$FL\6ARP9!T_CA_ 5H61<IHK8X*;
PHX]E\ICZ90Z7G7R]J?T0YL21L.[2BF)R]1T3(- ]&%]<2HO[K9)\\J\R;1-/IJ#U
PE:FLFO=<E[)>'1AO$?T'EY'2LQ,F/-4.NYV#SH-L9 ?#/1C]"L/S+/>N<E]$'-@D
P)%>A4('AD]B_*Z/&^*5P6QCGS2?S^9 [9_\BCUAM>9OR3K@&Y4 <*^_M['-K8(GX
PWV497\$F3:"$NH</BTD/;UX\L\/=A+O0Y"X4ZO%Q'D/:X\DE5638&=B)F3# (C1(
P(U3$WTSA4G.!CAE5_4:OG/[98D2</#; 8J[?\,A "B)#OUM2D_(,\=&L*V[UV/R2
PZ_,T^ \3DOH L/*NL!X2[V4D9.G<E8<=L:*I]UE1:.Y5W8KCVY-BBRTA:XWD7:<4
PK@M#<5DUZPG-]19<"4L(1SG7J1E!@,3/5T SA?YGM;>7'%)S'"X<]2F$>\+EHY[\
P3[CG2.#Y]8)I"E LR9\&$IJ!9LCC]-RT9':5\6%9UL!#6189Q5WS&?9_#OE)=R]"
P-@(C8XDR[D<HO\<OFC8<Y['-P20J^OPCI*SMX"><10T13!#&LGY?E";OD.,1;8X>
P3*?U\'T4WDS ^I^0JMY<]RBEBU!^2VT>GT#N_VTMD>BW.A))M?3V1E$'-BS(1_Z-
P?1NF]+_">P >TT:*Y2)F[]C6DK8XUY*GC/<$6V;<V2LGV4M8H9MN/"E'^R<0=!,$
PW_1&P92(FJ>#LI2FXBL.+ JTG^6"!0S<%43<(?BP1PS'- IA[I2_-/URV_@-&D@(
P:M6^HJSX?>7NF!G2(MUHU3#LN< K\0XUT\"SUS[/#YS"*%*R GN_F'_)*)\ST0O0
P%-129=P-:;P(NYGU4MR_K&V8R<ZF:K<2=>?;FP8R,+QK">#LD+O\N4B.EVC%SX)D
PH#]MAR]M&@Q!*!5E??(+0CN%S3<5DZX4#VR]Y ,[/I6H/CYW&F,_3H],"'#:H%5F
P4@GB+QB_.+LD]81DPFF!F<<8C_^]U\6T\J3BZ/O;I%51]W@_8A.>DF)I-PG4[1WO
PU=\=9O^^[(!MUBR_O"/(*< 9<OG,R*IDSH2%(<CUV-89IH["4#L+O,JM]&GTT1:^
P[_Y?B;B4 Q_<&*:I% 0<M@5\WCB)M)BL3.LBJHK;$-"655(N&9-,$Q79E^^_!(TX
PDJ+*GC24,E@8K;^*O'40P, L:5,B/@+V^]#YU&O?']\&C/VY_JCIQ&7H:R[K>O?T
P@LS!Z)QYQ9;*=5,6D(1RVX2E8%Q5U3F:"K?#.RVGMJ%(@".\X/]Z'5():<S$M$NB
P',)BHI<RGE>#!DBT4M'>1HZVGXEJ "F=B3Q[[AH$110&JU^K6PS+U-%9/8H_LOM9
P-"8U*, M04%BT#ZO=,&B"Y*I3W)3D^ #[?2PT>,[8V&J>O10BIN,+15]#(KLDA?F
P_&ZU\;]+!N:LDN_0L38,OOD,8$2*PY+R*:S*<0U9"][N->2RYDC$66G^>L8;)*AM
P\&@I\G-17!1*Q2SE/\TX:ZMLQZ3OD?HZE(U9C$MC0/YT2S'QOI^1"/(DR)O>'"@(
P/*&<8I1P?83.%G7CY60$X'X%[5B4\4P*[Z;JLM0D+]L&49>P8B,V$\(OG'Q)^4%,
P@N:0LP>0$4,#*#<6BQT*__-:]0.-B<PW&$9L7]0C9;OHB0O'Z"F,R><:D.,OF_4!
PN!,$X(-7!=\2'H^SD F.H0YT<XB\RNCL0/%")(3AR'2>I29.GV8RG2]N.FSB6/9/
P51"$*K5!4T^<07,H2C$>Z9:AT-Q-UC!+_KGM%AKSO5EL[=?EC'( ANHD<I_I8K$,
P@PV#2JJHY5#O>TB1!GL/8-!%7&1 I333@@E21@C^Q-/'] PNJ3O",99(D>MFS[#8
PML8E)K*!6BDX%. ?0,60XCK=##3 0.>)X[TZV9!T1MS! .YM+B\\#S+8P!<0Y#EY
PUK>1",:X7,)!C%@RW?0YPFB#K%JE=1E^2[79,V--0$#P2.5D-2PT QDB5/DV6K3?
P&GY**#:SNK>=L]L^S'/4P,33T% W+#[^B@,>J8!@ _.[%317Y0F0NHCT@8FJ8R;I
P&UO\DJ7[")!@UL7,0UGEO%H=N]2?_<#.&/[:R80RY5X9RKG(0?OKG*@OM79JG. .
PN3$=S1[WNZXO44FJ5HBACY'P\HY<P?"\X3%P(?8OG2TL2C?)H>W3#,2*;5YV@[5%
P7N,9^(BW^\HW-L(S&0\(\Y]6.!W&!S7RYPJ9*R] >;^<=7$5">_X0U9N22H$JOCY
P/-W^_FVJ5!O%J:DX$:2W6(M%1-BPMR9#M4,- Y;;7&@N1H8&"#KU@5AGX#B($]\6
P2O=Z\PH3K.0EV7-W.! -=ZV+;) B,MC$;I%?(\D/9IV0AQ-_V:V>9Q@_W8,1F?JB
PUJ:/1?=ZS(E)BQM#'M>O=#=R.H;^;I1@Y;_U!^,M\8.53,5VSUR?J@8.Q"M0I=V<
P3.O\GW=M+>4D;H,T?>J'?<Z-P^#;T_ [HG8=]^ZU6=(L>\#XA4B];@(J2$K4&=N,
P;T,_T<449@4X[P?7W\/?I[G'SMD656H9O;'_?M\SO0LPL%V2D'8GSH4SU?B; *PI
PUFNXE SD2-7:5Q.KWD_'IUU">,/9-_!&&N^Z8SS*KY^%US(FND:;+D2IIL'7TWSL
P4.9Y$@ J\Z(:WX5@ZJ.Q/?^=]?:Z5D+,55-T78^R!1^5)?!20YQ9_0-EETS&>"&^
PIB."XMG@'>P*IO7-*C E=J@I=5!XBU#[A,Y2'_9_Q>1M4%2@!WC/6OB<'1:[--D:
P-.QEIO]==D1P\O)7%MV-97_Q53F@FYM=4P#-M.^(R%J))]E)]B"@,"OMM$4J]G(#
P8]Z\#\VY4J6U/F83BMT+[ DI>5F>XJ9C0XX2X4SD&?%/6^U.IBDC:JH#&MAK*<*K
PD8.UMQD4(5V[TFH3 7Q+7FXFD4D(&M-:W$,<VT>E=4+$N>M\SB]J\'X5FH:E'TI5
P'FO12+>&785&;UR;71H[AE(99W.Y&0'1S"["]8"CN%04M\CDG=8$P^RK]B<K@BUU
P)*GO0.@<[],4GMT;"\]=07;17O#GM8_<,,*_))3:$R*AI APXV9J<-KSK)?ISU9_
PZLLQJ*]/MB@_P!06UB=(JJ9/.>+R&!B0_WY0^FOP?$TYME?1->WBQ=/AK)!7R3_?
PLAY6T6?E=(.8GZQ,:!9($D>L2$$PC'E,F,=5)C,[Y.K8OWQM;PN[-KH8RQE65(_ 
PD_5$%?$W\<C>'C:S,NM>FC !N:PNH23K/[]GF:&&%[<3&D4MP3A1,Q 6@/?9=I! 
PAYDC&MQ(<'QIC3*;R,T$0\@K6?T)..O*R"1XO]=^"=D!9\>:TY*;N&OYX_P#8D/_
P4_YG6+&33L9=Z%B%\_8.]J9/KJ=JU*;JY]J3CV6N;PN$>@/SEFZ'=[TS2N/\@!MP
PZ%[ZIS-9@QJVY/R=C\)6*K"";YC9\L(4.$HJUO"WZPZ,\,L0N(B;S$#K^2?Y?XNP
PF#X6"@D_0H4:U1>C3)$L^9=IP5J+QFTL>C7$J/\YDP9[HX*]UW%$#VSH>G%SW,O<
PV_4=6!HP]I+GQ9F#1L<%4S4/:9AE?-X'H1%!N23&!^K1$&_0!4S8*C>P28_8.MXE
P<R ;9XFV'=D;KH(YU?)=*%Y"PM(X(CQVPBO;VBU!B36DDT,24W;L\E;TQRG:%K$'
PE^TG;U@AQ*B"E!1A2'+1?BS=]UWD\B\+\NC/X7+.&BY#?VM].LOMZ>>. '^+IOP'
P>\,SCY!"E.ME=(><[Y)<N5F#B06\$IEU99VI?;[6KC,:I)./P(*VM;IDEU_G)'C+
P?UBR0=V=(M(_B>9,/'X7;"0Q+4/#/]>HA-/QGRI]JD81=O;<6<_8G;.$@UNLVF7O
PE@Y0]9#55.\*0& ='>M [WF<"=8^-N\!11CK!K**I4I#M<1T,BJ^&YRYBW#Q-I&\
P)N *N6I%P5$4B85*6JS<*X=);+KK*\47-X ,2H/?:?2,D*<W^%SM%C8UH]$F %?9
P:):&&8H$++W[5_&1,AP)]61Z2231)6[A7=Y&TD7CV*7U=K  5%D8V[,2[]!!MB-?
P[+HS/"!L3'JJF):9CC2]O7*O3X,4]7MUBLSM_[5ID-Y?AM:3UN8**@NR$L<-X@G\
PQ6<41^1+CG)\K$,9,1_N\9()2OTOE")%Y--56=*!%A,QO-[]VYP;\2^-J0LB23&2
P23P'6-L7AN&X>CP T7G2<JUF:$$=PHX6B)[=SV78IMS9)JQU>@S)5*O_E$5A4[JA
PP8X%,><6DA>DNHFA4;93A !MQ!1-0V8>:BL!FJOY!6"W,'F+76\R.Z7YE1>F:=*V
PW]/JMGF*AN6%5RXG?B*\_6V]%>/3ZSO+*PJZT'0&:>/PA')<F7]HFXH1=LRT]N8U
P9Y%'LZ?[H_?EP\<(RJDTDZ/(U;K-2JX/CTD>P;7^DO;Q9-<SR[>VDH/1UUBE:/H@
P3'0#42W*?RSM^RM>7P6I%#_I /0,:$X]M^N7J=E<%&)DY:9%+%]7=F]+P2OE4NL(
PKJV,J9I*OR@AG*C)S3^#Y?)RE]< \67FY/%X0Z8030;'K5)F#Y4Q<IW@'6VX63I%
P<R'@9^-;D\#6?&.@[)9CBUYB\=Y7/4=3V\CB;1 *\%/YM1<67V='E1@6MK@VBZ"G
P$,M F1(DH96:MBPIGYW1D /2645J/3+]C39\E\_NOGG=N46!4KFPA71? KI!9%K3
PBO,#4X.5\N\9S:]DKA:ZP)SE#S^F#GP%J'P:C7W6FY;37@>_;K+H/LK@R6;R9 05
PM4V7!XR2(T"TK;VR^&(7JIWLIX0<*?\:P2Q0#<R78#?6'5GDYPE.FN1VRJMUP6QQ
PQS04XDKSI]VZ)XTR28P42??2P>YX,:4Q>MT(!1V:YVQD7>A'$HVS_71T%(HI,M!H
PDIWF*$B\J6"L=A(Q-;U4;2:7C" L#>"<$+//1EESH$:2GJ+^WLX^FW@0IJ]2V4CQ
P]F8ZK3ME'&"&$-K7D6[I"ZJFT0)9R&/U9MTCK3URGV&;R]!S*7O]@G#OLG3Z)=C%
P7]!SO/1CT/^&I!T8B]UA]W;"YV80%0EXHUEC?]%79:H)+DN$BTHOM$G:^$ ,*7$O
PF%)JN_!WGH4)P YX)S(_$*BG7FE_8EXR>'&V&V*$H\60V4"F[Q!,=TGN=W<,X]^Z
P*:)V6_ RB#L&)7N_>O=Y$7H]H&HC<#>YE)??9VUA9'17!THY%.'!JMDWLM-8:3!W
P'"E2VX28(]+N;+!!]*"\B>MH6,(0_2T_0ISB=J!585 ?\J 3$"Q6QMAF7KE2/RT[
P@MV9T=.U-%G'%$;84/L@-KP(6>%[T]9!0?5"^?Q<&M<W4[V\'O)P\3AC"ORT075H
PK<Y?70I//&->?SK>ZXCPL Q _QOC83_KI N2(Y"U3FJ.>YB]O-OPS"L,IYW[=C^A
P>?IB24\9G"5[=,X\(Y1E1<U@7_@AZF%7:8=LW3Q9JY=D+*$Q%]/DGR-,&:4::!JW
PHBER4OJN\JW]UP.U*_?K=%\3=4J:IZ3>R??:.\R-2J[S9)/VN/<B*<(_ASSHFDJ6
PXW##(94&!748;Q[\4TI'+PGA]#L_O^_V,\ISHC1FE=53'Q)\^;_J6^D^=L:<=N22
P\*_SBK<$3:=:/!SSLOULSP;KK-SZAXQ,U9/!TCT7%P3&-SA$50L8I6#6O5AQO':3
P$)WW/K)@6#9E!BJSF6"G).+MKS MB7^2J\:'[<[./I+$<34(>G- 5:S70PV7 .HR
P9[^G*BB0AF'"7.K.(<''=%"D8W#*G9U%QZ9OKTU%*W+$ $-IK2N4W6),'!=;:VC+
P+=N=I^A\E R)8GAT=A&XCDU(%B?TT9-Q4&:)R[JFLDM4K;^5VV2H3UT*[QHBFZP,
P/,J@IR'?5Q3:X9 6I6#1<I5E([@Y>GK8DG,.4,9'BI[ OM\V?9*_&@]3W$-)::_3
PT3D3P%9Z%_SN;4.D<;80JK(?;U]2@N#V8*:#78:3"?R[\:,-A6%"?4;+50(B:L9(
P]LIS)IYKF93U7$_ IQ>H?/,)MBQJ&BVRH52UAUZVY2 XU=;R2_1C@U]?L%+&2$++
P$< #OT;.BRG&;SF(S/ +-?^DH39DCG2_HZ):D4EBK%6P7NP^JWWJ88CK]5>P_T)9
P@R=PTR1X8#'H_8\]5D;%YJTTJ'%*Z:-EP7/70)11H[W&:#8<_H9R%]EE1*-7J-]A
PIRD<C-U>%4/<,DZS]C5\=.(40G1L_51<83X1CT(\!TKKT_"WQKJPD 7$HRH.O1P5
PQ,X\>5Y!KB0YIF#Y1=QF_Y<^\ZE03NCAPM25? 6@RA;0OT9:Z_<.;1<4Z''KS,\"
PV"-C#L=;96F7>@A2<J*@^--V5ZP,0\Y0)8*BYFKCIIH<SNK>4\-C)J>5BFB% RQ]
P()3G:[B*CN8UB=JZ3Q/!3]I #9VD4[!$CLXG-;88Z7XOZ)(S72/CB%P7Y8(U:F3I
P?/).&VC,8?W%/XHI,,!80+@X\A\]*8$8B#"U/9ZJILI"&B$3E.4"T3TY0F\=Y&#R
PKQ9CD2./V5^AW=F8:U2HXWY:ADDN3*&5]XLZT(7TB(CGG), CDBA6W&"XZPN)J?*
P"5SX)_/6$=%FO^E>^XDLKBD68Y-?S$50YFV*PF^^_K<#_S41-%"?.:Q$8.4DGUY'
P]Z=MIAU#/ E)36=X-S[+?M!G")^!:HZ&%N-4]HS$82(GI! M8 W1#I\:M;D(W,1V
P'OG9$.)9Y'M,2'2YE"X&J;:#5%< &W/?<("JK<O+N'4X?C&0:&:L2!_L?)6[!)U*
PC$90+3[JGFZ#9137W '"ZHE?,>(4ABTUTA+-I"W<-J* O;33'?DZ>-V"+=NH2(39
P3MPP\%S![LOE=+_64!3J5ROS3-X0XR<7^+]YO4PG29<_/\5,>8'88&JQ"MM$XSZE
P+7G&RU76$JC'"R+WPP_"=O&DJ7^.C0D!(?%ENLIGWGLCH^&?/RAF]YQ<1RF'9^JD
P'\_7B5KK9IK_BEYWZE4FAN8<#":T*/62;B_"ZJ?L 89&>,27O8W%3;M=?H-7/MZE
P/!HMU4 ^'4)B$'^8ZC:H3IR2$7V>-]'W6ZS%./=0A\I!]&7PUR7@4;SJ86J8-7O.
PKPJV,_$N5WYKBQ872=B\Q19+;2O-8[K]W_P29>+[077&>19,I$Q_Y=93@9.O8"A8
P3&1!M=@'IQW% BWL$#+<^\[_TLE76:%15JGO035QXVE& J#G9$4HY(2"J,GV/VE 
P?1[+5H<7!?F>\N,AAM2CNE^IU6F/7YA]#>O)6V1)5;2;0[6U6_N!%O7K;JM\MC2<
PUVG7Q4P(W3-!2<UYBO7+-YSRADE<3;SKLH.)ANHQ"%+!_[M"'QNB XNONFI63,'H
P1-Z%IN$M_\R]K7@EC=Y#WA:$A/\C4F Z]_,1]O\NART +>^N-L\M?Z$'(Y$RN\%V
PP%0KH0#]5%A'CN7:[_:%0*K*KW0+C3+T(W087</(TYG(9%&%:RNGG,,@V9QJB'&X
P^1]DN48R8E&JX_2)S&^%A!0E^YJ% /ZF!?JVZR?1JINE/0LN&(R*U2];9SLG6C"U
PLDGY<:)EA/?7K27>',Z;$.4,X"8MVCV0WRCGX#*9AF0#*&FPK8SG8>K#=,U%SQ3!
PV\:##8RNEL+*B[#C<N@9P?39%*#Q4;B&Z)9AQ(3"7#%=2U&KBI7FZW'-<81*2YE<
P:ZRILUDEE7+K^<")#*,M_>M#]^>:&[E1%T@5?\(?8M>CH?X>:E"FTRR.WL][)\Z$
P%H3^^*?0=%6WHL%_QDWYX)U#?<_3>G\@O4R,H%$-=_Q:5XT<7T'[AE3MUC0_^I7'
P$VF2P-$.WPXZ-EH[0E&K6; 9>&ILC[/C&LQH2.81*3B;32J_A#%2(EA@$$(##_*+
P]TIA)<^(^Z$!1BL?$^,W[%)L+AZS65)Y9)!Q6(\>%P9T#<8(!)[*A B,Y<G9:_MN
P0)_./$<@8VA3$496T0IE5H&^Q!QPL4;RGJCN^8'DC0&5-BEIII'SMINL3QY+O.G!
P*Y1X]-MTUAKO=\!+\B8X05*I?&6GU&J-IH4&!'ATY*U]7 I@;T341H,X7.%S_+&Z
PJF$#H:87 :"LVICGY6H]&#_<"-S?<:ZI%0D'$X&#+OF#Z^!!N.UJ;NB?3"?^/M)%
P7X/BD>G^,T$*$1ZT=3,Q+JAF"\SE]5)/I-]@IP,_7<=O/9,XMO"GA7JP28 $@#=<
PE^@U%>%(>K.V2X&6L_14M7(Z>Y:ZAC#XEO*O:"UKKZV(A"U/>@DQGE\C26/T9H97
P4E)ISJ3C788D.02,XK%H27M5!0=FTT\\>@RA;/=**T:AB>]MN!#*Q<DYJWXS^=Y/
P7"[B1!BHO4CI*U=O&KEB=B1I1<,R>1:%@>%I'9\1*Q*^DN/62Y1R/&85\=(ED"<\
P[6F3E4-F!J+M7L)5[X>5ORC0K^7HK  @,I/JPU09H=OVG2$8YE,'YK"TUA@E6-6'
P&:Q%/U.91O31]W>9Z:F'+Z\SK.1C)#FRS?++TO1/]<S6-,'_P_,*?+-45U!#P8=2
P!UT/],IC$X==44M ?S6,-!K6P^J-S!PJ3BO"A1KFV#(:'#L8KZZZP+%K''^7;1I=
P6T;>>]QKL\+@RIY?FK';RABT5 @&P*M;9DL:'6(I.3O@L;N)_69]CY^2MOIKF3>*
P&_6<,1'7F&\0H5A_8(YK^-WCS,#,-B^2P8^H=$9NG!94-X4S/"$MSD0X:)=TIO0/
P1$=&'O,YN).D_9NPXL(H/NVO_'1H?UD-/,% :8260K%Z7:M;"W=L6X,ZNU%Z"6^8
PUS-%6R6-91[*4#RJ/1T3]% Z&/$<$W2LYF(2-G_0LQ\MU7';-45SZ$KEWG5#J;9"
PP'E'%T7&)BR_,.T+62#IW,E-\&C1IT-+M5)ZD9JH?>\*>(>Z!+,_/X98@%@S1ANP
PJCIOI\O7+^%J"DN-=+>+^"Q%"Z:AK"+!O6:5:,\G0=#?DBJ(1-9(W_1HJ0O&*SQ 
P//^>7K/F@&2'CVDSGB;31Z,UU?K&JJ9;+^KH<Q:U[O'(VQLU ]6IVN YPDSDK?Z%
P,1SV-_)AP46X^^+VXC5&Y?:I>^Q1(3/H")T!%S:G$[1H6IZA@V\F\TH.\2%L I&\
P"% T[7!J-TC^&8EJ>U]IC25)Y5LUH\-8Z3</$2KO3&GO#,T'J?IEJ"?-]3RA9XWE
PW^\ZP/,Z8]E!!V4G>Q7S#U>_&TO)J>XG>1G=(G%]E.K@RC,$DDYV83R[HA=0=9>,
PNB_3W',\-.9!$>P?S%SJV161=ZXTUS/4W$7KTW%X]TP6NH)RMVK%03()%J 8G-KR
P[+H*X[02K&CB>FLI )HROR<S88]9#1EPU1L4CTMW^/'&+W--7M%-:8H'!%IS][GO
P<X<7D<@P'H6\N='9.5>[:U[46H YJBPH_RN0F:AFAT1H@7,026O/Q=OE*US@PL@N
P;BFXL13CJ AE-PI==KHN\0ULM#.,G'@O?SIN6)[X&U0U?!T$"D8@F0.\V6>G01:6
PG:LS!V E8&ISD;C_I>4)&1GUPW6'4I'O98*M+"/O/H4;U7OJ];20XU(W$SRKCAK\
PYM4-GW+349L)"U:-]WL"3E&5;4YI_4[ZO"8YG=,CP&&##1M,2>1F+016U[,9/&O6
P0J) RSC1#*4#<<""/=#[BSYGDPVO2#0P5MW*>1!%Y[AJ:AGYMT(K-UD:)/J3B=*R
PGB8F!;&WV",QH9^E[KR0MA.NA*G=7%\H<AW$>WCM!W9D:QGDR5J_83)_UO?&KEDM
P9@>N_^4//JI%]O$\*4"I]$@#[=MP5L#KK/ST6#)L<BFAT0%=T9<E!,VK\U5XYBI<
P.,[TAT6#HA<HW37H62Y,[SIBW7R!F'HZI>$2%JSSC9T;2RJ%?[))GO7T*A \:N-;
PXP9D@<2X&G,E*,Z8I4]#YWMN>= HGQ[= D2,'#H5G)"PRGI-BY^&4.5O&Y-N&9F<
P>D@S)-1OI88U ,O'[P!]94!@@S(U")J7]*%)B_Y(\Z8HG&I-8@]$<#1@?T6R&#S*
PL9C J4;J2:(.U7\U;9/*6:=0]T0'E]<]L+J:OI,VF]4XZ. AI1R8Q/P6#N/%IOI@
P/@G?+LH'YMRE,;DU2F'18?W"/^84>J>CXB:R^%?9 "S3=SC<Z34Q4R! I\;5'WJN
P#$*WV1\L"]_JB,;._8?8'29PUX_[V6MI7_00V*":'YCA<1+>8B<M'!!1W&6U>[\_
P4^97<PPL1(.AR/=W7JLV!Z>I#%>YPSCH:DF<E]#4 P799JG]SD+WT674"]H*8^&/
P*B=.@:5J#;X^1/;["F<P&(Z3)V31WALV@GTP8W:W+U NNUR70MB_)_B3R/Y$A_<M
PF3*\#<F^*%5+<R#@)R#V WK, Z+]*0@$RS'GH\_CV=W87O%:$QE3W<)+EZ;:-<'!
PF6L/!>/[C>8S)@U?(LIW*:&YW6;_&:_PL:]'GQN6/6C=-+UQV/Q%CBP7[T<[)![P
P3.NX!;^UXW8SC&[$Q(25R8<;"3+%,9VKAH$VHSM_UF[N>\ZC+U@JEP&[)6J]G./Q
PYN__8$"J>%4UGA^YG/9J.(@85B-70ZV1/SY!*WK5"U+_UP/?W[;C:7B"7:')JU.\
P +4.@ 7,.^K_Z^N/:*79FN0TGU.@]M4Q+MP9>PCH(>@H2JTRHED&\7>S(Q@B<M#K
PH(^'AX;N<O+682%4W&<ZC/GPCANH4P'R$#+#$N(8>#FP2-N!CKL?O]R'?9C/>Y!\
P53TEK>2#&R'&G@%^YU-Y7<RE\8-]C<=:T-H99[&G8ZL:6BG?AWX$_F=>)D?,037&
PF;71M]?%GC<C/R_J8D1B:4N <. 6^RK^)L;/B=4K!,7> %-!RYVSEBF8*+ISZ;;W
PHV@U8FPWFAIJ7(A&D6Y^T"VXFGXB7NV!08,>*VR_(,=X]@'$WBR0#(P;RN*\:+A_
PC%-3"S/\QD6;GB@/C&;FATD V%]633?R).[5=2)&%J27GRX4P:6:7%U4 K2F_%I 
P6DN;HG7B>VON/!Z0_9XK)TG1PO;%+-IS<\FMR2!"(F;1%;)=,P/Q8Q7F1F%/WJFT
P!=Z/I'V5-;PQND^EBK/ 3^%FWY,)5;IX#/_[_'9<1F%9O=;',OL,E7CWZ3_9+#'1
P>?JJN3S8J?S!Y,35ALQ?J/9/D:A6-H0J0!= ,\/$(*Q5;L,ZO!.,FNONP5!#>ME^
PZ%2@/>9\=3D/#M:H9C0WPVT(ZO\DVF$R85NZR(HJDNDMTE>?S3< W3! 2X!IV8J1
PGW0M\GX>^!8""34Q.TR0+;SLUGVQ.SOFVJXQUM[-,UX.#KV/X>QK;*B:CZ0<H!_A
P.JFK:DV1VW!N5O*>V-!Q2,0C\ ?4]2JQZDE+TU'0R6YF3%^KHO<JWI&?I(]2I&Z2
P7SSN"P5$+F0I:FX@$6C4J8^6@EV4,_MQP'&=_6L74%!@$6ID3S5F30EO A2\]4^)
PTV2_&T?!&?G;A<&V1KSG=_L:LAZB7L3IE"D,=\)N<DJ86RW!?H<2X;SRZ03=Z>,!
P(T<%QJRJ5_0TV%##Y-H5'Q?:9+@'$$PFXXX^Y%9G%/VI<W"5[ERJ+/9P8Y&-JF&8
P6"3#TBO=>MG%HT;8D.W_S5AM^A44Y79(\U8L.KL<\L:R"-O)^I@;5 1#MD@S#<#0
PJI(H[%>7'$>2HATZ;51;@[5M3XE3B1Q?MM%=SET)VGS;U07?#1 NTNW "J"-SGDT
PL?MCB\D)XEU":= 3/@;:&4Y]0/9P*Z<ST:FBY0J<R-A(!8O^]0>C^G:,&/B9(Z (
PSFVBH1E]F@#[O>QO;,DF$*IXOT)I==?5RYZ59-G1*6#O,=:>(7,#E2?-]:@,@EM8
P6HRP0=:Z1)0 9F3%S&(@QBS9U_*/N2ZNE/"ABY*-<=3;8LM5<$=KZHC]3U)Z7,S]
P>V,E99S )(!AWIO1U75?_V>>@X!V/>,NUQ)!)D?F$IUE;&L^M:JJO*;#IY*3#_IL
PP\>F@.'(O6A$C/>)0ST7!."NMJ8T&>QA#*N"OYMO9'HN_OEGMUKZ<#8P6+8%9'/]
P.J3GC$?Z[T^.4'_.EOL"<D;. LF+*S-2*S/!8W_S(1=@O!GAC%W&4-_UC#LYJ2H9
PR4YA^0#0BVE6"D'O/0=2 5N>,Q-2H5(+A@V\S]"H0P9*PVM&PW/M.:X'>VQY#$4S
P<T!L@?SU89:2SV<@<(WFDXK':S?2K?ZJ@$Y[0O)EZ[>&ZL&+UJJ2I12>&,I^G;"V
P'S8WEY,J.)"]7&7X/0+6I.82O @UQKV5)^#KZ.("S'_CZ:\KJ#AIKA$E=L&D&KR5
PKVR3AP+C.,IR*8S8-<66IC4T,(;\-6*N>SFR\KGZS#J<A#C0CF$$_U9@T\.%:A[:
P>F,HH8>LFX8A(U\MD<4L02:-?AW&#=(7&Q#@$&K+.CV'"-2*%EZN9M,+I:V:38\$
PO?/9/"FF>>KFQ^P\H25J(=A3Z4ORV/\198WV/[J.1*_5L 9'*X1]0UFJW1/ZM]Y8
PWZ[F%9 I]QR6:2]>/ Z\5Y)!9<CSZS.L& '5&_/X7^ 2AOOSP&\PG>X>%!]39,&Z
P)'L84<B>,D):'D<&?B-Z3V&W\[\-0$4N*C2*4R<-OHX:)9%/@(:] 8BQE]>JTTRZ
P";DCTB[Q"H4Q$[#0J&[L/,9 \7S/8-@'.?,I,0,O\C51--W*V/7G&@K<IW07'D_/
PIX'H+7I2ULR7=]"P(CN;4=21][:]1E"S*%&0!UG+ 454,*KRZD5?OB1QX?R3RF,V
P&NE>[[H]JY%.! H:+8ACO*D)Q<%W4S:5<Y^#(N>*S]\%'3=_FX$IWGHV*RJ>\9Y!
PB8(I30;4@1=)EG+UFB0 ^&@6*=8X>$1>4%B)/--DI&,6KH4@7,)S_!$J%YT.95.9
PH9*N6<K'2U$$T5WB^ZG@,3WRVR9,H%R [)-;(IJ(V87S^Y4%22E=E==H)2<T>)CA
PX-T.W4K4*'>P(7&"5$1:42"9BZ*[-U,.G1S-/Z'M<L_>T&?(G_B.JN-WIVLO\Z5 
PAU?T*QC[&QD)6LER%:A@>DL$Y(B1@&\M3"FSZ[6W'I,#BF(..\I$ZNV9+B"A^2S5
PR4K;0E*V=1YW&'8VN[9"+P1)6W$!1+"B+I-LGOS[^_H://M+^ IJBP02YY6_W.^/
PX!"L<*Q[7H+!R=JC<_;-R2C@O B)%40.C:LK;8. "+^2OJ(*$N2&Y]7S(\1@2W]#
P^L*5K$;SV$*N7H0-& S%H=Y:2T/6+118"--R[.82$52- T!0X^H.-C61I\*^P8SJ
P--^: E$2$S_%+U?3K'IOO35EJ>4Y*EIG2,CI)4R=+G7191 %M;]!H')2*0L3S\F]
P';0(H2HX?R 4Y.Z2LFY?-P0;Z4J/B[*4(!V#2DZX*_TTSX-O7AU,J0)V Z]3@$K]
P,G4 F8:,K!.J;%=H/A?G\Q;=7W,LOTYON"VYPX:YQQ<...IN<<8Z8;:W%\M]#@KQ
P84A45@2<R%7I%S]O@WC@B^<'+B&8LRQ0:K-L<Y\B[MI4P4A3^^,. R8'@V5<@7*^
PLE[9ZQFPW3&51  [(5G[W*UDBS28*"^KG[=QW:T3\,(R21H$)]G<J;%H1 3H.:UR
P2EO>^Q#5)_N@TY+SW03\S(^JP:F4M&^W1<U@>S:\9Y!Q7+W!Y0[SG1*C0[0SFA[R
P;$98@)RQ91H_Y)89PH MGGK,W1AI9,V\?LUOZ.9U\!L\*'D?T*MBGJ>-WT/Q5LV-
P(E+ <Y#L_.VZMJR01P?.7\"]&.5+B)'\/5<!+KRBA-<$OQZ"<',F20\1<7MOFB:E
P*=9?:S_J"#7RS.DS'S>&&B+(67[)O!#.K]%F./XJ4HP\J A"LJJ,GY9[60%=UYWU
PY:+&%U$TRP%;.!MJ*M#7^8D>8=NZR-=VFV]=]BR^JZ-+-75]9P?6W98\;PRSTKOR
P.QLJ1,:=6UWO$R15#LH>[8!$ ,'R%);ZNX*<Q^=2N]HBG>2<W^R[%R41_8123NLJ
P3GL:E8D,(I8=DU/YK5<QP+5/@+W7$F"A@G,/76T= <@G14N)R+ %OA):2!G6C17E
P9M&%]#!A^Q"?&I1<GWO4PD=I3%%PQFFV5&A]]I962$<-Y=9KV^B,/)%7WU$:J+5O
P%K(%MQ90H24="!$:IIASVQ9(-,AL_:J,Q 4&0SS'\SJ#F?#>.[H3LJ',O#67,_@R
P-EV973,J]VV%'EM)!RZ4 T^/=Y8..VKE46+-W32E$A8NW<:E))"VTO=*LD^#\YT'
PMGU:0CNS:EO\/*-\NE1AOB>7'C9O1E%.<^2&P92  'SV45>[U+D"$8N#U?@V3#)Q
P-EUUAA4N,M&M7B^+<FT?!229YI BEP*=BX,(SX1F4OS6EA_G( V:$6%F_SFM_66R
PV;3+""-H"-TDE%O5&AZ#!R5 3G"\^ *S0DVRJP)SSGP4\<BH&$U,*U2/]2_O]Z"@
P 9MWT5?S@H6_0TAYK=CRA+:/1LVV;HU&Y; L"_,%YE.N*,DF) A.Z6X,A_(]V6L.
P"] 2_@0P]%O.-'_GC>IW(?CC)GP9W!%)SMPG CZ7L2Y(#(%*R]M'/8*QY)I#=AC8
P]S9%C@ZO'\&$'5TI60?:-(TO/V- 5Z2N[=V[W3<?[2$FFQ8NFED&%=+NCT&0&G()
POL6];KN'%!J+MUD*C?4FO3Q4G%"KX4OTH9G=MQ1^VX]>O"GYJEWEJ!=2 KI90H(K
PI_ 27Z('T<2,<1T:W61TB+3W<RD>ZS>\'X!X)HH\9=$*H74/O3RYN0$TZX!FDA:-
PQP08P5<1.@R5<OP1SG:YZJ.\%0V]1"\91E%-_O/D@DR+C9QR3 ++X@)+W3Y,IFN/
PN+*7K=<XRM?QPY,EQBL?%PA\&(5>Z?. 7<PA03_J:5MA;K<SI D/KR@D^EBRT0)4
P:!\K]@EK.:P+78Y,VN>F_CY_OIWYRIDPR2G@4==V;+->).KX@C>ZZ*$KYNR1#NH!
PYH/#C $C]_I)V?W9IE1J5X185#/:*NID?"K'GY@-[7!OEY*9GV#1(X.%J8I985@'
PQEX5\,^0M%O406/^N;2EUGD.[9A]$IPF>Q@B.3!0Q)+.FONN1;P6]B7GWR@ YCHX
PF4-?^W@QS@]41J4CZ5!)5[U)0RD..#?&JQYS\%2]LKJ!+EG!^"'O\PCDHAC5JS4&
P?9( ?OQ YANG6"FK.; YM48EA!BQ&JB"8UZRUN]Y#(M7BX4R)V]HTS\N-Q3O7A8O
P&.CB9E[K:NR0<A!ET9X%0%\B9 2B;FZ.$&-FK4:JD\"@Z:VO#>8J7+UT%XCJB(Y+
P0\)A"?1H50SX $=OF%0)R 0 )FZYQO H&7B  H(F5MUQD3;VMHJ4;FK ]:_KL 8S
P%QHY+73QK\:<M%>BA'H$4.1/0F51^Y4RU"P..O#%_&."JN^%G<)C-B=C=71K^-A*
PJAL,$/_UXFL6"V);<]F?N:"2P,M>:H#B/^<?[L*H"\2/P>#V2J]-B^Y414^R!%5 
P(<%VQ^:JBNY4G^LHR6+*MRM[.R^+2W,Q&EJL:)_JK6C073@VHZ^X5H"U,/S2[BWW
PHD.C_@(I6)%NM4DNY7&7F<K1P:01C:+^].WMW;PT8V1I%17?"89"J.2QN-[AM$$\
P</"B823W9P/#9%T$7#39<<DOD- =$(H+):/F$(S!#8F=T>VA+U*7PX[ZXA+H*F2?
P>L,TO@U1A*&G[ Z6AC&$!A8SIH+1IA%H@16W&Q;3DK*( E6LO>(YXR7_W7XMC":1
PG:2=#!(0P%N.-^A"*K-@EMS BV*8CYU\)I.2Q0GI4/A&)24<!H6K&A7R(6/9$[.$
P?&HYGP_X\+" J-Z6O1UMVQ3/08(.BZZZ1-B ^UGZ^99]:H?*50_K-< _@0X]/O,%
P'8P( H$= O4<M. MZ6XJR3+CPX4:JS0(LT8*87PE#-9(G!U/77*9"E,/O_$'0<>.
P9GB<?':)FTC!*P_>0=@ !-//BQ\GLX79>4@V&4;?07"Y(;^Z51(RK',DW"M/.,W4
PD4*R(VBF;P9Y14+="\),,H*3>4"1"4.$]=7YKBL]CJ<,7&J3 A\<O4A@.> Z&7O[
P4%C8Q(U]J2[,^Z@[@W;L1395THZ&0Y5!FBW+7]RT'V^NG62M?!.)X-^[BH9=7FIN
PSWXGJ^./S 9OQR[(/>FO-S<:!DV1)%ZC(J&K>*/ABTX5"C]*<K8)?*/6"\@9L!+9
PPLK_*M4[TQ.C,>^T2P(]KB?Y$ZZ/3R_?.5#.]0J$5]"8^1%L=0T_.C^'46!^4OE/
P58=:N"S!/=S(&<W=KD27@0?I=RP767Y2AS6+-0U.B,8' :>L"WR L/4/["%P"SS 
P;5&%F1$*\[\"Q287*9]&B$R<Q&WH@2N@?8E\JWHX)(!Y!HW<Y]!U,"VR+5B<$M&U
P"!GBB%5:>:$9D;Y]ZUXI2W.518?. 3=P@/'7_$UH36,L<1M_I;+Q1DQQM*M$OAPV
P2*^M)Q<YG=^4H8V-E<;^84]V!%\[T%H7TK8;L24+I[QJJ5MR?2XBMW0&*=5J692*
P<%8P@ X)QS4EH.;M8A D$;**7"56BWH!%IN<-&$R$<7&07J=EQLY23D56N')7&'B
P)GL>@6XR,4TGPWR)1DZYX_V+#PZB.<8HS+(+H3Z$$[XK[=[IO7-B98(X%@V&<AL.
P*4A\2I'/O0%O=EZ"?^E><00W_Q^VF:=QMX59'8O$,5&DZ?_%N5$\;$X^;>(2HZDE
PA#788L^>LYW72<K<#GC5O[K]_-KLZCPQ3[;4R,TW$L2O%TIFR<P)MBQ1]'F_SR B
P3064\+?!>)1N?@IVAK3-/<94JBC[@G&!S23$H)3I^&!$I8TA#OT:G<:.N[B9E<?0
PYN[ 51YO!%B<0)O9YG5&U;GP<LI])_WC3]Z%(I\PKR7:;%>%?"@0SH.V^6H]Y5_,
PJ-EK5TO#I%@Z((6KDC4YW;7^P)%T_\4>B&X.9DYV!TT,B5>T=^=*=!#)'F'6:Z?-
PSTMU;M_/KFPY5[(FLU@ G\VAYXO @1';E^#*--*D;,C7)M9CG,RM]1W,YS!,E^<!
P^7#QZ;&YB^#-0LP7IT+%V@NMXZ 7N\:1,.)M\60.DHC%S3 $@\^4B.?<QO&*./TA
P]O%KC;;X0SFY[]J[I*=((F -[5LZ<Q09>'I_9:5U-^?<3?;8:KTES8Z ^W<(AM% 
PW'%_8>%<E9[7K9:XF?%P7@""%?>MR<843?N(_8^SRWCC) ?"*3*H?WX"S^FQ]GW4
PW\.=BRF-L2?\7TSGHB#E3\> *#/@\)K:RM:K*:[P2?)P_QMRNH/:4=[F*Y7U;)E7
PBB1NOSU^H_5YSVKG58?TU/'2-#%<HJW\X:.XBNK/CD@<NXRIC.QD/"R #!B58+PP
PYBJGXF-M%_LFHMK%=AZB0GG8;+:D]CVGB($8RGG^B%O1C7@Q;_J(I+@U2?LW)66(
P>U+3;G:M6XW[*:)W'EQL=OJ6UY$"7,V)D2>5?%]071Z[/^,'OJ];@1)Y_5Y&M!=(
P(X1(VZ/?$Q'J,NW4[^?C)#Y51=^6P^I"7:&D3FY6RQ*34-)<=<!<Z))!@3D!'7QJ
PHM2P@F[]EZ8ZA-M$FI[FA&853K4'%JU<KJS0.J!-IS<6W[ZY+Y2ILJ32UAAQI#F^
PZ>*+Z0'VU<..#F #!*C1O^]BA=F IV^GPVKZ[LDK%Q%K*3ZAI^/FK_Q)[^1:3Q?_
P<YO\*07CF-!Q ,-3P]X4""E^KN]CW+A+1_8'4G^J/O$@;TX<_H 3/-)JY]HL6Q)$
P>,3A QWONI)8E&S-(&HG5\&!*1HQF_C8TE#3*_.TGWNEK7 \+J1 O&08G+HA%"N_
PY*7HTN.?)) A$NS#28M]@Y6L'\>N4@ #T<!+?0E&['9(IP$KW=GA8NFY'%N O0WX
P3A\CA+H!?ZV'_-60VS :Z2$&'%9:4_-_5^CB2V&-/7-8&1]FD79I\E]\7OROE]<_
P*(20%0\%]_#W@JEJ$*6$"M1RA.8AK@=PWF9<>0Y/H[;=%$?[&H\-ZI<J#LQZN$*A
P(&;VX [/+>.&1)@M$Y,C(F/,X7JB70KA>:AE+/O /UY&IEXS<KG94Q@(@*QSITON
P^5JTA8S?2O\.;<][<AGX9T3%91>.R\[/;%/=T0Q#EQ&DRMX<[/@P ;B>.Z"VZU5I
PL_;H2Y:LFB8# _4ILP0Y9BH;(HD1X&1Q#1CV;XGQ#5+T[+O\DY*RL;/FY:GDCNZB
P<04WXTI7%IN;3[DE+!I-/Z*?!%4W- $@'>X]M TS6"GM WZ:N=MP80)V9X^06PDL
PR$*=4_R;J4\J!#@^W:BO!:I"R#'N7.X'*OCKM:E(^R:TS=)_72EQ\9*//<44W7$%
P9UEUF#I2(ZF"WT&@?$6>(+?L+@E)=@ B.\;)&#UI-,1)H)68"<8S4D#<NYDWR+87
PG):A5-Z^W_<:7/G0!*=3J![);35<?LVR:2=R:/ 5)V5:J+3,H#/6_3*E:O#@)5K>
P:UM<]5^&DHYD(M,R -,0SK1M>;1M0LYR%;VK"AM?C&S_ZH_A[,KZ?+\G\W9KIZ[ 
P/%;9M<=?VZD3SK0QQY7>\!PD.27J+W>PM(;M0."1]-1YEY_69H$V/_=XH[#KQ$G5
P#^[S8RTL&6%[59EFQ\JP.K%\4P-L&"4IN- ZK,10/<Y)(1MF@IT9M"GMN])/W#2-
PQ3=II2;<]O /1--,IP4IAG4N(6%:^CMSV27E'2I\?-5IRTDE=C<W6S2C9&],;W8Z
P^:CC[N^P*LHXD1X3,!Z.XG'Q"QD1'Y<'+[^'L7QR".!H7%,9!P:D]<^CD$H9WE@:
P[V=(D'/'<7'7JC)NN;$?[;Q8038S,1,U)DJO N4,HP.'NI*YP[V]%\@]M>6# 56<
P8&GN?G$*>S'O!*%]( !1&%X&M:JG#%AQNIB6DQ*"HXRV0=!HN_QQ0VK(N!Z/&YU:
PZ^R/)'0$]PE,@H]KQ.E_'!)^DZ= H)381*S2"CU#@UQWI?[$W&1I&+"$U6F-21I0
P"@RJRZCTS<B:2M17+42Y\H0T=54@@A![37#&!9-#J !\:TTI\QH' T FDDS. "@$
PNW5N*)?H+[$)>2Q<VI;8-*7N64I-?VHE6_I*JOB@ FA&S0K6O&/]PQ?T1LYFQ<LK
P9J1_H_YU</<Y O@/K=GZ;)0Z3FA?U'.R^U18MUQX?.?![10C0!YU>7PX/,&FY+-%
PLLFI,CB0G1)Y6;L<=V+>5S29A\V#!I5MU4E,4/J99SY?4@&*(2',!\,O:0'<Q<&\
P6S"<KRF&?R>MX5)*-I 94-\8#H8*: C/!['[I6/_Y;=&IQB&,J29?-X=FF0)K<[\
P;*)LQ8)FY3%/Q7"+R5== Q2"8J#95:Z_=]*:-*,0^PO9A4O/Q,T%H(4&3I">>'JP
PGAM[U>W;7&&\#OI):YR?J"Y0TV::TBYVRSS6[.SBH+&=,J=\U=S\A&WHKF/[(CRP
PL\OTBXIS!#_ 9D_.A/5OY]$^[0"!5?AZ%4(X*3S3'^W=2)55M\"YII=U<-T^W<Q.
PF7QVCSN_1=.1CA) S\H5?D-BKGJ$15^!:<V;K7%R*G!W'KO?=LL%\TXZNOFTD&\3
PI?13_TRDF=1B+438A3BS*&.6NS"KX5Q09]=[1LM,#NP"Y!K8ST0A[UE4^FXV)L,4
P\;?^FKZ&)])/\FAS[]D\9;13!5]V5;$I_X4 \)&+#CSH"RG2)ZOI #EZ<.H\S:=S
PNB3(]YWZ=79_!B8[G,^R1VE)X"K6%7,*)NH>T2_W=N7GMAAT!X2\GN<7U4;_?5$^
P^_$S(VN\C3NQ*J@F;5<Y8(Y21! WWB:7O4"H!^A52BV"8@%<9R\<B+D!?UZ:03FF
PM>"1F%3?JOL_Z3B9S[[// ^W#D_B%UZ86IHK'%"#/[LLCG,:7-"(M(HS>)+J3Q[H
P6?K?89S45]AU-*S;^+93R>9=L-//['-\E,)%?WEUVI4]_;+RY$N@?B_2X>SE,9M=
PF7]-1AG)3BIU!450FU%RB,;F<]K9PUB0)TG(>.=82"SR\VW45J_L)G7Y^;,AY8 3
P %,VVR;/&*.;KS^UZ,H%Z6NAJZ;$%\4!WY)M#GL?>PSA=>?*754?>H:J[[GMB+B,
P>'@T_9H\_C>']K!7DXQ!"?&)R*3X;$00F0O"=O:YJ-Z1PBM$R9$E"/:.K@\)\?97
PS5X+RJO_0#Q+ZQ6K$P%")-0>:/B:V!?_EC\P'(\R=9_Z%.Q#O\?96$3:!!\(9H#3
P?D:BM54]030O8W163?S(687V; &_PN99N=\<0>(U=+]W3Y=3@Y*ORPWIM(I8/T9'
P-IL$@=8\MKR0];\\-9PG=![4'/08Y]MT6)8!C<!](]J)#<QZC#X+L(L_X)0SHD2F
PI<63D>:+SOV'ROYMLF_YP<]5W0?G6E#_2AWO!%7K9L@A>@9_F#BP$559WU%SIF"5
PR.%HMU+'89@81:Z4UMI09LKX\RM8F^U/"N&H,@AHQB*? CC<Y?8D$'+UXKO9I-O>
P_V=1,F"Y(^)5HIFN+7LY?)1CW U_.&4:246>S2L%G]+]2VGJ[2F&HUSS3E* ^!8P
P><7G]:( [B33SXF_9M^MI^.XPE0U<G_2%VB@U[W*OSX#.0RM"N67[/6!Y-%M2U65
P%V>J4WQZRZM0&%(6(WG>;:%_N4$6VW1; ()!']>!'6'AC;%6=Q(F U*RZ9?JBJD?
PP/9A ]U#;(]5,:2BU%I?D1C$Z\06E?V<%I:J$[JMU "RXM(Q,\N[;$O2 ^ #6QCL
PP>(DZW%69RGPZT,S"2-A'!6C21NH-<#QAUK0^XY%389,,*Q=IRLO^]EEEX7 0P>"
P- %C]54L( YU,*_"FD]1T:$]I$)$"4%(?D._3MIE/^F<U_\>6^G/?@RI7!/H[!RL
P4(F-K+]["55L)'6?"/!2Q9EQ)B,U54,FO\,+#C&#/$_3[Q&U:0!4Q^?W&=&KBTK'
P$<"9KK7H>(^F ^! 6N/6)E UG)%T&C4U/M)@8^2Z1S(ZX(%:@ZQ&PV$U7_N<:IX*
PWJ .Z<I>)TX3=(2;J!2I<;KN[^='"!(.I'UMZB9N2K\:7$FWNEXT_GT=GL>MZ->5
PAU)XIU]B1TQLK*-G][E9*8&6@0\_7&P3_<7<Y9 MM%UE25RO"45?AB6.!N61]Y&[
P29HUA^GIU_G/VRP,QYJ.!?>PAK5I$..#,!X[R80)%>%>C?F %9@X<_W*/R@] )H0
PXBZ)%U2,V;%,$E.M+,/HDNP'B$KA6C_>L#UC^CT[M<O@ER@H!2B$10^[3BAIDNW1
PR!WMD8*FBM7\=KIPZYWIWB,,C$XKM)M>E\$+>WPGH01@:OG%@=M9F4[ >/L+K\%W
PRG7R7-"/N6(O(,"N&H]=;]+XWXXH=7L#ECX MRGC'=QZ9Z5Y^/)8SVRA#?^A-3_J
P =#B0CP=JQ5*&K]F%RMZQ&B1_OQ_[3K=1YK=>R^CKX[0[^1U(20L48M"IQ8OZ,H(
P\*D# 0R5 L<['7_5L09?9=QN1([!-DZ4HQM3J@FYXC.LD;N^\W$*/F90W*6U((>E
PK! !9(C S7VZBL*U=C)&'C_[^95JV4L$4 !&-79L2;.9/AE6;>LZ(Y'R/;J.]2K%
P0? ZW=6-ZB-Y'Q9[IG+=WJ-J2\R15?\V5W[XMY1&]L.Q161R(P#=@#K.#76O.*_<
P1Z=FD1-O5\@2O]K&VB9K=F.$*E>4Z\8S1\U<<X6(PC,XMS-@@7G\1N<O4X6S1+*I
P5.M>UKP8%U.:!T??&:)S.UR)AQ"=:G0IIOZK6=O^, JWWI!>;CT4%OBC:""\IP'Y
P*O0/KLH!-'SF9*)T:[<+)L6;=LH=W#<G75+:)?:UF;G_@C998<EO9,4GEZ,R2V Y
P0@CV>S].8:@V=\/X%>$D!@5QJN[44R9WK^CK;D<3,SWJ=\_A@(7$'S"%TY3'U!*5
PT9>R!.C@R%$9\29,NE$LD\/!^.!I0]!=%P=FEG!2[QNSEVQ6-N+(4P:]ZH7%T;*3
P;%^3__WS.MDP@!^OANTE'EI 3R])2>5??AL3H_U9<#J5<PB^3.>RN$S# RQ'!M*"
PI/@/9).I(]([#I<VBX<3F^5__5=_P,$Z9?Z-R)9F &>R3-:%R.ON=-^*_&,^5*V 
PFBE(/H#T359T82>AHV"T1$S"1 #Z&3D^>J9<Z@9264MS4$2Y'0@:3HD3<I_T7"$O
PG&<A0M[?B)^]M!)0J6%%C,V9W1DD--P0\CBB)<V/:C@/R<."YCR;QYC_],UU-PQ 
P1X2Z?@O\"+>:K'Y.)J2@IGW@7(B.+3[)+09$. $45MZC\XDPMM .(BM?0L^1G3//
P,+<Z+[PE,+NU,(!M9%.-8GZ(.==0E4+$;W'S?@+N,N:56%WO(+A'OEW2200:RK;2
P(%^'1\9;&'<SC<15G-Z]5S/P:C)"^U4L>FCPF_^,A>(::LQ3&)AR34:-'@!\6KH4
P@)PI#P-8-"$./B\3A6=<!7-JU&LRLF3SZ4O5,AE\9[).2'4T-'B(-9G/#*;MR&@.
P$-BSU=3"=$\$()N_5DWT>AS.E[,/6RR>P]-1LDP0O(8V*&'H711K?4%B9?7S#&$=
P.C&C3TR<8:A,FB4IL!2;:O%Q2A2#8N+HQ1BBDC\]="11W)_&,$O!VJ&PP7S9'X_*
P?Q^<RAYX6KYD;Q5IVHE@B$&2>L5ZI9Z2)K"!YSG_(-N#FQ& ZATA/K@(=9XBQXJ/
PP07O6%E(>&D!,Z_*/$0H718*';;4(SO8@\4]6\;*-PTU<K;Z#X]K2'!$'=-I+I85
P]*S1-/@[UHO7/<,@5C4<18O&D=LSN\R3K-N7V>)I6!H#3'?DQ%&*K]IZP'S+S'W5
P\Z]O0>B['35:>3BCZX$F*:/7T[PC)(X#I  AJ=86X\N/PJ,%$BUO#YF*OL2E.CM_
P$1NPBRAN_T] 7_GG=JCAU7;%GY9]JM0%2=&!S53E <(8TC*EX-XFS+E-W/N/6-M0
PPC3*@ KD5$=\0#7_CCUX(;;$/^DB<G$!1_M$Y-$KI9=^#:N*DSRD%3I,Q?6<+8C.
PZ$Y=EES=!O0>/KHF:^:#:4%;WO5)5-ZX53R&B2]A(M\< X5U" LYBMF)C8GNP2HG
P%:O[P<7+#+P&]O68EZ[S*OL!6QK<GSYZDN' SPC0O?ZGBFK[?/Y473W ]K1["=Q1
P4LO!$BYR ND8!$L3Q5'T*,)51#J>6.Z13.]TV2L:3[62PU81%NI.GZ7"7=76^X)N
PG$.6DH[8CIJ4"?9=FGNZ:X?+6';L(A._XF1#$-.V=<+$U,W4E?R]=8)\'X7Q.>8Z
PYOWB4(-Y]ZS9+7\GG/$>2%!G)^;?X:$A9]KJ8B=%-L/&"<#.S0G4H"+D:<%&-Y3C
P]O\ZR"JE4]ICE$<0%ZAHA+!FW#*ZFPD+YO'GO\4@3;K%]U?]YST:4V0X!W__W:,W
P;QNH6%&E0>INU+\CIFO:WKO-WW];T)(!)(K(+Y"!40R)IUM2S0K0R[* $,L4BOW/
P8)XA>HR?NJ0@D O5PP$/_3@-84-O)&^9]F-DFP&3?BIVA:M?\;95JE"945L5(9H8
P'8E(1T[U654W4C[0-/C%-3?WZWB%-E-\DS5,#'U,']N:!-CX/_=V[?\#T25[G)/M
PS%1?)PPFCDB-]#YNB'X:ASA2R-P?[?D"775,/7!$2=TIZ;T'QVS2291/>[&@'GOB
P^MNW2O.X52-;\>AV]IJ"',H^RKS%H6AP3EG1+BR:]'P8FA$**NDG)[,T;#F;R7Q]
PKM1CK"EQ$,O\.>IU[*^$(= ,<_F0OK;"^OG"GQ?E8>G-9[CNR?DIK$I:0?U&6MV0
PH%5ZRJYQ^K>B]9SP<CC6>Y?@AF@B5M.R0:7%RZ$RR3JVM/P__V/LOLMV=BI(Y%X0
PH-RBMNFLM!G9,;S.H0QD@O_PEY9VU2S[IGX1ZVFB,7.2O;FU)N0)H\%*H&I;7Q"%
P@&2Z!Y[K8R7U*)T(#?PUR98L/\#D740HDBP%RU1P^*UE?5;V9O [X*T4ZCJ]\6U!
P3 S8^+.;NZ3&H"(P+&G,U]B#&8[WA&KY<@%EYWS)FHR>7WK+D X]^S!7WF[8IOQY
PXA"DOD1&9+22ND_F/J)7)4HX<;QS&[:/A*/^_P%G^@\DUP.B\3B72SF):A*C=LW2
P7$3S.<N3SMEK*B)O"TK.%=5)IH[GXVA,*N@PYS2$GZJ3179^BGJ'.\B\1, -7<R\
P&P[ZJ8M1">#Q^%./402Q>'@1<X"3EZIP>J1=&@A9;?5*$L/CA<!/;.CLL?EA:5(5
PM:9)R1/RUQM"L<\F'Z[I,YR9V%,_)49#'9:V3PL1"EDJ4R)>R87.]J5BC\!M'1Z;
P\94#!S32R>@\WRVQU4[+JM>?Y!2Z\".<:C&A1B)2;C Y;#CB)1"MK$.$@(JJ9H"9
P-G#-]]XL3'<+\(Y(^!>?CF)7W8RUT.U(4,W^YSM48.9\!&_U6X72 #KJ0#5J,[<7
P!N,4V@!"U&+-M<;_*Q%<KP,=&-##&V@HR(;A05F0]F^44E@0F":&^_WW-%U>87(F
P9WZ#CK#-789]) 6N*?+[\F=4L2YL3:$?K1E%.*WO1!V5;=6J4JO=G8Y2M3),QWDL
P(WX>DX^B<?*)=>!Q_)M0IF\*88JP10FK$?\$2:6R?#/AC_!P",!#K2)R.'#6BKVF
P%*"'*JS/S_ZU!1U108G3C[N+)*BZV!&9"$^>)@EO##TF] %9U2LP;!,-/@+$;#+Q
P4($5&4,N+?I!3_!<I))V5(:W3/SNRS/\5OTN_':A)%XVU)]'!AF@]V]J"QZ]I*H_
P2#[=]P1Z&&-\F<;5*#[AJA-](Q76B=MOGZ<Z,=!GC\]X?B#/=P\I7VUQ>.ZJ^=":
PUPU6H.3IT\)=:9MLM::Z2K>6W'(.>%G,).7=&\Q^O]C1NB\)5V%E4"FI.A>.;!9J
P]^)N L"Y( &O3 YP_8Q:PH._;3[]M,FDH+&S29\QC78F9!4/_HN1X;8F,ZW/(IOC
P$"+1U7*ZV+!QE2?1!3WG@[N*:+Z;6(ZF(M!D'1S--/+T;)>R"_7NL,;/*;1$_#8<
PY6SM1#OEZ@=RM\&WD$BL? PK1EAE"1?RJ8BZ2:[2P&WY8%+MRA/D0)VA&5,L\TC!
P1%>UG&F[+\,P"S5<#'? N+?Q1^U/"RV06W-QN_7LCJW=5W+09#=_>AA<^,NV&ZXI
P0C5'^>9%[)"4!D8('%1I*7YL6UWH1R_P^&J :KBKLK5?XMV?25^S,5HUDGA_TDKK
P-Q5\GT4GL[*-.1*U:3\^YWS=77U  L*:C8RT*T6)P%<&8W5):4XOPRVGF@&JD<E!
PHB]!QI/!_/Z,!Y*!:\1,'\B%QCG--^;@7O56J/ EU+D8WLD$\79<MTZE<?KR\RJ'
PV,#PDBE-4T>3.-<;6R1916T=?T:*W'8!X]"?#S]8\TC1@-FH5C=Y_=8XH<?A;_@R
PN69O/W4^$<WIOC^!IVV$BF+C9?BZFG3J*%_:^MEVP?$M[Z,>IUYP?##]&8@_P^\2
PK#]+/>;G/3 P]WA/$"ST6YYVN%.DBJEG!('?&0(W\KM@5/QLNQ*] Y)5U/L^RO&A
P87;RA+B'L@QIJN849K+U&HN_DE]=3*35DBJMJ0CUUM"F+\\EZ<Q7![/#%,*3MQ4>
P3==N\IJ=2<TZ4G)&BE.<NZ94['$]W;PU55O[6#7A7,X;S1LS@(67?3:S5;\XG4+I
P5;,$;^OST[73AS)&XD5-$6%E8YHXO61?IKKWH&:%8$!?5@6T1IZFW/G'P8H.7[+:
PQ7W3+GNPX7/=LZ:G2NM>(*6L2LP=VO]?$HM-3TC.!'I5;6<."?'N#&PHP-OI\]WJ
PWS.:2G @,.1,O;T2747^QFIT9Z%]>3$Q:-$_V-&4.^?V4B(AH6AF/AJC5NA;\\7_
P/(".0;Q+GM4[M,!J)27*:+"QRB[G\:F1W?R9^H1AX!XE/O,4"TTZC72"S<I:K:L>
P2,74^LS]S&>_IP(2_ISN Q0!=ZDDT>=\G3Z-56 'HS&(+QTU?*SD3F=UK!#\<1H0
PH*O^;^^S]Y9,:^O>KN>/I N?>]+R?:*]M!DVZ9>->YMX*B/SN(BSL"J>BA6"@)CJ
P3PSK;QO'ON!V2_W CD)T=7H*\L*.:/K&GM47"P9Y BG+ZXSH65RT/"P_*CUTC:"E
P[M&*VY$]"K"N%7.@;6]IW6@J1Z"5#O[XSS074I--=QMO&4TE[DGVFS\S('H-?ZH?
P#24$U7'FG.Q7:W0JV[.6^^PM+V,?<5C<O+?J4V5=R#JP@G0\00N8%](;0F3\S\=Y
P+5X^C-OVHN?!;DJSY730+_H'1/<J;C'C],W3_GBW!LP-&[UN1DG_QJL\?QC86#*J
P [#&M63A^D!LDR)9]'^OS6ZUI0=?,M64HM()JP9*<^EP&4Z<<T@>NOQ\[>P85:$&
P'#9=NK0U2_@3!.P5:1][AL3(K&^O9P=PYW]0/ZKUF =)._4Q6XDB%S7* &PK6AMT
P3X,[H:"3:\.#B%B]S;:B-C%$A"6;?1134YB5(B:VR9<BY$K.1Y10"=I:.JFDGA2P
P5PH-_:[?7ZB#D)NV6DK81.E/O7,XN.F:RFAGW-N#RTA%34+5((]9'>RU82C@;WK?
P?13!Q&@KRQGM_\DU14E>?ZUT_61R\2%['2MXFEOY3L(.D*G6E&Q!@>IS7R:$]$<F
PLW;ZTS<CGI4:#K'1XCY\.YU\-5$0] .F1/=(54^D6NGHQXO&!'-;!_?]$@S*,--N
P\'#7L)^XPQ+TU#\;K^?I\J9#&M_NT@^H-;GL$JWY:D1;;JK?7[RGFT8_R-">)[9:
PT<L&6O%;,J4ZM?7/N:H@V!9*Y 1*^U3FV-#G[_S%39@(*]9-1F>GD:TC*!00!T>M
P7M"#5\=6-3; NIRT%IF?-4O$D&9FEU74J15;4IP; 0<]>+T"7PW0&$>X^+CM$_3;
PUX.M++^74YTLZL6K+BT<,Q4W@9*PXF4IXZ&57W_.FFM^&Q.L_' 7]4 KL4-6JM'U
P^_E*O'=?:J;$N@!!QLXC'@E8<LXC4\UY$&:T?ZX=*A/3A,V[RSZ:#!2@'(M#D24?
PY<.TPQ>(/20N%VB7#2[F^NMY[<3MXPDI(!W/5/+&(FDSN_%CLSJA&C+T-P9E.,]D
P[O_XQ2Y7) _WR*5^SV930M^15>B?]_.-A/$A+ &N9$PW8ZNGRV'LOA*4_N2\4,C;
PV<T<VM4 /1I29YEY:'$AJ0?AGEX&3K@#IB#5DR%"$-:&\ F#UK?76_FNQT)8QU:<
P/$P&.76,Q@E0\8<(95)'TI6KVG' W3(G<I@::8:@!C[ N0;_4>ITK'(^)NV1'A)-
PL*]MIV#!$2'_2C2PA#^'+E7L]"ND'%G^0%/])L=3T>X1+?8Q;V*@G\_&Z9#(3CGJ
P2,)+7W4SOUANO\-@1SWVG?Y_9\N2UB30DT9EL^\\P*L<F1_3J;R.TC@QU; JM(*[
P&&10L/'-)X; JRLT+H>%VD*'5-N8/M+P;_OJ?1@H %@P1<G]!1J"23Q6&<T&5^+'
P=M,TEOT=. =)ZUYJV\RF7):;]IG>VK7.;&)JR*%EQJ=]8"[L1&9YB_6B;%1/-8ZY
P-K6S8M\W)F. X8D;8BT CV^*S9L?J^.!?-VVIT-,<E?Y.4O>]3$8-E@H_]J2A;\G
PR1-1E_9QSQ2^#>PF),; 08Y; GWKI0MAE\8\-6'V;G=DF\OQ$>JH^!H)OQV3;]Y<
PA/U,\FT04U-/V N^5% 40 LE8$:;3HT.RL/H I7X3?\!8V$^I?*TRJ_;R-\!5=@!
PSY(K24J[[B&#"LAG+VRYH[;!J?FDU6;@\I-HB?__+Q\G(97 YN=-#,2YYI#Z,+^H
P /C2$-ENO?9/DBE/OC[; %,X[V1,[^P*%["#6KA[J3V^W; Z?Y6OV=UR.' H@J6?
PEN5?2*++R^OE]F4O4N!D5-.'%U)IA(Z=T_C?Y7U>!0E7:(-D=?"'WVPG2BU0H:4#
PE5*(:@A2 LN@;&=$R>D].++'XL:8]K&Q<+0E00%*L+_WM^, A7RF-+S-LX/[2I;'
PV(OCDEP_U!GRG([KI52;$B@?].EMW^(%39S96:96>%WX8''$_'I"M]9,OQY?ZV)=
P'\@PJ+.*RAT<IM7]7*HOLA)<W3NB9,0_6PK$6Q/YNU'ITGQLVW1MKYQ'N*\<TAJ'
PH1=7N?'\3-4F[BZ3!28N8,/_C3URGN0CW:=<(00/.F0-)#$*44@[[[$1"Z#O0S2/
P[*X$8G^YC272WG47GNHT:C8VU2PK9X"8U6($X#/+@C.#6D=>?'PX*7[()KL/G8%I
PT%E5=I\A3<%:(L:-B)1=/?1[-<A%J%>-JS2CLMEF RK&)DV0W6,FF; 4UW/[4Q$+
PZ$^^%C*WI\/\NFD(6^USK9=;,(Y^ND&ZAN%ZD2G6R$LD1$_@I<0.PR7PSL6#-S[D
P;<"49)_E^D[R(G3;6Z)EC*_&RYUFL;6CE2E]M_:'I1%!:$8>'-56?!7J2B)M];3H
PL%;CH=SH2(8X0!)R4K\W)1+AL >] W<5BE\OT(X*@UDC481+'+P$IO#LT!]4A:]9
P.%7^"[<]#+2=^GBMYJ930N#Q%NL18&&"E]_[C=4HR76"-_VII$!B.MB$D'Z0HR;@
P@P JDL/:>OJU$GMF\1:)IOSN0V#LC03B%SC=/73KW6OZGIE&W:W[BD#WO37]#WK*
P5>R$2/283/Q^W@%VC3ZT5*^=@^S2W($4+VC%#V9"A'> 3,=(I*^$GKT*?9;]AX8E
PH$&W4]K\G#?(.OM23PF4484_ ZRI<NHP(7,/-?$" 7!ZWCR7+)1;Q[1O Y>KD_5K
PD^=.K$8IU4P67: "=KK+C'Y1OYE.1.SS<0M0[/>NP>6]9.L\B8HZ1;F5&'3;4E[4
P&/TN])NH,!SI1;41\-X.LW7C>) RGCAI9$?EDO[B<>MR0ELCE<R&;$/KPN?R!IYZ
PP2EN?+^_E$(3W* K+924(]<_[TL)GTR-2(@E9$D(%/XY-1%1)8&B@<ANQ[5U57C&
PJ-/$);$0PI.(;VE#WKDZ&BP&R%B)^;$C@:M)>H9>_Q'90281H0M)_&*W?1P WR7S
P-32\F:2HZH15"?1OM72AGA)R%5_([/N)2# <=0KN BMUH>&5+O*^"6DEL"*#UI/E
P O;!W)<1%FG/7M#S$]94<+NKF&"9KIN\=;\C]1R.E_$QH2LTY]_EA^OU88+YP#*<
P(9[+V?\9S^MKPQ,PX.D!WA\#&\/VD<6 @6EAF?JU4*7(U9WH0HL[=*>KY;S]8+-R
P IB"P10SESI$-&GATYACKWP5NS3*NP\JX/7;>'(P G5;:);C%-)B+#'O:C&47% 1
P@/T[8B/-9VNK*W8\&J[IGER**NYTXP> U!16-\YJ5?'1I,33-GUL[B$SRHWBA?=7
P?5H D?C:F+@!5P[5/QY&3I\I+>EH"G&PT:#*K8?;&,W(Q)E *3OO;;1SCT_BWQTC
PZ4^ M19"SX+/..L-^/[S^ L5[Y*E[69+;'X =@G\L>9//@^@;E(N"006JT*A 0G!
PQQCJYO!IEH[0!]@XVK44-H!PGXQ/_<RCQC0.77?"6'!)()GCQ3)&X:6@RVM01 >,
PM:>SG&K<*&*Y ?I=@>G3NM/ZI;OO?Q&$91@D:0)/(:^!UGQ$>/_K]JYD2]ACM+W\
P55UD4)ULD*-(,U*JPNM?Y*FT>HM,#4:657,B I" %^/,MT>^C^71,BQ1<?HC G\B
P$R?(&-48,]U>N4N% 5+2O',=+=;*C?*B#B3>39AD/$-LP7XJ S=09HB]+,BI<?F-
P1^F[]?8U?=2'::81PW]G37^&('&>/;-UM7]ZRY5"@Z F+*[<+*KZLBBT?/GHMIHJ
PS?#;Q^3TX-@P@_*K5SY.%=;A4QW:L68+2G0,@Z%L.]F1:YO*M+\BIK?(@:H<]<[*
P_VT=)GI"3*??BC*18.RT-@R23\I]!\;?[(V*V! ?'8IVCQ"I!X"Y9 ==.C'*J[#I
P^7OG(U^(PJUE+SB"1' %Z(]$Q G-WGI&+E9NC9\C+1-1OP(<<>O?Q;6#F>^!47,V
PZWMA^+XF!W<E-'L?;4_KM1J7\1>"Z0H3R@8_DLC39@J\L(\_ *'2@40EP>T!HQY$
PTLBUZ*O'#YW) 40P;X>8F2G]^Q)$*,$O,E]#*@;8F'Q*%G2BN.['-AOP9HA$EN^"
PI:>>-(.E-U)-[@\<.7:&R>7\(JMPZ1-GDZK9BLXHLO(.4"^T*3;,ACPTM(J_[284
P:5>^@47<*MH4#EW@:/PHDDRMX#G8R@5W^UK^&Q+ $N8^@DKZPQ&PLT^'Q>N14@+\
PDC_V 0"0]X";U$N$1S3_LX+_>$"*BPTS*MD8VIA0V1]"PZ*8J*KS3NNC.ZM-S8.Q
P@3)C$,ZCLXQ<MWM_NX>R9X_>_N-2WBM^^XHE!7&3-#7'S SJL$D;K4D'@!X!78SJ
PBFT6?;!"[;'VX/WR'X.D[9-@%0LSG:7HSJ%#DM%:WV>FUV&,/E3&&I^C5.=40ITL
P\5#0M8:[I\O[;V(L]?K>[^C$^HCS V_EBVE3@^ZFP4.N4RR,(/:Q]P'=3K5E11,*
PQS%OK_,>NCO;4ARZ+$J"L[45T@SSQ5!(T!1NZQ)1&D/F8DY[)Y:\=KAP[FQ-OXH%
PF<P1+&D>+F\]INA.I]/.%X0135HZ!7H-VE8.S9++M:NP?RR''C;W<YXQ"-3',=:M
P?ACQ"9.&9^+AEWBC\EU>6>3A((-;8\=-7Y27T=,NB6I?X!6E+[9)8I'XS1QXKY1+
P<^_VM:$+^G:.9HX)('9ZTQ0\%++]^M89]4]2L'Y$0+DJ!5'@"9>3)/,)AS8^+5@,
P;8AX4O2.H>]"6@7BCR4#4,3![_VM>OEG]=-5^=@2K*G3%8-B,0J9*+4 *UOV.]-G
PQAY]+D6^WLA;:Y+N,<$4-U[%>MI\YT"1).W<Z0'_:XM_S\U7Q7(:[F"=%\=9E*V4
P9\C9'=(F.;RF_!D. $7Y)]]U<57$1/("NER.:$B37IH->T4TK+-V5<P .F?%DMSD
PP-UOS_ N@59!8YR!5(B>?DXZ(CCK;JP$$\D;U3R?Z#A57E2&9!#S+9^W17?=OL-]
P]WV6#:.ILEJL&#?T6#.NC8VE4JH)V-6W*(7$';:=SF=X+/T994E[_7K#28^!F07.
P--@B#<,UVDR&IH1&=*00R$ 96V)&GE>2FC4]^A?8%)MQ>.5]45.- 8GV,_Y[B#'"
PI+K;P>I (Z<V4(5[<!F^P+DM8(@?JXS9KQ1*)BI-LBEXT4GN'E0J +:V*@EP/*40
PV@L&N] (E4)<>5Y!] P)AF]ABL[<%K=5LIYQL*4]GZG\HK-%B'2'%PGC/))UK]V0
PP_F+<R^=O 8R!B90F-PP:@6X9M<DA+B2.RWY&6I4/G))G@+KR$R==JOU YC3?T_S
P'L!YI>55$6C6<$UFZ!$O>$O#-24E$HF]_QZ7(5:C5T7;K0;&B<<%2HH9FA[R@7$,
PND?Z<<S FXP3ZAO;Q#%42#W..!7$7Y-=JZV+G.MR;'+-K8MMRU;O!$\VU%]UY\>7
P^W)U046"?887<VTTMMK/R?GG/6ZO]O\WB9U;^  #/@)3C,\EJL-AR225?[!-9Y8I
PZA_\%7&+]I ?@'_DV6<DC2!ID4L#:+$MAL&E_,"@;/9^@Q7'W(*_VE-HI.2$:L5@
P$UXFC>01^(GOON# ;U!@!4ETVYY<"_N/SF0,ZOY 7'F\,HM-7FE61X= 1!DK[0 :
PEL[BC[OZ3TZ"(^ULO<5GL*9F"FCH=_5%2?W&P.^02CN*M%1 \9A\)8%)=B?BP?KY
P@R+<6T#+["!_OZAS7VM\JN,.JJ6G)3[*2KKTA9O).H] [*WK#O;):Y@>T.$F=QW@
PAO)"4=;06P]X8Q'([+ELX ?B_L*A=PCFWXPPT0#=_VQ47FA-T_+_+/VVH:O)8C+2
P9"@A3!@62%; $8;5#+NJEEBZ38<UVEDAS?#Z3@4Z_[8 O^R\(^N$4G\KQJ1_QK#H
P^UHF*+!HEI2!2K.3MKP^_2*&C?*U6F&YFD?"0\U6P+?'J=B5U^_+&Q!JMZ)#W7@,
PBT%:*^1X+0+L:)-CFSB+@I=(WD2:\PM,)==C\:>:88,?ECT,./R+H4VI&JW>U"CG
P^+L &%I)]Q_T>T-3H]K,\+<KO-J8KIT0 #*9#2RDX/.(@=?5\FKMS/#$'X/9>J51
P]V!\OLF4Z^5O=E^_WUR0JRBY'<*VW%_;^1 20F\]!8=;.5):!5(L?[LJ4FOG^? $
PH5F^S>?S8XH7-1O"CVG/2KUD\ZOS[ SB WA-^C_A?^LGC#A0\,NQ,)SP*TA2MBS@
PDN5<F^)X%S/SS5AR72].N._WE96#.O^)!:(K5'><'%[00\FRD:OE _J=-$22-);.
PP.@92XK5AVV"<]&XJM$4S3%T>?/WF I)\$ ]?]8_2W'4D]>SJUK %L $E3R9LYD)
PE#*_DOBZFGQ=.&KFX58A5/U6R^D"<\HP%GLO>J;&)#H*P@FGFB2%Z*2QUUCI6QF3
PWC<KA V8FJ-C%O_%UL6D?#K-7SNDT+"C$R9-#'RWB=/EA5L\,*^-H;&(;7GB7@#;
PFO<<$<\)H==0^ORXB+RMZ\/C?/^75=5/3&QA81H6-'VNI=<&)AEP 2\F"_RE5%>9
PHY@0>@AR](5PQL;Y%1!%6,Q(Z^$Q$I]FV)VR4DS+_ #QP@$RM+,D._4OO#<:9P>3
P2XUS88:L+ZW@B?K-$VC';1=,TZYNCXU%T':\+[=]KY&K3^&P3S+OE6++60-I8CD^
P #B7ET]GQ7DKV=/7+EIMM@;].M;V5F5?BJ'#4LDZC2B,A^NKVH&W2N0%&Y,ZYP$?
P+$=3"VZD:)$;PI\F2D"Q0XR'TE&W!"2_<G_5E HHF@&775W-14:!VM1WI6Z7>W@(
PU9[AF +7;Z:TZ- ']1Z69$0'[C,X5A[2XU5 GOBA)@<H+%-^TVM5&I1009:L"Y2#
P>&HF\*T^K&>^<KF%?Q\P,DRC'(N>GH0[W% <)J;Z<,.$&E-O13,Y=-M;8XY):JU 
P&E3!X+P@2>#K[4#(.COE09\?6"2&_4HGS"@LS:87+1WGZ\#K:CV ?HXDX%P7X@0Y
PD/J$T<+/D2E_BZ\>0.G0XM9KAV/KTE?R+XVZH;=R;A%AH8_)OX/(57N5I76T'T()
PIW2WQ,OI&[O0<H*1NV$TERFYX!XQ9#E@X EH93!8F\8%V!N"4!!U?($$5^*SZ@WZ
P?,R+8C8"5E^^^^>K1Y-5X:@CO6CA5WWL-24.TAT@"-&EC9*BL2KK[W/^'F9<WWZB
PE,X"@W2CO29B@%(\WRS%G;A:4:B@?/W>$<1>P>#\NA:T]'8'9T^EA6B15(1J_I /
P1\F#&(*4&]":!5/D.S>B[]DX%N3)U/3*A:@';Q*/9Y?7/OF/MQ>W=2PC:/&+7:Y+
P?G8CTM&++/"KF:!)BPI[<5"67ERYK=A:#P5Z1& HRN-=,G!T!HOP;79D]#J#YI"F
P!4Q/ VH9=W26@>L&7MJ1WG$S'JX<"/8N+J6=Y"Y^E9B?#KQ1+S*/&M9!J=L!FD(D
PDMV\87/'^ Q%)/WZ"J=MQG"AZH>-31=01S/F$^QHK"@L;^[522J?F7*@96QC9K$"
P.\V0&NFUOZKZEU0K#8M7V@1@"QG<4$;?L!6*$BLE(_ 9KMI1BB!<)?,!$RK:QO/!
PCR++A 6I@"8>1B!,[3,V?PC,K^'&GZYD#+[2.8T8Q +VC2%+"[TH)RX2O1IX(*PD
P,+'NNF5U\5D_8==<58_$]M7D4C5=OHA$\WI A\N\+,2!R#?=@BT*/WS0RHAD4996
P/&,#>@^C_[G#'!#):RV7J2 I73*H#M3S3QPVZ:UV5R"-JYP].(Y9(L?IX42TLN+D
PZYMV0Q%,G5[2Z_6':>"0#3&NSR@E,7$@ZNKZ;RYFPF50*_#07TP"K3"GR&4QB;&F
P5RK8#^_I"6INJ,"0-LO'(K($YQ*.I+<<S>0=M+(2Y@ZQA>ZZ#Q*$5BJ_2$M#VH#^
PHU"TW"3%M!<>$O:+%Q%@SW*'O]8YE18+!+6KT]\K<_*N:5 /#R\AE-O=/C3,I5]B
POYCYLUW"::)P_@ 6^$5+B7=]=*02T/* Y:\@+,L#Q69MQR-SB"*:_YA\>N"B%/<?
P935*,#)KKCE&9T255Y,E[-/'C^&TO@3]#L$].+]Z((-T>R"D;&UZI74^0FR1W9+)
P$?_!O6(\6DY VF"/5F6A$J=U%;@95A$)<3N]X]6[T0M]2H/O@M+&C_Y*6I/V(.E(
P*<^T@71J2T3S%RU=(%"5=YRE$ZJ*K >. 3.6-9(+MI":WIFFM#U0M^TY>B")6L[P
P)BE&U2IB#$5?XVD(._;+,*].0E(1;(1HH6+8.>KG2]U2BH3F9$_#RE& -<IR/GEI
PRD+74_3_B[@1:\DTZ3>+4YXXLO(3[7#)M!=J1Y%C/D,7_BUS4 6.C[2:;ZE7U$73
P"  TZ%[^FC\7'7A,9:G%_0!JT5NB:S]>WC<^IWC0PA^U&3.,H9E]YT:KY2+VHZF!
P!,*6ZT7<[), 32N\'=HU],:EW3(I]=A)#YCLN;-MM0F1.KSU+[_J3SV/5/QDMD]H
PVKX=STZZ<&9]26XN+%)4@=DT $/\V8*U[K$H0'#<.QV*Q&/_7BS>OL6@KVX@4!J[
P!)C0FA9)G+;^FF4>U$#8_SV,8XG67I]2CYGB SQ[[1N$](_R5%<W?'U7+^: 2$/H
P@V"L?+C!US,K:N-MS[3\W.:J0/IF@,=R MUAI[F_SD'=R^Z7\,R$#?HU7CE4;_H-
P;6U!)GKDT);F1)'W'^"OI+E5:'0ICFW)[/9QD)1]YF/X08J$1W=,JB?SLCB:BA+N
PC$&YIK^K [*  ?)[?+D+\_SEN!NL"'[QW':K$3?>J6<'@]6PG!@(28:WQYGAB&&?
PZG_R3T9(6PT[B0_NSM&%KR3HH9,T@40.TV("P+KE'5./D_9S26'@NMW @"USN!()
PL /-\8\TTG8!/QO.@D"C'16!F)7+L'R%L2T#][M^68[BVT4!<./?=^A3Z2(<J)^&
PV\J()3B=(2O@AG,"]0=\.*.1[]JJ.];M9"F[K>WB^4J^.39)/B96KQB44YTN1AF0
P=OCE3=+<(GUP 66>"P4S'7UQ>%)Z9?=@WC3BVOYEE0+M7Z/P3R,T+U<FXIP_0_G4
P=+4PIP\4G@DCP'X8Y@$F33M=*6QXG2Z+Z6"S,;;82D9*!#*L/U,(/T%7E5<0198!
P,'*/D2T:V,+U\5$/ZK1>NER5@D?H'VE0;'&3>;+>/=NO$ LUZ(,XP#1GM(J$%!"_
PNJB3.LST$Y#XOJV/! (D6RE"_/*?NK8^+IL\8XVDR\OC,7'&JP,J*QNP?3_!Z:UM
PB4*)>%Y.L0=^YD[4SK(K.F.X B6E:Y3Q94VW8#X]-#,7@Y\V,V1E;NUSX;!$4JR<
PN(@YYJ:=OJ57F& H$3J"_3A,]K>REQID4@[;+;_.YR%_YFRNBXXX*JVXJ@^TXSXN
PX_[*=!ERU6-C('^MSKPHCC/23UZKL1TGIW.N-PB/4@A<<KB[+K3!6_(<^K-TM?">
PUPO#-$1[//:%GMNW"1HV#*/8R%GHI.PI1X_YH'A_6[S9Y/^<2B%@(CFWZ<+JT>Q)
PM")$YMB$J\,]G?!I3L_]^R3+V#F2^SYX<Q@B2786)ZI"?H?.3[C>B"X #Q;#)9E1
PRYGF"6,6ED=9ZTA6![L5.%,?1)D"N9#"-P/BZT48X,9#UK>51_F-+R67&-/Q<S*G
PE&IMZ6$'):+Y+X+BMHK+Y5EW2K-#"4K[^RC-I G"%WB'H3'XLLF$@FUPRU73[/#9
PQ4;N3IV )&0ZNH'^3 SM'1FI;D+%>W+L/,"1%4,YQ'<"<DN47D'K=V@SB*03ZV-]
P8;]J*G,UZTJIO6Z$K2?#A54ZL-;L5N:2>>6;5"JD$&&U*,NT@Q:":_I/MFH<*KTZ
PT]A<)Q]B#7P^(HNV 7Q;Y>W08ERI30,HE6GDC<@@=+ROJI9@WK^!>,J31JIVBBPT
P*V<+R!P-]%_3*KC. (.B:+@Z=O&N1,GKVVLC0PM(6]!;97Z7+_2I%"=<%O5O%++0
PMB3H-]Q*9_/(7N=7-'51:O%LRA3L>WSVK>)A]:(27E^S!PD<8_-,^#8!$= DQ8'!
PL=XZ'$8F'3.:.JZ^!C';TTZ1;+>1Q,"!M!BG+Z7QN1'4](?G,<]\K# 18?DS=U @
PT^0)-\ +QH)V#7N6A ]B^R#_G"?W;:>W+4LVC/I78W=V(3'0QC_I3!D5S6*M%W5,
P67]'!C*+V%<G-PA2%,$/_4\+O!3TPM*U*H@YZEE@3!9OQLDT%R<TY%<N1R:E\\=^
P9F>IEDB)H29! ,L6_IO9HY??$0/JLM12\4M56@E3QUYV[GV&P_ES,])T"? \)6L<
P,?W$ Z+YRJC#N4A- HRCT.]:"+;5S%1@F4[;$N HRGC/ ,PRLK *F?V'W&6\/G$,
P)RSN/I'79=93U;1S8E?!,<TH3U_XDF'2/5)/8R\&MQ5<$V<RK]O_Y@701O'+<J=-
P7*9UUT"/1VSNWOJ3ELVZ+W]'7=3&L9IUY@F%S^BX]&V.Q)I@M:K]CZ<8\QT%DX+ 
PJ,G92@)B?OC)M<2?F(-^^:-+\P004^RJI @R?3Z,69B(PGVOHH,%67GJU\WZV9_M
P&J4L:?=L AIH[I@CI%:D8"CPE>&*V!'F/^^6F_6C3'7CD(Z!CL8L:]< ,ZO#\1 2
PFN:)4'^!19)MO#5YB\&? PQ _HZ9LB\VVD)V37A3OQ\@YKQ"V6):OFK,\$DU_W!F
PU9W)Z;.&!YE^9/7 +G+,,,E8+?7=7Z.F+GLKYHC<0P"5] /22X1MUOW.?<A*6?]&
PX>%J70)9D_U^*KSU5NMO+3)"/+@V%0ZC8;P;6A77.J-.U([6)ABK24 )0LJL:GU&
P7O6\QCIQ>VJH0S=#D*?SD%IU#%0@%5F2KA!5$,?HJK%JB-L"GSQ6.DR!!WLL+8_2
PZ-!^K[ 1\A#)&[SG8P/7[TZD3-0>\."V[%9_"2>^\#8DOPLLL9,V,+]1_!,\W:7\
P(M YW<Q5,]1^ZD,& ].V I&D(=LE'-N]-J]V?QWC"&45:YFV&)$KQ]EANRB](0EJ
P0ZQZD-C"+YL%>>TM^?"]1XSPN@.C?LV J7%SI>\S-G7I$4:BXOS_&_RKI;^5%K%/
PR^.[N"S19-<C/?RK Q-2F,AJW^,K(YB AAO"'F'XX=T%-PW36;5S#%%;P76;9GRB
PN#:Y$)D!\EM?]3-5RH3#+$7OQ*MCU6.%?ECMO,+RX?_U"]^58IE%BEM;JKEBT\/[
PA1R/$L$W\F6*VM:*2N&:8I<ENZ/UYC<.7=V":A)"^AY+VE[.AFPH 5MY-L*;G#6Q
P_@7B.2#?&E?\CG-6"I2^816N0--XV>]>:M0IML35]KR"?BDH/MZ@4S<JTVQ/+6+%
PG_N^N*=2" MJF3,*-NU,O(QSP3'+L[WF6K3!5Q)Z3%:!J[KVO\[;!N&<7DLY\/@>
P&0]*U<D$<;U'GK3<E)N2SBLDG)LVQMZ(>E%K8Q*I,_<0%;$:1-^\!>W%IFI #PO0
P9*D"6@,0P: AN]WB14>J2R4.O2CU22(<7])7'+S3&N@A&_]CUA&%PTE&3D-3%%7O
P"K+%J.+9J27I91\@IKQ@]-Q&4LO.5:QZZ>9J/JLKY/1<D5[5ND9A?H2-+6^[2\CV
PS&%7=R )8#H#;&UM/&R+1,B:7P]&G?JO_6])&X=]008)-9'JJ&TFJG8OL)CK%"I'
P5D8<U3LV:@QA4?E;JLRH%7],G_,>"OH)(X8+^&=)'YG"MAD?&";7+SA2PU=[%*C^
P19CQD=GJQ;EA-"/BJ4X0@JO<8HNVM=@Z;P#5F_BJ*=4JME-+ ,_K?J@,K/4+P]0O
P,=X.<<=V'QZ;R@%5C0J!_%Y(ZUOC$'%%/^(3BT-$B_<S]=^-K_YNR?.V]2F(EU%J
P)(F(07U ;XKIP\5DV;0M,M?@9+(3K-%WW27J%<.0E%(Z;QH"W\9B.?3%RO220-\"
PQ!RMZ(_U,)_KLT ;-QL@L62E"O<X&0-1<R.";=JW<@/,=6(K_Z(.V/WTI"!$;J3$
PS&JN^7GF/X*W^C+H^J+'8<1DZC0[F_NG4+>O:>=9HYY OQ[YVA^P$)$?<X)[!SU*
P36?73NJ"30DQOXY7 8^*./"ERX(-(*)?,/H03S[;<DTNBUAVD. 1)Z:*)\Y8:H)S
P.H$Y!,QN/2@H/N?JM>,Z^FTQ[4Y]:^X#FR=^;>D%DT6P_X9T_N8-UL*: <.#QOI&
P[Q4$:%> %%720^HI9MD*.JP3"Z>Z #4<8SOK=5K\5M&.XZNM>!6@\\!>;1CL' 70
P?C%^5T"UGQ^.2NEK-C;/I$*;#7XX$(:AK[[E]3-GX#?B_1DF<DBO3Z1+SIT*M>-L
PNH%?*8#XA=+U=R?RUK%:A>%4G(Y_(99=^-K\WE3E*&W<>+WIO7XW(DV\:6P]#F& 
P:X&VS64K#+[E>J#3DZ5?5,?"G_)7S_^TQ5VY0=FW)V_1FJ=)Y!QJ.FB! <]R5-DN
PET:AIZQOX*:O6 \44.Y$5T^)X_&CZA)2&B>@?F17"Z&TJ&2\S;[;1PS3.#46'T,(
PHOSFGH!]E6=C48(MVZDE+WD^S$*BTKRV7EW[O=,W\-@5L6C#'%(Q4628%"S><JJ1
P\-U(RY.3QG@VJX,2W<2%GI.%J((=G8'>M')+G*,@7,DR^.M-7/*!&-"[^'ID8S.&
P.8J"E#GU%0_Q3V0& 0#410F2,9_=X;$E!II?42,>%9U:S&?;(Y8+ZMFFP#7$=CDY
P\#\]C=W4.8I[ES8EGYJ)%_S>.7 5@5)0P<AJ)J(A^L:5R^]?9:TB1EKHZ$DS&*ZT
PSZ3H()W-^[K!RAT=KY(2%A$P8#90/GB84[V@1L>LU587WP0:]A,%7*D<_N9IO"2]
PN'!0^M/')B6,U+8[$J;N>I!A80W+9(+C-_,$5?Y@W3@YOE*<,#=Z.OWH!.9!Q0X-
P*FTP8]GX^'J+7]-+IF5V>6+5>8ZR4EQI(U6,^L[.G6IIP1S<AJT#^7HK.^IOJXKI
PA.5%Q%)XUH&7H6D"#MY*]S/+X6G UJW+FMR!'[76JLQ# -9V>D-!?<U-TD]NCQJB
P422C45QD)F?.XQ="8)"*:\A'+8/#9A0V9=8DH"MAPNQ>78)[3'V,E\AV@(9$5K6D
P?=).&--H#7&).K$-.CTM_O53D\I$UN=& EJ<C$Z"<7*/PT>2#QOG5KDU/*A*:D\;
PX_9H(=;OYW$U$H$$' :W*'G0@ZS!P7;M/;]A,9G1Q<DL"*O;G&"M5SJ9B=ESJH0*
P8\@>>'ZTNIT7HD)^1K@A8S:*P([W!"T@RL"JN#' ;=3D0SM<$>WA;,2A*?%L;0Z4
P=Y>PP-JB :#KIHVC(6!#53X']LV:?#3 D"+=$B!,:%XRL 90]6.Q%&D$T.*Y+3BF
P^2!"/):K&I.JD9T$\C'66JO-.='<XUSCNS,!(8MR2KGZ**'?\5-&6@<N@7L76+T2
PLH%[.""4"BS\MURWADU@.YD&+]-U(4B_!GP;?J69A*E#-@_= 9'E97S_SA@A*,M?
P8&NL@S[-AX$"X:DI$!E(LVIO'?@;(GU?(:\Z6B:%](-<D=K]UTT=G29CHCB@40)!
P.,XS#K7&@KY+>H.WZ ]D=EN1Q(X2U"GX,] FODO\"?1VY;!SKCM4!T!0K1HJ+6T(
P]#H\I&=5OG]+(O?WX[@+B*V'TZ*U&H.'JHN"@!69==;W[*A/UVYJ%TXIM'[R&N)K
P(66\F#VWE8.BX&A C!=EOB_K<&)*Z('7:UVI_=O^+Z6M6/[\DHQ]K$LNWRCEG9\^
PB8TC1E>7,^^E*Q"4R\5T&#"B[51,WCFR4(A-NF,5D*A*4T.C>T-M"X$I8(^UQ[UI
P"VZC0PRP_AV?-]UK#$[$AEH5327],.FS4GY 3 08@*<Q!S)S,0WZ>IU<HHZ/3J8$
P,#@&:%]W/21AXKMN(NPH_!'S 4B658"(7*C!N+VW&67''F.[\5E?6&.*(B2_/+=]
P&#YLR;9.U,-6F=S=3B^D1LPY:I+L7X:48-W955W29/**J9>\[.Y;!NNK3=$0;#L_
P90H+?2WNQE$!@]>+&L%19F/'2P+IK]9G,Q^IURW^LS8^:IY/TWYLGUG F4H^C;WK
P)7&#>,5FP71Y>%WY:=- 9ZU*)7-&^0P*?6/A)2E$"0!"V1V'?%M27;.%((KBOS\Q
P!8\3K3.<BGZ#VD 3>).FHEG]8X9P:GA^%%N4"R9C=+\Z2[/P\2Z6<],CAYJ(T&M[
PUD8*O/D/)&/X7GCL%PY6L4J==4$F+PJU;/J>V#L=L.H^Y=EB-WP$(!KZ/**1/ZZO
PA4\5I;CA-K,&!2D*KR&)]X?#MMZT:@?_T)ZL-K(0"D_'4!'=?;G4/5,O"1JO5%\4
P[R[8MI>_69G,CK3+LI#?B1'Z3<CW^(8 KPM9G[6#$9'.(CA8L!1TI5H.5JNN7T_-
P?3'03N>%&A_W: 'B%[R! 659^@L71U.X(>AXZN^AL0MWZ!+<9\\5,4G Y=DYMG@3
PUQ>T5--!.3<I,.8XP#M[>!Y=/,5TIE\5(&L7OT.2?N:6^"IHAXATQ-RLYR8B Q@Y
P2F0OOZ&TZ7@59NW[,!OSZM/_?+F&;0> + O-68@+ZV'J;!B5\XT0^]&F)7>;"K;4
P)UX3H=>6@Y[#V-3VL6>WTL$Q$=1.^2RM^<8@>M+UV/<4I VLE^,V(NN[2%-I/R(1
PG$,K5!)'I9<%5=$24M]H&<*@' 2O9+Z&)ON3.?4QK.G@529Z%3.>OU+*/7,0'*:)
P3;2>P /:#/ZV5(! (\_\0)E9KRITQ&TSCZ^1SR<G'*O1D2"$QK3Q<RHIO61L[C0E
P4AW@ 2\"D';RSE7MCOK?::8V@T>^.ZRGL0C%':S(V_9%;;%3Z4F6%'\47LF[O[M+
P.D %PP$<$]72=K!V4!32SH,7ZVL!CW=M**A_Q>=99Y*D.*D0;0^'.2\ @>8@C/?E
P@#XMDB4>E1[&["9J1]5>CE"9/\JT9N\VCWFB(O$6X1\1I$] 9US:3VFC@E,<SIH4
P1M.B(Y)[,=;W.L:%"Z?.AI>  DF_2)EP!U_3H,'?9GNCQTE4<\$7F; 0R!GO8@BW
P,*@-BH!7$N\WGT^RD'&*7'D:+MO5V9F\3500(:SN:2HG5V</Z' *I>_+B!VB<979
PD+>/N5C;\V+M6Z<1#I/2.</V]ZILQC-$MJUEB!A4H_C&_/O6UVL-['LF'H<C#H)7
P!WOE0N?S>I[2KEAW%];KGB7&<20VKT.Y(JR4Z!66%7>9_H#%\6EDQ6Q FD&;$0FF
PZ$"X0TX%&LA.OES5+:?V48UK> U&Z2 5%6XB%M^K,VW5E:Y(M36*,SNI8^]3RR">
PN9J!TXSQ\RC;'!U@M.E'<[7R6'*H,IVL:<+E')8Q T*3@N'>T@ 2LLE3S4RO^9/<
PK8;GJFZV+M90D@ZSAIC0"D]_,RG6J>>0IP[?D.J[G]W,M3A[@58^G%AQ3X<R1O< 
P0)OO#,VF9)O2L'6=EUSI;2\9<T83(&OTAM-MT%*"!"X*^D!:$,J!M$GPBW!W<9-B
P;BSXXKR$)L$;"24D+3KZAN4B#DMJ!* &A-$A-B*R4NIF/ #W^*E0 \S4,,XO @L2
P)8S;W5RB^1?4+I*L5/U*7+JI]<%[EK"%<D)B7Y7CB=],'-X.*%3]<ZA$'$#%6"0>
PE<OO,BNM=ZZ5/!OBZ)#C"I("6[9;M[PE#&R9)/-7!F<T$DW.,Z#L',C2:$]O3*#-
P0\@O@Z/ Z92;45N+-?[N"#4,[^XL/@-T5F9T)V,2>HQD8D9,7(][M#3FCN_L9*5E
P.Y;M0J/6N((W[DW6>Q]9N=8\K-X(:>+#ENMK<'$,V.C\'E"QN). NUQ V)MJO8.M
PW,*0J$GT^V$PC 1_,ML:$6@DP+Y_O3GYW+72L>*PY8FSW18LS5PH_W<JBOW\<1,N
P#F*<@*P?3W '0WI>?D\X:&WLC&[\ZH[*P1MR+C[^%T??1D&83&WG!]<:-]:$H1+9
P&@')JX0'.Y.!W:D5<F$Z_%@1V^\/6XML[+)[0230F*V+<U-::'!PJ/RYZ/@6%=5P
PHE@NWW(%ZW-=H@U'4VDN?2);375%9\RZL9_T>2M,F8VDZ&S.9K)6#T1_>65;++_\
P/3'NQD62'6T,>EP5\HU^9ML*=</LU>\K<T.=U%+QB 0 *W0 TU*[U>_BZ]3QZ^.P
PK([PU'K3\-G^>G$!7Y7?(GA-&T+N/L]VU)V5N8J*.W"S_QNWS-"WJ.G4=;B?&1F%
P/A]J<6L,'BT_7C$95["/^5ST&PT8RM S8W;N@U9#6&J0VE_..N8AG?B[&@\B8X&:
P6M>_Q2@8Y_J3<Y/CW1& ^9GT*2@Y;ZHS>R$"Y&AEHQ[%#E=X7;=)SRE=%"..)]"[
P=UOU4TU%ID15>7.(KRQOJ.-$=&K29!]:KA ;N<YGBY'3],84+M6N0WT%RW^^?S!P
P,_2;P*ZD$Q6>F@U9?MO@7#Y3AX !Z5!52?"I$ZNXMZ=BN+1OWZ^$9>?:\]/]4@K1
PC-U47 # 0&TV,],V=C%$I"EX,B2*R]*)\D[S#P^!DL-DZB^Q-S:K[0Y .?O)2@;2
PC FC7;P1S[-AWYUIYZ#47M!G$J8U^NX*0THOAK'.3S!CX99FN$ZK\?.9<\C-''!1
PVJRMUYQ:"8"#[6>>K;^)"= 1/.A5I6A9G"E>:\6CB4]_G4P*QK@OM&1BF6GV&"])
P@".+$7C,TU8^"_K: W26.+4G1!1\NCA'^(:YK'?&3_#:H;]T9KP,R&I)K-V([=:9
PW@*0Z]O^(1X53&=CW"E5+<MR6"#ECSLV'VO>4EFY;B^#0IWK/:6T/$H+!HJ\W(1_
PFQ3T'B'L+L7GON3N+M "P2/BP4T\,+V:\==5$)-__(+E23*$D<GJK35O49%XPO%#
P$ *BXWCW8&A'"M%;Q\(%YK2^I<_VG$7KF)W:6(_G/C$QW=TJKD=Q)RP63%Z7O"(_
PMDB&UH)++J[^FR4&&ON0EI,8CK<9X1LR,%35#?6JPI#^L\#I+3Y65#Y;]6R:@#&3
PIQEX9<N=I"6D,8T_ZGZ9T#S2<J<HH?37&O7*]818N*6YBHKZ2[+O8DJK/Q8_#LOW
PIY!LCLNH$Z+5MF21!G3Y]4CSC,&^Y,6=533+3/WQO!EPU].E!>ZNYUUM,A37I+'W
P851]"IF?CR%7][@\>PSD*/?YMC106)6$]?VY>8C";7V$I+3K?:JJN$F.PFUKP0U+
P^7Y4\RAA?36>6#C(8[$\/^.0M+$K7DYS0Y2ECW(5AP][@FY%4M/BOH+1;.H_:I#^
PEHTHP.L93$+83V>A1T\[%>)PEFN*\GRBVOI08A9?X0/1^E[2>[I66;NA.MZ]TC/J
PG.@ Z$WVHURNHN4RJ_VUUKQ+OIT*OI"/U/5 =K<?X5DNJN2LV'WE7LVL3X#]D579
P1SX&-Q,36*R^>L8A2@+DJ\S="]#$!NL9#Q>>_T=:9-Z\<1OL[+G""F%]U:G\5M8A
P5QK6>X9J#.ENLXY20 "8R85[XJ?B+GMA@G(&&G(4)?IOZ=J #S$;]0=X25@PAG4#
PN0GC+?.K/$W8Q R.65_1,H$%C2J(B@K(B0)3$'.,IQ+@08!P*=.30LJNN.HOZ_J=
PX[J",K<%/5AAQ7S/\U"+8 0'.TOZ^<"T[L]"4=+23G]F Z\6'KUG'?A]%XW1I_ S
PK&@@3?G,:T"3/F7>A\9$;2+K/<C2)H^4=R+"K[]3O\[29Z)VD *QP"Z C.#4<N#(
PKK**:IBXWRCE_8"L3WF$G6>B_.67%,:]8N_Z!+>/(Q@GNWM3QW"_"-_(U$O(&DI-
PKON+UA,^;L6SW?J N9JHG\U-5TCGW -(JZ1Z)5W!VT2C&F#+3XYC3=^/@QVX/U6N
P<]0'J,JYV K@,S9*'=LL$D+'52D=!5ZOK''LSMM>[@"GW$6'+XMK@'R(0"*E%OU,
PM-R5JW5-=L?$%%OZC#$L[6U>R.#<)BXSRF"/SU971%'?3W-55SYAGFDG!.L7OO1]
P=]A'@KHRTP4I;TC@P/5_.JM)#VYS*A(A! $3]KY)-NDS[6$*S[O\/:M8 K&@0F,C
P91;,8RUU9JW]MB?<I;!+G@NKMKD5XBE>RGJC*T(6HX5+S^,.DT$?;H:,"-&/A+!,
P0YI1+#Z*.0J>J8.KK0:65*CTN*\BX"3R0[/E/],;QI<K+/<[@)$ ^^N.8A+)54O!
PF;%-\P:-@+I];A' ,%-*+1Y,?S6/VA2@/5%&8M]+'U&ZB(?1JR^ZL]>_D.Y;D/'V
P[%^![ /;8YL8C4S<5TC7?!D6\_T1Q]PIR)3<Z9Y"VN"0X*3_SWDVB:WM=J9F&!4T
PWY2DOXC(AUBKA8^P_6\^"T.0=\@X^55%U6&:*S[]@C&>NB8%O9FQ&J_E!*F8^YT1
P%?^B51'0Y#0#W:#)]>N_XE+-Y02 =VC]FM.$,["TCZ?1KA2*=BF@W=#.TD%>)K[ 
P^$ 8/C@ Z&,;GO=@?ICV)0NS:/C1 ZNEQ@H2DZP_\^W&>GO%5;WRGJE.4E"Z?_9Y
P!SN ^8Z%<UA.>#+P&;0M>@!XK%=EMQ>Q&E1\<5;Y:DTBCPQ#TK<7'!1K14;W2<:U
P0&=1D/B*RJ2)(@IJX9%&HY86F\B-Z"F_QK&K:EB:2L_6:M]HXKQ7 RPO0P/UD7PK
PQ<-(/SU3![8+MI.=JVO!0CQ7,*H%\;?$'7!CM$A"OSJZN#\J!^2\U#B(/S:E N28
P7@*S*,V_G7B 8-/R?%./B"HM$:[)\<&F^(Y6+X0TA8 KW%J8##*KSL0BX</A'ECO
P-F*OY#<$3DN;CN:XZ G^U(DK^,W)O<[0816%5\S90$Y:N":7+WFN85$\=4IU\BH4
PTYW)]PYOM*S*WIG?N'=YQ/NT"H%M]63O0V>+M>NSY:(B%X )7FQ<.0"V-I"X)6Z0
PO12.+:PQUPY5)O J2&L6-.#/?%4242K05;8^/YH/EE$*Z*@$:<(\V)3?4M)GFTN=
P113!WS3G:HZSADR$406^Q>IT/]GVE1%JGBPC"<KA>Z668("_8EJG>!Y$GE6]CC[<
P9#4_(Z_!K8]!R23O6I;S61TP6#MMF?8(5=@O?F*;U$P>VZFP,5'BF?]0ALC1N+;X
PU =Q(CHTM[<38SD"G$>LV^F$(%&8[*)<1BP?%E58[*+DG?^U9,;JS*>$$$PSE0\K
P,<=AMWGBE0V%I1:L$PR2B='9!Y5N L:NI9;[O^LHSZ4Z,4SS<>X5VW];[AB?J+J.
PCD$]5_$IH=#_)G)'(VVI4$"(KM("RKRA/QBY^A&_38*>0G^FX4^8/2,*7-MZ75U5
PX9 S29)%<-/C"P/SJ_RZ:X>AI80:*A3!V9$BWF)<! ]VS;-V6DN0QF?:Q.1K[8MF
P=91 7[P$-FFBE=L[_!<=@=>7QD!9RZ!CAMWWT+PJ%6MFZK_"0Q)&R: )H4FX-L.U
P0)%)Q>-_:KN& S[2D(RG4?^3%+D7?5SS,<VS1LRA> XIS2&(\MT ]QZ8Y7QL,NZY
P0%*QZ-#[\A6L3R>J)CJ:@;HHT-KZ/$]_O",]GUZS)MRMLWN3[.H[.1D@^_#><3]T
PU"L6" 00@84F#$50@V.JE29G]7X 6<I[_SY!L)"'?_M)5"&N0N1C?B=63\@SQ(Z?
P[_\/>"19DU)]YJ!ZAMG_(FFU)6&O.M$!4N#ZTJ<AS<4&P?26F.[@71+=%G*P35^5
P1BB5 PK?Y0X<P;O5><$!&[=8;AXV75!A@'Q<7/IEMX.\KW:$-S5I7'-NUG\/O?.J
P\YC"$L(/7>_L"Q5XJ='M^%R6F/U8JO?K_&,?NPOH3?)MSM6@*P7?%<D=$]O,MJ*1
PQD4[?D)3H^QB2N/EI7-TF,8<CK.)O0"_][S8J7MB/V$[72J*'SYTU^2&.M\2R@8G
P['P1ROJ0"Y+<92$+JW(>0D[_,QXJE&!218\TO8D2)^7HEW%ZC,JZ(+TPON)1YWM 
PP:DW<0'2:9:*QWF#=)A>EXVA?J5!QE0SMSI9VX:M=?0AYJ0PHTC9;%$^_$,G3U-_
P-YDN[U%()8F-G>TN8W35S)@/9G0;%SSJI9%O]QNAX66^,JCNOG0VODXC$6@[&5W;
P#S>8 I&L:B*(JH"8,Y/D2F*:V+5V'ELY:'ZEQ,,2-BT/URI.:O+9^%6E,O$5EXM5
P>.S>Y(R[6+(%HA2]<7=Y[Q&]5AM6A?+GF;6MSB  X1:<\7C2/ '*_VV3OB9O3X-X
PDV5AXLEJ-^N9DL+)6I?%27 BK>GCWK$08KS"!BP$!,N;FCL)$;7^<_C>GC->&TLZ
PT-QM*-.'<2$:KXZV'5;D2P"MNB4VK&L3%8XSP-#@8%V,"UC/&B6"45": /4=T7">
PU8];^[<I:G4APEJN=(SC_W;4&HI:)[NA5="[A@M9K43$*RDGECY_$W?C2:^L$Z?$
P,9%TN]DX[W6Y.1$[<SZ.67*=HRIR!L69MOH?D[Y\0Q=O0U$C&:<M;,_=N<+L&=L%
PP#FK/7W4R;TV;",,%A-4%??4LI(:!,S1$;)C?M9+]OJ6H4MSN>E]EMM.J@3D_ZO2
P@M 9-%UNJX/_+B_,1:L&3M<,15Z7./FP[$C$F&I2PT^1?F6@NI%9/7C9-FA;(I]G
PF7EZE96^4*_.U8"AP,$=O,&S LE4T2*45=SN:LR:RV68%<(O',E&(MZ=<X"\.;%I
PL3_:;SW:?X,(MI_%C1JK<==1&(>48/R<CBA<)(_>ZEQ-3@$4I%A[."@+L9X*RTMG
P@P2&)'LBZE_C\=/UW9T&)B;\"\FKV\]WH(PP<,SQ1J-4PZ*MF18_>%M7O)&QK\:^
PMF&X*H1!H3>'K&T+-/;=ZZKN!/_R@O=7H5D*>!WZC8PL'3^2GG5)#7RU3-<91O80
PPYMFDZZU+\!J:BHV P3_BKRT6YX/F<<=NHD5V!0;O44[-C<H]<BVJK??_1N^,.8W
P^( D?]7S:W_G2+D(GCJINIA;UF8@&R-=F$SK7TF=*B9!U$6 IT_"1*,ZY 6%2E45
P&8&^=4*P3E[->69@O@3=>,YFET2=SNLU-6F8>Y"?AN3_HJQDF--[#2]J9*+=P=CT
P@.(KC?:2UC<P5(Y^!S"WH$06U:.[@\Y7SE2WCQ'8)?.RT<01OA0B5WA^ 8/IX!K(
PH5M/2ZCGAFB<94^O98\G+,\$/W$X#FG\R,L9X;/<$*+R%%Y9<$Y)9'D@*#(+F"W@
P2I"D#0-_]V&77V6/0$[%96(4KS5484"R>#:9.:S'(KY')?WT6;_]1-<SJHO]>:&.
P6&3\OU&30\(OR"FW/;(7,,,W(H<N\Q'H'P2OQ3N/I6T5O^,7(( J4;_LQ\%=,&K[
P+'6@*TU[(7NU#I?XHT8)+AAXRW@;UEEN,M/^WLEBZV9(,/.I])GAV#NQU]..G)@H
P5!\^X8\0AJC%5'=D]H$^'$@B.*=<A&A[)Q.>(628@VU]LT@MO799R=.@ 73"\SM\
P&93FG]L]?+M2),1!E2QR:.1QI;*X&2Y$P]EL!ZX1H,G\Q?MR"'VZ*:XZD\2FWQZ'
P#,NU,,!OASR8VJ/YAM"6-UK6Q.9QHZU!C/'LOLY3%K8@^\"?>CBMD,@,Y:/TMQMY
P/E8S82^U3M(6?BL'P@WM626%O=F<J6W M"[2Q(=5RI#8ZY&JG.S@CW-C6'8UH3>6
P''MLA<KL#SG_Q:%7&L E(T4(V2)O.=<@ASNHNGM0@ML&R.7<_D#ZQC9[^/=ICGZ3
P\M5A6G(5V$.)I<(U+AV*:C>:$F8Y)-E78ER*3=3. KH0%11LIG%;F--U!5)&? Z=
PY+S^G2],]+,IJ+IS' XB["$R7*KIXG!'L</?.O%1%3(UD.RESD+4(^\EB/#90B<5
PPP&M$M+YQG&G(@WQAXS&JBGQ*!S0@&H'4DI]DJN_E2X9BSK9&BS-)=E^W!KI[>'M
P/=$U?':5D+WY-XE&'X?7B0625_LB.2Z!)S1U$Q5OA'(DZ91=08,&M"TK>UJ]1:#3
PVY(8)82ZB #W\C(R_3KI@0S6<%R(KYT$0"D)>5YVQ0[%%VZ$NW=+(I[*/ ;:L@M'
P^S.D@8)B'Y-B;M@+]P]**!ER]++&!A\4X5'KWW37.DET9@<7.NI1(BPI9?1693H5
PA:71806] +.SGZOC9LBQ-1!-^J<7R@HRK4^\'F!$<72.D;V\ .CJB0>6<][V9\$L
P4@4NELFK3I]=1,SZ#<1SC3#-[!LA05\N^%<"_H[0*-! YA]/AB71E1EPK8 -&O_>
PR*'.CLR\EO!RW?QTP$\&8"ME=+V$1-EPCJ4*Z69+%YHQF[1X )SS1"QD<BSG-S>%
PXP98!%-E,7T6?V1IQ.=\7/GH0\9C9WMUJ1I/4?&KW_(5P%18//\8Z-C!(1E<DI1R
P*F6J'0<()I1 =$+V)) E#MC$LLO@:=.AGJ" !AK)W=[\ R28(DT-&X16H6YA<5>1
P/H]OIJ3OP V;6<%[E36W<;_C(K+>@'%_DIG1J8+*;/TQL+(U:J*Q]'3MK\ZI^5UG
P&;=Z-]%J.@0BN^RY4&ZV3$"_D*N,H6\UY@$L87K 7CXA>;:]4>8D_2IRM>]U5H8*
PU7JQOKT)U[.W18 WN#T'$; 06> $LGD]#27?>VJ=77N!1ZXH".Q5!M'[SF/+RYL:
PY,@;P,?,0,;@*]I@\3UDF1T:9*)K$)T<Q](349'8%BPPA29_9:A*VNGC8;E$D"L0
P06I'TF%#PRF#;%/Q4@0[%X4UYOR+S,TPC"E]>4@DZ:<8DQ)<;+<@P7Y7>Q1X:"3P
P*YH7/@INFUU J?N#][$X30V*1ZI#*7'#=S7_3 93/4SHP"!\+5X"[S394>D_"D]I
P,;$I4X48T.G'_U\N42I<"C(?'\U V)9 IJV6VVF,QB&9[.5CBQKL3+3O3\[EC7\K
POL7Q\^BKY-MD6"84D;+-?C&=Y\D(_$@L>#!Y(]DK?.?,.Y&2E)>Q\=\Y(T]'*X1U
PO8#._0[[B,IVP-@'^N-)5.E()::D%H"#9*K"OV<&[(-QWJ&3FN*:@'&Q"MH$,$$Z
P>>=ABS)?PJR4EK]7&#^P.@!AO2BZ[3Y6&KT"# O1OQ_7ADLT0[5#:++!WW$/(\W(
PVT#'8_6>E0<Y0J+EE<!9PQED(MAWYV!D%>UZ:3<]-QE24;[BP#DK%/LQ!<"]M"@%
P(_6[,LN(<_9_4C>,H92_WN!&_SJ*JE>+%]R)[(]X(HG8$3=ZR#)O2+,]@)6X+%TL
PQO%-["E%Q4E5GSHV5'JE!;RWMW+.W'<T[7O;OJ P?;RXE[N]Y\OW1D2P3TY5PTIN
P$VI%-XO5S4@^Z.12%LF<XM0^%WW/1?HDJ=[V5^AS.B72N@>EAN-&_I%F5+J+=:N_
P&Y6@E//O=6\UGE]6#T,XG6\*QW:R6O<<"D1:^)3J#LA5I^W;:5&C8E#3]J36K 3J
PE" 5)W1^&'EQ/GK$R,Q-,1M?$W!,!=M:"[154^E_U R88F\<P)YFHGWNV4R%'+_8
PX?87$9NNU]T9$/Q(MK671<8*K?4H[]U->MQ&B-L"I'\3YZPN3-N%3G4/CH1#+-ZI
P;0FUN>L6/*'EFR-]-(;B5ZIAV_IGR]!PYX%FBL)M-)R:'<%N-"A$H_1-!THU#YT9
P> O8&<33O$D5#CKTRH+4Z0V%;]'!7F5:-+]Q6E7N N<J_=T:>?85$A4=T&[: &)O
P<]+1;O[\6YX6"'1['CRL!&-F5F*WF@%#UE?DUG+\1FX#AN"78,4AL.T4/U)2D.(?
P%/$-'T-:_F<SM3?]>H4M,A69E,17HE,0Z>EH7%FM,W0/EE+%#2W8%B]'1141=M$9
PRD6I'""0*PUWO$^;QF.4N\XH!AB-GTDO_B/&?9T8_3 9@T"*BS?L3NA(%N6]0\JB
PPA!_'9CI== "'NR.^-&M$U\]^V?/J;L+VCQ,*&]W,K%U%Q%%.VAO7[^^ <UE*9$G
P[WVQ),S9_!:!P^LV=!&&>HA>V:S6&NHV8[]6KL,B;:1E5.7 <)8@;<$/OV?#$;C@
P*]RU12)W786Z,EO>=@W:.><HJAH9_EK;7S&E 4U#\58C&8 !9;7,!%K-6]:X'U:P
P8)5"@[Y">:>0PS]D!/6\S6^_CE.ATYE@'%)]D_JRK\#1/17XYF"I/A^/,;.HZ)>M
PLL;^/>[+*AF.3T)=_7CBOZW*2,YW2^,- "Q9,@/5U#/PS#@!5 (XS-D8;P-2%GY8
PWE8.+>1^JEDRH^BJH%_:^&"45[NT4<83C5\*V2(LXP0/!+J.*A8BH[,YQ*I_TP39
P]3G@0'<>'A\DK.8;4,D$E%/KT6"%<DM*JG@-?![^ 5]VQ3<13&O;O1,B"ZC>I1HV
PU0!XMKZ^WI<<;PY)5 $^DLZB93[ 4AH.@ZG*PT,A55_D]FYP&<Q@,W<IT'Y8<D45
PQ_2(A#*?JI+)[-2'/B*?+KP?N$<);5<Q-2(D8EW! 5 XST-30'QR._&(!NJB-Y4<
PY,UIQ,YS(-]\XY%2[!#+50_%C<Q"88+<-]OD*<"].(ZKDT=H;8179!OG"A>[]]7"
P<^$@M-QV12@]K<!!;YX^M ?8%H,B'LS2L70ZDV2@T$1* PCQ)#,=CJI?)_=@43L"
PQU/P'8H%W2NZ.O<+%AJ-)9\$QW'=@;0Q\+=[4+CHMB3<$@P\D[BNA,>7"I\O_M;!
P?6DE8S;V?^$8]&-0S0'Z$W1G&*65%R%[SI.K3>A(=.)VX+B;J/D$,Y,7J@L7F-W4
PUB4B8G--*'T?NC>2<9<T2&4K16Z/71=,?1;,)*^!L%?33 PN0F^AE!4II^;[H%6,
P)>3[**G4B'1RD274[.96#QXT*-W<6JG.T%^CCLF*CND]18BJ!N"WZ$D]$UU7U5S2
PQV6MBS=6BQ@:FLA(N)GT%,8Z4/U0I8AP#[^HPW/&%[U-+69+P/7+7#>6C'ZKJA<&
P8F[C$-3$GY*K991 T6PGT4\4O:H!&:1< (/G@'ZUTBI7YG3H)>C&R<R=^T 7_X5:
PW?>#)S*1^(@+R1J<=5#K_955%E-ME9!:8L%*=0I\>>\Q:\C@1[L9**(P/157$110
P<:[=+E/"(2&7,QNBSUDJ?F<_+)E3T(20+<VR#>*CZOI7FM+T') I9J!)214+*EBS
P* D'.<F^63D\<.E(G70%4*6(L9.(F(06HQ^;_I'58,Y;8,NZ\E'A/TS9Z5GECRG,
PUCB"@9.K;#.QQ(#":RG!%U+W35OTGQ1!+6.FS:&9OSCS=?^MB[1C3OA_:?94G]@D
P&>=;; *-@4Y;^,R\>.T5JGAT,2B"IZ(UH1M_*<T4V(#_$OV^)^8O#P/5.'QP:,;S
P!.OFZB+ZSYKU]&+6,N:L;@RY+ZR*&V9#J\ZGK>[;!B:C12\9",O5U9RX,_TXD5M4
PT67)3"PU^"CCN?ID.U.(;:JP>.F,*D^51EZ<($YN(# A");5?%A 1_WL59 ,@/*3
PJN9@5_P.AJ!:/(#(3ZJDXRXW/\T9^_^>TI<CF=5_GQ6?2C$2_U2\KN^K9"B]91:F
P"K_$BSY&C6C*W5H=C*XBVZ[%.1R]'^NMG/A\PDFQQB:L>!<J_BV &H7R@_XK3_"?
P($>![)]"Y+FVLB(((NV:!Z.I'(;U*N20?_HHZLR[*G_C[P$ZV#SD$Y:K6#8 FF-6
P'%E&:"_-=;80,)TL)0)QHMRF5,_&1:_@> CM]VB?/A[\-\8?:3FMCCXC%XHROLGA
PBIM?4"X/> "%&G#?7TEJ:W();%SS:6 "BIZ06DML'IOKZI0=>7W+\<N9;SWGY7UX
P_2"4((VW;%(<[&T^=8%$;RN8R\,9?6X5]&V"R:(UJ_X&G_%O/H;$PO]EH2#5D=X6
PM?0?]D.#\/0;&RFUN .")C1!WZ:U!3_QUXAE\@M%S;N+%T.[-^5AF&R  ""9F#2I
P(1MOS4KU\P7LMGC@M-[",=C3YTR\F LD9S"Y&86]3]T2/@0HS-^1X54V$KX,JL^9
P1< :*)B#RZ<NCBA=<09]&Y[XY8@!L0I7=+1MU3I[A?DZ5+OG,/FUG7;.Z8NIXF?G
POL5YT&Y'6?^,K47>U9+G-(WIN.\E>*2.$?H,8D.._:Z,65+P-=^I1ZD6\;4<T&H[
P^E3:$KKP'T>KT/E;&N7E3E;AIFTG3'-XDG&EI8$F3:-K3GK*T?-_/#CT':O.5GJ_
PA[9'HK1HC;7]NHFDP FBY$'VY#4T1^;/G(<F"":H4#]GRY-/$AB\#\&M*87]9>=:
PCSVG)3%U9;22G80%ZWJV_5L(63P]B*HDL(V8/5AL<.^9'H*2\[7='#U"\\B%35AH
P;H5]72$DW_M:]H)C0^_(TT&@IH8BRV(B  Z*IRWOC?,EKIVQTOK$E\ -M]IZ,T6_
P"<VN#HX,.(S2PSP80*R'@7INIR-9]*JU*O$KT'<YFM<C'.@0_,)^.T8BZKI'HAZ8
P#-Q;MVMFP_)LDF4YU\_&00'8),B:G6,SXK#=BUQVM*]81F/U[XVP\?3,<OSRS'L&
PA@I'T>/3BGLIB]4':9X$!R-P99##WXE3>\0NB?--2J-G&3Q%@*56B['7A_6GFD/W
P%B^;I/OTF)7W5S%JV$BZYB93Y2O/R7^A\@Z?E!YE6P$$'^A['#8^3P6C+-H2Q(5,
P4#,*.[#3RZHH0T&\MZM-TNDD&A(&D16WM+)NLXY=U0.P07>2)CU$]#-=<L4AC)VI
P#]J(/+'&:'6/-:8<4OFAVLY=GH2@>-)<%ZP*QX"W)^T[?O%P>]I":)4-X"G7W:!*
PBAT0C)TN"U\DBUBZCH[3_Q19M#T&,FE'6I2,K[)NGU1L%C'OAN.N+05"2N7@UND$
PN6]FWRHX2._9W 2:G3'G"4"\@M^KYGQKEW*'?V%XPVXLC>@^U_V)/@$\$TEX752,
P9>H-D=_D2]AR,'.7!$7Q.3M#E"3%RVA>OL+0#@NW_VY,"U]@>;Q_"@H%%,^-K:%U
P:D%K?R&&CW(>;ON\47M\F? K:U_/KR-M&PF+!#6ZPS=U9/(T:KE;6A;;[RE?)_O(
P7-H7^$@C'#4W*.-$*4WF8SZW%6_/!E; ORD)U^%:#PC4,83!LF_VH;+& <!DV%-5
PPVXVV8RTZM3N1!?@T/+S3X]3G.^IF_+M30,;'GS#A3MQ/SFKQ:G,EROBF2.I3- >
P(3AY";%R2OY:>%.1)100XJ3 +F=*]Q$Q:UB#=N.8T70.,(6+W9BB H>"@ D5*]V5
P>"J*S.?#%1#::7I!HCY0&:@C]3\\/UF6OE9+KR%*39EN.M'4IX'F9O\$8_?%UT@0
PP/4X4BR/8J_%B?O&>TG@AA-?!?.@L.9>0/@#T*2H^5M]-:$ZE&3"=P9HGNH'4%LH
P2FQ,KKU014 'R$V;17J02K*9I@#?BI]+F$X=.SB &RU%%GECKC,F/.E6FE0=31\;
POZA%3FC$RW-Z&D%5K0>2^?9IOQ+6A=,P$W05O!Y[%=P+7FQUE<*YJ%46(( -P4.L
P(J!V\!+\BD!F&/$!-HL5K2*E=4T>V0DGYV5#.725I,2\RSE.1)#'^%6IC6T1[3[V
P:"F%Y1@21D9QS]N!:HS64Q* 9&<G(V41-]O=<7_5XM61>7XIZERJ[^-W)Y/7B>02
P@ ^'+)R"8T-W-%)/A<S;$9%KV6[G;SN6<G'SO YHJ@CEW:@X0Z),,,/HZY5V@:@.
P0])6-<3GA/T3#),7VKKF'C+\1ZS(+SV':93PIA^4:W#2GV+X[<5$N01+=ZH13N62
P^)  V@(++QFT7D8#,UU%OZ(#6JL'##A0>-H><=X]RG> !./H76KC",_4]4PP54G?
PY5+-^!?I_=X#>4AW1)MOGUQLRQ@EZ[</)&ETU(A5>-T;  $F1*F"O4#FWF=WY/&L
P9NFUZ#JK.'BZ9@XW::^1T@;T?X(X [XM&^5WG0I/G,DVR'26</Y^42+Q%_>BT1T9
PX^0IJ/#=K]SK@K><QIS[$#CXA#SY.9L&O[V3/CHOB.@$A:33RM]?Q,KWI[&M6J G
P]NYW2T>J58R$WCJ]!U :F4#T0U/F#M1YLS.MQF<E&[=G^$"Q>,,Z>I<2A#YTZL0R
P&'7H>4N@X$HZ>*,_H7+Y7(QN >K<1JU]2,;A^J!U(_Z/A%!G<B?80K?%\=C;(Y*_
PMNT3DEW>[L""!T6X-E)A]FI^NTK%4O387YF\4@B2&^1[D1]_DKC(H,B$U)08,EP%
P,N)Z*ULS :>)R_Q :"F_E[+'7_%PQ\:HKZ;&A[^+0OC=[X7_/="-(-(J(D%#\E1"
PSK;">N8OQ732+;R=BVY( 0Z=5B+IF/R686^0=B>!,-0=4(8Y0/H2&=;&US>(5MA6
PQ[\OD0!3D^TK:#2A$@+-*DOVW)&@Z+X%(QG7PG)5H%W '!_%M8Z("?\THB9;#&MF
P5S?&;FH6(H5!RQAIGKP%SVR@8E5MT-9T;U,2FKCG.'6*;72LLA%U;]XH>*8M4VN@
P^$S=ACH]-I,2L%!#_C1/LY+#='_V-4;\C1K\OCL:43!D9S4W_D1;!9D'ME)?&!H8
P@(K'G?X4QOA!Q<++G.ZL)3M_I<<2V88WOH.%<QZX^FXX7]Q",8);?%SN]"N!L()8
PG&'G5-;9WBYCR(B"GODO:>3FS9]>$ @Y:6)! FD5V&K@]CZD^I2JA!_CE2*$0B$Q
PJJ="]O?MF5;DJR-P$I?T,=MKIH409$"!2#00WC(DY#_-:OEUPO8L@;\4([ZMZMF5
P 5RBE\8_-M?5W.MVJ524NKGPP_F*\'$1R-TL8]F&1%T\.>=OIIB(.[<=4;+-WX5O
P$CVY]IX;MNQ2NW?1S0O:K)_$VZQ([/28(EDYTD SQ+X.++%KIG+ '.W %Q7.'U7U
P.=_6H%WF[*#QRD8?9H\=YH$!GE<<J;8"(<67EONY$O YR&2[ G+5(NJ@N2DF0+Z^
P,(G8SG 5WC;U5M3))V(]=%1NO= 7G]2\:ABEO6-?)*N:KE5)TLO?P#S^W\:LC] 4
P8VAK ER0XIR3&.^BA)%G%$'H\U[1^U327_[C+%/FTF/#J&7B80,93G ] Z J!=>S
P2R;Y#THW7=:S;Q263-8"41IY)#WI.N8$5LK-P^:[DDJ0828"<R=KG;, <'G/8Y+[
P"0-C5A:*:_QD[7N?S8X I6'7:%IZF3S$SH?-XI$#Q[S5Q1+#A^X0J)-1S&M0?4"K
PNF5KJUBH"X3[N%-N(]<<):_,1&S>G+. XM4[Y6-!-W $WU1^AB#%6ML!1=,04SZ3
P24949N4?48Q'?Z)@IN) CC42HQ(.[!=E# JQ*7_^+)NS_W<)S=_UM1N9<E8B?EG!
PA8RM9M(D$K='@I\3-+ZF JA'HGQW%O\-VP9@FAATUWKQQ!M5)3]ETYL&P(1/4DJ\
P\]%AEPX,\K6=CA%YM!"N%9+0.AW&SWI%1^L7D[S')%+J=35LQ*Z7-+?Y%%FD,(%A
P68E-]K=:0HP 4GOZ&.(=C,?XF]8KE+ UHVPAV+?63O=+&RW-17()/-I=W^L(#O3Q
PI#Z=E=QL%K7=(V;K*QB7,QXLEU/^M7"ZR-X,UA"M,I]HW:MPP!783W%N8@BI&"<'
P\!F.KNHW /%5H*TT3P?B-G-'DR(SP?ED;J6LBYMD$WUNC8U13^),3;97W7/EJD9Y
PU^ 5QW1HJ$$U?DLUM.;AJ%@[&PBAG32+QB?YL8D^]5].>-[Q5+X@_-D..NH ME\,
P1?TAS-F2S_>5*>[]PX7-$H3NA0?UEP48B^T(Q]7[O-5O2WZ8 @TBQFTIY]*;0"F/
PS^?#!#D5IXSYYLF-%6OHC)S)/Z>]T@@60FL)IUHKS^:9A8DO- .,3S]%O)(>.3!@
P*XB9+OFDS"N\T7N4(J5^IYEA[6"[#EM&X=->*TOMUD,J=^U_9:6(*?O0+3HLF[M6
PC*[[&>V#,O)7QO')SP<46&[*=.795T0D@D:)J<"\A*RM2X@TQ\[-$9=ZO4*4E(&!
P7I"7&/[93F+F-F_\> B+!C$8':/8X0Z\&K;8HER2S;KTLM5YHL62<M:^[0*^^$)0
P!C?9MS@M&UMT6[F%4T_>72S.BS?T[GG7!NXA4S-,['@TG * JV4=!TB#]W#E6[D2
P4D)L( [W#0W3>:-SZW;%5)A&H5!V2%L:0Y5&DS*A%+@R<(N(7R_Y=L> C@!%/,]G
P_7HFK\IYD]5@ A!3N!7V.";E9%$[U-RE=%)#F#[KG07?T5A""*^ ;CCU@GUEM<O 
P*H7VR,HFV_M;^_,8R;04[:+S@\NENZ/A9J04R!O7?6N9L&W$%A_O$93"Q:LZ&#SG
PM]K-TER5"?>8,3$2\)VMCHC,/^3G:I["\1&MN4WJ<;=O'Y1D\8@WHD>0Z_KPPY9;
P.:#&XL!85;^TB.'VVO?$-E/1##<)^>O:TSO3#WYBFDE#K%+:K)$RZ%ZAWENR2Z=S
PM5GBM[,O; .TH2Z->U5YO/>6,YQ42E#@@:G--^4-'JQ62F5&/ %FJZ<)@D'AZXJ!
P([J!@!L&  #.#5Q, 4A<NT03P27R"'O,:!D<,Z/N,>F$.2^'T[I) ;$U93*PX2#L
P-*2.PW>]$X[B16SZV9XNN*"KDA<K%$T#5&ZZBX-JQMK:L^VR>CLBG2B2?4T5D<Q-
PSJT PV3^8#@^F Z\M\4[OT100FQ>:C++]WT=2:,WK!OM_3%W/7TFJF;'!O]-6#;H
PU:Y9A7,Q=VJ!FH7W]1?OQF=1]YU&@.%W^1V_&/65SAG\E].RS8A3(UO\-74<-&93
P6CVY1=IC9Y1M$TKBA2IE1R.>MC[U21NI-_T9(, "H"[]H.PR32"/!_!ZI39Y=?D4
P?R7$9K_0-$)$V.*<Y1?,M@H$#QC^[8@)QJC@R==)E@V\(8.1\VS!_8V+36O^;=QR
P7D!)*AO!<GMY\)%JGN>$2#+!V?27J=4W]&_UC4-)841:!?&JB/B=12G!KQ7QDJG]
P=5=L/6*G) X\*Q"C38*VL9=X1/X]?F!(;,5CO13MV0HV304NQZYT\A:X>\SXFE%C
PWEQ%CT];%U0GSXE<!WB8XK9/] YO!U\ G");FR[?R$=DI!7MI'KI8/+VORY5U?(5
P^!.(:_1-V:J4BJ9Z=A#34..S0"@0@!"I?6!98L<Y7(<%_C$%*:'<V"$'+[#[$9YR
PMZB:*GH\T2?BG\<G(O:QUI3K+"L4.!Y)U0*03]CQI'O),:* UH#/PZ$V^UB/SS")
P+L*(#SDBK?#MVGJ[14UR\'<]/.$%5FKS8SH5SYR+IV5V=P)X)\Y342D4@*(4AA/@
P%,O9Z#4BU6\L1:9,4$UKS#9:]8XTX)ZWK:PGF63HRT'S)0M')_E9UTQZ[3"L(+E'
PT^]9M^]R3J)M>O! VE7M5[DO_&D/":@G\R\?2K2P>?,A2>ZAE_1J[JI9TYAY4O;;
P[RP4QCP0(++\RM+I$NI!T44T.@5P;KFW1S(V;^=3&] 72247*$517V!\-S%3P7>I
P!_\,"N.FF6DXRP:T'NCO4,Z#':SR\K)N@HZ58:(1-M"ZPZ/<%254[-C5[_\:F$X:
P=]577AKT+RLO;&2TASY8\'0=1N+72&\-X1&B$D&Y,=WG>ETH"6P);!^K,YMXU_(5
PO\:"W@PR9KL4-=L\H1]O9/.;A_&B5=SA']-S@T/0CH*)MMU9=5?B^%3\+A^Z!M/B
PR./1K;JB6R']A]*)<4OT;=>7*JNM9J):24>!O%$X2\&,C28@I\_H54[QX5>?=4:V
PN6NPR<OV3^\;LHQMQ+II:*&T+DTFC(9:4$=LYEPUMP,274F,>2JI.IW:U9$AC1Q+
PS,="ER^?!8'!9(0X3&*$\4RLA( %3Y^:"GAE&"096T]\CH:R&:IL)*7%]1D)[%F7
PQ>@XJ7%S:B/3+TU.[@S+U9QM$6I*- NA3 3 /X&@3YEC*F@CXUU-.VTIX'Q+T4];
PRK1W:P"NU3[K@FB14EA.#"YU[D-2LDS<;3CD6(^12]D>A\(9BGNV!4(I!VUF_#8-
P9VCAUM\& $&_2S-2[ :E+X=\RNJTR5!328V:OL+%J5?S]:4#7FX/5>RME%<NNNUA
PPHMKC@G>"C8V</EX(YU<JD6EK%V5BZM_QL3KP^CVV6D",^6A$TQBGV!.$E)BA?6)
P8R38<+.:$^!%>MN:Z=\;>?R!3%&'5TN]3)DQ,\A<T^-$AY,_RX>.)P*"@5'-!EW*
P*T.I7)/T_K-]ZGKWTM55-JKQ2(8R,?;!&"]!<7;/O0B6G5[,1?]*RIN:BB+6=M;?
P6SQJ"C/'4'UA!*5!_8F>ZG7+AJ3B.W@T^OIV%K[[U;:1Q^XC93SW)(4XIY*Z[?9,
P1]77X38#J0E% 2"&Y_YZ?D.,E9*7\*,@N%",?V*(&]PY:/PY[[A'S$,[*\M)\&W 
PLL::/1 D_)0BO]1R5\ YKEW=?XYC(R:[6"GH27RP[/"_#&_\K@VC&=M]W[*ZL[U2
PK,\.(30OLHR=3IKUHG3'S#-MD&J?ARK2S]^:HKN.*TSCFE>R*:EJ#3I>29.-")Z3
P)F<E1QX'52JD28T &/P\@'R^A^6+%=/3=95-I8MHS&\1=K?Z5H5FP%E]"GT5.)6[
P9'+V'>6VP:^5(0M@:[E9-UDP6YLERKD@W9/.<E^:=%HD/B9MA\[8@TPGFPMTZ9C@
PBR@)\/,'[JTRX;;.G;&J'V)**'U66*M"6#=^;K?=L<PY8$9TVV$5@\T?:3H5B)($
P&X<+<SE!7I' (JYO%R=^$C7"];H*C"RYV7(6'H:+? DF7GZ!:_J(#%#X.\3E0[17
P+!E#!ESC4]&I?B)'8T(Z&#3OZAI9NJMNKY]$JBA5CH[T@]Q/.!+2,5]!0;K@7/R2
PU]/^-!I8N5.3US]J3G4*1QFQ]^&XJ7(9I(,#+(5-<U_3>:V[S\,2/Q2!3]R1!S@,
P_HSA<)W=I8I'NJ1+W"QBR1AMG]RE9V!/QU_M<]TCL0-Y7XKRI9\<M+(BSVP.2G[&
PEB@U'+YU(-]0+CEV+X_@P)+]J%N5!&&X:Z>\UE/H(RZ()R_VD XD6I>1IRK^(BBM
P^)_@(,F<VWJ?=2G_G@_A5 I)JA[)PP#UF[Q[UI4)P%IE6*A@&8RQ&'T+ODD%4\U+
PW#,JJ'AW1F_&%$U@IF1MGBVK@V8\,DITOT0G3/X.1CCU1$8TE+#1<$_M,=-E,&LS
PW#QL3>] C.'GNM1-4ST(5<1H7TS=G#=\T16+2!\:^K^M(SR@&7+R>F5%.'=E!+^0
P47O;V_/H\_5'E8!ZPH(,&MP(7BO__36"(6C<2$+TT"/7<%7^*/+"9,O>=5Z$W4>'
P:J4QWO3HBH.*3E*#Z6W,LS!:K.+2ND]28?]\. -PX02!WYIS.&C@BL0Q' \R(^_3
P^ <Q?^K<[&28P##Z(*1%9L<> ,N#:9/I)*M8GFS4,B&>Y7([#]L[VZ ()7SR([;_
P8)C@U(C@_!.B@:N;WBDH6=;8!1FZ;WE(:X-UER221#.YC5NEGF+H"2DCI%B0"2]:
PS;@BWVFZ93:OU0//\41:X1WU]="D'"%?7@43R2(A: K"(-AO7VNK1(UT!=T-]_AG
PB9SHIVR(QJ=LL*W](6V;Z_!\G.P\Y$L :1DMC^P0%IQ79I"BS&XD6WE5D.Y#LY,U
PFD[)V=2I"TY M$FP+O&L=^V(/ME,F90EEVDQ,JV(=^I@8!,(J.G"L4A YV<B<2;@
PSB14<W@T/>/)^QNT0N+<(I(+5!\!_!&F5>8O7E:*F43Z/+>ZU>+<VU*:I\6!>?"5
PUB_- G?TH=8]::][$;PD%@[2Q["20]-G0=.(*E ,>LM.R>-44JTV+^YQ)%?8I+';
PNL9F(5:M:#"7M3+' YY<_R[G/WH\*[WH%T]EF0/ 4.=ZTK&>9%E8Z6V57EBMTX >
P<[:JF&RHT^[SP".O[<3;=N8?YZHVF]'?A2H9SH0_*U X?'I9\H+ D9'^#"'Z*XZ]
PL!>[/C.;6W.FHF@]992[!]6/Y+)IN*2\'0-F "N$D@O4DJ? (P5>QO0:O5:.(,]9
P8]8ZG8'GZ'8^0))^ 2H$WJF1I*K/H*M</92@)B6T)CD9FJ9AN--;W! #<#[8\0J8
P.6) T>U_7FLQ./;]X PY9:^+'/A,W5TVA>"20/<_63V,62KIC+)!>QUH;B?G'@3.
P9:^% $K7K>-E_9:C<4PASQ%>+)D1!)0 =F9GX#D_<SE<CY8M09;(^?Y)7FPF3C-Q
P2FS4!Y0(#&BWR+7NOA<N(FA@\!1&D56O,PA4YD);\5\*C18EX>\3*"+)<;254!LW
PH]+AM[%DWAP@Z7D9A3,4/,M#E>P"L@EWO]=RNO].R>*K1S5*>+-OXZ^7A*G)Q5YJ
PH#\OE6*/B:?>C9&\>6NXFXF4LLH!8S^E'_0 INJ]T+N]JMEZ45YRS4.-U@UA%I71
P?9*E_<_^W?G"1G9?'^6Y=S_%T,A+KSUZE9'8BP. _S=QVI=NZ;'F$[WX&$!=!3M+
P><$8)MN8],)F?NH:?!UG4SVC7O-3M]U)?J]GL/!&#O\]3Z9W<O2C^[V<=B#)B6-S
P2*ID'(J.UC5>63PP[/W_5TWG8-'JY$1CA8*H6R4$]IM4*4V@>0DK'<0,994ZL#_F
P?"=#L1,OCI-O@#5?B#2"=?M"(IT':]I%/)C40'M&^ 6^36.L[1VU\3^OHBMW\P4Z
PX$]'8"N#R/74G'"7)HCQ@O!/MXT:..,R;X@(MG'E,9\$O?$CBU 0:OZ'">B>5W-T
PW=F=\>W7_4CHIH$^1PZUYNZQ8R<T-+QNQ7)[0\9& +JMFLYSAD$S,&V%059 WK>N
P?NK<\]1W10(^2WG9H!QW7#?/'U,2FXG('A/&Y1QB=:+M4_$!@N6#J;:'+B.B?39O
P_M24YHF2>NYPQB&C<>8B^0L"A,&0>GCZCG+IQ_2-AA@[3](U. A!-_Q 5'L2$;;*
PT3VTY0+K9292*4"VU=[[ZXNACD?40\RQ\>9PG!4N#G.AZ"GH9;';7'5_G+;?JH%]
PB6Y^26'*J#?QD6L%^<CX667<6>M^^R.XFH@1G'ME4?=O>-N#!&^7T7D>&!NR$$(_
P#E6N(J.20DL<*STIRLRS+W^ 1"AAIK/[KR*(3IE#R8@8L=0K];B$7(%,XEO!^+6(
P/O]<2]XUFTTU:=&*Z '>P1L;H%*;:MH54'$J70X\2LJH@GRP7>H)SIN2BV<\8+GE
P8P.,9VGYJ>%/K&T\LE)(T'12HG@LBS2KZ2=VO9,V.Y#<^:0,@??XWU[0E($;%4U,
P[!:NB\':'=)%.G-O6!W0L&N\'EPI[5G:TUVVYX6[C@Q@)]+;"M_L"S?62MK>V5X<
P6>?GNU5NA,H_<J1#%V7RI5%QW8@-O-1LP8U<K.S-FDB-^NW8J)@^-6^"_.BZ0+HD
P?A8:(0\%W#_FR.UV[6_*4QOCUQY+Z[[MC\',9;[+"A(WFH!-STVY[/#\B'Q=T4A6
P1IP!A]42P&-8_<DMCN<OPP"K:TY1[97$'?UQ*4+_DHOI6W"\3]OX:^FG%*HA5[AG
P>D U(LVD2TSLG6 VII0L^SWCDPQPOK=D_=>5D/#CF$W"2UAD]J*/#G<.;U$O$HJX
P$5KM5I!,U:PF*CA-76"GH1@QB0U9N1?]^]:+7GU)@D.. LZT5RP'+QE3]T]6%NN4
P3"\:/7X6>CN+C>E$&@ZR0MQ:-XCH@#_QIB7.]"F4ZI[[ZB"C=A6^?XK)4_T%)@!,
P$1AQ3* :#S8IV-I1M!$Q =4FYE(S7>T/!A6]_Y'9S6"?8D7K>=\^L\3!O0:V9/[+
PZ22L2V9@?[_TAV\)&<^+ZT*0:UHS02MB!\&1$EN-[N_!VFYC_>>0%W 8RG:%1##+
P96$,VAB_D$%/MV2YP^LZGW<>KOW\[\^((1Q@+JR98)%2J635NOCS^4V<NC9W-M_&
P?V;'V5EJ_@[=].7X8P><,T&!B>.%TV]"[8*?J:ON@3U/,'(4)6,E> QW(<$U4 WB
P#,63>4W3N<]+J\&%RG-PF6CPQ%H(>4)%8>,A1>(Z( 4D3G,>_^6RPJD)YUK[>"67
PC1-%L9]F]A3,A5MJ0HT=Q#8W9W*_H7<EIY<D>_XY5,F"=L"U$9,/5?-5N50Z_P<1
PV(Z6L9F#,^C($UUKPGXOQ3I'RUM1!T-(XR'#FS=UKMMSL%0G.D_&?)J.36;AVED&
P'-R/21..6M-7UI'N1#()_#HPUI#B#$]U'%'R4J/=+X\49COWJ5@;M[S?NK[B^/R=
P,_8KC-[3@:[@41 VK:@ Q8\;L/='E#YNEYI#JRW>I<T5=ZM4*[D4M?X)Q_\_,[WP
P%0Z(2Y=24Z#YAUV 6V!D1\)RKEYD2B?*F"KL"6TGJMG>49,#2B_E&(_*[VY]EK"1
PQQOB]$("^%W4=$/C >?8%((4NJF&FLNN[9GZL<H]K@K;;$@X<<Q!?_L\9O;T$59P
PQT:J31]0$.T&\"6/FQ$3S:B  #C%^B,M$',C,/0%!E&Z]UM30J1.;[S17TJ9B7?Q
P5EVW1T^T6F-S(CZMHVL1%'8>+W&>OAMR87XZP*HR$W+U<C=!Q\/ZJBC-_>Z!L^C,
P/KSR^#637?V-(#I<D^[&W(#N_!3H1C?(T,LV>CZ*J"M3!!#S]U9CIG=G-?(:O#+P
P*8T*UC<Y:XPIQ"?<DOM=VRP8;%Q!->6 @> *@JI\?I+%T8[U'I.M@#3Z)LBT,D >
P'%E_H3/KR20&L$;$QX.^] >3)_EE_QIN,H?^7!!AY,?V[715>X&'%OJ7D+"3*-^N
PC[@D6Z.^"A\\,*7+L&8(&23@#*4R$8F,!8.?-?I7HT*@"WO>NN3=W#.8NN:9I$;(
P&?M(!F%.)37U?MWA'J0#/0TUT--2/(MG4/ML<Q[XFMC.P:4QOL*3EQV;K01%+8X,
POK*QEL9+FHP$<V#L952S>WK( M- $5EK8S14MPT8;5HF()IX8UT=&,!5=VO,.3Z+
P%0)[K']?R09[I\\*E^DYE9-V_N-!N.VZ69WN^=I!)#K(BX^/H+'K%(][^A^#I"@<
P(FCYI8;Y 8K)[U"4+Q["GH%3:,U,I52T2?T)X'HF+?."\XG L<5<M1K\:WC92F\G
PJMG_,U$B+/MH^7*,EUYQ:+5;4\\$*E5XUUJV44U(S'U/-X"B^K-4=#>?>?B%>AO3
PXZQ\!2(1'FNV_3B+K)I,9DGA !PULQ<"GP<H^;ILNV=J74IU9XB<(NK:L>A>UQMI
P-@A2TLUG/5)U 086W,DV+D[%<'"/M1O(P#\(,O,B[I;DY-W0B%O4LI8F7D[Y_[.E
PZLMS B8N+C^^%X'JP2J<P!VFG]C!H,ARN!,8_X)W=YFT!SK24OPFS<[N^[/YQFLK
P,Z6N37-&@5!!4\U6;LS8RJE=2"]B@#N9<$VB_!CT>D,EUHFC<2^[[KQVM_-;#!"A
PKA)DX]':U:#'\AC6!HPG!4W:&>!A2U>24X;>?3C5(JP*5@V996K?H:++22%(VG,S
P$BO>5N)88S+1UBROIH_)1S4(JS.)+WUXY9R!GI=&!'?JR00!F*7F10/Z6)[]J(%<
P,EK.\UXP;_XDS-B8Z=ZK&A"VG8H>#GR.URZ;'(&I1"#]FF;;E#8;,?UQH%O6\=]M
P=6C8%.S'IZF=WY1^^06S_ZM(TS[FG"91G.'.;%!I\.(JQ%U54<242&HB<6'2-&7J
P5/[@'!8:7K-Q]:CDM::0Y;68ODM3P?]O:\?AC3<C6XH!'[ON[PXNX+(7)<>+%E)+
P/Q^6"?Z05=6W=2_+IJDAE5Q!90I>'FEM!<XM0,;:N91N99\WOMQ\?.:"/14T8SHM
P=#)AZM";9Y%Z 3Z R&1967 D\<%Q#_95SX[FKAV66T%B;ZI+8 RW%&G7+;]")?#7
P03>X+IHC'_NZ5T+S9L%] L<5#>U1N0JY2,S- 5'69)UA6$0NE'-UQ9>B3^,/E802
P+%FHLIM3F7R%C:LAA?\N$'H!'2]Z7YH]#C:6C +#=M%7PD;M(<XK,+L?H%Y!7&\&
PVJV4-FC@1*7)\V,GTQI5(P#!\Z2T*\'=YD&%].9RVNH2'C)]"(LR[)6OJ+<4 @F*
P=+(!L30-'(;^%DHA,V^4-$1(D5KPR:-MN*M>0*MM!4:FAJFG0:O).RJ"R&YLND('
PUI%EZ]C)XP>UO1&2-!8/!1VW(:, *'IH<85OJ'^4KX^FWN@-#PR1.;9*D*]=0#[Y
PN_I3%P%3N9$(U)'>&%6,6X])G.A<L@9A&#$EQBK6S *7VA"\%[)HJ-IS>+USQ*/;
PZI\I3E:31+;.-6G6B:9YYQG)1J7F(P *2.H]FQM6*D)9?(4&^)..QZD))'X@CP)1
P835P<4$/JOW8 C1#F'UHR_<Q\-]M?3E<HA0IH!9&U7-H <IK897IS=HDCN+O8FD7
PBS-&\D*=FV1&8/>IO1$BS!9Y^@8!+=*\"V%S>.\PL]3]R&CAJA92@6QN?8AN-UM@
P,&60L_W*JOGYZHEK:BKXEN3()*\3T@(;3@;.5?GO=OSTY$ KXG36=!Y<&*M,;R=*
P^\AN""'P1=5&\BHKZ1J_.#!0/VNB^1$LZZZE_,C-OZE_.M>#D9H;5\7ZE[B$P*;!
P4*0J!1UYYJY 2MVX:Q0 L6(R@VUCQ%Q+OO/3\RV="O+8J+,/'_B!9. U.5L]D+]T
P6BO"HXD%F)" M-MW=<PDW$>Z?G/0/ >IJST9TS,F.*SQ:B8^FT&NF'T5]$((NF_X
P&$2!?J$>'&FA8M5@&:;^^?=_)'\-8D),71M0'=^VZC\O?7&9!2OJQ=)0"0V3C!*Q
P_K)=)>6@'+3&^L-"2!Z5K))BE=<'O^$\')5N" ZEU(96MC#RF6)LDP3-][:W*?KG
P U&[5R^NBJU$;O@+(Y4O()8[WN]VQ,-,A*U<>[>43[56B*]3G-C-[9%7;>#FRAGV
PR#J%!:FB'IQ*&@.ODU)-Y!4:^"R-.4;Z?68A277PN0!*+MG>!UJ,!HQK62+NH-5D
P/<G,?AF11H-0\8_->B] =HO!^%G"AMFZUH,/NS+WUN/KWF#R-1A+X<Q\&<HU;0W6
P:U$T-]V<;]!BD.[?;@_O#[SX8AGYHLE#$.;)6!H@U'K3RG?S4GK"*48&S1,!=_.;
P,>P@LTAET3Z$#$.;@G_/BH=\VJ)ISM)XC=;'B_+=%#_?O^K=@/NDS/+0+M\[D#)L
P3K!O&_D0VDL&L:&ZMOLF2P/1N_"[]5)D0QR6^V+7M::P,>NMVS>B$=*@EN%U#1@\
P5ZG>YI/!*;":@>Z>GH2Y+M:[]H[Y2@E1KT@M$<8MIF3V&Z2O>LGG-59K94=YWRI1
PCOW HV("F+"05:YO&YG6J08#^KVP,4$*9Y411*/##H[^U>?!_"-?HC9%Y#O@(*@P
PB&RWC-:9E_][E=.$$R.+ESHF)F@R:([ZAZY/91T*TG-)([*?<2JV;CO813>O3:LA
P\) -=N6 5P(Q?$OVQ#C>Q+W@T >)N&;QR88?WB@/(/ZM039Q0)$E+-+M-JIR%KD%
P0?@Q,&)_3\DG3:X,M.TY4!--]4-QL?(*^1,EZB1;M5WR-)I?C[KIL$QQ9W;*4J0Z
P?"OMX>Q[S&@Y$$(-MK+D"Z6'VC,:17*8_3L,/%F6'L[-_,:=W:[:G^ET'8!.SMP\
P"=2KW>UW72Z%E/=!+BM'G&L"T4D#O190-B.:_4,]G;=)XAJC&/BOP%ME1KO*+[!J
P!YL=6)"J<J^HAM"D1I"M>LAU,FY6\.$X@S^6&("AT8<3QH>;1BD_"I2'H@]+>H7%
P$YO4UDUW6TE>=KFL>'@B4\L;%#K;-^'W_,&W.OLMY^16F/%>EB,@ G4F'Z0%;0>[
P6\LO@C_(:0M3O FP?-/2!"3";OWBR]"% XNFI#NT[6-ES()ZCA0&KAI[$4I))YEC
P9F8'[4OT8"]DL?&[(7OU_#QPLW2P?W^"'ZXT<"_R56!H-MSYR>YY(52D2G/VI"(S
PL]W/3VHV!P@=#CZP(><0-^WSU?4/9+[X!1<@:PZJNKC@3F-JZ+/+4MH&Y51N+9D!
P7_8\2M1,"H#MJLXY?&L9&A!#H+Z5P^APBF:FT>;5EFR8IG$=UA7&-(EDA2+,\8V*
PW]?Q,GZAO,W&CUHQO/N*!YEI,+XFC[$(>Y$%\4D&Z$@ Y2?8'J4,=,0_ZG,9\]Q(
P@EA7N&."5P&',!T$ [TL:B:@Y@B+#OM0% GK+W:I+@X;N3N'I([O,6L-<UQ>>ZG@
PM%OS,6M.J_NG7A;1-86M9&7OBT1[X!Z[F8W6.*]3MPR2%O8>3#E1S">T-;QP&3(<
PYYV(8DAK7)7%J2RX]]87[R4106?:Z=PHE8CT*;.2_6,WL*=P5IFUYC*N*@?A.]IE
PXFO.:$6NAIT(L&O7/IJ&I?#+#-H\H4X70V.S([%T+,L.AN(6UBLHRS)JEX[15V%9
PP]>]];$_;# Y/A7Z2*Q"_C?Y42I9XW5KX8ADD3%@JLV;4P:(&=%W(-IV[9TQ_6 &
P5*(]QL7S)M-;)%D_ZM[UCQ:3#3.W"?=1?FT1V' 7CT21F6JUACQ\GD$1E3V@*%F^
PJL)?W85F.MS9,75)RU)G4?3P*[\;[T.F=^_8BHW84<YOM")A9PN,BH=<HHP$8?07
PFYM[KC?0NGY1;0\^*ZS@B)A[TR^LLK_.#508_>JU- (K0$>O1TB"2>TS'V]<L^,+
P$@QN?!]7)G'TMX+'SP)2-\R;1!+-/9TXE7.TLQK.S!]ZL5GJF# '^AP[531+(NZ[
P< !/8#]Y)/-Q7\\.R/2!P=K)L<L+8T+P/62$N\\,8Q7GA=O!F[JG$1@OS39Y9N_2
P6G-309--\-*9N0&&JLAK(7I&=WL1*^FOWLX[+).]S'VM S.'-_TE8[V$PLJ5#?73
PXODT62[-R<^=B\\LO1UACX\:XHLV1B^\<T_FD+ Q'H@GBT>$<M9?A'4]P'SQ4/5V
PZ6-[8RQ<0\8H'O%\ EZ!([03J(*F<H": :]9 ;W\?*0/88'ZZFY#^N)@X&O06A=4
P,;[LMLD!;+.1YZ9JXU\#TP/AW_B/P(*E/6I&U>/.\@E9O:ZU]W^T([WS#%Z+2=G"
P^%'G]U$Z3W; Z*9 795:Y-'(NDI*+:D8)'OA*'@JP7*[BY-U9'#JYVU",L) !SCV
P6,#F@2ME'JI9"QUEZ=-\PDA>'02IJ+\"KD<M*78&EU?YUA3B9*T"E?/,L-Q=+&F;
P_,++^1E3/I:!%HR7B6<V9AM^+\&]0"K8WAZ!W]HVCPQKN]RTO/3#4B64E,]8ZU=;
P&X2WK]PC91FFHQ;T"E^)=7VT'+J$SE"Q[7L (.6Z[H)SRFI-)-%+NPQ-E4@]"8%1
PL_K= !S3'A>.M?%S!G?N2'PXU0T"IJ[&0/$KVYOZB84W#LT;J63WL%)/\FITEN2<
P2=4R'?:TQPOZ;EV%^N?FF"_6*]5,@15U<W)I:F+WT6?A/F]5* Z ]S1KTPDQW.3W
P0,V%QNB/+Z;A)N><VN3<7RHEKRI9F_.92)8SUN70(^#+9-5%+,8FS!L682#X<M__
P$R%I><K5+@:Y)#X(JU[)H(-QY1!7S'LPTDQ"X<>5+:Z1]4N=[H#7[VDM,EP94NR!
P?H(V.!&2O00!H<+<M.-K?%'EC<)? &*'T)?C%+A-(^M!J4C"6@C?"B7R4W H%;B-
P=-R=ES]HD!NL]'_MDW*M6KK*.F,W:EN&%E\HWDBU=/3?E=)39$ 5?M]=GP3>C8[2
PUR-4R(JT"Q+V0H1M^$$NQHEXAQH%&YQ"0JP5=;]5=*<,;Z'M[N>O9D#=T]B;5RQR
P ^:NG>Z/UQ-^7,QX9C0'/8*3.%_3]51'WO0=[P$;V7"-O@(O@'I,=XVU)E?(UJ<S
P3T-PG-"N_L-T'6EZHX.1I5#25BU*]P;.)AUXOMZH>6UY5DB>!;Q4#>S"8%.8O_R'
PTZ-JS'YF_L<_WB@RJ'&51W B;J4HN<]MKV6C=8?7J-4S*<[W)S*=459+LZ&E=93S
P;0ERMY807KI=+*KX3G)I((J!#7*"[7A3%LT-"JJ$J_D59H;\+QG/82T:.WDGIK%V
P],T8(T?G%9Y(2SD5VVD=]9Z)@;'D6RFV1M36Q.6T@0-'U7F7P/I:[F,]2>DNF)MY
P%+:;6)<#XGK-7MD]=K\^6:_]Z);O1S-F0_M&.;*SIPMD?NZ4ZVX*?G3NF4=2 T/L
P,U(DT,1=U&C\K@IR_63[_EB>;E<X"8K4#]R][^%K*VU83:@E_1W6WHM-H$[;<=6.
PTW95@' _"J,5:415<-U!<LWG!(2U$\1(B8N7X:O"G%Q@#SKU*_R.<R6]_RVN$]:,
P"Q#E; >OC+R:N ,Z[/O-?*<SE8V19PQV[TU5/G\D*D6D"_]+R[2\"5RX3EA_A/43
PR605[]_ XFT7$LP>1#IYD)FBR<G'\C&XF)UXE3#Y:L@@.F)E^$>^F'Z,4V"[H,O:
PU?,.-;):J[;SZYD&8:(1.TSA;4'HLKS#?NHH>"0?QA =6FYJ22K1=>%K_CK7T79W
PS?_""!Z;.(\)A+*A,YRTF):"1@+795@]7O)U6ITE>4<N'D)CN;="V\ Y].V=VF66
P@#+C1/M '7U@B14&Y8LCGNQ^$?-"NRKNAUB?YETYTC[MG%.P3;7<.E>)[\L3\'ZE
P4=S3A.VOE!8"!3FM0.^9['@Y!BFX*##] DOL)_)Z[YQD!K$-9*D]2;!83SG][2,S
P !]5$^)D@$3Z[$H(:TNX+/NI(=7$_0"</RKXY+==[PT; $I4_39690]/32YSL7E1
P)IO,&NX>LJV#70&"OO)99;4 ^BBY%+,%+ "+$9>\QLYW(TS[Z9()Z)]T,B5T!J=O
P:VT_=ENE4P]=++Z!V:C;_8T=DW8)E8XIBQRS?YF>(K:]3PGH '*(<S4N+P>H;1&7
PW\=/J>_X6XZ1E[!Q; Q\ "L%M%-6,HE+7*HN8:,*^N5D(E@@>7JE)Z]-\)4"S*B^
P6$V(E8Y!KUYD18,JCP+2QRJS888H19#?DA*%7:2EEJL8EY:__CO,^XR7KEL\WS2W
P*O]6DJR7"J5*R/.NOFADGE(M#1!BNZ?4]IJXG6?<W2%B_-J2<N\0W#]O$,KZND6"
P'OX;$T<0U5[B"ZH7_- I%)F@N9UJE41Z.6++KGA&+@!U'XJ<'EZT8C+7_=?JWO[!
PF^6@<+&$1$+I-L7!R=S@P'^%:JT!8])4!U@4ZIR=@_60N\$", Q&\FV43&G]9,U)
P+.TS8H$:YO.B^7T%45&7^*@H/P/:O6Q!;&$OK&%2]\)I*V])^*"X6CQL#*'4(4U#
P7G!M<P&3M(/QF9X'GF ^2Q=M( %T8.,\"Q*? U"'S@\0?P^ITK*@;PO?M3B)BC^<
PK#_U"<*+'J;O[LFT"V"G K[ZZ$P BG^KFOR:VYFBPZUA(^//&#<@*(W2F"Y_<-+\
POOP!;C%A^63)5QDI[!I3CJZ- Y&[__P6PD*1J#: ^V;4M-(C&@F?Q18]I1ZJOMDF
P+G%+O-]%:RX<H$&\5UFD8591DD*/ZTE)B(V1*Y#C-IOX-'I*9\NOG9.8@H4"9E-B
P<PUO60+,"J2Q*C]0H8&Q5:OD[MJ[V56PX_3B=214\E]RY0+KM<W&/6[0HNV11Z7#
PH9W@1P-1)'.)5-7-=H)OS"X4["COO-HM3%.%IDSCFP5#_*ZWBZ_L>!G(A_&][5IO
PSHSUN\4M@,1IY)"U[[]N^<XZGN6J[6'H@UO_'*[08#;QG:.)>]1[UVZ1GQ-';%UH
P.@O(A&8"8,"KS9(_.X1=@L<<U;;&+-&1/>H56/R .+%V<GHO*Z.CG9-(@!+UXJ>F
P>$@ZW9'@I;+%NECQ7%.[?L!BE#A*3?]:XC1.^Y,*@3PFDY^]!>S;)@]E04%YO2K&
P"ME33)]H4PHFI"O>PL@:DDLF;CM4GCI&@_$8W&'BK^B!V39BRW434SFKH((2LDP/
PI0=]V?NTX6.,3AG79,)=%LN4XC1AYB0;P=_&#2LH2KW>-REN/Y#GS!+2K$'8@64J
PC23ZHH\3NV2O^]@1>]=X#.9/^0T23*<:DC=X9IP SMA[SR8:0_)\.?ABP- K(1 "
P>.VC:3P/..IFCF-278Z]Q*NZ=9*R?5@0 L70HG" 'RP(@@;C;)V=)28]G1,3EV2+
PXLM&KC\ZM%+R*C*(?=ZF@N$*08:2C6>8$ 26OP#1ISY)D[P6-F>6_;<OW=*5X3Q^
PM4QJ@;HY5;L4S-*4/YSSO_]1X_QJRPSN3F,\FWI"[&;01SB]&9P6+H \+D_?5D"S
P)H&#7"1!/O9W,T8-0VSA4[^%M0"RR]MH2A%@E7VPXUI_M^G5-I#21;-T\]EX%%#\
PWA6G3&W'6WR=&XG-_HY=7\3<1.56<,&&WN9YFO=JZZO5[-1+3 /VJ/6ER+!<2L7@
PGT\XOG YJ$.F]*5Y829Q#C4\NL7N_#![ &)A>\]5(VFVR[]Z;2;F<OE]'-,^?_CY
PA-[RJUX)O=+.@-9Q>)));^'=@\H8WFM^1ENM$S^=H>85>2+!R+^>9]&>8U=8,NY\
PTKT4^[<P:MRROU*5QQX=&]>!RAMH@''A<(]X=]3\3:LO0YK\3JW/L1GO8>_.VBJI
PO-3S;4(,F6XV))SO_(43)&*3UM_3)JC!JK 2I22:*;YK!'A>>C8\ 6-#W^-]W&_H
P2^0IW?!9NNB ?$$@7^_Z_B$6ZLPW1@YX"*3T=>@QGH)::=3>DM%R'D/0A[/I9_[/
P%@TZZTNA-O[=$8'*E.I314=?7B?L[_:QSX&?NX.5^%33#FY=]EXZ#9U>R>^ [&Z]
P*\!=%#.1S&'M<S,AJ24_T=^[=^XX1\0,H90(D&D.$3LM@=9[ZP!5LZ?<YC Z0W)9
P9DNR\IS]Y1F8],7Z(,88R1:!BQX%[-^2W99,=#K@@JF5A0S+T%PWE'Y^HOH.<3=D
P+._C\*$6EJ2TUH+UTH(+$6(7D1;PPF7W_W2+:GTO7$I77\I1W*A7WX?66 ;?27J0
PBH;2(%UO35:F^#=Y8.T,,L&]7O5@XV$+C#=WF6AIV49L5[!')$R/Y3@=\PV-FF%P
P/CO,\_^=@LW8!.LQXAGMC?:R97UA1_C1%,-Z4+DEV0%$U#G[OI_"9".P/J).><3"
P3P.^*U''UX3)1&]$I5;9WD4N"FND4WJU]3AZPXA%\:I[&"?BIQK2J<Q-S/08D)E0
P6E!+NQ:M:0AG!;>??Y+6Q&DE4HRC&\=CI0*>553\(EYAD/X"_^2<2EGJW]+[%[3Z
P7_Y9XX?_J\J*\M-2NY+>2Z+>RV?'&TX./#=(KO-)K%$V=U#4@P>%4ASFVA&.B$("
PV@1X.\I\ _P#NSLLHR?KN^A3[Z$#P'?,6 R_LQT"MO:E3E$K;B-W[F:MT055FAH.
PM$*+<K'<\04]YI)+7@*,>"XHG*SL>5<"(Q<SO5MD']_#5-V'U!2EGL!PU]2^4[T.
P%W"."G\C,D%C)-QE8*-1U(9]SU\FZ,P"'FJEPJ+CR%"=1%*)"5YO4MRS&J=N?*/?
PG,$/X:YXOMO6-ZN78U69E'!H]_CX#Q-+OY=8,U75Y^&CM<H^C-UFW5)RWL\HY7&J
P='"-YZK4V@%M;J%>G(&61@>9#V%FD9:L6M*+G_:&M;<;RNR7R&UV47A9B^52)N#H
PB\?-O+Q$V6&Z$(K.$73V5 I&4;"BER5!=.A;Y>93(<OGU6N8)]!1XSL(YJF1$_Z;
PG^]-+0>W2?.@ND14M\$[(L"O= :KB3&>F?1+>=A:.6*/%9?_B_<#+\._0--3TH."
P.ON%Y!XM-[QC TYVW#@L-EN)?@"V$Z31T"Y:,$/5BODWH]J7="9\S;[#]+ V)YY#
P,*3>:&@_+WZ8?J%J87/A)ZY-F8[NQ1:/OZCQ%R9E4'!]5W9W:MSE>.< TL\^_@S@
P/'Y2L)AM,K20O'DL7H\ 5-4,8/]4G^9)H,V\O2@\_TF'B2&RDF*B#H558.!;X7?D
P?)/"-\Q-ZY1:X@H$UR 7ZIC!J"C1&]/ :,$#A&NE7IT"=:3*P,I]+(QZO%#B*FO:
P-E_FXRYL=-CD+LJ34SI6!;HM!&^;EB&6.II [GQDT=ZY/&_=X_I*Y?@4EL-IEH61
P>QHH:T7%LH=!@_SQJ"E11W%1#HGA"8!P'.E/04O9[1YJ!.M;;GT;5O@]O13/>F%U
P^M!]:93-BTA+M:%0@!>XP>+CVA9JU3#G(%2H-^CE]V@F3UR6BBIHMB<! 41R/:B1
P5[I$LM[@+47BX"/',58%R([MAN2^U8!TT*BSU!&HY(7,!?Y^86I=+?E:;Y0=ZZZP
P2*_JI2P;A<'3'7?X8:KL+D],HMF#W O1&O+$WO-+WPY*K-KH]?"?6 R(H.J0;L>"
P6V*6(_*_&[?1GK;Q,Y-8F=R&N0%I.T&8UR!2578T6<$J+38RV:1QXO]/O]*Z\G"1
P;!PGWCY!Y>S'-)6*0E(/2V\7N <\)C1D+LED8!V1[?]-"-5$7Z,I%4+]4U(^K),Z
PIR]EU.OE2NE-3X=6Z>W)GPNS3VK +7:3V;I"0VW2#TLGS1JGG^.!"=L@S;?\'D^D
P%OP,ABOT/;I5P.!0A@?N#_ ""LU.GW^Z%P\>4AV97&V'X=$7)G2:':1>."#QJLSA
P.#$EH4>&EU_62.XY@=YO>$FA/=QJD%6</ZN_==OWD2WA M2;MXQWJT3 B4V:"0LY
P(E/V$6%>[B])LA*Q/^1E9;U2V3D$D7N=ND(3C>XT# R]H12M#9>Z[79=_":9)C8?
P<I*K4,TX.8Q5Y_]"^K_T0]$=SX4 HCBZ<4_.=P'U\*OS;GA([R6_\]CW\N0$F50#
PDRE3 DYO&V4JU[@NB'/Y]CW8XY8?T0PY-[BJ99/%,I!<(7 C2*1HQ\[ZT,#FYYHP
P@+KMS*:7?.I379@3NL'?C9@*FG49B\=1]!:([$\AGCR;D@M8L=GE&S&.TB/F.4-2
PEZ0$=;"[,=_/OD[)/G?IN_(GY5?I.2-7P/B[2II7? J\TJ0=./E"XEYE#T^ZF!M_
P-'XQBSX7^&YC.29F;092>FOTO?4'C>3+IC'QE:$>9CCI&J8"$^K58N^</["\<Y%#
P"-'#E%JO/^. ['*1_E#F8NC0=Y>YV_G;,IK<\DNY8G6SH.[2KZU8L]?M8@'JB,5Y
P37;QY S>3ZDQS?)W)QIZ^E .13_:DN)MV0PD,622/L8_X:T@%J@5L.J:]'Z0DSPB
P1[3W(S/5()0:8M2-193N,L?,X7\=4P'X2J?H3Q6C6*[9_C@VWIN0R)DSOS+J_+;J
PCA< 14<K<M66GA"Y83^UIC!<U1H,;!1@.PAO/8TT-</_FTEF=[3G6, !O=XPX]CU
P<#8AHTIA)1_@J*.7Y8&YIF+ B&/>"J,;QMWH[!G)ZA3!ZIJ4K]L! Y'$//C8K0T(
P0O,[L5P<5N<MD$&I6EG"M[,W2CSD,+(0K'\(R/9G>]4#BBB21,AX[(W-3'<'^U![
P2Q#G@H3/M(S\B4U#)9]$U,](AO_0=@@4!Q01(NN@3XY[T3=5B0QWO; 5"7(#,F@@
P$LFNNM*(OYC_7OFO4157#<92*@2")=$>D:G,4)C20#SCRD[LRVS6+K8--/MD"2UD
PFL!<_<F(V+V'P1M^E3LQ"\;'FZ_? 0!&S*TR'$JY@1AV!\"'QI .U[*OIW[9>SP6
P(%L_M45:1EPS ^/B>6H\EE1R?:HK[HF=%V)8B3T^47H/B%!>,"7$<5^["TF4WS@A
P<4Y'WV&2CS$LG\6"Y*3W1N87;SPYXY'-HD!;_V6(C'2CW7X'+YHG^N725SBI HE?
PABC15!)Y1>*[B,X,AF;"0L4P;Z^C_/0Z#"@6MLP&&FTPLG OS9L9D=$N^WUN3<[8
PPC6V>ZJ-D!W1XX\^:[+""_3WY<KF$KB+EG:,X:>R;U1E:,68X)Z4#T0#:_,XY0^]
PR&@B,Z&5J*(+M:R^ ?S^#?!2J*G9DA,R'7-\"4W:AR9)#^34./T#.YW+>HO,W8A:
PM\(+=DUW$$$:S*GLA.Y>K@HC6)W(RR-<B_IWI_$WUU9;W?2.+1VAY_[9]T+EX/KS
P$G7Y6&>,SMAFCAAGKHH#/^.=3E-0-FGV#60=[[VL["UPTE.VL9(U8<\P:5I0A*CZ
P84=!F4U;B6"@:1!;SWI%$PVD?.MWR7]C]7%^;,BY-E^6#K*+(=*^GM1BU;!&0Q&@
P"BZ5=8%89WV\]W?[=.GZT)!BQG)(V 9N<U7-X5'*A& ]=JY*F_+1W6:M!6][)#\/
P2S+]["H.A[&G/^,=$RYD2O\FQ =_]N_'5:[<VJ=VGP5][4,ZBRX*&QMPA$PKJ!,%
PYW@YH6ERM56$H<*LNIY7V2VG&($L[^V=@+]%O8:C2B-TADRE:0CT3-5+,.NSA __
PDS+[@@OBH9<_0?=R(P\T")GD2B(B7O7N.*5@?&L5/DU""2IWNXV:;K.JL%/GSMEA
P;L?WO^6?U$-5R^@K8_N*%IMS%(;O'Y BB+3O)?&[DI([?!UA]\,%HUO;L]"2@4SB
PT[:1=\LR)FA#MHK<K[#2&WV-:8NF>Q/'@F$4"R$*?8RS[>F5:_3E>C+T?)99B7;^
PPB#NXM%)I(D*3*#GN 5'Z&N9^&]"IV'F%E@&DH5,PD[KHB)R%;!LR2#=4PS/5>G1
P-L>6K[S#2?33?[]& 9]=FU63Z ZDTAC8-KE*4=JT\<9Y!Q1V"-V<X5Q;4+7><ECN
P_!X&[<JGUO=: JBW13^*,'+#R648?[#,/CW!9KZ&[,$Q$FE4KOQ\^J"%:1VN;)_O
PMXF%HS?Y41":P!2&K%581XGXB?+0BBFWG>! PJLV9FEZ[L91AGUM\>HYD4;Y8E05
PKEIK.^OOL(Q(  +8CNH%&BCWFO:"'!T*+.ZM#F&ZVV)6=)WFX#)C1^H^Y,5[)#2<
P(QZ_0J6DT+8[9@&ESV_N!RH&1_43A*0U(TWT!C@149?/7 %2*@ =9M'PZC&UX9/4
PJ9& '+P7G5@(2X0'380CF$(.ZM3:/_>481A>-*3.G7+!\W^$5&,^"/0B;A,&^3N?
P-Q\XN&3G_F65)+ZIUT3VBLIGJ9(R&C83CI$,2>]X,Z<QE^O=1TZ5:!4JF /5-6[8
PQ*"HIYQ1_CZ@MFJ+,]5/?#K 9O0GV.UN21C91P)2F:=1:6^2=Z %>;U"PL57?VAB
PX2&"+5^UPJP="4FQ*98P]3*+\<G)2T3:V@E>&EPMBMU&"B0TRWW-;H7]*2&68^<4
PTQ;"-""IZ4X=RX-U-(T[) <Y6OO!E3AJ_2E\<!HOGKIO0*"CXBBBH+I).&"SB54>
PB;E;=+8Q)6-3%!X!:6:J&4;42$T4R)//<?1BLWLYKOH[T?A#S$@ )BJ"M1W.[S<&
PP]5^,;=*+W1!V@?=!Z!NS\[0'YR\%$T^:4$=C$ ^^G  T,Q6D[&JX,2][0=J+R;?
P;]V>W Z?6Q(\1?5@%Z?T11AUS'+I\HUF!IJ/33O_43)8YH%A3Z6QO6H6C]^^3-F9
P#J<_^\Y"/,#VW=I%&&VNS&FZ8C#10%QC_,#?*']0G\Q(-3NO<'8EE;C/'LGG]O8(
P;9")6Z[H%$L;XNKG%IZ5=2<BILI4P"Y9@(=7RL#22D^P+_S.*=ED-@?25\98;J&:
PC:[S21+/LW(IH"JQ^YX/\PJC#5 YXLT/"!K,"[QBLTJ0:4[[H+O$_N[_MS<S+%O'
P_VM:IF!^=$37O&,?@"=V8(#=!W,![0$MOVZRCTM?O18Y1^?R>@P9X]O/YQ],+A78
P8VW PO1")Z5I$MDLD'41U6X-@MZXT.C1IW8L\C ^*!^TLD<WTFLK0\%02I[ER@-,
PT@S(E96@<D;)CD5NZAYE^3S*2Q?9<>%L%EQ4 \VA3Y^%8?9+_2O>^%#HIT'IDBCD
P8VU]-S=@B)P=E3G+7OI^H5GS[$WD3(:3I!E>MVJ@\YZV&JMU 30R'5"%O"[@C,#B
PY4V)H4*(18D$5AC>4ZHU^B+2?"NIZ2_^.[-<_#XF][!J(_)EY89E.I]Y])5*Q_7?
PW$6L?W2_R0.O'88^456]120.'Z9[LI%2K9Y)9HE$'X8=I:LJEC4$;S\N]>HX&?$/
PN*/<E=\:/SPJ29Q>"W<]SA:I!1K2\$+S1W@?>B>1\XI><%:$V<U*/X!GTFY[.[DP
PWGP,:6$6D69XQA [%I2E ;V5LCF-VOL,X%2<HPN 6N4J3GEUOC,6Z(-]'[W(['@*
PJKGM*>=Y.(!U UXZA1G$EX]*^,\/=$S$QNTE:Q *'=]S'YE&O52)SQSDA0J)[+Q2
P2/"5IA^EOMXW25/$RI:NW/%(9J;?3*?PM9B[3$9&:_F3<VA:9_&IT#7&N%HL!("\
PY#<)(G+F"UI4M7+W/J5Y5JW'.S>T.=G@8U2(0<;VC7K)XC-WHX\^EQ&TLH( $Q++
P&5C^D6[?#9#)D30PV8,T%O3=M,Z,D?7MA<Q0L-(B#-,:1Z0K\;2FW_IE-+.7LB2@
PIH/5DP0TMZUL2I7@!H#SXW0*W71V[6")C)EG^M&1%>'S5P@)C- K*_#^C&S)"6$-
P&WNXF4RD?%.@ZMDS'%1=_8A0&CTU3("&1A^/*["K=*$?*[/NMD2*3TC6LT3$[1[Z
P9M#:T3"L<$$P,G17SN/\I?VF.M&-'\*]Z;K%I'WUB'H/I-)%A,R'D*<\&\8!-\YS
P8JQM$,W[> B5EN&I<157 G2S@]V&^):OF5&KNR[N^;>._5 ETS07BC]F/9=&S?))
P=:^!U-QKG3I/OU9]/GX8X-4=3U OL$9VQS5V@EC=T'@C,EE023!2[$>#5Q2)NS]%
P> JZY].FX](0PPU]ZW3/0SAWBDU_0MK<Q,)4Z?GIY(351#4K.<,\[,U_^M4(2][R
P)\<G-KIG;Z!>']US5%MRL@LMDE%D?-K+67D#!8E4O5"^&;KFH"XT:RZ'V"\54<J?
PY3.\'.]-."C["L/],D[3I4>]\LFO4(\;@ES.I,@^)YU8=^/DE_U9X!!7\\RL3J(2
PF942Y5E;.;;.Y5ZNAXNBYR[.MEO6T,R,)/JJM0!XM3-10G>*GVM5?]"7GL#':GY3
P[WI+5.A=;([?6]%?/LUJ.XU23>7-@X770^'HI'JS^O,!(9W(CPDPMS7G+P^->K&[
P^'R=*M;1)%KL,>92+=5&J!HT6QJE6S$+X_H@6Y.[E-,B0M(4"FRF?(!4 ?,+WC"!
P,/6Z-1>#H^;_TH*@&_ZT17\9_%@O/R:\WH!YJVJ@'^&TH<Q\^@$]X]DC#@E233WB
P7:M55Z:WKITHIM+OA1AQ?"PD,PO&A:1W-(P_FR"C;Y!OQ[53@>>50YRK/H3VS[V6
P;W+#6YO.YU"Q<=S7)5N;LQR^_J7\D2SX9M8BP5%$OA&E0D/>BW1/O;+TVEQ\%H=5
P%*>-!%U#6C@\]M"ZU.&M>>N1SE=,$MX'/91.(\7\FI=_V0?%0@+$#]@DDMAA\I%S
PB39MRO8!%J9FEEIXD]Q,@>\A2U\#F:*\ V9_ $-_# \4DN0<C3P_6\ULHUV;FQC 
PI0LD[BMXJ7<6PO#J$SN.(:5$-IMBA';K1H01" '4<7T0]9N%7YQJP?9)4W4)&N, 
P!W>AY-$ 16-=]^R7Y(?Y?VWW$K;;'Y-R(;DR >@>H'P TZ$R4?FJ.60QIO_$6#DX
P6)^<N8T8740U?\Y2'O4V7HV[LTG.@)?]W^E9^T!OYA)P6SWPX3$3AET&_=H!0J/C
PCCQ4<B*4:L>8"]DE*/L+L,];R9 MXQ%A2D6*Y-;[LNPV^[Z\3T=^?F?3$S]%_PI+
PP8/:EL'U'F]5::BWKNY>W! ;"BB9:Q"2=U#6?<2\ ;/! WJFXG>A$]$T]M#E\D&V
P%3$ N//KU$!>'?#C@C[!>&U-N&]CM>1;V^H/VW@>QUPIG?Q>EW06!]].>8KWJ].I
P(!\XB#=YV]-N+_KL "T)C+63J[L:SE>)G\SQP+C6 <M>2*7:9'J;%ZPB2_7^V4J4
P@[-)TM:#L7:G)?\^4J-TD)#./&Q-%TWUL)6?DH&;7EJP^<BU6]"NIPE'3P(MW+D?
P@OTP:L%&70 @]RT8HA_77+$,M@Q]/=[%>GL\AG^ !\6V><#400IZ;%PFGO/DB.4S
PE%OF)O(T^#VA;*-IVW%K5!3DE7C/"XLGPWYI%^I!M=#@M[%3<ARG:9=99QKATN#-
P8=Y_LT7'8(R3/_<FD-.V*',/@(6,N"GR5PI/K)Y:Q+JS G?ZETP@\JGXYP;*@LQ#
P5<?\U4P>HH8N\HCAT9#XN 2LSBH2RE052%,3Y(H'D[>\G8-78P[S 2Y2V+<O9YE8
P,]I 0Z6?9M*D1M9Z6T<@LF^4.4=(UE%"I$P ,_9I ,$K6?!OHP&4?LN K0#_9,VF
PJI=;M3G9O-93D<UK(+U5[;,3*K7V&%YWP<6,XPPU)0SP+AY^OX3@EY5BPA 4BG=^
P?SDL*=Q5Z#WWTH<%A>IV9;C X#%2\P5$A&#N>[5$M=A)P$7NBPDCS+N*$VS&^F7E
PD4+:HC2U^3Q\*N%QJFP/H1S4PTCTV'I3FNN9)A&B*)[CEA/=ECL(#6YX39606>VC
P="]2_RK^-J06&>U#5M2DVV>*JJCBBWP)Y$?PQ1+%5N^!M'?%L7<\]Q:AQT"5J-BW
P+HJPKF"D+^D?19H%*AK#$&$FK <USP, 8P3.B:L=^BP4KF=(!AR[.]^17^?*[K<G
P'%'-6NQF)V&#TWB((R-@\'#)?I?E:U?++A>P#E9)HSBKV+C?;5F,SVD70TH S1I#
PPH?D&>S<_26N *@T;?ED 9VFQ!;" /\37V/@:B])1#XPEGQ"K28NHY(M>^T:-I*U
P:AUWTO<Z%=\\58G7#<RI93A,85KZ12H/2\],^(!T7-TA94/;>Q5O?7A:UR<D(RPT
PL_/[.#^^GUZH^54SGW>XDWN4,-#R&E#S;[C1J\O9,9'5Q%QH71^+C50;_$49D5!3
P#(A!^NHMNG5%R6*GE.;^NC0Q+MFAU^(][()5-U[1\P:"ROCV[D.)]&DL,)4D((%2
P.M"F$0_-X;[%&!/FY2]HPO5@>-<H+^>?939&R.:_VT*W./2-\$UVWE!;,/>G5T)U
PKM+_$V5+>Z#7\XEQN]! 7KL(9-5L+46OY(ZQ??!/QI"P.SB?<CN0PE 96;7OJ&F/
PHQ:,GR::E4&"XR+LQ$"IL/_/W8IQ;1M^KCM2P\$XC@13A"IY*8.=XNFF?K-R20ZO
P3$&_3:<\D7  ,5AHEW'Y&FNU_CWOO7_!(&'(H1O<".R..[O+G,U,!7J77#S0_YFK
PX/YR9^6%5"\\#^/'F2H?Z%2U#%"8RW&5UH9-\3:1BX63AG&2LB![\A*$I3^,SY_K
P.F941SH[[^TG.P>>:_&:57;+Y&E %4^>U*J1EYQ"P49_S^< ,3[.#2GW0G.NS#(5
PQOD%7K:NQL:1L)R'%$8(WW!(&V/(AU>NT$7=DE(?10$:5^[-[?I-.T*EH;ZK?3!=
P7LMA-"CPM<6L91;!H2Z7&9V03=L<+9*1%92"F5"C1SNQS) I+#V*#\<RXL#R?R.2
PZV_:J)!KW]MD1[@^V_!EBC%:-!W&N,W 1%&3@KG='N0I^[8V2@!'EE9"U#$:P.(K
PZA[K[YYT(R@W<;VZA@Z]8FY+D0/&,&MB,W*),N0K*N-#<3SO3X=:R*X^FUY134"U
P=141H10C+(.LC!M>[JLS8 OPICN2=TA]@%@@+2W["L<A05U./,FU QH KQ0<]"HJ
P]A=1J57A/2Y7!>RKEM_C4R0"!VU17]7N5*X,F:Z#-/;?<:@*P/8X[>JW/Q_M-/\:
P%&B)Z(+*=%M.\3>8+A8W])O^%>U6WG0?9=KEF'8+>GJY0P5.?97E-4*_PW12W?.!
P=DK(BKEGOP5M[%BM4;R.1!X@+:&".<D<+^;<A6OA0&UJ?M&_OW&NVLX2J,TR_2+'
P@=6LZXBZZ";0Q:46:6G7CELC(9$3G2!N%FU/P+<=->7^.1_:)J$N8@?./61E\2&<
PI=R\%R;NW9QSQ#'#@HXB;,$B+D7D09/6AN0+K$)2.G9NE(@\^M.TOI6B9\$()<%^
PMCQVKBN#/?@AQ623CT)RA#^ENZUQ2=C\#6&,Z'4-[<J=06<&HO_LG0<Y0B,RU$C1
PBO'#_Q,F3M3YY#&685Z>H[%0WCC4# TD@RE']I]T.E>!L<H24QH*>Q5+1]1IA%1%
P"6^&KJ:LIJ!FX;KFS;JN8\MB"E-+116]+,2ON==3+)&_(D2,B#IZZ/W.+-0)5:CX
PI5]@ BSU/4:[+[>*XN[9-8^]K+F50Z6,\!QD>S-NC?@,=81-_6JPUNB3SV(D"N">
PC96DO]U-??CIU"NN6;9L^W\IIXM.=[B,<@&!CSY%UOQL*'_AW<GH%H9=X;&K[A^*
P;.GLAR;\R;?3RD"_:D*-O%Z+(PG?)QFVS.N,AEOT6:H:$ GB41\C=(F%$WFSX$68
PMLL>FRY!OYH3/@059ED6#'=(YT'Z9:;0D<[5G;LHW <S.27J\YK5C^%%5ID.[L:Q
PG)70KRC6WY49M9Y 9'XJCCU8*UN)@E.!:<5IQ)6;^H&7IQIKWV+!\;7?$%'$7BU,
P?GI:8NQ-/DRS+3\_#+)N#2R<@1S%(*&%-7/).09.Y"N";-LVUJ5DX^=QB ;""X-G
P?L=F>P*_U:WMT:VA W.[@(2Y\0T0=]/9;<;\*(Y%*BDFIO[K>1R,U#EEDU2UVW]W
P;LG WQM%FP7;-E3@&MUW&G'1]L8@S/KM;1B3)8./'(L]Q  C3]U;%I S12XQ![K)
P@ 9@$HUMA*UBT(+ZQ-19MAJ;':%3Q%OD9^!^ XGDS Y0^&*\:<D>%?>@&]:J5LBQ
P?*\]JAYNVJ!&MX=S1YH;UYC,,T#6RI_J&<@)X41Y?GT>F!W2?4(IVIJB/7MWC/R]
PD[4X"\9 L YXN:/"-F:N/77^9*)BWBJCN_J04L*]5P# FQ+F^!RD2EBR%*LI<6:W
P0(:[Q1E'^#PD^]=;$4T5P$>M5.2Z<P"V*? <1%*& %T_1MM>4UQ1>%V%!^^_VYT2
P3<.50N'B1]WO\=:@S^ [,%Q@YAK_;@<;'T*;%PHV)HE.ICB_YJ\.32V/JSEM-;2.
P'0M;YC-^FL_N4SPP?<5!8S[-4 HF@A5L%5SGBAWB-,;RNQS3"'$#,"PPH3A_BHR'
P'(38.P)_9Z/VEX!SR,<U<BF57-MF+L*#Y7'GIC.97>9'SD@H=+684^/2260'6@PF
P6RKJ^EO-U0TY9N@/^MC(K'2"ZF8E?(LF\^G;?I+<#51[DHI(Z4#5>H2_<8W5\%\I
P8N+?(62693"PWDO,6(0>3*5H ]<U^Z-!+TI=:KY0^ER)XD%<HN5:A!M0N:KH3):N
PPC%.170UVCF6R)"I0FP6N$\3">M&0N^(\FN 2$S-&@NN+?.!"X/T P,":0.FU)[Y
P@>&86P^J,Q0HVP6_Y.)2I6'XGC R90B];\_$3%SD;.RP7 RHD[#\I$48YE"MV-[J
P7G?X!P-TB#VV 9Y$Z<T\G_T/'1H8+]+HW&AUP+ZPGZ^G?(:QA]*,&)OWCLJ+8(U[
P]'+SPY._$%X'WM]I*O_Y#(T!<@N@ZFM!*.!.;FPRI9JIU$X&AX3Z_LGK37LH/(.V
P=-P=3HJL(CU0V;%N6-ZO>&2J62>8DD (K:D;VXK\XPJ(J[P.SQ&NW#_5J%Z<<^9=
P/(@4(7GBNZ"QH*[,6,J+W%C\Q$VL"GREWJ&EN3J^J]%]>\%3XG< P)D!>J?FPY&E
P<06MU8H#7<2DO51VD3I0$.TF9\/A\?5>WQ0 2OZ:P+\HM'0Y<.'[/5\7E2/A-5<M
PGP6OMW2T<.QEOXG'_ B;_]],8(4LDA&5BW6'G4< U#P?*<19$@KWWGPJ!C#69:HI
P$M?F?<ZHQON)@6RUAUMC][D'OU%DQ <BYG",0 ;\'3E0L\>F=H6"M0/E/H]GQ03+
PN%N2)="K7D:7S[$OK*782**J-)(5*1/[(R@.R'M3$ 5GQ'EK*O=2E@_9E*904G"H
PE=\/5G&@#6W=>-#E#T7^]F&ONT""W_VU5;L($^NJ$2!9>C1BJ5$8S<<IF?9@5:)%
PAP_(J<EG5JA_8(5#I=^VR<'RBA1!5QJ'3M^S5>$.<O=BRM,J!8,A90(S@-K+/M.2
PL?>;;L)OG\191G[V)L2V_ILHR^/5Y W,A4R[VL4O. TYZH5T7H"-4LTVR.,H89'(
PMN17F>ND6CY'I]RHCN4F&!B-15 !XRA] /8KS]6"JBKH6N;/L%NSVB _P\^^\KV(
P..\:8-KI6\D3[<Z,RTSQX\ 1/51)_M[EFP,=YO"IDV_A?<WZWFRD@\(&.F_/;N?[
P;(Y4@UCS;I 6_.HP$$V=_*#%0,2-T53@H$0D*N$&RN!<8.;\\O-FO,)Y+NV/???H
P^;*"(PSV:W5N8C&6PPM[?,6NJYC*$C0<4.B+:68D4RE5PCY$]L6(*#7"ZW6UFZ\=
PA$^'B:1UW)ZFC(0Z4R@&1M@.,E%QBOT_D'L#3V4($B^5 OQ6D'HNW EAEJ"/K"PT
P"Q(/Z :"%G&7GY-/#A,0A DF:M"AY&]-]BECO-ZSMFSR3O<<VU:Z.6YE\"EXT4D_
P<@8\V_E+UIVQE67T!/U"G-,Q1*0R&JJVR6S!^;T'W= DOB +9&:$GLRKHM@#%G>1
PIX%&H2Y;;*+7O9XT67^1GHNH6(3IJA7,P4B9]/=UA%>D!TH?J'&>DLBT,.5.)":&
P)$3.UT#.S I3QB2&. M_9T7YCN1%W4ABXS&_P@C_\[+-THQY1T:8Z4$\Q4H96%>/
PF;IUV6ZX1MPQ#$1I,X+>Y4K]4C0QHJ*DFJ7QW?E@B4(OER,T%R=!+F7D<,)Q1I-#
PSLX7=^8O=41-*B%O7-3*E_>&D8. YDNAB8# 6D:..9G6@!I,4<NTAM%P*=$,_FDN
POOD+S<>I>M^,FBSXNMS0EANV]08,R#,9X51)3?0*KJBB7+V>4JI)OBN<P]KN6_^Q
PL'P#M]Y3'3+.)V40^"0D1/">YR901:_3Y7T@VWY7TO?4+V++ZL /,6F_AZX&VG)I
P[[K*.;M6ZG@MRSQT_9DP/"&^ZK[R(@CS?7$03.2\C9;D46*A',E"68JXPH%2SL<'
P*8D'9X[?2+#'UJNLWOA1Q0]\T@[>0]>Y'_>]MC[)FIV+4B<-*&V"=N7I 4]%EW$Z
PK20=!3J\"2-M^,R!4\&BW/X>OU$AGD=21BSX1DQ*:#K#A#R@K>]@ZT3O7'3?>H#1
P1%6%*UQ9NS:^&(IM0T4F4V_E@5U0#R.Z*:'.CT+;8:0'_X6^/:0LFX(ZQ 0272MK
P(SH"0]V;PCHYA<G -6JEP"JE^]^#C^ZY0B<U!T3Y#!GSRV>RF1]N-U!PD1<[:K6K
P0U,BM>6'&4I#2G":R4<6@!%T8,$<'@2J_@=J-UW#+[R-+[DRR/R+\K!)?H9%3ZF1
P!R2JN#RUTRC T!C*,'FC_+,A/9YY%1YZ0^/*5XPT';OI?,N87X^2=Z=(YBEG3(#=
PCV+J4'OYI$G4"=UR2J;^G^6_LXX7RT$\\(B=:8:O(*U+)#$HZ/C&>E/9^*20&KV"
P$6.1Z=VOQVC*[%FX=@C7^88@:%-=F"&>U':$[V$9N *=J0+7FI=M^K69K6ZA'0@7
P,K5["<4/:>9-5W:$4:]D9FWZA4:;])3/.%'/*(R3J5-#V%DR6*/S]^!*5* 4*5;F
P2";8K*2X*A'FT>ZQXE!.1>+U^C21<FS9VEMW'=PP>9<P(@XY35?5M.B2+SJ8QGT_
P<2MLQH75& @!BGE:IS& OJ%KO'Z.J M=5:!+2$ZE7RX*-1@@.RZPW;/Y;!_(9]9#
P$C<K@]6=%P3F$4J;D\,08?QZR0WDHF%S%C)DZ\S[)O[+-,2GS[;*;'$MNB&BZKEW
PL"ZB>M@CZC,6(EK*]B;0PBM$=92!XD#]W1:BW?2?YT#)1RXC.(W[ZWJ*Q%PC>P6A
P;C+ON;WZ#FD<69" O5Y&!@R#A2"?UY?>3@4:NB])R?[,"-!&]_G[QQ=CV3_>*[F2
PWGU?3:XSOH$$*MQ,^)9*VU^B2R\]W+M 1 X5S/0KP?R4F_08;?^J+U]<L+FL #C5
P&>0VTGQ'1M[P^W^!$C$<'5YUU-(A62$"A917$"]4VZ6!BOF]P>.%JS:XXO@C&F,<
P)74(+DL.TOYD?^A?=CU>4S!UGH!RH1-'0V0$%)-+JK .[6A1;17D)5:31'[$^P]"
P1\1#4L@4K&%'OPW-V;X2"/4DI\\ZA.%LIY/N0ZP;U"XO@/C+(=%OK[%2%,T':8,#
P&>IR/M[Q">)V@=$"0%N]2Y^M8[3K@0MU&#P16WG6)94U8K/%6<H5;D&:[##C>+BZ
PNNIIX3YXH1145^#1&YN0^F"K=8C]\HT/0IN_9&*'O\?>G51'9-C0CN1'U%S\/=2G
P,165(Z8>$4O6\E&)G2\,T-7+6NT5W54UF%/$&*:%"E2AW%_=WQ..CL+*:BESLQ(.
PP1S>4O]*TO>7R;J[O%?/X5_7D@J[V:?3NQ5R,V:#S&N+JP7L^OQ :JX[H3R'KCZX
P)KH,ZT4JF&K3!:9@?04X&XG<0X-L)^F>@*L@HOA!U^S3 JE)&AU*;4_QP 6$2#&&
P6@5=/EM)*.^K+4U:=NSY$\OQJ36:,('3KU5ZG-WQ1H\QA)9.[Q7U:TX8NE&&U#GH
PA#@OW1A6):'()W=D+$$=2?]73;UAHGQEM_R2" 1AU6.H[1>5FE1OBFJ@.@LFY@)#
PV^E&)>.SHSHI3)[^13[0+/8=Y_L0KID@JD^UGX U+#T"D.L?KV8[* 2[99ZPG\.I
PC:KXJ;H<[@ZL7"0#9N?F,GK([C;/-S;N]F/_SEH$BK[0)IQ1WA23I0?<69;",0,"
PJN=W%"0F9H\POZSZPQ&MUK(,9FTW+@7[$:S!&=;N=&*E:W0=OH1*N&#IC%A3I'PH
PZE0;(Y&C;5@\!WOI^"'4G7EV?AOT'8H,UZ<:C4V^'RSH_/YX3MW-)]9JJ$#W,R)X
PJ2\AC(1E0QB)[%VD935U")0UTJ]J#0(V$3JA#1X&H]P>K.?SI7I8WYC^3"!T5S=?
P_#RJ,/O9NX'.VVR"I>G\1K@ZCBXN$)ZU)DGJ7^W*0X#*%X8-F)10M_$:+ECB9U;\
P\:K*.XTT_]*('?!\?T+C#J6(RY K!RPJHZF>?V19D]%W\!;<(-X/(>9V&OIP+AHX
PR04-;AZT#=OWA;-D&ZAZH+34@+!$+=)UH\8S7=)+CH1#0J+<O6>78?23H[EM/8)6
PMS"**U+*RLE/S,7-]'-(T*";!#XL"I/5,)Q_YLWX]E/7^&64F&*,&QWJ&RRMK&K(
P!?^:;,GJ7%B=4<-!'J%6B%$]G5T9;/]$;I"BU8FO4'A#E)83(WL8*>4_ Y]IH.A\
PTHO4:MB0)L86:Z<QPS+VBOY_+HD5^RXQL52TWP['@XC0QR68%$P\;CB=W_"H$O 5
PQN/BG:M_83*-UN9:SX!],5-ZAMD-*H<'03SVS>;4\]#])W'O1\P20*I^:Z1K-[$1
P^,'=)]3%>4J[2:-)D@*Z/IW#E,-B-LH,ZMY^#+3(P&6EQ;%=UAJEV.5L-<8_65+X
PDB!(A]*E!\PH+&FU2%*F?+UF1!@J;2E#/Y%H/J&.BMA4.=I1@Q$ /;YMN[YQ\>4(
PB_37,E(&M]JQT-2#@! %I,_/AH48-NT[L?(.\3RAX:$91*0T"KTP-?A BE+F<G6X
P0IF4?O@'ZN\:',:+X\Q\L<<*/ 68#:_JX+V!?Y>1(8# 7LOU&WX2L'0M*IJI7]..
PO_OKSV7#:R64@L6B<D &:QA!&7N!QRI/G(T$9,["VO*J7/NZ81&]]/&'*NX.Z[HT
P<1I+=>"-E+<> N>1_FXXI4KOBVD6; I5U-]/?TS?0P5E[*\(\'N6^N2FPU1,#B>%
P_XW17=)VNY<^XQ-+[T9FH!PJ5+0YQB; L3YZH4=[[ M^69\]C;@\NXRS8ZN[W$Q>
P;F+%G [![M[;#8)^,PV#RW+NI7SJN"Z"B7)UG:R*(+H(9Y"I .@96%DY:%*5Q2&R
P=DZ89R>K_BN)J+_J?<-#GI)A@Z-C>3C LR3HJ#R#,$7>M4P!9T:V[]:9GC:!FM<W
P/2H?RZ34[8*4%]M((8_? T\*PP25&O72*&U.6]L:2P8,G4WO:CO(3/8(LL;!_\_N
P#CH2W0Y49KLK4\PF;0.),?>!B3/0(@[D_8,X#I'KUAR&PG"?_=U;-SZ%^4MN8ABV
PY/WMHXWJ$OCB0Z8.!/7PZON:A[K:;Y,0:Z )V'[8A4>^H>LS61&9!=L49]F83F.M
PU*Z ;PX6Q*7.?I])QR52-Z''\] X#2VO-,+0CLSZE>%*/U1?R.-Z.,*G/,"Y;'\*
P^-YPPM)PKZ-S3+5*&B8J4IE@HHH^ %4LHH1V$81<=C\?GEFE(N.!^\AW^=)5C@2-
P.&P^1N5ZTBIR"0O+2XW%T)\V]675@3[\[C;+K$[P\.M=S4RP*3(55A4!<9<&J_P1
P(W%T_MO'J!J8U@D?*<AXX]CX6<H'7C?+0?:)R&V&WM.8>ZO<S,2U?/,@QV0B&A?!
P9HJFU7JQOY.&%'VJYN6SZ8=[Z4'G&9BXRCBBW4@MS/@FR3)\D:^"! _+_SJ10T 4
P(J'  &?UEI/,) MXEZNNQ.&!E)7 )11Z!Z/M"3%*+QD#<KPXT%08B6PQ)M N@V*6
PI@$"HC(S9V(F3PNDSBHN'"A:2AT-";Q>XX@Q+N!U1(^\G])D;IRG9 NU@H$WWR] 
P R+4#!X#.^;G/R\_!E".W_(6:A$6^P2J0JCL"JO.JBO@ZE3KQ1DY%)=6_6X:SEX'
P"RHD;WD^2GP/83<1E6QI+"UG91?!OXD''5(B6@DYAOE".)U^W\&1 T$LX&9OJT\1
P"9>D,OSO!ME?UNY@?5;3-)>\B4N6N&B+HB(:.V:'T.=N>Q!ZR[BC,V^.U-LG,KHD
P%G;<0<NP_C.LB[["8P(S/%46VH>!,F0S5A[*(UJL]M;>;\E-V,3[WFK\E>X:)\9V
P>7=9Q'70L(U26FD!^APJ>\H"=47THM?B1CY,IJ*ASAH=T5WN#HH0BFXF#W#R]=ZO
PR(.#5\)A%4EBC>RB,CCH5L:M_ROC[Y\"ERQ9 433WW\%JCURR713DDCKZ+R56+03
PRTS*Z*#Y$,0 4L(2JF5;5H,,&NZ ]1"P&:4Y\Q)KW#"Y/IDQVU Z@G"C,5X  4J,
P80U_$&^XTFRP8%1-4D7B\\\ZM5NZX(R6?;;H%&30(OHN,_:M(43.HX0.=O41VE"P
P:B3TZD0H-_K-M#U23 <#!_ 8RKC731L(3M;,\.3])Q?/3U8A@\Z@YKF FL'PBUU5
PD7C"S"-ZXQ"]D"A'%-U =ODO7$$G^Y&W23!6S&F/^D'&]+_DL]WKO(K!M:[@J1/O
P<<2NINLIW8;?D*C4B)82S[JPVR@BTV\!E)WQ3Y6-@XQ"ILDCE_J8$0@XV[!,WOW'
P*_>#?N">&*^<DP@6/,  C&8014GG \33A1 SNDSEQK46*B?QUJ:YUEA1%_)*EX^2
PYKL>^.'&MX"T+*C_^(6&[$$/\]:TP=!_$@V#O:&=DDG#G<OG4%+?]=MD70J#+W#V
P4H1KW"* WP4Z\"I:,G<;AR:B-Y\25H5CY7AZJUP8GT*.9&(%T9";>Q6.G6O-+R+@
PR_JK?=3=NPE?[^+%3EOC=KYCY!90V4K5I>=?<W7N.(RZW5#M[X<^TNOHVVS*<+:Q
P?3EAS;CHOB6[F*MXU+33=VR@:3-=;6MM>C( %# \\<H++Q8I"V\N"QR]UIK+X&+2
PKW2CN<O4HX1!,*[;OL4N6M+N !;5).-V4EA+RJQG",R%N7(&0 0<^H[*; ET?4V7
PPS*L[TA)035+C1;*N>_6Y)(Y!&F=#WQTFEG"9MJ.N'6-Q;E.7G=))5;5S0J]L]2Y
P"_K5LHD ^H<OR<*G"A6G^9EIB&)@XJ05 7O-?62!%1J]:6<D=A.C8ZB/K404U_YE
PQK"+MW;(>,E-;BW7T"Q\!G6,QDE1K70GU6;QMP87NVQ?5ZK4.=/MFZK<8//%,O1(
P GI\>#!R1KW0-,3R%J)Z]LF9K2J,HF=[F05YA. %(?*!*(;9:<ZG^JLB<5=4+T(=
P"*0XJ4K&^+1NKZNGCTA6HG ';,S04"$;8'&D# $P5FT$< I6S",+X _K)P!(W"O-
P#%NXIG'4XP\L!CC,C*RMW19'==KFJ:7Q )T%7RJ?^I?S7KPTY)$=:A<FZK)FFR['
PV:7]N ;/<L8Y9]S'D>;-#JP0A!:#H..NBY8Z@ZXJ9-3]+'AR6?WO4CZJY!6Z"OZ$
P=6_Q8=<*Z !MG^OE! \DD6'ZA_D87E2@&?MO)T"WK?,RI]?Y<Q$U/&5R;+@^JW+5
PP*JJ.\J)#Y:I,#&I^B*K8!'QB28H374SKR[9U[Q'.+UCW(JUN?J=+IJ=P<DI3NM-
PU.#%A30>RMVKY]5S&7&RR3V"J5$HD'6PN3U'2<7:]%0F,O(QCU]',R8SHEU7=$-V
PH%I8\?R])64*W?BAQ+F<IBQ8G+A7A3<2$]_^=PETZ'P&^'(P)0I!FM1T=)3>N]_#
P%I/[4PL--=+,K:'^RV@IENFZ=O/TF<C<4QD?F2%7%;*9U.&$U39)*$OF&7TY5_[3
P'TSY(T5Z,'YWY;0 NV1/_6@B'=R7P4FI$N)T[QR9INW^.R,KC#N[G#YHPZ)J1H%O
PT!%G$&?FTS*^OVRSJ$&FI12X!BRJ/&[ZTS_667J>ZMA;SHUP-.D&,<#JA%+8+;.Z
PY1LFP>J%Q(F4LU_[@BV)^Z\E^W*JI)9RIG;:N!VGM8+?S%3(WVZY08W5BV<=Q8#O
PE$2@J^O/WB.;&UA.,%#1;=D"*J8NS+]9O<;N#S'*QP1TW.TJ.G*MH\V* +?:M\8X
PM(5R!1V.,(@1,.4$,32&_;<NF%IP0*$^UJZRI>WG_'/"[M75E8[LA>Z?V)!D%8(D
P'X23?(2F"^:WWA==[(Z=T[K5,)$NGEIU?A0+)"\7N+UR.2OA.\B?OA* X=WR[6*D
P;-M@:TM![',G>2[\2)Z8=KQ$U@?]0'L,R/)LMX@6KJ(WR*T+6Z/-S.M2&X?VV]MO
P@B>!O"32:I3:1>BF/SU5+O+))\2=QVOM4A,Q6RG5U($A:8R6#A\[&^(*6!AY9'Z<
PM"5/#_")>N0AG$!(H9#;2!+^_#'L:7M( IVM_Y9$R@_R^G8QS9_C:P+2-82RT?/(
P$0&?%V3-<]V>1?6*MJ=TTC)<Q7%80Q]^,G@&(:;8YK .2_&*YJ8$\HT#'1;T8.+E
P\P=I AA1 &Z@97."HC1[3XABR87IHUO'C!S$XERX5&K0.-W%0>XF<K(.I)E>0$KA
PG6:@9&4QJ=P9O0/F=:L('DHHRB:6SO]!#[B56&'\"9RHXN_0] 7E]1T*-=(?//3W
P#G0V3*X)G7K_%V=]P3D!+Z:W %@?V5>$EPXFO7HW!\ZE0%X^E,#@T[\IX'Y4]&3X
P"'D"(G0Z6?4OX0J1/@B<!88[M._NV^*QR>$&UDZA@=R;ACYS!96>K&D,;'HX1O2U
P^..55AXY2\,2"9^=E6I%S"C)TVG_7;LKBBO"\$Q!F\?(KJG6\"Z[28X\C>QR'V4/
PY*J;O$IKP,H5M-?CC^ >C(B4.1X_@_=%=Y6OS F-!]71TYE&#H?U:X^,? 8\-E"?
P77\C:YVW29J/:3[9402A%(M:82_E-#DMS]<WFV]'9&'OKYJ7MG2]EAM"(/-!9%F(
P9C*6H'9X-?;KAO-_H5?X,(RVA"QQ;X3AF4(&)N>F::J\:FOIP60+HX+C2"STAA19
P U]4;]&%SRYOI=E^^Q31(?+E#09L8;2K#XQM1ISI-;WTIO>Z+.C>0% 9\8+;R<0'
P475//_3/?ND9EX=J=IY?.R56HF9W853"A;B_\K;J5K(%10CB.Z#J:?\0/B&SF]+0
P97,GGIJES._?!H^BCO_%Y8,X&F7P]0IW>%@@O8>1$Y\!;5AD] 8;X<3CP)4Y$24=
P RH (&Q\<W&#.%0C:*GY=EF$P39W613*17JEPRJ)2Z+1/=C-::)%,1R3:%?.S#\V
P X% B"G>7^\6+;$N@F9@3[ 47V=NS3?U]E0:WH9T;LW<SRNX\D/T/SHM6"'9<K6T
P?]K"ZQZ"3P<B+;$JXN4W*WXI)=8ML9".]W_06-<DHL5UO$GR%W[%3E:' [VV4%H]
P$OL&DI!,??%/[X6 G\F[T]!4&O).")\A5))#"Y].=RU+^-]>)S'<U_B<3WO_X-H1
P/%^QUTA!1"M;W]SR09RN<5)4 ^:T!W<-R/7"=7#W/F96V7=_"ZH%BD/FE)YZ<PT9
PZPSG4M$TAO+&[ 5%4ADZYHH(L!&_Q-OX0J_Q=DUW+_BJCC[)/(W/H1@&U' @$=W@
P]F.2?<*ET[RN?_@Y]2/*"X\KHDOA"^<RE1<CJ/ZEP'UVE5;Y/8F=7BOX#!H!<7F\
PX>#%X@OI;*L764/5DC1U5KF[$0=T8"8'"0X?W7;\%"&?,CI0FD!)%_N:BXF6,CE)
PUZ=I8[.D9TN68J_572!QP5_-29$387JE!2B!W!D2/Y:8\:7A15%"A!ZA=$H08EUI
PCB0*?7Y\7S^3$<!)QQF$YI,EI[3<\R'BJ)OY*W_A_J"4Z_:C%)B%U.MD#WW6@5CC
P7K_/'B%GUF&1&\:B FL#761V+N&V! Q^HNK,*3TPL"O-&&&7:-L+(E*=^P<$AO<Y
P/T#RMGC6HWSI*N>97?\=JTM;CCG!2D8O+_[Z3$P,XD!7B3\*GAKYE49QU-M);**B
PS6OA"$S#S'YOLZ#JWUNU9.A(QEQ@Y5<T!<A"1'DH1S2"N7O[(\)/FVY9\$+?9SF8
PU399]6([RVH@3Z(M!?%TPC?-8N%\&,MVL?WA#'Z04B46,=X6<!Y,4^JUTG#N%?UF
P17J4]!OK!A:P-7R[!]6.]PR.?-FLTMDZCDS"JJJ7#;ENFCG&%]9UL;_D-2,@8)7$
P?\@;V%G2OP%E 4_%/JO\8EAMH*:_!H4'R>)56="!?6A_O@5]J5F5;UE8%UH<E7VD
PN.>C!@0$3/WI# 7:#,4^3]6?WA=J0<S10<,F<YBHZ8M>+>-.<S1%B2P_!0K@6##*
P'@!OWSM!E)1A?HR00"'.+HI2+]Z+Z'@FW"GQ*RA4DU3]/)\) #<>G"*E*OQQS.HE
P]Y%/(RA_-F&2E!]V_4/0U"^"[\","()GU)*E\'1K='PY<.AP1EH07]R&EI-1UA'G
P@:-,3APUM:B3SF77_Y2^69MZE[R4#?"GBR/26AY%RA287?8#,])&?GSH5<<Q]WSL
PE5^)%<QOL)EFL]!F">1$NG<,(8WYL;H(-+&$[FUD=]E,_DRV*#J-FAP]-T096X\$
P*4OV1Z7#%&+IRWBM!0I:E!!:H^;"9:S1$#[05,AMX7/=M+N?\(A0Z'M] !Y$P$/X
PW$U;Q=[^26\$_7A\=N234N3VB'9(<!X>[F/8WQ[T@+^5V;_P, 2D/5T%$I2^2TN=
PLBC6U18X9MW3K9T+@=DRTV7CO:4M"XL%$D46,)#,B6W:=+XGZW,/V(Z(3Y77)7VB
P)B"D2N$BK7LFN()'J./S:C<WS0+M.7$N!@9M/B#Q63(TR7U"G:SL6$0[E.QD0-^7
PD!NGI&^H?0>^ZGJ><F$B[^%>)=JU1[7S877 <<*5^>LGSOTD\B::\U<[L39?M$NP
PE[?:>52=)5R3\OH E9[71TMK>@BKP+3F2-.=*U!<TP!T>CK/'U<]J\7^U#^O]%"_
P,Y8DO@L8 A<_"&RK2OG.I9/7BB42]G+YZXK^B<#WG/;;PKM)+__:4NS[L,I'0:&0
P8'V#C6)EHIHN4-8]TRM;^BI4NB$[7S1Y"?[E^NAD\E2:QQE9&H.H1ZYEG&0% E@[
P]X-FO<*IGY,W<[5J$;+K"GP_K&UV=G7UM1]9?TZ>QNP-=^X0T3%S-6J @& X2)"[
P-T<G16W->KI;W4AGXBPA-SF@X^FG4,!QG.N2'-?2+S$M*<?@'0: QAAA(WKQ!$8#
P.;ES(57JY6)JB:I=_;K$Y4I%XZW"I#UI_"(C(C"$%\6]P>BLE^J$%KY;@OVW,]YH
PWX7Y'Y/TL0*+>,IWV0X53,*9V,=%WI7+S6NW26LRQ!&=[&MIRAF1<.TIQ7K?I+F<
P,X9O!H/*AN=%R%2WW4Z*D\='[:.IY'<1_3Z."CS'#$&;+EH7@#_W"'^ %]MW7$KS
PY\A*_S+!TQ88G*:;015QJ/SUJ=BW2\G3#4'/;B@YPY2LZS01)QDC.O0WU/L&W[:B
PK.\NL%18;O[;E!+=0Q9Q+9MZQH/#O%TPA-T&211W*QISCD4ZRS(G0O2E!\T<S)$0
P%^*T(W@S"$XMXLA5E3= $U,1+:*IEB&)UMRW'F"'OHWHN\W2"LN\;ZJ,[$N)0EB 
P1XE**!QTQ4$ 86PN"!W8G*T?=OB,Z(D,#99&:F4=S^+@G,6K3--8DAG#N V^^Q*@
P@=,^,D;?A^E/QGV!['V/!WL:[]L/=T5""*AS+]>1EF1;NUUK52/-=N<N?+R[O^&Z
P$2)QJM.\N7BKY];7>7+OOVX!7M#'ZT3](1JN%[N3G>P=(U4Q?8V[2U1_+J9H!+5 
P=])&L#0Z9.L3/!M7= 7)O:AJR0JY:96[F'?T9N(LW*O'@ 8AC3M"F 4;C\6?$US1
P_7TW&$;]VG0J$Z]^+25T<O+.MC]+B)3P;&B-Z/)\I47"4$&]WX.WL)51]C?TSUCY
P+;/KD,-N/03("XM-IU-H"5QX'.%!XON%^4Y5HY2$DD&X3/85O )LF7630^_,42"9
P2 FKSQ_)F'4M^!7+?3>!0E:N5#*#7G,HD%@JW951[/ECT('N-PDKFQRE4(<XE0V6
P'ZZ:1-@8"AM[>>ZF;]'Y$_G#!)(D?9P#%!D$Y110"U\YK(<J+.&^E4Q"]0:VFPV%
P<H&/LJ^.R==H4)02;F6LZ:<"%"/!7%F;?_C2G>^S8UK.[_8TCB1\=7P7D3)9GEU4
P_#)90W.N9^YGH/N9@Z]P=KV"S$*#)J75BBT 23I;7!F-I&\OK!PQ3;M"G!Y 8+DY
P#O\87,M]>G*[48"FYJP*%W:6@$^OS#78,R)?+=A^HX)KKEBKMU/<&7L#U4R.F%W;
P"3B EWB@4'5=,1C8%4IQ@K@L<]X 2(M</5O;70:9"Q,5K0_J6'\/6K\A1<&8"(3T
PP'0"]8:%JEA^#"HP JD]:JHKQQ9CN'TY&U1:<A+D,=*366"HXN\OO\EKS&>)8KUM
P1@LKL1\..E6Q/&%CEX04W_QJG-Y3RJ6Z9]J96\A;(-7Q5)(J4])2K CNSWAL 9HA
P]=^EV#H@<[,F&3$I?I%*@.EW+0N&ZR!-:)O^9@YVWFE&%]B.WNY0<R=D!9)OANWD
P0=&B??%']3[A*/A(O,=4U+1Q[K^LXW:=QLGX"0(JC'A:!U;S7S@Y]:_4N$ "Q2/R
P=)5&54/] N%8-<B/V9S^U\G2?]$I_I*&;&A,A_:,HS:YRAT5P#ND?A"?+G2?3SSI
P^!Z" +E!W<+@>>XD3*G(T<&O=@XU6E+C=K# UR6Q+U)DQ6Z=P0@U %>U=QA)U^:@
P?3&=</X6%5&8K#*^E['&^U8O!1HM0ZHZ2>B((E%@B+/E!$V_<?=*RJAH7R5U9U1H
PVV4#HT]F?Y(5&Y$D7'79-")QN^_Q+O$&>+S#%0\(LF/EU#7/CUS+"'B#4*"4<(W5
P[_BV5%A:6SN:]-M^LK7O/2LVJHM/:FXANCTR\Q@)1BW9:J]Q&#DEWDX@NAG/[]#&
P?NB4[.!_@W>;:_V@5I-G?M;L43!0?DSQP.-%>6Q")/:H\PL@$7J_8_%[&1( A(]G
P_:C=*X'F#:>33P+(J*+@Z?GTFQ-2)Q+G2FA]K>0C!=A/>5!;A"PR-$S5)Y5M?L3W
P4%(P"+E*&3$RT([Y^LN[G*OTC31I=TJ+>PXOM!*K[[R\/>22B#.*,%':5-D-Y7(Q
P$((BKI]!_2[=QEU[SFL*_?[+T/S5N#K;<4LQQIU2Z@J([^^3Z6ZIP%R+8CR#[I E
PA6=T(!$(!%=VQ5R]+5H;O3C.N)-%/O\6%BKTT2B'\F?#^JX"=RV:;$&[3BH>BLSB
PQ+AGB T5\[/M9:'*$.V,@;H<D<S^T70$ISGRLJM.$LSIU-<[0W42P!]^/@FT?(/@
PK?)"LHTI>O-4@/8>>8QVU[]LP&J1Y7)1+8@XTGX'=O\B=J\+$V$TFA>ON00$Y>+'
P<W]M>[WN*1"K0X>*%%2!NAVU6XU3Y?Q^*5)NX:ARE&7?S_VXL]H%;C:*WJM06#5B
PX3O]76_=^<VTG*1N V-#\,J1XYMQM)P!-5'#NB?GG!BM(B=@CE=RO\\FS0-8A#JN
PR !T5NHO*3GWN$ [&#P0P)\@)E&2N<?"@/"$D]R8:[(Q4QFDV:E =SJ!A%4=C/6&
P(&."3+W42KY@T&=0O Z9L6@$S!7]^E2]VY 7_:(G8:L 796=N@2KMQF19[]%Q+6R
P8MY'R+_-V4J6,+$M);%^X.XGM9$6ZH,-^KXX Z,6(XKO=99Z&>H84#D:6N5PDF04
PK3VZM91;.FAY+FY_XL,B%CAJ:O8M1P_[62/.N86=M;_DZ'R@4L-@L1+SWD@UART7
P/1PQ]L%X 7TES5 _V#VS<Q]F+Q>S:A;+8K^G:69)+*_;$C)>PEVQO0K(FHG73^/A
PNWVL_@EP9PHTK(OXYOL^ ?H>,?.#:RNFG)B^)/\-Y5.4@U>O!5 -HA8TCR:KO,$N
P/K8.L8;Z.,M<[Y:Y@;Q9=!ON\CM4P1]7D=&DM_T^!WM@6/<?;%L3;Z]S4U@V%:4,
P2E,%_559>-T*C_\96T!RD0DDJ(PZ';X?;&E,\5Q*\7)$<&]3>M6CN4L^ H6%E%]8
PWMQH0,CA[2A"! >FYL%P1L^"+UH*C82;!?-JX&"V4-9<K.5(0U;JXO)+=O5F</:9
PS+\%1()>^&XUQI1A(GL&DZO!T)!S"/< F_'5NR8.,TNY/7LES=3[<ZT1.,4VA[R8
P9M3[;M@%^T^-7U58!W1$S7FOA[4U1H0CRR$+XP6%:'_RB)UPOI1SC7E..A_BGM+;
PFSK2?*;BB7U:@FB2B!<G60<((P&=^JIG@ > MT2-KJ#>?@Q.F%55?1V8VZ-<1'\#
PF#:HG0>9\F!R<I0J <.S"R'B DDB78IT&VTWIZTHD"0"12=+W;5?1#/9ANZT>+&&
P4$H\9VJ9X$C;/-K+(U Y_<-0,UFYM-72:*KF\X+_"QF:3%,^?9)!;[@""Q,ZET <
P1PKYT=0,X-DDHDDM:YV-]N5C)=R]F_%CC(Q))ND2S!EUH!(<.O?Q7!=+F-5&)%I]
PF3=I3*IFNGQG3OLC^\;8S<3Y>^-R\Q,O9P3:T1;!+HTRTG,!MJP1_RU9053< WSM
PH+;'4!+0B=& [YD'12-+OAO]5(J=-&EUN&F-F9T/=@5-6T>>EB%"^66@0S474(H=
P4X(;,;N=PC\9:L/SK!U0<A\S1!V6ZHAF??VG 0JIX,='IGNX.'?)9CO:77$W>+%2
P@@&4]*'U J0O<@TC+U*+#C&N_0F%@: &Q2CQ&95.NT.*OFST/CP9S-;YN],PLP<$
PA[!]?$"&=[\HJ2ZJT&__8GB%TPML-K&WO)4_N4(BZ5+4I=E%TR3D:9/]N<H6!'48
P0:;=SUF/!OV8L)LNB;]5T_#[H6!F:(O]S5=-Q?;6+(Y=;;@*[38/"3[3?6'4&4'+
P%PSG=95I=5_D(J]?K&JA/<YY!%H;.9)6!FBZ@3PMVX@*.%P22."^V1ZC/!:U)#K"
P%)'9W63IR@2TBE5;//3%;H2+[)1]0/_*M79M;'0F6:7_*:&FW<+'[O<;BM%P=37<
PZQ[[(2C*FIZ5JN"P."Y!26$90!^U]MQ;<A37T:YQ1J;3+3L8X/O\-8#%$]P9HX)V
PTU"B@^ZH^K[>PEJR_\*4G_")$(ETUQ"+!9#UH;Q'RJJ (5C3AR+1?,9B[#17!DV?
P>JX1'H.U-/V+FMA[(FW^/-3[%=,-)V?JM>M'^KRISBS)8F_+-!ZZ%%6B^"FZ7"EE
P"]M-0JBNN8][;HOH2US E53I]14+-P/<S7U)1AG9$$)X!T]M6;JO8YH^T(P][:^(
P70D=@?Y[./FUID*$L%YP%2?P[B+[\<S+I]OZJC6X93:A('E<+J2\XF:3KO*(&\[:
P.[_&9E:Y%5NTXLR- 'IW0E!+ ]!9R7C^&XG;D^-N )%=?"\A@0H:>PLN(<_=CX"B
PR14X0.&F5M+&J0(KZ 7#)8C7U;R@!B)Y*=<;5:%U2:OC9HB3'3P!7AOKG 3$7Y=J
PJF3[!_R&)M(FV$@]_CI:PIWW_KP?0K+:+HZ$8/$0TD(862V_KDR <PVWMDC@I)IR
PN>[%KJ:^$MK>O#P4H2:=?3E9=N(5MRAC$B9!DB6<OIJ0_[&),0Q/31O.OO866VMT
P4NQ466*YIC]"#0%5=+%8 2G\G""A+B&KPG99>7VY*FV:+35>#?#%+)!52S;H3'KG
P!I]SU(-E-S&;/5#M-)6X1S_&G4"UW^GI7EX"=0BVG4P-%<(<$(D6&A9@Z"G26P/F
PVOFX\3>6\:Y HBL#MOOIU$I9MZ,^R.BVM HMC=O17;-%G-Z OH56MPH7IPM;S7,=
P1L!('S?,>(J$-&7!)YB*#@]B"B%H%%2U#C&B  Q>";G]_>LDTZ%6V\I9%?_2<72Q
P?AUQ*CB1Q<Y")3A3@0F/%/=O+K#L#Z@+G):8T;#/0Q[PPI\\QS3)8)90?8V;2V]#
P1%^^#L=X-IJ<IQEJ8K!4+5A)V.4!9@:9O,VYT7+*%GXR2V_M#XQ":Y]#S1GY#BPF
PL6N)\JAI[28"/_IAD%9QF?FA"8C]V6M@"K0Y2%_+F 2FS9?@T-9\,!/)%P&F14,(
P%YNHP>VIS7MI=V6)Z'0ET@/,  H4^QTB2:_FIJ[PV1OMSD@3:49-Y&2XQ(N_@WXW
PRO.F[RA.NRG&#"(=@:IS!4*(<^><K\[U52!V=H^P2S.=2RZ,DQSALO)I#^BK$N./
P7RIVRJ(VR&;(=/EV@I4=.,RMWV]260_P\&-&?KH:GZ:UT%'9M%8:]:TN-B<>J"T2
P5U4>:](C_5JM!MP0B4_,M5PS7!/3O]U?4G2/W"[WU_/HY\MEG9@'7959]Y1$74DN
PG%>^T:=JAZ)">WT*8RIUK+((2:"AND^0H\XE>9W"YR;'4Y:>+\[,D/-BPS,P?@.&
P_32 S#I\ PT7XE*IG4>C&*68'TPIU5M$D[(Y"\1929=#<<LR:>KBF)$8A>!P4K'+
P#6+'RRV?WF8Z/1^K9-NG@W7C97,B\B!N,L2H!<Q;*^SZUP:?!/:;!R(R^5U1HC$I
PZ7VHU*BU#S"-Y_#A_(RWHZL%1*TM^"LVV \'&FQ,B_7SBYY#MO#"E3F:3T!@GTJM
PWBLH[JT1L2+YN4^<F -A 8%0JMUD'-DWV&(7G+?HQ_Q0A^1K:=/)W_],[YJ@H-D%
P7C0@!*N >D'_5.--OZ%-]"?%HDU"("^B'*T$>\W):T=N_%.&R1T,H9!6.1R@6',P
PZ<7WL]T">*%Q=ZK[WC3_POV3''@SEJ#0H,5_1'A+^V:1G/&Z"KA2O$ VN6CSR;/U
P/[LX'3JM=XZ-I*AH7^@>*WKND&9K_/R^9O15V#:/DI21@C[["%0X,[G@UD64*9KO
P,_4;[0@3NG/OC8\;7SE[I/LTH6<92%8@FOC +)B 1.29_=,J5' ?CO/A\ 50IZ+$
P:9<QW(&/:N+,,RR-)S6 0=:P:B>P,OLM$AV*1%A9 DL]9@:TM49S$/R(HT[J!GFQ
PEMK>\L=]L?X,JB_SCVZ[17SUNG*Z@8I9T6MM+$+R?F/IA;[BB<K-L*".S6YI5W*Y
PL^ZN^ZHOOR95$5P8$7OYMV_V]"#'DN>HL0F]XW4CB8=D4XK,C/'W]GEJ_#U".N:2
PKN/(YO%T:M'HA]P8RK[)I28Q:[,6_;[[-UC5&I#G['=P?G@Y7+49B;<GYWA9TU=Y
P .D7HU<\&3U76")];!VTY&XN2PNHY]C(3)7S &G@##=D%$&0:%"G)EF.OUP;W$4;
PQ!'Z=EAG\G\UE6?@.Y5AR&X[FB.)'XLF) Y$X8R?V.^H\P5U9))"!@H'IU6>@^)F
PN,02 N,[I3ES *JNSR@5JWET[D=ZV97_.;V;M'Q=1<[^! U^4$OC#Q&L!QTM"1[A
PR.MG1>YL$[P')/1R]_:[2O&+3\\+NE93N(FHH2_Q$EP]:&F8+S1Q8^;EK*J7^EBB
PQ=%>R'2!!1W\"C>KG5#>WVM4M$7$^H1S#M^P1HDEPM5F;7AWBJ7QF&.]^?QI11#-
P4'N]5J&_.G\.9PHR]M%"WB(0XZ!;VU8;VP0YAO7HAHA@>*TF]*B$Q%I"3@0,(HEU
P*CT!C(=%Z$WHIY[ UN3Z-0B1D5 [<0WQP!XVF#8+A:(+THEX((1V^@+K+.<&3ZM"
PS\%#J(Z&$<_CZ-%34&[GY0LDUP9Z/U]K4#M&@50_[F:RS";T.RY@QK(Q8)?L+UZ9
P!! X7P O-P%]$Y4I[#;Z<K)K&UH5\4_L?$!Z3)2$5XGC7O]XX\U-3>9G:P@M#VGU
P0\^QZ&'YE<>=^7F>1Z8O(AEB&MK$U8O/,,O*KN6H9P=:A (&Y3K?-,?>G6 5=^[K
P4!)HCKR=#><(+P?CZ59]HS7CKF5=M9W!70O NO7G-?&G.GU9?2Y@[*4_"5C-2AJ"
P,ZU=J AO5JZD)U*F[ S"PK#=DZS+AG*#_]<V#T;;!S>YH"\S_G?#8<?_E'3EX]+8
P#N_0O_:H.77,N8$-H9XOZ[,FE8+*EJ<>+U*H:(IP[K%/XA!S3&?^N0&W3PY'R@<;
P*4 R.R^SKAP$"9G?7RN!<I\VJOHV#6OIA+(6S^8EE/(>DO,:#JH(=M7(&AOQY.F>
PD C0T>ZC=:*L"8DG,&RFGNC_+P7-G9T*)+''SK+'$?_+-WDC;=1 4\8X:H&88B5.
PD4Y+LCOY9J<BI\\[:GLXIN5E\/IZQK"2^>(M+@!:BM\E6<%[FJ)30WL5*6HTLMO&
PBRS3"M D\0[WJ=K28:D([^W6H)9)K-*GIKNKD.@:A<?1N3:U EF'F*1/N[Q)(ZOS
PL70&FXNL/#1[^JH%N(4*E2R-# $30POZ=?X97'*?[N$'36EP5ZG#Z .M@+BQ&^%E
PWA,]8Q:BL:W ,$'$R+&D HJ%W[]_JF#9B%5Y*=])5GA/OR<NJ"I:G[SFNCR5L*B-
PS 88$4LO^ S3^R*\G?R!=UL$A1<$Y&\89-=N#C)B$3V^0C=*A5G1[G<R8,R!L;6R
PSSI"_'"X*1'#JPTN#CWE3K 1@Q:/IRW@/M*OGLVA1JVH#G2#0$-B9CG/V5*?@>?+
P6%%.JUVU/>_BFO##H?&'' VF4C_W_W@/:ZN!/1?KN&IY5.O]<#GWQ[PF%=XMK.K$
P_V>4V<F5@A,=B[\>1M]$",.,75WK^N\: ,VZ;M;11SF(<K"-:$:%/AE6?0G_HINL
P=P4MT9E:N3GMR/6XI40NC$0B7YTKJ%.P&YD'>+01KAMK(E!7T?AG^A<*G;5OPR%P
PR;?PAS2'#<&J@XHI5D+&N$)V'E<*0P 'M\FM<<C%DD$PQ)/I..N#%1W#M5^0HF8+
PX]T!C+6A66UTH>LH#S<GA;*C:+ %(D\ ST=BN%#IHJH$1?TPBSQT?L4ON<2)>@@.
PJ)*2T&UKIIY<3>^)=?/$JM_4[)Q)40C??Z<@XH94G."?AGU/OI<5SLB+]WJ*72_7
PZCA% ?" A9*H[6DH'I8K'[A/3 _B19K/*<PU#8A;KJ7LP4=Y<R,6-N-PBJ:A(308
P31A X!8Y0K.4;R<>U;G'/ WP4GV90S1B;:5P/0H<@S/^!86Q3 \O;[FLB(L\$X+K
P"FZ=_M@$=KHU^E/P,.O#=M!PRMW([-O<H77(XD-N-1%!=9\A'P3A0(D!(BEL_+\I
PW"]>15W7F07%-P5!3:_*-I 923V\H/)8DZ''7:S+0JN@MA1*2L)DFCV=N>70GI::
P,(LR*4M@V2A@\S1CBHCJ8[RRE\]Q:;22PHWAY2\6S5YS#S7V7!8OR]%1F0(EG"7(
PE>#*D?ZD'S&(&XC873S1:&#\S$^M+Q*DG]I\EB(//6":@_3A:IIC'<K01:7X0%C[
PEP,;U9JFQ(3B7+^RV:^\+K9(LYKJH?4O84]0^I'2:,>M;0:YAZP?F%2,B6@H%ND'
PCV^I.B^"#9F)9N(<2BZ#M==Z]FG6KKW*".VGT^?S9K0Q3^B;Q6.U!':QJB55\T-H
P(X64<([^$=#2J@AG_Z(T86\58\OLX_]^I,1B5JW5[%E,26W9,CMH(Z8G*#^3GBA5
PIC:U^L!D7N.F[3KOFJ+U=W- ,C7X5REV -C8A*E*!GTMC#43M590DB[_Q5CP0SMC
P7OI*/O0IN" 1N(B7XS7ZPYC\-.2Z+CISK +#"Q!7@=_.>F^<LX&=T].$#L5<[;=*
P @76B,GXL4#K R>34RY0",,P1-P/S2UI0LX03VL(I? ZT?F[7'V.Y,44&KYXJI[Z
PD"5$AX?]^NJL^,O#MF-J;.P_60*D'9];989QN)-O =2NKX+2#LRZ86[SN%EF'6SH
PAFG.=B4?SU-%.4/I.#)$/T!UAN^FKV#5/ME)8-&)T]R*_ )M6!;"I'H'? 6I_::<
PK)1[A*?!^XV$I.2O2?VYFF?8:]&23>PA_.+[]KP=2MJHZ*#O+_VRL.A,YT/_CT_=
P1$*>,#!W<W;9?6?3_SOQH>B<KX705W>^,'/]TOWD'" I8( (/Q@014AK24KISW@]
PX3^^I(.E :YJ@Z'IE"FR^U!&/<;M[)<^;PB),BG1I)P3+WQ=_Y4\K@._OL&C(62"
PX$:4\2.W18\3F$NF;?KH6Z@OCO6J4\B7!KG$7A3.O;SWG<J-0]AUW 7Q-[#QS";.
P18?&\Y50^-F)#@<6W*<8]K:Z>QHJ'2VA5W^BHEJ]O"$@^OI 8YPC<W1T>+E%CF*I
P-_<J3$?+C"0G@Z>D$X:H$@N 0S=O2O?T>XXMIV0(@/1=2G1,P)G.1\JY"S>SYF%V
P.#>I"%8!4Q(@E,Y-**HY*+$#7H)6#%5TO?:5A4GK($\N:GR6MC(SS0-;?I:T3+,W
PGNX<=VBJ0(Y!.%5H:2Q-_RTAKL0\P3::M8^GPII"G+O.>?PJVU5*=\L==>>$X>F2
P$9/YR4UT#LKW+Z'"49=1@1O-O^J3PU7$4*!KFR6D!N9_XD%O.F?BM65\]&H&5E^.
P?@B?U!,73ML>0P@8ZR@]_<EG*=B*U4%:MQK!Y'OJOMR#71#^("ZP7]E)J%5W\N33
PU6?KFO4&MJ0/F!MMY"STWS3I_L?K*4"AVF&M3#"]88EV@+%Y<I)#] 5;#U+43Z=J
PNX(]Q#-_$HB+E]\:Z?K>W/EGJK38'P^:+D KW(ZUK^TO@MLY)-@3 C/)J,]0:M0D
PK5^'^)M?@;2JP$0PST'QRM5(,P[1?3QO4.JH7WJ5#4VK/&F62<,P'K&P*%$?%(>2
P+W_*!9,R$ARZ,2'I(7II)#= ;2PGMQS8_ADI9A6=%LS */:EV5=AR1AXVWP1/E"$
P.S?]D>Z$Q!EOF 8]P-99#3;6)[U+VD<JRDL(F=QQQ)NA:%@+&QK[^BO6(JS^-?SS
PN$7E0O2[/TW]G<[.MHW+7E16/DJ2#2?+<0A%C<Q/***+M^'/,W3TWNK,+"*'+]<;
P>9APT41U^+DO(!_RIP/+J:TZA).2/!YF3>:B'%'-+!N3>5KP!?3AP>.1QZT7H#H)
PU7"+YG]"+^GLR7-:LV)4MA]*[Y84Q)1W">1@GHD]R@JY/36#GR=R>8.2=.[2SM^F
PR_CQ?>T/4&_/S$[A,HA$S\; V*__/GMDYVV(L*X$B1A7!/\?$V:SFJ3X-WSBQF4R
P90#$*JT I?IZ=GS_*/%6?2HX4_S^^([_\-%%3P%ILM!]7@*RZ#P?I<YQLR8G2[??
P-L%/G30WK ;Z,3J0<MM-R&7&['82.*3Y'<DI5]/+;(=S;,";085Y#]A?J9&KYX)(
PV-5WC#BE]M$0#K6'E& <MXY]*Z2C"8$=W+T^O2<:A(\>-R*]&[)XD9A08=\%'7O-
P?$BB/H)-]CA^3 M,C,??=[3D;AMU[^'L^HJ]2$]6X?64;*MNM!(<D5\FQP/8_H%"
P)\%L1@T\ZS54\)]'ITT5-6Y&A?L.3MN']Y &5.Q!^E>>7^5D\^"\,29M0I[J:0U%
PYHT13%9I '=44YB"B>"\-X[[!0?K85+EXX77&_KZ(-*%./8XFM;:QO9/8DX;VMKK
P-Z_$_!<MMM#?8G4,E3[=J7&V& @5 )A)2E]L]J%4?A?YHDR*BTL,,OP*^B-0>EH5
PB_'?>4\\[:3T=?_QUF:.XMQ#L<M>TL*($Q;1TFQXJ=->\F[V&,:E%'QN6[1Z22]G
P!!]^GL2I(L4#Q^A:+#P7V%G<$8%>6N\T!XY#2H[T<+GEZ=5.4G7>GCRHY!<C3U6=
PCZ3G_'X4;8YV\(R:^G&PRY79?8<JIE4'.,\A18:&RY<)G8.')F!='KJ('+$BHW2!
PS7YR<N,F"@=TC1M=_=54QMF1WR."/Q_G8$+L7K/EPRXC0-<Q!F&]:&N[2V[1E/%<
PZTG</O>_&F[ZUT)A%Q;,UIOVO#KSM5"TIOAK1>#.;EX .?T1 3J]&6>#19EO Z/7
P[>+-W*K((BL1"Q?IS0W]0;BX_!^&S<>]/F%%SA6+W9R:0OVP$#V$8E0=9]8/T]N#
P4*]IVHO:=30FTC:QSD5G%"*G:F8(/)O>4#VNG5=6XX/EWZEXE8+9+S++>'/OB 07
PK_P,72E4_7<3GU#Q5/WTX4OD*4C4>D01@^1"87T$ "5AU,]J( [G""G-R3!=D\C!
P0^0N-,GO63Z;37L6EM+K;L&-KP[H@+47W E#HG1VZYT1#^KR^9<M)QO"+%J45UD<
PGLYU_%M>.[)7"]4,/&W0;>SCJNWSU8,!$1(DMB;__Z64>:5Q6ES9=^)9_:\?>$<W
PY UT^;_MLQM7APM25TACYM]12AD4VZ*<-,\^!2GEM>2GLB_^9.ABKA\36?$I!&39
P=8#@1DDF]=-7N4#5\4*M,S=D"KJ*O[,#$"K.V,Z,%GL%/,M.:NF\H&_B66<5E*V*
PP*17R*8I4<SBC47L%\BBFX].W'3B&ZRO5-\E&YFBT07P^1\"H"\)$6?#?*B:TL=7
PE=_V-@P$/5(%M4^_VAHHJ+V:!6"E=:;ZPM(*)\=.E*9/#(7$GY\/RO=^L:8[9A\W
P "<;2P"17^5_E%85#^K-:PJ! U.XU&BGEJD&\'K:[<%GH)T!-GOQ-@,<K1U3JK(%
P<A-V1+RHSWJT,43<39QT@Y2<0QO*%,;:Q%O4%'I<L*],)%/^@,^<ET!%$9B5:AYC
P[C&/!.&WN7'6Q#W[@=(I;"+8-89W;%Q1V[3H1&4VA"TJ]\]$Y"[.,E6N8Q"UISNJ
P"0F_/G_K%'QM;GH=['BBO8G,O^9Z "[-H(>CR0.D"R,L^X@Q:8#U!G5JR]HAPK2W
P5:R$!Z%/;<19)S5B\M+<2AP)613IBJ#.FL<]E*N;6@KWD5Y\.)W[#['E"76_)-D_
PEI9('V@.V4W^&@M(A_):*R1UC0ML<Z) 1&=NW->DM2N!0Q=M2>M$E)*&2CF9N]]L
P!SJ\ECN8$QM'XH<F>]ZBBE7P+49;P9MB8:5&ZST7%91 E SGNXBQ,K$9<%PAAXIK
P_QJ(&6\V;XVZ-FV9O,L%:\8\P3RGMVB&1>3/!B-!UEXBMJKT2A*@@?(=*-SD1--1
P0RS8'Y<@V!H.UWZ9+MVKTUAM+O.DJ#*0GE>'<K/-&T $@'?"N.DVQ[$0^ IMH.B7
PJ<=RBZ>RY>_Z>Q'EE3AM*+LD-EIW"9NL<K>!(>[YXM[^>MC7!9LI**'?G/&'%6!U
P)<A9L8JW*U;K*F=I&XH4$:=L3-K!<B'AG!"^T(!EZ6,!34SQO IFF#=GL$=3#SI;
P$2QVO"1Q>2G'"NDHQO]7+Y+%%P@5U(',!63L%.[S\0+MB,&AD@[0HD'/_@@ZQ(I8
P+7\5EB$W'2 U(5<"(ZQ-&#,WI_M\U^0G\7IC;[3,@?_5[QIYHY:VUM+ 0C[4L>":
PL6][O@Z3[KM3)!>U*XN^6"1VCI W>LI=&QC'4'\/Z?KJ2W09P>_(\R_;ML0'NT+2
P0[EQCRM284WGD@6F_F4B-:_$'QTLK&_L=?@<^Y]3%16^P! QOLBZ ]"J'2;UKW)S
PL%P.@M:Z?UI),N3WS:!,R Z=.!*)2T/&;G'S@QT=/?FN1I+4^SZK&D+5P*-%+O+&
P$<LS"V*Z$D0Q$6&OQ$C&M-&@>V3V /V'0)'U&L!D;S*OH."=ON'&8\[C2)U6N1U"
P\F:=K-)+A+5HW1B3B?./UIB536F6)9FO=X6?[R/P46<'!YVW</N\K=&^CS=T8V1)
P5Z)%N^V&ZJ.3SQA ^26:M:6'8#)6^7!;,6"D0NPZ/T7,_HNBN.\T@9P!;"VB@-NO
PGEIB0$Q3E]NG(:E;OF8%C(PU/>-*&GZ43XU(",R@1D*A\(\J1>9'8%#ILE()< F'
PS4(O!S.HG)<,2'V933O4'R)I$2^+HW'V]DJ)/_LHS_C6P7^9@WH;^;7ZRMZ,7P/F
PQW3<!-PE;:9V6=A;S"Y,5C,!5JRM90V1?0LE2,6_'KHK'*%,0\3NRCEH?.=NQ>.]
PO.\]Z((/@B6GW@<%##.#SA6 NF+.^I.)9W&=[ T4?95PGC44%3/QJN1;X@_6'[PB
PE":/]G#C92[^]:FZYA7LZTZQ1B?B"_3]&9"K@_G/=_N>91,X?=XX++N-T":CQ-'^
P8\9?6.,1P^3*=5D2_1;KT)M DZCJKO9,<%,P"YK?3I^*1!UPL@M2>Q>'-F$IEMLA
PK2BNC.KUX^OJ$Z'7 S-3>EZ_-5?[]?N62:N<,-(%S23)2P6#*R)9.9-.!?9LY$&6
PT5D"X@:2L19<\?@%.9XTC*$L+&W$E3WS8K_6/*-W^WF1",*8"W-DBY.8K%A@P\B]
P;;'.7W!R?F<X:;+_^BEOKO9R@1BMO:,+ATJYAAK!4J30*)YO];*?DJ%4BI5T+[0=
PMOR;N3B42/B<169:X$K84B::WK9PX?J =^$OE0DHR?NI*6#DL$)S-K7,E8"P]R2X
PKW^6@*&-,(7Q@*!I1.0%[9'Y_L*WMCD5^03?I8[L$AE.($D"-W6X7.IG<PG-^SSB
PA<)N\"KCW3):8Z+B2<Z[J7HWPN( )J8J U=93:EJ"<S450Y3@8-7[ YMJ9^UG%B7
P^[0?2^'_H]#H,J14+*."021<PVN\;B[A6M35\4\3,O\Y/*/@*<U<;#T?H$SN^-4#
P4C11<E+&3AJ_LW"XN3THS6DNK27[9#I8RJX6T*D0\S9)D[M&EK&D*MX3&@=)L@CN
P/!.CR"+#(;K+VJ8RH%FCR/30YH8BV:D(/E24$,087>Q_RTK5,@?S[:#,P (5AV=)
PR.M8=,[/Q?(#SLHT_-$T!YKD!$B= :Y/@?9R-/40HMIW>TDK>;I@)LD6[U9Z/;C2
P[G>%%OWT:=L38H"N) PCDP,_LP/TU-=;^WQ74]P%/_+F<%*JCS_G5%>&^/)\*\5G
PEL:+#VLIJ'X;4'K\]@S@[1)?"T^P3)(*TOKD6#)>G;)B5!K!R<; 9A.(LO M7]D2
PG:\#J-".@B8,^,D0S 9S"B-)N9[D<IPJ+US8CD(4(_FIE]]\<O$09$4D+3JYG63B
P?-*W#OC81?E'5SP>(U=9WVV"M!3YYJ7?BA@,S8460XVLQY>+%!<A"CP_'_H*^C^1
P,4XPJ:=61#WC),B);"T?A^V\E]AYQ/C'<LSYYD[:>ZNTKY<>^2&*5:G.$@D0H!NM
PJ<5%O;UTJK09+<6W%4\R5VW?249+-<@!:7%@$NW]\:)U2>]K9P[((RLET+;*>/[M
P/959\\COH^1Q^)QX8O@HG]7G0=);,&HT)4F\>;Z$)B21V+G[?AX&Q-ANK/BZ#]2L
PE2 DRF=$N,=+E5HF;>B<MB(UH@SZO*= C7U"F[C[F$.\5_[1U"MX :])HM_4D[7:
PVIZV1725GS&3?<$NE?.8(_Y3[<TM>@38LF5_>$8BT1^=VVTO80**?WM6CC /0H1W
PPJ!VVCCH;!K^>VPAQP0CTOY6(_7#WG+5Q^69GM42!2[OU;P+'E1;Y5R C!GY_\\3
P+L"?4MO4BOS#>Q:&'I/L3.0L]B@-6.HH@7NXN)*_K4OJ[K)I1^33M+_I82J\AGY*
PW>[V)]H28Y:7][;L^,!N&GQ:KT_XTC]^S?J[/Y_$; *:&%9TQ=.QI5NZ+!4]"::9
P--5F_(-DR\&CG5[_<JU#.[Z5E8.:4>V9X6I?Y6DF*A,*9V4A,TXT5G#&1A2#K)2I
PU]#82P!A*V<"01=H&#ECYG.*?8B$N1,WZ0&(XV$5U2WZE#N"'"Y\R?=\[S&MH-B.
PW4@<+U)4ZVE[V?V4.!*@6_!"(?9/-+*EM.OP[0GQ]<28 J"4RZ",R2E4[;:_!C$G
PK=X4J*D^3]\CX2+&'_,PU.OWN,::Q%&X[SZ>$^Z,4 I:82]>Z6-DS?BWY@$B[(]Y
P=.%^$..N%('@21T1]X]J(=_MHQ+S:VSF :+UJ;>E>T_Y  ?RT2I@8Q+\>Z,X$3$^
PD,342:Z<3>4I5V28@L/>O3#X^1[8O9+[+NP-!D\J-Q4^!\?ETEWC'.Z]KBO(_3H 
PLUROV)Z]OOQKE9/Q8U.\@N/M3N,ZDOE"3!YS \F,9";B_I_6OS^.-XD#&E\@X>6W
P26V !@E_\(A3FV(22Y2$YM?!1*1:&*G%M"O$K; J)S;;<O?^JZ6TXB6D+TK1%?/I
P+A,G0.(RLXC@"9N*5TO#1H22&]Q::S7P&!!YSRJ7#EV\&=/7D!4QJZK0+')9^]F[
P$4C4M!Z@&NKA7[U?$&IN'?6RYK 9FMHM]/O91!2HFY)\2:MF/9B'>SL5J,PQMQ=#
PM5]8BCV22^B:@6G:4F140&I(Q"0-3]3\>H<3@FKL$Z$8O2/J+P'%'[=_F=GZ-DV'
PIU9F<4F:W%4@FZ%Y;GLX;Q%@K<.S4U!]:VU'* A/6G$QGCMJFYUOC2?#-F94^'RT
P?>^Y=>'O1M6V"&:NNY"&5?3->E-KGRLVPOGJ> :M.$9!ZM)1H[4=4\Z\)!&WHV#[
P\AM@OLE4Z"K\;'^[;ES')8PM.P'7W$^>66FGV\S]L@PG$8:<C#IR$N#R)=ON%SW<
P&V[[4A&+WQX'XOTX0&8$?'2^(:<><O)ZBV_9GLC0JD<[F4CW#YXG&CQ'$NE1C=ZI
PK&/D\B0L1[J7E-XS,]PW.0N92[C55?Q9I(7E([+7%BFD:S 2 /-)W2?+' ,KP_XS
POI]Y61=A!K5?;@Z=*0=)-O6@Y(V7 UV87QX>5Z#M+N5&3#-%H#9'8UI>V<+2SZVL
P64"D\R30S,'#3JO<0&+X_:X$Y9H$G:]J!S6*?!B-,8>Z[U_L@WV>+DA D#-3D=QR
P^,G_#%1=CV:O7,SR @-=L%4+IZ#Y;&?/T2IMD5HSFL0EWP=B;TWFQ^:I>JH=  /&
P=LV037;>F'<',&'T,XIJA5<\C&1;HH(KQ]6/4W^:EG;><K;6K?XY)8CXPW;BSC-#
PM/- O[">L#@0N'/K-VGI_ULX?G/U)R'C -2>_GI"DN3T/XM%FB]R$AB D\^*'$DO
P=K+J&X:;X$,*A2CNH0DQ03I;5J3=_D7ABL?#)TAYU+]]!6XPDDA%QWX)8QK324$0
PIGB4#DY#601?C+T:!9H%)3#XU#-E!9WD7]IOJ.<V#-DR_JNSHUL:QM=NZRN(%;^B
P6%(M#QE"%P:_'XP[?;;MN6"RD(JJ5G%+%C5EAA,M.AC>4R$6'/IIZJZ1KB0"5ITJ
P(WX S44'>FVM^-AHU+IF.B@M/"]F,,K$^U"TJH= D$^WGR>(&<C6OER3*K<,V!_J
P%DT0GR3K>$P>.9>@08I.7V")[>M^?N0?(Q6PL2/!R6%=91SU'U87V14>TA'OA0^>
PM7RI^PL#J6H@JO4'K5/IET/(><TM3RM?(^%36@Z.DU \7!!KF@(.!"L^IKQ-#XOS
P"WO]P?%Z<-IDEGM#6V3< ='1EZA(;^M<X%9;LS<GJC0:J?FE^80MHUXOX;9'\!WA
PD$N^3]F1DD8\0W*MKSL6>B6^63H-F=8,->V;>>Z/'EBXY\!/K#SAJO8UHWW)_FKD
PK(_*[*ZU<CU[%&(LV:+?OF"D@1<0Z2<X6";[O'$&?Z9AD@KCLU'&*\LT/3 J;%6\
P,CD>N8'T<NPO$S*%L/;'V2Z9PI;,X*HV!B!S#'$#Q @\A?":O6NY,N':NT->I5DQ
P9&\Z7IXKNYE3$J=L*+\I'OL[)TO.8:Y\R?\ >UJF64@OM]R&/\V!B?$C23>@\%RQ
PB.#]16(E=;APC_OG5Y<S\?5?0EZ[$B6%6<7T4[?$0;X@@1M9QPP;&79U7U!B5]]V
P>$ANU="L,]&YJ(3JNMYZ35TC/S"JTY($X=CT:'FC._DL.X11  ;<JA@1ODZ#]':<
P-!374ZB7DYNK/;MBUL*XJ:H'M'(:]L3C7X&EJVLESY7ST>NL^XP*K:FU\J(T4_PT
P+_0>L8"314LKK8"8.J[_JL,MCE<UR^ATSV,33UWQ^?=@:MV.WDU['F'JX5[</?YQ
P/?TP+<;$[$\]\VQM&2=\TY+SO?LF*8F\N\B5.Y]:2()0%^S%Q_Z'SN//;7IL8_B(
P/-:_\"<RD],D;$FW&1,6TO$&_UU'[A3@DY+N_LO78".]BB^(,US:XR>\O;_CSW^?
P _2B'X]DIH.^%B;1U?GI?36T<^T84 I]?*8ES(#^M16$YQE J<F7V[YDPEI7J -,
P,*A[B)7_PK[B_59'9=)W*/ 2,;S5W;#-4/F,=,_M<J[3"!?2^F9(I&G!<Q.9<QV<
PA6A"24BX:O>C#::_"8*,LS!"VSQ(4<[:._VKPN(]H%(D9<SI_%9!&7$/N!/KPPEP
P=G#QHS64GWZ4-PU9 U54 O"4*(AT;1:&!*?&9J*(3=G=?Z14/L^\LFED>-OKHW1<
P'.$ZLNF=,=2[E366M[A8)D+W3'!&(V+W_)TK-5=S6WTBN)LGB6)H;1Z@X/*89;E.
PS@"F)"4V%0VLN4]K,/42%WGJ0I)'(T$3N$83-E'G\$PH7"13-CBI<P4[0!:#OV4,
P6N$PJCD3>+,S)Z>,@08%2+9T[S7B.)X3*C"8@L;]H?TS@UXZ^ $ <-\F:3_19X)N
P>4EOA(]*'BI$J5R&9.6*QYX#KS@ : DE W\99(@8.H,APPD;0R^:#IN)RMOP 4(P
P#5/@RX>)C"EL5B[=?'-<3R!/@7Q'[14:ZN);F'.=A2%40<6:1PI)V.U/4V+6EI$@
P2UCHCY?T_W-+0W/0P)7;.VQ$F38#/5P_)_9U!\ED$/E=6&M@('-C;3[D0HX=%=IL
P0ELIMN:SP<Y2<[EB$JDG2KY^0^Q55]M_FQ]^&/GAI:$3^Y/><=\\Z!TZ)G2=QB K
PF:>YWH:)._QA7  [)I'*;SH;3JR?I]F7!Z7R9:79>O,4"*_G+PS-TDQ _)WB+'A_
PF$ZA',3?+>6C^TT]G5AZTQ9.[1T%U'N];^^Y4I"3D!3^T>TN<N -<4O%/%FD%I$X
PU+N*Y9L&PF&M%R<[VX;C_X768TX2>\Y6<#]I<9MVA38_#"M@=?LC0&G%W])!%IAU
P].6Z4Q11J ZYQ"4^//1M;F<V($QA_?7!R.?BS909WA$</QR7@ZXF-!K5EVV -T//
P;P%N)A[I >%M#CPV*9<SD.J,63O)Q0!^.[\9-F #T[FX@Z*)99'1'V==/!VTH.V6
PN&J-&U=EJ_) R\Z=1JX>$^:2$PVO\WB_<P%!%2?)UG3"1;O+G$C_SO(\ZR(O](V,
POOMSU,%-[&LPI/LS82+=00#T[O6\3-02:V;@LSQ@_2YU!\KOJ0$VH@[KJ31-Z=;C
PGNG4S\=[S4B\IR9AZR/B3M,'OS_+FJ#^7PT+(3UY-Q_F<;4<9^0"Q>6S>1+.)S]X
PJOE%ELQGX]V[]O^/;9%.8L?"V%J0@G:#/%I\RQQC<QUQ;@G+#@8PF(Y_/J2%'![=
PT$NA/>K$N6R]1+-(:'PQIB9FT 41)]<M)\5$"IQ'N</ALB!*Y4L*TG6SD-DE2ASX
P=B!%0G-[K!J^FK OPKU.(RP@.UD/B52/0S^!Q.Z;G)Q4S9D^O*R*';77SK'!:E?$
PBI#"?;/C:BB@1-=6'2Y_4%NZ$>#9(J?!8"(TCE.]5:\]U;>G%M]D9>OG+0["V39P
PC]^&CVHI6<)G-_))[&#XB"XR\]]='ZG;BF\50YZSO/B0+2!G17/GUO#H\?1F,-L<
P?,V'MCN1:O7%GM'\I(Z@M.U\&@ 4R* _@BLYQ>K6;#IGB[*J6^Q!E]0?Q+V)&6*#
P94)R#-$KK+Y:6AQQ/+KI+)VU]5NKUS<19>UZGDAK@T$S(-0$!DTP@^1=X:V(W?#-
P;Y<5>>*2RK>5.C0I>B6=9J85R"?RM@ %//X)V5Q^-,L_8F KTY9^BA:M7^3H ?S?
PRJ0 .G'1(1U2E4W?QK$4.@R!7ZE2G49%S8-ZFX8E9R/+B838G1 AYGA!(WF2*T?4
P<,..CY5\6,O*:Q<7L+A$PM!81+!5.G=_]1=5HQT:DH;).M#U6HO- ?VJ_O-Q(86M
POQCZAOQ_@2<54L.%AIXZ3[FQ=/0C3@7GU/?P6/6+RGY8J!X8F['0+#S,@N!T@QU)
P'>;_ (T"8%HU&Y2B"LA-U/1$YGH@D"_\O(OJ-1BO"6D5P!WY^3M6FLY[0]'*76#3
P[L^V2ZEF6K4 DGS *XYR;9)@RJ@+0WD".N&4B\_+5># 4AV\_@N%0;-C*"V."T16
P)$P9I2W980Q.3ZN[V=T#(:6A&13T:$?>_.=.+&Q6^/X:I?ZP2WRCCV_M.(2?WX$ 
PER>$(D$H61EP;-:T:^"&WJJIPV[Q0\EC26&G3\2_!SG)$<)N.8@6:8D2>H(?O2U9
P@<'[_PGQ"@_8R>I*[^$A961<#[@Z2R*.(!Y1AT!>-R98"V2J]&A_]C!P:12_$Y2M
POKMCK9JD^VX5D*S_&&24E%PB=#7]H'/XZ3SMU <D,@'%&?0&)!US U]JWP_*+O4M
P;T<^=7G$L@( Y0[OD#E,36G23$/EL]=ZC\6RI=IW;QSS+QH%<]SOU&E,I/2JAF?>
P!/[BQFJFW[-GSH\H;^GIJ<LJ6HG(TF]Z>=_TYD,B(!0</#(#1F6V6Y&9V0P-6LA&
P1#/JB'J&B"1?=^G[_=R$0+ =XS!I]FB"."-1'BO%.'VZ'&CS!9!P^H4-S*>2U$Y^
P_)F6X<SNE40-, \VH&/>6' KD:Q095ZE)+KF,XM+@#RR-G"@/;.W >BY\Q1S<70>
P&/M5VVWH':Q5P,8F(-MBTYOUUED1^@Z"W$?!<N%1M<1<!!X/0R87M[_F*?A?X>VA
P7Q>_.4ZL>.!X53#4.V*T764D="_G2XR?KD2$B3Y$$Q=C0T6[(SE??_KBDTO*ZA8P
PU-@Q+/>HJOLS>D2XX=RY(KV".BRBSA0^$*/X]/CMI7X7]=B+R? ZCR"N]P'K]V2P
P21 PA%*BUD$K+W9"42N2W#8WI>7%>O4^:?U?APN)Y'(^#"71X)EHLI1^-M01=:.F
PO5B<CF?0MA1X<I!Z@VRMH7: N"OOM6(@B%"Q1[T%%^E ]95J!M>0)?M5<DB?"?:/
PJ&N#V30*:BU#2Z71FT6[438: +UHYN)\*$K75R9<5>U&='";;VJH(*\C-2 5DA! 
P@)U7/=PZ6ZXGM](XMK!*0AQ$X>]]IO:%>8Y;-T <#9/Y<#OOK.XR+J,3T8]G]9QW
P2B/281'%SW&M 5);<V,614L9(!3ZE2ZO*RF\<8$^A*@.\L+2H9]M9G>)9H7U;E*X
P+D"YNVFV67F?&-F.,JIT.XU+$.D1Y8%5</JG<O+BYYE\1/6\@+4K!LT8Z,FY.+#0
P<EA@[:B[@$&EZ(4V;$;.1V)\LL(*'#P$'AB,@IT O:!NP YA<+QA.6R$<2TW!671
PT&RP3[:CHNM-,>E2,NAG,9^6* [=C?]7F1 B51E')% #!WCX%J*3Q )P$SUG@@=4
P9@Z&OS](J9\%W_17+(A*#^:G"6N6KFU2&)&CLYB<>A%=H?DQX*(^0[K)Z+O.\6II
PO0N^S\B#0(^J"%[($-?2MQ\MSPZ:-$I3:(D($U?MN;IUW<+)&L"Z RKG\TM7, V\
PZ+A/6>Z8_?:,H28P?RHDI7A(>'T>>IR\C9Q8+M1F\(Q+=AX$Q3).[?XK90F25U-<
PN$EO)PEYG-\#N80=B/+,%-@EWQN.1B!U*G1N8>03!Z]/HX=E*JU6-DA/)!5EAI@E
P Q,J]]Q%D'$<;LV:_"4&1[ZSLGA!/H=A7ER::ZX$F7V1(",E1HRS)I3+I7'=J4=N
P8U>4X3-U9J\.Z8>SC8+H#WKFX@C8=FDVBXCV2/Y,;WM8(-2F2T#B+QT\0"97XZW8
P% E,U7^W$(#3]8?J3++_^(<&)[0R1'U!_E,"/Y=!!#.B>21MX;0.:J-5$#7';;1U
P3&_C'3>LI$Y[83<EZJ-DI X4LJXAZ<(V^][IJ0)*NEC65#FTZZ(9?N&3I![!3.JX
PJ\,1B'\YX?:GQP'"MT;1N$59<SU-SLM;V9'9V'_FC&)1)B^]." <ZS%+7PAP-N."
PQ(P]/FI1!N#HQ'JCTM9W)YK1L6E' LEJ,UN_IKZVQ>US?2:!,>?0?1;8W!FX24/*
PMU"_'19/@#U1@=+=N06,VHRGO$Y[0_;KEYO73+NI^B;3'_W^G9/'%WCS!=,[X*?^
P(Z J'X^9V]I!!I5WJ\1LNJ_B$B+'6W=/^@0Q@^@Y)U?Y;(&<1JC-FO(1F%G.-8)%
PVZ$D()$S 0\Z6N5H"-W>1$XBC]4:W#+#RO1Z?=SJB.P1==N8K@K/4_@\K5!3FJ@T
P:$D\(Q8_317881#2:ZN6Y4X&3?"\!)D-8!")W#& ]DW]5S9G6&9Y*!/2'.-L@3M$
P[U4QH%8*QFD]#F-)0X4ZV>TJX(G_"PO@1!^NEL7DG5I(4T*FX]IQ&OH.T2,+=-[;
P @?#WSF789\*1B0&Z&S!H#>O/)BQTK7-6K5^7V*5 +*\-6&":9-_Y\CL[H$^/GEH
PN3_'5I?\F7ST]WF-:T.B2M1?S$D&_=_4C)<WIT/T.S^9%]#L[WP*!-H?;WA.)%!U
PTC$]FY+$NYA.=E]&9A7^PHMFL'"5> =]'-#MN>%\10E/L\H#5.(1R_<^.M3]T&2A
P;$5@^*6U3;0R89-\C,78QD?WB]FPW[R8UZ9M=.7O4+/D??;F')P&'W//NI!EA3!'
PR+$&1[[*C;]_OWI&^9?*LR$>[">AG8?F#.U+[ZJ2!X*3HN20\RN_6;=VO@E^K_4X
P)>]2",+G5<=/7;5NIEUXVEP;7Z-WR>/;P](1[)<!UU@:/GQ\FBD-G8W,(3XVF-/H
PB1BKOL2Y#SZ"R:0()]45RQ"R#TLA:^'LF'C@1G'FMN+2*,IV&(OZT&B$7://;POH
P--#1XX@>;#:.[+\^K+J.,=[U3F\YD9HN;)NY RD%1(T#S')!>3CW(LY/1(U9]?@'
PSP8U(UJ;A4-'CX5_F]@%35?;9<R>+ZE!_\^MT+1?D]2?CV5C.#6!K\PD*W 1\Y4C
P8^,10ZU=!^[:L7*L\&_]/:U.Q-[FQBY=._-WM7F4I"DKYT4XE,A  &L69=)SSFTF
P2&47F)M3:]]336P,-FG%E_;U3F85OIITW.#50;0;4\B8THE-V_>+UM\;W;%$TV$7
P\PNWB[H^T)%NFLC\!Y9_/C,;I2*W^?5FG#/V3QE5)(Y>)H['G%$_B5,"(6Y FN[[
P?L8Q$'#(4$F0>9M0_(G6/&]O)1:[&';*B(I.#L8SQ[\/7 :44K]07^E2K!R'R!'=
P[9%KN.+IKU1@4'Z6,SUP)Q/@V$=G'V HL,SBXX+?F1C0+0ZS)CP1?_;!+-2!Q)B_
PI'SA)M"!H/KXF>C)-LZZV"\,'%4*_Z8\MYI]6MW6Q5-X[%6]96H;M!VNB/0*H</^
P!V@_GXLZ%BCPL F-01[;* 7^I$%[C%E.[IY3*!+UX0K<EZJ&96H]C6KO@A3[Y,M.
PA@/,VX%'C/^B_NJG"F0:IW;AF=;F&?.,;:V=[-W("WJ4\7:?P8+$N_'L[3OZV#D]
PC!AI]Q@UP?%/39;\+AZ/5!X0D=#R93SWZJS.D/=?P*Z77^'F3E9V]$E!0&:+V5,6
P5 =-]E\[GW'1$"^7JZ(QA]D1.^5X_Y*4J:UX&V7T#Z-(IN)R:FB%&?_9TCDV<L4.
P\L#86 N  =*-6ZL>+\#JZ"E/PFA.K)T>RZ&Q$:YD=$81"V]M]C:;RZ5S/5DEKXI"
PO):D(^RRK[\[B:OS:4;9W"2]C:OMA.LS6KY?NV$N)$DX+G.3/2'Q)H2@ /11(KD!
P>VT!7K;L-<7,XS7)S,U$"T9+6NDG!/EO_2H]-ICWM2JJ4/I=6*#L$/;>=)3@=QI'
PNMG,_5D$U:9-L@4IVW,2=AUR"Y&B1JGI(E="NT#2]I5*)@9=/N9'UM/\R9?>LS!>
P:M[(XD4 *'T]5^R*Y\>2/4#3[WM5X6V13M,$:]>WP==D*^=F[-5JR. CTK,QHHLE
PVLV8/I"L7B\@%J]618]<I^YMAAQ[+!W][S,,8UE)>N E9.RM2FNK$:.Z3R7:X-^)
PY_SW@X4;NH8/GG$12&<="&A\S^'*XI_W4"_7N3V05B29$>[$]+=3'\2V]D*G%H7K
P"9]RZ:44N#U6Z)9INZS._.OHN-+V<.K9:R_OCV?QKQK@:;[Y!CY#."\"^?6)ZA-5
PS=H*N9Y@?ER$H+1'0>EA8]+YJ,%JLBO].-T3$<OB3,'+5>:LS0[Y,!O SF570L20
P']=<+[J$L!3?9TAM,,H;_'=\J-X&ZQR7X!NSO(A5H]]DZ',$X_:9(:' 0V1:OD$ 
P%UGTZS4<_UVY-*/K6XWD7FE7?J3R+N\D*J>RU7$5]2@7BV$GSXY0;3GY7%_)9[ @
P;YO7P6G2J<G^8E>)5H6^&1T0-\\G[_M%:7?(>FF^D=CUP2& Y@02ER2,*'[XZC=K
PF/=2!ST?&(KP$R)-RC@BT_<9V^X7,*1;L;7_SAL=YMRW+DP0'K<!MRW)K TSEJ34
P#ER@'81OTSP0 T2&$&8=H"BDPPAS[PNY2U6[_#E<4SL*Q:C5Y."A3]7[S+^W3PA^
P(E(K!:Y_PS[-6!K=0SD]-O1,D@]+^CM!ME4$2LTCEC) WNP426Q[?@!)N)^K<Y&7
P%LGV+WH,T<:KR\LXM]>(BW2-"*T5OKCDBPH+,RF7*\T,U 4X*?Q$' EM:6J;C\Y1
PD1@KX[18E$$:<N1X-\$#P4P'SD2\+U#H!6_^6\[J+WBN9VZL [\A+2#7G#E:O(7&
PN@&Z!R6SF!5JP5;8VDM=0]OIK>47*/EMG. 1ECT#^%Y98PV)>)&/+&@2:H7&^;(3
PQ;4XKJ=<U:>AH:9&0B+GDIR/ZJXON'[JL$3&%&7"/L1Z[>:^&.U\ R0 _[2Q#<G@
P?]?HUD(-F]" 8%[CFR%H<M&&D_)E^[G''8(7;#5@&XV&W Q$!-S-C&#.2+20:Q9_
PIJ7'3+U?;6/BA,4!B#U:W[P:U$N44 ;2 ^U?!';WK)R!M09&@.6&MLSH=Y"N&+8]
P&:1B='QT*QT_A7/\D^%:%OH$'I\SI_D9TG[+P$FM"&9LS&. Y'XOC0RSX;09COM3
P\8GLBYZ^<F 0Y9-2/3I!:\2C(C?R5Y EI.+VOL RP;TG^/!T"_<K-ZDQ-RC/V/C=
P$4*C2V<('17*&CC,YOZ!,,'O_RB@>O_T4%#S5,B%G_G\P8H)@4LJ&\/^Q%*8S@2S
P+'#<TH2F >X*YQ(/F%.! :+ ,&SWZM/OL!''E$E:XNIBSP+)[MJP,W5?J\^XBM>)
PWK83@-9M #QF=UTUS)A.8"&Q_>M9WFEB _9F:EUUV?PC__U=>'Y.@"=NHC$W:OOE
P^/1*\< "Y+J$,$23C-6E02P-_>T*3HYJIB8'O0BVC"0?QK%(XS):R3%GW0V_0*DS
PFCC3KM/IS*0\C7(W',=.Z]>?,Z7TZ65*['W9\8(XOPMS2.PN*]/B<C,\![#[A3.8
PX'M^0K=BC+:\';Q:U[;F]9M<APE@1K8ZSGH=E7?Y;"BRC_# ?CYCB0[\\!#% M5#
PL2WPD#[Y,0L?UJ*O$8"FD(%F)H2,' B%@=HPTPI]Z12F*I#MMAS$L^)/S%I\#5C<
PC ::\K4Z0)XX<4G.=#F5/?1B7:I;HQI$Y_:O":A+Z_2%4&]/ON-N.P40XGJP'%VP
P1DZ1:]:0C2VAPT^2LFADPIHBTQGE=W-^I7"AZ;<I8=M^/7YB-F"<RF:+\GT#C+44
P"HYW?J\0K>5).GJEX!=)_ /$^L%>P4![WJO0"<XCEMB"R_?V.>G=2,)2\<&II"O@
PPZ-2 Z9PQ_CMIF XW&*J9IUK.\3RG2U @<V2V5.HKE^N_I$@I[]8-*6Z:6O2 J$8
PF$'G(ECUJCTT6$G:F)(?0%'/!8K)? TC;PNPJ*:.-(USV7(J?M.)9R[:,=X>5R'<
P7QV,V3-.0M(^23#9_,ON*ZR080@M;-H!*[@_W"!B(ZN0 R0[ 55XO]38O4UY/R!W
P)&K0/E&I ;Q73Z$,_(@6)Z](0;+WNDF0V-EW>4Y%ALFAJ8U&R4^#LT4PZ\AEN*-&
P^0;?:,"B*R8P0S%NHH2<_3[;BNE<*ML41=1/EH2'8J'>]&8[\X%0+48;B/3F&A91
P50CE9Y<968R2QO[L!32VANA*8&O,[(*R/F->]9GNL-)-@1XI5ZCCR8+LY:.NM2&Z
P0"I,M,7,"';U!?;R'V#K@%M;=\I;9(3<&,^X9M@H!P4RB<7=-'VJ"[DF-.LLA8B+
PZP$^UH[GV^)$C!:3",VL&TDIFSGX1[-#Q_PLYZ C/8\'@7]J0-T<XC=R[!%?S7?Q
P2TI.)V/RZ9X12ZC+LIDD$2?\;3)O[J1^%J-A8+%TF=#$5)NZ'9U_T>=[6-/D5LJV
PQU*/6LG<T%NX5&LJQL']0'J_0<9S5AHR'(@\FQH*Q5LOPC@\ [0_P^ S/Q6 %1?3
P+4#\-V;EE!97@[U;& M4:0I@26CMM24L)($P3=9/)4V1K[9*:.U9GF #M, =T94F
P$46E<5]NE44O0A+OYE5M@A-LG?K%?N5N;:'O&;-Q/D_LI>0C00;EG I@/X\&2]@Z
PCDY)*+$87JO+@H!AH74U\7+>-8@-<C^1B8<)Q^YOJT;W*J $<$HU&L2%78^4^6;J
PP#]U-8WE;*U,OY7^XF4L 413OORW8FA>A"UD; >5KT->+%38>JOJ4$8J+01EHVVD
PY<" '7;0536=V)$7(PST.<7.P9]V&6((KDPUJ 4/RD%?9.A^R#0FOT-/L9<OTK9B
PGUSS9H0\OB@#1.&DFGA0])+IL1T !2\F\',VFR 3/O(_3]+3\M;660\B,\>;F4@2
PV52@GS/O7TI.CI:_-M6-$H>KYL68+A\9EO:,@G8.XNSLQ?O'9E?"M4%1XYD2/SJ=
P8/C\IGP"'C5\"7:R&9D[Q"68858L>0.P><Z*]%A,Q[LEU;)!X-L7-(D5E4B7(>U'
PG8+U:\1@[9XTFEDU%8O"%B$"%'/O5CA4U$09Q\*"KHKUZW(_[)/5.+*. $G<,IFY
P2[#1.CM8)[8V@S3?S;KT5.":+<4EU<*4K!JQ25FC!7"1]//%!;+0:6K_5P'R)T.P
PTT *!YT.W*E /ZMZ1HDD>U"<L@?5W>B1*C]*I9/ #6D3,3(F'+=A^30.0*JSVDXJ
P"8C,&,'2)K/%QFVAVYZ+P4.$]E97^0=&MF",RW )63EA%1=MRY;S\P?K-8*=Z!TE
PT^R!F9WPGWXX% CL6N$,!FMMGL;II!VG DJUBR9<W^P_HCOB&4X-?:+8C:Q-KI9"
PR$+)9G'64MH1*GC2\O9#O#M(W'-; A.R*/7XFFAC1@<$I2(KE:%&\NY3QDTL1NLC
P[%M^2F0FVO75*:5E7+LI!)*3_RLW/;W5U":>2V)/L$4JA/.903AFA.<IN\XH,2_L
PN34(]ML@V4'$!47W"NQ(ZRX#5,W+B7%"@L0JAJ;=S?^/;LNUS1 0Y6<N,(?'8C+N
PU(<RMQP74Q#*[0WCY%"ZS>(J;7#DIF((C6*(\>KP+!EKC\$'!-PA6X6+M\E08C5M
P8PYNS755E*=OB5"!,Q-GJJF8SO!6ZNQ[UN_*O>3TFZ='/NO#B8?IG7K5^-=1G-PJ
PO1",^9Y8/#3%F'F//?#_RB%2Z+W'A3[(T1'&;.YL%IQ0A-P^8:F[E6-O7WLO#L&5
PRB))_*'T'2^H/FJ<0TC%HA=%1'(YV@_72B0VF+'[P-.X2CG"7M%IOENU"W^/@V7U
P<&L*'-24M">2HE"9IG5<D)!0\,".@>@L38/N*W6!J5E1]HWLK#;$WIOW&)83U(8;
P5X#:'IW6*^/JOF$YNJ 3#D(*A25?,H9T04R@&KYZQ<-@8 -'#WM7"!:,]A,W-'_1
P(T! =%T6"W02(1VZEP'W_P-[0_7>-9WROQ'5Z#99H-:^#>A/>M99(AVZ(/7;31U]
P1<#8C3)IY;+&9"EY(O0GP[)I?.[4Y,ONM0V[VS5YUR-!9Q$!90?K+ZC>T(96ZH-Z
PKYFRR(D? &=75BXO=F5"M1N;%G;!_?V:9'!%P*YCT##2Q96WT.)$?U]\&F<B=Z?!
P]N\L%CS).ND<WRH6CAGV^N7<%Y_FT2WP.]_3;1O?"&'-;0[8Z*?N*T&JO@O\S*C(
PE$XQGH<=,=WV)P[32@7@Q0S)G(=F8T'5[+ 8=W,<# ?(.5\8;D#06Q$&T_JB!DKT
P<,58*B)HX_W>M[NJ?AWGB//0 WHCOQ":5]Q^PM7!Z"8;)K[2]=>8\'Y"5QQT0=JZ
P,*8YW; @!7:G6T:\DJ>-H9KN-"VQ7SS\T<;PU#R.E]&9&? T^!SS:=UZH7!PZ!Z2
PYM+^%6GP)3[FK50'(4@C?+Y?RN(AW'G^W=>[3M9&3%(ZK2V#>^V06*%[4NWU%YG(
PZK7@6HTV+\YR5XK%U_$\WFX](1O(7*DB&Q7LYGXSFT%_Y49XGL4KD9<4"NA]UR)>
P)((4.W[;'(>9>537->#8LN;3R,- G<(;?C.<5V_VJH!FA9 ON]0E:W*(?PHQ0$LQ
P_^:74XE(W\HXUK170T$G;&4JXGWA1C1\FDR>L=*;_5/8G::Z0P>&4DS,;&P50 YQ
P0C%JHRT-KL\%"O* /0.R$-'(UC->*I1;@N/ 3-F,PS6HN@8O(H.7HHQ)VT'[R6'\
P[072R /W'.(F4[::X0*-C& (.?\,='*5#NMQ2EJ4'!;YVBS??'B]]3@,\-;Q-%XF
P>;1M +YJ8.J*M2\DKI<0S<D-\8FY!R&4'[MNWIF]C9;LU&_R<9T:QPQ&->%1Q]$/
PX<O5],6MUT(96LFO8%W']+D0U@[=B+$<94FA%JL#2LAMQTED225-BX4^U,#?QZG!
P2&=;FZ.*2&^WI?&R*4UK*D4</4%\'T/HY@AIEN.)W))4U*H*5[7\-<X_+S\3@D(L
PN1R*UP-8JH6&P2,&5:EBB?H)/7O[+L\%TLLB"M8&RM/05GO-5#G^9-* 5J QGWI:
PQE(V$#N=W$L*V'70R<?DWQ%S@-4O/E#'!%B8QWX\$X!"+%C>J*YM,Y"5ZO4 TG; 
PO1RH,LI[[;>/H;B-31N#MI$/*O\B]-NNK\>[XU\C=:KY!M(%-=7T/J"'_RV0LTIV
PFZ"R%<W)93T>B+#QD!U'=AB3OI( 'W<C8X2(&\S-FV!PT*!E\LDTYNV/'0T&H.6I
PL]MV%70J9N)>PUM+VLY'=O&>LM;V!:K[I%N1+4LF0^I='VW8JO%/9FX4!Q49S%E?
P:=FT7G%G!_H61;Z*JL$J-;CT@1>>?W:!@RQJ"="5"_1 <*'T>F+7(#'3EJ,W0?A6
P;2PAW+-<(!= M4EW[XMP#(\-C GF[# ,*'/ U]U1PH5X"U8@*(E@'##BB==@"":9
PQ5N.,:.KK>\3'[N.=HR%>[/^OD3N6BY\KLS3<@Q$.]P-)8DO0R^1Q5>'([\M>U@U
PWG?PD?Q8D]XR^)*XV6.*24A"],$P#RS':,-=>\0872&FR,>XXH31?+;.K-;OA_"6
P$+5^%%?K79<X<M$FPZ^ P((G&<6O:9RCVBO679L<U)H,,G7F$H?E^T4$YA?+%_>Y
PQPTOH#HAU,2V\Y4 #!N-!3:+%?%S^Q+%<VF@(M/@MGZ8=)5'9Q$)'BJ_18Y6725%
PDOXT$,8XAN$#H9:%UPXFH$+R@;DJO]P*]O^3W_4H^W,B&,;ZYAE+L:G28>>_L6D4
PCU+WV;!K88/@<']@(H'E!CG@ 5]A.6MV._%,! H]+1@C#$K4B1YKH3?V*!F9#"]?
PF7YHR&[1IU +7QBU-5"8*A(,MT2PLY5 UN$15=B\AF$#4,?MBX)3)A0GU$##W&%/
P:D1A]<C=MRGJ,1@7N^2<+>/^_!\[BX\D"J@FTT9Z4M4]-7A?1O[J1*W?0;##DU#I
P0[PD$E'@*R:&^(O"U#:",6R+*?8'5RJ>I%;Y3^7WD ?KHH84H+DF,<U=YP]SG'DY
PE3PB&5"_!&^;L2:]NRQ>OF8(.Z,DUWH#LZ(&KA:!^K]FD)0@Q2BKWLZ;,G!Z%+EC
P]J7>D)ELD]!8'<7].XX5N1LW_)^C-U('"5RZH_<(@ *W=P"BAD\G@J1.;>)\]H !
P;1-FRYJN8)C(N!G>._3>4;YXU1&C4*0"E.;H*@0S! (.:LVO?CIKL:P@-PK2KPF,
PCC+-_/>T5?/6Y(),V=XW[F+* ^*>C)8_G^KSSAN#"7T6:M I0R&ES?A*+8DU_RHS
P@$HE-QCE_+GET5[!'>M7]-*LR"^J#+0\T4+#.GPVR9P@/+[3V*"0W#KN!)+"C300
P(@6W*F)(:=IID^/$-+8Y-O#(-ED@VNH.Q1G47]RNA(!%H+;+%[]43-X>TP76 K5S
PJG_ =),Q]$Y(K=JT5DSSYL\S&J#C4$6*F[FG=O%NNR2>,N?9)^*/Q9:Y;"$8+]B8
P (UHG]U?RG>^W93/X_\B>M-9I @XCV]H.$[Q$Q!BV\:0QPOP\VJC>@+Y52ZU=?)G
P7I\A'2YCA3^ !*0;"%XW/>MQE_/A.73HUW$0R3GG8'N"S24MQ5KPCR5-0SNCST"*
PFW]EQ/D?"4;J12;=LB*'"ZE)=4M,(M62][6UD&< C2:K*^]'LHEHE;8'O&<RV[69
PN%:&C:.GSZC8BL=FA0(FO\L8.>RMF(>=OU(F-B,'9:1CB)F%!OUL(CBC;G8A2(TJ
P19XZS:7-X4FL]1#>')+H6X2NM]0_%)<T'?//!Q'KH,#+X!PM-Y(E4&63KFO:MQVK
PEMX%65U1L/= +VJ*OTZ]"XZ:C!?JXY7(M-=G>S*&KRK*1=KDDY^YLV;DXV*YWHK$
PP>#(BF-?9?AS5E.PW-856I>].BG-WYFWY=;)KX>V."@]==0.CG32Z)IB)BP/-5VL
P(^O^_$=7HDP_8U(NZ]L$,LPG6G&TNE47;KN&_;X]B897V17[PXK3EZ/P7"JR56A+
PH(_-]^!_*X4(AG\:,O W=(*H/3:\ZFA99%J /+!UX(7HTE^=YD79RWX3'J3;+91B
P_&1F6/7U/C9\X5>6UV< >=Y)E-+_5%!D:88C96^&0MC^6%$"6U\NKRDJ8?X8;FTT
P8>.M._>P;_'P,6]:E4J[-YO 1R8IUR?T276-!*NB-PP=%/YOLON+B2TU2P'F=7IW
PEG@;P$W&9*ZSR@M8G'N4H[6 =I"I!B'_U FF4I[.//^?A-M&H0L0S4/>N]%"AZ__
PU$*U8$/<HQ+Y,W6HXXA1!\B0!@TM'4 M'HU:ZW\$=M_G!4G!)0B;E3"E^%2#"07%
P6V>H+@H"J5CHF3C@R,[PT?.H^EEBFPX:\B=CW)ZE5EAO>;T\&RA&+L_R8JB-L1*Q
PP39F%$^P[]A47WMS5&AX*3 0FT?U)]A.])'S7+QX>R+LQY]^KSX%)O-/9)T<H%9W
P\ _/K8R)]SH&:^^ZP1MK(SNQT<*97B\-W-GGD51/S\)(\O8\X;EI#+ N_QZ9)R&$
P/Q["Y.&G2\9X$E7"@_BI:_\Y'T#.<=OVXRG@MOCO[I!"^*1W:O"@/3@N8,EV<K16
PI;9W!"KQ*Y^/(P"W>[$B20=\%D]IO,ZC72'Z=!ZS/+\M=Z2X/3-7VX(CCFF/CCMF
P92\!$$>%IU:OZ&GN/XA,LS73_1"R8^ZZ<"$./>_10\GI3&W*%%M(K2S55=#/<5^5
PA/DGO0HP$0*8?]V:;7)K5ZJS#=&!GAM23%_TBIOI#BI0E^/<^3"5_/9.RK]H4:=*
P@IS<WM 4VO*L-H#-#_66@_9_B&3/S9"$N>R]4\+GP+>@G@+1G5I@Q<QIEA[,Z0'V
P[H;FG<+YCR7W+P"@SHLH&,")M#)I@KG[R1X]\UH6R_&"NBA_QU35AZ['!Z9'TT!1
P1ZZ2UB1TK&Z8-98@)$]M3(+H@;B(T/_BY _$WE']6U)8,U)^]JM&@^]EDK[=1!-B
PSL4F\1LCS4$29&6B(5KMT;/R"PRGW^B8GA [EOFL*I'5)2"%($!;T(F\?SRMM?V^
P4LAI*U- VEOP8*(H F U]IEU"R<;L0S*$*9N1TX%1M+N_FW J5()I::N0;J$CWX=
P;TZ"(NUU7?(@&?^PLR^;+K4T:E^CBD1)RC$0!)-^)Z;:/F,=KW\A+6NO\BZKPQ)+
P)DX<[-1GK*K4*4]3/Q.UZ:6;;3$W @= TQ\Z/M%]B?J&M*L)V#]I"%VOUG'3!AH^
PW=0Y<62%HLY:U?I%#"7:OUG3>G,GRNPCO+5_=Z0 (T%WF]N@HEY[Q>@67D>AU 7P
PC0"72:3N%KB$_@CUE:F6:M?3OPL]$5,#LEU0%"%-^GU]8_QO_C=J"GLFL !ES)LN
P<I8]U:';4'TW(@==L8I6VB&?;.Z/IYW6@9TQZ:8<)O*\G$H"[Q5VUA*$@W_V1JX$
P?:R5"L$W/IXV=*V;9:#AN4S[2X-R.!N-B^!$\:JIGO#!=5=X,(?31G6D^O:9N$6W
P1#*E2;5CCQN@\Y#K+8K477[VN_<T.6A8-23&23J:V\)X^LZHV%9%?\(Y[S"EV3SU
PC5CCCZN$[0M>E!\#_\1N@#0WOQ!0P=KHZ2(X9&@T)F'E7I7<"IL]+>+A'3('O(9>
P-EW"9 6>6W H/GD\<CVJ'+*#U![RE<F6;'^;N[[0,0DR]AI6^ XB>$=H:"-U+?J\
P)8P1W3S!K%R#$OX=*88<MEK^PH*7Z[H94=W_Z36\O7%9#M\(WYR"7_VDQ$*@NA#S
P7PR,?=D!I!D$CZWUQCK3BAK$16:2&-(<YD^#V-"7 *&:*]/1PG0B:[3X#J]2TTO$
PRS+(,>8L)-'8!D^;3JS@"(3;6(1NTCD_1?,28?1$NX[W?-.2U^6OW+MO=3"BZ- _
PVQI^:I-W&K#S209/^J]TR>P:$O(5STB!\G1-LM5^S**];9B2^X;E,1:S\K(";O4D
PM%X"FSH-F_0O 2H&0@8)L<,J@0&*1T$2U,=D$,FIAEOMD#?W.^M.4'59,\%GRG$U
P9.T!Z;E[:*C;^T+95=.LX) 9NU&KE?H78X(86AC=_SN0//' //#@E3.4<="IWA=[
P5;&"8SM/N\0D5$_8@:&\C],H"V( 8B+[H%5UY0&CN=E\V'\:O7-?<W/=0C&LM.G^
P,[B#4"UZNRGH5L1G.D@N#@H/'B8+J.G5X=IP6NW_(5_;SV7,$^R35+M^Q;N#Z(TG
P8V5.ZC89GQG)ID"I(6V/XH4/]=^"C(;E"GN*$BM3@!S]$)T_DP[V7U98-UGQXRT,
PF8 6+(%=908L&9+![.N<=O'0$&F+T]V^N_K;C(,#& ?Y7<8[B\_^Y\;Q,HBA@LP(
P=6I]QX[\-FM5' DF!8I5WU+I6@%&UA^;OE8+,=%?T2QZM%$,4;![7KV(+]P76=?)
P621J^<G3;X@!Z>WEV0=AMV32*M)%UO%&8@RKIH!8I:&W[(S(JYXHQ\%G;FW1M"=H
P@NR3L+>1QH_WR[&&&L38A:,;_)M*/> \K$<K76!L%F'(NC5/(W!E-FH%* )[P5&@
P.B<GZ*;#.Q+]X<A87V^%\07HD.MDQP^SOJL>9%\O<N&['(-LPLA+6Q"$7J4(Z:DI
P S<)PK4(K)#UTZ+3J97DLOY9,]RW]#;+D$=RRD/R]@#)>)=/+;8L+_!6/>_'*_0>
PRKL8[;5_ ^*MNB7$N2B[H2 O<I:: [3'/CQ@-U7H0SQ_A9'%M/%N'*@24+/6/B3>
PYX0\F6U4GD'K\>,/C!+/NV9CBB%VW\?5MW:OL@PA5Z4QWM^'*4@.F*_% <CR%)1C
P!#RZL>>,46+9(-" /]_/Z++,9EJ@H$J!'VNR7LE5&??SZT,9$HV"-HT@F2K-FC!+
POO\MM"*S/&_90M\WOE339\!=/KK+XYXGH:Z['XME=6,=L8K"">D"KX37F^1%=8ER
P1,FJL#][UY=XRFEWSXW>C:5\\0M9PX?U^XX$X)7..&MJ+>=?%OZ0R01I0UA4#EHL
P%1?&Z>@Y.7F?<X1V4JM_5;]@E,"><K0Y89;._Q#%].JQP%>/:M\<BEFB7374=[VM
POJR@8B3>J TK@)C/HG_:[FI,O%:+=.=@WMYDL$M%5A^(@\YCXE=>$(8\Z<I.9/;J
P3%%+%?BV%=_<573+OJ1HDG;XFHO%,N+ME<%,N(>_3J2I2<$(7R-\/W&C,H5.J_" 
P2;5^2#7IH]E?N\Z-:HX9BT'];OD2]M?"HEK1Z?\&*'L%NYMK\'KEEH93'Q=HL%PO
PO8;5JTX!2(:P5^XGN1//WH;$,5WAVZT$,<K?>;HIZIF=TTT$FU);+Z1GQF/ZLIFF
PG&,:">1!7(GKN(-!F+"-[.*[?H\\ [)9YRUNF]4VMML>2MB+UJJ2,RMLU[(+2BL<
P/0Y=CB?H$U[@TY<F(9,%^[O^?()EA=UQ$%"+ONA=!_/NJZ!F0R5^A7/Y%,>4W1E]
P]_YMB[G5OD1!I4UO_!5 E*-%9)2!2O>VB.8"Y1YE"*H))!N*<#J(GLBH]N5\^S8V
P6#$E5&1HV!S\8JH6N4"D.&OS.Q5/^*)/;E)7U5(*4SJT(X':K$*^XN:V[+8CD$A.
P7PE3O9'CXX3PI\X#[!"O.M*FFBGB,]1+0^\Z]O#FD;77PATV)";I\=B1I^W^-9^&
P%O_QB'%8G^/=IK=PLU4>O:67 ?OKS$U6;1]2*#A[2$(S@]LO-5S*P^QD96_IIHN)
PWU>F*<B22)GA28E(43&!%_E6_5&"=T3' %A?^N'7[#W;!7B]K\^.$1"H(+'2&BXO
PP3X835S#!5J:O\>I+0D!OR6^2+Z0 TN(2LZO&\.C!X5!C@UPN^-8AA%%1Q1]HGER
P!D_QS$,(7D+$Q3Z4O8?UJ_66X:G-&;(.2,41-H<@(\_O<GF'4KPN7[%2MAN:6=XV
P7\X!8&XF+^=YB!.3L50#SX:.YO]T=9?"EUT(B#/1$B2Y>Q(HN?1<KSB _OOMJ'JP
PJ[ALY*-SPT8W^+N#YI&I) A7'Y-F!OP2)Z&T0WDH$R*%LZ0&T>'8!9U-_\5M1;EY
PQ8XNXY J%NO7C1W]"4DW3@MDO@2_5@;IZF;TV],7][G7JIWYS^BBD -*L?K1:R;,
PMBDV%9?!KRR'-'*D8*=GG6BMC0HJL^)GXZ- UXOJYBX@YAO<[U!@/\A5N%H4=>@-
P)N>VH[E=@Y.@P"F[8H-3<> 2%I)EI\7B& YV<47\Z1#TU@N/B,-E"#'5'6&,1SR3
P/7!:09RNF<-3@PJPZ(HC_34(IFL%V 29/>^T%1#YD/6'E*8U?!:(HOEGM*EIK6&S
P$%\DY6U:SANR 2"2QDKGC,$(U5;%:NL#2GW+>!AE6.PT+Q(FNS,>)N49&;I)%F3>
P37/?P2MOLZ!?3?!\J:@S1BJ24,CD#O#1LI'F:;TK+N'UY]=I4]ZM:<EO#ATJ:&0B
P+O;A3B+_H.#[MTBXREB1BP]K4FY2OBE(&9Y6U9]M86ZB7OF<%UL&&U)\50E-FVA:
P7^)"SD<#C.]8(6&#8GB/JA2[0G(D,0@D2CKZQ*:ZOY"A BZ]F]*M8CC$_XDZIZ2H
PB*!A&%5)OR;36I1J2S>?;/6(\JV:4&CQ=ZKOEGC)N R"<#TLKYK4L,>S]Y(I3@MV
P@JDOVWM3)&IL9$D$P93,2IDOGVZ]H8O4FM"R2!DQN1&+_,"SA2S;:3(5_6B!+ K:
P5KS5I/(">1=!?O2!KZH"E-GQ'8<FD8\507DTTD$9(0=I</RAX'$48DDC3Z;7Q?[/
P@&DZND/D%&P]E#KH7%-JB]%ZX02E7Y[>NUY+Z?MWFHG5W7N5#'@GQY=D!Q?(W(>]
P_X-\8GYTLE*9,59NM70]@]K:%)ISI&0Q-70U(Z=+3I[4 YJK@F[O,PVN4S^+S6+3
P8()),Y7X/*[YBN]/]G)\+Z@E&]X;V<>ZS:;((<T:[Z>I*Z#,"CY%J9G,Y+[A3:MT
PLL7\0K&H58'D>=VH%WMR(K]>47.!!?IJ^1Y@7KL Y_=$K'./_AW"$B]V!"'.94R0
PD<%R*R[HBQXONFMPS[(CDF=SP2P\+AS&GS6D[06816W9/(AJ/V=@$#RC^+EBW/)C
PB2G#=?7+-?665C2D/9BDR+V=LGTG^1  %%\E*LH]/OWUW-:CBAY:Y!9+].#]L.P>
P#3=F')YG4'P-.4_T+6:X;W=NQRA6G$4DZ,4')A)^,<1M./T[(E8(SR4%J]FI>R73
P=O%5+E>.X:I,@LV*T>S15:\$SP7"4EDKNH8Y9^ ;7BEQOZ"&<+0C+<:RQM1^0K1Q
P\G>4<')ZLY:'/9\8NB6Y*(9WK 22IEM*!EUY.BT/'8IB]]61]@RSG &=@UL(C08#
P5839P\P0'^.P(%T ! GA?V\;K^[M;\]>3BRB(7^.Q;"$<2WLR:XB@9?@IX3+C=;Y
PU4BVKR@XF0GGFZ0YT2K>6B(ES"VR@9(6@YR,/,V52(0-)W,%NJ#I7/ N9F(_34((
P2_X=Z-"[\B%P3/D!,G%>W&0 S_I&TQA\AO[/&V?'*")\S[_5)X_?F"HL&I9P7CO2
PAD!Y:QX+A/.XKXVZ?'(D2O'L"><#-%Q#VQ%LD\9\ M8D."<J1S5? K*1H4'.1'Y&
PPLMO=(?)8(LW4C3R?O^^T606 #;-+GNA=.2PARB8-Z?\"CS'9A&^_O(*:9"68:[:
PJ,)AY&K!IT?EA-RO=W6!7:PW'H 6.@\WJ@B>923UON/ X<![>$6\BC0_VDFB.9A;
PRS#H^WGS/8D<;D/.BJ>*K^VR*ES0T#=:\(,/%!E;^XGV.L:4_!B3'R;#5<*W/),P
P![<NAJ?^?X57N>C95<0%8LS7H33RN"V7 T[QK;'LIKW_4O&6:T\D(]6$$[ ,Y;18
P\[U237R_\V76_5DDP[D!$<2KB88R7%U?S,G*5SL3AQ_:XWYGJO::[>FNHWHRD3&0
PWB4U":1-%:\M+^HWF=0=@);CD"3N*,=(6@+I4(T0M ?U>WMCP=[2[XU4R1BYALJ<
PW,<3.0?5) SHPDB,/8_O;5S)K"5ZF[K)7N-O57#%BYMZ2Q+K'X0-,C[[(N8B^O^S
P"TBDASBI>AAF9A@0WI[AIYRE].$5PF^=Q3)W-.VF\(-MMB/QW$))FP-;.KD0*@BH
PINC64\,RF>"Y"(=(UR "43&K1)$=SQ5/KK<KB6F@#+_8:K&S_V_/J>@=P8[ZK.>M
PE)&.B:KB"K!O^:JWD#$(+#]V_"M>QB^>!NF:Y$02T,@OJ&!F1#8OBQ+#7,OF"PH@
PSJ%-&%(,7 #;H81J@$!X3>S)U-@YACT;URNI4R.T_,TU=TZ>G1/SL1;<\>)XZ@7P
P;;%0'N#JN-ZMRFUCVW>O8WV;N63,J-/CI0#S^S82<H7GW[1E*/!21\5?S=/V7'NN
P/]E8+/15=ALQXFGH/P%J1 V@D5$R?5]Z7W4YZ!IK/KE9RB/B_>AX$4*5P2<Q?\O3
P?5SJG80D^<L9UD&7&FY3X<C]3&2/Q!O[,%(6\^=W02A'2Z2XP@T[! NDS90:32__
PJE?/V#U<+_-WHH$,O14_>^V49SY6M8]2:: AW14D&0+AX#L7041AN"\ZR8F=H*?1
P$:FK@6H547CJOD9X:\U<FJI4LI!-V/W87BEU7,IZA^YUSIS<O0&P#-P\#RH U+/X
P\I&((=H.9\<EM@V/KZ.-.@N#0_WOD8X:<;)%.I:-$QAC*>84:$=AR@4 .:>(FTXR
PD(ZXIWM8"J4Z[>,3Q:8B;X4G"VFYX>??YWR-3KMK_SSLV-.>LQ832^G.^@O6D4<S
P2_B7[?IK.RH<V!^K+RO9[D 6V!_H"X!#@QYNH<K</G#>L8K)AZHA"K3D&30<J?U@
P^ <!S3RJ *"K_RR<7V[L+<>K.GD]!V?+$;NS!+0:S-&NE2Q64<.H<C*9V?.V^E P
PP$FM S?N/--B0Q9KT0CDUGG@:]1Q[&+(=+#D1X[,]#^@0'#YC^08U_<G[UYS0'2M
PZ0GI1))?A16QNOAYVNC6SY0,/\H(W& 4FK+-J?/RQ'E!0@>'LAYXLO_' R6VP[6.
P1L+VY,UA>9UWQ,4K).<#^HZJ-JL)F8MD88L722**2B]$^ V8ID=6HDGS ]B:=K8=
P[R!-1I/<O.(MS4W-!>(&Q?'B& @SB,W'>>U3X\P5!!-68(RK?N60>VKBEIC E::4
PH6M"2I17;;]=8H9,+O1/)+2(Z5ZA&TYCJO.8*JA0<1Q"H8HGQIU7ZQCL G%@O7_Z
P+VGW;E/6+%^0B$*E@<U6&X9M!XE;?Q3&1YAUC> '(,11B'X:+W4Y9WU-84;/AA:$
P-)JQQ*NZ'=NO\)4+W>"BG9A'XR>$'C;49$LVR5XD.R["Y0-H:Q+%N9HR#W+X&VKA
P:TS*SY&"''E&<K!V 9!/M#1IA<IO3,H=LAV<M+.YWTGO*2GPAH>*OP@*%IZ$16,-
P"L(?L@G)AWC$V)\B1V\Z+..-Y!;81_8TW"&:\O]_$U?863XW%>&OOB#XN,@TBJ'R
PVO 1M_K/^UJV'XK.T&.(BJ[W[:P' <3$+@]8)^W41R<8%94B?1-5A-^] #G=*/M0
P(_+LA/+"'=O$'BZ=4!BC54(O"ABGH,6E$)OD.3"RDWS>;HR$(5I'2FO;M<RI8@E8
P_&-C\: =Q#1*9R/'BN8.F<,,O"I2Q[]37>9J]KM(UPE-/_ZN6CL;M/(:XPLI,?&X
PAG-E0POFON$),#BQ9Y/*6D<D-^-K0DODE*U2!W/CHU[]<*8_X#8]+K[D#EL/,?DF
P[T:$SU*E8[7H"+V;J$C#L7&6W]8,Y0-]&D5=B]D 3X-BC;K'PX>2G>7_3:^Y31RC
P[7^-TQ>L$1_*6A%["#ZN,8S=3(/_*VITU$?GR&?0PG$R /F"JN 9E]OSR?/QABIP
P))KJ[%W*P>!K!49I>UCG;5WC"8%(AZV9.-.)4)2>"#4ATHKP;*QWN+GJ-0MBCB-G
PG7&1O+Q]@6%N1]61EVRHV/*5@I>S*;KQ4 !0;3:OE3!R0H=2M_P0#6R=WHR#MRS=
PO9J;'#5VE<Y7,^2S?6M-,*FT^[S=>O7OF5FJ!$FOIP;#N7_N9+*FRA &5PZ0Z,!?
P\>,?"H_RV& AG;6T**^D;0R@*1*+1KLGEZ<>7_&&A:B9+QWWE)I6H,WF+[4%W%#%
P291\ D-V_PH[W]1N)D0G'MSC+LH$@+48):5JE!.Q_K"A0J[V.@2;4%LO9=Y?9\]S
P#DIPC-*![%GNB0,&S,[/"]E)4%AUS6X3@M _8.2BY!-W\$T_REY>,%Y30&Y>?.DY
P<U7_$"GA]:P&;E^(X1^\LH-^$TQJ^F5KFJ/C_86&\E>IM:K' ?$&ME'/@0),,";0
P*+<T"P:JD-TN;&NGJ3]01":ERB6@ILMZ)"B8(B1@RH A]_)5D$EL*1F\/KDF[J'H
P IKV4[?'<SRO4E!,;/BK,N&+8T0!Z(L-MX UZ6I3ADF:W6L(Y:2T4U0J WL#0F (
PW2O "G ]#LU7CK\" _WI:3('J'$?E%^22G$@-G*1"FVA@AF%\70TBK?<U><0ZB^0
P+2I)AU+XX,.,!_/2OFZ=1+"HB(%ZQ%]8])\5CYR*%WV 5!X\B0])<Y#(_]5[4*RI
P)F=:>)C;3N??WD!S*W9K(K% LB_(XNY%H(Z^=[J83=+QFN_<PYC)^P?Q-JH4\CO:
P.*&?@Z?ZA>9(-9->[8A!XF&/O4Q]5&T+&K9B\99Y/^U>V"H^:8>?.,'F4ZMP?%6&
PP)_\+8/)B+%;IV=O*'RP;)]-=C)OFPF( X?J9Z51CA7L#*5'N"+D%\6)MR!IJY1O
PZKQ7W#"WF#M.3(D*P9TEY-V80-E(+64, 0N_1_T/N2CG-=G72G!+GY/72K/XU6 N
P--B(XESAR^J2LDK=E*;:LEG6WT PLA$=4+P<=H96"4P46G/J"%\O+,V[$P*D^1EG
PI" ?!)%',"'?VBR0E(WXF6O6('!E97P@$S,5!<S0?5Q.P_71L*:/5U%DIRCA NXQ
PYLY61!%;Q/3HSI\2&'N<9K%6Y^'T,O6%PIN8=H@T,.^VZKFG.]3CY1S6IWIG7AL8
P05N+%JIE]AP&^4<),SXB&.W+([VRZ;0;87&-D3T(9_UQ:L^]T &0?I0\D"2'O3%+
PEHV5@2N@$=<KR$XT[&]M33!R"S"(1U0$Z\KO60B??=@R.8UR16RJZ.#0'O=/ZD-G
P^TL-2J*=!6,.+],&NMQJJM?^TCLADSBC1YC@%D"_F#3!<&AZWU^LH_<93M6..'Y?
PW;KM:V0<%Q*4.%>R@E7?0WHR7$OADQ:>?(7BJ+$[=)*%JG-OH.1WND\!%B1J$",>
PR'MO+K&JI!;91D?<K$G@IP4,-S3SYJ9Y^"['%)]=^H_$2*0$J"LLO7UVMDRA9BOU
P*E/'P-U3ZI'=%"O(/=B1)> ,AI31ZA,&AO0QT!X%R:300C2E@L*<;V73F[0IE?-%
P831W,,RIV@7"\21%X\W</?R=#@6&1K[N#VYX5.[)QM#\XEW+$%M7AO%X=>8D0J--
PA#9?KWNE]"6]>)H=.Z8D$4M_U-FW"AY1%FV6I**6I-RG"6G1\18ZB.C GI-.XO-J
PN<*<@IA9CD%XFIX)7T3POQQ;O8)4/UI,Q3YC#4B>3DS<NBW0+"VP>;#H?83K7 $]
PA>/*Y\6*"=H*54YQK3CDSO?K_Z>+^'.7!+J2X=IPOIXI'Z>O(0+74-:!8AQ[V>(!
PC*>'$)18 YZQK VC"F(5/N(R++FNZ,&@TEPN&"$2_8L*Y^&P_0Z#/DA7BF(@."Q%
P"$M@(/]X(9Z'461E,;"':"(\X<;*:OXY"%WB"EOHTB$ <*]T5CUWEX**$<&NP"N/
P/F^<"5?W]OWJ&[PIW0OTW-LY8Q%>S5@C_T] @#?.OVW./[N9D]!!,N;="&*(YD'H
P_SC[!ED;2EZW+3QS]Z%S0E0\KGYI*B:;L(@J:BH>T%/I(R^%"AQ<(=_S%%D!%'VR
PW3G6\TXP8%B9.>GWGHHZ)U,'#_%=)*OXK>GRYJQS:6!)Y?6,D>8(AB)*LSR"M#B"
PEN^Q:M?50DL$X_'QR^7>>FOBLG#5V.)FO//+1HO/]FD#K=#**FLT97!9F#A-+,AO
PLB184;<^3S;/@HV!K<&Y5SE63\-=5<4XA.5%T_)J1;M'7X9ZD/>NKR3HYUBV&K$4
PX<1C_Q4L/79HDZ[,>=Z1)-NX&O-I+*F$$^0PD"40^!K^&;A#RP1PQ2 UG="/_+/_
P[[OW %V&1;9*3FO/7FS 7)K_GVY'I;9,Y\IC%>D:+U::IC6JNFH:KLA>'=:[I=O'
P>)>-X2K%0Y2WXPU8IC20,0YG+&^(D[D#A00)(Y;0T![Q\\#8;WM.W^ N&JG>HQS=
P7Y02+Y4+(8WK)A:J\O\OV^B5] ;=5AX?/ EB-<1HFL0>\6 \398)+"D?.!I%)5K-
PCF4-;!2J+)BD"0G.R*&YT)U>"%<%]9.@DKR7"Y:[9_[F#GLH#\&;JD98=-BW.?5-
PZ:+M0/^HZ@&!\Z09;R.^&OP,R0!&08Z>+2_&T?RFE4%]<9[S38R!!"+9R)83P]/<
P2-368+@,H&4<':)ZYB@.#[6X8;+AYCE$0!8,-(6U[_D[6R;R_?RQ(\I;83Z[SK>A
PH\QHH&7,XA[N+Y"-+#L_5A<8.G<:XAJP'\>M99 7N\YN[QSZ=2MMOB=_'V7#B+NQ
P',3JT5M'&Q1%'\X!^[ ^<C:%  A'DP!4S0T8@K'8<(D^)RO4#@6?R._2'ZGC&Y-P
PNTH-6_&/"!*L)47L@:8>QSTB&V4Q_(Y&+'B>]*SY+6,L,PB8-&IAV&G3/.%$Q8BA
P6)EO":(L&>TX%,O S?MV3NJDY$*,Q_:#*XX7,@9$IGLR#"NX!NUTG#U++HXG6'^$
P]R3 \)UA8YM[7^B4P(L*QJH,BT&A'R#5C(PSTX'XJ("$:K##5X?JUP:<YH#C9&O;
PF2LU4<B?2J^D?I+GW'HTY=RP>X>1VJC,A#;\= -)<8_7#>IK)$XJXC&Q6,Q4"C)D
PW3OJ^1!7;\EO%9C7RAY[K$@,PZBFZ,4BN&&W'T5K3/BT=-]!WH3SG%]7 3/9-L96
PC^AAJ(E/TG<H:4^1N0%NHXEQ"O$7A,,V^ZD(LFBK@V^M&=:)-MO"4 ?C9,(O^2-.
PZ%V2BXM1/W5ZG\M.(_ G&CTF<! 75J[>I!:3,GPNE_V'=RU6K/+6>X)!A48_T_-)
P_E'MQ%!([(K7$S2-CU)+/_=GM ^?-,GAVK9(&JZ<AHB:^,.8VY"LO=R.2=IJ0^:5
P^!,G^( 2D&!_A2CB<"1*7D6=)#]GO_629UTB^3(6 > @CWS^V\SVI#8,E0ZY^+<9
PM<^&S%X7?XJ>5 KLJ3Z-.4G!+W745<$?0O76!7\2QOD=RH)'GN4JX/HCO<(09( \
P2X:[]<NG+%:A[SI%:]-7?&63P3]AN:_]//.5\FLN66:T].V>].S%+$;2OUBB@#DI
PSNF-650@;E76JYRD[,>:1>5D&N!HA.[=T7"YYN:+CYCAWV!NDITJP,_:@2/L1D1L
P19W&&*B?=0;'_A#N6T%Z+_QX,[YN\A("%IOW(;0X]^*DU'5Z\!,^@;"+ @B&$6/X
P4Q%I=:7LUWZFRQ#>7ZG"Z'P2C,*8.1M7A6@MDZE!5O1TZZI6^OD%;6AHHFXP:Y _
P-P\E8:LQW:"<^%;Z-<MI_IY,U5[=+?!M-/KU'8Q:>Z+B\]NON^,NWG8]2'R/A^@H
P-.I9;,=7J#AJQV\H:VHS(LYPM@XNMCJECS+&<G]S:E!6TA7MKW'4+Q9]CD/$2HVN
P]B>5P\G_X>.WC]$V>5*7;\+&4EJZ"JCV$&IR2V%PCVD U<)[X$D P7.>3Z14;.'J
PN5:R4]L)S4S7--7&ZVB"5VE8I77>=?%UW]BJA%,Y^-58X\-[= $K46)?GY =&QTA
PJNQ/X!3AA"VJE^%-_"'@I$7,$R>NIW$/#A&H!@DXKX.1<76F>GL(!Y\:7;/RDA&,
PYVH>9:F37B&YNN3!5[L:::+TT/EG3Y@KYHUXH08L0^*03MWTD<.]\02%NPTS]*7"
P<5GDF*YU)STE16DO:LX>,NE*R0=F<)/4;, (><V?&,_23:KZTOL_Z=O+?9T4ZBI9
P@99@0A^LHJ=-J#/3;[UX@]]W.Z=%6WG8#J(<F-UJ?LPCSAWD'/3P)$7RNJQSCWCU
P"^V(K+H0SUXM?F:H&F5 N?["5H1'"^9,0"^9:(2):HA$IJ)8<'>& !IP3[@_=H&/
P6P/HKQBG"W__!(X!:(BS,0QDI4:4R\)7=5;@_2,R-EA%VH5/_+&$:K"HN/4]J\TJ
P7/?ND"$,=B(R3-Q;J;-6EM_.XK8E*]2)H]JO2=Z+LH6DTZ8($3\>!QS-%,-SXX!;
P_RG,T9G<!-<A_)@S9F8R:S7?=FT7_2V ';9B"T"L@;G?K*%;__4[NQ**I<?7,B" 
PKW5_][Y%!R29E0_EZ3Y,=T*6O<Z?.SQ8/("4@6F=DP MG9UXE8P:*](E<VS,6_T6
P"+2=@@C(#(!TN/$B',CS0G.8E%U5B*#Q]]T+^074@[#]K_J7,*ML+1WCSHI-"I05
PF"\4_%D8G_Z8>]ZO:C#Y/;1KY/!UJLG)0R"T%.EX@ZD(6Y!$C7,N&M30PV-JK<@D
P+>/QX"AC?G7U7\X^NXAV++.HKYY/I7)*D6F;5:YFNPYFT<6[/98FL*WLT_R5]M0R
PS/+I0ZN"YS#Q5#<W BGAJ\L:D/LIYO*60B$B-_UFD,JI'/-WCF80IGE]_S$[((J9
PT^T#X=JA&2PZ;808UP*C>!R7T [E 'M+DKF"2KYQ2P8:E@0S>A7OS*#M!:);7ASQ
P%D#2*?55:C/2;*ZY*[*2L9C/'6[<<<?,EEYKL)@9"+:FU;*9< T5GU<F!#MOW9_Y
P';T%DH+*4U&[9=N<G ;W2AUNHKN5B$]T*[0'K20M;Z_[%9:UU9K.GH@^OA#>"#,Y
PG7F1N1Q.+%%S"N&N\G'=JG@<V/,*SP5"E6;]5RDASPS13IP[<GN&84DTJ3CT5X85
P3=PF,#^<JC@;[KWBZP0/WCUHL7:U8RGG+FZWI_G5D01\$'-QGY0@E/$O.43)1MRV
PYR"'JP0PY<M>ENYLTID.V5._#YFT)58)W>13\8D/K5&_A(6V\BFI/3/,Y]AUC$LT
PU#F'4KQ*Z@%Q=I![LZ7A!"^]#(&,*#C%0$5:>IEJHHHNOBV%KF)"6)%KQPXHL0[4
PR;;BD$&3RFCL'\E>M$,[GE%A@ F!1$[]3>P%)*S;-(M[/\(]I%N2%E\WL)*6!]LT
P9N)0L1CL-^U]<+T1J3_!$:!QK.6\%M\#U:,.M>W),A6&D4$F_7K<Q&QW]LI%7JP^
PX]@\88\, \'(.!X4VNA</=81:LO&;_2&$$D@TIFJ *J^0E6UFAWD/3?-T)H:*770
P X$ "HOS1+KJJ?C3F6]5B"U1K-M?)IWIM:4X(.K<F3//YH>ETI9A/UHK\_O8?9O[
PJCW/?FU8/S >J,(!U 1";VX;6W.!YIW.:*TP7WCO%A6(C#),)1U&XD,&)OCOT!MO
P1>8BX/:2Y^:LU6&J\4*JVSM%\H!0B@ .!%V=..=0.$82$'6P> 2HH<$T\1?ND%10
PR;0")SO =>%C4.. _)YV%YS(I?%T\D:+CG@Q]@/?RCPW[ ./"<ZN6JTM9J.!=T3:
PF\5'&\71BZ:5=!V,%,$?9M +G<1)HAIG A;)DB]7XBNI"=TZ:88Z7(D2*7O]PDN>
PAS)")0;&DPZ%7-G8L[$+S73WX@:(W''O3-F_#S-=3U6,OS,OK8G&X5\X2LG4F]D:
PNP8CC0J*GU)?^>W);@C#L,*:I5+7?RO%PZ!CK::W0E<NM+EE\S^\.)04XU@+-#Z&
P*+C!!WNNB[I8,;^YO_Q,"$P/2<AT<YPB]= '"9X)% $,[RK/BX++4;YY%TW$.I+I
PLQ2 _'83*!LJ748O7.KAS=_K43!V5!+@9M*%O$#8 Y:I?+*51R7;@9(CR),?R7+H
P9KU=.0(DUA0Y&LTACCZT)'_/:G\0X<,9[LCV[G2?S,S74K3O@E$'L]IA"'@5HQ^C
P_9\,(,Q7PL7JY";.45%#!.S@Y<#P25D]$YVN(GEGR$?PC[ 6ZBTD26OEBHZ!"7A>
PU"LE6]S^%AL2@*IQ@$3(*1#7<(AO,PE=_*>NO%'L#.U[84H%Q?'= Z&T(YQK!,5W
PN24G,8%NR,H\42-LM%WLC<_T8<")5V3#$SS\"3V;H!1,X/IYBD+4NH4&*.3_@/C5
P&S_ KO5A6%JA(%8/(+<OQ!H( "[[J-2]_;$9VMB4PLND R[G)81VH9IH:LXC@F7$
P[U/N?4J2 WG(I3T:_L+2K,KY?1]"_2^ '^Y55<(+I&NRF^0FWL"*ZS^(<S_B;DWV
P6Y(E&N9Y0.,S/,%,U\;&>MN_-];TAJ ZB"7QN K?^$L58V]T I/3N98KA#]: E'+
PA$=Y)=;F].TJ2X:VY69((UXPP3,Z+&\HA;Q(*,D?P>6AAPG*:+]TP$S.&+ 4S6SM
PY1[P=,\SJM,,<8]&75+&&2O! L-?\Y,830Y\/A3K42T[7)MI CU8/MZ"2SY#.GAY
PN:7"YGD!\1E-+*C(--9&!5TFA#=V7'#OP$BFHH\/UZ/?1\-?C\R(T=S(C0^O?:D$
P>@C/-I*:(PVXSN984AP6RO):*3^*G+7O+Z=;KCM_Z$/YI89HY$CN8M0#D%Y*QB<=
P]Q-'028GY9.2Z9_S:T5/=G?(R#!;/%X^(Q12\#&@[V::$E$[QG8]7/KHS_K.!#RV
P(E!4<SN)E(>FZSH;^ 1W ZSJL@NP9+MG#]164RB4GDY4<>QX3BW*Y3AGC?X^60KV
PO$GQ+8TA"?-X'=$!UMNSKFS$T&]0TT(]PVBRC*65_LHX[<QIJXB/;D-[T,])HH[J
PENJLUS^S5^\:A%CSE[48_A5'7*9ZS2>&H#JAI,]<=94AN8L$>@7MA!2/O((F]H39
P:E3UM_A.?&O&;9PR,?:G3"OTK@Z33;;12]_6+G#N>#?BOD-\/OR=S7;N\+E%I-^W
P*$6H'6$?0+"R8=4CR,(R>0WJR!;XL!IB-?OI1.#(5%3#FY [_#%-E5WS[NN"TF[0
PJ'5L05EE(*:Z0[;$$7!GPLMT!=:Z@-KCX.21 4:("=DQ?R.2;*)2=]U45)]J.7=O
P(;N7E&8]X=@5& :*ROAK*AG9#Y:WL!H.TX"R^4W)7@_2E3OLYY.0KJB.,+2+A,AO
PKAIFEM;'$,$I0]T2']%_B9E/W1L)+P53F=],WNV8CN1^U\FMR7<%:YOV.T(J7FX_
P;?G_@N!<Z:,#!=H>$@]3BO"GRT$.#0(Y4^?3 3T,+R7Z@<X7RMIJ2:G3:$P0@9B0
P_?V@+I/.^A=/P6BY+TIW,MXJBLU..I"?Y!\2@^/O#E0@W3/R5!:)[C>,7VD"%WSJ
PQ;<>EML=H6,-VI9)' %]OKV6&NA^-&V1X0==4BOX<?C?QR=ZNO;N@**ADID[6KG5
PI^BW'GB47%M15@T)'0B:4V&3AQA#95A3#+HF^>[GHM7^6;-8X]&G3->WA1/.@J1*
P\"&DPQBTW,PO,!'TBA11'$4>@B=GGP2WE^_'34_>&[:% 64V5G:)Z*GCWN-+A?Q[
P4DJB-B8Q79U;2A5R 8R&+ $4!'&<('.@ ",S)&T,XW]$X>[SOK"(!B.IAD96/'2_
P:(!#P\1Z]OO$(CDOJ/#\M]L%^RT6JNZ?G."Z=439=)YA'D?I-)]FB\EGZY#K[WOL
PNBO9 -,M<>@X\R\%>LMM64",QX4.O_T<H]U@'L\MUE"%?RR6+44TL(BWY"@G"V$H
P',HUCJ5K*CN@302 Y\ 32A!)R@<'2#3$PJ 5:7KB"F)G$JPG6$06"_;O9?E#9=HX
PP)"D,Q\&ZE2FYO0PL]DU[KUS8\C0-J@VF_Y.\ZK6P:4+BD:&3Q<MHOP>@&Q?T<NC
PEH9V_.341 '?F+DU( -IH<)$O.L$-8_D*:@@5R)(L1U?J@&V>'<87E:<D13EO^%^
P0AM"L]?)5?!\_A>>\9NY+^7@[]"O ]--\\5.W]9I;&!U;=ETJIPK4.=9!_Q_-!\\
P$L=V\3U+_P4BV;X)AUTCQ=/YIB!#P#C!?F,S<315 *R7>4 M35E KB&C.55L6;<6
P/;(?%7UD2HMH;$%.@.@#F]S9#9./.<ZET?J[/6P%!YR_7C.$J"_SWV_^7#^AXS+6
PYL1VZ $SQXUF)3HC]($LD=Z\61'<-DTF;8QE20J@?%+ >MH_=@%\!!"B5O 6!2OM
P%4"->!F9.O?5$<K56!#_0ZA*UCS""F8=DE,=-6ZU7"G]P0H8#BGJQZ^%AN'1#,\!
P[<[=)13'O(>0QON1*(^EV%XE8C;[[W'A@'5CM^C.*B28G1G[#<6%QO2J7O8V8U#G
P73 ?"C$/=*RJ N40FHP**A@*CPD=CO=;DDW:!L?XUH16H(5H=%$SG.ZS;9>>2]!9
PU)\CBS&!?%*@$JV6\]1L$Z7ZH"M1N<PQ7!&:23]AF''8,0\K2S"YK,E]YB4ECH'U
PN-57 OL,AJU#'$F" X2S><E36!&B 8IR_03:3UX\7#$:MO2%\K1Y,)^<1;WMZ35;
PY0%(XMSKIL;:T%R4]'E-9?%O%#ZE&43C)N5:8")G2MQ+<13NIKZE93WS),; FC-U
P*9V""')F^Y*.4Z\%[.WV>X4C#$\OW\RLMEG5EX 9H#DCB&8-6\/"8BJR!PDO[6P7
PKOYW.!C4R[/7I/JO'-[B*3SU?JX:96'.USU1ACHW]"*AB.>] OZ?AS8#W'PC8/LG
P[?^S(+/ZHAA'!J\*7BV65.P5='RR10/"XI[%MET+6\[&G3 $"X*D09.W9T<>8'G@
P\!A[J$KG<$2!88 QY%RIDN@7P?C@!Y$![9D @(HF+'9KNMWX,\?!C23H2(<< 9S.
P]' 8&PP$LJEQ.A+,R@)L/["'&)^\6-:@Q-A&6O<8481+S1]W]1"KV0XSR0=(Y  H
P"X[:<ZEJ,'#MKB";P$SZ['!IOA@J,UI6Y"*#)><2CV'@9%4"@&N@Y,SE\83'1FPF
P,W\F:I0D0RUR5@TWQO>*"$VH!%+K,0%O(?)OSW;^,B?'$)=H9\QW^+6"P\@LXIE2
PB(;DBT4)9=J0C(1/:@\:GU)AE[Q,WQ> NF)NN6<>)#DGU3B,3,$8Y9MMRY0.KIKP
PZ_QB=W.S"@@#S$C@PI&Z;<$2<5M2.[_4D#A5>:IW!'U66=@VN[8K#=-H4BA6[^$E
P0QM[*.$ROWE0K# _Y=H>.X02B42$P4^.3OUL+8%3SD3ZAC'Z);?Z\>2&2I98VFA 
P2HTX%7%^GC$Z4_=.")A1H9!=TMO:K.U7S:<X09-YB[]K#.D-32(!.7^XT])/U&O8
P9B>EWTS/;<NPR6G)VEZ98!L.^C9G,@NBX>-U)K]-%1<5?('__RMC6US:RC,1\E+O
PS,N4_WYO"]9#VW(BO3Z=U8.Y-H"38B=2_09<^\:'-_+-W9R+'Y!ZD'ES?KFC)H\8
PQOC69@G+E;"0\GP#[YKLRQ\X_ B^D\3XFPP+*_+T8OV<!N/2K 2+,Q_OA%$<#@*?
P"V?PG<'$#P:?R^[?L_[8DN\0O;@-?XH;?H$V=L5SGT]@#(\&/K,V#"JF*R2609@=
PY/-0H.Z:#IML$3I]'.T/C"U?E<H2L/<7;O)4*Y"4DF9M "GZ5 ;,0Y@20'(AD7&S
P3NJK,<8]VCI_HDO9)$!BBJWAK6&+@M%A^2R#4A1;=U()]XT8M&I)R[6!_XLS9]=]
PM\O4=)A5QKPHM"@PAR%@(PXPQ>L1J(B4?Z\-/J@+?MGX[?Z'#>7F9I# O)"[H217
P:@_7'IA;%GAN '9%1FDU*%WEMK+-<(8@W-RW/ A+PYYHI PZ</X]B(5B+'"0(&ZW
PK?>R%*776.D$^J6^0'OXU\DX?Y6^T2IP_<J>5XHFR&\XMN!,A=X$_DPC-%TMA :A
PX/1BV1]JAN]RG#^;7A%I-EAJ[&^Y"M,TS3JB;64*[BIY_(E>@6UX%Z5KLWA]]3,&
PEE/^K5P /FWU9\..&BK3C?/:GS)S+UXD!+\1\V5+J_6^YL!M^^F1X"@,C-BB!R(<
P6IO56^9O(2'^L8-/C%2R6Q)GGGK9L%D!;@%#C$7 >3"D5^O[;:I*L#IY#$R&? @_
P/ 6E?7JXF &"-;?+OK%(O#NT]2!_*E7"FF9%_*1>>:Z+)U,%6?CZ  Y%_-R@.UI:
P*WR_49F<'>Q@[(7@M:V\Q&T"<\6'HV54$CEAP_Q4J:4-]54F31&+3Y](J[[F8M1U
P'^ *Q64@T 0@8YTG1V4.#RG(C(#VZ1XGBJD4U68*IW*4XB;F)L9BEM5\]'>#-D6*
PF)D/$U4XM$ZXH"]<D6FQ\Z[L0TC-HFZ7!J^>E#RZ<@GQE,5P:I.$Y/1Z1TUQR>'"
P_S@.Q4W:@ 'IVLSDM+K$71CCW)DTO] PV %0KL?\@^V"Z\*E [-0:1.X$(/&!C%%
P>'9+2 3)(=&"@+8C7_8AL'&S"S#4!)';OK@$(P_8*KPC>QRZ>;IXD\ #AZ.2<C>)
PE?@H8., &.A!Q.W&V,L?21.G%Y9WEL%J"R[FVI1W0Y8=9[1S/P& \9'/40%RO&W6
P?I%:W0?_<*T)75B+0F8X-6,BUHQRMOD#EY9";N$K&3<EMX\+(/K&D%A(#)J@/M4(
PJ$%NRJG@>S;\;YS=]L)_^-C2')#P<4/)^D3A;R-I4GNDAOBI(R6UIVM.F0C""ZW[
P8N-#BM(:)[UUBWAG8!(0]7MO4-F@!7Y2\QVX05JB*NZ,4&OEN?]Z@5JWJOT3;#=:
P2Z51W@T7R!E]'G-,Z2I"I6P)2FLQ7+/@3"X"3_1?YT> (V9*233HW+U@K21<09A_
P1P8O,BJCVL).*=/DX@;%$,W*;?E'<R7>FVI[+5ZTAY^O=!@F8P'6/"L"E1Y+AM13
P"LY1(F'HA9HR NWQV1]78N)U'D=;O 8"H*-*/?,])/N6]7)G3S-][EOR'BP.82T4
PSKY7'!%LOA#-)*NMK5:,"2,-FC+)ID6OYI8Y'OLA)%;[]YE;4J/*$L:<[0G3Q<*I
P/8AD!&M->R>4@9):)@IUM6*HYI0;P2F_@+=@5&33D3@%)%C4C3Y;W#>:HA1WW=+8
P4]$A+8.C]QEJFK0LE%Z+I7)XV7>\4GI2ZME[?ZYS\&S,_*D&M,I$G3>_+A 80J7F
P0TXRB%\*;A3HV_LZ?H:N#P&9=9 =2NG1CG0@"HEOZ +\#N1H TL*4^_>:E;U_JM>
PFXQ%*S).Q81W^AZJ8(MEI&._7[J;&"+;DH$)_?F$V@B?<4%LL\4Q$7O&WMM&CT[>
PV$<2^NQ3;AKIWR@8V+M)XU[IOQ?8B]#GVO#&!6 GQ[6R!K2.,U<;R]&&\8^+\<,5
PYJUU?6YA6.1MBA3N,EES$]E>4+NEZL^6"".E/=5PF48Y0MN9U=L9#HLGOL';%&IV
PPO2+^:X6\36KVGNP$2V!S+I0MN)I_;M)B2*7GJT%4-[D_BWF\/WDINZ*&R;Z65GD
P0!@U)4Q9.T9?$_A],;_%Y:0A=%/K1T/FQ\S#]'T<DPE$<@W^()DW%:P!7/S"[AIN
P93SGHD1Q:#W9,B2J:KF5LN%QAJ=\@5(WPN\IUYZY6W ";*)LG7O)=<Y@J?YP5>D6
PH$P:&"N1T[,*%[]Z1DAB@ZWIS@0?]N  8@72 ,VP!OZ](^$SYHKUQ%>ZKR@WD2?<
PS+R]N&W$KTA=FK+9<BF1?W;9F!BJ#A)T";@)B *!>S]PRG#*%)$K2D#O]#+G.P\+
PGS&F,A0.!NHXWQU4)3*<@7:QLQ29)5M?\CA2#,LO#^I5TKN;%9K(V,<$+!\6XKYK
PV#!&SA-"J&YER6J. (.^&F:D +EBUL_#:U*XPUU=VY,/K0,V9XLN-=?4FI.;65>.
P''J"C&ZY P/W84@?3);E@V,J'S6-<ROX*\=26\H(K90!0(#T+UNA!<7ND,]?%.QZ
P%*/]48DRT2XI5TPA&PC-)REV.>C3B@U]L]"">42D-PS$8OID68]H@KTOREJR8[=[
PU,J):,8SU"&9$)T01TBGQ?V/II5U7B](*?M/74U7@+FRH<B69@TVAIA;=4MD!$']
P>,!TBE9;8\2&H4QFK("D9U^W*!A-KI4MQ5P2W@MPM>M2/-[["6(R33CY??/T<7RG
P:31P,#R=0R4?:^R\.K=XU(NYT?FB%85DVO>5X\+:BS9SXUX'.NU"L"4#6'1-E1B[
P4.).E":RE+3;%-TLYL8.(D[^"!7$JK(M3P-)\WQ(13CXD@T(\;"(ZU*(0B^S8F1&
PCR679G-:5EO$SHC#MJK9A6ED*O'< V4O,FZ!3MV<#L*7_<9'\K'X1<NC^V"J4ZR]
POU6_($W\J/U"B6RD1 -2.%G O.EP4.1AH/FD6[/\X-VGX-E8>#E'$O7UQ1)@6MTM
P>_LM@*P)ZQ"_3<8JF+[B>A) _?CS=[Q(B,$&4(HP8EB<D( R1HQ'SPZE0=/E0=-E
P_@^XM5')_GYV19.F"P"L^2:,AR@ PU<SR-8RH  <%K+6.#\8O6Y"<3=&4#0K4Q_>
PQM5&M[I+!+Q8&S4[VK,GOPV"N=RYE*A$,&-U:43VPI%2L;I)X14[KLR])4$D**3B
PJ]R'S[ES)Q?MI-B8XYV@*Z)B,"$MG0ZM;OGBS%VN0>,04Z+()?ONT:-#]]O?%MT^
PA;>8855:J3CUV\SH_!6V<\\#AVE81N ^S%6YPJKLKO(N1S,R'G'?KP?E[12>D^F_
PAZ\&,16P6NC@:R)/-C]FT3?GK7;3)L+$-TM'Z@+.VSA2M $=/IDLF8 AT669*3U?
P^PP+OU9MO2J#Q;_;](-UL*L3Q;,[R/;XZ&H5=(:<TO;FU?S*9,/)[W(^YL1&W;!;
PZKQ<#.?+E9]R0C03.CZ>2( V<MYLO@*[+$ BX VB;6O [G-(<4%++*69_BL*&,X-
P@N#,EY!TV%[%UU9^6*<PGD(3*THY+?DU[XSYL:H@2&((SRQV<QH19N'EHS"$I3TC
P#[=+%&<\SW*K6-066*XP[T4WP+/$G$Y" ;OO/C!"[!?%+*O%9NQ2<'%]^3]")0*5
P]CIV;ELG3LY'-BGZTJ*[7J?(!41&,'),[/R6!*MVP#34=GJFW4<AY<Z)F^_@4OWV
P ^Q0DR\=I4ZYK+! I=W[K1.!9\]756,_ T2BAMXK%G/:"DA]N(=;1!_A1#F=IJ;5
PI2WV:T\<E;64@@MRRQ O*9%&9P-,PPT7J+_&ME+VEH)$B8(6L\N\?OV8G7IQ@X7E
PRF>>T]1P6JAI\T&VNJ1OTY;B%XL NPTK=G*VRV#> 6:7(J,VW6CX9?V5GKT[2<3:
P8QA-+$\SA"MR2.7=P-%:!N0'& (=0?@45S].+ND?B2+0X@Z<4^/"UI/YKRS>J'V3
P-1?9=<-3R'2G6T7<9\M,#)RIZXP?@RWGA"R^I.&L9/%JX%* /FHQ:K6WLL?X&DA 
P%K-*1$/BZ<+Q[_H<!*SOU6+(J1Y;8XV#_M;QSS1C#J+A(JM75/T(,<M?.=3OHOK;
P;LX'1[*O"4J'-B^Z=)VVJ2\.&\+N[C?1I_;<8.[[B77=0'$%77\Y, PIY7E6.FS1
PN0QDV03?'/U_]<'#HVJ 9B6TXX3QER0A&@@Y[5*X'ZU&2>>2FC6@Q)FA(+KI6*;$
P(BL0'1XNQD)BHUL(V>@@BP#'5ZO.2+-LR%CAH1<[4RITF-PP>M#+)3,82'Q15Q*_
P.<&P(HD9PI]?S"@GD*VU9K#&SXCIH@=89JIRT]$&'W-<;AF5CK9R!3:&.\\"$_Z<
P7;L7U'+N^*9,/'UJCU6"3-O@4A%!ED]B3R%DZ]+*V2I6$5D"(DB6.R?6]QY2U$Y7
P#1BGUI#HGAR[..;3N7U"M?&!K4-IAE6CQTDW(H?R5@X_AC&*.H^C])BH\E4U&JRK
P:MT7D"D9!I)C!.,7RQ 0&0LVM4\H3"L H^1?\.-2^G< %,.YQJGV]@?T6I6$"F(2
PBNJBZ&I#])YAETZ_$Q_J<D_R8:J"&BNNUEC8_987Q4DI<O!0QV;U\)Z8H.HXW"5[
PK0 ":D8$5H%B@$V+DE-'O.^Z!1FS>L(M67A5Z/]DP=1$G#($!,2LG@P!'2FP-V\E
P=$FPLO@/L'^"M*(0*OL(!F1 0&MMWNK^R.-TKB_(:26$_M^:\EW']H)=Y)'!PP1Y
P/'XK)Y$/HOBC.FVZ__9Y$HBNB]$T1>5L=:_R@>H/+&>Q03A&_\CRM)>;;OOG:7D5
P L>Z,M1:I\1,';.5ZJ77>ZHKHH_K<2U_CI3<XY?N9UGCO^N=._ 2U:V>P+:F^N.$
PFKN^A!31/1*474*\X\'N!W3+M?LNYR:TP3$3085PE,H@"2$KBFO)-#/@ZI5A2^BC
PU4:K/GM@:[+YO_$*RD)".]2DXJ'="=OWK@;:ER89PG+KY]*/,^:=<&I4'#1_TZRB
PLW[ "D'T/P_]9:S.5;'Q-R@/7>  U!AV]N$$ \\';DH)ZK_' 12U/4[&CE(VZ)HJ
PNHBDL+'W="5 NJM[#SB<#@;3HF\ +L85 7OO*VCV:.(^!*Y.VHVBI^,;U%3&+#SL
PL0UNVL9BH4Z#/5.RVXR'+7]CBPG?>H[IL(>^ANEP<OZ]R,X\95VDQ82;8^E8$RC*
P8!FC"=*4TEIX_4\4>3-HIR*3_*.[^'#K(]X([RP:94YC=5VHY'! \U$NM!0UB8[.
PP$A 32H#'F7NJIL3H(M2WR&>RHA=99T+/UF-OL!H<[Y%/$9,D(!D<Z52MW;4G0:)
PN/GJ+#L0$M3C(KS.<<%V<,*Z^J/13:.TP\OK'R^T,Q*'V:H,RA_UZ7W'OXQ6QU"V
PEOS)C#U^,47N[B"NP(%OG^DY_=-#%ZVL7N9<#A^FSR(8]7ENVRL -=\7/Q/TX[Y$
P]UO.[U2*:'\W::#G:[BRR1'AYI9&LSD*6AT5]6X%,+A^BDPTVG,C9:Y3@\D%S")*
P"%/L!A\94;Y5#Z5\=(O^U[T^C+3L"O%U@QM*I1LG:9I-4'*NC-R.,^8-#)#))GK[
P;F()^7[15KG/.V8=DN55CZ)F]*7X,EPV[$OT(00EF_%8(&HTHJNT>?2<RQ*!RI% 
P.H>&]'[)QM6D;KFI*?OTWMWBQ$&+;WM[AN]>6C"8!]D5Y04:&G:^DE9++8.,.=L 
PQ@E:H.5<,CE&>R4Z'V9T75*DW%"*'!DU2_3=>>D@TA\N,E/>.=HX9&_1SE')P4WQ
P3Y#$C86=:I\3.VK+!*]5:IK:V,QV^.X\*D"F3HY:UX3\WS<^*A@8>>$ SZ2C?N+T
P]%@G2+)-#N HU0."BBJCW-DT6^.?T?#;@?7+HV> SNA<+XBUB=^S?C\L!V&3=@;^
PF[&L8/X"[?9I55;\D6(\$ZCZ1'3D_[ V E(Q2)>Q;[W JO(=)*,EJA>7^3%1V1 R
PU'P33O?;VN'4>*'Y9]73>C5<-D'(=@!OFV09SH')4J;V^]_YJ^&*P\ZF;!E,9)7&
P 4? 3[SO#&X!+#90,:1XWOM*T@!/'IX@<]HBOKIDSOJBE8I>@JZ\.NN2\Q2JPKM 
PY^>W>9UL=3G*6L7SN1!<E^8 F2'H6C():>#VZ7D*E$1!ULWC/IROK)[#^9;W/UA.
P]LL;Y-QS$"/C,RDXN=_=LS[;GJ8:.K?\>*?4E<.;/ZS7/JCAQL+3)0Z;DPL00:5(
P]YA (TP0@*3I6656"J0"G4J[&E[9>0A@VVTT2PMM6J&95M3I"FH#.$RAI@*7+=/,
P"6V!3/,5=[G@=B5)E7AT>]^D@"9Z]^Q6>8NY6(54&4]<3 O8S-^@:%JAB!EO58FV
P1Z*@IER/_/'*#23N<!]_[]>8#!F2\/HBQPB:LT%',>@W3 @^0I>-#]@'[S@_89:<
P^!PZ=N@+ZS;>R<GV%YGK3X'MQ-8Q!&00P,@@'W'B<1\\S P0L/B3VV/@/?S7Z/%0
PC_OQ]].2RK"(C?KU1!;JV25"$@&7TT(F603*=FC9##Q31"+VZMMHC=UJ]!>*21TB
PD"XT-?,K3Y$#8% !4DP!(O>US&A]E@_;AN_OR=:YY^G?J3<;D1_#Y-4"T6>XK!#_
P2Z<+5P&_-P)$MV7\6CI*;/[U:NT LF\0(AE_J05\]R*L,G*H1V=F-+>;?$IIKGVS
P2&J1^NG@ M0X3APF%>1GSG19Y;KF7"04H42GA-BSX)GJ1T1P0MX'UT/.\+Z32.45
PD/T8HK=&Q3DZ]+#^7X^5RY7,^C&P6P;'T*10K]+#2W'_\/VOEPI-XLL:#=T*+/;T
P9UY"J3HB76L:%B%EP%BY=3A9F0U0"**^H#RN.#"(HSQSSOAO=,?\+$]2 J<N-6!_
P9&!3D8YQ'6CX6S7FW.!^?.(30A@/(_F[.%+TL3Y: /;KU)NUDAX$4=7_KK %R>\4
PNV1\&EA>(O&=;;+A)(8#I( 3LPS_OQ'][ ?B?>G2V1>T64AS5DE9 %DDSG.J$,)S
P #]]+<>Q)UJ&KN[9Q<OJ6U M8QZZ<O02;].REY1F(#!FZ4;!?ZH%\A>1WS3OKF&@
PW8$O7,,D7*65+Q0P<&=LOU&V!=KL%TXZIO+Z7E?X3(N?G\\> E2;.;?Z8<7WO'W8
PEBRBV<J&=[\,>].;_3<SW(:$/8GUQF&V.$SQ%E[:LIWN:I7408:HSA9VX7ZA,56L
PZ(='14O0J";&375,"LS@-U%EK\A=<FM]Y5'Q!,2^C)M/MLE%[YKD]0R34'C@M(#;
PF8E)G8<OC(=FB5Y1K!Z-.1YSZ'X-LC\M["AUH>&@)T%KB()&+[?Q>_.]\+S,!?M_
PVXMQ^7'-UT%O)H%T,]V+A,UT;@5M5C6<;'52PD1&R<N9LVL3-P(B^P%6O6-QI'TE
P+R<O<P=8HT[]**5HAP?WW"+T48("7.49_Q$N2^L,,[=5&K&;THLVMJH_*R+<7+@G
PE="&5-JDSTJ^3U$3G-N;>8.)?^E&.<<#"P=1#B9%4X"U ^Z#S^G2L=-T++--SIJN
PL15)VE31F T:N4G*D,M+@%GQN/ M*=\@8!&RE#X;D$6FMYITI#1 A-1"[-GO]Z\)
PPPU+_(87]U+1W'/^Z %(Z#D^U5^#]6F'-B6+1''JH2?BP@1BTD&4<SEIG)ER@\9+
P&6 ZGH39U#2@3%+&9\U9^K06!::B%JKZ/P%+0-^T,[B5)#IH :^I5L&<&6>\H5O2
P4\?1J!R3PJW:BZ)5/DG9,;"6XH47GJW(DL>H-K]&=#LK)CGN5'PLM.(0CBS3YX/3
PXO4B4DC$TUSM3_ZY-,X;W1RXU&_M"SH #7RX4<DQG]-;;A^OH('G^^FLOKAU60WN
PSYAR(G;5+XU2Y42III49 DO:KT(WQ::ES?6+O"7EDT!!RI&"$T>WI>@"8T[[PPFL
P9@?Y(5ONFGSGAR*/]-K X34+2B"9G)HERB?X2F3F,PMP*(*8 /C&M!5M*1;=(!6.
PHL0X!ZF]1;I3C)3"W%35P?#TI-"U,0;4%4(="Z)6*-Q;:Z,NUSB<ZT];5H/9DYY)
PTYAR.X+/5*6 ?TP.>0XVKXX4(FUO[#C-?3'WBUI=WY#)@2,M:_(DS]Y_4;/&-U30
P0&#T<@SY+A-!">(T9]]ABUKJ4\X72=^;D!.ZC]XIN'D@J_,7^E'YO7GM,UAZYFTW
P*W!+7<3N\#XXB)<8;AX;+3&V%O+'3[!9P$QL-&V3L01QP.4EC=,PV@9H5W+V\>)I
P4D#KJM#UQBSU #_E?2,&)'_W:/'\0EC71\O>LWP!.]>*RY8VIIM[?0?>V1$;@!)$
P"D$03S:P['@&#,"/70]@.M7#VA#!55[(#CWJ-4CE5M$;(;V=JNGO(M8'=N8<ANQ)
P3KV]?EP&ZFA#54+&F>[V::TH\MHX>5?>5K640Q7$DDNJVI#^HZR##DAI^#+#VWBM
PSBZZ>8@*G%;'*/>I=0",2L+4<*L4'TEL64$-QBKH8CO =J^'AA*6<?\W=F=!$AS]
P@"(OTH)LG0"$^;U\\>.-!K[N'TGDOCMJN!V%1P*;+K9;4PT9G3_FJ"#GE,B/@4.;
PMSB WK+%0Z4HYZ<+K,1^)6M?6>&D*6GC>8(X\B#X;YWN2(B95NSRD/"C",D[ -SY
P9OL5:D-\_M()A%YA(DV8Z6.]PST6*E"?<N /UZ/B?_!>!SP4K?G<ITS$XA>RW3D+
P'C>%L'^%7,[L"QO,.V$)CTX\O<@!ZFA7YS!9R2<#G&0ZP<5SL(97R![9CHM/ZZR5
P3%30$!PV9(B3F_ 3[C@5)]7Q,:E9(Q%9()XKG1/OM?E_%1:9_7'>5ZN]$<-^]KNM
P])%B<:I4HRZ&'3<EIF @@&CJA#U=MW6=4VZR X5O_+2V'NAQ+W]'O:K.'OA"?G'7
P&@ 4P,]#II"HMK_';RY/UTU*>F*?$^F0S56 Y)H&2BJ][%;20_O,J*EGHDJJ0$6%
PY+P'CO&R[=H(3S%:N>_%D="]7T3A),O\FQ5[% _,TGN;/NY3Q1O33YSJH:\$")B^
P/V6H=1$<C8SB8I;H+L"R&G=+^A9LJ/?7SM%X1&A.F(DG#]9F6[PJESJK*X@%1O^S
PR2%M ]W5>D:I6SLH_7WI)S070%+FT_'^S\W%0:CZ,#7K$<^%'T5TS&9MU/;,2K1G
PG)X^K6*_X)5<=.J-FWEM(RFL4&='SSMP7G!Z#=5F!QP RN4]M("T;=MN!6:-W+E;
PZCKT-(*-%CI.7;5#CW@+"6I2W:A(K-6#[ ^LU"[B<\+YKQHNP8V)&K>A YL"'0JY
P#_?"6M"HW22(^=1"4AQH'DP0K;:W-0C8UGL%!5[PW&,H:[+DJ'MGZ\.14]$[\C(C
P3FP,;(^8_%H=PV+5WG>8RA!,K(^OSXF$O6R+DKHF:29H+W1YOP^2T\@MK9U.99]T
P7@H\QL-GMC)@J0WZ[X.#Z:K1BH^+J,O'01M%VK,$IF;81-W>IEFZ9[MY[^C4NIFJ
PLWHRN_ "/'1YWC4<YJ$/=8"16^.>?'DMFQT0C#G5&^J9@S1"Z$4R_G"7Q<%0+HET
P]A*N;& I!.&-EX##)2I),XJ[C:>UEUCD!>2Y6H)7GP5H<+?.(FP41Q=CLM5S!9"1
PZS!DE1\2;SL5%U?S(7;X9AH-BBUWAM#T4P%H^_.E3"UD#MC52\#XEDC%6H%[H^F7
P<'QHD<L\)/YU*-M<F!>HR*R^%"[)ND),;[$.9N\( Z4E%J+#"83!++J%*"IKZ.9G
PXQL5]Z,S6>11G1R'H:)-X-+6!=T +02!135"@8SP"@(-PG0L)VHBR?%S4.>"<=[-
PE%EII/S-\N7SH.]^M'\5[2$<?^^W>E,'W%4,-?DR:"!6S=M*G<'[-:_P_7MYZ?4#
P5_[;N"=6?SN.IBFQNZ\_R3[>TE\^0U+@EI_0J.O%>'.@._P5^Q>GO8 0%/YSIO,U
P)AG(+FXV2HG.;I^BU,J>^CQXT(]7X,:2<PZ!?A0!?T3&I]9QU_ML-P$QC8&W9^G:
PT[74=O'758O#DE+[+HJ<Q9Q]9<ID]-WE&S/4@261?D+:EV&YUSRU$U1G!5[<=F1F
P]]Q?]Y3^$9F3;:')14,)^P4>.O9( FQ=:3VVX4E5 *SI=\]IF5D!+EA2P0L0FTSP
P_$T8,^"P3%FW-U2380(9#?+.4-2@:LC]RPX793'NTC# >D'26X_L,;1DD37LODDI
PTV@%2?7!T7U6*,-HD:ZBQ1]&##BX]799 @A'TUO T]KWF<Y*DN0%3J>@WVIZC-_=
PSN0B*4+X"CN>PU\:@Z.7,5.E&]=D=X?*?VGV$LWM<5;T\D?_N/;5*G:9%QZ"A/\E
PB9L3?/OO7TVOLWOA/*(?P *F?RV^97=,H@+Q/ I(!'LA6\[<2RS.?!]WX=28YE@.
P@6&'UW,LP _/QC(4O;O<LT+5FN<VRU "#\.A&O)QGZJ)N(>CV+ S:U:)G="@F.0<
PH<AP%%@C$Q6IQMK-1)(A[?Q,QN""PVCEE:,0>.,V=Q2D_P?^$^#5_T!,MZ#9;IOK
PEQ:E'MD)Q+[8J!A#D9X/ =_^D0SE.DF!*_I\?D P/%5/(M2*^/^[H[/80Q2Y6W4#
PJB!M@GK3&T1*!Y1*!2_::N@F<[3NJ#-(^E']M&18@&6+>G)8.Y3N)8NU'E<M@;2W
P*U]]9&JF&/_^'@4+/_2S=*&4S_I1&IRR]OI=Z\\(_<K,> #YTV9B$+:BQ>C""IA)
P<<H\]X!5*FRM:?"5W2UO#3_PTZY!&M?SOY1[U&9N0JJ<:EP2<[W>$SI2CT42:E*;
PFM5 8>:HR'QP)=>(#1)$H<U;=;Z3EH[M3\4Z>7<2M<Y>MZ-7;;N8F!/#5<Q^-$]O
P+RX^U50\4Y:)D(9HO&XB0JT\;C+TG_+]*Y?MIN;6T/?,P;G.!.X"'-D-0W&8C]U%
PK@BQ>XX/09<%*,^ D<B'JXOY,# G69VWO=F>D_U#^ CU:%,$\B'J%++[@+C[3M]=
P6.9E@\$;R))ZZ<.XRU*"+XC:SUEPL0&3>?(ETV _M #ZY?T2P>CH.CMUB0!%-,(Q
PHOJ<MA[8-L/-0? ?,$?ZBUHB:0M3!<W-5_-']>I^5[CN_^QW(UY/YN^:; *_U+-O
P"48P<*WJI )VQZVI*^P=$[],^DY<8 "3?*Y\87V.A.Y#P?'*=2*J.C9\0Z(<9/+L
PPTBR!E5X>V.XNHHL9E6)0K:2U"E[4H6ITQ^=]# !:P13LO.;H5\[C3)Q<6-"Q/%0
PPA:U19U+D&KLY@BLSQ/Y.<!X /P4"=-S_2INT:E&Y^NO9P#>.I+'[2X7%FO=5FSI
P3^_4=^>^.RY,Z2:4UUP>A' K!HKVC!&1X-].)N-;P[_E69\9</(S(3)+$!#18'L6
P.TYKVUA4,Q"GMBVPL*+LG6 =J(3WRDQK%Z0_+K9LFC@T"H<@;FB0[J&,+VL[<GGS
P*CDFS&0D#U/DU\P8DN^T1S#.&K;[/19B7154Z3=7EA4<,,7V0@[X-3SA7*O89\)"
PK_,"Q/A"\[1XM$+P:-IS\+1.B.0PS^[%?S"ZJ;T1/W),F@RCP)H*0W< ?#@4FO.O
P!@L,G&XKGSL:)/H99;9WF867$OVNTB20=FJ(*)T#U&LID,MH\)44=XO*0S$2M%UF
P&_?VWTM4Z[R("5BY^ONV.WO\8 UP)("(X I 5!XP]97]WK IG)J@P$61"J.WW[PG
PCH6J+XRH?9'E?N"[,XDX$#J>7O>AC-ZU)3@2:\\>$6H>)'29M[]CX]$ZMGA#0\0"
PP_61L\@[$GZL=TJ4P1*B8H%N4\/RB,+K^81#BM $^4YV&:\J]WV=YYQ7]ZB9"HE?
P[<A0! X/OW-G8GA<:I3< _K;::HAY]()M&3-0;O5+J-KW3A>0QMQ1$R%QO>J78J$
P-ZL#/5ZZO9D7DC/^!N@Z."J;LZ[ $.-D" :$=2I[\/-;; F$$OSD/';7L+^:0Y6M
PAX9!6[H_<JH\.R[UQ47$UT:CJXW?,M[*"Y^R6-B&^68Z/RX >] THO*OLQ\0D^(=
PV<<0ZHV$NL!DT9-,HYP ^W]N4"17 % 47RE0:'5OBE=)?D<[&T  030F).0!BY. 
PYX]CCXAT<+5K1OV%(R/8U,'#U\C?G6 $HH[0(\UG+%5\"@+,O#X[&6>C4T40J6ZZ
P,Q.(@+&M%9@!GS.R<(@I$U!<\K;#'B _U3G!TW6U^[[\-:*='[=+.?;H1_R?DW&S
P ;!$I>TZ>8Z[IO 42['\K*/9/*:4+'^ 5CTU.:,:34!]=&1TT%EX;%T+><ZWTEI'
P-;OK1"W+9U/_T/BD48Y5T[=,L(XI9<QV :8D >2/U0X+M$PM(DT:)%,W7JJ<<;[5
PW2Y-X*S>[B8G?C:O#E9\Z"V1 PA6!S!17D[.LT?4 E)0;<:A+Q9(:+ZK6!B<O)\<
PN!;>IAUV&  H8C-;,8<M_X_LFZ7.Z[34.TN@.6EI+]P?XWCH>6]!ER(,OFNM\ 3+
P8S$^5*]OG;A6 JG#%EN%MN:%$+9T50&)G\BO4%KDSSVN'SQKK&34$JL;<54,#+_ 
P\+IOVQ6$VKWQ&$]X<X9B %1+RDGUWCC$"\W99>_2SC]TT1WROF=Y4OK^XW&F_(34
P*"^SSA4W'Z:\!-Z:%G6JB/ %F?5,KG=8=0'E.,=NY<4&Z6L^'8J*NX3D*]L-\AO%
PR08><"=UL,$9,K:U.K%#TASVQ3L4&#W@JN+">(V2,,;:MZ L@/R9JM'_(>A._GYR
P0JS[[U'SM;CN:M,/WTJ]=EL+?--F=_),XA<* U,&[U!H+GW@NQ<D;T;!9.R;C%"B
P3[MUK4L\6:9&Y*:1VGI.X@/I "V4-X47O2R=(26%I!4B?F%7%20XNPVL=&U1*%7I
PPXMV(/SIIF%4IQ6_(QBO@"[$Y)XKU[(/&57M'JCP@WR8Y]&1;9+;2/0=$$5$+:<F
P_P(Y-[B1'=4TD).4(^4,V_*0TE"3[ER1>'"N6()G@@OVF$7A!MU-'CX%Y 3H QB+
PR>S-)LYH:)3QBX1"CC0(ORM#*-"'USWNU'"J,QZ?!@D5/BM7>GZGW=0SCXVL#6],
PMF(E14%3G'<$I-REX41<384KO\OSTGS\8:,>)$.-Z"3Y&%NKKE*W]RD_^Q:5('(3
P<&_Z?1C/UA#C8KRL>Y0CI7S17K6/R<*DSPJ\DZI[IM&?RG'U _E_TN6Z>,):Q<^U
P5\L4V_.Q28CL;]S$8LISPS]*VYIH-AJYG-QQ?Y^OG5U.Q-9L%=72==F:."FJKT1:
P5TL6\=RMXJR,FP7/[.";C8[.0MLL''-F]\/[VN9=39 2+A<=%#:(<T^EVS5+^$(<
PZZHT]B>1*2_PAO^'DL SG],]=PY\%[+L<-N8T8YM2EN\Y^='0\M5*'?%(B'<SYFH
PX0Z3H-RBH"LAG)MK$.J5_=-7_Z>PSF2AN>>Y?L=*$21_!QKFHWV/8!_%*G+ S+?'
P;Y LLL_9I07K!@F<U$Y+WQ3P1TIZ!XT?B3L!%'7'V6,F[2_-D>*MA[U5G')[J[>H
PSFN[JI3QK\T@M[L^ @@D<Y2ECD>,LM.=D9]#C5FL*V)@"8$IYT 2F-G6.83A!_IR
P:1#0I];%OW_/^J/PC+)3(+/UUXRU5^.=4*HF+1M.0@#:=OC"+GALY-=6&KS]8H5Y
P#&8]2G01EKNO=1QV)KQ9Y1!Y00BZK6@CITIDZ!*;5:$H_LA6T'89\R;CP9M0INP\
PPYBP3ZI^4\/5H7\5::[OM7, !V0"GNLI;+;F_O;/-J*23.:I3O+/Q_W BOJQVSCB
P&RV('<FDCOHT$5/D#WD(H\1\HG]4P3/LKA ;.B+.L?Y")38.ATIFR026YKTM0\BA
P4@4?L:PW.L6-R$<!1JM$/-R7,CM+E ON/8.<!2LZFAQ3,.JW7,X-IQ3?SNW0IAY8
P283[V%@^DG&"T3=I*!4]/I_[^5X%GAOG9!!/OA>O[^S9K!(>BU81@P&WI\BY9"H$
P6+S:X8B$%A/& ,X4-:[O]S$JD1D(YR;/VI<5_<WI]5O029P+"XYJ6Q::AG!+T(-%
PMD3T? 5\.=G.;!N)5?Z"5]TG TMP773S IKR?A]/$% \(I<M<=]7RK7KIUDAYR,%
PQNH4W)M0 76=6# G7T03?]DUZ/^L%\;S:F:M$#7Z9%:EG-?BI:FW^ADZ'K/\I\?G
PD$:W\,B<KFMVV*A0T;Y"+X89EI018>BU5O\V5 ][6-7X>MYH)WH7="?SM5>"" PP
P&(&.QYT9I5-3,]-G4QA@+W3.,B-2@G'SW_<S!<E@M_/Y/!JFF;TAJM$%IQ$-3&;Q
PKOM)>7W71:?(/:ZI\TJL@<R, +3'C!;&@S$5D7H1F0,H%1W<_TVIAMP+&5\R,KJ2
PON?LJ%B<R2_!]+X=&:)=RB3<F?*5D]6V4(820.>4^Q<QMY<E_UZ0S)83=XH_^AT?
PJ[/6G4Q*4G)J7$>/@3QW0-Y&^X'#O0IZ^,PF!)=%X,.4DD?P235AUA1;<A#KVAS-
P^;?QO,<=.1%=9PZ)9.DMSH1J%4NA)W;)$<YH8<(N%E^+J=,:19BLLOY(12(R_BK_
P2DI:+I2T0''\KOXE7"5HWDNUR)\>GNY+=I)YB>FK<IB6FBAVM \X$X($M/DEM)T.
PBG&/%U[-HI3[8"H,[$.>^XI0L$NV-%%J].6N?ZGE[G =_>/BZ:-\7H.^_G3$&9[5
P*0"_ULM+B,=(T3Z*CD<5,F,[=];"RI#:"2.@''- 'T^CA:C(C'PB/DII++?%T&AY
P.MTY7VJ#&^VZ,CH/2*?"":@5$35[V%L6G)#6]#XPB>D6#H7:_)[_<S.SB^[];?KV
PZ$^<M9SV<1& >YY95\/C?,Y'3(:@3 !A*<D-^ ^I"(U]5:*!VKK92[_)O1KERMB?
PE9/KK@>QC#Y4UE]XVQ>C"4<!YB_G>?!RDUO!2F3P;\!?5KGHD*@\C6J'3RVCA-EL
P N)8J0CT5\P/\VG,ID>54F=@$[F.JYF41Q$[)6:#7D01RK+/?#]69HF:S)1'27+1
P81^#^0#QHIV$H0TBR>[L^'_(9,?,YT]$2MJ))GJR6@M5UW4F3O%^<6B49R/X\K=^
PH+;ZENF(>NFBK0V-G)AGMU0A$A@=$-:Q&"4\&=?DG(XVOYPP"?QR-ERPJ HNH% &
P[9J\FP;.G\A1L.8T^??%J"H-FXR;-!)X+*@42?S:VN#'F_NQMQM5[LQXHE\*1:"K
PG/MH)D]XF[Z K6C=L]::'*T.V/8^Y^:USKC!+=OV$4CR 5F4#V.]BL&_Q##IOXF_
PZ\C')6V3GJ=,5&@$P4ET]\Y@DNZ,WMU_$D**5;;Q2ES=L'4N7!3OMC/=UD/EIX,J
P@Z/C7FH[U7C\XJU4M1^$H Q!#C5'$.^>5EK((0L"]?Z??+TT=S7![9OUHT&[R.(N
P->QE</TOO:[4_C_# '0 )LQHP3S(&E I]DL^06J\YFS^H 1"5F%:,RFZ E"I2/'&
P++#EI0/G6$7$[N]=.(BGM#.)!@#D=%N#*_S,=&FX-*XG05S2FN$HS?6=,R=!SH=J
PGJ0BD]&0UUH7,8852Z4$5H74A9B9X2C3ES.,VJ)+LNGY=I7K/R,G>;)%$N]!\-3.
PR(R=,\Q1M=$%,M'FS^)M.W@V4[0;^P?P2/,I<GNT\,?:(->+.H:3%9B='.O#J=SE
P0U*]%&3CEJ399/A;L'SQ[_H&>^_B7M6'*9WDGE)N^^2_KK'$ZPYAANSOIF+S'&1X
P:3>^2B^#!4SH:$1PW*@7FA1)N^LAP[\#Z)%;X>GW&U(+)NE]0:6(Y.BN!_.G.MG8
P?8TUXCNO+@C+-OY[I!GY#*0/V@K,2LD_8\O+JVL-2=BAT9&[D0YR%I"I&,IT@*/T
PB$)52FIRHBU1QA BQ"OE=J0%N"T'!$\G7OV5VW:5 G@CLSSGU0OO75-C*\L+9"78
P-"KRU >^=>7 >8@AG;"$-O9I&X"YAEMJP#[TM3??=[H=W)-0LF\0=NJZ@)6PCM!V
PE]8JX2&EZ@*5VB=$;5DDD>$S*;8L$GDGG:L\N#L 5H5Z;?GK+=>\"*%D;]7=ND +
P309V'KI(S]H3 J?UFZ$NA=WN7#2;>!.',9>BO<Q^97%I&D!W7)/!(OU2JWG*4<A_
P/74!XW'<M66RA^'02X?[7A7WV!>R^J>O#Y(9'=<LG81SOY\P0?5J.<#5,(QN0  ;
PL@\>L]-G=B;2\R"N@B<O:S%D=Z#$1,URY-,D/0!0MM/^EG7VAB+U6>4YH!!:3V1 
P< WJ+EB5IQ*T[15'LVZ)167F&F%#-IQU]'J/]KIY<#2I];UC#N[LLWE^\A]W_?RB
PRZ$[)K_[8L9XB^3NLU[NIBND<:U/E<&A!+4"G%!XH^K<1X%+_2P^R%W2&,(])7-*
P E/87J\5^!VL)*,E3#_&O*Z$8W9LYZ5D_V<HJ8F"+%4"\$I;BB]0=]N4 ]/!KR[M
PNY74.(/'GK_;WT;=; 0E\.<G5I<,@Q1[37;C)D#U&W]\(U_\(CU[I#;:[-;?4<K,
PWH=P-VZ31:L_O#"H-':67U1'N)2L='PGDJ:AS7+>Y!V1G2MU*'3,U3YK2[--F[;,
P,!:&;((FU[P#@HB_V8LRSV /0<HP(?:H :U4=4)>FGB=\>JDPRHH'$VQA3+@Z,A'
P[\;=CTI%H*OCDIQ:RY&S4Z,',N\10-^:O 2'M^*ULY@&0S389O<4>J$D7 ^M)F?I
PM>>'VZW2]-$?J=& P]1D35FHN[4#6XM[-)*WCQ,/W@,&4,E.;JUX3BHSMTW=%62H
PO+-.+,*]0RU8+I?(NC'?UQ8.?L:JZ_U0:"<9W[MC:<D&ZB(  &:-!8\M-82.Q[CK
P91[6ZC>GD(2_D)(F =N1WE=R/O[IKN8M.CE.M^$7_]!0#L$6?8A13HCA[/[U6,)F
P*Q +2K(SD9,K7N%:/TXN+;PCS^68 >0270RBX!L#BEJ)$=^84P\]5:-<V#YCX"H-
P0T+_@4KSM83H82\%"(9-3 398WSA:<&F XY51,)KCGV>AZ!^@1LXT-1;WF@2]9I/
P/):^.\7Q43U[MNS[Y*\;A/2@T/W#;0Q,ADI-YX#.Q,>365+[LV*L:5+$%JK%[PQ_
P9J^^L3_):HZMNSWL/C<:BSGI_#ULL$(YTI9M9^F4<]$3#-SZ.),1$<$%I+DWM/_;
P,DDN'0*CQ<B5O7 QSF,+@X1*3T +<H]G40H#K*;<E)ZM\%S5%,FH<8GLY[G"(+7(
P8..(Q/!714*<J=8>[FZP'O'M <?]O!&W2JK.<\S+!.=\2#$Q&SNC_/.Y KA\8F!V
PR %0@HJYU6+'N74:SWLKGPVWX;F5@SVXEX2AP!:?HE<H/9$'3$MNT^(+(+=*UQ96
P2REI\JEFK>>3JF1-D_RXGYYU<E-3$!6D&/&L@4=?]=3]VK.IVOS2*!_^R)\3\+GQ
PWQ<E\7L'Q7CJGU+,*5=',SW1;@K88+4ONEUHRL>69,6E^]9&G[LVW]I5H^<89/'&
PU4#*5TK-560VOG@9;E]PEX=.OZWR?1'#&K9*:A6LE$E[995H#1M%5(AQ1<#\?5RM
PRK6-<T=Z:&'H^OXZ#+'6O&LK+M>D[*I%B:RVLR8=/\F1TM*^QW'1J>0H]R\17V-D
P5^8!B&7#;XL2@N@:\.27].VI:;$=EBS$6]@30%A1ZXV!G#0W2D":XFFBWH1N:/#H
P#ZM,T^LR./PL'AOK6;=?@P%Z,Q,(YRU*(77>)(]MM>:JC3Y.+>D&R!FLO(@89??L
P+-\.V<.;.D8+HO Y8CRV#1,B*./%(L:%RWS9?:J3([&$N.(G=]N'](":F<D78YS*
P<^G#8/Q?C9<D>95.2_<"\S5GW?$>:IN.QQ,Y:PG8&&LX550-;NU3+S ZS:U:YS1!
P -L+,C0W[,$EJW2Q:#I\N>)F)M)3,HD.:W<I G'8AJL'@'O;.B+;3+!J6(TT#QFN
P\$-IN+)\B1Y_=?BZVTUJ+^1WK9A(4O1/Y'3?5P+\+[I^C%O5ADK?#]9VWM (@6<_
PWIG6A$C2[ 49J]42EI^;#O\\PDWO& OOATM;(!&E5M]%E/6G^E47//)NL.5^B[$"
P.]M"7C0^^V"*\G;^\UYM=Z/X1#(<P1?0U'.[Q3M(63)/R+%)S6)VV23X8"SQ&07?
P U3P)K:1AB@7NFZHKC'6JQ5*?!4*-KYR[QM/^7O\D*YQ9T&"GW[R#"K'>0WD': %
PEC)$Z$,,S;8FW\4^#4B7W$#'YWM,??E_>>;: K \ 1.:_</'#Y 0>=B#QGJ^C+)J
POZ7?$VOM9>85-#XMBU3$P,3<%VP ?3VF67+1Y?&-Y?QMY#7UZ]O?9#8XS*+33B)0
PYZ\:Q_[M_SZ'QEG*R@WRC2%=B.Z<Q76Y(3<ZDWM0H(+Z'0W?X&#7JPI&S$_X>;%;
PB">/ FV!:JU'VZB(F5/6@.D4B.JU*9R#W3[BI?>8-%=\]:O]?1J+VY@!J+.SI'GO
PD^ ]X&=3).AR)EJ84S1%<\NH5!B!\9.P(30YXTDPQ$5 L1>DLQ>5SK#AR$JIBTV3
PW MEMX!CWV=+6.?/UTN<R4ZM'/0+/'%<EAV31*?8<ITKF*PZQ%X3?_]CT\D-S>F,
P'F2L>Q8GM$Y^09%!K>S=@V0UURN+<\\*]<I"^EO1#.G?OR[4?Z+6E4Y&7:74M?[,
P_TQX;A4ZF6P%C]: !EY)S.:DE5PS#?P&FO&=5\<R8N^1(D@;*S<M])[1D!J&E\QC
P_HOABT8!Q$(9$.ZDY%3TAS-FW>/S,>8^E3@T'OD%ZM9B1EU*'D'D3/^1!&T-J5N0
PC$6=-9L_X4T>I&-N.Q9/42Y"-8 8K=#SV:$IWJY>G%7UI,,$B\3NA3F=?EKG)>]M
P/93:YDF_,C?[M I55O\#D#S[Y#EFRW6F-E-%DDC_>D8VCD4P_:.Y55>7?%8=G5(,
P$>7K^6&00MR?&>=]C[#VYNW??'PM=(,+C#)]QVD]N X941>7P?43FKZHB)*4_\:#
P-K/T#SK+RQ>7FJI"A%.C). [>VD@<[QT+T&3.;0.6]3IN?)/S5V7<DOQ7;.=KCAZ
PS8N836P_@Z-?\F@7<6/GOEG"/AS:,XJ%C+V-1W$2;WU*$W7H IO<+M67>YRM0;>:
P^/2@\<V/*EW.,*JONV6I*I[ EWD_WH/2"DU]#FB 6N%Z7I0!W]",2KN]#$?_81?G
PAO+K#R'$*W_)<,/3#].'OZ0Z)S<!"T[6/6RI3E_&M:'S#! AQ"#+TNJV>Q'TVUL)
PU,7FL.>HN#%8V*&PY Y32%[C?>\.]C5F5BZV(Z@R;Y>$!X3Y_A=&HN6NP$^B,)S9
PS9R2=_RYFT]?PA3Y^\#+?!)VBN;.TQA=F0&&X:(O^@@2NL.)HS+[..WT+"FTLO#7
PE20 /0Z0![**<*QO %#52-LXVU:"QDHB&IKYT11^JS<BF7V(8JJ?MJDNPQRC])ZK
PBU!^G:?]?F/<"\P^]\1R!;;B$HH4^;&\)OR93[*K9:<(E!Q^!YT"#'VYQCJW=,^8
PE298VO>;-XW*;P'=4UI^69Y76Q"F.0_YFXW6")\F..@F])R&I[A\E)P^7^\(C@DZ
PC<HK1(#J_>>G(5LPQO'[,"2))V]:J+HB5@<Q/CKGF5W90+7#NEI Y*+#E3RKPQJI
P OG!0%%>!/_B:9J(6&F*A-[@HIEN@@0R%!^$1:?V7'>W8U8V7;08J!;D1TY@*,SR
PR-O/5)@IR3O2#BCI*@ =IMXY:N:U=J9N@4&D(A$.F_:QCT7Z8V=/"^LYG'&I@\#/
P-=:9D(AL!U#4>.:)Y!<*?%I<,7G9L?T-G+H,_+RFWY\6UBDHQSX5D)QD,<@HI(J&
P:RR)K?AI_/U>Q*F*/STUM;,'FGZ#6G+O]DL6UQO??M;G5UYD\(]/*#R=WAD1X*3\
P#!T<-.+Q+3NT4]QK0<%9<!&1--\8,G$3=8UR^%QC)CSJ&G[A1@:5=#/3;\A=NGDX
P[<1,]02I\N:,SN:JZ7S_80:W*;[IK]J-T;2C"'E!:G@R/(.M'Y978$,&9I41I&6Y
PP5UQ9L-]1%AN(=)!4U?TRL%:E_\((4$7,<;(50:+XI)J]5I68J)$.XE'?!4@S>\W
P%22F["J*ITP9.$D9,_SZ5*Y6;*7W27B>L _U?YV(^R.3.S'BR1MDI-_U6ED:WER^
P><UJO9PZJH0%L-W'!J:)BM7&*'@_ABYM"\07_:RB(4K2&34!5#7?S(*/5ON2HY+ 
PRR#GJ2;>$* 7+\3:HS;P=1R4>FI5,R#E!F& S<:Z[@48OY/2+]^!- >OK+Z1X/XS
P"HE6782[I3;U0!QNS[_Q5SU<>#%NI.&8_?9W:@D88R\)+KCJ70.M@V3^G4EB'+" 
P1W:WM13'C0-P^ZNQ!]\Z/B4GU]BL4I@/5<^0MH(=I/="[DK^-K&&5T/\B.G)>M "
PN\J'TO.**!,RL1Y>QJW->EC802?X+'DFVH(7*QK"LTZ16/)34*MR=D@VR#J6%58 
P9B4N&49NTP98AJ,#190KJ NJ,V-_W5E#:Q3/,^9CT41S8L:9Y&@UH+W] SG$7/<P
P\"H%0:\V-24JFBX(9.(6M%L6&FI=1BCQI%BLXGINR>3C;KVQ1S)N]SD<J)Y\7TXR
PT21MR8_?R4+K(JA%*+#W99D2YJ9FYU&8)'(RD9S>D9KJ>&XN#3L[%PP$?GRV^6>+
P>_F'0@4P=\:8,3F]HVY 4&CVON<L&<PZ5I$EDTF.^2 <<I:;37].NOAQP?":K=/:
PL8\3FXA3(8O]I#H_ZI?CG5235K&/93/Q2U"5'X;_%R5[CRLQ[HA%M9Y\5:?WWNS7
P07%7"(IZ'4%'2AL9RPR_7,7A;GQWURX1QJE_4:%>4;S**<=^H>E,'8>M$*.RDI-H
PC2DR@P5@2 J!$#NV$S>S G+;@C\FC=-V4)A@MN?N@54I^\]D[#OEJ$J%0,1Z'G-B
PN<%8N,'-69^)66L!H:Y6I'S_3YQQ]S'I0!8PSG5&JXA_&Z(R^0'3S!-9/G<&EL6'
PB3%-+1[&**12' N!/52 S"X&+A8#T.;@V32+C.$9BP33HGZ"#,1N155&7[1^PID-
PM3EP=X=%K[01-*B0+ KZT#B/QE(&_%3+GHL^UX^]&-(+_DPW;Z^8N'[@"_9ZX9OB
PX>V(5 F,Q [P+]=41"06NS2E=\%ZZA]EIH(-A5/^D92+9JLV3K*DV7"R.T@8\0)R
PF]!N(EY:$: P[H^8:L)M-\J1M6,-D,8:]7YJTS-?B1Y%U^)$BV#^WW^H=>50'YNE
P$3,2M^!R:,EU4!ITNA8HOV-IO(^E0T'16,CKR!9[;5HN=G):'(AJC0I9PL5+@/K>
P ?5X1XRFWMB,ZX*?*8@]DX;W&2I\DO^DWWK]J': Z(RD>'Z-R2[U7"8N&+(GK[O5
P3\!HI-BWP8<Q':T2@SW.(X3H(#8=-Y)Q1M>Q\F<(Y1UHQ><Z- DYTMI569.66]!E
P\A^TP:N\Z.VZ<>@,.KGMCEI8R O**$E%$'MW: #C-^B/\#R-AS!K>KCU1958W:U/
PZI/7\" ^[Z&O(3+@26T 2?1V;,IL;XLQ/)6@NECC34;*Z3Q-@,E$&KFPO_/JX6_U
P+SG([=W!Q\%BVH\3\7"QO&#9\RRIK[ HX3NH[E%,T#( G,Y%481 U[;YX&/N/:"@
P,+I=$(?&!BT"9K?'_@SZ.+!W9\2C2S_\A\ 6BL"S4=>:O@WIT^/S70PI;)#I"G\U
P4G2PV0&:AD8J33&L26K)<4@L'?F7F8,]1SX%QB& $@OV?'&(6#;I^O'RF1O2FN0N
PR/U!L^@2RQDM <=I@9]W"2/M$W)G4G3=]KESY7?%DA:P9=V%L];7B,, 8X&<.1A3
P1\'].^5R/'*U4V"J%S5/AAP2TF80:/F65K:C?A!C-W=B8>K)EMPJ.$F:O-08U^Z[
PIXD]T&AT3N-)[+5X$HD=W4P<Z*]WNW ^U^76Q99%$JK<M0(S -5:WTC'L?Q91%[S
P?<XC=?[:E?N#6$WOY(.[H!7_R5MP;<8EG&"/=M3Z7_EL?J4ZW":IF]6!AT?>J:+!
P96;9WC8*373K76.I$>%R>,UF(O+&=H^+?65>H6JW,C!\8;W/(V  AC852[=-LFG[
P@Z5&.O\,1NYK_T531FY&$:F@?E.Y8EBQ-X!L/B2_W26/Z"L!H1C(;]-P_Q=VLM%L
P^A"W^+>[;OE).Q@5IC<WC9*WW9"6BQEOP@UZ8P-"U,1M52^HH@=D .F!4]&,S:K%
P*89-KX('J*E]R<Y>M*"%6(?COA!23IT,?R0HCP9^5'U[',23WPOMM>PZDL_0ZFD%
P)]>P,)T_*GX<)2AW?%N?^9OU47RZ% @B%0%0^.JCO[FH8+KL (HSJ07W%(GY^Q=S
P]S,H,1Y,ZJ1I"JHS A^=!DKOVF3V8;(_<?P;M(JX?T:(^SU__&D7-M2.BKKN2%V#
PJQ>)JB9,4;2W^.P3T='<3^X1#T5K@CAW"(6!-_$.QK+DY3EXZZM8J1("_1)ZVAO$
P#DMG7(KJR<E* !SGJNF;3$Y!1B9'^XVO%*A*$1TEC$:"NI8RXRI>?9[4V3; W$(4
P,U564X#0O+"-\[P<\G1W0PDD;XJ[9K+5U*R2N0/H4[\2A;]YX(%NW9JLS3\/[!5K
PVZL$P^6G6FF3W(!@RY]Z6,@I^\K[Z" UO%3@L'T)]KHG41F@JT0@\)"9BPGV8^2F
P7IZ9YP7$0RQL.2S)?).RLGE8GE*(VR%MJ;JF59295L P8ZU.5X9L\&"8:.IU@,+K
P;T+T.>@:K6@7XMIJO).$GMGT\9VC;+1H,4K9^)&/Z[T(=FWO\U]D@VF*V8/ZS5-H
P==,>J]^(2LGJ%^N . _T6+1N*=;N'R;X&7VL0N.?W!]A3PR8CBONX9/C=4?-BO&>
PE*N4<@N1@L ;I<]^QM_2E]-./\KP^46O3+U=\,C_.;:AD7J\$"UE;.:6ZTLEK=-#
PCC0[T7W=DXIUB<8< Y@6@_>00ST1F/!MSEX]Z^P_XES-D5*594EJ>U78#;X7+*"I
PO] +2D;6)[+\' "6+Q&590'USVJ_U(%#RUS3DAZ4[4NA8L+;3QT(7 T(X"%)F1IK
PN1\ 4;C:AT[WJ7'F,]P]5<?!=$Y:83^6<O_8WX*$K%7=?5:EEU]5134W-_2#K9<:
P D%#:+8.O2;$V>DF2WMMOQP-^A'/+F2 JLDP&F+C>\L:G*3[#.C")ZI ]#Z,G2'N
P K+3)57<^5)D$2F)9@2G)P!NY]\'(<ZHRG:TER)99\<DUP4I,0=6 JIU+%HLL#^+
P<!K04^B0EM3R[NE!=5>-%Y%($Q=&H:WV3< Z X:2\EK,5<308<\Q^'FB=<PW2+']
PC!^LVN;N_JDJ^L>TVKPPS_Y*5C_*X&9*UN"QWWEY*1V< /DL'IA4N5\)@Y* KTB&
P/NAM9Q)M)-\1,L?69N&:V?!^2;<"EH10*<0KAXO56F=96HH<W^Z==;#E\R&2/ 98
PGVT"C)2B'M0J OQ0<#=I,,4N[RMU,2U S074ZG5N^G2I<8_!3SOPE_5Z6F\0$T8K
P9P8P],>A;HE.@#Y=JX!V@SF ?"'/1B08)@LO*?0*2O7@_%]TII(; *%W^+.O#W44
PY0T)2+$XWJG#[NK * B&5(PX(R)T>3U-DE)T8#O=YMA_CVPI6L=^;9$=%SVZO5!5
P5="/"Z.7#'T-+IDG,=*GKLQ'I W\3N[#?0[7DM5E)=ZEMU*:#?%5=#@ M=%KY%R4
P!%PK,B#B!LK7'7O\78F[3":UGY QQ$L&@L8@1OA:&(L?TT,VW9?YG[ $HRNGX$RG
PB>\1B'WG)"0DC*T8A/)YCBJ/U;VA'87.!(<;[1%GH+[":S@R4<5PVZ3(]E-N<:3J
P8*[-NQL'?)[..]IH-4[OVVG4_RH\,5PMQX/8&^]I&IOO*&V"Z[FH,HH[A=*<81@'
PJ*JY W!X'/V<3'H>9,J>P2?KIA&D$@@ATQJI;CQ+P@<F]/:[[&L73_:'%%%"6EN!
PA<E9@#,:T 9B@]F"1 HJ6_K;KSNL;(I?'J1\3S-'9N48V V/43]P,0"C-U>83BO@
P#:G5F2?@5^R]#6.,:[[Y-6X]Y!RA<G25YY;O*V7]N149E6U?A%?E 35NR*/XS[FL
PE)KHM>N$IH44%?2?,,?@B.01H#K4?^HTQSUVZ?I*)#BX(_+/8("R6R;.3^K'[7RS
PBTD]H[H-;:J>"^$'A%=ZSB@PF%2Z(3GM';^ORS;0N52CN#%RUHBH!*7+1<6-^J@7
P1-SSJVU:0K-J,D8J5/H 8P=Q7AM3 ,,'$?<"#+>6HY3P6W%-F9WK2=UV9@!5#>+*
PWBO-GMJ$:29+"? "*%ZXW X.XEX_D[ 4#(Y07!C7;RB6KY)ZBUF/RP22,W<4X)ND
P@G2YPN!Z_=3J%1Z:!-Z6 F:H) L9Q=S@P60,=E7[,4X3+$:]SO)B:NJAOFB"RF]A
P+OW76?0.=$1_4,$T#5NIR;16VN5;)/6+>R<2*[X_:1Y4@1[X+F/[*)WR@>+;'ZC\
P<+\<H;^  D 8X5^+*GD)R3,M/9-8WM9OAW1^JSA*(,I09$A\- JJEI0-)[T_C:,N
P2R>?=P,MINJ\S\(#C>R0(^.I#5!N<2H_<V-E]-O#=L38@L/K5G _H;*/%,Z@<"=M
P>+?3:N57,A39SJ3;BY!%/[*M.F0TM4U1>\V6)1M/AD?SJ;371H=/%!(Q&H_SJ76V
P,#+*ZYQ%J6I0U_!K?_PPM=AK_=_^3Y+?ZX &.1XG4G/IK>-"GWT2W# 5R-;+^7;*
P].Z*/R[*@>X6Y%*XS,BA#8??<D0I9KGN@T+CEVQC;G]O/,/X--; :7N$*\^O2DJ(
PE/S3&@CA$@"5BM<\VK@0^1FOU@!V*3C6E_F>>14RM.5M>U?@+T,;<7GHW]&F:=,Z
PTM#6X3[U]9J"72]KN:A?8)9QCF8115?>],^D)#@1OKF)&O&2WH1@L!:')+J$"],:
PY+>++Q@V6SS7N+\^/"H KEY;$RF@H>@=;VGV*$N!+LX6 ,5O#P@F$#D=8U,K/IYJ
PQ;%16T,J8?M ,R$>QI0+?CH*0<H:ZS0K ^OJ73$J:^_:8Y[_&,),=C/5'\O<H4.7
PXHD3[[;$YV6^FEZU'C^$$D?1^/P/?(_VF)\!+'5[BBZQC0#-!$FS]59<>Q4PKG;_
P3<&;!LC"Z _H0P%O8H,\_CVN?:[UTA_]T(XGX^H%8[4#O=#::L+MP< $:![:@>%6
P1[*4=L"7OT,EGVT\=X0W:]GR18\L'(I2@'ELOA]$;#J +&L_T!!U=X8"5!)]D&9#
PRF^U^T"_@*P[?RB;D80Z0?(_V)WS;<I1V?8G Q/Q/K"* AQ5%$\Z>(/23<&+R]*/
P#"AZOX49OYK\Q%P,L L:#@?<^\D U*SR3WOOC7+%]!]XJ  $/ODR%N\P>_?HW;<"
PL-H([.B&#HR-LE+Y<X,5"6- M+\HY#E !,;*K"V$7IO("ELN9&HYU89*6J(%+8'F
P*2FZ8_."M_N'!=V.KGFXA]9F+N#<X@,?XH+PO&VSX6'JQ[#\^>,I-5[H2%3[SC@#
PT.H-[V=\O-#)K1MAUWLDOB,%S$9/??9N(U/[3[@1LHHHB8 S-9B>X>^1GG2&BPG0
PMDV\*4.0SY].S2@P!NM34E3"!OL1,;B!S'$A[?>"VI((BG./8RN=W)T-A!FGC9!F
PO76Q(U-6R&ANZ CZ$QS.R#54>E/[6CJAH'E&W2>E(L=A/ XK*Q9FQ&/[($61MG<!
PTKAF0H$'UZ_0K!\>NJW2KA[M]]-ETZV77_EZ@(O'R&NQ^"N@KDR/-WPN"H";J)\O
P.WOE[8='VN"R8WS^IGS$$\<0 <$_N=A6BH!E<0U1IN$@.NC9X_;4K85DW(T="Y4L
P0 [Q3#^+2"^8VGT?=M.@IQWY7']A;%(7'6N!/Y]=;T4..:YXKN@MOJBN%VRV*'FY
PJ%/\@T?;[>S:$_J !I)8,'5QRBLB&(GL*KE-WI-E;,-;KS&(&OY1))A^R1KN)L$C
PU:C9'G='-KJFU<H\ )%Q<K]C"!SJ'WFSZT&?X!L?]7T) ;"'<H.VIP/(Q#&\($;'
P!$ <IF$$BLXBT_S#+<%VQ?F.0XBZY0G@G/R8STJG]VHH_>2J3PTB$V_(KW=(:YU7
P50*D,]9+JZ%?)P"&QUTT!DZI$;.-^AIXYOG1-?SS4T1FIF:_X!'\RPO)I6DK&6)<
PHMA3_GWU@T3%ODI2L*O=KEB/<(PGO(37 Q#OYER>BF<]*?.=L@1ZJP:4GDUA/D #
PS]1FVWTA8ZG08X;NY0N'-!@0+:__^+_RM#FG;$0"FK6X-1W@:EL/> =ZUI\'(4VL
PU,X9EQO_# 7!QW[M30+&XU.K>*_<W;.=E(YZVBCH1$ #1B^X),=?;^PDV21NRD*2
P/#U9YLHW7U_Z1ZDI^7?H_ZAH(/SX4)AVW'H*6X6;#3Z>&+SJI>>B[P^ACQ]3:\+-
PA'??BI/+N?>2 (U_"1C][^4'ZP_>6==BH(4^HYTVY-, A#Q+;"@)J8F)14>;SSH!
PQ-+5O4=P33C)#YC9&.3:$W4+RE8CI(#*]U@;@U2G/QZSF]U&S=[EP*2DO&;S5LA:
PS@-XO;OOG;D+L01@O.(\$4Q!/M/I_4LMJ6UA(UDVS3FV46,\?;7^<C)@MP%Y+$3/
P&4>#^-B##F%KY)VK+&'4@P/9A[4%TQD P.N(YT:PY^=*KCG+E3;E1#?-#L-=O5U2
P?D6D(]J2*0)VW\/*H=(BWT[+VFZ1[+78:E6<?P+_[)_<N/1<GU;TGGNVB)BB+80/
P]>'2[A:T^JV',H2$UM."F:U"EU-(@=5Q,,XM=F<S5!4XJ1 YY5\#:W'^_P ]!D?G
PDJ=M/S6N'G6K 83B:&>WJCEOE>DO&*R.$X]T;.F14.HW<R"RQ%1H&#AI_/"%/MOG
P[<%;R@MR?E@X(;'E"0WP2\-JXR[\?YC1BU2MV2W"2N:^2[W.D%;GK5]IDB8I)HI_
P(J.V..V'F9$B N! BN)I@(IZG5_)LO;<J^;7F4<*E;66L6&1'I(0!</O*Q$5+\F>
PY<!&;#TZ^@TJ-"^ZS$EB)+L?CS1AI"/@#D C!2%?_[B)S'@+O:Y #&EKON;V+IBX
P!KZ/Q;'T=@70;.ZAR778U^J Y[<,Y%*N@+3\L_=CR4;4_[QDA&Z<ZBG'!OOBYJL>
P#7N)%N8TPR"?-7#S:N)Y XAJ?LS,'X8A? NW$LT@DRRT5(V!JJ> ^-LA_IPAFJCJ
PHD<3YU_VA<\X"8K@1I.!(4J6#'A%&UK5I>L$S@:DOD/=S/112VLO!7NA]Z(,AC[7
P1<1/1/Y/.\<A7C)3%F[@P<9_NY=((M7]!],*V5 <1:)36 [5(*X%-*)0!%[[X5G?
P,W*$C.@/=R/4L1ISRR1>TE0T)7^F@9O!V6TB2+::8Q'2^7S7V(7O]T3#6A_C[U/W
PW%ZTX&. )<5Y(R$J=4JZ$G+;(5C=E@&/R,K"35H"49.:^.PJ;7GPV39MC-(<U5".
P8GI._4.6@?]-6"F'/G;M1UW6.V^(]N +\"//WX<8RS[]BBLGGO!ZN0HX).N9N"=!
P@^)'_,+U6'XHJK:8</#]5&'F9&,& ;ZRY;6V* WPU@A[$QPV.<R,19Q0)<+!XU.\
P?[FE$PB;P3O$/6S)Q[WC('!+)T0N.++<]:/C_*-7@_T#._ST9!Y9ZE-F@N[TW8X^
PQ^@+KQ&YX(U827A*\S%WQG )U>UI16'EQ]I&]:?5BT<($*R>K#TX",Q%B7E]373,
P&0[K#B*2SQT/:Q+>T-BW-F^UWI&-(5K8X]Z=$*EN/(^9/P/?$'I]O'F8PA-?Y+B(
P(7QYWKNF6E6-3"=.JI^7NG/F%L$+:ON>YF;%T\08RH =_L7445IA>,S I[S]ZT^:
P_@=-"&X3.SJ2*_A%@UOJGHQ7L:K&D*U6@!*S49:7/[? ?D2SA+K2FX'FN.J))@H1
P<GD4JB92;@B=E-@*OW.@5QEA4N4YT_JJ\H[4_T%*6()[@)S28,ZAFGED..%5C?#Z
P2V2:<*)@5Y$@!+[;[6*^ #'0",I$?68JBC]9/R9].A<MH^-74C+FL86X=-*O]R8K
PB SFU1Y?%6#A"[\#)/+XNX*SS"ISE%3@O6,AJ4[X0Q=]9FWM%4BI8\LAB)QBHLXE
PSCLY>YJIMS.%]FAT<MI\C=?.6:/U'PBZ:.T-$I'3"67'<Y\;2$!/GV!0YC./K6M\
P?H:\_*)W;VM^;DQHQNP>C"@DB.C ,\;0-8UP!TDDOHGTAF%1:;EOP@-)MBM/)X93
PF[>1V/GHRX84XL?1+L9JPJ_3RKJ<MY,C[9,+NSY'E]&:RO(73G/R;Y_F]P\?R=VU
PS$>P^C(4K]W/4UA7ZWQ,M2C+,WSYI^2KH.NXD8[,]K;4#N/X6Z/*,N_WU=;D)$FS
P6/?85#!V10'>/(,63^4Z^;H$-H%J95&&&F]T@]A+#'C>2 ,@+F*Q5_N9UU+X!F=;
P=K1GV0:^R07-DW);@!F\,".)&C#%S#QU*&+7<3)O0JIIW3H80B?>':C-U)@O-VF!
P[G-+1F2%[YKNNE(!*T5R-?L'#V<.@'Q%MHN@(861?27T386*XKB[C&[84(F$OA*0
P@GI#13MD+)[[-RNYS@$E7PI4L,C'XVS6AYD 9Z4,L?N('K?\9-H3X(N :F#H9Z54
P;3J$U.<=XP1&# 0<Q$G+?;DW=P]M5"G!/\Q V13O+62ZV07 1!C^ 7;AV]<?DYQ<
P,K:-7:1H,  -Y*=1!9N0-S8S>R)3>J]F S<69"8H\JC>MK^A+6J2)OA<:^J.9@$J
PE-*Z5/+)FX#'W]U"XR2(#LE%WJ 'H95N"W4#$T3&%9:OZ,>0LO=XS>M*>(8\&/#J
P@6GQYI%Q44'_BQ OJ5A71*+]$U?X'LF:MHY6HX[Y;S3R[I1FNX%XEV>9MA4Y>+#L
PF)0M&_HJDUSA:<)1,XO:Z(-V[CF47OM )$Q+T#?!SP+S)&8K"G1I'Q1;475"2>8<
PFPVX&S&;6Q>1US@M3L&%(NX XQW"^.P\^T4C3E6(8ONRBG'M&5@@M;C)PWC\8X4F
PUS! /A10M(H[]U(!#VMZM=G4^D+ HZ5V&[/1F@V&-I[8T<IQ%\Q6E\VOCV<[QS]$
P'NL4C6.R- "<T3O/Z)@XMO+F+=!MVC\\_?[*?D 0.=;_7J-%@OPJ""Y3_AJM*UP'
PD"CT@F2D<R)-]2>U[/YFK!ZV;.>C>'?)WY,#W@EYW\VB-GS8S0A^0I16':9)+8Q0
P#:F=Q?4HW1TF9*M0RDVO[\T@DO<V_L$+PSG;SLS3=$AUGS.&69&UIUS>E+50EN61
PU=.+$ZPX'LQ=^4C?TFLD+R3;6( B/1V1YF/)HYT\*X8._)FE/#HZ$(MB%=5#+E*?
P'AV)"<0A$I!A-Z,:7)8+AML_Q$_F+!//D0KVVF[ASW[?,J+M>L51 S^FJP7_&WH>
P<J>1C"#.-NKQF7 B==>-8"CJ96T682Q_[WDA$T9))4]MEK.E9/6@0K6"&[%JT40+
P3;.EH7='\*W@&?]6O?A)>;5 #[1,[=]55&3L4%@7(N]6BJ+2]D5+FD1#>%"QN3U>
PZ(ILK^1HXNP]0A;<6XG(0(4LU?PB^%D9CBB]S-)DX5@R=KG#O^X)B%L/#HFWJ"-.
P;O$.;!=G.E8H]@U8D@BXLE!UQ\<!%<#.!XD6 WTGE[+4X$;:PIN;>8\S[FI&1A\C
PP72R%0HJ+D!W=5?L';)$!ZL0EY$6V;$3NU)$DK6>RP"DX&]VZ <=\"]I$\]^B6:O
P2,W\;6O;BYG0LG5,7+M?65E8P1=;;3KL.UODQ'2D$WP0RLSLQ.7<IL-7%SM_JU@Z
P:;N'3N1%2)A\#XQ26B0]L4+/C_UU)\@G B4TZOK-X8F8X;5;SNZK$BC2CG%D6+]O
P^K9?+)PS86NI1MB*) 9;YF*W@3ECM-<S6^/*(O%1N:@MC)II=M?YO $+6_L4M.\H
PM@:YHF3OKZ]L7*GV]W<%P*N.3Q+/$3E+W[5C-?_X8M_GR6'!8N<66M-"4#DI9U:M
P8)ZHM+#V_F%+=1,+J:V/=ZJNY6G*:J$A)N44'!^ZC)$M5#'YD0!)).[.BUF5H*FD
P)GJN2F?_UT4%UE XT["X;BZ"S)')<:>YEY$.K@AEZ_A!JS(-:,Z*J?394 KCFI_1
P*CH84CU031 C%7EU9[%7ML>SL0%CS*Y.@?X[W]WP[\NV>ZY#4TLIXC6DQK'2[>T.
PLY6]#ZXB]4*??77SESWFE=>P QUA"W_>83/2\58=Y\5LWH03J!^/(T$MA?6"6KG#
P3*LC4!N1YIXP'PH71C @<M,_J=!2]3&KZHE ^<6WZSC\L+N]*B/\U7;5G;!H/VPT
P%!YY(@\IK!0$>1 =3OI8HY!I@FLHQ2CC92##"RGI(S7?WBAZ^2@:3989L+^0K_SF
PX_JB'E=^8F<1]\\J0';1C8XU?)X*6BPN&^D4]!@YKH)H0=%^1BC"F)XR="O!"PB]
P@2C #A'\,=88C4Y5_SUMZUM]MV ;OYMG*%!WYI1K[Q1&CS>-#I:NH,=0^\/?))78
P/>8KZ%YL,0)?D1]?Y!4_9LX7&[L39'92P8VUWPA#N(('.48S@.O@OQ,OPH&6[6N"
P O+OD<9#3%O3H%DE49&WBZRM1N 9/I2BW'I4",4ARL7A:AW,DXC!K3N$:*PR%#)*
P !JPL34D+$370$CO^&C!!"'<J$;;TT4V4!5?A(M%B%&M:O4UQ4;O[,$]DPA-:(,N
P.T$CF^NGZ*SCTI;2!$^4EW&?]\RH!ZEKZ6'I4PG<)0*9(!XX9H3F,,4R,3%JN^Y+
PPV>%(UX?!W1?K3=U4C2>[O44 /<_/OXRY8*@@@'3[QDBR=*.^ZP:UO/Z6;\7^YZ&
P^L"GM>R>F4CT5ZVPPVY&8G6'_#RRUDUY9%^JZ8^U*68R+6 K3(U6FX0S="6=D.LB
PP"B)#5\EX135X0'WF; R;';@IBM'R^'A9,;>T<,-I,,-:VE684*!T<&-A*^I#<J7
P6SVD&E)7;1$219<[0KM^5,4[LRQU\JO! 0_2IHW!Q>7A8:OHM*Z]%65",GT#H L\
P\IU/&%DLO^24Y:);ANC4/M"EQB5-[""WG9S0L_?R"G':KGW)NHL'_E4#E7;NK2)V
P&07/A&D=;;LB_Q>E<O.1L=2R8ZLY[5ROYI24S@R!_CGW?7W=7)M8Z*=7_,+K7D6(
PX+Y\Q6JTQ-7_%"*XS226@1JLQBTZ3BR/Q-??8QWH3-/C/$'V#U! : /]]V2&D<O6
P6U2<795L$W]+DY3SL?9E1 .6C)<KU=D'Y1VA@KBG'E&E(=8/#X2UQ^4J'&.IIDG"
PV.G2RA@S[JUIP].;^L'S!13 5,&';94D&>B[ZMYC $OT,M:GX'9>&)ZX%0K_=7PZ
P<Q4REI$Y:+]4Y [_2CFF@5/J\%>*]H_X A8E[SYCF.$1-OA!DC3=CIB_A-K3DX.V
PP[%#=+6P_^7NBRAR>6:?JJ6KXV*Y*&JZRC+G33N-NQ4ML_;]VP,.YQ0E_Z21;5]S
P.!3@015PB,%.4.B7>;\0W/Y%%8/[/W*83$\^DR@D;JZ#T+!-LWMC:R:TF:XQJF!0
PIJR2W?]#,,S]SY^9^<PF6O:YR$C_&"+CT^=A%@S%Z>K-_9+_^OD\JK 9M@+;)13*
PO@$L8SL54>!M,)Y]B4BLL9'RLB=Z2+)6>ZR?]!:/YM3ZOK:H]7<UKGI=E@,$T\O5
PTDBHIDN!WTY.LE&  L:*[^EL'ZEE?J@2*Z"J^),:UJK="!3*(#0['9=.PL'65%2"
P;[1 V;:IA*W^2BB>#6A.RQX)"3Z(1S+YZNY0\54S.SUQLJ157X/'5 35]?43M?97
P9:%D\WG3-FEJWY ^@U7+;3.1$^^45EHFT;"8MV]6VJ_EF"S0#)I"E7B4_X^DI9+D
P.M 48^M;&K;4RZW'8E.TY9#-# *,A9W:RX52=#8= /  6:):XR"XX]<.I^<FIJQ]
P8<.O2YW_#VZ.N[JKE/US@R)9>!>IOD63M-&W+E0*G5W%;Z8D!Q "\GR5$LW:_S%T
PHG 4C;WUTM9D/HQR3/#2NHBS,5ZQV0 9J@E,&666W6Z+! 2=%6A2)<T>T/-5R55D
P(.?F-M7SR\C+C7BB9Y[/CL%PT@P+1)(W=B9)NUO$!7!N2T+1G-#]?5.3_-MTQ(Q4
P@T(A_APP2>PG5LRTDL0MF&03KDZ<P%OQT9^]2#:PI9$W^(QD:(7;(1;XL -N]/#^
PS& :5UI&5R/Z<AWTQZ3Z_D9C=6]5F_+PLZDM/M0)0]F"/00V]J<%QW4CQNBTP(18
P1C>L1]R5E/8^#*=;41FK%')R\=X+++1P)+QG:GKX28T>EW1;)1/VJ"D3\5WA#8%P
PMGHT@>A8,60EHXF""WFK2AYRB=!,)/6\Z6CQ]&V.RU %D/UE#HS.7B[U% (!!(,F
P$9Z=%8J4L+ ,:J><MO.E22=A0N>'0^PW2X>G8]=][S7/BTQ@6&1=$4;=K2NF>+<_
P&%R"2"AG@:ZD]=/>%;Y3JWZ&79L-*L((53_U>RY%=P!+E$#RE$^5Z_BY[*Y6S4 C
PGNY-,#?U+?1YR60E8PQ6,R#&3W?XPLO!=6=H9#Z'!2:/^A*+!%6;P1,7+@LX:&L!
P9J!NOYX[H"IQL^BY0-65UZYL/B6#C@EQ;EL,H,ME]/@<0Q/P;6-Z9%B'DW'[DS@4
P <#K,*>XQO/-0OT9B7U96,9A^5:..VX^Y61?XHAA7\JC4!/0/0/C N4IHH-"48!I
P0)8Z]+14ITX:V![\%&P+XC>8>9U?;UM10T+F4HES[2X5.U%MMD&=-I,:&RVTB3<;
PW H#G&+S+7^Z2IGOW3 @9;+C9M%TY ;(UZ^Z72RV\Z&F/(S%T>1@=3R"6PQDSJ##
PK+(I<]Q\L^)9?9S/)= EMH'S:3H6YPPM^:+Z57+'0OPI+/]<UH)^KG2U(9=U[0W:
P@[T$"?07SAW"\O"!F94TR,AWNE57?D ''/$W\5GE>\E#[#CM?E*.&"!WL>I K"Z)
P9_HM1%4&.=Z@AD$CC'3Z? QZ%AEWX-*_'S'\\%TM$]ZLVLIH5=*8U8653TLL8#B?
P=L0HR0H,V'F</SV6W.0MG="2&X_ TD-7_I>\&$:=S1DL[*C%O;@Z@M>WBNC)RP! 
P2'R*MD ^B:C-#%GVY*,0-;M%")B)6KJ=E&@Q/T. E=5%W8EDF7!\#. 6C-JHS8.,
P>//X::2P^3<"!KPX-NB<S5L$,+1\(C^7,K-D=YQ31SC@KS]]%\)E>_5I3;]'CD/$
PD*Q&2&:3>831OGM<^GA*'W6-3@_GFO'\E>M,)'ICKP^>-#*,ZFJ""G9J.1!\%GS_
P0>AIJ-&'J.ZP?J^)D]%@-$J":.BHGN7J$3BVOZAE=(6!#W_#OX#Z7]1^7WR93L%@
P-Q#'M:V/6(1NQH+.^S/KX7>88I_9;OKA[C6L@:K'TP/-B: :_O?C&X:Q8S!-/][X
P'=._=7:[2^M AR^?95#@;R'@RKV].W*J:L%*J5@FZ5"V[,!TM<HR=<5(X''=DVCJ
P,K(%2=CF7^'4G2@AQLF=<B2)?ZKR8MKY:N#QD?BD%X^FJF%86LPIRIO=[K:A(+\L
PL'=2[DY"6B#K,( EV%W1M0]"L*2SL&,"#&<*$G E1NT?R># 8V\;@?0H@NW)KC8D
PN:5LZV<[W0:38#FXQ/ )]>6:?#J<%!JR=R(Y^G?<4<VK^; _\FPC>_D"D\/MZ/+C
P>EE88:NZ&\/7O(-*V>^^7'@ZD,#2 Q.TW7L0*F%C%1^]=D.OZIANN&U-P=*'$M\?
P @#AFDIGF5CWRMC(ZXS\>/]76++X!J4%IWY-\VO@+1\VE,Q.\7$]'7#*[Y8J*(C/
P1!O[Q_CX8&G!SIHC/?NU2*=!:!?O(I#[4K7.>\YV0I=9:@+/M8MZ%=<45AH) G.D
P#>QL.?4(_WC$9R [WW( G^.;!]Q4YF?:X:&"Q8T-[*F@ S3=*ONK^1FSZ J<:XY#
P&A'JVC<Y,HC4)6.=&1 (X> 0B<(%#6\.?*N!M+Z"X+3[5WVM7T=LGYM_42KC.[:O
P@I$1J5-+?Q.B8Z7&SV*2IX)^-^#!*]ACOK;)H]>G0;_5T%L<@O<[4>_7\,^,FW@?
PMF*[1,A12;%\2"=?,I"W@%C9JRC\7>+$;O9AAOS/5IPTYUU!8XP1"M,FZ0.Z]@+-
P8O(YL@-I@%7_&1EH9U=+$JO[N"ADEN+;K^H0+2RD/K4UP!&E,ZJK0C:TWZ* 36<G
P3:-?W^E/NORR+E:K+S#,(=\DRMKN2J%-)@&Q#MQ 7FUDFM"(W61=X7H47?V?2>X:
P 1!8MLD[^.:$Q=1+$ES_N[I>&63LY,BTE3B&L<*).]V519BM_M7\&H'3"3J W\!D
PG?_NKH9QV3'B%XQKA@\1NW8H+Y!_NS7<3B]FV#6_/ -Z;^&LIT79[4XDLHKVD!^6
P3KR/:<7>G0Q\*'E]*2V"G51TP#"R1LZE/$X-;2X]& -@7KR?=F](OP D(NCE%)>T
PMV%'JS;I9HEHE=CSCX?E4[0II?OIW:1N .6LSHQ(''"<%H.*(#]6%BX>U_?.^UJ&
P@Q R%J^SPV"N:@0?[G^FXZ2;3][OQ(O@U&A:Z9]A$W1VGMLD3-H.DD?WL;-:O?*L
P4@*C"E-MII99:9]4Z%D _2.WP(77JI+9]J5I%8U#+ @CU"X+5G>S'5352A?>(PL2
PCNG[V5UCA"-(I*,/ZH](40/VV')3N<Y6BK3<]C :Z<^J4AC)4WT5JY9=M(3?(I'S
PDK+2YR'6<>>FN$*%+1LG<?C)':+SQ,[!;]/>/V;*K)L[)K+QV,Z(T?@DM! J-<U=
P(*(XP@>M7E^.2B+%/_7W>KLC1ZN(Y%A%XY^0IV(XW&H+3%,S84M%S\V(T(]4X<N(
PM4_'?OUW2Q%*57F@]&K+!$11&JH87/WG"_+[%YD$<C^VQ.R+I[U-M(2D'FW0$/?7
PUFBB]G]G>7A#:R;)DTLZ=!2P<%G5AS?90O;[4;CI!10_\(;@'84.WOX2BX$R,/,W
P!T_TL&N\/Q=!YUCH+N#CENJB-P.&:ICQEL-Q3$$ZQ._3C$$@@[O3PEVY3%'(T"G;
PBH.)<F[)3:LAXC,K<]UT82Z5IV]&G R3FMQ+"%0)4]4=U&IJ62EQ<J5W4->@56#F
P+:?::%27Q?Q3IQ]WBMWGR)Y<4V-QB1&)T5'9D?9H@EF*%A>H&<P><A!E-X4(T_H.
P\=QD,&\%E\?=K3KW8/S9KL)JAN-1*9 WND.D->_-V;=^[6U-6[0R4J$-#(,#$IP9
PP&HT&?UD-%P2@ ABE+0CT^!W8_BLH27DY.^B[$]([M!)C.LRL9>E7N[J^JKY)ZJS
P-RZ1^B![TXA <^(U*WVF/$,G\&GX7/DN9%N&L/&DM>'DX"$V"(H<XQPCZX!IMN&Z
P_NJ%OG*.9@+$]C@)KT)O-,G-)-#X!]>YFGDE_7FPROW)F&?1/GU> ?M*XCA&&O7*
P?(>&RML)&^3]HRM3F>0&_G9NK99&:%NUT.9!F4+C2[DP;,C?V+"TA9/#ZDS&]OB+
PA;OE;:"3Y$1,^9! Z<HD_9![GZ^JY=_5ZDO[]"?2.*&@B]6#&1(T,PCQB81FVT<5
P=,R447>HCOLAWG@)E\Y7S:5+JS@Y XV6]U2Q114R$3Y$7/FV&8X=W<N2A;M%<.OB
P(R;FX90]X<O,! 9W?$6<D_Y#BA;T:+4GY7*3X7'W!&Y_XEZ+;;=HB2(_"7A#IYP9
P0&VHFN0F4,Q<,)^1IHG+@NW&LZ*K7^<+V&WJ$V6T-!W4=7QJXB%-]-3^T02S#-/P
PDS@[SE\ 2CA\LHZEOE+J[MXUA!27TX>8F3'K=RT?W3V23?HC*GU<Z0)Y0:3\&1.P
PE=E1_N"X>WO*6#Y%CL%(J]_!:M^$D&I^P9]S +@/T1^W%X:=E<YGD6+RJTV?@G!H
P '];4QU-<Y[7U:S^"R@,]LO4Z1RS.V>%VJ?S?1(I?9\XS[[61+Z/\T5:Q^LZ  JG
P S-T:Y6$(+./&0\$><J7<!6'F2I>[L/' EHG"/+PDVF*E3<DY5C;/&."CP[_RG$1
P9JAKXV"A[21Q+HMB%G[C7U-%XW?&@977TOPJ9<C">Q[SM@GTV!>5 V7K.O&YAZ ]
P%Y2&'7F,Y].I6$"JM'A?"0+VK+VKDJ.0H#5]G12!<30O7RDT>L)>%HKU(9O@8X8H
P5P0^!C/9EOB"5SR;0QYZ4A.9T9:1M#MGO%I?"4<VVOKHB1Z?S]I8Z@E2 AU-B;R-
P]GO*YSK@H#"A3A'=_Z'TS^/E3'L[7AKC'P,O9HH@55G*F4+1?[1_4_JF"A7"B(9M
P(<R[RAQN+D O1.+0,!R0883%&*/(U#I,OK5]7+<CQ(_*_M5712]VRL*H3M(C_V"=
PP>("JTM@S@Y3RT^;&5_Q],YSF\$@R-93KB$ ,$O4-PAV-/?FR5S["5#G?\RQ3@OM
PL"N5_,=$)CQ^TE%W^$0\4+5$_7@;U(XNW_3+&!I&%/9&1=Z?2!1O8X)_9D(<)3WV
PP?[4DD;=8E)0[I*(:0"N41 DIMY;N/'^*=Y]X8S^[\I,*BP\+867[8?EMT9X._98
PRH/./"VAN4BV4&K>OV46G6KJ67,;!T2"T\_=^/:4NDE[ZK\HLI<V&![=&87SZTNC
P/7Y/RAQ\"JOJ<HFYERQMT8*EG!SD:W9H?__T]@^TR3ZTE4(=$<J>)-:>*@A%4:T_
P/M+TH=%71MI88Y>Y_Y4J* S^)\TQK4>_=S#)Q;T:)>"*!U)HCP6\,[YC2.HPAN>%
PF!T,L8'*!U?PB%UPC>Y9RY :#@P%YVYV?HH!V&.HW4LP>XCT=82+^Z"1A0'S )8W
PZ+%'>P67C$OOZSSQ+UO\BRWAO"Q!&F\+9P +>DCN3_WQQNL$]&S*X2:[HK&X5DTP
P>_18,@#S[ 5P[!(]-R!\/N(=ZP%V;@5T%,KZXVX@^C)=7AW#C,0V!ELR<WL2F:@\
PW\RD8;5;6 1@J*HB"(L4@!JV@5HF3+$3(3P_?DBEC$/,]C>+?-^X+A%>6H>;\5E+
PX*C\U>:VS45<,YZ.VH-?:D@S.K+()=K5DIL'+1T\S7!.=4;&==]XRH=';V+TAEH+
P;6N568/5[LJP!NI[:8=0+A*1M-#,?%3OT8G9_[:S0R [UMF$?,):2V_=YSGT&(OJ
P_3NUEP>:D=)NNN1O($!^Z7B4"K!>7&Y%,^LD>X<-ZW6)39A+-Z.19GZ7 UG%+[E1
P2,34YN+F@LTW+1MIH#9#3N%=+DW["L"POFQ*,E6L!FHSB['7-^):I9/(I8YU-QU#
PLM]8?2]F.H U9)_7P.YYON";122K].*6KJM.06VD8O,6(R0Q]8;=)FY0+2H0J)Q$
PKV'^ U"<0S"MA^S$S7&5@KP<DIE\H(-8&#I26/=<Z8TK8H\2>^@,DQLQO+<#$FSG
P0[0R+/YD*=Y ]U[&UD "QM)^+7YQ8H^:,>5I\PH)VS6)'#DR&G;?2XF^4M'G7CB<
POF82=QSU=9>"N($JK\'Y(T8,QH<;3R97R*L\O3=Y$G73-7%Y>4>[BNK*GDA\U*/Z
PW90+^I<Y;KV=Q.Q1AF@=K<@3UE=<[+/YB#/?\V*'PAL!H!RM9A[3_OD@N/=#D_;C
P[K]S2."WXAJA3R.MFZ"213_+5W[*W5"%=N,@#Z=J+O^:\H3>6M3N="0-<P;_A !D
P$(WVT\8*%1L"?1Y" CNCMRM6$/Y /J^U3KP])QB',ZL;!Y%!4#,^B0%^FI:DH!PB
P@_"3*O1UF\A R%1[=7[''W70P%DUBPC<F2TJ-'PO"1EWE["),<'?]D5F(W4UQ/=:
P'+>.#LGFPC)_5ZZ^C6\S4'RH&U0C+#53X!,LY7RX]NW0$1G2_/=AJO?UP.]=4;6)
P2DZ%!EP=H9LVG@^RRX,E*,>'6V,41XJC5ZJ?N!_FLV28ZNRT*?8_#!B'JB1*L\S.
P43RVUGFG8>?E<E3+[]ZM_OU^EC;00AS>! E*27<1V#.-PKL+2[+V_$$;#IN*B%]R
P>#82&RAO)J_P^&-PMXZ\.1!Q8P"15<!!V[Q86>A'FI"W"DXTT7V;Q0+:'I<!#Z!B
P$^@5ZF]LERX#MX6'[A_]+8960W1/1KWC456P&1@41K#"E<9A$WSJ#XW>3X/F:-L&
P Y<+AZY$"A>XHSO^J%.5B58 "U@-K$U0U2Q%DJQP[#J'X-'3$+2L5PP] ,V8ZD/Z
P 2[QB[",QMU,=N@I'N3_M7V5GRQK>9<M(0]A_4IY, 1)3P;\DR<5OV7P?=*F4;@]
PLCDA;DY@.W'&<'Y?/IGV^?M.E7&()ZW-PG"]F06%G]!" &)+.P@K$%49M,-*[:F[
PQ"' NS0S!UL9;15L<6!+075UB>5ZY^36QS *.CQ<3XQRAF92"\&""D5#Q?KH;9LT
PU4WYX_C!J2"/P;2LKDX=*))??2W %0KS&^"[ ROEO928=>651T"".7-!>LNN"O0 
PE#VAA3O+\'V@]*US5.^J^><2+QW/?AFT(?G"H,A2.Y^.)@E!#0KY(I,#F<QRAUG1
PLL<6-\/COFV)6R1E:P,E5/_\2>DUXVC4GJ&J6V9DP#"KJL*KSY1#5"MJU=5[J3+.
P^ZUJ$<#2.P\=3"Y7A2X3O/[;TA"ABU;RY!VW?5/[*&59,C4)G"[+QZC=W)(]P1P6
P;/Q\\4G6F$NHG'_;GX!&\L#+%/%R<%<#7>;!51D>Q%>&Y*Y%D2-*%\H,0>!(9QY=
P'4T'4&E,VT DGH?,)U%2W;[[';0Z;K=NTL1,?_4"%3#Z'#2 E[8S;1-UYG]@[>1M
PBCU8QAJ;!NEW-1#>#ZC_>U&IJ(U:)=(5?Y1 B)P9U,$2MY!NR['^?:[BKQ7N[J+%
P\W(;"!G2!J@D<@CR2NP.'F__K4N^HD7'76#\NT'7ZE $)HO\U;5%"6>:NM?-+*J<
PE@9H>H>*Q&JC/)Y((*TACY40-/6Z==_XTVK\"+:N$R*9KNQC?=?L204(^6&E#T.1
PNE%,U2"KDD''$IBT;\O>8ZJ)R*B UYPPE,XN*T14? M)TDS<EGR822L^'1V86B2%
P37<1, ^#.[\WE%RBJ'(V3?SY5^3&#'V6;GX<8MI3Q JQ/"C9]-M5D)E&>-_0>%U=
PN\,;9<UGPGI$]-[IQX0BST]A9)6",,2X-"6[5N=&%XR#'Q#/%Y4?]#?F^AP5_UY6
P9KHQ3YA'\$,_UX4=],_EU'%YI;VB/LE54DG<7-D-/P/$QL'U[JB N$^@/F8?/#K(
P0VG4Q(=-@&VKF&:+AD"(N SKV;36C0[GP]O+&?Q?%V2L$6B)&<(\IJOJV4&Y)4XB
P7%%W5()OET@88TMNM_4?^*OH+V<OTJ$9S)R '-;X 2?E_T^<'%CZ-B(Z!CQMT#S0
P%42UT5.WSOFW6'0@!JOA+X4Y[-JE.AI6CN@/A.A6,?80:93-1_ P)ZX^@D458%?N
PR7&-N3]MF+R4X2"3<@@8\WBF!>]1D/[]&U,FQ>V+97?:9'(]30L-A<R 65EB,P,"
P]Y2[16/"U@MF1YSACFDZ145$1N9 2^2O&FKM>:X,OL.LX,T%UN+R0FBV4*;B^U[\
P/$6C_&##'JV*R,:0/:,-!*=6)>U53>?W<)')XXDS%X4G+M350BR5P*N@TW4(+@4,
P&$ZM<S -X)TN7P,47Q+P;EN7>8"6.*]$I8$< ?IB5F"YBQP26U4)XLQ"5S$[!HR<
P'Z)5 CDW+7:2HHWGA=FSCSXCD$9)F;SW@2U$U'0@#HXZJ0(U )4*[HCD_ 2N-YLU
P;\/A*"'45!-JC7WW*WR>WG!,L &15Y!$\6B[^UWN5UH$'T+>,;N0U4G#%-R&DU\R
PZ_$6LTH---37JD ]6;-;A)U(">WP=M^?0,>H$BIKD#'?Z[AF:OA;@V7W-3P()/P"
P25A$MFXO+#>EO]4@&NW6E?,4]G>&2V4"6=C*X,#F\=(OIQ!GF3XG4>(PH<R8+-/2
P563+9^94 G3(_]6EI9Q.0ARGL.?IT=I@<\0@*>M\(PH!A"\L\W:Y*JFB@VS"DKXG
P>T,>($[<$6?+&;2-FB5[.1L8$808%?O\XD,>$V>G95%7J1M0CAO:37[ 0#F[?X2*
PJ'HD-$0:0H*)+AX(M\8)Q\2?$]<9)5R$@MW_(U<,AU,E4"N3S!)]"X@+J!G0 MKT
P0<KYN L9O4+D:0?0,2HF-,*GHTD+H[C>I097KXR/%K.G[PR7P/'U;V1S/B6/U3N>
P@:L0CUD,#@FS7;:CF-8]JHWB$J1YWH/R%@[W=KDZT[Z@NITSNFDY4"$BPBLYC(*8
PZ+FS$4=\Z:C?P^^9)EB0!A-"^_<ZWOD0/Z1874OS10>GFQAW-%C#N?'/=7B H.$2
PFT2']^Y_#^_]69,(D B#XI9EFYS^5G1D"6?,!T TT(^U,;[YB/X!GWMN3)T/-=D7
PZ]0L2,*/>YLX;;E>=:>P:K+U:CQ:6'U;LT6]'AP>[:_NH1"+F< ;]S0RIXHQ9S&H
P10!+5+[;SU3R8E-E@OFO.3!7B"@2W60DJ%E+_OB*_'D240TJ><G>EX_O!&HM6+JE
P=/T_4(68C"VP(1&?B94TZ1(@Q9!H?R.Y'"H/B#08K./O 3GR:I:381\?G_"ON3Q$
P#6(EUN)1LR2G3B "$C<!*A$N>B$!4C6()(@?K^9<Z5.*$T_&AZ55.J669#T4@H&:
P:QEMXC1$4\:B6_O>:N-JU.9M&\?W4B_^LG9Y7VO+J_1U9TLXHX)GYRTT  6@D@MU
PE5<:TZH3HF43$.5@A?J31%:00*Q ;#^BLP*ANK=*XTB4W-FK'L+# 7'45O\D5*6F
P _.E,3;$9E]PVU3K&X.\EI;:O@LA!BK3O-Z[B-<>;DM<VS #FDB&W1X:#O,:.&P 
PS:--(P:NY*9"TS\_MRM232;:"^^1S'[NIEHUD%8MO4W2P&P6OFA- *3B)OZU &A:
P>SR9@<@XC8V>GGSR,.)'L^?$/%Q,9"7?!LQ \EB!@?!T1$:CJMMP_9(SW'3E514S
PL[Z*%S;F3B2GSHUB-K.X"GY#9"';JJ2^'AHIB%:CA5[?'"V6*E@VDXU730-^V)7F
P8RU#F@W)<#-,4[;(\2>9Y+QFI]U@_S]#25SE-FP5VQ1M[=A'\M9U_^X_X&$&-ER@
POD=WH1-[3)7$.C-)TG/GY"X;]UPN0-V<"H?O?X;@*.&VZ,V^\9 L?,B/RTU7,X0:
PN25_S]X5J6+ /CT _ILT(,;!,=#M*NB3G6;S<[P&H'Q(KC6OR/4#;_-RJJ;@<I@<
PCC)A56_H^S)N$]XS2=WRHK(KC=1*!!PK[5QPL1_W72MQF<7\3KDJ=AR\ZGKSZ,]I
P]^.O*/E-99X1KA_G0.LV+Z8C S8M2XNN'6R(Y)"HKA4#XQ%!(=U&H**25!3MZ$#Z
P0%XQ$]$UC1KE9#AGG5E.,RK>W.^KJH0-1]<72=^!Y2FNH80&FD5ZL7BM!M+VI\Q2
PUJ54-7?>7J:'FI(ABV*YJ4Y8B2;,YKJ:5B/C-LD^-/CGR*9<44L;Q17%8WD!UHN.
PT\&;[EDW5SYP1KRD"XQ6/U,';AS"_W?"'Q&4[4"S_116V ;K)*Q6B.*I!)?SWZ\R
P79&HL=1Y"(&4V#X8,Z)J\7":,HG5+19B8KBQKW4W"@F%Z)1(.QPQU)>S4(0(,4U,
P!_;"A2Y/?^>7M;IWJJ(#[_,?&/'*0&2*FU@[7)4)N,4H@2B!9BW75)IW9]?,H&2O
P9]V+B[&/0>)]97WO\& ,[F)0.T'[;NT2&T$KUI 65-QCIL +FD:$EE2%Y:/4DCJ^
PQUC'+N_ "'M2-LDV5;UABF!KEZ.<& -!/N!5+P6V@R?UN%:V4([FH^0<!YL"9/Q[
P8!)FC8[L,?21EL?(X#RJTS"W@B:!;F1Z\CW>FBRR#=DT9IEP"79:<W*)%)Q(CO64
P@&4IB83<?KOC*S)A41Y"9]DUIDJUQ!N&RKVOI):W6;')^^:[\V!EO/ZD:<.S=XHE
PKS#SE@XDR(J5(]*9:GQ6V(O]7QHDEL0TF+?0/HOK10AZUBN=.$<0I7.IV:T]G.7$
P(&$)L0Q(/M*;2\!1X%T8_-=,AS :Y"G.+,O.GE[?VO216";QRU;O2=S#(M8:A<Z_
P-/^<[B(<1Y_C!3Q?IP69?'&'QC=]V7N^,<U!C$/_Y-T^RQV=,CVY)LP.._*7_!(P
P)CFD\LKH+XG)AA1>Y.<1DL18A%H2!)0VSEXB0QGZX?/#0#'J; ^$G8NK#W_#11FA
P*]);D&/Z":RO8D:B.?,\HU'?&;&-]]78(2?=H+F.G*@S,:;%NDS>R*]Z?,$V=04B
P2N9:<(XZAO_U@L7ACBZSK7F8@5[[2R$X=+=AS0?5R*3["&^=O(VPBEO_F)3PO]_T
PUOP73%12/%)O?$W_<P2NTJ4R$J*00@/ M<I&TA:BNHRUU[T'>(9]B(CS\4:<,>Y+
PT^3:W"G[0D@)>3$RA5P2M2QB2^G'ZF_8A3"DV%<G72\\UY_Y&TKIW!0N?,(;CI%Y
P'N]YA"83?BZ0H!3HAU:_#/H/6+IGM*<J0L'JUDD.#AAG_9;*3!+5TP8^J'ZKF8L1
P?4LAMQ&#3B&7Q!A!'/FOE"NAHP([KG\7'OCC,YQ&XJ#9./?9 6PN3":_)%CI@:9R
P<6AORK@)=LU!0; -L]^&IR)@.'\S;LCTC2R^(9)?^=!AM -Y-B:-RXL@F#,=TGW@
P\#!87Q6H$#<4#GM;$]Q\&2M\*<(&>F=6QZ2Q@HQ=X<?V7+I.P&/KESVB.<.5.0[\
PS!J3&O<)9FL<U5^O@D("WUQRG&=#Q.'\Z8P?QLH&]&H&6CI4N"?8WAX@*B<40W\T
PZ1U@BWFS_.^4-7;G]9\1.)UDM:8B8T)XP2CI\Z)0V5\=5OKR=0, ..[9,:#8TFQ5
P0-<?M-D;!'[G(@5AM?3>)Z;(\#XF?^(L4 1R$1QVEX!X' MFNB**,9PRC,1I\/J7
P%?$:]<$S#3'1W) :>PJ=V1?D0K(D"7'91+0GO20G1?O<8R =@G_Z91LI)OQ9P(T6
P>]& FWQ6?F\&$GVV>5^K4,YL(II8/U#M$8H\%B,V9RR%W_(RNV.J50&ZI:5@:R20
P10T&3=!?8A<H;J43D;V-\YZ@[R/Z2*O"Q-/";(&U#OP50"=^Z!#^%Y5V##BJS]%/
P>-F]T:8^P0J,'DW^#H'PQ8ETF^(?NJY=0P6U2ODQ %E;D@;,A001/2"87\LE.=A8
PW*RW=<9DH^0TV :=\J\JPW1*LE%@#EZ3K]DEL^YI;,3O<8INA"J,B:&B;!SQ"LA-
P_PI9@$M(LB)<^._ELK$X(99KW[CT1G57T^&/M^M?90X743:/#F22SN@ NSDX8,AJ
PH217U-F-:@7G0\GLS\),24)'H,4CS(]DH5I,.L#:A!5CZZ3]VD[1KJISV]V&0"7B
PIY4-@*5P^?GXX8^LV2R3#N?R]WQU-1#Z,^5_$$6H7VLX?D\)3"*-BN#,/)KJ=09Q
PE@\<ZR++P_D7_N,'W1.$M;MI3T#^K/^6;"!IO_<9^0?0V@-3&TJ 0GQ.A&X"ZF=S
PPCCHOV6RI6#2G1R^ZM[^R=?()!*_L<F6^8%9[:X.=;Y";)[GW@1(-_ZL4;H(]&LD
P-Y"T=N/G6/ QM1^B1VY1K>7 :K!4 -W%H<N:$6CC8V8,KY[?8-)S$F_6 0_6+ZLO
P>\TQ0^0SMJ&--R)%'-*#'94DSVD_J7IN(4NBD-MCNY_B3?@A^>[$; @RG4\7(F,0
PZ' %]T1E/G418$J[/G_Y=B'\":B:/Z6,3U9WA6'\E2WL =G;[7$9]9,/M#Y<,2'?
PQNQU)>D^_<71<G(;7[G*)4=5#E%(GU!^?WS([KO^[GZ?),"F?3-JO&F!'VQ90#HJ
PL8I)^ 934N2H8TDG/[Q]Z'7#7;#2D9J_ EC4*V@:Z0 8@<6W 7>B=R:7-&\!@6-I
P$!"?@U;F74I9*3FBE@0..!8ZM9(/][N4+H!I&V/ >??3:%A=_.9-5R4F(][?T5L_
P*7K0;D$#CD_4D5\ZZ+*.B-(QT,9$YW$QM1CF,3^M3CI^^?6[_J$, .0_Q?9B6I1\
PL*IGXSG59U]T--AQM>EW/X;Z)"H&G\=B9@N*&&[Y$PRREJ9\?>NG4)D1"-<_GRN#
P(Q-+;]^ N>DT'A&_Z@2.Q15[7Y2)$7(3TLM4H88*;.279[.W T1S(BSB$^FZ^7J?
PY#$,^0?K@Z9K[L=_R1*QZ(;.35\S6N2J>(8/#CL@%^0D#)%+Y*!=PT_L<;J.$0U2
P?A[UIZD(U4(I:4("G0Q._,.#=K!7#58KQ6W>?1\3Y/4OAD?HY#<ZG74O^:)/;SRF
PX?24+3G/5,F/]"22%RG!34368R-A:S Q09B4S3IR_K(8WE\ZF#>$TV1#4[\TPB?,
P@F*T/54[Z+\%JW%)5GW$/" 6H9(U%[)7?V47?-Q2!>^-!-&G![$-]4.Z;=2-!D9O
P_-]4D!89:3,MDAN-R@@'U8"?&7>"VU7&X#^3P4I!8XH..>#O+4@E-1489%C,N;K^
P)8UI*'5="/USE&YI(.]\F82'CO3"Z_G1UJ_]\P: ?A><9#1^W>,=>O^M%RYXG\.Q
P6^@J_8"^GWJZ$J;S*\32!1NBLHSG\HU(@)I]6+.P=<&_GDT#R?=6^FF5E7!YR6^_
P5<,G[IEE9R!MAT_7T!ZM%<U-*&S[WB4GRMG"*L]_/H2/;. T[B1#2(M1F7+S_)_W
P16JF,:*BD]]1*;^*MZ*/6KUCW_6<"!(Q"%%C*W(]09+G/P\@B+L.1'DF<%=BEM*B
PU!%<'_X?I[YT?C[J>HS,10XBKG)F /:DB; I8)P:+LYK]U4H$-=30B:@,\^DRZEE
PRC*&)&1S,G"]3_3)P2VC:5$01?MZC>B&Y;:YI.RN)CU>Z!6B,_N,*ZAL&+@:6"]O
P4K\]\ER*N?@'G<+KXDO_Z%+8\=W!6W.WQ&,AKYD1"P;3$T\V,@_P[MU>.DF_<@;R
PD*46YR/+YO"Y>I4]FF0$*H?EO8VD_N0\!(1Y*7W_IQY!][)D 1A0-:F;\S66(53O
PFZAT9].(7AOR&CZ;#]Z471QY90F_YE ALOY[EYG%(7(>AF9VA@F4PW3#(J\ 87< 
PDI.+9*/:-0185_LR3"#%(1)"I__(9K'M>JDOPAW8&[ODYBO0/ FZG3O]!.YR:BC9
P(=(MAO4-'C=MVJBOO!"X724[ACQ\)ZVT<2 JU_]C"+> *Y.[%Q^6__?RA@N]BC]$
PBY390#&M7<,C#5?)2JJ1?YHZI'G()")+78@JVVM@O'?4$O9:]__DLTIV?O4(PM\%
P"]DZ'-K;/4P;MN8AS01-++ #YG;'MDAC#BJFU=WA"O:VDQ><'2ETTPXBE+W6*G^]
P"HN,,\5,M IFY':O>R'NJ3'2RX@#B0H(O$'??>42P8BNX"T2:_B"*OU9W_D'T4V#
P0-R:T-^*?2^1L*;>\<<$KS8B()W--P0>'$[$+L6"E_0X!C]I3M6@$^6QAJO"_*C!
P3)'::K1D7.O6E5PY0?\FM=6QJN?@N-3U\*W\68_P$DJ"P@QSBAOG\L2LB&QO/%;T
PH1@9!] $L6@A 8:;Y_=R"68@.\^MTGWT#=S9< +8)IXZA"D)Y=*.O!I\060[DNS=
PH@5?Z;0.#5 T\%:>S!K/W(7/_V182UCC\C+$<0E:3C+*3#\ 5]G;C21\MD:^QS-X
P%Y -<J"F9D088,,,\67G3_QJ<J$>61@P\D]_LPN*MZC7B3ETJ#[<%K_*S8L%)]:P
PRM[X_UBTQ!,0&IP]T($"@SHQ$<\K[KV\QPK#9_P^X>><O HG*22I%%:TN'PK'#@V
PWT[1?L/W^;.#6>ZANXTB@DN/RJ_,9\>Y;]I+G-78>@UQ,-?CKXK!LF:N1=*[3=20
PP^DRL$*&Y/MWJ9=HYA%' \)X8E<01/%:1F_SR;9VR%LWZ0ESX-9_J%E)J[*R8WRP
PO+(K:HLXR+B"BLS*X":O[<2^,12?)/?K5;"[](LZ1Z8TE,@>JO54MZ%!8)M<=C8)
PA" Z4Q]R#>?H&#.YX>@YY1%%'BVA'S!GP$(,Q#UC<\8#6$TCS;/)'$/* VEA#!$^
P*D*+Q8Z2#%-@6E@06TG%.F@#V\<652,Q&LR#.=L:UV/W=DAM:7)6(VNM7G$N5A(A
P!!@717RHNC(W$WJGPJF9;4S\E=,C*9 @,AOU71*X6RWAK,B_%LLG?Q_R@P[ XK)K
P1EFY(/6O8-3PZ4O;X&_H[*BE.8S:[JR86;:\#,].UAZ&X95*EGQ1?P).C1D\VQJ$
P5M5Z6!+W50/4)Z+ZLS.<__/%514T*K+?I )IM&!@"I*SZ9WY$Q>1U:VRX@2HF_0.
PQI>*WUCM]@*9;X% 3U7W#J">0/?Z$4=#";L O5'[;*ARG!&+ >LO52%,?2'  L,>
P\DCM#%[3._Q<701>H^:G@S=!\)LA$)\HQE9>/U;[;SZ<D4*!6W)?"YO5-._<D'*7
PL>HEO,//P!"'683W3@WQ;$^4H4F4=[AN>;Q.RZ!6-4X77_$Y8ES*+RVAYMY7J3HU
P6(ZGFYX7Y:R=0!>M)8%[?L-HGG D5-P7\'#HI]DEV<R5W#HS[B<1FADQ_/#5A[%Q
P3<533*WUKV1^I\B_G,73?-##/!F:[SA;JB'$TJ/S^TU4C-;:\95(%0]KZA)5M_</
P=IJ*P.;R]3Q$U*(4QNNS2;L@I7(\:V$^ZH]%L9*N%2R3,5F<S>-96S6..:0+)"N<
P9[1@FU$8&EA7"IS"Y+/1:8D5(W HR&N?\Y9%C@\),_>[?E*/Y3?^*JAEPD1(U5JG
P"DL#,:OV-T(DST*@U_[#K--?%S$LO)E2&4J5UL_K9]R<P>JJ,MU:_%TG> \Z95%;
P7&2AOX@J,@)[W,%@AXRMV@D;Y:&)>$QHH$\P<0:XGFGJ,\.G7Y.TEKM:?-YG?3LR
PNR+BD08J?PE'7/T$?7J6/,C"Y6 XB.Z)HD)IZ<Z8I3'$Q7]L=5A-(W"2^7Q'3>9W
PB-6NH(O_@H#@?2($VD93QWB@('3*G_3#Z<A+(J3'4%#1$1H5A=1ZP2S5B:^NX"$#
P!I4L*4P[TH_=SVQ3L^@]':G8/AHCCR!#B-_@/C;,&0& //X>T)YTF@- Z:D<0%G_
P4-_/UJ3GL0&<71?1^:-3YQKQ6 (#7RH[N4V$E9#HN)J@*78&H+:KW/CPJ4VJ)^5<
P]H]@/KXJ4J8R_P9Y6%Q=(=%5J\Z ,5C#D8Z#%^')N'<.V=OA2000W8QQ-5E=HZ#+
P;3>T])OEZ.9E'(:A"*T(+,:/R/,3WX:7C[1-/[K%;& <.B"ZD"K.HX<#!!2.+Q"B
PM &@-NR6S]AGVG!3"1MS?4+$>(= QQ)H8Z6M1Q=3WS#+"J+"D%S(&VQZL#N#M;+[
P@/:KT-:#)^+A@.B@%?&OJPP!CAFA%]^7E2](PWXU&" TTL%1]<4&W =IH3[%F?$.
PK11!BP\=S[ H"!BIY#P4[Y&]);!;X'T&:#X/_&6UI[:FLTZ+TD<4'OSULH+2.\"'
PEB&I06+I\[O?];A'NE.4;/OQT($\9RT@"&Y@?@"2_:H0%HD2SD2*O>8',\$4!%6"
P2D'%[W) :U?R[6^''0EN43J?B@(P>QYB9FX5IV&K -6NSKN>!;"B2L>W)^=FGG]V
P$.NE%!D)/"!M_3)RNLCE=Q*ZQ>B_"6>Y$>74_)E5WARWRW[#8CL'&QF>Z,7NF7MG
P70<(F-A]%R\T^RUX0HPME!I#Y\.:04#JU."O*#KID=]K+]HM&<W,F.@DZ('=PPN@
PZ,27>OQF+'TR\YE@OMO!TN>Z/WCD]>ZF?"2->/^\*3VE G<IAPB_>2WKJ0]&[5F<
P:67Z9S=HXOYN/-8 V-:(Z@]JL,;S(0=(A10JLNG?B&I'OY1-L/E1RV%BM=TQJXN2
P@Y=M6X(Q*^B5>E_O:0'/35B!.O",,6-ID;Q ?P:X$TQ&L7?KKR8G[AF]DPF7!."Q
P@0*()W==@N$Q.Z;7T3\FSEU/JD0KNZ;6K1R8PDM!T^0QEVPI#1P (ONJ</R=B+E7
P-^DMB6N4'^ZR_T^W;N9;6T(*;B%8'W)[_7^57@NM7[Z*6I4#1M5CU60H"T-PL6HC
P%"!1I;"E0Z'_1>49E\Q L-7O#$$K_.F=5W@IWRITTCA,HXO4CE"))'((8G+#?>'^
PHOE!1-SDH*X+-E&85%\J-@H83H O?@RQ<!H*THHCPFV18A_\['*0MMPS7G* &@DM
PPW\6D47VV>Z+I($:+L!S0V1X,._&=IU@--^QJNK0( B#S4LBLE_&*1TI/9M-E, -
PQNN%!#R!-9.)0*\:=JV'NE@UK4O'"? ?4;:M<\Z\U[HISL2$.5OE?\=UOJZ59X=F
P%ZHSW+-NP Y(H%_3W,LVGX6N;M3D Q$TJ;!2WWHRXD;P1%?&"*"S,Q-XQ_>4*A5.
P_P/-$W+'&7M+08JX1>=0^1K8VL8B?$QK,Q:MI$^U&EAST1H2KI/8ZL['$VO$;7\]
P_X<_".=T@-)@_O'220*-S_?]E!Z7LJ%.:I4T-0__*5BZ P*S8LR]D)3B#^T@U=K*
P,:>\T$[GANS?)=BV=L]&4!W@U2(H!O4,_X8M^ 9_#6\_%P[G+1(<T#'MM97%F@4*
P[<[WFK*9I&, 8-6JTD12_&LCADG#R<:\%?1U@ 5 ?R&_;QB;IP>)%3%%DP@/1DYU
PHN:E&X2"WC7T>Z?L#G+P>S<!EKN/A8[?* T44?L<9\[4^AUX*RQ,45TU[=0B](=H
PP*#P*K/HK;!%8]$KK]K5ED!6]CF5EVC,&.G&(^IQFI&$!>;;U=W6I7*]K0V'Q);O
P9T*45Y8+M)>KEH7EZ;9BA]QN1RG5<+D4D*LK2;LEYX[]QV?,7QE7P_2@[25.$JAU
P=U3\'NU8:\&U@PAI%0B",3,)*5LPWG%NOP5]:&;IE1D%3,EADSJ ; 66F!'G'R M
P=<(E<#S#J!D<U\S'&&.K4]SKT-K<!;MEOL8A2OL:IO4SG+>=)K0^E=UNW2T6YSS)
P>%\3E6^'I \/B"TZO#,!DT<AO![94I7K@0?!BQ;"%]^CN<^I ,J5?) IBC-R\)5:
P$':_0359N;LEVOEMW2PEI3^,0IC+"#FW@;QJYE<7DD6G6P8=(J@;R'A%Q1O:\TL!
P(6UP@40B?WT2_U5SN8)$C9T-E'K<$)"V,O/-U0OB$78!C#^A]9TDXB50($II__$G
P>,&:TKGD8CQ@&^!D1TT-ES^)W @00WZ@X%4NQC<KL,.QPQ67:VPMD4NAXLFQ77F,
PF/*DJF<GI&0]=>).FYH;19&5GM*%/XZ><57MRQ=\7&R?\<)4+[?K(R699H[[$![<
P@J@/?*1UQC'.$Y-K#HN)=Z40A;=*1P##UYI$,_Q%:K;-;9,^)&P>L1<41(N3?,S1
P6.=@PT^F<HJQ_1!_?4&WR+384S;@9-P..^-',E*\NOMP5%AXK&YG@MV(@6R =K*L
P.,ZT^KK=E%^]*E-ZK<C =BF'IX*:\W^/ 3:#MNZ[;'+&K+=1([X)9LH2*LJE$T83
PML@$T>Y7DJ\FYQ'86QB2E3WRI/Y&%_4G/@KJE!FL[*S'?AR5Z:)R9GZ\6?/240EB
PS!R8F:UXD9#[\56609P5K?3(7$&!83U%]+11B&9(G0@J6BQY Y2!M'YQ'PJ5,2^W
PW4,*Y ]DI'$:3*'2LIOL3DNZPWOQ2,9SFX#"8\_NWK\_]/YS]$!S@VR5VX"M[Y7G
PX5''?;8 -CZ8+AV:H\O"\MQBPLUN1#F88L83FR7WV^?SC[Z$G+731D@T49 >T$<X
P/;!%XVU 0IIWTMX;B&^)2E=&^M0'NOS-&5*.>IZ&+3DX)PP&ZUV05Q<Q^Q=(D079
PKOU+ILC[UR>3=/!3RB$Z2P/5 77R@ZA",:YY<%<:#576)P%U+2SMVZ.]RGN5>5UP
P9[>,57]@A,<*?0,5@JK&XR0RNVJO'5?3)=0P_':P-^>KQ'H5C#>%&BFEMZR( UQ+
P?KERJU8NWACH4GV(K;K%]]X(\P/ P(H#7+,K+H=]^#_@S-I!R8YB5Q/YGUH+?;D+
P79BV8Y1 4% 3]=%K5_IMYU</N-,CYR1-7D>^(-5W77BKKIUI>^1JJYTU+/_*3W-T
P^S6-. -A9>:OZ:IZMZ$?W:)5S;W'.R"7C_"NU'KFV_E?&&DJONF[J6TZ^%R\+5T1
P>05Z$$NW/?<(!4%E@[.5R&L4VP1=G)O>O?<S!T.F8[%M!'V6P02<0?C'_,CR1>HK
P;"A_2"C3'<)*OU1@-5"$V^V%ZW4,T>K#1JF^FX:_S@)DI(,\#6;2]7$IV$7#G<"4
PU\UBWN;+3+F/*.F9S<CF\<-G#M2* V'L*716KZI&#('\>$[0D(@SLA/+JW2FTZ8E
P3,2 N%2FB;[^3H)YWR4EY\@)^*+=,^.1#Z/''&DYR4)(8[=>+&>-!=7F(,WSN:WM
P!E+Y!%2=N3_^QSH:*4O,"8]NU-)Z-U/E.'^\$1'=L-_(8#PLE^WN8C$.E'@]S<#>
P(>G7JN&">'$DV-"XBDRX16'M@2=I_M>CW'#"<Q5#83Q(8U]AV(QPX(-28K+_6!]-
PW!YJ9>Q] B[(\<Y_7%Q7XS6HB:[A&/B%/L+4K]=Y7B2)$_KAF;"7U;P@FD[6RS"Z
P$N_CRKE#*1I0KI5S71+!7_[J55R=K!)^TN+\]N1+/OZ?4Q7\:OMX07H-'@_2"WS%
PWJ]G9?!R^^FC3B[ZAA;7@>QU*$E 4CH&P41FQ<S>%7YO"+=%9QAHL54(FAA>*+,8
P&5 V)V@FQ4#:[0HX0.:JC!VI'PUNS?2T=&J.,LBNO8&&9&K"*R&@_/%PB@NLY<7G
P+I<A2(3EC [AOR>0H0;<_M\L^T;DU?]:AZG?DGU3@,<U[^ =/W% ?5N[L0(\F3$?
P7#1-'#]N@-\DH(MV8/.=!>&M:=[(0TV;(1/.E55/\G.UI037X)UTJ_F5[>]TSVL[
P/5"V@2G0(?,1<B:"0%T.^LTTH9A!EMCI(?TK4&%#E%]/^X01K+?J2$!0L@%8P3[P
PDN/[8?Y^NJ&6A.I5_G@T3CT_T^[Y%R'QZ_]6#@7%S<RIOL02Z'O_"NO&"D=4])F&
PZAP$AR^3NY@[8RX+FN(MX10-]P!SBZ%/G508.>$OI$(-6(-J0#<7P#K;*#G\1$X4
P\+SQ5K$@D/N:O$FJB*JB&6:0TXXITT2<C ABP"^[0Y82Q.G=@[F[0):_;@\?O-)[
P-ID)4-)C15.-S^ "*9#Q[=[H%YOM-O7-J4#KDB4OMH:+9%TY><.30PK#8;/K!8?E
P]$V34J=WLIK2V'+FL6RH).$Z-2/OB+S#SGSK;>[/+9/KJU WDBU]<%;BQJ7DO [J
P6=*,J[P]8D(#'48A)X#>AMB(S]0#?.73U1L5"NF>4\DS R=@DZN<=OCSI\ED],[,
P.O2KI=3-3*0"*SOZ6US%^PTI'(%\2XE&Q$0O>RY,?AB"VB[51+NJ.3W"G@'M/P+/
P@?V6?4TJE;DC$J'#V@3 TV:0XXI8).:Q9;SEUK=0.XFAIVIG'>D<W:ZCRV);(54 
PVO/4O6,K,AV0N+4R7]PC'KOU3-3C]=O'6;OU$2[QX0\.0 R43(!B>CB,Y'1_TG>(
P2O1)RQ=.3.?!!&Q"N_H!G].XG^EYK*0KPERF0D7T*YG@NC\%7Q4J.*=O@BASBK Y
P*L+XUYR#Z#*Y(R^NY"[" J:!W37$]=L]&P\ -*!<ND-9WE;HK!M]/C)!R13.X:W,
P1E@+?3T2TR01CHWC)F:+[*;*B'^I$5NMVC-O\3F^!K$G>EPUAY^;^M%; U(V(_=&
PF12JW[EN]*55^?7&,6ZG>]/HE=<U,8= [EU>%>N/W7<D<E\[@^'P6DOBOB[RW\2X
P@VI!R3#4Y5 @MNUT_%'U+!<38J&41K,]IS3J^97[.KRVL')718PDU)N\H!O0Y]!2
P!-!@4E'57DR&]K3-L0*O[XLW$-#)T?=;ZXB3(D1D(TPOQ=T_AE:L 8]79=M:XZV"
P](?).G5[(.6P]\G>VA(CJGC2I<_.[[ZF=_(7AB_FF@51SU;U3&<AZ9^LKJ'5/T+U
P4MUJF+9$S\9"=4@@5!DQ+!QJY&3!7L09[(H\X&8]!6C92?_^FEX;2$E3?D;]<OP6
P+/I,+C\]GN;Q].TT"ERDHQO:%E-_<HBL5K T%?G?7AH3XT]"=50U\@ [M99?2>*=
PV2C_T6^],58S&OT":^205.D2QB$>OBT4C%%,7F#<LW9.I54SQ9=U&F+"%]&P/%[9
P1[AU9MQ6H97*J;(>V #O0NR 6S+&- >4Y].Q?3;*TDOE2(0CK<!D*9-&/=Y0)?*_
P(&XWH%]&M1$"\HZD*<9T^6":<*U*>?MKT.Z/I5:+%-98-@$1NE:4M!*/V"FBD<Z9
P.'ZYR/A6)@W0"AIR*!3=<) A49F+6G5!CN$!OCR"9_0WVPLQ79); \$+BC)GJ@2R
PX_P!CN>\%_^6I_O2@Y?;"J]Z/Y)RDCT/3Z8L%7(&OKX]#44+[/:@= F6AO1R?Z':
PT(IE[ >5O+*JP$,8:;3C;A,,$Y5J3?T.Y #B-O OZ4!,E;<AS2Z H_VJZ,5+&AP\
PVC*D>#.JBG24?>"4GCTP!JI*R\>]$:Y,B)6]+&HFI2,[I*&G9[XY=9QWF2?="*W:
P7NV(0NP%/\P(S)-D1GN^_.R_S7 !F /+_>D.'"4E))$CT(@D,CQ=W0GQ[36/9<N6
PG8O\^L<*.MX 7=WKFQ$I":?H.8_R-,C&-R'GC)AI&N;%V :]$C^7)^<W,"L"@L&5
P3Y0?,DY=8#';UY?V/Y(0I$<N%C]TY)[*';6DU+JN09'[1M"J@\0:%8PXXF>(FSU[
PS""(S!W&*I?<9SK'>D.V><'+JK1-8>NF7M7,IYN,7&:T@3HX:Z."E9AOXIO)WM;1
P_'!7-CH"O*2D AF8O7>;4W?OM[CSB":S?\Y)M E;LZC(^W@[)OZ:P7+Y "B]_ Q_
P&1]-0[,ZD$)<ZM@/46DG=VW/X)V $]V'DIC^/FY02LAN[!L#2P,#NOAQ*B4U2]7?
PT%=+I4 *.T9!X['4SBAX,I'5<#X)Q2N]4,084MVU'/+08&1 "-Q(EBB.BBN/B;C5
P]:Y:) <DHQ(55DZ0J;$VM6DSV>P71>T8Y_4E=A0I?4V"CE66 24H)SPA*:#&3N1[
P"DLPVR%_?:,U_&S*B;N<[O!G1Y;(W@&'3UC*M,&C@)7T\2G*$_C[/)ET*M>ES^Y:
P0W[XH5FLVCWTX8S*^"Q[^ 6XX:$D6\.IZ^Y*E;'8<V/+S'WJM]9VH/HF9NBOK6<;
P/@Y1!F!KK_JIBX>/>X4Y#0U CBE0DRG@S6"9@GQ(@6/BXQU1L;.SS2/(3VLRY%CQ
PMW<[F/9]?5W4$,(*,@OG,XQ]KI7NU$&(, ;KB_]C3[HRZ1C-J<G;<ND@'5#@ <T=
PWLC7EN"44Q>/:+I-AA C]+) G:2_I:>J$DCG\K,[QU;^AX'((1'WFU.D"%!B2,I6
P66!8<FUEYK&R^V7BDZ3Z%K=3OPW5DB&H5%RX^RGNGBYW2K>QJM8?#%0&-;P!E^&0
PNGZND-?>064P0TE95VL?O[643BV&B)@8"Q"WF_6X(W.\:7^XEM$"(*J5J&0G?;LX
PXR97_:GCKB[C*RR/5A2_MN:1K+4!X4<@SVOIF 9<]NB/.%/S_P UYN(@]XS.H!%D
P)HDKA71/Y 35?^:)A#@%['?$=T>-GU[-8K3RB<?;O#EK*.N@_I,>[IH?DHBH9!1U
P661*/@AV9,/3P6JVG[)RC=Y3RD^X.0H8'(#R4+LBN!)G*^1<COS06+J!(CK$OFP%
P)=G&,X'$#QG>W)S/TS\BS$CF[ZN.#6WE!&\L %DNTV7HA]]W?="U)+F=93I M#XW
P:^SM5GN.$8J4-Q W*L>/2T:N8\$*>J+M=Z.@#Y%PO"B,:RM0P+3M;H.9_53KLZ(*
P99.T,EPO_<N.P:(>T(6^@VO7!WKW&P-6T#+U !YT\Z'DNG,R]>LL5^;G;]WM<#FE
P7OML+?5]4D+>DI([B0UDT56H'PLYU*CBHQUR3GLFD"@%T@#**3T?.<A]?32;8@0:
P*HN[9GD=D.EA>UI7IXTXZ"C5MLB\VE$(\A<_:<=)UA%E(:>!.[6(YXYFV3MMN<0%
PD:&?"[:)I:/1QJQFIC^0/*ES1F/7+\>-R2!2'UMO:O;+5DLQQ.4N,0XVQ!XNV<K.
PH5K/DA_=!SD%T+;BHA6O9\%:\@UC)',@AC+F+&KB3=.E:D5/;W(.)<O:[(P<B$UZ
PZ2'#VCMVS))\*#M0:[V=FLU=ZD#7#,@Q^;28"97ADL21U](=RL[6>N4TRJ:XR$??
P6]H-*16\8$$.AIVA,(:%DFJ>4#W04KY95:65:!<0+&SGDFNW:,KXXH"S^>%+=Y#/
P7P[=5ST%]F]:NO4I,JT^+]2KA&>F M;J\/- =^[-N<5A276.Q.9CTZA5^]<ZNB);
P^*0N[0C#>-HVRTSR1?>LPHZ_,+4PBI1(%$G+FF1O$NF#&2$K7<NA@H]P>TT9HU6D
P2'<0+_?;N@,MK"A2R*S43RR,0-X)2'WQ=GB3AF7(-@0!VOLR\[YC8JCQ QZAU'8'
PFYQN5*X*D:EGX")DS22+W>]KL^G*2L&G30^$AY<AO2V$']S^6UO4AS8,N$//XGTE
P4..V/R=RYM=X[,6&.BM()O^=.==/%*SX&BJ1@EW\/&UI4= $SO1;##_+P[E)66 8
P*=FA?"7CV,*M/RN^HV?4^+]@N'!.C!(WQ+WB+&5DN8#4*("X$#LB=-4TP&G!(JD_
P3 D$+&8-S1+"R953:RU?B$%'E1FW^4SG:KHHENLK%F^E=<R6R 4/^>Y6Z76?.>Q/
P;>X;ON8F"K%WNLNF<*;3D\:#5P;N\Y_J?LQ<JT;P"07XIO%E#0\5\*,RHAG #25H
P1J5/]? !&Q=J^*74P[MVB]&;F87N3YJ5^KLR'ZCDNOD49%X.7^_D;0N;BZPT"QS<
P@PL3M<\]&S65,:\="7S87R(-X%N6SR0(@V3N<%]TEYY4C!MX%5\<C<S'#MMI2E^ 
PHX=8Y+VK8OWC&E OTE_=G*?:WT&IOW/".M"V?#U;ZN.WNR0P&HY37V-A3IZ?(QY2
P&$?!KQDY-R^+#5OCYSV! FLM$0VQ\A 5%-X$(*3'48JS)0$KP/4B'V*6NB0\':_/
P)%7^%&B=.I-JPI* ;KYA; ($RCBRY7&D=:L_Z@\O/^/]3%A)IP3%I.NL@L0XW6LV
PF!@W+/=E*648&7-\CI]_8KCPTMJ4#:]-?-H7\"P?\EM#[6XOVN9/A$ZKVR]\S<Q>
PQXW$:6&X8>^AK3#TZA_(Q\[KKSOY2F]GW(+1D\%@;1 ;I-X3@,0]B<;56W&&K"[Z
PGX8[O[-6RT<K?TWQVH^)(B@/28)S.*<UL)Z:CU:UG.\(Y1N"KN7#U'AY]Y"XL":6
P(#06YHAES&L.HA R)'C]$XQ;G="H(DTH4O'Y ?J7*"*^Z^'HS\3"FH$-D<<$FS0V
PX@/40>JA<(!N-,]P/=8?V(I.T\##;?6/.E=A9(O:Z1)T]*_,CK-X2^E3(*R'.\1J
P!#-&+)B2)M" D&YIXS1.;$:]Z8I'P#H[6%H)@*_@ RUA@+K)D.^!,IL;"7L ,V-<
PL;^*9IO^(Q%LV\#^J;(R9@M/%V8D>RMS^%N'&VV!F&AQ_\/A! >^-+KS:A&;MDUH
P8:'_+N])+[C+&5),FQG:J'_"W1I,NDUH)4G2L';. N9TV\&,P(>L?$6E/\^YUN(6
P0(R:P;_\M+B!DF>.8_PP,U][U-G]7.EL2.KDYFCZ-/OD'3PXZYP59K@W26]H4^J[
PA.GU94[$294NX .9!E=-T&CQFXJC-7B/2ZG(VFK9$NJ !>]#9ZQ/^Y\S>'?$6TX/
P/H7+6O[H*$DKV "L8&AQB 2\)W*B;H'F#CGL29"E=A,*1'P\-3Y!O_^CXC$SVB<E
P\R/C"JIS/[&=*;TXW;^ [":PU1SI.O5N/^RCRLJ@G\\;;#CDZG9750TY'T4+09M)
P[0>JP@:UEUHX3E,'&Y]WV=7OO-FH*\'<%_;([96?UJ40JD?VQMLUE\>38!>+%R^G
P[Z39+SP\HHI3(RO@PZI<5.$A7]X&*H7:!W4A(Z:QC/6>F-S;Y-;M.;_ /%].FWH>
P'A Q[4 D3"3(O?0]AS*Y9.FQ#-<XSG=.4+ O&Y$R87/QE!!H-+>VJE>M6HX682\V
P*M7<;[:+R1N=B8#[BZ8A4Z/_K4&P"Y.E/&H@NM^^+X7-6&0P3U1!L<265,*B%[<O
PPCB$#<BYQE5(_4L9(S0Q.P%:S-L/^4G;PT@OL&E4S1 WL':,=ITYI[+"O<\U&4M2
P7AK$B-3FC,8<MMUW/6UQC[,/7?E3899/!01+< F0+J0I\QS3^D\0>5,8-\AX-/^6
P&/0%Z+L45%Q$1-S3HHRB&_Q/:R:=T,*1DC"^R5A4@.MI4-Y,#43[;$C3XVB\X+#V
PCL'W-58[U%CVL:=A)9,;N=[)8:KN_;4_G=>[="B;3.$6ARD0TF#]GZ0]CY:QT2+$
P=Z356CW\A%5O/<Q98&U20) F39W%'"P:*M8A:U-G'N#8R,,K1+I_^R7QEJ]LEJ>Y
P7[ '.^^,JL_7D-T[>=&VY7PV[Q/EQQIJ_T-!YW !())==6O7**<N_ZD>6$ODA.E'
P0>633LYEX%R%-SY&X=1<KG[<'GT8L?YA2:;5UQ;1I%B@<C2/L"F9%)ZOYEK+R<PL
P8N0(AG?+V=]I1DA*IS></NYBG$Y9$NE:%NJIV\5"E07I@%J_2(<_=7R#D\NZ%@TR
PG!4=^>/I_&$.Z^L:PS7$:!H[UR<=0%B-,NQ49R+?]71R6'C)9TA"('7.C!A>(!8Z
PU&#8#5HAEUI"@V_%6RUE+S'\P3L4W>&C/;_8J10IT>^3;R.:RZ/-U2=>M@ 2'^4[
PH2-P[)@CW-2U+(X7?>[_D^C>.,:%&Z[[YFZ1GLUEFCTX&>TAK)U:@L>!"4'5;43 
PW.DGQY'-Z 9Y?B>M_@1MW3]N;HY#8^-Z6,MJ!T*.+!:YR+++@+\2%X G/PA-B1J^
PP0(N!]-V!0":L--*$A:YYD]M?0(C7X'ABV/<%$60/Q^5L$OK"5XX:7BH<BFZ%R]C
PB1&!]"F3D5X47Y*L3V^L7P4Y>73$DZXLY:D#*DG!GJ 86_DE;5(@5Q0!$UJ)M/N%
P3FVV)F"0?@>S4LORS/?YQF65>S2!S!:+XU,7K13K:' (I@Y%@0%6?+T"AP]+?Y45
PONRSTT.N!FL$Z$DZ?432"<;5E)!VJ.MA%#P6V(Q]669YJZT,=>/6WR/FV:X,8>2%
P<!89T(;KFD,$\"9@PQ6N@&U_%[UOL:-I7!B0J'K,9-V5>6QBG*DCJ7*1>FH8%L5R
PB3KAA!_I2R/= 4]57R: PM*#Q60[4ML-ZD@SC+6$5INJ*!_V 8FSA/6PF*;4,&?A
P(EPE*S2>VBV[\0&&F=',E5BE8F+1C-.37X'D*XGTK0(4BL+KI1;8!T*X;KW5,1FH
P@Y;+*;O#J]8OX"GV!CDQ501],%GX#:+\R.FL2.?1,GQYTO0/51A]JI9V.. \U#B=
P0&BR\>7Y )B,6-]*4(.-_WP]#)!>&*.Y: 2).^=<> >-:0WTM6SW0SL0 O3WJK^4
PG6I*1H"+/.[LVN'E=BT+40GL*EJE+/<7_D=U YKGT[PP&YIQT^;<_OV88$)^;\8J
P:@"64V0L0=F^;D"_36)B5H9]B>)W<R6M@>V9(I)(I/J_L6@1#EW)08*&6)#BK;AJ
P1/90&_<2YU'1)-!SGQ+T="V.KFH_:B:Q=6,D?4T"FDM[O(4M:.5KK*WWS%JD($3/
PF+C?^B@A%TM*Y'& T?S4#I2$I$'OCQV;!$=)*-TT<;(AH![)!Q$/ZCF\0@;I*G&W
P5L\I'  JM6W77]S,)6Q-PN(CV8-PM<AA$,EXC%IS*6M!U\E\$RT;/@GDW1= PNW?
PF<.MK'[B?OTY*G^H_@PKS7]$D_:C\,!J3U/A,ML<0&P0UL:*K21W,453H$QC#6.;
PG;B'KI*)@_"VLBHJQY?U&F,MX4^@+@;9,U:.%Y(76));<^J"TVO#*GUM> C6R>V+
P#C9[+]<ZPR'95OQ;,0_. =V7=[_7FW/\79YK^AB!X/\5J6:Y1FO$\BP Z>O8R]J^
P:Z?6TI)GH,LILY%9:RX\3N>O_3B9-L&4N0WN!'*1MW9H6YE)JJCJR&-EE>''>I];
P916"#$C(SL90!NK$'LF6 <<>TSZNY#@)#U/QR[8&"KM3\I%QV+8Y>PE QZ-JX-2A
P= :A"%O>PF=>24>BSKT8J"QUHC%1<2)%;K=(K'[H7MG6[./D>6QKN5^?B5=;W]!W
P2:NVV!E(*E\0AF%9U*BS>TRI%^S'J8H0X69/S42T]$];NR2ADWA3.@_H/?,/0J]<
POPP;3K>?+W = V%OZ:'"F.Y.*"/V =)1[,@B.MAT(QA?C37IP:5C@0>;TPC\$2R!
PM\X[),NCXUY2[A >.34BA5.TC1?2"Q8']^N-5GE-QFKV/;E6V[[/EV(9%"Z#M4QF
PL&3 >-]R9RQRG&YJ#FIWZHN'#-P=?@?@_$4)6J-ZS*D;@%\"\7.Y571&F@-6LFX(
PCTD6,^C4YS8_4PR[?J*WL=2(/;B0#V\N]3")'8*.N0>W!9;D[G^D)!:DELF-5L::
P\+3Q=9<KF?A:_A(+*;?AU[#P<..?[W@J3A&2&G?J;C;6LJZ8Q7*MN(V0+.S;-Q>?
PFR..9V%YV>'A680!>W@X($&[0P2C57@@H[<W@$+'P;_(=2QM* ; P$:B%(:B5@8)
PELUD(0!W!P]G_)AM =16,(W ?WMGX%2OH8,L]@DNYTIW<;"D@3WHT90S"+:Q"X[N
P;Z-,RH=.?V>8^B^7)#U;+K;0 ^65$LQ"_O>]%N7NX3H%_PE3)*_8=08P,NT9YKAH
PE1@>WF(KQ\:S%121<8R.IR"@_S5X0A3Q2]^'*0P^J&,7JBB<[4TIQ<7R<VFY^JWP
P3?.%AZX,B;U8J=Z@<?/ \/S3Z&,*]T_@N*:5,19>[CM@&_U;13=G+,.60TDF*3%!
P$I,,((^A0G3"P?[MC798[D!2P'114>"O-;(FFQ&ZV#RQ.N]*C&V.GC9.L*AU9BX0
P?_AMBZ(_L:IA?Q\,Y2.DM^(AEJ#7_LL+M<<3787)KRJDAIVK!$US@0P<0I2%M,':
PKX(Q8PBI$2B!;H)(*J9GYC-DN>V=X9GO=K,M&9ZGZ-78>NYEP#J&HES@9)>S;!ST
PIU[HT]*$FKSV)73A^[VX[4;9U1"PW8!'1$[VC(*WJI!58)GH!9U+X_X#,[0!0C=#
P JB]TTP"=YKSU)PQB\LB"\L;C4#P3PM Z"ACPR1)+T499SUT=&+*1@TY_:C0&37\
PX6/FB(BY- 0G,,\J$256N:\-SB7VEN]JC.L>+DQ+MLSI\%<@M<G49Z^YD%3OU\PM
PO'*Q DJV);[K3A$#E+77\9,&J-=X7>1YR?;&#V1?>?Y7T9=2,\!_7 X+#3.+KI2M
P+)\6^F\:R) V?!>O!QR\GS7&(05S!G4W'FHW6XHY"PVW<6)._ ;8%$#EL0L218S+
P=.VU?!Y A:XTS7[4)]%T;HK%UQ#NX4<>CKL4XD_" 1R@!BS#B0RVR!8V]+:6_0UI
PAZZ=7W'X[?&DO,#'9R)OD7;8AR];T1%*E=H>\3*[3TF>!T(61%<2;M*O-DX^*H>1
P'X%+9BU<"+!/![VSH-^QP-*8\J1=?OT2L1'S2P$N% [8;,W;N9E&]:39W@DQ_JD_
P_L4OQI$05;<//;%RJ8A08PG,=?)MD00GW5*9SLJ ('UG%RVYWNM%4:E:2HQ+KPQ6
P@MZ,8O0:EAV 0/<G2==.:!UR91"P0LER"(G/QA?X< (M _Q+&]I@5[Q(A=I<6L)=
P++@9^F0HAZ4UD]R&=Y*Z923Q&$?];"*?Y,[2\B28MDA++I2BY$'?,'1C_<Y'J_^&
PVAQ'G/(&+HWCE-/J&I0(JB&<&%<0T.\-;A'OJE8:DU,W%WHR.6%>SB6:;.8I?*>J
PN^JZ/+52LS96T<O7=8Q/1]*"2CAIUJ6B\46=;YJHD S:!@SX N[TQ=E1]Z'V6%L_
PIN<#MM"&#IN/U9Z"RJ*''"S@)D@&$KZ@A8M^HR7Y(#KIN2H7IIA\C;](QM)262J>
PFQPEYU&C#^&UL(4! #[CU4-X8A#STY%8IJ_9S9\_0.W[PXZT7;!K#55"78E"(,]G
P*BD[F5B(S$X1L-.,[@JC#=+%(E=R%*)M,]B92*>,<-+2"^.6$TZSYZ5+D/Z$E@RE
P5/];WJ]+%RM*VPM@"XC?B(4E),)2ZT,YWE-*:T+F6[.NT&FIS<M7D_2N90H^^HL=
PBI:LZT_1C?'4YF=^I</YT/@+^/E/%,M$1"/"<"2!LF*\'4!3U($JELT:;!G,!0<A
PKHP2@Y?K'4>H$##]+#^>_BIY,2%(_'MY>@U1&Q@]-7%/,A\)\J]$!_CM)Z+4GV9?
P2V!'*+T3]K3AY ]YHO^..'4A3\ C8?2&!N5"43+*-!I"0US S[&KO/+C!N164/'>
P @PW\>AY-2PND5UTT)2I"S<K@9+D>6L+-. WW/&!$E]AC*L< @>W:==; TY_,46R
PD</3RG_)&[=BMH)7>GHW]KYZ_HAP+!2(8$F.4KAA<KT4^*)O8PZA55?OQ^ZS#S8)
PEF(H;=%@(H<HLB4K$:T%,)=8*N[L!\C<LV/TSSV6@3^NU2/^JC^YXEH$-(Q:;T_/
P%89D0R<Q^)V@$@+?JGV\=\^VH3[C3NZ'FVN2>DVA3+.!.A@F_D>N$?[ U);=T8<+
P+,RJ %>=9YK_?MH%L]F8'RPBJQE,D:NM12K_KBN)7-SWPYHL&I;;[P\;'8[LU:1#
P[*??*7A)<$)\]M?7PY6_<2(FR8*^66&)769"%:@1K[<'AM.]^'05%[@R1JLV9CK?
PURSM^7D'7B@A8R/ZP2T?U)K>,#=^7'8%(=S]/-,"W2V;6_WDTRAGQP"5MNV$#JV8
P'[OY'P#7NT!D*?!MR6LMX&?45Q/B:0V[Q8"?QQL?"'<L!KG2G>(K UPROK];5[M\
PZ'P.U1:@A]C)XL"IQF@U'UH02P8;W3"5ZT'HE B;76FLU9ZQ.G6IIP=U# IM>O+9
PU79X? CFC,@QL[>+/N1@,_;MR1E%&X4^I93&9]:OK;HV:!\7T&'C;3Q92S_\3;:E
PXG%)K?9_C?  @6=+F-+L5L 2W'W61E(L:N?>7O64IK9J,<74E2=J),'ONF:QMP&]
P*78X="SYS,22_I>3;BI.'5&Y$R 3,.A \4$/Z*/"'@*V/=M0%RP(/3[R&QOS$$&F
P.T+4\>>!P::5.F<[:W6PY_8RJ4S+!*U+YVLWP+I-/YV<,\/D;)_:!85DK-Y!]C>H
PFWHMG5V71 8YREU>WE%3K$MS49E9A:#]OUN# Y^]:J%]27$Y[[]:-$\.UKS,]@50
P>], .#I"=4%F)(HZLRA/ O41!4>46>DM 4@ELSE>22W)Q5"1Z%)^QQ<YJ__TNAR0
PRI"S^EH%;J47[0.\1V@^7:(PH+/1%,\EAE]EU]T_A[:\QN%1VUO;,(I,?-.I&,V\
PO7F'_.ZIKZS AX0+R?VN)G'W-8W+EP.ME*9($E9 %YU47F&M2AJ6J+ 4+"U&0?7S
PR(ZQ=$'T@#29DO0:MP][TVTFZ,H%$!WG3)O\,4-J3!:1Z U*0^F29':8'R[ ILZQ
PM9 $\XS4!-ACP*R64U"M\"$7!"!3E7*T"?.2K%9U1 K/A&WP6S909&M"W@Y2I4AX
P#I9T<3#<L,W N0\(QC[7+$K-EVOLT8<5]_G"R0!ME?  '4C<N6K &FG<T)'K?J!R
PFJ94(*((NQM$+QH:KA$KP^QJA5P2&C"[U"0]1B\_>QM>V1PB(NR.91\T <Q(YTUA
PRI&6HK.[5KI-/)V-T [#3 +[-AJ/KAV8D";I:8A,T2]]9O?(-_!GT  \RY??;5MI
P&$7K;:(<AK#D"R%5JC%#JM.,Z/F]T%J%@>=ZX*@AH_R.'J,'/["F:\A=-'29+9."
PPX$^@Y(ZSTZJU2]E4"2;%LM,H%?"6997@FY ]N2>Q^_F0BB)'LE];I <#WB^B4=>
PLOQY+.@2N@W5Y?<B%P"-T8"$#^8 WE7=LBT:'+KBKD."8NV#JO& #]MUAJP8M<@G
PV6C'+WT(CF2.K!,-F,=['%.^FD*('7D4VL9;SR2WK_8:P^ALT)(YRH_TU%!!OY9:
P209A!,%1^+GB*>YG8(&9.'&C$!"K+XL)?G&I8,7K.*,OR+?)@E 8A=0%V1KCW>+>
P4K';*V?)314D3D(='_VL01((K3[78K;U^RV?L9(2,\M5ARGJZ?Z@?(J!;%S^%(Q6
P7\NF_E65;6E-X%PGL'+IH?ZY;"5(*Q!&!,7[4*XC!,[+2PC&7'.I?H&<?.>"C^]4
P:VXY>!Z#Z'AP5LEAUBEJ7&9M%Q3LOC5$K HO_53%1T&E%PA1XZCF,E?#B[39H_^V
P7CN"BC98%L-.Z]><B2=0@IP:G,0BR*DO@ K"KJVX?C#:PM&F/Y:WXV34Y$)NCS?'
P/PKPNV3H>(1//&WPIN\8'A7;\A9:AND8?ZHNELWS,J!0CJ#C8DP2L&Z!0:G8I5$*
P8\"4B[(!S(^RC&@4YF?1L13A;CLNW^-^Z;1/'7R.A'&__.YC7*89&>W5 3]9NV5'
P*-O'6;K5A'$,6]*_$5R>&5ZY]MMIVQD][4FB_QNWY33F?9Z.S9TH[T3GVO\<RM:<
P:BR3-XDYC1/G0G];=ZR$%GM;*D[BL8E;ZD_G&>\<K%VW<PRO H#.LZR? N=DA\=?
PK$6IZ=-=SP,"C,FN%QY9=N-RY>MH8BA<FA.YH.S[5>2)B[)JG#-L585Q0V7<VJ7H
PJD[X3Y05^U5$6(#L7<RF.6^NX^2S8!_!L_.Z@\97J;:.3089OBBM_0>[]CV#JB(3
P^$ 1BNR'J[BYW3[4^T&2XV5:QVDV+,Q,(?8X7QW/KY"[<,64.@.I*6G*\Y2*].8<
P%*AFE/*>$J?=):5356O&LM"U&L/S:,X/6HTJY<_3=^\)P#+655$Q:1='6(R>0;95
PSG8!^F)E^S8R:E."  QSU/E%MA12RRP#&*M'K"2%Y*\]KKM+*@NJ$ZLGA \E?\<\
P":,60$_CE+GOFE(&YCQ848K=Y$56%7'K)JAR<C[W"IGM7A0D_G)#?2\.]O!QI!3X
PK(D&0^ !)ZUZAR6N?&,X;Z=D"\M6&:T4-@GT-8?V5Y[6SFN'K^#U5C9O4 OW[P<X
PA_9=[/D485/5A3KPYV31%S%,P,; 22?] (K_+$ 85M/NQ&JW::8'2)Y!$OGZ(D2,
P>4I_+LWJ3@RS91Z@?;?-?:^O!.KSM2L]=D,!%ZAR,I-32I#RK%B92N;HV@L[_ACE
PK^$A]V0(V*/S2E*$O6?YBBN-"FL-,U%?4QS3V.'MW9W\)+!8\S@3"<TW.M  5_7^
PW)>L#U"V [Y^R>\=.W Q*&>UJ7'.#E7E,&S1YV!\VDG^*S\W"WB/([D<MTYMC*E$
P'#")?G3<<)J(M&QLMPLL(^,L.2+_MJ=VHEO"KD[O]%K"PM/=HR5,PM1G\XZ6>%_R
P/LT+D3S -WJ<(;0+9I(5C<*UTT"A=/*7-N0^W+@8]U)O</P:CJW=@:>MG>V3=/#)
P>;:_QF>0;TFJD-D**"DR+\)Q1I-R1\<^N#IKWW59RS/=0JX+9EI@&*OQD?,82HRE
PK)^@E_,J<'VJJL(TA!K]"K*U[&,PS)(>U2C&+Z/2V="#70M#XF8\ #]$X$F1,Y8C
P7!G9($JF01 O=^@A1PI&C.JY%S2[FC]:Y$C. R&:/N<(8:-RV^.="V=^&TR=+<7K
P3ZY,6'-V1=(, _LWZ6O+B3Y!3()<R$RO&R?ZO9ZP1#]K^B%>=>,UV9/BLM%*-<A.
P&6-VJ<[.7K=NT68YWXETB,U!LF\S9T6(6#HI^01*GV6LHYGRQC:%HMTS1#:6E&J1
P%C+#V@#,Q\1+Y0(__4[BCMYC=%QO'^=?$8ZLL:7&W?EU;V@I00"FB.$\0%$OD/K,
PEMX!\CN8Y7,QKS:S-B@U<5S_O\XWH_J>6)2K+LMM5NAVQ?1CO:L:34&7L0)U!"^,
P-M8:?& U&S:HBJ0@F'V=H,\>K!AA2(CI0<-S1>W.GG-3&]@#-8)%!,E-M9$'9(N(
P2^;&,#!"%2%8^O0FB8LH/.M=!38+E2F2HK=I[63E;E+5;Z:#7.2=Z$9?<2O]=>2W
PJ\Y^]2DTE!-&R/XC@!1ZK&NQPY5G6+'Q__9U6PUG6T$IN'U1/*F;$-N;WLJ=.?"'
P(3N/"Q[@*QP?5O7(&9,L:8@+.[@H7UF;\9Y @/;!"<.%R$M4]( XJ&DMNQ B/F:U
P#!>8G)96!W)(VS79YY+TX5/RWS6;JL9E(F5J1BE<LJA,1EG6'X(J.Z7',1\YQ=[J
P&%(I>!6L'+( ;^"8BO ^B3%FOQ;<<$6>Q34)^F<^48.@.\(I,A"O>%0Z1@#@NQS/
PKOBV)>=//1Z(ENH!GT:]$1;<%'ZOV:XL@X#ZQKFKM)S]'IA$+G*Z$:I'9A",#6=9
P+QN^WP&6$[N7E)#30OCY9>8)D0LF8^I#&XW9KH]B_DD%V9\!+<!J.=V< * 0MRB]
PFA4#VEEI];\ B75Q,]![3;>IC-CR]"<6_84#'Z+(RU_P*.IV(=3K<@7B2;0T:_4,
P;T*6501$N?AU TM !B#G"H((YX4NEF6+591O8V$R;-4T!/N<']?4&<AHXI?''SX#
P__@OH,'B2_A"(;!E(BI@J WP47P<K.QET41^W?+5(NOI?V?2;_#& [4:02IKU-@;
P[ES!IO@TQ'G\EHBVR6X+2AES,;:3J[1 F!SG*(]=W\9H]I3J[)/*B7Z0EOY].&K;
P[,QR!B(/%@CDJR[@&WJ=MO#0<$Z!M9U[4E<Y!#=/]QSLQ!W?)&3Y0H=Q'H&R"*,5
P,]C,N8O2GHG,>Q&'[Z_;%6W'2'<[/A2Y@%;+X*1BAD6ND5);.\/50<<S1K>)1:\&
P%D\^:BSS.Y;PEL3>O0"4#?EK 6"- UB9C3,A$CN&T+'_,?)KR)8.>N__M591^2TN
P?CR5I(2QA7]8?CY00>>AEZPVVB+3,0P$ L-I&@K?KCLP"JKFK@;6/&A_?+D'Y(GG
PRB47RZ1F49#2$P8N1$VBA=X3.1:  X9JD_#:;@+YISA9!SZ\<4D823JC!]>\G]]J
P<X3W<5OX2)][,;-,8P6G-6J7SDN'W=42H#5K#]A6#V^5A2'-(H9E#:(<]B8L=$Z'
P4^&)Z?_,!_:34\T=72QL C')E#$]0K(YM; N;:[+,=U"U]CU+"SWCR5<2!R+JU8[
PIP4$,5A9T':-^@T-D .[(&.358\8@&_736]4@:1*I^=M%S92M38KR$0 [PBS . \
P$.D#E0?,96$K>IP)(R[IN?EX^B5R"E6 (M)D4YUPTXO2G(6&, L-;?W2IFL#)9PF
P?;?..#R ]/8<UK\SS@ZHZF(F 0'!I'!LO+-^U0:A[":0NULUJ8+=:XM:EVNP#,7T
P9S5&!# 3F\&S]8$&3F33&.%0Y$PF1)=&T/R4K+3R3DO0*))O^AG2%NY-Q[-B+S,5
PPX9;J/!;8F:\WX&*X5TSQ6UXU;0:6G<YZN9)F,P&?!.:FM%^@"ZS;10 ,(1%EF9)
PT,;+_Z%Z4M#1<_,PDJHSKYV",B4+<5D//3LN<UGSQ&Z63\.RU$N(,.$+%"I@?K!+
PP/RG.:YAO_L$;%_T/H?-:?_ _-F?"TQTT7KI]YQ>PT&IGV3YC*2CY*KJOA["<<[_
P7N_*?+BK'V8MI[V8 !=6 IN2]3Y631TM J8B=EO3XAF=I,%(I["LYK?<.&NVKO M
PFR2K9O>)?FPRZ:-TF3U9%O1)I"6:4EQ(0U(%<@7HB[IB*$X.).3>MXLY&J0,J+4C
PZ:#'OE+C.5^3YGU8!9EO?@]RNU;H-7!SAR+!R"L%5A0AQ;5S*$U=)L=TK&.D#:_M
PE2/<^;%7< 7CL>P_?K4+)/4W12RV@==P<6F"J >7PLT@:)M1J 6R_5CM-K?9&V[B
PFQ?=C67\O,;./!HF"-7@]V-W\H6D_6"<F<:M;=O_MZ+&[_>S>*+1<O T>A!7OZ (
PT:H9-'Q%SY! )\E)A7WTI*S0LH!\*0-YLY3,:/$/)U%N>!]I0$R66=PAV2/9H28)
P2D2P<WJS=$MZ%_[+K;%VX1T1,#)#3=A<GFT@\2 D]T(J5<WWM&7^?H!P PW?&U1D
PBO!B+4P8WG?])^,]4@X 1!=*?TB1,07 ' SK3IT;1!\T\L"*:&%%@2:D!")IW'(*
P*YW8:Z$"K?X9$SH]H<WZ]W4#768 E%7Y01,'F)=EB***K.RW8VKWF)._YP!G>YO_
P-^*:2$<=H?D4T\O-5R?B6@%)-^]JZ.N\\=?<<JX:UB];3J9ED(4$;];D]7VE6.X#
P6_14N16<_EQ6*@$V]5-$*X7HY_@A0GAPT-8U>H>T:3"\4?TDPA/!4><7JR9A7!9N
P5#T)Q?)IUHU[MZ55M+=QI\^Q!"$;6R^YZ8CT\,-D5K-/2A'N(5@'S_GL8HBER=*P
P[2R,C%:"T8D0O*TC=24TJ[F![0VC2/]J,-.SCG_?A.)1(];GL5E[@[E(?!]=J-XJ
P.%A.ZE!=4 E[,BMR'8T0JX.EE_B]:;VPG KX9,S+H'9%,#0=^Z3>"/@8'Y1%8?$M
P"/Z2]'HDPXT%N>-5'"T6J-II)"]KV,XGK\@#N7#PPM)D,!YS'!3#=YPZ&%T@=$L=
P-PI\C@@7Y%M9;: BB3;#!PBA TM):&T#:D[>!5AM_G@OD#@NFPWGX&J)MF0^M'.C
P?KDX\)HG.)+P_-+E3$7[_!_5I0[.6?<F"G&J#KT6AG$--W:!GZT\8,2[ZJ3XB1OW
PXV?@XT'#;+S._,S(AQ-IR+(#<;-=K1/2Z>Y52$(8B\^Z?#_JIA'P0WE1HL]9J:]:
P8@9ULB45I$@#.F57M:8_LV D=GD-.JKL7IEI&GB#]&SL7]=IG =&A/E7P\T<-%+Q
P=+DC.F9W_TVRL!IET(I@J7ASS*"7/^(&"^(910XYA.U",.+1E!:P@40 X^1"61I"
PV3OOR8#Q>\#1\PL1[KK\OF!_9GUVHG!_!*AC)*2(*]D_W916?NP6N1R%@IVP\.]G
P@0GTP%#)Q?/$A!4#@&W[5H'\I)GU/+2I7 1POTXA*F]/4$91+"ZL%_?EO=1F2W;*
P#C0P*NVG,H3$6]EX>05B7:)I[=L_,(.5?F,;7J?@S6?^L,0UQD*F1V3P1,63GG7.
PKBOSR?,'M8BNX^^U("#(;'+[+DM/C5UMQ<A/HKV;,;#4*E^0IJ7N!)&S.JU[46T/
P4K'80A_2M;.:4M=BM##(P22RP4@2!7?*MF^S.BZ*)6 G?\>)N73,.,,%EW3HG3[N
P=?5A.+[H,@I-9= H1-LD]?P.P[A?JO)6,ZD,6X"+$X]0OKB&DC+JL4A'EO+)"N5=
P7W]<A19!T!$OR*>2RI- 2RRVR#'2CJNGJ!$FHKDS6DH]9\HQ!D3#,[EH(X._-PC_
PE#NG#=/L-MTSP_MJ:EC&4;=B.N;\05GD0G1,R..2 ?_NGO'>X'H8HEL*N_J</:X1
PS,USB<AKW:??OVU:E'@PS<FC3*AS)R7W$&5H GV(Q15U,(].D2CK$9=AVD7P]G+N
PF+U39)AZL*^Y$+W?3U/=TKDOD5'"Z;P4TC_7+PFBH^6 RRBI'$#8@J55XS&X6843
PQ*-&]JTNA4AR!C&X$07L4-<P7*K"ZU/.\]\9GH*6F$GKC5&FAS+O7X]+[:$ZQE @
PRBT2T68+RD>_*#@?4I,914\)F8B(P8-(BJJJ]T#ONX7T-9&Z;NUBD\%5IS*]%_[P
P*D651;GWWWC@ID  ?W1T-/"?SN*[:(<;Z957GYAJ,V[W@9BQ,KGT+_J)6-X_@C#U
PH-4Z,YL9AUZB_=(#NIL_<M+X[FUL8&IS%1\I5AV)O97NJ G.P0ZJ.8:V0ULK!(PB
PF+,47]G\$M#2\Z/_J46DN*O^D)U)U.G_+;6XZ'@MBNH89[SU0CRT T>*IR=:K?X.
P88D2);9PK)>L>3.-><,$PK>R2;@:&O04-OZE_<.;]Q6LT<%M\E*#7Q"=^Z(5"$HI
P[#M#R6^%4+T%-I2(2!0MM]?_I]'[6+O$Q5K6F>M^Q\ UIYB8.["/UNFA1\R,+1"H
P\>6#F,-TX_5P5/XMB'-RHY^8L>$HK+"H)(-&0QE:[?6N9WL;'R64NH. =3E.5'KR
P9,R>R7W7S]KI&+!P87_KD?N._$>O>"J&.(O+J7&[_EQ^L-7GNCW^K)J,0 *,HUA_
PE?IV[]-F.<\-3J<>FES4T#NUFJ/7X,'RIIS,M$O[=%XC<9GV9XK! V <O&) (;:V
P%6[P%K::WE.D%<\%;7E[A"6E$*QV+9:/J,(.%S?HNAKK4$?U.@,+9X&U8.TT7MXX
P7&89M_]\>H[WT:?VV? 7OW60F__5MHQF ;%FJ12=6-'Q-^[19TF\A)M5K'30O+VB
PY_.NJ82&=J[J+EU[F$Z[+W&?NLLS:?+3@>A(1B*UEX/#0%;.-@V%Z$[E#VEHJ;ST
P.)@?F?'[-^]FWQAP*/["\;M[5F) ]C2AQ(@Q:^05-TA L[%X;7K)H-CSQ-85U%6]
P<+&1W5*IB3AJ*:-?+F)2T@CC?SDT'&^J<W$2Q$5W[DOO7I4;\3=$?C7I9Z4DEW#S
P"+P3RVQ3Q%X7ZCQ>H)YQ1*_D!;.AUJGAN?="RM?:G$Y;!OP3=\[PZ/5HC 0Q-RQ!
P&^*RSIHCA/30HEPK)1(\\;4]2VU$'P(\2VW@C2\K;'.5R:XNW;W)NN90YV0=T6/"
P2VJ&4_'C=V(.SJ5PL: *B5@B!W<H4S]3I">;,^:',>>[>*WI>S(I/AW $7TOGQW(
PB!]7M[<;ZA++2O8:O5Q.TDW%*$ 9D;LFYJBC86$?!0SF*408DZDWYN_3HN#/(^AY
PZ.ZM>\DU+ODMKG#05B@KJCDXB4K8_#!-^2A* %)[6RX?@&MS-V-%.'(1H?&.] @<
P&#..RG&HLHRMFB_TH\6T_!3%V^A?G*A$IGF JE&$.N&UB'C"J+882(.>Z3N>7V./
P9C+":,+0X1;@2I@+F,E:>;DL=5U::E62;RM1U8)5X?J)8C1UE_E^'W&C7NA#;J(+
PW/6T@]3W1+A:%_9Z>0]#C+S15.@G"8^8SK2MZPM\BU=BLK[^;=*YK)==:X)B(LJ)
PS#OEE^DVS,^11?D/L%+X"S#:QLL]?Q=Q?=1*;&/XF&TH=&ARC_^%AVC'%'MAR\YG
P)+I=Z6UBV,4,8.7Y#1&55^@3D6,@&SAY/>$K.7*$F.[99P)DRM9P71R%OMCT6WH=
PV5/G#P%^%"7YI4>*'CD<+LD!5-APZ8^<I-)S(@BI/H_R;[GD" )2]3/*%E=YDG05
P=19R3KWHJ&EOS7=V7P\_Z)($6;Z,+*R.<A5:$]0B7Q^.:,; A1OF9J7,P1TW&X%]
PIHJ_]Y7UP;V8E?BK:L:: 1&+:NC<X&@&;Q[L&WIASLRWV_>:PJN*8FSJ>I>":7#;
PR5Z'%'_;K'I08D@J+N9L($FB/6.4$)K%C(V>3>\=FA0P[TK=XBC:7^55>A."#79H
PG_C^G\C''PU$L-S<8@LWC.ZLM5:B'@5)1IN[/P*>['.[?8I$0F&+$$.EP?_[CQU=
PIGF/DLVG521_%%!FPTF28XD/+?T&EP6U%X/B?3^.$/T35[D[FH@"M)93D;Y08U#D
P;W8'2P!+'/A.RZ/P5+K;MMAWBO[$_BP;]N5*$D7+P%\<9G@+#4/B:?[+[-TW_!('
PH^]&47?25UA,I'"W$,6QQH-E)_O7H.$JLN')BL"&E0//10+%5$!I>BX(4 9&O,%X
P7%7CKESSV F#2TK32*%<O[ZG7OEM$=H]#@Z2];6$P> S6A"@6/PG203YJ*Y 8'8*
PC[$V.WJ8KJTX;2YE$%N!]>"/W.)DJCNF0<( C$9? J@_HQI:*[2'^ +,YK$8(XA+
PDFWG+?D9MUJ>SK:RC8S?%I"H_K6M(Y,>CI-$GHEPE5)#EZP<:0D)OE+R^O@'6)I\
P?JY3ULR]OOC-ALPL7YI;JDL?'<=*+:.&6,I"DXW!R7[RY[D(TTQ5$OV:BW9>C!JQ
P<CXB.MKKP>AJ)$. $>*Q$9?.,VHE$&PJJF0GZ:BBHM:$M@.:EOF"TL=;_.+L9%DO
P\W)"M3-3MD6H#^U@@^=^M//N9(.X(7CF^190IXL0/S'^29Y*T(5</*J9H22S_Z+M
PMM-$62]W#YH._._YK5GKS&S 5<>*/ SMV*9)';72?W?C]8JS2#U:U#'R0AN'"7:5
P@@'K5Q=T.94B+<>'"+34C6R<&/I<@$?2X]87 KK=6F,JR(?=PBN6^K7<X\*X32OQ
PU%;:)7#]ROP/X<X,]!6-[ZRY"7Z3_3E].?H_].%R)&,>SB?&+0NS'\'C:('")$G$
P\*/:LER;7 7 IU)90G2F3U!@L.9K@.^H75^U'9 :P!R_\CU:$A=I7<. Z?8<2K_.
P8A@Z,%US:F7,C<@H;\8/RJ*^^>P@4QAJ6;Q\2)O9&+:4-Y=PSE+].NI(;E::=6DC
PS=MTD5[KQ)^']1OHSUDBH\\ &/(XQ_@WK@TC?JOA.FN@;QXZ#Q(]+QJ0]7NK7,_\
P.8#^S/)P.K3#[DN'1NL1<ZB_I"5TL58H\66\!_9G=NYK<(=0-<AQ_<;A,2<4A%J&
P7N(HN1P=OU'W%L*R+BD]V2Q+@@0#8@&,O.N\?2) ._IK>-TGQVQ9_V&Q6"=VT,:Z
P0&0@BF4_JLA-7MM.A>.<- >/4DF,/%RD+RX/NG1R,V.["X5 1Y8PN'BDZY8.-B]9
PS%4\MKYC/*!;?*NB(-VK^:1)*U7T],@"@%-?<(H7,DZFL6Q^(TJU%IB->\[\<<1X
P2^@DX2 A18?B[4K6EM#;&EUEY,0H4U6=NF6Z'A#/"(<-B-/R^QW? 'B\G]!-:U-C
P!.RKO_SIZI"*/^_9%8[,%IHXJR5H1((S+/A@Q'ET-=YWBIG[4VRS<\ZJY:=<D8"N
P5@K"+WX;PM-RT?'= ^G%!9RA>E?9;^YS^J!U):*.0&:3.H\HM4SW9LEFA&:$Q_[>
P7D^Y45/9@CSE0T1!:^B),0-IH8^@ 62CCJK(^T*<ABD!)-R2E//E"SM:/%H92=/:
P>AG4H.@I;H[V]QZ>)\$P'M>>$OR^)?K' H;,DAAV_\;1\0M]=];CXFO]@BARA>\$
P^:0!WN3EM#M-BC7R.>!3I!5[6S"GWJGO5EQS*%>DB/_RR#U6GS_A8#=6EYY!E+95
PE2EK./$_'7MZ9Z?CLWG3@QPHP;E\Q8J!R B74G'MZ0"@+!;]XE+I-M':Z"4*T:"4
P[.EEU,/SIW;R B4/X==2X5:D0HVQ\H 43)D%A/ )"LXX;$\,"HAY;SK1N:UEULGG
P]I+/NO#%,@HGI=7LWG\A^6<V\M^;\)0QS\TSU]82\'J@W/"@>Y6#4T-BG\'?=/'*
P2J/(6R1M_<1YW&H<7\-)3B@^"V1=X^LPT4IYPG2Q>B39;$> 53N7#K^0'9.:*'=.
PBOK?N:7LSAQAJ56UM!:I3X7KRC:<,JIP==701^5QQ(&UH5]_WHZNSN/ [D&>ZQJS
PV.ABOQ*V5M@!Z=9[BZVE26BG:Q>FC6WY9CO!7YKYJ+KU3[W#DJ9\IF;TWYLM?/$T
P,S&7]:LO^9W=I?L2,+&-RJ>7HJ!#0T66814J8WH5MTN65S[G[;4]LE3;D6D]Q:O3
P!T@LUI:,[:J]L\BEDAOE<IH=.&JP3/M0$V8)U<E0^AN Z3#N\ A1OZU/]'=<R];Q
P/]G1!:<+6MYF$KJ1GOCX -P9I*HDJ^7<PG)S4<&#^=:EB^:2UX!9SJ7,LOZ'%34A
P88OP>Y5'N_JUNWC#*W2NR^C3WDR"@8\88UV<@"ZO/!327R4@7H4>>#$-S;-"N4',
P)-JSO#M5V_[V)D'_F4N[*N(=,.G*H=YMX[-0"1'0#D_%#CH"(;$_!4D^_:8Y'R/$
P9\D6XL%2JT2$ JB)@BON=L+(C?;BV=&Y'I:A. %S>:&TV6!041>6)2Q_[VH8G[B 
P(^'WL:>JNNN_R%V]\(]YQ0+!VD>;DQ-JGE(E_>FX\=CRXD+@>YF%^VV,RK !D(\I
P<-)BAGMZWP>T68%(II #*GU\^>O+\F)" <?><;B/?O&2!U$8D)9!B!V\M H^T$^;
P[.A1QSK7UC75,?^+0G_4EO\X9ZE=M;%8D#X.T'1+<HT#%PG]>$["%=^2]2:42C%:
PSFN>SWFF'S[P^/W$S:B1?TD'W!8N6N+4_<%J&$6ON&6_,!EQ/+DD/UA8++(#K_&\
P[O5(X >(]]\C NM2J*@HH5@Y:95'A8D1_&^-*^J8?<T4OIUGK,^9-G;EI(JH&'8_
PAR-3@UI:)1.X8%Q#B^U*.968QTZ\D[+B __83JV<RQ9-#&Z\^N'73?7C9SOEI0?%
PNO1RI4VH3$[R'MY)^LR\%O6"!62MQ!=96TS+2&/G")#2>^@QQ8$#UDES0ON"LO8$
P1#25??! - =)J=E6/CVS 3)5UD<86F)]2PB<ZS$'BB/>,0-6EQLCXV0>JM_<Y7Q3
P/%C IO<6-/0[N8\S2?U_<BXYX>6\=[%2H]I,P%PC7$;$R'A<!^$23&*34#V!O'ML
P2X2RAR2?-5OT+C$8<V=6$G]A+WZMBO.75@D?#GZ>YNS&Q)=GQAA<X7W&RE\R?>&R
PQI"CRKE>@HP4J+=)951C8(D ##=>X1C'8B80?^BH=Y@'$6YH_14M O7#KBNOO)22
P]QI0S%T 9).,2M+V<="K.=L)J(8@:.8639F+4"-[@--ERS#0*%3:5-&QI$V>1-0A
PH"N9-?CXIZBOI;;E@3D+G!/I4'1K[$KSXOPBV.&[_S&\O2-@X^A >[^R_V?TRTK 
P]4! '],<G0X"(-1M01M&BG]KB0I =X!7HCZL;SV>Y,KC!L^U:XI7[[6WR+#!.ZZ$
P9JZ<5DNW#DH6&64+'5 HWTD@[QK1=@YQ_(F;<^#2_D1]G98C9E&?W7T.[EB.'4B+
P0$.NR1.W\:TR5I(X&:H419CF(NZ!?(-=AG]C$[I!9!$YE$N?*Y22>N*B#-:1V,XN
P)KT+L(5/>55?R6\BHU0"RS#MU]284.Y.^ 5.TN9[Z[!Y92]TQP@18CA=E? " \P&
P=JP32G-A^Y/CG7#<M<OML/L?]\PQ<U;H\\M $]J<(I&<W9FM+52Q "XZJ L*?!<O
PPC)DQUFKVA/?O%6 WU;?UN./'H5S9BZ!C_/TN&Y*"/7[G<W\Y"PE, -"%H/?X^]E
P_I_$:X;9M%;N("3S6_4P2<ZL]26'-FU>L;>I%A*>5(7(*6CQ%C4)%_,E 3Q-$R=T
P%/O.!AZJ6Q4#+L\NY3.HC:3D]\76LL.)^I4Y3?8:^#2::0T.<69K$@!NY64=+.X]
P4=C"5 RB!].=@7AEL&^(1Y4<&JN \$CKR1BV13V#HTTR 2JSIY=W(R@Z.PB3F(AA
P3)+BHG*#&W[R;L$<WC>S;"F.UL1E=?G[R>?>B/5QT4"2+4-C_J3W&;Q.41!W95$*
P9OK)A;?GPWBTASIAU:;LA[S_$W.J]!4@)Z9>KA>.K]XA@(H&(_(V,E(OS44?9#<E
PH OWTQO]S36YE,R]R>)3T2HD \ZICL07E <IOX^T>$AC0J$R<W E#Z)2U7TWG.P2
P);WK +B($1CO-+IC^.%"T/(0F3>(@<Y<_5-.9IX=(8TG^6UP51XM?\P,/YV2H:!'
PT[)B/JM%#:>$KQ](IC<[!E!%#7JPFLJZ'YGU7F):CC@H4\\JNT"8E>\R@8*G#RIL
PI*;E,/C,V$''IB^!V-E84/4(.0LX]L51J4"ME@%BW8#[ #7X!9J8TRLZ-[6PZX\C
P /#FA\Q/AOP0G<%@69>6;M1DP8[68"W"WF6TG0XQ'(,*7/N<UFG^#M%O:&#AQ?\Z
P=8J^26)CUV!A=?XP%?JT)B1^].QKLLET7V?LS:25@=)6Z([.BRMPL*G-0K#R^*+H
P/C'L$.SF"98SWB33;^9RR-&]K<.663;K8<4YC$"<&[?.+$/2LB\9#4;L_B>C,WJ8
P=-F?;C)H6H[DNC0E1+!GEW*Z4E/OZF,.Y=8(:1JD<N $">&L"S AV2S?K^C%?9[T
P/!!N@M1G(RK@0D7T+O1 W2B)#O_^/X4J$5O8+:_L$(0]=C(;%)DU,)M#^YU &B3&
P\@PRT?<U&)U?M8M@B/Y0BGE;KA\H7+$5N62"'B)XL@UG,[L:?T1C141N&Y, =LC&
P0G;VFJL2!8:G:(T4PL6*,J+ GB)_&XJ<+CE;N]R;GUK8A,OAX3\;$+G4P+#N@,1O
P%#U(4GFYU4N>G285'$L\AV*"/>'-67"8V"E9R\,F2 (.V+I\);##VQT(M%J..T.8
PGY?K[?M\OX67E&[A_!"A?\9+B_D(R?IME-.H#0'Y9&/H3+5.OD<7B;Y_-Q,9W-45
PGY6M=BY!X$)*UVL+42D;6BS-WNPR5'CQ#!)FVL<!R[<@U*<G,+M@@C9K42[KIJ=H
PR;=+0L5 D;71SLE5NP4S/1M<ZIYDE4Q_&M[K&/:8!&\_+4A;:L*W>G@#U&:1#Q6+
P]>OFRU+VI.P5FU%$<U2HT<9$7#C8EFPRT(X.MI2"@N.GTR!-<:O.ZAXM##^M+FRC
P27*HC9WCZ$RC(&#%Y(F=^FB($>!?3)WJ2 (<H\-69_#86XX.?BJ<L+SE?".XL">$
P9Y@('>8&"O6!<\+\V0F:[,;CI[200,EB F/5UOSVI/]W8CKRM\\BJN-Y@J SW$F'
P?/1\K9^&%NO@*L&4VS.L.#K1O54+XR;%7%@I#!-&VQW:+A*(AA8%H<K*X!O[,510
PUUO@>"ZL*I0&KHIW"@H70ZZT=H/T0*YS/L-56FP]HM([U8PC_T9> P.E%SJHLRKP
P[LNL6%N!C)U%"L4\47,^.BP<%[A[AKH>_(Q1((A"I9DJS'6<Q5,%GPELB_TCA+A9
P*$PB>U7>^V5B^NH54D;8A#HLV0^DS9;YZBVYY"WL=0X%":1420F97T5FS"8!=2C>
P9QVM"%USD5EIYYFTQX+DT[(&8^S)$XO!.:T83]X =?I/1V!]S"4L@)_!AA@;NU%9
PM3K9QJ.9FBX#.)H3HAI'U(+NE]<.T%143+Z#$:&_571D[U;E'&]1,KU8("[_".@T
P9XL=4__+MED_J]J7K#N.C";HG0#8(=E9.2&SMBUQ-YL/I* Z=I48O)I3AMD!^7.L
P&DE*EC0:G]#C^&W.KZ]\+](!; 4MTC Z[HG N9= %[2*5<)NWW*?G6^8Z9YGSA9F
P12GTHIZ*?+/<:<M0HHSL#L2<C&9J2L^?Q.Y_W.PC5_#F[(UR3__R/NY!5FL4;P&&
P2^=3)/R0&SFDF,FJ?#<HWW]A-KU?*G>B>0#U[=AC.1(#1(P5EFB%'?M>Z*<3\YB\
P,=X^:1M#T: 4<9YP9P#SUC$AG):KH& *0 ^K76%F!#ML(@:R,,TOLWB.!O8KMJ(]
PQ+P;1(JWGA$8IM XUJ"MFM"(Z?1W#'^89''S2_=;ZM3<K1_Q[ \*Y&]0PJA7EC)P
PJL_G"N+2<@8[!X1&+5R:Q1"K(\>D+Y3M^D?[ (C'$U<'1Y\R@VQ!N2)4=*E,5,KP
P])\AZR6M0%=Y$YGC!UB:F&?TVNJLT%[P[1"QDY ?F9V>)1RA$.N'>2M[!<6\[*?H
PG%0>$K/U7Y X N1B3R.%;51K56(M8(6G]4FYDG=(% 85!0'[NERN%&TC,KIBZ(05
P;T&+"TZ.)(<M8Z0G2MB^AJ74Z7X!'?CX6:A#E(_00FA :KFR2*M;&+JGW O8S M7
PX;DEV)_MR?*C#$/[ B]0%&UY+./T\GGS,Q'[;[B/@T $L%F<VW="3AY3?7@SD2CQ
P17OWP[MHR+$OQ\,<IQNDY,V= LZK>E++K"QH[8JGX\[Y=/Q%75ZOMIS3,-\9D 1E
PQ(=1B@?_A A:Z(2L"PL>(^__VD&6X:]0)E$AZ<?POW8XA2*U7I$N1@QJCGY76GR8
P9Q=:<O"]8Q)&WZ#P9V,T_(+1&;T3#XB7(/9Q%(*\Q9IM$;&=3KCFS8?!#<X=MNLV
P7>N_/!]LXTDN]U#2JKWS\5%H?-#':B>ES2RCBCB3)X;_G(EJYX5))>6C&QK>9Q!4
PMB!/.DKI?5BWBRX+FKUDR37&\,IAPE;!A<6 ),D?F#06VWKCI6;B&+8[72M"-YG2
PC$'RJH<CNO3F%S:?X(*[@,36,7BMM/7KJX C6)V:B)4#8R917"E)3&P VV"&C6%,
P@R$B<UI 9^)TL?K.(*F5/"XX<]%K*V]8T16&F=QJ&$P7W;?0#/*B]2WK!75&=B-3
PRYR81=Y!VNAXOTRWK<N59P.LT7/9'@ 7[*268*"5K4<B6\+(;S]5:IL? (_%C_Z:
P+\%45S@[ H-H\J63'8%V.Y(-_;$[)> ;8KW>"W/@LI. ,GN38J[O??08$^")<XZ<
P*RNB#EN[$:!Q$Q?;RM7#<D'$67Q:Z62\HV&@P-G9),;#3KVS6%*XY/M"()EGD\W!
PL&DXYP_CE':&2^M888?NWL$H8493Q##%37H_Y"%%+Y?7G/U$N3X4VVR>#U0+#5S9
PV!(G;99_DP4$UY!>Q<G0?6+'L0L=6N1F!PNN#(GN8*.^. 3R*G*(X)4$ ;G4YA"8
PE#N/5C%N0HY629= /&R7ZDVR/MDMBDC38PJ^P'1R2O()@.4)O>I<OK$\>#-.?H1@
PO38R66 ]#Q'_FGU88:O+ HG>%![!.S,0:#2]!XA)J-J.*W)X\:1YO2.%[FG51\D2
P%+MOV#<@9W/H<BI&VD7K;KZ&LNQ;?Q[2ZU*$;"UD=F1]D9&7C)>QS=Z8<BL=( #<
PQ<N-(>'06]U7+?FLD#O!\"_Z5</G;=\2OW/5DOAU7@9M;B\4F6S[H6D;I<A1V^M>
P%\%-EL82,;6E%]!9<W'=;\91X!A+>:_XKD)-?,)>T4B@>\/<-AC^*59<+F-OWNAS
P)T*#=)J+J8X4[,'KCLQ$]6.0C7M1*;$Q\2=L/31BE7LW62>Y)WER,IG"9;&FY[$N
PF#Q*2IO-3V/_DP.\_>5* ?!R>^S)J]:DXK2U-+E<L'V/!.U-RX$W=)T3<QJHOGBD
PMA:75\)"J(<%V]*.ZE&L8/9'5PC[QV$4)6]<^-"P8P:%3RN2)4LR\UX-0S:VH(Y3
P7I1XT@G4BCF57WV2-S+_K[ ;$.8U-2BF%N[+YI:6T_V+S@ ]5Y5LL"XW50WFP#B!
P#->YU185T"A=9,:5P.%A.V4;<1/AOJ1&'4H++$AOZAX:WL -8.$*8^@8EE!#K6Q?
P65)=GN,T$6KBB(1*.X"G<KWI4L(;0G"20BX@7]>+3W[]4AG)(E?4!^6F"L/6!\^9
PG*Y1\GZ!Z!-BNZ[,9+U5XA\?D%!61]DJI/3RP%S8BO"TK997T%-CO:A'>Z*30_2;
PF=LO.6(T:DCL,*V>R@"OH"H07@:U3:Y7:4TJQC?,@ ?N=,4NEX+.W.:V4=X$KVWJ
P_Z.KMEH1$6=(FQPAQB)DGGX$A'DA6*.SM0OOJ*5JU9G?+).7U2^2)-L9HY:R9L4 
P.$'9K)78U.5;Z]=0&T)\QI9\+<PWGD6^H9)YWIX#C4HK[M?,6L482)6BA_RR("4H
P?MOVP7POL,9["G ZER]._?DU=[K<SWNZ4F0481V/6F>E0W^S[IY,-G9J":6CIX;J
PTF0 8;J" XX]#LY>Y7UE2;1 *4M4V[^+QQJ-$6+VO<J#7@&59#/LCS:[I]ZSVBT;
PN2FGK9IJ"&,8\+0NHLC@ !>0!#SB(\_3/W35>*AB,F>!(%KO%Z%Q=/<.,O6BLP4Z
P# H7VN3S?![^?]<0&[#.;Q32467[79&3CB)@\3AE9T$'3O![I)PU@Y\OKY)P/,[=
P0WPW,1;1&3>%^2:]6^3\?!%WX\9K"Y_^JK_.@@.'86\R$3!0-@4 !TWQE,9+G<KW
P2+'MA VY1M20OV0/YC,R];I*FRT4DO$MBW%P,I/_MK?DE=@@P*_[BJ A7DCI0_C-
P<RO<H]J>J./QYP9WQG"Q7J:E6].QRDXL05%>G=Q@O35Y!VG<)F=G^XA'=*.G:1U&
P N.UXC/"@JVH[LL'@WPVE1Z>44.DRBB7\5@9[R#@QY"CFNA9(=H1.57UM1:_+J(D
P-"SA*+EMG-.*Z0N?2TZ\SHSF29%,&;$C%GM]PX("R^M/?$[ Q4K;CRU1XU[;&5+<
P#FZDVAE&YDK4\QW55R((WJRY388"GO7;U$,JF&&EN[J,^Q"_!A-,!CSOJ:N,DRHO
PYDQTE\AU9N@4Y)/TS%YM!_?+T<-Z,N]THJ3<$=BZ<JAYT2%VP1DH#*BIUEZ%"O2>
P#UWHEVZ/E2GS(A@I\+=U/ OB##!ZU:I8(*2$I%?1]K5K;T6(!OT;48X#!];;=I&H
P?2!@UR^@'6X;_B8D1V@/V_4(A,]/?3#4ROJJ*R%]D:8$SU. *@IRC@?M,8/'9XI/
PM2L]VZV,2=E!]84KZ'X56NV;VLWV EN^L:Y+ $$14.8VOCX!.=V>R!<*CU,?!P-W
PB1]TY'%X!$82:P#\6A/E^';0H"3E$Z^MTZ;+OF(8'WFI>(:Q&])/;VI1EA'Z>FPA
PW'38X[BN@CJ),V>0Y[A>*Z@T7FS2"\ >N2IIXHXX%<BY:)+95]B6-1T] ]J&UN>6
P?%.H3G<*X@RIR,WX_!C 3=SW)D2)?S\K/3X:F78>2N_LYA/9[&Z$$G?P#*?^S2+I
PF3R!40\%JOP4Z.)NZP(*]]JPP=B5"UZE4-/E.$AV%_K@MQ1.B$3L,Y,SQ:<F,XY5
PZH.#G&ZK?BZ"/Z(Q3\LY\LN/M]4UO5W ! DHJ)6@+-U2P'<E.\#\E.U<@8!0P^TF
PA&%R$,3,]G"5Y-[C_D1HF_JZ9)E\+O'#P_-GW@-_HT9#_T]*V/:M;7[]\)X.=K\_
P4 $@$)M?G$.)J?S0ELM+.E6/\T#.BX&=+:(?[4E3*P$>U@I*PR_&W)$9$.\B,_&%
P3')^$-'U$"1;XSZUQG5.!6Z(V% )BBA0+Q )LN%+ES]5_NPOE-BIF]=F,IYS(NX-
P@"HK)2S:?I\DW)YNC0&JB92M_.>Q%",%OA.'"#^IKW^N&)U(JN^@QTS(LMCL;YJG
P/8NMF<)^+&O)]2U9"1=>\ JI\<AF-2</6UKL+>!_W&QYFFL&'N&(B*MS"BV7^WD!
P7^VAQW$"UF'#M7RC9X^+L=351M#=E'Z1G^UEPOK@.Y>,Q26$^''[:F I4]-6SAZ/
PQ9%,!3L8&\SBQSB-SUBK6;FF\-#5V-@HXRDNC6P[-)?M'%H!UX1[VPPQ2')# 0[%
P<Q%5S#,%O]]Q<[-S?PP0=>V\K&V??%>S ,FU-LQ&'^EK01*)D_;+==71':48E(Y>
P0MJ=&E=?3L4XXPZPEUS;FY-_J$^!D?"-$QM_ $)L@S,2=*R-PZO0#VBO:80G%SX4
P,,OKV$:525>[H=@[O..DUL/T2BG-9QW-%>'!125'^AN[+R<.*&E.97(;20S)JQ69
P+=XFMVE!^HY+L1M:CMV\6F2[)6H\C<RA?M'>;TO3].S_^&P6&AXA-5*Q2H*/D*4\
P)4+!UG3T02(5M*>;O!_^",\NBY6-JAV\.::T6[:50#+[T0K+\S1@*/[6J6$^+GBH
P&8''HJ$?%=Q0,A4(I.B[.#7I)E.PD.E4@*H"ET$0A"ZEKTY#0FZ[NQ6S>NG"%#,]
P9G0B-WO [C&)M7>!)MK-SA^&5!=NI_Z$S(,J4COIK:II'/DHGK@]+X."J2N74'VH
PO 5LH]=UP7E7NHFLBB#CH)5H*<J%=+:B"YD3MB^I/S8P\6L<#;LTOLC)IUS >BO&
P4JI=Z!80Q>Z9[V383Z'62Y:-OT*]L(Y1'DLN"2\AL'@:>D\U_1'5+,XNK&G/"WB3
PN":1Q.2G/W=%8''Z2<R)X@OR_<24@[BRCWM0]!N3W3T$DFJK3I)GZD3L?P=S9N[(
P0YV#$8$?Z-*J_RS\O&II;D[S4I!\U>"U:1:L57M_<ARN#DA3#::DN [?&.'U<3U-
PGT4_K\?G59=.*&Q0K]"LY;12H09S>6PR>-X$I=8-6[R@J.Y+LBF<-B YCEA@NV2Z
PD=.!_Q)W^6]V<JF%C*];$/KBJBK'02 2?(*M/(M;2,"K.!.QK#5(E%F6)?..%CIW
P_A5FM3F:A\#*]B!,#2W*,MG_%SQB'4^TA7APN+IP6MYLIP.1PJ+F'GX8I)Z6%.L*
PN,ZK?['\JQ:!H-B'W*W22)I>B7,OVK;J<V:=;7TW8/<J/^_2/RXD91HC> "*N!3]
P(]:",ZS%WTW!%B<H\J&3CRKXO.;?2$!H%A3)SF-:6&4  L!1_'Y1#&$G%B9A%G+C
P<%4%1^"8MXU=^@AN8NB%N-0=.V/A"'"LOH?)^R \U@DRKWTBM",D/QX-PRL;! T3
P-Q#'!QX,*,HYU7Z2B27XA]$BA\124-<>+,D*$ZUNK-DPNO:J("9. J#"LDF1L.*?
PM__XRQ)*$>8I2OHM<1B>+;W1)!P S5CKR3#"J_L9AV'[*G?D#-44BUH>MFS*A=I#
P>:H=_3RC<[P]W[_FY=H^TGT]>9Y$WB#=RXXIQ]<S33#;\\?]<HG(W0$?[*M8O-*@
P_"//BT.Z3Y;%DFI9!$VU>";>7V$T08K2:@RD7(^K?D>#E^BDB1C%+02Z9/.C?T"3
P\M&TJJWL">;4[?9T_1*[R#Y[G _>$J#X7QWFW_ =]0\EO [F6P19^<%<9=F.<0WC
P#.+=ZY3'E+O/.>H"I1.H<@AAPNBQ@J^SM486;F#%"(Y.ER=TR1M#-?[5R-#5MF/W
P]1? ]&PHK[;#T:<5_%+7C]Q<DOBJAPK#W!DQ1J=1KK5^N/VK)<(9M#)$N2Q<ZK-!
PN)99P]Z,K]JBX%(3!K*YJ ZM3/!#P7K'6"N6+3:8C59EI)!O:*D<]=L_*%E67AIM
P0F@D)&98B"X@[BO^9$S.RJZ,+%3]B6?VPQH5PD&EJA%(8 [LHTS;/V7: E^#0#>4
P]MIO#!\PM-T\D?.98%<?*(@Y"(^#%;VV'YBQFD.]X_KM.X\"F9HN4;H$Y&=K8$)7
PT.(N'[I<!*>"*'1V(O32^I#1"3) 55SWTY7; 800?)4M;XE1/F!LWT6] DAM#DL8
P83@:CF0P>_ZLX0AW;'TR >%1]2&59Y)F3^7YAUOC5; ^+ Z2M'T1QZ(J+3J$V:_B
P72/Z#FI])OO$B0 #6U9\[@6</9'9  %&*A?8Z- #5D?\?419F]_W4F Z^>, 9@P8
P1G .G\BI^M@@EO?TR;K@>K.&$<)R9WO//3"IKY_M5B;7>P(0K]N*NQA0I:]+@[@K
P(O+,KQUAM6^KH;'?O&;!-J24MT# _U&\+L2\IWY3HP%/)TPPQ!U4,=3"!F.YWWEF
P<)VD7/7U"Y:T;G_AI*V$=E^_*#N)[J!1N![^*"!*%$D"!26JRGXTL&Y@, <7>,(Z
P_3J>@(E0(:E#T'?$%-G[[>Z'$ ^&!N0!76(Q&3 ,4-F[(Y&YBO-:S*_/@V"W I5:
P+&-_>83WS)%T/C=5SN]+\Q87,E0"35+^)29U).CI Y781>G+06N9^&P?M#D7R5,M
P/,,"/ER?YE^]F))%:>T.UP7+ZCBDHS%JTB;V/2-MJ7K!VEL$ZLB912;:YISN$S1Q
P M]IED#R2YZF5E*U8P\4VH)H#Y\21.T?.*H9$TQYE443QFD5$R+]7.TOSV^QL(57
PJ4RXX/[+D70/H]#[PRL,(W,<)WF/L24@3>.&_B1!S!J"05,6#:(@E=7?81"#9.;7
P;AQ,/X1H%+B3<R3]0GN2:W0&YPRARH&R*\Z'3=(I9WXS'1";GC(5O:MXJAUH/)$)
P1++!H ]6^(U"R?S$ =@U:H$1RT@YTOQ>C5%G+DL.*+#-&=\V5'+X-.XKJFGVRNI5
P U<)+) 9K##E#J0O=2\IRC;**>'>5Q1%$/I1KYNKQ0PA4!T1>M[_]G3>JG^1OU8$
PQR$^D]-RUF::P^M5\<Q#(UDS;1MD@O!F]U)U,DJJ=L"G%L$9QPDU>98VPK6?KH?[
PWS7)KY&];)-E@\4;9X&W-"SCW?0;5!HH17T?A9#2O.KMX=C9,75G:+:,U?U*G77G
P! K59!2BX&6X"Q@,JT"C!%$<:?\+/50[@E2"*X+L\!,04&;0H4ODM2,T4E:D(T8P
P@QO\2:XJ/WS"/"Z3H$TRQ: 7''*%J 8FUD>A:;"U[7V-F,S98PKQ<@&:(&7F02D>
PT7._C,D*UL76T^XC/B>SUT..5P+HP/C3W0K4NOG@SWI<-[6*TSQ@:'"];B.SF!H7
P?))HC+\ +FH366O1+:X6"MOCPA@6L)J,1!<:G<>2U\X$WX>H7WEGP@[!:(FTOVM#
PZF]3_';1[=NV2GB>:NG_1(W>,8N_F+V_:U_;BT"#.>:B>$@,M"TR?-0'$M8:M+33
PP_)&X"6C^&6L G@M87+FC&]L<\2-_@T.]$A\C>:)=PP6]$XR+*@>8YPE<.HY0[!&
P&.":/,7442)TMZXM!2 < 3B\7'GBN*V)C^VEH"W:DKHU\]<7;<K>TI_7*5_W&6HK
P4@^X:L*HI&OXT+)DZC+F+7H*$@^P3C"%0K,AU:FX[+S]GVFB\H?J3EBA"HY:J #&
P7"E8JDHUU5@4/%QIBYH/G/#[_JE$*CZ<:[%8MA#L>\>H/#=-70$V+[L7>0[6S"?G
P#J8](7P!#"4 [8HTI:XG&;J!83M'A<_P<8$_5E^\K'(2IQHZ(,8+W!B$QCZE%7EF
PRX[PR/X'")R<HY?QM#NI_:@RY;487T3PWTB'L_SWR@![V#.S2/2>;[3QT@$4<@'P
P65Q+TUB VLJKD^%@#2!Y&V-D/GZR1^^Y8?H1;?PE2?;9S,)N2#U)'M*W^'TW*[.Q
PA-)G07*'%0./ '?#5$VI_.YP P5C6^C+>G@N6_\4Y"T$G1V02,#?N"HT294R^.? 
PRX8@G*4(K\-@*F61)DVN2L\-150G%_O[="+*S'WU5.9.R3EJAC>)1A+28TLZU/2+
P]CW]2X)$J=9_LZ4F% Y.1VMRE!@?BUX1EI5M4$HJM 3#!74Z"CCHQMQ'T(JX#HY)
P3RE=5S$8E?YM\Q ^EQ6^;/>-,UK_:!'CT9'0JL)PLL/'A:?+H9Y]R\D1<PL%5?DV
PR@;!Y7AJD#_->Z3,7MKJPL)W[D;^/H1AQ@&3(HS;C1X;&E\20H*U<B097:3FVB/'
P9_/<;0<.I2PGESSS'Y"OZ!MG"90L3V*Q<UA0FYR#T!LV/S5Z/*;C_Y@..X[RMK1^
PL$1.?B?Y9]JMI%(A!,'*PX]\KS]_D 9\.KM";>9E%, ?P&7MS?GU3Z"C!*1?JP$5
PIR&^GI]-]8>VM?M\4/]:1C%><G4[CF^S#.0DP4GF =15=9_0[4X\$;#QLC*K2W]$
PN9B7/1A\7EW;?U-C2BU^*7Y.A W_&BLD(BYX#\_RM+0;B]BGD(3)/HBSI:=]][><
P9LW-N6O5C&A5?O'2Y_V]%)#,T!:WP:0).<Z'I!E:E2&D17IT. 4+JEKO*2V@/2U<
P'<[IR7*FQF>:S.3@)0?B;E@<9T@\9QBNCSSLE'[9@VM,&OO'.8)D@->7+OO1COZ'
PFL^@9*1IR?M2EGP+84)Z>3J^DH%X!ZJ"49I)N1CQ)DG#*0'V7VA%1)+E0<^[.,VW
P]OF^-Q6VS<BU?[S<- %8&+PL:*?5E-FG[1MJX$.7C8TGMUMZ+Q9WYXC^L84S3.E;
PAHQ(+';&Q]FOY5NZX5^,<G58#45X<'1K2*TYS1[E )FCD[+G"V04OU).H>5=5M!@
PM1/"L!H3]C+&3/P8FJ>D*(V(0;$H]6C!M2X%YSN=G. \PT['/M)X,!!41TO6"UU0
P I'ZD3S&!3N;408OIR2<-@E=/#7?9X$N4A_,Q"LI\+*W,3*X<P=:_X9^(J$8<>A?
P?'!PT!66T"3"2?,Y>7^321+_EX,+^$>\GL\_Q@N=6!0=0Q'=@Q7'*M92*^'0VR8C
P<ZNY)IL/()!%TF*$<:YD *X +%F=5^,TWLS<V%]9ZD#D<8% A\=1#3AM(G(U[;QI
PBK(;"%^0LM5$=H\\?F*!HQPI$%XX+"F"B#Q-_L5.+&,5(BJ*2F5S=."$V'Z@_7Z6
PQ?N3QCVPT9DMS_GUV#V:LOK/2%#":E0M/;/.)\/FN'O4M@LOJP\7/3I@'YY?2:NF
PAT27Z]_NJJ;0&N6*H=@=2-H34*#=M8[[OB_H4YW7("+,*I-P-="I (EL)DGD/J63
P6*?T*Y^YX3X"5@)$NK[K2Z3[W!%!+=/I_$<5CBN%>[D .[Y9F%W0Y'84/5>&VU54
P-,L&]PO/:PPG(&ML1@O[W2C"$:VB"W2M9A-/-P!;4%2EUD'C6-.N)4$1KRB+BS?S
P[Z?TNL,^ZIXN\J*XR7V1V EGX48GGVJ(99M0,HT%OH=HN,;Z$,H!^W28('0QD)GD
P3^G15 T@V#\WK^?CUKE>9:NRZU0=X*5+3'"Z#I1V&69<Y8JM+DZBV7=\RQ1^TKA?
P!H2DXQR^(<P*AM]8+=CO*'PJY@P!S7J_9N[N5\J$CIY&G+6^G-=^L108?8+LZE()
P<=S<"B6%=5DS*Y]K\[1]3>QC,"?2]F;,,"&I3DI_%5BV:YZ25M RNW)=W:8A&F'E
P>ULE2\6-!=$WA26BV,]T1HQTCAFJ2/C_U?M@4_YP/ACT) N>18,BKKA3#*A"^A>[
P6)(\,9I_-AT+LBV;!Z9RN5GW8"[IO>M\"NH+6,8PM*H0![^[ACEM1 @L5Q2F^QO;
P8X0!ZO%(NLJJ.KJ=O+8B*PDN[("5#ZR3Q?O6JPSSRG+X@X'>[C=7>H-P5>1;*J\U
P-*<Y"*Q"+F(>R#T<<44R7!5[[ZL E8NNB:+](#NG5B:2^(9Y<Z[K[S@> >+3.QC 
PSUUGL13>:>](5&$2-+@4')J\Z77).9<Z6Y[=UB.VVL,+EB'GPN=:[M,HGV'A[-FP
PAQ?M>1Q_7M O/@ H2<!J4OOUN<. CZ+Q-01OW_ND71C_V/<CO2/P'R9@^;38GCHF
PN0P8&]..N"CQLW9+'Q%^K$:CG>9!6R/&9PB"=2=.'8];5 ^PU"4.NN[QSTYVOFI(
PA.OLU4I9ADHO,[2E_YU#:=[K^;QT29,X S_J]1WB:'?UO$[HX#CU_-=OBJ$G/%K 
P?%4 [?92E!@++%]8/3R!#5V3W YB_[%3BQAUTZ#15__G:YTX"A4Q07W9<J[Z^MO7
P*;#@?%NS#JK#&0^7?*")@45W>-+\6L+>84\ B0E&(5*7-1HS'K=VOB1NI(\GP 2Q
P K&+B_9^<L&5C&= ;MS<;Z+<Z4=;A)Y*XP]F-Y%RODRF.G%B:OHY(?M,Q@]DEB>+
PFO)VP<XY!#" <*MC&W=[C5L[(.JGFINM>Z)UBCWO<%25&8!;MW9^0NLU[/$M-BK,
PO09C$A'T<P:SHJPE!:)0_;/KI@E@: 2T.CS!!VAHA7T2W/X$DB<;_3;AN;D]MQC)
P7NZ"H$=Y56#'W!2$^J3=QT&CV4S;Q47?G#1$DZ;]-* ^L[V%UF%+*27?ZFYF8SV5
P-TT"QWEX%!3?DL4%VD:>@4/BS1-#M:A$DT^OMTNK;!GY8H!;-(GIE1VP7\15R_=X
PR*>+V+-[/AG@;A]DUL;5Z3EC'\3 /3Z0KR(AVLD:+<N?*3YQ3F6NG/V@OE:\0GUV
PD?^*_]V8N$=J;9A,=3-91](9'JENW5V7P8[B)%CO]D&0#=K433G["M!_6L&I=H2P
PF)MO^VY%3P253KZ)&I-]QOJ*YD?1\>B$,-8SK #L":J_UP).R#+C3>(4V%+R$'57
P$99W?!6,6^B#B7NY9LE$:Y,;3Y;]1A])G^ !'\#H8:I71]8CL,:6[S.(O^;P_'HN
P<Y#"&QMSAA@%OO9\Q1C5\XG%UT8'RAN7RP&-/U%7[>KP-=9/"*'V#$B-JJ)S$"XR
PR O"W1Y#Y4 T7SLC; IJ/@6'W&_L&:%'S6( )@UQ@/C=G#O\Y#'4"@P^)6T;K=!3
PEBY-80++$Q<P3 D"HK7QR)A,,#I]%-%V^BVRO4E:?D@>!E<PVAR,"1%DS/M9<\%"
P$\D95&E%&PL8^+"W*Q3AS,.J.&O+'$7&J,E"/!__ESK":W-Y-J*L*!B\;5RRFQYD
P\3'O*%MAJE7EB\D04-9NHBEL>>3Q7%2),I"FVS).P]JY2 C%?NTP,VR#]*G^^A]\
PY&"!_,(?W-F8P*&P6WO=>GZ\,VIT&0W8[%YO9#JM)7XH&\*^-0=#7JT"!#PDYIMC
P1*FW64[>E4J0*7@=D"@$:#15^IA+B>MDEI22Y(K37CK6EVKK:/Y@Z+*;9WR@PKS"
P[C>?QT.7+!0)^-9XAE]L;,QQ)T"()1SJ95(Z(@.=RPO_Y@+) 3W:7!,5)M%JX0K8
P>@7KWC%9P-Q;43<UZK8ZKS\5(,(\1020^,ZQZS[QN^7C2"]/!WZ'N!U<H]8!&J]I
PS[X+F3<@/VZFR!J1Y^?8Z8P9.@P.[=\TH/TZTX1FOPB1BV[5G9II597N:F6X!2@)
PBIFV^""PI45GL<)5C=TU]J^3J3O:AE60_YE*ZZ&%Z&98>@,HT)![AI;)OAXG4?^<
P8);IM.@&&TD7EBR21. "!T!,WW_K$3]6-H_O0&4P^"O'7,HQ697//>\:^'ZH"<_?
P@PZ M4$[QX@PKDUR$L@(DC<3!##?:O.26W$O>1B1>;Z\C6'FI>!UU&_3Z"MCBNC6
PEVY>K2HMGTBN8!QP/K@(1_YK_1(UF&V\W>$LBWG5J&O@ T4ZX*+ :YDN>@& F-'I
PO:\;*#I3N*<B^3P9\?"(5'I")TQTEA^'=\*/M.\LK.KSD#AKFF'#_S!Z*_<XG]3%
PE]?:VD"P \LL;I[)E+8<^!#'_^(@<Z*W4C;7X_ZH,63,G,/P6/*8BEGGP5$7O_:"
P;L(B;=#.^?\ J'B&* K1:I-L!RSH_ :E^ZOA,5 V= BW+259S(7!RU:03S10%!+<
P6!<N^/M3UMNOZ0W/1X;P3@:!:EU[/\/[!G7<7:FQ*Z=KC]>*79[7%/=?>Q#!+H #
PEM%MG \AL?@#-:_N)&3'Y.\OCYVM5Q7G4[;SX^^)<AK\TM*['VYY._P"\QKUZ$<:
P8R#P ^RF*:MXBJHUBOC@:=9^2#H,M7;42R@?M>S7<*P5J^,*K/Z_V2M!O?%3LI%L
PY9J+F4K XB244S7\V[5&OY_THOQ)G\+0:XQ50O&.=^2.L<D[DL/!G?I:B1FTU]0)
P@\7PWQ$!]L%47_-^Y+XZ.( >29/0!XV=.AG=94<R>N&Z!/[DC9VK,;P7JF%]2.EQ
P.$TH3H A/43:9__DU]G_+RD*/6QT8D?[K! :3A<86E$^C"%R-N/I*T$/ ;**6<X"
P-YA^Q !Y[S:9L?_8N\0$M"!)HZ9!+U\I#)@]6>*Y^Y444ZIYXZDJA^SF89JTFB+1
P4,=4<)W7!@>]&>6!([4DU)Q*];5"&*LY&'<M6$5YT0LY "F=%D_X[\^W\[3]:X<*
PX"YGDTK*3/G5(7"/?A*-:SR;36O;1(^%7A8GRG7AROF,RPBMPA\!O%<V@<+T'A<_
P<7(;P\&A8IK&ARGY"SD-K7[B0&JNS2S244G$D"4@(]>H6 Z [#<-*JA5W/MK^@7N
P5\*!%(\)J[B"+J!GCKWTT/[-MXUI2^=F,;!U'+Y25[V7).5YX1&P?7#@]7>?Q352
P_R?YW,SFL[@HDF>X[3QRYH!^ONUFU$ @[.UM'#F>XSWL@0UW.29(J=R.$68Y_:?&
P4+RL;VO-NW:\)A!-GV'M:&FJY!L6@Z8(J.7JA\ 0X'W_7R -7&:4C7]11BJ+)"A3
PIPP>ISO<6$[Q=$L]U4G,&BK?E[(],=^?_/^4M^HY4CY[QM4>[0K>=.P@V:'<\23!
PRV0'JV)W?0Z&Z?X"FI; XDR@6=UN*((<&2+T[6*A7,/_>GSQ0.RRG$P?3?;.;:\,
P]B>:I:'PB<UQ1Q>;&L\DIONV@%P[4%XY)),(CL^KGX.$,DC7'L8G6]2>49'=XJMB
P'[/4HY+[Q[8!L']M%[]5NS+G7[BJ)O17-(@(*,\:;JA,.']QA@^TII2.^MII?37W
PO,]*0SAG%+43M.$1-0PO$7SHEJ74("*V@+I:6=D))\D=/(*E*5PK5"XXYV2J,(^'
PS(VDY2$QN$07/'L^QD 1AOIFFHZ<):95?/=> U HGY/ 8 F(OY'O5"_2A/BY7K8&
P7ZY3]JR)(!<8PN^I_+P'Y'>[\&L4&:>4SSG*X60G[HOGB1@%D@]R[+U2IW1R)"JH
PN9?DT[BY0-ANY0LBCXWXY,6E51^/'13]+<FN I>BRUYI=,<I8<-H&9BIU?*TCYU3
P8Y^J)^VGVIL:[4PY=)I68/VRI_/2[7_]5HU\%/S<ZG@MD&(ITQQ#68</(5)+XF1.
PN4I74%*4#!)VX 1X9U9:P;4#7[U\S<'P,0!$.&I,0VY;PKVECW'49XF@^Z^N3 -I
PW."JS_,,5(JJ32_HD T)+L/"*L<61\4$%2)J="B0!+#O%_%V!.\^$WY 6^MA5<;)
PHIFY^2A!&87KAPDK]PJ,>"E/Y@1JF$4=I]5X+WD#0EC<%"_DQ=PEK27,,"PS6/3>
PW#!B*SQ\=D-W:< 0[V=M!=3X@!2,)$5<R3:#(/9LNIE:E89VAC:F5F)7F_0:<;.L
PL+#5:>U(@%&!8QFU@KK?_N["J5#NH-G-'6UXV5Z.TVY]%.(W3/JCY61P1L'5L'S:
P>KS[R6]!?9Q.G<T5MRW&.V+R'?OWX-Y)H<S?O_-IUW"?-3YGJ?<%\KO2V6E"VY[K
P'A*WEZ0:Y!!\ZX]#A=";BD(S+/;4)DX(DFARD.8K)R+8X<Q17?\ZAB#L<_'894  
PP5I=^H^AR'&QUG,$?D#,/J.H#JHO353'J[::N4KHH?<:0)71NR3%Q(;3M*&*M8,F
PR'MW.3CG+2:Q3THE%7+N6$5HUS+\/\CMHT&'[C+:XC5A9:GE''1 0(N4\!)\ 1J7
PG?TI\+9]X&5P8[G(KJAL$+J-<A;CFJLZ@(%=BU@V2BRT-@9MW;53GPX54N_DX<)S
P]5:35JYMI'ZL=]$2R_GG\SW^)/06Y*FME>+S#<Q;8BX9HX,BPT.>M\RT(=E2VW5+
PM4FM\$G3XVE63GDN+3D7*,VRZ! *9<4R@24"!AFS874]Q7F=,5=A!U1X(Q;P,/4W
P]F%P\DSZS93/B$*([T#K(@4:T1.5D;93^-#@XK6&'4%5[#G45&"H:<WH#,(HK UA
PW;?\[6ECLA)_%VY2;O81NQ,2C3#9Q?Y1*T*6SXAD5'L0<II5=)=.74Y5J#WSSY- 
PNY%)NXJ3FR&DS\PG@69?S+H^@\[K>:X!AN3OXLGC\KT4WSJVOP5/MK7*QA-O1V/T
P(($4._ AJ]CV/SLL=WI\7M,_IY+?F3Z6!P(5HA/-]S L/KQW= OP@QY@)&PCJ24?
P<SIV"1L!.J6<URYWRWZCS&@O+CD=JD4.JF;_-1U!A@S[P3[5[NG1G[YOM.F$&\RV
P+JM&8!LWG@B\0N OHJJFYM:A];Y;#W>Q<)NVOA=!P1E+;OOG-R[TMK=OEO@\6B4:
P'&'/S93;?H*!BDK$)-^X9EL!$!76:WO^5&D3<N),,"#'NG$&UFM-*DT]2';XK&&0
PTTRO[@(UH/[*!^H&N<_GMDVGM>0%)F31)J B,1UN:[<O+ ;JVW%TMKYF%RC@E1XF
P+_H$Z_Z]F'**=:8R/OM2^3X"[HH"=<65)W_SS^S8YV(K6 AY&Z^[=TV$)+^[CL?+
PBI[@)I@<I!$[#M8;!Y9VS'%412ZI<'],J9LE&;=;(RP\U'^W"V2,/,OZGW7N<=;9
PX;+K>E]E?VMT]NS!X&$G_WRB4_GTWWS.0I9D@*;JXGE'W3Z.>5W&NCM%?]V401]:
PDO=$W&1?^+6W:=,XHKWOO>"EC*,92 F1'9W>@H/MA-V6;MG$^ ]WL,X_M&2V4?@Q
P55@;:R,^AKT:;OWL.W..]B!6-0WZZ;>^H ::S+BZTI5YYH$V"&ZSE/G;>&%>]$',
PLLI)>ASX;W6TB_ALOF&V9#T0ZU[BV+Z?FWTHP?1,P5BHT?EQ>80<OQB8"H,<)(L6
P<H1=2+"Z%+Z-E[W'O]YQ:9I#"DT._64P5Z\/KU5+>$'N)D@>4EMG=QWB9O#'6%."
P 5M8]?)7":$;,GM?=N.R!-E':TL#QL=&?1092<U+ZS\@[+&@,/(7Y?_> 3[7Y4IO
PO##P,T).+,-]4$,H9VEM"PWFC*BI:[/?LEEG:D2S!FA.%;=3YHBHLA#&CJM,9H5N
P- 5BBT!UY6.CX*;>L<$I\5'5 Y*+J;_,"]$V/Z6Q25<\<*<VR:M6O%H<;T_Y95&.
PYDNP8,)>K:];E#3P7Q!$=LB4E+>56P/<G(H0TA3[&#JGB3>X0>6](O?:(DG]#U%M
PG-8N&"-'+,"$H%3]U+WOQ.BY6%.ZT^KU\0;#]:W[EB)PJC"&DR*/D._2Y?6M/;5"
P-,F91+J2N.2!=O(0/,G=1;63BFCW36^II"42%(_/4@,'4>,(WAGA*\2<UV"J.#]0
P;GY=^K2Q36ZH8?=*+XA;J,V?3URARV6*H Z*JY;V[6PJM;(*M-5P4?$2O3+=-1,]
P?B#H,<$HA%GH26WR&.49$I'>R9I!!O//ID4I6I.Q\&>C63/%8AIH9R+&H2W]?]97
PG>O2](5A.>#!$]C(M3)UUO''W7@+!K^N#_([WND%9B2(4C.Q6OI #>Q]L592[1U3
PG^Y*Z 78;WZK+W-HU*+;DV<M->&>7,I[0QHXNYNT8P/E& X%AE"#KW!^YQ:SA@(M
PS0GMY #!/K'JS#'TI-)G0!<#/ BZ=HQ;Q@Q(GN$;9OVPU=L@F(E\HE'E5SP-N&?C
PH]L[5'[H'5B5#*G>R6Y8MC"7C7'[=V/ZV<4Z#FM%86<5;S@'_%?\%5W.T22@>.4@
PZ)E,E=L;?<M\R2;WD"^_3W6\NSTZ1"YUF&^<F+'QA41#9H>A7<<6^V=3""I ?MM^
P53.M'92A-_0*KM%%[EEZ)N;@"*591VU_RSFNQHJ+9Q+*;VFH=/+3!Q>?0F?O#!T[
P((:!")OG$8]ML3.Z"G=8V5,7U_RNRU\/,/58'63Q=@GA=\'V0UEE2NJ)?(C8%^F:
P=F6TA"4B5*D\&4Z/Z 0%&V=NAN3W1QJPIJL'T1DR0E9U\R] 9^$7P&2#N<TUY85J
P8H"6SQF!+#?LX^H3&Y^:&##8!-\SAR&R"C<;5][#OE@*]8$TSX0W>P%I(XEA@MU9
P[?[VQ6>IT\P^PHT ;.^HW[DOIB!B]]S!\A3.%#N)CMKX,@]"7GEA8($,M<P%S "@
PD8JX4Y>77J1&<,TE[1'CW#^=A,:2*E=3YBJ%0#%FK2'.<U2F1BGZM0<$;_!XWARW
P85Y5<#T.;NMK5)E5)#'NO\A19S1K67!)T/S9N7"J&[)L80AESA$8N)I-HC>0>X$C
PC[K2RU ]?J]"/'[ B ?J7L!QD&M5"8_1/U<H6#%/I<8L;&JGH^E+D(\+)NW-]<>I
P#V%3$PVF=(_>4(DX61ZMQ3N^MQ/']]DIEA$D4GB@693<(G6YN(4ILBD<+^,M#6*\
PJ?$9G-=,6"KTU4M'9_J+-!N218]]#K.X]*=4NNL!24GN!YJ-=>6M=:("_5K\4#ZC
PG&=]=0=)NQ+J61_BF.94*![7=E4("SVM2&+[!NZB"W2Y;PB(Q]!N+Q[ !)N(HV9[
P+LYJC'\NJN:AP/Y(7K=31:3?!11J[9,7%8G', J_=WF#'LPCW7&>@CL_ BW@I%B?
P!(S(ZB/T"S_@B;6@ 84'6S^SV6%'$/#L-Q'TI\D6VA%X9&,_\'NBRT._7:2800NX
PG&E^"X$OW+4*H']F;KTD;C\5%[KLP]KA9_3##VV5)X*0B%W.E(5A'!^D0)[[3UT-
PT:N!/-ZOG/JCDA=Q+AFN^F\^NO&@YSU/WGG5H,KE[BL+O:;S3HPG\(O*L.[<').B
P%\<SL'#?RE1"&6/J%_S%@<K$(Y/MO6O&8=[K_U+[>:X7H42:-(<$N]Y/Q^Q#[$LP
PNH_M6"MXUX'@E&:6;;4)N2^JO]!BA![(<,#VZMP#,S JC,+)]O*VA9!V*6_D.$UG
P4K^^.2QLGAW)D^B6GNXTANCMO59&&D3<]T0.A%J4B*G_W[E@K1(S5T6[]OXV^3I7
PPO+3X:%2A!IV>Y>Q0Z;*_33[]M;4""?.$0<%'^++'J)*(P]V@F_]>0(-FM,I(2QA
P1( =[]$F8;N?:H(OWY50WN/8"A*NOH9>2DS%)AB1(&UB8SX-5<T=@GVUB,^1D2E8
PBX7NP.@29&,7DWV(Q8+5\.G3N0B0@>?M=N;W<I6,BCW%L$-SW)DF-(JD7,#&*?C&
P!L= $#(]T$&A>=FBU"F[S24"='%I8R,N/TM'M$H1DC"%!R[#-A+R+KK&RD$5*%"B
PR^<SSW8CA ;#!7-VVWD]ZN&<(!LNK58N%X^]4QV?#;!N0[CC%OEW7!]-"US33>ZG
P\JBJ"I=0K/[(UO=:SE4&D-V7T)$[,#NN%K[".G'N.'65*O"I2@E!:=C#R;CU["_;
PQGK/"%5HKUT@]^I_O9.(WRVR^_L)@S"URG =2TKV.'A)/^C]G]D*E#R=N-H[/HR1
P(V-,"7C'?Y'W@";*@S\?DA)=<(2:/5!% _MQQ77N^!?Q!55"IX&N+@"F)H]2Y9-)
P]*<>IC[<V5@UAQ;\*R/ZX6-D373-W=4RW=*F0+AAUR[S^[<34_++R;HO0DS 4Z*3
P(1;/_$Y B%NI\15N1&+W/FO3/;FKM2,L6CF80R#G4WDOVQ F.RAPP_U0]/6SQ4^W
P:9Q=,9/X*,I8L_#I>G)J6Y@?'1HL\>YTA_CF68<X #U\4WP2/ZS$ /_&B.U-KT@]
PVS7?RWP D\A<@#MIN0!=,-4R8(-RKCGCHT["&@3$?HY^Y>0NG))*XF:TNRS#B-8B
P!V"*\AAY0$NMJCIB(W/;<F_2#ZKAZ)V:+O=+8#8@UJL?_VK9+F2ZXMY@=CV$WM9N
PVML?3WE!F)XDKW*T_F2;*(C5H:+5C(3Y1]@?-D_3,AC($]6[RL>F2Z=;R=C(1?G-
PGC>F9\N(X1C1]3W(G']S4JFKV8J(."^\7IP[)F*X;^( =)UM!J:8]G:Z]HI%/XR!
PVFNXX-*+2 ,]0Y=/BSX\NC['/KWQ1C>$N$N$,N>A"KX4<7&2U#ZN(&MSZC95'?Z#
PC <F/"N.P+$,8=,;%N%31BV#4N_\2N9VU"GQ?;73&*V&0DO%X'7[LH N9<UG]4K?
PQ;@>@\T,=JCS5=M4(LCFC2Z:%6+$SD8$AM7$9=#TYT8-'H;MQ(9449YB%J#O4_**
PO'5V;OV^DFCK?JKRU-@EHE_AHO'F$\.(P3_]XZ XGGS.)!@^?"^8P!>];[-)[F][
PCX\YY';G7WC:;NJXD3(Y:<)?=T=O,>"!Y45M85R7-I0AMU;E7'Q'U?,T3J1SJ5#K
PO:$S;VM#*9'ZF0O,!HOP5Y&3&7?(KU)'&A[E7*,9B8DJ.+!LRA1?D9+:EWL7@R]_
P3)*.O=U-HG $67 +\JRI[F/NNZ7QF960NS\5Q].^^G@M0.2M'69OJ]/EC?/(0-=L
P42;GPT=LNG*,5B;4!?40?M:"Y'PNKI:0,>Z!HT=A9B5#X<3K<#?V6MQ7^.24&!$4
P W;(#1Z(D+:?+*IZ2-/!)R.!N_4V@+IH(K3-,SV:07 [VGC]?E23$+Z _$?\).?M
P8ZKX99:D3/A.6=PZ.R?<(Y$P)?<\'^^9P2D,Y$*GS'RIGVE-R.LFSS:CHC+G80C.
P$R5^NPV<%>51>V5:BC>ZI3BB*@!\=3:#SEHQY1)T%+K@^:RS<5;:<1T4>N>=%#3X
P0-V=OAPS5K;.;XIO\#Y5% 3!'B?7USX<#^L2!W&.^"\#P^ <IXLKJG5W4Z0%SO6E
P@K>>&_29JI/V)U A8_B@W\5R=_<(\+$X9<5>94,M_-0C*;P:T5=<PP1?HPTHCM[>
P($2)M9L$4,+H; -V KB/E?X->X(_*<OY%G^3<]4+O^L!*I<QW(%$;H#*XFBA'(G2
P6G=A.MHG-I\<3!9)^N.M6%E9=7PR2]J2BAB!N&6!#7J*M-VOE:@FH*[%A"*&\R"3
PDK)>L"7N7+\DQ2?]4 L,W:'0I9Y'441UHR2F!W\LN@R_MI<8+[+/^>%9%9YO/Z^P
P<?45G^<Q3QK=!F8"@]77<*9U$^GSAL;<C8$<S@4R2/2J?$EG#C)4)T6]IF5GQ]D4
PMGLA8 ;)Z_;<O8+-DSMDMI:1+FSXO419+F4@Z!Y: DO\2G0;'V7+76;HHMG3=Q<+
PH]= RS[+?;#: SU@^>4C>3L)ZXM%NEZA((I6N16F,#5R%8]=ZC71Y#+R]A@CUAO[
PIM U_PT>JDCM24SL*+^X*V**L57890%0)EWR7E@R-C>^Q$<GR%7HF.\7J^L'1#3>
P8LVFH\E]ELE/.D]WC[2_],4HO'M9?'*[(X&<WN +D8+[G ^"K?PYG#;:O 2E*"*$
PU>)EE:BUKWV/]_3C=:J8)*CRR[)R57VVZH";>D4OP-&X@(P%(']9!ZT,,[FH;>..
P"=#'HD7><2E:48AUXMX#+.B"06!0O7$)OB]VD(77]Z1F8V+V.!+*^-\$1WP-$5\\
PWZ+!#'"KG:EJM-KB/(]WE'^7PRGA=O2]N-A&I!K>_M ]D6B#LQ6I0&F5_+U<\?Z\
P<*!!M!O:#+?,N'@TV19W%]I/<J)GVKNW_!#:TL#G[FOI2E"M^'L\T6EUQ::ZAR97
P[(6XR*BRG8?>EY&C2;G);<D4="1482FPE>Q@?3:;6+BI4U&M VR#]%BD;S&@=P7A
P%F&1QRZ>$;'THX&#:(+:^4M$*N87R@P1.3<545L,PM+ NEI0M")?E#POKV<M$J97
P3:E&;#@>EJ5"!JV",X!.=8TG\ @E_Q^K]!X$KX_(>..T\KA02^@(V>Z##9 29@)V
PXOW&\]^=DB&D\*U^$/4WS3&D4HFME8KCSY2R%IRN]U&7:9-:2^SS"T,1[@\?T[L2
PN_MS=/*;%\ZXB%WGFL4YNMK?DD>)U9'S(KUT Z%R/ WKQ^^IY2*?/0A1G=>E%/>-
P4,*&56J?^%;&;.CR,;E[/CU=L<!B?QZO&#^GNL_2)!V7EJ-)__AG+1:&W4?\NGK5
P)$%IV?@V4.<#S@%[G$B%^8^]K3V36@"8&IXP[3[XQDU'W(,U:/2MD)$H*0(2:@GS
PKQ][W)GT]<N#QUN@B&'XAIW\R_-[F0RWG[7^LDQ12CFIW!!,*&;7J?[QE5A Q\@$
PJRP&$RZ;P;.(-@H-5@,1,PYE87@#,,LD7E^L4+1L7V&)PL$0@3GC=Z4BTIX^$?YV
P^*T6.N2*Z @]K^TQ9]6^)$JX78#*Z2:%TBP)W!H=S-!9Q<#/-ST">C1,$9)D,+G$
P4-(Y$AV<NP :@&YV>^=8SIE_^_^(#YUXN=N]M/.@6P^*/XEC3F-3#$1BF];Y.W9*
P\)6Y?:4I]N3J)NR$B=#231&CED7].V,/B:Y,.RQN.^A)_Z%8J6___NPL=[(HY6Y?
PWF.640>?VDNI#(@BS&=1%E"Q>L">*&:@?UU:5C5X'HT)2C7,DM6WD5XTB+TVNB+0
P(URH]7/1!&DBBE#?CY>'V*7LE2 6YPCZ%YYE]]D,:"#@;!3HR#72TL3G^&X '=:\
PO*7J:-!Z)CN8MXNCW7;D]D%\H'$[$BU&H,8.+$"YLXS%M5+=%QI-XHMP.7ZY-=U@
P3JFOR[+$'WQ* TO",QT!/NJI$1,I)K5W.)&-"2)6-T3XLVRFV[$\>Z]_/1NR5&G3
P^K2V799"8U 3]0'ZF^',W/V;T4]9)=$<Q*F&F05I3,XZI!FUWOBFF6<D+5"?;?N.
P]%V7,D+,XQ$#ZST2#$CTO'5E]+0,=6/=/E-2]!+MS_GZ]<T,EVOZ:EASZNIU;,+ 
P_?&F&%DTKH/I.._DT(667ZT$;#/\%@O&HW$VT.;=B?F#6:_5LHI 0ES%I6(F]+(P
P@[-;PT->A1,;(Y.^?=B/ C.R:]V%/S[C7DTS',-XG'L_".*I)!!H7F,RG1T3JY*-
P]6/KHRT6T;\62+"XFKP>._;#)0;3ERT@3I)@7#PGA(Z/S(=G2D,9JO6*09K$L/BR
P5XY)8Q>IG/$P],XM!^" YV 1#*><HV@B8+H#Q,L*7C190"L610?E(30%7C9>GN..
P7F7K^WGMQMXBD@F:@-X?"CNJLL[+U/T5:WOGW4507[RG0I=5\"P?;Y/.\Y0E?]/Q
P$]&1E(C78"H;FUKO'(7.% 0_^8YNNZBE$.0:&$HEJ<W]'0AI9EMJ!GGKMPS4@XFU
P?!F7=SQQ@OBE"*T+9;=6@7_#PBZ]-EG960"E'VRV=5!B!O8" 7_UT@= B[0=(KCK
P6]%6 -+XVU<\E,\@7J)6HYL3[O@%JBZ]IS>,4%^79<03-J^GZ!0E@.D3?>4-5#"V
P,;*%11-N(6-S92^J*++A'!FR* 1[AK]$2T]$#SKN]N%+RX;9V+E6ZD)H81D75XYT
PCEF/#UY)ZC9FXX>GBA23H"-'JIN6A*A_Z=$C$;'OC>0NSVMB8] &,AB1@5H@2Q"Y
P7!S+3++>3\;"+_B:EM*(KX4XF!572V\D JC[T!1K,3$XEVH(\P</'+&@<>:)38;/
P*D%JQHL1#F&5J:<'Y=0L(S@$:Y7$-8OA1?= ]<Q1:*F]!EW6!9CJVLG1==ERQ=U1
PZK@$*,->H8DZ\#Z]@\AF&)B]*'GNV^XA#;CY <P+1G,* 5-I\YC0 J78A-'AG:F>
P"K3CIA14HM8SS0!PL+=)!7+YS_V_!T.&2G;^^L/IU[SN&_+[S,JFT7Z,!%K;" :L
PLO<84DR<J0$:<[CS#B%Y06O=71R5N<@ :\"L/^I^L<(%Y3]4/*@U7SKI&N-#I\6U
PLJX)_/Z?Y 1WO8):FS=I/ ;;7!N;!(!?'#<<&B-D=N=&4@DEN_/\[RC-LO4C)O6W
P/_*?/8L BE;TL2K'9"D>UL"_@1X:'H&&%/Z&TL9YZ%;H15 ]KNY1N'S& OO<#8P\
P$X5K#+Y2(G"]^Q<*5J#QFV@4<@$/:B:,*@?BA$_%<P@)1 O?A-#BZ>?6D]4;!]G@
PA?;W8:FJ5 4Y:,]PRM%ENO5*2%=+(;2B817/4V%:A!&,+3R.]X/XB9:W8O:9.NVH
P4HU@^J4#2-/3#1>5QWE_PD#<#@5$8@!DWXFXUIP_I;RKZYO#!?%P:Z9)$'T]^[@T
PV@@^.!JQU$R,4)PCTF&21<2WW%+AJ-S>IY+?9%D--XC5XS96S,1 1EXN":(4]0>@
P_LD'HR)!V$3E5SJOXS\??*M.^<GA:JW20765'@S,Q-+@*E#CYA:[7-TM%2D:4E+<
P$@#H#]&[0"EZ&XW!#G 9$?F"-_^<E-WU1P<P Y70;\P35"'PXW*X'-^/C%4.,KAH
P$#E/Y,/W]40Q%LBE>]6[;#)!D3H+=>*_,57H+KQUFB8M<OY/;EH$/$A.7#D!=?S/
P&XZYLN5#R(]!I<),^23;@ 86:HJ<^AP/..&=_Y;L3[SM5-O89EE/-)Z+\9%BT7DS
P^)7!L=CJZ&W]^SYTRV%_\+[G"? C@0=EF61:?JP^A!K;M%)=<8$1-1B =@Q=#;DY
P,,3D+5Z3C![!(5G>)WL1A#[KLU)!>V;GW,_-(L"J7,.J0-^6 V.WBO9><:4F6"FB
PJ/]>K]D;;K/=O=DM*UCWLPS2-VK D$FN+V+G6<25":,7B^D;;#<-G#!8NWPS 4\.
PD>X4#+6YP-\59V4/>KSK@<!0'MF['N4!X@J2JZ61#?R_'V'@Y7TFZ6ZV4?OY<3TQ
PHWJIV+$#F 9JBQ/'#RUK).;&J)3G$!H7\?@'98\%,4P!_$KXC$K,!8^K_@)0HA?'
P.H__RU(0(L*]<6#AT%KZF%KAQZ#!H2X?FZY\>&'*&Y:"J\%_> TEXEBD$\OAC0+.
PZ02N:= 3+F+)C1,9GWC(:5)6KO&L*-,;J4PI_.?< C.!U3ZD72I;7<0-#>Z;/3^1
P7J!81</'(ANB/,B;!F&,BZJ-\(+\Y/[PU:$ F5O9Z@B,IX]O*1MR0OQR8:W%SRLG
P).!=-5NB.S0S2.:^Z3]V"7N\911\M=RCG:R,L/>5AMB4&I?%8U!O7!HZS^@"W52R
PZDQDKD\^[)VXUJ7?Y='\+)\5#9$]?3L^H:]#QDGG(Q,MYWEWU(("#Q$:=HIZ?7M)
PYS(5+*:@_*4K1HKS$HN>P  -@W* T.=_K29)!RQ'?LB@S4-JQK#*.:KDQS"[V'23
P2+I/@@_?&&]T7>XC,%I3\-H@'+0-YPF>$5H!F#(HZUU@?]/&S8V-NN VYBN'77SN
P4TL^'H<]'B6*UZ@JG\)%&XJE1 2[CK$OR&I\)MD+S:(YH;+1#B6L^?8B[:'+K("^
P]%E^..CV\JJD=4(A3"(\9E;XV0O@N,C((H&?[W>BC)B%_^@(56.*Y1VHWG!FBV88
PWC ,)[@(]8VDJSL2WWM>M^WL8(_\/!8R_F7:)C<[_=I'IE'AP3L>J$N8O/],2'FM
P/)=^V&4JUGZ\-R".P@D[%15FR.G;!N*Y59CFY1X/%:,+.BG0J*0,\E9Q0;VY!R,A
P3C:8%]N?<UK;*]-=$K0#R#0)>7'P] KV>TE<\AOHB7.R5@0>XE2_I\]50;$5D[IU
P_PX;QE1**N18+1=[D%2:KI@<]AV?+ <XX0INPYK+A!?.]1Z$5K$GRSD)<UU_\Y][
PP3 R+,!C+_BLHQB00[Q'<IUCB%MWOK64=!0('%?U/LM?&J:GV%Y1^6U(F+$^^!>)
P3T^!WN#)F4#".(+\ET#VRN^DCS-K'A*WPOQB<;-J21"D:E=V*@.:3[5B(]+Q;1FM
PU''.0(#_PBL#9'%SFY:?>)!UR&2:T592/1@A7V>J(@*Q+N^=K_#7O_'WDRCTGBO1
P36/F,^YI-7;421 =N+JP'#8_[?#9\XL!@&'-I"N[9M;Z(^$483K&OV8\]/SJ;O*T
PTL@UH;#\T<%OTYCWD=9DI .V0AI1S6&'.^EPF[K<C97H=+NYYC*8L <&R:*$?0GT
P5B1*^7^3>)WC.APFP^5=#S/_;=GNVX/W7[<[9J0'=4G@R6ST8UBQ\/U5-?\6 85]
PY6Z6Y9E<[J,3*Y\ZV$69<M>'+HX(>-"]!@\LO+/O]8Q9'Q?(V]%DB6NRE6*^6\F*
P8+WZV/-WYS43%E@!5E?$HV\<'?Z+6#?_=7.F/X,@PTVJ*@?0?:1R9R<[+<X7V-P/
PL/V'V[DUJYLPM-7%\EJOY47E>/;6\"IJ2^OP00PV,0_C8TB3Q>+?Y;=?V9MT5P['
P-7UE@M;$@6(R4WNVV;YBZ2ZH@5M6<L#P,7_-OAY;,/<4=^*D:1#I?:&#JQI#Q__.
P2NSHZF)Z-QVWPVE7"CE)/_AN)\4#>?%=I^^&D !'^'5)G\E"9;/U4VV%7&5F':T>
P!9<'HRVL<JBXR1W*/7H>K9)0K^4#+/+Z^X&K,D=LOT_5>_JA(V=2#NQ2U+;.F$3*
P@UI Q)+HY3.:YS-V=^X7K 2UZ6K('OSQDH2=CLJ][ESO>G7S3:!46-1..SID:44O
P'"7;7JU 6MLR+FTR'GPD6_)SU=>IZ+^IWY9\4L"I+U,D(M:L?^6*8NJ8B$Z='UBR
P;5=AV%V+Y.>'A2VX7,&7VE 9U;O(+=U*V !'A\P7)SZC#4*!'!MS(8HGXXCTL"9J
PRPBA=(JPEV8S0)5:UT*WLJ$)8 6C#VI4=X?0C=F&X4%A)[19%^<'HZEG?#S\'&^Y
P8=-0)WMP/RV"I'  :IU55NDK=YL:*UKBLF%A9K )>5$-?* +;3:7R5=4/R5+G>4_
PUVX8\RWS&@ J@15BS,6*L(Y&):QZ:M2O:V>\P<2:8G4 U+T6TR%6'JCWM-HS(XUF
PKUW+'K<)MOR355>5"UZ4X[XP()/VWISO 8INWJY*4)#8R/N>"6\#,9JKT5(T?C(L
PFUA+4>6E:;_WT<U,%EF#E M$17%D&5E+IRK6*U[!P"1;1]7\HA3T,)A+]Y]6C#B*
P%7UH,B%.U9S&O(&]%?-3XU.-*^=??8 MPR3?D+P2Q6%S<4=KK.62!%D9[ N<AX<2
PI9$_P+15M^,_HSL>JZVWE[E]Y+8]]P@)GY[U).Z1_S6M#W>)B<F5I<QQ\42<"=),
PKF,E#OR/$?8+:&;5[[R'[:YZ9K4*-!$2&MK0=F.!\2S-#^0 '(DB[$)Q*'&97V#*
P)1]XY=) S:ICH;Q5P54.?L;DR8SAZ0Q^V"H:U2/JN(@.T8RC"=4AQNY7<55$<AP2
P+Q[_-7+^MG^H:44RMM7=E/A%N.VX1))#XQ 2)AM:E#Z98MCJ(D@%KP%>,^FO,$30
PP+0.KO&N)IJW \2N9NH!./PPM*%I/V$-Z2X=ZT7A9;>+NWF-R1&9T2\)'RB\I9? 
P'T?8X^<O'<2JY<;&H\P UWHVP\:R>@B9P=ESVBMF<3-)7ZV0GWX\I]N8?THV,K-S
P%4U4>$"*&S::U\F45G*8O0Y)KDVQ4T\UO!4U7@N)U0="'-:I(N$JENYA*XK2MT8K
PIXZ(K_!>C0A\1(6I"VP-%SCG3) 4J$P;UC]8T09Z!ED[R\U3D(Y-2"BX)=(QZAU 
P=I3M5Q_H2W/98NY6K$&BD:-1>O.T]2.5XP%=QD#X#8,<=[&B.,?&!$,GRF'IO"5(
PI)J*H_7K[I+UQ9S9XHOQH"RX)S_)N4_&#Q@$VDML0+9'[%+Z,T"WLLWA[-L(L@Z7
PR>NB-[]RE4!QS'B(@/5ZJZ/Q,GGY!1F A#IM=L53\NRB.>\>)(% +"OKU&-_^-RS
P5L PLG<B,;NJNFAJ8R"M0U]OQMC0EV0I^%(9F_YQCVF8)IW2CY+& DNO1'+XQ)W4
PA;4V!,(J]"*$<LI_'._Z9\2U)9#S5E!;-]YP_OR/F/8K4H$G_N1MS:CYLLL7*0*\
P$,3OYD%-2LK$5\"JAF+34 V7%-N:5T"H17T865\UKK'QW>K_FY&Q1U8%L$Z,6S#!
PWG2N_CY<X,5^YT')>TW_*;?+E>?-H90#HM-5A(#@?N>4CR#EK*W=5/*!*HWNR<LQ
PE6(TF+U#6<(107==M'N*H?"_2GIP0FN=='&5J!?X9R(1VF+[%V#S0IXLN*8,)A+K
PH>@(CBK"&;2H_R#\9UCLK2J&/WU,9LY8N'0])KAZQ<-N&YCTK%7^^G)2J_*V1M86
P1YZ6J@HCAH7W7P12;2\4DS=""&Y%Z<&;@SIAD?&<63B=??U.S<=*'?IM/AKRV0?.
P?6"VPY,=MH4MB 9G>EXS^]=6?+!H=NKC,&NO&=>"KHL':=BPT<)8;S_V*+[!(^YF
PCL*0NQ9)1VK*:/WQ/50M/8!8%''2E2.FJ(P9DE?KDS3A_A#E $>T]7V.>W[[2KNV
P H01[09XBYB!K76FS92Y.YF>,/F]S]XP1, >=+:1@[ (=%PU @+U!C-( 23LJJLL
PK::766I],#@!D??"N^'WIID0J^DP:>$B$U<3J(-IID],% .=-<79)Y54[F**#./U
P\6@C>^%6.*B:@DZ?#53K!G*T#&'%P],[L+!DLUU.()MC2[>=TU^EC2XH5Y%R2K&W
P:L\"G<P9V>4,C849N13MKT6,JS"I;SX^^8HYT']'94Y@55TKOQHQ=MMY\O]$]>"D
PNZ-.7?%<O41RAW*L 9,T=(&_YX[G]J+?/A&AU%[<>TZ7,4U#K'V HB%$N!PEI]9$
P_>"/YWQEO <_2_#3F,H3OE,$<\/OE X>],X-=8W"G837B?V6EOC?ED(/'C[">Y3T
P0IPNUWMLEL]KW8>B&JJU\3./=_)PW+MV5$\THXY0/JYFR>W<8?].GW*A46V+DAL3
P\FS(MQ'=*GFR_H@<RK8'L$VA=+L5F#T@2^1$#CB6E3#]Q!'*QU&O@)Z#E78#GN,!
PY@$&9HLE[^XBO9.,@$#PZ"M-H&5^+X+1[I-NS9[$U>.1+0N:S& ^=B.<8U2.*G.?
P))B/?' F&"ZM:(U_7M^Y13C0=E'[)NF /A18DX=]+;H"&8UC<$A633SJM7ZTMU'K
PUM%L]$>!O%]-UR=D3D5_.<1\ULF^[/Y5@J=]%Y9E\5U-]5%E<LF&6]>S @P0,R8!
P8#1VL<"9Z'"#=IND*:LVP:S:] YR%J$>GH(?O5@5BU8!0]JXXY%@9B*J#I[GZEGC
P]"M&_;\.5:RW8Q&Q=JI7V&K@>Q>6QQKV(RQ=BP>ANTT7Q=JZ0R8J,-F47I3U=_]3
P.(2(U4ST5(I*]L;2RP\\([_G)/A.*F--])TW"<LQ)K*!B_H;'GD+ TWDJJ!<G!=O
P@E-A=VMS51_=)1U6ZYX4<))N#Z9M$]?WL989H;!<)M7:O^7SYT6>!C?LD;C\XWM?
P+D3T4W5+3D6AEWJ:,R&NO@L3@@/B6%HH"=H"JAMOTJ?'+8OHM2Z,K7=V+W%U'.<*
P1AXE._+_8.?VCQB[C@/"%VCUD/T^FY^-') 2R'R4GV$;CT;9OY[&KF[Q]=Y9XH%7
P3*O@IQ%X + UWI*>5&V>4S<31,W$U:80T:8OSIHLG 7C;[?O)+BZ8GV*(4T!)59X
P!X<#<W[)8M1-N+NXK^$@Y)8S;O+V=Y<SS($?Q(,YQG<9D7N;\55[NP*6W==X5U&(
P491.<(3A7//BY)_)0F3:5$=BHYA.288R+>.45E#=ZX $/"35:2F\^%FX9'\(Z[$ 
PWHXW+5>2IL.)Q&Z2%DPS$="DNFQ@,%5?D81X1^()3Z9R'SY'@&K+\\-%N!B&.P_2
P_JQK%!Q-K62Q+99E11YI/JHFSK1LLE+?=$<*3B?ZY%$J?/9?M&O6FK6_*YKD51G0
P>Q/]6;'*[)/_L;;MUY6V8,T,FTZWLGGA#G"OC+5-8*H)M019YBN/%!@>T+GK7?G%
P?$BL69O+^FEZFW(I#Z9.DY%/('9B*C*.7'NC$#._RXG[MB41<^?]A)C&P2CO]3^L
P!QK1!+KD/B^^SGP-?&/Q:];B65-O\'&(/-?\#*Z29\(3O0%Q-YW78]>E4_T\%V)Q
P8HEON@<",\49\8I>DB\)=LRC-('7.9F7"0I^(!WPX12Z\+-9D'"?29.5LB!^@NV0
P=,Q]X1Y6."\T#K725#=UNT<OT$%'Y8D-UXAX2UH"?0<%M*_&0/AG_A[2A8(?O_E<
P&="B_!CNHL72_R=64G;N(Z<9;S>RV@+)(*A=+I::622%C@!KWM,R;M&,IEBM1O\5
PZKC4?>)DO[*&MCJ[;*T0I3F.E^_:'Z/&=Q]C,4*Q/)462D#CK,3>0O3=(!G#PM1W
PT2U7N9&\*?XW'U0.;@&]@ H/P-D.Y%6Q$#+ .29Z4KCHTF6^\(&MG9=NAH27U]P*
PH*)X'X-#;/?R$7D8N7@@E81V6QG^V$GBT<TIM$H.'T_MX*2*Q=CJ@=?=*O?VOY8%
PX%V.W/ :$PSN7@[(8@-X.#Y&'YB.GI90>[A;2?R-).E+P]DW1PG7)^_TQTIN',].
P$/]13,'9!)X-"2<]9+C/"";176[2S2HB4!.X2F&-J8(QC)9V&WY7B;+Z^>"Y@817
P[#\V8;XK?Y$WZX;Z@FOR7L:6<+\_O*%Y1I_AS 7F%6_>]-S7_9H0:MLR'AGX=MJC
P\@RB'CR2'? T66>>HA/C^3A<Q9W5._H_MRD_.)0=( +^1G*1*E9^-]QBPPU@UF@Z
PE-/PKRNS>T!+XB0 *Y2[1?&C9*2@J0R2;+PEB41PT<^N[!?)J+'A$BH<F3[HY3_9
PRNR'3^EU>[4FR<V<Q1%ZW-<N:;?J!1*$_!KL-8%,K8'P;=C,><5Y+AOII.>D3VP6
PAVC'>HA=!_AT7GEFPW[XLW\9DG/H47.H@CL70;'E@:^UPZ[8Y0UW]><^VCMB/5?B
P'Q0^DS;0#;JP"3D%K(AU?Y*"!>$K)S>II@;!S@_$A0$FG@PK@E\&OPE\G4[4UH/\
PN59 RHJJ$H[Q8TY]F*<&S8I%#'4X; 8);U!O*N6ZYB+, 5(@\ =!X&_1)R#HFHM*
P[7Y:)B=OY=[!;:B]GC>(!=EQ#IYTW:<Q\)X:98@K'"6?0F2C'J/HI&+89][JD(#A
P)&+Z=%5&K04W3KXM5D X7:<\\1KQOM9&J\)R!W\K)9<L3(=0!"WU-9FE1E9'Z1$]
P^-$QK99.;Y\TMJ=G?+T)+G6*]=CA 4-0B,YNZ$',HT.8VWV@]@0UNO!7GTN0A,&#
P1#QFX&0KV@1YARS#+^O$+03\#?-E2H^1S=-Y'%_O"8A>)6(VI94BUPII<W;Z:9G 
P?)K2RL<QA]O;\;9$H#-0;SX)L,XK12+:9TF<B"ODBUGM<O1P]*H^23%:YHR$:_M5
PA(Y]IH"(T3'; M&R6?NL)K8)C%Y)I1(WGE,7?V;50FD.Q1 JD$?Y[RZ(^$E95Y?"
P"HR\AE:]!JT#NR=.M?*:HW7\PODE7O.NX,"5B)<"3J"X E-]_.?406&D."2U+6T$
PSY:<@;J^X:)QSR,AWFP+S!49;<@L=YGXQK"4#V79O5W^]:7:AW/M]B<VT@WG&MDJ
P=;BE6#I!MDKLA(!@':+^J4EWJ=!OCY5#>CLZ)&&! 1/:RUW3.^/Q89FL-H5-G1/D
P(YJ&8M4=D5JYBVB,W"-7KP)/Z3I/!P\FD;/=?E261[7M<$MW'"2&$2Y4\R'V,3N_
PE25K0I-+=E2?$/4Q_1Q,(@!*D=GV$9:YG']V[2!#6JCE+E"[VN?571\=6/[LR]M*
PTP=O:<A#_%=7 I8?8 [3!>C"R3F\!/)\YW8@Q#*+X% B7?&+W%C0PE@&P&Z?<7VL
P$T2)*QH?_-3W@-JEP:/?.BWN4(A +NL))F"&7C"IG^.&=9VT-$2X%.*?/4%.TZI'
P42G_RS&\B$Y^\2W-.SVS&$_C&9!7P" @29!Y??%_F*YQ#_2*A/^.]<YYVL.\?H)A
PLGNTQ=6MJ)L(#IZ3 +^N[0YF@;C?>"CB+#B$V OET>I8D2M3;<#/.@7"S<:519BU
P24^'TH7GT[7<FE-"?/NIO0P2\BE=_LX_V],AA ?"ME-1JY[UO<U:;&?6];;JF%6_
PN^VX6:C GN5!O(@9%8T%DG;K9RYK-BMN77F*2=S,?7.4N9.''B3IL% XRZBT6YDL
P-ST/D*Q36(_72@=)BJ<(A"%F4V^HWN)#6EFM<X,U./N]7S7M>+? ,V<)9_Z-. !S
PBMW=R7^]+Q*%VK;7<=/BD5.&)C75G2<ZT]-08>%7Z%[8LIU/GW5,X$UUV1D:KH1=
PL47GJ=VF6/SQ0:QP]FC'Q[V.NK.A!1;XCX)<[N]<HLNRW(M+VC?HR<\![\>J?/@<
PCVG@U^X.)]SI,ZE]FV$A0_E$) !Z3:(MQ)4&?A6 -H!Z6_8%K?0=!9%T?WA,""EK
P'#8L\AW_X7.'&<]6WUC\S@5D8 *L<K^D8ZVJ58S)*<TXUD8\>#& &%U[CJD?%R@O
P[H(H=H3OUX8V3P64D?F36H?7+?3D&P._P<H&=L2.D6W2PRT9S?XR"8JTW_EE\A>U
PY4X"WE-:'RE]O-&VGMTCT7LIU<AS'QHDIL4#:G#\2Q^'QFVI@M ;2#W(K8%T/1J$
PWGHT3CT1T!M_P8+5B?N7-#F5%+$WRU-9!RV:<Z6EQ3G+3=R[_4.A=L&L4TJW\=6,
P:".UL[UN]\^UC/?D WLVI&[BX6Z,+H8<F6 VJ0AS[I5A$)K9IE#XE,0[@;(IB@X-
P)A(53]=<HG.0J",0 !NKTK>#]/(B(TZ+!TN39DBGT6"I7X\5R5^V=MV=IQIH#XLX
P(0[Q+,!A=O-9;$9*O) ]+F$^$JU;4P;X5STNL7F*9"JQK7)R<0P$Q>'^U(_U?&YZ
P$5#J,4AHCG=28AIT37+D"&@R0$@XV$C'5/')RUV\,%AG'<?S%HCR-;UHHE'\5=EP
PDR[Q;MF+(>3RC95@_NU2\V<IC/ ];R[(3E&\<=B8SY_%?/F:IO5 -5RWQ7C>I!OO
P.0(_<2%S24XSHI_H]WB->@#[ZDP&(@J/ET#^W)[6*K9]3C#HA3BAL><3_'YJ6]6T
P!8P"AXQHCU)#-9L9#^W.W[E[%>[S1T[3/GQL<@N(WV=-:QC+6#57<0.OB,P <1&?
PT;5^W7$H^$7< ]3=-/_& ;0S3^*=RCU^U@#QXO><Z]FEYR0<O^(V>I?64(KU&/3>
PMPG 6LFF!_^#CQG0RQ4#TQ$Q"/(I6TDQM.B*WR!Z#5E^).X$AFD+=9]+I&)):@*9
P$*P==!9&<2'<@++Q/3!*0A$8%_'X,GCYJUX%S]_&O-K2PPF8MM25PF=+@*AY)_0Z
PL[6/?0$Y#N<A@+:'AYG$4(_2T3E')V+R#[3U7H+4P\H:AH3BT0)(J4_$)O(Y"M7M
P7?Y:RZ&5V4-D_=P#G_\J9#=>*I<6I^ #]R:/+/NN$59R_,<[JKW(/B0[.W(].5]Z
P.\&6K&.8YI9L; XHON"&S2#:_;:=5]X.>0P>OR\@#;GY=B\KH]-1A8$W!O;G^56_
PG8'&5EML^"N<0-N6DQZ5T[V^KW['M1G2.$Y.#!1SLO/1;O^/_7P8ZG"?9PR!B0EP
PG)MV)I0RRZC[02Z/@O5D]K";1BY:]#ZG9[!(0[F!I81RI0K^MI78MM"(FWRF9G88
P#D4,B!<0HH-A]68T^(Z/(_B+A$:GIWN-F4 J\4HB.:;A.D9G!S+E)=[0XX=4L7U+
PTP,IY8=+/%5@Q#<L45!Q:] J;ZV$5AB00> >+],.QE<(9QS5_B36S%"JQT)U>>P\
PXXH(L\1Z8Y@A08 ATA,TD>A#74'2>N363^CUS6W J,!4/2_)(-7?!FG6#;E]&0E6
P&.D,RZJ+=TB5EF0DNDYO JDIW\-;3D"\A;XKSH+:N\1##HLUF)XCO*JF?D444<SA
P1\?TAWS[WF(E#GZ6S43P2,*;,+V-,AA.2H1O$#[O3(&KSQXO77)6SR,<I? <>#)Q
P@5AZA0@HJ)3Y/"J=S1'0*+)4O[HVQ)SF!!BFZL<?6MH7-?I@*E'D\L1!4 /EBIRE
PR0T* KGH![+H37I$/KAD3>,F!XD^YY"01J5N14NA^&O"8%0/6Q$+%EH.55E7-/$<
P?/4++#8TQX/%F:1VQWE%?0#"PIO+!I',^Y"B4S!"?*>(:@*4$I#450F^J=RW^ W(
P]23-.V!BD>U>B; A>&Z=-'/\HJC\8G-[4&6MY,9\4TT#\I8+,D'W!@!27H_\V;4&
PE4KM=A\8"9K%^;83R4M.D+!"JQ9C-2K<+_('R=5)+P$'89QD.?BNFS0; RV!N)+:
PC63QN:/_Z0M31I/\1_NL>O423R[H$JTJ /5>1GN#BHH:V^[8'CM=#O"3)E,JMZH$
P#:UU";3Y0S6N5M<\!_5RG76.7K\4S:&]\UQ:\\8S?-Q+RJQ/OT_>#_&!<[ZBK^"<
P1ZB+RI,1;BDC!R2-8(4M;&:!H-@C&GOFFF?9X(=:^;NY=QC>M9A,K&G2HV7SYZ0.
PX8$7IW&)U/T8W4V:P:.>4K\22R].2]G7DXLX1?I&R]14:K6=AN:SI_H][E]?506S
P0C,:1;/#QQ#G.?7<#<)(M"QC2?.*T/]DF]&FH1,6]8"1ARD5.D8<82ZY(:09[U??
P*EXFY]41!3Y?ZPC2^W>E;U[T0((24E5UG+!QO%+O-($#<?V?1MV'V,=/9D#=*<"X
P&==LZG2GCPX?"S\&\<4#_HMYO-RDZ^_NEUSO[P]4D*<_L#O"T8NID45U4Y6KLK;+
P%JWWAY+)^HS!MB]ZJR('9)8L-1T"0>9:XXH_0EWB18$$HOJ1UP@C'&^*A*5F<J*I
P#"[K@4V8+#A4=8>G/UK]TU&$C_@9RZ9K!U^:(62PS*T2 Z%TR,@T-:Z\8.N>9NDG
PK] @" LACH <5<X_?<XSO?B[ZX%?RU5O%7QFJ!LK]>\9ZKX@H;Z\4KO\<S:8UE4<
PA820R7;5Q$ U>WG'J/CV\'UA.$?LLEAM%K6LMG# ;]I9^ %?B>-1/2,7:<RAX**O
P,PI^%:LSS5#Y=MXU1Z'^GK"2* ?U @WE/F^Y( N%D+N16)I:>(_&3V6[,7_V7YU%
PKGZP[2.LN5C6YRCX-),WT48_!291%!66Y N^2=86 S:[%\'ZJG48CC=R,\IRS*A8
P(MP/DO%635:8]XV,V_B+%!:\YJEND2J#7C>%V6 B5 V*=KNQ2$QBRCVZN0/ZT+R2
P$:CP?Y'A=%:\DM-,E0-1Z$A(7UJT1I)239"1$/5_S=9B(B2J];GC25 XF9I?-9N8
P5)I4CZQ;<+HQE@!?_\II?@RY%C?!\6WT79+>B(#FY<@@GL&D)SUB+)3[R ]BMA2D
PJ%,7O<DI"$TL[@%5';/!RH^R8K\VN&OP_;/$\+UQY=T@VM%C!ORK;F.O%();O6JD
P@# 4.+A7-H;-PBAPB;/A(#TX<KSQDY5RT#7:F610-D*UBAK/V=,Y0CR52>Y9T<^D
P$8(<X=V=#47TN>JRU6[H<+9F,H9F18&O$'MR4'R3ADU^K"'S" $3TK$/IC$"#;4*
PIVC*,Y;.JLX+YOZB;3-U27AFU6%3#V?I8AM4A[Z9H+L=7TR+]H4EK&PYA+SZ.@,/
P1I 66WKE33!3[@7O 8Y9(O38.;S1[[[MV!Z57C(!CB(2RF'."';2_T.TLDL'I"PV
P,L7'BY#.$>B".QSY5O_<Q=O% (=?RS':3E1,@\:Y'<MY<2-DL\I36H>JDV2J[-!T
P N-P(Y!7U,Q"3#^57P_7;V)) /*"J(K@+=<JS:\7T@IF3 \O"E#L?CA4UN5^V/Y(
PT&4KW]VO5X"SZS'#5I'SU>#]^FV'DPI;8_<?U'OE<F]&!D\ <#WW8ML\(W3R=-<>
PZV $]\)>#>8/$2@";I(&$2EA6HH<"49*/2X4/Z2;'IHYND'=R,22X\GM>,M>0J<D
P[?I59U1$!('B<60ZBGV0_>HP3^,IQ7!I>8D.[4OF3W=50=(4G?+SH&7![I'#B'OK
PXE<U"$8\A\Q4W^'WK&D+_D!%FCW3@2A7._\JL.FA5]X =KLEB'E@7!@>' M1IDBE
P+DBM\%4[O#:-]@@S"UU#N3Q8)V7NYX[-!1L?I'ZA_=2A4SSMCNCERV<G@P_0;DWF
P7H$9H_)(EQA1UL27)G_'0>W&%5?4%U>%1*"$>=I1@_D-LOM.S2R@/8FI'NX=\AE9
PTEO\31S-J1Z)("N: %&'+;UQO?]/D>PS%Y*[*<<NHH[G\.7S637E=-F-EN0Q3.?M
PM\F^CRPY>4"CUTL[IJKO>OU^ W"4PD>'%>B<@?1"B.4A\F?M&T)AT[NZ_MU>HL#[
P3;*>'@W67WO #M' *I#$<&%=34\F"B,(+,H^19\;;RG+C!HG_P63P9)@6L:RW,E$
P(ZB:_OI&L$KZ;-3R-:O)2B*2QFW/\5&2;@+54ZE&YM<V.HJ2)F[Y=& )YW]35P]Z
P-Z!H6/&A'<I:7P?@["OCL9Z#@[[6)HZ(W^B!?C9^W9,MKUV9Q1R5Q<PP7G-7<  ,
P'$Y8$N=AB2MI3PW[V*H\\N+?UN,NU0;P^,-:&8E%]7L^?H*<WPOWN4.D]!+O8V=O
P::Y%<E%L&"9RP/=?@,_N3S7&V#]C<73SYDW)KZ B9ER! \4V.+OGJHZ6D6A(\ZH?
P&8LU)5!>:8'S')MU(6>E'KGWZ"DOYY[A>[\,FCK^">Q.-6^L*A#7HVA'-(BQ6?(3
P0\GI5]9.@VQ*@0H?AS)-/)D6=7G* (L]5Y<RW&_'/DP=[)?[VU,;B59*,5R!9904
PA'5U>A=:1J%2!M15I#;RT1U/CXNB]%S6%7;U.\FU?@9H 0=/<CKW,R?'[/[:LRK+
PT&3ZBIAJ9K("4FY'QH/WE .)$>_S)V"!Y!1)E< VH#)S'BC5EN)#NOI:364.W,V 
PFJ8L7?>N+LM5>1 -Y+!EF/4PX'1L=V<?%610+D4BX)<^+S W14BXRY7IN%5"!! E
P.QE9!X#/BH$GJ&TTUS M*71Z+]%)L%N<)#^2ECV[)S-VHND9=;DAP)&%4W 5XZW'
P/8DD52'+>J[JC0(QYC=G!I,/>2&SXT3Z33& &\NYN/9,Z]KW1:=K.\*I/JB'P?BV
PL0W(XOUK(E]X HE#I'G#;@KFJ3;[3ZO Z2?6B6HH EQ.J&_5CR;]<O(\83B=AJ<?
PZ9LQ R(OZ'[#E7?Q?M<X!0H>NI^@]),.DI<EXM5IG'/8=,,S@S'>1W(E[JV+*A/G
P^'Y\]J<(U8 LT''6'JS=DT!IP0S\XV+U!>>ZOS-CMM0UZ0"5M")O8T+(@0K -G&?
P_S?EX;[CSNG;+'I*ADL,:?J;#+1>]3Z.EXND]I#(P28A*-U) ^"(&@?E8F(=Y,V!
P*CDY4$Q\4.5X#S%YU!N+R+3=Y\WQ2?"SBA&3;5X/VVF8*\0K1^G/H[L\;5K1HY,<
PT)>'<]&/FUACGCF:P>P,I[^/E6J9VM(BBO=XAFFZM3AQ?)*&5;):/LC!:60;N B_
P[ZW88NKAG T>V(6N"PUD5# KD&JV*;I\?<XX3IQ11AX93YCW.'H/R8*:-! @3B3,
P3$/7A0/2L*>J9M@W3:HZO#@HU3*V-BQB+^/.1MO6: MB]1Y5OQ64^7M/C]J6? -:
P1<N* K(9R]RNG)&%!9=" 5'^OAG<4JO8BLKMR OYMM<=5K]!\;I;9!Q7=!DP OO]
P:PF8'/GUUE'7V_!Y/(FT;$]>%J^UF[HP8:@=R[ZV2<=6_OQ-3V26<(UL88^,<<1W
P=*XGV#""JX"<Y>'A<"^@0HG X7K]4 3B73>;T=/^<_GOK/)*W#EG?!+QV/I:[8A(
P3>#0J\D=&L(O?']G4B1XNY^;]_.BV!H"/]$4_^K]7=0O]W\F%#7R-_37L5V+5BHR
PK4C.7)>F)3>V@4%?";FRUCAV.A?+WB2EV.SY)/HOX )PE[N:)YF:S\U43V4<SR.1
P,(Y[96J*9(AW?5"AV-IZ@#H4/FQW-VK),78B(='OF5$V2'LWJY7.?T+DWRW<1<N9
P%BO6:\<BX'O@<#"8>D[N*8+7$,L*%>PZ1I <?V4R"0HT/C$.086(*:4.7 D?ZN>3
P=HBC+[\R^)2Z8'9IK*%->#4$[<V1M:2)= 02T: 3G35 T;U/G@.&^K,6DKHM#:))
PD&#P+:2(.R7@@MSJ?OOMUCIQH7LI"I9(G$!+ <C9"U^^W^+"%1CQKJ0:(0/<?EID
PO&IV*ZK8Q4A]15@_R9\Z_L9LL,+:CTKN7RTA8O0@[32UF1Q6WB9Y?WMM)6>#Y"KQ
P[Z>?FC!,7?W<2MC5_.U>@>'8!S(&>T:J3RV)CGIA)&+4KS78A-[32T6['>F?0F0Y
P%0NS, %K$<+9.Q_M 9FV-5]-S)T7'-Z[)\8)JV;KJPS)=A@=8TP6BH%*?<]&>M%%
P>2X6&$/++%ZAXRG?Y)W*@^&*AW(DB0&A#A(:3SS69="C[6>H2H++)_\B19I67G4X
P<0P"=V&'K^#\]'%HBONSK/K:^GO748U.U7"PR!)F7+CS1&_*Y6E82$,%+#69[L!;
P$H,;C$>3*?N>WV&*(F\ 3X+MLA_[_8/9"5'?^&7" OB$$^9:9=6>T@D+%P#&9A) 
P0\@_[P,D?0RXTE0ZH1Q(XI[^&TNZR.KT**W<VH/K,;H!HT\HWUG$VRE<EYX3FH$J
P(^GOP>_'*K4+F(QGAPE.WOGRA*;?L* :Z!H<YLX1?5T5BK=D;/E1D2S G-C&=L[,
P0=D+$#KZH/^?Z=[2==W1FTG!A=3X*'[=^;7W'CD9^MR#/[_9]: 8K[]RXP!=T),B
PLE3OJV+6D&ZW1B_  ]6Q.PZWE=5(Z.(_5Y$M<()M;L5(N\*(4LBF7/H94!H2ESH#
P-P 5%,,Y>^C-E-*%@4"%C'GWGTO\1SZ3,17A[P20PC\Z//;A&P6%ZL)\[II[=!VG
PSF$N<$KG_B;V1YO'NUQ#EMB7S$&LX_O]J($8JF3<1S]8F#XW.;V?3P+^6)-,$6 7
PS0.Q$LD'JV) FC*2+"Q'EFL)JP4Y*U9^#\<^@?>JS3F3KWH#@&MBG)MFL]@:,_6#
P:,WPK8V\4H+((:E*TH 4S4(>(@RA2>^V,>ON&3R*:L%7PS)L*C5,L8)[.+K!PR\X
P4*;8CP4A']#=2^R*IT.2 +OK%2DI'NJ+T(RI=W+U]A[6'@)CD,%O='!3:[_27+ 0
PZ W(LZNCLV/5<8FRFOQUZUF*\0K_08"/18^++>J7T#]Y!.@B]VTIZ1Y*G-EVL5EC
PR.Q_X.GMX*1'6C*/@<6E>F/:DTE'PVP]Y5)OM2D9=A+Z!?&E-EY@4?C?%HXJ0#WO
PR>4KV]!GTC?__QJ@PI<H-0FLU02L1Z\1-G["8]<-@:-S7LHEG7P":_RX P3*FL$Z
P4=SH@%50V>IX[)08&45NBK,J<!"O"G9B ^@'N]7<UA1I:[O)S04DC&_<%FJ,-?UP
PZ=^1!WHPF/2TO]SXO>.JZ*F/!=1EF%6"*BMAK51!/VP! BF@U^D^EM8//%@$&"2S
P MF@.PS?7:6UVOLS3LSK)=(K9X4WG$15V=KH9^IG';>\L_;C!11];,)B9+W](J".
P[GN[^D?HZ\WLC^0)4LA- EQO^\[]QIH?\R^,N(!>6CL /.5?T5-5SI_DE;J8T>PL
P%6KB7WAP[C$R1R\;D]H[$I?0LS!AR ]5G/RL!!H4MMOLOP-_(8L\,JR8KK)O<%+%
PR+)S8VX> ]-#_92Z3J(R,.+3$R]/OH=!N;0D^>(!XFIUU%.3& G*QB4I4SJQ?XC/
P#D+N6OEX >;,TW$^!L%<$8)N\W+?5P9PB!J@UQAAJ-MI74V<-L19BGL"V2;'=MR[
PG2LJ3@QT;DE$GB,UVWYZO9>J[<-"W7C>#J.&+!5F*5*WR#F'UX[1=UMHTX&>6D0D
P8F!U"$X]/O9L@>2 PW2DS?BJ+=9)HY14TT&_EQE22?LM(/SA7-"HOY7%6TX3^\-?
P1LGD0@B@JD4RCU)I@!3\;+-12<<88P]?);S@>53JO^O<V<[+KVX)/D]<O;PN;.Q%
P(QR1S< LRWQ4U;6L/W,#03IRG50WY)P"]2BY),_Y4RP9'<N8AZ9/M8F4-V8@]_$G
PZ!@-D/0K%+O>IYLC,S>+Y!3)V_KD5"(!?/B0IPNQ(H !SU U=FO9'B6XT+ZFB9Q@
PU(Q9+D+4Z,N;H"M'%VY_<N]4Q$<BQQ9C81"<%Z@M[QHY/O&V,NV]&_?SR"U@:[E]
P>V8HG !MBER![*K=<\T> ?KTY2^(CN6N[JDB%U,6N;P@8#K9YR'DXZE_)DX]%I%_
P\TO^/I:9C0MD*(=CMS](N<>!U=+#1&9;'7]>DL]EV_T4W"%NST;65".K8=6^>[TP
P=IISH;OSEP ? VK%Z=ICL6BFM05)@',23,*!$&&9_ Q='8W B__^P0)'([7G3E$^
PG[]7X[ X':J0Y#V7/(D&JO*U^V]U)G#I4>)'>E?H+WJB'.L[3HJ$HKSMD635L:JK
P]XYN#S^J,7^^FLGH-/,CE3D!V%?JKPZ,:EP#(P[&"/-!/XBGC"<<D?K6#^5D_N1!
P5./%)!K,% ?WFET;@P")TW_WC L*8N*P\YU1#IFV> QUH J(0Z-$6<06+)H_/_P3
PX3*I,_EZ%"DSDB:P?Z^G$;9^(?@58$.U3V,GUC>!@@AQ5?XQ!A!Y !&"J:,,LQ\G
PRW*W5B CJLEOI"G0T"H),RY':A[@:%#5Y[M853YIHF0L8H"3? EYBK5MD'(-:?/P
P94,JG,H7K(A_P0P!1(MGB[ID$2B\>X!^![JRK^U9]Z*>FPA7&_[@W"B,!PZT'CC@
P<?V3I6U>*(%C@^#(('H11O\7HH:'DAI2BBU-?+2PGVC:FPCM;$M:K; $)X8EOJ[V
PO-<&?BJA!70W,:[2EJ6JM4/TB>%;B-G[\B. -+:L%2$>Q>N!A)4.N%G196H4 ^:?
P+@IHE^V?CSK!(W9SE9+_+5]GC>! \C'T:D A?$^%N:=GG%QWI >PDQ!&U<#^:ZIB
PD'PB]L#>5C=!X^=1-_(1;%&9'+ZSK)/F%(EH9Y8%40KBH$?35+>*2: 2C]B^4.P:
PX8Y9'8/;:LW9Y-SCBB!? SIF XR7"%"OL@K7HZ'2WFR!,^X P<R4S<& .V45)FV'
PO1 *XX,ELIJ.[W;1JZ;0\4Z:N9"+QB$DY<@5.<$^[SI7A;N@-IU$&AJMGB4OV*B/
P^84#IR=J3O!X4Z6+M@!@RU1_MILA: /+'WXQ#>LS#0XV>4>A'M<6*H/X<^4(*8HA
PR<Q4)$,@<?]'UO?FEO 3^(>&$I'AXHEYVTHNE1>5!%^:''D=]4//_4[K1^@WA^<2
PE 'UR+&&Y)T*9WW;F4HCIPFVD/RL".:BI2%H$5<P:=/LZ)O9Q[.*P#Y36)$M)+##
PH$^DCB;.B>#IK_X8U,Q.$%%5I]QB(J8,\D.?U5=!)?>"!#V0JRAZ\S A6BQ30)L:
P9"5T+LM4EU8\@!CX&"^XO!YBG>]N3@__/?_/>J#=#.HA7^U"#2%A"ECYAB_)68_!
PG@R2(>2M/F-[\L/V2K&,VYIY214<T*#1\V=;$FQ9CE#'3%1M&HP!O6#: GAX/_Q=
PJERDS(9Z<N9*G1/2<RFS*Y$G"%RGZ'7A H!2A,HL#B)$^?/,7P N$6NG$:HT2+=<
PJ.F5 )6G)AO<,;!J\**)*BVY>_B]I47*&,CJXA'/N2'V<IK6(HC@^?2 64RY;KS5
P#\S35ILH<;0[5S8C>#BTR,C%-?P6:W"NTLGGR/CE0ZJDH\9_KI<@U?I3H#\WD;AW
P4AX"9PE3JS=TJB,/[&?00420N)#TY^A_063"HQD9KUD^[(6@JL.FOF"Y9 UTD1.?
P<-Z20E6!I933@. 2>T4H-CP"?LH%)V3*V004 IHC@1("C7Z=H:69LZ[5RTY5=!I<
P:?-Y83RSZQ?(0CY_B]ZM?WF[8GK9ZTD?MO!  +&'V[T6024]-A>I\ Z"4%E4%A#O
PF9OG>7C7T@8D.( K"=%OIL5%5,?9@'(O"$WEYBUN'G?Y7*%LX3_XOLF-"YO0$F'5
PG[96CHT!A.6,ZJS./65KE)UN A_$9 !S$O%-$'U2+4)U+TQ)EF(9F/)P2E[<YV/0
PH0LH]G<WNPPZ2PV_D\FI1#LP=C:/?])K%5N'R4@J^'P/\YJT0F&2R?H?SC89.2AH
PNQN,XR<,_9[./A1&GH;?+05]SONQ_%B@=342CAE.EG6J&&M9\PP[%C[*KFP(UJ!Z
PGP*$#7";J*VA>:&_H+W+1!.R.S9$JBLJY,4I$?L@37[,9"(=PHZO(.NT%HRO_J\Z
P86ZS,,=M[<&!F=!]^"-@+@!U04 8:Q$S/&Y#N&$%=4Y"GASHE]0Y>;4];O%@G&WF
PZL! [N=N3,Q<5D9ESL_$05%1].EI-3_X*.,OF"&.XA@,(C;*<RV_O&<X:-(;,<G3
PZ3 +#*<JH8[4"9'C?6^-EC$51XW(-9!]F0A'(O$^":F6"="X>0"D ,^4-V*U-:;R
PPO>C:,T@V=XSL9>9WOXJF62^N'M;SY!:I0=<"?O5FYN0U$!(=5QU0F$J:IWW(WE3
P!6V1N&]D8KI/$;S_N0QV/C^APLV VS'<WRKN0%WG+HF#+A]!!^#2A=-FT*HG&,UM
P#))UP)@MNP[!M0S-%QAV>[]_H1X&GF;3,#'TT>5.KDCV/B\I*.I!K8DJ@N9TOT;/
PYXSM3=/+-M[NHZ^A.4N#YA$2/,S!]M#,-O.&3RG6I8?%8B1O(6DG2A<VYBL>CU7G
PTEH<^<RKY<7WG!MPF;VFTF/<JYP#_7J>%==_-4*<)^'=@ZJS CFH,_9T.=ANCA2H
PU8D<M07@U2!>TM_2=K_JB,!'MVQYBK5_>C-B=1=(XD-,',<1Y/XM>1Q20XYMJ-!M
PT A[^#PO\H58OXSG?:D&8J&-EN>7)8)>^D(G>GA$3Z4>S*P0,N-^U!L.(7HI<@)C
P:"7OV@AK&\/P]XI*'L?ZGV(LNE4$A8PJ(M1F>']<;9MO-J]OGU(D_F]MZ,^L7>3(
PC,E8O^-A.-$MA[(JFLL014$TY. OW.@C#3=70A8,1)[*FH98(H@B[W8J6!4?_&VE
PL26<&"HJA$%1"L::9;CRZRV\&O$!YH4K!,S(HWY$2RV>K"B0(EKCBOJ]I4,M',"G
P*S/')@Y.%K=^@;"4X+QBY.0QIH2X^HFV.K 2VL<\#P3RD4@T4&.!X'J,@/#:45O 
P /ZE%CJ/TM_>RCLGGEQ+6=-ADP#7"'>FQ2L1:C3.$NQ>A9.Q86T2\/718D"5&8SQ
PAEUT*A)GHLD=WU]J]Z<;PJ+,<+<+NS9ZY*(4HIDPS6-XU37G@FQQU+Y'&P7H&,,,
PBB:AV>V_JB6>1(QW\9XOXN2*PE_9@7N:2WGMTF'XI>K 0KF"7M4[_HR$ R";=5G>
P1C@!F;=B1M!N5YWL)\%R1?2G'50LUF)80*/X G(S>A'X1NE$7YX_32X<I0>0I]J"
P8(LXL/R&'/9%QNFVYOO2V<9>XS14K$LCHBX\-5S;D*^CF\*BVG^K?*<Q9/.XSMP'
P#RS#)^/7N=)%).UOH8"'-(L2J6.\#P7V<D2H>]'U?Y5W3J4B<WC^G91K]WQCRBTI
P\]<)$C!O]0P4+(4LE$0D=4Y5I/+-5?(>I8E.CW:@Q,CTQ92=B3;B]&$2T6'OP&3*
P=P$YR(9CX9]:$MY'FV<P#-,: K-N[&8619\/']I06-YU@JBG1ST#[! L:N4<"V:I
P! [_&4[*PD9S6\_T0.WA\_=F!4#\6E)1]I>T,T'OO4>8S3E]UABFD^3-I,UT!_)[
P^;>0 6:X]S[(_>:A-;\*=%BC[7Z@@NF6=,Z.(E">45#0$8Q">1!TAZB-^O^?1HB8
PT9B)):;2/8[@;\9B+36O91D4"-][8<J4UKFWX4'TCE%ER&H7\^R4]X$II? OP6]+
P:MEP9R$',W'.PPK10H=JN'H<6>=GH!N*C)I?HW7DQ1]VDY(BNPD*MN^T<_' .O]U
P0FEKIO;J<_D%6EZ$U.T67\RB;:L'I8BI@:=ZH&*EW\.AT5#IFY89NU66N)JIG,3[
P1O6M$&G_"$*_T6VKG'U.@L+S.UO3BF9\ZP^@!SG=&;)OB]F(F6D[@@KO@\XT0K;7
P3:*XMA.7;Z?:]8MVX8^K(&R4-.V4+#$1N-T=#ECEE-E P$@%0HXIAXL%]?_&EY.9
P,D"!H QR [.<:!6F:X^-@N!E/N$J*2RM+SY>3738(+(YF"0ZT?#-)<B^8]'=#.")
P==%:..,=$EQM[A]]I_^BVJ8$2G'U<:%@NWT_GVK&/7\/1B2@?)0_^#_>6.[BX7V#
P+HJ/!TLV^P#K^674;8RP0LJ4G\?/4:%Q)[E!66P9P]Y-#N06$V(IVK:P;#JTS^S,
PQ 4R!" N#] -75H@WZK199);@38<*9PN.)DI8>IUU0:86-:=1 (?5QV17UYD.A:1
PX4MKM#B-3*JP3MT\X;Z22V1X32K2G[Z1I;)FXC2<5%;"3DG/BR %<6)QMF@E[=%=
P5L9Z2W&^TJV: (ZO>"_;#W&R;&8H\/B0G2SDL&2N 6R IO*]*^;[VZ?HW%7R)+9_
P1)HK!B_7 0&V?E-*$[7J0@;7E]^RDS@JTFVG R]I '_?@@6D$]R:TIR.!DKP.84 
PE97H>)^X4GBQ@(K6Z535#I)FLGO;_,YP+%A*?H%I %%[><514#2.-32%>A?K>0"!
P?A9JA!'3>0_!H%</4'K<*%]&RC*C)+90R3ML0FQ=X:K9=L3A:7_+?(QD6XH%.*)2
P%N7KL!CN='4102M BFWKC;V U*0")<['>$+8KEGH!5UB"SC($;9FV*G+Y]Y;6.UQ
P=YX87<."$"@Y1(MZE(H<;]-P@?.6^@\$BW,R10['=97.N_@T'L(IGAC1FP_^S;=Y
PQ5B@)'GE.VU]=85@948>C5E00(+P!F=['Z9N^POCQX+$/3&^$XKD3^HTMGG@-\<D
PO/%5Q!,KSP<_]VK@6%QV]&0J9M[;;#KS5:'7&<:LK2VS%ZT*N"]B1VU'J#TN^S;;
PLXM?U:GQ]+S-,+Y ]:!>Y*+5;:23S:CE#23,@W  CIK1I'7)8D]R#W#GT)>@:+T6
PG7?>>8\()5[9FG/0B0N\&QVV3RD&M*O^KK_$4?[I-$4B+7P'%!FD+DO)"2!@C&7(
P$\W$ JPXA!Z$ONGH6-W)--9$%+::=T8"@<26_"!F/'8*M"[DJ 6E^WU$!R"Q0R>I
PE"YVLD4Z9%)\9Z+ZH#K!'GX^*H>@"2:/&P$JU'IRG)D)6^+;W4_J<7(KCAP[CZK1
PG'IWYO[P-& M/]?9H'"SW?=VI>B3XNJ!MWU_IW],CDY?RE9[-/+:P1CAW@IO B=H
PCCAC==^H_[K.[JJ(8;M7*/=#9<"U0J@TL+@4V#'<-'2M)<G.D[76Y'7>GSTJQN_)
P]<GKVZ_G3*J3EP+JYA9MH';FM&!!4^A+C4?9&#V3+[H&BV,Y(4,K'V4JGZ'D')_D
P"6^1MOTOI&-,P>H%+3+UL'Z$:1FX )TAADN)/.0T*5<"QLI(DX0]P)W8:B7?+01%
P>L(GSJK[*)<EW:P],.$ZLR\?GGKW MA\F*5P*RY?#FXJ6T?D11U[2MI8KF?"%I*&
P9_^D$46C;*@C(6#YG[RP/4"=7,\*[8L[.312N$<5]9X4 J\GJ,1#M$7>EO(]ZZ=_
PN,UOP*(/I-(O1)A[ZACB_JU7V/<>4&C=1U30*YWUFFTBAN\Z]2U\J$ZY>DSEIJK7
P)^R#XRAONGIZ&S=P;B&/&L;G(;$5]D"),3AEO4OW'F;]QLW(JLZXCO'SM)JE4L(,
P0334ULYSEF;-[,04)9B^EV-#\8+FI-N@[GK&KEC)=V& LE>Y[L;N>S.-&68 [X'M
P3/8XA #YM^)$TK0;I,/T[UXI=A%AF$L'GL:62 9WPDG[UK:Q4F5L8$82&QUIT9D8
P>SQKD_$I0T^I@^EJ-')6RT1>'XB16B>,_,#VN_J/T'/S5D#<C5DIP]IYZ.+GV)V^
PA(X6[5'YM&P6>I,SW>S>\DH:JA*(>$K-DD_H!%V]*%&:K>%-JEK;7_/R_UITY")K
P.G#6"/P5FQ(0(,F>:>F\@2-=N@ K[S,TQ0N C/584;+R517YP8KM^QK5Z388Q_P,
PX$C>+=F2A[9ST+$;P"2MN%RR/J-Y0B(J:P'HS0KC<"^G#K0BX0[ )D!BRV)1!>=7
P,2T%,J+]F5K':M.C^VU1(O)@6B"S?1]@Z?H6?/:OC(\O7$9[X.MS9JFYDYJO&3#]
PY'Q[:86]XZAT-](:I*74HKZ#T!)CG<;N5H)'S[O7'E&G? N.&=(2C<1W?.7*EB(P
PFDD]"2RG\#X!R5XR"4TVV;K:_!//BF^^EI6%A^!9N-1FXCPY9[ZPTN:?##*K,T$J
P+N\"(>8L"^+UE+!5[,O75;%KZG-BI-R!JT[?L5JNN6.,A>]D[4%D 6B]\?C[K#7*
P*$9D$!)@N.&[4IWV!V4T&C[UMU))D!;W:UO:8O"PPU%LC@V\N&.)+;&JS*!4(SC,
PY"5D,J:(L$07V(ZGD*5VX<HY5E/JA&YVB4<(T.9RH: Z,JGOTIVND+U:V*B?A&1&
PPJ>F<X)\Z [)SD0PL?C!MT[W,>(GF_&>P,:*G_%-!C+OH" '.9XL/.Y'L;IZ"\($
P@Y^S*O7UV$%>!Y\0"5"09Z(5&D,H0>PP6^N+6DKI1>T-(H*)WHL"!^H+7%>R5>L[
PSJR[O0!.I[O*NE 9?_W1IU_!:=&._I<=0&\J8C+']I4'%/35S3SZY,\A)0\#E50.
PSX7W=TI6S:*3S]6R\Z*2F4N$13;?4CRG!#EWB:\FL]B#GGE7/U^J6#0T]#Q#/VJG
P%Q#VYMU(_P4!(4>-'YGG;VK!CDPM9N0$>JVN8J;K19<H6(RY[4FFU.^L]>..++H'
PVSS=%*L[I:A1&]ZV)Z-?K#0-PC7849 P;\GQLD2Q-EW/DY<;=U1! !JH$=$=@_-4
P]@CZ W.NKYY?K>44)0A#(-')<[3%22YFS,D54'9QP7>'8U$Q4RI\)BE?X'?]C&H:
PB6EM0E&2D4<V8@+/JC=?SI$C/_Q:G[T2CXGLMZBAA5\2LS^F+[?QD#^X;-($K\5V
P ]A7EXR&9JDURS+:'7=P?^=[5U#DPO?G-H1%NB@UWKRVY RG(W7;LS-DQB_,$!#%
P5^&DKV<FB*YQHL$')MJ\5'_"5@EN.W6AMJH9T+^"&L>I>]ZC;]W>)DT(BC3"JDH\
P5$Q.H27)(1*)"_YQ;=OG/1 H<2R8IYW_! QC/SJ_\:]WNX 7@IW60X;.OO)$@?>Q
P/IE?B%NT/R6.\*.00/UCT(@+%#,K?,FI91\M;-I/=Z<H7)@T[6+I3_N=$7VV@;2U
PA,B>0OQ](3)I 9NX^LE\>N&%3DQ+V*_2&C7 /W^(1->#/Q<^M9.@&8TDHTR/23-G
P/'7#'SU.*GBCXY5M,&4G<"Y5UNYHS5?93%5V9XV\F$>.!P,V6YD!5I/),SI':3U%
P_N\#SYI#<RO_IT4961U)KPW9YTD9Q_'(L'1 R8;F7"M!(_FD"7ZT30CS!>:<CV4'
PN90^=GAO?J:^KH_\[_?[M!*&EZ^6#O<L'4]58L# ^I4/IR)]_'!^B&QC72D$,>Y"
P(2'*F  =&$:O 5::RDE:WCMQY"Q:THI8?]8K;1H/MI=#VC8TS;F?[NQD@V@'Q#>K
P;:3+)/QU,GTD,!VG0LEG_[FL817AK,AI /)&]S".$H/F!.;< '$F+4*$5YT]KO+[
P-<= HN>2^>[%F3'*XX: 'JS+YUSV[6,WQ4!CO]F>'.G(6O.33H#1HJL%.B(0#V'%
P3]V9!.,UNG_"7D^,D+[E(S]W96KJ E-4E]F^XFMI@J!_F:J(WHX_=]-5A Y8W1Z>
PR8!Q*J,W-K,7MJA_K9CFQZH 9_VH]88.HXZ+S<.B-S\DA&/G,=!-.$?.I^X.S('/
PGOLD?#ZO\-'D^=][1(]TM.\8'!.ON6D4N:95F/F0B86P+;K+X$&%:TCH(:4>CBC 
P8D*%:6!4*+?#;L83S^P#J4*S*55/[2?CTFEW/*/6H4N:7K:17+TAKD]7WZ0?;_R-
PX,$6XN1MWQY"G>!<[;';VP3W0Y]L4UX$A ?IKBKP6K+X$Z[WX )@Q,YT,X#$:!3C
P/^W>J#3YQ"=#C)@[!M>S^T1TVLV^**-RH=UXJ\,,%IO60.&WXP2)49HV7R+V>.:N
P^$MP](R.H/KN7MZ9F"'<K1NOG)W"QLQ]=Q?L^25'JN4&LQT[IZV!FH!4MS?(>P&:
P?_?&5-?*T2BX4P?G5\*S811H/ LGVS/(+Y(F_JA5199NQS[!//D2^M\2:RJQPVQR
PC>PT-P9QS$$0P<)I;5NNECB7Q\L)\I-O@W&P;EU9CA61QY,A(*F&5MO**D5]W]_B
PG?4ZS0'R'> 9J0BBWL'1!N+\MPY&>W?)1_0O#4'\+>@5S"_B5JQOB%X"EM3+1A_I
P86$UX()--U-\E=-,53[8<&FJ22%20G^C-""HQJL@/PEQXA?."1G2QX+;!S'](<%.
P'9P.___$IGP2EKQ9]FL7;M@.*6'<V9.2[U?ON[JD9DRQ;F<X5MDY&N466D,7PT]B
P_K!9"X#P&A @']@8BH0\5\$/0D_(6U)#R,G1N=81[4N:%[>;<X(0_S*&=4Y^8;=5
P JU#9O=1I=WQ>(I%W.5U&6;)\,C"Z)\(.H5CN+N>%2,%=<BO\J.=Q:"/VUUA&$L:
P@PC0Y@/=64^B?E1G8R?Q_9&/&X7YT8G?^"G?N.-PZCE,[V%!9:**#<@#+>P)_L&^
PX0V:,KQR<<B9HN+-CCGN*5^G\$7)J-(D!WGQ\6MZI+>:ZTBY:1LNHG)_54*]:3C4
PIU>Y(*7&(8.GT9V]I'$8O]LL+!ZD%-$10-Y'08B!*3Q7:J/*K?=0TT#<<(\ S6.(
P?W8$TLL[;,4I\\3 $,]F<C.4":Z TI5JVG'PU<41ZSD%H>JJD0R:&U@9<:\&$>S:
PHVA!3P0;@<DSW\B89F1Z=Y!J,Q/9.!H;L)_\32E>[R,398A=WZ(H7Q]Z3 =,AJJM
PB$X?2+?W--;NS8C0!RB?>#(]! /BN,LH[CP,N($RY6=)$3HXS:#I<6L;_4-'*7"7
P# HR$/$M;-O^2S:ICO>!U9MF\G0O6A^1"7-[*%O=:N9(^6PPW8I&,*2L9CXV(F#"
P5G[LU&\0.R,.D39A@>;!+!$2'>37L*_HBRU&^&IK"N27<M])_C0$]D"+1V0Y@42K
P;I[\N;L<J197-D3&LV/EUU&=G-0-36DG4&^I)@)]/!)]JFEN<'W4F2NGR3AI6"VM
P,=[DQ,8PO>NLM[#;Z47N: [#Z)&<?7>2ZSBL*KS"L^>W*\1^7,UE2*$:"NQ^G*>]
PZWVVA4M,_<@S!=RUFD[1CNW.\>6Z3\ XZ&0AFX#?Y"ZF-L"-<&E!XH-,0&@_AY/6
P*QD%-S*9E]"JHBV5(-<4 *9%YP'MU#/Y2]VB3S<S. U28\M+(]-2*ECRI.29)8;_
P)8#+K-@J#AR6V^"3(6URG4EV@"%NW$]$+@-C#(7Z[WY5AG&TD3%-T:.((8$PTE;O
PJ846P#EB[ER2]YGEBJ7%5HE:AOL,1(X5/M7[6XG1^7-_%^M82WWG49UQFU.-]GOY
P_)O'3< _4@]0&U*)KC99$?LUVCQUE/^!TS]+H7U_%T$70:U</\*EYR+8H1$+ 80'
PS;1(^\4572+4Y:(V0?<K^ $WA!,$KV*E=!G\RD@X;Y?%G1<GNNM9&32=%8#\S#"P
P9ET.'/?23NB\4@=XS(LL91HT6(0&IAT):]92PLCT1:=U]^<_1=OO9"BW-C?)6 -/
P/L"LF 4*;U$YIJ/7V6T+/0(\/:K8/I'.,@2?/5GC+N0QH 2\*)4WHXY9--&!+<4<
PMFDD_M;+8=!C6%TW*4'XZY5+\+K[@#,()S<M /]?J9QDXW#&%X1DK:,^;D'%WWWJ
P/JU, 1K5#7<Q!3)%T];/:--#.>?[E;K.YV7,"/T6F65.)FC?2,95WIC#R;#;,+^3
P2)KB:=HH5R<1%T'-K[#"43 DMO!6KR@MZ Q(5OVL^7QR_C'AUX;CH6MC(<U)B90_
PGHTJ\4YDH+\'?H$?3"U/L5#%#&(D>SG(ONL!;?)<D>IX1+?7)ZY;F7>QZM+C3#ZV
PBU:W-$UEO?T?"5%U!6&/$ ^A)1U<4*,H;UWWAYC'B:VX7R2SPY*OU]57N U/(]+O
PN^^[KD0#JN'!8VZOU*+Z[;8LQA0=0-R+EQ :*=]'IF4TCJG297=66,6[ICPG%69R
P(=UT;1)TCH7CS$U.2FPP07Q!K&^48\,I((W$^8'JN_GRW!,R>:K"YUQ_KD._!_6R
P)#.R[9>I;:-M,R(%GQU2U1(F%+,2.$' JO,T;RE8A)#/74 7<"Y_SS:XVF+ITW@:
P>\Z'!-781^@/BFU!\'Y]\35+E1=#TA<LU_@N Z*W$59SR@YRVY7P&* WC89@-K7Q
P$U, Q-[KM^>IX4NZJK*=JERX+FGEJY(P!RWF>3*<G%?WO2\@TD[F34%83ROGGBN:
PI%*V3E%VZ9]O7_V*7L?TX=_@_&RF2L.4!YG7)L;E2?L>5T$=F&4^)A=%R*_90[%Y
P3$\<?=YRK$><B8#HV%?\<JOP5912=K*WQ@T':URC $SK#R21-X#*1R\J4==UO5C#
PAFC=6?0A?DZ&">5A"0CVFEX80VOG\)K?=CK5@,2><K;MV,JJ,I897YOL;AX6&CAV
P51"[-$4.@&D<SU8F'D&GCJ_<';T[VO#(0X27.#+_HPDI9CY'4\DWM"WXQYL!$>BJ
PA)&(WD^TW**8DI+9[-@-D<?8K_>_[97B>X5#,I-(6X=14++L^XETN>[$0N]3 '5L
P:@#:HW4>U*S$$KW4[[PW1EVW,^QD92S7J[/T;8'UI\S\ =D.QPJ2!,, [*2B?<RG
PRX:) _90T\(NDGT29-"I:C,?^\])S0'/]P!<\^V+475QN[H1/47&Z_/9^3P*8#_?
P"NK,UF 5&DM7# ?X^0_^#N^@H_VR?TU=38<)M?B/QN&8&W/N"T*MV""8J5;$.KW(
PPC?OY.-ZS-O\ZX6XLK*"KY1D.#Z%C9!$/4QVEYBO,=/E.;7>ZTJ1[?5\F4+))GU1
P67Z&#<'+BN7K" 2682NZ%O[A#7YPL1Y5HTRXS/;CX*=1=6-G-5]G:A+O*J!=@G!7
P0!68M33I)I-$?A;.F?ZCXXWTAAJ2711;G2A.=E_:2:*P)[/MR\@#U^GG.].:*VX$
P;9^3Y3Q:X[^%I: '&$A@A9I+& %QW;<H']X0@.>9?],;O9$!)]\)8:]-7M.?NUM]
P&V@_512H:UU!GB@WK[K8+1%!(L9'+(WN"$&UN !SKWX(H2Z$G=H42V7DF^NA 2'B
P<_ U8CB"AMB=2ZKSJBA''ZH%?@!"'^(A[^,96CG';<O><=R\UH:S'MY;,NDRQJHS
PQO\?1--D>P\,<LAS T<X?]IF<4");^()V1LX(ZR#6+?[F0\L3W-XK[C_D)?-9,$:
P<9BMBM,C9@MHNM'E-^+'B:-4^'(KO=I5(3*<&GKO)>JLO>_LB>H/T6977U+3;/;_
P6"$R5DBH1N>U"S=4<6+X40!F@W)W1%QGM!T7HK%,P)+X61C^;AVLH"X_/3J2XW] 
P/$O"R'3]JPXRE-!L%FD4%QN=1+YOU2JU.1B=N/*]NT]Q3$<,OV$(OF$;Q#M/!VT6
P^*_HG9DI29UNPGC1S'ZQ9EHW?$M&!&..FMJ;)FDUM["JW%AOUNE40+;QWM'&C:F4
P9NWK6M%%(@%)'9BW(XUK^OW^K,F- 1LM_(I0I_J$.;?:#\@--\USB1*!(T'1R^ U
PH4^?M'!J41^<XU=J&GC&S& 9G4_X ,D^.O!<V[W@A3Y<WP0)S8MR[)],2+\]MF@K
P1C#*[+Z3UQN,R\O'L6C]_HB3VMYSWT>:-D(05^+O,#TNO<Q=;Y9Y59=R$K\!%OW/
PN/@-8*6ZJ&@Q;?8-E_LN1QY!-R] 6QN.#ZHAD.O27NTZBQUZ(V8BQ!RJ^T >$4^X
P8WH5KMLE1DR!9*XW>=N#08=1&S<=DR&LX!3F;>8 BVO8R!<I@A(B=N_>%"%M"O/T
P?;1J)??N<U2#%ST'7G)&(+$?#1'HB2*,PD,&O-XK8!,MJ>WT83V";C&U12#867]8
PM ZH*NN6"E]/,4UW[A!)A3\$-B2BTG4;VAY8HP3R06^3&_DJU__ZIZI!9:[J>*EP
PC<R1 (&HK%?O&\\3,KD!<KU].Y>HBNG6X;4F\5][R@7E=D>:*TV"_)Y!JKR95#A!
PA/UQD=:T"X_P7 T9%H:^C -E,L_H*[44#3ZU=PFS5I@L_LFXYO)H9B-H =5D+AVI
P!R:]F@G!@X"U]7G\EY<;O@5T"V$RK[)EQLS68SA"HDNC?%P3:]L*_,B*5*9J[G&G
P!J8+TXA!Y4!"Y>G%(VLE:N^ DB(V,J_2J8I/*VQY$(D:CF>_3G9(K#P!/HO"+N3X
PO.Z>Z$INDBB@-I?T@UW.U&3,VG7C0\MC7NUE@+#-^%"6MZG\V>F/DY-]%G2P5UBR
PV*<=6;WU69&\_L^_#A[JD@&_7E7(!VTHF=R1B?&N:>F<;]!-'T8N,/+QL&!LJ:@,
PWBW 1.(&LKUHQ!B$TKWX7,>?-X5<364\5)3SI>!"" I(BEG]]GCA %#(35AV?S ?
P3Y,JUITS>,.NVD,ZW'U;(9@ A98($5H12X%4Y=S::VA!@^60[@HP]5CRN1:DZ:)2
P=*SE&C<$^LSY(W 38D3Z()]QU--KL6BK?WO2H<;,-XV"2A\B_L(@<NZ $4@+$'R1
P($O<:OC*:5LR:;-AK.5,R<."W5R.X2(B]VM:DB:C"H!]T$EO7[@G%]".I@)=+@O<
PQG,F5+L K*L>=@+KCZ)Z*/ZI1^DJ26]TGW]%;1U$&"%QL3JN+^>U*\N^Y8"D!5'&
P'2V]-Q/V"?FH6Q:YN_2CUKA*\FY@C-Y X AV]M%5%SX^:3/-O21U-&CJ"5K#0;3-
PR0_GD8H6DO8.8['H@8VTT2=<-IBR"\Q!+5!^::<_817PVB1&+!TT-@;,88O=V0ZI
PA)^HYH%A^T=>V+=]K*#"-;8SO/%4N% IS:/]V_^2UERTV^ H8WL^(6;7.HL0R;'$
P58C;(%#:(6@(DXX:=\>KY9XVA M1(Y?Z \;^D&7,)OY1=\2#QN'2\;;\%$4WPU55
P<23U:X$0.W9Z[MIYH4.O=!E> O6ZR7I'58N%XT\"@D\%8TE,ZSJG_4W)O[5535#M
P/V_6T/WEH&G] 01JO*5X4387@)3;?X!RHKK]=K"+)"$_[=XBUO_+F\J;V^UQUIMN
P*,9RDMJ,A[R(&]N4Z#^*XB>X?,^A:YD1*6*84C\)./'BNR>LM;7 ,$0,"TK]?U%N
PTPVD@_)+5 A-^QNVGN96U*^="&WK[,R>M$F1C??9O_">MH*1H5DS-<%+3F/JH YV
PH@.\GB)]*PT0:LM5*FA25A$S*?_^>_927%0_.7)V*CHX1P $-F ":X M/YN'^NF(
P2*6Y$A:V!"=ZMLX!B#G8*0IX(?Q>VIX:VZ,KC5&&W7_'(X6N\=PYP"%E;@QG;U=!
PJ45>\OE(?=1X3P9P%4RV^JNXTW$WZ5Z%:<([R5XLM[R2NMYR0Q<)1T1JH!GN?V@5
PC*7VL@TA=.?CA89%2") R89QN'2 "!:_\8^=GJ%SS>O7,)GUO<MADFT%&%N4#YH 
PN;M9[%*?;%"U4I(TFX$DXFA4W\Z4NQ7S,G@$E52)U@K.>ADDSI^JZCS#9\.YE<-C
P5B3=IP6O3W7WZ$!.6  PJK7369E?4V)7/-[W,BOMUD(5C;7?M=&QX',/;F>$'5>Z
PAV0#BA-G?1.[WU^3WO(>@&$9\S*,!TJ=F<LV:67)4..CS+<B1-]["YV:"=13;" J
PNY%W*_@^-<767U^5\*+/Y*7NE)A^WW]=6"JV'+62NS"KKRP@HS<'_914O/OVTS,8
P6!#5->K2Q)-U1<$Y;M#Y:=8+T- "V#>2>)")_C@^"<@A+#W5Y*!_NGHP/Z5;>$&_
P!HP<;&MP <O3R+R!V ]B;LQ_1GO]& 2'\X<^]@ER=^76!67./*&*TNJZ?WP:E;L,
P:'0EJ6G@I10ZTATE6U"-BU:O-!<0%8DE<-&5TY=MD2UJ(CRQO_A]E0S9J2^Z)^,N
PA2:.JVGOXS5U5ZERKS&9_2:4?#$M^55IVQ:'<R]:B\4&[L.<+))L7G?V#APLZB]4
PC@:?;P]4E0R[+*S:3=%IO$76?Q&U$0,R1E; :_,_.PKRU>IJ*$.32CLA:*EZC/)A
P-FKUTO"BG @PPF3X6(.2'4DU#,)N405HK>R9U:$<Q8Z@X^9,&-8K^<]_$)*:RWLC
PMB,D'3,O:,+' :G,/BKA[JA&B81(>?XH63E>V5U"07G&QLR(N^0550+FJ(+U"(]7
P%_^='(FA(T?$T>#CU0O?SFZ]9FR#2]QFMA"V$G@]D#:&%;EPDFWXO7DE^-(SP-A!
P8?OTB[OY,^%55VM\;#T>'U!C(L1)2!<>CI""'RG;U6LB85XM=MS</#H/JS;>D';I
PR>.)K16\W57VNHO,T.7CW-,;)U:OI'/29>XS^#@Z=@G2T-,EUR--WKFW8Y9JD+Q8
P]9STDQ6UMQQ4M+7!&$8W"_^*=Y%R6!18VEE.Z$%\!EXHAV XHS8@D_[SLU>>- (N
P50AO:G>UM@%X@(3'1XZ)G"^$7#R\O=#N,G;PK-<VN_Z;035C*PWKE0[VT2F@D'ZV
PI0SZP_U$;[K8ME<E9U9X*&L O<<_"'IY>(-HN9:-D:ZEVE9W9%;%. *WO2!8F8XS
P?A3SB?26I/9]4D[V.M2U#Y;L56BV<5I+$DC4\PY.SV.(54(D2W'-4\+%8"?:+N%M
PA?X!T)Y$GL+57VFL1TWA4CGM=4_O#!<P@U,M?%1-'=UR_A.OZF'_*_]%M6$3W<*D
PF5Q$$%'>L#N=IZ< 0:4FR1WP WC\K-1/10NUY3X\A LYUU /Z1M!;,\S3X3OPT^O
PK9CO*HY2KAB':1Z*R.Z<;48@J"3J_'12POF?G>%7!OHEEP;X?F=[T?E @)BA<>G\
P]*@MP@MGY*&G/2S>6&L8QNIM_Z.L:W/=ZH+.Q-\!?$3CE?6$5UY;])I65.0_YHY/
PIJU/L*,Z^FU+-)$H:RFR3( ''9QQF3BF6#+(0<O"<52#26T\_^7XJ\\Z2%Z0'$J(
P[]& F^F@DRXDB=1+!AX3HW753G":)T.GKRLG'+?!-ZGRFU-R<0*!V/3].5B'K;NU
PNU3)?ARNC:P_=X8/<D3\7J2FL]D(</:J3XHX(2:L?R/AFE^U?XCCI3BSA-J&J<*/
PQ3O/+B4_!>JQ%L4@YNB!.M+^18:I]IQ]IYK?%TH)9 ]XN_P&Q5NAE+92-8-A5 LA
P48[\]EP%$SI'(']$MV>9GRS]UT*%N Q,?#OH@<F;-)Q%H22?QFD^ND"G9!?:>>PA
P]'5*W%4X)WHC2.K'4EG19TWARLXE!7O$1K+7/.-B])8J3.>/BM_T+A/%*2.ZJ-5)
P#9"*"RF*V7_X*.:R0RR[_)F.N+8;R/W+]UX"30O\F](BSUT2#'#SG?U(PRO$;K55
P@3"NRVF?AW<_UA/8XQT9.Y%<)MV7*/CF:T]YSQQY6>MD@Q$8-L$P&W\+$'ZJ4M'B
PU4&1QL<($$M.!,]FLRJ6F41T+85/6XCC_HJR6D8S/&KA6!^6.CR#DH6@+:IE*!(:
P]T 2FVT>+'+-PAQ$W.T<;8X530"R7-55O&'WO%=P],JIDJ$9Y0'?K.V'=3OJ[NO$
P^'2OS_+10KNR<V6$9?E%STLL\7-0H:TTWJ,+KUKF'!37SYG>Q>DLM'F0#8![L^N.
P,T2/V?B9M_H?&GO7=UR<;?1/4U-0,40YR_C9_(0"E)4^LK B0HA\1(?^M69@AQ2B
P#<FZ780\&?(#-:/+QQGCT.Z66KF$-5 XZ52.=@A:T:?JBU[W0;>NCE'.K$RM;PBM
PK.&F+JG2[>Z:[I#W,;9NF1V$W4XYQBQ_9JD(+>Y+Q,&%-=IBLDP53$L:9#J-_\FT
P<6VH=+P*<T191*:<^83K*_'761:%>A[!E:S%[QO)MQPYHZ2AY1;XHW5VW9X=%R02
P[G!U6W=M[[!PPJI%#+#$2H0!=3)!7)DV'TKK!V4SR6WH(J$4:A<RH6V&(E]*@O87
PT^ALA<8C#V\!73'M=3^.PK1Z$7JMIQ@@2^TQ9-?K4@Z-RLR6(P-0Z4E+NWTW=D@?
PP4!>>V ;D5Z5GOJ1P=1P;RBHSV)\G4]:[3)%FQN^&_:%_$EJ"/-02'N@J;7</B*&
PO6/7]:Z"J&0D"0#@JBY8-W[@TQY&*KNT#4*)+$D^0:7%TF?.Y>JF*5L1-7>?:2PL
P7W/K?&>U5TH0Q[)/:%9SEXH2(TS0=4PP@\<*2L1.&LTN]KS#4Y)[(^Z08VP5FZVK
P-@]^W,=Z@<HR=!NN,VL/ X:%39X.D#8^A_EQ</\1RGE^WQ&6<1XCS7B0#=LSSDCE
P=;7%P-FSJP\!(O%\K,MSXSNP0SO3);8QX_2#&B[H%&G+'L%54O_;X(5!Y,5GV0._
PE)L$NH,[9F$?)8\[!L@578IIK5VM+.2<OPM=H\?B]JF(U*.N12\_ZRNTYO")G8JR
P.J E(9]AZ(@!UZ<VO2XWFU.ULN-4;OU?H$ 0(NIGEB[>2&@ZIDMY@]+JH>!E(FU<
P/!JKO6@N Z.(_8<& @I:Q-XSA!*^0.CI),HO1C:W *'X'76P:*4S.H&NQ*W79T0U
P$ =@Q[TCY#@-@Z\K/3VN*P#U.KVTN>;M(H_GT"7!FLPO%J.9B-3%@N>;:!?0DX'6
PK95GR0P(R;<<. .GB\,=_N.-?6-*P,MV.\EGMD/#2-_C/P1%B.&7?3_TGH%_1V9&
P6%HH4I/J6'28P'G!FOL3L6]T^99IREC"/:"8@\-,L/FQKFXD-:;% H^"6\*GV.CJ
PZ!_-/VGP9+[J9#ADBU:TE9<!N?E 'Y<#;ZB^+46NSM/CK&]1?P/;&['WS=!&C?--
PJ;)KD\+T*W$ZWWN%?,_8;93+6\6D2Q&>;558S00S:(U(T6SW@J/-W5E&5/AWH%;>
PW::-#@1_XKS)>5JZ^.M :T(S?O=MFM-[.TU<WE/4,#VCGH8!LCJ3?::9DN[)]"XO
P!:B]CQ4810,NPI\Y"B:0V;?KF:%D(.ZONO49?$S2)<CCC\E7?)\$J=+$!-+51A>-
P02"AEBTFTB5ALLT1)5H31FV*AZ_X"B7C)Q(6J)$'(J]O6A>Y9;H4<GMGHV9P#ZB#
P@T4 T.]W!]"?:]>X?X+B,D[*5@.=68E)BZ&@F=5K@M>IWD[1J.!B5#J<I^L04I6'
P,U,]LQEB%!OYP2(-?L4YVM.DG',L&%0)<ZENY:'PTOS\P5PAV/O52J-$HI[TR6^*
PU6#Q0Z<",)GOJK2&O$ 2V) B/R:IH)9!P8-#:>HS!Y4(U7+,,EORP-2+J(!G8LP@
P&(?X@C:)[CCKOVPYV^4IYPF&3&TW,<#\X/>9 JI$(S,&O%=PU1QXYJ<BO@BZ^D^2
PJ/^3_*5. K[8?GO1SR<B[D8Z(RA4O3JU[ $'R6T&Q=41JMR5_Y&29+OBEE]OH_.I
P PBCK+,.#$>#X^1I-)6GS51$\/;:(29A(C6ZXNUB1]_C(!5V4*N-Z7]9[.?>J1Q:
P#)<D<Y>!IRWYL;WV],AJ@+8'?KMUQ.MN]H4$@P1.5928W.I84HKWPI46X ]KS;4G
P;%&IL<AM!4!3BY /K@-.7182;*]4W:6&%B7'JU0;F?&3U'*P".0=;(>MJBY$ ;M 
PY(O]C0U%-TJ2%US+]1PA %7U3;[OP!EXMH6H^>4ND)S 5-QMGM^._-E:=CZ:8^$\
P;([2:P,<S57Y=#[;B&AF*.RLG\<ZI+8;M?>M OD]W^NB3<@_#A0:8GT]2B%QZR2>
PHVC'\_-_+3^L!KGI@Y#^9I R,I W(XRQM'ZO)SX:QS[;T65+Z)U 9,9 Q-UY'ADD
P7)-0(Q0SMP7*@:$5=6?&+4EMG%XDDI>/\EMM.WUW3MNI1Y[9NL<NMW$XBUG472Z9
P!,1SHLI?/I]"(!7Y\1;UV1^:8-3JAI>->7G2H;M-GQW RC(LBK0;D'3[[9OE&[]6
P"T61IN]N:UBO;*?H5S8I9*T1ZA1NH$=&FA?9>!SF,;W[Q..B"BZ[5%67$QK9?-)Q
PRZX?K@$RU1 8$3CLF5EG@*.7.R.&8"8BO8T&Y.25/2Z774QIIZI(L*A%?V%=]@7O
PT[X:*'1OQZ+7"IW31_I(%8W*D?ZC(3&5H>:XF(T!"[3. E\@9#<-W5RM7PQ*-X/<
PUNX6$M,M?,-T0ON^#&Q==\?\3<EI+KF 8Z^'#L#6:; Z_9_<9;_8O:?6UQZE/?G9
P>DH.)77UM5=W_00&.EGHXT;\///&3PH/C4\T].,!'QU1-NT8QO[IHYG\0([#9WC3
PV;!0'(J37K]XQLX*)0,2OWB&C]_=M[O6OMJ,NP+@+61#:O],(]<I;VFW&O2CE:-6
PG6C'>#^6XDETS/OF&NS%R-#/*P8R:O&E:[\16+*>;ZS=V+$69<^SAKN61HB;2]WM
P?L*$UX1U);M<_KP(!5"2#AI8:\YRPCN19>(WI9F6I<QR_3'GFE(L_NHT^N;5YO$;
PD?0A]!S= MU*?8K$&<ARN[YT%W!,S0[4ATX2[TVD!E.$H-E*ZPD^AIL85$1]2;QR
P^-!*JD@&)OTP&"]J)TE!Y&3_M)G(36T)*^06M="P5ANPS[-$V0,8TD$#\+5MC6?#
P%G+F[1:[>;WN HO9 M?P B\G?#@;N(#?HRGTPD:R,_C"\94E5P-4B=I5?;TY!YB^
P$_#(+P)T4:P?U>#B.6D@?_S]-A*FZ20N$\KYV;2PTTF*1^09.YDG/$!$$X,B]2KF
PL?KL/$4[YAXFA*#$5Z>\/=.-FG$)E"@#1E\:1]!8SM7/:A*7^^D'(#(WP:+-B(N_
P1WMN9'W&HBXQ(%FT ,C)C21P[IQVY78^SJ@=0Q$ E6:F8B_1:],^71@[^+,#_WQ9
PI6IDMK;K%I'BE3.2N2;"9DQRV^DLR3R]92W-EN;T+_$+@50L(25\&R?<=-UQ((H*
PTX\.JNVW&[3E*R0,(16WG@-64V4$,;#()FWM>SLUU _^7L*&:O@0B9=P]9V8<5])
P3B>4GA2\LXW:-V\0/X0V:5H#E20GP)/96ZKHD$YJTLB!]^WBX6 =6LQV+YJ:Z$:H
PC[WAJCP@0@?R,!XD$W2:B@/D8'^WX*[8H.SLE^$S='X7(HE&L-?;L&A_PW4'0G 6
PZ3GVGF&^IUU**4 D:(\"("%[G/&K ?4I_8UV"E8.4\&-_1ETLR(A"T!.U5[9(0UR
PI&8NA2U*DWJJZ!;ZE[:\!?.$I< V;\M(%44$9_J06\O;<I0"WJH'= IL<I/QBD,M
P]K>A$6XP,%1_MO3)MXF7UK(RT@KIGJ=',9Z[*)^[O)2J#[:-JS"[UV>)*;$2Q']8
P8>RA'[CE^C,I$E$YD%]0@4UN6["7O$@X93ZXNM@*!AW]0%D<(#CE.3AX7[27TK2J
P,CTQL2[>25;;XB[XEZ4H65H7K 'M(]D[?=PG(:558H_))#Y;Q02;5N].,9I!^R)(
PO%8\!]K3(<.NR/P!]U99[+EK.C<FJG^;RM(N@P])4)X_U1CZ^,DCZ[[$]G329POZ
P>'CC#3.9OY>M4V\;H?.N="4T-RYJ5:&(]K4 A 'UQ2B5X.V$1=$Q:G^O+>+6.K4#
P,K)Q U)83_'%/7S2*2L? DJC%7T"",LP&ZO3!9&>28-)B.U3B+.^*X*1)*J"S0I*
PV^O4)U)/^;W=^(X:LTV1),IUQHW:%7 )8(B+=(FY$+PLF*!0>P/I-W/(>*YZVANE
P#Z01?930U1KG ]=QC7Y@VRO:U@YV)T9C2!EYJQLCEQ,MF5U1@I H!N,TA.CU9FQ9
P1?KHL P\1)VB]K]2P(;].+7T$BZ*1=$^%_\75QC,&)B#;2,BPX<[^APS@DFLU<C4
PW6V*^4T)W(6D]?Q:!L,M4++M?!+>G779".S G@K!%UR? *; WG6/:^=F/X]5YQC(
PS!"MWMIZ) (R(>#C)\?L-^]FLT.CY<HZWRS$^RL5!?72Y%E;I!6,^B?'$P2@.].5
PM:4*2YD^<>;]?KJYPZ#Z0OAM6CM:Z8&#O/NPX"-MXB@$C-97*8/H/:GB3,0BM*$7
P_\%U89"9)Q_&;OMVM9BNI*(0D-SX!(?^Q?[)K#CP&+9QQ_QE\'VX+Y;.@?"1:66*
P28 T>+W/<8)+5K?3N@CI-ZX<!NK_G"7+,SC$[K"^[*SIKZPZ)6J;FR"B6W3L?>C&
PD 5@M$I8A)W <FK?6JU)>@_']2,S$3ETR+1J,["X1"RX1[E]W3EZW5+^JN2/ &\@
P:60XA)M&5*B5N\Z1U.?9.J?7T/F(\\=-"!3NZ34 -JG7D66C;:>\5J>N549*/\?X
P>/SVK6-_&H;R5"3LU0+_C_>92KM?T_&5(F=@@8#HC5^2!@M.]OYQ:JZ-1'S=1WLE
PR?7,/>[+A3E.T)XA"[U*CN("Y3WM62:+8<39W&;GH/I#7XH:+=4L@RC(@X$ON#Y'
P-FT)P:!VQ-.Z;X<+:"('\-1P":]V6(6B=18YM'QBM#VJ__?DH,OU'^,)E%D5J$@G
P,\7+U':E2$_DX#;U9,\.CUC6)=SK45P)XRKFXXO5UV$S8,ICWVX_3B3P./_I>=A:
PW^Y]/-6Y(7#RS@<]"I"D>.^N G>TW:W4I])/3BY!:?W@+W)QOA<P<9?&#5O8SX#X
PB)Y1'%,26M_92+VD:CK&>D,R:._=Y\J%>0.CHR8&*S186:_/'B#1>U3/&C32B=N[
P__#H+TTVO*5H[,"GDG7"K/);MJ+ ],/, /#2U_QUVFWMUU8\!;!)M5$)&&=Z)(6$
P \_-)8O4AY]-K2X0DYR7ZRW\SIZ6]FK9OXR2I!#B@XQDJ#-N?:8&_N_<]IO/Q.K(
P=4%4UC%8L:J/^2/K;URM<T$)($VI.+OUS:2TSK;0*6WI1\XRJ]Y2IITVMD7D&3P/
PP+WT1UQCYG/AJ]:F+K^$TPT2]T=NAWC[B N*^\[*,72'M"WYWX^I/):7>\3 5\^N
P-HXEXY+'$1)B\/IN[A=QND<'"O#7U^W!<>N,(N5P^(+?@$@#>Z0S $P#1,[$QNG(
PA_P^M=PZ/H \EK$*I]Q5*ZE$G&(JJS!@;2S_MQ\L(!]\3=,I4^BP>PQ>KQX%P9B-
P+S4,8$_#I3K">2;7PCE7_X+G];IE$9'B@<?*)?^IZF2,JK;]]U%^M!$>'ZORB'TD
P.!S8E+%SJJ? KICRG5O;\WR:9?QGHK\\B'FZ3\VLE&T30@\![O4%[&J4T\MH@Y8J
P B7.2B9V#*YW'U"(=DUG(+CZYF!A7TF.B&:Q1@#EZJH9#X">1VT47'O5W2\V%C3W
P=_(B[>+:MY DH6E0._9C4Z&3PR$UK>(Z<[ \A.WF-,]I0@TRU\L^\I&A4SF$=+I3
PY6]F7PY8I^N(A*Q;VQ[71W0(S;K#"$7=CA./H\.ISC'YF1PQF'=T>61K])?W%_6F
P1?^(SNI<;YE40,>_43_,;="R,\?GF'O$;*9.CEHO"A:P:6+Y^1^Q]_1;D&A8R'\N
P*(RCH+P#(\RDW5:H11R;#XE&BSUR&K=]H9SB)OP+8:;M+1X2V04<@, T!%)N6EB;
P\A:H'T0:>O4!QNV-RP\EK.J'V0,)0VQV'F!8/QL+:B%@VG5FIE.DK]6GOHDV1/57
P2F#SX8!C,W;O4%E/4$/%"AUQF+CFFVLU3/_HLW%ZT5 CE%+Q"4_6&K[_N0U'LD1F
P;^(ZA.U)<V#(\U?(LV*?FL5F\7W1P[>U/V+D"BR]$S\-8#W68AJ8YI1G C65>:WB
PK5;$.U>2AZ^5IMY</5S.)S)'=JPV+ G<D-5O^W1*O.0/<](%NS/H^IY*^!&SIGM[
PPOBI@JS!?I[8S:DU_GGG#SYZ^/KM1@'?.!>R(_/%3XMQ'HB-XJ'S^*C(]GYBRHC;
PMUKU(4FHZ''8L!/G07K_R[4;95O?I#:S=O43338'10X*Y[OOCV\LF<\K&A4SJDC$
PLO6S4F=S8TPK<?Y"Y'*NG\519YQ[X,3]'8ILMW9=>*Y6O??889IK3*/C?_*8&XF)
P-S;UR2^MC%DO/W1.9WC)/NT.X=J5N?MXN+<N4.'YGA/4HWJ!NNM^JR;?:M)M P2V
P<A*_$)LJ0\ 5M5$B33EELYV(5<%D!*H2^ZW^CC]?!;X&$G>>TFF/PQ*&;)(->.&0
PL8"+2.9!9T?XG>(@%#P@TSI+??ZS%8<D;:+7>A.VX2LJ$,EF'+)MF-?YM)"M(^0R
P5X&UX*0DV;4L$M0.,G.%@>/"91_GKY2PK>SYN9&+NH0C@N-]<*X?P&:'/C>%H,>G
P>L(5#JI?H/%ZCT',TH/$?#X:[>DW_JARFL^<GJ /+*_=45#65O<&T]5O$;&;?S%.
P\BL+:[-4!B1(_&5:RYR$*R?."K6ZCKG_+Y*;TBX6A&^YBA'!7^0,V4B]7%</]WL>
P>]>*Z=XVR_NGS1%$J)5;Q1BA$HJ:8^=> !^P^GF*7Q&96J:3'WKJ'V7\D%QJIL4I
PBCV$U6TUMA'0*0BOVH.0[;(3A>^,] BWYLGWHJEI1ZW3I@F8&?G3DTK)")@/HY(/
PTA@E]0AB"0JG\ILY%4#]N=F>^GY52&1M8_>XB92D3Q$,%@UQ_:J[L<< ^#M/C[SD
P!3@"P%6[Z!\*O]G1=%P>HAO41L8&<+,+PJNW8"!N.127] _[7DTOLY1*LT6;(IDY
P[Q.S/ L_'OXFA91^9K6T%[FA1B6>QJ.2'&?<CZE>LRO#WO4N)@_(]\,-&^:19--.
PRAD<(K6Y;*48\>B <<CSH,6Y_J2U_XMOL:BQ97==XM*4<!N,._N'7["^JJH/5.[2
PB0MD..RFCJ.SU'&/:?S2$+C[0GZ[#EG:G1TQ7$/=A ?V.4DQN9%V7_/-SDC&F ?A
PK#]])6.1'V8T#=O O2PHXOW0>^Q:@E?G<VQI2 Y7< HC3G.CN$1S2XHGIXU:^I:M
P[)(A8XKU=(354(P$U;R_#\[P[4Q_&^B";WM>+T)\L5'Y\5 D\@8'43;]SE<_^+$V
PGL.Z!O9X%[:P32[ %/!5J8U903S25L@1R\F)HU&.T@^5+/)9%[@)5)0H91,Q$4';
PV!)&?J"#*U;B($"L&@26/STR-@9C-\NXYI+X)^A1X/FJ+<0<B35R+Y-26*E81L60
P:/IOP?@Z>WG.X989I/ J>:#FH 17E!L5(.0'#E_5FOEMAF'C_#HMX^!?88'-VH/]
PQOHLQ.@VI;A=3C2.#PN#2EVE#^NA$G4OR3K*?L9RA<J#?@3GJR[P2 %*'M9S_*?H
P\U[4!X2AV 2&W*1 6@(-TDEANSL%&P&O$!P9645I.<F"J2:+BY#Y[0B(\<*%ZKI9
PK'."&^"$]!8#OA<PS9,!4<1K,NA7;W^ZZ(TETN]85CF;D_\Q2MC!-EU]S<"GFR N
PC4_L827#=#N^(J8_BZW@XA/<_?8E?)OZ:!:RJAL,GLWU?\^_2RS)["00S/Y-/P;3
P_VDP7@.N[A@4##&N$/]%BHVE&3YBU/\/6#B-1\$PPS2,^K7D.\X8M7P3*YS"V4XW
P8<%,/D6UQN] <C2<,N*71HLM'.<:1G&E47_$L8YK=;OSK]HE,B%UV^,G]')G$)W0
P;PW$MGGUK-O-K6*S"VUZP'9%)>>"!JTA!V%=E$VD>*6UIEI&+=J.VAD2LMM%HE(^
PLO'UU"M71;*-(B5 ?Q,22A^*LLZ] ]_XH>=7E%M^1UI=?::@N#F\)*Q^M49M8.)6
P)([DNOA3Q:ZBN-3R&;M+M[:[QU=C''O_:%#T!,M-VK-@+,CN!3'Y5&.6WPZKHJ%2
P&U6 7;O]P*1FUDOA;!E.5OT((3QPFF_JG(*V7M(V=PR):S-C^R9I67ZI#^MB-DML
PT3\^+E^+H!VF;Q23,Z\;T27-R:7E6_XZP17TY19V\P<V%]8CF%7JADE<"WE%6H.#
P\?._)7$W.= U^+&M71[G1JT+Z;U;301.8V$5D(*??$54VQL_P["C(\+OI9$YM0OW
P 0Z]Y?%+[! 8>&>E9,D-*[\I]:([4T:U.P?Y!#H$8: HC>Z/PNM>^XU!I*LLPRS4
PU@AW/2B636]3H*YX9(?-MEH(K\EYX*%!,F$YZK??6*7#M==PQ==5<!BT5(5R3D7&
P/=9N9I<A[X-PT*9>*HNXT=V)<S$HW\P.TR;LJ WBJO-TI1MRX #V)_:?V1T$X ;)
P[DB7I:WP_!Q X_<*KAD.]5=CB$K!4_P-3<</"]U_A_"JT=X[2/MV<_54;#=@/U\!
P_%7$[V>SVW);70*K"T6;BAR,*V^O<V$L+JSHQS)&#BJ24@L\%O6Q+"_'=76*@'@)
P0DHJ:O]WTW!$XM2XRLEEZV._&;ZC#<UC1 F1:R9P2Z4K":7>ISX@R2CF W/7/=S]
PU-:66;X1)#P?3F:LV MKF(D2BVBF5<VCR3ZG?LM-\W*E.L_9IG6")T'*SDNJ8Q[L
PN#%+L7XWI_ESLPX-)P_2E8'Z]C=6(46F.&N'?I GI] /X#KE%S'LS:1VBI>@69RO
P3N<47B$CT+<T*^]#$\R]O\LWZ-7RX4S\?"DPT(@MCZTDL@NV])+)(?"#>%=/S"H8
PM"C.2.$$WN*[CB9'#Y%O,M(T?U(/D9/FCI:AMU@V0>Z!75DQ)%9,S$Y&QMU:W4SJ
P_V)5(5KQ"*:QF!MY0JJK(L_O <!;DO#?6&?MLTFP6W(;;6"WOB59?Z+)J,XV-[R1
P'. BPGSA7SL3GS1 (S]F/S5:UQCTZ;1<MK+"3)YW$D DPN;V:FH1Q!UI[1O1PHUZ
PXRQ=4=.N7@ T2T)1*LXSE&A> CIV7/-4*W6.?W Y"QX+K)6&<*QF5PAN7NK[Z5*4
P*^J:[RS(2C^5#+ $*"+TM)M9&POJRN1HRX%(K5N.X*(5X\SUEX@JODU[-S87T6'Q
P-9M1PMB@-LT5[KLNL-\X:.57 =Z7LZ$+<?2[C8MLC#J^G@QCB):.-@Y5!8R7MDLL
PJB#>_<H.=;P2/W5*P$#(E&0-YZHW J&K'T KG@4]&CI_77T<)%MN*;) +2?*72 Z
PD U1'@X$BL9Z4#-$9J$(4"GA\:C'$:UN3!*>DN=#S-#K'=WU@XJ[X Q?SML'//+N
P$IEX<CN)BW0U<?J&ARG(25NEN_I]BL+B6)+,4A;GW%M!(Y[#Y=<,:P@<E@>^KS3F
P1_=<7 G6IR*$Z4A3ABQV&8<KH6(_=VYUZH$Z(>AUN=*H+^X6@'7%STJNJ0Q^T@OQ
PBZ2G,.N7MRAYAA)W)8(!")!8W4,XI):QW<Z14_"(N@TIJHKQC;V)A$G(18 P<Z18
P7T(:1(RD,+_I]KOY-GB@#U_!#OI\LUCV*O^>%E =;&'CU/399H%HL>O!$C".\S1"
P52:2(''S F- 1:B/,W:IN[PMF2AUY86*72Z3UG-4.ANEJ#A)9ZUM'PO'F.\80JGG
PP(RIOMH$5#I^9:30M:Q$!.(,@'0"$PJ#S8MF6/=H%?3OOV!NL[-?Q1OXPH].TE'2
PZ"^+-.O;&QX?I_H5T)6,9"K/JL6UAU#%=""H-'L-49,TJ?O\PC_QML,CH9VC_H*.
P$[4YSNT+,(YR^[7O Q1+1FF!6,WAN/R+^ DJH7C(?!&OJD[ELY7Q32T3)$DOT=7.
P*8(?1)LJ2[+Y9?]MM+,N?P7+D'G,BX=ML!2<X/.6U6RW8N"8>\: ?$LF9QJ]<QY8
PF5I!CO;84(8=-)7?&86\AC)>NM=J)7ZF=.V&1.2@@(H+I2()O/O.UB^0P. E2*63
PW AG0NJ*N[ X6K 2<SK&#V+?QJCW59VU,FO6 /JC@54Z5A4Z--J1N2P\I5&:OS*K
P.^,[2*B@>97GCX?%D-*^7OKX).9%OR?53"EK2![YN-48Z2C1S5TV.\G]M_?4D2<I
P&^2S&%WN&W$EC(9L5"A*5FXBCC_$ [3>#4^L-.(Q[>J6>C2+V="5S#VHHQ7I1,R9
P5TH?Q3>2QSTW).*%T\2"WF* 8;_[ZWE.639I$9F8=HX@?M:);,>;_.'C1W\G*0RN
P!FEXYYZ4"&G? )6EMZ'A*&F\!;X)/"C5X>_E3QPQROJ (V)5_?N,>W9VM*KN>?E3
PW]=_NO1K.0@JE]@)F11TX.M&#7/OP(1:94\2$<Z>-J(H'-;F8?*3WD+PT[Z^@,BN
P6V$"\;A]>1T%FF<&X-1/\IO7"DD!_VMR>^\5B[%'E+Z)W*@_Y,X^5H\L_O6X\\!B
P'F9ST:D$,=6F:&#M..1+K.PK+2>3-PO;/]Y7[]8-#/.V\$]0'?H6R*?G!O43<"AU
P9?2I\7XA8C2=YPQFY*URH>EK=!_@BP* D0Q[6> *W$Y;%;O6[D0*>$!G(74S_3:^
P^X[1?1'ZC437W!J<+"V--F,-1\;-P9]Q]_(-M7W]WXAQ 82I?-=XEIH%Q4<Z]IZ9
P]48N#4C>DSLW,:JE(7"1OIN8(P!'(TKQ>H=&G*AHY2:U'$]8Y\J\YW4=.VFV9=U"
P\'?9[FB\3" (\)W^&6+<QY"5E!HC#8%87E%9:QO#DSR.96!PR8(RD-9\;IRHJ4'+
PI@.+B8(J'D14_+>PE4'BYY8@6M-Z'I^=B8)$/>UB>('.= M2%Q,OFP--&G&B2X9L
P)C?LI)B5Z;.S>+OK5*?+FTAYRBADZ$G'.EB5 +\.7RCQ:D_:T!3.\4I-V92X63!I
P-J9\WE<T"<//L]KZU^QKN)IH[;*-WEK!RK7M8(:M01@L8&L]&[W?GVA.,#=B@7F,
P93+FZO $,$8C%OK*0'XT][^.V+K7>D8/GBY#@& KW&9JS1"HRZ)4DC"/RWTRAA6]
P[Z^R#02./%0%Z& >G-#[C*OU;:$]7'T@46YM,>YTNS18(\['I28G<<2"X*$3?\&6
P@E?T=C+2=4;NS/ 1JN?QX0,OQ1ZSUBHK_H?,6 \ -\SWX_9-V; &?BUU_2#F*)M=
P+U$^2[HC"5LAC<IXPQGH0N?GR-5T^$\ILWW*3&?\1I>!7"#Z0S59DD/ 7J'</_H1
P;%FS:/BQXP+U_41=T1?"EJ%B?ZK09MO^=><@:":&I0Y;#!M)VL F687%S)\#*\B7
PUH&&2KR$_9[ARBK1O"+?=:&C_30HXE )&>G)VC4\72B7CZ9NQ[J7YD@,0;@"V4>+
PP3?:%-9$F#>W?.0S&N<*;0XV@1>7HSP0>OEVT)4\)W?JJ,$ARX3!AZ]T=N15LDTW
PC'7W573#=4F;/4#G-["]J5J-Z@' SRQ9?\E$X7C/(.Z_<H:CF3PJEA8Z<7 WKWYB
PIQWR)*8T1-?K?,&\[=GD%;(]\O??1K =AE>I^W)-C/,,9!OQ; #J^2?A*E"M5;R%
P)?LI5=R[<L \<=0!L*A8;J<W37U/[[!HSJ$7RXA 0$1??K+UYT(LU5E,*KQLB0B:
PQTCBR>;4F%>IHG_!-=PL4\F60:&#AQ6S&-DE?GJ-E7-7H?3#>O/CS6%7Q0"R6E-.
PP</]&7I"'L;-,:=\F82&GC;!5^G2S,'3FG[;IF7?"Y0!BPXWMI\WK59D9S%6Q+I"
P;%9%1&">=J)PW;/09;F()0Z^3GMYX^%!K%_JW60N-GM)MO?L&+@I1PCD//@-A6@*
PG'T-?5DT^[C%0M<"N3!>0^%&K',7O8T&0&S;-5C#+(CN>T.=4JC+^3BW<E[332!4
P(1SCL99?'@]+S:0S OTE\BPKIWX[ ?%HE=D]S:YM=Q,Z]J6O$%R/8<T/@=FR$9O7
P-7/^)UE8>".R_E1N+NT>SD+,<8PL0E1V,'R(!O!C;-)!Y;5-XW]K8JIT$HLU*6T@
P)V4!?M.@+U#(65O#;4S @-SR=AUB0I%._0EI XEXNL#XVXUF&RU&$]J+H5<-[7&E
PQU?[!AII*EM[D&OJNPV7J6'9ZWS <1MY@8^49V*CLKU8'0//^^+Q::]9B+OE)!.R
PQ=["_A50I&*;P"F@37VBWW2A9X=$P+5JROUGOL^/J5*G(QUIB+NL<"?'P=+2&7Y;
PR9SCT.FIJ]S7$1ODB>6FDMN-9U)3.8P-?Z1_I0?2+0<;=25Y3R8ZB0W"S)9K^(LA
P>19=K:\8P\1\0.WQ+D+^^U'UE.MJ-6"'7 _A[S.B1["J2OX->&?.&-.=Z+[U\"UV
P3J#<!H6X/=GTP_K,T=Z)>4?BQN6F.U"X^8TKB^??ZWQ#8UHHZ<\KPIJ4B0N@4A5O
PZKR[YL7DJB>/JY>GX'IC1S'L]'3.L048DA/ RLR34NK6$:"T[3C /5QQ5;ZF$FK(
P=1-$SK0X>\]+S'/@SW_,8X-G1H8U]>GWKGYXH)1(FM#6]G\T<+BO%]+$8)U?I/7S
PYH1DQ,N"0^!(6.)BQ,*P;_ZO*K]FC)F2W8W>3YL.F*[U:ITBM7;[K>#2,4/JCM;#
P&!#\N;(CEFCV#SE4@B7*V #BC!SPB1W#Q*:I#O1Y6*H-M-,H%VNR 07$Q4O!PN&6
P47-+Q -J:A^BKB(8),] X\O-QS9:$+<=230A^MB>6E9;_0L:FFN>J:K=[X$SXNRA
PX5:$1@7]TA9WN>"V-SWCMX<]CMHK$T/T>C(H2BCUN47E HS<.UP< K- R.DLB:JW
PV>-KX5-S5A.P9XDHM.^B&M.N:10?#Q_[SHL\0"3>3+KS;INJ" <Q='3Q [@I0U3+
P3=RR\-#,[PD4 TOG :4*QMX<??>]9!S")DAX$4P08>YE<@*Q3G09U2!Q!S7$?'*?
PWUM0=*$UOUP4A<<.L9$96*Z]4H;'CHL+KPW3G>A_2;=3KO@ 0"='?=>A9-H"-?%B
P<)C-=/XI\N"N .R/\)Y19Z!X&>C8-[D<SO8H9M#=53H?.$'%]8KS\KPZI M1C%P*
PXC'T'!6Y4P\<'[T6)SGK-#G)7<3N](:/+?WV;B^!BG91LIW=O>^::S^2_K0 Q*!*
P=!BS$+E$1@17[>T"P?#1.Y^E$O(VW_")^'S/]&!+V\(-AY!:<+.*WY![@2XMT7LY
P)Y(,KE5R1#<$%+D]NK'S[1#O9;2HV8&!D/\>:LT1'V1]5(B7#HL&*K.-W>-RNLN4
P&OS=UX>:@$5UU-;/0]B,/&F^G5) @OIKQ,0ZRRS"$E%U@4[OP)#NG_GOGM35P:P*
P05<Y9D-O^!$E5GH#M@5Z2LAW[]'FD!EL;$(UXTK;IC(S2L4981^I28RO0= (,+&<
P3XJ+N7&_+<]N>7)I>$U2Z"0\M6]00O-@&DKHNP?5SY=JE%?6--!-#E"'A07?Q+;=
P+)" 0PVST0W9C:YBKD#SV"HX*O#$3!<60VB;V;4HJFK]ZRNVA2:IG;-Z&%8/]7C&
PG%R#:%<#''1%EIZMC5#G^_6.%4OJ1_HJJ],]5T',P IU^B&HS\8UKF%?U;[TI;6$
P@B/#2&%7?\5M;PW+;"KCN<;K0-12=A/DJ]!XYXJF(>C5QBZ</AA"-A#0R)/ PJC?
P6Q-:MWDT2Y(]YB$%=34Q-1Q=#19,&\]I7V@Y\T0?D[BZ-=GWKS#\]"/5L2BU"\/=
PM72$ORZN;,)$P?&PUJ&7H.'U6T2Z-;G^^6S]J"NO%KHT!S^^E--.H' +S1L+<B08
PQY"2C34%KQ=MKT]\5#9?U3<QN9D) )H1Z:>*TQCX<0=0_*Q[Z$G#88UB5KAM:IZ1
P=33'Y9G_:TTBM,KHYI$NJ>Z=(.LS2!2>L?2 B?^9;>RC@/D6+T5%L>89&SFWI^>A
P@@P1&;+"]M:<MU;%6!^7;S5USRHBZU>">@2EMB/#D*$H:R#6KGQWX4?U?TTK1%#X
P[F=6SA%[;6P_CN.ZT>O]9(1SNH/.;S--1\9,F<R>MP81\LY<=<RSTN"[%A<VD")_
PARFS!/(=-Q$1,EY4$":HW9K9N:>AF74?X19KSK>0!=H.I-=3H_1^)8=VPY/H=?7=
P>6;+X.W-"!'*'W0=6L&%_,E '"RSWIT=WI(@7 $AV;<>&CD8_2!R\JXDRR*<IH_Z
P<<3G5L5637>I1+ \DJ)8@=FP.Q7!K]Q4A$A!&MCV'A;=9C):7S!(+(S$_(R(L[-9
P/7FMCJ?O$0E-&J:"94YJS%L6L#.5B*,:BRP_CK#:"=CG2)![3]?-T$J^Y!:NT(55
P<<I-X/1UI_/(7D!H!7IL =;?YS9I**YLC8^B<$8E8Z>9RO;#[]6%M)1Y8X4@*L5.
PE<?WW8'K_NJGK+04:8G$BG08,JD_>K9\Z%!4 [7VH>@[:"[0,M;9O$]9LY2";L\>
PW1W&Q]L%CN&(7;,(\V.O5A7TU :0F$X(YB]>K7=Q .:/$"X@F&TH:R3X=JH?:9 F
P3.!T0H+%#)5/$N4CX/60LP]^*2_MOG.\3L'#MW7_")[!:T\LPXG4W4RKY#[6LUD2
P=6X?3?,VQOLMC!0G969L%9NL6H1LRP/42NJ?1&+&?G@+)4/5AGFI'T^I%Z4A"U<Z
PUJ\/C2.8L*Y*SKZ9684.URSX\\K!=CPL?/Z/;_0DP4=8(':OT)4MR^)P!^1_KJW!
P"0$33P9S"<K;:9.(@/97!<M+*'X__%@CSNTN*YCZS-KF9AKPK!Q@^DHK[FF*4EX!
PP^>,FG$Z?<)!-JYLEDNE;.+>CLQR4'O7OMYOV-8 1%MVD/0RNH<9+0@BNM(6EN.[
PQBN3.R2U[=K+HFYGG&=/#F^I7G@A;IOJ5@@P,ZNSMNX]CC/>$?];W^EX/ JX,GQ<
PS<5U;^6(')M,7=&+@"M9Y;I/>=KV%!HOUM2&Y:O$D(=B. I_S_BN9C$88YC//"K.
P1B"\W"(MQ[(F?,'A_BKCW"1G<G<]]BW$HO*FPUT;#'#B ?*,F/!;!WI"=%YGF-7N
PPH2(EH6'M)@\RE]1W:);OC9+J:U8*:LXUA#Q3(&3RK%U"0$9!Y*5H)Q[>>;=K] +
P A;FJ?,0)Y,<.Q"XH8Z1-;$KB6+P.@],!@A) X9@MF6_P)Y0F<"+E9X:Z<:S(:\^
P;Y774T_GYO]PUHC]>(L I<%6*9M%6UP@Z1U4%_LP.>(/.$@M4Z\_7BZHF]#3!$YP
P;X3")1Q/KL$H]H22#-P^BI/1AW/U!<IW15!@NC^?";=!14\C[<N*#C.PKL0@ ]9<
P#^).!1>,N(N!G6+_YI;P\>.GW;U?/L<%3&9C^3NUHXD&>#V]\ "7\+<,FLLH-\ZM
PSU+B$=L;[/>1>R(G4/W+#$H!:\R[=]>PH1BB<$3%[N[D)&WYY?#.42,#C08@=S]K
PH-*A<OJ[Q.Y7WZ_Y;?I:PGS;%4$R+V!]KO^JLA3&!5/ J!1W<P1Q,EN-O T;6>%F
PC2#PMC++,8D\*\>_\CG.I+H1U^"V];??LN.%>G$$,5>(-K]S8#60B<OS9?CJKYH=
PV4 .)Y=(S",=1P;Y89U!F$#'TCJO/VH6"C-3^DGF\Z!7OQ?E-VR&5C&6*],]!U+L
PW*BC'VP/9;P?JPM?SHYTN"AO0E^DPW7=C""X0'WCOB#\Y:"'80&-&SX;6C4?Y9)2
P!O,+7$OU1&C;L*9\Y]85P@D!%J&'P.WZ$VGMG*7ECS?8$L.>PW==^8SED"#0J1UV
P:YQ;1P8G(LB@4;-[^LV-9=SK.*BD/(W/'P:J=HK5ZM;Q']ZP!C9S;S*&MOG)'01@
PL?AC^W&\^0$5=#S\?5-"XM WW$[M.UZ+M4E:.'V(P(B5AJH=A:C(-+G!5SIMW[J"
PGH890M6&&>0@H.V0T*<N7IJIG>ILF$BO':LQLN"8(0H'&KLX9+$'(JUH?=<@43<"
P+>:3@L;F>A(W7_41Z"J6CVZ5*2*K&Y+"]L.[\1;XB"!9% 0#[-*H>@F2^Q*3Y'LB
P.Z5 ;*RDJ.K1+['-@.<K3@$PJX9Z4%F:BLH5W4!8ZAD)Z=@HFWJ*?<N[6-(>2:/4
P?IP3?:#I4 ,.CL%-B\\M=9&JF.3K_"3PRO230.?R+6>&,JD]" =*$JL$NT@RU9H8
P*W/?=1&16V'A&7B9OWRB'BOF9\,ZRQA7S\.-%-9U<K!P> 1CXP@I8+]FS^T 0MNN
P1@7/U\ /LQ)&W*<_&$4&$$]-%J4OK%PCZTLZN!>1M+^2+C@/^Z0INW0M^QISNXD;
P.L=X7>T- &+H=2!2X7\C&(*<Y^9,=PZ&92;@9E?%7 Z$YQ6=$4RH32U-&Q=#(P)C
PA_\>@PCT/\_$O5$/9V-<9+1)UEK*6:B/C6=J6Q^I&HF^KF0 $1([C3L>MIB.Q^9V
PZKN:VXU*Q (=K%BNEK14L-[8)^2(*%?D/?H7Q,&_B@##:81??\;7T3Y1K?619<B=
PC70UW"^Q/,3Z>.G(LAQ:+BI3HOJ["!#P?HT?CP"T33E9XL&DP"D?VHYWO5/V#;I9
PRO\VT-L4N<F9_?NR=]/EU^YX^0>'3F13O@^[9$+6([\KOA=RV[:SQ+:V63H!!_V1
PMD/#X$#M=/$-^[]C(9=\DRU:O2Y6$%9$Z84W?2J,631QAA4<\Y1P_*L_6]ZH)9O8
PS6!H!DJ3 L]C+EHDF)^*FU\TO+VG+M<G^SGW?JOTIK6<N"Z6FS/O!$PS72(L+!MP
P4S,PTIY?%"FR)9N7761&-B=@2D3[QFMRA# Z \6GEZL=GTP$*N%9J@ZZK[@E5WZ)
P.#_U>OJ$QX7'F @8K!ZZ/;Q\%VE;8]-6=E,X(55FVH\.ZI]TVW'#-3K>Y+PV$BI=
PWZCK=A#E+DF?S:=?L7<L@,J%=9?VC"&]F+S+U]52<@9 -WPPAX'EA"F*MXB9"\[K
P%/Z36MD71UM1&"_8^$8@4.MQV"O%ZX)>3W$]./%?XT__:C>?*=11^RU3Q3WX BJC
P/(:I2)QYEDEA3FMZ/_.G8R!B_)T'<>XD*O5=PKP9_3+L>AY!&0;*8T;W,-9J?'F1
PNGPGJ?%4]S?LC$!^<MN7G.;66.)/^W_/I.S%4AI@[6UOSUV!AT&\<0:K"_S^M5;N
P25B2\Y;1"R^@YD5\EM!Q[BRA''%MLD2SX$LSLM2<NLV=,FOOQ7U<==F.GHBI[O:8
P:,]%&_:VNR78(Y9'43]?BSLRTJ_K!#+ZV1K(_KVB2VD=*KM$;JCJ8?ZU;L5;7D7S
P>"0)76/QKXB%1Q-VFW&1+[MX69V&^;1:.Z7I#UP*V&/"ZR;EEC.![@2&2L@>E@-)
P=K&K*=_4B8G@L<%"_GXJX_>IR#M\75S0[I"*TJ'%7T#FTP-RK9N[0VFB('4D(S>;
PV\I8!1?;@\Q0_DBT=J6B4'*S7 H0.C+L:V^9$: C:0AG)9_/+P9* OL.1X"OW='3
P+8#.L14T]^($JNQ@[$G!')>X)0FS/%XLP9(2F]6^-F>C'6S=E*_AD.3I!\*II*&[
POO:45%2A_13B@-;[EH!ZKY(,:$IM4")&7NZ[(51'BM&=!<Y 723=2V>=[V)7;WUJ
PX$ *N93C)90T*A6;(C)0NX9_F=#TU7RT>E\BMX<X9_@/!3LQRT[1UVWL+.0#O<6I
P@X^P[+0JAB"/9$*IXH+*\P,%<OR;!/3WO+ ;J5\]RU9[VY'LJWS#+3WFE6*]J+@5
PRL%I4]FN@VQ!C TUPHN[/#V3H+QQ+K;;!XM*>MZUQ0R+;JD<"OS,Q )'4>_;UM_<
P8VB:@%KH"$=>%J16JB)4D',6T):SY3T2P?$)!C_NE-6*C%CB"&%XC=0F@O=+D1_8
PA^3TNJ7IXCV*,(4P\;GA(FE 8("]"C&70I>W54&5&YOAH*2MNYPR(8#]^*@/9OQY
P+%%IW:?LL-N'[X8,,NC@!W.+1ZY]#;K 'LDC:,JH34BJ-VEZNZ"A&E=*!Y'K&@>]
PUJNXE-Z9+F69ME #NMD:!/4@WFYNI)QG,'M:X(DUCQ(]+!J-S_3[%LY5(?/ZJ>E-
P<"MP@N=16EW..^T!(/N*9J$/!9\7VQ2=IMH4?[%>%+?E?]2OG)" ;J8S594[TF"[
PI%U)JYSE2#<?$#W.JBK!SK>E P"R+T7:VWW0%9-ULDJ\3F+G^<4<]9T'DHC[9J,L
P*9NP3KM+XY:.73*8=?CCA<SC LL?(;/STNO.@JL\-2G@:A6XG@,-M*4$# D/_2.,
P>4DW1U1FB6T[@?J=P[A)R6 +-Y+D_0F?\Q,<149-\2>SX\JH1:?M&#.71*"HCA4Y
PE3>XVRDG2:\7] <NCEJ$I1V]@,EEMHCK_[\V]6 ?_A2KYNIX/J_[_5B052Y*^YFN
P8+G6.@Q8JC@!X_>@ 4-33HKCB[U:TOI]_"=I4WS%T'E_DBQ1"\K<Q]=.%G>]:H#V
P=1J*NC;(HE?\S0ZT%0^-UUHK5'A"846K(R#9MX.0&A>_*7Q<9:%$5D:)K@"<T%L0
PLE$Y(^B**.[Z_$.[4K/ S))-?)I4<=LEM G4[63=41(\>]0J]^5%+.5$F=$/^GS9
PL/]*+[D=.IS4Y&![4L*VOWQ&>S]F&,88C FMK;IBMQQFM L43(^OL^@!4?2GX>^F
P>V:PK<3,R_S/Q8;(CT0QC\CMGR'VG?EG\ 96HPSP$RV?JQY=$_\I'LD/HVB1W]$U
P?'1L@CU>*N[1\YH,'VABH_$^'%K2*8$3U@]?NRU$%=8'1LR4_SKW>D%(;&UI$C=+
PG.8XLPQ&V/?2+XV?3B$HZ><T,CB8U3;OH_ U]*>:XDL+%(G%39I1P0B,]63\ >OF
PEYAA_9DI+6DP"*[(V2?076+]KQ_%G-,^ B?^4M_DTVHN%'XO8)=A,I#]N-*34."F
PRP*5NJ9T@E;-\+Y0MRX,"#CVT<1(?+VG2N$,$Y%UW*,)4!R8:\X?E3@.$5E1P4:,
P>IX<"_96>/8.E87+=IW.+"TT,Z0_(9Q4%;&GBO#5!MAW3"T]?;[1=)\%)AUV"]W,
PLSB6JHKJFA@1S5S8M4=^U[PCBKS<DL%L)": 8\CU,E:">0_)Z4E7[%VD,X[2L:<P
PPX%E=2:4^HC;=43@#0H$UAH.NA>G(8,$_$$>C[RA@M]HK-JX%]B+OK<@9F 3I=Z\
P)J^SD'6B_^MX*%J0+YB,X "1$)=('#9?R8<T&LOP'TST&EJY -)&J!H M[J5)5/=
P$*0)AH=#AQRFD?GO=PE^1>)6:_R\0>J)WWI<J>7;_!8"['.%MVM'@\KYDV'V6(>E
P(. '$"SJK&T2<9M%CV1S #^TX84$:F-Q*SJ'GUV&8\Y<$'EU(%F0$A^M@E,;6_@5
P(_-2QMEV9X?9,[ 1KKF%?_;3.=E8&3@%BWC:-& S9SNA(6FR-X,V0*53F_2"FKB(
P4^L"/Q16=_J_/+6LA=<Y';2U^,F2#L5$-*#B&"7)D4S@/AT!<6$#'6&K+*(:5?^A
P3L,!S*$>4JJ'R$TD]X]=(+,Y^@:?]HQJD+X$>J:L-6G"QQV%J?Q<ME(']BA'03PW
PVW*)0\E.4*E2U?<92"7JD:X1A001('TO>3)-^6YP0M%+S31\*K4I;<[M6(QC>@:5
P7W-B!B\5$;X>N]+"";U<GJCL+V!3LC&8+\B['W;:D7H,XH8,>#10$5N^P,Y"(N+>
P,CUNYSL\47CX*?^'/H7J= HPC!PW VB$.!)@F)W8A\=A5'<;_BEN6*?%GRP0[[QL
PC_CK%[SCD1T1I4^2TGBZL9K%SRW*2NW%K7,N1_O.1J\SC,08&.ZNU0@*2W!XFUMC
P3T;6,-\V\_K5)U+:HX>I_D5_=AD:@M"7C7XB"TS!8F0I.N0UUZQ#3>_GAP[K9&E!
P VJ":Y2 42QSQLIL/<OC9T$GQ78.ZNQ<):"3X13"NR0<FO@M(_:!2X:N.79_'F 4
PN05R@)*ISOY_*S@US[GJ"^,Z0OM-1Y?,R[X?^V[_>O_%S9>A14C+C'N><_Y;/\%\
PO4"H0'M2;=P+_WA/_D][^?U-'5%U^W3I5!+ -MSIK<H-3@V*N*P9/=T%?@/>-,S3
PP"L=36%?BYE?_E02 K/ BS\[MS$9L\TTX&+(DNG6N#WK573P8_0==5'W&D /'-*T
P0D$D"E;55WT:3(-\$YW&-08>\.[;N*245].EL+^U@)ASV$.)=1;G9@&N;$*6,?6-
PO/ VW3QV:=W$"TA9R&FGE6"5XLA/T68W$EX9'&:3#]%A0>.4P#,[4+^9JZBV0B#/
P?X^RG._5:BU;O@-Z,,:M?"K\7A^>WQ+7J89KB5A+XM3]>D\3]QO-1"':.?O>E.&D
PNB0#S<V\(1C_[712> DK0\S:NE)S_1@UZ#=6!V!F]%U4Y%6XB2;"YR;+@ GYI ^2
P2N(GE8./#*'_0\M"53>'R_ ]?>8X(3V[66"EZ<QYAH40>8UD.[L\G?1SF*K>!)BZ
PFI 24"SN/>P/G1J%%Q28?N8?_Y&:[3BZL [N8Q80#IWL6X^D22BSW!YE4H@U(GM-
P_S7IY@P@)U;-U]52TJF\R?CT+QSMPZHP]F=J)R08$\!VD+46=T#)(<@N(9#U6@$'
P;>UF]/NX8X(6E>JS[['57V<>55Q39X>0 \6+OI=*C61OR^M:SA%<W%?$)&I*:KV8
P2B.$LG!*(VE;12AN[(""A'BZ9#E5;@(E&L^60&4UU5S]R(<&AG$C9-!<46GKK.!2
P;/CC#BQ1J%J '*? 3=+K!S&D*E3!-<>7-+TL/!,WJF\8V[8ZW5KE&_+810([D/#5
P+%T/U'@3?T94/^!'!;D(J^JS8'RX($Q-ZNMUZA% :)+)F0"8>F#\B;V73OG5,87!
P20W)+X,C,^T0D)!:!,'9'P\#P.VL25V"HY7]>LGEQ2.&C$ VPD-4S=+\05W&OH2 
P7?P<.@BQ9BNY1HQ&)_?$2;#8_ZPFM:8)IF+!U+N^)">+^+<.ARMI7MFW--P^3^=[
P1[:*5= @$Y;EU!<K7TN(-7 6AQ<ZI>^MCV20V&+)O SXX$9SWO'Z,+EL8D/@3,-]
PC41BJU!JL[%WUU+<#5.RX(X<'WEV2T]/4Q[S!$Q13$VR5!2G^[''5.E[]U^PW,8,
PEV[ ILT'B2WEU:.UM#S(;SM^OEJTVH,V_$&@>M3CLWJY$8Z&9H7J'QD<2$J@H5SA
P)@OP*B+7-0J?&J-3@S>8J8MY:F[;#,ZR#_"UO_4J9:/9)5(!P3)H,>/I: "4TQ>D
P$1H<7\H,>&OMA_(G78&O^QY,(YS@ZDI)+PZ&39-N_B%WJB1=3B2F=Z.F*^;."=31
P!23\%_K'5/P-D8 <K:=?7J9J.WFSLG[PT;@E:G\6"=(M^B#D_,\ULBLE4UBWT^;!
P=IR$!+DY9U:8*X%V?Q!M12Z?S"E+4Q>P((-^!VIL@8<7R*^[S4G:>J6Y?(^@",W*
PU'F^>4,Z.A?N5IHGITF,5ZYSWJ _!MG.Z_1RGCISB-AX.%4?\2Q\EEHM2GIT3%.P
PY&:%T3@3;LF_&U?8D$\J,6&OT^GUJ.S5!WBBR*ATD6:%J;-8+I"X_%7BU#?ZX<M(
P,D=*<?6?$IQ*$P*D5.G2V7LGU;7U4XUH7")Y4LD>7$)).@?7AM\!,?X!%U>YXP;"
P?T9-+.#+-Z.[_(H'W45$?D@]M-IL)9=;ISQ9Z@!%4\<VY1C]^X.!4,(;RBUCZL:2
P6^9/_$=+;0M!PU%0F<@;[$+UBG3\ 3 #2#"UXV$LO8EE4*7<FU<Q'7>LPC0Y)(]X
P7P!AG2^W-DEG*TA(<4+@)LR$0WCI,0?'5FN??9R#6M'G43;"&"&;)_97X/)#)3[O
PM1L9PV3O$AB\O.9 Y)S9$[R<Y>G[@O&<9KFTA0:)X\I;T7*;JX$L'PQ[]-0MS3XE
P!-')J;[0P[[,P,I*R+U]'8DO3Z4>BTP-/ED<=Y9U63E5)#=\<XNR3[6,TP' 6NR7
P7GXD3B0N2K$9$I=2R'44<-,6UW@;,8^7Q'W3<%]IKB.?&)3CPQ0-BH&=7K,-26/%
P$K<AB!VDI L$1P@N'DXS<*9V @4+6:)>--8 IRN#V1$FC4E!),?-@W;=$ZX_?^NJ
P5 L_4QT3KUS;*7"I!^)'2M,(3?\?<["A55DP9EG@0/-+E5K0L_3]JNDAHUIOZW;1
P@.45I2,(0+UA7_FU5>"!EE8S5C+\G!F,C;;BK[:.44C?C]J+OE_!-C_C'<@#MS4 
PCML-Q^*2#'?T.'R(C_# BP[X*J-)<\S-/DK%8-5Y$G,'$OXK JAKTS;U.^I5N_RL
PPV[]XGBM,G9@-9.H1=F&[YQF7OV#ZT:X\'2@7.!-86 %>*JAUJ=Z03J%(0XE*%RM
P$R2_^DK:)B@V&?8H BAB4\@$1XK^.1Z=K_3]8DH26W>R1A2H_F5TO8,=RDP="7GQ
PL_PF,J)WH %*P\?" @;"9-:#<KW@*R ^-ZY)0^SH(T 'S6/CMQ2A^UDKN\NK&V9-
PZ)"]>A"(X.\#2;YUMGZPWN%@TC;CT*K-HV))C>M'BJ;M,(0#(Y:ZP^]HS\#FQG'%
PYR44_-35%M?MCFVD'9/9JQALUS,31^* 33N_V46WK7OC[ 7%Z=HL:PMR\>V^QKE\
PM$T2O8B+LN2$ZNCY8;55=5S\<X&R?UY"+.UXV)3$^ADI?]N<+MW H_!$V\)FPE7D
P!MX/->>TO,;#\R/<WULXSF%>!L$$%:DI%,1%)A*TT_QB@?4_S\D16!8B6I\(2QHL
P@[ )47\53%:++,R[(F<)*>52D7G9Q^Z0CUI-0C,@)LFW*K%16I9[GR1LBD' !!%U
PNY<Y,#@)6PH"WG=?:;ZP <',]:_!L4 G9-FAX'T<[YSS(UK]&'Y5>D^LK%[,AP3%
P!@'$K1XD^B[UGSA+K 56>S$1D"4>B@^2TX#?>F%SJ0HNJ*3N+';%OW3T_Y"J^0,G
PX-6"S%[4GN0AW4:0H1,@NR[N&?5_33J-:+,>,2GZ"/89C6A2"F38[I+LMKT $C5^
P+!=.F/V*J*,!UFJU96T3GBL1J=N@FW[QE[*R#%J,#-\88]MO(<1B5Z[R'D,@AK@B
P;]9>_K6\04+B-9J:"PKN"H]>,<0;)'CV@(_:.L6^9/+DGP,QT0C=\7=8Y=JYR=K8
PXKE *=C#H-3???I>GV)39 THH%BCN3G-_,F20WGQPT9"&<U- 7.*%A"(F_"G"<6[
P!@I2.91' VXM-%0W8-A$8$CP@GCYA0,+3)X];)J"):CH&?GG-.(F'F VJ)DQ C&Q
PK"*Z)IRV:1-5OH_@!$_-;[*3GVYNBJS^AJ1WHMZP)?Q368\QG<(U^XE;/]X3@,@0
P#*.<0Q+-4YY58\ZBJ"+6";0:G5Z4"%3G.EAEXO=%$HXA&/'P^/E%9)9"6\4*4'ZW
P[,N)K8938L*@ UMT[T;^X!NE2SU"S=M.1C&?\),<-6AKN1*7P;U%VY;H56C"MQ&R
PO.S,\E-$D !=P-B/UVI%?W"!=,M!U>M:U@.0YL4CN[O:I# #^PA>1[% 2,EE0&[)
P@*8@"L1QAR]34S".%@X3$G+:(C.V6!02U8'>QYD\Q%7:B9V! */CVW'#(SU3CVH!
P]>K,&Z&W$LB%:]BEQ.G(A-(]\9X/3+E6?XQW<:\>C<2IEI1U#W!*R#S.12NZTLO"
P'?"O>K,V3]XO1P/CFBV!9,65+#J'FPO9HHN*GWI(\^S68XSRS=OR6S+Q)3U"+\-<
P*['8AB)\!6G9^,#Z+1.[&.N<*PR2_)>"#!@N7PF4:20U/L5-J]50/HM*<>![27BP
P>9*%U8>'&V-F&EA+#W+5%CV=]>^CQ4R@E_JI[K/,2%RVQ_7"KBI.>(QS&244E6IN
PS_:_3"KNLW LI1C>,<]@5]E<%?$\S%(&^IH69DN),)Z)_6Z1'WYZ;[5NIBF$5$.S
P>+'-*O@H1PKC49ZH9:R+V(3^8&JC>9W9,]T:0E-CYA7U2>1PH@]86WDX]/L0:L,9
P!J3^UWXJ3MR!6O4MJ@9$;15'K=AJ5*V-RHJ@>B):K+&3GW[T9I:^_5*(I8S=6/+=
PBJ=IX-K!0 7K;XB)=7Z1$*VL;1ZXX">QYM$3UP,RWM) V-7M8==%DZ]?#AP:JGF5
P,96+&/8/ D+_=Z/TP,\\TSDIKI>TW]*]E>EX5H\\:8&*DM]A-P??N;W_MR&V$(>#
P_CB@Z179K4B'8(:0G$"OQ2KJ Q,_XQUAORA*1!O$"!?7X-<CY$^]:>=?-_%9 5U$
P$$Q RB.*HZ;,HDB!$.Q%=GZDB%(_LEQ",TMK@Y!J-W3&8.X!UA0A63*(10N+ B$Q
P6KU,.7_N6^+V7<D!ZQ B'ZF5Q)QL_[FQMJMO_!Y"*.PC\1.E^4>;N,!G9REKH*(5
P>O>Y$A'P!)E%7)C&35BUO?:DCG&52L0L%<'1)_6AV[: 3+Q?5VVJK_)+E*9TC-<'
PB'W!RG$,T3W7+8HX&V9*JG_7E\66W#X0ANL X;>?G!DDD;5D_T>&12=4TRC6PW5\
PO6*_\P*T_X"N3L];2*P !Q3M1/PEA:$FQ*6$)_:LT/7\CL.4-Z=F<M*#$-A<RZ0_
PY)>N U0<2:"L\(65_@9 %D]"T F'[MO<+P<^4PK3&WX]AWZ\+CR2"!8>7SC2BF"7
PA+ 2%P.HUXTZBDXW;KC"\5+W,;'-Z44[I%^) LH;J U50BUB+4"U-1J&"UJ..TW>
PA^IR!DF_,+7J*\%)$N&+\312><U)(/CO= 95@NBGH[14=[*"(""B)IE+(QT$D]2/
PV= V2W7V%5=AHV-K9U=TUK)@I#/'%^JK5N;/>55A()?34?-'CIV0#%A?42  662-
P',!11C=;GR)P.N#N5$7RX:JD4V9E$A5#$&^'0E52M3 4L\%]>EKX+*;)(H94!3SM
P0[W@;KYHCQ^!QFKQD?D"C:)J>PDSP[D_;D^J.*)A<P\MY/ ]FY@<]6G:,)']R\G9
PU:]V&;P5W%(F7=A=O= &S]0VVT_:9WF"IE50A]'J1C133_WM#WD(VKQ:4!/98/&0
PCQ$JE%SI7@CJRN$%X&/BDLT-YPG6W(=VV&5?TSNKW#6+O/9^H?WYZXZ13,!['D&A
P]-*$H'@^;;K[?79DS93C-*Q36=3V]C-,/Z=/.(F1H89YK; _<4_%8J!TXGI9$12T
P0<(T$/+VWC7!ZH#]Q>UV(\ES'U+ #7HH!*Z9*4_+>_M5RC043!GXFT+8@A$)]: K
PG8G$)[O+?<3:^$J?YQ"PAGJ)T3F :B@F'P;@^+-Y:(B^I\-TW[EC,JC#?/]'J- >
P7A>9X,ZDZ>&-S?3Y?3:@8*3^;^5S<DKLCEUS73CJ)\9XTYTY=0G6@T5H\V)8H;PA
P E&,W0;9U-65(G/=K^]!Z!)UNN4654#JW"[(C!GS;KNN4N_6FXEQK;0L]3ZCDQV5
P[V.DMS/Q^[;D&\ @M$T8$ZT[\JYC3$;;K?'FR32[P%:ZO;/E]>>2@=#UQY^G-%[!
P)OP:9A@-O+H*)<M"Z"A^JM:_]/)EZ/0R4$QQ+=3W+[,/S1KPL[P7. H">F9$<]]0
PF+*<WY![*VYK5S89"VXQA,'UV/I%1/TFP+&='Q\H5'TX3S )8_F#.;!H<O1=P^S$
P68'8N>N*Q!M3-?GY,3N'IP7S!E&MPED!NSYKGV$KPFBUF(YJLK=?M(J9$CSN',.X
P!,>W1\K->NWWJPUO78,2(OV+N5@%SO#=;3)S\1<6VJW\MXF\0V"3"K"N[MM94Z-X
P_ QIJ?\V^ 5Q'VHE'KO+V"._X_,J%G /7U=DJU$?&BT3<R7D#^\ 0T'V9-F=:"W 
P/T@G'#,YX8R!L-."+WU/GK7-+#IU>[KOS):.D!M1.G%6\U@O*1@JYVJ1IEXK0GLY
PD #3.6<B2#9&-.(6_PFICH<POSP$Z*0!(41IUZ>Y#%.'7/(NIN),0USF9!?+P/7;
P[,P(6>V"6O^\>QDMXBV@>SXN&W/0_E>86A[A $B&*V0"%+R$P.H=A\3WI+G4Y<J^
PG++M/'=,$FK2YY=4JI7R9YI8HH?=D&/&3VW#_AQ&KD\5%!XB2ZISXLZJ"]+YZD"3
PKJJ:,B-CH[9X.92EI.36:VB<88&U],SWV(=&3$Y,V=;5B*Y?*<NE1ZO@[L"'YO<,
P2ZZ18=LMI3B=F6#!_%LY24L9N!N,#C!!OC<3;I*X\CVF3*10"6_4&S-$2?-(4!^#
P:+QKQW1=IZ99O.88^N \;HG>Y#ME6T-?;C[R![GG)&<')V.,L[Z=A1^#>UJOVN%C
P:"YF/(N0$%Z%!$DZCSJ(W4S:,8(@UC"#K++*N;E^9$'^=S%R'/,5^9&E!'@[.X(!
P6;QC?!SK=<'!WYN*Z)*T(@GNSBH&]4? FM*]L-!!_U"F:)'2^7H!#J!3F3\=<;&&
P":[3Q>_0Y'KR9EZHY928;&P)JBB1FOV#<@IL8LG+LO\O!)3\G5[;I>+*RJN1?:QO
P43:"*H>'%PR.A%G_UB#KS//] Y;YMRL;WP4&2$&,4YG[/*#\M->[J5J%;V2KK?<4
P"4.W4Q?.@*UG$12 OPX^*\ZOS*R]#M+7]E^2,_NH=&*IS>R?,Y<1W[^&3CCXSHNZ
PXB08;83,W4NP!]DB0VM@7^$-9RKL2!C;&?5"3P#Q[PW-GE^@Y#D/'BL :?2PTR\8
PY;W3;VGT<@W;/?S@JL.)Z4+9@=S6ACHRO!; =-*S<C)I7@$E:<!_X@?\<U30FJ8\
P)H@Q#K_1E0ZS]@I8?$5?<UE70WE)DAQ&DK;:(("4X4D"P752BBT6R8"2E'!?\V!N
PBL=I*B9.P0=3CY.N<2\\ZOI[J1*VOOC0@!^Q;;8%JL&]]"U%6',J4*M(@Y&YLJA\
P*,QXP3%JRRL82_J\EG"6_-W.>+HKH+8 E\X_M_2>L5O:G>6_VJU4>#H9?[&X-H/ 
PY_]HQ!^\$ES?WAT$5G"3FO_O::%+_X=H]_Q&<2M)L*D6XBR^=E=97^_AD1R2[.[!
PO7,1P'?IO$DY'#,8H$H+[B\9G)I%+(D'V11JI[38Q9L*%Q0HO_#Z@8F0X43'AJ81
PFD(W.L99[)>;59!<]BZ=F(&ZWJ:>=57%K_@J8(?N@IG(N.??0H7^WJ,\0,(\3(,B
P.TRER9L'Y8#]'$'WMXH(=#^2FE\; 14 P!"NV+=6[,O0WWC&1SMZ)O<A17OA' Q3
P75Z;0X0@^S$W/3!4;NX#7W-W1;\58$/#_D%$DWKQ0>-(W+B $O6"IZC^,OA7NTI0
P11T8=DJ<L?QIM[!JK&)@['?(UH+=*\2X25 3?:U 6'5U^SL,8%9'7$:N5 %J)^V>
P*4?M'EA8'"[/M"XJEULD2GA&G/\=Z#^ YI'(A1^Y23>/*_ZO8",O^&TT<4JV-HZW
PRB\LB_I!@$Q',NQ&2/HD'JUOGS^W0J_U,G=4^#YD=D9\<KR'?$-%YL(X#2ZO^:_O
P4<I.*VD@()!9_(3W3RI7W5>K"+92X:S!_XFK_$D)@$U+]E7B4?O+%S"ZN,LN(?<J
P5!>WC%DV@SF=L9>3Q'\"%3BZP**AO+>GPK;_7B:X1A'DN''C;'ML)B,9-*N<0!NY
PIA95&H/">TDS4%A.M'N"YS IWFM!H:Z2BG,%;WF_FR@+@B$9%'P:>$DS1<%_!PW2
PX%:X#P6_R@PC_=HE07G@R[VY\7N"P@.P]$=8R ?_=/'G#\@:5PY* 5:B]/36]L'\
P*K$+9_2BLCJ=UDNJO49UX@C>%5AE\$D94D0=Y("""(459-;WM14_W5<UE/S,UU%/
P!/C99":U88!Q.KD9BMH7>%#PG >^#&(KGH#)F/>. W?=[0-1(]Q,[=7W))ZB-8^/
P\3K"]SS$!Z#38B3/?ZJ"NRMG]QELO0K_Y@[MP <>,MO%DC.:PRU0>7+6_U(S[8ML
P]82H#D]]=8TTX]O@[M):V!?CG?N*I[#CC1?HV<FN'XEN_"*32OQ!G,!^DH@9C2F)
PD87.N]>O?S<$SL7>SRZ'%;;Q6L&7L\!E2IXA6;34ZF:FX53UL7\0*#7)HU8H!N/$
PV\KEIZ7_S*VY2-@-LYS7?MW"2L/\9JN)@[TL4>BM/UI<H]2P#)19 P.'.ZW?*P)]
P^&U6[R8!:_ 5JSK<E /V?GZFPRE-S$N9$ZD$V;M6*RSOCS+2)1,*AY%WAD72-ENM
PPC+0$\^<')^W).2D8I .ZPV[L=Z[7L+BG@8Y% SAVVVZ%>HRATL W)Q@K*6"HL>.
P,O1,SA-C]MNL6#A3PW,GK@KRL$#?PHLY++2.=/5K!*\Y$WFU7S>BM[KWC<%EI:7M
P48D]P-VX[C&-]QK84;T4:ZL)/KO#][6H3RJ63,[N:^^1?YT2+MGYV)(_0E?%BNQR
P9]6Y" 4K!'5^Q9"$(<DY!E13TLF<4$10BSD(C8ZZ"-<Z:.H[-;AJ%!-@V7-\)T]7
P[.D<I40CQAL"]2U]$N!]XM+3Y[BP#-$96Q1)]=^#14>Z#_2;A*Y#.S5^G9&+#@>$
PMP#-7!GNU;:],Y"=Y5*8U=^:'?=J$?%4@X#N2[7D =:S#L%_#+8#!92[ IVF=R!=
PLR]QK+\,)+06]@]7BGV[T%!HE-TWFSVG9YD4]SS 3N!NWB:"-VK3'N5?H^STTX3.
P2B,8<\ EC$ON"MBAV[QZJBG\D0ZQ)VW>7-J>ET4#?D"E:F]'*482'8K-MAF!<E[D
P1$ KFL10VJT;P#G5+KW$VETQ[[Q)O%\L (,"2#!'HLI8GW_?X_"##$)EO5ZOK98U
P*RJX3;E+"9\Y-X^[W$ R.!>6SE?0@N4(9&%+?O(T\J<EA5"(B <F+@&D43LU\CVD
PGDC@M%JOH[[-%I5NP+$;W4IBC?\8J92C[*3ULIU-KQ8G9!LFH(763<<&[4;BQ29&
PF91<RM>7[@1 >]28Y#2F9,#O1)BC^SB"$47A&WJ_Q@/[E(H.$'[GW6V3$'W_UP&!
PID&IKR4[,2HY4A,HD]S@AJ0CZ)B[BAGEID05X@5,?\?_2H77&7WEU*?6!=1P3N;D
PP[6\"-I:YG4,U+$B(69]L$:1+A@4&)T1<X$*V&=8646WLWIN7J] NIFP0,3=3Z)^
PP+&B/LU)$Y KFR$1!O"F101AX/J?$_TI@4D=@D3P9BU-;#CW):W-[OR4_",5.X>#
P+DN:\GDMHE,&'<5C3 ;S(-;A^P&3[)TDEXHA+@3TK[C3DIP?Q&^ET[!F/XK1V;BF
PBY@WHM8I7%,"Q?@FT3\QVSB)5!5I"YCE(@9:9A4/<&>O@M9XUP;)EN_W0!+I=H,"
PLQ8 @@S:=T&$ *3]6@)[82\!B*QY(&I<V03+D8B"LC5O&T)@*]+5F\]9UCZX/7I>
PW&HB-2J:8>:'SA/Z.#^'@ I#TYIKT0P0F+?WVMK/?0UAN*T3I1!,]\#S9O.9L#5X
PB5/4/?$N:UHQ"C\TY1"[KYQXH[:.KY[_1O).@!0D?FL?U$';<P+)NSBERWO?&2BX
P^0ZNDO11OS%0G/K/O_;*)D#8$8(]RXJO?[@&?I9=1O.&5OT1.G23W@N14]7$-6QE
P&UI8]*V)T-([>E2*9Q^7I?<>#DY'H-##Y.TC[Y'?/3=U!V"-R)VNZ\+6F1;KGSL(
P#8+CM#"VG-;,+?O,/0LAKK/M(6*4-V'!TF%=YE%R!VT.5/3>;&+YH$:J2=>^-8#G
P<(NPMUOOEJ"E#W@\@0-CM+,WF:<Z1#MVR[[<]16FG>,EK;R%_80)V\.?$M-17V=L
P),#C$2>G1<0"MGGC0F-HCWRPJ+F!&=;%KOEV%J^K>,@< ':,1"/OBJV7$$<\6,LF
P4IR1:6NC,C5$N4JDT JR]->9%B'E5$[M^"$S.^:.+4+MS^0Z@M<]&MR&G(;2]T/*
PWQ/HM)K-86V0UEE48H 6N]QJ3!@]P%HCOA!)^YW'<O;?WI?<7A#XJD'KGO6"![O6
P$QDY6\RXC*@0S(S'AT_AY7J)/YHZ!D)[7L2Y%"GVK8D\V':2$7&K0C>XM3, %7>D
PV28"\L?M,&WGA7K$AO81&O?Y;3EJ,_R@X'[^?U7!_#I1D$,FCDC^]O=$9D"02D?V
PL1FU?C:<-M6M@69KA8:H3=FJ&M&,0.D?"5=7Y(H@J+Z$5_,F:.3=K74WV7$=@@R0
P-G5]C#B41L"F-I%/KS-G+UEA[J3I"IQC)Q(/I6)NO!,<"&@ NL>BW2SU5 $1;\#Y
P.;-P"[OIK1(DDO.F:!'-/V7RT,+LBW<?)T]A=L%N.X:&4VBP(D#8'77EU=,RH4:B
P LD,-HX=E""5>HVGM/:+AH7#'Z@M*CW#'"M<+5.B:D+LZ[:)@PD!T#%?E0 75=,9
POQN>$$=K?18>5#HLGFW#*?8PXB";9E_L(E?_Q(:2!LY!4KRP;9E%')9"8P-YOR34
PC.KYGR1V<Y'8T"UPS#%5]NT!G+$\N_')];J01(Q$KPG0W=3D]JRZU,KKNXG5F44_
P*&/GG]>W41P<DK(4;ET=9560)/-2$(3<-9$G=R_KM965ZHNQ047#!P^DW[$@XM"C
PFL=K[X\U=.%R]:[84]\[TW)4?;GT9'1>.W5Z.ML@^<)?\GNWC]9M7[5I#@K'#%*S
PJ#MUCZ=%DX"W\]%:(Y%7>K_'LKS8W1'O[O>H_**(#'4=QVL_Y3?&D\3RQ\&J=PUK
P>FU@<I-;:T_6,-D6@W'Z<3/GJ7'DN=%T#]LB.DXC5BFV\G9BT5,UC5/ ["+)MKFX
P^F@FK$">M&0?*'0 *L !HN>UNY4OAK\=*LJ91M!63-_DD3@V+_:M<HQQQH$+;IX=
PJRM84P?)3D>(]QNIX/B#0 R1<O:I\"2,[).N_8*WX\;B=<!3450XK,=+M:\E92@E
PH[:E,=?]N+M?4PMH(!$TT5; V,Q74=< <\\X5*0'K2_G)O5G 4Z8V0^[[M.3NZB$
PLX7.UQWV:)\WY)'O:,[U-P,5U/PC1Q8O^KQ;?EAAO^93:V_AHN (F1R\#]R30B;%
PTUS8WV!<)P-EF]>OOR=PT)W<J5$=Z5A?Y*H2\4JW?WBA5B"QIY=9.O\P< FJ<B=*
PI:<\_ZL@:B/XZ])?'6$\D97^_5D*4<6AN9]<KA-R>56FD9"(A3?[/V2]S;;.V.?$
PWH.BJQJ!$XBVH28D4I+;X.1E?<=([)^LRX1 AJ%-$E1]9_()9B3H"^#X*J;%XM<'
P@J0]&:B<\9^#&-Z6-CDN=?^D&"@0+R .26W (!J-ECF-:P4U'+7U([<5L! #R]W,
P2W_;KJYT%/60S1.J6E?',T@?0^XI.;H(#_T/KUD&Z>0#7+ !16.TAQ=M]KWRA *$
P.UK5%!RL66E:BAA? #_I%1.H*+UTI5KE,+KOU>?HG05]SD-10T3>[M/8<BZD:F5J
PW&:U63O>$Y^TCO7@SJL+MW!8RCN@V1,41E@!Q$X;-\N!! \EF-[<M3B'H^J$G;H8
PQLQZCU@&Y9<U='\VAA*_IHJZ/W##@Z0QT,[_[IXJGD\UV/"[GR=1(V=; U7YK?)G
P729E>]PB)G^\[@M\,*![(V<]!J\JC@F?L<!9]8X%!JA,%W>G_J+48?[$6(:VS'H$
PNJ0=:-;/K_O.'7GE%GDNK:)HK/+5QHEX_=M/ESD^3_4(XN! S,GE<_!JQ1-,8S+*
PQ/=18"T=T#H/!H0N@_!N'.6^<@VTP$I*W O_+^K0IL5ET4%%Z]/WS7L?M'&,7#":
P,*=1K511$J"JUMS!/E0],9_-K3O$*-OD'H&OW$.@[=80E>?V*877,1U> '8,5M71
P+GIQ!8NP0*L;[W[&R&]=O/@:[=BXJ,CVM$H@5?$1L-@Z;C+V@L*F7>?K>T9RO!6%
P$(W+SI8L1*T^9KN>R1JQ!%8U*[$D*/:RY.9:VCK)=>&AH9YUP'LJW"*C4W\_@ ^F
P5]/4N@#BS))GDB*ORC?JP&]W%1(-09 (Q47SBQ-9CSQC.12($/H/%BXMAD4[<J S
PK!GV!,)V,2Y&%7PZIQ[)3!=6AK99'P*5K27&+\X^A'S+'+&$QWX;9%NK.D8UY$9:
PP^IM>X+T/>'=I60U71\VI,;YZU\BJ@NZ/"=-&O>YA#1:G_-Q7"(HE"0N]-?/-[V/
PH50HNIQ'5$&B^KUV<6IV&3"):/E3)#=1\E8<0'E>O*+?Q HQ"(08@OL],R*'SRY2
P82KDOR"+#U\B;JJ4N/M'3?%:H-?]Y1JR#4.=-<XWNIK;AG0U2PE+NDG% 0A9*KN1
PZ;Y"B87S%/9\@4MN"#6)S'X0S\Q;PMY1(,F&?!])+?8..ONM'H_,NB8QKKG%;$XO
P"G*=3LD87?R[^9H<ZT=-,"KVO[.'GN\$TZ* KJ<[5W9_+-#YG!U(E22M4/N!<>/2
PF)>2-$Y3^#]/QT@3P\$U% 5ONDF)C3V*O=NLL&K5   /;P&J+6,:.ZB#NA>=X'L8
PEQ'D+'DH?=?E]:RB*?EZC*7LVN!8F_R_,:^O2:@[!U?+^*_:97J>8._TSC>IY"&D
P=,34!-8E6O@&KFHGM<IV@0+86]::+0$:0M6O_ 3PO:^15SR#KB?&'4T>BDXTBZ33
P#5,-#4>6QQRO,>2D#=NK7T5*H84Z)>BFC#[Z&?$F1]AWWC48IO0$N?F(?VI'5Y>K
P#H'3*ER:?E63LW#7MB(&'L.O_N(W^6=W- PJ5NS/W[Y"<4*WN?T$2+SGBD8 Y OQ
PM1;5/F=;QNR&M!+@V&4*COF_?*K7US[H:\L@ONH.:\+.9F0.]S !O4_%E?'/I+Q1
P44<;HRB,A<^$)9^VVL($YMH['/MSR1Q2*I/_)E2SZ!')?->VAZ-J^LE#C99.0TOW
PO;E_(^YP!4S4P9M^$=WZAAI-VWE=VS'<,3MF[[>D,MXNT01@%@,[<NM\U(@6LY'[
PDD_RUHZ3+BIZN!@U>UEF&@R9@;_$S8Y(46N6LJ\/L.UK)>5$;";*[Y=8>L#PTMC]
P"4*FR0@W3,,4I)3Q><3WH9;:JR<'TM^UF5+Z/_C(K_:9W.VX_]!1LOM%:_FP(O0J
P62M ?6!##=.-O=  UJIMLKE!>&IX[,<JD7>LSAX:H1(*H/&#2>"?T;7W5K\:*T7R
P)A-U\!%H:TZPWV@K8Y>9 L\"-HV,@OI8&8(2NF4?7S'_.2L8=A^^,+E0$AUET=A*
PT:XI1+N:QB4:+#\!7 *$6O"Q^NBMJ'P:+0:Q^B3#VV!9:^6*50(0L:?,"O30UL<C
PT.',(F5BTB%9JB4O*0HB4O2C?%L'M3.J)S0@&;Y3-J 45\0)_%0=FD]:\<;=7DMW
P_5%=' Q.']UM!Q-"Y8)*\=?YSJ$ &=<5%ZMRX9YM8J./JW7K\<L2$)+(_25U\?D^
P%8H S8DC/<:8G0#B[ZN#/@(NM?06%-R(+&:")@6G5U79$>*"2EZ>J06]PJA%6YYC
P$AK03+O1S '9")7VF?FD//URL]3+F[;U[=_]A,T6L,)GVHPI;5.$UN63GJ+[R&U[
P]DP&[F[U Q_SUS=G'6-$'_.E*#J$E T7]:WQNQE!\ ^&H@T>D)J0Z8[MVRI$- 2&
P0OT_?_?A=;[6@3C:!\!,_1>-V*,R?%CY+P,=*NV+[915=Q"-]9 ")-C,B;FM;E8=
P"9,:<#^PKDU4U#VOAF"=&P<F&7L@?ZAWHETR6QM03$STYY]?JX&C_;!&6=!83K-'
PMP9N3D[DA\XC;)+DE]\I-:I0*_SA<,E_QQO/03 O$[S="-Z7EW$E;-E!W0_G.WZ&
P\-V[]6^Y/W0?DX,JN;L>^(J2<+P2;$+9N W+.-WY*V](_(R&0XCLYY^MWSOXW5 ]
PN3[&,QEVU1TT]B=O2CEFO2Q@:,!@B!1V3YN5LN4QQ=W16X4UR<$ID5%-?D,RBG.N
PR)4(N%!SEUK\D8]:VB"2K("[_ I"19_@K6X=3:B?5X,;I]$-==<(U#]WVNZ0&/:Y
PDV;0[S.^G?=I767G973$EZ6;#KOB733!M>8F!7.?#M1H(A N!CJOM\>PY/JIA.'<
PKDHV>U::XO[QE%A($-Z1/ZJL37UMIS(T0DC[+Q:_O,1;_#YTL\C'@9]U8J<011+D
PX7LA<$8[X/VQ'#1>R7OZQAU(049X"%.R!U@'0#T[G]NNF5 FP[)L_$]\(<&Q#N]*
PJZ@4KVLIB>5(W/9Q#Q^E0%L=H[@52(\\^_,;RVY,U;&9C(^>HKUT0#0LC4$:/)/!
PTD? "G!:5\(?7^'YXKIP"V/'&C]H(OJ5^J%(0?\ZUQ'K](U (^4Q>E!RDF%NVX7,
PVEVJ'E]CP9GSU= ?Y&8Y(,L>Z,[51<\'AL9[_"\9QS5L>B_<95,H!]JF@!/8??V=
P2RT1>41]WQC:#DK:70HQK%D,_=5A)WY#>EB>:FA\)QM%>;R1EFZ"V  $/.$3N^<B
PA"Q6D3K#WU"79.N0 PUC=#@4MW8=P-U= =<_K;-.*:KY=4?E,^!VC46%3T[U4P/X
P=K%YSJ*;5*.7E/TE52"B-XS5+N4,SQ[D(!?'>!I/5\ISOM/1DOT3]5+WR8O*DBV@
P=84G-AD=[)MY&P+ 5'E^DYKHVX1X]F"=MO60U?(,&'>+X+91&5;MVM!K<>YK?1K 
P-)?,DZ]JM&&OVEPLPRYZ>6245]LQL61X53T)9IJ]WB5T620 X^M!6]^E,>\ 5YTQ
P)H+I.FHT00]<=WBUX-$\<_08*TU6#.)1K+\>@Q]9XZXZM%=L #FO,&1=K7]V=P4#
P3_OG*2VH;?=M]I_/9BK$7NJ/'2Z<9NF^K1N!U7GI>XU&@53@1Q-FT65WS@Z;.& X
P?O]3UEQPY4X'5E8@":R3*V[9I:O0XTKA12=/N6Z,)2=(9R0OI<)3ZO#WW:I5_%[?
P\39XMQ\S^*9$ZV(@1)VE7IJ&JUTFS"'))V=KHI:%!?@OS5U"!S68X:2%@*PS9;K1
P-!C3Y;L_+AA-87P$<)9A&\5B8.\O<:,O/NFK#A6_S;APSYW-(Q"T%^(X3#YNPGF_
P?9-(D?_E**P["ZFN,9C97><2-6]+"KAQ"W:($2"P=+F[,I#E3[4\@[-M9E?UIL[S
PAW4H1?V<(:Z"/H"&^>JMR2E+P%UZQ V8ATQ16FYJD7XJT.CKWK,ZP6G8)$"(2*Y7
PE"L1.';,"]H3/M4J?!H:H7CKD?<^16,J=CSVE\'VC/ #.45.7#U1*U%_V%^5;>HM
PA^+-1_!^<4PPZT+7O[(J47EH<"F6Z9O8ZNOX4'X)9T;J))J2#IRXK+AE^\TZFTG?
PK0,04>=^J*=&@"2+7\U:T;7).AE(::0>!T9=<S51^&18M7V54V1II^_>N&D!Q7DQ
PU+[XW#WO$CC<[E:Q/G$/+%J_VT>,$#I;I2LR3.O/(?F+07#.;H0WBL#Z+:AM\!6E
PY!I&;@IPHH?'NHD7(<.RLL9 ?@2GO$DDNV)*[&1.)P+BHH&AMHG 4G$&6W\F]R[J
P_^U43L7JUQ#[)(=7H\!'VUOOD'-NN'@A0#D(4VO/1(V:]F>W[; :^ML[828Z\W/:
PQ0&!Y_N]99YH7VP84/["4Y)[/E76[:>YK:MS$!MV?UL[O8!*;2R4MCU25M5=6Z._
P.@-9O?!5=4WO^W#0=ZWU][X\T 7^0Q=@NBUJ&/9'<F3,@0)W<_XAG@L-1\7-8QB9
P31X)XY(>LK]J)?8)R;(]S>W/MD]X-IG"JWB/F%9=Q+<@"M]\!'Y9PMUY+L]] ]O#
PV)]$UOK+8 N*%^#-@V3BWB7*ZER=">P-"2 IU^R?3NVW90*S80+QR70N9NL?;BB'
P 5922<,J#O>]6]_B@-88IT8*J<"^@R35)/7FCM&RUY/@LXY//5,T*+N0E.JHPU8!
PT\T]6P6RSO5E!U*D7O162VAQM0S]Q4QBJFZ6 D[VW3[83:@SG61@]BS(T(#Y!;GE
P)UVB5Z"W7<79EYWG.P3EHSC1&;3<+9S+-1,EY2/]1B'A=W.&LZQ\]R_H*2=]O<?*
PGACP[4C,3H:R+3(0;??$D"2J5].:'Z?]!)-W,[@PR%+@8-/4":"3@2'.U/Q%(PQ[
P!R%)<-MD3K=G#3PJ_@]U#8:I.BY_G5:[P;I='JZ!W"&P*4GNY6JL_;W:ZX/F4IAG
PCQ&'I)D+%"=$W*P;DX17[NWHI\2MU$.M:-7;B-A3T!=QDO1;^]WV)MVH\K8'X9BE
P77SMN&!>1"RP+#%1H::0J_+-3>6 &;"A96&H6I\L872'S%S4HN%9;2H;-YD)J]#7
PE@_1H?.90,;UJ]J"#$3,8D)O.]D7ZIJ'Q.0,/=/%AA24@11W=%^#??37^:0_N89L
PO.7X2F,C\ HPG06=(NOF&$@5N8?10=>UP>^LR\XPH). C@]2-+%"9T<RN_*G+*1M
PB&?&D<(/@)94)Y46E]ZEHX9E1,)^X*&-W:JPG"^W2HD0L09FC3^S*J+3XT-R=/W?
P67I 8\(ZHX[_<T9ZD1*D.,?21-TYH=&=P%PS,\7_$]0LU@)D:M]*D.1!VTA43C6.
P9N9=M$3VV"?>>6?@0L0R00'<% .M'NHI/]>$>';[*Y,:(5')RK6K*(8;=A.G:_UG
PD7)1,U0P0]6=\\96>1[$L'F0CP#N].Z(#P1.I0\6V6L880C4RQ8!U<\<##NJU+<K
P"7I)5A15>TC0FO@O]M:I>=DD4^JD$NV8^.1]7;_B"Y$RS@9X- AX2DGJA<,*G?KX
PYIB05-,YB:<Q^?16@;2"3I.A#)*0:.0<29[K1\_"Z:QW:YZ-39<\JC,3/X:-E6^E
PBJ0>]N3?@'/P*T0P$P"V%=Z$[EM\AUOP9,]:+;=%F--[PSBC'P7J21=M7KZ/Z[:W
P-13,(MH',ET=2.6G#C]TDL$Q1%YVZGKN1V/Y<[Y0MC?J[@4";*^U#UXAG)C#S6AK
PE8OGF=?.^!!,N?O6Q5Y3Z 07XB^JG;:@T'*B=K/ZDQ]E.MW;""PG74YHW]E/AI%M
P(QTME],WV*9_$.4K+;R75C ZJ1$!0K _G$*JL)5*YX-WG!5]L$_&3/TZJ=U\AM9.
P/]^_GX8/DC;;:B#%\<&W:/7\"#4X%:BR0"(P$]TGY4+?')[I?:W4)P*(-%YEB$0Q
PS,!=D,0VZKUV>3D=*^=FXVIH4<:V,:!QVZ&WB/7A01;V*SX4LZ[3&0$5N8W^KH]%
P[*GRM-"Y.N)J NL@F>M^HPD>0<,ZO/L,P]_3__P7=L ][12M2##I<YR3A#X"($3>
PDLYF:QK @\)^3AD_I&GCT5Q]-F!W_#G/4ZV".BAVVU/QF"A3 DF$,9)GJ .X!>N7
PPZ_\N_R3C*8?&7\G68-UG3DP]R;\V.MZE70<[\/1TVO8?5T#6W8@J#:%Q^Z0\RD>
P>)_GEV1,5F,F_X"0PQ^2>@&+$DMO/,M0V>.UHI3E<<8FG<&LQM/)%BU2.[,.2!X/
P<\RXW6KZR'5:M?S.^G>'"Q=N"W,UEK&2(_DW;M#F)BSCM H:S\T(P2Z7EO!Z4\(D
PD-KX#>+9:.T-Q7*UA_N9IZDFE@3Y&>4E:36D<RQ\[8AQ!::@\V(EAXKYFN6Z;].P
PD@/\9GG@%4*?QQGT_GS2L]I-<>G2U>$TITC$G"(,]O]G!UV.A!DN>]4J#)/]\6_N
P'8HX,,Z6$YIVL3C8O-8*&MXKX4\)=L,X^<,N)FF'>3]AAM ]H>;$?:MMM""-K=EK
PUKK?;N#F*#5=6XA<GQU5#G8V$MSQ)Z2[&@A-(%M_&*,5_JU'M?6!H5]I=H?J'^,R
PF\/3'5<WQ-&_!-@5H*:A7AU@J@V [V4_7"WIR/):QG1.+FLP+DGZYH:2KG$J.J7M
P7X.TDAS,Q,"W_2;^RNVCC]2AO]F-_Y0VN6LH%G">4'P3\<*L"BS]=(.B^O+;&22Z
P!BGYRC6]+*^'G)B\]B8:FW8*#BI_.X/I&[H($#SOM9GH/:2GXE\XQ/KQ\-@RZNR;
P81*SI!2IJF5#H/#C+*:4A$QNK8JGTIWF)&<JVMO'F&N>%(K;-4CE"/=<TJ*8RJRC
PK":$1%$?\)M3%D[6'G:@]4Q_S]M@6NO4"QK@(^"#4[0EOK,(?:#Z9YZI3?;ZS'$T
P3-6T^]/';EFLV#5F?HATANR.->&J"T&@0.1(?*85MJA(GW?4=QQ^;K5DQ."''>K0
P>O?C\E=HS$<J.F QLC?!32%_'.,NZS_^B*A_7M=8G=1&X#[MM6!>U+<6)2_1A\\D
P>2(  $:,5S70[75_MI=_[E"BB ]&#<6NPIP+1Z9%&%[JZM!0ML\G$4L4?UB9$F8K
PVT8.6@.'9 3"YNV:H1M77 *RAI_<H*PLH$(S^C;[67B\I% Y>1K98Y ^<U7- SEV
P&V%?WH=2D=[[ 4)?SKX^UZ>M,;<?D=L7FI*6C;A82E+OIF3+UONLE=#-6D%V=8S#
P!@2G5@:A:(L%XEVMJV* -4Z%HG9^(Q ;WX&C;"2:A[CC%!=W2W(<7^2+($<A8/%8
PZXRA!^OTFBC,CD2I+'3?XD#H#N5&^XREKK>YJOVU )\$U[)W46GQT+_\?R^N@'A8
P]H%$XXPS7PB_@J"G7P7<DC&S(^>YO-8C1+3%V;\TCY?4!Z8D'@1:P@WHLY_;A,AA
PAK0-^EY- 5AJDH>2RWP18M^?6UGK=$O6P8](4YH:/H 8F7;(,Z5SD$+P4SMW6@[)
PZ>?A"A)F9+$F>X'N7S[[I:0P)YZ"GP#K$PUS^B$L#3&C.$?@!KC%2G#\QGSGQ -S
PO]6@C5SDM=*Q@-ZSXN^O9U0= 0*AEJW;X_GD)+7YPK+,<+THJ47??;)%WBIO^(6X
P1H,)\)/;]2B3N+FBJK2H1+469!P%W6@0I4,L"B%L?SWJ[TT8!(Z&AM2'CTK.G\R[
P]*N'@PS3?.[7,LREG)0'#E8Z>"YL[=@,K89(5_#OZMV%8_M(V'EV^(C@%;2=(@&:
P]P!54H^\G\LGW98ZZ)=B]>[F,Q71CUSC#\"CYOYTZ)^U'_L4+RN-6[0BMV--NH&F
P4<#H)H3?GT\97]^.*D8QCY( $N3/=1QGH=$LTC,-('^X%3$H9"90\>,Y1F*@G$A;
PL@0Z$CJ%>LL0X:ZU':$DSAGHQ:N*HY-NQJB_USI[=&/H2D^8AF:;V.0'R;R>LR$=
PKL";I3R:*"R[VP*Z]5&MA$$!.A*CHU?! A2_%T# D(XS,FBG#9D;!Y61/)=:HB)O
P<1ODTN9"AJ*4>SF)GQ[_B*+!00]U-@KX.0ZI7+*F+0<G!'FE]FB5/R&N3;*_J*=.
PTX4NX;YH:/Q^R\IUJK6 >5>"#ZB[#>].9+H;-P/<P:Y;]L6[07B.A39O+0!4\4 G
P#TTA(63 7Q2UDL+WL.L\8$T] 52; R>3-!65G3TI*+EB6??/^9L(O2%]@V(]("42
P"U\X:A5W&I1##9&/<('-H]N')([Y8+&I (*3S67RP E5LVO0^,+/<RGQ XO[87*&
PWS5EI ^<B9[# $B^=:8-T-JDPXJ 7[#'-5;>"PQ%J6VU.&LE] DCAY;U)U?QR1//
PV-J3E@"#^L,J>5^M;1G:!*P!OG/MYO&&1G]2E!Y'.:*=0(X-A+U(7!3)U:F._"'.
PBOLC0IIC;23]N1 "8$1UW\+R'5D-%*M0'2H&_@4M+_;0\[&R&%KY'(Z]X80<- E&
PTLYP^WMX $@O6U:&=W!AF_/?Q0;:R.!MW5OH>P,;'Z1G>W5TY/=G-=6M#AR8#FVH
PA:EH)U5S P-7!0^9E3]-%KH4 ?=8_$=T59^W.[3>J*ZL]S?*,.D*?+/_'[P*LGUE
PDS0!'GN[K_[BT0PB--\]E]3I[DUE>)C]<M\W90!W==WBNAA\"E?Q7(B@.)5?;\]E
PT+)MDH8AF5K^(ZD#,#F!36%Z#-)E\(.K"K($C2XB-SM_Q :B_0_D)8!H 1(S$!)U
P[R^I;?X2'G+>J*AW[VI!@3@W3^ZT>-0@?:E_,!*R-O)SM#L@D, )(42LV''OW'R:
P%1BVAUC)?%I@X7#E(124N<SO)8$!?* RABH.D*D$)-OMM]M\""'+Z(*(1P>G<A*A
P>8?'K&3Q9B5EU(QP#?$]5'O?-:,E)/P>F![1A.(W<-:IV;Z7AJ/M=', J#WMUTFF
P+X<$#,%/MX1144*$IJ8+Y)F"(C=P:$]TR$B4L]G>#7)\X5!^XEV41C_6ZC=-F@L;
P&S(MR*'5!:6YX%6'Z"2A40J+MNMEM&\S?21F59)J*L,Q BSR*C'0WHD.2M_;B?HO
P17X&;R+87^Z4LK,GB9L%4YX\#;"H^*%<:9"=0:?_C"L>(I4W,&+OUI5:_L&K+?A+
P=9$+![6TAT_^Y1@_.EP7L@]@[!-WNY*!"XAL9CK(L2-)/1YV29<ZP&&[$78&UJ09
P=U,^V- 5FKI/E+H!X^Q,;!"_A<9.[5\<;N;8E94;337MV'9G>6>3T[7-H2]3,U#8
P+:"!JI)13*'H["?+,M%[ .*)O21N(T[=R>,QKTG4JSIH<#JCA*NNE7?WUNKZ)U<V
P>P+PV2DD>V9# #TF7;\],^@8D0$X+ %*>I@B.[96&F98#"'D#E-"Q7W-W0>I4ERS
P56M@7CZZD:R^ZX\61EX@.KJ_*(PC=O?:@P7KD0LJ*#>52EM0:*GTC4C_E<;5#Z9B
P[KYKP.*5Q F(>/%%3?T]Y YDRDH^]P[AI8SHNZ7*H.SD%%)Y=>I<%<KW0O-;S"=4
P!RUHJBA"6C\H"=CB)JRI(UO& [9_ZD"Q;R7P'H5!5G$2/&:;.;G0R2KG/R4W/@V]
PT:P2* 23(_W:02Z3)?K/*WME@)I  +XKAPRIER>D658HJ*<[?N"T((G4N-+%.#4&
PM#Y-3-%6@X0B2JT],94'EG+JA8VB9$?+'WN549FTF<&]%^QCU?*'8FUX;_?V;@(/
PP@"PA*0.YM&K1-:VD[9GV? 7B(@#0W\B;;^1T0T%&I".#^M.27)A"/#O!=)70$7F
P5L,'MNA*N/D K#NK23)?)8(S89!O57&CHZ>D4Y(5R<0-1 J5+DE*@I]^?+WWPWL'
P;+\$H*IJ3&R@V.==&OEY4E"8*J*?L+G(! 52[,;W2=(.R4XQM@97_5C[0U4E3,/]
P<72\D59ZZMF!9ZFS9_K:*XK@X-<Q1B#E<BI\]S7VK)?E_FJYHXT%(4[_44Y9=:KQ
P#U6Q',)Y2#HFM9N9%V"4P,P+/9(,O>'GE:Y!@!<GTMW/=?@IA>E5"]%M5JKFJK(^
P9?+(=85K IQY/@<IAYT#M-IL::"!9?,%HE]#/)='7'[/OI0^5ZYT#K0Z?\8&MWA_
P;C^'0B>D4YDGPA<5'BDCI ';8#1==1F_VHV_"[-G+DTC5"ZU4.<4%%R%C)B1%G9%
PF +C0?[])+RLJT#%,)[1--5"B'0'CAZ(BY##+3^I JNQ3K\4/%X7HJ5=_@\I$Q%G
P(_UR.J=@)&/!(2JN0P"F2PSBX, A.D@5U/$,FCR*JF;34+*C*/6@_6K?&5_Q*I>+
P%2],Z#YCRTB%SZ=T-2<W5"%396&<A12#JMH'HZN!R:L'[QZ>\\34ADDH%1=+/:=,
P?+FQ3->T0:/]]]1NKP>X J3>E&.7/UJ,RA%&B5] QD<D,*O)&I&J_]09JPY;91):
PV18]3L6>D%Y$@6XL?JA%_+.&/RN8Y; WU/E_!##CJ=_;(@C4'-M*NUP(!' R%4&O
P-C.3JJTB]M5$0/&VGT['AYNGIAW_VL;FH"'&L3Q=^OF=$[UD'#H9S\.^?NZ@O%I8
P.0L)KKDWME(PEU;=Q3188?VW7/0!=VK"",<SJ1XDY. <9G23"?Y.8.%).\>Q@T=(
P<*V<57B%9BU>!&3Z+>0L8N?(X:2D^C% $Z7 N5JM^A9OANX]8@^D?GD0=Y.>2NTF
P(\V2I=.2,+&>/.D-?8&-)N5#+?U_@?%O+\9ENCI;/NOF7F(I JW2:4NF93M8C"$3
P[6'%^D 4R%^XDNQ&GN4A-;_DD]>)"']SX5/QXHBHPA9R(#0548K'HLA/0+.HUW.0
PE-@>(/U7PB_)8:5KHA6=WSQ(+K:@Z\ON(%;QOLTRB!8EXI^1H"H%"C#>TA@BGLQY
PM_A6M P86!4HO&CT'#EGGA1]5-@TJU-<9*=?.$6<#JH\#\-37FW,HA7\8+ 8T<_S
P/WC4C?EIF(.K*D=H_X<)+1.\]MF,])%/855[I*;<:)Y,'8Z('" 9Q"!'H9;=J/*S
PA$7ZP@K?V^U1&W5C!.>?RU>);*$7DKX"WGPP>[[7K&!%)"W>#8YCDRF%XY(K*D@N
P^.@C2\'.7//7[JP  XI5/$HQ@(9\ G8Z7BX\_%GS%"GWI[/<&$N]=XZE;^)Q<AL7
PC1@@[5#59L$^)&UZOT)1>6O\4U&A#C80JCD6 V!#P84.A$>L(L)V?Q:OO]"DDJ*E
PY\DQ);O0%7P_>.'O1H<?F1\MBHQ^(TX/C)$+_,#7$-DG'P9CJ*<=*P'Y$@0LI6XI
P^,%.)X8*HKL[AL*M;?1,(+**CQ!6I<W ;MCD291K;3'2V4>!71CE77A'$Q"^DJ7]
PQ/AT792C7=2K"DSD*_P6UUW"]IA#&"'+V?\QJS Y^I2B7RR?6CMJXU)./&J:QI2$
P*P_W?>RR3:Z/3ELSS85OZ'+GK@N=$V5=_B"'^W8]X/N?)A;/\13YN5&MFF<@!%,#
P.C/3*XVY/N/+NEPA8ME(?F.YINJ$TN^"]@M[R W/X8L%W_E5887/8WFH$T)[TJ:>
P*\R;8M.XO#332SDM&.''ANA#YP.2K>*'52^?DJ@=JNI\>LONY==G:AS=5<$/U-' 
PT/C"%IQ*3+6F0.0JW0D\B>(+DI42 :]WWW(!RFND6B-<M4;LAGI%ZW1TO@)$,$.P
P?D"+0 QF"6QLR[DO;<QHA6$6D^S+43&'>OYZGO%,U$_J[H7Q_[E:SG2:N>".3*%Q
PB.:0\[1@!/R^!M[ 4PHXB0Z;RSZSN0]_","BDZ[=I0"UNPUZK7*DHJ%&CF.7IO3S
P8MSM.O=P<:TOU4/)A?W4#X8NQM@W0;K;BG^TA[XCX]'VY$D=TW!DW'!&$/[=@ ;:
P:,C?#=C?FY.=.Z$/;?<RPX/,09^<8* "F5)GPV'7M#E^5SKX#W!5CX=]X+03]C^\
PNX$YL C;;KR"N-V68R@6^Q8=JZ.*CM$$EU%M X9=65)MA:Q@P@\R=U Y@,SWN'WT
PWEFB,5UF.L=N?/ZGE%W*K+K-N8RNRM<^+0WV]& -8_,)PMO8B!UZ0^5\E>P?X>D+
P37Y!Q2#QFNEZB=,(,%;7=N=/K.M+E_A "3=* UT)GKEU%C?K>_*%?;\WVT-Z\"=@
PA^F=+5DL86CK\+^ERV/\K@/_ZLP?ZDM?;-NI[IP"RC3%7UD%;*RMO>GL9G K:?''
PH29''=7R+]."HT0F!.E2DA\<+2%2D;)+JO' ]%M7!V^\3(M4V4NSI,!R=O40PVXT
PP.ON]);\^%:O%+T[= 6VCH"\$M$?6SFQ!D,YV^(P]1A%R9Y"897T>X*NF[]KB04N
PPC^6#"*!B,E%^WM]>F(YL-.Q)_S(('6U+ULJ(!G.6A4M/<DM]F'URMG&0J9^H$:>
P'JD/;)6/9+9;N@L!!Y('J&TF1]QZ/HH2'EW&2UZG_0Q$3XQS*>SUA[(@/XE $:K!
P/QY"T?P"U=0"P3.>IJ$]A=+<%Z7!?$][#"PE<W%^,8=<.[(MI3H4<:'JZU(R&EGU
PN37<#[B014!Q2M)\2HK(FCYALZ7]M5Q8V<,ON]VO$7<7C?&[@126*!VP>JZ(E?$$
P9C/QO3W&]19#,KAIQW(7Q5;;.$D7BOPQ-QR:8I*4%:8^G#<@82I3"1+#)[7+JRK$
P1/'X2')$Z5AB8V87^0M54+K.N C1&>LE[EOL/UP+<CV$OV_X"V!\^JY:__ 0_$]Q
P40HK22G#<ZS('5S<M>T*72&<'",0CZ:BV4$04BAZ9D]!D=YX=BY:._P]#3X[%F=#
P:#W4O'SWB#M9V 2:>!WM?(ZMD8K<'K2)& *&.>&I(#D(&AU#> L@7[>VVGJ&N/-R
P\KV[&)F\0,X3E/'"Y6ZHK#\*J:'@F#--.T@KR0OC)64.AUC?7^\KC<^'C@64!^36
PLI<.JQ:G!'K^"%)E+$XWJ[R!([B/O% YBFB@:;/KR#0!\B![T'(9=8%/S)P\(N^H
P<%.C?CD!>!7\:E6(C'8'\)R8%5<S_0R\&D[2'ROKTZ60? LW0T]#?']: (&^C(A)
P:OBL)AC2K\$FH/$_*(\$BS$T #3IFE!D/)['$P46IP#EZQ42DEH6Y*^U"@OK#H&#
PPKAVB,$KL42ZEAZVVL:G]$?J%_"BH@88IGLZKYY+#0+_#.-_<V&COYQ>*-%*K*M/
P_7J=PI;O, 12))?ELD;%T=-SX/Y9/=_T7M3K.YTDV)S'/-<AC/PVIB%'5Y14G*6I
P&5*IX<K$&#JD)&]\C<WJ<*<QIX%SK[T/H_]__$8KD*.K%'YGN(Y-4:<K$P/.[LI8
PQ0*TEKV>6J6@]-AU36,GR'KES]%%8L\UM9G(8G;+%J5I6?(77*@N\-Z#=DF1/3]\
PC#BEO,:MTO)"F/Z<POE'_VB:"7JY/D-%WNNH#^3%;E%;$Z@D?I%H>4"<?X2!:W<4
PU\05X0">Q:P1D#*,KM1Q6^3-XPOQ?_\O,8UH\Z=^R:/@C'DKY,D=]3"VSX#ABRSP
P$A%YA[AM<U0A[U[BF[&*VC,'#YFK1R<-XWR(C*/W?9[D6=6A\;@O)?NB'D=?5KJP
P(B2DET_F(JH;.;+].*1\D&W(DG/WC7'\]8C?&ZDO$4H[,['V"Z^4&:&K"!2W,.$]
PAF1:%L4,-^EO?@=H_37D0D,Y68N5L:+"^35%#T1*FPZ^ UU'7-UDZW9(%G#;HJ'*
P<9X<U$:@N%:75X!5!HWQ>929,]F!*WKTV,#;;9::Y>^3/0:8Q* /GBP+8DIEV_<_
P#&PWN RJ5>%38[7Q7ID$Y92>NEW$LK-BVBS)+CA,,P+PBVN9F2F+;KWZ/J'9U-^"
P(^W]#%02S+%);2:(Q(/\K_L=].IA).=H>>!']3>.2QDQ=8),?V%W*L-2P;K@!SN?
PF5:4H$*IKKOBH[F,Y;ZY,\M;';RW*#_'-9SK-%#,I?ZJ+D!Z2G(1-1@]O:Q66(U*
P:/5'!-68'J7HQ[8ORQO\ C$#Y=,^,G[GB,YEUI9O,>D+X*&U==Z18'L.^[>N%[F5
P[* QXM];ZE!:#X!$5,]'9P/&%.-#S.S/D,/"<;GQ/T_BHN'C#EI,C%L5BS:>CE!#
P/[E(S/B5C]Y\&3BB':X!HIX25CUQ*$LLYHD@UXRJM?:.:;<A0R>8U\OCKI?^]=_S
P0=HZ!6O)T%+:KV:]X97SALC1IS"7IN1B!IS4LHPGFL[4N-\!ZM+5D'A!5N1T7^N=
PS/WHP7)?\0UNS5L?I]_+BNOC",FH,#HT4!Q@"JN,_P+'/<W[7K3D'A#D!:5_V,$>
P&J8((+K0UGA8?WP)IJ_?/$BT4K?GN]XY-I,<NC,'4C6 UK?*4:X%T2IV;K2;4%5)
P?@?>_KT.'57EU/+5'^5?5.V<5,'KZ9/U&A=.(L"I'@=H"AW** [A$UE=G+)MVRDN
P5?I%O4O!12ZL7#CFSX/X1SU(QK)9#G\@W)4($6(7D &7*FVV+O6_P=-/-/N-KM[M
P!72K!I.-$/D_\\V&,H%.<%F%XI(U8)@W;$-M]_\#5.\+'?9.YFJC9ENSI??#6H 0
P?!=IKRKAWCLK,21?%@*L$!6[XH/'S2S;=U*3<'DO$ /1/D9 +)#G<ZN^Y )>,:GJ
P29Z\.3VE9DX 8U@^D(2<A7[V<FJ3R"45M9G+].%_&<'?<T0O1AV0W\F#4K9=R6QI
P=OUUN/.W(K2:?.,$WQL2MKR/PIOV<8#YCB+YJQ!::_O"PA07C<%.R'@YQ@*OD>6N
PL"W2>JPBX%?CV]XD8QE/ ;G>7TN2_$(]*9W%A%7WX#M&/]95J="*AI?:@P KD:5C
P4;,QG[V82,Z\\(FF;D^5V L9!:$-D=F+UR,SNGN(YDPHGFEDAB%O1<U0/6VLA$G]
P##+F.+I3)=D*O/ 8;P[H(E'[:M:P.1'\S&@>6(*Q@Y4\J+P#JM-@_F/OKN4FO]KE
P&Q-^&!OL?54]17]!F8OP@]^A="#!H&LKTAD (P3>09%BD5U?5QBE UU#K+J"UZ >
P$<EKA:#HY>L1)7\"K^%L.MWD-H%Q(=$-R;*UY0%ROAX8UWJ\)1":!#XMK_/GU<54
P<&TBTTL3S06<_\D$>VN_X-S0(2YK]5\<M<07;E8N%LH'.6%6/<[=2,B=900(3>B-
P%/=5NW1R,5BQLW&[KKX_)B!5D\RS-[4^(LIFDLLL29# 2R8M+!$_JP@/J^2LQ%G+
P<E(H&]HWQW0M["9%K=$Q \I1O9');,3"]S;/-A6<NVV1BE($K,O+/5@H;[-(G(F_
P+*["X2Y[Y4#3(\>. 7P*JZ71=0EBLX3_ANF9P[&!P(^;YR^VC/BJ!_ZSR8T:7F))
P=]R"8[58!<A^0#&*I(^3$$,&NDYQUG]D,#.!NPT^16C**^Y:"2]3$2WK< $NN>CA
P1HA2#(6^M-[&1SSW9V :)>&Z;:*K6,>GHNU<@0_2TRS,(O$^RD7]5WW&(2\? /CF
P\Y<0)]-!LEWJL]^CW5O?.$QSL@>XSH["GN D)1-!J %:0C*"S;ZM+88CG T/29]U
PRG]AGO/A/;H>)8>4_3R#!H_QE8<\43:LC48[=:;[U#'E@LGH*87[U,FH&A&,/#+M
PRQ:NIRP<L5&:P@K4\)O)=PN(W'&1;ZKOJM1S*9#"XZ=-;:]*YH@8VU+JJ9,:!5GE
PMOG>*.90VH&J0ZN_ @J%O;KV+*WI]7EALOH+CBT1([Z<*L4".-2?@PP(Q^<&73?)
P2WJGH%H(790#?GDE5P2EE&M-C$ W'H1K?8E[G,3!2<\$J<?<.G931RL-S1P@$Y?U
P<,SK;F:1^315S2>UX\2ZLG6YK)W^Y@:.J49#[U<%$":Q@7M^]^_G'$$Y\A5Z/#);
PD8FB"]0JHOA6R&I$O,XHD7#^)<E?8;".E$B'RTB1B\".89O[RT_S1SWZVE1$N\CF
P:=C]4%5)'N!PKR<I[/VIM5B2B_D*A. %\'^G=><;]F[!PY$G'GJ/=T058KBYEK>P
P\O='/>.A74PI43;@KM!]8_X-OK[32.&\^:K&,C$:XQH+L@A+P23R//X$*IV'^*G(
P)+8L]'J(B7:#FW0:]#6-O48-[ >I(Z7F+;/' LCT]T.KC.,CH%?^7R'L/[L,BL\9
P.Z(-:_RP-WKM^@(W[9]7+,*X7+4[/F;4T#@T;7C1G.SMYE:M*INCLZ+\8UW^A"<U
PL&<:]J9P-9;&:.0;Q_RD ?0U+I("+!Q:.'QSKM>:ON7C_K.[6QGU-G0N#0[^N%U2
P('G"4^2TIAGYU$BEJRYN!5@K 1D?V'F']H6#[7T%'!D K8-;+^GEAG -D5.+D3Z(
P$Z/50/_N41,Y(NYEQE9J^=0C,L.=/4,(:Q*.H,CA(FPX**7K9DV1KKN22S4Y.,?L
P1;HL[M7T5NAN&/-CIZHBZ7X4;6-P;HNF4(XD+5A@2&5J/0;"U7==_,Q07:F?5V;!
PV6@]0MN-UP>H6#=UPV<;3XK=UHM0^C5+_A_*!T'YI^H15'*>[B5YM3\Z1-$(R[V*
PLCN.:4+(Z99,7"]U-/M=(5'=V-TXEZCO;7+!;5_(1'**Y_Z7FX=7[U2[*:8_5L$'
P82Y_^,KV^WS*W17D^=F#;!8AB#Z*I:PF W+5^V9;T\GJ\PF<A<4V['L;QF7< ?$^
PY^&2S&4QR<!,,,I'0?IV8UEJN(?,$\;2<:#5Z+*]:MGH18>N00JK;2(>WTYZYMB&
PQ?@Y%(\'_DP1@.&[=.CU,4]<I71_?Y*=^Y%UKA]X8CYM5Y+(=.BJX[5*4"XW[?YH
P9&9QF6&^2/KFUDV"\\4&<UB*B,@'L T$Q%QZL1GA[F<B<C[ U-H2FU,'?-%8P]FP
PV*MH05JHX6Z!>+IT8'?L9;KMX07]I+(/G5MC<?0S^UN[N[S SA88W_7,A=.>VM2V
PA?BB;SX4X$S^;@HF"<9 81#% @R!EMSGG4H&(\[]V@6VHM\K_+:7$P#K>8%QKD(X
P>[SEBUD2?R+D3:R]F:["8R[(7 >W@F=7&2^5,0%E!67'-=ZDE.6V(1WI-D-'[#G*
PUNT").Y5WE69.>\=RX+<[F8?HJD$"TM2=0MP=I]T:3@(HP1]%%4Q5_-BNCD-X_.L
P,6J-A]K'2698Y%C;3[7!NH@-@N>E+4]( --S@NA "%Y=YQ.F5? WEKRZ/G<J7)Z6
P>KNP;@1>3\GZ"HV$]!KUNO8=X3SW#P$F61,-VR:=UVR6*/DL@[_E;'%@V0/'8BK_
P<,# U9]ML4K)[FGN+N*(&X1.0'%5JUCU0^IQZMZ@EQ6]978D$\&(03ZFGB(A,TW 
PP60TCDH+)K2&6CW8^2C$A93U9<M*=IXAPV[^@D:ID;"@7NAAH7 J LATA-?S4J<S
P_JY#1IPXQT/(DYN7$-<H$DGHR&&VDN2.@ G=:(G"+R@DU8!%E>DN4-;IRDW>["X/
P1YDU]75RK%DU]/K9]+=;<U=E-;QRVCN'TATZVQ>_+YETRI&:2:(_?,?[KZL"XAK-
P$_#%DCY:#+=#_5P]L)91AYU279S^5T>#7U67HC(\AH'F4))D@9S^=*F<K7P5-$YJ
PS]68):5QMV[]UL]K>1-Z3I/3T('&9(SZ,T@[<>-$#=V]N]XY>>TH^MR"["XKN4[L
P1('ZK4E#&BT$)1 +#2%]+.B"4#XR3^$= 1!%E1V/5AAGL^??U(ZIUTN2&9',*],N
P9R)3CU+&^QOBBDQXVBX>5^5CCX(#E_5@1[2[6D/2=@MCBNPO4]3#J4L23/3!]'Y1
POZD]9HYV9(2B(KFN/27VZ%PX6GDXX;'$>*^^((NSOGQ5L>P^\$ZB A5I54)XR7'U
PJN\55&16Y8V:B;LOY;\)6L$>P97S!)[0TD-W9[3RL)G(9-!MJ3RHR!9P!0U/I=DN
PEJ9S06G1V0R*-Q^X3(!5)EE\RR+Y5$XY^^\E;(_.[:E0&TH"1BIK+N% S_\W)9#X
P782R*UF1U(9(:YT"Q#R ,3U6I6&3]N5N]ONC>S5[2+K+IQ(IAJR=NY^O[:1\(E0B
P)J\<%GV*#.PAX(FA%T!S+CEA<_G42S$)6B45^GP^#T1','2O4#/AX=89K2%FO;$Q
PUB4AD:-ZV#OPFG[W,4,-(8XE%17:4OC<!&AGV,35P"DD=,]CRG?HB];5(9+SE79E
PP]Q"?Z?HAOKE-*8]*1@2+:1>M*3")D_6UQ:IK09,RD&+D'Z.0>:)TKO.U,+B#J)J
P5+(==9?X[QN K 6=#F+7KC3#6'+\CJOJB;ZK$M^MC.NXP=>+! \%DHS7G/10M+<D
PDJ]8G0F P#1H%R!!QO\?*O>E79LJ ^P02:G)_:E\F<;XI5_MLRHT98GBG#3/V*7)
P!_\%A5H?PA074Z-],?,W+U<%7\C)D*35CQFS'EAK&=4CY(W=KPJ']#5H>52*RV$4
P(6N;\VP!Q,-!>@U[?P6 1P.\CEZ.]:8[T>-KN%HK&JE("] -)FL3OW).==6$=_@ 
P#/*;"IMV.C%]9+T7\U?YV>FB]YI=.BX6:NGA4$LDT^*H1AJC','7;"<M5/[(F64G
P+;)<(I*EPKOI4VFLQ>,::/:K2@F2)ZMZB?T1.GYY52T5G"[MQF3]RL1/1BS5)O-A
P"7R] Z]TO(W"Q/3/80=9>)B, NTR7+4@;#R_,-SV:_SH[;P9/H/0'DH:8J-B0[H\
P8WP2ZB![O&3\];]JW@ZW\(:'T 5_O4X*=1A79:C^<'F#I?09L*]_)FSI4OQ."S:*
PM=))6=.B?ETV>6NS;*0*Z/?F;GIAE\$U-X1R]W@DK#HX@>Y48S2@I:1F^?R4,;F>
PJ"GUUSQX:KL_E#[G&)%S0;J6?-9=3Q"_]S*>DK(QBM(D@LV)L6]W[T*LC) DR%"1
PZQY75'D.H41LNDE/#(R84I#-]4#61FD4$[Q3$S$\L=&N*.7*%[YZON46UB%&^">@
P?MUH*9=M,&ID&T#YZWYR]'!,H&TCI&\M&:@8*+#%.#8DQ/X@"/8/N!M^"*Z;_I'5
P$43=B2M<H/4O3#1?FV!\669<Q[WR\2!:+0<3[V08Z:@!9Y?OSON8GBS7-BBR[A3'
PP',0Z#L55AESD&%7=51A&@_]?>4%EL(?8)8P7>(@ 1GJM!,2Q[82I]]4%GSL !$W
P D6T<FKFZJJ,DYN@GUV+*F?'?+;?KLEW&%"O4.[SK.BN;;%SVDE_MN";U-T,"&AN
P3POFK:TATRBYZD"_,[VT2?IV6.?;C2M^(TOO]'\$U4)1?4JH>+Y%[%(6/A\B-0_;
P%VLJ<O,6U];Q76@;0KXT4'<0/RRKRKZ9L#NX"I/R6Y-E/FC++G*Q0FJ6JX\=H^^#
PE^V5/L'\\("62957 D[QPT8+IAB#(K-LCI?\0C]HW'H_-SE!#(C=6CWEZDHV<)]G
PEZ^UOTD^HI7%6#010B[6?M2,/VVI'!-;8MKU!!SF:75$WZ5<^E#=VW.G1W)N5E0L
P*!7NCYF66)TWIZV\/QWS!]0<07K 1O!_1:FJ;X"3/>VL\$=!'<A-3"S?(5CEG4&\
PZAK,X /?4_8U 1@1(@UOCO<0L[]-4U@\2_/3P:&-AN<?VPU>.Y"W@-,=F<BF!AK 
PPU9ZF=/ SLTX]#5A$?>A>182]F5G+@S9;3CRBYU$=S(=^6/H; )5PED[*:WG$&_X
P+';,$R5X%H_625-X:S AX&L4HA5"-BT0E5G42"JISY.F-'"FLI+Q!@&3EQ\ZQE&N
PDU_]:!H5%<24E(O+2YY^_M<_BC@HLV0V$"\7J2#NLYAG0S ?LMI@_:6.0>$P5!UR
PP$[9O]5Q#%6VR[&#IJDD/22%+Z3T1(AXM&0L.@HACJ/KVEV6IZ>\6\U6TP+X(0?!
PBI;NLE8C)FU6OY 5:3Z]D'Y8'+ZM66K#V7.WYMIU]S<V8?3-:_'S-2FQ!3(]-O:H
PKD5,6 W#.KC:@/@_!<IPI5\K4OHKQ"P.E?E*R'N=:X>G_7M*F#WRGA7^#4@3Y,@*
PLH?U04_K1E!\8&KZH'-94,3QI!BHDNP#B<(^7[]8D<CYGW\B-OS<*"])/118;SF_
POH *,#2&8PEJC&1AO,&P;WW1/1OBP[IXM %J"V(3)P!RKH#"_6BH.?\*:75#5.F"
P%Y+#+=@+@@B>YARJAV0KJS?>ZKZO-IKT(( WR[TYMTX(7*GE/$9B57BY.Y50QK6T
P3-R'6VE>.P!:!)MMHA1Y1&&3MMX:O17Z6I[^989PNN_%]SF8?_$M&(1;:;D//;B6
PD_<AB%[&:25$7B/Y1V&N8_N\8Z;FDNCOW1N0R"FQD2R3SPD#MXTL';Q4\4[^",IC
P#LB?!M/4IDV164!HZTO 2YUK!1IKJG] WO%TXZ'>K,J!D<BIT&4"/&@=6]$!3S.,
P*0II\<? MQ/KAC=6 X=P//?@H$[Z\*#"(%OH=22FZUX#%]-Q)I4QW2K5'M"3#%'I
P[: ,2KHJ)71"%W9$9)E+WK#W ;]H1V&EW: NLEY$EL?U':U"HAJM&8#W!VY3\G^0
P[E *77/9)7LM"DV6N@>=VAA%PH280JZ*5: E/^_;I^A).%=JQ<X%+!BI/2"RY57^
P,\RX $O1=7Q@1)DP" V&XD#"G8TUI\B\5]#JC86'TU671%IE%(8@(/Z@:.U8\E?0
PZD 47*H^O$;@I?/P,[1:_K#G.T5[&D&U;;[\7>OB<L?CF=A5=L(_UP..;OH%YE</
PU7,A<PAM4=$$!5UVX=2@N' _%NXYES]]E#'=-A9"T9 $/RX6$62 (XCYCVK4M+FZ
P9-PK%U9KV5R\1GIJR,GRJF*>5];?LC0VQ9P-T^2- RA,^KJ+K( J3QJ)1:IX\_X:
P#008Z4.9N[#OY@MBN;)>C99:Y!!FS-FKB-)QCV+01^7!:*7 ]J(VA00 .< -H:??
PU4GZ,>O<A$HB9O1IOJ_?;U8IL$("&L!>"LMR*<7&\0W_+@E?%1W](].P2U^**HE;
P^K+@Y'H+&=:UZ6EMCX I)T.B:IM#*P(D2M_T[=L/"0(LU,4_+/4,X%$3MZ1H?[%Q
P.D4<'B9.;J4%<-,FWZQ#^$J8KP(W!\;$K/DOFK<S2J9HS*]=_?'QG30S#>,Y8446
PF'P=U$;W:S2S<P),P35,RB0F2Y97NUI1_^^L=V7,D;H N(&)E513;ROMG;V;,K;N
P)/4TT'=CY:1$L>N%RFNGGSC4TK)*Z:0'I@68(4=_8/:T$S@Q[I+<[>2_VS7;'_H[
P:MTOK#59&SQ*A46$X2.55"#1[3.?CV>3/#1-,R$9HUFML9W%0V%&UTV& [)L;A0T
P/@U]!:PP@]OXI, W,MTRB2I56 53.APM4T&?46&)OA$?8L#FUK1S />,7,$D(H.N
P\)_QE<NL$6QM;[[#<:$M4[]:K[.=@YU(#C94HN*L=*%X\BT=X7'"MCS[MKFW,M7B
PS&DM8O!NOB3^))]QKM08U$U:U:M:"ZVO"K0"6M[6(OUM[1Y[<^C6D>&F/A 0HE@$
P&G6## 6DOTX5.*0HYC5VJ%D;Y-/LW#%TP7ADQ;+S^O"U;"6GD3#QPRM)I>RZ7M;P
P<SX(C H,+-Z87CRI7D;C 7N2QZE6Q@[$:'2BG>0?;B45EM0L!7J+%G:?NTQ.66_(
PF60Q#;N@D)6G%V]$BB#U?EGAL\&__6\'MZ;DIXKW))8HRCA#N !U _6O\>B9_=NA
PJ'JNDV>F()?G8I!WBB;G:0^KF 6J]S.7=?H]7BED ]F#R8$-RJF>T GF/PWD;N5;
PKDN:-^KLOH2^]B'*A@-_ 1K(B',DM*@?_E8+;0I=%T=":7R++4)K^[.'EX^3"S:T
P+*A^L+CD9YR]I_!L)+;6@?VOD$%.LH:T&%?PI(IUJ-;M-M174Y4K M FQLY^+(F1
P(Z6<8M%.0?<HI";(">"Q,Y,;D<!R&Y@*K8:B=P=U$353%/=A.6_Y^Y?K%T&8N11?
P:/;2;MO\^T/%+N=7>N(MP5>%GXN'*BC6&*LOB-"2"+ 5Y'<9-+$Q UN7J^M144I^
PLLGE;:75R!5&=IYO?T184$@"Z8KA9^NB7JT@&-('HGM5.GN^$V[<@5"*8L")+M5.
PH&LB?%?*:S]?_9KY+^TD4O_.WF\M<.H.OBRH7VGU.!:3JR$0'$TL=B ]"$Z@2%WK
PL"SR*_#0[ )X8>EZ#$R(?@))K5L-R:@[B2$OV#BA-EVD_#,UQ=E$*";N!S-E\H+N
P74=9L S)S#:P]QO>XIXWZ 2QWP /E!#K]\ALI!O6C1*Q8,)J9#7IJ"57*B48\.23
PV1EF?ZJMK07<(^&,!='DWWFB0@S2F-^>I(*HO?HYV90NQ'2(QQ7#LCG23BP.EMHX
P<N\=V:9^0K<KX?-?,U#ZX?:G2F%%OK*2!^#/8)5+=ON8KXF&!RD(MB]-F:B]]V--
P\B>&DVZ>;G>1#G7]W[?VJ%J1'N!SHY\7@D##Q>?A63*0E$);?IM'1YS,EUPQ<8CS
P]822KTLBCJ< *S_"?IWGQ1B+#M+G(]KZ&0-PT=Q%WDUXYRHDR#]GY$N_>!]O8>BA
P#!K1GS#3&GFJR\E9Y!S5C9?S4^XUXG]IJQ;)EK-JM-*/ZM/9-JT-%,I*JOLC;AL/
P$HDC&J!7[\KE[RL QQ+W(SZ]_41%WQ&EUM4^3>MY9HAX6I@PPLAPSXP[;)T0!'0M
P(.P6!75L:VV_QUANE@#HU"=R20H9T!*[C(<[-T)3\^> HQL$HWHZ1G/62^8PTRW?
P89HE*KW!*+:NXD[D4/-T7+)@>A]6<NQ3/?8.T"[H+HR7#U_904KUKO)()O=S)_!R
P%7#?&W^;(BK"J-)'\ $QJ+2V&=!2^SQ467%OTVA!LA8Q0;\*-='A=&&JI/B$:V*=
P@HB'?=51H0F+*!=S34#)V"D4FFQV/=\&[J<./T'+"F7/ HZ!->Q(IP976BRQGON1
P-1]R;K_HEVY^T72=/07!>G80O('>;LUOFNC]#M9 HS-^\@ WA)'JVK=&PEQ%HI/(
PAZ"K>$,IK[_,$\U#XAIV;J$$&$\&<A@&X$T-:HXHQ_D4AI S[I5:%.$!GF/&_1^"
P&1Y0W-HG[/@]Q #^\_97!45*WBYCLUEWE=[1'EY(51U"/J+TZ3FE]KN,EIFKQ'7W
P+IJ-<OZ+DU*%1!7<5#H2%."7EIK!=9_4+"(],'+,)X^#"L_<T&-Q<@X+(73"7."7
PE5ZO QM*X,+1L-AV["YFF&^M\Y71*#@:H@X3_CK>IB%PP!+)5H<+@D( DR=C4+%@
P^)I9,0A#$)Y#LBPY1^YCHOY#3?4\0WA4M1?%^6(8;EF\[2HO/G;T#,01$H@0$V5)
PQ3DPV:A*!Z4V'P]@18('39-HBT=%JJ\,L*ZGD>_D\4/-45A5R*X08@^9YN2IC/.2
P=CN'^YACCT*>MNB'+WWX3^"C6DO$[!S;F2&R_H&+"=^31,5+Y$IEHIW.UDV624^#
PLCQDW"V9GDLM.^[(M:ZI?K_\Q8[93W5Y.ZK?(H1*\-$('XKT>/==0\AL1?%0%S1H
P1<!Z0O>#%3[5:_VE8,(;S"[FZ[QJU\VVG"3M.Z\ZVJB%X@.L:*ZX<'FA*BA.M#1V
P4[.&>YO*+.R=,NX#*QH=C$_G?E,UTC+3[Z,U1#4ZY L8,M'K-M6)6@*N=VXSE!=)
P5![?T\.+(C[1JS.;A7"-2:+7QKY!-K_UX WGIU$+W$.F=QN$S2&HWV]WH(::UGZD
P(XRKJA_B,>&G9^]OHV/.:Q_8H@KJ3 2$<.*WPWG:]6"KQ-YH% 8Q#*'$:4H,*_>N
P8O/C0CL!B,^@B7V"Z58S<]:=R3;NVA1"S<0'0$"F=6BU(3.QVOSB$SS4"EL;USPU
P&)R=K>UUZ(>$*^5'TMSKTC$5IJ!+Y4H"IE'G&0_B,0UU$2E?U0I>"%Z@/3F6HV9I
P6" CK"<_$D_G =Z:\"*6_76="3&M?,(<,+H@IR:7ZU0.Q(J++;1Y:J504TMX+!:$
PY4F91$3*,RBQ=1CEDQFBZYQ7Q:N\2@YGBI(V=G)TP3V!<(#UOE9G;*6Q>Y;O+(?&
P=7B?#QL:<S&^;A;EX?YEPL:22?JM^.?A ;\)OD#O4!BR-623LT6*\]T0^2PR65G3
PN]*8N.,]TB6+2T33J-VZ.EQ\R$!S_R@GO)76FSN.,S4A#6<?"[.).  \0Y(2J6?%
PQ=_G=:[4 7[.C ,6+!4?;N] D6-='9LYZ9 &J19CO3?Y^>">!Q5\.EFX$&O$W/S"
PX_2702* BX'2JM'.IC']^@?.@#Z-K:#E?O3<5SF4R<%I"S26F"@8S-3OP7])]-YF
P\T(,)D2#%?NB5XL?H_V<H%Z\C]V\S=J@^W!S'IDJ&NMWOPB";N'8.)T$1*9]LT\U
P<J$]Y5/;C2L'8G]CMK1)9(]4 K'O-L N+K#;1I"99N5KVN+#+UP/F5L)Z:Q*1-E$
PMQK2UF+,YWY'8SE17W:O7"A6UIKH'30PVX"3=+JW&JGC=8JY8>I\.Q;CYA;,@\C(
P<R,R9TA7$5+ALN"*Y_4(GV>/SPS<E!^IJH-CP:FI#S*<K$-$G8R B8=YQIGF-F.4
P@5=P(#IU);ATE^:\KUBPT0V*G17.94/C-!K8(-T2#R#V#HE>OK8.5$]_TN_C[50M
PMC*S3EM12#]*#61?NE%;3)$L>?)4M_JM[XC/,3# .;BO>PWA?)02W'?'8/#O!AZG
PP(.3PE5@6ZM\XX!,H7*@8TZ0\I>32:;>3,>UR+).*\=APS]#&X*OM@$S5J0B:X?A
PH3==5"Q[BI)9,ZL#_?F3HLXQ9GC_JA++SRU?O&@5Z72_CACC0R:\0XTA^*U+GG)1
PG(L6],R(W;JLJ\#W.0MQ*KTQ?UF'JU<Y]T@?S7JK@RYLC!^0_Y+Z X@716NF*BGY
PG9=;S3!+L^"QH>HB6LP!!N1[.3'@V:HPEU_RN*I91F;X/4Q@M,E#K )IH75AH8P#
P]:4F!=705])O[M_$;G P9!2X^5OJI<ZA;9N-Z8W>7>IOYL+A2*U5+Q-U.]%-&^""
P:1I<00M(3K-=]:>SZ]-J5=,[>QFCYXD2M<5Q6!AW)"[NP]W8W>?[AZ!3O?'^\T*+
P/G]]H?(M-T'D?@\5I#[1MYEE9-!TZ!) Z6@(OY0-\6Q593G@QEWO#%)4!ON&P%\)
P]"!G(#\9!EM);O[4&SPRB@1!)1E5O!KAP]NWTA%G@)I2Y]JH$AW-<5S3V? \S]I 
PJ0Y"19MZ+DF@Q*TIN/;#$GX6Q3S4 ")\ ZZN-84S6"7#N[!T39CE-)B6BL*<')J7
P?BA<6J"73+6I,H5CWB.K1_=3=1&W+S!T:"R!*!D "UV^3)=B.ASBJNH2ZWN]=SHZ
PQQ\?<Y@:(7EL!F6;(?1FT[->?&:/ B$>OKNHTI4''/^":>UL+<D/>U^J.H97EMHO
P[]5[*ZR6/TH;Z70+3:\2.U=[J34IAY/K5F#QUSM35,4Z@H_V29TNU,IP)+Y+MJ <
PZ<FB7OD-G<$802OSB&')%X!)#$F:9^TJN^X8]0NO3]1 60/C[%SG??]V:BG'UCIW
P0PL9591LT+[E*FLU_EX;AZNZ/?*^*B\8\)]ON@XMKIMF]% Z8I )9[K S;!:U@Z'
PC53_ J@;PY3SQA&IAH9*X(ZL.>&>#H AJCY1N%O1A<6E%%"6HPT!#0\P<D\]<DE0
P'B5Q<-\%5Z_P/PO0E]FF?]OY1BF>4Y%:'YK(Q=3HYZC]:P =\WI@-T/^>(JHU6R;
P<RZKS-'3WO1?XX6Y%$F)MP>H)@;Y-K#5 IAGE/??87PL*S4K*L+#:J'O(%FZ]=8N
P2S-.!)A@N4$UO3"&'\#B('=5>UC(*?@3D'[DT_/1K>1 ,)Y@=3&(@(*N,'F(^#_?
P2FS*8PJ(EM3O6*T(#W*U^J?/G=/]/J6?,0H"*05Z6S=';PI:E/5/E^X=MM*Z*A'E
P>%GIY!=M:XCU0MKX(JBJ!K5!1^GS441M6B>F/6PZ#FMK\;&H/"G^5D$Q*/?7>$5D
P"#.GP792-C7E$YR7$A;W9M(ZA6"!.I5M*UP%"^8@*M]<W;5-ZLO?<]POB(=CV:0X
P!OJ<,< J4'G))_!13;T8;,)J/0"\"%XP1V*"VI>R:\*_3=[!C$C+P"OU *ROR@:4
P[N7TDD=WTC/DZ2IQ'?'!H)EJ+>&!^PD$G?^*1O0+.7S%%AKBM)["F;U_P6+N[@RH
P4H0[##U;T9K!&L_VIX_Q'?%#3/;][+I248HC]!.5]?_T\5]&G_\(2S*7Z77EKZJ3
PA5L+.=S7O%;2SO8G&6^\X7"7W*D0'"<5X:DC-P,EVGH02+,<UHR(F6K"-V7@+"FH
PX[KM-YC]4T_[X]*)RB*CS](C ,7!9.4Q7]-PV0)R$ZS_N+<">/N3^XQ\5#I$VVTL
P_%!Z+R CN1O@!^H9)YA;-78TO[@4/?>_99.'+3<+%:7PX\DB$=IT]"MW)WBRKBD:
P"5T,4\N9LM*[S$PSTZN/PH^H[2\)F!8+Q7TFN>DE.#2\&)9T73U$.&221GIM6M$]
PK'^)\-0F]X!Q5IER7++ Y3%HJNV?P&[H4,)O!ZCZ4?4&MQB3!5V'I\S&M4KC)/IB
P>ULTDS,D_W?VS'VG=[ H;Y_9%A39N1M0 E"N](K<]FI9P_B'LN&]R:L6*!P%8Z!;
PG@[C,0S2<O."G+1!=?!V.@O*&D:I@0V^#?X194VN](.&D7R@ H:?^YKJ%PVP(7OK
P:4R[74TP2:[810$]A,@ST1G7K+8V^1$F5+5;>?%U=_B-52!.''_]L.-W#9DO2A[F
P+38O1_=8OTQ^M<=D..G>H_67509O=6V@:P'*R'.I:W1."6T)I+-PR'=*/@Z_UM5'
PYCT8MAA_E1S_&;\9 DF5HF4 I&N1/.NG3J"C393E;;+5 Z5PB#<:*>K]32\%D3G=
P)2CCL_K][C>0FW)AVT7'GJ#B_#V9854;NZ7<BA=.OR+NPNL1ME>3S7"H#W_T1]>E
PJEJI2BYE5=^JW0X)Q99[B5".R^T4 X[R.SAD1WA8[>*ORU+Y4#*J*L5@.IA\$4XF
PZ[::A+6JT+RFZ>6UT1\8G=N^YI=)<:DW%%<"(U)$%ORW=GIRUF%J[Q"H_M?IQ95T
P",J;%M"]_54MSG1Y=*GCQ\*2 '\;?VT39NO>]M= %I*195+2!VZ\JMD^#W,(G*FO
P$P4I)'D<Y\$=I#>H6ZTHLDG13RT,P7MW]!AA\A:JT+EVX8;UB\Q^4\T)>\>)$RA_
P*R QU\M=RW5<G;F?E[M.0I?_\^_1?!L]7 O+"_T")L7_9G8BF19SDQ= ^[F)O8@.
PE.!8B,8]6P:MA%Y$=DP?SQGUKBU/<WFP;]S*$K@?,Y805\8:HIAM(629 4*^/LN1
P[*5P7J5,"*$#_; ;3#V 6)Q ,)B'\_6HFR(.O&0'I=?EZJ+BD07LV#QXN7[F)K2 
P-(DY:Z2,)G/#8Q"K&>LE2 =Y\3Z.MKVF>QP,;WO9-;$I"8@&^,</;GOA[BW&(Q"3
PI81[1&P5%[E9P-VD0)8:SE)\'04MRPL*H"CO&"Y:*.D:7Z4KS4IZXW]# FXTWGC?
PP&L:8LJ2L;_\#/ X.-G*[EO\Y60QDQ\H<GW;S0%MX!G7,,@5ER"90;4GZ=JDG[\4
PUY<RJ>+##(\?5-.50.Y12=I8X<@_:#-EZ]_?AF1"BCSV-3;'"=4%ITSUT $/[05!
P:6 #-"QG6];]>'*X?6!ED5IJA*.'"EQ+U!J?/S?55]_5#H$5 CGBB1CP1N1Q?<X-
P-Y:F+4_.I#PD=-^;7C-.E*@>J\D7.0-,G&6\#T5THJF")'A*M[97^R4D78OWO,2/
PRFYD6YOW^Z!VUDDX.A<O.UIP9QLWGK]4W9 (T&>&$M!9S'=G7QAB,QS=@B]*T1:7
PEP\BCGB$? @&]%D>(U4R>=X0%74\.;A<1F1CY'3>O*!/09Q$T[P.%9@I\48R<'O)
P^ 0&G*E0R_*O2 &79,H]"HN,&Y%*,]XC* M'>&V3\+S>;WB#2P.05X$Q=2 N#7C3
P)Q(Q+!9X+$5@"S^M(1)CT,3>"#.\]]X;J9AUR8FVP!9JF&;+1X.S#C-D>R&QJGLC
P;UQ&D3YP^F]?%UHA?1$Y$";QF%(EV\ "B=<$5(TWV8VM:V'WX;.$,U<Q0153FFY!
PD\@1#30(D8)7C@ FZ;MCX(E)CE[L+I3?;6$AA LQ1K*5T;#K=P%@KY5* ]-*559H
PX0HYCX)=K$TUX,HQ,ND^T*EUV05'ZDS)V/WO9F$TN::T.+5=);[R^!?)QRP:(UU+
PO?G!$W"U]6HQMG$MRH$(AP^^W@=(.%$C;U6G?Y:YVFI>^Q&#6I[^V[JORJ6>UR_9
P(RPB[OD[A=#&X&8\'7GNW/CJ$I]'JEJQ:=IC.L*I;?4G=1/,RWQ!\; ,Y(:0M-65
P!_5BO:0\'0ABYCCY9+9GYEQ_;R0&0VN*G^U:HDL-:VNJ2RDI84NUN]\DQH#$N%?>
PBH,[^"]*F>?=DS8>=$*1@#678+%MH2+FBLORN6(]'TI"1>I40FCC>+">_/QD\\RZ
P\<."0H@-HJEH_<<9S8Y[7K#M_9D0GI=*7==QX<'P+$ZM9C\E]'@)?5C%2N+XE4K5
P<DQ%-]U32%_56L!FDL@#UH<2J>AM*4:<2PP\6_V3.[J4@T$<*;>79R6G 2\_89;_
P)NHR$3X^><[TB J+A7PJ?A;NMI?!D,]'MRK/<TW09VXL@NK7HV%2;>H36!G*V>U^
P /0W(E>8H'LQS#-B!.@N))?@Q?VR'__^T9ET7A"NS74&CBC@X-I?EOE, YG]9?_Y
P6I&3<9AL>57,&L:GNDOCC= !R&@7L)W^\ 6H#-UE>%N7FC@FAN-^L T1L?<U;_3X
PDT37>>P>))8+EW=EF;9WY]CKP']#4.W=^/UGL7GO8.>P4UW/A!P:9PX)AV$%L1K&
PG87FU9\R0E#C7''2[$*<;2F>)7RZB$0\>8F\X4M.1B4SZ,'@M"TXOC02\?%U[.7:
P9*0JP]7Z"RDK+MCW^,3U7C2UIN3>"C1^Z>S,25;;\?-RNK/5#3!O/ATNA@__$TX(
P%N[6&K>8V>$IWYH4T.+F9X2][TTBT-8OH.ND[I*MXV^YULM'NO7W7"DE4PA*X]W>
PMI366L>%;MK6]"A=:$9A!3'^Q<&\&4/++DI0!Y&?<V+&Z:Q/?8_ZFMP;PX D4QX:
P>CS<_\85[5#QZ&FPEZ@R#380,4KE(9#.:8YV8]H!>;9'[#KTQ"O!>'?G%QT-M[31
P'7C/4TI!'5H.?TUBANK^7PU<;RGP$ ?M"I=YU=9$\>=>Z6B02$Y^!IA+V\1D9]YZ
P<4$ ]V6_407XHQ*PQK$B%ZW%)GFC&)L-)2UG';/=KO<!3^[8%%B.CPJN1VI=!G6U
PG3<. =7: [S_ K=RYJ7?-"QCLUN.R@V!K!&6+!FJR;C^ \][7-Q8SQTSM%MKXM.!
PJ?3-J8^Z&3T,L!'2 5M[T22OVQ83/*HRW*](0:4?XU+ 2'Z U^.&>:2EV2UW'9W&
PO2EU"1 8ASS:EUC\'A=W"3Q[WT2C.QLN@-(\:I"T?%;&8A:4/5<SS0_6=!N>1E1!
P55%A1^C6I2ZX?P& Y&4'QN&V961KQT8!5P_\5-99%!^,:%X5;)@V6Q%8\NU)8<NK
PF<F$A"ET@X:_V6V3T_<DY*U[;G8@>O<H1G#3)<NFESGV Y4^LX/#P\AOC6(U5TVO
P/Y&L5Z?NF7!F^?I?$(^"::',@/P#-N*RHSR:.YQH$_\[<?5BYT)$B^*.%$=$[7-<
P#F 94JHRMBI%]Y6!(N!M,:O/;U^8LOK Q\FMG_VKKP?Z@:SJ.WN4WUV\.[YK3<E*
P'F=_(/Q7Y92^7,+V<Z0Z;MA,\H>=(IL< $JF-+TFDM!8!7L?CG(@>9Y',F\FX-T6
P+3,/AV\P?>/\:%_]I>K R1&)2HFX#B;JFP= <WM-.)\4.PW=0:(B0L517V^HD#KX
PV%D\W>"=8#K/SV(Q?QXW!33MU;#3=NF)24XRZ54:)F3<8E7J0YP2;>2QS:<'2]#]
P"U!5<P;L1JE!QSS<6QMK1GAA0F)9#?7+3*D^B#;_JD_O/] #O!;-E#$>!Y5#YLVI
P*;62'$!('<S6.\Q%AJF($2< FC]@"W_W'SQA(]=ZUW, D-W,OA3-.>_JT(:"IF*U
P-"7-BQ0I=HW6!2'$E\$'#N<#7SF=_RS04&;IK8'CACLR$8L-*PDF#=$;*^6K3]KF
P[/O(/UA4\D4%;9DTA0@>5%H*7KT%I-_!1>RT$ 118TIQ/(DL"LXL_*32*TF85K*/
PG@Y@D292#!L4C>*U.LPY#-J3]J!/1%Q8]I;XQU._\Z/(,_CT71--/?E-PW) XV7 
PR;&V&2-NO*T:[]/>(C+KZ4%]FR ,$W>_X/K9Z8SI =N1?$UW:1Z-C$"R2QW&6P8%
PS[Q;\[(>Q 8@;D9A'U5F4,!/9GR$538P7TS66Q^J$$9=E/3*5X1QN4J'9QG>\7*8
PA(:J_, '6@'>LD T"$=OT33J%E?)PC3X$(\^L*@?+'GLL%M532K(+P5,4RJKWG,M
PJP7J<J6]5J\OP[\0P$!$Q_I/Q7B^SBD]CO-5IJ,**RC_7LG++Z:9-"\9FI,2&G_1
PPKZ@=GQ1<ZDD"6T=DV0U?:E[(ZM9\^D-A'?.RAYP]O">Q79+H9(5VAYEIY##<1@5
P^S1FU,&MX;_B:!.A%)@9>T?[:?"TM=XL;U ]9SQ@W%YV.(F3!#3<3N7?;J3OW9]Q
P7NCZ MOF[;;%5CXUBZ?,.5!<5ZB->H&+6A 8PTG_*6(Z%QGG\;N"-2M4YL)"MI*!
P_7H37KFE6"17I(&%_I%5+_0C/7>&&$4C; 2^SQ^8E^4Q\<*RJO'K.BNPM?EC_Q8A
P.EF!)XXIAR#/_5IL)T]. 7KN=(I85>:L7Y4QN$WBZ&_0_A7_$D'ZI6SDM1BNZ<,;
P"]DI@9]XZSEV2Q@KQ$ZR3G$V$E?IQL=Q$V] CPXP-%*[8A(3:P/>QU4KO&C9A4D2
PH:DW<Z-9M(TF\,Q(!=B_"03P%8QYT/]/[+OIQRS^DGC_M<)6RI<C@6!Z!WG]W.7(
PN^O4ND->V46]A:58X,OMHY#"$4T'O2D-2T4NGV%'8BGNJ)5!ZGE<L+]&/4KN:K!R
PXTEM^O(>2O*0&_L@-^#]WX]@((M(+IT>+$F\DS'P&!H_X*I"G]H\C&G\L0%HBGD#
PCOH#]3BY86AU03/OO>&>?S\4_?J/%\W+,R 5THM4Z3UDSH4[MSQDM_QX. $'$X9L
PNS\+3W8#>#&ZRZW_RM>9KLO9@@$M>):W-C0.ULA@TT9,;% F/_?QA((:K#N>-&K=
P?( 6 ,8$H&0LFPTMB@G&,YEEKI^(\4>(I&G1*PG(N#"!U%TF7CN1SA#*(=Z<"6Y7
PDT+.!]K=J(G0#V+%44C ,21,;A5:[,!(= )=M$6N P,^O@P4T9 BY;K$'7H^?/M!
PU9%S*$HP2QXSZV-GL>$5%N5>BF^]-<QY6HNL U[#/ORXZN50&4ST4A?PO(E1Z,D_
P7,<KLP$GK^U1EA# 'Y.$DJ,<$3Y",U-$XQGTW/^J.ZI*JAB^\L6VL/W[7,D;=B/$
PKD4^U4C$6T&E^[QU$1BT=TH[;1)@<5'C0TO0XX$$"'L5 9G;YV4T%]27RV,?6Q=Y
P4*[9Y'<^+UT#PX$<J<#:> B_@OW-5SWF)1'*]?9&:W#*PJ.]N[83B"DEV+-DG<=K
P(6\3% -SLHQ%HVNLG<,!X#Q2Q,UM[=&[I-.)Y<HEDAJIQ":&? ";22N[4*;CQ8=T
P(DS!F%#9*O[G7W!O/M,YD\D"3[\,T]_^@WHQ39XR@:[3]<8TW=>CJ>"2G=EA\$E0
PB6RE5E4FS_RX/W\/,B=UBMVK<'3RPBW$M:VXPDNV+6(&X[>KH0;5#R,OHZJ)T5EO
P\U/?EWOP2V?1IZNQ6AYY,#(@F-E-%YD9PK^^T9QSGP!T5Q3N!M=)@("E$85 ^4T/
P2! 90%)S!T]DU0QNLT,X/A 96)Y 3$;'[1?PK^??]&1MWE';3<TUJE26;HKEQD  
PQABV'!_CO<4V>-BM ]E11-;+8?FEV*9KG2@[73WXYA"MA!+[J3B,!^P$D7\JYR88
PX@+U.Q0GUF+1LM>HBDIVW"1WJ',[AEF6R?LPA?V%@K\)G3FNK,"5@D E!"MQP>*O
P9][I-,/IT_PT;_ \AN4OSF7C '"#>/&3!$ .B"6A%DUR:P'$;8'H<?)L<"-.$HJK
PR0T<0EMZD="%&=6:P"M&!&^__K,QV9LH0\#^.,Y7IO$)<0:0OFI$8.LC$>@6HNU'
P$U+/:%'9[W10F(+=OS1(9AR#89690M=:QHN^L&ZUV&ZZ*/@3E[\35U+YFJ!9()PV
PG^=GF8F$>L'$=;)#S_ ]$A9 BN_>U?V**;75$%0$MAXK7G.XY[,JG)H@JJ7K5F A
PYMOE_YX]WZ\;: 5);6(GQ@:?6Q(?4^QZM@N_';A0@&31O2NI1Y$U'- YQ.#XUY+2
PJ PW2=9]])2FCJDO[A!Y(RTKTRI,["']KA127^[-P"<Y:Z$K6X2G%7=41'0<=K8$
P9/M9<K;IYSA%=TEJFO9E&1BIFX1C2/<))TA&CB^W\/2V&"G960:Y)F:G_Y+#API2
P.D;ZE%QW[78#D3=UHJQ2@PX:@39BQB+TI*N->AL6@T+$7#Y)5T=JB*L& %2GZ1.(
P\(BJAWR">"ME*CS"48P93F9X"P%'?W[FE^"4C OK>B^CN=MI2=SR^2?H[@0*0>DF
P(&L@U$?-J1RKU1=5DH27KQEP_/OPZUSPG!5([>MPMU:J,*$AS6":H++<:ZO"B5%0
P=[CWK?@E43K/U=[TX.*"1:XB-PT0X+R8[[,.WOO6V_G3G.-[>IV-T<L<%=)R@BK$
P3GLK$GZ9-^GQ/!6!&H\R6^KA2 K-NQVD;?X >W48VT^EFS!7B4^V]1]]C)CT??PA
P.]A6 D")T7^%W5#J_T?$+A#AUB;]0J^S[LJO$%D:Y^RTUW7Z0$!F/@0"=V)PNQK\
P@3N=]'6E(+::DF-JY=A,PE)2LKCVMW^#BQ?^ ?7_+RW<4P'^^>-K6$-1+TM>0\5M
P6K$QL?0CO;B+$ 7J<R=;Y$((\X%_!L:>-!T1+K(J=7,44IB4:CI_2D189\$?U +N
P()C@(;!U4*$06!TW98.B05LR;W%N40E=F@^(M;I?-[8B<@0G,"I=L48J4CW_*V$1
PC7+VZ!24H?JXRD_$9.7X<!B#/1X[=>-.C4H^T],MTE_4XFUK\<L09AQ5$2L6/"OK
PBI?9II9 #KF& $R?CZGQVB:E\ K&6Q"B'8')%Q-[MU/.D(XM*P:,RSTPI$/T/7AP
PD:)9S0A;4IE7WPK B<W=A@:@_4FI&$]7CR8PQ4G.4Z_KB$X_P"P55H7(!T$4;^6]
PSA#()GL.Z\Q#GME]W9$DBPY\#?&TUM%W=D)I//VUX[2>A;*>!.QYF.6$4:C='6C,
PQPW&$KMF(DPV@;WX+D797G30+E]ZN:\@JOG_WP<.XW-AP4K%B:H$8&+K46<T#PLF
P"3Q7!CU'^S5"WS#)OA>C^W+<VY9!Y+DPU"5?VU#:V(]T0HCE@ Y6=+'#[O=.B!C1
P/H\/\S&=A$]THFX$*QR%92A<E'S4[P#A6H*BQGFO_;B^8,8VCYSB%0V3$EUZE?9H
P"W*0T0Q*SVD1><,2?B$34_VF/2ZHVA=!GPPA7 OL*2.%I3%I*4 /K,L4UPD?_2UD
PW20KL>]X\#V.[#CKW*#7FKA_(A\%#K[]I6KK8M@FD-$/? 40FD=\Q*7V<'T&SF65
PG2>R. _OYF,#V[=V6I1:*E:]]8!AXA&3Q\V9\6,PA>80OCQTKJ;:%P#K38O9=X@L
PI!2,W9^Z05M+Z!4Q)&\VP\L'J[P"K59$/FA1:- CA\+:J+RDL[KCV2-@N5VE<VH0
P?>0V#T7WJ541+ 104&>Q>JZN,U8H=P@J]E.B;N5+E-X!&[),U@SNWN@LV^VX"-&@
P<OY*<KO8+?76M"A(&N#G,(+I6QVDCBZ4$MK(IP>F+HO442^836)EU@UTB_[F:],-
P,^(@$ BUT7 "CA679^YP4<#:#S75 @W*?ED3>WO9C:KJF;$J\8<AB:BGD79%?G5,
P<^JEP*RV1GFP#W(8#$E2BN;J/YZ'E'NPNL+R>X;:7K</,"]G!?.5]=;7-A8DQ:%W
P"_0/&<BJM5T749*KP?2);_YI6 Q!6A([MZX@-O%@<W$=VAHGOHA<E1%)K5L#S:+T
P2E%:ZA#(R/2,C8?E)RH6&.9:![$\7-]I=AD?Z1T&MQ=^OGG"RD9\K;FQ,4\,ZCLY
P',VW7>&P%EF;D9ZA 6HH>_1ZLIL_D:^VJZ*H2'*:R.1_MN\=Z(&Z=9PG1'%5@HU@
PSNM$=]4M?W?LY9+.VX&?-SA0_K.Y?MH0+"5O.CB^VVLAXI- R$*8?.7/WC :@?)M
P[%TP8"3HL&R:[]B1]DGR:=L@BZ_X;HPI$:-]@H'?^.E<DN15U<+A.%CUE^I&M._?
PE1=.HRZM+?/;ZNEPMT,9CT5---?$]'(C^X4]"J0FP4ZDT]#^$4@Q%2P2HBJH^R(C
P5';VJPF(H73T01IU>;6NQZU7U&:8*07\S#@?9AAZHK3A?"L"^QK9"#<G1FS:<WV\
P:D&K5-+7Q^#AB8^BZZ7A3 ]/KD933BB_3D624GC.EA-NH-VG;;5!YV:Q7"SB 7ZO
P\E4<&__L?L]VU[L6OJ'\K4/)B;Q84Z'9,_/8?U4\A$>=1B**PAJ-Q-4%:X5F2C9C
PL5U]M?%Y1O.:?:G>Y&# EGEID%U.EMW@L*0N3^XAH*9/BUEP_BU3;JND735D[MV;
P5EQYQL86YZ_4H03GW6P@&15J2>T1*[ <ZL$=I\K<$QT"8:]Z<]-U\%. H3\'3%L]
P;,2_IK2K3CT<V.?:SU7Y:;)@;^\Y *P6D&A:"FV=BT?18A,^@1]%*'M^3H64.MI"
PI7=QR$:UKHO6N&6+!WFFJH'L.BZC'LY,,?^BJS,HH!A-'IH+8R[%39V<T<FZD@;,
PZ3,76WD.$([O/TE.9ML<#5P9C4NX-'Z,X =$;#]>J?R8>NS$6XF-36"VK=&9#_0/
POK\(?5V$KD1[5 )7=?67\GE1N[/1/<;&V6& ]HP <& OX^C%A!4./N)0_VC9UXVG
P1G[8>GWI=!N)1VT!.F;R=+3[^YM]YT*0,2HAS@1+U^)W8>F:/SA1ATS$S:&E*Y@5
P<X6BY^P?FEC10LJ<*4R0V,8NP19\ZF-H;XFV2=&H:.>_.I8(J:AS-D)0G)$]:C-&
P?(B@0*:Z8M\XUEVS5''P';Y]"\#GP8='$P%SOW\<^^P/Q (V!]I2*19S1QPT-G#?
PI9UY$04*$72H2@LS/;% K?>BP'EM0!=DNYZH57<!6QRL8(S]#\5)W^#*?XR9L-L?
P>$K5&F39QKOL10P9//0,M8O"$'=*I/[WHX"3:3A#1-"S#)65?C'VM*6&['&G1GRS
P$H>'KE?Q=?+T. QOM5Q7<22))6LK;6.VFY-V?#A[E4FU:[RO\!3SQ5V#AJ(7C%&Z
PK<JRZQ<LOFBPSMH(]3E_("+#>OU#27XHG$,D6TZ'K:;3VFQ4TQH?'BW@H()@LT=&
P:]$Q8!&,S>%R.J40V\1[R)>EK;HEC>7=J8*#,1IJ%TCACJ'/]_C4)^$?>,_5D$,J
PP]- R0(2Z>:0?G@B5@K4>HP4(6UQ9.V]25YI -A^B$^R=HYQ]>]PCJRX)JQ/+;R$
PE@^&W(WA_$EF8>%(EY&S@'^-_JB/#&WL!"5PJSUEWE'-MN!'</3LH\Q5T0MCE&#7
PU*>UJB:!)+%FKA)]B*2>?O#E4WG:3_)GLE&@H9^S'=EW%-45]GG$."[JMCBGV%IK
PT>WGE$"K-)#HK2=E<=O?:&7Q 121%EWLQZS4+I(C]]:AG8U\#/ENKY7]\+#R[QSR
P2?"_0C[M<@I>61D2O^/X()TEZ$Q3@S5(,&PA&WFX_JN2+E[XN2$HNQ8M0WVD-O66
P;KU73^2-/C8&R5D.\A#;&[,,@Q0^\^=V.N)"\>G3P^MJ4-P45R_E:'N>N U.^&*>
P@'"8<]HBHYO/."N'8KUMWSZXQ2[%<%U&7K>?I+3#-PHX[H**3V7,:03Y$&YX)J&J
PZ4UM'%;O&. #\=N)T$7=686E>YC57KY/?3&K?;K'6XHQ'T%'!-0@5]]IRH7P:2@F
P>)CTBR;@K@@%AB[BS^D0UUC<6 0DM$@CLQ^C+[]V]9#"HT72S1HM$:48RE800":Q
P$9J/K9=4Z-;Z3I"6O^](NL+SA=!O-HP$[Z<6S8)$9[OZ>?=%TX">\0NB-^U9F9DK
P*U@]C0Y&@%40(U5,FX34@=I>:;<9RTAE?T!&H$)XW_$>MME'1ND#HLJ.Z=/,.5W/
P1P)<V-HHKB5I=0H65GV,*P^W!M)AKX[MN+U!? H O4%&+W]X.L"@]D\T. (,J;E%
P8QAY,VH7%]"7)>.\C;*+'X0S#*Y!:-D!.D$&GV?UE?"3K@X8R<$*J.6VW7#<VDD&
P]+>1+S9QMV36RYM91*]B"G7/K[6@_-F<O@=]ESB>6Q9\"A3K9#K0:]"#9^-=!3A0
PFY0=U^*MG?XQO_A6)A_#%K IWK]S0&@A<R1&T&6F;U^2#?;9)Q-$!OO-YG#IX)5D
PY\??W$%0L'J,;F3EW8&)$ZCQYLI W3:6Q_8JVA@F:8UBA:/:#:H6.IJ:%:%;Q\7I
P((!Q .UC="^:]6MEC5UF#(X1Y I6B^5:L?/O1N##)MYVGK^,E*BY'DE2$=?(HPNF
P#5A^,]?SP\YA+2K_3EL]''F"Y*WKMID@T?UWPL\!#GZV-0^\M:#<1NY 3_35+Y0'
P4##&(V>IMQ[ QR&-#A/^#*"%*9G$(Q#XT1O673(5C?131A>+'BF*B! ,?3G&W6N<
PY'U@25_'M+@PR8-7OZ7F9XG.K,5 P_UIKCQA, #ZL[U#Z#\.;?FB2D1DHTLNTM_O
PT=\DQPX53\S>D:51/$=K^U)[8:5>_K^0MB%^*)D]I,!EO &>B @%Q]8)NDV0BQ=5
P!I45OF/^%?&(M+/U(7_X[GSWMQL6PQ:VGVK"R[T41\@&C,AH*Q9.#*)&9"W^9#9C
PS_[H9@YGG&%H6?FZ;2VFL936W.X0:GA6(Z3_U-];&@K,S$@A.9B=?T(.T]F).C/+
PZ(T@ZJ8.@+F)U\>S=5!=7S1/DUM3&:>C98IO[M-A188K(2E@AZXAA-5 6"^Q\?0I
P@KF34!JM/Z B2 C-3Q%)BG-I$PR0.L9>-&: ZF@N6E!#V;D&N4Z$C"UXOJ^KS3)S
P6]R*<@+SX;QX$Q*%%+B8'XC[*IM61QT<VG?OKJBGL"=@'(U/%2A>1I"W+!GSW&<G
P&D,M<L;8_;FE)]Q7TB5O>2!4:^1D07\M@\Y/L<G7 P^BBUP*^<R\V$1@,MV]]<=C
P:%(U;^"(LE_G,S"!/8>0P>["'+)<Y%"8)T5Z1#= GB=\=*#Y.,0),WC8OC8->G&$
PX+98P*^O0%VAP):WQ/Y&FB],D)B/'HNH?8?,A;"!_>%,W6')]^+=8WRWJVQ98(7'
P2UU799;%<L7J9B?_MB,ROK7WO##1:]@[N] R\@<_&CCQ:TSX7^\L]MZV2*GR3H1M
P*J)W>GQ#^J@7[^AJ!:_?EY5*U&DE[PJ.Z8,G6GP;>Q/=-^4;DSF<-C#1]T&IA<>+
P@P0HN5P$%< $&!%<))?*L^L5==EJG3>4;SNUS.:3#:MLKE8_J^'SIQRAUNWD$3:/
PG*A3PG\S+;AM(VD^T6Z^7WF9O:HJ#"%:1SQ_R'W*<KKEV.;7N'U(-'C[[(FU=JT;
PHG5_&5<Y:Q*4#RK^P_/WZDO)((EJK\-/^ 5B"E7V 6^?."-:&J57A6O+O(*5)@S'
PD5V(;?[2+E'<2J\.,) =M55\_AFCH).:#O"*C1QZ[PS)D8UP'5E+^-E181M86*@C
P)8U2UNOW2)ADV;@N/>%ZLI\Y#$.XH$I T0Y (L6G.QKW 9>_9DK3'A_]PG1T=^9&
P/W8S?TB)H,:6MY'/C=_R7>23CV1JJ;0&4TQJ*?T\33U(\7RQ7[[0\*((!V%R!=O%
P>;6(:7XQJAT^AWLV70B-R]3Z!ZK@S=WL</#\VS:G7]^^..J?IL>D5)\<18;%<DF3
P+P<=HR/I L/[><&M!1J[7,N#>)'1!_0/Q'N2INA72[D^V^FUR<R$VA_$BSJBOZ8K
PAF$$!OB8L)WZ=Y- 3)PAN7XUZ#2\8R-+9H+Z]BNPGC3"&7S3V:^W,D/=_";:.9R\
P&R:^9<+_%N)Q;/]3"#HW]XZ.:(#$*'M6ZZH(6S:Q$+O:&7Y^99R]3_P ^ZV87K9?
P=52Z9V+E3$G6W/O=<]@AKQ=OG#T\TU0=ZX_WB9JJ'K'.P3G#$/P@N6O@G# Y":/<
PH*Y1T4_>KGX/#=+T9C6SU]S%'(38["T/7&2]0IR*L=F,.WC#I%POH3X%(*?AD9I9
P:&81OO9*'40PD,IWP"V<4I(RGP_ZRG"MDU9C.;(P=>C%$(+ 6L]T2OBXN$X*:7S\
P*\^T51&1JKQ H0FECUR5R<T1-]C?2O!\2C F!L5@MTVH+2;&[TE"CNP/L4QGK*>_
PRM;MI2_7$A,2\R#5@47I][HN!%@^^G]FEDWH:>P=6+:)-2BEFUZ,/4KS,K&A=T'X
PHKIZ)F"(<_PC&WBG3CYW^WKFX1)(]8N,X]K5*'H]597!P3P?TQ)0<N0JDMRL1_-9
P#)V>X?CD9_X=U'QC4^>GT<1 D$^DY<3&%)W#<ZP<="T$]ZEI\-F4;'W\!2_FV2I[
P(\26XD-M-AZC*A(N1X,027+.$]#?O*3E**N^7CG3#$$1<[NOW^A](]':?<-GE)&?
P;FC>\N<$#;7R:#&2VVX81S]712SZ16;EVM9)*7-G,#6-A?>0B@(QV6UG@ R9RAM5
PSNX*T3U\/R4#$""5EB?3MQF'%,@(X>Q*6E4J*+2G+YB/P-^J5A8QND<9MD!LHGU[
P6RW3Q#(L8X$.A(7#)J[!/X QJC^"IG3T0M&@: (@+9O00;('$!#%: \^R)ZQE#AO
PM;9LZD/0BDG'6O<RQ:[DO,%K_&#70R['"H< )?>23^E8=8RL,4$J7<4;5C54FW'2
P1VV>7=JUU.>G1J,2+&M(K8J#DC9:Y*M',#9S"U-VHD\P%'11N:%2\X]+P?HY00>U
P/?VHWKLOSFYTG\I,OMO>BM2%S/5U<OVV$"X?RDE4/(;)?;'Q, '9/WRNG\L@8?2'
PE"S>(I6"@9*%9^--1 L0=>?79;8B$ETW0B4KT.:,1C=G'?.H"C0I&EA.U/-<JUM6
P1^\(]0<N_C6QX H(I"CQ 512Q,# G,>BY<8)<0V7\LHZBZ6M"(4:"(7;"JUCE=2#
PJJCV8"_/!O+>;I6#$@3ME.G:L\G1YKA3#)TP77OH1#7Y,8M"##Q-#R].71XU\6HU
P9WPNJ J8,!X/G))Y2M%,<V%Q=Z0QI.9VK_"P([4F[*^8-#BQ_)SN=L682U"@T/(/
P5KLHW=L.E$Y[WKDL0X@V"!)=F6SXMV"'V=5<W"JFF1B/4J6$PQDS:^&5Q@NO@_#P
PD>/!^>$0\5;VIM?;:PS>O%+B:%,4Z&(7?N4T(D@\SK[.Q+E8%+=W).BU;+NGW?XS
PWW(L=I*9+=N2_'PY-&E[7LCAYN3Y6M7<Z>ZLQH6%0&OLI</N<CJ2N!V3^.7T# ^A
P;1'V3/[CH#TJKIJ[EC_!JXYU'T#[(T3C3@-#;G,P).Z.&*-N8N/-,'O^P4KC4)/9
PP$<R-HY_".V-I$U(!#IG??79H=Y7ZXW1NWW^LTL:G"682*:PI[4N*4!6ZR<H!23J
PQKT8V&AGN]W$GKP=YFM)R91F1TLU@XXT$[L.5:5\*75*9X(^\-H;0ZEA":M"!65P
P!3,QF"^B\^ )^-@\V <NR1%OAQ+8]0;M^+3"3"\VR,::V,N$4QA :(&&>C! :YQ&
P8"09C*O9_];>S15^R%^B[HA1[N9QK#.GI9N"O+TNX0?XS<;\6#&7!.2'EFQ"&&>/
P+!6>F2]<^3BWX5;DN3_?GUKM?P'"_VJ'X?*17@AA!8.P ?&6C4QMO-EW%VX8H(R,
P<!Q$PY[ZA+&$&C>5-(1(66C\%/X,><"&<-K@KPJ0Z?04!:NB"XGRDJP,FS)7R%/C
P\^//HAI.=59]RZ+"K<9)_D>%08)43+S#VA!X_:TY_E-6L,%$JPGT-PW",7@-;434
P?K/,+;0NPT8E9!1B?<)\V2K@[F]*8N],/@8RT.47L>L79H\DWT-9M]\$T+U50I0P
P8^2'8/)Q:2P4\0:SR<XVU9/1 _FLS_AT=?M5,TMPD_53(3#Y^-"VH=KH^F^8,'+D
P^H^^_'KOWOA7V($^F>T-H\3E<0 U<5VDK_RN:T3HALFX_+F<;X2F_Q-0Q8 K@&0&
P%2*NRA,J9APFNC6E3G>0#/<]BU&!AM]$MD]#*2QW8J4>C7"5J1^FCRK'UH/[(KOK
P"JM'B_W>R<>@YU?4Q.S(#$%)O'#=^10)Y. -;>379_\R"VQ:;'W;QUK72(XU@[%0
P)^(%9N$ZA\.6;@A&!R X 5:FI=^DF\<2><KA,QEPI<>%V6"("5SD3L;)][J5(>-I
P;=?$NCP=>^8)SM^RV-.R\:>8"K%Z7L<U8=B&B9"KV@]*FJOUOCST8&RT?<M1$%W<
P$N]6I?,.VR*W>D1?-&'#>"0=4\+ X\=_MT3Q*&$PN2P.23&8G!T@"5V2^@@3H5W5
PFY7OJ.POL;6, +;S.SQ_+=Y3_K.QM?EK2:[D"5-;K:8 G\^F<;(_AGP[8!LTVLW-
PC1J<VJHZ<&< ;. #GK>R$M1J6Q"DY8LQ 7/JK_JKEPB@\L@J:A]7]-"L7H"5#(>Y
P!=Y>"5Q]@H@"UO_HO+O!=)W[[;;[T>HWP55N_+ @^/Q_N9A*Q: [\CV./!C#4$FZ
P>92+W9#DG ,M\@J8,M?C2Q#BVD% 9HKS>?AU(F.YQ0_*$U1?7%:$S_8_()R4)<0%
P2="W6Z^N2E1L2Y.@3@ ^43W1-?)\7R2-TNLRIAQS2X@#\\B/)P>((H/V &MG]''\
P'D<I[2C+65([7P]YKLS9; _QCQJ4!1(:GY\<D/4M5[JH_M._>M/T$@:I+<2UA99Q
P8!;%8J4-J?8>-<[E,\*-/@C+]=L:=*NCC3K]I*M+^B6O#^Z/#EDNU(WWI.4 2:<Z
PJ4<GBBLB);)+/4L\/(3[#HGZQ^(FA\<[F!ZA4  U($5R3.9,LMK0WJAN19AKI8NK
P-V[('.6(Z&_"BPX2IXSVM+9^6%]=WMWH2A2D,I(JWD+D'Y"QG(R/O>7T.(;6U:1 
PJIO!(SN;[H["M"^Z-'](X4Q:%*53ME\+I@?*LA(R/.6XH4V!IF-V$'. P\^D%OLG
P3,-D"D4&N"MC>A%6?LPOZGO"F _*ZATU&NX>5AR??@F4=S\?.%UJ8I._MK4E06P6
PD_P#J_ZM'(WO)H8[E>WZ2I&-!HGQN*UME2O,I_KPN;EMWT/W!%PU[W]F,\N@*VJ=
P&)Y:<UM)HS2!3HS(1:BGG>0B &>>UB]UZJMO\C25?AK#OFQ$<\%'0A1RA+!J0U<>
PUN :?<8N;KC]Z%;%Z$G>U3'W%-VP89CJQ14GB2-]^?I0)A>&L9RYD::8P#489D':
P\D^8 =E(?/*CG9CM>I<G0ZI-32^J&P@VD!^CZB(3I-FD"6#GFNUI%@ZBK/.+( M+
PUAOKRYL/;.SE\[88-X58&M#+ H5'EFA(^[(L]%G&,>W48P5Y+-@D7W['HH8JA!G4
P>G$R:6<IX&UGV=/O"=F0(%X=KGE)$$&=P/=M5]<L7_]_VF, T0\9+C($25=X*JDY
PR(YR1[A:(D2%/D;FHR'@JJ^OI'/:KEUV>#ZS13C[2[QG-\J="^6#ZV\L$_B"L9#.
PP:^A_'I<?W3 D>5R9)1]YS\1R6'?4LUL D-D,O8)%?C(2")H:QM>2*.F/XO8%%I*
PPOQ7->3Z?1)TF+1KK%M0N[^9/L5^H.T@L0)J0*NRKUE\\R$#5)FV+AH&)ICVK_,5
PH*!&$DWW##K87+;9!'7M>6A/OT#Y'P_/Q7VXN[%"XT" O;ANL:DIL^/FT60P3JST
PM[?5VVECTX+(6^K]1]UC. /,;AM5[>MTIF:5Z:&0*B6^U]7>1/AS0% $1>Q=_"Y6
P,C!6#QL]^S]2Y2C3:UF8!>!MO^GL,.&=[T%=.U<>"<.01@%<A3AM -.D1@<?RSH8
P^0O>4G \IIWGH6U'I<UU1%9^=]7YM2#81.I[SC@L9WWU@FQ5CX_,LN=24S@^&]-1
P>2Y$OJP\07U>D9Q]"B+A6:+0RUZQ\%=]2490*$_O<S?\A*@P9X='Z%V^:8=)HASE
PN=H6+(6*7!W5?!] O^++)%[7'LJ,'!Z+@[BA#17'A7>CM*KGKV8!?7!E96LA)2S?
P;-9+AH[[:%]?,-DWY.5Z@VI>%UX(_^<]-<I;8O_L@3?(8[!3]%^D&Q.PMG=5A2&^
P=.'+W;J>?"N;)+[7W,\"+U+>E31:RHSDB"Q"UKBFWF%OU4V;/P8&M[QJLUHO<QRP
P@ X+RFTAX G&]CVW)XPG\.=PNR&#V@IIR:NM(,,F3T/GK";\T4'W] *0PGV\\J>0
P> 3O*@#M])@?N6YM8 5;T\TN_HORFC;2A/Q#ZP[V_F7^%G\<Y;KTIQ1J5X<0WD!Z
PO.1N,<<6Y0Y&>%HMA?,OD"^+$C! AV&N&O\#R4N)P[54!+T 'OJJV6-K98Z,^:)>
PM)G\ ';--N_C"(%?6IW6.6539/=XV)F%%)FM@?M[LQ9#E $%V3\YRBPR#ZFCA'-[
PP_89C'1F0';P\W #$A).1K>(;:U3U$;4[ZZK5NHCI04IS56M<;U^R%IQB[ZH9?RZ
P<]$@C7I"";/>YSMQJ'OSA:;LP]F*WZO<"9D8!+\;8%$[^1BB^4/W84Q4/#(M;VER
P,ZQIGQ:<_P/+!4Z$*6DM>HD)@N0HBH0B!99X P:WT5QI]'5'<Q'<4LE O'+"0UO 
PUXI^]V 8A):T$L%#S."9'7HDMG, -,(,M;5*X]C'HZ;Y&,.YJ^SY!HWZX_$"8W.Z
PXDGN7J(TH_0IPO]1^'7%\8J0XEY@H*5V>V(!\^NX),M#4JV^]?PT85X/3J9C*#E+
P$&N?W%/#Q3D$\!Y+-1T+SAPRQOAYX@3\PJW#L+KRA#%,/ZVI"_%>'4.^M*I/_!R&
P9>9QN9!I#J#^"-DU>0;:!^D?P-\@[X/.KP 'I:_ 5G%^+;EI^U:GU>C!#*57)]76
P4\IQJW.'4ZFLL)LHO7N379:ZHLBT;DU1"Q87%$%?&-X8F;NL__)-NJR-*$U5 /'\
P4L[5U5ZC<-7JO^A]!30[M)KOA]13A.>YP213Q_,<EBWD/](\+Q&9(OP2_'+E[V1D
P/%+KH;6)V7\IE\E6YNX>D@3*1 XP+_JSRP#E>L-,ZHA*SLW)GVA9@.1"'Z^K"D+2
P9(1!0E/1*08^\A2HO(JS )*'=A>_8"S[89F?3.OQ2V<9MK2A%N:)*7Z *1#^B%M:
P1L G/,3Z5^].%5L#,[K">5GU,8;7G8>4C\>'IG*L9NV8BAWP UK3#2\T;W\Z4I6M
P*''>@K12F"YNEJU!*=ST-6DPBZL)7BI3#VAMMYO^Q,"*)R+]1+;&/W"NC&[6V9D4
P*BQ)XIA *G8R-&FW_@8UZ6$^IQV\Z,7:,?;L86,:9I$I"&^'7JBDB4N?/1E5>P3+
P&J?&"XT+[+RR*"!O\2J^5$J&]HJH%=HK8_"8EUE(Z*SN6(V=F1BP"BJ*"1-=SEIJ
PJX]W-B$Y_AK3F^K;[ZQ:$LXMFTEJ\./<Y]!%G!5(_#U%!@#RKV(1U11M@=_]%"]A
P@5VD4GWZG$^Q\Z9HLXQS'E3Y>=.MU$@%UJE3:-'NL&\")VQ2;U$=&$MK_=KCTAB\
P>8.BO/8!KFQHTWU=4A J;VNGV-,9T*8[T:YSA@*'GG%Z9.^J!!GLB?QGQ 9R%"BH
P+[X9]<:H94E0GRF#I8L([Y9/Z.1N>DUI:36'2GX(*J2_ZBLV;7%1\J4LO^S"HW)[
PKGG[MEOEHF'W:O+>3LZ".@V)K-,[U^SG?F)&Z];%"B#9#+-E4M(HXI'$RC<VRE.Y
PIB'@G64!AYU[(8MTG1%LU+@"S7/6L<(YD8K+\XUE$EB[7$ ]P">I^<+P=Z.RQ<5'
PY2[$5*D]"RO/CUE_6//B$\6*2T_'VM+[BDR=<F@>4I>S%KJ[,)B3NC,%MJN_XPI9
POVF$D[B;'G4$T@H?F*WOB@Y\"4M(N(ZTU,1EN"8??BJ_G:?19'*I@$Q&&#0&A,8*
P?;%@/"%SZZ0&L!F.ID#U=*]_+:%]0HSJ,E]O-N^!O&)WRSFF<F?+MM[FT+G:9#L9
PE"F.\UD/1!!F_4388TO\:E]IT4G@9 E=1JBRN"?%-JCT>@;NR$ISW9L=?HQ-Q7M3
P_0C%%8LE%O6]9/9PT(V0Q-RUA[)^.(K-RZ+Q"&X4U+$?1Z%4MTO"<3/EQ3^OZ9)>
PDXXM\J3=+<_\[XS#*'CENDS-[![CS>Z.? SRZNTU,'\JPX^WS.16Y/[T+Q)3E=I@
PR-$T0=;C 0MQ;FV M1EB9C<_/ZZ]\X@&4Q/B7U]?J#[@'ZRS[.B.!O'2/MHD[[, 
PTX#"&S%5/!A)8$>M ?B)PD@+GQ)E\9U12F%!X9/,=&N[F-DAZ%:GQ[;P5&- 9G!1
P6?:!FMM0V:N2%P=+8K?-1B9!!&.$.AZNVI2@]U0-V:&1F:;Y3%S/,5F'!/RV&*A-
P_.L'L.1FQ% WRNJ&SDU,',U5<RKLNK@OS8A!KN9U-L(4%H%%I+\4)G=4=84.?A.L
P_W3D.'*JKX7,#K649&%\C\EV*PH/9(3. OPPBQIT^716WLMP[;RGBK@68<35GS14
PM28L:$;L^!X#O\LKH-9:&&&(VD%F*M6+&Y@S$).N_^=IZ#/*9Q%N7K=R565;N!.W
P-51'FI[7%\-?(7!E@A[H(9P=3R7\=I4_G.[.@,2^PUU-' D#TZ)Z@,M"9;:VJUIF
P'WSS8S71M!8HAA+8#EIF8T'!+";>//@PLZWTGY"WMO019N[8&=N^DB4](-G'@7^V
P$I*)06^?$30<_!3WSAX).S3!_^64(LO.Z!L V=K?:]MP6?P5$Q_@1*%W+3C$.:L'
P"P&W[AWY8M"<3T25 5>[&VQ%5\XJ)O?5_WJ1W0NG:;=+-E<MK3!;!"X^VL+848U@
P2]R3R@73@27?A*UH9.>\RV6N\9[IV:7E5P-]!U(3'[<(=^JWBG:9^''F_D4"VO"W
P"E/!@X(5S;B-4M=G<9: )^!3 B&A:7<**JXI4@%W+[?=L<P*\_RCP)Z.O;Q2&;WH
P?)8^5L\USK!!F5(X>&14,TRBHTS@<^4J!(G:=7#Q)R 4XOL!8HCB%W+>./),T>-B
P+ZLSK!/GV-ZNP8"QVVQS?VL:1SJF"P(O[SCBZ[X]'>U!4V>#']X/E P="AUNP&N[
P*?3LQ*&..7LIU4TU6PQTT#GXJ#<Y?DKN40:AW.8YL#)P.5VDO6HA<,(RVM7V8='O
P<G^47U'8K!9T02>_!EU]G)*D/L 6H6>4,"PX*JL8_FO:I2 %:MK#KDJ(#&W!"9*.
P2!$P8>;PG-"!4IG:O!N4H"?$GF+/\HH%*#-4?H_$R_$R?!S1_<M**.1;&DP7D19P
P2'86ZV(QOM5KN3;"4;LK2CS]? K(@>C2]Z#<>>HQ3<0_G$0^B<D#Z%>H;4.KJYV\
P2*N.^O(9A$=GG>\"+"LU>1[#(WIC%#F>ZB=6SF>RA+]64!OG](</!YPM^1XM4 JE
P++"2M&@&MJ:+ Z!+C\%H9:AH9F'^)A/L-Z 7$PMW^G-^T69Q X?-=]G1X[0!_C@J
P<XE<"'/)+!*6=,N;$$;QV)!"Z&2P%8;#(E600O4VOMS2] 3,? VIZ$29D17X..N#
PG2O"R)07 2I/$P*D6))H;_!]6FZ2E'S0AU!W?' *ZZ[[FDY9Q430CN("J)F(F%D8
P640T"7!=QJKJS[2/TGG)1L)J%5&BV,OCCK[ B\R"9\T[@[N 9&%A)[S+P68XU\#8
P6B#HY#@0):Q6**;5AY6R8K)F-A2MRS96J3C,51)/L/R$>H.NR#@QAH%]O_S!$[?3
PE(<-W7%C<9R]((N!)D7*U^3X?09*3'*VV,"&EMLL$M^ *;S8-L-MRIL.QF69;VM4
P0TR'.B3)S.B&/#,\N-EW$M E3.34P4V^*@L?0F: ),-(@<W[*B?)!%(#H9L5@.G-
P$1P.ZN7M'#@.FJ2AH-QN(B&K)<+N?V,(E0MF8E&I>DZY$1CBA[_I;Q -\CFO\#IV
P5?+SM6=*1('%C?V)/QV>SN3<\FG'<,8*9'U+NLZC)*GI8V-=4.6\SP?X8&Z/STV/
P/7TZV52;*_ K*8MVCI0.,+A4),GLJ7B/G0LMXLFHN.<)^W$7[E'+@9O_UC4>"\[(
P)^>+$RLI_E=@)2#;60J_[M=>L&F,SM*VS>NR/GW0$8*TDU.P:PY/(,?SZYH+)F75
P*F8^5Y__7,UK\'H&A[>(JN$V^[7'N4)](XO,@PJAH_)DXW]*LV-4Q:UA]D5/H.!L
P.8BGLDZ/"CN' M)*%!HW[/K@0]%Z5)V30'@FG;U%3&RH*"#*QKR-<F/+-0S#"Q1 
P^!=%Z8YD>7%"2-#GJN8L2S#A!K(O^3-#=AK\%>_XQ*-;,::62;P;PDOC%(0*N_0&
P/GD]O3SO%]YR"D#$AP@,Q"OW]1<C_8LL1/H("/A.9M%@E<=)>+2"?N/?Q=NV:9YH
PP.M*W'CA&$[,Z#< FYI FW4' KDG%=9;V2^E8\WKE;F[-D7I88CS<; 19]8X_&Q 
PSV@RKN*S$!!#03[, W@2KLYF%Q<,$@V^DEY:'@=QYR XFR%AIL=9*RN?+@-Y]I,T
PPAL1SM3<,22AJL K>P^[/XL^MU,'D@GC7AS:OW77+/26?];E"=L1G>ARU:NO"H_C
P G+^B)[>=2+"DOOKPB()>BF//1:!LRO-1UUG@L5$Y415.K(:B=*.,&N/3NFD=0+O
P8-@7R!)R%4DF_HTU9OWYRXRJ@?W@,4_!700%FBF_*/Z(UT:.YJZIXO:M ?C%AYS'
PR?DQZ^8!G-\1X)1\Z-LS"HOP/T2^/:MQV%:&:^\%>8JA ^%TWWM1#&WZ!<JCR><#
P)YVT^+XZZR; 9NG[\RNIC,RGO4'7%*O\12JH"1?AE/73%UKS3$$H4YAW:WPPUZ>4
PU[WTW0CB8VZ0TG_0.B!6:QGQ6-^2G/%E2#+(..4J/"1_UXV+1T5&4B*P8)R,.Z?(
P LW)/[]>?@A@9:>BD;TH8H6)^<RYP='GL#Q+*[\L&:41H'!.?/5((P6<%C>R86_X
P?@@T;X#KF[YJX4WI4?DI@G9X\RE+4FC7!8+TRC?C8<#MU6G5DAAG7C!@6B!)9!!E
P.95C)H2#&TJ:+>>+'-;)0&T<?$P5F8II"FTBF)+IF;[^HF?LLC-9,FI>ER"B#R-_
PDJ:EB^T0VO2>:>_3EZQ3[!RN)#[;&_2RPAMU:%+O.N"[=[";TNLNDZ6'O)Z$1M W
PC43>04(&D5\77!ZXL(,N(L<00*L_/=KJ8[K!$LS2R1_YI@\LGLM$I=B571,ID.VH
PA".4MVR 8&)W@AJ4DS)CV9)E<-10QD#,7-*6%R=3W-(<[?X&/PFIG@D3H7:<DUI^
PU%@L#K1.G-GI3EAS-&^B$VAO >-E^)3W'&<9M^4!7HJ(.@KPANC-\QQC.D43"R5A
P&(\=3/L-,Z;*_2<),SN]E&&EJCMA[1:97,_#"Z.QMJ.10\74Y]S!)I^J^+ TZ?_]
P2=0NK'>/BPEG9 4Z\[L@=CF8R_&DFGW_UU58>#-GZ@H$T(::)ZE;LCC"H%573(U@
P,'_5T:_8R\?+!JYN2/$=G[*;NF"<L*<BY4>8"-@(XS ;Z*7.A9&A5USQ6-/;+KJ7
P8_GJ)'NF]866:N'*&SN,!0#< $IFJ)*%:9T"P_NPAS\3+.>N[YIH9 KZ-_LORF]/
PAL6!EV"ENY6ZU:(7+:PR?SL'&DM#KNH C.A^7SQW+O.-5Z+03'X3R?/L,U0MQ,'9
PPGGYW +J(IT%BA<0>H1/IU=YHCKH]8<T^'6)SGS*=%G7$%9%AMMWX9W^.%W19"JN
PL-4^,)M6-3%DFL#X1^FNF0I*KJ2@VM#[:KV:L#M0Y4-ASC=>"GXK0\N"5;8XSUO1
PV^J^^&*R"\QO%DFAF\W>0\)ZQU&V=]J.XTU@@MP[#-KBJ%M%KMDM=@[,P<DUC\-8
P5K.(C.D@3X1>.#'2DHG<TU\@+:$C:&&<WY!>>@[Q4 G[F1:[-4,F+0_;YVWRTP/(
PBJ>K=Q(JEI<'A"MYZ8K+8P83 =!%#]C"K5=36AU:KQQ]V;':,Y6Y\UN0$ &P<(!'
P!HS:&A-/Z&:2-_CQK#X3G^]LE3+8ADP9+F:3$]G.6 >\J3B2G8S<:Z'3)_X'^76%
PNWZ![=O8P3O'FCSBZ+(1#:R591'0K&X_]ADV^>- X_E"'L!]R38OR*K2;)^\F'C<
PF>:@\Y<V,LKXI!) 7^*%@-7X1-(^X<8ZOSMA1A+091)S2_9-_4:56[RN05[ZGUS&
PP%(HIPRBV/A=C2A"2D\^7[M#<J.J\:A";NI!R^^Q=AS(K]TKQ/:81*0?$-0 ,T0Z
P#/G ?M@'KE/<<$K4TL7OT;RL-/6M5_S7;U?()U*(HOTZ+5_S>4T,?B!*<N\1]G\0
P8JX)^OK\)5Y88E+5YXG%)GZ:X1E1-$H%XF%"6F$)D  UST;E4<JNG_"+2K9YYN6R
P3FVCH+X6; G9>3.""5]1V_IJLT$:_&R-+6!$X&)KQVCT;$Y\FK-N/4%9R3%JQ+*I
PISGBS[;\KYJ!31.1Y_MDT*>,6K>DNP9CE@^[5VE-N+=@FB4E8HW"^N2>/L?7+&[*
PG(\>9R$]B?&99$9N)ZF_L^DGMY=OL:Q B;EG)[81TZ6>;A9B6L)OW$D AH\O:(0%
P7#F^8@O[)<-;J:.\V0RL7/$H0E#T]VVKK-M/BT[0=; Y9:B8HDY0$/^HE87_%V;"
P75"2X&%X^<;+V10R<%?M>_%)I$X-^C&VCE(F+K:#!/8#UX1]>CR?4<\U;1X,<:MQ
P@&O0#[Q;XB*-N<7K<Q"0/M5"]<%/,?-/H^;')KBR?G$?$>0!F;4C6@$-W]4L\R*F
PJHWR4P8B<N"#@@A!+ZL7+W%P=#;AR,387.>-52]?SP_TG^3Z%R=0K] -8@(9,6CA
P3[J[#^%,Y;\-R^]QV1V6 EW)I256(J([];9ET/I\*_,) ,Q;ILI.TQI1ED#^5*(7
P4OE$V AR0JWM$F@]5^U/@?)>FV3M7FUA%B\U58-3K<JS /6EY3M;A:+U8#FF_<YF
P'983 =J]9@;HBBLH[Q,"M;XKA6N?,W]RN^GAU?XD6E*ZK9L.R7H8>^H]PJ<Z%<]<
P"&QZP8(!M?!J-!P((".,)@YL?V$(=(##O@*4%,<[1@AI$9WY<\BO3?<0ITQ[#H+[
PO:*DR\BG%E$Y]>U'1$D,FH+G!#K46K-TI?V<Q2]X.8OOOW%EX8OX,S91TP0%M./8
PI^S4K^$AC&$!1BQ)WUE(V1FK+87CA:ZOC&"VL,>YI_-:=&;U7S;]_ U?[Q++F)TU
P#*"6<3N-=%_C[/%LNH'4V+(_'CP=FSQCEGGFP?OZZ$'\Q0)NH9#*HDANO%] IMG'
P! M;DLMG I#!$(W 0''C-W[73F+.5X($J6:B7G+7!";7$;^@E7]S)+8^8MN'6YD\
PPYNGNIM>FFCDZ%R5\_F"XQZ9PPY.;&MR.P!$?#OS,?EWKR(07H%>4H_G ;5C\8RY
P2)B:53]%A![HNB_WBAXB[2@ URB]BL(0XNI%^K<4G',\8'=IEO%4X.3UZM?=_>9*
P!($]Z]XC:7IE735V)A2A/-5H;TFA@O/NBEDR^HFXIA-QB0\QO;!_4!J$<A1V&>96
PX4]YSPYS"G"(VM=,[%;@W)6:L6Y.R5ZO]/\VV(B/,;%GBW)/*Y>&2=48B&%$7')Z
P8U[=W]I@A)1X"V;_']0N^E7N*0G[NG%#"BS7EEMGG@%QW6QV$.GXT8&=R>8(2"?(
P5VP+X5_VKFP07X%/RKA^>9)=^7/$5&.K%! )YCL9:8>T0TBC,&^8>80U,EDE20*P
PA8?Y-UNZI0-<NG430]&)E97@8?6OI)"16I$*HW-:4O#86ZBC$(I9J,(?T2AJ-\NG
PPA-54V.1GG@1<+?TC,Y+9@0NI85#](JN@*#SA:*?.S#<Q+*;1"12'HQ=;MWXJ%->
P/UA3^O]>)W1=8O^)X^]Z#,!R?J"*]'_SG"$PE^1P]LQ(72<% P8?1+B#.YKR;MO'
P3Z"]3G07UP1/7-+G8H]7'8.ZBX@V.1)3OK+\2\O4?[M!]1\/N57UOA2=(D.+[6N0
PJ4>O(T].[ZWA9C.\&*8=@:?6]:IRO.G2P<!CEV7MQX]^G%O\XFS:Q7N9(,$O96._
PI\<(/O^BRP?KV %5/JN-B=Y3DWQ@0E89&C W+V^S$]XDSR9'2*"4,@%Z>$9@:J+<
P+?FW<*FWWD5P&<+%IN$MLJ,EY<OX:"9@;P);S$1_8>M/F+-Q]\' ?>) JW_M0N&+
P>([#=<7\V]:<'Q*R+-]D83EU)B3^\ TOXDL^@ Y>P]KY1T1YW7 0IA@KSCZ#2\S_
P.]#0"S=-K@Z]T2-;J(X!<KM*]/W0.I>1,G^D"=N2=D\^TMWMF]ED(K]F]Y02SZZ7
P6==>7<E2P ,YC)#(,5U-0@ /VB1G+_4.6<2M4VN$>G.5D;\.2XM)RU[7E%B%_%*Z
P-L.R?66)9U7G 9$C+PX^PY-3LRFI8G'[R!GS?A]48.,0N<P'GSEVU("C"KJZA[6.
P</.]HX="SKA7\KPH2'C&/@UL!MC'4IH7/Y6,2VWWXS9*ZQ+O;JY]#/!O,OPI5RQ0
PX0FE%,EX*[_^ME00#,AW(PI#*N3G]4ZDC,2AS@+S;%&%3CET2>*;GF*@:MW;;;6U
PXI=,,UB!A:0,U@_N#S#GUX;TU#RUYC=]@P>XZ_T_$/+8\7L&;)OB E=835U6,=@-
P,28)W>)]/$7(BWN,V3PN?#++AKN+VI;9IC]O@5]?%W8YJO9%S[K[*_F?IE4SV6-D
P+$ZFNKP/N L'9?PA D[*]/&O>A;0V@7:O(]5N,0SM+5 .SH33@\NAO2"'[ > ?ZS
P6:^$1F#)Y[L/+]*0[X<<YY_R=$_2U^I?5['/2+P_YUU!(WUT"R21N%/"PFAX-!+/
P0CU'.2L/BJQ4BY#D4Y<^2L_H -XR4GZ[_XD)Q=XK\YO<B!_?6K FCRHJ*>2=PZXV
P\?G(4U."E 3[U?R/G.D=1<ALJ6UZWO!<PU.4Z>J;JZ7?[CQD+_L5_9[L(YK.5J,N
PJ@(V!6WK(0.+E!W_'U/;/LJ9Z0 AUKA\UD@T,%(]MO$SW)4YE<J6PC)::&'Z$_(P
P6>]"T 7I?#E0Z+??/RE>Y]07.+NG-YL@^F9+16CPX(6P@LN )"A@[.^T*,.45?:#
P\WKIF,,5$'\RR1>+(UTLUC>F%9*XE"\G$?_3$K!:PG+O,<=BHD3<[.S/H?UL15N 
P/LU9[;Y A.]PQD<EN>9^^53,Q,'\ZL="OAFKXP'B4@?;5*/"!0]WVX7\NT;+6[5V
PYFF#"4B[GR*+;''-(GAFU#R!N'Y:F5K5E+O08<15;6\DSF'7_/?]XMU"8(LUZJ*1
P"EM#X7(+)+&(9W0@H0P<@'MB#!Z0?&0Z_"[V^;BR)E0H2W05U%?8EJ1SRV;7P/0]
P8G<5(3>.2/%LA!I1);Z"V(\?3F"5:G5_Z\=B$?M3Y09OW[.0:[=^&4UZQV,759IS
P@6QTC!\_.4M<ELM5>9]&V@(C?N"8'(Z7/F1?H!'E#]O&#S+%S/44R9:VD9^?)ZQ!
PA/^$X49M6G+GAGDD,M)+%]I7Q5?_;HGES"63H=[]2,[+;G] N- [\^FZT'QGI#-D
P2DS1F(ILN-<"/AAZ*51&TB#Q#[AK] '0TQQ5A/B[B#NI$L=S[C=M\_VDX)H>$SXB
P,=9@?+<8&[Y7S?U*ZC0>%]C#"0,DM8JIT>F<0"B$CPD_&T#68M(@":Y?8J$:LO35
P>.BI#K'D?A):M= 7:O<@R[RHUH"/X;"#_[7I5-$:86HI=LL@Q/T'BU$!7:,_\I([
P5KD2%-'0*28Z>Y'7T;@/QB+UBD'[9;V)Q\>B'2"H<RM(3Q6)*.180*JRYHTF9HK#
P)Y0<\)] DB4%XIPQCRLM,"TQBY6.^^--MA:N@"$S UCD(XWLU9FL3OS88VM,.1X\
P,+R"2&."7G<*A(KGZ_;-+87'%U]9SKUP0+=U_B25P5M?8,?IJ_[(0P)JZ_#2Y, B
P39D *%Z>UE.@+OHR0$U9/#9$'CA&2^N20[2WWFOTG]PRY>E_VG0NUI0_Z8V6/K93
P/*E@2QF'1R038M#)Y&A]1&C2+A"VG [C8<6U."HKU_YJ*#::"4=(<2C]K$;I/$N>
P\B4]U3G+YA[NS4^<AWM(=SY*!G)[)E_(VX_UF7*82.ZZXYCQE%5%C0CRN@X9\)CK
P& YNC2E6GU.L#40K<@]7!K$X<3!PBO.6H F#:R&!\/M%#W[_67(2TXCP+ZTS.;C>
P!;#N7G+]&8OSE0SE(D1UKP4[U2C+!0B_'@9 6Z](O6"K6P+7J\2Q@64'$0%-$1[U
P:6"9K!YURLXV$:ML7,@+=TQ"B7_O;'JD>\J']SQ[<')%\.3S73!*Y=* [ 73S*8)
PH#1(UC<^Z +V6<HF?."[S,*=/'191&'K]-+S><&3*X$W.TWQ[X/.LPL@M>WB'$((
PWE4)O;QE]]T:1?6$;LQS8G]'K(PW\MA"\C@LHA49OD>!=5FJDB96F_JM#+.^-GV"
PXS%.;6$62";:H68&J/A]G0F=PU^[7=LVUU7X_!"-M\O;;N&69 !6(!XFH[BA_XD6
PPGC=7>4KRN^[(R&IJM642F:3V7)KSTX)Y)<XV!=>Z$J<EMM=:HFY["GF&7&DR)$!
PJYA>ZA="Y.)/V1')]^K)CJ/6,J#+RH/=N*FLSTK^0U63";=5"-R*2L- ,62TT41&
P+AV?/QD6D9_H4?M??<CB_H]J[?>K0I7%V,V2^G;1GD6_8891J03V=&T$57Z80KNW
PD"@U,S?]:!PR)?#HM:(C!=23'H.R2&K>\(!Y+ 5WP_%2*:N0:V[E$S2F;9/7*H46
PDN$J2*_5!174K*URV2C(/"POKF;Y847QK+B\ZOC&BG#M.^X@@7LP80+7^?4L$$6!
PU'+[[>>A[U5?KWS_&SLTX84[IDT/70AX0%BO5+LJ)?\MZSN+A[&.T'GXOXMYK.=H
P]N ",\2,L9>_5O\Z@IS7!$KU+#69-_'>_JQS V;G-T(\+O+J87_VI622:3MXWK*6
P@[E&)YP*J/WU0P%]&X(*ZP$MEBPJ(.#'4H:7L'#VM$E#?4%*0/#\C#RJ,Q\59B^/
PY6M\SG+;UM#_;IR0MCUI^[((['"'L-T:@K^0-[?'ZWL"'EGM$U52-0N4@H=C="Z 
PBK:AR#^!;_ R0$X/85^UB)BK;0%/AOB#7(,IG_N8WL=N/L,8@@'WO:,R;/L9\$)G
P7*L2K4 T)QND6E/IU%2T@J@B:5X,$^Z?_(<A+WF8>C>H$0+X?;+1P!J.:0DRV!WV
PDQQ,%(O,;IS9 YJS>A.$\B[<<*Y ;D(N1[]990LM!R0Q45<^.GH^$SZ-9DO25[NR
P8-Z/\OPV586R4^%7/?T_G8SCPXNO<B)-!-#34Z9NA9K5/.+[.!.63I:4WD+\5_N<
P$<1A;+:!:74555;?>'S7H$6>4@P4@V@BTN*P8DR@=)4U;,'6_#U"CL_-'*3D7V*Q
P.#RHOP=;(39M<0I;+7X^90ZF&.IUJK=<(=,BT+_!=R 7NH"GR>!\V9!:A6[4C:[#
P5)WOMBR-L5-0S:6'F[F[491>7%]J[I(:M*[8.[6!*!Y9%,_CZ4[D02<<'RB^#2*L
P([=(#HZ-.[_K&;&QR3EY(3-<H+FJ BK,)64J;$_(?,9_"@BLPZ_)=DZ*!?%9''$=
P&)!*YMV<'J46H(PKDK.]WZY7=/_]V&1;'/>MGP]#_4/'2S(R3@R)VMJ#4>RA 6 \
P9A34H:&M>OPT!%?33 :!Q<B\W0 N_U/LB<E6OV=+1=/+L"8?7"*GM$*N&VW3%.EJ
P%C8N9.N$$[11I925AKS7MLK,HM?C:1]@^#"(9"O*.BBGL77--H%S,!>K-7(23.:X
PC5\$RK4[:/ .Q)4A@P!,$$+_=S+#*G*&Z%Q)/A*F@P4E8'0#^R@^X>7NF8Q!RU%0
PGU-(9&87-EO%B<&G&K[ZT_\9 Q)ONJ95*4/Q'OFK@H6-#W_30U1&"U="@F"TZZY%
P@U<(-5!#Q2;L/LDR4\M7.(S_]$']/ Z/*"SIZ<0*$(JJA7 ;XSM67G-F#&'5>SN[
PCVAL?QRQ@Q]S6<VXJL$"SFY"M,2  Y-_8A<#>10U8H )CL*K&R&S&F"0:NNQAD6O
P6<Z4O>*5F \O#(V::$$-ZTID\8WZU\'Y7;F"I[I>LJ(8,XW?!6)L,-07V65Z6/5%
P!]>1-N'G?R\6^H^V&:Y?_:38M_B:8X(>VK'_9Z@A[11'&\G8IW^<ST+L"X8@I!+-
P$(.X4[J9^W85(C2!\@\-V*M#1? Y7&P*NKP9S6>?6MZ24STLRU[9!O(1AP(_OJ68
P'6ZG(#:1*V5N:&& >.3<[QUUJ4: _B*9*MB0(JT27OJ;E#Z]@H2D=72I3N06KW6&
PSO6 ->DWXA]LUG9XV"P3;XOYF-:>9/LX!,]]5'G,VO==<53L M"D@,E7C8Y07 +K
PG^K%["0/5!)8>G-) >OH4(]2K/+V>Z-'-]RS*DP;U%--USRG\&9E\]+T9I5' ^"B
P3Z!Z_<[5N6_&)BL=G?@B/')^.A1*RE]==D%R^R,$H I+YA_+OY=?&3S[,?A4VDL#
P/M:1&A%6U]HT<1* %^30:,9.S\A<?JR@,@,88NIE\9@X'2%9LH%WY=B?M3S7F+VG
P%;>2/4.D$L[$#)RP99X*"[63'4:+=S_GRA$W8<R>@>[T9@2^0;&?8 X[9DBW=.&.
PUT!&UPN:>B8O/YO@2>=[W0\6:N8GL?"->D_D.Q$9G9<R"P&-!VXD]+@HX,_X)F4V
P]!"?] (A$UV70B;RP[1K +;[@OGV$&_(%X?&N6A.7^G$)!BBT!1+PMGQ6I5Y]IN=
P"!>*%-L%VS633X+6WH\N_"*V3I&8ND(369IU/XXN]*3:'"BMSTK&!]Y\ZPD.I+"9
P'UJ-LO5"YJHW^44=8P3\CE+/5[Z1BQW6;P+ Y8[\\AA<)'#;"?/G1XL6.=I0MB+]
P,]0N8M6UF]DOY9<@M1]##5XJ))C,[+.=WD@$,>48C0NFK^E3WMW0*=Y=?:"@PW]!
P:>]P0A(V_2SGA*+>_=KZ*X"454ZD5UO/7AL8_@EB0>1 5.7,/KMS/NK3Q&\=E7I)
PW6S$[N+S8F9&WF!PLE \.H8+$#W)(MH#S!S:*UMY5WLWX+OZSQ-#-'FZ*3WS.G7U
P19-+D=8G)97^>2[@[Z"*=/%1T P$&E!G0YTIQ^R1H8$TIAAA8OYEBA;#=@=F1FY#
P<%N!S/GIDPU"E"$8<K2[[7@WNVV*70C$-^H:J,E!0RUVW[Y@C1O&$J!NBI71@G:>
PA?#9W,EN& '*$:!C1ZKD%BR*EU3>&#0+6%7XZ88#&/#:5W. HV]7_(A@ ITV2]TG
PZ')XV)6=PU(N=708/E<=WG]HV:V[&"W'MFS2G9T/KU<3P6SS%?UOSE;VAWOCZTYK
P>EA[OBC?H BW%J+T//8\Z50V+ZF]0Z:[V2V:%ZGYEFWEW@XVT/R?/WKOS)G;=!<;
P_-[_PJP, WI!/>T-M30-Z?9%V&G>WI#6J/2H%#QR&M#/_Q)^D3/8F9#F[V>L/\=H
P0'=;U2J(%OX;/?V2BC1J]I=R9JMJ;](]4AMICM5HFZ<7FI,PVX2G$?J)Y?"5P>!_
PS^@+N*IZ]BD^6@-]C_H:83$&!\'2*$S%!@W".'Y1PPXD1@J<B"^T FMF-Y5'B ([
PPB=<7L&OS2IZ?@P^_22:,/6C)0_1:%-\ $)NNU>+P29EJV/6%MS&P+UN9[36I9(3
PEUJ(HB?!<XCC_B<#@>N82:=YI$-J%,]L)BSI9M+J7]#S*MH&2KA6ODL#QG+OVKJ]
PX/#5<,-0;)O7&:4<4VN+%)0M[G#8#N.(ZPD 35E\K(GNK4E1&.BN-RSQ5(=1#,9,
PX)J.AX73O;.K0L:5V,.QP6"T H[JE-)ZV@THH#+P4LFRU=VT>#L<KNW!W@<>)S4F
P,J;D&%=O>V>IRW!B <F#F6Y--4<CS40U\J=BZ+@<XYA* 29!1%BC))#\!#!#=U+^
P=&R8?4@B+VMN!Z9_;8V><@HA+'%4'ES+Q6_:?TV\)M N0IILZ:ONO;6O.4/RM0KX
PH'_A'#.3G>PJ?7=RVX4ZU$,E^^Z2:0/K2SZP>[8P&MN%3M; :V<WZPR4!.;X/KP2
PK,2FRXM\=LH%7SDK<H"*-$S^#9()>SU8&_$@Q1 \=?IG<D!G2^Q=BW4>Y0 );6N3
PJKBZ3*_N.%L/J3 H$L2KT16L$ EAO-3-A%D%@^$'W?@%I)+UC_@;Y<D&0Q_F5]%0
PK+\3;^#8Z.3Z#H;Z(E3YO1B*#S217T;G][=(I/1N.L(0Y'4[S''+'NN:F-T_Z,?&
P@A9Q'F1PABV1@TBVW743C"?8DSW[?OV44S\ED^][8^W>6*?4\>^O+#F,(+]M%5@$
PTPU;P?,@KD%_L,-]I&==(8'/L<KPZR&69'&9]R9VG&6':_%V\I?5-'N/PY\%.3HB
PN<ZQ[/7#+J,".7B$'6(E4YFF%*211FI2FR1 .@]\,2R(C^/!R*UIO@LLMT]%Z.A;
P95.:L'%#]7S/R?#Z\A132,RSDZN_0X#K A_40IX G?>46;B62?[C^13KY%'&45AS
PI/UI&HW1Q'!C8&J;9*F-X3?!LUMG!.%%N 6_Z!C]4-M];ETN3CUB8;4>/=2&X.X9
P8H?FCFW_6(GR#"9CBVI^CZ:;4_GP;"&N%N?,Q00_[(H7X9V@D/P:MP_UHN"_@KFX
PU* -Q>K"PGN_>G\+O!.)DG I5IVUGHV_4XR-6E5:IAX]MTSYA#LWD/\]6_A(^]Z'
P)O#($9-#')H?Z4M/2HVS[.FHNL\8^COAR MB"[0F<A:P:_\>[27F4K1$K9PN_;KN
P497RP<!P',GCS73@1KP[0AW1)XN!4Y][,#"9L<P@8CG-F[,R@!"$56.#U'SY,Z?%
P 2P3T&';MS<K9)O_3[Q'"H%]+I;AKP.Y\(J/[XYWVQCA;OG;]+!A\8*??G4.U?.B
P]J.0D $Z1<E54@-:[_UPJTZ*#@'ZS5>@2NQ(.< #ZF>U,-)>_QW90)'?G9DPVM"9
PZQ8Z1F'O) /^MEX61K9\,B!U;JY=;DJ"ZO7D'/0[@,.6]OLAN&Y')N?@#A&5X0"L
P_?02 X)F:S[DDD9) WO[J'Y8$?G2'@UM?@Q#_RX/[&%Q\2X%EH]R52D__*$O:J4;
P3I1IX[NBQZ#3>)&+1A-$G$1=BFF<5U$OXPU%*FH4I*K7S/QQN3\LZ^Z[+SG84O,P
P\_BE\4->FNT2;OE_!/RP3)'0?$VJWJ^V$D_Z5%+)PQX8JL#3>I+$G_T3G\5(M;8!
P71;D48B0C#B^WVONU!B2*0/IYX&<4V]:WP^7A+!-"(&05%NVJ%A/(MNFH6F'"LE(
PH>J4C2^8Z.:"Y[\RJNLTPU9*"  #CNL<7F(&!_*(K;!VP;M([QNCE#1U421VK#NR
PQ*/9$_X&4:A 25HA. GW:EE?K4*$1#_&44<E#?C.O'F9CUV>/-?\/S#W*^HIT!/&
P'JUPWNNC97P#9"O'H)/T]@#TAPCC5='O)UFB>DQ2AUM2&O$9H(I(WZ'E2$Q$SFIW
PM+Z&!S@&/&I*+V-EE3PW#E>_:Q"\[%*/'Y :*@P,KO.LOZR)3]OJ^;MM_X<AQ:4;
POC5EI 4VC.(I3C)O"'@<0G&N9<PLI+'5>C>\YB3Y%;RP(..7R$FUB=J1[@LN0JR-
P*O@IU]YC3H8\W)_<03-P*F?$OM?EP2QS%)_33 %GS1EO@7%_#TQQU 76C1TE)"% 
P*4KD@2=@A"H.*L).=X9G9^L>6=FL9,X)W/V>@,=MRL;I$R8#3VUCKRP\5SBP57B@
P9'O4$GX5KTDF?<0L99F)/G7W4\:@1GJ#PSH]+OW.8/42<F8[A2P6O<@C3-)XH\2C
P<&>L3WZR[>/"NT-UX7-@TJW?>IN5TANS\UED41B8N^F=]ZMS01T*2TS\_P(3;.3M
P#UE-;*RLQX0ANJ/-W^\=:1UG^0"CYL$OGW!0ON4UC^Y.9PGKMVK<>JS0_?C<;M+9
PAY)S^ZM'LA3 74D)B.'*=A@_EG%Q8K_^DF+O. .EVO=D@3R\D"%-S707UQD&7!,3
P,OO"</DH.VQ5?8#-%8WN!*1&+2:-1_J"]LES'RXX<3U#7;/86H?F7[P0\3<1XL-A
P>$96&L63"\KE6J25EE\8D@?\^P245DM"AH1;:V/ADUT.PC;NHPU?F-*;;\OI,P: 
PV]L%9\/W\_CM<U0S[I!KS+!HY16RYNGL>&X-#Z#!$Z*:I>3&]R8X)^3@E%FA57VT
PXA6I[XZ6Q_T=L!3D-@VXYWN^ &T',4HPR=8YCZ=*LAXXJ.+$UI@/HO.UM5 ('VU[
PJY.8-C'#OXI JHC;86MRBN&U)C/3<5E1F9']H6%F?=JMU!7MWW52@ZA/@+'&%V,F
PW;5,"/]+E&-]U7,;S7<E="<:OXA;M2+>B[A'^OUNAS^E#- -?<T1RKTA#*4HEJ5*
P;]JJ!R'Z\<R7]Y]O(W8BLJ-TI,U<C<+V7=(?5JV89*RZO&JT K./U- /B;^PX\G"
P?I^3YZ)!L=C#T&,^T4 R)PS#<GXS)!- R<LXS$<@U3>3_.K<YN+")]>\ID7G! 8(
PH(9+-HG-H!*#V OC\,:)@+&QOO>4LT3($_]5I?1-?HDU ^WV24I*8GK/+N4F_8/3
P42$-"P@5+L%4K4D^F+]MFUSE: WQJXWZ,TS\4-6<_V(_D=1HWYBV><(D*VQ*\O9,
P;S2G:ZG^'F2/+P),4 6]/=TW@[/@1'C.=-LTB9B5;_*A7CWU[PY"R&E[I(8PEO5M
P3P6X=%$W'+P9+$9L,]BIY3?T+')@QCN+!"Y-X>J6450.1I!Z)&6K&U_E9)'.%E.+
PO%*76F,:H,4GFS^+ZIX"O&623!\[B[.P=J$BE_!7" =9,.D?2\M-+JTK$<$QV7W^
P9$KH%4T4>\]3GP1:(CO(?8W1F69?UL8B$:73_EB6K73@\T*K(W\22XL[(,&"%9O@
P-L^E*?)!3NG.%3':&.P"HH62H#7H,5A718W&5EUBB9+3' E.B3TCE"_ZXY5"!*N(
PEZ=J86J#:"0?N2_+<D>7_X5WZN87F01!61,<FB-L3TY>/2R*0'8(=TM-1-6?'>-"
PN(;]CGK)BMC432>F%>2CXN&WX"<-C653Q#>;=[;*+^&VQ?E1/G[._8C5ZE+W6*98
P%OX(Q*0"LS9NTC&8IE+<\253H9'$.+*U3K]"9;L<)/FW6]?@(YI/Z+QRYR :EV:1
P?_[^J[T:P4^9RO%B3IVO&1FH#-B,Z=.]CPC@WQD#BK]Y,-K?H)X@.T5#\AZ"2K\C
P)%^BC<3U\6?\B171W#MK=FB9]">Z)>FB3#3. H:2=1];2".+8&7E?"@R@0PGQW4+
P&KUYQ?CQ&M,DTP&>J]!>1A<S@ (+U+FTIB]@%!R[FKEX6R8LBF:%?%HF&.;J]OFP
PC[['[Y* W4)B/L]5&8:20RM*EO<1FL/.OH+ZX1\V32GG+7.$:@6LOY>3$S?4X^^5
PI!@EZGF&#P3&]VFEBKI'S$82$FT+^YA0I"LR#4WN9"Q\\_[RP!K,BI\_R1['/VF_
P(\UTC)9/9C.Z:>1:]X2,21U5^Y>:8$4W)8O0 #ED39/?IB]D)>E3M=INFV2GGNJJ
PS26D9&FPW0^MGK5B!K(,$*9PN85AQ BX6B&';=8!+JO(&6,*EW[9)KMH/YKY2K+0
P@[=3"T,\OD:BQOF, Q9Y76O*U*V[8/_27%K\!!J<H?D1<JG!L368^YEYEAEC@D2/
PHUW? 8K]G1:M12_/"AL]7\]RY[/DFW42"R&RNXZ>_I8.'$4.W(:P0*3NM'IOWT]P
PY1Z;HO#0DHMD)74/[O,:-JH<@K+HN;OQ%TI6-P9[Z:748_*Z:CFUZKMV._5582Q1
P)I*?03Z1!U6>BR;Z<1>1LEO L47'$T?'J>A(A%B&RQ\E3;)X ]YQ,#96-E4BX5]2
P4L!'BB*LY90R%6BR?V>6XU1(*-';'94-DJK:8[O>&77>(;6/.HB,#"DU''#@CFF&
POAB[!&T,!RN,'8H!EA1')^,RI[MLH].,:&KZ6X@ZC=F;PM\-BD36_W+KDV&-+%QM
PRK6$%[T=D<O@E0L3I8V0$I&P3E<MMG\;.E:@%&#OOAU-(K\JNB;,5<T!*.-QYT0'
P#>")FBG!>FJU/_P6T2F6'Q ZJET1(\!<W<XE'<Z"2QHDC0KV@7PHZ0C(\@[!0C(P
P)TCF-*DI/:!?'?:'*O;GS_%[$J0:KY@"#BTVO8$.F42*0NVG('Q3K?["!MC_#,.8
PM)C-$'3^NNK$4[GP/MS-4UN5R2(U]I@ -23 P[AYALJ!%E7[!E4J9N/3/C3007BC
PX[?$$7KH3'[/O'@:JSZ8$-!SU;QPF]#_N;36PPO*M?0[M!U,(<S@O)>81.P*T02&
P6;&1S,]S?.QJ1E1DR>=AB?@NB?N_7I%[:=4U >(HCZ7U2=/'74NU)EL1_(]I8><\
P?/B,A\PI9E^3N*>>/#J?-DU/09F;.+*2^WI!?UT^SG<!EG<XE[;LD+ZMS?0LIG0H
P'QSHZ<ZM,'5-.9B_3&\FBL!5'\YGF"MRA2HOQU1'GZ0>!$R@10V_=UR>M6%=@HSK
PD6!]X)I#*M%,$NN^]KEP-L4[&^K.[:I<#RFZ\UV[\0L8.KVSA:FRK#=%&?"[L_6&
P=/,@FA*YR!^Y$A-&EA$US81C!-R1MYBCY]6M-%*7 2UHRM\E@D0QT)%A733&&>#T
P9QJ7S/S-P!* +!3P(X4[T=RDUC*UQSD9<P0-$91.RDTL]\=(1>3$F-*=-ILM W$W
P.F13B@A+D1R>&8TM?M3 \':WOEYN=:SAYQ='RO=5BO* 0O<)M<V0&+UJ1=C#<"H"
PQY*0(_;["F6N05!2R0[B_F]ZF5 LZJM2BYT&Q7?)<3IDG[695%-S[*,^]Q^I#0Q8
P3:SQGI.FT)FV3[^+CW$*\U]W?'J10?XI%)7*%;O&E)9#=7/-5NTQG:;>IHQ!/7DF
PS"WN5/)30]N2JN'#D-9+ZS>KB5I"7>XD7/(0!D%YS&S$D25]&[582H@RQ@!_:P9'
P_0W 61S*.T[@_+VQGP1E QM]@\^Y1":6,24(\7(O+P9ZTK,O!]RJB][92#_6UVE8
P.J,8X.1.N,#^"OL2N<BD8S?JG;?:)DB\N>!@\?%>2%EXI_LQXAYEK-_#[+>X-\H 
P.^YJMQ0XS#\#F!7/^>^"I6B*F7&T#C))O0R< :OR;<#&%]+7B #X 908BY[;C_J#
PS;8#0*4Z509H NJE"7XC5\/;.<4Q(RZ>CC^ .=>6PH8U,<9 ,!%/L&\#8V(8KZ1'
PGZPN1AP';E,9.99NKB3Q; 7TJN'50SF+G-.> 1T+(@EQME"BL!7A)/-(ZIE[\6/G
P#^&KL:2D:2^/80P002;2^K):M'>&^[\CM3DTJ:O#0/4!:BQ%6(R(. 5^LIJ:T(J 
PL"B_9 I]#PQN0&>1N16.7Z-LY'X7W0[CN/5-,POXM7/^=2& .6H-+R@3 _CB]1QA
P6OAXR'[TQVF79@\9+ZX;;!)$=>>Y MK<MRM;!:V_J;B Y]C]"1(RL>"W69<0V-LD
PZGNIQ$\??3DD^)OT/ 4'5#@/^Y;OJHKU_L-&E,+!\]!+HB60W!TSRT);#0*LBP0E
P]6P9':5)7HA P>T/%A:(L@JL"E8Y&[A-O10JPI7OVQ1%^DY=W-5.T"Y<PV=$0$@<
PFIT_0:GP.+K8J[H#7^6BJ5BJ_-*!GP!&HMNBSYHAD3VFVFWC&G:BB9\%RP*=Z#+A
P>+Q$[F0Q&="XT##VTX2>TD<#4WPFJVY9?9LZ%1 6"+/F9)A0H!6+TB[[/M'1D6]_
PL"/]%KAI'"6)7Z QCQO2]5NK#)D=ELCA4^0<RK;)9M,(W#86\*6NW;1*(-!*(.2I
PJ<04=76UN4T\W\87Q&7M>^3TT]I<6135F\1DP@9B")I@#$1IUGV+ +M( V[/@R&9
PPIADQ==]OW[MN(^(B(T9,+PZ(*C?Y* %[/B^PNG#$>=0;VOE4%\A=(UK33V-@N-Q
P2$XJ684M%L4U.[&(AC:7*0#M))\KY=I?]U62DHM_-,H 0BRHH(7I[R]:Y%Z\*$/"
P>]M&,QJ#)9\B8A[J$O2GO?2/058'0$_'2_023R_4:*0P^W(I[N4A3IIWP1*>O29 
P\7O'>3RI0$EY[,':4%N@YJ;X)*3-I8<)/(G'\*R9R,O"S.&'C@GABQ25/2?25^HH
P,0PF1YM<;;^_&8F73>_+[8PAST$1WU!P#+(GO8:5'<_8+%N4VF[%,'Y"MC+;\(4X
P9X1D=)G!DP]QB*_80K,Q9A:F>U8674-JJ/8HPTR"0"W<OH?Q373KI"*(,U0TI6BZ
PEQ&OA,ST?4U6\3*DTA8_S066$T:Q]IF9A(1B@/\FT7!E%'C),6USI1F]A?_"+&0O
PO#)J0CEPH76U]/3CM;&ND. D'IZIL:]\3KTY:;AZ>WK +O*JF>TE\CT]&*&+X[!/
P#B)!^ ?4W9OWO@=M6C/ESG3$&Z!Z8]L[0/:?[;&&(#,GWHQSF;S(3MVF./V##PV@
P]2Z@CL(R C@#H-IGL*CN1)7XB0I-.1>AY2^D,AELCT2SG8! &KU-K*2[$?KQ.5J2
P!:??&!B,[&2]S/=YR)Z58UF%HHYM]U\IW<L:W#A!0N*T5O#X=O//[&'$']K"TVZ<
P23J[;*?L:\Z?,B+?A>E7RA=N<R" I0>W)FRSC-.1SK:.?O;*)BO(H_/$(_S(S,J^
P/PET[ZB%!FFXX3Z@OFBY_B^8II93K9E@H;\E*\.W1CU\SA::ZB0WL8][XT+>^#-H
PC71L\/EF!FPUU\AUP1.NB#H1P:H8>E]BP%H*HWVK/="Z_J'S7?SRY$'<..QIJ4^C
P@L&614MF\4>L8)WH93]#UJ$\H["%@F-?U*H3 ME^@+DO('7FAP2WBQ/7PKPVDE3'
PV;[T5+#=9J/H:_^ER5RG14^607!>KJ@:83S;0LV5I(J2T<F(I*A52V,-_3993R.M
PSMAU_VA(Q,FU/+EM8%^C-6QI?/998C>/*-47MR6'I?Q0X0CN?='(7%L[2$X$G7M^
PO4 C2.5&2-Y2W2XLK55@+.@>T)8Z>;+-NYXV-B ZPL*&D ,^5"_::[K!< 5-%'K=
P/TG<ZPT3G ;\)/ZE=6P7-U+^X8-$,5L<QX-$2"0S^N5FX_,7;TBRWQ$5^^UWXC5E
P]>&7=O0X_A0CMSVA0%AJ>.'$A'MLD_:@/QI?=*.VH=)@2T#1.>EKZ7TF#ST,"M7)
PZ -AE4%?0X6 Z(!"[A4^*_5_J0E_/1@5Y0R.FC83&SE#S5O/DLC4^7K,K#X3;+"C
P4Z?$<F/J(^JEQMQ3E@&>^NP%EZ1,,70BIY[C95>&_29;8^.)>-]9-+.$/""DN#32
PCP3\GU^8AS[A2*1/ ,*>Z*I[:,=.T#5$O=:4<STU71ELR[#&)-;;3 .MWFC3$0\^
P^$F*6_;MMT D]NG2&8$V %G**7A8<+<H2S]L,8B;/EC(L0G]DBK$*HQ#;//3;Q&L
PNW6[76HFREG+8(_<,ZGW 2.D=CI5+W0.^K1S0%>'%$QJUAQ2WWZ9/VPF+&8*$9@Y
PPT[-+6DN X'2JK2;VC)>#JBWFGGZT@"4*I!Y4-#GX8^4%I]<;S!.:^ H)]3(;1Y3
P\.-#0"UBZO<T-#B4?%E])C5HEHFUT$YQ7,IT-X22^C:9\B)\YV\)35SAMHQFJJ$$
PQ7M4A;P2 >>;TZ2&($55QJ?C[_[.O%9U^<!&&=(*$B4X+R&9X"__ [VY-?W$M^0.
PT7#^Z)WE-0:X0Z#!9QE^?V'Q!6?(41315K\K;)C]&/:B'D@YFSTV&M]WD?GXH$$J
PYUFLL !XZGJ!2#4V,A9>7%9%  45R4?SJR]/_98!&SR6(&!F2/53C<GHG$W[]=<5
P^I:BE'KG96F>,?;*B\_:V![JLQNK1"U+]U_HF#%_$IEKYL5PUYDW3'*UWP*=8)M[
P@*J) "M]T0&+VF-_ AT&(+/3'OUC[NM;86^_3C+;YF[H2L^["5)')J---+]3G,VK
PAN6R  W* G3:C\DK)_0W25(8?![X[P$*=3A<=,W%7'KG:RC:Y.0<GF"O!-^,4KE$
PDVU:'%#3LP3=BHS>59)56.[7"[D/#-JI+!OE-!I5*[4X-D<E?<'4HC9OC W,EMBD
P2>J#,156<\2@3[="B-'T/]VN+>6!D#@8_"/D@M1>_(-/'K\F%W5;2[@0QU:YCSQ 
P['+/U3T3Y4!PEAN5WG]%Q?R>^CVCZ+C@NM&P%ZX(LB7CB[0D_Q1$?5[44L63D2-Z
PRMQG9)@Q$V:E[3RLG?OC*:"UM&ZJ\EUN:.J(BW"GPQ'0;R\@5=*,0B8FL5Y;=M=B
P;C(%!Z=NQ*7AFQ[Y\PID0QK FX9#;KH#:)P)V$/6$ HG[?^NIE)OXMEX+'4=?]A/
P$(HQ/!K4<H1AO04).[8=![O:X1NK%H8R7&GG@Q[N40M[M<,*ZA&,-J2,HLK'?+AA
PFF &-_U+5,G7UDVE<Q2AX,F&C@10]@X-/@@B;&L?"=@*=0G!S-KEE2)$##H^VJ39
PM^8M0:F-!IV9"&F^>+I9F'K,N<JT+"A;S9^+O?9WRIBZ#D 7(!N\VRHT969\[?* 
P(QX6/MP"+2((#N^<#HML@T ^=0T2Y F\-91DW@AKV$9 *+5>?=0ESRU?,3F(A@W!
PP#E67HVA5(>TH<=\26%K6&*,-?.-==&< "*<D/ZW3,,UF21.C\!PAC6<[UQZ4%36
P\^MF1#Q*D',3:]FPVQV57'45='7J'\=1"><&OTT(40*LOH1.(>NKEIC,C9@7-CUE
P>)_M9@MNTFM4WM1L0)6+L22A58+*"-?SO-&,5'M\V:^1D-3!"."Q2*]9M <G=9VS
PG%O,?P"8K/M8BE-!K]A()31:W[1G-&EM?_/G0G3:?HW_[(4 ,EGT\&1C1:/=US,P
PJXE29,&3.1"V$T.-6-?9FS"[<@<()9WMJ?UZJ,@1^\J^!<K:PN-##ZL05#4.<!#D
PCE<#LWQ9 Q]0Q#Z_F6J'H[N\^>/:\A%Q[2CY8[PO$(NH;R6A5[S P+EM.^XX/VQZ
P[$7O5L6W_Z!OJIJQ%3$@X7!FRA0<^XR.@';1G)R6$!\(K=40M=!G?^0#W8-"=X%1
PK=Q 9Y%J]D[BW4U;+F'WLK?#8JTX8I.G/P^/?"E,G%/+*_)9 #40QDLW&0^Z!$B*
P'EU]2],TLH1&5SN[4@:@C)'8\>YTC%8IED#ZKPK'2#/-Z*__C3H:$N>9AAR8Q=;7
P2E<8*'V(38/<D^%,/1*MN*GL4E<9ZI-NI:Q/[N=0)G8D1?(74NM8,VR?MKS(@9E7
P5^WC6&D**1 -C8S6'7D?LE]K?4G_U5[(O-WWAY*\!A_X/]WU.39?RE,,K&%KK[Z5
PS2W#4,"5.[D=$NGA<>5\>BVUE(+5@1WI\(AJP$RY)&:&WF43C1?UT''+*BR#1_V^
P0TT SK;SVY=1!8JA-N52ETV=N#J,.=[ M0)M7$&E%GP6!*8=Y"O2(?6F\[+)%';Y
PJ@IY$53ONMO$H8_6OZ+..HB%BS>#SV,W.2>R]LXU-H&&:KOE. R7:K>#/JI.>(AU
PN)NPSV2QK7"HQ^-H0\1"H=1.1-DL+W!UY&JN+Z6+QW:DJI1ULY"7\O'OD;=9Q/O<
P-]^_]$E_;F$0ZW@@/35W3(,PGN?=S[>"^-DE]FPMEX3G92>N]+-5FHOSW7LGRL3/
PLA?0E?JT_&8,D+N$[V[*$@XM37;D(DXM 5RGG*^XH..\( G],_PD#/LGG>D<.I(T
P'Z'R9+Z>.]TO3P[I6 %XUTDUW$:#B/1H^J6161P+P7EM$YV**;Y7-<)!HUD"YL?=
P:^[:<D0D&>)D)SL72*]4L@GAM%P\]8UF8BKZ(EK:CEF>VH8'C2X O]4)*QV>(=Q?
P3@,(P,;W9Y->>8Y';4! C/P&AU$,$<?.Y")*,C0[24Z*^83^P&!T2W)CQ6*Y@]'?
P):TK1/RLH+FV/@HW="G<*"<&UI2,'A:*"&8_X9V$\6=K 4X:+F:6&_I<<(75+YV9
P.[ $:4WV!9VVJY.+"9JFO*+'G&\&;S,B5^U0.O)1_YJP<WSFPAIAFQ(_(YZK_ QH
P1I'N)/"QNW6LV)\=LX<=R*2T8I]RK+];0FXY^\-?J?$E&OEMV&MJ[%%?(=>C<::(
PP74KJ(\4 OL/KIZO\^3Z$Z@&/='$ZT4*^RVG-9"=FC+RK] API^H8 9<=#&[02@L
P:1U,E,E0X))(#C2,^:55#=^X1%6<GQS^0NTQQ &NEHT??X290KGS=G=@5WM'X)^[
P!L0G%]Q.\%PH*[[,;:_PFS@@.$II7]W8FP'1:03D)G$NEW+H\'#KDWF-OH[AA<*%
PJ] 2.S-0BGN4+FY=@J=3\UW,V,URD#&\P.' !#^K0\24QP)G,':"QCX16A5N3L(#
PT*C)WU@3)K"/';QV1H6P\.PV$?'B&RW6&I+/!#[OYFPKF3W&IF_,?0:I>">G&X\<
P,^+K5 *=XK'$T2T7V1+9S[ZU(9K!+N2T;B5-OGAQ6PX8<*CA&C_<YB9N&*+9;YFD
PP$#70UUD#WW2NI+GR;\/_>P4,T%0CT+"UEN>0PO7ZUJ=,B9Q)>.JG*$8;VIC48RW
P%Y7@RMRW';%%54K1^M_A_X39*5BAV?@8ND(D0K_$/U'&0($<6O-CH%_W[CV]%\)_
PS?22!B;1- 2T=OS6L(I@+:D5 FM6;;]H]8.E]Y4OHF:A+ WTRV5O&LH-BH/5<"L-
P#&T<"UA7"6Y0%QX?X0837_D7I1:=\GL^B=&!_9^73JEEE+#5)V<$IXM<BG\KZ:NB
PA:4]]O<G1--BR@;@>H/+JA[<UI+"87O\7H#U%AV((>B;,% /#4"GG^7'0!WPROEY
PH/%E<6NY2OL>38VOZ'0G%JD40M*E!!>E[S3#B)(&(G2)HPH<,AI0-JQ/JU&N>?YE
P)X:XA0[<+U31J4(4>>;V&D,M8;F;+F>''PP>-!R'"-XA3@?P@=CB+)+1!O[ HHR9
PO6K=%C=2:K5Q3_ZW6&&%^-2?I@T!N HF0S</;FA'\W6.OJOJG4&)YS&AZ>BC(=[_
PG4249_^8?VH;#.P+K&$S1-L>7TW,G\Y9_H&6<PV],!?NPTUPM1YKJ19MWA@9<7=Q
P13PYUG*'-IQ-4I,*K D;("'XIJ;$WZ)V IV."PY4IZT[8G".Q\.+7R2\ IMYZK(U
PD*_LGT[1S%_4@+U<RLO0@P2^LF;5I^_K%P%.1K+SY^P[SE"I#.T0KKM3L0N%?LU\
PVTBRXF#$S8BU2+Y1L&C86-_(#866]ES@!KT<N*O]\YZC.&LN'G;CBT,]"U]_3IJ$
P'OV^S'J#S$_.2B]02DOM%>S 9L)!>5-U[Y0V2/<.2]\'-I(1L0QS.LK9MD%;EBF7
PK?0M:E8<)V^6@.2;(G#+U&D9G')QOF-'-$3//,6>QXHA]J1.A%"<MR0G]05SA/R,
P]AB:P-/@;'S#5\K6 MC2;\2<_.'C?\]LNHU.[,:Q)!F<X?I.U S<#<1"?K;]R8 <
P<0E+3H+H[T51S@/8[6J1LW$*,7^2]TF9O<A;\F"9NXX7?MK['O5_"@KS]=2B?61!
P_F:G#66@^:N\G MU,E#'R&MTY+F#MU9H'\6B#+NZH-!S434[)*L12'T313OFB2B(
P:NNAEU-XS)4 Q_<A.9@GNH<V-L:3B9I.E3@-5XX*1*XW-V(GCZ%SR"6[E"G96L(O
P@:&,L!3B\SF>_A0D=U3O/,)(I#YOGX+"!1&V]8';,^B.WBH3$:?HT0'Z,;3-=]IT
PM:M?T1:!\'(C)\6A7+=#T874?+76)STU@>CR^Z\Z_)8. 2DZTF>JZT\J>"B#$8_D
PN7I"%]226Y:BE7)YH^OQ1CU]_\!P,?A-!<NF /K0O(8F*BUJUPMY"[2E4!T_"(2:
P.3MG!C_L7^GP(FS\3/]NDAEZQW'[B 8$U",W*^H@:R$-F'>A)Z7F<VL_7J&EHQ='
PVI>/7[C\W2KV$8CF#?G<E"QA[AG78Z"!C:/;C=',PX#SWHG^P/3AH[;:X:&U=FW]
P>YV E,0CB6AXCYL* GN!U["G$.4:$ "9,A?:=@:W7Y8L7,_X$AMW<D!]2UI.9!\[
P#[@90H28 +T)8(*0?Y+QK^$/H^;?8CF6I?7_A;)QY)T>#EZ^\05$!)XU ']QJ4BK
P_[$;/)W^R]-5(=PBNX4\RN*J@L(BAI47L8MP,[K[1BG?\CJ'F&\],N@DD#'*Q9HO
P&&6$E0&1(-]E& ^D,[HV0Q\Z%TAB4M[Y_;@K8D$(4-^ODH.J<H_M+_">H7"1I><4
P#QO080B]LD%[CH"_VV=+GQ:Z.?JJ0KZ/#/ME9PP=ZX/N$&B03<9E$7JQCA% 7-C-
PGBPMNI;,6':8O1!EO-DX,5F?56F,.D>C>)RS[C0#HM+F[8K[T:QO4E_\>:8ZD5U&
P4:G*A%91"MM5H,<,7#7IK4I4L/*$0^(BK+>#8UA@OF= JC=(\9MK,F^5V-77/W/+
P9 HC3AS^%Z VJ(?X<#*IZ*AF021>86Z#M\*(SQ..4Q!: *6ZKK.E[KMUO*>Z %O(
PZ>6:]D,#'O $Y,=BQ?A\6HJ[W[_ZD< 0F,:WSDPEV)RK3U(MT<MT[2O4OBXR=E#"
P/A*XB-76-R.[BY$'U52F<9802NKVC[/<MPLO(GBP2_F&HUQVV\)$QUIMDP+#T#2O
P=U+]GG&[$?4'-*17,RK.!(1/L0]*=222&P/@.C+H*/I!K*:K9A+/I,W+*31_H#G7
PTC+F3:S83Q105ER+3RDRIN&FI&3V>/C 7<"IR$FBJDNML;BE;$F"79S'Q.'FB6@1
P-ZGXV620!@].MKT+)P('=33V/V"=;?)6 Y8[VE?$FPB*1?FI@"!%[C8-*9G4HQ1-
P.5;HU"%@,_UFLXXNX[O_SA<IT*-!-#4W\L Y#WDI]LREP$QBHKJ<^/0XP;-"#\38
P!<K1UFMU9[&"1P#:#= N6R!7F:YV.D.5CK70?&:\X6KF3U@Z$B\419HOS58;&$6G
P70^JK1PC?6S5YH3>2[]%$^.!N8L,_JAGF5%BG_SNL=1.LA9.@T+NM@!WI9))M<#1
P]^+L/(_8"JYZDR)A."Q'V,GBFAG05'Z3(([> WPGB8O;OK:E;IWHSN9<GA R#FF<
P8EUAA9KX;6%36Y(;*4CYQ$O<:0^ECFX%^5EF1HY:!2##@? L)5S"4$^4;529^):,
P0,W>Z/B0J2RYS>/\_6N80_SRP:0XE2NC?\T7IQ31BE[1PMCY<V>='/H)*/T8>Y5\
P:EWK@X,NZ\!QB(Q6T=)(3G,]8<;5FP,4DL0ZM&BP;);6QA>.:\\&/J30!9_-G%DL
PQT' CJ=TJ@6,5SN22\$A17KZW&=\%Y0PT(](*^W#*H/*:]W 87R5&E%<?\7[K=0U
PIB>GV6\V-S(AK5UTF9S9U(3]@1L%<;,82VAB68,K3>K>"ZKF*.?EKJ[6>)AVM!GX
P94*4%(RW0M8=]<@VB/Z'A/_81>,O 9&,?E">)4KQ=UXN05HVOEU0='%&0)E3_DLD
PRA&*LZX9&]7\U)=9"_9_BC'78@*9QBW[/W\=*LNY9H/(P[_D\T0NHJAA-J3ZJ?(9
P#CF_N>C!5_6=$U5'U%RJ+IP:G#4<ZJ5=&5$^Y5*/%7/V7K<>3#ADRC[O(MJ0&:?#
P $HTU1J8Q8ZNX9)H@O/6TI4'P7U.U[L\&!;Y!TCW6.IPNX.O;S=E#;4&K<((JX04
P/;2SAD[VWD]C68C2,_!!GG@SU?D<#CV -$)^@HD!"JZH]&QRW1U3Y_)U4FP*D;W-
P9Q7L?Z R7EZ-53UH3?R&N:&4/J#(FUSCPEE^;.EPX/1S[&P_[M:Z#7C'[JK)SH)!
PKM]'B":&,D?+ HEYZV+4YW G0&NAE9%#XS2;<ELZE-$E=E28%B843G&&^YQE+V9%
P%0P[(CSFAD1C/+7=OZ$CQ_I4;ZMX7)Y [ZW2)E%C>5_ <2S&?4++M:L0Y41RG\93
P*IDGA'K^K/3NX A+MV$T-5$(?>_OZK1)HY5NB\_.'BK1G>*?F1>2*M7I?=B4;C]+
PFZI>2"B/:<\IO0^2HF'*1%>SM;+'=CJJ3H%%H;<S\DV4_PW02,ELGA;2@..O+;/A
P@AFB*Y["-)]8<'?TY.X6]U7]9<5N"^8KJH[S5C2RLQG1X",;KIP0 ,2/'".[$X+F
PA9A<MO^DANW!-(KRB2$"V0"EA5V"D-,<<@%MTWBG[?9Q!49L7QG0Q S!WMM\T$R8
PD\1U\M0K,KVZ 8 %[+_K6I^!JP?<:2!+.-MU@UA+*H+^,090)4QI/5GWI.R&5\SA
PEQ2.RB/[#"#&!Y3) L$@[P-FA:42L[&1C).]Y )W$T_0KM0WT<?6R%FUP)30&OM!
PD?VI VD#^F>H&EKA0K#(266@83EW.7&-.['8O%01 Z#I"??QZ'*W\IQ)L%KA"2SU
P)?U03O7G*+6MJU2 U9_GJJ\>O6O]\V22W#I!^YV"AKZ2,0*9B8ZS]Z)WK\7+X?;X
P*9LVX.]"O$;,O [,L,<5.B]O+L3H0U)BD24\N\Q;1LSN=^%L@'BYA.=1928O@2<6
P98>",X9$-]>]^ZRYC4/)GY;8G2].1"7>NS>H@%O1F &$$NW?0$S?;J*3AZ$N\GV%
P=/D&Q8#JQH\U%R/TEE'MWC[@X=/]2E6,+0VSQQHIV20L_YVX-,4[JADU'#EB6+J4
P2##6-+@4G;KP #8MTY(O$.=&F7Y)#HU,KIJ=@!#GFP@FY:#DVOWDS4<PK$9(^K]Y
PS[ K,5IGBI6WN&)3 DIB!8<;02/"^ZH(45L2P)BV>:$"LHJ,,!J]KHY_ZTMKKU,]
PIX@/!7%Q4YAO?BB8E&LWER+/0)8Z,EXE/_!I0IC<0+/8M%1L7RQ^K-%5*%[^BZ47
PP=X+L:$'7"J7S7)UG?^=7+.DQ(BKJA9A15A^&TU_[MXD :(C^UK;U\CM4ZE=+:K#
P -&;$4T4Z>"<:BYLB&E2G7<)%)*5@XI,/:[H)? ]+/Y\_J_\+V__F#G@/K/EZ'LB
PN/ O)7V09\7:I8MOPQ!F\/!;58<0I?S1@60@T%'$FC$EG#<1X;VB"#>Q?L.]MYNM
PZ2F<0N)U".Q\4EI M"5)N9H#RL6EJE%STY0=S'*"R\V9B:KOE(G\@",FY*J.Z%7E
P3 @P!8"B5V)PQ-W.\5'KQ.V)";+$:WK@,\E081MK".<7M-,B,)=F<$X73S3,2[,*
P/*9W#D,==IX7=+T)IS?1F7*,;5?<4G(CN9_]K@4.H,B4L^_'":[6@!O+3-PGI.8.
P@R^J!@;VOWJ/MCM6U([CA 3U "4#&G7E_(Y?/,X5Z]%V>8A)!#-!# PZ0WPG+O;$
P=EML*H(O5(D0AH5E<Y9B/V@H<A[J'LG:7\[R0<%YB@O6_$U#?!V(E9[4T56#N0M#
PGS7WM!]I%Q"6>W1LTR1X7:7Z"XL;VX+?0HR?@-)[%(J;JE5IC2)D,"F[-K_;_:)V
P1RXQF*0@"V&P!9S<--;T!U,)SWY(3=J%,<Y)<-W&/:5V ,#%=4L$T/Y(J' .ZF-G
P38S,(M&=Z(Q)8#A+8U:R1X8/*Y12>\N.\*%W?S>L%B^F<B/N\)7B!Q)HB@8"!M/[
PVSK,JAC^%X5N])Z'VS9.Q-0OPK@(3XN.WWC<$]R?U6?P*.-P/N>[1+E0-\%OWN<9
P:ZJ8ZC*9@_GGFPA/Q]<&T*6>//.F;$&W[E:9+1Y=K4^V(:BFJ/(Y2,CO2UQ9D= J
P9[8#B6YHM,MU8@>I789^F-3C>S*UG9!@<C)"O&FG.1ZG7P(3+W'B9J?2@ 0%A2<=
P(F3G3W:OI(Q,362E.R7$XG%P&VS%=%T[)4%.&NBZ_Q3]0R]EJCVZ-C/JL5";1O.?
P,J)W*@S18L@*X;W$"BH9\ZH$:<ISXZ>JH6N'Y6I(FP]Q;VRT K_-)>ZMS$*JWG[X
P\E.W<32K8S0@47WJ'^P>G0]\U+_5"_E1W3V48,\+PW\AO[X#7,"0+R4O*/J[\GG(
PO<)J;SVBK=$U-<E[SZAB:/>*:]]  /:)#;I4EAGJ;E47780+@QG'BWPI7%=O;W%Q
PGH=+1QH A[C(Q5YW2D*MQ8)B5X+D44RNB@.A+Z2HR+C8%T>9Q<#8;1PP#N8YL%OT
PDQZGSX>DVS<*'319RA4(U.%U$.CRP589TDK?-KTGX+FX!GQL:LSTE];6_X#&8KO=
P7IF 2Z/1PN-:DQ?3Q[]!0\(D)>2.R4M1 .^-59XM)Z&KWW<U9O#X>Q*<>_</\I"Q
P'1J&P;&FV766SM_;D$;[_>,_A]QY^^85+M&PJTJ88F93YLY-IC8R8T^RQ)L I%H 
P)7@31:;?3*2[NW1ZG=!O+T#:<5S1#SP;C(W\' (L<<.$K"9#._A/2,G[9C)5EK"P
P%#KI$KVSH#C9N.(C2>%T#=0FA&N!/]L&,RF"C6PC.N%S9[W!X"FE88^W+XC%-4]K
P</.V3 4?ZW"CA)5Q#<4%4!*XT1:"G5\SI48KP#-D*^N=D.IS6[SB'+RG"G)6VDM_
PA*;IGL<HNN?X!W+/K[=#$)<<N!V'J%%M^ROX&3O)5>:0$EPK]BHM"A(+<2_ZF7'H
P:R9M[-:A/-!C;WTWB$C(WACS&^4SZR%WT,X\@LG)Z1A%:]Q+0A3 \U:=R+;7D>R8
P]@O!GCA>4T[5\6D=UQ$;J99P2;*0I@0$XPIQ;V9N!A.-_,99?+U'G@#9=^"\(_"Q
POG)0O)D;(Y9"(^XK@YQ^QM?I+HBU\9:AT=&M0 N1;]F4>]PYYHJ9B!6^;H<.W+S/
PU28#G8UD]%(SNG%5Q^[L+Z@BG<G[):#E5]H,T="+43K+UQ=GJ#K!(8VAG6XV:P]"
P/ZYJE]Q<-&WE(@9,Z K+CY/Y8NI35\N#;=><O_V44RSCK<[1%51%-F&#M [UIOIW
P3LPVL_(B'=T^M/LOHD9C;4[J0,Z7(,0LY\A<-B?@&\,?BY/H)D=DL("63D@"HQ>#
PXM'@/V!;@7@5BONB1W+BLL!@X[28]*HS,ME)^'FI_L?")R.QL2K4)@GY\/=H$_UK
PTC(+3>#DE&=P;3?(J;"\+FURE$U%[8G<SI$-/W:QJ:H8!G[/'5)1=7<S^I6) ,R6
PC9(:Q]V@E_,QNVRMHHC/[_$#K:( RP]N.YB7$I</NOYVGY2L+TF7XS@@2[N1C>]^
P!\\^OX*T1I$)G&0X,M%QNA5Q)0)$;9S3MS$<NK'ESR&5_S!%Q8:J^D=P*W@< /_^
P"XK>3M%<Q9G@T\.@Q>0X!_OU]OF>VT@<I\T_<_T%T2F-SV]H*BY5%V *W])LUS>2
P).!*1!?4*>8E476?AKO^^7ZDC*R6/F,N/I*"<1ZNQ757,3<E-0/6MWT?:;57YP9Q
PTX-9AZLSJC&NU2?,;B.'Q$!<JXU7YR-;+IR<=&W0'?&77A@R_WT#@Z]OAS%<H4$X
P.G:[:C%FKFS\<)^%19.$'O8Z4Q%U]2CJ5/K&&%.&I!M>^6>E&UZ(/A+*E6,2 R[^
PTQQ2LV)%9SY.7VUVYC:/7R'X4AU6J+*^%A(X,Y$>.9C(\K/'-T>3&TAA?B9NPN_X
P+Z^'",;\A /)7V&*A?"_W,OZ;HR6I$S1A0_T*0%IF/YK?,.Y3&B<'S[(Y+,S*=8\
P5I@0_-6-TL @!$R!:\CS5 /*YS3]*AC^*.=)A&J&,46H0*_T.A1G MR@@*G'>\/\
P8),0Q!X!2F,R+(_'-T=48Z_FDIP9*.D90M3JA,"$+G,H"![F;?=0.IRW*DFA>/(I
POVD]YZC5UCL*_=.9"]UR+O,V&.95#S)E%M/N=%YU0Q>R[8:AHX#XAJ7\!UZF'F4!
PS,4RL"==%0P-,'G*2SK1T^+7CYLE>C%@&'03+8'KDEX"Q_LCMND\@IPJK\EC:@[O
P!IX0IK5\^\Y,#-(B,?&2>6UK+8<V=!/3B"_-P(9V_3<]1F6A[I2[$8J$G^Z8,)XX
P%2@U &X\\EP?B,^;9QM+6-^;O@WLI.189W1LV"[-QQP,N<94BK@T!,:W]HFR07YR
PZ<6:8,URM@<N+;4?=EBA\ 8O!I]YF[Z6QKGN^"L$F&9)BIN8:IQ,2-7[W;QNE3\J
PM;G\IS9:S=2C=(*6(8ONYK\T+8P9GS0SI;.35S*I?0 *;/>V\H!A?&-[2 D(]W%"
P;P%AKXEG5NJD82"3?BW5.3\P,B^AEM9=/,)"M;B' %#0H<-3PZKW^ 5/$N::[ ?)
P*P^BDY)G['0X*1IL"]SHMN12FG9JYT(STY# #X/C/ R>63UWD2S>!OKJU1L2P?V[
PZ3\5-E='<-ORYH4T2N,\*0.JPVMJA@U#S,896+'Y:VA(;>;,2'5$8O("#*\RLSNB
P;5K<#53[HYOB?"D:%SX7%^C0)N67YD9UXF!_@Q=5(Z346^Q<BO;0C]P97GZW0@1I
P,_5%*6TDX\<72#<_'=-S#+\Z,\HTNJ:#=>U1OD"IE5*2]K+$[BGY_'^,P=<^/1HN
P[_*(!%EQPKDQO4 1\DE5DBBRDW4G[<!#87R[,(#_])>FS^1LJ^JCV=@>E.V+UTNN
P(7"&?W#+251:1.R!HN#5/U^[S30!W4I+<-$0X'J.:M?I2N*599K[K!F]\TNRH]KH
P<F&HJ!\7MBHJ@49@;[_>P)[T>?75M]1*4;<V73-'QG)C.@EL#W\9N63:+.BZ42=U
P0@S8Y-5+9EFGLX#D\NO18AW?6G?L@QL*P]J)I#/3XC+% [</U&)SY8*^F<#9640W
P+<^*XSY7R$E]K$%A!F//T;JF1UAO2IP.=</P/%NQ;\*3EWI6)8FJGR=^@>5.YC?L
P\\0"C1*354;G)LD/XORF%6M>/H?ZWS?C&<#Y9R')XG&'A2DUW^_D2#VBR5)'1_(W
PL(;RHQZL;2LP)1_#['$3F   F71BQE/5#9VQ5R^=]G3*K5&"3LT.D[.T!N"[-]1X
P3?2V'72^#U'><[=+Q#H@Q@8*T+Z,+1B"JX)C#R^23!!PXQ&T0F'+N.Q$VKR1X&>>
P(R.D3C!^S#SR:;I!.;+##OVNTYIM@&PIUW&Z<#=L,"DAR'*A*K/A/V,3@TMY+.O,
P&?%&3>7\#0GLC[N.D48^^->0D\]:S"HRM-R@B>A\]&3#I3WBMDVG 1KF^S:DW!\3
PM(M>):I J:2B!XFI[/_Y(YYE:E!R[*$!=[WD<$ N+6*7SBSZH7%8RD,OVO)2/T'0
P9T++AT'<GF+NKF@?9FL1^%YR-#+N^\AHIUH6_XJ+5-;ML4DD]!1@#%@O^Z<"V+ I
P%JPZM$AR:JCO[YU)3;"QGF3J7@2(!H.2J>G?SVA)2ZF=7]Y%#H$,W[I7X'E% 56Y
PL,?Y#T]U<0Z-L=FT@J01I6#5#HQ"63LHV"O(I^@<,=#POC=8^%,/9Y)U8*[/[18&
P2RL$P*B6<PG&GM94,[B(^]&S7ISDSR5K*Z=)51@Q/#"96>;QT'FK! PZ^[PLC4M<
P\2-LR5DL2X)V\L+ZY\A# ,YWH&C/MKQE!0H)V@25L0 ,/&I&#6RP-9;_T\-X<H>/
P_^K(1=83$>V]@P[\!NI8<U %<=GD.;PQ;78=05G."V\.HHLDP[WR:@X&?_ORW 4X
POCY&607DY]QZP%,F,NFN.&6;Q![=!#675/$_5?<&=&8.7L@=Q/YR3EH2)G]?V7>@
PB6>WGZD>(^*G88T/U7WE@2L=)C.X+*^4\0+)X/&M\C&YC&U)DQM0,\> %^]UM[&M
P%1]SSO0%JYD5_-P0 I0X6;U9B V6F>ZG\ZNUUZ/R@^1H(/N]Y>!7>X'V[<P%\E.)
P&1HUFQO"-LIMA,P5#U9]7VQ[N4QZG7I[Z8-[1SL=0G!Q?^8.RNP-V0'LLLB)UO"1
PADP,#.3L,5IHA:^%J;ZI>N@X59RP#XNM U*WD?V?1L<B?[4S)\=4T?U^X$K05J^!
P;AORF]\.0#SD;QK..P&?B#2,P*V@A/Y1_[L"GN:(1_$M#O!I=,K5_QF_=Z'\3B_>
P.10XCQA ^M_K=U4'#0>9;\MF^'9'HL,?+USN4NIL&"!B:,W7XI;D?_ZXX PA+8C*
P0I0L^N\!Q5(&!YIP&[SY9A[10IJ<EP(XT:YG47FL*9LZ$P=!2>9KX15]=Y7;IS0+
PE1+":G*BA(RYMFK5BX@$2344$@' .$<R^:N IO"?Z7*A HU2.J,HX4"18T[GQC&7
P<@S] %W?S0UE;PT1<OG\J3D&FU;T ==//NS!4[+C59?S:4JU'F(3A(;*S6D)*M16
P4\?.IA%"8H.*0X58@\( M&]R!"[6A-TLSQ1@>_^0EQ?-$%^L"Z9!Y675\IMJS$="
P+8X1:[<RW&J4'I=8-%207P^E(<1?Z_&M1Y=_$K)7Q[?!N'VJ;K@M4<F/[H!YMQ %
P4Q\<9?CO:'3QVZ& F?UCC\=R2B(SB\3XKW_1OP2O?&=[*YMK81'<1+!-,;C[4 >C
PCWM?=;B85#3J?L>040#6L$SNNHI2KL.1F(.Y>WIG4!:;M2<8G#E4D.7/"HE9=N8;
PMP  #TY[SEX *OGULF'?#-0N^'0F!R Y\@+S:?H&C$U+@];KP(B)!1U*2GZK5&L4
PQ9^2!^C_WEEV-F4:%)R:2?:2T(9*FOU-SZHL$P5TAU"3XLP;3UHJK)\:/J-4+,!U
P<_LH,:OET>8'G>C<\0GF9\%P!&V<=<_T>A.YL9T>8UZS?4R0Z((R@?CE[/72$%9 
PUV^6.1F9HP6SKY=_]1)'[C /A*&JNWKS_G,.Q\IQD_E1^^P_\>K)@]F\5>FB?.= 
PXJ7/G:.WW&[*G@%E903G9]/2"G^3:6IT+HKG"LR]K\=FNA>J\-[> :9B#J+7KTRX
PRO&> D(ZQVLDWJ1DC27[(A"'-7$)D<M<QG<3;Q=U?J?Q1]?)'.@4*LYX=\1PX>'(
P,M-.")27O&0@2;Z84<(;%C'1C _()B[)H+=E <>;8K3[<M3'YSZ->4D;V4COQ]Y:
P(\'"%!3],,B_E\$TQ(K5>B$R215#AH[5=YU!H8.&LPRS$>$C(5HN2\5$27*W6[/5
P@]C]QEWP<;O73:;*MN;WJ6#4VZN1Z_<7C]B$P:WO7E]_C:T "H_+]A>NJ82^;?IK
P:Q1H,PPS%1F[090ME'(YHHDF!)M>\F:%M.I58H/Y5W$8>-)=[Z!. =4:8]:XZ+S[
PYN=@)]@4$J""I_0K$^\M-\"]Z$'QJ^]6GTY0)$T=JOP")R\CZDK?'MXWO%$7*@I-
PO3_[#C'@>,@/&DI0PID'[L%U+GEP@P.Q$3Z_(^YLN(7Q+0N!%"4WBA\TGMO8)DRH
P";6$WP]LL/RT_S4+1RWW-Y;I\/@5>+?,5/)9)28MSW<RM=(]#85>@F^<Q5;>88RH
P#^/DT\KL'HFAQW#0[WMBPP9+3F-1\^D^Z0N=(S]*,L>&_YX*KM43$;CYM:H#'4#C
PML-ICJC$\PT %6<-V9KTU-6++A%%X#5;F]"YOKM[I]V2I=H2[ 2H/2%[<6I!='2-
PCW< 9U$5XR2E?0H[!@:+V@Q ;;NKU?2[ "EBB<6KTM91(%BF5^S6)_'F_[>OBE<5
P!%@IH<>5]O0 ILJ6(0_&@D<(#^CAZBM,Z,TG+YI,L#EMJR1*G4')4P/_*>99:,!>
P1O<O;3445EDWU%9ZTY'OBTC O2M)__(9>JZ6/;JI/M^:RWKI^'CU4^#DP$5-SI3:
P9NL7!?DKZ%M6%!)=J5DY@/"0FO_'<6?Z.(+;N6>+K".\I RN'[U/Q#'F!\#954]C
PD-MQN7"P5ZB'8ZDMLUA"L8RB+I'9VZC '<MZ]QF,:3E[VHC6WM#CA7)O9I?<*W[D
P3JZ/8<&2:<SJ4U=G454E,ZY)WXVY3?B],"Z#;AW9-)Z$J)KIJHG0B, H5I9&N8M\
PR_?14K*)^AQ7F%07&%H#U2\H&F5_L(CV'&UU_NF6M0;_P*-DB@KH.,W4J*42WY=A
PMO46=XOD1D6!_2$1T\N-VR#6N%T!E7;:[NA'DA[N@V+\Z3=4_?DVJB&\/SC$!E^,
P#2-\P90[$@1RE&N$!IU[TCYEC @D2&HGE]4XQ</LOP?Z:P10[>M[6R[CL_]*'Y,U
PG21CJ2WBF/Q;LT0IY1RX(+3YQQX!#KG,VTLWP$,+/ ,S7@8B3GVSK?Q8U&_6O=A1
P?705ZRK,/JZ91L]8$Q.FPO@"T=:1U5HXMDD$$ !NWA)#RZ:%,Y-LNAKH4WM".N6$
PTO2>LCMD5R69/?,SD6"K1"=.Q9H42K*PEG.KIA(:S5)YSPL"1;1O:E*VM\1E9H'(
PIH+3)]Z8$]6G5[HY)JD;5-P.L4BS -O"M=/'7#"8W-<X)]WW@#: K06.('VA/M2_
PK-2 _.3TJEDJ8P[_WT?>=Q!TR^/A&^<\7BZH)[9KP<_ _@/NBEH>&^/(OG,/#B74
PE6$BDY!9:-4%K&P(\MUJ-Q57_S@)=OJP5ZK=%M<U/Y^\OA91X-/BQ9*%$7(C0U34
P>-GGQ.\W69Y*9_J#I=;J*AS4A-?*?&^6]]WN<O)#P=%K(E-3"E,L=[>)7?H((@=,
P[BV7XE9%& [?^S4E(KT3$<T.:A96EG!W9^G[.HOLZ2/VH(7K_%I5V#L0V=3HYRK^
P=ZW!OJ&>GNZ\*?'J=UCDY+#3KI^E<>S KMMOSZSGUQU.?YJ)N/UJGA4A,].^:J4I
P?N9V$X ">[=.#C^H\$>RT\LX)_E!$K]^\U J/WX#NA(R=+VW"$38;S"N6X):091-
P?>KW2BMM&YC%T_% '? 7[^G)?8B#P+5Y/177=SMKJS^="U;3+[_7"A[Z-79@)H*R
PQ]F<HI;7."Q(<H#KO0[(RZ[[%3'D5@.K4MTA-)-40(&X35.\,PY;%#NAIA%C$1^B
PV^%WN]./[N(1-V(VGPC!G$[)1^0^?4;H]8;$7'LTN>CE-JQTJW-$L4JF+DFS=R?%
PE-DV4H91M=8BR)J0/P&N(7"XW>[5;E"G\N=K+6 VZ1OYG[,_=R)JV25%+2RF-J\L
P"F5_:52J_JS  !"7"!\$WXY9V?./EZJ8D$!6@VD4+EX>$09>27++]P3FI'IO50%[
P&_,3-&/XU"CQ()8RA>S,N5@*Y)&C\:K=Q3*;:/GT'4RZ:B.0H7164L$5@_ $WTSS
PRAD#[Y%>*_>'XC@6 A596VX"05?@UW?-M01K"63?4!-T$_\GS'8=H,0K"]AV]1B/
POW>IK3!=%/P^@40=8K R+&5!HQP3:9\3Y]TZ:+89 !V1<^4;O4$]0C; ^HXWGQSR
P-IL6NIF[HL2<_KK;Q5LK+P:C86J^3IF=]4 JY#X"$KF&SC8%@_ ,XH74DO\SGF,%
PH49W!E]R<< (ZRYN[CASRVLM%< 0\ZA^)PTE\8V]<"Y^MU3^R#&0:_9[&H5M<P(;
POJP=4V8^VV6/,#=,KMB[YP5J2G3F#P>A!/=C'("3=O,=B?;]]L)L3 B9@AX(7>&\
PB8<3]J9\WUW7*9Z.DM82=8_6-Y?I/3H9%\7S/X1E@5Y-PNA'.*APGT4N+-@J:#ZY
P?38OTO=VP=P0N9GY8)F3^T@Q,. (VX[6Z0SRK1OUI;+<UT=TI0S_./&U@E'J5(Y?
PNT"[(*_Z>QMGIHN2'PR;0Z2%660Q%>7[8+;*/V"2?-M,.N3F6HYR=I(>=DR\"TO[
P_G3JV])N6 7D[OTZ/U+.F ?LQ77JJ4R:S<O=/3K8WJTTU883R.O8WFW,Q,PY/,OL
P !'&?)9K48KPASF>FY>_D),=/)JHVW+'VOI&5.OG)A_-/:!>W;11\R4M^(ICY@38
PZSFHQQ0;:?,:TMR.+O[F(_V4])?*;M-; $47ZU;0NL!SQ&L=(!:]TC(.^\RZA:HU
P]-RJ(&%.X@&.S,-GF%XZ]SZ<7/3H!%D6H0&$'VLO>E'GMUE>SQ1@9[948#C_L4JQ
P[3D-(YY+I7_W*1+A/0T,3VYA(U+8Y_&C3[<3WM,=7(II(==4L"Q\N,OD:3/PVA(8
PZJC_0(2;XA@DEY)![ 9OF_ NP]SQ)EE!%G]?+L[];Y0E'@?%L!:0F;;7V^Q_D*HX
P4:;:E12D>[F3>M0.8\JOK+5\YN[-]OW:A(;6^4&F1:<6:E*]][W+EG(^T_XX.9M#
PFO@WP!%.387.FM@XZ8W/ZZ?N7S[)V1;'D1<PXI,;ML9700MB<&Z3I' '#?!/@K!!
PZ%D^:%_MQP\3 TYQFD$COV,@.  ]'RL:M7D9\X4,T!M)3I-!3$>>C*EUW&\-R[1,
P3"[,BR\?*58N'R!$60?T'N]7TH"P6!3$=,,>K<05YS?07\CNW_")C_IVA$/HC=?/
P\;.#U:B+V*K%E)ITO,M&[3$3]$-($Y[]W;2)]+?^ASSYBR#;K,# P?1$UQ[XI)\$
P36.6:'000)/RS1MW^(&V2;@@!&H:G(./-#H+]K%4FK=-=R!B4ZFQF).3-K:_GLCF
PNK>5M.!@>\+FJI'_9+<9 ":W#*E71:Q)*#>&W;\\@ E *@]HI.?X@V\G!XP"TKS/
PP]W KB0\GY+C\2&$-DT:EQ%!IJ9MO2H&DZ9Y&HB[#K7@!;KPC)/%,Z,"NYMQ/8G0
PG7>GZ/Y<8JIX,M3Q%"B'JC]4D1%G7R'ES]:\85'G(L6[01-A;;AL[0&BI!I^VN#C
P%",2&Y3U!,6G=$*[D(RRZ\UV_5$J;2?P6^$ /QC%@[<7+WG3$O9]W,>G^@)D<GWL
PYB922H,87&PDPIRV;8Q'C8G*+P2WWPJY4$K/KS9<_)/\AQ]7D#DEVQ:/P.Q;E@[J
P'4GST(/^">MDNEU$3V^=_#>RR%-WV7DO$JY9D)>,P->3K)BRD8JO )DVLNSODR@J
P?5,*5QJ N<B[D)*E\HN>NM"3:SAW#S6AREEN)1K;E4.X"<<:J$B(! 9F2Z:@=R< 
P,!2-4KL.4V8<*#MPHT)KW'D665S/:#8\*X5Y.Y@6M"F!NZ.7.<D$"(&4'#::S92R
P_AAIFKO&!U]#OZK++O:!&:/IBCNL/CQNJ8#JFJHC&P/3T*&,]D\BH99D<GV'6[@4
PJJ 781=>E@<HX=.+)W(A+=LGPP(9A"1G?<0BRGDMM5>Q()T:<N0>P&>2 5'#B&2)
P$%?#=*M*&%=#DVR%LA[3%TD_U7KA]\X0WH3ZXXD..>JG;WR4Q/(;<//H;*/@#9W"
P+1-720QO34M=2S6T@H.R8^9#0^CR2_$B&19+DH( (I:V=P-2,.8"0_Z9VAN[O)]]
PLB+CH<U.$N @K,_"6$Y@A DJ/N+"V,KY+QVD$WFEQ-L\_+'SIULI@9[1#PS>[K3$
PX,L7#^:O*G&]Y/!AEO\,X\>:U'TX62<3 T1MGZ\S PX=-AWJGR'44\'PM!H!8MB"
P_520U32K^?B<PP89O,<573U(\]_)9G9O)AT+_.@X*NR]]N6I'*-H%2,UT@!<&7X#
PQ2V[N@R7FLP7U!=I8%F\U19!KXT'M.V%]6#YV1 H0R42_=OMGJ1[*\RRJZG1O08,
PVV-38$:(*L4\_! J2>Q!D=C!2&*V$]03B.E -@NBLX=] W5\B\,ZKZ-?)PC.I=<\
P8+OC<("CN"T+SV0.!$CT+KK43D&KUZFI#P.63HFOT'68.\JJ]LAK@U[2;3B*,+O)
P;51_B +CJ69_3OS55<IWK1E<$)>4;[5JXIJ9":@S\ E^$9/9/>-<F!HFY*FXP*Q1
P<4MT'Y&&1X"?*>@%'A,L> 8A85G\;Q4LS'PA763C2VY\@$EYP4[#V:F8;4QA\4\L
PJ$$ XR"58FW"/S<G48/ *&TK9[!Q"8P%X''CB+HN4FM8^.(GIW^AX499@O8^Q7WC
PSS"N2]Y-!G7X)!I]I^<IT1_S!K+4TDP^K!5-UT@2KE&(Y#3=\KWVK!UIM;K>XQ,^
P!%=+UB']0/A!.9&;1!V'Z<L4SE?P[AOA/=:(SAPW#@AGTH)"D-AA0M?&SJ&E461[
PC=N?O&=].T,E;F!4W _4[0UA3[79DQ9(GR9X?*G\''L]I4Z8&3"7RVKJ ?%[$ W_
PGRF(NS'"'ZD3(J<D-M^W &T&HW2^Z4[@M/067MC+P<:$KU1A_!)].'D_EA?J1KHJ
P6%A5KV09F<%%ZK^*[(H:? 1PY-4QJ&?2_+V<&#NN>WAC7JRDZF1E)1!P6I2$=\-G
PM#90(^L  @LFV)[8M;2,1II#%I<H+$CW*5+\+SN;8KD'<MY1"RM>#,Y" (SB]N?(
PK)3_7(]@/Z%2H$20VI+8=MQV>AJA$Z!,X0 Q^YPV21=KN65T.;PA/2,@R6[S'T3U
PN>]-HJ,4"_7UF1,6;MO.$,Q!O_@!6B3SXII=MMQ(E7EJ$85\UU9IYQ^5%,D'$0 /
P"SZ]U8$$HK'?^F:C(>C.)U9@%H',[*7W$YTWSKBO@&'2Y(.F 'PKT.<R\&FP$S?^
P51]=#C.QC YB0WC4<55?A[0FW%AS#WR6I"",%O0; ";XFJ,_6DA/QS:])M&KTKIX
P*3(%+QV,"_ ;&_L-!U.@;6'T.O096%MY(;YFLG?Z@5[(7-1?;S^(CO1G*'LS1I^H
P1@5;O)4G*W"U+.+Z>VL+60]V3G-2K&A[?:$/>TL :!'=]F?;<9J4W!@Y^'1] =^1
P^*FJAI@H#\_^,169^$(Z1U+]2R2]?<X=TVW#!'<B.\Y[C9"C5+0A;,-TK=4*$NOD
P?W:^QE5])7=I$ VP(]-%A&<=X$JQ*WFY%YE#%=N"5L=S^\6T;S;@_U(O%JS/!4ZA
P;KFH9*IL&8&6&Z?'FI.I3)ICW^[NS?K6Y[ONP6[D^-E5S@RZ7FH+OR!--.E8Q=.%
P)9BY!PBVMQ"&;\MLK,5=@T!S&S>EWS=<$QCS)L,:N+5)J,H_C-NJ+W_[^\RVH?40
P:'U;8-2MB>+(?V4,J"2WW_>V"RT80#Q>IDX%HKIBA2S1[>"EU5B'+)<+OP[A[Y%V
PI1OTE8"@.'IR9<0__EN RO^:#:_<8254)<H!)"-W1(6K.&M#$! U0_5Q>!>:C7T<
PM;YZJS"V.6["[+2.N^H[E4Y<RFGSO7$]<+153>+'/-JQZ5E&XT-6Q2S!MB!KBJPR
P;[LWYW-?Z#9QKO!9?#E4-BCI%GG\S,=^@>L1#]!]O: T3Q[K\\7S'4G<NP3AN^C5
P&5MX>+;.U2'9)/1OWI<[&&)I/?C4W6+:FLD?_"#:+Y$Q/">#R'VU@;2%@ON:GP(<
P7R(Q+9H]6)Y96<F%UV-3Z851W7YN/LDKNW5BJ*@#_2/$7[':E;*!Z3.',1754]B[
P[BF6^^UUQ2C^+/.JDZWQ8:34!0LZ3+AHW1?'[1Y(3+'T%R'V')7$&'46LB>L^;T=
P;=BFY-6&1#"T]T@4EXR$%ZZ/.C-^4O4:+FXV#%Z.LZ,I12TMAGB#V)&"-?X@@^DM
PK) #70B-#[ !()21TYQ!(SK=#$$VCZTPZ.8>XBL&;]29"@Z)[W2@($"DC%GH_-Q0
P!*%_OM,'Q>Z#M'!F!3X.LL+^",<TO@&+MZU-?Q"Y]CQ!]G(S;GB>"):-#8((>>SJ
P30^!["B>;'+K<)<Z0#CS4G57UUD 9906IMVR_B H(WCWACYQ?-FI._+@UF>L_H>B
PNL'XPUD3%)R27$W3@ >VZ=+EO901#*L9N?Y-+8TPH?QC2@1LV;OJ8@_/6Q"WJH/]
PW3_+,$/<)  /_K_1];G$9VYR\'/+D>9#LJGS9%%B>.]8?Z4J<AB05U7\J-_E'L@%
P >ZA)_8OM3F,GL"+&/2#/RK2T+;VU=TH9GUR+\:#ME(C][?P/T'.FEM  Y%63#@R
PX2_=1DIT15Q(5;]KZ=T0&8BBJ?IA@Z-,Z4BPV[GU1O+GILIFF/XQ)CB[5^EN;0(&
PKF(6F&XJAI<A&DXIW-[AN@?WP-=+31=\Q,9#"A!AQA-$B1.UB_OZ,&.Z\).37TXV
PO<&L,4DXT*,B+@UM(P&!64J^JUU]_> D?$RD0;5)D&Z])B/. 1-JBS6H?KB?J5!P
PD*OEB^BI$4N?BC4QN];4ZD146"<77ZK@LJ[6F\K>X. KX/6ZD(HH9@G_O_"UZ@0"
PFR@TR2^>59JX<@LV*T@BL[*HM3RG#.N670M8%OZ0W7B$UFO74^/[/PU95!4 @JX#
PWL$EF9WKY7?G1L+6 PJ"D(W=?:^92[3#D) X2:I70.3PGM^5M_I1ZKP0MZ-ND.Q#
P'YDSZ(6&KOE8?W'O#0#_IAMI[_++@*<E\3)_2N 0]ZFHAO;5HQ;'&FS)[76>49T[
PCTKH7[G&;>FT[IOITCSOX[ULG6XS%Q-^4BL@M D6;-#3H]6 E#]7XA(2)#N<MSX\
P09]Q>&5/8/EKG)IQH_X\.XW>K1@*5EXS#SFY^_I;2"T%O*'.L&9.M^ _D;@BK[GR
P*&6?R(XGQ63%7%!Q%AZX'PH].M%E2K]Q!&;;#0^47HC1YQP-CJ"2YUQ&"IQ:5IX+
P<\?B\//&N%FPTWAD5W+1QBMJ@ '9P>JH,)[)852J"\%OQD4C? !!2FE[^>8/_,KZ
PY_/97H-"6*D4&DO 5ZKPE8W-=M4T.V5B,+:(^SJLC3@,&<A_+\WFU>5?&Q(NWZS2
P:@JC;\9_(:\(VL5UL[OKYT537JL,I7F#X&\,YW)+'WN)H>M;:!6G&U=VM-P,-OL>
P&=TR-NOY.M:V!Q\53,OLU@%A7YVAY5+,R!J(+%*C!=Q&JYAUU)YX&]_3UEF%_@Z2
P"IDKJ?"905OI;'E7VRJL90R:/HT89NT=(G.!#Z7&#_SE3O'XIN#6+OL3C!C;D8K3
PES3[QQP<EQD-#E^RA)EH6*P)%_T+VJD]-J:^XHHG*$D"^W1 [4C&J.24+LC4JT8%
P2E#QVE@9+^2#Y" OQ#>M'V6Y\P:6\JF#8U#G?2ME9TJR@JP6L^'XLP#[6I4_H&(R
P6)))ESC/[XOK*XJZB!6H;)&8"8M.5<L=A5&]!O;8-;(^MUJR:N%$LBW&NW5$6ADV
PY#T>E<<U3CJ% WI%@5O!H4S#NV4=5:]0C_Z@/4[OI#J,4%EZ'FZMM+D%0^@=H2#3
P?;F)C&V(H\U\@M[Q0XPWSY$*BIS>=XD81-;7/T1Z<L<C7BBGJRC\OH^T_$N<M0.H
P\06TYAIH^-S(39]Z9:(\8C3\*'8:'MSYZ++(C9#84H&[Z#%N.)EW"3O6-6O"IY2D
P:_6-K@*96TZ GMYX7"_ZA_REF-'4BD_A7&@S'H]@!;R\I-+6U99V%9'_2,Z&D2%E
PE<HO>JM)+F_P*0/@:L&5ZJ18<$)=1AYE55J$I66OIDV"S6E7E*G5.ZT_^_3R-J,+
P!XP0,$R4J2]!AQGGL?XR(>UF.S8&NIW@:XD3Q!D%"QV1WH6?;8^.IWC&[2RA:<C6
PD;.ZR>>XZ,MI9G+%$I'9H6."=<KJU@A1!Q?:&I_ZQ7&/MA*PF;VL!9&ZN!14Z_-V
PB5Z/.W=<61@PH;?K)ZWT(-=T!;YJXK?T) G-:?+-/H%S8_&?GBEX&Q91JRK5[;,7
PUC ?0)*E/K-_=P/"<)[*PA]<%Y%TL=*2&L6%?(SND.--D$ONS__C2-I(=FSLSM<V
P^H"N$9G8WS8C6.D+^T(K;8@<BK#UL&P2P@']VE::7>R<N#?"70=P4/SDYX@,IV&I
P[\"B(-HWY3&NU)[-<;J."?LG"4+.?&\''7$F>Z2.I]L3IU"&SSB>8=R;O]Y!G=4$
PY\2F3ZS6])CH"?8;C7G:EI[KI,NY?,B;88^=&Z2J<VH1G#=6&6!"(C6$0KMS4[1$
P?=%Q0*#,/?32\A)+=^?-:W0O?U2"<D'J(E5V=CD 2'#3&"6*Q.%KNO-O[?X Q'K 
P?7KQ1JZ'##.YE_NM??7*\+"UU\1]@FXO'7/BYC\:>:V^H4<9D[6!*]V 6YX%!%Y!
PPNC^I88+D@UK;>H2TM'E_F[=>VTS.2V!Y :GS 34HW5U/GK#'!XA4.!%P!-QO_]4
P"4F!_$DG)_NQ?"[GMGP:"3>(9FVLK2:G.&[1>":6-LO5;(''SMYR975%D\ICA>X+
P%;4,28+#/@!WN]! K^6B1EOW0HC.-D))-M;.9>9(Z3Z6?J1%ERGHTB^I'Q-(,$[M
P+T'VE/C[K,1K+DH3#.1:"I&_PQ7:GU%H",R94M<U RPSI25JJQVPA[[7VB,&L/OB
PA,;R;+284/H>0?]K?,W_*[6MR7/PC]A!\/\DA!5^_5@;<PNZAAH)OD,=C8 .XMXY
PW<YXO,=:0W*FJ5O#-:4/M[!7MP#'>DV(5.LK%@/!CY #L\5S[41R)MZ3=6H"<-W(
P-[Q0DVY0VQM\Y4BO:O=Y1CY-'Q_0"(Z]@%=!V=_+_6]1J=0:5H&&6;]=XW78V@K]
PQ#)UE7 [%O_\.HOBL I.9;7B;K.PAZ<$GYVH8 *H<B!4M!:5UU>J<'@89W-5',F6
P)_-&B5/:X@>]12Q/6'SN=QSMHKU1<9ME?78^5I8ODI(X"6CMI8J[>%+^&9S:>+%E
P6/]&.0B*[>N.P'ASFNM.P0+'RE&'2^@Y9OAEK\*M?5]M0QYADS3=/KJ:&J[R+0)<
PV./J2%\YCXEU;OW.<B"6\9H54\@H"2YHT&7\4#]K\2AB/JFT07\)(LOG&';4M]N%
PSVCQ2>.SY^E8E!9V_ZQ+CP8M*TL1C#(&7\J7HK_K'LB+/X@2-V2(MN/7L"AFJU?:
PZ5Q($;UP=N(L$+K]OD)Y)->C(HX)E>L*MW![W'Z^*@U[!J\SLF+TGS3^1NL^<@^5
P<,]QJ.B2^^NRBKVU*K\D)=8%Z3.*I1;[<!%[[CU[@Y_$.X(AB+)8UX^^\HZO@=[/
P[KK&+3)I'E[9HVEYC32-NO_TA-D%;8@ XV_$(Y:Y9/U@H4Z#GC? A2#H,A.1U.G[
PIH>V=Z%^(L(?I_O,!5%E5(<3.0T$?R\#!^::D0VW(S9OPJ9I2C=A4X\TF=+V>+3/
PP!8,%:\+34]7D]JVY;?:#RR\?W6IZBMG=P9"_ET7H&J#]S)T7;PVMMN2)+K S$E[
PG"UPM'P.O%M(>GPA3B&_G+,%7,4D';,$Y=(%#;(Q.&"P)[JEB5:D1&L".3A:U%3+
PW,=]<:Z*67(H!=7Q.PBS^SU;$B5<Z:#2"L<F**)J++[;QFY'>A;NO=[%M+)U!FOJ
P\S!9OMD"#YG"I49:@!IZRL+08P,X6?EO^'2V^,AT?.$U. $-@> _:XV\+. *OU+#
P"V3[L@(S#$\(M36X7&]YZ_VR2&%ORX%PN&2BH^V:1\].HL.ETC=(Y5KN;[_2'2SH
P40%?*<0:BC[PD[>$P_;LSQ+]T'_#:I9>K\1JOI2S,\A/!_V<JA2:2Y&$:EY04_F&
PQZ2"%9JRPF.MC2(70=C5@__\RPCU)G.\L*.!A^2.SJ-J6U[:(:\6^YA_S+2X:JFH
P,$7VIB6DBH =7([CLMP&)O8*#[V26\Y%-^E1>01H>[U1Q &AXNJ>PK#W+$/>53^U
PIL38_V,H8HTV_4 Y*9DS7NN*;C9Q^&&&K4'0PUWM&Q6S*3H7N=.A I&N#O(/,'M6
PT UEUARSZZ!KQ:.8+'[4^^(>RLO2:1Z9CAP;TKQT"Q!_\;I2>*>D@,]K"01H%OSC
P1JSL5\3=Y[2GSU.;RLJYP\JX@[T9^^:EEAVRS<SB@7L<1</[]V-&<6VXO5_<TN[.
P0RV"(&J92"LB)'U&*D==!E2%#[V/4=I.C:^]\L^_1NEW3O-]RRH;#CKLLGWYS_90
PFPS[PC%V@L'4K*XH4!R#+(.!585,.];/ @N&D DZ0#21CBI2*PMEA!\A[M3+L:?K
P)B/G( 4;%(&D7/54*)?6M]O ;!W7KQI\PC>@"HI<?_'P'V,YVUX@!^:TXMU#A2BA
P#/XFVIBU&-Z15NCE(,(P% #"6Q>H-=^KIQUKX5^IAJUNO.KEK1AO*E''<%:X&W%B
P-WM(,Z7&H#B_BZMY%"%LQ->?+&BK)O0M$.*7@9XJRV:TYJ5SE,4Z#4I(&DHG&]Q;
P!R1+Y;L)D\%T'/U F!QX4LS^E]3*9HJH$@VB"45%;_[]9Z'OENHCY%/][^Q/('I@
P9V^Q.^8P\TI7YEFC(5O%Q@."9 %(>AXX/1M]N*'$ R?21RG4-#^DUGQS 9 OQ#ZW
P71OX\%!.1OD[4Z#FA"TH:N6VZIXAE?46MGI<T.?C.?H5#+J)KK??LMZRHGU$D0#@
P?CF8OW$KQ=F2]\Y?5C043!]AM=<Q//0ME$(ZYZBW!X0D>]8_N4K_JL]0MYQP[D30
P S4SP OQM4-.<0'$3Z3XC>-?%_74H@6(K-M= *@ORIAA*"VWV4W&:Z=U@U8-(LD4
P.66RPH^)?*U> [)=-!T^5KG"/=OZ!0QQVVUB+KT#+ODR0I]9VW@V=(P]022ATD<\
P@@H@G\>J9ZCK#1G5L.L<*/GP I*2/;'7-%*2;'T+[MLH-Q"7FTGOHH*X%N"QOH)!
PA>LM#: S$8<<O &K:AI??;&P_C3];ZECM+@>BDVE]7BM0^G<OS3]XQ7UH8I8WQVZ
PDU?FD;%48W-D#IK%?ZG5;5 YD:*1:?EL6S"VZS&W2<"']%V8)'B$OQ2XA+$FX7#Z
P4!]=)\A<*$WGE5RV#>-+>VLC1Y5@6TRP7^K78DS'* X*/,.F05'@,SF^Y@56[1=S
P^4,DE@G?<@D)Y"VX:7GT"TQ/T!Q$_@\"0$I.C3K9*1]Y<JK /HC-I(3,D?I^^;#V
P&,WV"9#?3_I3L!UX/M43/W80H*MU/^D#PA6=YHA3%00@_"6R^(V)Q_BJNV6*A$8;
P1)$:+8=8$-?&,8,6:H#Z]_GC5QQ.L+>IQ.\$#"J)D?68C:]>.>RG9*0,O4>.8RN(
P<XC.([8\D!LWMJ5ZZTPW=I%@"8%OW9_$>-> ]\V)-SF?J/9>AU47Z%1.^%*4@!:<
P$A#[&4."N>X(:R!\)K2W%2FD/R@CUE,AP.["]]NFVD.K(V'F-_T!9;FXZ+4IE11\
P)JJM<KW1-\\5D2?9'/R)M1M?[-#2*_-4>0E)34:Z>4%:M#(YDL!A#CJDKH>_05VB
PPX<H[;GQKZ</P^IO%,<@L*N8F\JBYP/PKT8"N;%[M:=:+??;.7[@H:(LD*F"<K\3
P6I-^G#TYGGG(S_5^>=*:/E+MN^_Q/LD6I@B19)F( B_+Q7HL[?/S W>E1LSUE )V
PDP:<ZRA;G*2A#+(" DKZ R&Q26MH"P7CS9C;?+S<6^G&'G2C;*UM0TNO@'4)&(2S
POD-_$.VVW]5$09"Q'(UG:N[NIPANJ@&>J$%GK76\)MWDM 0UFZBA\!UAH7@"[5)>
P*G*C"6^ :!VMY'K7 U60FWY0G[_56C9J/86P6_O5H[ <PT;QG5J63JE;T#%6Z3]J
P)*5>[+JGLTW_D%JV(-=:5;V7GJQ@VPA,.F%R'B_9P1)Y/C0SPD3.:?]S*<\KL\^*
PN#-XW;&@;?1_;))SK@\\):R$Q%[K.@Q=N?]CC]FR4#Z?F#.5%F[NMJIB^&+J=);]
PCHPTC:"L[MERW3N,6.!FV7<%Z[8)UE^86HH$5?!Q-N)4>8\+WFP6,^BUH;;_>7J6
PD3J$ $S-9UT-+;9Y<AM'(6 (7*/'PYGJJ_F[><7RC%Q:=O8-<K2OWPS#4W#;[=(^
PRQWD&0?7_<?$V/06,F=D30@M;9F2R4]5'7&L%GI_'_VWC9YR+R*L*'O<]4I.@G*Z
P?78UXR<+A9O 0T\,JI!(O2LE>V/29DZ4IU40&\*@EHL"UJ&\ULI9:;VX17+_+0T7
PP"&#D^\Q;.E8#34KL(G7]^H'\L4#-F7?Q-I9^>VCE;[H+_R(H7=;G7/(M*;G_P8U
PO-M?_ 5_WH\F,A1;= N9!H>!,O1+5 &I=Z_94K83551TMI^K+9@VVD_LJ*F^3LQ+
P'_C1SM@6*$#!NO>G)RJ3HYQ5!HHVC]6.)$(4>*^0-4YGXF)2H]%9DU?WY:%58@9=
P(! ]]^$ Z4BED:R/!#PF;E9'&K\;@\] 48A!$W6*%/>QYI[I1UAB$R#-<()O3NN+
P)'Z'0T<7\-(,374?) P^GR!4#)/PX)U7,"::5VES$-'L8TW0>[XPJV 5W4$N1$SD
P#:-%NL&\DI*#"+L!*8ZW,;UU!^1 <798YKWV5W9G$HI=?MO ;'EY!.AUK$?RKGU0
PL&F<F)R@/*[P[4!W^%YW7S3QGG!P0J(S3OER,!LM72J.M0+K.=#IN(5YW-FJQ7KZ
PI;[GF:@00Q8!:H7%<3Z+"0O<SV]OT/Y_J)&=3!)H)W3@D759/M-.FCD 1H'EI5W?
P(.4W=P7EZ.(!"Y8V>[_:-T[:4_EOU-.!BQ0G0+]T/OFVNS*#FNSIW%<9C]'Q>&QX
PF6ER#]:JWZ.KF+,T=QN0=0KZ_Q5X.A46N\:O)]J=/.__CL1Z(Y#*6)Z7@*/Z6;UF
PB%,Q4%5+/CL70I+YK6\@4VP%^/\21?Z8E@5!<A,3DUF4@]M.P1M2\X"VO?;5SEBD
P'LQQ4#%?%_TN+16111M=C6&>3*?D-Y(C^NWXX:M&\MJ(G^=?*V=/R5.81LE=;K.C
P+H_1/<"KQ:MA=RA]Q,0_..4JS\WPGE^K"XD16!?5=V ",?-]_YRGFA)*GW;N-?NI
P-0,RU]A'TBKD*KF!R Y,;9E:L57LY:K>_%^=%/(73TG#LF"\2"?JL4T)>OOMV;)/
P@\6W/L!,M:ZW%O[X?[U.OW%6<]*\"Z9#"10G)DLF*I]:]OSD')C]?].Z?M<4PO9U
P3"^5/'32  P:/X9_=:WFDFG"Z)5*,A)9Z1@.@W,II1&6+8-\-=@;E%&^<=1$7P#9
P7;'%A.'F556%!X[Z(^^\<N X,MSJE2IU-L+8)**C$P758P@A]$&3OP;-22<[Z^>C
P*R0EI#90][ZC_3?1)+[)\^X;"0=E E:LYE9_E@TF9<-J15/)L8E^"DQ2A>K6Q=KK
P#8@5%,^LQ:-[/+#>-WX*A"W^#/"!V[BH=9% .,$C_7"^#EUKD#/"577V:%IXD:#^
P=9'-=TY2BTOMB/&[!SVT&"JF$C*Y'P? =0K ,W-7WBA$7\R0YELC4'RH_4G\3[+H
P!4%]+&8-<6W$[_1?Q&3):XC(S2N_V^Q E(@8@Y>BH]5L3P FRB*UWJI6MX+_ZE'Z
PA\CSI-+0M&.?-/Y".7*]!>I"Q2_Q4()P99P9F8L5!4]%L4CMVK,OKFAIQ1V8@HB%
P?E4S$<;D>UYVJ45UMS?D(F\)TR%,]!./+:<)RF'Z9VE7# GP[&>-&CGPR)X9)M3+
P1A-S!AY=:FC*WQIA?4$*KO9T)<G>ZFYCKK4U"5,UO5;R\_T&!2"\\_AHX!?WPM)-
P68.P(ZAG": SSUY$ ;:2'T'YPEE>%49D:0*L%D G]SI((7J8B0,AV8Z*6@W\AG=8
P/UC6JVG$8?[+,3N!QJ-2 DX)68&)*J^,_G*C/.G<9%B1R,Y?O 2!I,@@T*F5N<&]
PZ:RHV$Z<6(+*43:KT*!BO@Z%T$@EA,&O]P2GV;_X[KH]GCXDJK;$EFYDA0;MW$"I
P67<QKLN^7#TRKZ,*384&3T_;CI:6-^_DS$3HUML5Z3;_GP\17V_C*_>N=M%L\-/E
P8;%6<)<2"+ G4LN.4='..M8O8(B.J!91>P&KO<GS.F7IT@[NY0P]XQ@CSY)F$RLS
P_#P9 UB!<#)S0I2D10<Y;"B^;8_CI.O88DVP [=7&$YLI=#*T&1%+TZI0J(>H7BJ
P%,-%X$;R[=WX45&2O.90Z^6.41]C$KG? ]<I=1SV<T2I45=S8O&,QL@ O,UXJ'%%
P%F(K4V>]> L1F(Q]%&R1#*T!P@W&:5-N*OV[3+Z/V'0N[.'^LMFY=X6I"R[7!.IC
P#%Y!J>\$)Y]O7?QHQT/;KA^Q$)GH-*Q/N&)#4ZG18SNI&=$KA6:"^V$*NXJS$-<E
P&^'PSTCA[A5&#R0C8N"YW#-#]:)]$N"597H_,L^,?VUC=*LJ>9@'#4JF<W"F2MP!
PE4P=S:[%XMUM#F:&.(#2VS3($*]VB_5V940,HQHK,"56)#=.L9XNJYVGBO]-*B2/
PR[M_(NK'-227_/'J=R?*3H_N4_P1%F:+WE@3M(;^'YVU+%\SLR]+(!WX-)FY8J5^
PN(DZDLF=N1[8BR=GTN&<]7+=;0/"-+'MK&J""L9=>HEDA<XK%*J68)?FG1>1!K0H
P;IM+,[CL8%'!8FGH9.2VA$K^?=22D]5'4:#DQL,:7JRH(ZL:6/7;CEWHSKC]Q=4%
PRR?!(,A?4CZW& 4WV'!_E30;A-S@JE77XP66U(56&B>_X?H'@!5O/4"<_I>ED6W6
PU2>ZUS@KC_L'9+LG%"T)S-M#>Y;'79&B;4)E7G:8%FW(+[AY-^'6EEA<+$Y?I">D
P "KUO>&@N8R=/=@Q-CL:WS[P![X=5S=*!=!$V(LU .DP<^H5X_F.S[8&D,ZWL;@J
PSNOP2C ,2NZDCS5\QQEZ*^VU#R(3B^8> 8(=F,_K5HSW]86U_&V]O@P*%G]@Q4:-
P/LS22EJJ@@/A5RUJ!!2M2\P_"60K_A L/9;1[:V+*="'ODYW$F[BR=QIN=Q3P8V5
PKEC\"(36EQ++*FI\L6GL)Q2SN[ 2Z5D-Z @B5Y3J>9$Z];IS2+F/'H.E:BR6N,ZD
PAK@M=T%G",3 4>2:F[*XI88D/I6I!GS+K^(&U# %H5H5@WJHXW#U/S'4D223$.G^
PJG %#_!F3 X498F_-BC8#8QQH_.%5MPE;(XW_;@92&@[_@ <GTGZUD@?0;; G<BG
P<00KZJO[@;(=$],=%/_,E98K(7"?F2/^&/,) =LDP+:!A0?/ <IA=RW\^ "Z">+O
PQ!Z6+U12'>U<VFH]BSU3;"F_D)/+OLZ;Z5&YJ@*$<M5[;S EO%W=J_]38V5W0*"U
PV.?(62APR?,L@<K>7WNNW^')[ "$SL;/R=2>&:;*RJ_)I'&GU<?=-**;Q)=>.-?O
PIZX(UZ+!9>;L'(=\##*?WYN;C[$ .R&\6A:N1(LT'A/2S*'FQ)B)R1R#J\CO@P90
PWK<;:XPP(:1_N-OLJ5]ZZ4E&M0_</5X<Z93I]#EQJO9WN*\]#S#D9WCD^6XF%MV)
P_$KQ(KHZ]YR%SK\8=TH>ZA QOX!X+P.^C_WPLAM*_+^@KN-)[*S2 FZ"%!2"@1_>
P*TKBQ@"R),NFH;TK2XA.!17[.:AMLL [B^QO693&;'H6PQ;QM"8]C]CJ"?XW_4A\
PBKH>DBEK-'+A[]QW;28&7)5[X--A0K[:9Z]V)M^;-!K4OFH,VXH>M\>J2)KJ89;A
P&J2EAH+G/==C4U;D&3K50T;^1^(6R'0-%\2?3&A)=<(MZET.A=IF&X,&EX'.*'V5
P3$KA^+X1_6&;H[#7:*X.IK@IZ",V!LLVV-;R*C@FUKVPY83EB@,(E?\A6F<48(&$
P$WF-M%1PAOL'0Q-1M*1[8\,L*')&OB>[QK;:@ U;.W<9[\;M"0-]P+=E!)F.!;D1
P 02'Q.N+TR%8;XTTY3WX"7$C=N8!';9EOL/(!A1PR>92+7_1: 3!/:#&D8B;VA9P
P[0MQ"_OQK_^+O)&,*2^E<T8%4O@@R_ *^80N*MJ&V Y4IS=07&592P%YDA&YPNC*
P-"1F!A]]<&F;!1I2Y9H"[RZ[=H61KMDR6N7+J&!+QKV,L?"6*R/>8J"196"T!Z*"
P>*%1@O\2RVE% >K/QL*[3B&YO3AC\:@'#+IMP!8>A+-5E).! GNR9T)N!><K/AX2
PHVC$EVZ[Z>*-><C+&R>5/[Z.K1V%\\&Y^C*' U \[78F)P\#"<EP8>LXD97/DCNE
P)J')7IP"UP:SC.AP#Q]I"$/1W5U]<&E >AP1;A?-6G#.0Z$4,5U)N3K:SVBRZGX,
P(0U+A9U MCI%G^FAR0FOYEK3_S$&-L+&7K3B$&Q$"Z#>%LF6:H*NS[0NJ\JFC()/
P8P0/K*\MO];B]M*Q-@2M^!KZL9(:'3J&1L#\!C_49RMPO2&^+D-F8T-:>"8&7/SY
P3'J/1/:SBMM7%3$-WUP@E%-B6$ @@K+5O9^DN+_>SZ(%0:6T6\0CS#YM7=O#P0E$
P7@WSRV!-0;O\NC4<:&2RDPIA=3.H3E!F39M1X/EH,F.>1CM"=I]DK55B,.-^B<[M
PHN9O^[>!M^*RQE&@\9S<&JJ789*''3L]HWCK?QYT-SYV[")% >\;,"0;P$>[32\6
PY&7IW.!@ (=BQ*:9,4%>:3>J3:&[L0:#.V[;2?>P<JEP#=6NR3EZ^BW_R0=U'5V!
PB#6HF5@);S)ZZ; C>WE%/E-]-031-I-_UPA_0=)_BG[\W,]S%Y;OZKSD@*7J2/;7
P'<Q'6FXQRG%Q9ETJR/"?\]U<,NN4ER\'G)$WIDD=1HYM#2- ]4G\^IVMY(GE)"@^
P]/$\KJ;4&0%([MHJ7Q/0#DHP$;&?(_FHHKP(G5(;57V?G?^9OL,>1VIX> %K#:2B
P(>+JO$#X?8*[6@!*:3M8SL,!@%5P3T [8P[?-P0$I,<U(EAOU*8+@T@QLO!SP7>S
P1\+QW=!XKOE]BB"!5%&.S/@78B?+Z'CE1./,I\ 4XSK$W_=91G/F UJ(_1Z^'?7J
P,1E](F"T$UB;5H$9UOATMM:SM7 ^\ #R^7B\S1LX4M/+\C&ES\KV)?U?V8"""--"
P##CJP()X6_\C('3S B.-PIY]OT!<*'+-0:?:[!KMH*D!\O"33 T!&;.1=<1XZ8GM
P=JPND*=&]2RCCLUC4,(R+)SBJHW._5\\?:&UCPQ5-5B]>N1X05-B+\B@EXR;(T:B
PYE3]UNB#^E;L5]UC.11"SJ<T7=S?"!]6]F:M6!;!P2":@4/!-%5I[>V9'<MFXLX"
P,2/9GAD09=)H=[R9JJNBLFXXI>,-BHF+;U83UB.1V9[N3150?)K,WJRJ2-_;B\GZ
P <)FF?P"DLU3:FNU;$#<&"\9CVB&:>A]_&_0A!2_?J.1)H&9'[&,$^Z@H9(@OO=L
P90:_3(&)UVZB4]W;;U5^JQ_@!CI/;&7"RGW)=I[J1B 4!BMD='?_283MJC:Z-TT7
P%)0"="1Y@TO^:,AG!CM+6#MENYI=OIJ7S_1SX;^166>E!ER1\B[K!8D[C^R('B75
P(><*-SRI5$7+\;0/ =ZQ^BKELO1]>,5?,@EJJ^20XJA8KA7W9+VI^\R-S#@@M PO
PR]@BJ'C&N_$1$T9H37;7KT;+%,-XO4/31%/#F$KS]P:]@)H),9&T^-# =[$BP%=Z
P^AA)Y+,@HF,"6Q'"I -#7F/*<":-E0XF0QN[:AO1:C"NE!9^IE<UOH??4>7H,XV<
PO;\?C';ST]N;,M$W"@=1=_-:;MEZ$R"]J)0J.F])<'@'SJ+U)[ZW^X;%"!R=!*6E
P(]N^QV4<7;4XW"SU=N;CO0\QN$1%"P&<8\ZL"S.2>SU<9()9J3T6XI]")H!$140L
P*K.NA42O?(!B+_L#H68!/-NG;I%F^RI)!?^=)^'4&WQI8]%<L[6BXFVJEW@N(8XC
P_D\U?/^4@>'D5W.[TX=<266QR5I[F60VN1VVHYC*G%'E"A*-+F0NFE&LSWQ6UVD)
P P;OD;+PM<]+9(B#_ TQ=("$XTUU&&7H:2] ?7SD_3 1/]8!MN>$3>1ML^:\[(4&
P^H]ID#+>=36P9<DE$<WXWJL]-3@O,8>*!T<:.THS"RRC3<'<2SGZT)E1T-[L>#HK
PUR/?=W3*-0:J#AQQ&+M%N/O1I8/N:@SD-N5JQI@DV/%6Y2,QZJ<K=1DRLUU]^:."
PL!!*^Z$_=&2J")R"MQT[B+JV@!0/]5P2,F/O<;_J29?Q9G*^W+^A"H.%G9G9!>Y"
P0;C-F2HQ$PIY<6X\5<H7S^_F>QV)<V+7SGN.$KTYU2#E+K;3"%]C5+D[?[L!7]'N
PNP$ %R]5*<DU!TTR_=K$98NA&##RW: 9$^?H[G50!?N+S.^FN&.]MTK]5 _.L1'^
PMMWWTW_[F7$0]0+V E)U6<WDGVT -^TK^)3$4V?8Q)8=X.'.CN)OWQK)5> CS*ED
P; G#MK==_7'6A3$AP!EGC3LV@&+F&W@DIYS$GKX1KWN5B@^IB%=Y%1S\#^E8HDUU
P22/M'*]X^85/9:,5[4V,@LK+2;02U%U@/UVN=UH?1*(A^*L$BK(S:%F-##D5:)"[
PMR*HGLU*O./H &$<ADG'>,[(*4?W<"7\]1>"9<[&.=W%S'&^2]U]L0)QO2VI-;8"
PD]AL P_C.(*\E,QGO,>ZVF-V'[SC2B_S7I2?IN)RV&'A>U+$TC#[' ZZ/)ZOR,-4
PW5\I?1!CNK)@?UN/*[C/T7N<^&D* WKYR/-R] "<QS%)CR@&LQYR4NL2;>>*H--N
PQ;D/6K^2L*YS:T?N-[^!I( (Q73W$.58BJHO=X4UC(U0AA_QCR((E'H@FIO^0^HR
PQ%[!"4N_'"#]T..FAV)L^]A"@?TKHXS@0%R<5^TL#7D6;A#VH9A/D#I6 .F@I.*>
PBC/J[B*.'J7^[;VX+*7%02S?^GM6+DL$G-7@9P-FQ VB3;_];U/>\RC \JL)D!<#
P4P=WG5N@[64)YO^KC+ P:.8ZH7G@7?[,!AEN&0A=L5,7#E;^FF68WCY!3K^/RY20
PBUTGKWD-D*!Y\]J%W_SR9$(+5 97B]0P,VEAV!(&)\4'#\NJR1/:/9GWEJTC<SS.
P(>("SMN5]<X?DM3KEQN2 S0C_?E45K7HC]*N+ZN=+K1HK]FAC=(@K4'300HHF"%1
P\&WBE.^WMP4X$1K/(H.%AM_+-J.5K4NC6*V,+B<\,8@BX-?,Y+4# W4VNE/2M;4W
P LX[ ^,PV$O6K/\B%MI3_G+3NGL6%:K","6GV[RZA7% LS=0)[&:0VN#PYZ4A;SX
P><<%5\U@#";UJ$2!8FIH?_MGS%'K!M8P].GX#)0+> 5U18BS""5OCVM/="T/?.K7
P#?@B/[2*55Y+L:]#;C]N'H[I.8^KX#7G%8 \3#Z/<L(9/$;0DMT=(8W"UDQK#C@,
PB=WDTOJLX)%3>:)FAB?%N@%)>>NX67[(D^]7"P.#IGO[*YC'9.W@QV3)2&'=&Z%_
P);:1S+]\K^2F\GVF(]SA?147 )WA[^'6-UURX*2LBBLA7I4XW"@8Q;5JR"1%M8[<
PDZ51;*I<U0+5E_A'9#(5'+>#@56-T1D[6<5I=:8/G?$.D9!S*B]6BY8:A_U7"64Z
PH#E)_C,^7^7;AE\P?OSKJ9(PB2<UB_M],!(-22/=F#9IZI9^BI4$,X!3"^J-L]LX
P8Q<7Q=NI^5((6OE"WZCM ]GP9IN--CL=OO;\/NR6:GGDXYGL@/%$V$7 $P*?G /N
P(A<O"R'-R%87,0\Z3I >>L' WY#O1BUW#WGO%!W]_]/_$-/M>^$.F\"RX/].2LY%
PBD0+TA9'U2GSI$P,')]),0?7.TG-2=&CG[:L#Z1T:4@MK%41%C.\]1Y9SCJ51^M#
PM.UH?:A8I&=>/45/6=;@OEXQ!Y2W?*J-$X;'Z3PI]# U?XP%MS]/*40NL\TO4KRC
P!TE.B<,GHG@7OVN@"%AHX:?M(;=8BCWR7Q'>A%>2C$;5[3[N?UID2,/3S,,G0CA'
P8*Y45GL21*F(S("T@7J3+_D 9#EW*4<Z'QHG>"'MZ9P2TD25&SLDGP^ASH/[4\Y!
P#R!AKN@R< %$^'L3F3&3MUT:V F!!T5WW+R9+[*&PB3-(K03&IHF+93:YB=66RFU
P3/7[M"39G>0+JK]GE91!=5 ()M)O,^\KO=0HK7:CXJ=RQ2(#RTT.3,#$GGV(7@^[
PC:UN^.M.N\(N']736!Q+B*L1+OW"+WH4S"L#ZFX0XLEPL",1<J;P5>R#9B[^["+]
PA-\?(.; V_EI/B_2XX2S7GC>N,8YRI6)1QXOI9DM(B"Q"B-V4=GMAJ"4>,:,+@W\
P5^*[9$^]KG4YU'.2AZ>O,;W<>N$I+4O4YT+1,2DD+GAG?U4WB">HOLN.#[S6(+V\
P>)%:(B0$  1HP1?_X;19FN5M>>#]$+B1?"9^>7,T#XZ.XP9P(U4V>)A,?YLQ:TUG
P (L)((B1_<22;JUPF%_>0FYH#04:_PV/&HAKZW<2?C^LF!X*QY>GFSM1(5MDGQ@P
P*<S@A58U;[1!C1C-:65N"O30>?_I!]*IO!KQZSCDA;\I;?L4H4*IBPDE;^@+X9X]
P<"Z\,UN:2RJ>1Z.7TD#=YC172V*P>%I%'6JPAVEP^)NEW"/1<T!^FIM(O1D,-0;>
P%?#BE%O 1E_Y9IXT0*>NR$7J3XI:^IE5QM =[?&5AE!5XNFOV<94QS-A:,**P'F!
P#Y-E'+"AM5G%HP=UK84_D3V@R9\?O)QZZHQC==U3'>C:JKE/Q0:F>+^1\6FI.T^:
P$@$'SAD .UI##AU[5;$YY7G"V)V;3N14Y1R);<MENK!M;A?]Z P 3+ ?^.;$J"56
P9<;8N%<2$U3^2+]$7"2$FBZD?D97*;W''*D8A]^*^G HAI5R&JU;>&,Y07IE:M[N
P+J<09$8U3C%BF6=S%O?;C"TM1<!AQD&%T^;%6#"GG V4J$7]\SR^(ZLM)WTC4,BX
PH5RY-!CYD%FLNMWK1&A#9.C*(5J*\Q3'RF@'<H(]*.0/L27$1"W#'V@@M(?Q>;+.
P6_[VOQ_$<SJ6JON\M3?+,4MT;S5_SF_;4 DA:D-V2QHOD9V/9"!]\?N^ZF,=T850
P1T+]H:K3(L<(RJW2WON$KSNX9A5+:((3_[JK&;JXY!?7L9P+U+7I/2="+0=C@"A%
POUEU2<%5)5*HF>$>5W)K#J-8:[];!SK%/ 6J^!'@4DC@VLRMIV-IECXS.0LYR_C%
P:XP-):,4'6*KLP2/U3&8^?2/3?Z26[3LZ&/'B=F;DR'219CG(K+Z*:X *@$B:_@H
P%6W%5%U7>G)!6-($I(NB@YJSWGZOYH%PW?Q)N7CA^X*%N..1"6P/>@PKY=A'C 8&
P//Y/DOBF;E\IHJM":5744)]SN)$17 ([UTG5>ZVT4Y^/K=HJHVD;G5X%NE9$#E6B
P89$1:NF!G2G=_($3V81%!P5M#D:]HT#-4</<-G,""< :L+UE E/J?FA<0-/")?5/
P?I!M9#!^EZ"'2WV)"[,%TWK,%C;<.8>._??:; QY 5%GR1\@!/?E3Q?92:2^+%,/
P8>>T:W@CPQ/1>#(QW+WWUK]R9EEJ$'GCT17(X]?_):<W5U:]22Q^=50US4$RPK.S
PRQYES[].B_^,%)5&:X53Q7C:8W&I'C42*928[(J-6N$J,#=XEV-VG3*(^KB#"%HJ
PTDR&Y[<>=+&0?<U1JT8D*QEI%K32='!OC#+M,=*4N%;1H)<54^D&E@GPSNS_EDG9
P=[@(E4IV# *Z)\Z&NZ[NJ\0"\^M9*@R"^D59.Y?>^[V EC*$*6U;&@.7+6>%9T>K
PM);[4%XM.Z_Q,!(AKC^5.(P2^VNXF.8HJB_.L)+8E]&/#!=:$% ISEL'&G?'XOE\
P3<0/IM1!E*3Y+?]0B8.*Z,.PI^2K)C8=R1H7CN')E+PGA8/^O8\UTG<*'FAEYQ,R
P[]S><.V'X+9"M!GD(9NY/W1OV)NB(4D4 C^)]/'0DCZJC]^!G,QQ&Q[V!U4:F$8-
PR@GZ7:-K/EC1RS&$PV,]\AX)!%J9U4@\@W_&#V%\WH3&08MBN,):$(]WV7\8:CF#
P U'B L"O)G.N;3.>H Q8+4[Z*_P42ES[C5G0.B2[\E [!QF;YZAD8(146@6T'"$3
P M*GZMTY]Z>D> 7Y)W'\*!&Z)<\BY8"95A83[K-RBQ13"#0[ZLGUC?P,-K&/(O92
P('GV+S*Y/E06K:1=:-$NXP-?Z;3?<^$A$:_!E;#XS6G!@FO,V1TSS-%Y%=8OM@==
PXC&:HJ&M=$%VL4[ 02[GS-=Q 6I;XJ:I"/4]4@VR&,5PB?&(KU.QSK?,A295-JY6
P:JC)24)32(RDQPLG*CATS?*E8F/<@#)3;[KUNUD:R?/EDCC8VC7.%S]0SWW_;P<-
PUS"2/>^2IO)3H4[WKE&$8$IU590E^>QZ7J,=:>R4<8NA $9Z.!BU?V;*?$AQGKY[
P.*X+?]N:5(53!0E!OZH[)6VO.WYK@2(-49C7+1L\-V8^3;T&"I2 [\0\3[F"HMNF
PY&?,ATDH2\'RUZ*E:I67HF%.*%>U[^PL#/;U\P"0FQ_9CI<2\ZL Q$%Y--K)H<<K
P:Q\^!I0)7=L%-G\-A <$*JMM$ ;PXJ_0^707?8<'C>5XG_W=EJLN1!^C3'N>S(C<
P[L#9;6([;!^@H@Y56AK],[(0^)>/5NMF?+:#Q\%8*[1A,N'8V%*T  / J=C:@WG@
P/S$-[IBB1KR4YB)BW?/P#?V^HSE.-GM'GQ]]<JQM]D]'H#BW]JNRDATU6@#=2-"2
PQ_,O(;++R0MDYQ37PC3'E@P[MB(VL=2I"OM/5R!UC7+4=2@["A ^!C28IE%-&LP8
P[\&21(P#1B##GMX. ^!LAE_Q@9?OFQ*ZEF]Y- *9A?1C[$2N_CI:;/Z32JJ[-4QR
PDF[9^T'A9!WX5['1Q<A_9-]!0$EB*-X/L:1G:W?X+W29-F(X;Q'M5G0I]I(5N;\7
P $[<6KO_^N.H!=854W'2R,V![#ES) 8F4GSJ36_.MY"/<5AZ*\-L[;C-M/S0K"A)
PTNWWBFR4-FJX5Z0CZLC(MZX)<)?K$9J-8X46#VOK>6IWI&?AI1#M&<>CVQ0Z3++0
P]O]<)1S*.0! =1EU/AK9%L%;%A!IGC\,EF.QO!YU8">9=?KPJ.JZ?G64]8$$22)0
PKCF)TC+OC"8)!WSC+T<YXS?B.S/. 3I R-*N\$H<KTW_9&DTTNGOL !Z%3L[YJ7A
PP@SKE&JCF1$*Y'D?*.7D9 <PG#4O0YAHAV)N+C3='S/XW<<TSP@O6GB+Y@]LP.G*
P%ZAJP&=M2'2ST)#M]LW#$)7IV)0F>:LG&7<"-9PKQ1#LU8<:P,4CM^Y/NOZ,HBV8
PVR%P_BH+9O_OJ? P:*@O[;K&\O;N\'PNP_V_&03Y>-'+3,N$)<'XI"2[@&[;'IXA
P=,ADC4,U9)J2&0[J%]H\&**C859\__S_<%RV2A,@$8V4()W3?,^F:+&XNJU;4[<8
PJ&K8(012';KTN>DW:/NH# S>>U1^@$,BTY *("-J'M!B:A<A%:TV'/[:^&3AP8H@
P%7MI?&R"X2YYO17X#P>8(+!I4VS=BA_SUF($AI-!+=YQV9<*$8]K$ET-F<QIX]Q@
P4+'JY!BYB4M[L7A.K-?VAIX?]H'J/,SCX<#AVD6_Z9+[VW-$69#L)J8 BC+5MDG:
PJEYTNG/R&MFTE6;G5_]_/897_#1EN54U^XH>2<O7O6T^6O_!;COX%E\HQX[,]<M!
P$!@K93B !&;^6! GEHWGQYHXA.D0"NNH:%)5J.>GRP=XOF@R'02W$O.\' JFY;V9
P?1*=(MLP'CATN0F[>ZR!R0!P!E'!S2<:_[R.,+3?.9XX/3'D(YL-<,3J#B\:[5;]
PRX=%R;@;TD94+_;U3G+'?R=>OXNGRF*6J&O]N;H21KD!WK/-6)C4R$9L:T@HPD;T
PC\GPG8FP"'TK6IAJ*L([7.^ARGM2?"545G+%A[(TT+L2CDP(XP :9Q%TLX<VS@?>
PF:^;V:R^&_@@[!K$ZY,@F=:TUN)$8$M<DW.7C6@/S<>7IM_""5H[JUB ^4VV.4+&
P<@2"&=.>E5@09*^L%D^>O\K;F/FLW%IPZB?/'E,+];@< TIDS!FDKQW"-$.YB\L>
PU6N%E<&#\3G^.R+&YG\;,,Z4I.3,P.HRL.4\(TYZBQ4IO6V\E8A%DMYOHEE_U?UY
P3R?SR:>E!;DX_..!M(*%]FE.Q&+P^P/UVUPCSZ98#A;C5;]++ML]:@W!]GPQ2!T!
P)Z\^W]9Y@=?XNYSUEK,)3.Q^^$2C!%,X0?!.#L "D\\-<9G6LIR :8>^CFF['[#L
P-/J>FQW##L1UN]'B?"WO-"()O,AQO3[40@;8&KTVSQ<3(CJ.B+'H?'N>L<1I>&D=
P,T-IRH_GM)?U9!9/'_3*5!1A/= 0VTE&344)>HXQ=VHPMY]3#A9T" F'A>??!'HQ
PI^>.CW6^+Q-^=VLU/NT%4V,>*G\RYEIB'7+20..+"W0SLR*-H_.+S-J3P-HO0W8(
P73-E2);*G( FVBUVXHT:8"*"=PV'K2H&UE$+P>3K)K]:(=$6*^3)@2$>IQ*:$SVZ
PNJ4^ANEAO+8NQ$[K#WF+,7D^+YQY#TMK\Z>9!C3?#^KZ8]D.F?Z=<-&P0%7G."IL
PLAFK9+H;WY\FD@HX'_@$]J\B/.K&GJ&H*@=R5+BJ'O"_0-KQ M";XN,X*G@W:$27
PB$9XD;9Z 7TE_3D5W.&0KHO)6HJ O 5R1V7L\"RQFV43-Q+H3K6A[B"'#^@"W'6>
P %WZP,\$.]XY>6"_^!C-17C3")S%PPYD&W$J;;<MD,^1JT@NN%Z7LT'JX4_=[H_O
PPN3#_FR;H2W-)S=/1)W^=?281J=OFC-?NMBC)CHH<F5F/. $]-!W<F_(!=5SI2!-
P,$MOV<R?.6FM>7QAQ_$_T)D38:O'EK9=5-D[V%=A!<@]'N%NFZO4F]IJI\?-ECK=
P_>"(I N@^@!W$KZIGO$#Q<:'DB5ZG"D^P2O5-A:^R3?L&:N_T *'6/\E '?H*Z:/
PYM0V:A$B2&'@WT<UE'W1:-#KV^^=>[C&0RL"/$1$8"^\9D/2V^.5,A,9 6:"PFSQ
PQQ.L:\60-I)O!!BFM>A@BCAB&+CH-N(Z.564@')^9M5E'T=]A1R&21%0D(-S%B_)
P'2OX+Z!P-G[RD7W&4I '<&\X1P2)W\@,&YB8>ZH4BN$$'2V7C-X 6MB3-:FJ79L"
P?@!"R[I>YST8X&I5B+96&[Z[5QH8./YN XZ![B0A@)]4M%'Z",$< &*,_7&M0S\-
PL%CN\]5ZT%XUJ6>?M+//CK^P2P9SGM7@7! *E:]- []4ZXH\ 6GB<7E%L(D)NJ67
PJ GW9PPD($)UH:@-=NOF22//B1/66;4/W%J<Y^-Q^Z3D/,=%0]_C*-V8]4S@,(:\
PZO!^ F,[L_DG(GA^29-FY-9:=BI!>O:A5KY5]D J@J7?+V-"/?O41+G0/?)V3IX#
PO!*D3O+DJP?X>C(@,,3V\.2FSNS'_,K[XGKF$7;'?+[L_%PH!PAWAGA W_\>0RE<
PR;]*SKY:IW )6#YBR5OTV2R44,U<I=%*&E/SGWO.WM]\\_OH'4G5B_!=%5!B8"F<
P7!B]_FQ\&""D?O>3L,7,+8Y9DEZ-F3:2'@G!J- 7H**&\B@+6"R7OW\""PQIH6_(
P.:XQV[#756O,08R;>W,RJI3@(O5>S=T<*/%_1DO9V]VU2&+QI]SL?PY,R:-=.#^8
P1_%UBGE-B9I-L.0K(I[1\#WU/.SJSB!U39CKF >-TA/BY'_5BY\/8;J8@R[\$J+-
PMH$7F;&C)]?D@NT!P&(J+_C,<R[!6T$%Z-:!>&'^;KVB;.<$3SVO1F[YB)^#LE(=
PU-F/A M-Z<5]PHV_[0P#:*!J*B'FG+")S$3:U3<WFMR+^3IN[%)K.KBL+OX6XIEY
PP"=/I24MG#@2+QBD]5*"7&L!9O^L\Z9KE/'@A]J;$. Q/H@)A;U6S9HOHJ;N1-M/
PD1$2EOR3?\@(2$W6LC[J31\7JS^\@/-E(YV&KDHUI79@9,&X\.CKFRS+@_ I2JSW
P%#SIDU#30*O.L26($D>SQ\4PRX.+4^<!2'B(#3 KH_\1WZ!@>,NJ3:AX6=HDCIX^
PZUK:>HX^],>1:Z#>=&WPY[2DAMK-W25PKW:L"D?(*M47T)31L#840F1=OC\;BRJF
P91L:8PS8TKZOC^T77+O] JJ9DWF4X&XP+NDGS[N,#5=UD0./**01@F@6S=<-ONK[
P'*@-%NNLAUV2"C>)#A/[OLU09X;3-0+?S_P7.1;%+!4;$J<$.RV(8;V_1KRB);AZ
PC C@V@W"WL)K=\OZ]ES9K'^!"[STAXW," V-.9XMTHK38P^XH_?A+J-"O/V]+-"=
P^([F9OL4X CEQP<@+!?<SS_[B;+?A6OZ6,'"T[;)HT41QN,S,,',D&//[61<=O=F
P#3OIVT'W?_QE2(ICKQ[&]312A5Q4*BL%5IN]C 5BM/_0'3Z];4_?V29<NJ842T(I
PI9-B# V]WT._6HZ<E^J^6SS/\^H? L_?8RT$:+X2(N!S7A(9U@BN";<M9&U+.!&R
PC\=K%O<]A%/A\]WD'EW7@$.+K=MC,QQE0<3:"D#D0KE0,ZOV&@R#T]/G=A4K_!E,
P:_)ZE93]%09"Z9FB&Z2'O#1X4$;B"Z:\/IZ^'SU@=TK%17P3#:9E=M/:TC8WU]+M
PXH74?EG%LO@H8J;%?;"'].^_\Y!F\ Y/MRKD&<]070/OCW$_V[QR'69K*(-U.(&@
P!<L$*S5\65XSW\@,!(-M9G=9]84I]X>91%-#RNYAO0<E/=4L5]!E52!"[TM3>5U5
P^D'>W8,JE,'*B>3N- 5P"ZRG6:SNS.HL:#6IZGB\?W.BEFSWO*>/=>VFDQR5;[J!
PGFJ [S\2"+/!7B?[/O#+&S&'SC$.MAZ8.<";K_'O9 !O]2T,A2-?CL8J> 7)>DOM
P50WF2_R#I'$?=UINE!)T66D<GFM-S[_7:8WN/D0C#U;VU'O[?>!)5T_4WG7/.$O:
PK,8X1I@]EK\!5%W%?,-#,]X(XAVA^\X_>RZ"_OQ: <0RZGX%#C(QZMX$M,=Q+PKS
P?Z3NZ?5TM8<_'RE*TJ&%D2^P!:N[4:$;C04O&\HFQB6IGO(-6Y1?YJ(*]?$A[.$G
P#Q32.3O1FB3_^+-#V+3@)(I[YB)4PZV"-5WROCH95Q)".>*6XIY99>>Q!'VC*BO8
P48.C;RS<#T-D8'*L_.':+C-MF2A#"U/#K&4ZX_4)XG4V!O/:K(_E6TW-F]"J824R
PM%3S(]F4_CB46G?XRUM<O()7LD^F/BWQ8-/Y,WDC9E>.@.Z<#NH 2 4MFP&J7#;'
PQ,X<2I1(43YDZM<Z,%GM4S$F E;\EBN (@*'<).>P@/#H=1_O#S/7>? \@OYW>7H
PCC-27CC6XRZT7VBP?K]N^*FN:QO<+3:GTW,?(/.ED5=& 78S&K9._IBJ5DW39"+F
P4SXLI*7]\&L_O1JO'!S"*(&C^3HH%V@K:*,.::(G8@^*&G&6EI6ZJ ;]:G1%8)\/
PW.]PQ>+7.6ODT#V3#+N3F<]7(E5PT8^<U]-475.(XYK"*U-J$H9K8<G&PV(*],(Z
PJ,P4*IL[UM86LT&)%(J'3BNP>\R^C,[H]7:*1M$"M+'O2?75\;P7SO')]&8U+82-
PAV6-0_;Q(X#'[U5'?X[]<8@LKZH.^%$B,7P,YQGZ0-O6I9/O1-9YFREX%BA:HS![
P^%]:+]*AZ@+A4GIR8<*KGD;/+R3B_$.3%55X;?:)OA?,<;C(J3ZW$_/>!8X0O\/.
P+XSX"X6KLW+-W1726 %OB/Q?%ZYO%UM8LOZ\<,2Q!O#,IS<(L;6)F49#JR7- ^6.
P_T/<(5P$3_;B5$1ZTSZD=[!A B/J4CZAXJW]Q^LD>F<JR4ILXIYJRJ0Q]S@V$87&
P7)(X@J.2%9<!Z0<9&,9BFLRK;+XJ21ZE1784X136,:-J97B50 .'PW>&_MCJ"I[>
PI\L=K:HH=V+EYT:R;WNJD* @D#_4,![P?SK?C))?30C0JMM.^%/P[]9"9V<,C4\T
P^0UZZ2K3?Q1,L:1#Y@12H3&YP@UL+\?U5MZIG5L&%DN"<[3( <>F2&YD;(1'TO':
P6,)^+7'ADM&GQ\&"=@.:@AT,5I*^M(S!G+^]M]]OP+DR^:>YS3S>Z PI.EQ#&F(?
P$C&H)9\\J_BK-"^)+BX;/N%V%)',-S-I=IY:?0&,,Z*=DLE_Q+82X*!XH'G8FUM(
P(L6A*6CL:(!_5&"*OBAUJWJXXT@983^X[+R/5<6H58!116K3L67I&"CA<23\#];T
PE;)LWZKPS46EZ1F&#GPEN[J<!U2K3R];1)-E0>1RC'7\P(56RD[<R J[S W<RC'T
P_*ZVIA)5E6M".,DUQC:.1W-$15'YY9*LHW^Y8Z>XQ(>67M9*3SBH\ S/UW7E8/&2
P3Y$8NB0)F,'G%Q^@;5T\C!;UK@+^+#7 G("FDO 3_DAH27!&G$7= CETF7QZC@.W
P3WE->E7XFQ\[0>Z,O+SJ/ @V&R';/33_#!(P2OK0=ZX),QHI'Q@K^#6;0JO7/@%=
P<4_X+S4TJ0^VF*\EB,8,Q=(:PH^:$_W'C>0NYW\=C0$RND0D+M<G[=A--CVN%;CP
PKQ89)0>KM&]_P9"N[F.C;W+8ZR$L+;:Z+8(@9>*X<+7<KJR_(9MRX3AJ&>$9&OMT
P5<>E@F^$DW 3SX*$=C]OZW(24E4KR=211O6@N0=4(E$3XXW44*BMIVYGILQ2PCFV
PSRS((L<OMCLMDS?&!$SK=O7ZYB>H=.WH:"<+"9(>5<OZAE8,":NE*[?":F-E@8GM
P7@MU_CJP!5TQ%/4*>Z1_.//7XSCHD6]H+HS*\^K$Y LE+Y/)ST<]<T> D.JPME$)
P@J])R\L?L3)9EY'OQ7*,AD=L*__;X:7R.JWRT6]0;4H&BVU>MF3;?_$K90(%VHUY
P;#T]90F0'*9\Y4;,&0LSIHUOY/B]E(SX:1Z,4Z#_4J)K)FM 0410UJDXG2?5R8%P
P*;L:RS3\<+6+#J6>6?QPX1=<3ZL@=?:R[^4E4263PLTTJB'@OI4EHN$P#S#.PJ=0
P2PPIC<)ZA*#< B3*TC;W6IB> .0WPY5;MQWA"0_\B\Q*T#9KIA'B>JCJF[\T,OK7
PJ%.VN>%UTHP?I;[9?1*HR1T_J""#;;0":<- BP'<H*^Q N.P/Y% $Y_%A2Y..C^'
P "#V;2QEY7JT<,E7S3\KIMR8Q@>W<7J%ZQULM2 >?:R6A()B=%-#7]R%J;3ECGRO
P0YSQ5@B]9+*%N.2&P2UXS_@2KYBY?L:,VVQ%955=MWQ@0A5?3*W4N^<5.XA<TR[@
P6=\$IAK*7[0#-"W<>@1OOV;='G7I&>LFNRH_R>Y-LL93#C_JIEGKY+=/F^</S@]L
P-FJD"?X,-/;N0J9G%?L!/_A%D[^5' J^\.?^DB3+52="^E[D4EPNZ'T[$R,0W?NS
P%;KFSTAUW]0^"GZ$?EW[SY&#9?;\V0*?T(0 $Y5_3!;NW6@0GI4D9&@U!36VLXT<
PL&?X8PG5^,;([V9>^/9?/V0$JEI;GK%;S5@>F<*Z8ORI$,A>$A62KQ3/<)5F)R:T
PTU7\YUJ[)X7#4:QSN;?D;04,>9OL8YO18=</2=1":79L!9Q^)"%5O9G!->ID1O)S
PB&'(*_:Q&PNV ?YX,FJ"K+)/,,<TN6H;<'BV)#FBKW+*6/]\9E>T66-LV-4S)TB:
P<^ M$RA@E7+R<HHFC#/&W(6@GYCAIFB?_035_@%0C<="(D":R/Z&//#S[;B&;CN2
PM65W*BHU%)&>4FL4*=/!##AF)DY02^XL1*"IVUZZ>^HU#XQJ[PGPP)UL_*^,W<;R
P!6\?^/IFSL*^9SNU@*@<0)NB:YT=&^2U@ /F4+'V^X[&::U[P6Q829(%-K#JH>C@
P<=CN%@J?R_'C=H+0*U(C%@Q.77/0>C'-\1]SM6<S2+KNU_!G=1U*9R+]_D7V&/1>
PGL #_XU6:I#=7>^_&1UA37G-/GI&[YI4+%<]R5KDB/=?A-SRZ%%220PJ?B"*>E<5
PVF%.-4V+I6P2*PG<[#R=_[29EY?2;/4]PJKB2T%5;R@\@LJPEF<J='<YTY >_YWU
P%'6!SI_]&S(PE:R0.T,FI1&8>N6#9 I"\I@2153,69>0$,Z)[#5[<NS6%F44T,ZU
P^6DF>NI38!:G 15#GZEF!GP";S'(VQF+!#V1*Y-0%U=0,DTW'%V]I,PH.?@9RXW-
PT"U0-99]7DYDEH#;CD6S>^5(N7)3P>T&,TA?M2$B/#4IJTJJA;_2*QER!;,CER)H
P(^><3<4![[2C:\T-('RP'.2JL"VI>'_FTH1B +--?GWW15H)TE%GP<UR[:/="[&6
P0@:(QN%YV2]!'2FJP*!I6CJ\5*HF!I9*D9:,J2J=Y"$6M>+"EX'#Z=GY?$5B_O@A
PT<IU_ZH$<]D)3$2*OW-S=;UV\A>,?=!N"7SB->T;Y@O<V)!.@JU$,Q&V7*R]6$6L
P)YR>:1>XKW(QAS9EG5<>JT?H,]O3B>D119SNH4K!VGI3,>,@"KP8<W<A2OG]'SB(
P$#7[3ST2&<T)"OH],8UB.+WCA:^>GF+>>%)&Y8OU+*E&?OL?>#;&9_#D0H^8:IH5
PFXWOH('ODV:=>WHDM*<6J0!)!+FIZ)1R??2N]9H&4E%YO9$[7X\]S+Q<&>3Y\QM'
P_\-*X-,V\NE>@*L"RMZP.="7V\0N@J%-:K#;S6_'MD_>LQ=?C%!V=I]11MSQF#48
PF$5VK'Q5"L*B=$XUP^RB#WA)O9:@G+C)5</XP/0JN66(+SE.\EUNZ(KNR)2XBR7H
PM+0ZF6T8N2M&+\]015?5PUS*&)(S6@]0)>ZI96Q'=S_'"*M?W(U,C@I$QVK/?^ 3
P6/;XV2F[A.V8>GF(IL4PF3\LL3RL,[]Q0KY7US;LN*2N W/T\4/;TI(\0ACT[NEI
P5228R&!DP99#T]DW*:E[U<R+JE;BF>(X!(Q]!J>.5'I^!".#B>)C=W--!("OPI2+
P^2HZH;:/4!@EYNU6:+5V=/AYCW-C=NCC]/@S)^4K[5&-$5=?_MK$$<=8+L$ATV>V
PMB[Z7. XN2HI;I%ZN=&>.)<Y@AMW6Z):\NUL4P39T7*XY,5;;(G"&*X=NFS6=,TA
P)<9@ ,ZJ'\D;9L[A\AJFK=/W13)5+-&E?/DT0DF;2 ;DZ_ZQ<<$1\+R0:JN#M\O,
PQ7.(!IU_Q_7O-';>$4?UA/$WD<Q109SFE\A!/ LFV(D-(XA*.$,(0T92GB$ZQ#-W
P#4J)4\#S'-R.[6:KPYGK<&M(A[8ZX1)R:/>.;-.NZ&(T8+L;BF.AZMKU=WD'0(*Y
P%\W\OZX79'*[CA/^JJ>YQAW>K.=&U<[H!IH=FQ%D*G[65E_UD-%=;E7<*C$%,3[!
PX;*AEA\&;CC<,%<#2H^^+GX;%-&M]QL/7!PUPLZS N[G#Z[!@Q;/,.\U;W"'*>:V
PW=]QXC:HHQEIRS<ZSG$?*=[$/A4N?O$C<=!P'CN'WIH9S@J@FXZX4H(7&9:7@9>H
P8Z%9QQJ<A2I81DWSI4,/O\BV&E#/C,L5&I/LK/_0BW#!967B\Q^Y)#KP'((!"W]2
P\5Q*4#8A;ZE!MU9=[S1D0"0&+K9Z : V>Q#>AIS=0JQ4:$AQ=M:MT!)#XD"@.C !
PB@?N(X3;2^*8* &WA.O92RI-KBH8',TA9P=+$I1=$128%(E%5 ;,H(_*--BLZ4@C
PRK^]K-#?@X@381CXN:/:]3N'+IXBY;""S!)>J2_7(V&7!:J^71N!-^+Y\:ZWN7FN
P;1MF"/2FW/0(,%/Q%=#M&H@XC9+M\D,*=^0@4;:D?H1E3Z[+I>_,B4\G'JKPN*T5
P25(:1+;N+/U\=8!*IU4+RP'$]IV]XVI[\:-*:\TY)P[(N(P)W?2TT)64:-X3#TZR
P-?!GJU1,)3BC'TF*BIVXFB7O,:=WS_S5Z5RXZOR?E6'&"X5T9* IG6&6=NQ>"(AS
PL_\JF'+()!?O@+5KDH:[BT_1=5-3_A]66RI0"7Y34*S4S-PZVE/;"YYN 'N97[)1
P0V,0'3C&&9&]P#,*+W7^9-]K0\UI'N>HGY-(E;;S7A$N JL.$ G3GB-H^8 ^VGWL
P68G:>PN= 8+QV RY"ID>1.'Q$DU5P\-:)N UZ4GW+([<HG4?O WF]<%Q U/M$O6:
P,\%YL[W8'#4+&PW5* :8V0((5^R1O_-N T86+#VI0\86Z1R3_:C7T/<.RDK+B07-
P 0_/SP>/(@I%-]SK[4OL_%&<$GN:W3V %=4U5607!TKN\7GM.!Q_K_9-,DJYES]Z
P/DK72<+??9U -%K^V4,[!'+L!LDAA\B(T2>RQ#G!QB_;O:IBY=B\TV0S9;21EM/A
P(*FFWI$WJ]BQJ,/$AD4$V][& P\^LGA7N33IMB[N=#UU",-VOER:D4(-5IB[H<-$
P]>.L@RB^%[8?A/]QAE][,I:NB(/$C;WOQK3FH),9?M1YH6CW<H;W\DK8V,EN0]NE
P\H?L\^)V21"8=BK%3V O-O ^B7%B!J6NOZLO/7MF^:<]Q7H5"*W7AU/Z VO_7JLF
PH6?L+@;W?N6\#Q'Q'=^=!R1[C2AR4+>D,2]+$4H;&Z"; 7W<&+Q<^.PJ[(XYU=PV
P8 [9@EIW2TOY+'+!2Q?,"=3"(Q=-4 _J^BX4YIX'Y2Q6U#U(/L!C9<+L:(EZY!E0
P V*77<U.1_[J]1(?Z"\R3?X*>+8B^XXON)C4W\E(VZ,\P-5'K?">W'4.;O=X-?B(
P5+I;32LL\KF*ID9TC<-\<$6@M#IAW46$_20R)WAKA1KC)Z^B[*=7VQQ89\02X\)?
P339:",DKK4O#[KO;[/%H+;]>&ZXN3J?]T6'G14B*QOX.G._Y%EM6IHA)T2 0@:=:
PX8YBUK7:_HG*($(]=<4-6$W)@(\P9E4P&,EI)DT;NO^&MV>SI>^5>&I=-E=\OZ:B
PD!(BG;KJ2^Q+OUCFMHD\4D"Q&)U6,.G32I(@%VJ[+*J@<M3 $0?$O&3,&9O8!6X^
P9"SR5-"!?KO';P0:A2DLA.>=79 <B=F_"DGRN*S>2CNFV^3+*U L]H<+/4%)WL0X
P@N<D)2J5$4J"; X0E<N*,],Z _S+ZG"%X0Z_IY[)F&\8PZ+>!RDJX1YI38N+RY=X
PQ8.GYL0!3%4_OD/H,K2)*HBDWU&;(BQ$.<"0!@_*NLPK&GP+B \XQ!6HT2A"6::#
P@P=Q=E0O VPP:GX:[Q*G\UVB4HWR>$7>CUF"<C*+:!V$Z' 8PI%G0BWR5BM!]/$Y
PPA_AK>IK(:Q"JDNTBDNDQ,"?6C]@ B$MH^8.%\FS)5JW9(JD"M#B33<];.@BC:7T
P'\D"OS!;HL.8LT*SZ1@DO+K)FAD5_?MW[KD(D'OTB3:VODF("Q%;DZ"?,L!5#CWT
PQ^7<BFN(K4/22;V_LI<'U@:7KAHOP:>@LRW45EU5!?ABJTAF]AI/R']XTR,0$)][
PIU^JZ8%F)YY"UJ1%-!OF,?=4/EQ1!HL:V\XJ(U=Z\5MMV0YO@58\U%@'*KD2S>P2
P]#@W=%R,G344;UL"-D3(&L?K&.77_4M77D&5U(I1W]@?D@@K WF#E^NDCU@G7TR?
PBQZ0$S$MWQCE9^R?N)L^B(Q%HPN*+C!]+E/=')*:(P\O+M#OI_F-UTSFI@*(;P=M
PLJ*FPK:/'0A7M<?-), 9!6@5G_(KXBE)S.M<@0!%=XZ^B[I ;Q#,_N4KG0:HS"5O
P>9"+6LVDJ!!FK1VG/*"QG\E$\( (AQJ<("OG_[BT0QF=GC;,E5!*;[G[LY7.;(&#
PY<L)5M&)IS_F2S.>&D==#X>U..[YB.&J![9Z#5TSB#:*5)TN]?S*.W#<0MM'A3;$
P@+8ZK>O8:&CA%Z&M-6'D^D%X8EY;P+'<*S\])LB['Y6 5XO9SQ$PBF";E&RU=?9\
P>@_O!)2N"JVDU2B*,I]3\RJV66UU,4]>/%M-;\.DO#YP*RER\A>*2+:]==$T="EX
P8UWL]PMT0QC;="WL5^B$!H^V$%G&I*%4#;E:#SA5N:.;"*U8.DR SO:E@7M\(YUV
P?]_%.&MA@2D:<82I(DF50.YP%8T7!X&VR_--%K!)#CEZ99T"';N-YR^^G^T7H?MO
PI;(-]-X-]23?(4(SH;</MU,MW<'?Q?[?A[$_V3FA:1LC&! $%31Q?2S3S,>60@#'
PH<537BJ91RD!E]40K HV B+IPH]A7>HT/.\6D(IR]X -Q=5!<$(D"!H8Z0Z"/VP?
P%4,GUPUU2;W$T%/?Z/^)S0:$M&CV\;'J))VT6982\<T'-KWWB\ \8N;Z>R;64T<C
P"L$W.K //2=Y)Z>Z%)CL$K60__$"X,9Z/<3JG#3CX['H6OP0' ';_@K.S)_UYUD/
PL@OQQA;I#JCZU<] ZGF+##1-U;!($,"AMT!;PT=GE;5I'9&5SM,X4GJ0"0<6:ZM'
P_W K?"@>;B\?#X3SHN;>7C!1'+Z+XQ([3Y'\R?0I5FFP?P8%JC;S8^9J#]:4SHME
P?9>;'_#TR.OI5D[8\_*^F9>#9>)Q#!V$U>&]&GXX4GDPT_WRIJD#+6V%/A]C!C,W
PW]N.LO[1,<$3PW<DF>>LN3N!L;S\!\_2 6S@IS_9S=KA4Y,1=(0MQQLUF=R%'6-T
P%HT9UI>[G#1$286QAB*X\*9; >, "Z_MY!S0-,($T0=D$C[C:[@[$GA[M9>'70)!
P![L J=&:[C:\S(3:(=4X"T36GK*NY:@D1_):>6(3B]7/3T@?,M< E$Y#=+]W.L'X
P2KV=]"T'-;.Y<?!"#_/M=%=%1.'-2$[=K_1;+1W$486<&8V8 YPFAV-;R?=60L52
P/1,OL5KRW](YI2T .5&TIM9A?:TX:[F"EW6S%[,-'4P2?-RQ[7]_[FZ3V_"9F$5,
P.KY/2<F VI\ML=_RB69]<>:P?E?7,$83XKG@8*(^48*3;=K%O@7VIVFJV9:/8@U2
PJ#W4^4[!V]OYM! #!+NGZ0 7F)!$9XS9/9<UW.*&:Z#5)\ @9Y5G8X#EPK[2_"@K
P8 K+X&/=E,^@8LR?^'*F8AMY;@<N<B[L"R/GR&KXVBF9O ]R("9BG$ER_Q.:$%>*
PY"ULC;8<5\4PQ#\ZQ2!-=A;WD2JP[D=J_,;([[B1JYSB\DUNQVY6Y-"B-U)/M[B!
PH7BC^('$O(*=BE<&C!S#=14C+5W=Q"]YT(2;" <-,KF"A6WJTK!!-U0HZ)P1W%P&
PRO2F2"-%S"3!D$RV6;L'M,?9K4A<S_4X&8^2O1--GOSU>,CA/>NR=,FH.:1ABI%_
PK);,Y.>EMBL[-FP@4P,9HK.JZ+?LP;4!RX&33E*$(TRSF/IV?].>_^P%,>IH:H<:
PK[;@?^-6>,#BHY(:95.-@X&)0WAU3-G?3Y9<CVYG!9-%3")CQX8D$[-C07](U67A
PGU,UC!+\H>1-FE&R1C-;A-!2-"SDJR1[))PLY<<$"(@4B'+669U(M^1J&"H)C00O
P6[E^UC=4"X\5P8R#</2.*.<^8Z9)J.BY:(+_<;PVYZP)3@;"N^_*L@"'H=Z= 5<S
P8MH@""FXT.*TP,B^.VH@!@H-K1(VQQ50 8Y.@LN&IPXA=+T&P("#5\2J3D!'&OV/
P$LOS3DD'6N=AARR!\7@WJLA,GD:@:5^+<?THN')T_O"/WF(ZED1HCQK(/B?XAH'Z
P#8A#+]=@_)9,M5.3L$1&0U(.Q3<%-X)OAS7FG\X[5Q-1GI<3+T]6:[VB/66YE<?-
P-#S%<9CQLU)H.EM8>B?GY<UJ4]G^)P(.(*(HMV9[FQ^*,O2@"1V"'FC9BW:-,RH0
P%K7^R85B$SSK:V_:HEW?5HB[O!J1+5Q!0AQ@VW>9D(C,D/-/R?17\;"M0.W51I3 
P-"1DXDX.D>@J_D[Z= 'U'DDU.A-LFTY]U@L?'96C5]SPNL<T5\'<#K@#>H!/O\4L
PE^?O1IC@)+=<1TG8\>1 8_H\J_/>A;%J^,/[!N.GU1QV>1*;YEF+/GN->G+@XA6W
P#QY089\N):%1L",%7D&&)1..HB)4N=NW,0 *,&-IH"7$#LQ>FN[ ^B59!)(A!@$A
P0J)TG9!KT68:$KP5X7T.8'S?LC,.$370AY+YOET+%:'X()/ LH&/>6"^UCW&,"-[
P6EWV;GS#^-+DH>,!@#[!EJ3Z2R!_HBXYTM*6KW<H(RK,_H_!'IU%BW?Q+WLH1@K.
P6$@ +MZKHG20LUG?<UMK4Y\HO!7RT/U?<,\Y1FIV@ B@R_W:>4E9&52X,DS?94X/
P'"H4N^6'H=!16%U]* DCXS]^K4./Z3-G4V[TP]G/^$;992)>2Y_(-M6>NH182.I!
PQ+>79#]W$KN97K;Q(_?M&=(^N!"_MHE=*#SU%4*RP[>LL\$)DUO$1&)H@V".-]_5
PA]#H Q]9?;-^M0'@X$"C=H@.2'4*!.$(T438 5/F[2.9N?;KK^IEJM>%5]-2N27W
PG-(""-+[MP)U-92'0^(5?^+A^@B@8V$L900X)E!1;1N_.?'ZK(4*J(?8^OLR>RYB
P>&%,4X8$<!);.Q2N<E*NGIVU6U9(R$!H7D* F8/L?>D0I6Y7PC>;0<)N;=K#J?7M
P2W2(<1+'&QG".2%.$PN!;_6(K*2)E+\]S5Y#L/#[#/'OODAXV+&_#!8V[P;W:*:F
PU1\L*13XP!O?+X%%[1':O:91H C2PA;I"VS(ES"D!NSTF:Y\2B0AMREJ/7T00N*/
P SRB7%(J[AN, MSQ@!D[BS&<NM=$0]V-+8TH"EK+Y#G=VIMQI+WV%-E7$HIV(9C:
P92)CK#+IV%F#7C/R[HC*!DB!(?!9W;A,,\+4+ Q5@^R9!50Q9ZT60";,_%5W:^_=
PW"^>U#5#\^NK^P81_<>B>W2'[:G@QLR+Z9EB"\3 &[WF,8Q=C&EV;<^1. =:7/XS
P=$R;,BJP6<?A@KDH-%<\JIDGD;-J%^#U("U1=0TA:+S(YM8Z\"WY DIHQWS;X*!)
P@/T*D5>P0MD>)5?&_V\HA-,=I$JOEG$5Q,V3F'%&^LDF=:@:T>+"L>@-M>_6B';F
P[NS&@D[6F @H7KK$R/#N/9N4";T2_M\H*SLLYJ'^?Q4WOPH"*GJ<0:0#]H]/E5Q7
PK4:.8U":;*2+@_>D)\ATVP97T]QV^V1);!G6)Z4QNIEZ'E!$<)M.S>0.469@_!:&
P[D%?>+ S_<1$.[I[Y(TW $Q5-&ZGL)N;S!=B4@@4!#QWDEDP/@_[2#//0G@Q0]08
PCCZSJF0U #.<:/<0V:A:[A.XNV8PW"&6Z!N9P8Q68F13BD77'6<@@&1Z2TXZR<.9
PB='N2EY?V"=Q0P-T-+H;01_XAMS2#[ Q;2X&0T\,8Z;^I;785.E0V);X=]8$JB:(
P7"A,KN&MR/PGF"R[,IFT036Z9#;*HZ$;]0-KH?F$(N \'0(-UTG3:@3GX.%Y ,.E
PT_;@<CNF^:U1<7")1?F/PH/,HG^$CF*JW=7\Q1,A.QMY*=<>!\<.VY:JKI\&ET=8
P<P>O!(:&T.Z+.*E)G+Y<RB[([%J5*;?@&A$MY@"=IVJ3>[\-F^O:#*&^6&X#"0+G
P%.N\Y^J]^Q](P&#I2R$AYB<Y5<LAQZAH11>45#A=1.2\EG/@^LZ*Y?6G:JFUCL?J
P.FL-AC>-O^@;0M'8+[%8X_R#?/6>U-V.[*)SC/)D1)& E-6(R[K:![7P:IS!]#_,
P_)G"8H?RR::^R8S*"HIXQ&#I6JB!6\'C"_?2[N.N/PJI-B<^54AS&9I6N0KR\LEG
P"EEYH.?@=&^,A($A8L8FZCEU# [>3&<M7-,&5Y<8>S'-'#(U1BL&_:##/%8U[WOE
P*<P,?%IU+5Z[WHJW.Z'(3HW";>BA>+)IU)V6N'9MI#QGF"3UN^7/SSBF>(/:_\X 
PSGAKN=]QN__L1.61X[OH91'S*M7XC7S;ML@?5!:OE8S8BE%S:TWW-@DR_)Z61_$1
PDS9.V":T,-%2*UE-T&E-L%,EIBO)VE[Z=!L8F1?/8!T8]+F^Z2;2[VZF.02R$LHI
P8RA2-_!(36H^:=?8&/BL"C3<+<4KQI6DJ,GF6A4[%FS)_K7@]DY<CE"LK>@9>+75
PG9^N1Q'$;P:1M"\OR#AUBJ_@P7QU&$EDY RH7)1H'>*)Y'B.$8 'EP(?7+^6QZ_I
P*]Q!(@X;D%6J5C<<FADSY))B4F35O% UQRXYXH]#0NULO+^-5_*/Z2C[-]&D#E4@
PH 9#)0!;="H9=0D KV9VN>RW?H D4S[\ZZO%]NW>F*=NKS8E2RQ*S;*#Z9DSE,M9
P>90^(V$BP.\49!'(6WX#_U-K(1[HC8( H69^@'QK77-H7&@=%+3]ZT$DQ>?#6;N2
PN0_V8=FRJ<D_8E8(GB2RL%M)<NQ57J:(! M75)0\8I0?YDC1SH(0OHE#K/R)]D@?
P=$G=R\53[Q78TWO&"0Y"+7R>R@5%(1W;+)PL>G;A!/TJ:,3R)9]-P?3/5Q +4M):
PA/[.QG!+S$_0QZ5O-@T/88I5F'M!"39UZ5A2B#X\(T*S=\7:B_$H1P,;)CC>%D>+
PN+*=<S8NJ^.2@9I]83UN<PU*54'1+G0R>P[3&9&X;Q/84J9;2I8WQU3WW;;8ADNB
P9\Q>QVFM,#!]:*,;V]$S49@.VF7?:U,6A..*QWF5GON)B():/Z,%C!X$]=+'=[7D
P%;%(&_G:5DH/." IY)0DV2[O"6E_\"NS\UREFO!@.^_Q9J[O:6@S ?V!"CVD/(+Q
PZVSDT.M<558I#=H8U'E)ZJC'2 EH;\U>'6BDTB1;GCS4!VT($\:S[) #QQ@&\L3!
PXG>WG:NT-[#S--4\C*^NCKK$JTV(7!!0@I8:;5JP.KL+-H41A)NB"C'4"CG0()(+
PG<$Z .DF!*B4=9>1=%NJOO34V_1<\R>]$QSE[Y(O02YB<%.8\6&8&2NJ#=:_%:17
P'8JF=$*1/VW'FX*91W:W2<N=4=8+HAN5&EWUY1?1./%A,'@KV$DJX!;'>IM;36^#
PX?=X X#0"[/$2]X5;&'V:G\[^ <K!FNNJA1M)L1T_A>-EI*BFT:>+BX]3(1THT\;
P0/+\YL(!;\S.7;\1B6 %HY(0->=0(.RV;K\]6EM$5EL@J7-/NP&YA+\+B4YJ[VEQ
P[%]4:% K;FY89-0J3K.@V>^AW &S[,!MPC*0<64 @=/7[%V*/;/OW43)?]L'LZ5,
P%A+4C^HT%'D^;!:4)8Z2-:OU/U=L2N8P3."^"+JG"*B'Y\I:U>1D8Z.5YSQ-(ND*
P&BQ?):X #2?&Q@#:(G;BTQ4@O-H:-*8\^V(RL*0&V_UO@/!2K3TY0_JDTO0!1"$K
PN$(T=,[HP,/@Q&*NJ>1,($-<N0COC+EC9/ U)TN(OXA9 =SL#[BZ7] DN:^5\4M 
P<[QZ<QA#RQ17N^,Z>!X4RC\,\S&KJB1D79>C%-+-O&]KWPIL/'%.OUE>&"6\KP'#
P<I<SCP6"_F/"(*5\*/Z09I/\[F;SN'-+H- N%%2 +TP8/H:9(A=$<SE.Y <3"#&J
P1F.^ZNAC=[_R_[+,>H,97?GW3O5  N\$:*(H7 <Q@;'SM%CHYQT'>^ S_UX9Q3CX
PR%_N"7-O5*3SJT"+S65)_UVYOV,.F#X],&OT[HDP<.^QGY^M#!QZPNNZNSOH&\B\
P1@W@9C3 TT9#(IS\RB:D*UA1 -@?2K>#(>\$,"7NM&IZDT70=X_-+L'"M[ES"S+/
P!6H;OJ%/UQPQ=H2$&ND,9[S"NJ="9B1LS,7OV:C3V$S^DU@[K6=4C,YC1#03DX(O
PJ$RF AK1U%=RQS90BPTDS;"ZZ<'F'-ZA2Q,#WGY=+*>(2;S77IY7Y\C!+]D4.PW#
P'%&AT)2Y*YSO,SH+XL ;GN96#\#+^CBH5BFU.E6DH_W>]HJXAX@FGJXT<=KE4')>
P#-S]W2ZF2)6R($A?[M--*[RNX%Q7L<C\Y;M;ZA]O$+N/V*%@M*ZU<^[%D5? 2-B&
PF8G0R"T66ULP*2*S);XY*\21/0.:&R?D=T:W-;WE;#"W2RLWQH,XGS.2?5%+M)_)
PJ&[&+C-$-\CV^'!SL-?)0'"?=:-P' )> 9I(D0B/1-9E3/**,V?U"@B%2]_SZK72
P+$0;U">%"D\WVC>O5*F]22:2:?]0U#TUO0EK#R]7=8I6=R:#3[L,N+:5LZ/G*?'^
PL%G)90J?QP]T #*PNMO6H"*,QZT *NN@Y'JT5CP3))"RRY6% [*BQLQ "HQ!G88M
PDA42TQ,$RX\NU)F8@$+7R\,Y"-(#'40:)I\QA'KAW-:[MOKSCF-M*[LD"8MV/T*T
P)! S338GW7GAA&>8ZH@:#0AF&\NP8_N--'P?0T@@&RQ36J*_MR,UWO&##4PQ1/9O
PH0GPD&%+LD,3<#.V7)26_,[(<>(>"!%8P4(3.5@#&ZI$ 4Z\4IKZ5:Y\R_'9C=#Y
P3][PY?Y16Y+N VB5'U2RW4H]%Z&)C\75A#G\9]-29=&!EO&W"W@9==40:+4X5-6I
PRL#A;;DA$AC(04S%UV R2P.FS4!5/@I9..I<5[Q.$DPRXFU,- <E+H$Y7JV1ZN+M
PJXW\)HC6)BCO!)FT$<W;-KM5Z$IX-MZ,NW06^6"J%?.W%X<]<!"A8Z0"5KWXN40<
P4X+78>QV)#U@!>A\K%Y%#^3)QCP &8V14)]OWT&_1<)B7Q,+:6/M$(SM4'K7RT%*
P:?T!6HLUPIZF1YR%]MK_FO +PT_X===9L?7ST8$:4=NAUJ%5Y#9^Q)@OD<L7;]_;
P>3&498,^N*$.U^D@UU>T]*W2!&BA?V $T1I$#>S6$53ORXWI;48<!V%1#5*KLQ/#
PGDCC UG@M )=^BTCE.1:(84",N *R,LS0^X91HA7$#R[SLB/E.<Z^PN[9#['__%*
P!4,#@B$=R"A^^UR]\$3@GH8[&9+&4C<=KJ"* 'B3,U)]H"C;<,^$EJ><+8$MQU9Q
PI-,7*'"A&'6(D48P4?TO&,C K6?B_VC(M]\ 7BYZ(G8I;/1[\;*[K-,\<0Y>\S8W
P:DD!GVG!_#J,1R'II'H.PO&LHT1T>CZ/L*F50T&648UQN_!,O3-?VUDG&JB2,$D<
PV+#=E@PPC5%8L 80Q8'!NAAK8O+$^8&#&C#4*K,;1MPOT(!FZ$\3S19JTC$A]PBN
P<#N[0L=T9-:3VA?SKB5/W7*VLVW;>=CXPZ7R,-O/6&O!_!NC;2YBYLJRP@2<TB%,
PG%!D[!<8J/L9^IP]U#.X87?,K"R\I 6(GA$GKZL36&"6L3$KV(0ZK[(B>L_ $0BK
PS#HD3%I8V\7'US\&D$<$&J08==*_^-&>^*$)Z=F"+^R#%@%^K _!42QN78Y2$J1B
P$ *<#AZA,]200VL6N%3LUJ$Y";1,?@7OSW0V<I\/+)6!,[L:C8"2(M^-LJO%>'0U
P=I$DP)0DG;%9-Z'QMMS68L;.BZ<Y:CDA+O:7]VSKN>*LX'"@'2CL'4Q2R ^P'(;2
P;O,=WB8^V5#JC&J@O8CO&K%AMDG^I*]XQ]!\%0P"A,X>[Q.D8)J%#Q8[,,XC_7>_
PRHFQ'&5"#\VVY]'P2XK,>^$2S#HC$XB1KG@,#< (OK\[.=TRV&XI-19K3 8B=^!:
PN<>_6_>%#86,:I-HV_9P(6P7C\R;PLF.ZKJ5G*UN0MBNXC:4@9I64\S90\P[%XR/
P(!4\%^A!>.;&+O4QZ^[:/>@&B_Q':P  T=E0G$$>!4-6Y)@*9 2757-:=/$F.I-9
P#>1SBMX(!&?CH/@4=I4E@>2<-3-OZ,45M5_AUU**OE"#JJG4]*YJ<QT[4V<9QR>7
PIAC#/FV94QZZT$:H"K2Q98HQE?Y*_KP34#NZHIS5E5CD2< ]+*R''BPM[NR 5;F%
PLU=)- B 1:.WQ]Q*7V-O4>MT3?%1NA4A-$TM &]-VJSO1+'3!9KL,;<MD+W*>J? 
PF(U ASOP%BX=XA)WWBJ2FN^4>88JMP7!4P* 7.!_8/#\, 3Q.!<@X?$V*2_:AV,S
P<*;[!/)EB%P'O#U?RC3+Y2]FTY2PY+ OASV(U^5_Y@"6"$Q#,:_O\45/0M $P8JC
P[VF+($*WSHQQ>7%,J3 A?G59J6[\N.0Y,4MDC0Y$]0B7.IXY<>2(BL*FN9: 9#J9
PTHA9G/3C70)SXI'>WEG[17=[BXLK9G)5@A[#O>JKD<]MB5UWZ,[#>J(F?L_?1^C;
P+\W!UW/:54QSP&1>A*V*$Y;R^!>\V1<5KUOCI"AC]J]R:=SCM,D8VIG;?JU?DX.2
PFET9>XT\73@> 2J&A0R54 )A)RL&>4Y.O]*^VG%,G[AF=H5#Y+.<5PM:S\@<I&U&
P)K*J2JZVU.A8>"<A 1DEMT?;[4*RJ#0HY.QO\^,$"I@SLMM#F=,0AY:IS++BM+YT
PLX_$G#)Z.C7KMD(VZY.^]=/7BNYW.E[4 ?&;W\JN(.X9J; RT;"5I_R70,ZE\92)
P#[(60N_9:HR5B"Y#05E@C@;9A5"A.T4ME7&G^*BM!E!A:VE 1.W/)TF4!8)NK3*U
PEH.GI.F"A>8LKGA2,[WHD1+!XAZU!SAO\)CQ2A_0MV4>L/SY<-UG+B:6V?47TGNC
P1025?I4=;]N!K3X) /(8#MWEWU[/2%Q;RP1!6E]1^'5BZ@*!KP6-D"0UU+-]<W7K
P4QR>O$+X\=?#N^WSISG?G3>D!@'[<N<5^?L7O&TYR(=?C$,*K,#9458-T550MH]>
PRZ[&?^O6GDLH?,=WIBM?C_+1$Z4/9@W2'15=89ZYF%S<,S=2.[R4A!ISC]URXD0N
P-+76ODS[]GV-IY?GZ.ZPD161T1/Q%JE1Z,YOS0__*N_\#Q'%8%OU5\<:CU.I-O;S
PFP)@@B'M3K=)&>LH,;H?NF1_'2S!N[P3Y$"J4E@**V6-RA)GD<;!B(1E8T>RDG98
P$6@%=K1W]!1,RJ)]>@ZH*3R$P+ZG9[S7>Z@%4V)UBD(H9I/OH@@1(QI4MDC*K(P'
P4D3AS62(K:I?@<8FN3M+J4%YO"^UVE.\5^CLD4CL#Q$NNG U]@NR?HO4(/G,T_65
P ZY2RS7MCEM#Q0!J(9(XPO1+.R:LA0Z/T]"596R.CF,#& \:</[5:)=:)+DW#PNL
P2^2$5SYF(9VRJ91&&:?I"YMU=Y$O$*90:!(MCI^LOKT^,5#I7//*B@\X,ZC5,L];
P$O7H;,ZA53E3B.%I6=2-?9%QKA \G8%?K^>YE%4JW!NRLI2!/:]:<;:L%Z3OEE;Y
PLHK*O^T4G;6L7]&DT11"'^,ZV-%F!=D(2+?R[#7,B6A]:DT#V+)8,I) ,H-[':J)
PD?7[E"V%ALQ!.W/ /<IGLLG,9\:"!T:ZO#&"1[(O9\3P1J0I/M30B[G/8IQ?*-J@
P!UB^(-+;>TJR3:%>TT#ZRY[<^>@0X6;.;)"/]Y_J6I-/Z$[/2%_QAG<Q$ X>09>T
PKGCUK/THUY%$EX&O\'] .^0H$--@6-:*7>4$Y["WB [B,=RYS/]<G@,EV%Y%'7TV
PVDF"&P'"$]E0F$1)D+YOO^<!IYSLY\H0=(2$20?,NZ"[UGVZY\I.FXC8-43[@,.=
P[QY!,&U%6=2/)QH 'I0R1Y5RHZ4Y^ZGFM1?.64A9 ))D%)7].*/ZSZRK+5>\=<SO
P;^1IU[J\FH$>0""QLEL_3-60'F">W4\6H-T-;+%C_B\,1NP75$9F**7ZAF='@!MJ
P7V;"<:HH;0M; 3AT.>>F7F *O=9%IGU+I@IL\,DS<7T2V5?U$_3HCS,[3R45!10_
PV>&OAJ\0B^!&VH1M,' >;#ZRG#SMU-5P*D]Q>#Q4">=1]:7:WC"36U++G_431^ 3
P/:Y62BDK>S'0>TAJ4HSYTM;/0762N[O2Q'ZC02&EJUPLZ\Q"/&+M:3),GV=D2*,K
P],Y;I]WKJ/(/^VG.AKF&+"K;+H;5GD/0_U>-FU;GK"=*<9<BT&WFP4I9P*DWOX'>
P'UQV!JD2AIK.KF9B&?U2#-,AS#'_!6MI+K]0^,JZFYB1^(?AK[[F_W6?GJH3RIP,
PS?'=0ETF)Q]$Q"\H&P'*WAOSN_V9=CXC] "K%A@;U;)O4[C 0:S=_L<QCM+*J-E^
P1$<@#J$;Z]];8P:-IF6QO^5G@M@OD3[+.\66U>-E#D.^1LSTIU4#[8W2;DQFOUF+
PAAH&D<WI'F':S > 7JQ)ZPC4<B0RKXDBT57(?!(00YQ>*PH7_D,&6!GB+"MKZ[_=
P"^ <ZY\*6I/Z4-I*Y0+V>9B3X=[;"UB3\'YG4O%&;\HR1R:_ RC<9UYMH8)-EJ*"
P7P*Q+!9 KH<^D<L$,HF'%<^*PZ(*]G ZXTOLT)&;#6I=-#Z#O%F-;4!Z-^DA?4--
PU^S9_8"Q7B;4L ./HN<]'&;&K &AH/DQ$!]8R?DRU2>X/4J3YOWN6(@W$UJXS((+
PYNV?Y.<HUVI@561$F:P -=GALG*YX(U.@UKBG=/0B$A,+OY5M'3F5ZP%P.@;KG,_
P+4<X ?.W*89-A'L_1Z4JC!.PQXI)#E71XZH)MP+B#4LO48OIE?GY3QO77WX%US?Y
P^/4;NQC%CQ::30,EK[\U-*R6KC,>[Q* FJO.=B@LB/N[Q]^93#?RA=*81_!X:WH]
PBXO55ZGD7E"2M-' E"1YX0Q4Q #(5=V<?XLI<E7.N D:1##"L L]I+#4*/8.(W@+
P=+%=J?I7Q+46TP2-MS!EB%@<XG^)/*@J$L11SI]$AH&;L=IFQ:,W&72U"_4"FKT;
PH!CS']K#6!&=OO>(*+X:5!XU*JI1#>R^:YIWX&@#98%552J9RH,Y7C* !>17NL>O
P4_XKBV."3PYO29X7^ZL=-F\:/%K1BQJ/&6'1;?Y$)71N:_UIU4AU<6G\>E6)&"$S
P(2IK]+ ;[E-YW^T'9=43%8;?[AO"HBNL%7HJZF"HWN]=$_VV;)$DVKNZ R#.(#AX
PS]8E-6177YBAL(\LFF!VK0O9):>+AO9"N-8\4AG6G;X(.*+>SG'.55.'4+[C++7L
P/+GC)#BTD*#:[*%!%NR<M54/:5VY..>)OIZA%9(+2H6'%;M**P[8WC:!*'$JR<?<
PT%]SNA?5@A<(')'1@]OVA79;O!(:3_0^JE1T9B;W!N!*EWR[X3GFU7FW%J772)3*
PD5\)^(5VY%P540=/&;&!@9W4]=4^RME97[\/<10=,;^(RMV7_%+[Y_7C=>GD&+!M
P46!5? WXCE34L 3XPE_HX"(VH'V!N#TPMS#/0FS&%(F,BH-9;Q8SM IJ+]4QBDI/
P;>D\&9>%W)*M7[%C*.%!O#N&E;8&6E:!8*'A*&^GZ>>UQLEP:))$,9]EP,R1UYRL
P/,X(LW7BF-3S+OO**1Q@ZTLYY#C6T]345.=+9N4+=+1MPU_YN13=$>-+QWWBJF+5
P/JNL.O84<*K\S9I\_GBO<;OY$M8:%EE3![6>WG]0SQVN8?BF1C##+L'F[\O&H*0,
PJ-B<L/8((0=!&5ANI93]G-<45&J+7D<24E,XE8=%A7 ?R=+5K YAP=%1&JU4W9I9
PWQ&?3BQC-HIU?CLTB1KJ90C_9_H$RWT+$)*ML=R_CHD974VBKI]#8E_,MNC62/8H
P>?.?W51^/@PM5>HJ/Y,!\907^BR\>')3&4=6/=R$&UA#WLK/LRNG8\-+QMPZ:U26
PNB11F3?#O;/'+5Z7KI13<OMOE6<"G5N&GN7W4.I<&<>(Q3W_*QJ$<QR1;_J2/3A2
PSF-.+D5"4T[/P:%E&"_>F-J-@K7?X L!PZR $P(C>O/[P3WJ\&G4V+:[F:&_^/Y1
P]K+^/)B<!=AUGK]&\)/\X;]%B6D#11U1;:YO=SJ@&:?1BOY2?,H>93E?SQO0(4(+
PI0(G=S16Y=HM.@<HL]8<0_&/!GNA7G13+$'-J,3_+V%R!>-=?#)BY64?0>0^$NEU
P;RG6P^WBM=%Y6:OCN7_7/:CU8XKE'ZY[/:J+.D1#?!?0O3N0(-!8?,RA%*9;NK6;
PDI !?/SXT=1-XOV L](;Y7__&L6#ZZ<:HELV]X+%XQCA52@4T/=82N:+ SK! ,@@
P8D R8_E\[+!PGYCM\(%62S;0DWB53<30:>RX;A+6#)FF X#WX96S/&N#B[<J%-"$
P Y&>K(#DNEYW8S@3NU^R=I*,9H_1UL0'^C*;6#^$'T2)RDPZ\ZS8WWW%Y'2?Y2_R
PF^8X3TUHOZ"*2<2FC>'THVY@Z":+:Y_V#%MI-P>3=L:%D%-0#84G"*7#B(\H)J0#
PJSE ZQTNZT,)X;V-Q6@@%HC>]AX;XAFJY>8SON^:UC!N=YZ%7]:4\B^V-ZNOMOF5
P9!5GYK]?ZM3T6[X0BTLP1'M/:P[".7,*,DA6BY/W5]Z(TR8'>B0])8]EW@S)A=3,
P )U?P0IELHS;:GRME<"MK^SLHO 59XX2,RQU;;[V-\$*#7=@Z?AG&C9/6$F(P6"G
PIOD\IE8'U'%4B4MM1*76"U7$T7#UV,HNN%T!NOOO:0C ^(S_5XCL>)33UVQANW7O
P7PQ'!N,?X<Y33)F'T9R)S*/ [2S>SYPM\A(*N^=":312H?P/ZY<@ZQT-?+\Y#;.W
P%ED9<Q>_FNV]\J?BW=Q^OY%(">'DH#A\;-"C666<I6GB=OI2 ]R6X81/NQ>J],8T
P!*M&T;P%XX6C)^L<G!,O!TT]KBE@&IQ3#K^A+,KVWH,ZF452 K#]:2CB%>PZ%U79
P/V\R@77F?A"JIP>Z@H+ZP"B_#-<TP:_U74JIO'00:)=>+6R]^2+L6QBPX$>'F!' 
P)0&"[T-BQ4'%=/!\SYPGP*FHD"<"6(G\\$O- [Z05@+QX#%C\"7;<!\48L=4RC;C
PWQD/FLG-],)*[EU!_'C1;E"AD[Z_\,Z^ZE,'^!'Z.#SQ;/'(R<*_:TD?O:@$@(&"
PG%^ $;1G5F0[.["31;NO\/Q>$B1IJEB;212&TP$9B: )TJ'@(ZDBTHO*/Q0OMD1V
P(MC&YP;<GA#DZ'T+_=V.0?&[KBZOD]. !^!Y=^ZOV60=EN"UZN(XA;6>'Q(U/MK<
P>C0\(>\-BG]X<;QEYK4U:XDVAUKPG!=L9Q]\D2>)%\)CO#8=)@Y ['A<JK&)=E<N
P; #[V@#]W8!127:3$8H3ME#$%0"<6Z];)-]2 ?0A&MV!?;[,Q@!"^N;TA/*V_]['
P$R,BK@V#@0N;Z.@6QS>P67E8N_I^S)[V6?H+G6\.!V4$ MHY/S^'AF\259IN<__Z
PUDT^]G31'HBT/LY)(O/VFZ==):1C@[@*MEQH%9DW<9L"$K2@^-;= L#LJ"?!(HF5
PSI0Z=W?MH[RN<]KUT?..!VD&2$R[]\H#DVS_WH*<F,Y(N\[L/Z3-5!K!CB/T5'56
P563!<>,_11I/S:C<'F7R0G9^U?S0YL3MC?%MN<!U[L&\?*&#[JP6]*8#+Y+XLC3F
P#P'FX)"U#H$+1QTJ9$-4C-UM4?#4\3YVMI!%"AW[>&DCB2S!L%:]-',[SK."JN$X
P;T_O8Q\V*; 4YFZ(59^1=YXJ<7I$/]S=#1/SV;?8-ZAUURW]#R5'UEO:/OY?/H7>
PDNB[[:7&E[6CT!/L"4D;T/F^@WB==8<49.X,#8SP6*^Z,>6LZ#S7),K+QZ/G4D9E
PA6!0\(".4[JA\_24*FS31M?3P85&"^48LFG!I_C"]4T4#P)M,/G:4+#JA6GK1<8H
PEL8'/ED]$XGD*/*BG_./3<XP?*I?NDPCLZ3IQ&[TVR]\7-?*C/;RIOR*%2D+D,RC
PK"0S19X:T>KI$](KZ)\IUXPV[M(_&MX/!UZX[C8^RJC'52Z*X%[ N(>1=^#&O9#0
P\?;VIH.._!:^[<:<C/CVBZDW7,3(:+?.9*ZP^O^Z4I2W7^/,?.69A'0KGCDU?(]_
PL$Z+1L\B<Z(X8:RJ.I(.6J\(NCVX22<FU_0O3/\JO^M0A.7OYXPJ%/$\(%)8B&NW
P^G)"=BHJBKV^PMK7I$8,@#-M]-S)FV#*'[&^<M<Q2$J;J0K4V-.^8INO+*FR["(?
PIL4=C0TN&1#,&M%VAS)TK)_/!U4 K6H*'@.M(I61G](42S_!0=$>=R(I1H'=VOA>
P38"D4]P',?.4^?!\TY4V J1//GX^#7SKI!D*VR'.PF4&,4"(7IKWBX@.D,-?/=8P
P6FSQNSB--%ENB)5VBB (@+.2:88Y#YX)B[W)NE'TF'7.-\(^QZ6J,<P;>Y/21X_$
P[X73U'Y%9XF2VJ4XX]*C1JMOA'M9@(E5C&"TZ;@X,1OK]B.)H-WHFX22,0%:7[V 
P=GBC $=<_7A/>O( ^S"S/@NT$SGE)>Z'DOM*/SS.![>YE8/#!G.=QPBA-S;$3+!@
P1__S\$]G+S<EZH5+:B/.-X:SV":>!<RC?#B_8#AM-S_22^_H%:>R;L&4=?W3M%)?
PX 86?PC.ZQ0LC%<MC2'IA1U,T,I.:4.:L@LUSZIXO((EAC.,%!$Q>[K/(I90!S3Y
P;D^DT)$T3NG<7!Q)D3%XQPMR0F7/M:28'T'P*[;O\_F\38B$IF!.QN(:=?J'+.A)
P^-)FFU#@EO%;N:H'#7!0"A@Y7"R/;X1&G>\:&=HDRS/,TERKE06&](!8#SD_';+F
PT=G6%1F&^$74B%<-:V C4,EN)I'CZ=[SM+?D%>QWT$>U'YXT#ECGZ*A2CN^=:[F]
P:QZ3:W?K<P-]]B.9S',B1%@J0>\>X+V0)+QN+HUX49V54&E)H1HA+Y?]3E< J_/(
P$R")D&FX(HLF:_B:T!+22"D"P&\_>HZ&S[+4GDB=R);1MF$(JO?5N^ D!$FCBC%!
P/4N\DN.^O?5:SURU_1'DVJS5[W\(E!83<[0XN9Q8>?732X"/XL!(&,G8!BY0U8HL
P\IK]>@QW,J7Q 6"KOEVT,5=JS;C_!+L5!."_AN6AO07;]3S<';5-7Y,K@%!.BCIQ
P4AO@>7<LF<$3T)P6&D5#GLU920QB9OF2(R8.[N'W!4EO,J5/4V\?>D-V=U\W?8_)
PM/$>;*#3LO^"9 UL]34P(9ZU-!K\4"AN9ARSTGY1*D7UL3A?2PS7W<V2&]NS4K!;
PG+P*@9^57Y==P2J%@KB-@-<M=/9_9.C%D^@GJQ&XB4D.IV"-^SEKV0]E0[5RUN40
PH6^HOJSL+,A\G!O[E?=-=_\6= ;?$/KBY$2$W5U]*"9@\E4S)AM*\*B70W-98WN(
PRM0@+B+/KB%XV.)T&Z^C4F=X8"+OCT=XUJLG0?%2 XV>D>YEN.5>>5O^;6EMM*.9
PFDZ49(4_@N1/)5+UVRM9]2@Y"0UXZ+HSV.Z29PQ.*5 M^T)*0P'#,7%7O?KT+][*
PG1.V6)I+I8,\N2U<3!'01\BB[:7JC$2B .^]V^AH4A-;/5D28WYK$BRF3S*:=Q^^
P+(3\UFD5X+O:7TS1.7J-;196W>(,P;':;N)BQ4%D4,V7)_EP6K1C=K8+++ J87O"
PS*N"X;\J29X"4:KP+(AO.2%X (KQLQZ:75=^1+@% HW*]<\ W$"[TI$X*DS#1(:0
PS<GUJAH;RCA2N\%1L%X'/N?PSQT,T +&OI1'"0G=ME?_FX_Y"^OXZ^11IV<OQF].
PJ)ZX5TB2EXO"CUU)'4ER/[2RBID'GJ8BTCG8(XC2SE!C3]6]#Z+(V29S(HBN'S,_
PA;#3MO5]4.$,COOT(H]!\')O;L7.EP5/-V[&(Z4'&<^K+FT.U,VTE?A" &V\[A>F
P%F[B1>8IKBH 8N9>*"T'0^!)A(CEYRE&X_+S]6\,^1B"-GHR A@D8+U+%>-JLSUX
P'O%!KH>+44^63=E 7@5=*O?R5)P3J-R<FYR.KL.W/ 6RATK*/"X8";:@IQRXF8\_
PS@Z\KA%59B5>:0&&AC$*$K/ \S0LM2B.&STO\C:7_&P+)#EV_*/7?&6H0+611>?=
P2WSQ N,7Q82?,VVF0!E ;'%U '3;1;&:A  NI" TZ^VZ?5,IP[NPC?BT%[UR7_@5
PWOR-V_9MJ4P(WDV?&ZZ/3-%$U72\L]%SCK[S]@B2ERY"7?XGTD^@[4F\N+<":K)6
PQ]C 6<H;$NYDU.D+/JN<\R8=$W$"RZ43GP85$,BP"18IZG78B][+B]8I5F:+>O3X
P>]4LA#\&K3@Q/2L_2-R2K*4\<A\&:/H'TLTAF=";^')+DDDC9AI&^I%1+G;3-:GC
P,.?G,>+!G>U5"/924^8 JJD0JOU5PJ1OPD<.-/]DIOE._C$U==Q/_LVV]FOI=ZC6
P,O1!DA^$=2EG$5DS*="0(E@45G-=6XVQ"!F;XWG+*]8J_B8@WL_19?]A$SB7MU.X
PK11K8QCAGV>>\2H485).YF:B:KX,WWC-7=ESBK7+(G,'9'L:]0=&>'=JFIS:A=Y"
P@Z=R2NI95[AA"?7W@:D3_64O2BBP][5SRD!OONU.=H!N,[BW%I88-7Z2UC'9*'^B
PP+ZRA!?L\=7!B!W^"S^]J7>![B_ ?<.BIG*4NOGC? )NQ;>N4.I\"%%\H%QW67>L
P]FGRDP1_EA!H!%'#!)'L&5P!$67=% I0WX" O4CFO$DJZC_S3M3/J;FX45(5<^3*
P0VSA5S%;=LJ'W;Y1XEL:P,ZZ9UB>I[)P[NX)VE*HU6W<Y:%)-"76QX2"Z'S_,N\(
P \C/;!!!DR)Z'1JCXF1<H%TY9]\75AZ\=\%[<&0T![N5[A3^_QWH7S_J6O!0\_C*
P>,FKW[@B$Q<8#CY6TFR<Z&"EJ&["O?_JP730X[L?0HFH7OHE_WYY@4JX&>9CUP,Q
P=-M=^'6CZB ?E@S/LX3L^PRTP:]GKU<&BRMPN@4M.1!+^)]NH*1RK&C)2/#JXM=D
P!X2#\/\"Z:_AO\7?HX60(Z]H[=VGB 1*W/G9B-_TK(L*J^:>E__ &$)4W'BT$V7R
P#_XQ WR@\">V$.%,&.S:"=P7/[=TU4:C3/%_J>Y;^)(<@R6@YGOP#C&:W# <O6/F
P9E2]%5")OB#TC,$5>^TVQC%)R8_+=%&-J$FE*%[,=L/8H@=7E=]]F=//Q;6SZ&4Z
P0^B]Y^^UQ6A_9J__]5^H;B9@\3]RJ9<1Q5O:5!SJ+(Y4,>@\)& #PY,4*.96+^%;
P?MQ8E]P"$"_.^N.F7YTI"7:EKCO#9BW<%D+,#LD%*AI0;\7%3@B,\AIA7>F::96P
P'^ H1I<:28MBV4+P1Q]ON7[8RT1PS>$BF$WCMP#/:-\4_K+]X[W8WE "BZF#:I8+
PBWI)Q,YQQ$R5\#6?8G%L\.B?5^B5X[&@*?)^M*H&;F<$=H+MJ.#)1TTT.&&>SR;H
P5</LX941^]IKE1I3F3%8C1W!/]&R+ O7%.A0:!B'%9XT7YD% R,Y2P\930$W!Y^0
P2AE<TUCI.84="$40T2WL:^)3#$%F?18&QGQ)*%GY)3;I*VP%/=(T_X?4,6*-K1H[
PD*4DQN!*"S)>68?C:T?'GGI.F774R;?R;0RNC2$\^ )(+Z3;YQ UU*[; ;%6_A-,
P+H>JHU6*Q@#@C'#X&#\6<]T&=/F#TOIA;G/3N!3QJIB];Q=HE?*]'F77$ZDC0(BZ
P@B(PX3%*MC"CX_*^Z_]9CM4'&7YL')JF7I55_O*X+:ZWELBU?%Q5A#[V>(RUUOMY
P/:W[G-WYY2O6PQY_=5L4,/Y7AH5H'7B-]G#9$?#/>6@A*QDR;<AT6.WBGK>PK%EU
PF23LO3X#+S^T2<#T2%ZIRS<L1:,9L%!/U+[V'%ZI$H?>HUD+J"(P*55,S++T2JK_
P^.T;@^N>3[BYT(:NZAD\2[+KLH-_;:UAC@Y":G[Q21)]6-]O!HN,ZXI:JZ_7G(;3
PA2 2 1V&W-PCJ9A9Y1CHG/SWF7-T59%62"Q8IM6=0FYOO+DE? #^#GZ5 SQ.UDY*
P0T]!!?J+&#^7UZQPF(:C\BAF'8T"]X%-^\$G"BR,&DIE_\[4D/AP]ST=7"+1UL,%
P,0KT['EX_;C@YB 1H:Y6'#',^ +KS"XP3@!?>C#0OO\?QH66,I>WY2,6.LM.2 I:
P$H^C&VH+\T.CK+'%Z-&F(]QJ5C0QH"3[$Q8 B %L%#A>>H9AZ4*],?%77>]:E>H\
P@MT=Y2]4:K\M'%/%')2\D-KY:"@-GQ0DE3_DVA)RE@D\Z;>Z&?,SG$2K!S&L*P Q
P@@^&'J5>K40 "J'&!@9XR0DUWD=IO^K#B0RGSGNO9E0*N$[B<JC<JPV1\IF;M]^(
PA85(]"!0XEHI8'R 1H:/)FRV+&CQ()6MT4K"5.\*3T9#/E? GW[NMV[P(-*4$B9H
PC(X@+>J_.9VK]%7BP=2SV^M<C*EMP"O8(C)\Y'.H&8 $Y&6J/Q;B"%&G26*I1^K$
P:AA<'\#\ZY_#Y13WT.;4&:^5L<O[C1?B3AAN5O=0Y"M^RX^L[<*5D@8@:YMIZ]ZC
PNL;"'!A39?;-CEH38@"NN0UP[0QVH)>O].>'/]KG0)/^=T",6C1/D#]29;-U5]'N
P=L$>5\8@S%_BM7P8\/^^96LE-P:U>U#G-YW=99B#KPM[Y:[:#.=499-<C)XL=5_C
P%6<N\*/>,]7'"HQC'GW& 8PT"'U7 K1=J(Z5W3C]%-JV1[2A)E14:[:[*CQA2'"4
P658K!*"N2K82(Z-%&MQ7M4)D#P3)L?'/^)"1"40Z5ZNC?^QJ"#\[6.P$S-;E/-VX
PJK8A+)ZNG:F.QVD219>)E,*D>^W T8JNE+WNV:,%6Z?2R(Q%*#U9SSGK-&B^!.Y[
P57 1?=2B8O7\E(0RSK9\R='K.*0J$Z;L]3^Z5S&Y# 1P6D9P<^L5OISV-A"EELX<
P]E73]H*6U'',[=+>\E+9;5[T1)T@>-'S\%:.#,>*S6")$HA_#?V*I 4CK0J?&=@\
PD 2R8BACE[R_3J&TC#)'<V4&V2"7A34B-)CT:).7;(6]!3'LAKXZ]@-*W4;(?.''
P.J7%283_APWEHOV7);_ML%D=B3(+W$,W>><IIZ##SM;)V5ST'V>H Y4%,NQ_H(KH
P"$\2=3R"UQ5*%N^=U.F-YM)^F/GD/*=EA;^:<O$),YWO K-3A,1^*^?N]-#KK&JV
P^OPQ&J($_G)6V! -"]HJ6+]FU#NKA-M$[B;^9?,W(V%(-)UH\V/G<]/R?/4I_PGC
P(WROZ^$(2EO0!KO=S@KC_[F_A2H]Q7PJ1F#H/7GB(/D=R%NEXS EQ$H.,37%;/6!
PC\4YR^R[A.E>KWB>7(\GD4IL-[CR(3FVVED\ZIXRL^,6L3@4!ZZ[2%HO,'PID)RN
P;Y&E(0U9R68@]S.+5):T\+ $$[R(]>FK.W>Z[7_M !\3L> 1V3WY?BJ/<,= )K^8
P2Y FF@,[^/15<$6DO?=KU.R7 UT&_=29KGEBXL+1/-YVI4Z>8^G_JLF;&.2VA_:^
P>CKU\J.SV]RM:K"B!ZIQMTSP5ET^<Z[;OR]\;2\O'&;*8("7B1JS<DQ79&@@?]7 
PS-GM3@SL+X6:6JB_?&T>/"W0:\[(MU_K6?]'-R$[#NCYB(N)MA\B4>D>U'H\9P\Q
P:\6D6"2RBT45ZVY-UBZ8IX7X!NPI0";R%9D-]H.DI8C5A 5 -]?K5JPX@8X(VPQR
P&6O5.F,">VGZ]UQ$\.A6GAH_LAE$:<@ZTY8D)WH)TR0G&F= #_+H\7'GY4H.^MV5
PJ7N\0^FS_PK,=R$KB/O;W6R+=IK!>:B;DFJ1N )F@*B3X\PV+DW?=L9 7/_:%WK<
P("F4I)V/'0]X#,/7;+EA1\&&-<;(M_8KN9842'+.4;/D$CF_IF5>RVX(Y(R)ZCUZ
P4VQ?C7?TE!ESZ-6SQ)?P=[*5 \1]<V\%.A"@_/D+0%,@;4I/#3/4N)ADZ!9E&U%3
P!SLA:%7\ 7#B KC<)'+;*T:)4RP'LH=\'@?C^;&VLH9?D%+94VCZDLJ7)ZHCC$5%
P^7>G:54MW6@O!5#5[$C&P^+?,A?O:;!5]7E%MI,,*DN6I.TM7[&OV\9Z95.=3S<!
P..4EP\%MOJ:_]QNAD=Z_9][I7$[P8\US'H>Y-/_YI'2 U?7O@6!;\3:'7J6;HP$5
PM2^;)829T26>ZV@L?97<9HJ%V[F,BZ8<MR8XR 4QA*&@8>9YBQ$M=EP(%L=U;W,?
P0=>MD&C3J;F?V$KKD_)4'$"_XA7/+&4^XCK+VX'Y*O,VV9=B5C?Y/$F$7N8E.T\U
P# O]%%20@'I@[ER^,DAYG.6YO<&JTNIX(9Q1@ 1MWV3:>+CZ?3NG5E5I/#$UO9UA
P/Y5."<2]V;@1S>Z-<O"<=+='$8C%Y9E'&M'"7P:_,;EC+# .)XJXSV?&><T/:VJ=
PK?@A.8&U%F2S[.?XD]M\?J2L;L9!/Q8'UT<V723_+:> KT.ISHV=AZ(ILE[T2OOS
P-%N6IXYNVX/;8X2-[.@P?Y#L&O'7=V 22]0N(W-=4IF%*<B;HX'@#9M9Z,E1@].+
PYOOH.Z?;V9\@BX\<TLW+Q@\R=GN=##S. PZ3_Z&<3W(?7?2<;!M5^Z !PU+'=#4)
PD4Y^U@OT045L8(PWAY#M-7B",.UV#VF;.*<;X"2*&301%U=/S$+GGKXW7AS"C@>!
P15P=U^(560E'+#;MSDM_W0IM)*B6,ZP4H5K^?J@X$N;J7AXVRFISA[QZ?G<9_I$$
P'&B,KA'6%4E?E&1[+?LV;MCQ[?1W 76;%C;+#8"ETY9F,7.!]\BO^W[KAJ?W-6\S
PC?@[#SI'K.5^TCIG%R!IK]W3(M:& 2^1I*]+3))3A"CIXSKMITH/NH0X]\QX;KUH
P$[];VR@')_X;YRR8#BM-HZWT@@"V]H1^A%WY^T\&KB(#,#! )#R^"RD+Y=.Y>>;\
P.GSEIH/TO':(857>H_([T4B) 9+O.Z-X! 8J63\I?)IY35IUG9L,].;J0\O]S)P@
P8A>71S/2_*<]IHK@LODR+Q-D"R/G[?$FP^](K*F=2<L-N%NT-6$A\6 U VY,"G&G
PHQ!$\0L/[/]N,=!:+G4/ X</#\*B;N>^M#^-=7HCMI"1_)5:#*2,,6"MW),U1#6Q
P#&EN'#*M8]T2_C@QTD>K>^^ M;YZML\CL4<.;]^6";Y^1!"Z"-6KP':/,5'P]2VR
P%<A_N2<:;"'7 -%3TO)[P:?M"\*]Z2=<7%..'LH.@^@#[6,#_JHM$FJ8_CSA#JY<
P4,'B0*U\YBA+B-P5P[/@D369[@RLS'1+*9) 2 CT#&[8>YLHPU#J901>7@T<&;E"
P2W,$R0)0H?X5#NEN94 A ";-&)GI^/7O;)L2!$Z>_ZD7+]T\D0HI&\/Q/__8D,#%
P@+,T5=#1Y;W?;ZENQ(,"Y\$"%:<@F_VU**5O(J"NB[>/@9"^IWOF,+(_(]4 4V6I
PFCA36Q6R(CWRH'L+<X>  W+2-1IUMVT=V;@B+YC ^YZAW!Q]9'^+Y0.>!*HAE)S'
PI:=[#4;5M[&;:J7>*,M_S;;G:7Z.OM.((M!M\MOS/= R/!"'+=A08@[_D,5X$OK?
PH5,.;QRG<)O?:>L.F*:$]@1TA!EI7@6IO318@"D.O<2V'*+,FV=S5; SKNK*$RS(
P(=&0A6(W5,TI8]!GL.<1:AU,ZO+7AXU]D4][&(EDM?28)AL.Q L:UA[NP:XM/FD$
P4+&%.&-QL7$I-W57N)=_M+PV!0EI$ ,:.+==KB44>9TLYD:L? :CH5DF'P3F-!V>
PXY<>WT$]+D%J-<"0,]=)7^:QDR'CU&(M :DU=5)(Q/-<=^LGG'^E01KJ-/?+I*F2
PSIS[_.P.&+<V_W1@/6/NDRSANU%I,7)THK\;'89[_]O&L+$&5H6D)%A/,WOGX<5Q
PQQ@\;XF)*@K-!VL$>9H86E5TP<^C>8AE4 ,GD<5.L2;(GGN$=!3XQFD.&0L,'!0F
P.<DFII2H_5?_XM240>-LONE*VCJD&X?%JP>&J\ '@:0%Q:7'YD+:_7'*U1HL:06!
P'Y;!Z>Z@7?G,\O"?,M+"W>W F;AE2XO 5HRJ*-H.XL:.*0=5@,H)X(W!&)" 0Q9/
P. AWWZQ(1_Q@W)';&(QY:W#<Y[1+N41>ES8P<_1(1^=69G_Y:MPI[9 I*%8Y"SJ&
P?G#KK";66TSPF2U"F^K+HT/2L6(4ZIO@=CJ]WJQ5DX"TN9Y4^79_3$'Q%(O+"[JO
PY,(=IN#[5%N$63*I5<9%>'0OEPH[KG9&=#4'1!XC@DR5[!^E\BEECTF!0>5@9G32
PVN/SEZ5N%,K._G_)5&&60$/KI.6D,.=?JK@I2PG>"_9FE,6V<0<=Q&RL9TAF4HPX
P%MV1X&$^R=R,UKD1F+Y[TF6="+I.45-O1Y\G5VZ[(+>=+$1[Q+I&NNHG&@ )/FHS
PUQZC#(E @QR8,S>\9"XKZ^U9W3T'X<L8DD1=6U_E*3_)A?H7<#%BNNSJI4Y-4Y)F
P5VT_/Y4T ?9]XAOZ0JC4,V[9X[0N?OE_/D@>KC']GTB:A?J46FB4,ZW.O@'%8,C5
PXF6QJT16W,HD!\]](1!D8A]K'?7K F'Q%Z$%BR$JR 5->6;;(D4TVFN.2,ZL:IN3
PXL0S:AW3P^MD($%D]K_M5O?Z@PJ;L% VG6-CT!>CXPKW4$*RO=OJL,Q+&UQ $NGP
PG[;B1J#D92>A,%5U_N8\I,,&>$HS_HK+6$2Z"C@3C%3CEN#4PXI*,,P_!7#%:$F,
P6]2<@SJ,8YW@9_&]%:O=IYH)Q&$>$?I'3I_?G'>Z=1R_K<N=KDG)):RU6C912M/)
P7PICLO+/Y>^8!*%Y5?4,B70MJ@&$\&-$+GB?$63!5W<0OOV6_((;_0CSS\?J;P96
P[T2J++#<]<RW2C5<?A(4$>^F_A!X3DXZB1;QSH]WJ'YU&,Q0<F^XAHA)19.69'8J
P4BWS74 H@04&4TRH?I79@^LP=QL<FX!I4VL<)4WN!%O-8%P(-'  "21 FT;LY7:F
P#"JM1B-" /H?^Z67\LDRJ?L_D,& IC%RBHL>'8>'B1X]5*F!C)^QE]H'J-"?K$<S
PE.[L!';FSF,5ZC6.CMJ$A4Z# ?!,?I9()I0( BW7X/ES+$S09?ZCC1.C%LQZ;U7!
P%-]ZU.IJ>LO%AER-W0^QCF,^&^04D-;0590X+B/)RV4PY1KWAPRHP?RVX>[OS%.\
PBM1TL.4'QN0R\KEYA\C-PJ&VFHVH2=T\_]9L:F^')ATZ#&/B5]_*09B_1NBMI^GH
P@45/8P*;P-[=7Y1VW$R&# $2^*^&U]A6X-YTV7!#,;H3=%&1+5QJ>R=?47USW4= 
PB#YY9&0A!/@BI"R6%EN^^-"JGM]GJ"9=[^>A(G3U#"R\8;"=*S%PG39O/)]ZP1LH
PJCN$:6#TB^JF#T.;NK^]([9M#^5-])SO+H'WEVJ(:7640F)$J/C=T<WT#2EE4BS$
P!_[F9\&67(L&\)M)U"&R-0<JB7<$-6H)%I (E'KPX%-2/ >!*0E6>D3@IF.KL$!Z
P6=SUMO>C;*!?[(QY.5@?XIV^(WZO*1=!LP"1]@'LJ4-?IL:R@=SJ$EK2H5>?C4\K
PW (=/J)<I4RJC,@X&<H]@64;.MN<V<X>C"^2+Z8N@N<'UC7%3B)'8G(00+=S=O^5
P:N6\>7F[?U87Y+W($.SQI474<"@CI(<&71=''2SVKD")E,DU"H8KEKQB/BTSWRF8
PGZ9_,./LULBK_^@55%1PF6%ML_NU@+"C01QW_ ZJ=_-539%7TNW:9L"V]&ET"<Q,
P5%WK=EF$-]QQ1(1X9T=ZZZ]D_D"'K^8*'$-*GSKX00O0)*9:-G[,CAOOF^XT3K=1
P:@2':([*_+,N2@5Y%G#5>A /UL2_'*IAQSIMM^]T8^7:<5I,D;;8RR=2G5-=R2Z-
P9"P-$SG'_9QO488L1^E^/C_)\)U$'9)X;054P.3V'EVY$@QI:>EV(IT9D>" 8](B
P"MX4%0_O!^-R';'5'^R-7L#:[[8AI&+D@6 FI\N\<VM756G#]"ZND$?08$!1VR4@
P7,L.4(&;4R%1;RI5'%Z)KLL!H+XRB>/='P/@I([E*%A["CSZ9]\<N^%/BMB8S1R+
P%V.P(/K]+Z>[P<*XV7-G'/U"4Q!X#7!W@UWL\@$"(3"7S%O=\/;@10AYYQ@44JK5
P(?)'1<&11RYUR7-U><2M5'A;.-P4Q)1S8934[4TBJ/SVV:JC&KAQ[!(":H)<2:K=
P)#6L5ZPN>_VH5%C15;J*;[N6)F<6EI> :<MANQ'/'6QW-0KL1DWDFT];TSR(@X+-
PC87B/?L26\C3E3F=@('';D$\$Q#OZ2WM>BJRMJ?A_&,<+#MWN<GE]&DX_9%=CF/9
PQ@A9 WAW%FIW(KU&EBCG3H]$@7R]-YI, #W8WI6V&)/G+WTATDI2F4[%U2062H!$
P=H @Z#3Y30WW;VR5#?!:E7="BT<W!:VS+@93"A!T\Y-Q2B5(@H)"XC/2);<@NT.M
P!C%?MCKW2)VGGAE+(%9NJHM_@,%.E5\K<DBZ\,I^8WRP>*9X M]^YJZL#@ 7SHN=
PJ"I24&<+?<:/9"V76CPWA5[.[X:";TY7*2P]2MM@96?CNV%"B\-U-SI.12(FICTP
P)8V%O,N)QR;"<MZ >\V.35 T.WRL7II!3\_)T5931(+R-A)'LHD'\KM3"F\P.L9S
PBA2X$^E+1+($,$0,,/'/U>=7?MCSJ/! 5V(=*?$.^9Z&3G><@,/!6%IK):'Y;?'.
PMPBYPQ;</=<J6UZ?)_/M 5BG5CP.[) P0!A[T-3$?>D5G: (<5G+-I7DGH!;MZK!
P.BM*/ZMJWT+G1:KDYD.@G-9K\E2L6?[ /RB7-<%AD1(*BA.C$,JUST(GG'=^F4 <
P,Y>N\$Q26!7\+]T) 1F7-F%\249GHV@SUPH<[^24O"UF:]CR&MPVG/PS;[O!#7?U
PV5P2$_!0S90"$G>#EXFN"FA\!-*B\#99#@GR\9)/&HCKQMBM0B#W9OOII@GCR8/!
P]TZ[12]#NG$>U:]Z%C!!/6Z<,R!&9=#\NG1SGLR_>J F#?]92$&B,S0 ]&F_4%&7
P>BA'%!WID<JF5S(.MLU,J:.+K\O-8X<HC6H >''.[[6+F]6)6Y9JD'M&KF[6,KE8
P=CD?J3!@I81=%K27/0W:FO!0\X:_P[EW I2'83&/!]53#[$85C0B;AQ6X>]UN_TT
PGH]Z:X">2^&0B'23H'CNSKVA71^Y22<W@/IKV"DO CD&SD#_C>X;+63\ZZ.YE5L\
P*OA=V@_^>^$VVT91OEX/1*_D70@GO=DCST5Z( 5<\ZCU'@_K;WKM<57G\TDUP MC
PA7<=_M>NP7-^F!?>#"ICCW"@H?!@D ]HB&@3#FR'^Y^D4%]ACZK[:Y3I8%7>VR_.
PRFT*PGI[862_5HPY(K(BHLQN7Q$I;ARS; $5G(_O]M=F7MXJMV9S\WO3$\Q>^0 L
PB9G-6_*]-,N^Y&T50V]71B#B5(F(WVW9T)8^C"TJK]AA,P&*GK5:7W/[LI"VG=%;
PKK]/XB*= B69Z^KV$GFO:IPDDD&?M(AG3A'\F,=@XZ94$#$C0M5<P\^]#*'5D]U+
P@V@P,NTCUW.9TKI(1\U1=KZS.J^,\0QN#P5\)0# ,3RJZ5= Z>"1F?NB6BXV;[@G
PI*ZMCB-- .M4<Z4V=2<U^# 4-K+9Z7VL3<QGG&"<(G?:[ U2:36K#1*0Z:@;Z;AW
P?#I!ZR_-!IVU]W#F:XN$Y[];7N)^?&DE%+#(9G..FS0O?WH6*<?SX\Q>1\//U'JC
P.AQ*04P8."EA%<6!QA^"/0].!(+=X;Y>]\J1?OU];X.@[T(CLS>U8SIWF?+@A!9J
P84SW"KP-$J1&3+Z-Z()G@!*P$4T!Z #FUP *2DR&-[3,!96R6KY:UY@F?3JE:$(@
P0B8MJ&99+'A"V445%^H@\'SGD/TUVE1L2@69T&.US#9U9JH]U:8896X&X"<B[CN,
PE%L(KSMK7;#5CJ$E!65/%0]?JB,T6>:ZFKS'3PPD7)[AHHF1W$O/3Z'SE#'H<Y@\
P/_[5!C$2--A&E9=_HB]KVB=&^QXD0HSNT"L*NAD,#CEF'\4[D<0C>Q-;GXEGFJ"Q
P-<+4EG2H%)2:,_7Q3Q$$.*26*?5M8VZ$J@QDYCRUZUI/XYPI.,@*9TD?[YO+\53A
P;.SD!)5*IU6039:%L!$LM+ *U'-?:R9L$JY 4;B5L^,6 8Q^^)"M5.R=3.[/D">C
P:6FF!H1X56T[I]U$QV5Q4<%%%,Z%"XN%2[P"U)A3G.16J07U?@FG*\+[4&[D4$PH
PG$-@@8VM\BM@I8]RX:<<NE\E@3?!"2BK[=<'[O@-SS"Y&5\=?'T$-U^DZF<.9^_H
P!#*B(8>&<V:H1?9>$^!S'0<":*K5;W #R;[\"#\9<@'LER^<++7::SI3NW4W"]Y<
PB_;R5999Q^5[1(XZA]D>@9V[;SBTAUS'L5F[)G"%/<YZ(U!&W  /K&W6/\LZ3ZXC
P3&-T\WUB;46=29[%'-^"E13+TT'H]5T/LM-E.<U UF5KDFT?AXV4U[%C"CM&R-)F
P?R#</@\5Y$K^*RM !S]U]9-WYBY*W,=K:%W9Y',>@1V8M2G;2)8&>&.KBMV:ZUB4
P+GMN1 XDGZF8V./4P:G?)=09Y@8XDL B6 <^?:X01WN8:\#5G<:&@!LPS?Y_ 3:F
PC0N"S<,K\YC.8JS9&PDNK7;%W:G$7NNC1GPWE4E6*&=X?\"V$1,O2K%QYV*J$+^F
P8BENKKG>6+P@OC-2T_&Y@+WBKAGP61)RFP^+'OY@QBM>K+M3@;^ M?+?H)VX(,#/
P>/B #9UDJIKJV4:8+18F]:SRC(';PDF 6 -24NY+"W58 0;K'ZI5Y% B'DY5')NS
PNY3/CIU?/+/@[O07T15D/0@I%]$!2T0FW J&Q5J*J&7)X9S 9P;E3WG7H@<&LYZ5
P5;=0-RI\TGP8-- E@<*8'>)NYB>[AB@]T]/Z%15,A)">TK!C9ED.F]L2D\<!'M54
P*FLB3R4 IW:?O@!-OCXXIFXU$*$=>;;2G.C]@*SE?ZWNWIT+*,B3/G*)RDS:0Y5]
P+GPR'?6^%@#>G)\T V-Q '*/_,!, 9)Q,5@(!KYVT(/MMA2AXWO*CJ5>Q$=0,CC@
P;C=VMF?'/MK0CU8B"S?G29?X[FC5C.]99NYT? 57;=V]^9@K>(,/JM10+P4I*JU@
PKE1G33F_%/[YORERN,<H<U9 XY':=4=YYDT1@ /YOCU8RDKDP8( J.9!;37 8X4=
PN$<);FEXY59! _(!J'.P6J764KO5DM)T:"N3[&2AT'.1M>S>SJ=(LQX"6%,.2%N>
P@+;BXE<@KX\I"^6MG# I(,\">G@FH;1>1IJ:_I>M&?2LW-Y/W@<C.B3@,.(J:T[>
PBTU2R<KCDVT^+PV'(^@@(3T@I4I?&-CC=M]1'3'&=(IQ5]$1W]3TCU?H(F&R9V(D
P*X7C7ZAQ:AP.15?>Y&#DL1^X5N]]CE5)AZPM@&U.:XM-FFQ76TO(WK@^U[X)NDFV
P7[X <L<5AP?,TQ_W\KQ)Z%!&&:;=L*-H7R$9>*4*F,ASP&9LBQ*\/IDD(_@1*[-@
P^?D=CY4H=B*"QLB8TYVSBRQ40\1#&!'QY*=Q#K7JK1L=;$]>=HFU/-@ /%V_GRW(
P_Q]-R<H1HW#W23$LC-]7\&GSU,'U$DX0M&^B/ZK-/!N;'T'?F8ABS.7NM&OY&2,]
P1LR;S"X':X(RK"VJ/P6%RY1J4DM>4BQJ^W\GQ_=/M1=!D*(6TR U.<HRA4 $Y]&/
PGN?N6;?UE&@_VM"0%&DT.P 3NN/#!96O-Y'0M_+_=#ED05V*[I9'*:P-KY)&"--0
P(8Q[("8LL^S*Y"[H:(58\LEFCAVCF&)FQW-EHSSNC*-% )?$%/@!:E%I6?K$B5N\
P(.^RJ#IYYP59#5:"82$&L'EF*4:8S^.%-YUI)L?#3$!M.^SXH2<_3:PB[2\ 6[<%
P)> DJ;:X-BG F@E:*J2?:6!POU9$,HD@/E$,CS'U,GYNW6/NE_/:(%YL)AR7;=:I
P5!W-4M\GU@MA7^NK#(/7KSC5S#/3>NM8A2>0D2NP7=5?)XHB=IUS$'3"BKN$V$71
PJ:&)H7N;'$S!U7"CA)IX9'J'5((V;RZ7"A!BT3 YV.'ZT2E^C(K9PHQ&HSW_R2ZA
P',*:S=[%2:XR-AS+];!QEAUL>[F6.=TRH\=C ^W)<UYO8*86>$7G=^,>\60)5."A
P;4^5HD(W+>''4&O=?(]XN;._TYD+AT,?'109IA(?E6=Q-&W9;REL/7\^#P9P!2;8
P!OF-]/R(:Q([WK"B&Y;G.1,!F\;CRA-VW 85QP0'2*_G]\%92&5F9G,7,.H*=,NR
PEUN+X),K,S(!8'CZ1$OW J7+W#?^B\UI?Q+SRP"/K[EY-PC7'/I];G*ND6Q> P*N
P'<ONC+(QJ[.7-3@7LLT:>N[;%/,=:IL=/U%$,%UC%E_Q.J;WF(<_2YZ8YFE[UZP/
PFL#M+7Y&H[P/CHT,[/2.&3M$Q0' =TC(,S994,D7^H,H;C6.LG+X]3;&*MF&V-7+
P0/+_KU ^%Z:H+(9Q[O]L'7^$,V-EYX$9)D@U'?,@[-7D\,,NC!><9\7]2I$>]-/7
PM8\0@NP$2CY\WI>4^3@IKNZ[$?-''%*-NM,U,L%6P&D2-P"R?0B5?_+3!8YY]_6J
P#):#KBWV0C%S?O3VG/8BTI=0?<8KW\PQU8G(FGY:U$M@ 1PP_(8/LG/1Y8%"!#:B
P8+,F=6!7Q2N(?^R%^!@(H5 M"\O.V/L[['$F[:GU:-I^R=IA7V%>QQK[@P6U'BH0
PJ'*)Y)\$4W'@! <&B@JRZ(*%J(2MU!?QWP:/ 8[<K+T:ES<0,,X<,M%+S5IZ[8"H
PL)0?^*#5Q&&H4N&]8;)^9]O_WXH!.K)D;(C:2A^^@KW]QUEGKPL%1<_!N>S^>LMB
PZ'O8O$\09JEUE FM6-S2,,2P? ?2S%@B*SGF],?C&-4#%X6OVI=\-#@PCKB7 _!E
PIE6GF9:4DL4OGXP=MY O$2=X9N, L[Z+%IL40M2=;FY!:J)/R=@G@&HOD&NA[ZX\
P6F@J:0#1^0-X9 !RA3HR>!/'0/B#XG6QY)XVA"&CYL2.81=[^D_G"D7.K"TU^[%K
PU'TNU">VO*:KC8."=!"GF9:2;J_X$;6<D>2,L"U+.P;@54S>4DT\^/BY)[_O;*OJ
PXJ/0\K4B1,H<WT7RCP^+HXKA8_HYZRE=E_F\X5K%<E3$?_#8'V4,^@1V4UYV06>E
PPBA2-\BMHC<5=QV> 7#+X^TRFJ37_*'$W%T)JMF@HU# *6-L+CE)E_!YTK-ZN.YT
PINQM._:@6DYT]@Y+*OY&>(,RZ"K+EPQ-" 651/.!MCH 9+VVG:8=[P]SAJ;' O=D
P32<*Q+#96::A(#&W4"GC-@-AY$D5*Z'D95COLVJL\0M@5]H.20-%<.9K.@3*A91&
P-[HHPR#P-X !'VR"7B^HHQF)5U[1#P3;I,7J J?1IDOU1^KT+JS_^Q/0OA[85*0<
PUSO^/!*G>,S/=?(+;WUV#A."'P=#&M^PT!^LK>.@^8<E!DY'B!+I_#PAAW5;JFW 
PZ./?Q[M,IQT4ZIH_9/8I59M90]J"/<"3;[>,:0*Q1[?&NAB<#]VD&Y3*WP"(JL_A
PJA/RZ?F$#@J@F9,: ?P)EAU#^0MZ)!4?E8#IJKK/^<B1!+L;20B XZIDFVMT6@&\
P&;AB7F0^:3;+EO7Y>N@,O&O0>_/%R#K3B63JO(:!YZV%]8/]7[[A"X6L-NS^U$_4
PM']\_%+NZ[YV$ZJ)BT=MT K;$;%C=,KO-1D,MSR?.65M-@D'F?]EM0(05#"&8$?J
P;Z_TO/"R>O=O'R';*8L0I]08_+FWWMJAE?-FH9DO IHT2$E-3I*4X ]EJ$;-)8ME
PFAF\27YVKF#.@2DC/#XFSC5JVLK/ITM('L4Y*1*PV9!^0&ZJH&_>G<6ST(I.X7(I
PE2:3]%&#'>GCI=C<>R9 ETST%]^C7'TC>AUN>: LBE(;7F02<K"6]9&'^=ZFP!RG
PNGP!G6/3?"#V[II2;TWR* V'7"-#VI2AJN%DK(D&34L-9$S.8^/) 8]Y%EEOIK@^
P[VAVM4]K:$9!@]MFZ!\3KZF1^>#I^$A;P:TX:[1O4!N*G?,]V"QK&[RA&"AI$LW7
P#.-%T,$/&/\/)_V:(:H7>S ='A'Q>@ETZ,<1\P/A#C!*10^VW<Y)#D7R%JB.N\2I
P_-&G*(&\N>F4O6EQ8AV.MQ9B>0B=^K]>^%";'(9.&S=]:,J+<1B8'W:G]+J!]=;U
PI0&@>CDV/" VX$&X]9D0<@42W:AG5YB\-H?(;QR22KK%N#U)*B510_"X 5-B!V$Q
P:I<EWK1@(Y)T</<C,(;>SXL<Q\DS,E&\Z :2:R^,=S,*53#.PO/(3AMQS7WVMS8?
P_!-SJ2![*+0DM_\D1+BFRTZI+U)3MEA@YT@W9W[CNY=>,2=6A)^DK)FARC+'BRT(
PVU!COKB^_325RU97FA^ZW=\MZM_S'%K@,>&0MT4"A]]N*&W3*9=HZ5(U@Z_F(L*K
PBZ+7+U58VPPR4PSC+GV !JVH650.G9,PL;:#[MYP?^_B.G9>=TWMFN4-!>ERG\W4
P-92#<PP/%LEUXF]N@NR"IE(70WZ\\)QC&@ 2ZQ'_S4INSGCETA;><;KNSC5YHB@)
PT\0+79 ZO-14][.GV0^MNZ9>EP."JA@Q>GXU-6#%6QCE//MZ?XL/I(TU+N WH/])
P@-BP#4@/:+,L5RCBE<L= R'Q'(0<P1T/="U[3NHY 7I <&PW!8]$T-^IBMD9]J;T
P9W/^12+_>$5QV8# F#Y09#L@.82B+DI-GK]ZA%Y)^/$+,6=H0U&#HO$+.GMDDJ-_
PRUL>O@'/>50=VSMD?92Z/,]#UT%AJL>M:O7Z&X8F;-;UM"B&RAU5C1 >5"6 I/1*
P(,07ZE[]%R_=+YF2<VMOWR=$"1CEK\Q-0X; &>[G 6B>B7 4O^2*@E$V>X.F-RSN
P!]4K#2'$\L&ZS=[&('G:MWBUKPC@<LEZ+P_HK\..$)_A9^]^9Q1B(-IX5]GS@-^F
P+[+SE82!"0X1D7^)['P]_-VO;'2G':8P=Z&1,O2X@_ PWK_4<VDP7DTV[2E%.SY*
PX6^]XWW7_#\*QM-CK0$PQNESP$D.P^+ZTTG?Q02#A]AF8@S@R.+:5PD"VM!0IS&V
PG#1@8[&D88\\YT3_IM]INM33ZU8!3+'41FW%"F6_H;(!,+K%W@SU62;D+*7$ GU3
PFD+S&P#Z"B &Z.(K?; [&QHIQN+L+WU)_GNRV7S4R-*_/U+;QM[R&_0V]0-8?LXY
P:P^JY2,5JN;F1]/ C"?5!IXWHPG*X8?IDA2J>[LAM.^)Z-",,JY2XS%D<@NG5Q'/
P)3F.MS[;(!"G[=1N2Q-;?:TF7JK>)/LQ.%$I_6WVG^Y?CIC_Q"3FY7($Q5KG? ];
P$7C08_,4@F/W*0(S2>5_\RHB)\20]2,9$A"[A2$S+1/\&0,0(8F?PH/E?Y_WM1Y7
P:>3KG7$$VF_;KV*CRB*!"(=!78C7SR*;S!:<<9DPAH-H7MPQYT[,_Q!DJ%I5P*&&
P,2#E6#5?[1+H&]9*+Y4B)SCRLW"\R\:5!G3;=?_ACCIP9R^J6$XWGY%!0#S70\+'
PF9$R=O=&;.1'[1<L_ACU$_ZY[H+\ OTYE;BSMBR_!  #]7$&?0"]=,N:]&")\52X
POX[M-88SOC>V[ 7=!1W3AKX/)&Y'S'*Z-QGC_)B# Y=S14'0J$PE]-I(GA$LC%^I
P+W&"QYFRR!NOFOWX-!D)#Q1X-=$B.=9^[0?5_7PRMI@4X$&7[(8T%F6K.X&_[DV!
PEL"T(^?K7*N<N=NA0?P+]!O'(W[X:!!$QXSD<X&NJC]A4\.CIR@W\:E&B?Y9F0>I
P,6-8O8!$UQL*#PVQ+8QTD;OR0E!)L[??U)[R!Q@')]\:<KU->O5_TFM#%U6_76+?
P)^]\*W2OC9)DF]@R6">^2I/YNS%O+5*]5<V+CP$_B%&Y?NE(_?*I6N&?8MAQ@I8[
P_7T3!P#.M<NT< HXNG]G?5CWK94]>-W//6?%:W2?9P:^)&=\SXJ)1^OU:YZA8N8_
PCW ATED![AOU Z='*%GCK+'6XWH/76 I%5,0EVI<-[+O[7&#@,B(R2Z_("_@3([K
PM-I4U=&P*9B3^*ZR&FPB(A8![]E=*"4SJ>*/IY;T53J8EN0VVWT0GR/@NTC DO!,
P0+))+-"_>O/ALG)?9UFC(8M;5;U**54$9K4H8<;+[]G;!%@>_,"!KJ"Y\; 'JW(%
PHQA[)I<3Y:%@Y)UDTJO%L8;)\HQ+C\@+TUM, [C=X*8Z_[]*5,WFRD,+*O83$*DS
P'/@&8Y+UH<D;00)V5A[M"&+6O='GV])YUT239KW.5!)OT4U3J7NTNQ&.>IJDM+N#
P:+K0&VTZ21'[QO*+'*XY/18).X'43J@2(%*]Y58QOZU;"DD'0L"\ZS\^Q0"!CB**
P2P88][]>9+$D K7C>U=TRBR$^WZ%3XQXF7$>+&>71@HO!9LQMI( 9O$+F8(:-++@
P7!P<R,'P#CTGZ>T%J7S,$L L=>UR.\62V<+<@JD6SS>S>O3M^.W!-)'S6,J&5_#O
P"(#'P<SR83@L)^RN@3&P)7H![VG]OF#O5W=$#_M:%1,^+D-D&Z'J0[XW?S)!"BM=
PAD??\X; T"L4#<,*A5CSWGNC%%# UE'T[IEF):[<E6D"<*!::\;'@3 ].>T<M#W.
P3W<.RU&K%]Z*5GZRR90J<$A@1S^Z_XFLU;?'\1E0\;+_8<?A<8&7NP86EQ.KV7'Z
P*=SG_2Z%*Q?K'T*_W-D3-P#7\;7X!SU' 1<>%QVWD)3O);:!/LJ7XFO 207O?*D:
P0HM!<13JW:X0GT:S(N4*#*V4"9%%,2+*#A ]AI'A- FK@.B035!Z(AW=/B3XOQ!A
P>VHON[>92@<WZW?SK0P8$J??O[TS_Z@6C&PD)/9+G=C:! AM;?IR*N7"<VP<9 GL
PI_4LP,[1!,9^AX6P4IROA@W IEFF^"/0G-[BKIY%MQ.S.*.WPW1/L.H''UC,LPL!
PK2]O$P R3[ID^ [O_!2 Z8R $;Z^.8XXE6(^[X%>B2(-?P7+3Z[GR;=91_/?YH\,
P-\QP'[2J@*(@(TC0_'?/:8.?]D-\':+,H^GG5R0AVBX$ELS)(=8($90<Q06\S: M
P2C62\1K?86#\G(76>,(&Y8PNUP:>>K.0O8V&:>%F)2\EA9Z/Q\0<GO \9R@CU;^ 
PNT"^.S;)KD[U(J%C2O*&V YQ;'IH4ZX5A0$]Y@O46C<#^E^Z3?81--Q#[LY%S_H0
PW4O"LHQ)G(!I,X9)/'61?<RGP)7NW2:^O'ODA:^ (4ZQ+9G .":2TVX]7^UDX4O)
P!1$_E*&7GG9@FQS()I9*3DFJQ>-[?,GT('<RT):;I)]7#^'Z)4(NLI\O1:QG2V"K
P)_HT%B1\=\D'G9T"/H<%#' ]_T<Y>1>9<_ XXA=$=C#.QGC6DLTMWN@G=U*P:L$:
P@AJ!:<SL+VSZB.K676AFY_3-%:3=RTN/<*&=(]YU@W209XJ6>35MF6B, ,L[FX<7
PDN/:4TK5 JL=Z64]RX5RMBQN55*=13R#%"B"#]FL?8A1T@+M@+6TF&7.4XZYI/!2
PL?]!7IWIQB#2 ZK>D4G;BA5I$)+-@PA^.J_1P8*+8FS]"_&X8$ =F5SB'\32MA$D
PBR#.V<F$RQ,Z_E[-R.LZZ7LRPJ>K#P?^^O$E1")!O(Z6^@J:S&%8KXLQD:\($P6I
PI-35,+$Z=";*L%^[875W(J.G=#+;6LC>B]TI<=H5]TABQ?'C [U=^(Y;/?=C<FE)
PVK:)R[\)K3#A"JSX=(3*$INMC0T&M/R"@L[I3+DG=4PL$@41W$E;*O21#R+)%K@-
PTHB51+5(][$,^[.A/ESQ;$98NA@_F1X\O#S0Q)Z",<0NR"?T!%N'2XPP3+'>E3S0
PT;C.3OTE2L.J+*YHQ,9Z,\-)$LR35H/_?(6K=+9A1@UR'-JP1B^8;C).?,K6E.ZM
P8$49HJ(G!;THO%%VYDT';NIR5/76.D6$9CYS^ZHB&WSFF14%$S"K9?5&\RE6.BYZ
PE^58(Z=F; 7.<B$N"JN2[J,9Y7BDLP%3<9B,A9).4&.)47M_-U=L!;M$NTD97%3&
P7O3%#./H$'JKI,DMCTLC<$=NDI*8E2(4==ILYHWY6P+%NA'K[]F!!,8),28K[4C7
PE=/"D@AX4NI61/VN;(U)I-/,2O@100&XXQ^%FL@5!%E<$M3WDV;-'_?,-"?+!#J2
PY[4Y/[)-@!"*GI.A^#=/ OIPFB/:&AMJ-,;RF,6Q,&+_7U5-:N_JAM9NB[0,FN_9
P,?T5$BAVM9)M%U)%E2RXOMWX<F<D_/"V9B^Y#]0F+>9(8OM3X^A8%0?9G;2>F[]4
P^P#TR6D..G1@7 7R RXJ':[!1#6HXG/GCNFQQ0D>+2.;=<5>68L8@4GXSQ]T?:FL
P*1Z0J:^U/DZ7>4\,15EBSF__X+^8*16W)S\IRU (1?*(PT[CI)W"/X$D#KPWO<:-
PHF09A\-&>B#E%(P+9+UH<\6(<<6VY(Q4CFWY,W(I45ZZ?/ -GM4[NN/#12=6X(O\
P-<W]Q>AH"3NR#9[*LL".KQ1NLNQS,Q7D#))GUBQ@<A4<Q&XB$FEO^JYWC!'D24<A
PPV*1_2L-5VJ-<L$8N/4XTG'P.[7?D6+#7@E:H),$/5/]G")9JY2<3&(!.LBX2ZAS
P&&5X,+2:0K[7]<YY]3BZ!,/R,,VV(#[3'2C<E-)4!G<I] 8C@)7I:I\O6[0:/?X]
P#FTH_4PM]*-$A/BQ88-,;$+JUQZ1UR5NH1$F-FSV5GH4OOSSF#-^%R8NAH0@1*(W
PO5N*O@PUR+U%&YQU/E5#5YA3Z:8&T*K!60A\MVH9=CDQ)G@<TZP"['U61*Y\P*N'
PE)@R]T".Y"ZLD9[$?FG'7Y0U-:6):[+3!_4'L,O&/=&G:JSQLTHN=L&%Y= *\]/S
P?EM*D@2N,<]+C(*_?A!/[IV[H7FWDELLZL/!I!3.F;@4-7V!^YJRRYLW07&T!:@<
P= NBY5DIE$I^#^.J6U<B3X.Q)I:*/SK/+/_&GPQ,M!:_<#O&,,]E3B ] !;(+7E(
PY'7\86?6;IF#84DNY9'QPZWCE]K*:JN=5F-E%(U3691H<\%PBP=Z,5Z".?<^FO79
PX4G^P%"L*I8#G]*AW\7?B(2>ZUD+W"]></V_#U&,2E2H$(5^P\1IN&\68@I.@E-2
PH!K^A,S9#2][R"LGSV*HM^NLI<-0YK$%"M8+L]@0 -C[VL($%:.7'*5DV@!G/8EN
PMX?4[RSL*#ND&/:N?N1 F0+/B@WD5(M&=PBCRU Q "FPVW=%!1K\$/X&_(-'+$Z%
PQ&O#%;N:\K<;M:LEJT&2M'<8*@/Z?&<0%D(MPD\@=A@Q2+.^6"E*D??+7:RE&I@=
P[!%W-?\69Y$=R\1MAXIOW7>E\(@8MY790['&,0<RC_'EQOR:#:&!_]+MHF-BO _-
PGPA4%5!V!>?3(?$MT3#H!3%(YBL;_<[0V%I'V& 51&5!<2JKS5OEK-(U)/.V9BTB
P,(2HFX]TX]AO[.*3DL6Z!?@Z&5)/WE!M-4-8#" M1+DZK]:V*C:CFGL8?Q/+#^7D
PEJQ":TJ_(&!PI2"<?-:=$#D@P9$ 3[/4<*4!7]"B'2R!&1;44 /Q?,RDGR^'"PO&
P]O/Y#@%*MP_#>;T]!%C&&WY*:AJZ7:&'_#8;5$-WPY=\NZ,;*3&.8RWE(*9AWJDC
P^5EB@1,4(G9%@W/(&S^#1 ?(RW8N?T.U2#45^:526#U(N:(N4A,3@ 2F_GJ#U_@#
PQ+/J?J@@BYYC9^O)JB;W),'Z/^HOSPS> I+.]M'Q\PPY='=]>:(/WA8#A/(>>F$^
P]W%?+%<O\_4<PO4<@=S*]?G:A'HYZX>.)['!",I;)\&^42M\MZX]N@I$SV8(-@N\
P<H/E;S>]F=-B0#/T'VZ[8*%G+RN.U6GN -@[],=(W$F\9/;-L07@L0C/!?;?@#!5
PU0G36#/A >T6S4[@81L)';G'MQ\:P$\0D;\Q@8\D.J=S(2XIBUE#C6@*]DBVCDP"
P3L](! _)* P@X457/$VA.MC9YW5E(^)A95 PM\RR<_ T'Y>'R]GV?<@7*]FT172F
PLD%_9^[/SOM#_ LE9E/8G.6H!EM??W!/@3-<'FQ"AX;4C(4M(D:%R2-/)Y,?NH)C
PK;MV[(%@*@$N3(R]S0Y340 CRG'/O--N\3Z[O/TM^AT'PM"MVQ58.0"FVNHHKW<S
P'M0QS9^I[^\H5OORXY;20G&F$5PVQ*B%4NGX:#'294"# %9SI?;L"#[;L59B((J+
P$K4%O'9ZF#9YK R..HM^*OFN[5\8:[XI!*+TRR,+>[[EO3:H&[XHVQ!'KE]4P^-/
P#99CFM"X-E=\])1AOL=_58K4;[M8$X)&O#R77@ TB#1.[7=!J KH#VX!!K\)7OIE
P&W?:#9^D>8@)P>#_YK#$;N*K-8J\U6TG[_/L>G5B[D&*W5ES+SY=Q,)A6>+ $U+?
PI*<[\#+$N1(5MIJ?W")I]0JA:>M&B:D[KWG:3( G( @Q:WL4K(5Y$5W$:*#-34E3
PD\1]UIU4O)L1CZJ#6B93 @0_7LU1VN8\)_(/0.Q"GF9_-A]#&K4+(,W/6S!./9_=
P_P188O]1RAOLZ/:'-X>$,]TW/^Z+[V#PR@FXWBV3/"YY#Y(0"3B<X1LH[_-K80R<
P=!UKV<EP<[.77=F9>!%FUGX)5W9U5?XL:PO" T\HW;V%Z63I5#CA%\@?9;M[])B$
PAQ/Z=>1":5)?03_53+K-CKB8U;'ANX#)B0N6I?O>W$>';WK?X55U)W57AH+>SJ->
P@4E+P<OD1]+Q+0 U=N>8Y.2C":OLZ7!HUP]ZH.B<O_K*1(\/=Q"72+QW>6.I]-)Q
PEM0:E;OY&LKMV]A <FI)D2?1=A>RQY<VCR$\$6$FTY/T__N)=4 H(+&\,=W(W+#&
PM\_X?^ >HK8"1_.2L!:(W!O0C8@(B7@<.EG06@AW!1@LHT0:#_5X3$MZ(I7R864'
PO @P.S]AFGWUM.X126I(Y3%H.CVE@5[(/1GPVXU>PSL5($-<QY76_KF?:B1=-4:F
P3V_ R?Q#N(7:@AG&B];7Y(>-#/8R+\N1&E4J7L>I\O/"@AD"3)G!MW(C&FYSL,$-
P&33@?_/8UM(>/6?>R1>4M[J4ZZ! _VQ5@_&S_"B7U4LCEA0 F4[+5#&8CW6_<$2W
PO#]AC)K.47</:L$ZE=\:^5SMX3JU Y&<7?R3-(P;A_M+PG&]QT>[)4/U=(8O547F
P4\]XHBMW[*;'U8X@#J!%]%L8+ S:6,U^_'B=.2J.$BD@1_,[:I]SV33.I:DA>0YL
PNULQ%NEFZY2*^\?I8 =5@6GV+0/&%]$-C$E2>,I/UXB<+#F ^.P&0T  :J7!S>.I
P'<[U4;9?M4/M2%4EDI*47;-^-(F](!:-:_&CG>*A1QJ3!81!,5B_ $#;?//M/6ZJ
PB7I^S^Y 53 9VZK7P;GIK &>>NA01T: K\L+Z>CW_2^!J?Y,KD5^<N?LXA]OL+#N
PT5H$X]O9V/1"?.VBCS14UK@"C[)O&<T26ZUGH=C S6:FD\-DIP?IN2S"47P1KC\W
PWQ<@6<A_>@.Z6)W>YQ1Y0\9BS.A_2\U<7J[R&'M%!\)CY/U 8V-2"":V[6Z*A*AU
P-"B;\T(M<&!2I:V#?U ?EDJ)_\Y9<4VX]ZBNX%D%EXWR']2"$H_L0XGCIEZ1$KK6
PQ,8SI3E9U0<&0!=LR9MDK7C0<7AV+VK CTUK.O\[F=_&V$:0$/$;?E-W6V.N.=7^
P/J]K%?U^0LACK,DCDYN:W?M?OQ^P5J5S3P@R6/]Q>!6<&;K"O-G08Y2+QAN/TB.M
P[6+(N;F1K-A"DF'W.FS]5R1F1M0.6;&*G4U7D6KE&G=HM(ND51%$4ZVJL<9;MZFU
PAB]E! MTU;8?@)=D(\;[4:E]BF3>UW>#840(>*]>?^+ XV!6Q>]<ZRET*D7+?7,N
P*;QC?=,KE@OOHL,N6Y_@"3HD":X:V"=#+*X#G:72QP'Y(P<-63ZP^/D 4/$7^:VY
P+<]%8B@QU9A_>)*!PO3;H?7%T:KR$_8A;T<GPU#IV%3_R^H\5GL[S*<#OH?1PQK"
PJ5ZP*^''0>K6"6Q>22_==L%L 6]*C,P;6:?4.)AH,$4>T=)I@1BY.>MF":"T8G.#
P/^_GB U=ZK3-4"/,CTW'4J!SPH88M;=:*RP^RZL_2;]XWN]*!-=LM3V^.-H(.1*>
P5%]HQN\;@M;>$8O8&0W'&14N1]0M,=D0P<1?H+A-+5'$L)4^!9>X89>*!>F:<[0Z
P<Z^JCK@\]P'!?.K;R!*Z(S\F_W2$-311,?&HHKLMDY4DJ0L#30J\;83[!7@NP1F3
PQJ7PJ\.K9)IPMDP4]O<\A6RKVKCW%(2M$D!P\"WHZB5N+L4.T:3Q*" [5EWND*0!
P-&UU ZMEC-V!W>CP<@S\R+'F"=G+X)_R,H-%NEKPU+K9)I83\;8<!,,B!V95'D1P
P0^$CCW_2]/_(?N1TZ?;/&C#K;0%:PJ=9)/@HREWGFJ3/XFFHJ6H@/ .$3LL/8MM7
P6@+9GKE%P5K_E3;J/PM.WD8X5C6U)<JF_AU_.YKD%^Z260]>45&RQKW@&R?_2V_=
P.CM-<":4HJ5WCH 5F JA=$]1&P9,+C+XG:;Q9<!!4P1(\"9X+L:)WB89%@!'4I4H
P&LPFV%S$?[WX)(\2"LAI;S 4'6"4T"!2FR- ]D)5.Y]V$*7:U4CODMN([RKO"^8'
P6*@Z@P8KY0C\6\H)_,^&Q0IN@;I8$7,;A89EFR@+ H$@X#^B=?X%[$L7O:-&E?5_
P-?.3(/ZGWE5F$QE"N0A##AIG#X*KA9]';N;[IYOOG'3^=RF=B(C@U$0O#ST@_.>*
P5UWFL2C=^Y*N*Z*I;BZVP*R?4(FGSNU *YM$YV2;0#4N)*.LZE.;NS2H=5 --HL$
P(9-<_2859,&B+4E82P!ZV'2!??Q339%S:L#1+'56TZ=<6 ]H#5+4UQ>QX("C1_5<
P)&'(2':A4L:):D'@E)V;Y:#-78GM)SF,K2#Y-)5=,+%)PDX7G#$?M?< [CVE7MIA
PB-6C8S.]10L-&/NGFZ>=PV:-GU%/37^AHE&H0Y.KC?J-"1]PICL6==.7ZOZEMV/$
P:*?JN5,M1XRTQ@YO1\<71;#P=_;]F.3WRI^KRFZ-B/R,!U#0UY%CPM".<,H# E5G
P?RPI2 <2OW>%9%-4E"%L.=H"3.?[91-6IV_:N42"";LCCI6O_P,>>[.@=S(7J2@>
P$] ;22A.VQR9#:-7D+1O'81N/?5E^[;(+2T$I-#G#$&I>1Y/,>Q&MO.O-%;1\9"S
PKU#G),Q"C%:,LJ9$?+$ZJ0"_RLEY5:.;?.X\X"O.K[YJ7I'L.[MP1F" [)Q4VMBA
P\7>10!%A8'"<Z]3MKZR?CL]36M9W8NWDG"XU^W1C$"RW'$TB<+IQ\%Z[-QTU[@4U
PWNOYT;5T1UA'>*&!Z'/2IUI#;'#F,SMKQ*YZ3K))(&]=0?021=*KZ>-DPC()K?B^
PPY <99!(.R9BQ6+[PHVSEX6N+SCC"M6&.&!Z8FN[%V=N2$;QY?&:CVF\+]\(4&D3
PC/.DL+$34+&*Z0A.F8S?M^)N;&?,]QY$!S[U91J*9+-:>M0GV&M@?]4SM'Y./IA?
P'0K#7@0.VU'25+4PPB\''LBY$L@S_Q(;*SD8E7=(YD*ORP8M>^1<R1]4Q1M8='<G
PG%/O]4O657S!(8-L6,/ZE9#2E7M"8N:'X,,:/.=1  PJCA@AKHX704; ?4]=_.!5
P@,SSXUL;P+5F5/PFI1&C?$)I!.F^?^S7-\KR$R%NR)CJ?]!OEDWD:49K]Y=Z/+@)
P:ZP8I]%XMPZX2VR"X*E%.3Z=>8_:M9FD X2]%^1I/L8.UPAC+?DSE;HJU)&<QX>%
PW:R-0;O_Q4&K-5=NS_3!/6XR8$%IRLW4T(NF;I:O@O; &)Z_W>-;P#ZH;;#.W?FD
P!'?H;?@,^U3U%^2(45\0V;?S@WK[GW**JL]!J4.Q:N(1T;@=^#HEO>Z"E8AU"L?H
P7;E$0F1O&/;LS;&E:6^*^"H.?N21PHG(L5/\0"6U0LO/JVE:])J3D#=6(B)>5"ID
P<(9\Y--9)RQ6HQ$,0+]J^8_O8>6S' 4)NVU5Y#F!19_&>"FGZ9\%V^RD(LTI=8GO
P)#:B+_N,5Y#^*?_5!/L))T>W2\ Q@8*::I2"3TL/:A>0CP&NBN+ +X?X!-+KK4SV
PNRB[#?/'*9.3W&'[5C-1SYXO!M5LB-J(!BIP-3V:XO+,,6F]\V%1X*OGF%7B'L$ 
PC,M8R%.B%,;\?L]M95A+DT0Y^UKL=WQV8LZX4O;D1@C?*].KG@EML:;BS]7**X^U
PKL6U: SLAWH0_Y'1K.4NKW%E?TE> DF@0DNS[FO0Y[LK?@E.9?D&O^";5>HM$RZ?
P,&=U, KL9?CTT,NS-+,+)>WD*M-Z/&,AH::M0E0NH-ZDE'R*TX3< $B!P"H!Z#[H
P("E>J*A.T**;Q4H68^DSFY$M.I]=/C<BXOJM#!<\1U(OU&@$^+/Y(HOPH)3<B"DG
P_K>OVYOUV'S^ 8B,PQSO^[#, '=47(CVO,Q/1MB)A\LE?#D1(X,3A0[UN";49>I-
P ++8@5+ @OG)EB)M@%JD*:LO5[PA./CM:&'*0S85PGB[?FS(>4@J9>?BK@'F"2WL
P170Q;#+,V7VX-.=?!-+WDLD;6<G*2291H_#AMJ\ ];W%82G1ER*]LOY(VK$XWEOJ
P@Z9SP,*BV*$4:Z*9CA<IR0T$Y@'*%F[GA@;>'<O==Q$"=!CLFA.*Z4F&&*#[&!]<
P4J)%).&)F,#A78XEX[L[; 4N1]5@YY!]2Y#ZOC9^91FDAT/ SO%'ZYEM)GTQ;7R6
P8P 3&.GV!5#<>&[AA^73$2V]DE30^9*#MSH[+0%+L>..^1,U!OB(O!D2D\)H/7L=
P?U%&]=:X!?EDU[]+9O',WR^"E5O'G^;VWG_ILX*[ ?[)\N,%3D#).M %&PO'SLVO
P>W>,BCC*SHZC@!P3E7(24",_&E:R7M#X!&!6+5?[)A?N&U,MR[QB'([5ZT)H^"?N
P%-Q85C;Q.J MW(!2?W=NBSIS3EV\>1/?5I >(*#=RF0F&^-$S7Z2;:Y\0U9+CE$\
P5/J-^16^D[!OB8L[)=TGI6M.40CL[,@T1W(*(8HM1C4M G-1G[6@TLC]V]T&BSAJ
PBF?MO\0F2T]$K\CG7AD4FE/3\23_P_#POD)N8!C,S*PF]\=VTR.!9V+I#<G'29\%
PKT&*^Q16=96T\<%)!JQ5!-.*U#1=J<MC' ]$F(4[T\,?^.+)6_W^9>!C:A0 :J*8
P#Z/=HQ[IQC,DQ $M??&HV5\.$!<%3 1'K$DD*_+E4>-WC4UP=D2\+<;5GF^$)UL:
PZ!^.CP;QMH2*2D?*J[#AE.\2>__O1XMH,KDP(.'+G/=/^?T?V%21MYZW8T$#,@ _
P,5B:>^2;XVA0(P%715B(G1*P,DX]JP\*K1B 67B;;XU>9HIDJPGT8^+61^;-4H*]
P)3E.9[.)(R2,R6\Y_EN>_1XU4+0_"XOYXQ3]OD 6PUT :0YW_  GW8$S7!5M^:I0
P-(<*/Y)M0XP@>?S:>#2ZKGXE[!)L;Q<]5I1)^A<FXN,;2B-N9"LZ)GZ^FI7P!V1*
PD/UYDL9S<VXCG&%8GKDH?&+^B8= 9/7UJ/B;L(.B5>RSO+7>VK6E]XIZ.!8XCE,X
P*.-XDS3;5[88H<"4CPW45T:U1J6YZW'#HCZF5U340I5(Z ,=N3C>Q!2XZ[6S,'_<
P0V<KOS!9M]U0PW^H6 -\SS+J1$NU]_]"(E!$!C\&]Z2M(J_\&I@^KTT[3SZLPN]P
P<:26URE .?6([ BV5!+4U9$N"()E^QGWW<)ZE (UJ04N6NOYRY':$]]WF^0,-4?^
P(4=+BOK60S861SE\%&>HA",RA=1@H!1!_BTAN<CT)-KIS(0XX$XTL+UOT,G[ T^3
PX3#6!\IRQ7ZX)I&HR@W%&()DGMA#0=E_&>57T[$?*$NSUJO8PH>N/#99Z\MHN'*-
P".H1P$DN_F=@UON4E2S=AQ@YW[G]B].=V20%W;(-):8P=6M5&DJY(,4J/7K&=YJS
PCR88+X("++7B_E3%4#QE](QC&9WD#M?AW.7T5G7D_=]/M*B$?Y6^))DV*TW7L'Q_
PRL7/>:QRJFL#$+@IM:OEPQG\72[8M)_8U!5@'I.Q61>:"I@*AS#?)<A!</KJK_4E
P;K02T825!^F2\Y8;IR "WRFGI=I+$3$U(*,=MX=_F[=P%BUXC)E ?2D&/OP LYG 
P$9/E)0%\5*'-HGD\.K(!FP3P)%6I07R05Q N?:E?SX%3_)7HN3$"("FJND-'3BOR
P,AL.82#]R!\>;\T4DR1"#;!A47B M7Z28 EPVJNZ;':>2O0$ "7). _&A2TMJ5&,
P$QPVCK;6O,>0WZ:(Q-#O^G&Y9(HLS+E*0<7Y[C5[Z61,F9U'&W$6\['(:YOD#BPH
PBSNOS->"VU1%-?$Z22Y]0$,/$V(:77[SYZR#397E/68D%1!KD#!U-9!%NN-T=ZO2
PS7JBY^+$Z0E .[]S -4]1)7"Y!SN=?":=NZX&>M?@2]26X\?J%,7-[K2'&Y2K\M\
PB3B&'M<QX3_:XVDZT!!R;6#"W$YY(#'C=:Y_#S7;BO@,76HY'-;.OISQ-=^K092I
PI7':4&T..B&.-F45*NQJSD??S]P"H%["&4_DJQ;*3S*7^44B%RCA0G&V&ZH"V 6&
PMF:,<#IGO?U^/_'AU;E59D<%P_0-K/^YD)]O^5G:$G@FI T3DK'/B$:*V(I"0*,Y
PE=?Z;'=B5.$PB'_9V6@PY'@?]JYW8\"F?"O<73>U&LI*([@;MTK?_+PL!K9TL[)D
PMIK1R6CK($I3X>"#@+XCS,'\C&G2EAQ&D_V/GT +4SR&Q1,Z%M1X0SRM>CR.43]\
PO 4@T2SA 'DO!W67>4;GC^78=:CM3ZPQF!".I17ZX'ORJ#F 9\\WHJR%>6\)*AS?
PH&\6>T1&>?7RI8X6&C[9N'C7M#''XS21;V1PSV6M2^O!%E>A%FT"!RTA_9FK!#^!
PDBNI]M6,I5M^>]7[WQI9XR[-CSB$?HDCP1Q]@F.(TM8S33*?Y$/T4(BK4T<O6U:1
PDWT_[L(-< 84W.MT)MT-]RS6QIHN]DU@M!&Q3Q=K$4,0Y.&86(#QV)1&TD-U1CHE
P*"\9RF&.=G<4!&F@-+]_)Y6)#M*#Z%*G]JR03Z5^E.@_C,@;!HJ*$*L;9.BT#R+@
PWQ=P"'KG8M[9;E3W;$/.#H^!V"$ 9M.F.IWD^CQL2PXVVB2I]4MC6QOYZ3(8H]UH
P6SD[?5O2AY^1>*3R?W>=XB"HA4<%1'$@=6VOH>$*#2'^C8WVN\,R,]R[2N8ZM>&,
PF5[6W+6'AQP&5;.Z7F?W;H!\:M7))_?8MRK:Y^4V)T^Q,PAA5.' [>X+4J\V@W&\
P3\OTFV"DT+.XX,<&O\J$,DA#'!1OE:)3/5)Z.$> 2V-LVC':3D@>)H;'4'$_B_]:
P?5R]0TO?_QO$GH;D^ZP5\62X 8ZR2VT&\QKVCC#_.M=@2FUSU=E$CO.R?FBM/X3$
P<()M)9P5_^^,F!M)UJ1H**AF-:Q3^0BOP_(D>>J3N<O0]^]D[^8MU/"^F"7C^*=^
PX[2BK.\]>N6AZ:^L7^4._K]$.&FKME+-A*D_/NNI7XW?(+9[ZQ,FFQO+(4YN6F" 
P4VY>3  B)]QFX!,B$D%1F#J0OLI:VY&C:;'2[0R"#]WRSS"AF@K%'*V4K+HX*(;8
PC5?='8>H\R4*,8R:E%K)->T)N+X['KS@)G5Z=6O*J*BJ6HI7@+H*3,>7RPQT%U"6
PWQE:K3CA"%#QS29@+V9C)]/B5N7'K8\RP@_[#;]R*P%$"^1P&C;1)G<_74%@W$G 
PK533J*O*I<B>^I!IO .GYHU&3.#WCL-B._ #)D#OU[F(;M$ F>L8/MY1D!UY][K.
PKZ\,#TE)F$L*B#,VC_6(O^5?Q+OTR_0L!+/WKKUW)_#\7JQM&G:6DRB;/CNU1+# 
P $>HB2EL,)$/G>H'QL @MM8/8P/V6DP?V!BD\1C#[O$KJ'>$+7Q<QE!D<I7U$#F$
PJ#^)RO7P7ZU:[]\/0MF/^8H .<NY]J^-U=MHS ?I6>C8.$7=;EJ1(:> W.FU@&^<
PS9^(ESBJ<=ZM"/YR^=-.RTLVP32-[T]Q'?-D]6IV>C\W,RK64&B/9?0;+_<^,I2>
PBQ!>-_"/G24SF"KVU3EFB8+5UPO"5^PJLXGS.FMBW2X<3#0*[#8*0!K3INQRK6Z<
PRU%4@2^<">I[>^GGI6 Y$Z\B6S;T/MCK?$CSB]CP*G#\4_TIATD"1;7C[2D ]]E 
P,=71D6F)Z+^LM/G,+'LO,EFC0D]V?-1C Z+ANB9D@F>!B_*GU "ZVJ8G/EL4VS1I
PG3 <K!8"V0'>%>16MT54,BP_0-4YF! 5<@P0C^4+!?$R!H:^%:>X1YA^VT!&I56#
P*;<_@&]/WE0Q[4!J(^:*G*2Q5F."ZZ13W;%:^\]3M,:_X$'MIVQ\0IAR3V39V_*;
P##DTI^#LL;UYS@,,_>@ U9W1O,X\:'/"96=+HRI$N/"0RB#IXB1E([Y[>LZIL.NF
PX(OU,>K'ZA=.;1SCMT"69V"H:KOOZ^$!N)721_'XK0Q?RX >G%&7?-E6G0OE55JY
P:C:V'E-2OK#S#%7$N^U<XESW U:M'+:0+(F JN.(Q?>@A(%U'0-4K'G;/#"+<5C+
PPX@)0B.L7%>F:+4+A -&7J[_MNC.:-Z-6;KU8=F5S9"Y2\QR8'? *)?$A&JL>Z';
P(181X#S]CX=>9QKPF6T//,TL@3)I@@[%H!2_!4\$J5&IJ!^/@!2023+_)O7+O$0-
P<4';AS6[2:N$EFRX<'#Y@$H>,'?P;H3!HP11*OO!86L/9RX"([:@T7V]J DLQ.@N
P] X+0]88,:JAG*GI^DZ___]<'*P-=U%:;,P$K ,W32Z&M"_ -#2&DU*+U734N\-H
P86' \93+[>;/YT REN!11I3=N^?U5T5 _+FP@LJ3^&=W@Z=KHVHV>?V/_Q32#?X2
P>_"4LHR0P5$7* YX8Q?&T-CS]!M GRS)?;Q%$]:(H/)>QLD!%K:.WIKB"61CK4+"
P]27U2KLE9(DUV>75V:/&%.[Y!$]*790>FHNZ7)E4L+0U^7+'Z)0)]&R,+_8^H8O9
P42+8M_<:VE2Y WP>$^)G:PL@?6RN<_\HX!'QH43C=S)B%(YZVGD;EUB%O\>>O6U_
PWC?B"A)2ODU.$(:(.6SAW%-/(!;_TR>%T';;&)OY#FMG80[=%:;7O(12LD)X10A8
PA"$'4NE"R"^>OZ>)QSWO!GHM7<G(351,+)=BVQIC/D6H9Z;1B!HZ&,2K70;MF2@A
PU(Y"=M6.5"PO)IX4"/ !R/MUZ5VS6/4/R1,D(:I*=V4EB&GTZ?V;-[6J8#W!7>6N
PV$VY9>Y+D483S$^E7WVC /2>@S/3I.A<-O_97=Q8(Z@' O)5/0YP]F64(M=_O%9(
PQEFHO[;L)6]$G5+&#=MF91=N1R?2_*1<.0:R\J&^I J[5-]N+6*;FS6I183CKB#R
P8YSAOH!H6:L^U[9<F!JP[W-TN]" ,^K@I;_4<C",^":SU[8VO&8CL/__3#G7#2^I
P&"<5N*5E[>5!T?:%B1Y17Z>5_\E>@CLPUL@7P/*LUUVL^B$N4N]Y$J49 Q0_?13=
PMH84H[*" T&NW5(X9FXA)AE"IA.ADZ:(,0VKAN3HF4T>[X<FJ.SH>WTE*;ORSA^?
P]HJ+ =8B<=JQ<!TMO,.OFPK\T23,0T.1-QV%TIT\.2?Q4F)\/<G\R,8>5'Z'( OG
P&*1PP((KNHZ.E5$ZX50P3E-H'Q-!68TI5#WW227B-PA8SGHP U6R&DMQTMC//;;B
PD87'XSRL'^&^.28;%W'$!]X=+7\>9GI0Y-6&AND&(%"UT"6[2[>.9UK8^(O5"^4U
P6A=3?>F#(U9%[0:NB-<K\] '6&ZO6Z=/F*_\6[:8YF^9KY7OE,(+NRK.M0<0>-#A
PPT*9H;HZ3R_=#L, 4ZC)8W:U#SY XR2(1.9E" A/&JJM/P'&P;BS!/2FH=Y3Q[VG
PF#;(>OE.%R:FCB-5KFZ_;R$JZ(+DE'WX7(8&=EO7_WLBI8,O;A7,S)HPX;"RQ)GY
PR;=FA<11<CQ'?'UW'NEF_'F$$5!^>OY!Z%T<:^P^O\M9_!)&#3HD@L2>ULVV/XUD
PEI;_N.$(++2Z5MIXXPZ/7\T#F,U4?PC1A(5$AV581$B9C[=C'PG;RX+$[BP9>Y2<
P#\C,O5A.(MR,2N(W-E)\3V1G5ALWZ1E+S^6SA9&SIF5?*ES.JF]C?V >+GL2Z,;Z
PF"RM","0Y/DVA$[%7M%M6T&!:69N>7*G+1(*6=<1+Q#TV)O=F\0T2:HRQ-/7!34+
P!TV,G)_,1W\=SQ\:*RK3SJ7;[@N*,7Z"#<'=0V NRB4.&0@9 JK>*->:ECRQ';"S
PW^5 C,N@F=>G;RG[RC4:]#+$]D_\M+ )WW8JUYBN9PR7=10K#[DI#RAI;J-B;[]]
P=/09B' D:CSV9?)>I2^06D"2<'^E3(,8.^IF5;$A40ZN9R\.A9BOG5F<WO"KG]XO
P(%CZ=,!S ^#H[WHB0*;V;X]-%Z_JGGTB.^TKG_^YXQ7)H=?B*(3MYU1(=S234,Z8
P#[LO=%NS)OX1L^:55TT.!8VJIUCT]RG2040X94U]1^D27TO3>0R%QJORW(>M(UJ7
P.,.&V+BEI\NE+,FY3(G_A141R(+Q?A]-@ZEWW!=,N5%$I/)&/G'QK-K(%W;X@NX%
PVEH+ ;E>76?3#,+X;#GSPTX]G"3N"IPMQ:26-&0\[1S,]*/)UW[^^H&VP<6,X_O4
P"O#%_$NW7 D,5H=4<(N;>!,0(5')IO=3?]*^?].Y!M-%/;(9_UZ,#YW+'O6/XS$N
P,BL_67W!T]8<,4QIO2#'SOY8D/*AXZ7(P5D#A=%7N30 5N@B]0@"5E$4\Y8.]$:/
P=(9:2$0,KG0MFCMH7",4)/]Y'[&>>478E[K9HLVN*/2<8AR5^,32O=O[,;$.=^70
PLV6=W/5*0K$'*'J^\W[%0Q'%:<B<MJ^;K('B1,=M[<&,:_Z)+A02*68V0,/@/D.U
PJ/RR'JOK,5&1'UBJD-O VX1K=;O<J= ,"70 _03D$5H1KH>MB<-BD2;\N],Y,-AQ
P RV/,@L>UR'EO-=N%0Y_!E0X;W@S$^G2WFX.Y8SOKO[J@^/ZN[]!W_>F^W^62"*@
P:5O"682J!%.N-:.75D4ET'PH15.JR95E?I^F:?A%HT*"@S^+ND6,P^BR=-R85=$)
PN,-CH:R#P2Z91O@6$3*ZAUH+1,6RN:RQG!W2^"O@&<8;^U(+>;PP2/62!FPOHF\-
P')VX=?B"X*6.L&65D-L/(I\=?P<K9EX"@)L U0!5[([+,(] AX5*')_S18-]U'(9
P4%V DW@,OH$J0$PBI_9UKV%^<MYRWZE&3P&=0[W!Z@!<M>OY^,F0CNKRJ)LWC,;?
P'3\\J+4@;@?_C!7WNA?<$^\ X&IZP4MEYMO,?8UE25/,9,.%-MWZZ34BQ(69Z@77
PB,U0+[#VC6N*.4@[\DA<0Q:EU&&Q_OEB.Y3MJ)Q"NF8F+*3V ;H0"EK?9<?**@E6
P47.T7G4EC1;2;++5-$-U[*[[19382H#N('2P,LEIMAL!4D';SOKY.7"]DIGVIDV,
P?_-.-$-*%868+PK'7US^0<$:XI5")7<2.?UYRW*H[.J,H=L'<6#PJQI\5$4DL9EX
P(JM^9ONEOU+XB4<?F#KI0!JSCH\7YC!-JF98: ?TOE#&>5ZI^0(,?-M'"U(Y;3^Y
P>Y/?5&'&3TR6O)@!_N<PO1 \$-2OXASJ*0%%:@97DGTX?%EGE:=F!O1!RZ@(3J#,
P7@F\ FC.'QG\!>+2J*FRBDUM;5*!2T^DMBM24N-]"(6 , IB-P_;2) H8HVDF\&2
P_0IFK,%BLH#:"?9QV!%V.=S>[1<7J@/G[L*Q[_HAK3'RK+D]Q2VHB!) 4N*^Y/W^
P84;/-?:Z)OX\A#TW.&5)KY^9=+&JT%B<8KE!O4-[59DWK^_ .+>?J)XK>93C0A= 
P]R-*I]_UJ/JI-HF;'7?Y'K5$A1G#?I3R1 K8N[VXWARG>U(+P'15G87,O_;:?J0W
PS-SQYM1/,*<K-Y5>>.B#+O;Q?H#7L5H/1>R&Z^"JQIS(R#X8%A!2-"EW@V8*605!
P@HOSU$,)"D)IP\G7Z'PB1HZ. &\Y)#S=P^A"8M=_2,1.V<P]0TM8#7<SEZ_3SHHQ
PP)E;",V]VEN5CP[T__-Z=F !.A,;EK(+6*%8L*1$_>I?Q7T<]5_BLD 8RA.;.V(?
P .WUS; 53!N=^8LQD+/\R'0Q\]A0Q+?X*5+S8$F&99HD$EKK?==U'PJQ@#53E?IW
P#0T.)QYJ*DM+W^$X;._"PHY\VI"8WU\IYRN[[P__Y>?$SZ\U]88A<H^Y.:NMX=Q;
P*8MX#_K#C"4/3Y!^8D91X"ULOJ=("]0)75@_]^W#R#B=3 B(Y(@9YSO=^TZ&G\>!
PL>;8.@/;'=T<:+IX8TJ#J?J?$U[PW945'*JO#'8CW/$^@G0+3P&$[ @-6$;A,5,H
PCXI]R\2_U5FX-%\> ^$K<76J8GMX#T4ZQP\%1*EDXE4K#MYR5!>99C;<!"%J Y;D
PB]'_I<KI=M^KUAE7.QY32B;;M+ U0"(\4=_(:K^66YGPO,Q/TN'& "=I"(?/FV/.
P2!4M.R1'\-FK7<27GB:Z5,IU<9F)C!**KP"%M0B=V![VQ'GZ280FZ-@0M@ZOTDZ\
P>0S1:ZY=8V9BI7JINEU\,2WWS#9!>J+\9]O9%4%_6FA<A+T\*N96]^3U 2K!GQ:H
PZY_A5-L>[GC;>:$N%<,,20AD;F%?NVWUX#(^;B8M7,]$&C^VX>Z-V!D@0+SGI]EY
PV  S-:V.EYS*CLGPA$P+<JNX==#H!$@IKY3CVZ?(B4%#5BLE.MY?B)]M.:[A1[Z!
P5Z]CV@ "2U''+O-H1SFLQ#J;_XMVU]-(01*U.5ITP"8W;\A%#+NJ1;3N *MC;1FT
PK>2O>_;=P/:T\O9W=+_:OS,/;(W^<CQ(  *OSE?Z+ADX,N]/_:$COZ&<)Y3#=6;[
PAOKAUK078-=7#>V8&M!/[&UD 'O Q, 6%V/JY0B!Z[4+>EY<>FZY2/T)0&(*Z*;.
P1Q#2G#YM/3T@K/CBCT'+)AJ:SRVS'!#ZKJ@&_&UGJ8OZ"](FE_WJ[,-O4JH7>2'A
P4.7O&YCF?GF]J8%=.BR3FL8_H_<_EJ']Y*2I@1=T:X<0(H2K(2>'UGX@.J7TU-X=
PE?5E2UX#M+2'&KY2.XV^5#I*+S3%"TY,89BLK>FQ__][C#4H6:N7[TZ9XB"1-.ZP
PQ(WQ>3RSO*%^X-C1X52MESW#;D%E;]2[KEQ_TKG(QZ&O2$LKCS/G1A'Y-GW9Z>68
PP=M0EV=WF,BQ+,6R_ F% <]4*AY;!-CSQ*M8=P\8Z6H*J[%0@)IWTIH*,_WN33[S
P_N9&^E 3P;+2-MU1JOS8=)21)S;9BYI&=%.$0GELSULAQ'5RRLS,.+'U*L1!C$_;
P> ^?J:XH10EON/7E%'B0O!I9@)NW^*%7*YG@)34=./=0OBVYIJ&*>(-R-P[Q+HCZ
P/'0\ASA&X;)AUO%;-/4%?J(GSY+NDU)YW^22IT.(<9&X:T@K4<^U@<!!PH8E%;HL
PS3)]<S';[79K9JF_GCWSY#E_;"X2WZDDK+@,8)9>+E:I)"FXU3$W(<U)%W$ _5CM
P9YFW8N-4]_((J20GJNY*W\4=(](Q&=;MRC1E6+/G)Z83,_;0]B0LW\O5;8-O^<2N
P+N6JU7_\Q)5B P.*!O0@&;#3'B<V[?6L 9NK>]<<E)O*,R_Q37'/$9E6"+BA@$'V
P=>=[,N+)[BCNOE,;S01JK_B1&+EXK-/3FH3U&@;6K1 >1ENFV[,E6,+Y8='/*Z,[
P-'0;PG MG^QU@)' #ZOIX$O28C+Z.J]T\LZL[OZ"9V_4A_-X\C97R1T7YB:##X$Q
P^Y&I?SQ3BDY1T4#Z<.FZB90,,2]H^^XLU+OJ YH08*] IK1AJ[U/V9P+V&3B)2QE
PU)M#KW(K?HWN>0[1E,A]GNC-S"J60-)MMU\4B^EY-FIEYG<2G)KOR,?69'&U181A
PC2\Y5)2+<QD[[M#2<4H(,'N#<\^"7F11,\V&F52!(C#O<8B3/NN@3/#6\;C3VE-!
P>>KLV,\ SH68Z?></A%34.#!53F5C?WNXGU<:D^)R*]R5_!U?K@#<)JL[3"TA1%2
P#V[;'A'144RWXDCB'A!)O_+"YGTHQ,>4@3&_KCY+U)(B'NGZ>@:&ATII\X:J&O/%
P-8/$"M&DM'JB #=]'<F4A3Y5N&7=*#@9+50^*]:C:TP+-NA!BC&E[ER\OCLL[*&*
P6KS0Y]E"40<D')$P_^C_TO\*CA[\9+K7//7D!**0KQ7=B=Q9/?.'B6G&>5^8Q[:]
PUX15+6$",6V;!%?NT4FMQSLLNK4/0H(>X0QE3.=6.%YDD<_>>'95_2)DF9UPG+Y8
PW\6YAL"*P;?51;"'@4AD&NKG1S+.Q*40/'TY^.%D+JH<$WOUJK9I%RHQGNAJ38B 
P"5WVLPE.*T=6*G?5^ )AR1:PEC?0%17H%6<QZ 12DV$Q[AW-FMP%J]7/.M9=>KGR
P$<TM?&2X)5DQNE$C4F\<( ?,38.GBT;<ZX1B>FB;PEI.8/BRQ]T/Q#E-0#0W]FB.
P4S$9]-K+.[)MVMM$@U>,E_9('-Z_J#4TQB=V+D8@S?X?/N':=U7<4 ;.',A876W]
P@)G(*1F]J$WN94.XTD7.7'JC;R0SPDMA\]'Q'R^3%.V/^.2F&&9'TP0]$*2U--B4
PS]/P$T+V)]UONQ)XS6!:K_)5]*ZN_\J3IXTS=9M]$+1$1S4+ZQ46WM'V-[TS]I.7
P<VIOX?7Y6?>'::&"*#G,E:W7G_R$?&@,4)7[N(<4I00U\)M'N:&2WS97C.?58L*F
PB-6?[Y\-^4<&^_JE[D-3S54#H!T?';XEB+2BJ+NOM\*,B;RH\+@HR7QA6$!15[)@
P(9DFD)\N(_.3]3[YR [6=K3FP&+26,?G,XZ9A/W=['B^# *.'DE#Z%>J81@=FLTC
P*]:AGU2J+EEX6;%M@#G\Y30N%O.;MWZM6)1GL:A^B 02NUM)PKT@4?]G:E^=6TKS
P/S?D-A34AWL]#FKCWVS0_]@Y8)C1A&=(AY<XL!PT8X]!43E^0&EMJF#;@$<Q79?B
P8/OWKHDQWT)BDJY;587RWT6&L_$]I%VGYDU+YM#-"@&44VE8.)==G]6]%UGVA[&J
P)-RJ61"I+BQP66>CTK]S5L'9[Y8B7[EDZ[L<9<#(\YQ%L*Z*IDVH#\JI=E@I;,2I
P&)V=P"AWP$OFBCB\GQB?//SC_>?&7A.A\M?Y=-A*<Y=I1<C%&O_%1:JR;D>NC(N&
PJ**J<\D*VE#>4U$?M5/_4FS\SBOH8Y.Y' D[-^B 1T%A7N-9M<BS^C,#$\RMDM3K
P !1^#;K\_A5X\MI]S^*V--:'#;"S Z&.(0(H60\[]_$(J!(Z6=1ILT;B^&3R8C)8
P!U'  <H#L+JOOJYQ'J%-?7-I:E);OE,<OWA#ZYNR>T@.W%L9#+1,2V\T@8."_'U;
P,?S^JYXFH$5$%@%TS4H80!<X_.A'RYJE1\NOFBJ:VA"F80RB#$%JU;@V/I-:_6I<
P(#'<%F]>D>GQ0!%8N! C0@F+$IE";)=W48$RY>7[46I*IFVD^!,N<*7(QPQU1>BG
PL\B,99 :(G\5#(K+X:J:YX[H.])W[W=0L<S$-R!9-Y:6I("=/"1!U=H:%2"I^037
PKYW/)A# W&QK_C )(X40.EH@BXKV 'T^GQ]0)#1\FISXM9.,''UM<'L[,0)J^31>
PS0!PH@>\GJKD9GHTJCB$*J!RXEJ&15LYZ]\E:$:ZB?3*0*8#AHQVJJY[[2E0*=F-
PL<:!B)/^2>;T#VR+U2P4]0UC&^873AI(/^LH$#@N=!=H^PC?EFIIR!85N"+3+*MD
P\<*E2>^RS]O>PYU] =GEE-8F <KE8P)KD6&'JS(@2_J^F>.&H:[I]$I$,D<AA(\;
PI0JENB4'K65P$L:[IE5T"Z3[(CZ>M6<1R9M5> AS;T*6S/ ""H::'B+_MC@404=&
PIZ<2YZ@&8[O^/4_>]$M(6YT@YN^@GK0/,Y<S+ZC[6<JX*K"=!2./[=,KR23F-9(:
PWP6J1T50%<V!I+W:ERXJK5GH$9LDU="AM5I:BP5NV3$I2["CY;$]SC>R\K;M@7UM
PL$Q0SM>,@!.=NV!__4*DI?FJ;L30RELID\!!Z]WYR-6PI0_>/QT')9L\-<K&-R?Z
PGL;@F0$NU%KT11 6[2D<!GZNPB!HDYY5#E8Z!;%<#70S9 VOZJNQ:QYO>MO\%?\H
PGBO]FK,7H$J4S$C=%+A4E]OVH^B;BIZ4]VT@99@@$26DJ8R_A18S!O-1M349KIR3
P(>5))"-IE^B=QGNP7A+7E<5F>P_)Z?7/WA!X4]$%1X\<'4M&NX]^I S-6K#>SF> 
P,\14]!C'4/61FI9GPNX'='EU,S^TW(' "R/DT.GAOF7$W$MCRR2!0!;1X.3=<UDQ
P-.%CXDGV&L%*F.K\MIYQ/C34D W"]SG6/QE*', N*B6Z<9OC36"OBH!?0DA.PD]7
P2WX,_B^Q8#8>E'1,<G^!^V@(?U(/A5BD6^;#K>YO1HOPA4?,T5NO*N?,GW,2:778
P8R.5S1-11-P&N?B+&V@C/LICA5MR'66*.9;,L@,S/H4Q.H5G&OI2-NV]=E-MEA;[
PS>@F)[*YJX@4YA>(0\L4VPVRV:C:F-+RL7IM1680#9HV< _/"&P'HP^7[HOMO(T+
PI)2QJ-\S70GQ5,Z=FX3;JTK2&Y)&=0:LO9>*K"QT3/6O2K2&H#A%(T2PQ'UP:@=$
PS?6Q\MWIIN<0=V)]&.CFIV._>L@]FA;SB81ZZO5!C@3 B,"I1S@2;,B-R&@'XVC+
PXH@-Q[N4YP;6G4>"[>&XK@B\/8$AYV'7J Q59?Z:&$@QU]IGUX$3@84LM]L>'RAU
P9:1T&$8K"-ZD:CR;KT%4L98!U#M N[VST[6+2^&/OVM0?_AFK/H]HV?7N1Q<DZ"7
P86@N'#,YY)9B9Y??EG%L-Y+-0FZ>!G94D631K@)0R?A91,",M3>#)NFU[H%7TNG\
P !M5C&<7O%_1:[5#$<<VPZ_664ST2R^[I![[V/N/K'7S3'SI"=.FP[$;"C&V+P@J
P1BG/K35FJV!R%S5BZSY:H_8KB%^A'OI,HFDPK%V1.];CZ5*&H">X\-J-:.7O@5DI
P9>)TU<[(V!^LNRX ?6JM36/Q0^):PBP_WU8;$1J8V<*Z=0@YF;RYW>%DLTD^RQ6=
P&0EYX4M6<DBUY="/V<)\?O!1UP[^Z<VY[CLDO"02:$>-6H.AGTBU>_;[D,Y81OP[
PE4CAR1$]3UE03RRW;=)]A"2G!\*,X9O!6(-9>!;[:<W%(8F .P0"UG<(3G2PR%XO
P(*Q#?+Z6@E'&T3%+:YSAS?N5=T@A;\LYPTDS= ?6_+OY?PZEU&CJ"><Q>H&.JF&A
P)1T>/0L5:^5+$>25<$1^/PD%C^JB\NMPG$'[-DZ0I2I+<6M$F!_2+OC=#PDF7^_;
P-$<P ^9KQ:QTPC:3),6NV2@55\+D#-[KHVARP]VDC11FB)"$F/U^=D#MY0#1'P%G
P_+&Q<?!9Y2DEG%8JT[@:GM7=:*?J,^]QW]\BMC)+KH( G<K'& *<PK>/*U-%I!L!
PZSIEH=2+V>4-UKH.]?&!U68>.:M.!.WFKSQ96/JKCK:$]4K0W"O60K#(\6B:[ETP
P1'.CE2*^H(>.G@+Z3L!V1:J)MW#J^F=%J-(KC?A)#HV'1L;:G(MLDNJ>9U(<%FIE
P8@ 0;U*(R><GV!%,X/]+QZWGC=W4)04@:4K&"4T\M,1.%/+NM96@#<$"^L6-[IFX
PJ!HH7Y)&G8/,6B3H2*(FIG=)P&2!L=9LK9\0\XV'738HC' 94@2W82TF[R>7 :./
PT]I9,R]]UC.FQ"G2F)Q]KVQ=T#"="6.KMR4V<X(?0^H&FX5_XO68%(D9<O- VZ?7
PQ3UQEJ[F">:R>N="F#&$"[CS$<.X$XV^[A,YNWQ:L)>[_"1NC,TGZJ?6#SF,OG7<
PACM=0/866W2(1[8Y2MR8@1<(<J]I&)_5UPWZNJ6EZJ<XQ_$%^M7$.[ +5VXZNJ[?
PK,4W9AG-@7Y87[E,-'K VWU\<GUQ=VK2,&O$E:QSFVJL9#>YVGK&\O:/?XSX/_[8
PY9^=9@<W&T3 ;>UL^_8EEU=$W*P2;#?$P@S^UQV:/KN0[\J%! =-;8,LA0O#ZWA8
PI("/"]++=[30/4"?.&TV;=)2K>_;[\9P9V\D"BP-!.$L;VG[[O,@]?(9(#8!;WQ>
PES4D087(HWD4@_W!=_2]9&HPPSM-I2R#1 "[Z3@1*O(,"GAJ$1]F@$B(JZ;;%%&G
PADJ&R(EFF)/Q_D^Y7G0TO2,./&BJ'>K$?%,=VC,_XIQ47J;]$UX!AT^@H.M;5.Z6
PEX9F=D8&(,!=C?I_A^0XYM=+5)!PMSHXN15&\1TR2.<=/1FE_7PD5=H2*1W#Q2\@
PR[*UK"N\4@R,-U+CM9D0VK @H/%?K<P;J#F3?Z(JOTE'?P_:O=V>S!O!$?($ +:+
P&QGEI7'Z:LGNP8LLM,1:W3O[CFH]CR%J<.C1U](#K8Y!=;E.J^A"1=2D]6F+#"\[
PM1!>PVL"L2&J^3$&PI7VL7$P;>)J?,Z,GF!QX^(UT(^?3-)&/+68Y166G)$ .Z_M
PB#X2$6/#$L7I59<=2L!#)NB6A!;QO,6EJ,^-OZK!5VF/MRS7J<?;IP'ZI+,4O#G7
PBUEU&8D "2?+%!,\WX@QZ/<R6RR(*C2%89E^?_@KRSX5=IC]OU1H( A2KZ%ACSQ5
P"*>*$8:5Z>0<-T[$ZC ("T*!KP[%4V2SR@85Q0W@"W7"M^1R6I(D_A9*N6GWKGT2
PH&%:UR13ZM#S7M0+5"T*%N^L4VPP0TP&E1PT+BZ'I^$B\MHJG=L*+"BM_?SI5&Z)
P,00]X/OH\3G^%IP3HWH)$DY->IE24LPSM/5'WUY& "6+'L!U!!4K2;VTBXK%]_EP
PH"(*D6H7P= 9<"K^#HEGL*\J+[:FN+T)@ATR^Y,I^YD["&8I7,@AM&6N /HR;7S4
PCWF3=:WMEW9#GG-WARIN$TN%D5C_7!AUATQIA-\$=K6;N5&+)?21PRT';Y "PH++
P/HWV":S*S, M7&,<N-PN,.()]7^KIM8E>ZZ#/5?:3K4O\M=D@G6-4.JDVPH+EFO>
P;V5?<9,'=)4X96'NKXI>G!1FVUB;J][Z-2T5C8CDU"T3>+*HL"*DCGAE(IZ_%6"8
PV%A\595-Q&6%6B18;037R#E@)D2H().9@Z[R0MO@9=9WI>G^/5&PW!@6[WJ16OFM
P'I0%E4%X&PXSB-[9@H\60 R4V&;\I)(;K+D%N_DAJ'\;(! QS<I)B716%K @BL3B
P"I]7D]L%/@"?YH.Q/XFV58SW#]FG>B*%0@G@I)H7/S/4=VPR- -^O?6S10RL08QG
PCQ@&/F]N%2CLI:KN%6BE'Y8T$[;;CR8$DX>1E=P3K[,G1>Y,0&*7ZV#;2VU *=,L
P/0A3Q$1'XTNX#AA_9J]"E+.56T&"H,%6>J10I$(+%?G:\V"GM[AS:FH%%7PB7PR<
PI,XYY.S54PHNR$YDM54CZ'.U[T##2^PU[=HT"CIY#.SB)>K:66>S8R4RFV[-/6H!
PY;7P>9;@Z=:RV^CB58T(OG%PHR]T UC.Z7=FP@#K2>2T<T^V2 1?2U@%"D#4X+(T
PLY<\S6A)5X$G-94,MJP1'PP// FR:MI2<_I20=74Z2LX(1>UGL85>F)N)H &OR/U
P+B^^2UP5<4;08MV#/LH,6Q?C$?EO24R<DRZM#@$,H9G7B%9+7HI;KR]/:99=IHFQ
PJN87$8#R^3MA1/PJ4F 0L=WRB0I;9./"%K89=-CH[>@G7)Y1D!OSQ6 %1>,EZ?,"
P3XY>&0U40=/A7N@?I#TA8TV##YEM,["<I]MK"$3_<^K:A2\T<X6>U0,E19JV,E^6
PW$4!CJ!&!@^R4 \V L^"DH!,_M_,XQ@!>OM:3E741?4MEV\(UW*7*T908G=/5VXK
P@RKY'TN2)3[KUGM+LDP.(;5C5#U, P"[B\ZS<]^C_J@TE//NL1DLC@I7+#PE2#6B
P%F,"7?NC-916\Q36@E1K=KPSI?\("O=PGQA1=7M58GA\I2GR2]&][E7@]FZ@4.1O
P?(F0[&1 *' J$>]AA7OG3@]R<L;&)BU9RTC:?@]) [R22)3X(=\Z$2ED%+PM6 RH
PM1X>%UFGC-&XM_WLU2I*KLKQR->B6\6:AK+1Q_Z[UP*A+>MB[:!:?#=5(2Y&$UF5
P\*_WY=]UV!=N9K<T#'3RKK$L$-;LQU^EC;[!-*S!E@6W3?PO78&8D<N^I1$2\H%P
PB"M8#J\7J2]I8Q1^D^A5@ R&,9:[EX?SG7(8)2):B#(7\(,V&,5>9F?4"6X="<9@
P72' O!NB(_3U9-6D4><,N25C'XY[--Z52V'.^6KKWN;B&W/^_#G&8\/B;'^PZEVQ
PT<=S-$@<DII[T6:,0GE:D :.'?$ C:QG*6#61]BOMK_]G:4)HWR.-,\5O>AV8Z=4
P,76(E9(O6SDN1,[\4%>LJW/SS[G_RJ[<+60V[D(YFD_:R)<3BK2XQD1Y,ZP/FNRS
P_; %]9O"H4X!75#.JU_VOCH,+".*3E"0]G'%%<7<N%QWD!!NSR_9C3],5-),%"$\
P%6E:7U@VT L8H!+>T+HHMKMPD]BZ?Y[(R<YD)@O_3F^V$AN.8ZYVY:D#]Y9O1;B/
P2/]#;F*XC] $_>"W^1_+R>E_\,"8/$?I^Q*&_PV?VAD#CXP1Z>:$,QNX\[E[XSH8
PZ)K[:X%A^D<<&N>\&KH[L13]:1NI"F0 PV;_J"G*-6(YN%+O(."3+4,CAJ2W_+(G
P5H^%]=GO]H\HEYI;O^P%>YC%G[K-N+=-JJWH41W*VWR)W?ASM2 /7%,CNGA1W-=L
P(3A^"[>T^A%G2;G[CB([Z8)R_A'J,\( (G'.=_H*C[+.Z.T7O &$ &\5B@:_?AU>
PGC2T=[7AT]I"P]ZVI#TEH]UU6]-^U+!Y:6+3Y:Y+=@]!4P]Z;XX'#-BE:(D7D(]S
P1S.#L7%9"B(]E36M)/6KOA<FTI :&X-FOZ44XKR+@FF,?^E2=)@W #:9_'G%.Y3^
PW$JRC/MR:0ZW;&(DC3+>2E+!M3(9T>8^07=HYR^BS-K"#BK+GV-6D!Q)KS$!<I&,
P.P0R(-"U;<U U2G%#_+GYC^LG^N!Q#D;C+7A5PGZKXS+JSQ1_FG\Y^/R[C8",4R=
P<:W$,\!%A$:JD.&SE&QVMH LYZ(5*04S78E8F"6 Q[<T!PI%S71J6R5Q4)%@BK36
P],=-:\@8SE([2S)4,;#>"URFY?53"PH'UO .R5\EUTL8Y6)(?@0,[6RH2W?,)YP]
P0>&.(S18@#&CS%A9(#78N5@/O$*U H/QNE:.?I/3]=66[T/C@=ZB&5:<MDOV9.-!
P19:KC1&]UQ#F\*MLW,"SA W/NTP/%W(:I)E28)[&GA]'ZX:IUI4?X.01*<O?]:O 
PX\4X4X93MMVQV#XD!) 4+2:.Z-P#+G5$]0DG8&F^FPHH&12N>(<QKLZIAC(;$OJA
P/5=>D+K;I29F]FAQF@=V=_GY#2<&O@% <JS?<Q@*.=91N6J]0QO2S9("--XHQ::G
PM39]U@9P$?CRAV[OIB3,(&%[C)2!)T2Y&.K@.]U6<R,G7$K > %SK5U;0G,R9]&?
PTB.5G3R&#6NU&$.T"6H'QEA6W DGXY87M0S^LD2C^)CP^!9D)[%K!L3BID>@A' 5
P3%X&%=4$.F#[1&N!KRO%2)C+EIG%.8\DBYH?VWSNC[1.8U@9 ,KXW;D&Q37WS@PV
P7I94W: F%+X],(5;3D?B%I73FLL+!@Z]SU87C?8$YGU Z5K5,<!@L2?!5657TX?)
PQ,5X359Y8JM]0HHRI&7 ?C2WQV'"D-_.?]""1?^7))->9\PIQT?]=%?@IK!M9J_U
PZ]S?5V(AJ7#"&4#D8<C%(R31'1P9E6$A+*HZ]3=?D8B[_-9H>. J@_-F9W?%WET+
P;D[L6\.?!>O,=8[4TZ2%V"'HT]7_IRW98%%+"^[29U([-U@Z"*\HG@7Y"ED#QI36
PUJ<)R0];9FJ"9^E #K?.XALHH#85J@A8'V6.IX$CQ#;:NPZW9C4W=(1?7(X9#F:S
P%(81:150\UQLK&%[+(Z,P$%G_J03?V&;]8BDKCJU;-";!/J-YZ 2DTQR=Z0E6<B%
P6X!F$RI&7-O39WOZJ4\D%A1@9-7G9;7^"")\'1^[6]_(195S >GI)/BUOM7B,Z*O
P2/7!NP6X5@BRII"<P?A)WE1*Z>_Q4%+=<9FZD4[4Q;MF.S0?Y+-4_NE-.GE)14P9
P8*"<OYSV6_;'=>F&;9>+1>,KR1>KNF.01(AF<E1GZK3IU$N^.M8MI!!R&N"*&"\ 
P @CB^N5M'=PGL(6H%3TZN?Q[*N,Z9@$2+=7DNMY)#5=$R8#M1M#&%&N.W7W;0795
P3+;@Q=2L&CU?X(=RJY,WZ'9QY+0R ;9N<AYYXC0913%_$O>_*PX,]WZ9KDWQUUA3
P-JVJ)U7!NU,QM6J@--U5@(Q7KI0>5WESO'SI;ZJ4HMZV'+L5DI4#+\Z(,4ZI2F%L
PA^:52)*1C$QKLN3QPJ\,]Y#H7#1#U\("F0DWZJ';#J3K.@N_^0<*D0B@U%&(%;-Z
PZ>1^M'$N%GQ#8.7H?J]/L1)F%5&&0/YJ6\W_DMDCW"I@DQJ9/;4F.UC-&()@:XB/
P-J6W"L.#<9]1])(<OGF4(=$)KAR51[JHC-=OE$@T_.Q?#0N9,X=^#8M5R?\L;IQ1
PA)7KTA%S8J^5(-&:T4&( /U'IBCK\#\^@H^N\Z"XFM[O<NWE:8<%>0I%.RW62X%"
P!EC4HMJ<"4;KAK280,WBS&N%#' >838MV:5:YL%)K9CY##K5;QG_##W?Y^;VP/<U
P[E;A[MO9,H-GJQMKFGBEB9S+),'6H6;)SU9*8:_\D7J6+!'C%,+SGNZ!(:2FH%+B
P^[.G(DST#7$O-YX+!6>7"S+3T^OU% =_COMMU,&]*HW^K,JF'+I-N7%M[ K_L&KR
PN%,M1([>)J]W>;/@T6N_B/EF XVJK>J[24XD)MMZQL!UF?IAG WTFTO*>20]1GVM
P_.GZ*^V]ZAV%6D\QSC$WK,F+<4HRUW)%*LS<^OT]^QXQ!YFTK]J%.@_Q8Q**+U\#
PR?>&Y[Z59X$8-+8,X]4T[,DSU;I'T1G=UZO% M(5+=]8PG^.A].%^,*#-RF9<N2(
PN>RJ(Y056C)/\ )2 !D+NSC,VJ=J:_0:< MZG;L1:\'LT39)L<\](%->L@5UQC2[
PDCU EKAEL5]DY%1#RK$TN7_38F+^QJ,,L#Q]A)7%MLUUF54O/IP@U6MCQ6"S<&GK
PT5^JV:3=@Z22>&#TW6Y@^^/Z+*76]V^7N@<?K$G($Z@7\I')^J?)*E'G]-1D[-2S
P29T/2=#/3_,I7G))FZH)4J6H#:!ET"#JL%':I2S'^;WC)[9OH9_/^U2.R\^W K: 
P4CBB0/8D_@MAZ&MHZ$=@H=!'.<F^M<L+@G_D+6(TEO)\]_%F>;*""H%1?S2E"@O0
P"<W*35A:.8%4T>";MGF _%J 5S$H9VGSB,%&I\99=JMM1.8X/]A,+],^@=FPW=<C
PQ'(@;]:FS0TWG=]K4SI\]-MIN&=]YJZC'(Q8 [J6*AV +Y?_)XLXBF(&KJK)BABV
PK +EN/ZQK6W=&DINQ)#D<F;R"[*BV=4T?SR8)868XPZW+VW*?7 7=B:;&K\%]9+E
PC_W,Q3)Y040W0X98P0(2<-Y]N_\V8);</O3)2O$CJY[9C*I@6OO!Z<Z"!_9>:/(F
PF_23@]T$W\(U0 GR?-V_06!T774Z>.^ R'M?4&\F#^@D5="W;0+3/>FL=1I"-7K=
PPG5X$<21$L)).H$Q@X<?^,:U-?^=O+/^Q810:>,AUE6T^AM)L?O";0'_0!50#Z?[
PVO,SPYDF+@T=')U>^:?DN3;;EB6C]V1&W/G<0M<^W:X,N$'>2]TDGZ(XS/_:T:Y&
P;NTG>=-QD SF'AJI$S%X*A*"5E"08@]'O++ZN6-4.(%-IDZD B?0"5%!B!&O$F0W
P(2/?R!RBVW@2#9;?0FZ?G/P)0Q>I/!L6&BVD$L!Y#:\GC< %WODP2KS8KHH#A/<H
P>1=/%O77:LQ67GT5.<>0U.94#C])ZV*NL8KM"JWADOE* 0'CC>_ )&FVT<MS2S*S
PO.0-$[_]O95GL16?"*+H&U))2$L8\@B)(.,Z;C=U#73WPAQ3,W!.@/DEZ$9\>]5<
P%(+6,H$JXB)\-B%>VH_76(=6-@+-H"7_R-_4P([^EF_K#F#$\BM>@Q  IFUQ*>5E
P$(OE1D,*A0:W08&/Y3H!&%(+G.&@Y&50;>*S :1TX)E3M!6ND3Y]2&QRPL/Q$;O$
PQOO%TEDBY7?O3Z5_+*T\C+G/TP]"S.!1/E@Z8"=L;@K9]<["ENR5GR=-JWZ*F+=9
P@XK?''^JTSN";M*!0?!AJB>QK"WJJDS:^2GK!Q_)$?K2Q(^.2J:G%>22=9_MI.X2
P4;,/#8<!\'I67A3S*MZDL2I7 4=ACRS69Z ?#N?6%B/$Z@UO/;;P1ZO NPL**$BC
P\?R.NYUC?G-<%M9N'.&FWDM'GGR@(<6Q75OZU$4[GR'UJB&,*),$7N7+\7\;^+9G
PE/&L0AG945CMNQNH]>#D$J;C<"6Z75,5=Z!$'6P>F670'*NQ68DO2E.Z,_KO#&B@
PPC7&("6D'.1LHXLN0*]T:O/[VHHO$13;1DUUL?0Y2CXU&7?HBFT_.A>#;"WDK!<O
P<Q]VR^9O3]YR'YEK"$)9EU'!G>4F,]DC917]&)Q0K@C.W#U&\#\WBK=^DN^T)L>-
P(]>4<*;T5"/&:<^(?HQ1Z<.U]3G:^+0.+KM-5T""V0KRAE#A9=IT#D=)1^A^/54O
P8<<.&9=5%C&>;GOUISS]O_""#JS4=P;(W0H+_<'X5]$'\DJ+$=;9-I),?(,/%$?8
P!2.U^J*=I!$X>B.8%\(=Q-'ZBS7L=:_$N(O-+]R@S1RXOOZ\M)X_S\A'-->O,RG)
PB>31G!WB_DV_+JJK>E&<@C!2UP- Z..156$?KS_]!,TG)U<@.C_MBULXK/!2JL[,
P$_^[P/':=C3+$GR@^_I?X?3=8UGX-GUI'C=1 #\8BV49)L'<:ROY,@;3C8S+X<K2
PS9<E^0YI)]%QUM./!F3P0WA$9TS7]S> WR9];VG$J=]4!7&)\0 S<#<L%RZ)SS?R
P8:G#(D<E6&N9J$T91GRV?E9[6PV>)!9VGM^C<4(M6!)?XV37[YD@N:361YG<N@]*
P_+4WM4YY^Q75Q>8>Q#S(WFOI%P1R[;3!#FG!#9#MN686WK]ZG,J&W].00G^E3/Y\
P(7^E^6=J 6K<C$5I16D\Y"5KDW'^G7Y[COA;*GIK5;>5);G[-EZ1S*[)F7JT7Y'K
PA> ?$4!$G0;M3_*:>E,1L#D*]A[7(AS,ZHB.LY?R]L6;MQ^/=8N0F)%N_0_RD19.
P*OV<[+EE[C%I70\I%Z^I8^"XLD5V_UQ"D,VF[<;TBD"5AE')[P^@H0=C;XJ]I%BO
P?&YX;2$!S 0-NGU_3&HTT;,((*[(>+E9( &T/PY<;.>.0 LS0_H<L!)K]H YCI5(
P/P)8X(\@3'M"(X&WN5-*J11T H 'NIH :AJE.F=;.GYXO!*EPV'41HFHBL ;\ZG]
P'%0HN&P437J"NA+6$I&P.2;Z8V32!QY5'E!Y\VN+S853LGT52V</4@VE["IO]_IZ
PDY55N9_;"L'X_(>LHJ.  %3\U)D%B"ND7[IY^=RYUS6+%QBE&HI?N=%^9U:P.H^Z
PFSN4E$_8&H::4(C%9.CST0"[;6-TJ2,4&\_ #FI*B)>M &DIBN#N!0R;5J05A5H 
P#A6MQ)!-O[.6XA$BMY:7:@S1W]^V*%"D2$.G#6L</E8$I/63C<M_LN)C47TBAP(?
P=^DPX="<(,GQ 2!L:@D<X"*OVW=<BX^C( J3N&)Z?_2%5B@7GUC- Y7X8S[U=H!L
P-"BB%?FS6GEZE:<WW1T58N>LXRM,"RIZFPI6WI+-,FK2-K*(R& G\]W_34]U1X4[
P7">_* WKP?!)5>*8W9D72*DQ"OQXM'OTV[ ]&--%!.KJ2&X1$DT[QY26<R^6A0L!
P,*:4H-JMYBI"ESC\[A\_2X=LS<B_4)RN.8"771%D,OJ<KOWXW)!A.GV3S5-[OS*!
P!B8L'TE=IF0D%9ACG2>#Q=\"6S1!BFR8&]8-+_P$/]\7@V+B(1+2$\TH#>$.\5W7
PM%/_N&I+P3%;_SSE"E#:&A17(0=:Q;=UUTSA*W-SFU /$&,\_]06Q3%S1V:MSRU-
PB"T6OE8763EH:D@P>.<'[-'@EXF;3JE(/8VU$!E#%>$^00D)71+T9LNEAI0\C #_
P<SZE;VO.Y+!0 >8 S@UK_I-KKZXSR.==B'!C%/D<[Y(;MS6E\1U1B0*V*+UT,G6Y
P@X(A=EI/Y)A,7OH\M)3,Q5_-*UHZ/U.5  :[VT.RO"'N^-!L2!I>X9_[5)7OAU=,
P>V?F8UV*J\GKJV[(7['??XB0-9KMLYH<2#8>]TX8KFC$=)\TU[;2XB%7?[]V:!-K
P3"!K(Y4!D=C/Q6;T,")CQU/03.##C]_XF+"CW($^S[0 "LM]3/S\5U6,]_P2V!(6
P03DV#A+N7LFAO.J(<U3LVI@"*U1H)\J*<(OYN_,,6/$@%=73L\O:BETT;6BD;_E:
P8O%(:O_8KZ.>92T>*B^25X5=ER,'P93!KPEMX4LP:>A2]AH($[L)E'AL6V0VY?:'
P*Y_@O89T^EB2M?4D'A[:'T!V@(S)C/N?=F>9FLI;"#2OMP[2.9.$Y)5^_D*XX!0O
PW+/$36U+>L9 PF]BFQ)Y+*U3:3C.W<94'9+UW=WC[E0?-.;[_336F$[AI2M95CX\
P-9*9FB\C75M.F8?N'?X.._R20")O7Q0XJBTL^#3IM>0/6]_"O;^"?]'E@1G%!9N0
P!.\[+@(!/6+)_@GLAPQCYN\KW8D!#>22+.DUR'[0Z+)+ZH@=W#;5;NOJ,P;@SA$V
P:IF/9VP<_9G;0M BIDTEN#GV-W8R@[YL9$60960[0NA%U/\K5,GEB@<&FTLZSUH>
PWFEM+^4_\"0ET6 _NUG0I:O--8C<%;T2*J((K4GSFYA?/&45L)<NMZLKM24['L>C
P/0"\4P5,KM@+N=L@Y1[XK@UF>1D<$L"H93ME^-T?B'/>N]FPWSB>UL[,("?>MSH]
P/3 NRJ(?.43!UXG>K=3]A]"@Y3%>VP L5ARW:(K1"A,2,KT E,7:"9F3)%):37;A
PS**9F /O1>*,2*8I_W)-L25[IT@6J;5'1=3K!V575M\&+JWN8@U'K;L!K@;S#&C2
P:]Y1:1BS2S%:0?M/MG$%2V],_B?N"+938PA@VM9D\YTSYR@+? 52;# 3I4 DM:M"
PALF%S@CKG?C)]/ L_VO5,O5"A^ZHZEBW;5%W_GST]9DY@\A3_O%?$I3@N=BE&< !
PS4!C;2;QB<X5E;HBV"2+0QYE:91B_N=>'M(IN#AW45S-[\254I3-?O[#8\3"_D=E
PY6\8S;L[KQ *.EWI]0/,=$T2C3JXVMW&8&*E7Z(\$C)=?_)K0.#<0#JE7U$!G&@2
P)U:/9_[42% 8S7/H/OGTLJ'ET(A<ML;;BY,<F#Q+(C*[.^#QB7EU#O=@C2%AE\CE
P$N2[OO_5HP/#U=W<5/C>.<GR=?$_IU=ZOH%Q-AA _7)=Y5"]#$:64*^.8Y<.5?9Y
P(TVG#0K<S)C3/V'X$BQK8'E$R>#O\22S:"8AV*_(R^:EPB7 D3%'V@*G&=&6C*)(
PT_^>BF\1?XR\D[NRP9T:ZN]'69O%6>/5W"Q,9FGC'?]=L6FQ)W/M;U2W<FR'DXU0
PG)?C?:%]O3\N/Q,^FV1HM+2$7INKA50[ $D74@Z6-E*:,%&ROA,O%]<B?:'C7S_"
PE-_CS\PPFDGR AU4Z!N 9K"H?B*HO4S;&+F[D2PN%Y4'(?!)"7ADAOY)/1E042!#
P*=OS1L:<M33X B'OP9#< OJ%644RJGN+8#"B>[QN7WEF#Y+J3&W2C,Q1#477LZBW
PDV\76HYU3]RS9Y=#C"VZB1? (ZLXLZ=5S::"X=.)U[%D)-9;^H23U(GQ)?7)7C;<
P<& LAR/XK)/D@I:*05%V)GI&2L _S.S%'6O9,TIY$2A6?[)!YBXJ,AH)Y@9#$(-D
PJ9VE<&C @-.()<H8L\]!>)G AAY\TZ:#B&LC+W?&28NM=92B47_STV2VXDOW>;0W
PR8)*1EW>CME/,P*]N.K'IX+T].P/;>"DV='3 4Y5CLH,@Y=$R9L*"S=C3;'^1ACD
P"JDG:')4/38:\0*6DA^/V#BE]_PKEY;ALC(GE*12!ZW7RSX;G%*ZG60HN*W"$3 0
P0-,K((!3EJQ15RCFTV:&KNE/#A"]#:1RVG[@7 0ZASE\SX+I51E^3.?1CBEA>QVW
P%"/[P'EN@&&WD53CQ_V;.FA)6+CAW 4C62A%+P<Q==D@*T,ZI-!.S"]]0WUX6(A;
P7UE;O55U(!<WG\(&W/UILJGH:^B^MB:*]X'+O8;\0-IXYX,6N>=R&F_"[_S?DLV3
PJ;[E-)#)C1>V?03%Z<W,,!W%2 *K[Q!JMN1D]BG^>O=KQ=N^%JY]81.?$-[SY6QH
P!:BU=<&5(_-?\I%)HD.!LV+G QH199BQC/VYD=>5"Q7<OA9V/O*H5JUJH4!N(A \
PRKB4L2-NOO-^[X?H4D )4UXD 4;XX&TK^>8^?,7PQ8"K<3U2DAZN@WB_]Q"\VTR[
PR^[ Z4;R?16JF=O"):9$T*5FM>6#(0B@A4'G';<O(.GL(/JZAEB+BM<MB@<PD\N 
PII@#@,UN;Q'E?%>8+MHG;'YNH#HI6#4I[:.9GZ!8-/A?J*88]972]=PPL@2TS+@"
PLD?\WS ZNZ+.J)C^;0]Y;X<B&,=[DN[F)C3B6S+1\V/O0;L04Z7A>A91T-8MY\E"
PSE/(+&3J4KICP!DU"RIANC*FNG=?R&NVB$6*_']\ /%?QRF.XU2:G*:,Q\_SEF^R
P_\6^;R8]3^E+JV]3J_A+5_'DFF(\*O 4AD'C 9B]@+YE011 8U@ 7(>,)4#9M[)=
PB"(!3H96B/>!_MIMG<PHVXZW%>?7.3_V[,8/5V)F4IOE@H*G)U@*F1L!2]6IO7X?
P#"02CEWGMA@GR(7)YG3#(TDFV;8-F6E$/=T@8J]=OKC]("YU$^BAK97!$83 7"Z=
PF(42(\,L4M#VMSG,T=SB]V^%SZ-/,-"<V]=5I8H9[ U'<Y,[98/(]C'DM*'4X 8.
P/-):TX1OSP[0)0M)X]0C!ORF8-A/=?%>1Z$C-CX#H!:7\8]=&]?.RRJ'%22#3LSM
P%SM1FZX3/T(0;-1M2I$B&NH4-;*MPYCT4ZTQ*8.GBYR_7FY1%#0W F-LZO5DDD1N
PJ<6FXG523J(CN/N/99@!;;LG)/0,GX&SJ-[+B.'KYC+\F!&N5T)NS]O6FT%)G.<G
PF%%G_$%X0OEV=SYK:*AC6R20:9(X*,!C/X8 H6NW: +/:LKK;2>X<6Q:% YDIL-L
P<RYJ4,/*6D3\S&NE<@S:WL[18WYK=#$=$.IMJU/K'[D0 E8I3-$[$Q38416*/5_S
PN]=\RPG[7X\HG>_;_TXTU:: &FK^'JG#7A:WNRFI#N+YP:I,V 7/QO"OX5Q6RX:W
P/?:*NZH<?&IPFE,*QH-%5?)T@/ 9" >%C(:8P[S7#-;6ZUH],4ZB<"#WS.P04+A;
P$*4'Y'+)<81IO:1,3VNF(,G[1Y3AK9;01CA$65H.&SG]GO_Q "3RN"AD%4D9<\Q#
P3=]\(>/?<]K?@ F:"]9%Q[@+U&A=[%!=$V+N'9_L&RV_9LGU[\)V@"B?;7)O/!;C
PM-.>\;6=->P;H[;%,:B:,1CBN*'I/'J)I5ZTPG+.4B0,D9^2^:L/,:8G1QQ;17-]
P3S9T/?E]SKJ8FH2:CYVU>9+<#KW$2O*Z8Z:?F7PK09-1V&8IH\FOD!<$"@R75H#+
P)NO4^,.!@;.F;@Q4PF3["5,%UXZ44KJ(L=!4BT+6M;1)&TS,@HLI'=7FRA 1S(()
P-!J-U[+$"PJ:_FP5G4YA1O@@@##E&;UT[(UX:4(,=OSPQB?TWYOM0LM1M%FZ#<GI
PDB]RZGN,2,EEWI ^<T+HA^RXX=F+(R!.Y9U&?3B:8]C<3%EVRW 93#W$S>,?LA6_
P(ZEIJ D8X'_BFU',:!]Y<%^'Z=.!#^-9TJD2M^%INA4?9'DKFCO7ESL*%G0H)0_/
P?35;ISY=0($.2OR)!WH3D%C6LJW^1.:G_S&QC$[YT(C\C7C1_PAT=D2'ZAF 9JC.
P*KEN^QWZLL@VT5MLEB,![(YA'W&0Y-2[>3083DD55;WME;$5EPE>8_,UM0:]J'S:
PP:F8)#A=#/^!QULC]@VK7"N;1U:,^!6E/I5]DH**.36BC ?L\5\,P0'?V9$NC^>E
PZ5IL8X!_0*$#QQ3;%<J>E<4A0$*.\6TL('@F (4<Y2,DN[C1:U4^@ZDJRF^+0L[)
P\V9FR2>1YI$UI7]]C@VM@K6+QZR6$XKO4Q6@=T.B>]94;'AE0D<MCE31GN9-A##4
PVLN.B5=J$$N<=D3E>(#=TLV51\M$KHJE[#$7T\@8K KOD^:,U=AQP,1A2R,3SI.!
PB_3IE?>4%^J8"BOS)LR[KC;N7)Y"THYK%V'2X73)/JMJ NH=C-']Y&Y7NQ8A(V^*
P2:H@.[K,5I>I&FBW\:07O^8/?/C#/.PE/V0@-G:GJ&E889- Q>.#Y<9N*JH:U<5U
P^^^>0_4MH?-HX5GDRR:<T[0K6:;J^0-X]MG/ OEGB+J^C*/5O&W)1=Y,H &GPF8*
PE*>)%56'*)0 +=A5I2QF(4H^+X=$<V6;[%\/ CCX[/)2J<%U'@MJ!M_XV[P$;5P.
PP>_[<_T+#DZR0A]ZVB[/3XY.I_@ZI1JYF-"&^*9"T_DR%RB\+Y1Z:C/@O>Q9K1[^
P<)TD^P5813PD*5M:*P#O\ %I/3V%<+Z=^E<N[QC6POF-UI<MXF5)"*X3-WNY?#'*
P+A7VF;PAT</9&R^4E>"X9#']4!S%F&,A=W%.4!5:*:38/JE% 5C;^7X?WI[(F/^[
PVX#IL46D4+4"G?^;ED,,5!!<Q],L2>U$EFU)3LD?0.>8^.&XHDS Z)J%+S$\\SJ^
P()WDD=[DN5HT%'ODC^IKA74J>4[Y2)]A@.F82:RK7RT^"_A/<IFO2KNYU/"$K;:Q
PJ5H^,CK(R*4\JH?1*EDF93C3U]6Y*36MGA'BJ$38?_@&,=M&C"QG\:C=I;=LZ+G%
P4/KW819G^6R1$6'@-!".,;-E@WI$:9-1TB))9:\+0RF"_02&J6/:+7(M%NED9@^_
P7!^(ZIZ?6Y%^#<&Z".N$!ZBB7?)P\-H5;=;1=+?G(&K9'_N,%0OQ6/EQP3M^K4?J
P64K! C,D;^826=#O5 G1/;GN"MRBI@42P+=5UD[GJ>2&SJI<PA9[5XISHB[8IC6H
PMR;46$:1]2X.A23!W6JCS/MP!2%14Z+;J&CGU+J^?!DY6.AF@(3XC]1DO%6/PZ9V
PD$Y-W_\!\.3EPX/@"RQ=S:ZG/)O_\)^@8%>FR]U([_>F;&2:;%?9= %LD]\P9E!K
P1$%6=62FWC@CG!XH(:POLQ6/5E=_84DC4O>I3@U3O"W1M[;BPR39V7O]TP9/;BH/
PQ>>SMQ\F#XWF$-(SQ*).Q2 &$>TC3UC6II\BB<LF74N13<RSGS',(]9KB@\98;90
PCPU>:F1>Q*KIAN2%C*"],Z4INE?D!!LN0ZL>*:FY0,DGW[;.WU2/&-E3/(3,C%=Y
P0D\)S7UW3$090)CZ\Z\E;>!R>X1B9?*PA"!CS/DHFM,$\BL+L_=E===(DL#!5VW1
PN:EX_K\$L6'<>;7-DU%47*.)0UKP\?DL))F_<%^WL':7'A6@QT!3F= 0)IE6>4]^
PV 93BM1?!U?]SHVTB!99P40B&>>19+QL*F_ZKV0V5SHCZ *=G#5XY=C,_%9AO_LN
P,8QJT2A0+$BRWPY@"GS&8FW2,^HA+>X4?Z3>?1 3>;S?@PQPYU/'IL PD'H%TU$ 
P;WK^WB"'TT(*?]6/>K>4YQZ$]?+SD<ZJ0+SVT=I"U7U-;CQ&>PE^#_AV+-]\!YP,
PD-CK,XB-N)+Y< 48Z-;T%AH,)CCE91P^I0)%.].#H'3TRF9A';NY%JL $;3O*_=W
PA6F_YU\1]\<'E9::9&]0M8)A-2;^^-K#BHH*Z(W>V^F$:<V8$)1/^W]J@R=-!=.:
P,81;5MK3F9*GSHUKWO]9?+\D_E;R)/YC'UYL8DUY_\(8]#[<\U8SR" MD7 6^_<&
PQ+7<M?&B(F%N!)$R@/73M')WQGT*?:%;XZ2@GTN5M!N:('4\"3!PVM I5%O>Q$EH
PU9G3..AO]*06">K(N0@V#T]_V! 8^D-!>2C;#H?%[?>C99B(&6EIC7ER /LNT&60
P24W.]+Y(Q]#X2!4C=E,I:]MC) ^UYW_7\H_1U>ML?FK;IR:/!>F]?=@DLQ (2\UI
PB^")\(]R</NO*(K=?R(T -I&-3NG]R,D'NP]09 R-;9(U+E.IE2LV*?M#?0&0N.G
P4R)MG3J-9.7M^+N7\!9J"T\#"=X&U?',HD;]4)7R[^EMM@S@:8WEM[38W?(0_*76
PV^K2-%M:WHR<?=9<4O90P1-7U!>MODLL,W:"66"*('W>V0@8:N,)A!W=FO7]-PRK
PNOI6 NE=YR+(T5VQL(0@(836'Y%$Z'[O\/:V88>.5\A]N"HA@%.&W&@H-6BWKL=1
PHS"8F)[SO8R>X8$JDD8%"&H385NC2-IPVM)[FP]D$>Z(6N?@OX^%<PMN>.=>994R
P]\YY+33,_FK99H\-.HC,N;-K[^P"C-ENALM$S/3"M2%I/G2OS$R'\?OH&]892'5<
POJY1<)^H(>QX[V-VH2-=A>RQ]O-^]FPWKBD7<PQU=NPJ*0>E,2'$P]+IB.WZUD9G
PE+DD"/.TF[S4B!Y]83T:"WXR^Z!X&^S>W CIH" @*'R6\HVPGG>#][6\S/797F58
PC4CT8AZ27'NK/H)')%VW4.D^TLZE:9:GW/6TQ48LO!X$1;M2YQUD<3?,T-/0QT;K
PIJX%?6U6014B9P]"5B)?] S!J$82OOP(M3:Y)+]1-B<TT%BBX8%)7^@&S5[X519!
PU/TJ_G:^%-P)/07_L:XE8HTX&D2^?AW^N^CH LQM?8'EICPJL!'A..HZ8(:/AGR+
P*?Q#3X&?G_6\79K=U$_!5WFDB;H%G1*]X)U!&77-F^5K<G=DLV_61XZ#P>BTH(!6
P#M"IG*1_E'PY?%<MI-],P <>8TE%VW1$?67Z9AN/17>2/4I2<*B+S27%UVS;1 P)
PSOFX':8'IF]#JG]LK6_$>F&8/B*/AP^<9HJ\A\3OBP.">R'\2F2Y^Y(1"SM:%,^Z
P #+(8LO#_TQ<Y7Y$<ICNZ^09#R8;P"TV46;?.H)ES-ATF?5[U@OYR:@HMYG!+@W;
P'*9VR>^!GB2AKO\)F J:/_"YPLXBBL A?'Z0-ZP60BC 5W(ERWP<O$]\1DK?GI4D
P*PJ/O1E?!G)#8Z#GK%!QL9J,B?$YTWD;&:@1 E_3HF!T XH.:_:H&R<]#_L/"+BQ
P46AAQ_R/TOY RO2+ 9@"55AYW&^L)A^W#PQ)O.)0<(V!,:A+W&&*.ZHL11"M0'\@
PG.7E8U\54NV?H0AH$5_NHBJ.8M@)Y*<K+K1J;D#"K1%9^+"!@_V^AM!%F'X[CF$L
P>M:['472):>56A\4<">HZ*.;>\?U/(FGM9KE"'4/=/R<0\>\L+SH<FPXU+L0^(40
PA*I R4O20.S^RS-5_]>U'GYP*I+Y9VW0WUOH:WLK$0@,33)B^%T)YTCZ3;<U>7ZW
P[\ WP9--H8@D)O*/,O>C_(TY(/F1DI1>JS<^+C /W;_",+QHI]&ENXTR4B.ZAY7\
P(>_LN)Y@'@'5MY>?HF)PEPCG77@;FU%FK@>)@]14G;TFC&?SMOU4<.)P^HFQRC\0
P3B.K(EC]I+WL? VY_!D(4#LI@422DE[IF?Z>.LL64R>B/75W,-R? 8&E *DH_S2T
P)\9(4U.?98^( V1?NU7DO_5!)@V,^ACC2,IY-R?/\53 @/.#?345=K1@9K$RS;CM
P*_=O438KZP._ASCQUK634%&5F)E!$]K-B 1Y6_3MD\3\])L#7I%B=5V+G*J80XP4
P[%RA R6X6&6P^CO@T5?U=6:=_ N+N93&\BDS+=D,-!-SZ<>[2A7N2E\JI1Q_(E2#
P=@,/(NYG8>U \DI4V<$[Z2,B^700<](W8H37-\Q+ED]<+6MVWPR^&%0/_:5>6P((
P>Y]XM+:5)M!71M752;Q6YGEO1^NR63A?X:).P2,4)#K?HR(H]-C+(%)A&+0P=]X2
P+0S.]!0Q9V;-*YA(ZE.8A@UG'ZK99PE4(54,$D07(QBE\OFMF@OQ_$JUFD>]!'R@
P>[5[G^/K#UR<[#\&&CJWNSC++5Z&.:4D/L@!A8VJ0$5@:D4$LV2$#QF6\6^AR8S3
PP7&2BYAT"-RSC08XBJ&^CTUO%+8?Y*5CZ*-)Y4\SUZ/JU(SYO1@3L&%TQ\14A%FU
P/[?J.</[?AGH11+ZCA>^-<[H/7"VA@3;826QG7'>HI_GHKO@>_'6.,0B]] ONM'O
P"^2T= ;^*?=8Y2U=#Z=^IR)E(@>K0]D,.='^2H<28A_N]Z+70DA&03GE@]%R/V5C
P$(3*,8LGS',LXNNJ7,#HAA=K$#B<5_O)OT.02U$<DDJ>UNQ G5[:)8Y]C$;T6LY9
PV%81[0F,>>N'*N_:O\=>';VV=^K2)0X%@^_L_X.R57XSYO726Y@8GR>U1J+KZ^5^
PXFC,+S?OD:S7Z!T EM!^04L&<*\9-H7-M4'-GY)['?*<0*&J1SJJ&>M:=H-16:7U
P&5( 8)>%Z*RS$#'^JBK(]=W[$Z53\]S$4#X@#;JQ=A6PW09=BN0LF6IZJX#]+7\!
PQP<I7&35-T<1?P#-N=)[Z'&49WT&-PX._WO8IH!U$81^T\%7LKO5\G6V-RE/#>&$
PG"E'#&JX _TX*6(52#]U5V WL@(V!5:%)-+CMLO\G\_0ZSFG&P87UP20R'&[*_5D
P@"GM'$2S=1PYP2MLW<>^H]0[PLE2*G7CF_20 S@8GH#8EH#\-R ?=$-&<8K-:>J)
P0 #[&N!.X())N//D_2I1>87-#;Y=PDDB"J"\P(D'?\!RLI;U(K">&.*'_&SF)O2L
PFSX/12J!,9FI52@1HM\6VCX?;A,IU'MS1'Z_N_0 =@)_32'N#Y$W*1+PRH\9,<"F
PY_LK&*BJ8'7:!.',!ZRA,@7+/&T M4!9U=5:,>:<#&&,M^'OV'?"]DO+3X06X%+7
P/_XV(88>SL"!\-5IKQDPUT30I1"7XE^ QE/]K=Z2 3JM(H@D(5HM^@"QTA>X"4E*
P=+B-S?FU9HND&[>.=EGM.=:'LE6D=3ZG;K(.:5,Z5NHSP8,+0J=ZG,F\L3#[5P;<
P8!Z#&.A>#-%<EW*R&_V+-S-BH',4+FH3Q!0^IV*^(+DS-IT?67V%.03A,J0C\.O#
P)SI!B.4SYX>E93[M!_[??N 5?QX<<A)TP*V4<ZZ&Q=74Z *N],;(TCN6P 2!3/<I
P1  @C$-HPP;QVS'[$3]A+;**=+/U3.<>>D?6$3L*)B[%>$SQ#67!S=I104N5*N.6
P6']DFCY[?BQM-<A_6]*:XJZ=OAJ>A14!9T68C3&;4&D/6JMA0&.R1:KY"JR)^QWA
P G+Q"P"UF1&F7]ABWP,AG5-L8S)[KYXI"WPT2P>E33?]-7[RSO92;4E6.&L"%\^:
P\C0@R(9F5>-5!<IVP'C'W0K_[EU'C-P*"+FLH!8?RDOQ&4*->?CK8W6\QAT +>(B
P&+,YW^#RU#0\WT>.F@BB)&2OT>+$RH2*IZ@KMPV]LX <,R6?@-FLM,Q)%%I^AM6<
P?I=$$]&H=0:"!*S?V\CH/DSAJR*S@;226O*Y6B 9^38@$0/A]B&$(+#P-M$,;!+D
P/N/E;%:A=7?2>'8#[[-)$N]/,-69[UC:WK%-E )H2D( OH-%^<V69J&6EGHKK W<
P%U7LEP'@:F:YCFF)<+^^KZY)86KFU7^)[8/[Y24@U]D(V*1[,  O5^$RHGTI&%BP
PF",=7M,?TC:PM8;<#JK0'/J[-=UJOD6O6$O;[V=DM@:J%#ZP8F 3T=W\;I#NU\<I
PJ*_VF!(BI61M  >8P-G2)R?ZQ;Q4'F3W%V11PPW_RQOU #K\KF>6M[0ZY#-+PYH3
P2LIX@WC6)XHNU75 29XVJ4>>:Y3QU#>1I.;'CZ>*I_.9Q25"62L=-29"!U_&]!=_
PL;+>I6OB-A,-S5C[Q3PR4I$%+/1J(,>\D<&S35DW/PHQM!;P^LX^1&UPJ&M?D5Y?
PTMY:'%-T/#U6:1C_)BE5!**(^+F^0F$M0,.2/ABO%0;/?C*.NQ&^S-+],A\0^==A
P!]=;HS7;*Q5P$R6;\;1.A<-2915W/$U["#4A?;/D&^UFG]R#DL+15) 5B&V:E^'[
P*OQ(0?=(,=_:KX"NDYV5/LSVV#'7_9 6J%$OTQMK4>:D\@>T*FUA55@X4OBE!23 
PRS% CD,FUNRJQM98 \UTZ9U$*OG17.F0(%9?)R>>;-ZIZNWVK;9WM"<S#(*6-/^:
PD)?=%^*+D=-*=;S.A(N))B%(\8FJ5\"6WTPG#Q,/)&4,@[HC6D]+4%SATLK5S\K-
P;ZU12&EC.$9#R7<9+D'^C0>F\'@N=B0T8OF"=[/KT_3_7 +^\H/U/>JR_NLC,0JE
PGY#"8')]K#RL?8IZ5 S/E^>;H[EEG=@NVN7JH;2BWDS_,-[OO;Y<\(U?=(<:M//%
PTP(#IE62 M#G<Q"PXHC\5O :CM9VS<@Y],^(LJZ7+L_ATJ7_['Z43-M LY(AKJ#N
PM%L<BJH$F!8.5,6]HIV"P:8YF92VF,J 317=<T8IECJ[0\,^]H?4?*0Y_5ZDYR0K
PW,'TSP,P.X:R+3XJ %8+(CNV5 L;O^/Z*N([V^'PG&^"Z@(+&4!PL$Y7&544)$4\
P+$#=KA%-E">)>&+'K-7N93*\ZE<)RNJ#DUD:#EL\/HD=O.@#A9/>LX<"D+*6%LX+
P22=O)'?'SQ:EH%?9S262MR?4*O/= VH)X#H2P'=G]2#L<0FB>?\ _DQ;QJ,BAA+F
PO0(BF.?*Q3F&.J1P<0@GU3"ARY?H$JG5$R_LM31'G53TNYVNMH2:8)68+12LOAU6
P3=Y;@<67>>=KT$7 OFC&DXU;-.Q9?":EK%I3 0:#6O#!'RR1(V+"TN9!4<MQNLK1
PE.@65#VHPX%D2_V*2*!R=NE*CN/Z2+<?<N!(%X/H80>04@[<1KVUE*T[\_8#O&*)
PN_EF>7W)!*2+;T*S77OVNT@^3(U@)3AC5J%D&H6--.,)96-6T_>0/L>S$1@\WM^^
P\ATC7!6ER-V1I+8[-W7BW**Y<\)YUB_ XU94=U5FAZS[^]F.9:*9IR$BTTF.:F04
P@5^Y;@$/OI#M@J2*I:0JC>E:V:.1^,HL%F(O(O=8/7C$K<<34D("#'!C/AOU3&<K
PW#18.<ZF$?ZR--WL7&_XWWZ6A224+/>=G"?O&F#5CO6SJ5TMEZ=CBU?Z*^QDH(2V
PWL#0\LB=P^QO=WNWVPGQZ&-7(LY7,8N#IYW?6:MX,71Q1^B\C4UR02JYL*!@$HT?
P#K&\1_<Q5DQ:AR-@0#MU&UL"1O1(SY*4HR,WDTT5[>=N1XUVYC#AU=J6U*>Q/0N4
P[E<5E!A!7RWQ21?XVJG\:AIDZO_Y#,P0C\]\M^E;!TZR,Y#%1BYX$:K2BRR'#$A1
PU&[D)),,!Z*1%047'CI <#[#8NH@M;0-Z?.U6);14_QRB#([-DSV8L#$CR5J8E*A
P-HQB4_)8K4.09[835X//:IJ")X,"I>X8=E>*1GS*FA<!?Y),A7RSZ>2'Q#AI;^LD
P T'"WWWG KBWTJHP[D$H=>-VN2B+]VD0BZC>F"!18$15!31L.BRGC\]!70(%X7,"
PP3;\C[[J"<GO0I]2W(U:Y[-,M&LRD7(X"4X!%^FI0UMMM5RY&OCL5[(WD/_W>HW-
P8Q/IF'7$PD[!U2%,]6'!^0, !B-,"2PY 00"D7$I6U[I4X)9FOM( EL!C+%,35F.
P6]-%QDC=G#"%M?DX^1 6T<Z_UA-_JUAM2#[*)'&:H3"-_O\ J7#"E=H[W!.;#45=
P0=TM[=H@"HE%Z'K=>.45VX8P4GIA 0QM-OIIZ84@(_EM8CJ4:96P'"=3SCMFS3'Q
P#;I1#/^R$][NH!>R(HG,(1_#"+7SG[I-L)'E3S&)/@_WEXRV^NV JT?(NOT4TR&(
P7Z!C@X!8?5=WE;L#:O_->M;M"[.6L;[Q20*N4G0BYKB3*BS] #&<VHD+Y1DG45I#
P2;3H:K33D"OT%*O]?O2XLQ]MN42C-'T-42#'O[G,Y1YS&> LGZ\PD&I[TE,RP3G?
PJ>*O%NFBN!6O(E+I4J#-S95%]?6UE.Z:6S=S$B<S^Y/>*#@](A14&>W'?_BQ6J!U
P2W RYD'CL23.F>D?T$; %FKRY*AV?![%9$4^/S*#]:Q#G 8I3*IL:G'F6C.\"\+3
PUP*5ND,G[>3.:,AYV3AQ5+<BPH6;"NXXZJ.O4E3CYR>=:_T>3T)/2XCB>Y]#G0:L
P-;I[Q !@$W_G=.L?[8K#4Z=OGY/1$@M4?'>+1=O98 L7G#WC+\/H36\-F.3/!BG_
P#-Z9PFNX24NFX[:HX0]-@(2L1'\^ CQV=[:\G$731!7J"]S(KW?'<)M>SW9^KC2U
P)"_=@CRR-;I#-P%^=WK-X8#GY#F/E,[!W['.0WBF@;P4W'8SE%V-.Y2JWAPPR'I0
P\L_?I'=J'O&RBR7.K-89Q,R%$,4NFF-)-YO.7G&@":#A;$9RS^Z%6C*B'E//,O)^
P-?,&C>:ZHD6F"W$I!#W8C%OH?QCR.ON)@SJ^+4 879^4Z6?\D($FFTF-D=#$,"BM
P'F]_Z@*SXLY]DX-\.Y.=-]?;2(+4)]VO7]^K2NL !-!2MBXU%FG8#O6(52JK<H>>
P2P_.N@4COF:1)-2S>LTN@%X9UNWG] L6*.#H[HU\[H]("OC0X),$WX)[T^6Y'(*2
P"Q" )S%:)\$OJ;/S,@+5R!.A"=9!LXMX^ 1/*J=U5T84=4/#&=R 7ZI]]:]UOVU<
PG5 +4_1ONN.=SOGD,(&P8,96SD!["$ZD/OEDC][R\F.VPW<Q^U"-*1 $7-U.9;')
PPCM?JNVWA<%$$1+3Y^1.-CE3\-+>5%1"1=(F(;VA$[0KH4IB=H"XG$PW%L%+NX$2
P^C?!65@/AH5N55D0,X(*)T\1]"1Y&7,B6+2X_Z[("S?6[IK5JBU4KK6DTA*;%/US
P4TZ/->]R3(QSU-0UP?+B5H-\^.E:-W;=Z@!1K&A[6\:+8)@\YY?ONZ+4WC;A$PH2
P$48S^+>F.:MGL))JF%YE,\$\;E'PW\@48X]V>7#O4,4R8_'@].R'4KH+KUGFQ=II
P;BPX_&$80Q5HMHM[O":(:'0N6F9O<B0_;Y)74P]!H^H1Z8>Y+J.U>++\F0'7X3G8
PO:B6&>?E^]F-HG\131^3X"-8Y4+5/,*PUDP/R>?1:D^IP=%AX36:W,N?KY.7KS,C
P,.A*6DM33'MFS18RL!:U;H8ZPSP<(JAKT*:S6O*,8,G;,O1 N&=Q<[/^#M-BWX0B
P'XAR_P/.E8A11A<%I:"38$_#9P9T:IK.B_JB>%;N%@VHP.>75H_FF!/YADI7_3?B
P8X\)?AN<BN,B]]14!XZR?;68\LHF!1!L '?3:-O.4\,+E/RF[.X*=]>*_!_KP67V
P-,D]%[D^ VSP36T I=&!#MPJ]"/[ ,[L">WT(_;].8>LX=S')I>;1'(!FAK6;>]!
P<D>JY-S7]S:GAT)07W%,I!E\!:8)#ZHO2^,@&:4;3N'=Y<(QW)30Q'A@:2TR XZI
P6\-9B;3/HV73&)-CQ$DV=CJ_8.JY;.6)(;"*6+>!W*P>&4W9<.GO"IZ O2<Y>MAU
P(1?V$<3!F <(9$E1N\/>:T> H$'Z#OEFP5;<7AE"K8/>_6!?:871',!YMC0RPOGF
P;Q(<!-H;6T:#:F",^ZOA]J_'\UB,U8_)&N40[[OXPVQ]*)[JF:+4X"C -<8: UG^
PG<1G_#%$7&L2W1:;@5V$B5(\:'MI^:E-EA"0*[2%,4T8E(^LV\[X';N?X@=5X51X
P:]_>#@YRR-LA68HNM_P/[N<^+#H:WWPWSZ FL\'W;WBW<><A4+Z5@-MSZ[BUO.<Y
PV64/6K+HSI-,H7B4'X"7?4W+.&'XR['$&U6U)&-/02MDRQ\&\ZDH3$'$]6J \%_N
P_J'5^5=1W0J A3L4HLW$]"..PC!6')$V2F]3IP *TY/[XM0"-'_<-\#$CF9Q\,PN
P K:?CM2;9454P77V$-B#M_Q953OSR$?)?A#@&$Y+6 \:N@8ZAPBFYI]PJ@MUQ*<9
P2,(@Q#KC!67NGO_G$:0X_N&#AI<8VI+>B)O@^#WKP-V&/=Z/B0_?H/,S"=K0[2@)
POPQP.JO;O.+QB*1"G@9WATWVGY6&4 O846)8RYR_*^C7MZ#*>W+H[K*>+A8^L!\#
PE!S@GF6H5D=^^Y8B0$74\:((;]W^S!3G?R[IJ%RML">HW3_:VTLBEB<@#I!%M/O9
P$$)U)T3U'MW8>,__982-9S@+?^^LK.IH.$8RL=&95[Z(U&7I6!X?V0%A[W@1$M"5
P.+X+OI7<*WWN6UN8#>;9L5]<AW&%/ 4P!*'LQ^/LP_M:F>_N?T2LCK';"P:]&/#Z
PR<SF(:T.\;3SD7DV,69P EO(-)<>E9D]#KAXE\R,18;(&@;X6N1@P5!5[$_I$O*V
P* !$C?" V* BL/0KPKN]*H/'0.'!/*54ZZ79F7$CL!1Q$D4M$4TOJS>6>@6X GO^
PJ]+@?,)4MWGVR&1@L:Z]L(MP[3*[L;RT>H6W.#)9?9N1XEH0VT,AQ['].5]TR2'U
P0*/V:O8\/Z#;!PUE45?:YR,Q\;T#^Z14/4"/U"/Z/=OE_O"P N+6V?&PPQ_KM=JF
PL/0>0!G,*HP<C415WE5*D%W_.3/*A!3^DJV</2>PM[KRC$<6X%G#K-\2Q!.ZU1DA
P&F5?+"R;>6 D83C\8PYU.VV9C88HTE-X!XZS-U:HSC\VMO/SL"9Q!?]3]&PJ"->@
PF8/ 41&2[[XSA80:#MWSG\&CMY-#MCEB=J.#$F1L>B.<$WGX%B=9AC,0\ONU-<7L
P^P^L+T!)%76AX^-KO1 1Q"+*ZPB#;R(LTA(2HQ%M@'S8,(45/6>J$0O!#S7-9Y?P
P?:)6546PW36N!G4.N5Q^WA4H4G57B //(;>*%4?OPLS7;E8A;Q"+=K],=JII8;S*
P:)QG&*3H^[&#8N2[J#QD-=XN%B?<,*@%;W 398SNU)&'CD<[$"^4 4@32U@M>.;Y
P$8EQR))RBATFSB9/3>ICA0;><@,4ZDFV_C> 627/-[MWWX\2;BAUO]0W%;,U1@0H
P_+_4,D) X:^+[E<@7-Z/P!*X<0^;X@BR\T GA;O_,";^] L-S";)M!(B\$NAGMDZ
P)>2IOW]HL 6,<GVO!O-G_)LR_RK>-EP-UO+CHC_7A-,=?R=J5&<U2)R8*(2U_ X8
P(U(MCF^U%-!;,L_0&4>,"!!XE.71O[DV7+^ZW6+%QV2BFWRYE2UEA1! ;BK%G"/Y
PF.1%7Z;)8'0G[TN[MG=+8I?1@B2IU9PPHL6GUB7ZDI$IQBC:WED:%6E5F8<%6F+4
P&S(N8P7V;(ZA7PF7Y#[!C"0(@I+0@@NZB^Y#WE=GY$8U#E<&_6'(=WO@E35!%]D]
P09\(!X9&&68O-AWPD_2-.=D2Q>:4E3NV:NS#YB B6?!JV3P;;+.<\C?3E]TSVRAW
P\\@F<W2/?>0G61\C18)KSJ6YYM)CK\!&VI K?B7[/_H5S/:>7?:W&NV^+S\-1PGY
PS:LWW=8P@3F.V2"C0TD08!1T2B9\:+<&R<4=?2D^I@M]U5<I W(($FV(<J5#@4E?
P[;MT#ABP0A:7W9R)L>2AY\J*A.U.^HIV7W_SG0/-$>(V0.O*9 ).H@7@/FNBWNCW
PU.;3],]O@.\YBTKLT*>2*(5=VW_8OWK(39M' $UW2\2&_?COD(N'YQ%_)-R>$JAF
P^#]]U9#6UR)VW.M1]Y$]*MV;LMY-U'X(K5$4\%ACWO%-Z2\T_BB&5\M]<Y1.V%0\
PUB% @\CO,'%9X$OO#5RGRBVX*7["O46\/#7I)0  "-"ID K&<L9_4E68BC4U2S5=
P9N= ,$]TJ8(V\/1:-K]E5>G8\D&1_)WQS&JQ1HV,O/YTT/;;$@,BO V;:?[ZR^0_
P&E3ED+T/'ZMF_7/WBF^7J<E;&)61B.+DVAAPS1HLT1Z2#"#[!:EA\E4L]O/&%UGC
P&HP>\I9MN6:,R\OPD;PPNMV[0'J;(@GCRT2ZGF0OC$"'OK'J/V1<2LDH+_<QU)AW
P9%#TLR :*PG3-GI<(YD!&6#2J/$W@.9?;3_OP\">_8G5*4.^J)E92G+ &!F>L^S?
PVKRT6>K0G,7#_Q2/&OU^BWS/3<+<)!E0 WG0SB:9CWBBLS_F22OI" >%M^@[NVL8
P@Y=R+WD!2-2EJRI.JOS=G<CIM2$&!1H:FGM:).W5_9S#6^_QBW-YUDHZ.+!OG#IK
P<*!ZCPQQI%;/C+]G>+AUUQANC#BF0PG2]('Z.L30@.2LI\@\Z>"[TTY^J0KAJ'3Z
P,[$.C]MD.YL1K,ZP_WGMZYB(6::;=51$C%)YT,9%>3]R:IR9-FJYKGH% )AK@U&-
P^1_UN.7ZJ8C+XJ 7E4\, #36,>N]/5BS5H5W7ACVJM 8-*YZS2".M@B<?0F"2AY:
P_X#!LM%^AGLS4TAY,L@U6?1G9+I6^KCGC/@'K6NM39KP[F_@6.]*KAYC9Z;9$?J@
PJ*)!K'V0GA_0P<YHR_ZKD0%!O,&I#?I&=B48>8_FUI.#> GN<)?Q@;18<WRB[MLH
P=]5I%5^F\'H$7[/\W.+GK @9(<Q(%4#X(YMO[.NZ79Q<HL TE1>;##.DF)2.Y L'
POGX3CN;$4-S&/X)%*GSW%_)L!$C1HP2W>CB?LEWVE_K%1GT764EI7U3=^.<.8Z6O
PMGB+=D(*^NI_N(A$TFJS-#:4QXNUQY_&*0N(#]G<^8@T]/<6#*>AE<I1X\=)-BQ/
PO%F6R)84ZR5^HOG-CA%S2(CNV,$BP556Z+KV<I8 W416\OGJ&(2/'9:*),, PW(0
P6]@5CW^!9[KA.F7N-ER;CZN!TC%WCH#8>IO.QX2L[#Y]LHB6H5!? D TMEG?&C=B
P]KZ)5[N'UDY:_K+OZ"6B25.HWW@:(0U^6LEW?E/(SLNB1O9UC6ZTD@34A7=[= LI
P$3;+H^F#5[!#C'28,)ZF-JT='HS7IA"JGW[W ECM9+O^]8Z)"L#Q$];I)RGFP>H1
P+(IULML@0T9+@7*0<."6OL1N-/ +8>3JJKSD;)C,L,(DU3=]$5Z(9\5[==T<WA!,
P4 H]@+LJ*9UCTD,#G1=9HL-6P!B\AUT)7YW^<*TEV8DU#M!I/>&TSQ9[AA1<D3E5
P3M, _M'FOG!G>8+N@GL''GO,Q9#V+)8,F4F#3?,9B4&90Y0T*<",P7<'JD,_4](5
PF@!MC[UU346ZV:99PO,5L3<OBQS#;!:H4U*8E@"YH@I\Q@>O,E=0JJLS14L0,Z'H
PC\$&@><YUD/+(6"R/^^.BK!C)0;4S(B%/<TUV.J62[+B^CJ>=RD!J8HZM'VO_*#[
P&!RHK% %TH<#!QX'5W#K7Y4@FM-*N$!.]P/ZV?U"7H&+847DKM#[TQS3B-+TVP:(
P%K.J!#E%VLVTBL[.\9!3P.Q(KLX-: ?3^\^#O9YY G<7E=!B <<FU^!M!50_($S7
P@[0,F0H['.&)&^^?"#R+4\C:!F"SK#AX=>X;$^ Z#";=0^]%- /GQK#7[8X AZT 
P;=XR'"+MF@D73L7MGNVFN($R6HFK?1'(./TVIVZZ)!F9MU@T5,RHE3/P/C$EE N%
P\>%DS_M0#LBV''!Y"A&/!#7[ES\AQMJ&0ZAM(BY=R-@I;'B ?8ATP[)83MAY?V:<
P#BTX!L /J_W_4HA.U-\5_F,8B_&CXZQS'#M5%<->?[DU]V>/543LMW;M7-S5X.V%
PT7>VNR=_H\B-&*WFC:-FEJCV ?6%4#&A=$<975;I1KQS8S^*XYB)OM<N#U,OE/%4
PW7K-$SNX,L>_TU#PT,F*%K)F.9;.E=_MR!A4VY$IP<L]LUI[FI3F.H5-%LH:?>MN
P#PU"]2"Y-"6)61(3[4=F@7D;MZ8.=^,SM*? F@G(8OA8<QX/^6$-IX@ ,'^BYEPW
P</621]EV6@-_?=UGQ]753]:R&X,&X<_A)M)/70B/(?$5D>@O00TJJ5?&*>:W'0J9
P1#_^NQ48HSR3^_+X+Y"?Y;TH[DI#:XBJ>51T=J4Z#02%J^D*.:^!8T%O$-^$'H(2
PGWC$C"RH9J1&=Q"7E.4@AVZ.7P:-D[V)5Q6Y'7\9I\\@@9M/:/76Q.CVH=!:&*,1
PX=,:KVGZW"4+SR38C%8]R6C>:IPULIU7&]_)CB\*'2YL!Q.^S)\,Q%6YKA!/:$].
PI L)"R**(%X4WV0&.E&CT>N% S*%\Q0R(3$V;UZ;_B'&OX'DS2ISZJJJ+*Q-+Q9N
PC:#&I,YG='TAZL4A%A!V93'Z-HIB6RS>X_]YX?\Q LH9^O:Z?*LW)(LYED'>%W:\
PGW@R"5U8S305&?OP$P$%D]Q]R#_I1#AF!_U[+AD^FA%/J J,14(&87Q\5IQ?X'H<
P<RX!DZYR>YGL$35U#%H #7'18.S84?XZF/LKZM%YVP+U5=G\3?:XT.7'9]^>YU-N
PU]]NRGH@NT$PKA[>&'*1K(P.3/M1DP/[!>4D+1:<WTXU\69;^V+;:=<6N!/=<1F\
PDY]CQW(H;LZQG NJ):F^AS[M&MTX%2,TK[,/.J:,CQ1H?EF$YR"E'W^^4CJ]V[YZ
P4AX6RW&G20H.$NVLDELT!R-K3#CSZ)Z8@]H^1V,#T<$"_YL@ !.4E]CQXO@Y;XS1
P= _SYN+?0)3#O-#JO5G[&=+>]JNU):7S4!;IR^*T/09 "O".@0YJG< $>NVJ[B#]
PZK0_DD%#V*[U?!F$#ED./T_V7R584%H7"_P0.  ];VB=;N\Z%5NW:;W)I/ -K,ZT
P# HPJSP%LPZBGEV?QM"D.8+[8,7NERHFJQUJ?:9LF0!XW#T&"4&._&7-D=X:UK*6
P^D6G4=GLZQ2Q.-[:!T]Q:'8]-8A<(0K(?]U(,"O S\?$5IF:\_7][NI/:E=4"R98
P=*D,J%K+3DX7+7 :->#PT8^X5T@,S\7,B=A=N <KE:U1BLB0=&@K/.'!A!\\";OS
P>6DDY$$%N RCEM5ZD?C+OM/BNAG84"KR;RSP=U[AUCQ'2M7<Q=PZGN(&C9E-A,(P
P_*2+S!NQ?0\"DD&X4N-2RK;2_90Q &@N5;X:PN-V&A3%I:9_QV'6?F&O:^G34-[1
PI)2B8\2#,;A)TU/U1T.36CM5_L<)SMV]8TB_FKDN%_A0)5:]PU=D)UGP7)]@)KLH
PM<':*GH 6&1N*6@_AMO//+ $O_OO!?]R]GUBWDA/(MTX! (WVS>P?BCEGD.1MQAI
PH,)Q%@OP'UI<25NN<"N\)91X"W[V05AN07F#;Y&31./>EL2YL0U5,,'KXP+^5#1[
PF-7,SHU#JE'!*Z-"1EK-93AZB'V57!3UHW^$(5\6.Z^)HQK.>?VJZVYS.Y$;+JB0
PV>96$A6*NS\N^S%0N-!6!K 2Y<Z)LAP78;MUB^$?Y99E@YY6PWG<N,JHJ="$K;/!
P$KDRD84B(Z9]Z*VI/B5OKZDJ$\I'PP6,S+7=#5RA?H_6[E5@H34/QO9FH>18 XC%
P!_[H,@QS'/0?ANE3  L#\GMAY=(SGRW%Q^2YC0K$LX_M=N;U'ZV.'2K[F"<_%'TW
PX#Z0HG@-J I.6P#'?;Q)?:$<NP[7_IR\81H(B^:,CXW)R&)T6,+#[:I(@@)D0?/D
P'L7.4+*3_KQ&N?9M22$MM2DAW0]!:CC6UX!Q)8!\BOUZ[D+I<MR'/RRV:E?#J]'"
PWJ'5HOK'?C3>]6Y6W4>-V!1S!Q\D-K%*_DL<6>0LFAR4B:#0U8YO*8CD' EYI3D9
P 3[CB\@%]0#B299L?HAC%98#@VX.V*@Y6,(=^]:<_9X@H14<^7XX"'RS2, 18N"L
PC+3$M@+'FUQ&F8NE;ES<6Y1@-["0GZ^DIT)^JS7BYEUD-\K_"U$(F*4 686#6\GY
PQ&%CS!XA?];&B*I2$QB.\@P8>^JSPWQ+-$G30_SP)!(#'\>BI.?R,F+(I4>23?AV
PWKV:\VF4>@F\!++H(-!E%D\[H[L#8O_=_O[C]!7P&>\6S6"36,Z>)VKCJRP2=BK4
PFAKA6Q9TSBZ"6U!#W*F/XE^IW^4KUF6;@*!<WDEM@O![!X87QBE+*S>QBG(T-YE@
PGS6/HA<:\"UAKN2I+G.]"J0-E2;8L[H9Q*0M*!?JYRYZ(H3W.FH>4!S)S^+B $8#
PEJSC_\;-7K?-FH5)*Q0WG\PP$ZJX1HR*#764GYCC!_0AG=Q,)/*:^73ZE[AVT>J#
P\@<^8=0]E?WFKW7KK4N6$9Z7+XJ&3<#I(.&+M>MG'&L44R-TDPETC<PI(>HQ*Y_+
P'Z?N &IUEG>6OB"5ZJ@>=S=^*ZC(,IYW'I<>OI8@E5QBX.4A/_-;_Z'5Y_/$*MF6
P)WG19J/4I\G?Y,PNT [0I>#Z55^$-)JXX9,["V>EL?WK QNK+.P'RX>DZ]>7QT(S
POV(?W:6%]/?"7!KX6\B*C'+1GAH"UH2^ R7NCZ)[KNTZ*]-@Z3DMH(L2B-2[-2%?
P!'R4'!=(3&HJ64;_/]0ALC[J_LUCD)MBX =O<3?=[^,IIA.]P8"ES'751@7>MN7/
PLQ\T^J,Z2+7+LDE:C08SY#,_;6(66]@'FHA;)"G</U&'5_JIWUM\ GA'C53(A$\P
P"J'Z$#28^6/Z]_KRSI#J#2#W0#NS0P72;=_)Q&.WL$<6<T?0VK?-Y?_^OXV@L==S
P._:BQ[-2_0=//[QBZ0"SCX^6WO=;[#]=U1[QJ"07<W7QED'GSJ7[%9M"KWSJM^/C
P;O3GD7]/T'P\QBQZH,G%>8G@] /J!L6NEMGT5(76,S<9H(F>SG^SUNPK/V+02<3K
PZ=GNM1E(*_8A1?*.:?3VU[)2/=WBWT_88=E'1]C@96R@4P7[=T4]8F%^(]H3?Z92
P!AJ(ZGXI20]G!W"'RQQ%\ZR9L,^[E E?-%V"Q/GSR'Y"%%J]34Q@S)9KQE9&3A 4
P*003&Q[0K)X-8DX,IOZ'_!;W7#[E6PD=%BK50U LDP%AT@/K6H6=84. 3T#9YWA-
P1#%"#C+>5)V16!<*9" 0?(]&@KL!F:['4FL3-$-K=V'KP&=]X;'?6VY=3,_;/# :
P>\YTMZ977!\XF*6;%U$2*I$E#19X-]Q(>I!>H4/L3( 1+U1MU9UTEXI$FQ];*K'B
P,9V'MS'R[.%.<]Z S=E-(;5K5$2-!=H,3J@P2*?.<8:O'A>TJG];S5WM/JX1KFQ[
P2?N:R4EXR>%T:-P2>=+/WD&P=#6KN:@.3V6K-D<9H=EP#U>A8-N#H9I*OO78*+JP
P@5[Q&U@&SK%:%1WWL</@/DF4,!K+I1P5@-HEY8;Q?XZ4?HM_-%%(B(Y==4<)QB N
P$:]Y'P?9#BCB=_S&QWK'NE$J:=A+-W#P()!1,1EY=R97DG0C\^OLDC<78"'UJ) 8
PL$-X3&%\.$6;>IO +2E65%V%%.&M7/>F^1U^?Z8.0\-J/NE/,4U$+Y+RV2U:5IJN
PT'&\J<W-*D$18(_"<S:#$</)MOI/0:->F03V3)[N 8,I+O7GZC0 _M=MH"B,9O>H
P-]GT,[$75.WVTB8GJY_@!'8+&/"3=)#!T1;%$Y$*!^U(OWF@JN@2%ON/7S?X;W$1
PIC7.N:,C)61Z_'[R>5DML?;S9A1->MT9IE02(J):2=-VZE<C!GT:IYRLC/?9&!NG
P)ML+QW-J1=00( -N.0O'"$D7RWU 8-7*:J=1E64F8'-(^H%V@F<?AP6N-,[^58AB
PQT7:RXUDB*214.3V N2@LR-1U]!/17?E0)*&]'*P+70Y8BS9E/T$VT\H!&23TX4\
PT@KYO+1];B@*1JHVFZ4/=AAYH*Y2%7)M'*T[I-U$8!/"P1OM]>4[[^U[*"?\+VJA
P0M5;\48&^<B)F]&G J>#AZ/8K3C1JJT)FY>6#%Z_7'Z5H]'FNM\VJQMV2?(Y@>DR
P/#&-?=GI\J+PC:IHN:IBR'77#3^9H)*4F3SVJZS&D/D%^[DJQ%:E:(3B<)<(J%$;
PPK+;UNB'>]K""CP*R9I73Q*$B(BC&Q0)UEC1D>/O[\0BK05<0/^T1S:])2==Y2\<
PX+U6&TFO#,-X2[R)A;-C_3$E=E,/<"BT&@N@QMYKQ^_6RK+BOP)#45(-VVR->Y F
PV,V7[_2SNW6V;BF:8M%J7F@<LQ;>^>W9\@\%/$JD,#IKU;<ZKWN5X/6GSS,B3:$S
P3D(C[!)Y Z]&&CR'O\@+ECUH=4*'C$/$E*PV_6XW-R>]+:X^HQRVV5E%Q+-:(EO 
P5Z!M8%6*MQP;>D1!*?+6"*>X@>?EO<O&"BWC%\=@)7_BE1UHXMI!!+XD/X-K53E4
PRYZ')<K&?+\%CR#,#]5.<^M!Q-+)Y?O\AHN>ISMEN'&I23A/01/F85Y7S1_40;)(
P=>BF&;TJ9;%;.]R7R^Y %FZ7.@5]!>'AAPJ$E=QW7=F/Y5F])6-GM8.82 P=LX?D
PIM\Z5KOKIA\W"\!3P+@!V=%?;_))>:8F>$Q "1+D:?*B0K0]>#>[JZ[D1'A-P_%/
P,%0^EO0?*_BSQS\I:"L?"?#Z^436[97I XBH[=RC%]*W'+L)'!W]A#OHXB1<]ZHM
P>;)7N6YDIH*5C5ZTY6XGLRMFDB<\=Q>/<)=OS%1=)REN:YAD@F:<L.@F,65BX,3(
P1 %Q/ ?SW^3D2I@CL9R>B51<LNNETYT?%B*V04N_Z%%)--0T=2 NDEMM 7I <X>6
PER]$;P"C [GH+?0(%E0<3#?F""67#0'6>X,P#P#>GCRXT*1KY2<TYW@IS0P_202$
P)O#0BV[71L=QMM!!KUV&7\883WXPB\#O,"%O;GABYM&\JN?1"Z625G@EUK? PB)V
P;6!?^+0;K*38:Q.2;'HK80+IULJ8[POE0VXY6=L>6C$_L8\59_D<=DT'QF <C^9>
PT9E:552V6;.BQ_DOF@FE5/W8J$%0W)3#%U0 1\[9KHO#_O:@-U(22PT:4M<0@\1Y
P=*9L"\0U<[1^N4J$_5+',8:JXI^+?8=9S$B9"BD>%"VK%)""?:UZ/G!Z9".']V")
PQI (\YP''&ACBVT0.M\5YM54Y!LBUV$;9H6X8?9#L[D*9-&OJ.*%YA7T2M^R+_M>
P4[FC9[IN#QX6D*/MU23V]4LU%5#M'5-*M?+Q.TF6T'/X*_[9^ 7SJV_TG@=5,669
P&"XSR=E"7O*"_7_%"VFJ6-UN'Z,%P,SS[_T<G.)7']*8N48Q/8-H_3J]>'W8,N3A
PW[888>NO!\9IF-ZM2*O-[V#FO2$=CC^J"05*W5M"E<E:0&DEQ+.Z$]%_L3&YN^H8
P:#--8%Y6[>?BJNW0*"/]N1"XGU!ELA=LEHF/V<0@R&VZ+C(<HU(0+!"H*@^_@A0=
P6OICJH^=;]CO6H\D%C@#QT27(HA^)TC>)$Y;,BS\;=NA="-):M\+<U;@)DJ-,1V3
P,=[O?U_SP\,_\Y,[+6.[5%(;5CI\+2M FDZ0=TE/E;C 8V)-9F7%N(_ZE-5/?D]F
P)?QH.AE!U>6.5M9=A/N I@J^B' &QQZ4=:7.3)BV'FC-S+B,Q-;;/O=:@3IB_Q2K
P !L4Q+3(,;[015_QW3?=*<J]QCB3#; 638CW@Z>7FRXJD9K;W*@F7T=,=+NH-+ J
P6WT-YR*#6Z.:#]L=Q2;I")TA4&O0<D%7!FV(U9 OH*-?ZS\(49XZVN;\[_\7 CT1
PF>/++ZW[L&+/BL5IE<%>SM@;]_B6LR:+8]T8&JBRQG/"'! !W:D=[MY]'Q+TM7(T
P0E\:O!-WCH:$E41EAO^)S*E<A%I[20H,% Z #M-^>@4V[&_X[^6?WD]S=G.%SON,
PLU4)9*F)F!#&UY.OJI--S1$G0^>6GM_;^DC!; ;%OP03M6BR-.*P6-7O@9O>D7T_
P-!GL*@$=<N3)IO>3H5"\91WO^)=EDA/1$;XT>0E4X!ZG#+XDUX!)D@GN4E!([HX6
P*SEC5Z&VCV;9"94%ZWD#L)#[^!-NZB:>=!9?GO:J"$@&@Z-UK(XNI_@>DFQN>++%
P1^# @!&K'X^&1GNZ(F]QR/%4:T^QW3SJ,K0AMC)UF!;+UDC#R$S>%>WC3>['^Z(R
P7[:8>1-(Z"JZU$V39M=;#[LAW_"U&KUS?V#T=&W]2E1#H\\S-5'>W0KHRB)1[GY5
P78BCB)2YDQMLT&>KPWL1XN546;+<1W%5V(6]6F\5E*HW&2G21;[_?Y@$48J.]$RW
PR-+GINLP%=^2=ZP4\T+'NTA[7#2A%+Y/1E++//9H3KQ(.2XBI&]WS#O+E;@Z WN;
PF3%V+?+^E"AW5,6*"BHZK?%+!:=CZ)<V^?FOY5.TF+&H]ESXEYY:ONR[1]Z0L18>
PA=JDA:F$_?E(V*UJ4DJ&H *I8(AU>*E=)Y"\JV(2S]HN1M/ZZC2G\Y)6RN>;?<M5
P^@T5A*,O>:>+OE5[WDM%A(",7A-NH?'-M3,+D6G$\NO;6=5#1P5FN[TGQ9ZC(?FB
P!-VY7!X;3F?9%[:<6<LV;563N8V,Z)? OC6)EN: ;HB-\/2U7L&<; -0,@@#_)<,
PF M/"C.TZ$*X>=C^45@PK-KY YI%:;UU^9<*$C!Y%X^CI>@E)B_281*Y7E^%GTF?
PV_LP]-KC +ZSL+YH;0^(<LL@EB#L_($T<)?RM$CK^%1.+>G]1FY>'-/<&/"UHFM0
P%Z(K9!M//IEDO=9ZSQ3VI?P,C.8WCDF%8Q-> ;7ZK;8#V#/> ;IM8H.5C8;ET!8S
PH%9X][#)R^G&<07IXDI->DQ,=?9B3E<$=/"36]%F;/5R:Z2VLKI5X785)<IT)LZV
P\P /T6<)F/[N,"):!"5Q(YSG\5Q^/(U9.CO&DJ9W<:_UB73QQHEG@CXJI]E_"\?*
PX!_[($N#KOV)0J3&I^K_=XCR1/9D;6(6%6^6:[9%T:-.2>^^P\6HZTPP([X0P&I,
P)[F$$,5G8CR>]B=D1D'JW]0O=T^TL?MFA1&![X45 N&2DU)8(F;J;>$W8T^64X6[
PK1S?">*OCA <D02\+1V &&F"^L&7'48$O*T]KMP31"!4I[;L9]3'-DI:QJ[X<2K0
POD9@<,V2,W7@VW>YJ6MM_^]Q(.,I50GEXIHP1:/4*+00JJI$Y.N3V6(?*<7M2YN*
PP#\J^(<KSHL/P.9XCX%C?$LA+Z1\$5 Y&(B[YFPXT1FK#F1RN-.D#?29:MY\+*6<
PF^I=_I'J%*<G2)D,\<5ABU3]G$"]GE*5=^$'X$%+%R>\&8!S8Z8K?WXW7_M8FF^C
P_A?X'V_X5*T6=[@]"$33?@42)UXOLO@YATI[EO4$;W$"0)E)<\Y0%!*^NP,/.X4>
P"V*[K60CRK$UU7]@'VQ/>@I4S:!@R0L1(%&/!MK.Q8G\4"<>P.Y:&PY!;-"_V#94
PT=>AAT/__#MGHL"^1ZTV]32?_PP:6%O2KC2,-X7ZW[MU /Z!0,".2+YY[;1--Q:]
PGI=;7)=2X/958YBKZ9UU9)8K_E)P,F.NBP?P>9XQM#=I,3?9A#@'DJGU/"I[#JH>
P2YG./1H\M8C9N S.52X4+H;<0F5/!:#CZA]O*J0RX+SG'E4GW<P7_>R:G#[* T@4
P"V)SR"I@HH:[VIPB8=%+GAR&T&PV ;\8>C"1#;0CKI6'H)W!WD<IL?T[;OP^W_F1
P[-)Q-/>^;R:H)\^_/:6.T4S6JF&_O:M]GXCY5O_38]O+BKPO=9R<SA;*68:;SS0+
PE:QHD+OT8G4HVX5./3_Z>3[4!D/ 7H5?J-F4VR%Q*[2]8D10\7!8J%KYC@F'_>U+
PE,;MTV?@8>6U0HP4D%]O#+JX>[,8I+ ^,6S\-TC=C",.YLN_*7XBU(#]C /8JOP 
P41]W#_!=E%H[YC*^_53%RV<L^[.Y6#0>R!SNKD?[+ZO4[NU7& ?C-.P8.;S?*[RB
P Q#S*ZV"YMJE!1BN4!1H0A06>VW! OSR(+%^<-6O%Y3X+/?;;H/N)1#ZYVJ[C'5D
P!^DL5+#7IASOE%X%K6R8ZR(%&5JH DV$2EE&2_#9ZWPTH:L33,:NP)3[XG6T#8*6
PL6AQZ3XART'SJEW.KC]P$RWG5@P$R#W4X[\$"C8-L&62JRBN]I+<0CDOP)7^<&/2
P11M\OMR D,!56]A40&%V[9R,*&>76[>@47V_L; 80".!3?D6GB0Y^K#-.$C[XH8J
P[+!7>HU_FY;>U^('<NT1N&T]Q@1%![]3R,0%>H/1+JH@9O\J6,4,65.R*BV^X6V0
PZRF=_-FBHS13(U6E[OYP,/VZ02/YUC2OJ37:R2-T8U\?-?%VJ5<049:*$THA.KFH
P.R1^)H8<+FSCI<##$.TU_P&%@H6T?LV  L!H'OB!Y2"*'46BB(36W07Z9,1#9L_;
P#4/' M(O]N4J\MBD)DY([<@"G6_XD/A:>))\>*1R,G9-7>A,BIO</&<:V U8-J.C
PY]RI*MTDY9 )]:A](!D]->":);\41A/C4"B3NWW_#X*(;>>F#S<E+=.&EE>1/UV]
P>C>/O)Y3M656QIS8.C$TG;:P[5)L<^*+4TBTM PHE_7\=9>L.W#OM4,# /8CI6^G
P''HM,9"^0&55/MG]U_+Z?:"_?6$G9PQ4O0H.[N_"XT7YBPH\*IGZ4%)! KGT=95!
P-2LPJ)'#\7#?REO(C%7\T'@+/0%YV(>Z!Q(<9?$4V"/,DA67QJ@P/%"PL_^U$(#^
P "4P=3@&)!D7^:O!MY+=A0&UPJYP3?Y:V3Z^T+PDVB4.O,83[UH%Y+HF^&T;2X 9
P"0D@@>(UZFTPS,I8E[+3)#V,N-N0<HF3R Q=<Z;$?9Y4P[JT1SG5;W8O!1]YS[_X
P2FQ*%7AZ-\TLL]*U\RL6@M"LWC(0=.!EM-MS@F))SZ\$KE:^F:E?B8;;3@'R.R(^
PY^7YL"E\'B]P#]7R3(, U7ADS"WOF/P.\9HH<>@_M]"<T:*3@&?I]N+UZN[4@OP)
P89YWKL5#C?=.TY3/>K7YH=3'<;.3Y=W.8&ZD]V?D[5.)FE1?"N^X[\>4P9*;("HA
P,HA:XFU1^*F*3JJ$Y$KGJU,/^WR9?^.\;[K40'0WK9M]YO-R#E^AC*0U)6O?%4(M
P8V#Y5/,=;C8I81/[V+R52:<^C4@:?D&%/'.XY058%R<;5VG&-NI>OBCMJ/-ED0U%
PJ-6 %>Z";' (G?(#"FEUL$KF?)EC!+;A<4=%5=CTP/<BY)4DDY&NGX'Y&GOV1_#3
P+99BVL96HUW2?%S97-LX= SO.'G5+N(>MBX%%DW8C24CHJ@'ZK]IY !]-YQP^"T#
P1^9*POXV+D!/S25/MJG7>@L_<STZ?]<D^GE5]N]5F$\X_A!3@7_LKZ-Y^PM"F4# 
PDTKJ!?,V -/?K(1=JAW7/C,YNN\-SUPFP99&'A;'E5FA,0D$9:0_ND^U7*W=2GIS
PLS)[7@E363KSF>.Y;C7_]V?TX*R:O4<B/4N!580$N-/;-IR8LS;7!4)LZ]+F[JM<
PN&YB:H7$*.+9$GA D)O0?NGCR2R9.-4.J_^TA@2XL128V>MCA+\T:+[RC<^8?85S
P1BR6]"-3\@13L&1AIJQ//2VS9QC)9O=UY&D!"8N[)-)<K-03\:=8, &;W8D';,2B
PQ;UTT@-J:!6W.*D)J"\86,-<&G,WOI&;(^%,[[LN/!^;<9)A'[*'<4BG'CC@"!*B
P-61LFI2N=U=9I3X1D8EW"V/S;7_ ) 2( QP-O]D;IU@!FC3ETYEG0Z]$.D7HL'.V
PQ* D?4S$,&1L+UM_>9IJ2'H5AD':T@P^3,+=,>YJM/$&NQJ?;"]:-6,PKM45%8)H
P6:%K/ 1L3_ =\< AGF!PI*:&WJ;IY=4<VE<94:P+IIH2KW[D%(EA2 !FJ6)&E WL
P@?.1Z+Z#S;SHGSMV*D7IBV_5B0'1N)RYM]G].D73_P:Q&PU/W/L4.]Y3YZP$L;@0
P,"8=BD3E#J1[">0T&[9>W%3/&^0%.Z+A"2B%$(#,SSUGU\<CUN,;+Y)%@+50G:1C
PN)(,-NFXJG?N>K(!^(A)5Q1Z8#)M CWMJ*T*E-V<S'G[:]V5[O[PZ4RZQ@'+41./
PUHZ<FZ)5C@LZ7/$#_9+,YEJ:G12<4N7T\$?#!E(I0*RW"T(G[L&#4_V'_)9&_HG.
P?._@KGQ[!AQUMQ?A&*%](+'15FMO@CE1^E>'/&X=4L.RVMX(=) B<9_,4]=[0-JP
P;52DLYAU'_LYP48YX=/_F-98I%*GJ-V%D\@V_DCM..LRSLY+M.XX\O.5H56AU3Q4
P:K*"<FW,#E: 4W1E!_<]PVF'<6G8ZA1W'(US/]4W582=/"H/M+HO<>% S$]BE]'%
PE(%6[Q0QTR5^R51XSD)&4!&-O*5#>,GR@C")>9,$W61M01YXFOJ@PZ9MX42'_K[A
PV0!JXQ>G+3(=AB@<R+ ":#S;<KFU5E*:%,U>A.)9NJ9]MIM2S))]VB'OH%V,E[L3
PHH7E1RB+ET\OS0RR,98W<Y#";A++>L;6PO)J=_+D!>@@TJODKKM5E.M(^*MNHJ[F
P,^N!_=QWC%IM&GFM]RY176$XJU:#0' 0P2:PP!<X/N:(Z ;*:<(4P<2_1"^.I TO
PA@2V!V.N]4=1\N*GKK<_OYH,?GK$2;?6/\$W252,+0XW??Y]UU,'KPY/O(?_/=1U
PM_0?.YE_;.)$3#G"I/[;GTR1ZS:.<>[V:Q\R@&O>D*(EO6\ IH@\_O([WEGZ' +N
P<+D-5?^&)_I&#!6\EJY4\'%PDBZ)H0UHZ48CJM'S4ZLME6O)H5HO6W.5>VN]CJ>A
PK"4*)9"XFI?,W LU:,S2Q0<+ZA< 8D@=8597YZ3Z[;X\QSL"L\\$21@__&*HJM@#
P%,.'3O%H@AQE(--@\D!;%:S.\^@^M/UXE'I?QL>004_[SB5%._%%IN$_S22ZJ/& 
P%\6HS87VKF5FOIU%/U?7A.UT?$^#3WH0[\"[B7I6\5-83"L[W'K^#VPJ3U1?&S/J
P:(6-#OK3$K,-D\M!'L5=9DP('7]HS%@!W9'2R&Z?=;(7\)/%)"HIV&V$$H 24^M)
P/1MJ/]W,!?;@M#1_=DQJ%X-H6=BN!&MM"Q!9=Q6;2,*":8F+P+Q(>IU@AO 0=2/:
P](N=-H9!YJK5ZML]S-\0TQ0F!.@Q0I <0:4E;ZI;:5*N%FEFG*:AY[:'3_@+5?'-
P'G*J.EL'O<T9VQOFN/A.61B[IDN6Z6V9&N)#0BS:'3DEF0?HCSN4.C71C41Z&E*N
PX:BQNQ=$3C9"/K&Y-H?)!M43?#QLALSRT;>2.1.[?'JF(<F)9RYS26@D(XC'VENJ
PF\]^WH@2&(>>,F\;SQ=)_D=:4E?H?L+,.5,:PAA%,7ZM'(P-!R-K2D20DI"O5(M[
PA!/O]K<.&_V=U?9G=FT\EK!Q3E9):.\I8_(%7Z<:Y5<8\E<K,39L&]@8W=5<EDI*
P=>4\<N-7F9>%SD32!N"HP$?&3O:.N@E=S^BVBDZL?"@@ 4,H;/-KP8?_>VZ3NT<N
P8_1<()J1A%]D?*'S] ;X2P\Q+&)]=RB4)%/_%TH:TGU6N3<WV!V.G7)I$GEC:.2"
PAU^DJF<50L%HT,3.X,JA\_YO9LVDRP@3@"YH^J9++SBIZ0^X/!K%3OMK*:MPN;$X
PI'RWYJRBN)[EH<=UO_82;#51=FP'#A\O<701M4L.,GUKD\16W"7ELZJ)5B>MC+P!
PQI$:U$Y?;XLW9<Z6DEANOQV_$!K,HH?D):_T$4O8/?.;G.&XN4,M @+#429.8NDC
PM N49N&S^@Y_/^2@F"UKI ^V2(GZO1+_+DED:9P%.H:&<0E)_RCG(M%.IROXM.8%
PZ3*^%0$,*4Q$TXW..B7VQ)*AZ]1VN=\1MQ]%<W2YG>!E<CL[FLC@%#@9YP>PX%PQ
P)T+%DE*;X *%@'-54M7XVI_H?D>(+,S>X^HCOORP,4_G''NI97ETRQL%-PQ1F_26
P9(*"X Y;R\"6\BI4UJ.HFEE\G>RR"2=TLUFZO)7KHM8?HPA04O4:D7&-M>01I,\7
PWW5<^+)#^>".*5$K(#4CN 1<>@NQ9-\QLA\BF<>27T;UR:*XT 9N5E(C][*C^>>+
P(AG^!SE,YT8R[?W.I9'6NS&&,1,$2M@_X<BSU_W@C#_I7 EA3!C,F9G&<AU]TZY8
PIZ\;;'/2Z=OR@[*^%SGL0]#&=*B5<;S\ECLW_U_$?RX.XT*JRVS&Y57$ '73@<?_
P65^O6.R&QZH &+-3VV?%E655ZWG&H$3+E=&/.G$^0('CUGQ2W)/HJM_NOO]9LNIX
P)2A!WJ,R<U@@^JY*/J*[I#(I@3=SJ7YC[]U":7@Y^PGFM@,#EH0QZC2NQ-&5\SHH
PDVI!<G//KXZ-@W58 514I2L+P;EVM,,#G"(.)MKU&Q#K^TP8.C>3($"-H)AVN-3%
P1UPM+]K<.-07GEDDC3T[V(-8\>AC18KYD(O?!"(@>' BF!QG75VC+6") ,41CRCN
P36BWR FHB4P1E#N*Q,<^8FP2=:3<L/Z8D.LHMF,ZCX(8J(OZU8 L@C<YCW7]!";D
PXYB#7G'0^:)<438+^H0\O6T4 LP94KLSS;-2]\A$SW![.6\Q$.XOJ@H1O@]*-V9E
P! I %^8#0VW5F'4W/5?V5/'!A!;:838J@':G+__8>P)8?J2^[$ZC9P/$G"^"Z_DX
PXX'6A@)CZA.\V!^+PDF1RC<)Z0%HDJ$N[S2+A-2BPIOD"L?]A9KNJ< '7(WCQWL8
P[4S'PH<AA.R(X/_SR*AE*VV73QSEF^9+ %3'Q4]H<UY=[/1F!HK_[&<="F35A#EN
P]B)>X/NC>%JS=AWZ58^M<9>@GTR,E1^$[C4,;?TRS"H^+2ZO+VRY@6YQ+A,L*_5#
P(5%SLRZ D/C=5=7/+(\EX2M$2AU_.-*2]HP*F)))(I;VKPH+5_:DZ&OH?Q4SGMUW
PM.R>*DU.NS=BV:S[[%2\3,%FYD_P@R:WK@MD;[X/CY.K(52)&O622G:"&C7*,!4C
PC?;4T7?!! RNG)Y9T5Y%*A@"J<%44.(>HYB!(MQS\*&(EI;"+]L J 5L')&MD1?!
P!L'LMS@#FN:?:KTO%5MJE):L7="!88%M-&0+G7G;D8]6F"]"<LH],F-FYODR*23Q
PP>&+R1B?!\&LH8$+?QATDP0G%$DB.&1201FY@L-&[%Z_]@L/-XL]9&>\)-:+%H0W
P_XQ]IZB4'MF0F%>\66&=.63M\>Q&S$1$EQ]>W]NG,KG]-Y1MZL5]QI\+&-Q2CPW>
P/-,=Z,E4D@NWW$4)PPFL=3N':74_+2FE+=\"U-3!,D/H'K4S';CXB3P[]O'E':#E
PGL$YNSX!SV6( ^$>8T,#,4T4",_^5@TX/V%0[)4?K]= ^/G;4^$8/\YP^^NR+-Q1
P?_J$_7*Q-JV-YJ\YR4V?3%@':K>OKCW=JAQYC-65AIYOXF^P:(145F[""T.LR$?X
P.;-9P"$TV-+B7*5#86*^_Y""F\JPAV]JTQ 6*M=PF1B#9@N;(YV=A)(Z,5AWR4&C
P5J&C9GB'TI-:TXDZ6HFPF< KFL_9".,*LB**-_)#4<&5%)F/]>?A:GZ$[O (81#O
P2[P0-S"K!W"%O!!?5B7MLO\]S8&M)4\93S%.,3V%O%Q V*D*9FPW$<GOU7SZZ?E1
PR$+N:P?PC\/&"0FSCJPQR1Z;,M9A1\6&_Q>CD_X)@8765RL!EU?NUV'&@[S;$!^A
PW30J&8=R<^DROUJ>WPW]^O,./.A(0.18/UF'106)1";_(FT7EZ3CTQ+,_\..$0,?
PG: '+2 B<M.=52_;PU_T"Y._);_Y =(+19GR-:+RIY*,J#MH%<2QV&,B(C\D\*K 
PTH2@7:(NXPFBJ]N Y,LH0J"YCW6P^*9$>9K%!-)$";_DJ6N+P ::KYYX=0@>E'8E
P%O&-8^TGZ[QK"^64C.4%T>3"S@;56O"PP%'KS6$4I%HC+'?9"(F9T0@_\-JSL-=5
P3.J=4OJSV["NOQ@'XPN61C*_JLYO+&F-E##YCY+ _TMU82Q!'5@4.W@M4V'<&3PM
PZ/KN40P--;@?=\(TO&UI#&?&T$&DJ-R K7K)]!^!8V(<JE_&;(/6A'<0.RG;>O:B
PHJ^J(9,5 & VZ64]3VFPIR5W0)Y-"(9Z(YGW^&9MDT(I$"5$O\/^,0X%TC9^>_YH
P.4;J[JXB35F]F?09OB*-KTGKBRJP[84DX4,\I:WIVN?T"FE'^4B*@4L*2+2T'E9 
P!BI\.(H#'U>" XYQSU\&@ML[:L!:K4BCXV!V_MB\*UC55@]CCH[]_!-HP3*/\1NM
PF<(S_B,UCI#:>7:1>?FA&T\7[IF:&B7H!:47\*/MV%5U[I-^[6FQ#P)&>?UQW>3J
PE6B\GX94AKIM\OZ*[:*D]AMF",8&47DO#V=/  8N1Y94X)L<3[]>BO/_5@<"V!7>
P*_<%MUMHIVF^(IRTVVI3'[ZD<RP ZQ]ICLJ>1PINEDR_7!7##S)QU]%6_.:S<HM?
PI0@-[P36DMH]0MEMI8YE-6-FG^S)LS@ATS_@ ;92\'E\%J4)&^.L:27'U3*"H?L^
P86>*1"HAQ%J!F$H$/A+\HB49%F6:_(I-2T GKR)>T%S0^V3!7O>G7S$$ XU>@X'Y
P($P.RD0<L0C8>.S?&==/73F'1:M'<@]&F]0(Q\$M(F3$[XO5%-BMX3<G<A,'==:"
PE^]LC=+FVK/P6<5\1)A=WT84B954()?^&40<NLR@-% <(04^5SJ:D,KN<E7L"0%\
P.71[L)_!K72PJ,WZ2$*0RM+D#30R3"\A=C;7<.AS&[$*0@C(CWWGC!"=SBKS#%S.
PO9Y;B--=I*]!.Q!,3LO2W2(V,U\ZSJ(_[T](NM0Z,5(<^160>.MT',@P>GQ2UTFV
P=I0B99/)F70#?D@N__GF/,X-+--AS5?IAYS#)2 :Q9=B52,O1QM[\\&17MU5(W)L
P<M\J^&VLJ5;:_'%$H,%*<!2SSO*2 M^26[E(MGM3K>\_^D\ G%)WJ+%6B'0*3@ <
P_'$TW2DU=D+?*H4@H/?(9?6X1R\C(M0,9\#.0/2_ -&9"#N1J!G+>GBU$ASG]& S
PKUT?+C^K][P4B#AKKY W$5Y'6NF@/5]4Y5+55$9N>;IVPW64;V4>MPTA]= $4&R-
PXP91D028HO[RH48GU)"7\]<&ZA3I/P V_G*/,$"PE:K1X=)></D2OW&-WR/GVJJI
PL.5/0LI.0E&X'IE!N:7NWT_@C< =XB)#V>0V[UX/;M&IQ4 :QRU*-EY3;T"3^@YU
PN$6&W^_/!W.$U\K(% XN$+"&&V3<)!^6D#:>!7DI-V(H%TN%H>C-?;GD\"D," /A
P&B%?/;>N#S&_ZY)3X6'\L,D23PJ0C".U[7GIPA1S'G7=YN4<_K2FN1\$##57 ,1@
P:B5F.?96L+X@A9H&"S)D2=)*)_@N;^NK!T$/)"2GK&(O=E!959ZI.Z1*&ZY1\GML
PQWS+/O4Q7XHU,[,)@!>VC1K<V!A-X?O[4 Q9'[':D<"IEZX=MC43*YF#LPURL9OQ
P62I!T&:4J6:V#4EZS9B-"M<NY9I15X><A'-$=39W^'@S" 1I)LW6%"^SN+([FDX[
P&$-UF5)N_\O#ZAV.^D8C-5[:E?I-_SCL 752IW)ECP>HO1FIF0*B0[-USG6-R178
P#"HFJANP;" OEZ)9U$2_EZHV5EQ:4J,O16\Z==N"(L?4[DM0;2+D&NI3;%(4Y[O;
PPV"O.R)5@&,BZFWIZ5 =%<T\$OGR*(4#I0Z'V0/9!?V$B]9N!CY8.H,;($,)GY]Y
P=(4L1U.C:4P\$>?@E:PS@/? B][/J9+ ]]Q?%X>/%.GN[PF&$*;Y3,T2G;C,-"/W
P(?>)]IM+D"M. M+2T[P6/C\DW)(_C$+@3^D?N0K Y"'O!R) \C"Q%=%%MW$P +"N
PF& VZH5&X3A.:4EQL8RJ!C[L."BH^?^D<M!04!#!TY'AH"UBL!).X%(F$(,W]6LB
PJ*M0808H,0W9A4.MC454.0A/ZS-!<(8GN-3^?? F(!ZY%??*BIFR/?YVA@1\4@;H
PBUK-J[NR0D%";]($FYNV<\/$YP,Q[\57LK]4S_"!^\6,":+Y  4/)=ZNH"V&M.*P
P^3AXDEMS/Z.Q5%U'B?=Q8OT#]9EAB4O5WS9VJ6:SY3AU[%*=>M [*Q&#_0MW:!/L
PG,JDHZ>0H!G'=KFFN!CJ6%4:?WAV]WNIC=*^*?4F4FHX-'UH0R]\5N%6U5".?$!/
PY *"AY(:V\*?32&1!Y1$VK2' :SFJI39+2=>(%I1GWRN\!HN65%J 1OO80R,MP+J
PB1/O8*1RQ.)Q]E+Q=6[SP7SGN6 B3O<AT_6)(#"UA46/ZJ[]Z-O3/]Q6 @[7S?R:
P+;!:$RT,,"=OC2<B<# _,:Q:FDT7>^#C[(HA#O(B7G7\AHH.?^8C4H:ISV5"]M&I
PA/*D1\U0T)!1-"GA]XMU],NC]#_6:;01P*J3]2&F7>T 1-2K7;,JSVA]ZL03%EF3
P#0<PK;07$2PFK^&:-^6YTV<YLSK1/UIHOF)OMFI(3JE>$GDLW1)+^X]^KHYOX@AC
P%PKIY I7%U6H;SR-&/X@WGIIBL0DK/L!2L7Y#*R.0UK"#"YB?N_G]Y9KP*HU$&.Q
PHQ-?BRH[P/W&6U*&I4V3B4N6>]5W&>3IM+&"W131O@2A$$+- G1@;"K(5[;J55AY
PPR/PJ.=3@\6%J8OO]>X!97+3RW#_3;5^>\R=U9*[CPIFBZOV33VS1BN!JMCB1L /
PA2[C0"#29VG##EV 84'XCE90=J"#5M$$/)HYY+1-H_"C(.E'P* /(L33=>'F%B##
P/YRS?PG%1A%^#5Z\YK8DRY!?,+[[4W/Q5S,,&\%$L\RU=W16^ ?G/7C1(1;D?*C*
P 4A_S?62=?_ZZ>P, D1G[WOIA%E^>Y,L$:+ZO!((38Y/T3.F92L$+A=$RCQP,$-2
PZ G(K#"6<6AEPYM=01A1'^Z>G+KR(&Q]LUY8'EKY&C<\59':'>1JR9RP.5Q @+IU
P HE;DECBZ2-I#QKF20@#9#0&W+?D9"7YB*4A1A%<LVR\S@J)UB+?7D#-)5O0KI5\
PQE(,WV9(D!FHA<R$56+=*@K0,E"X3U>\5ST=9&]WFU.2M%4CI7XZ;!.HG+/>2O.P
P^EOQU]L:5H365SVHV\(=EL: [BK 7?FZYA7Q17(;X11[W 1B%N4J[QV*O&)UZQH"
P[$-R(82?4@H.@00#0DMB\T;(SKN)KN^M[(3_-I'V%%5+"L@T((M$"/UHO-$XDKVT
PPQ)!?:VLB @!@3+?=L;P:W!ZIY)<)A&6ZAMUW'L\S]P+B)XYVKA%(SN"+7TT'!\J
P@H-K0O>K\2K8E1L@%!,/P7ZSP".'.!<"R>F8&1S6[:',(.D1W(6B&QN"..5PNL &
PDE3<_810U;O#=30L9EI1]I 2*'WR@8 ( =V_@YYOHLHX<M1]^IZ!_N@C4$]C"1'<
PP.OJ-U*2^@B>2#-%\RYMX+N4(@WY8QY>B-$7E2@((J[<E1,;(V\2[<.]-$%E,Q7C
P\U U& GQG4F+B2$")_!GN8"X+<N07]B'XTV(^GV==8:-:&_$/]G=:S,MR?\Q%2\0
P%53">66+H2U.FC5'->SI:&]!XP].J[$,[$$A^+L"J8X7WY0<050KGR=Z]%_FQ<WT
PR<3/W&N$R6/\^&N(G'_M_IKZGEVVO"^H!C-Z]Z.] ;J2I1%Y 'Y;5E*"AP!O<#"/
PX?3!@G7)+X8:Y?M'+-B.4HKSU4 616O6,V%G,"&+I?R MPDCY%TZ.!*5M^7C19VQ
P7T?G.?\<9V<<!"H1.\';XI3"6&%9JANF97ZJ>'512GG%\E$P'+E3PXU^R>?R IQ9
P]1I^=)8!&,:[;QJD*?$1O&:#F%!MI&K8@4H& B)RMC2)=$#4  K5)^Z;433<"'5M
PO?MT <P@"G>;88QC+#-R?/!LC&;C''P?OPVOI1(>1>6[UPP%X6,_WO49D3RL8 !)
PI?;(VTQ+6Z;X2XD@Q$5S+J?VM#?;29>W&8L%2&$%.N#U>%)[OV*S\[ENB'YDJ]6_
PXMVPXB65K7'@V=8JP95-K- 37,/+$D60-RA1YL;AIA"YRC+YG\W89<K%W.,ZB5ZS
P6O+TJV!KL\!]]MD4ZB(5TF-U? 2JYEPRRW_F**SO*S.QAI"J3;)23YJ0/37G3,%,
P,E/5@ 5ECC5?CL#Z&4M0!*F,,,2=X#G41+YV$B99VCL7=V7]@9N;=L_R%!]?$:L*
P0,58:"W4Z:VL?W$N:8N[VB8=CWP @]4&C3ML^K9/:'R-#3"PIHAK75W )<JP&(TM
PL +94SQF*)P8T*Q8]0U@^P"K>BM$Z#52,?RU/V.R5TE,!$%)52W3B]S/)_XGX\<:
P2?M7).<9N];XKPC,_H6.+$_E^ 6U6QP <UA0BLT?HD,AM@]\&O&BQO;M/F9>%@*;
PX WP#DY]J=IZ00"MY0':[^ENXJ\UL:9"XP9[A"+!JPH]'*!QS*:WXK#@IMU>]F$@
P!.?U#?32C?]XZO%BEGB=V"M*7FN,T#RYQW_,:<!O7/IR6$^I>,JFT? GOB]K'I9K
PIPBV^]GN+1'!A$$7P_2'=^1][E=*;]>&B_NWS/GT.T AMCMO!%!PY_4T#]2Q.:1-
P W40&/<'K\J^XL&!B755V2BD;V5:#CE.!0%9D@]XE9R3@YFH:,Q<-*<]Z@V3<'XY
PPYO]\6S1^/M"XU/5<?A@GSHSTD+Y/ZSMG32CH.>&:G,FY)SQ7F$?N/'-[1>G8H:<
PYUT4&99A:&ZGN$%YDTZJQU_2(U00PR?Q(Z,,.%VC#2"N+43"W:-M[^T23P,K8)-+
P&0XCP>2Y=XQ]55=6+B@D'N*,(?&2>,O\!0&XQ5!&M.KDB[H@8E:.[W-^YX!Z4">Q
P$A6IVQVFE-4PT;%;/Q23E5)6;T]DJ;#>?8L36CF9+P(V552X)=.-H-4-SI: CJZV
P5&:XH'M9#Y6OQUZ5MN:QY]:K4KS/3N[@XM4#%%^N(Y#)V C#$1TD02O\+\:\G1$K
PU_N9I_%$@+!B7RRWP/FI(1Y)? *SWRY/5]49=4?YR$ZB]J^5SO_&ZKPHX,,<0]^Y
PS?NRG,GY!G0W'EZ !^8\?WSFO2\<1@=_3:;)RE#()^;Q X$9C3 GFE>K]?0.=2)@
P=_ZY:$IFXW'9R:#RN"^N2+)D=F)N7K-W:2+1>H-^/;<?B-,52US&.YU$>>07^.&/
PH;[2U34$F!"KGT&L?2-4/ GK[S<CXK(0D4C$YZ3BRDFUUL*. ?2=-4]!!3T$V"..
P4,BZHD\&9YF_I+]902W:"2%;@LM-,7$S;Z8^\K))CO["SLF;=W"CMP0B(%K:>H+R
P<JLSAH"*$QCBT>M.4DO.$(IQ,ONS5]9-HM&([\5?/I8HS#(Z79V>)MAX-CTFI@7/
PG5:(P!U=UXQG@"KSO_:H%(+*8I'&.[-F26 <K+Y+5?(^>[<SU!A$P/N] DN4:+!<
P=0TO'&'AGEXV'7G4:S:GADLF'$7->53D;T'0-A=SK+!JXB;BLM U*RPG8/(SN*E7
PWC/  =1I0F\4\_K)^UW 8?(>+^1#H>,/2E)9.M61P^I^8!D&4S)W5O/HU!OOQ=(/
PLM5L@\=>"-"7?_B/@#O:9K)$F)WFI60#B7@;T;S[_<._"1!PI-1,ORC;M>,R45DC
PVDN;,Y:$[K)#N=[+BCO6^6Y5G;>S>*Q2FJ@3/0\)49.V<<3"W<N(F:\5AS,*ND3R
P?=B6A<!VXR!J'G?,VXQM-NXE>P.N\I=%G75UG<4*DA05K(OXU+1<?>V2L15XLQ?E
P-=TNO=#G_%3B.YN_9(Y9'8HXKZ8YY0?:-(Z0K?8[Q;M(XQL,/\\Q("'-#\8X*]1(
P6VAKNT:1ZP1$U!Y'*L$H6%BS_9%IU %'9[IY?\.XF4%CU'4UD"\F1KS#'^3@5_DZ
P)8(3<*W?X]KE.T'YZ<:**2K15(NBXFN"A:.I!SJ>VRJS-LR@\BT <1 @P.ZXZ4K@
PB6-Q-7@*Z%I/I448KP&:5=K=0E>-).'V+!K1F +C_;8$>HVE>XJ!OWKX/KI>6)&#
P.=7]5Q(R[$';#>_8_&SI&LG.?#<=6-?_&$_[;F--(B;L[]^K+"U091VY8\-6#!(&
P- $X2LFK"IGGGN:PW @X(G<:N3/*8U$EF9UV/V%/P'GCK#3[6(4Q%YS@6^-OOK#F
PMWJ]1\]PMK?"5#A,AA*R&U$&XIMOPTA[!HHW?[5[U3$U+#)>/I-OT&MD*2%6!P>'
P>#;YN)H@3^[PVAO.\1PFYK+0-M7*-ME ).#5CMO<O!,B;#FHK1*+P89-[3?N.2*I
PJH:8@56>9:CO>$U5QXVBM JR?/^R&_?>GF[1^'U]2?$,JRF,$+[4G0@Q^,-F#HZ$
P9@K]8DS"O9'XBWZ!Z3I=LI&OH'T@513W4(S2BZ.'\D]U)0)ZSC5(8BM88BL)NU1+
P0(\#I) SE5VNAI9\_W>6_8#3#M&=M(2>/JN\PUI'PZ*";(AX!.XG06>@Q?*[LDB-
P3]GWTC((\I02T-MB*+O##*@UR,BBOSAQ[!@B4#,8UZCJ\L2@9UJC,-BA3.X689'T
PV8AEC4O3@A8KX0$/X49/-(PR>$>C@<,!H.)&?K>IZ\]EVV;CIT7A#=4_V>1,J2>4
P%JRSBKH1-N=Z*GB[88I+L 56\PXC((]$=/JCC^RBOT0R+0$2*-Y7"EH++T65BGL:
PZL4>D=4,TVH_>KAN07A'#5,N7(;@VT#/>.P4C=AQYM,3;;:BQ7LXEQ$0K^+-6.F_
PT.@M9S"!O=7_<3!+V'@O;'>@M!/14]KO8C)I@6V'?$:P39P?+=\F!,-KX5M*O'#6
PQO;NXA\?[>_MBB4?#-%-'6CKTK4NK7G=*+5@:@Q55X.EG]MH*B&'CL(@  $@F35^
PIG$0OXN^X.&95I*V)\'A4S&W.%/:;S7;!>$9"]F([$\JVKK@TH3[D"@)DCA-BYLD
PD R_-&IT>3=IKDWHNG]TJBULI#7,\D1.!R2%'F63>N!+ S*=]<=L%,K1W=BM=>&0
P]T9(X<[00:X!_%K<XL>RE+N4[=U\(1;H>[3!K:?,SN#H+I.AV6[\K>.13066U? !
PN'!80<@ZM[SJ9K#I'M&O-45&(Q-V[*F!JD%[_&,'0?RGNYB[DKW:'8;38CP%X+R^
P;P8FL&5\+>5@8LKO]_K3(:/2[;]6E;GGVO<'CRO*T424]28SG5Z89!SKPF1JRDGO
P.RO\9N23)L0&5^JS3H&(WSB/TAPK@0$OZ)4K5C]H&JWG=4'O?2SQ2,8DE3#N:[=J
PPFR[-#%W%Z!.:&9UFN#2#7.++E4)R^9UWL]H*JDV 7^D;-_]E3X?*;+4;:POB]JT
P#6/LK6HS0]<;4^B\PR,C>XOWM4RQ1J GI_1_A>Q-F-ZN!6NG1$N5'45Z9(N]31ON
P7Y$<%]^%?N]P&KSLDKZ/#[?3W^IQK^UJ*^7:I?0[@ '&>2970!&:)&;QLJ7C?1U#
PG@<]^YXC,3I#GZ6/)RQ:D'FV T1*)KAUID&T,27[[/AZW:C(:Z#AP8#NCPQ4"&F*
PA5C)<.3 4F'XU. @^MXKJTRB/^RT;8QLX+"K&'%C"E2/:="KZ'R?@9F-A:T]*#BJ
P0U 8T,9:I?Y94 'U'\$-GT>Q/4&3$SY89F3"E\P(NJ1V=D*:#):V[G?A6NJV>Z\/
P/OQ& )ON#61(36IJ6Y!<0!1))9_;GUSH3; #,VI4H7_37[&5'%\[QL*VY:;D>Z)L
PITPO[%$_Q8 L>[ZH"_4$T.D+=WT,MR#%_:&VEV(&%Y<E=5D);WM1/]8TUP=+?FYI
P<*3%WI!P_>&4OF>RH"M.214KB"F5HAS-Z+B40?AQ[1I\5A_I7((@V#R.$<RT^S'(
P5_))C91W@/914EL5^JO)$ZVCB4?IO-.AZAVE3 (,APNUAI)OMU<-AWH.U>%<_DH?
PR$1@2]07T$82\1?CBZH@W=@^O\S(A0C(>PWT/_.R"L\&H&(>]._U1F49JT3P^]21
P8\D9=:8&02?N6CG7?1X<9>SR;^L-]UT\VH<D _OUZ@)495P6_0WK:FR9O@M$8(A@
PVFXRF5'55&,:3V@H]H'(9:,SJ_"_59AT(\HH08IB@4K*7B'2Q4JY.DM(G_6J.9XX
P"'. Z(WO"2(N71>$E/[&1"UV93T66FPZY WS_<V-T7[PH%'O"^%=BFH!ZKILB](P
P0Q(Y8\2A6 %DN$C:5B]X9^I?&&8RKY[C6M-/%L(>?"=*)HT[*.__)EV.6L-[J"E2
P7O-_%+"C4\V:+2A16"\(2[2@0QX"8^8\ K3I3(CU C+CZ)BU#%IGNLGGU)G?BX.N
P=O( >$QS%I?,#FU'9CTE_4"B?-X7"E$W'EM#9=WU/S$-:QBVA@*G!#M!3 L5/^6T
P 'I_"25%>V4FDW1<Z8%(E,;(&"[=%$8TR2-"G(^ UC[,]W#0M7;LZ&M6+@D]&RHU
PJO;D^@TEZ<!Z<B-%-.-<-V\1>[;V9X*GM10ZV19B=MRMP8<?#B&Y[C]N < 2SI"]
PB4(6H=7G#V$0 >LI&<8;$QDF@Y!I5;F&DGW@[X2E%QF_W(<?0'<8LLVYY)9P?$68
P=P9\%G/,1Q-CO1[D5YR5&/D);*,E'9MW#3'> =/4GV_FYS]/Z&Z$]A#DWVZ4LS$?
P?\]86;""]%!]V+H1DV2D1$O _&..]%.P\VI2G/'.P0*^;)AURB0V<2[:5_(N>&D^
P1#TW =2(/F/Y2*OLS. 6%"?>W\!/^HW<678S6.UF9*\6[+O=LMPK8\G0.D>PSV(<
P'-$&+$$H1^@96YA1= %V+5T$%_]\9<O$&VLDQX?[=U!+I2F1VDY9 8S.UJ"8@G_U
P8QQ'*%0DVAA,E+-.@;!A()V,RD)+U(6\<VA&G6\_\%1-B65QK/$L/G@B_!"OQ>@O
PV]>\+%]]$>M%%E*<"#H(RP!7&[0.JW%;7_NS8%=)_XCT"!EH2F9&UK"PG>(YPXB(
PI7BF6IB*<(VL*/\BD77K&<V^: 0W>PSSC;9C7O5A"61SX&"CD3D'.0P\WQ808_9E
P/ #BS3)4<D(P06N&L<FK <.L&]!>G(0LK=I"QX= 2CB+X+RV:NSH4O;]VOIQLK15
PA58&2BPZD"G\-IKN97.>:@Q8;E\>SA=1)G;U=T2^8Y3D.Z"$/'38$)Z".*H8Q@1-
P>8X75?J24('X%E2\M0QDT DV("BY @_"?$(@;T V\P,U<)?YJZV(_>XVR7(OKCIO
P^FM;5T<V^ETWT%_L\E=%H0Y-2TMAS.YZ2V)T,G>)7557G*U4[R[^.4=@0+=]&$XN
P@A"F]ICT]D>"WOUWOM(&]&5( :9, 2=@?9N$/%%W[FL&,-4*-#._J3W<44 \0W>2
PM)MD_+M6J]AHFY>@'<+05-_/I'X:)4_GI 43-VQ3J),P5_J?'H@AL?];SUN)KZ^*
PIJEM\O.\038U29NNJKKUZH^W+SP&I4YW-/-WHW*I%8M(QP'#S>BYV[&25#XYYZ$.
P1 F=GCRWGRI>X5VV_;N6BJQ1-XZUU:4/4R13&%\Y ]G.E#UJ$!Y:^-">GY!9*03@
P?T4CG1I ^^).]9'N7/9]^2P-B? J^9'(-^IJQ?CG?."89/HWM5L1.;E7#EFBT147
P0$,7=<G[3)Y5Q%3%S8":^$N(/CHND;V\O1@:[)\3(&VO49</1%$3@NVC%X297]UN
P4P("E=E./@^O3-KY+SR0<_("TN)5.);^A9]%^LL[1C20O/^0&* ^L A0M4-*QWAE
P, )_+$)2F6$&.S+'Y\8S67@++6)^D?*^M&'V4=EN/*B U8Z9':<NI,Z;O@UZ=QC<
PQ7JB:RV9OLH9HA<U&2/[UN(X:H;K:$71$*X<150S$-T&L$Q+R1Y:&[PR:L*X94+\
PYF#Q>3IX[W58) +J=5],ZRZ("M'@!JRE=Y5+BKKL]O[)&(Y,KTHJ)L:3MA.>V0P(
P568 X;WPL<9V/V!!O,74 MV?;W^:L@C,O#PYFTILG/8J;%G3<!\VK&UGO1B),0VW
P4G\H-\E.^L5#8."=1EVE3KJ .)[ -OA= @B^=_PJ";,<K4[&/C#R ?\425@:NMV0
P=E93+\65C@,?(0OFK-7T*:C/DGTQ\)DY#8R<F+(!\$B%B^1<BI:*573(B]M6!2UN
PYW#@13?7^"9+[W&]1<,]<]^?#-Q&'OYUYEU7A\1U>]YT=>'F2@GRA<8<@] L6=7!
PV-ZJ=L@H=SI< _Y5FS3_AED3/^9?%%"UM]JD":A.A')L>R;M8L=CV$8"8$C)X2'H
P,GMT0FU<-?LU2 T!37U/_)XP2(#O!?G(JY9-AIQPC/E S?O[V+59Y^Z4$\3/4CQU
P  2-G1HGIRAZK;?1(7 -%K(J<'[>1N[/D*ZE/*ITLLDO>$2(^GND5'UIFN\>>X)7
PFT4R#9URMA!S[%--#>! HYJ#R^;)NA"A\R$ELZP[)L_S4, .TCC\Y&0[E(?;Q10U
PU@'E7V4)3NYZ&EW=M=COFJ+& \?ZLE+H7HS"[E^#CH=9W_[0>2DP'Z]P_" :0KU&
P*\ L)G6'!NY]1AI.[J/%/C],6A E==0A"(/1&]O+GVK+.X+GW;_ 4B8RF3B#[%^Y
PHRP@R2RXF:4CUI<:9_AZ[P;A*=#R@O&0O917.J.FN;5)O6)]U8I2IT:0&Q1'$T#]
P6M(X1.!I)W3HYKKU8^E]AKK,G8?0&G$^69_5HH0$BIF"C?GW2="F";)"M4)2=.BR
P2HR/3(:(WI7BVF$WJUS_C@MFL/8LR"&'M.5&](SX4I'KMW1J M9<M$"E6X$C#9B2
PEP:\^N4+VZTFC[V9=IL3QQQ'Y 6/A3$*;AZ4S>:=3@A)#UDX53H^QYV;=8G'; =[
PA=;X1EBJ_L?-,,B!-K1'=,".R::,7QUP?6=4Y]H2\U<)#.BAN4$.K%F+$[U%IB4>
P7BL20E6]_P7MZNZCSH#.@-#8G$*\8'YC+3S%(B";IZ"ZW72:="P$+@7DSEM67'&K
P9M\/L%\#.'\5*2AX[G:WE#N'+K6Y,,@AD&2Y:0#0\8-9'66Z\]A]ZX^;+'^=95^5
PQ;Y&JG02(@PKBR Z4<U 8FAL)K I\25^GIB^LE%?6CYYU3KQ6$88XC(6"34#6$,<
P=!_BA7U26F\$(_',R5H'6=XACY (8'+F)W+S0W4F"#?$,9&%RO27< /%7R/U'4)Y
PAJ-Y'%2_APA_4Z_,VTR3 \IA;Y-%M-F=WL .;%5N/W92R=N_!>$"4P.!(QD=+<@K
P=*+O=7WRU']YT2+K'C@N[S9>C*,%)P'R+00^:KA*W&-].43F-/E/3BCIK21W;\"Y
P_E-T1ECVE/5X]B*&C].X&JT%6U%5Q!K&^>YK9:O&D%_^UZ5FPFCG(8,B?[.>L(G+
P<A7'&4G'&X3)F+=U8;D+2)+L.CY#,$ =X9\YV0_PMD^Y/%2HS!#2T.9Y-E-V"%00
P7DZCC^-*19D6E  +;UFXEC.1'MD[JC$]D,,@V^=>I 1"PB@OMNH;1#-PN#NFYK?H
P>XH !MI" P47!X#'^;OEL:;=L #,NP%!'8('_)  "S"0F5T+1/;R$-I''OU>MVDD
P; $J7>9(FYPHPS4-0D$H]P*LD=>]$'?T$U0-VTC]@ZC1N YC6>\R!')'0$5'Q)Y[
PIA8,L5 V'&*#C;UX6@3^GW_#0P5[^>P=NU[%JYN</M5*2(UU$7B0"Q_+.PF4IC>(
P@>Q(M\+J'C@])64GM@@HN3OD=BI+T-S ,2K(_.D\9K1C%=CX]FJ\<NCD5G]"<9D1
P5\@]28V83X_C3Q)QL?E <5] F"*&NWR+@K\C5$Q%2[#GCJK1/BRWGH+_8*=BJB5*
P4$OZ]/\P &Q^0+P.'G-:]UB\PA!+NXLK?O_:"F4%5(\:&47HG.W[R<IP/S8)]H#Q
PE&,"!G\ *(A\61.[RQA\B%S*38*9G&+Q:+.$UUNIY:K&M<J8P5BSF-VV\/*Y_["X
PR;"203&9E\OZW?)_^L#4K<]0E8O CK&H1M1HM,)GOJ2IODD!(4RQBU"48M#/:E@[
PHT4;<+NO#\GY\!HP*O\F0._Q=B0:-9[Q*WY*1\HLD_ZF">,T&V7=4X"P9CV M<CY
P"_#0LVN\EA4&7TE^#=W@?-W=8M<>#>G/ZRXF,O(;Z0T9P%U,XX#NI;'%<4_[#XE$
P-J,:119)KVD.ID-PA:BQ/8QP-O!.+V,5"9"D-E$>)E 0>K?H+6B.^.QD:YQ=ZH% 
PG80]4K460IM$@:C&0D3-9P[;=*VG'$X\C+<8Q^U)K]9]%[AL19OL-G[GT0'T>SBW
PBEK?T."@0.5!68CR_ ;[*2PLP&^&8\'7@:*Q3ZB>Z&RQ_LP[J1-:+0S=AXI6@>Y;
P#XM@;EDWG_I9S0:/N%S]V\\06+OFM(L<NC6RUC#D C2@G]TT&W8P=N3#5G2D=KT5
P8A-9RGLS6N S_;@[A6/.4M0T+JU2V"VEH9H8<O?NA6]IRS&4<&&4G6%@E3<[^EK%
P9VY!BL:=>_-.Y%0CH>(S+QG<OZ] /<A\%.=,^HO+48%]R)O.;2[TG*4XCX@<RR,)
P/G(;U468Z?"T4<@;9RI2RP#(/BEKI,-6_=$!X>ZN,%0'KMSL8TPR>BI$/%3[$M+%
PB=HS5JVTZ9],@B(25P#*2::9G&Z)\NJSJ\[H0,EB04$GR)6%MZ/.5S1B&SH5VE"L
P&CK+W$%@-8%V[K_N,H=]!7%P) 0HL/K.'42^ @YM)(@18%SRCCC^UN9ZGA*3+'2I
P V6&T)S6M?HX:5H['N" DSMZM2Y!PDB9M.,@#A$O-2PF#&^;[,+B\#T6#::%2JY?
PXZW8*)DL/H,  L ^94U:59?E/JLXW3M\S0X3BH+!RY.P'*3&F#]3),2QTC#)E+LB
P@?-  @OR!> .>]L)L 8LHIP.(-MK22_>\T .WC6G@*3Z =,K\U+\ZM"]N"P.=Y,&
P+^)5M?T:\;4(:T]7KNA*5'!0YEH;ERM3$YT3G04> ,#"$_Z]51I[I,-:/$!=*4Y_
PMC;\ZXE7IS>XD3X)YW^M]W8"]CZ4<WN@^.5\I79.I" 3%9D/S"Z531)A%\GS9*<@
P?"'(.BVX2=.PA7:EF4G1983M5 U,M*6E H \ .:AWO:%2,?X6SK5K<,QXK6SB/H(
P,[.$)AP$,>6B/9V"-0QS0G'2#BUG+1<P<'_5@&T:8LXKEF*3;J##,DZ4X%TZB>@R
P/_O5C-/+K41#-S$2-=]%,T:E?+HI\Z3+6!&)?=" $E%RUZ3^/[SJ(YW;=(-YK1^^
P<P">^$)7!U/;;NO6=*HPYPM:5<LCR(,Z%&TE@CP[P?3 #=D(VZ2HPQ<4(D2E%Q\$
P?#\34<#_)A*%O0F[-9<^_;&:IA6GJ6]4NX182I^WI<__$W'H$6_#5V)%FYOU.+.M
P8JJ0B2ZOOF6K:WXC2X#F]@ P,P(0:>2 :!@0YU>!H+G8TO W&#YC)?%&446UP?J5
P[#T-@6[2%D*31G0E+ $U;CXXZ*1," A_IQ;G!D^H4:VL_1B,U"_W:; I"M^/>+1C
P].]5-^Z5TIM5A*R7*:\T:FY FY!R$ILU7:"F])9^(#A@&?//7ELHYN6G._WG5)T<
PC[W1^674?@F(I&'CQ)4_6)7@U1#5>I0&Q7__S><W5R-)EY.$\- $E@QB<V> 6J!)
PD+^)W;CN>(757Z(+K50PF^7+3G+&4D+EZ)VT:K<N.-B."U][_--M@LXDN0-04D.G
P AB=E<+1X<^"AV*03KR2:W-(."@BT3@HG[>UD-U%YA[KQ4H"'=_&5L)K'+=<OB=+
P"102F'4QL _V@?#%;(JY5.7XQZ57?S]:U9A4HW6.ISYRK1$?DRSW31"CE1\)YC:.
P=D@X;9 T+^6G4)"-N<7*24?JS3''%4<6_A.$"XT@H:<*U2,#T5!,RI\&1#LVL0,B
P^)BH-TJJ &N.K;JE%DZHX5.J,:28R2Q&;,CD D?$3%7Q#9R,OX86.HR$I,'@&JLO
PZ?S_P,)ELD/>0['&M9 )SJI+W'D>%=*1%_ZV:8CF=2DFAIWH2%'!48W=1OCWL^6@
P^MN/^QITN;DX+VN<("OHKZBW\S_UOKGUP,?^ 2T\\,J\^98E881*=@#6$?NO*@.V
PI><H[U-+!B:N<JJ9HKZM-C".->R>C%.T<.LC!.82SCX(G $7:K^ZDX./'YQ64TCB
P:2\IO@ R6\<)9Z0+=+G*JDN@Y&HN-/B^^!D5FR06902;"V#GS%81:9(G G:)>"TZ
P#.'U9)&G>@PZ8.A0K],EC=6%8Z9P5,2,1P BV/YOT;"H*@J);A1-V-Y.W(Y41G1_
P,1%D@,ZI,C(<[+!*!8"2/Q>\5TG&-9ZC^_@])E?FDW]>_=2?FTY0!M#L:HA?'DO#
PP]$X+IXI2_T;(^,1=YK,OE0$T='OKP@A%U/9>,'WXYW$*P* SU"E<*D>&4F%$:EV
P<]9C<ABF)]:(M9A,@4Y' 1<.ESX"Z0O^]30CM:ZD(U&Y%X-(3[UCH#!F@W.4![/O
P3>-4MH'/K+<,[B87HT%ZT"!8F3;[Y[HA/'MR86H2SB]>?[U+=1'I <L"K\> G%N%
PC1X+G(O#N;>)JU-Z<N\NC PWZ+A"B*<I/1^8@@T*QXY#([@TI>[J[0.%T-C$D))!
P$&2#C<R5T:(]Q@U%8AHM?U'K!7NN&)0!UFT%KM].B:KSA<.4B.%:1QWVWM\\_>:*
PCE8$1^R^>.J-6O"08^W_^J)IV@4=3(.ZMM)Q63!C^9<M_0G-FA?>Z7L>#/[R?CB%
P&HMR##D\4'MJ*. SP:6,:MX[PR@-:ZM(=8@KHFL3O^-A:6F(WZDLZ(KCW,R\G*%R
PI^[MNYC1IGJHI\P O[;1Q+$TN=K_/BW1(6D=T%N=!7!Z0%=O@D\D;6-'5>ZY2/$1
PF_$'TP\*KUG*8,/QX#Z+_;7B5S_<B7?3K$>. CUPJVF6@;7/D C$%Z+1".9IZ7ZW
PC:Y4(@^T0T%V)=P,FMO>!V!\VROI[??(RXH%$'D4<33Q."M-!Y]-H"*1NJI=4B;[
P#R-(Q:RGB50CN(@8+N(L>G^</"6ODB\W>;5@H,A[()S7G]#/B7 ISI_X12E/-L,M
P'*7R3(7CF$M\<!8:575&#>7+DZ^L\,X/4:\D%U86)H!6'CB& 48_2)/9CN'Z-)B;
PP=J(!$N[L**LR U1?NS;BEON6]<R?H,82 R&Z28*JZ$^DMC(_2 C )UJU]_<)!%W
P(FES !L:;*@; R(T[6]T<2.*(U,/3#6"@3T4E:HD@[B\]O($JW?#18W+%)\#=T.9
P_@MNWFN$)@<RB!E[F<@\"7FVET:*84F"((.9?:/3><DJE6'/?"[22J&ZW!R%DD@[
P8\W%[U0Z/.^3B-VLF#Z_P" DBS]"%P%?W6(-VL9/C/O<FZH*)I7/5S=GBD4"J.7W
P&H/3+EW:(YNO&98FAZNTWVQU=-KDAAEZU8<Z@G$]+B@6F@LZQ0OC3?=<J6+[KD?>
P[?0YG]6EAC3$V\^Z^7!"]3ZQ!F&^2EDK_.1/8['8D\B9NBE$*D%CCIT;EJ6\<-# 
P[V3Q1YP#7]?40Y.-GCU]0:\XHY3'04&^D/&=BJ&WW<9ZOYG%O88#J@UNB"6AD/'5
P<0!=9V?\O/LITMUQPY?P#/+4L&H?P($/,8CN37\G5??,/&?E53(AV#$A"SW'X%@>
PU3ZT"?U_U@D F\6E*F":P\+5&A(D)33%&#WNQ7)P^O?3RX2>W;H829B0HK+@2D2>
PKN10!?9-+;]YQU2GHU]0D43/>O3,4[$[V^ON@H4\55]S+=%OKGGH%97P[*3 I=,8
PU\P.Q_WJ/0[\!A+@ ^[Z%0)O0JOW*>,S0"NP.#S+CS&CD[G&7!07_^:@*1ZII#?_
PO'?98G<TE!,/!IE6X' :V25WDWE36'L'"1C/F%MO\<N(E"Z0E<FGYA_N=.?*"M?J
PG9"U?EZ@1]NFK#9O=V;PHP,19%$B/+*Y0;=*< ;GP]^O2=)MGI?^HL.C1JK*T#+(
P^),@"F_./=4,74SQR-G_XL?&(X0,,4+'S0PHW\7#V\7*W<FUL(B3+D6)M9:W'UC"
P=CK3P:>^0;*T*9#E0I_N5)@TK9T-=!&-0KSH^];]8H3?_FLE-52>G7<[H.^XN(E$
P;AB"'N/,>][-FZK6OD[/:42Z&9(\SU.R:\GHF/S*D@F^@.51OOW/]"^)QCM$C\[S
PT!RXIWA9N8$^."AB&[=#[@AT!^ZOM"X?^<,;4@BF<1L:;:OS=>9.'Z4=7T<1"UR@
P6/6,GQ[$K(8XY]I!\6,3B;WLQ!%;&S7][^$G]I":TNFT5P$]U ;!FVR0TG]03;Z]
PYCB9"S++R3K=C7P&Z5F./1NAPT>XM',K\[$.[57XZWZ*?4?Z:JGG2XBW@ B-:NIZ
P:D==XHZ"[*NS"O6MSXDPKLN[^!61M=8A7D03NN&RJG\W^&*IL22O[4I7JI%EP\N7
P.H9TA:U4^A25,*OK452L<:.YN]8F8]&!#\YQLU2R*G'T4Q_3M_BVP'O0C"53)O"2
P)R*FO6UOPVI>K6+=F*XLM_>(_8U/VD?60C.AV!Z;BH#WZH-#@J',O4@:Z&M\$E-0
P5MI6$VW![7?4J&?\A-N$R#\/GA,;EM,7;)!OK[X*VB=&XI%E.(T:MCD=-9(64Z*U
P>I0'YU,8UL'I*M&@0:)N$=*6^)7-40G@0X]YI83-3J-1$3O"O\I%/]Z$B&2P*_%-
PD'M.E9Z!T\+#E?"APG]L=Z+'9,Q'YK0/FTOA4RN(#]"*B^,)J_]\7+*8'D9 0YH6
P:0"YDL6][B2IA3DJ)9:"H4:.VZ@(-=R>\^,1]',%N;-=6ZA]IL5!PQ%PHK*9MTCS
PW+V==)_WL= GP['749L*]:DH/W^Y6)7!1QB$;@G]BO_Q7H%'O*NU<$MLYKQV^1;)
PW1O@,05254%F.=Y"S6*XW#>7R0(8"G=[88,)L1F?<02B\6XX0>!UG65#%C'"AAWN
PV[P2V\;#3;UN!3)2[U7(Q<U8[45!=0NJN]S/[SOB3(JB7WS38V@(/:O&]E&.GIJ1
PR.PW .5:M0@>C^+\XMAGEE#H/^*AI"@W51N8B,GJCFC]MU#4N3^ISA! -.YB98>O
P'D,ES$VB?"'A# \ ;1FM:#1/*YNR%UO#KN,,,J^QV(ET4E^2:<G$3F/*^KCWP[-=
PB:(2%Q;!38*>1\?2]CP1R&8%NS69.;E6*FN1L1;W<$L%D6"$\WY#WQI2?QOC(8U'
P\->?,D,0*:B+=HKC*&\&UM:KU];]L8<D' 5@_3$_:68%&D,1D-E.U0\\34A/OE+T
PSOBHL/O31 77G2.1JJWN,][G1EQMK\ @FSWD6GW.^)8):??7>3] :#)#82-68+((
PSQ_[*Q[B0"$.6^,+O3X;V/[!WHEB=&S><&14(=FB HJ$<\_Q2B-+)"8(\-F<X" U
P;!KG50X*L"PZUS16U?=B;[XCS2;C9*=-B,(E*Y 7BTROCW/&*O5D@JT?:Y[&B/6^
P..^EME,.\D[YT!A@0180=M[_&)Q/%CM%-@?.4F@X&.6,2_E=)Z^*W>0\?Q9,JPPR
P)]>O5'%/Y,SS5W7;"IR=JCT@BY4#F-TZP(9O$M]N7 FXG#HZ8!<-R9[WMPV<+/3[
PY6:EIRB5"N2[T[J]9>+$)&QWIFOP!NXHK6Q#(^;#-VY=>ITD.!/P&75+)U<M'R5'
P .(; _>;$TQX+68$(M8G#=67K0=H?40"$%%@*,?%73,8I 9R)3P)S2^!@S8T,_PS
PZ-FRIPJP'<V.]YH@\,F9=7IQN";?ED("/L5P*V?!@-.N;48-+/ (;'Z= ALB7O[I
P+L[LIZ.;B8\$.DT$<NZ2C.W^0J8<82YUS%.AZ30CB?U7ZOXOG!@8;URAU)7?5@ ^
P (Z\#9R+0WQ===([-N:FBP>*PK+9+],PL*Z:T#<;(Y'C=JR@G((^@S*"$4 W3R*^
P3@Y.S:=G^(Z=4FP!G7;66VL.*GFU9^T$1!7EK0G/Y;VQ\*#Y+>!5$FSF9;(ONSY^
P)J080:]&99?88ZT>_ZW^22']4J]6-?C);2'9.W'1"5X+4IB>K+6R';/>B>>VWSS[
PS5O&GUQ/K#^8X,<B(8]TP'^9658TEDX?S8I_8P4&ABP?+N'7/N$U;SA8/V%@T2H:
PO91CN4+B#@H7_D<'%O6N4?%FB_AQ<\Q9$Z-&YYKD5-XVJ#*_7U+GBUBPTY<I8OED
P*M_.,8[[SJ+<#F.S)&]W)H#==L! ?A3E7=,HP;H0S@X][!%(9'R3N:]N3_\5C=[N
P^-EF163WGL0^]!#P2JI;'^*O6WU:/5AR-*"KJK@5'*!H">743@RJ,4X(QD_IC9=7
PM5,7#L4/@N/4T,-A]9/T'W65>6**!73D4@Z41&!#LU!OO]B3A-R\P.0^ %))_B(@
P@,6(ZY2&VO,XK#K@&CJU+NH\()!+32K7')^L,"WWY )@CX5=$-#B&!UXJK\'\UU.
P)0CZ-D(XTA;N=865ROQ%JX%I799?[!@5FXAJ>WUF">SQ=DU$S?$N\\XD#0G,9D(6
P,&R=^P_2*3$V-$9I3O/6J(735F\ZUEA ,1;229 K10EG=YZ86@F/.S2@>%S"^<<:
P[KR6U&81;@K;93!R ?()(!E5S3_^XR:Z>VP]Z]^$=+^HY"4NB"R.WM%\CI7C.[PG
P<I3PYWD2(_N9X2FO,P#,>KP4QNL+D62IQM4@@XS.X09!#HHSY'D*EWYNDN1@GY\4
P@3Z@XI=J%&2NI7QA'EY"64/-43[FPY</^)-(O9%#:?"(.:,#J]<W/M8LOJVDSTZX
PDX]$!C,^3$*O"FA\I<@#=.Y"1@3H&^H257>09\X-@!D!W8N8^R<1;NORFDXMPC++
P"5::'=5ADR>^OX85:^D;&,-[S>C0@S8I+L'[K]PH$%)>H%M=+V'!65CU0&<M_[6O
PK&N7\1=$E;-\L%[=@'K\VK[+/5:3,<-@K3N%@"8(SCWH'N0;Y#;\YJ<Z;2.KABC^
P&6*HQ@HN+C?P3U(W&TI$C1I6*P]PS,\&K<-+Z)W837!6$Y46&8 2I5EL]S8%K18&
P(*>AD.A-*[\4\!K+L_(2#_LR71_X.%EFJCXCJ:/!)&1X3<(FZ( QW<<A3@@HS]>$
PQ=_)51Y=(JPN?O1HT](A$Z7LCC_#7R(V\@>TX=9#RE?;2N8?2+4,T+GN%)8&:W^^
P\_[N"8ETX- .$Z[(P^IPVE\;NFM^C*4/1DG=!SOZ+?<CLH>L<,0!=UDUO(=5%=ZO
P=Y>8<5E0$\6)*8['6O'O[,56H&MGDG$S!SO%M<9"3Q54[V7CAY)$J?()6Y%/#8O3
P/>COIP=AFM!,31;<MN_Q]!4&Z'E-(\ZC;^J?1+Q%_X93K?>#?VZU1XL@SJ"<LFV=
PQ]P7&'EX-3>VZOA8EG-OGE46!.$&<LG;;7K'TE6'JQ9 #X7Y5PJ:$T_Z,X*!J)<Z
P;.A+9MPSNZ*Y!][-I;\'.?EM+% 3WDVPCOZ2W.E>G-_%[;PJ]&5N>\Z44(P;R/:?
PXKT("(Q S]@=C)#=-:R4PNM.N;4:6,ZZEBI&K^*G?.?>O8K3^>D_QD_+K_,]?Z!Z
PV*?ET/I;2[PX\=?3?[-,.$)C:".NE[.I#8$A%E^F"2,\Y#D]FI?-QTTDZ$JC.9(T
PI (MGI<=(9!;@(5O#BSJ%S(#URSZRR>^+,&CVIDE*DVUB_-U3\/![B@AM.;Z]#KQ
P[N=G)F4WCW@4J&]:&=D82"+$Z1*IN_YB[%SZI8<>/<GO"9=[W6]@(;!.#46(K?MV
PG<[,9+SHI0J^O"N T2W[LX_P+"AJYV8*?$-SS3.+%>48GK\OWK+V Z>QJ!O,;"'C
P ,S2+7G T$Y<,8GI]$L\EQRAW5M@L^$+O377X+N97RN":0_/TU1%)<7-1&Q48Y*U
P.QX2>52T8--7,55\&ZPT6PA!A;+;A1HS.O?+AT&8N.X(']=$9TQKR!O]>EN'"^+B
P7T.KB5H]3 E)0!K28/>6I6H\/-ABIRWO1P;\_X_)883!)*IDU\J1"\O8QL=/HI:H
PO@OF5?6R/.8ECK^*B",QJ'G.)K->=&UD,"L+#D6LF>P,L8/!:+&T1U]V(TT4F@T7
P@7M,_8'=O2AP5<IO]-H:'-_R+K@CB[OF#7;Y)M$'PS)?&[^--4+X(8V;)J^AQE!L
P8'U,@!+E(@Z+ZNF\.<GY" M-\N4O]##0.19IZ,Y+=/%6/$GII75NXNJ@'-(#O"5Q
PG_ET4+%2G*HYYM>7?'[E)GL)81!.P^I@8EW.3Z"8A)?&<@30'B? YUJKD"8R]1O(
PC >'I\X.4YH[/V$U*LS, ?D9F[:2\3_PY5 T_##JA'QGU(KX;N<2YXJ*S:''!76^
P@9R;:IN<UR4KZ-,KD^-RR8AK;D0YLP6VK[%RK[X!PKL8]]^:W5NHB(-@8=4]U4[7
P#5&$>U@*>X1$N]G<#M P0%$[2:V2;4U,9MRFHWXI]NQ0<]?6Z!=#!\]90OA]0LBF
P]L*RHF!U[=7(#?<N$V.ULZ+L1Q)?FW-(HPV5AM3Q1IEG/@[?C=V//57[4EUU7D;3
P;=;)B--U5DW2' #;292H@_Z/VM.X20<VU-D(6(.5&H>*ME17]_V825<5_$,#0R@Y
P^=VO&1502<$#B:Q ^0-\C@"Z-RYDK&K7^(06!UO5%2="59=D7K;D&DI<%&(N<.$P
P)U^R0=_)FB_.H*H]SB!\*GRUFH(58!%#89K9Z[G#R%IHD@Z?W*'^,=\:/^TM_?]U
P 0Y 2%Z8>3C"0IH3&#T*G=6Q=(.Z<C3K5FPIX\#RHD;C/!;$U;NP6=$/<&:#MJVK
PZZ&(OIKG)%OWHXENS[!^(0NJ0I2&-/#]F7;1Y/K*KH5>OWXFJ1]G+RU74"F)ELRS
PO61_KP/I?.Q>4E<6*85I"*U!@=#32 W\JUIR;6.H(J:->1H?IO_Q5^IK=!UDDI!E
P,;P#4QU=+;0C^PE!^&!\M7*SA)[[+:<5R^*SW=<%N[30YB@GNHK6!E>(SE^URTIF
P+_DPNQX)#8T,5)V]"@9N@W/G[%W0M6>550A(2Y =-)>J/))#5Q%;,%IYIEW5]6F3
P[(<^79-U&_",V:\/:.0#V'KRW _\Z>1B:VI1H#5[7$,%X8^O[EDSG_1_PX<E^.;^
P<NK,Y,2A_SZSOISLHLA9"@ODP=_]I0)NA,H@KO\4&?2@G)D- X\3N+\6B?N\!=#S
P$ V=!5)&RKM\A;4.P?!,([LT=:B?UC9&S7P6GO\/&UVT)2R#_T3!+V0QI)E?'R(I
P*4FN=2-K)11J!&[LVXE8_'N-#UP/J+H)34HIEQB-,$)UMFL:%A+>91S;9-(>L.$A
P%[,8O6%%>:@Y>+E5D \TV 7H?"LP]'M&XT9Y$9+*$J\7:>C7&O6!<T[1N&17?KET
P=\]'6&QD1MI< Q)3L/AONCMT(V@U]%1JG73JUT?S@>UZ$..57XR_E)UA!U);XIVU
PO>ZSE-4&Q9*%2^Z:,]!5=Y<;:]=%@V1W#XSSK6U!G4#+%[ET'<GQN.$OXB\!I&),
P-@_G.^!.I9ECYBVUI/\'R8IQ]'@@PDRO?3!A>Y0?.38R'K!$Y\O'AJ37W!Q\[D;H
PH&?_4G(7@S)L!VO; Y,,"C)",;J)YUY^8Z,J;P=_7% 68BBPV:&52Z_USZW [K@U
P+'##<>?:BVU(%$1(X,Q!3#L5Z<'Y8V;9N*99S&\]=L]R*RWQX"BOWA8 B$^*8VX+
P!LBRI'7R,+#9';:/>FSD1J2NPW7[SI3S,O\.Y*>#[/NS-M\]X(S)TZJ_BT\=9,TJ
PL-)B++.W':P(4?5*+KV0Z\8>'=OSAP-;QNL.T,(3-NB.L46H^QNS:J9G*=I*A>Z(
PX)<GN"L TC8P;<T6G,Y"5LROW,AS/X$$C'A0'@@!LU=^U>>.C$L'Y&EY7ZQ 0;?^
P$0%M4A(2D -JU.T+V"'F_70(5>D#O%V84O3);XT;7(')X#/:K=X\-$3\C[7KD@12
PM[>'8)+W8H5EHZ*U6.6E1H3PE,V<A!_R-/+0>S!5B8N-28K[IL;M+'(0' #F?PW@
PDU0W(I&DCJ9V7D*NYGF.=>7Q#\$I>C:(MJ1X?U"_-_!HA5RR C0Z!;A!K&5%%",P
P8MV*S42 (PI+BC\[T:PK2IZ+W4>9*A[]=<W(IQV"A/3 7?'EZD:P=,#GFH\Y &79
P6*+Y/.:@8H %Z-S3XZ%X27(=Z<S;ZV4<4'Z00SX4.OY?5SH]<]UX+MUI9R/WPT.^
PQT?Y*=/.17HL@QJN;6]8 \\:TB*^1JCK>S1HVT#QW.*;6B[83)-.BOM=]7QW D%R
PTAN#KO5S]_XV!5%\'1T.[G(N4?'6+'H]H6O6T</*4_!V#C@(UJ#JIBM.Z'H>_BPJ
P^=\-06I^#5KZ2]4^E*OL,0R_+69EU81>YLF(7C_9KZ&%=4???YH"*!<]Y<2GX>BA
P_I3K_ZF#/=/5B8?1Q6<CAQ>'JIN@CK'[G#636CM# >.?4"A+K+YL-( \$&*G04-<
P1!>++5OA4G;@W##*E^_+?,X7"@DAF*795QP-E1*[S'IE]0J$>RKUUAJ;-1I)7R==
PKKZ=JQ:2IMI*^>L&K:*#;9J:18BW+C'W2X8+<<Y?]WUXK90&YW-LULQ'+?--91&D
P!AZCBVX*%6PP3%LZX+T]@&=JV1SC847*5?Y$3*<G9F("A5Z4R'>K]9*YBL*=56KH
PG]QSN!('VEF"O-'EPP7=O"TS+;VG%*1<F$_+)>YJ[21Z("KL,AL$#0/$OR?:PMF7
P60*&V $+Q561_=KZHS[*B('K; #U_A&!L1/Q'P(I@*+-A9RTH"!%AF$P6>VQ'#(C
P[S+6UV1M19\#QV01$B9<#*2R6N*3$!/$D RX(1<QR'T36H7@@29R$&<0SD[F J2@
P9&)V:8WHG(\=;%;JW*<B?Y?\'Z=85=,"GVX)O;OGR%AUF1YG#'DQ@QOVS\:F1<2'
PA2X:S/^0L&@6%^V UIGS==CC\LZ(VDZ1,9L7:J<&?_>S-(ZMNI=M&OI%O/+JI5$8
PD@(0HW0J<X)&I9E1/NWRY+&N ] YTL".?M#L&\[6)[?D@ ?PC5$U@1F.U^[:X"?=
P/W]8N8D;O2<":3A#<HQ**R-_Z#1@9-Y*T(/DF.4V7(5USD[??MT+'0FQJ%#>:D4N
P"$F7.<TB;%MK>O P6K\),M2+L=L3X,FMU,FBE(D)/ZP,&-!&=A')O$N%38';@4 +
PNQBN"U!PA%JY*<4WR::<SKT]A (8-]R-Y-_SGNHA;5^]6>X^GOMC<D'#6H*/<YLD
PWG\LY&56R@YS"!"@Q:4SMXU!?-S\!,RX[ <X2?;*&_VFX(TGW;250,<'<YF=%1L,
PM\VC33N,9.2!ZE6-GQWGP+JQG$29'!6)>Z@;FEZI+4UV1M68*/97&/ _NR(T<IE*
P JA\W]/8W!EFQW4N$CJ:;YSFR_0&]EL=)3>O&6@P"6*/N=U^\>- @'#.U"IR_Z:%
P*W]? '4DPK6YAT8FSDXF[IZ@"5;^6]&HZVMRQGUY%(MS5HCG [?O/><9N#N7WUM,
PT(S=@O^-(N^@,0U1*=I1S^)-$8#99HIY('<+0]J<_$I5T0-B\FXK_<+[U'O 8MT=
P':]*(%MX%6KG(_N).4J%3G>*?4NDYTDP]0L">&J4?5WPO_TLB6IS)@2-SQ<BG:9J
P+W<6IWZW6:[/@OAJ#J.H#PNW'B>3T&NT_^@85!'$M0Z1.T<GP3S^S4!+,#3_D&CC
P'\0-9[Y:3'R!?0]RLVK,0@B(#0XH_%YF>RNA!VO?JLGPSE>S&:]B=GA-Y "B=QEO
P,0_=R/L>2$/SX*06,D-;BWV\86?41;I@((;9A6('Z]2;LT6?5/8E*O6<&26V!C@>
P/\/KEV\]Z(2M2Y<?"MZH=<AX,A)4J/]<]T#+2I^&]8*!>9Z&J?0'E"N'U93;/,99
PY\M4/MAY5(XO]R9)^BE+5^TKG[J^!!%^U9E!OJP]7^DEP0^]F_:SQ6T\F(B$]Y*@
PNNG_FX\,:@5IM[7,,YXI$4P>S*=?I,>V#F?E_T2:F/^3/TP\V_@:,TF\M@&NN;7\
P<%.[3PP!]40+^B W9LU$UTU,= XIQ;,01?BV$H=,^WFLL-ZS<T%%:,NBI/2EOBE>
PR=,]AZN)T)$[; 'H&\DD9Y$ETGKK!>D>U0 S^<[\A,TI#RR65H<V[/R[/UI0ZU.C
P'66W(V +)-GQ?0JP7DLZ8_29/NH\Z0&6'[F&(5IT>Y[>&9"[B%(]6_,,C>/+:7Y^
P0;B?WV^1E[B8;JIOY_DXBKX6[%>D$/;%5"SH\4A05L;4\[=3D7E+]:DFR)J+F&'?
P];/D<6H62'&$37N9DL6 ,=1Z2O3ALCJBXV=K57@-B_V;-V>AN-!A^NXJ0*RQ.9>D
P]K!<9H=\C9__M>1(':9;KZ?A':=F#\5C[0/%<%(*"R%W<P@7?\#Z/^RNN=WYG-PB
PH=^IQN%\1>KB'3A.1>6^#<[^,?>]*3?!B=,N[\'6TH2Q/1Y.HQG$,4&Z>,_OA_G0
P1=8T7-=XQM<*+-Q) %6$!\;JAC?_4;+NV-<H]'TD!6H43C:03USIP6;Q"5/BB4T&
P4U\LDW=E(_*ZC!>"L9=MATF<M2H)F5? W8('04.LQ:-YWBNGTB-P"UOV'KZFF*M>
P/TR:&AKI#H_/RI-TADT]ES-CK9$ICL^4O_ET(*88F<8:43/"7,)_\F2K5=CCZ'%;
PF*Z/Z,]RSOO8Q8*I0,N_!X6?Y&G.[+?-=R__GUN%6+6V_\XJ:E%('P\ D L ,'^;
P==UH@T%>']5:VV5A1 !!R<M4R,:-SL2PC,K(P,EBGF,\ CL26,8>!"7:DZ,F801+
P\(A,1F>P\=>;U,[3/3Y>8M 5X"9<_ >V7"A?^2"8 02GLG\O$+9"VX*?OCFKP4:J
PL78( LB JLY WDE[?&T28S/FH>_"OJ_C8W!) U'2Y_OG@:S+]A)CHR@FLD -J\+=
P&HW*R]T,P-U0C8=-'MF'%Q?&^@[;_K.*OLXKG1P/A\9&VB!2FS[->EZ ;=OZ?D'\
P#WL4X"LO=%@J\E AR[O(E9'0@^&3F75<X)QUFE8I!//G2-UA0B-7HX1"%:T5?0IX
PI M%:D)AI34\Z#<=LM)L;KYC&:YBVU+4SL;,)U@!6M$YR%['@_6&C'Y.P 0!+GM&
PTIY^J>\-S-=#()T)4Z5:0*1P^(P41R+D\ZXZ,/>1+;"&QLE]+:2 :VI6BQ40LNJN
P6=V:/=(S,CX3PKJ:K.'!L+')O7!<RM\D<9 0%F.9I[B6-)>9&'JB"3MDYOZ]P.(N
P.+@6^^%X12,+IS6SE/U3S,A1$B"9R!/W\M:/5<1J>P &-JKS@T_,3]=KW<-UCX0@
PH\.>[[ D\4W8<8_?@T ,O18B^F>"L<>W@0!8M7A.[/D,+!J7/,=D&L0\DDK$\<=9
PD/@CN,$4LR]]7BW4^;P;P\UF+5!^38=FT@HB)<!S%3A!D:I"\@M+0IFSP)*4\6H,
P&0[U9E@WAYOJN"3\\1:%S34'F7X7'2]04K7W=NI]"0Y4?0G^=3I7<JO9N)RRMF?]
P0N5W$_B<D<&T4S^@7+(V<>L4-"KB0]Z&8$;RU+<#WZ6[O[974X)I@GJ"I3[,""FH
PA<*<BZ!1L#8C0/,][7L[R>9R%XW Z*=V((HLDJCKR<=_<?7+^DMKV5^P$T)BJ@9/
PZ8*F)AT*$J#N9_O9FU13C5!O,2:-T@51.42.0;GJ=3Y/7.X$8MS84S?#O$2 ><@(
P"E,# 6>MG0Q-(=HU-3\Y$I0\4([Q^_:N."8U4P^#>3H_E(*XUIV5?;[2!A[?]ZSC
PMZ7 ^_3PR$*D+Q1;GGW^:.@*\FI].%[5M.Q/(G(ER P!?/+N 5\,G>\P4 55AJ]&
PL8:>K(I38W7U1VZ+9^^]?P)K.<1VL,BP8;NC.I'O&N':FZC?SGD4[LN/KYMQS*Z6
PC05($]N7I]BT<&U:D[=:L>P%KZ:@*^A6"R172-PW?N8^;=*@J#"(:E^7)G]_Z4GC
P(8C4&$_U>8KCI0<R )"S<XT3$55EF;QAZA7,R)?26"9#6)0CRCO49.M1:L>(JHS.
PBEAT;'8 T54CYVM,45Y9,'5$$T(&]-D$+K\ +3A >@@:#X&+6.NCHAE(%]-'JG#+
PKW6X6$5KW;XE W"*B2189#VCLG;PP6".QG*8L*R-CXXUR;U/K>N[.]-<]LR>P&$4
P*#&HD='$+8L3 &=I+2JRSR6S#)ZN3QKF*3KV=<^XTY&B4\= 4["^Y-TGCW?#NVL5
P8!D[V>1'!\::X%Y,9-'EVI' ==YA_QTAN:MJ7I6&2?MY568*(M.:2R6&CU >X9C(
PW6J>(K@2BA_#%+6!L28PX+^)H*BYQ,F%8W+?9C+.*+8B]"M$C\3^@F$2OGU+-_Y=
PQV*'O0"M:^-==796]F( $\*M7TO)TL[<"G7.?>N.,!.A,M X$I7\+KK)J.C5M+[X
PX@D",->>A!EK_PSMJ@?)1]?9#JB+H$.W]+]8A!YAH&7?5R3>WEU23\,K)CU]9>2M
PWSE3M'40U;N?40Q/I7JFA3?YW"T)V1Y-9V+9 (*M[9%^*QR?;.?KF$-4LVWL1;L"
P%YJR(ZZ(Z+M6[>+7 :70.LV%;-LW%,2/6R)A#)]5_##(FWG[&;OXEGS LY"L>>\@
P\Q<.PL)B>)[P#R LD85;+O?T3Z6R""^*&$]G2$@-X='V-@L6#B2TA&[,33J*^Z_+
P-K"K>F0$F/';P0OO^5]'-D8:.P%VUZ#\6_E63"/&F/%#P9E^#^-DELY6,+9JHP\1
P@')JK"SW@PKVPA*2QM^]VAALECW>/W<X5B-&>V[1!AP*R#^IZR3QHN4\M^@;61S[
PD_:7.*IM=>*5#;+\J-H:JWYZ=6?SA U_ZW&1I6UVXT:U8:8YG_I<WAHD'-/(YOH2
PZ:%ZOUL5@&_WM^,4-Q2\4\<*STT2!'\#I.%4Y7ZAKSJ\V&R&\H:1++X4;$"5=HH]
P2MCIXFG+60=D'@42?BQ>_",[UV*R$</=R;- CDM-(T,].<$CQXX6&2'8)MZ>Z@,J
P2=^.C;7(I7942*0LU.>X>6PF\B0A#R[JVB1BKLOT0LCI?8<8MW]V%L:$"073-3KH
P'_7LX_=2"+8R<MULIQYOZ5;#=[FVFK%=S5& ?0$PU<VY&,"D&BPJ1TV#8*#L0X99
PG7[#CJSZBWMB9GW=?2O,Z3=7^TY0CER55\%\!XW$3S0"Q5#76NQZ>SP-=P(^S@7N
P51EUW3/J%)KO<LK'_09HX!1AY*!_9C-T<*YX1S61OJ]8 ><42(#<?T*J6+PX%Q,>
PRX=,4STGD5%]D03DEN'GVL8E3Z X[G@UTROYB@SF?]8Q/6K1.M)C^>DN!$1>''@Z
P "GG"YW?Z&"T2E^I523I]X@$$H41KA+6_4PI7O]AQ S:)4&=W4^? D"J1EGY.MM>
P>TW9\UTK'TUQS2Z)Y5TNSQ^(_'2F=F!3".U)9&('@=92HESO'@A^/"P8 010K575
PISCX9[>[$XXQ%F!5Z#OZE+\3<.*"3W]O9#&=3M\CA9P]>:%D([=-'M;@KQ/2GG/.
PB?4-TE5CX*NO'HX!MFWNUN"- .PG;9\ER$+78-49PS<X3MA1Z/[_\ZW, ]E[A$'\
P50-V__WYE*CPZ%.Z?K/CU";ER>?\$9<ZFAJN6W\OM'LK8JJ\SED@G9J/RF28 DR*
P3->.BTD$F%=HD[L;MWJ![X;)_(]&11U5/P-DV/_@\!;1@PIG/F$DR-F[2+U4V8&4
PN]YH  S4]QR<IA/%LGXK'L#=JL#5K!S?SJ5J]E;Z10(Y6!N2G?U[$C_,TNEMI)[S
P;[GJO)AR489<?D% T(9VA3K5N13C!7 Z(D:NE:N()@8$'UF!-1B!W*9)ZG5=1OBP
P<.=\C^::T!OY#"%4UP+'MTS# :K>7?I+$V6:#SA,<.0:V=*R0B?X5Q"%FJK,G!W>
P[FD/-G C";O?6<@,VJY3"G4HH.8[S6/OZ*[5@S\)M8JWK"KCW6=%_V*]P"(#*V**
PJ,+,8, R!ADW;1=P1N@E3\TJO>[/@K6K6RX^+TJU(\9Y&+2H=35PB7:C_U(BBNYY
P;U$O&& 5UHT1K26XG?V,5$ZRG+5-=:& =1=IVQV*J$7#\BF89'_PBJW+-S3!_:,;
PNGD9K-_YSMORRC"4-,UM_1F"YXXVRQE0^7NPN<7(+)%#CA ;Q>(B7R=\R? I) +%
PQ6'^9NB0.K\O/%S_$TRS(H]FBLK!-X4;P$J9LHFYR9"/R 8#>H L7CSKT;0QRU1G
PWP#B^RA&_CM@9N-.:ZS.+]6!7&ISYISUX\+LK,BY<<%]DHND]I76XG,#:I0"+[M/
PS8 +P]8%_>_XS+[J'+XM&'@@9A?/"GQ%P5HG4W=O344B+TKGZV1^GO:\RDL7F;*P
P69Y:2#>_?S*1N]ZS#C<E+DC;)>6JP<$9LZSAWO=K(]XKU/D?2O@KR@ T^\;0K*@P
PR5=S\IQ;&9FHO>9+X7$0L&CR\$"SX6>PDHIES.14H]DX6TZ*4KH&57_Q*("8T&3R
P9G(B4X0C=7'SB2?J4LK=&5 LK/;&[QP16OX7]4X12EQM'8#J\TP5JL1".(PS@][Q
PI0K1]'\*I9G_WRU)K5)4LPHS2BOM+G<J^29)"[H8T(BJC,+DX+<L1LI8$03;I 3D
PR3KEJS]^&<J?6K'G%3Q@IRD'W=A$'CD,!'6N.NUEBVL<TV8,I[?]&\0FY=ZX'SY3
P]-OQ0QP?D5QW7'FT5G#:R6U/YS[R;>HP^)TCG_RA ML')RQYO&B$2<=_ID)KGEEK
PHIH8.V:5/S7++VMHA/*)O< 672J!'!8L8\\H8'=EW3F<%4^' Q*J40$3P2?'6F+>
PC7Y4C<T;D?%OJ$4$GFBZ;:C._X/Y>..N0P78L&3OU:C.*;,:QWAKB%<*)_&:DJ'L
PSE,/?]E8E5%WGH4A M:^Q3:I-\E**<.>N=MF?N>!8Z1%5ZB)EQ(,Q\GZ#"R'J+H@
PB+AM2Y=D<4(_L03G)_.$S,@AB%X\41'^W=*D4/QW_'YGF%7,R>Z=Y 02J(GG2!._
PZHS'?C;N5GHGYZ]=RTF3.(FM:&TZ+&C. %(3K,[E>OL:5M>IZEH^BAR+2!:^L))V
PYZ\=T[8H'S^5%U;FV!4^=[=<6F/RN?#'V>[9_]\/P&5,)L3B_ 1WEHZZK9ZL#*<.
P_2^(.BLO\=]W:U<RY'99D099I39\:6)T=BZ)EE;D1!24>N*#  P@A&O?FL7YCK[<
PZ;I.VOX=$AR3$PDB44&BF/<X.8WF= /!<-J/%I8"'.*O):EQ[T RS$4%GQ@&?TFE
P[<JQ2:UT1;*":(GV8,IPAOPI:#@CD&!*?':+(S%^+V*"R9W&DZ4QE.T+F!X%CA.8
P9W99F.9[@!-/*TB155CI(C']H(1Z1'DAMA-9>0<(^W<6=9$W]SWV5:HOQZ/U5!B$
P'=;*[3.;GLS]O:DZXUCD-MYVN]:O>[BF'X+,=H(SPW*(PUO %KJE\B:K+EC%(9%S
P!(.M^5ZB^5L*T2>V&,;5#2=Z<\K5*+SM^3AM5SFM ZYWFO'H%(@XG)0/O5V#GKZ+
P)?-<B#QZ(&!W.@@L\4\*2GI+G1B*K*.G8P,P^4Y_>S/<$&\H#/WFN;/G$>(2?*."
P=$P H<($\.F@50,P^SB#FN7H?Q5>O*HP%T]0%9X!]<ZFPXZI71&-$O8BV7%E#ZIT
P^]>>96$->KE,%COP^Y[E;4:).MW>VCN+DY.EO(9@X_^7^9[)0O62;G:PBLC_*]9#
P?K1ZC"(KXQ[1+53<E-6S(,SBTB+*QO&VY]7PD8*F6%[*7P]7[*%#DB)]3RMJD^W*
PQ 1TI1<)R+X*65)+/C0?C9XH94!*(R!+(88I3X52H$8RC-+TUIGH!0LVG:B:EIB0
PQYR']0M'6XQ-D_A-)TI'#K;+T1@45*J0AZEVR*=.YBH *WGY*=SX]J6'*<"2SP':
PL@'YR1^^YW.,J&^9ZZI%PRM!4J/ 8R\NPE/J?=-[+;OH*BQ[Q8]/YKL(X2$/';TH
PGK[G@0.1>NRO#L@QIN>'F<-)<<(_$M%E(?I!M@,(I4!/W[QOG@G(>DC6Q"@X,3BD
PWE< H ]4]$R-%L__XPU+A;%D6*.KGRGWY6FUP"]-(IM'^AAS#_>=N O@N+#\+'TY
P"?Y;V=52_2-&%@J//4B?-+:"-,698/FR<\Q%0BTZHQ<MS4'^*XXC;Q=PX>]YLS>3
PJ2[PB7R0O.7#:)++!+ #9&K@ZLEY<@&D+O3(VG*[LD!PX?IC%5AI7LHT&472(+YY
P.9B56>G]^6@(ELG</<E;(H]?<^[$W5EJED]Y2M"4B]^KWTR^:AT-+'OJ<+W'2]OZ
PKCBQH&="_\$+KANO=4/EJ5#KJ=K'R9JJQ_#1)JZ'XVRSPCR%%?G\<PA 9)P:K!P 
PW488L69>I1:BO8O&_>=R*V_M3 SK#RT(_2:A&:>$_?EX/Z_]]V$08,?1D3N=FB\]
P;!,?1P(_E"R5P\=2XE$B7HU D>L@G 84Z%?Y U" =]0?=Z+SM</<8K4QIPWZHH[X
P_':VKC2P-%QEK/,]ER*=Q!0*W8992M!)&<N\3QCA<M?=C]%OPLU46TVA>LEOQB&/
P<->7.;;72 HJ:Q\V5(XPG&E\0-,2P<N?4QBT\S'];H&'8_N$!=T$1+BOC&VY$</Z
PG4<RWK3D:"YF=[]F #RG'%K&/CUQ#$K/UL%C(>8U,.%1F?FS+- \,T_0U:+,(55G
PJI02M2>V@X2(>?]MCTX##\?PKRLTBW"ZI$8>E@0@Q81>L3OHCD^N;->>4Q5-7XO&
P!>O=OYS*Y6[71?N;1:PHTGFH,9 @%:[\%:2><X3_95MCKW[,MM3PO+YO+X(FR.J3
P2,\Z+O,!ZY7T[MVHR\"_6O,N8!:$.)!77#/N[X$3A8@TG<]@2=(/J(-&C13M&02G
P,X-DS4)=^S3VA)PP>UB5ZR4LCA/D>,>NEJM)Q*?PE(U2CQE9TLAN)MW''3&00P,*
P[NN84@Y=:P+.OC)A5T4FMXV5YA_V@Y/WL51^-6GDA[!*<UI0FEO&#Z8N^G973]'<
P#0&,B)1^E8HG/WT4'ZN]X%"Y)!8S>-+W,HZT<_-CK%,MIW39QJ),$;%-1YV*]83#
P*QT_.#B^#9!*ALD55]FA^NBC;::RBOT6<5G?VR_1*!&X3GC9.6+P)T./@NB#I^% 
P3,C<X3"V9'\.D.&((""U72Y)_@U>I^WQ*H\6!K0*NC]V'A""XWJ N)[&RD_C!1:&
PJ%K4Z9\Y0<VL?*H8^HV%4,D-X_#*C=A/TM@-WI2ZZ)8E#]6O$=[Y3O<C(+.C1(W=
PN!J&1>@*&36OP@[FKK *"KFN2!H*0VJS%]:UOXD=+3.P1^8,I%*A^L"4@I^0K <C
PGLD\NGR%8N9IBGO/^5/BPCH39*I[5%F1[#K203#1XT@._+?KO?4]Z<UORP[AB2*/
P1HQJ146ORTXCBGP OJ,)>5_($@>*EM[_PE4%0>)TBOJ8(K4N(;)K%?!@0>OBSHEC
P&Q\BH7D41-S:K133G!UC ;:%&'(O=>$0#VY4E6A<!5B66K!C:XUA:)%7WMM14FD*
P2Q19U\RV'PXE; [R=C28__C\11QD>OJGI$;W*?<S!'GPE:C<M@P!WFPD=X!$>3&&
PA2>&P3Y@U0Z.%=4\DAAXH*A85>.N((,<3.('ZC3_:2-X&%&+8M0KN+&@T/O<=34Y
PUA/Z,0S:.Q3@0_OSWTOFG5@L4%KU!OBE+N;<78"G 1849*Q*;0F"IKQ7QUJ*9LS-
PUR],S,=WFZPB+C'RD7#^+^-3DP6-!#=3^AR:4ER4W3),4$*QQYM#; (Z0T&94I;H
PA!RQMO4)VZ;HV@?.Z%1?72F75&^4?ZW:ALDN\8*;"81%MCO.19/O4A&X#9\ZFB&#
PRSK1T[IO3>WU=:2<#$+DTNF'A$#P$(^\C4H4&=(D7WQ?[DEP"'NU]#S>SJ4^/K(W
P:>35AI]]^D1=!O!IB32_",Z' VL$6[D?)-/&!V%Q598_G#\;,6ION?'XB=%R^O:_
PW?\GIIIW;%*(L$6 '/<7L"P"BF4QUY!R,&[Y<*%*WLZO#U79,+=DZIT]FU,3935$
P@HF*7:+8#/]L>YR!X[4+E.T+':O*\=&N1)_L3.FV9<>'FB/&F;UPO[S8>< &1^08
PUH; B6RD/Z]&O'9M_DHZ^O9M?X7/ER0 =:@ \ ,EJ97A("V*_!7+"Z _C[DZMV16
P[LI8L9*EJPV#U-M1]!-:!D%_E7JRQ/+1/I74O>Y>H-Q..@C6$.LK6\453@8X1PIY
PORD";?**^$BX>+(?WAK\4&G3:D<OK7#?2;="8$F@JS],5\O,3P1[,J>4NLU#4=0#
P!2TIIJ@QZ^$\LE6F#2V.CD^/?AL;%<.,8?$^JWL%1GB538O/5N6/4@[:PMT#V(]U
P5@+1ENL>X#JI) B-BGMG2W)N>:O&F>6OU+;1"XN -=^MWW[M+OOW?:X_#Y30D"DG
P/EI)*HZ UXPOQ)!AI3GY:/R=>B]<*NT$8/D%9VCR@)PTQ@ZV7R]5/D:E66W#8J00
P=/SV;<=.*CZJ-<4#FNN.ER.ZK/0 'D5[=@T""S8WR712GZO6O7@_$=#4"R&N,'_V
PJ[EV_Z,6P QLJ]5F/6W)!I(/ :Z)1NC9$X.JBZ$N\4=[(G%-JKYBC'D#6XL^AV@T
P.3!8BM#$#G+@E5:10:&9KNAYO@SDG$B'YN6HW\T2\5\3F^5_JMD6#XQ@5A[0K%+ 
PD-4;'B]F-!9PD^]^<^1W9LE S'O-;+''*\UO@SN/QC>C/+"'H./13*!O_^-)@DK[
PCB;F$,RSO?3#>;!,6EH%A#9DZ0\UMF$BAF!I,QPHX#>_ U3:5!Q3YP?>98C1(7AJ
P[*NCL2Q"K+W0C88N?^N&S:2D=?6 :%DS7W\XVG&*SL>*-#[P7.!,FPE*'5:X)ZX6
PV$+=;CZ3JLI(5$GCU"!*(4'O7="V3@5[Z,5T]1O6H@QEML+_K3&]TD4)VV[U9;_@
P#,M;$D%!_M3#FN?H"H;1W>RUU'PT#X0 *<R",<(EK!/G%/%FT$O/4Y_=V'[+,VDJ
P,(&Q#RWXN[1'-B#]NC-OC**8<^1*DZ=\<5[Z@HO4R"8A<9173*:=19&5?7UR580V
P>HB/SK^,4@/ 7PQ0M>R]IK$_DONX\@YB"!R=R72#"22-849<>^@Y@8:""?_6$QT*
PTFU --W!\.AJXH]D5.=9BO="PS*(%)6NH._@Y&G7JEH'F@!(E[ U\\IY!-R!],4D
PRL0K4>V6J8[!^WULHS&/'G:/6BD DZL,G298.IJBTEX%73B@:FW#G2F('+K8@WZF
PFUCGOLR9H'J/ 48!V4TMW%3V4H:Y!<D@8(N&%5ZFB 086CL9L3:83AE;^" :?@'S
PW7O$RB+:WA0N.0.F] K[$_!CC,_2I&P,<+GF5DK@1BMZ4@?0T:GFR'L*O%E^S,RH
P<1J0+5J1<CR#".@1CY>_+;AT3F1/RRJIMA'63F,![%^GS=EG3BR[QW$*7WZQAUVP
PNF*V";%U5Y0P]02C0TX=#K*+%H:N<CH2% -,3V5PA8?"/ZT^Z,ESFD3K\6@/)W/E
PO$WOHL$&_Q>O6Z<Y@OC0.L=S[@_HU2MX4"[LBB--I6^G?#,2W$K.MA!^,B %H&43
P0/N&MWOG_D('$(2W0KED"I^S+'O"$I-.*);%QQ)%[..!W'+]"DP5F,1)[J#D+HVT
P?#6WK&N2,ZE7=OU]7@_-=,('Q1TTL2T=\+&[L_X*P#?<:3T$E("O9KQIHR: -.VE
P-QAIH7-/',HTE[% ]7?56QL]/ X@BF:YI;Q5!T&3B>6H7ARRB:_W%%$;\J\05<:J
PN<HG/HA?_&XT./L.->0\YM#X19<:2*_"P_G75Q&OP4K3[Y[XF1PEZ2+A3!4J4()^
P\+!FMV/?5]NV @];G5ZJZHF<#A9MQCN69'2#DX"/216OA+92T2]?E7(+;J-HE0M/
P=\1,6J]BA02$O_Y[*DBI^%-;D"6^?K,\)L"<9][%*DN-GY%4?D[&G6?0GUI_MR)O
PDPLSH@'WC^M#JZ<,TX&WJ<CY?AUB]?4B LI$X @]K%XW/).$=H[CAB'U<5X'4]X;
P+'CUS+?E6"Q!PDLZY,P;F^\8;Y-_@)//QR40N=>0Q/BJ8<O!E+K5L2 _ZX6,31_,
P%F]<TZ!;I*9WCO@7:1%M/LQ3S1 ^%[W1(4>#="^3<,BN#EGB>>+!Q294,SJR[]UU
P:;0!+E,C>+_'93#%HTS%4"2P$,MPL]V1?9L9)6>H.(_61]!Q90"#2"(P_)U/H#0+
P03WLARLI^R (6BUJA BJX)5] A5\KG=%#=J<?N'TLP AXYE9/.X:K@ +!EAX1J^9
P388B@P76VM1LT12WY;2^2CR+)F"D%^/]_ECVHA\@[/*C2>?/?V;D4F+!0^#'CT.0
P:]:J=\(4_SL.".KW=3;/349KE6%H2P#^D*^.VA.<$H?/!S_6:\OZ06 P:4K;9YME
P;TG:)G80%H2PKC.*F,54IZ4\8VMY>E!CWDV G9>=3O,*V$A E0KJ\ >6@>(H,W+E
PU9!GQ6HCB)+ .4Z %N8E>O,6.&X+K[>)UU)1VD0&BR>HA=.VF,/56!#SNH-6N^%T
P0H.PJL5Z:BWT/D30'SFP,N!D6PQ6/OKH8H7]'F18?9\':(>WC#+DF@7F1>2[Y_6*
P>B3^Q;O:DS\&#T/\4!"TU6<@(Q8;N>!V(/.#H=J/-3;ES4 72:'O&M^]^4U9T;T9
P?+'BP$1!@B!2@DD%^I4>G'D5MR:0N[ \&XY?(;/6\,!5<IK@L@1+8IT^%Y#'^+_E
P9TG6I'):W"330-T:)$%!_"&[,IB9Q0;L3&0B$[Z?RH4OH@B9.@C@V-S62_TJ^+LO
PW,U:C+KK$GP$-OSJYLK?NBA2'1;)<@&(.!"-?'S# ?D$@C D0HFYJ)!T^WX;RQ>>
P%BES9)[V<><);?[-MG&$G>M$S!@R+IUTQ>N(4GU@5T)>)VO%*T(0<Z; (3C$<$"&
PFY2>K<9"082]C$75@9-=8J%X/#%0S*Z5":*5'!H\Q $ I!WY(]&Q1BTFUO^RQD%M
P"\;%VCQZ[A55 VZ$419L:CGKAC>.J@2JXMS]6;/*H8&52+YRX*YP5ZSH9&CJ*\_M
PVUBI4#K^+G2E1-H0?>-U9W>Z]'\K=(,RQ"OKV +9'PYQLF"?_,F78ZB\#EI;3( G
PW;PL#XAY3NK7H;=G^)&$;W*IL74(_G3_[%'X6ZG9)GWX$[8,,&W $ZX4<M([U2CP
PXRQ'<CISK^%%&(8,W$(3B>4*UR18'].-\";50MPNC];N/;1O&3<IPDNJUF'K!8RJ
P2)6^T?0J#JTD%$*/^1-2A;!$VAOI- [>&QP<K9P0T>.RH/P4::OJDV0F.2B<(FCU
P.3E9,;O:IR]"$%7^PLCX+DMX2'+*ZD!T])(6"'EI@'CX@6@!>H=VP41,65(*@Y= 
PQK@\(=QR,+B$@D) #*4;!8UN*:NSX&:*7S]HLB70(#SKK9HJ?)6W<3T$<ZYR5:#R
P=*'B%;.&LKR]2OV;<#FI(['C.7]!Z*G!'*[FH% +6_I\8KBKWN=J;*0'/E-[;)J 
P5,ZK.8[G@"7#44O+VJL0<1[FX)&HDB_+R<SUN $ZYUA$,OIB;6->(*DKB;2Z?LMT
P4>[ P?>1[\_>2(JI+03#<+7/Y "1(GI:T\P>\=S+*I/K1K&Z\<5#)^OCFF=/BVJ0
P[7:Q858A>ZJ'Z4128KEI)L9E LIJ.S4K*#F4KF2P>IA^AS6/Y9&]8+;YJ\""4K:+
P3N\G[P6T4:GP\!W1$3'-BN ^EG+8RY DG'^>EVY/^P0V,E:]2XTP7;EA?17OI=IU
P;]%+)P0Q7HFQ^>;>4+0NP)%30,58: S-:+:[<UBH]L'[8!R0<=A#S.<L)UHT0E4J
P;USTW]FA%R3KY-M\T#0N%I^*;5<&64\'E,-GP0BU1U0:OB(2JE(\.!;_CVYS1KR4
PJ"BU>JY=6'P;1N&T. QU]VPE\:S>11M[6G#."?U1.)N*JH E%#&MR^;0J1W=(.=C
P,!IF!2&BQ(8,K5WK%YCM0/D56#AI< #OL95M@FL!=@CL"J8(%-V3=X+$N/H"6Q!R
P&%'6_ 'KIWF/G-.;49_6;B:F%EA3!-U-"A+($ %_;BF6-["%!8FC&Q N(MZ<X569
PW6,K6BKLTKUT1<;ET&R'B_8)[GGKQEW?;4EB\,A?BTEG.^*=0$H,U*6_TU8>5@PQ
PC>E15!4\\$= 9'" 31=>J81LX$0S 9U,&!!W^>N:/>]Z5\#[S*;+=B U:K(&X#[)
PD05XF&QO#:EJ\/G:HT:%H!2WK@?XWT08ENUK .RH3+^OB R=B33;[*0\@',NLP1S
P<4\4<OXU'$#"7I/@UGM0X31X2H=([;]AND@271S=[*<5#LC%G0403CD@C4<+;@Q^
PMR2>B3F<%@QPQIO'W,K0Q_L<7S4_RQA=^V/^KSU$T,_ALD%-L,#F#5'ZI6<QI\^,
P(Z0([)J!#PG +6/3?3?.N75\.#DLH@ 8^D[E>Z.(*%S)?.<IL=0\!S7D&>MIV[IS
P<41UHMTQQ@V3\P &^^ HU0GRHLYQ$!6Y?=Y5:L^@6#L8!MB-;1:W4'Y+Q19AK3WQ
P8YN%T=%\A?>:=E%+D4+CQH!+TXA,C==Y7ME;$7Y1UD]S_H:\1C*YZ>NTKMSHA(8U
PW03^]0F$'@%$(8+CIV"CI9-($D;1PH;!AZIA<T&ALS_3C@^Q)%N6)"C;&5*88"E$
PMC=H>H47-[/Z^3$+\&LE"B>3,/I)P>,BO[6%.H%KMCO3DH,IJ;- \<[KR-N?OBH/
P8AWTF@U/=^T0D_Q4%+'>&UD#X./<YM#/%@!_6<&"1C'TS)^C'QQ^-),@A/271K?"
P;\H%MCM,K)C^Q/Q(SNIJK_QG@WN4+97QQ3BU9<['ET@N/J&.,>/B(X,5U*[H9)\H
P^NFPBJLF7%T@#LPECEJJE=-;,C,&5'*=:6=@'=,K'C35<_5_@MBH3\UR\:FY+!$6
P:G 9_C*>U\]FU:NZ&BD1+ 7'U?J?->H2%?,ET2=P;E_:8((RO'3P-.\A(OBX)Q_4
P*A[2K:*QR.";V9^EGEJBB<2Z,U/;+89\;7A- C'>(+=[A+:94TMOW*=^0[73XH%N
P90>SL(NQ]7DY%'D>'F7JX##?PA^*6><*)%KG+]]/BK;0=X*9A[A^'GN&VG,"$7&%
P"Z1C%:EM$E'3NH 9>!!U+1(AVNMS.[.0+%: ]4_S0=R):'R;N/0<7NM;JL7,TJ1$
P8+$*,Z2QN(*W6\#2/(@WZ\L"[W6LNI!1^&ZZ9!@F]WS"K]:+3)0\QM-\ZO:UZ:;!
PM@;U8PYMP[9L!PX$T>K(4#/?TO\3+YK]B=]#]?T,;?K[LOPG8$;4V:B1I VL\\;U
PMF$_:?O=6K=[=:_8OMR(!E;8,X?E@-R#V.77A]^R I^_8W;=]P3_L"CN&N#H3?%_
PF\ 6/@SZO'+4]S8<0#P&":@CIT+K\ZE&XD3@*HY2@VDRRK\<1$(&$\&.VPZ#X/O]
P*= &=R?1)SAGMRTN\LBLGE._YA?V"AR4I:*:=V\QAJ7SA.BI4^))+Z0\EEB:!>12
P6MTF9<N](%!P;?R@V\2 #AH?SD%-8"9S7W,]FPIB1\"X%L",$QN^CM@]L2M$\*J(
PZ.<Z%MM0H#_B@I?GR&,E!?V2JBM1XP<&*2?:6@##?U9"@8+.V=.+WQOS'AF(\3*:
PO@+)U*$.H+DJ^XME,-8(2^_9#2B)U,0$]VW(@7QJU[P$C3;D2Y5=;.?C4!TJ,P7?
PC>G??:R@-K5H:4PMAB?C/KL9YH890B?\91N !3^FVS35ZT2GI?< Y@!!_R0E#,YB
P48@_/3*.6C$8(OLV^PQ_H57F<F30SP)%\X;=C&IXN83BU-'J[N*5S$V&\5\RVN B
P0D8OT"/-;XN,24RWMHDB[1;T4T)\TPTD[* %9:O!02NT-]&\W1-+Z[,(_ ,I"U6O
P#L/IO*\F 1<A=_<DE_/L,>)'DO(JH_G=K1O.XXFD-G -?0KD.]*6[AQ4ZD$'_U^,
PVDG&U3N92LFO)1;')40-T0N$<^65P730R"/[@UIUP. BCDHR(\<_D@B2A(DW*&K7
P-1= O%\=6W:0<DN[]W3W07KL(\9P(HP5(",4*O?P_\O'YQYK?V9^<HYZ]*CO[-,E
P.:;A$@_\/=F2-CMM<BH)7(S60B@9VF1U!8D;E!7$?X+R>WP:"DTAER/!D7V'I68<
PP%N@:\! +8NQ(Z ^%T$$NBTP%2F\.I269 ?+[7=-NS_[B7#6TH0QOV>Q;F'I]P[<
P)Q2^0D,F-[K>Z,*IFJ8<8!5 ,GAWFTNWF@U>N:=6WX."B&?7PR>@#=-N[^9K/MEW
P$#G20G9"UB](A,)M\$S\;H_%DD'Z:YYXRM&#.[1/P.S2NLP+8JV46_;<HGN[ :4 
P+VX12 K-C]Z9FEK2C!-@J9^!+Q3\)X3QDU>MCRO #WN^Z9T3M%80$0T^!ZY%QY<-
PV(ZD(%* 26A-^ZU:E*G@JRH#9MX,WTB^#-=FOZT6$<AZD_U4YL,Q4BC;5R:F&^/P
P929 .<%5LS"+P@5%RQOD+VX2N3 AKW3RB>*(D;@<-0 ,-23 9?*ND:+)@:62EYI1
P+6@_$4)&X;\P,0  5_JX* *D87[[F5C%"!9W'<I\&'9G+Q.$A_?X4ID3<)J&8%QE
P;9>C#0WJ]%?#"]4\PW=>A0F5AMC"*D;&'<Q&X[##'?!HU9N+##=]G407C<LZ5OJN
P%4>/*Q9X$I=6*TFCCV>7-Y/$,ZR/YX2:V0E9!:10DT+B%6_3<U;%&X!W#-@8@676
PRSQ9B-UO^T.9<ST,<JC6VP5 ^H9=9P!V-,)4?I/>RMPPN$F^A^'%B9'*O>BZ_*IB
P>DX*49&--W67Q*"PBYP$?GJJ75[=<_=$?$8+;D?\OL:2$Y[D/0F@[R#',N<2X#R[
P_I T^'KR]D6NJJ):@Y:-3N[UKFD]"BO3W@G4>94U-CDMN+@YN\M4?P"P8_HN#Z1:
P]=ULB0-M0X%VI@.N4 ]M+-WQW7 $"_7M"87^^$4JQ^ NW1&8P&AA4%EYBMYJBEA\
PK[N+2W$&ZUVK&E9YR'1($?-;+MJ WP 2#(//7OD_2L(_5PO1&*!F/(=<=N*VF8=9
PEOS]8ND#*;#HEZ#L[U+U<X'#XVB 9"0<$5AV>6->09$&NN'W4D$@"Y"';V.9PQH*
P :)U--=$57BFRWIC(VEM7"3K0]^>"1DT<DG&)O^0)J*1\+M3T%[6<VYT$T4NC*O=
P3@D"9<'W&05;]1@8/(4HY>@10WE9U!4?I=2Q?X,DF(V@@9^0Q/F39 ?--[?&1DRP
P_1\?V7L2I" \1:LT#@C#D[P;(/HZO2=*"GJ&[HI LY2"N&FP\"7VA^5W$G3[6$L1
PN;"^6L*BM=K (<W87?-X;Z--Q05 +.*N?,)80D<$N0Q_"S2 :H+?"B"@9%HR/;*V
P:UYNX@J8!+AP:<-OUZS9UGGI2"R;F-\"P/M5>LV5NA%[SX)1OP)-^^;F%(EFQJW5
PV3##[KC#U\P94-7 @2PB;[0]LIN2ER(9CSS BFC@(>9]WK6+B WU4@+OZ *#1&$P
P!AE S;H37WT0W%M^(5#D_&]+;?O*!SRKIY48MIAH=&6C)J6875M9%PIG&E/K]R<Z
PDX5@)/UREBNTG7+EK1AJ!>G7<>:)#F:#!(N\1MYS<MIRM6D7#X-.K3 *B2F#1HD3
P%%@R#M]@@%[YTU5J(P9IB375_QG\-G=@TKG1:;K6R\/J2V#>+BGQRDQ9=)<<WIS/
P0E.%ZEE7^';;+6L:^7:$@]\?GHNJBS'8ULJ9_-!3D!RID[.PY-8HYS&@,5B[^'+V
P1-_ $X<_:O$(IB>VO8"6E!BCJ511GK'P<^.W5N0YB1IJJ01-7*]A+QQ'^@2]2890
P=,#UG5%T>$/$\'.>@M<?=1P$J-4/8&RTNI4;<T.CDP-.):'>*Q"2-6T$\=M1I%:4
PC66$U6HT[[;%!Q.#'NTP7JI4NN:K '*V+T(+VOU/1I;.ZGK!8-#4]^$8**V+RN"^
P-!WA#%&XHKSHZZG=0;RH^XU-:V?,YU6E.1 2%N(4 U\Q1"-V*&-L"_:Q1"95HCMR
PY#)+MK2>J,,JG*H\I([\'KZ,[8FD0,ZN?/:M(%\H7&_=K=C6KNU&\.F$QILJP<](
P>]2Z/SW[QX6&="'IIA:045LO:%K]"PS-=%YSN-K>CJ3^3N1@@'30>6A,5ER.F'D+
P/S1(=)O#R/B.4T'LU#<#!PIT_',(EGXH%LT]#[F*]#X0_F&JLO#!\]@38BRN]0P8
P@[>UZL29/DIPM1K5[."XFQ.RGHDAGD4<?5VIXU#Y]7@R@D0^B3"U&#")?_;/W H'
P_T+PULG*]%R)-W77B4/5N/8%6NMVXXUAXH /6?L)/C%R!KW,:L3P=Y]XR_9\18_7
P:D5:SE%0X-8_DTW[K,6WP8WJE\0/XO5X7T@@ZE)U!@*4&+W#XY]T@\D&.K/V2^]!
P03-\-9A0&L*Q7;&P.LC4P4WUYR >P54BA_ XZ2'#7]3W5)C$938P' #VT@2"D:"F
P^84*>4_IM(N%#FN1&QLPJ(ZV:IE8LCYQ68CO;I0$%\#L0,D.%@U!TA&[W?BY(X>_
P9);!P?]S^W;6'OA:$S7)XNL9MPL= P>Q*&V^FSZR30U>8PJ!F/4G <)Y8FB;'%I*
P_R_($5N:2"5-QN'[?^9R[! !N'-)PEF*E]L"<64-B0G[8<&105'6+(\%@GXIW[V'
P,EHRG>$Q:@ C]-!PG%AITRJ7FYP\0ESV'H1GC0'$PC)-[,W^I74L_+EJ1CW!JYWC
PD;\BJ))204SC6D\;5OEN<&_T)^I=]@9Q$K<"V9Q*N"]MG2,47U'TAO72>GE30-J-
P9F*7?DC0>KC (DCG!*QQ)\A?X_,7.5_% K"[M3;G,5!;3\$>DI4X2=E(OF33:-)"
P-F,STX&5CJ"+5MCJ[\>F!XQQ'4MF6K"P(35)W:Z>34DFP)3*T32Q=@7=LK*'45HN
PEC V8R2UJ2]9#DW3V9.;-XW%LY-D_55B0MQ;GW0(G!]CQ0 ^,+<BF&%R=V8F_ QP
P IPIXF_JU*4H,!VO.2N27F1WQ?3RA$Y-82'2%ZHUCH6=<,)%<SGM FG0AD8GG!ZN
PM*V>E0<D X4-M6F0H*3QV V,+2:3&IX58]F@H4G*Q;,M(&N (NP4]MQM].QWA\)7
P-\$5M+T:P-3SESN*=[T<-#[NA(OT>7.WP@)(^Q(R%.I"Z-RXMULO5J,I;[S>.$DY
P_R79AP-CY@'M98/LWKG&#UTR8,%-O09AXOG#\9'D!-?_,6SZK)XI!#7XX>9TLTQ:
PCE',+72;\Y=4H<)5S=H<_1:W)<5T7VVJ"G,]D4[KJ0RGE2?)78 &AT!%0WWF6\A$
P&XOA+IH#UM.T? +P)ZBA2KZN'Y,T5V$#SF>(7Y+Z^2F\JV][TBQ3\@X2R%HD]4K5
PUNGD0/<X,8DJ20CRWU\ F]!4*KUE=+>\/6.[<"/X(2YIIGC[FO(*%:I:82R^%+E+
P5Z+3'E1_2FIZZ  3820V(;E'<T8!(BI_-ZBPKEF30OUF[DE$ZI==!LXBD($.U[8L
PO*CN7P,PLKL>@,6G)*M,,9FK$N9G06<Y,LAVT2OI=?E &]DDP!:6Q NF]D5B4WQ,
PE4Y+;$];LV/##[97\QU3ST3$+R+;66-F9=OST'$5O/-P$83I&UP^/_0I';A_1 X9
PXOUKKC1)9BMDMO)3OY-L7"_TX2:VC"@H<C9+H'#4-R9,U\9Q.[E D== *W]"$/?+
P;.WJY1YY?*NSE@+'G%9@%:2V_T1S_03%DY!AL[7;4MS#08GWE3^$=I<O3 F+^"9S
PG()EM8F]@2W&34AN55F?K;?DW,9'X1X,Q;,6FURTCP_)+[3G?DF8;;DB:=W@8'Z5
P,]O%QP9WTI3.$IF#1%F6F1W=:&B)O/=$*4T/A7*"%XA.GL>2:[:7:KH1^CMC!XX3
P2P&,?B;85=K&HR2 NJC4U&Y#&27.C\73SI<\V&6"AXMQUZO>%(0CCZ' .)F\J?[-
P2]=XE]\0.R?OIG2Z)9))\NN3E0\L'6;/1"TI%^7YO<.ZNI^)6.4GDI#ANW(!?D.3
PC\Y33+R=0V+-H*SC<$FVNZXQ0MO.+64,H$JKTX4VH:?^/&0[($C.Q:@KL_^3>Q/@
PF/8<#5Q'L#ZZ-G(?D4YNYW2@4K_>!N*9;Y-8Z0&;E8X<&V3WCD!X]146X2<+3L^:
P6F(U\D!NS7ET6IW.FU3ATP3_/)Y30>M%SJ2Z<&U!P_--4RR7HI1)@XWQ=Q;SJ!DK
PQ.5B:$1L!P4[$K*NC6D8U#3&UB8YEH][)B58W*!F:)8  .6 VMU>U:!C/ ,?'PUJ
P:@3QB=??D3PGFH%V0"8.A6 7_R/+]B><\M!\S$ 2\@BB/V2F 7[^L34X&_ION+84
PYRD[@5CMWI8XGSFLQF^BE"$RM7N8L;;UZZMYXH\WX@X#!+=@GW7QP2O'SE$-W8&G
PT:IH00!27V8AEPQ7FQS:(.PH5!Y4-[)\:/,_T\=':?WGC%AQT,9UI<D0?^;& \SJ
PZR[-B. ;,5"/S-,BQD(&NY5:T62@D-T=0\=;@52;@#(_1JXB3)=$9=)QCS7V8/X(
P6?U#_SP)2$VOQL"?\'LL)=%IG0H!AK59!T*U6MMBCS+?35DJX[3([U(+%O*9ZZ99
P+EFPT2G:%V$(\?DQ509N#<^J62C8JN'P^G:X> JQ"NXX+;1)G-XBTR*P?[\]+^\\
P(5R33JJWFPRSAG8_T]&/&;!1\?J_6^EZ&0>\WA[X\<C36C>\MJUH?18Q!U?B.A"O
P'_4O;L"_5[J0&XGRVG7BOBPE8::-284:9WRPATR?6H.8L^5.Y,X$=DX^/1F HX1/
PV_HU@1+3,&*JJ$%O<.H/VM<C_AE_"UU -&?Q=^SX 6O;&&HM(^*4W3C&,%QF S"T
P*B41G]>M(B Z.2D/ ECKV.^)M#7WI0 A0R\EI?PPOF/B-E_/\'BTQ#B9J$$F9FEO
P;Q 7* RE721J38G9CZ'AH;P3B#A'TC.5=("GM8A$!/;<:3:)9#9)FUHX2>-7<-NX
PV)/!HQB"&B@#2?##%@KM"IU3#L($V?R1WI5<<8O02D@(K%F#*E%\YB',1CQA28K!
PVE*< $F4WO[5RCL>;6?NN@6(^8MOS#;"QA.Y9WBBMO5V(Y*L:^Q;!;R'XG5Y?9GB
PO%^[X'2%).GRP6,5D&]I_/H\'E@*B=H4S89GP$9WSUQIN\ K2 &2J^\41)$SM)9&
PHFTC[1QOBR7"E:J]PJ6)\7:[N-;AW_R1/F2(0L:+Z<@:K=-<2 @QKUT9HP"9$FO_
P/,8>D'HR@[WOX%G[)?UJM,VZIS(<F=W&,L4HGFS^[(JN)&:9: $SUP_*C.!_FHL1
P8L/ 8]F&LR^,SE4P/[.-CMK(<JI@@$(SN6GAALO8%U)[UMJ\V98CX)Z,4SV;*3Y1
P\F@SZNP&Y?=RJKIN0MI;9U]FH_&?M>W3"W#+3XG)O&$ANJ/*H,,%7\+#O1\#:(D9
P8 S*5 7$HZA1^^E)V) ?"JYN.5*49['VLA%LP64VV(333\,:8%E/-+\/JGLU\%_<
P8J[N(NF_VAB8-NFYIULX]N=$OH'MW[KES9%;8_(P85F[HW/KFJ'./[K[P->*(\7S
PTDN-UX"YED%])>D(X#@%<6?^:_6@G;M.Q]W+X"[HCG@\\K@UKR!NJ7GB>@[VR"1L
P'9!2!?\^XYVW4^;AGK]E/_T96 ).:5(N!%3USEDG)!TUO4K?[KH-;$2MC_;7'YNL
PCW]U3T_3!0\#]82Z*'7&N3#6%&[-J6-MY_$^B,0VB8./;'QMC?#P?T@NPK7WWS04
P$TIHN \C2(M2+WMO*/I5\Q1Z:T9WOE,='N#=Q*44EMSK,!'5YT9P@5GL8G17H\YX
PI53<N2L^MN086%Y9G(17E+#\_-V3!]1"OL'$P3C)H5]'LFM'.++\$F+BRQ=NA[@'
P;J:9 GKC.@+V!,'V+X*9-)G6;<[DU7>-*MNRFY!5$MFSVUVFG08H*4QQR<,-8B.O
PO]FJ>[H:=T@@G3))5$38"'+&AH15'V<) LX;?!%':;1G)6!]BV<&26 &N"T9&$U!
P--<>V;P>T?ZH7'=B XW&%APJ=, /ZW[5&RW'V0]VCQ5QWL^_1L_6[5%:D:0::9P+
P3&$@"C/)J_Y*NDO1Q&2%/%2='8ALOTK_<1_ &7046[U&"9JKGTPH%<F18LP0C4P7
PARD8JG-MD9SK%TG%UQ)]W6A7* #WCPJ&N>?$5L,X=O*H];J?7B4&'S."@[<U>Y':
PE-9@:^6E[H4,G"B5Z3UFD!Q5EI=QO^-7<99Y(G((;LVY:GD1%J2RW3<O6<X4:Z8W
P[>M8CS4AEF1G%I+>"UB-)4;QAB,1DXX+_QB!2.C3ZHDA'>6@)'D7)P!?&29^\RK@
PE(+3VK,@H'!#LDT6EP.NR*4TL%%YTMRHPV^GBGRB?:XK]!NV=MV'E2CL3>Q(EJ@9
P^8>EHJBZ#MZ8_MG09^&1R6)X)R]#\P +P74"RDXX#T#P]5Y$15F*8V=3FK,@+@&9
P&I40$RZS.G[?65@D&DW- 7J1FDB"I0;;6O*@$=I1*!0IX]^=2XD7H<Z@8W[%"^],
P%@.<D_W;&*[?7O/]Z37A$;7%A.N8CDY]D2GRYOXSGL,LM5XL?SP!T\1X:LBRGB%A
P!MN(%VO]-EF;<;T'+N+[:EG!'&'F#P4KB'4ZB=7J%G-J &2ZCV)W=$]^ CDK)0*E
P=!N@DLP6+N8OPN0S*BM,CW7$\BF4X.M%;N*)A)1$>MQ[4[ 6V[?9. X@OS',*?SR
P<+H4#US7?_'1W2F-$T91XNU0E=J23V!US340+L,M2VFVE0]B)0=2GNJ&DM1+>X.Y
P%C+IO;E>'KMRWTE='V'3==8@[%TE<&9 W3O_2]E(N$?WRR7!P/&@.HC6"7&$QX*$
P4&E[;-7?R9QFA-LM0E_[@A5Q/%7E)]I>(0P5 :^-W?#3ORFD;E&&Y0039:=2GC?T
P9%2*; 9DLHO+#6Q%\V/X?S5$.FA2EM)(?&"^8D&C7A+8V?90"[6$'_A[KSJZ5;@9
POB$UK0N/SV["BO2)#2ZA=U?8%!KH)\+<HGK_C,;&V1,P-AZ<B/F8_)(-^I,\='S2
PK\/J>P[\I8F76%>L1%FMU5[@I^#@R(P<\/:7D9T\+F>$G[H0A:_'S+>Y)P5(8?Q1
P.P7H?17A>"@#SSL^^FI*)#G':E9ZYKDIZ !,: (;7.TU\+L[6U?/ JF@$BZ^%<O"
P7=QT-4:L%APA$94,#>VK]IPY%V5/AT 1X4A&/Q,R>U+*S@W;CS8DP7.BDV7%[<5>
PV;FBRCXX(Z8DR+6TFG00+I2UR H0/9W-+A+]3^-*]!M\9)FA@=T+_95 @QS\N2P:
P7E^1[&T*X,SV?1D,?TQ]*7F6_:M)6!6_EFM'!F^]4:+^&S8:DFNXIAPGL])!#GJ]
P3#AV;;MHBIT1X$=S='&0^] Q CZH5*@YR;[T@S<@CO!9"<OBD&!L'/T3_7& HYI]
P4$FRYR'%%V#(V+R8%'EW9&##$_I;&P@?MW>)SXNMXWW^^E*@9+9,Z",T9CE96MZ"
PN.LX\1^E%)4VIE@JY0'/ZS@G'X"1[XL:YELB?!]!2[FH!M,?E4T-V4LAP[*D],Y(
P9J(J$R2):[:M@>"9N<IB:5JK@P? A=B?%&H[D?!!$&B<TFQF?T7B1052F.SF26<%
P;L:$QD7/X<8&GEBF8[_ 9+&'#9[D%JP9$5D4?8,)V8*U/)9R12W''N6:'_O2?2-.
PE^/DJ;99J82B.AP-XX,TPX!B"-2J9)S7/IK^,B8;%=N1@"^EJEQ!^\^%MG2)!G)$
P92<^*:',EZ?;4=H8>1Y]=@.P"C?:MJF=-^7-!YH?.;?$ '/M4#%H"32]L5#'U\QL
PN$RKQ\%VT3W$</"T_ #Y24)5TO+)9JEKZ/6P<$>2>205^&Y8#A2,H9^_0%)801/X
PB2$,OQ=K.-JOP.=MV>J,LD\JO_W$*JRM/ZJ-@#;%T,W$4^CMB5QB-+'-W=T7=)^O
P*5Y KA)MS/Q8BH"DRL6;H._,REYM@]=^ Z_B8!9U" RQ>PEK.P%324M:?PF0QH=(
PUA3@3%U?)E HB*NS=GE!TG*90]Y 0V532=R)O<XIPVX=#SD+^>;U2%\H.%I_?^RA
PD@")*'P7SOA/ '(HP>]7!;B<Z@<>D,TNI:2";\X6Y[]!D3X$^+K-<*+(%]H*SIFT
PVHN#/% _I2R?7G8(ORR@N?F1;8PIY9G+Q"?=I_ )(1$6)=W"0JFS$MYD=J23$J'2
PK#M3EQ1IGP9M]-D H"Z0#,*QJ.%C@^C*]J-3*80?^A8%C5]'8 P-0&G7=[9O%S96
P@#X;@ $D1 5JX&F\=W-H0&.:ZH0\QP4BDU")GO<,^K44<VM8 KRX0!,X>J7T5AFC
P^[>RB09)&&6YVJ(>,=P]PXA&'TH%[EOD-698::#0G96$H!XD>=AGU)3<^-4"0FZZ
PO7A7SAPCG2KE/F:@B57/.L&YDRH.!/L)33*1O<EKVAL)6&=JEN1W:>O9H\J ]C&K
PNRW,>B@$R9.B.X6[CPX3M2 $H N3>ES'RNO:6[+G=&28HY]--[5(0Q.J":IR,%X8
P5#5@I\&84[-?%\ 6%9%B5CUJU<RRW4I46'UN?MTRYQ=@?39</?W3)NQ$3!0N6>9^
PM04NQ:P''8S8LZ1!*2RB&0]G> LV(73P,%<K>JR6IG; X40 4#NR'XIYI/F 9X(T
PD'Z0O9OW 5-L0B9?Q.";..3;M_$"VO*>_^ +MRJR)"2 VJ4>?PT\Z]>%.U[#U_]T
PPS(O;4Q:/H.PL4%1O>F:M5-3/<X\*RY_]SNZ/*?B=)@(\PHX<,?\Q#')6@@ KF)O
P(DX,V4W]\/>\I!P<M-GQ-]Y-!C,&2*9'3ATNBM&^+53M)@.7JW)':^BAV/.H^28A
P?-INN'!9*4S7PU_RH%]9;SD=_E^$C54F(%REU1IU90@^L-49W:X,*E\S^AB-2S!<
P1RS=TP4W3',"*2;ZN%4T>'+S@P3=^/)EJK9H=A-L8E$40E> P<(E\^DZ1BYH3(&B
P+0*5C20?^/@BI] 7=3DN(_PB)BAIZV,&AB PKH$3R?"9Y7Q>_4AQ1D>[Y7P,7M$Y
PF!J&QE>WM. YMR\<6_1<VCJ8( TJBDG6HD/XK5*^Q"ZF'AGS",$OP))")J3-%ISH
PN1G3-P5)NBJH"G5,]Y%"8"="WU-4]>R2MEL Q['C':?K\.O F(W20(]T0;FH=^7(
PGB9L"-7Q(I&FD+-;BS7JC^$$*C>/ #BVSI!](N,:%EF)?@_$WJW'P!E5K'<3T)"C
PG*=C$&,?^_M&-[F>2*2Q0H."W: H0]F5IG;!4_2;SD=/(E%) .#:EXJ+<^_2G%9\
P4$]=1Q M]TL#?NX5/W^?@@)BT+5#@FMT7[8#)=4$WB4 K8,?SXGN9O:0.(EK&R:E
P0)K "DZZ9/Q7<\^F4B"_Z>66J/ ;TXMFOIE0:J%.?K$(O(6Z];@97GZB,,MB)@'K
P_S(_.4U6?TUQ?K7<T>]V3("I>AKZ/YK^$F ]"A9.SBGQ>G1+(E]2#$(/4%95P6*C
PLWH_F4K,>_YV5A.4JG2CS#PE2Z0T4<DW(W2:10O%<),MK8WNWQGO^_"TK$,4 Y#S
PLDW\ZZ7U).B\;=N<<*O58.:?&E#>5!)9V0SV0KE&UAG \EZDV@?.[VAS0::Y6DR<
P.'M:JN<SDG%5P@D?^3[S;HTBN1'[T&DQ&TK7+>DL"%<J6B?HC'@XIXXA\\P MNQB
P_C*CEGV67+:*"1:8.)Y.F@2O1><3O'?#60J$AQ7XT?,09U\<S+X%1RB6\M'8^89(
P8ERDJ%<J%5'/-G]!_&!N@;.NGQ[=&&.>O#Q3^T6T5PJ&+Y9K"7"5RB/>VC)8+OCC
P(,9(J^25\<^KWC+N=\G%YVV:[L)UN]^7$9<BII2AY([: ;>4_ZB4D:LB0&%==A%+
PM*!$KO4O/0'-14]YL%.7N]YOEE)1>1@W\&$]5!4;'\E^&Q0HC=!O;?S2,/Y@U)(R
P1JPZ5Q:0_X(.3/MIQ35U3JT++>5/G?+OP_,E"X3\N#*M-F7@F'&5JVI!<=R8>?\Q
P8,L[N]0A8N;+Q*K!HH/]W&-"T,\*<)LTRJ)R3IMK2$ ]< UL67OJM?N>;ADX/H8V
P-@')Y#[.GD;5R&*]EQ%L25?<L*&M*&E$[ B33X\<V&"T99]^9L+SA>"5)D\_XQP<
P'8--<D,XD4D5#$SKFO.:W?NRY#4/#IA G9'#.DFN/F%&.V,[-J&\@@^=Z"3Q;#[ 
P6D-O4A@F=169X\3!VD.(;\3QQ,)H^JV^^A(*5&N+.RO9%V@]UU*J>H(5Q_?[AY7M
P(BZR- A\0*?W,TM#8'N#*0E15I_1I1N[)E3CD%1><\A^IG%!BZM%W>^20E;1@Z<S
P#>)#$TB6[J*!$YL_":^PI@W:J=66$_M)FS5*LVN^EX.VTK?:$1^/L5/K]2:<4_=A
P5]5-#FA62VZ+S06FHZ];//.0"SIV-5A\[9FY#(:G Z2E$7(+LU]?#.PW?NLT-X(_
PV:OD+;?2*D\.!<Z)_5G^IL)RF4*HK6=9LLI5U;8\MC,I"1W/_?Q= CYVE.UMJ&I^
P#:-:A+S%J#K)>L,E H&L<@#BU:G+F/6U>)4DF;90S=,+SJY7?V$Z"]YM5&K#8(A]
PQA_74\)7=2-18(^0)JE@B8CI9]ELCD5QW+W Q:RE"_E\JS37A E7415-()8DODN 
P6L09@&I63HS>6N&>'KP">ZPS<PKO#K'%'!N>B>&-+(3'44@<)#C!,%7EVK\0)#[6
P:O6JKN46D$RLV> )R 9@**6D* ,R)IX:S*-3H-S">5QU9LW'8CA?;LY\AE5US"^F
P,&>*/;_'FT'(CK/LQCY._8_1Q*^3M,?"H'#=1)6Y#GHMFT<,7PA@B.%S*3\HMFE_
P^^"!/,]?,3PIO,%DZ5RXS/T]TEX+?9I:)BT_=3F*NMSAF*ZVQ&^]EZB7Q%_]*M^,
P*5>.L"=:D)#AW0U</7S\YD_FA\#?NE\UI5>;5D2"FNX%V.!]YJ0A#%PVII!CZ_&P
P$#:"I=(@G0O_DB(;]'K*$'7(+HDVXH!?DG8@*\F@1L\@9QH^++U1#&Y;F4WT &PB
P[_0\8([/+2_0+\?_/>0!0MU]Y-DQVU; .7L<^\ODT$QWTJ];;<0J2+QBN4QSNZ.D
PP+.<-6^E=0^JT^7?+[%=,^74_Q7.*?PM<#Y)W$"98)\R'&R]>D90'TWZ!HJA#)VH
PA326;/U@2++# _4#D[3/\Y61;IY=3H0JP"U<5BZ>?SUF&I:WR,,QVI]<#Z[?=?50
P0IZN7N)GJ:4A%RL1NFRA'==#(])3V9N&J_>*\AZ^MRXCS<SO.?B\4$LU( J __AM
P7G<3=_6+A65N$ AU&:CLH(W4$0B!,!^2DU]%9.35;E(9;WM>EC\036-3J)\D&]-K
PN0.X</E$.+")V<L+)5,C;(V2(B05I!GSC4>V4?A?QO@DR*5R391R0H2. *T@Z6-?
PBZI YS2/(<EXMXLD=;]\@C7.%N[?$T1CV=3XC-=?.7J"P7I07B'7]^2ZK"P5 Q*W
PL+?J->B<"<6A?N37Z[/([MN;KT (%*==0DB8#HUMLMA.;E9<%C*[>Q9%T/G\#'>4
P7]*4QJF7]U4/8EAUB0>%,@U*(2DRI <?[,'AO=)B ,2?*P;04_/B0F4L8,H.+>UW
PN5H]EU3=Q.B-"9B'7L2F+(YZ,I_6'"\Q&I^-%\JOYB9F,MLC"Q:?&+:0!GX'T0:Q
PLDEW2# T:;COM!+OF./W8 8,RYU@TSS[]F?GWV5=C<<J[_]BI8-[V,JW]?\WNV8I
P4A$+1$?A(#Y QNJ;7EYF0<UA1UDJ.!?#%I&6@7A5[ZACG\S;R';E<;VEG__3R_C*
PKOT"G'>:C+\OR"!K-]BC4?8>JQ0: ]7J>?"D$S<8(\RR?]*9E[GT?,IBN%&2T*RT
PRCP\J"#NT"VEE+71-2'N(D5M,ZQW'1*4N7D< =3U\RQ2%9^0EK&Q#B4DY?OSE$-7
P*3?!N0B2U'-AXI<HUB;9!&DWO*"$53)MJ2U[.^"@1Z &N'9<XW.1Y,65DH*FTENT
P=44@^^DU$X%J$%(9AK_P)H%BK5%K_T0K#[!%R5UGIYWT*=GO+XE^%J2.U OHJ;@*
P'CJ@M>I>!NM%]:(9D)J'<\\5Q[;?3P0]TA'(IL[]=-<Z1;73LZ(Y#@6_Q=_Q:ET-
P&$'M< W5*N= ^%L\C1[*IID+.[5?NG#,S/L[+^QC<Z.J&/=$9J]61[I2-6+6+*K0
PBL.3SHKWAYS<90L= '912!TC]QW:TB_V0QYMW%1^U>\_FL"R!J?'2K?PUZYM6CX4
P[L-^U$L<:%U:!7T5%P$A_30C\J4ZJRP*_R($%SH[M81GTW@/LI&CQ#'N1JK6P;W3
PW=66A F:D[UREC=?KS_"*S28H$)& F;9\7(O;U23\TI0%T*N2N'Y'$AC4C=*G@-N
PT-QTLJ^IGYGNL*-83)S#N,N =UW6^W#Y?_K+?6=T/O,PPY:.Y($3,_VF]MFW[,[M
P*]01K"C8W6NG?\;Q1;GEL(Y'5;<'?U^FF^(!#^\H1]]7PD^]_9_6C^T4Y*^-KN_'
P7#@;J8.W_#A$*O59Z- 3\3U?IT%C/X^%%&7^7$G]GSY@'3]VK7QOPOG7T^G5]X\Q
PENQW\V6TK]VP9AV>)$[0D--;:UA04)3Q)1)YXN7E89_:]7,S&3$H8RWB7>0ON,(?
P[?OC1$8GUT,(9#"SULBV0I(OZ-R,.SD(1L_VDSP7>)XF:XQ7WI6H<FA1M:+)$CU&
P<A1 9?OJB)M.U.P)CN2#6W@JX]W#'V6YHYWU>F,?51+37CO (A//1'_K-\(_2I9O
P#K^5GKQ?FE!GEH,DOFJL -;\?"8&TGW[NG_8WWI1^M,N5ACC:V95ZX(^$4T1<=$O
P;RT+=!C]U1! _36#A&:;M4+[TTB\@5+Z@X .##XL.3FV38!*8<0=.$8O8D(K+6F>
P/!)A>K6]9F!VQ9BXW&ARBTF8,BI+78IP&T5X;B98+>#(&8H22TI3>0OGHVWLAVR/
P&B]H0_YL.UK/6^,.I[&G'P7\HD-P_U1=L1EJ,<1N"Y&5"U%S(72K8X=<KH]6-25B
P$V!AM6 3$H*<\]U>84'\JVZB:S-?^Q? YG#2 S$5J,_,'\^W_*'9I)D+PUS*0R,/
PME*N\X?(KJ%9+-W&C:F=9:V]2X<1,R44D2/\\$M\NOO?F6NO_1@_51J\*0)Q:NP9
P<JJX*DI6  ;EP!Y;W=]+,+>%IIB1O$_8<I\5X'*;U9/?3/@^0M/#*[_TB[.@UDKQ
P$\F^M,"!PAZ4M1VE7DY!8(6-%1"ZTF>QAC[*M5'!Z]QBY1Z,_"OEB=CR<+0*D8^-
P7/XVM,XKJ6%.JL7+";)&DENZZJ)W CS;T]L@3L]H<52;4N:]1>I?ZF,&?<^B<^T7
P,4HC]A;*YSYXN35(H\F?W?T6"0V<F;^(6#F#%=>E&[QUI\$Z=\[][[GNKQ- M^ 3
PA!9A TT@7NP_ E%(A>86B5'CO &<:&3!"][C'G\H9@X2'X('.M,%C=Q;%>]>OFJ(
P L[MP5SGL+5 +ZTLEF8%I!7$B*!&][O6;3_VQJ_,4+<,1%@N_=DBV2;I<&W9.S#]
P?0&X;/G,+XFJV&#9CD-;V#URRO6+Z*!\^REE<&4'P(F>4-O=Z1<)Q'FF&N]_%G.%
P;H4H-5A>90@WK)(*') 3F"1&%,V6</(!KTQ;>P?+TDL9)OO+[!3O75+>0P&)9_E=
PE87T.(8UYQYT=I%/K)9N_9O&G3@6?^OT21TN92C3^'EZA&7=YHBDX&4SV?N<P/:N
PZ%O7"%5PPJ-F%=G"_4EK+FCT0@.WR:=<C?98_$_O4O=95%UM7*7!:-NF]/FE?(G%
P5LA71^:%7/Z_7K K<']ZG?G9T0B9!WD?J6?#_AJ]?K8-C$MG?BF7U\[MX3X#J^[%
PRX%;Z&ZN/'5ID,D" +&/1^.[HBPD&&$>H/OXTLM4*1&1 _#1>2)PS\5RM#$9)?/_
PN'PP8IQY'TU@^.T&O@<_T:(1+"=2D8&'OC&:#/H_./<(=TV8?9E6:NEL/D'&7"B?
PSHNU2F.V__H]Q%7MRU '*^N$M,;&";4$,@5$7/$+?9<;C'*%%K'*9@CLESJ]_5YL
P!06IKC:,I$$'+<O3"5T>G@]WDN\)&H2K@E1J _[[:7?VW-)0/],BCHHSY?"[M:_]
P'L<OP\O*_G0H-W@!I#<IFTD2!G6C*<;_=6A"<A=PV9O@4&Y]1MW'1=R=DL 9&++=
P,<5B='=RBFU+-6E.D%B/42D\RQL=>6=,L7&'_U]NHUL9LBIHPST]I)(_PN*;3DCX
PXNH(4\U-0G_Q0]6F^"U_=&3 I(]JS)4QJ@LJK_XCQ_^1RKSZO_0US&SVC6<?_RY)
P4W4O<-I32430L':3D?U^K%412^,*DJ[8<^_"06%IB:]#P9I+(?X$ J\+%L'PO[02
P,R'P8V>8"+H(69F_"/R7V^=;C"I19O:S*.L/P6 !OE*\*C>HXUHE=0'D%T?$M=T8
P=37BU;:[M]]%FJAX5-_]$$#C:(])T&581IV X;^)#V^Z-^'>:7V/!&TQ).\2L^TZ
P^/9QYG[%XKI_8$(?OQL#P(OCG4\B.X9APLT&52UX4J5Q!8+>JN\F6^4@,:YX[%TC
P<6TZBXX(N5>^=MHZ@=7(9 6^L=QV;Q471'/FBB.OO,6FS3%>2NG!5(2%";N3,A?F
PDU($\ U*RL./*F3]_PE25&&+2UV0ND[4N [[*94*BEO*?WL&PR>J91RDH%6TLX+O
P]Q8SEBM(3,QA9I_7T=0(]@&#8A$0I0^I2R,8.<\O9/K&T,(WZ@A9<*5@"8>'1ZN 
P!7,>H0P.P4W*BJ#1OE/931FQ0<]',UZ8559<G%#=L=H,:NWB:U.:93_(;!Q#9+X!
P50_J;4M(;3!'_:_/KFX:NVYU8!=KMM]>D>JO$T?4^0/C;B,W&KVV@@?HJG+SMH0D
P@6&/[]?"RU##O^8C3)'5BMV^?)B>B.90-3CK\,I96C6)220M,3#434.E]\XW+[2.
PYUWPOOMEG^.2K?!%LH14 F0"&+JZQJA>TW3OT=JUR!)9W[Q;HPZ..)R0"2^.<T'6
P6!7>Z%)4P9D:%$:E:I6N'G7&0<5.$_HW$2.7>#_<:!D&&#OSC/,+)(->C/E0*^'P
PQ%"2FZ@S.](U'EJ&FY>N&_RP+=>I:LN>-@(+;BG4- QOFO2JZAY#^* T 8:^YCY4
PC-</)FX3,4WAG I,)L7N&(9('L=HXQ1TPU&?L.]'G="A-)4^Y<H'FH4]C,F]T6V_
P9V407Z?;/N2"NNQ2H0Q?ATVGCJCX1M<6$':4'B"@L $G39*34RM9Z_<[3J[N$QQD
PO$M #LT]Y;'[G/>&BO$%-;IOXSH9_D06=*&O$@;O P2M7'A1?4#/\F &W3+-L&&9
P[NRB3?_Q,=^:.N40BV(=%'Y*S04R"2GO/!*""(%VPW:?KSG@H_/%3IR13"'<0S",
PF@A(V4!@VS: J?5YX_G4R)6P0K7@+J,:9X8OIVRYQ[F;8:#U"PF[WC\J#JE*V'3S
P(OU0[1'4WYG6:+#-1"#=?9=K"S!>!)^*:*@_$_U)'6YC?E3$T]1ZI;$*)\Y4+F_1
PUTZP6*<3ZZ;N2A!L08K$["1!V0*QI>!RCU@@2@)5XT&^)+<).JW29'?#\$9(^ OX
P2 :"\?#&ZB[R<M>A;IV$/CT@)F9H,\-!1@BH6UJ&/XSYDAKA<?HH $Q/@ VMZ.V>
P&IM>E+,YMNO)JUE?"N#5P /5%,0^*2KJM=S]U3QG2PO[M+0-][H9D7JK/>BCL,?1
P1Y'H =! \G:*7 24%9Y<C5OV+,\U6R\_\IGU/'0WG$:=.+,.7%YA;BIM_<KS#<CH
PD? "4+2A7Z2$8Y:;D93 M;)FIU6W]-H3>I:&AE9$#&^:_5H\#> =EH[$22F,S9@-
P0O[^=^AV8._XG,\PM8Q9,F_:(4<#0UJV?D/$PER@LC/9? # KNVFJIV(OG-XK.+"
P9HX^*K]DEEX5&.W$+0OO)BG-VN2 \75_S.Q6R2].21NN'#=WTW>FE#V5(W%PV^+A
PV>^0%%F&DF,KV)OZQ^U3_<F[9MCM:2=L)SMS:^ !_J?X,V;FH4._#Z>M8YG3"'Y5
P?!!_314=!NNCD*^A#_RT6A^]IOJ]<ZH_L$I+ V/)2:$:AZ ># F1.)F#,M1=R%38
PG!3#AV7U><8GJ* N$HEU ][6*GR#RD(;EVJLWVCW-"PE>!,4V N_PG:9V&+MR+R(
P_WR;6#_D):GHKTB5+&#V$^L&I:N@UT^5_*\'S4^%G7/?7Z !;0H2!-6+Z71-N))>
P].?HU*3UX342A:5DS+YNTQ5YF7.'M\(\)H);_?QKL[=HA&^ZD4O"A:R9#[<IE+I"
P2X_EYY1%C5/U<8UNO:%/P*M\+9,! (8EM96$7((W#PJ7\N<QID0 U4J4/GU5OYO=
P\G)'!#/\&O5BKCU9ZIR1 SS(^U[IY*3::?W_QZOJFU48"I(%N2PR0)8F+<KT5/5T
PZ/QL^ZTG:(NSFA<K.\*"/;)_M4,!C5-K]Z>&=;"?DNF#.VJ'V.(1B?3>&;X8'3#6
PCW0[3O2J;XF"C89J'P 'ER@%Q1M;T(+ 3##>>H6#Z#1A@$RM,.C\\0+O*I@8N8\-
P.>IMVL@V/84-D0R",=S;9;MFARIX]7M\.@]R?H/85_I4/(0NT +[6H_'@58Q4I>G
PGZME[W[K7^Y]==Z]H-_5'KD][8NC@.B_FR"I11CN8B%T6.],H@_U=JLQ9[**I<=J
PCZ>6]<X2*8BRMQ$9Y6@<RA\F6@0KQ/D'F$2GWQK9D4;84#HF(V =-.>L.8CNG%[&
P\\97)U/+N0)>\#"AQN^,UF&\>%$499/_"XT93J@/EBF[*O@^\(JLU&5![\[OI($+
P.FF 7(YTF+VL,+CIFPF-N89C=!8)SSW[060[;V53P!:H8,7&^+5O,1GH3LZLJ@SW
PZ-$9#.=P.1/FJY\/D!\S5ET<GQQX- S]RUX,"/=+$BF4PE1Y\&4#;P#%Z^&O$)^5
P3")>7F0.YUV_5OXLO&193>BJY"47FI-QBVLDNOFG!$\&@X(AOW3>=EWUIXX@F1<6
PIRY. R=N"?1#D#7#=)68P#VS]].I0$J)/5)!D2OM98176TJN\*#M7O43XOV6GG2R
P9M>:E7Y)90-?J*T\#H'7P_'_=FOW44O79"I1R\QY,47W8ZRR%/6;=;2,GM@"Q6\&
PJKPG2R5_Y$X[LW3&SS.K&DN>?5SS3<N7KU>'%<I=$J6ZWE1"O@3H:D:8HI37>#8F
PK2RR5Y%BSVS2%R,/NOXID1IHI*#"].79H, UN=$+066W2I_E0IX-09L($DGL9D9O
P87N+[X1!*0,NN%:$$MX#]XS&ASA#LHXDO6]V#Q+>DJBCR)R&M5>A=LS?@F-A)"V%
P2YIV82\,XPQRS;E.?C <+C_1OIPM<*-T6WYI'F_F8C\H'6LNZF)3 !V;?2'/ZQ* 
P :+ZX+G[Y&GVRL$K6FOGK"'<>MBGO7TL3-W$<T\#H33R>.Z8*9 JS36_-Z!S&?AO
PT+,Z&NLL]IA5XR@)*,^3YW =H4H%%3L2:<0]W)C(XP4\F:L0A+-0VMSTUR3$LYEJ
P^LWI! XU!_9_&P0[;P-9M_^4@U8[W=%#'DPV[,ML(D2+SGERZ%!:"+&L*E( ]#>"
P\G%"?>VM@Y,_6$#SH0D1M%=7>HU:JNP/&3W0S?<_>1\'L]Q%="_ ,T*7_%AK__^$
PD/#K\BUE4PH/=]L --,6AE^A>P> 4CQG$A<@&XK^6%,DRCL7B7-=&7(4O:IC5DR8
PAIVB(900W$W7-[D+@I=IYA-4P+%4,S8B%9F"5&? <Z@G-5\?W86_KK@QR&*CN&*#
PF<4N)4:-]LAK]578I]M]^B-M%K^#2H=4.-?9A-4?UJF_O\P\A+D!T5/:#B#['A5]
P$:6W,*OH4J6<X_0/W(H+AI':E)&Y-D\ZC8'@YHV53 *3"Q[+N3A#U=<)_+;1,IY"
P=NYN>P60=*,K!%G$C7!RW&%XL<6NV_I*YVK$3_?VTNB. -=/_3H9ZK7O1M$+ABZ,
P:FQLZZKI2O&"U7T^^]G:XR>+SI*JZ)2[:;=>*AS"F;[ +.2!)$0!T]*YA8EOIP!W
PGP]F*Y6#R6>W;+VU00VFI>N(_K'-ZQZ<+A1>.UL+(>0:"@L1LBIPLE7>\A2?#AK+
PQ#(1IDGC%G*!V7\9D>Z")&_'1&SO06F^@<0,%)YJ&$+:*L F?-EU.R_;F/&ABK86
PST+))9;@;H+$&<(#C'!EM ^H^H4J5U3,(L"XHZSHD@@_W45+=Y4.68(2&O:\G ]*
P=[9>[)Q:&)N6E*>",^XJ.Z6%K!G;;8?]H2'/95N-UGYTT?KBE',&Z >MY&*%!Z_B
P9NQYOD-_/US2F&;A4>$;*?['T1C!!@1=B!@G2E<0>O/?.<[HZLA8AB5)!-^^AC\5
PV6_;$/W1=(3@PJ"+XPUJ4C7";ST1^-$5Q4OE!9;!&&K>E[AS.TCT[W7O5R]I&7&%
POHFC1.03K2JAHUBS5 %]6V6'H^7.5!R/IS3VG,:RX$%BG]*GOPM7O1_^A26K6Y6,
P/Q;N<$9X46%8.>M:ZZLN4^Y;25SDA-",\5PH(?B@?;PMV\)IP%"X)AS?*0N6J&G1
P=H2K12%7\L\JGKI@72P2'#[R?W'>M:*MYXZW 4*.L'TDRYD;0M?E>ASQJ<1&=Y?T
PVRV];_AXN="5V,\7A(&%^)-*_$(M-#7QZ:9F" ]87FQ-P1T+=-G3.SRO34KL]'!8
P1>AP(Z8"/^E%3/WO6XV263C>[,-?T#=/J4);)#+'IY70YU2W#Z<G\#>>BX6GF'#6
P;#(:-^R*Q4M60X9EW]O.AKRB201[X4F<E)5$?>8?$8@A+*02##8U>;"HKS*WCG$:
PW)EO#ZZ*?"=&$9M-9/LR0Q*Q<A$_&\-R)5[:EG7N[-MP2:Y/B7@I'7:[]FH# SAZ
PXR0S8ET$-?(FF1E.6"2Z/5Q6W(2RRA6)LC1XYN??KU]##PRL,,R!3U#90H_?O;QS
P;Q0Y!\36? >NY-IP:5+ K_AYL6AO;/^B:J @9#B)DLC9<)%#P!:)CGHR&7=0NG4^
P7&3,.7_X2$TXU6<8&U*/M+3/:CEW )RQZR=GT@OC@2J+ENF4P@\.!W8)7W\^=+_A
P42'OP9YY*@ C]/,Z%'\#$\43D_C*<D3:NS-KX6,>I^UJL.N!.?^XNNP<:5W '--K
PM>W#CJ00]Q*EA,<A"E:=!7S"1S<M.5:XCQ36 WFHAO/A3"=> <0.)WQ18?Y][IT_
P.\ Y1)6:SG1$R%7R&FZK!)DQ>G[E$BBHD'[X##P7[6B2,L7BU'.87(2KUR+$S_7>
P@T*FF@W93R<7X"3V%4Z,\5&P8.:<VR $!2^WYK[RX(9T=CST?LG]A:L_NDGUP7#7
P^_QGG\>H?%Z_)_SDS\*6G!C9NYR-8X_[^)=@3_^&1JRZ8KDI@!'^1>B>EZ?WI<A&
PS0LT,#*=S'3+SO?#(0]35E@6@^-@C,DWM/L'RE'/IEP:_@D$&)_+D!4!RZ<D$/$^
P=Z;.S]>LK,,0Y,)&B4S5DU/HHDRX;> 5W=1?*)%FRB4\G_Z<)/I20Z6-/;RG!+1'
P&\$?&U23_8-4_WOPL%**XI''4T$D\<-29+; KY&M/AURVU?4ZI/7R"%:N+O978QO
P'S,H]-*M0_'81(C5NZ=I5VZ_*XIOU8LMIAUU'TM-@@QBE+<UF>EST0H55HOU3^W>
P)6V,K%(8"[BOI/(H+/D=2U#^TM9B9)IS6S_X%VG<T'H0+\6F!2I=\I]A5\2T9R(8
P< >0,AM=DK*INYC4936OBY?M+>4ZA8IVK#8G<V-#=3P]R+0!H8"[@2JN#D_@=0KT
P>BL^+F0?5DVP!6M2M^0:)U#CL=,J ^9AWC2'6]YM@)1TRLIOOIU?>T1XI)[;E#?#
PP.0_P;MC3O,)@58Z@RMN0*?<>L!-?QL:.#6+ U8*-\*8E)+1\3-;%S</QY_#^G* 
P.712//1ZHS](G!C#5ZF";QP^L-"7ZCY'">4C[H>]^]U1C2PBPX2V?0MC6HAHSK)'
P-3;O%+T&9U\LN\1JD!?5B^%R]>J$G<SNSH F4A2^Z4!A,"5X2$ _\"#Q\4AS.5;#
P]_\+K5=&(STCY5CN);.#T^V:RV,S1 ;HTE_IEG\AV_Z*SQ-WR1K92S\-G9*MU4!D
PKHX8MT..Q:*$/EL^CN).:?=QJ] _!RX<J6^^'CTE+F@&O@W)4.=D;KKU+%!BU*,=
PDC!-A QT0QA5>)%J,'@C88-N1PD+<<<-AUTP"7F=&+$L/?-R&&37-Q$F?$KOMB;K
P3X$Q-QKA;<]N:I,1P[O>5".GA\/C=3Z,1$^E#.?07=^):3TRO]L@&$0:6XN$=O'N
P;?Q>U(\_0NWVI?@9%E:,SSFF1-CI6*?D@Y,#('0 A4LA5,%S^@*F T"-53,L@CJL
P-J7T#"9U-<)Z%U&KCEEGTUAXR %*'']RO"K"OY%5F)6/89,H6'Q'4I8-*98I]:-K
PG; O)=S#J$ALQ]\>]\=G IY&^WJ9D, I:I>L87%,#N[I5]P\L'?:=4GY55PQ .$,
PKEP3FK^N>8UP6-W?(K AOPYK@2/? $TGR!&I47?H^C]RO@I)D!Y9W[<A8X046ZM9
P>A]IB!K&IGBO*_# 2"4/C#V?X-4H81%.^8W/4W- ^5BO)[OP/SY5V_<=(9RG]'(C
P4J'V$@G0L/J%]=>.7!D>(LIX ;S4'^&T!R347E+G:P>% ]*< B16DO04Y!R7,F4/
PRD9E,E]]67&-)FX%+4J0HVWDA!W0^1EZ0]L=6(^*G#3HIV:T*27ISHI0- 4%6JG#
P\LJ@R8"RY407 2[+FV)E=H60!8LGWR$?+)?21X#:@M;IYU,,?AWF3Z+VA8]H>C(.
P=^>;EH+3MY.")+HO4GCW$ EU]9+H*\9TE.7DD=NK[#.X%!NM9&_*])@N&1T%>X#Z
PK66W#KQ7 A-*^MBOE5N%DM<J*MJ))X9)@#<4B<_MM!+L&DA,SO^Z'/$;M+IUV<EW
PT8NV,1JY/+Z)W,8M:U-W&,7RJ^0JZSL'4YUP.%[*&396#5Y<9DO&_4T5F3,'7^O8
P:V^<.XG8G4:,O*+2H7CCL$(!(#RF)Y]10,Q3=F)BLOU0LBN.1C*FF-*K?\*3!T*:
P?E$HQ9G_@V<=J27FN?"6) /0.@?SDD$;, 5X4&1L)5N;U*&<:"^OL$9LS]*SD4AE
PZS+(0(+J&QZ!VB\KG)2[3V-^P>NJ5WR[E_%3]]"5CXSRU#NVK&G?6LH>X14ME9"M
P(SK<K 3-@7Y-_6VAGT#CGD1"<I#__&.+;@D^\;?B(J'8H(CEY@>\I)G<_TOO$/+@
P^<F['?:8?J*GE./AN9[/WKQH):\.5UQ,#*(EHG9U C:)? -$9ZNC*R!;9/4"&;3(
PVFV^(-?!(#HPC0=&CWA-^.PT_V)R$[X ,RRA%(*@P9%TC1.!.2Y4#%ZW0U>?Y[MW
P[@DF+!4DY0!89Q_G4)^,PTJ6"CB$Y6"1$EPM#>-)*QHTF;R#%MS5AM"*0AZ(SKB#
PD=]R5V>A.TI<9ELUX T!@IMF_[]O<]CR\S5O\4$Z88J^51'T-%P^)/+-DYK'#<^>
P7X=S")@J6E'S@.&#.,&\%G%((ID<T=*8U<T1"U-29AW9C6O6$ L;3+L!I6&N@OB<
P A2\=F,T[;T-./GI!7>LQ9&,JS-A,<HQ,/V)LF]W;C3XZM]-J=Y%H?B,O)BEI2GK
P'$BXH_!?V.110J_1B6\KZ7E%NQ>41[A/K["72^[(-$]0*QJY53'=VT?G333!IB;S
P[!6 C KIE&?XW219 ;4K%9YD[O!P<C1!&J/C"MK>1NMEM1GHRPC^7VVCOX5*Z..A
P67BB(;)Y7 F@!YR(+6'@@@A8-$VHBN11"F!2;F[RI+_I6HWQ]@&,]VUP&PF?4QY!
P9<YQ;AF\^ ,5HC%(V7K2];&!M_)=*O,(@I[0:[$0<D$)6FN;$1H*P*JBF8S:X;'Z
PHS<EM_71R_SC?%S699V:LGO=B=6EJ@747;VV">+)E3\RRK#IWZ"N!=)1N'2UO9?U
P5PNUBQ3 Z]D<;79^$4-;[G/[P8_)F9CK=K<-0%&ANL$Z)FF<3CCAC &[)OJ8S]P.
P=IR%I\W"]?Q&G*2$9+7@*59@C85\I]5?8M^I!&<B>S#>=.;+\'*!4E-U11C7U2),
P]T[7^PW.]AW[L;?4$;_ZY5_OD,/>U3P+)CES;FM+M#U4=FP[_EW1@-'<K5J\[B_X
P6.[;'/\#HM*_>_H[27DN,55YK(>_27:#D$F@3)XZ6-OXXIN ;2:-YO]K\NUKCY(@
PRE8R;&SA<OJ0]VPPBLOQB<B6F0Z<Z3]BRF)J<V,0/332-:*9LI;O & KR,B>IZY,
PT^-OP(/+J"_69.]>E*Z_PAFQX$.L"H3I$8E0\EHK5ZT"V8?'#: RZ7XU$8 QZ1Q@
P)J!^DE'F2@;=9T)]*&,H4Q8?&%M<.''+3ZT]Z44P4[KT@R434ZV+RPX*]'SC=%AK
P&9OO7T8@6_A9,TPU(X =VCAVP :(]VA=0FZ]P!&B2?6IF'L8VNZ@:MZJ^?]'*)_5
PDVCO6_YTVVHM+L=2<(@0"E;GPG6X/SC]A;QD+(5Q,P=RM(+!K,PH:23QGO-1-=9T
P#&Z*3:TLMWN7P1(G;N[Y74T4^^U:K. @<7HM%I.DW+VYAM^O_1B^?%RG2Z]-0?9L
P0@+^K'@_E40L\0KE1\&JT2CWOQ9:#<FO\87;>)35%5&9X:G'<-N(D\!9/RNMMWVZ
P/A6!2L\6^/L2B_LT#["$ :[#K75MYZ.KX]%]0+YR!XH!YMG.N9%X_E%6,!,O?/?K
PU:(3V,"T92BMYA[?0WX<$4_#DK2'$(Z6CDCMGCXDK2GHTO_^WG/)M7E(XM-/P(/U
P[+0* 26;3'T=HF>.]]P::,8LI E#'KJ/*HUH,JT$/1&"#S-CWNKF''S,4!U9BSH^
P2-\8F&59V?6D=F/4IJ)&130X&4JR9#LUA9ST6EHX+! -,,T%K9%8BE@&/E8PG*KJ
PUD6RA2LOV& N+4;^:QI,?%6B3LD$L[ "F*U2C.(':XRZ=:@7I6=$LG _'ZJ:G'.H
P463RBR'!!H)HY2.,,>N^1PD^V2CIUW?$N\J]\<1$I@B'RZ@>2ORXBL[8.8-/I:E!
PO1GF&@SV]7?I(W+A_AYVABVSI0L_A( GL&DV)-OWPI:Q/73<;5-2RHAD<#XO'>&T
P<,3RDZ5YR<\X;9824YH&Z4CE B<EI4I"#(]UH0XFH(N$F=BMYKJ)[6?IWB.\9+:Y
P(7=4?#_9^7EB$WI$;X<FUJVB-C.>QR]8)DX:.RI<Q1I\)];PT?G;+J!Z!R66WWYA
PX&0C0$,/]5B+Q/WX1(\1*>ID5!DX\V*F8=O/S'7;^#WP8B5JH"2HKIV"'?"8CQ^U
P/85G-9?C^PAY49;NU?/Q-#N!-._^W7C"W!I;,#,Q1H"YKLH8"SS&I!B&:G1&/5-/
PF>CF0CI0O \JN_8N<\AB+)0K?\6YT3?>I\[:N89<??CK^DY<;87ZSS[Y7JL'TPW'
P7/^8\I_S;[D^9%R>)IM*++!66QHGUU_.*]92)F$C(86!PYWU9;FSH#LI!0GEPU>(
P/CB3ID.+XM. [SZ74HUFF^(RAPZ:T712M:WD V&BKN32JM+_/F7OP&5AMRU9G^O0
P@+99@^;<LF/)K'RVHF.#,1O WD3FLO_C&=K^,)27MM%&[K?QAJ7JT=OSYS.-(WDG
PB.=K:Z@4(9%O)DP0^U'*.)@'20[[YLQ'S2L()#YIXV@-_KV,YE<]QD.);V:O\[&3
P7Y+-1?.ADKQ440;"#Y]O?@5/T[L$:8@B"4".3 %/8B%P.ZLK3EAIY+@\.^48*6'5
P!2F>7!G1S-D15[!QJ^/V_P^)LT5O@><#_",6WW1]=.;(8\>IKXH!S<M'33!QR@?1
P "'N'67,P!"'Q@3Y_P>ZH"EN!T >\6L,")Z\R!H4D-A+-##[&ZQI"Z_=8H=^3@9;
P%8!EY)<= \NL?4DWY4[EEN6N6@-MLD3S\,;7Y/P(5 63\P!H?.23:N>B"VKJ8W:*
P!]00GY^*_@(,2Z:<N)R&<'XFXXX'1"S?^&X*U"M#2VIBG#>!93V'+:4 0CV>0P_?
PK;H6%*DXY<VSL;!\K-1;8Y$ /TH+A[6B M3U>!&(T9;[T_*39"F<:)$Y>P+6/M!+
P5Z%.ISO8CD28A?$!K[S"RV(4.*]A[ 8W*_%@4#/&>%RY@NGHJI;US7#O] X(!()=
P43 &")]<"_R&ZK,QE?1K4!O?[:DO'A$L$RFO COR#E,LBJXC':WMFA*YX@MMKMIS
P/I]+WS[*R[6J'BW\2&PA?HO&W^FLBOZP] *FX!R="5AK%&:TVN;??<TA^_+<><Z"
P!%(WV/0AJKQ$S+GA<8A1.<N@Z]?^.$88]G48&)KK(GF/', :T<:N^6Q@AA:4FZA0
P/Q'+#Q[FIY;<3T> K",.QJ0%RJ_T0<087P.-\3<Z^ )\XX@)OD\TJ).?V0,#HYI"
P$K'T^*$B/_JU'0[W1M)1U/ @8-1'%%5F4J"A\1>S/PKT.PRA?'#UY0HWW25Q&&;2
P:8QF(O S$KD*DR].'2^QTLBQV@B2_6M0+NVEQ=2A,NH #^+!TN"C/RS$#K"KOU1O
P9J=D&0D6,3OS%\+JJ#<,EZML@[Y%L;69B^^.=$:##+CCX#2#W[>+4%[A\'I__@#&
P79!)IK08L9";DN>E8/NR;$SGC-6O=@91:M!O=W)!U"T-X!-77=N<\Z:6$2:4T%_!
P%+Y('!&"4_1%'JZ%%B4JWD$^([NIS+EZ+1+_BC"R7D)LC>P-*\4(^_ =F["@VCK)
P9\K02F$=0T.P'1[YIQN?38'=) %BD:L$0SDMKH$3R*>.9(T9=_0RD\^G/]_=*MNJ
PO&5X2];.FC+EQRR2?XF53TM\$W6&R*R%8YW6!*K7Q!/S*.TMRB3.&4YPM&^8+Y+M
P-")N6?L\7 %:(!A5(7OFTP2<XY7P]T+Q0WPUB059X?-GYY,$LU+ <$]U;K"KZBG!
P2-?T.9P[B4@K8O->+U@9E''WRZKMK\[?LX%RC.DJ7V@(",4'$"JFVEV%!ZL!SJ?:
PF29'-UMD?:V&&5=4)QV6H@T95^W6[RL]($5U#+C]"U+U6/ ,M(GNJHNZ!O"H"4^E
P.Y'["[K:R?75E;&'2%PU#JQ6-PMX=#)5WG=R%EQH15KLDYO\!X.H.F^[_H_+;('3
P5 "$U=I0F%%[^Z7-:VZ>5-=([J*JIFI2P=P4AA>K\!SNO"1E.0J?:%-74YI>N#EY
P'J)EKAW-4#G&O4'NB5[IH8!SU^VB7^;9M9%Z7-/CT]V^5; /XBFULD1T/$$ZWP39
P+UO7KZ>\K_0:>,3WD<@8[Y/[AJBMT7_UIDP+<Y^>5G8)"B+9Y&+;U=,OR#S&A'.S
PX;&)IT*8[5A&(0N'2?YDUWX+D(=,E0LM(BH9XQ7W468:;S9WLSD$AH)I@(?57EOI
P:$DPE>=53\0H2O09H$.B#Y>?5!O *0\@M3/39'R+:L7QZ+/FT;B*?%\4M]NZH+'H
PF1MDVBLU84N>AD\YY5.WA//GEEL0\:SF#\:>URD[^O/D.ZUPY@TJ>B5-)!XMSO23
P2I&7[ ^'5.F8AQR<.<Y:;8\!5 Z07_4AC'DO=2@V0=%3(UW5D:T=ND]\+5/2SN2X
P 6?QSFHXCU-$D=R^=PT*%JC=A9SV8&UT>Y[2IUN1N[C.?__DS, M2QD$K2]RX2-(
P8U/:^+U _U!9/E0WNHL>O+;FFV-5^@=E;3/U.\>%178KQ((B7@A.[:'0&!@]'"1D
P]#5HJ0K(307(Z W]O_.@<01/ 'N>==QMT"$*F2E@T*^Q2S^BK77O6AM&ZB-;W>&[
PF7WRDJ8O'N@*U\$3TC.-M+&..,K+IC@'EW/HN(/A34%4!'<\E*&D>Z"_7!06'9Y+
PF,CCYSYGO)FXR8&GV[AD(O%^ +S)I!LX-<[&MUY>Q YS'@6XQQMB&(?=C2>//MUF
P@+!04Z]HG-]D'\S[9OG+.["'T / 3,R6TF<62NNZ-L=_4#]5Z:5'C A%Z=V9$('X
PPLU5!$TK>T2^EO%D2>P<:-&7^<^9?:]5#R$>G;7!M<=P5CCUF"#O_]0NQ&,<U-.3
PJ!BY:O4<;GBN9L@J@5BS-NA4BYZIT)@/N00.XX63MP=.Y=F*)%<I"@*4>T=/@1= 
P+.VUBYF>7K,385__;8DEFZ<430DJL[=PTB <K>.5*G][R\QSW=6VN5H?'T)B3=5K
P-Q!#DA=[ &W2$0&23FWCJ2_0A>KDI6OAB-Q'_"H<]Y,K=N:$I*54 [5L8T<;PYWF
P_/H6M%PO*$:Q^%[0W+ H"[QKL)K2ODR0M$.KJ:WT@T-=2;-L]G<O,'MOWKZ:'^G8
P:LZ5=-M26_FL1X I!VH918S'MJ@6(<I4MO'VD>;]FY(K\QUH#56R8:]376,[0J3S
P@Q-O;,&:0-#9D!TJ,I0L /\7S:X[D$32C D5Q%MR;T-4'AD"(BR.E>P>MS-F QJ,
P6,P<:D<K5J\JJV5?J3LF/O^J(B-FZN1KT*LN XF0(3PR$D4Y[[=!;);4RH!!FN&V
P^]3,=GA*'?@HNSB65DP['L.X5/(A_+-;IZ#/GJ*&/Z8@:@K(S*#K;X6;@LK@[FG&
P?LM8E?Q-U@TJ"'Y_ #R]C3:UVBB0\<?BE-O@H[Y=!0R,1:M1A'??[SC5J7#GP.;8
P#04++6U7*CHE<6*V5:"I6]63LN-UESFU\9XBM*>6.R"F*G5E2"P//$5F0NR-A6JB
P9[%AM))P_>"%1AS60W4)-^W#.):^DY;R,/B/.Y)G;Q:>DE4%QB1S1GSJ[]OU0XBR
PPDHTZPQR/R)B\:C(&ZH?5#'2Q!U167N\413W9UH'T#:H$!'3W:!IT" %LBR:^YT>
P-[(K ^.,07@U/1$%Q8O,1O1ALX?2=,<JDR(J66 XJZ, H+W9KU)*?'=7O>PT581]
PMXE"EF$'BUPARIKY)?))('5[EPJIRGE<O'$%LJ**=)Q-+EFUX(/&&E!@9@'*9&6Q
PW[0F>VA(C;FS7U1H!+C.?JUL..AR@2#D\1A0X"Y%A=H^K[M(@9V1^BQH0"0=#S8R
PLEJ)L,#LJO 3B=-ZO_K_UZY,CG'EXE1%Z1*<%J_CF90P\QT0*9DM>U&4D5RQ.QO#
P_5O\3FE#*I1?5>5=R]V$I/7?5&X# NJ9IG[QY/>27PCF.9/-J(^!#7E(R6YV27R4
PJ#C0M"5%A"LS)ZLG7XH[2L1!3>(C%W;]SQY[! /I8@&WY8;[?;XBI6SU=!^;\2'G
P]YH)=3C%"UIU[8M4[XH!(G[W+/+YCX[$>DW:(3YNH$FCRI:7U>!%HC1>O*Z H3,W
P-J[MGCGIS>.;8]JA'KQ/TKHA1QL#HIM#_Y5=WI]TY;_DM+>C2C9@E#>2H35'U#V5
P-LO%\3W-Y9+]71;A[@087>N3ESQ@WF$'/([[_RK48Y9/ZF#%FU-59H<2?C\NS.YM
P_G+6B+R$/B0@Q!J%"(PFFTEEUF,Q?7HP%K7#%,ZH)Y1&?)%QNX^M0K@X1<QW<Y9E
PDXVI,)X!,9L0E9(E>YSI/%I79UFH-+RD$I06#=R8Y@@\69SW)K9M2(N@HV?B$]L7
P7VN1&RHC>6TG]PEV^.<*2\#[GW@BGDGI%M'UE$?V_2K?(F[<JFJ\)8RT.OOSF?^_
P),D2,F!R:CVF5/]9C\ 66%/O5>FN:&,? >EQ8R!D,YS)^.+;\BT>@7L+];*P\9#E
P"U<W.5SVA?7MAY[-83G51]Q_AOUSP<V-0\;ILSZ^3==W5;/M#=.(&/W&R(5)R+T3
P?DK(43,6".#I;^;[]DDCLJZ:!N:5CH<./P@JLI9WT5W<*!323A5F4+O;B(CU<4NH
PFWT)!2C5&)G9,TBES_/4O6$I9JZ!*##ND"'K7.'NR%+8VC,Q2RQT:NXX!$1OTT27
P^XO:D;.)&!Q6CDOHKD+!H+R <W#? 5.T''LUD^!TQN@[9OF<3K3HR&_FTQ6-+U!+
PL<6F>U )-H5O]Q-M.E#5<BG0Y?+S-U+D^[)!,-HP.>\R8&NTU?"(PL-.?\C'B,03
PJ>P2.D<=?UN:MT4C7K)N?_3=7F2\@MMM1+2S(1IPKL[L=_2.<.].7:3UT(?-^3^8
P'V-5?]24.V 2$[G-@'2"L[&9SQ>/DI.3IJ5\C$)@1S)89X4IC=$Y^LKS;=N$ UC/
P2(# >L0RF.XAF39^A7S6E%1&S9'W16DCI^@@,O80TA=T.D3X&U>)+MDO[YE@]-P*
PQY?+7A3HQ@A?#Q?EP[)VEYGS+15+:6).\&+4@^1IFEPZAUOEV;5[8PD6)H4ZZND4
PM3D@8%W2,%]#./Z#]@Y*U.A)#44S*%:I#X2;K5+H(DS^#,:@?9,'2QIT[0?M1P&!
PR3PH%:]MX*2>@R^2P\56.KYGKY.9JFOW"6)- <+=4#[1 \O:[]/4:9!?O!ZL7ZUZ
PZ.)+^C, Q711MZ>V0QTC^[-%B<[.1W9+,3H^;N?NER[[J(SD' 3:%Z.E?>&\O7TI
PI[;&T(F\Q(2?8U$85>SIR#QD8CF!H1YH5B.<VE2S9('>2A&J/A&="T,%6+HJX+D*
P"6,IU4=/^ P&C4$I18(7G6,:3^ 2DG S;Q+ZXEK-,>1)'.+GJ%-GE@1+I6_](6.F
P&: [HR++1P&<G'6:,DH"&@OB>UO)*3G+*Q*FS)/X\:EZHOOWBETRTNIU,5DM^D$O
P:D]HG1$E#HFUY2..,A2,>>4)8((9DE[L64O26HAM8S!D(J779P7$2 >-N]'O9GRV
PI!"-=SJ8MBFLFKQR%=]*\;$=^W@51KI%>1Q&4A*$SKD+0UN87V^OOE4?U$8&#T+D
PO\=&#),7TF^+%ZJ5;O%50@:<8"75.RJ(H+/6&@2YRJBXC25(9N$R6F$!E[!KS^+D
P6Y@"P7)JSQ4W6D.5#,)_!07N&A]?_/V%CX&>K%4K[W>)+A3R7\F$]8E)9XP=5@R9
P'LD1;"^#/ (E-<E_4.+I8H?Y8.<73V[/)GGKAQ]!WJ%9I:KAVQRV-/5FVZ%J,OTP
P3;0>A!_4<W7T5#J-\^'KL!+W_X:T.0</38;9\"/('9$!JG6X[1$WG5S%K;F)#'BP
P%9KM!/_LAHGM-T%T?(&0<J43ORD7IV[J-CN=$EKEPHXJGD$;X4ED:$ WMO<"D%U!
P*\AC^AAYL(9= !=5.E&4A-* P ONO.X8W2+0B)C46#"94X0E\U\)SAP2 M0/S Q?
P M(%XWI]6/X^%#+&MVY+UW^Q*E5^K>MPQE'8R+(B:"G:=4'1R%>NE7%(*=&>%Y%B
P]JA4&!4E#'_TZ3&%_M9P0FD("3*ZEH'IAGMM;>=AE=_J&P+.G*V#5T%]"PUV>,)P
POQ!J,4Q?18>OH:_#\>UXKY(I4+(D\CZ^#D0&.9RX<N=)-LI$D)E,X%!-9V.P7G8E
P*1?*>G,X]'D6JM"LGS':_9%61$'\[ORB'OQ#(+)@L^N",YN>8NI4<B/L?URA@4/4
P>, /O^)W&P1[J@T_'G[],\)+CRCRLVFJWUS+A8KCI)NFPZ-*W+2]F=2!D'ABU5CH
P8+52>;>? JE1!JB-%1U-V 0)KO,R$H0O/X@4OKE-CDL;FNW8LHSJ>[B.6F(=[BCY
PZ6QY AJG9#U0_W-I'@GXI_7'CEE[WAE!)$(G9$Z<EH,NF.:Y4F(?U-$+#$\_U(V&
P4TUY';.@J^*-$=N(*UJ$#5Z .L5*G=&J!D'HP=FB+>IG"2ARC$)\+7!,AR?)W>MN
PE3^C^M*90K3O<&WSWID'N=X](Z6$05I:KW_A7IAK>LX$W^OCZ@$SR$68&&Y'64P2
P$Z!\V&G5ZBR9!>07+J$!^R&4#LM?Q9.+<9B)U](:I-M_-!E_)>=VWKKUQ5Y&PQ<4
P2#Z3._PY)4_\#&D:9HX0)?!R2C1;UU&V>QZN-25X:RUI&YY:!M9/*:3B&%A*FE]S
P1#D\ZY[R@GII]U@2E:MQM QX[0%^B9'")KF-2R9ML]"RQ^-.3WK)5W@^=[JAZ\-;
P%K'V4D)RV6N5(XUU&L8%0AD@(7OCU?8GX,8WJ$+$$<IA4SUHY./I[(QZT\]^F:G5
PN^C_K22R5B&\-7>4\BJK)T(78Q[)VK6N8>D]#'"W4^Z>W%TSN6]57)1@E/0ZRF 5
PVVBT]*&\8=GT:#=RO_VXFZIMQ$CP,\59,689'*_O?0Z[=35U(]V#[S<,UHL2BX<=
P14(]K"VG2WYR3-?7_"X&EK'?]> 7\_O$7 9(Q^CLJD,V*GW&/?_S+PHS]37]-XH&
P:BL<DE@\C"59Q?.,#+%&GJD4P!)\Z]#L62*ICE[%%<AE<1U&8F4^BDLA$X\39(_M
PH '9^$7,.04GZ^8XN-BT6HYZ06$IP?  !7-^8GT2*/:EF^,9Q&DW<-^(EVV+BG30
P0('NEUUY,$:L,\@.6I_'*FS/5/Q'%TD +(2ILWH$'9C7,&X>:!]SD>I$YVUHY)2>
P&FGJC\:/2:B*3O7-&$71*M\@BZ ,OYW,PPLEP98Q:[W:G9]^JF9Y3K@>U-$^E';T
P /-O$S/WGM7.=_*9"7<9-P\938"V$,R[%=8FFVY^2EL0'>QWE6T"$+1P.-%9]#B"
P1=/LQB FISR'T0E,32$)/A0J;Y>*B+T=;"8C<K@U*3 HR QKVL=WJ&9;7CB3P/J=
P>>,Y@#NF5(%";.0.POZCT%L5+1WWV^G=Z()7C(,0]]>&I[UZB&:8I,(G--5-T/.S
PA<SB-UL6WFTO#3*ZN1&NHV5=VD@?58/9\=M U2OK^UF>T#^=9%L3&WN)]VC\OZR!
P3:Y1QF]0>6^4 ?*Q>V>EUZ53)?5OH2&@5M-WT3,^TMMS_T"LPCRQ;?W]8$1N9<VM
P[1BE#M'1ORA[3/>M9= F,KY O'W8 $!$LDL#SY,U1?M;@0%%I)U<X?2TO>GSF"@/
P'N,3V^CYMYXG<@A?"9X-<T=;^*^<-U YW#,Q>-3_;F)$=B#M C-1?A;ILYNXF5;V
PGOA1>%",2Q6HEWLAZA2N:M\G)1=B8HJAYAT%5"4L0N<DN>PB:RB![-H!!$K+NY!S
P8P4JJ)NM14?OZ:I7;,RI!WMZV!?\>UR&TS8R0#W*C_51F2_J5H9\ES<"UI;Z -M"
P?!W;H],-R-+CH922)(ZJZA+5_5^%40F)'(Z/ 56D52)5@/1@8"50H9"\@?D&Q>L*
P/%0N,?"T3;&Z!]%X )"R__E6:+_KDOKOD=-[<P17RH\A-WBPOVXL6]L->\%&;D66
P70Y;QYMY)#1:7GC%:C$9!T$7)J;<Z?"5E^4TC"A]XSYF?[,0.A_Q'>\_RV4":#OI
PSVK\/>78"5YYS+]^>;*@)<[JRPG8)==&&YMO/<<-> =,2@T]!%+A@+\9C"M:=X5W
P*8UM3Z(S5*0GLFE-/Z\NZ25\*[KITSF^3*1SS'JKN27V@D8YS6.V\'"29X::055Y
P6.P<%55=,-8<LUM6?KP5RD30+9!)W(4_$?NV40T5338],)L+<(/ITMHTO9AKFU@/
P133.F&,6LM<SF;I'#V&#YM-3SW8H,-?848EV6M"6M_&<)07C%6&>I'Q-'&_?D; H
P)&EJB<7VO*%>G6;C)J:(0FDH<C,+X.<\'1KMM^,51OL0CB]Y:DS@3 B\?XLU/-/<
PV)RX.#%QX;+)M7,I><G-4-Q87U;XVO%/G4>0@4"T_T6.Q;6^*R&2H0.1SIE/?X/@
P)FKW1^J1N#$# 3XMLWJ<GWF1:T][EE(@>V4Y-G17[C$&%^$%1\1>U4E2U;I/^ZT[
P[O.RR#@H8:LP7>['%S0[+VD@]SA;_Q: 9 ^:;>8A?6%IEU$XN*0LQ)"VC(>YGVLX
PF_2CE6\O\& .CR7W-3AR)+5%.Y5*L+PB;H,U6??VOQT'DX9>[.(_8'-A58_MBX6B
PWM&1<@YJK0S,P]8!U]4JG]OZ63IRH=]_EHP(W@]%,+(\@J:GYWGZ?N.!_6R[EKC)
PDW?ARJE\OM_?O%V+]NU14X_@@BRF7V3U%04$[".B[=&(X"M)J!RA3!:6L]*H(PDI
PZSAEQ9+)+T .G];MJ^@F?LFM.28+.^>#X?)?% K".^V;FC4S8N7M0&=[$ZG7,KEX
PFZ@L">]YHAE] YDYZ=A?#0YH')>).':]A[RXV/^ I-TS40SXA22SL.SC%N'*@"1#
P.0"Q-8J5P7]"XJ4V'!I[P^76_-4<TFW/M%=YUL^4Q3[B.H\<DY[EH(<F]H+OJ&1#
PB">K"$"6'<OP8&)QC%2Q=LP+,4]-QO-)476O+2>RFB7J1A'1<MBY*\*[)GYY$-',
PFQ!"#;1;KGA\B3Y,^OB4@!M'@.MG4A3()FJK)I++,/4)VG 99-D: 6+UF )57V^;
P6GD5[D'!4/;":<B))YB]R[%JBR'1!%@,13#9R#')70/!78"+IMHVB%-%-^R>ND;,
P\D0WWSM\#A<&&N91AEK7-HLQZ]SQ?<7>%LX>?O(9A7^SIJ$;88[X5 1YU!CR=(T2
P'?GX+0$8 N?22O"SI+0IJ+YB/\O6N'P%>288N;&RNHJMM:)F3B+;_2'M L8(;S\'
PA5=W]Y#%-PW1/$N_[D-&T:FAREH+E5NNED>=9.!V7F!S?66343$)Z(#POH("9.]E
P! *MAL+P/5\U4"+%:LYMTRB#)LCPIFE_=FQ@"NV>OQPIH=K9N""008" F25:@9KP
PVJ%UJ\)'B/59B(6,:%,_2*F@3 <M('#9!\"N+@\-P[4Q2./Y(>AF\TUQ4I=FP,IN
P8XN\9IYEK?=3RTIH9K]$M6RW[&V:9AUCJU""-5(31XY/SA/,';R,]VS7J:T8;0VI
PJ>!H$.'5.$7-FT7 #7A'CU )M4E >I/^BX,J>K=W5VYN/3<S.YU/CA1449HFOZ^_
PR0^U.9I*@U\W+C9#YWI7)1(;1PR_ [MWDCB%8N5'-=^^6/!%".AH0?1)2CXB4#[C
PXOCY#M=3;B784W]2[>_QLT!*S+7O69,*=2+OE10]3$V-1JXZ+667.?>45X9___R*
PE$ 1*KQ)=0(ZJ *>UJQXMY@KUK<D(SHR=41L?R8$$'0=8<NE\(WA%OC&FF4$)% B
P?L,W7S\&$DTXE0A3B@'EYN.#Y<NV4:D+G.%D&1%/R'(KN6M2.*MTN>JS%]&E'->"
PQACER"P[NLOG!U!/ ?R#9I,?'TS ]GYI<^-+0'.D\[:19?++.P/%/?-1@O&"(@XM
P20O- \D^[)-(7X /%F; =,U( 6;YZ:U,WXY)C!1^F8=GM9H6I!F!"LP3.Y)FN"1A
P55O)..S;;H$ R."5H+;9W]DFU;?I=XX@K'A)V7U-/"80)KX/5I*LY4\-GPE[>9ZI
P\Q?O]:%(X.HS%D X^;R;">_SM'DY[H+N_97TIT"]K7Z% 3,BU4P*,@=ORG*1(U7_
P^JNK.K.F )4&E?7!0;@(-3RP6)CPX]M(C>F67B5\)P]0FL1^WI]9@*GYJW_.A,DR
P LC=M8!]U(?[,JS=VNI$3LY1(V)G[;V'/F7!K&J(62BVJ8QRW,N-("<PABH.7<+U
P.<,=GSI <_MBVO:'F36/5]_K%-Q"BBN-\5K9Q("/APY1PKS^3N6K>X=0_\G/)SMF
P!M#.IOR5^*RQKK2M'@TN()<X?<0PP%S+B-KEQEM'XAS&.E@ZT1D'^7O70ZOFJSVE
P"==CY7^0;$)-M>J&VA'-*%G9MP[@Z3&L^=4Q=@NP*=2PGDRJE <RS%=74(%PEN)1
PY.!%N%5\F<^,82SZM Y*?>M%'BSXFAS8  [C0/83N4<!\8_O5_7!"#F82FCIW36J
PTC>>C(W5)'<Z@AW:M_MXJTE(P'&8IT\@:,"K&%@ *0Z.2LV9OE4Y"D'R9\PUG(/,
P-;/*TA%(47CS4IC&LH:MT9'809@%Q/5?>S$RNNY9986RE*YCNM.8^/+?R$0N<Y]%
P>B/_C:Y(ME0OY'B?HXM/7W?,>%XH?2D>85*AU%T;!(MV;9  W_&G% IF9$3(7:,J
P!4$=\Y.JZJC;-%-5?.1*#GUOC3O@D=\VVG=7DVW7_9I_??>8CPR8^"0:@LD,<NOW
P5AM;EJL(CH:X(\HY.%[EI>U/>9UB,/$I25=59NL#0GD#E#!%$HI>@S01=][&D8K(
P1U66Y@H"35P&0=3"N6J$8 >FFL7N]Q5%#K.-7;STPY'LJS2 P;_MEGH Q+;NN>D'
P \] #A1*<.K4:''V:@O8,B%K9<?H4UO5="!:__@JB2+\7^+P]>]!X2APVVR<G+A9
PU\5*M,(R?=&,W%G6X6V?;#&7$R_-JARM.W*5:^_\=%5^/5'W<#YKC?2UIF>SN<DM
PC.3UT=WXC)ILL\_TRP)1L)Q(8U"S\,,=5)VY"'KWZ#1[0QU=,3MJPR&EM(W_38$&
PS:\F/,.K2"T:G1Q 4NWXGU%!Y+ OK080CZ\81TONTLW]JL5U(G9Y#=1L%S@EFG4T
P.&&RE6CY')".35R82&C,"HZ;-Y*B[7+-=@*_OLG!9"!<-MA'*4KFUN(5VYI67)7Q
P-KE?G%M7NT QH%Y:207ROE<1W.L\O4=&9_TAMMF@]4O-:TX0[O;J>:-E0#YEW7^U
PCJD'OHU25LP2E1SP6**(D!'U\/;DB,Z6KY:1.\-KYOBNEGF>2O#1P360LM]ZD9^!
PQ)]P4(01=*N? 6%,XM8H3M JD5!<BI*F' \1_DB!(<L[JL-9;AI\B32NI]RK>&>6
PFL]T<)1106?<H;#B:R+\DE157@D*!HNLV&WR]4\;=?Y+"0'JH)=IKJ@,FQ028_:>
P"IW^3.2B.ZJ2ZU&TW:+S&3#VPVW+C/T3DDG-$P"O8&>VF=QY1C/%;^-L_H0KP&GL
P/!JDQY]I>UI8<FL]2L[=3[?,-IO\[Q8S#5E^A2ZH__-\6JF7<NY'LI5NUC:35+B:
P^DPF)OE#O3QV2Y3*L>5FTJQ:U''P:<B+EQ)V++@G)L"FP2*<#)?_>W3KQ_!I;%++
PQU&OGLCK^[++C&0?FZA82(-G1 -(0<66_-Q?UD,*Y>!T(DQS2$XBZXEXIGB^:_0[
PA4LR25A%0C[41[TB[7:&ML*1][6MEQO,<U5[#!&A(T[MGIWPE>]]PBW@ID_1+]"7
P3<MJIW$]5'C7-K$=L#(/Q<M3$1V% ?ZS,O8\9U'.CZW2J5"$D99+^/V+2L1+<F4F
P]T:^=R:G\5K#GQF(4_?\XT>E;LDD8:&<Y/&V6%4"Z3Z;?$S?=92T#G#N6'Q:%ZN)
PTV3L7!!PW8I#L!-:J2.,; X''DTWR/U-G&O/1)56VB5M"/"C["E)RSW/G\;%]'FN
P(U-3X3U1*:_M#)9[=V;O_PNOEF>9",V8>#?,:,O(FM!(D-9ZSSC&(I_Z9*V"L-]H
PV6U)_>^COXPTPJTS-+>$%%O'3)6V)/3%KY9O93;\(+K!C^\!"L'$6QD3)$.S:SME
POB>:447HWHR:1SDUCW1LE$!E+C1%]O 8FQJI2$G@S442#0B1 (H0>3? W6)GGW;O
PCK+D]T_LQBDL5;2BDNR2+SZ;B2HIWXX0??E52D"+L>/#ZHI;_K6HNX4T^7X'F<]1
P0APZR"4+2J<MY_FV2ZV'$-L2"@EHQPUD8_I"/:1S*W-*R#%^L:S'5^C.ZO>Y0 $>
PC(Y>;X0IL70#]F_J$.NJIW!$RX)F-"NM]Y+* W_&*7"!LW#!)8N1>A" @&W(N/O*
PF=*AS"JP<9TAIN JMO:6HT\7@D*XNP?H-],[G_$-I_D=?S283 A8_^:_FJ*2U:K?
PV62PL*7619> %F])&@:W(._"<V:2W%CQ)2%@A@@:,6IK)##K$L2+$T ;7ZCQG2UE
PE1)9L :"GK_'P2#  <K<621NS^>Y?J)_\R+/TB86A?Z8P='I/X2Y6<>OX,#&;TQU
P2 2J=&,I@A[BFDK0ZE4B1;FFX>>E7JV=6[4P1BH\).>2TIH"M3X..:K[<<PKQ5&G
PN_G.F-<_ILNB-SS*491[20$P\B"MM[L"#6^;G4!5"DY[>X(8MDBU7A<WY< #E:.'
PG1'KRL+3)$M5>  2P_0Z<NH>3>1X[ON],^+[*[+G)J?_TDU1%1O!^4GVPVO^;H8@
P0Z]GXJ.\M.TI&D^G*A'C U%[-2Q9,5MALQTK;-QRI( 6Z_()57.J'[VC1?J4?NU;
PXS7PN0X% Y*GY=2(P5>A,A:T=ZB;)&.]C6V28Y'O;@PMS23([ )[M7?QO]2[S/:8
PW =C=T@ O3[74%[/:,@Q<Q4*RY$(EF]:H3WL%2=,_=2- X6X3BETW4ZN<T?"\_CI
P]KMY4S25)):_0)AKC)C.Q8_2PT-H*;FAT_'&BU"][82;,,[E00?*=7&"F;-E^V0C
P=]8L\C;A4NS1G[H&V%%/S+^G$G1VSY-KDPN<1I,*]K-O2SY#^OHW#_UFZ[SN6#J(
P/LSMAE6FJ:KBHG\B&SSL=GF8&R).=U&1 FB\6V$2/GD9.P:Q )J%J<SV 5!)](V%
P$E)H<K:)(/W?&=U.\.P[N9&@:8AQI.5#WD#5LUO($7YD#L2<?C 7Q6YMIUA8I.QW
PM8EIW@?TW=[1E3L@3M012,5FNL5X!-K=YWL>P4OT=\)2][M.(U"!TUX,*@(!P<)E
P0^W5@R$\TZ(XLPWV5S=Y3+\8T"-D/5%R)'!ZA(NW\B_@,X3-D2*0#A7LH>:&'TT-
PP@^U(7=2[5?'QTO-N>0;JB;6IC@<:2D2X^1I3+VST65)J?P5 \'Q,O[#0DZ/NRLS
P-;Q]L2EK0K@7%]FY_E98CMR_B;I0..(7WVW*4:(K#/N+('C#X%HF+I^G7,9H;< #
P"BF: 31@O^)JD#\H1K2_0PC0CC#:,;K=>RESA0:_4<^=[<FYKTH/PQN/5\]Q^NOA
P!R43VM>RJL"T37-.!UT)6!7E_P8\^A#/_J YLO#F0GH,_TY<)L(X0])N8F,T/!UM
PUT5QRRRA4]28U#N!,=.&39JJS^2S2^$&H*#_MGH"!E:,,;;!?CHJIC8_*:NH30>]
PF)DZ"5G/77HK*A90Q'Y,DR4K2W\%&.G1WLR#T8RF;@[:JE$(S>G_3.O1,B-8R69^
P;Z6O<#G4BL' '5+6@%>A#LZ!\>*@VIX7Y"A!>T>\^CCJZSUC21;!==6X'M/?21TQ
P(+&6>C8%@NKQ>7IU6:W[1KHCY 1W57K9&*5\,Z\=JA,5XE&GS5E_EUVCGK4QTZG9
P%E20*9&OEV<K/6 X!68F64V!3S+0-/Y0V,FAU"<\!$5%DP7)QM=#?O 44 [YSUIB
PN_HH%OO/G] %(CY'O*\[8D+! *SR8%%5U:\!5FM\ 0>;V?I*V_!%?U][8:O+1 #.
PR#BH^#:H:$F]_J3.7C&KN%KIHIW^8K1)6'OUBFF=W6"PI#)ELCN;#AQ@S\?)5GZM
PT$8T:K96"1N'CE\3@=9F?*2*M(<1X-SO0ETX3]QE^J.CD7XOH4P^N!P>8@K-V=:H
PW@R"T2HE+HY-,B+P"//H%,A(K3R# <5Y_G\YQ_!% Y7NA:O.4Y^44R37NU]B'MJ,
PF5$&LJ]0 <  #IO+:W2?,IW&>YM]NG.SH)C,.6]BBH/(E:U-#,JXVALT+C1QSQC,
P#73C44*! 3BI8/>Z\[@8^_J5DG\Z12:Y5S5T\$K4U)M!5 \]80YIN\5(]OBU\Z&C
PX]GHT0I"!C08RSQ] <$B^9$"\!=CN):BY"QP"R#%]3@*MZC&8E4C:O,[$T_\E-*D
P(D,V1TA%P^/",ZF%M)?XMP)Q=:9RRM)CS=N%2HO&(4TW.3#&)]"S<D,6Y9#]1!N2
P\AV<'9)",H)DF.'WZ+X3!+K+\"UI78C3N*^L",1Y.[/^;@?\9=/Z/3A&<06-=:PM
P4+=(F[Y0H)YBCULQ]LKF QQ(2CQ,85T20"%W1+OQ)8IKS.'9>^8T?4K-1<"2%N19
P/&%CD=@,_K$+7(PW-&BJ;AM>Z!0D!G9]'>B^+WX=,7LM_TPYI ,YE8"_1SA0<G.-
PYAE]N"IWX:1 BN!TU^4BX9S $(M=PX'\QF/)R3VGH9RPNQ;%:KX7704(//-Q\ZX]
P,4  ?,$D:.+HS_-6UXIF,8IY]<UG1&*DEU479=+M'">U-Y_?,!8E:QQ#A^$TQG8>
PD<?A^O94=Z7=6R"ZG<"88_OYWRY$,WN7''/%JY%GLRT3E7MY;CW /-V@0E&W^%-3
P&$^UA"O(A=S<RJ;96\_/^..#\SNWY!6Z@Z)M:YZ@H\C* W\V]J,AJYS<2F2Y=]8"
POL7 XVGD&ANM9O'52N^?Q9?!9B$?XF3MIDTE*1/MXD&(F:H#9RM%;/ Y,IZQ?+A%
PD.'+1:?6W-(:JX?[\B1'F:JE*&ZB@B5T L?M#I-A<B?">;*X8';SIRA!._$)2X^Z
P;2]+>:+2*)H"#T0^:-@V(Z7E$H:Y:P)!@'L@HQAX8!,8S8;M9O<A>G"AX\(?0(>3
PDB])3^N5VI4U<+TR^]< +$MW4I.LAZJ#S;%]'B6W2:P)#%QQ*4525N28);C43%2X
PX>CXC*0YB3$MU\H5&=K@YQ%ROJU</4^N2(J[!W0BW+F7;1MA<A),$*EG7?"%;7+7
PSZ!KY/1FQL^M? JO&T-_=6?IS*!7HE% OKM3,GH[$(8[Q)QM(;GD6*)G!?-XB662
PV\7)8EY7X8-P2537HEHA_BG:-)AZ6,G!_YB*?V$:! 0Z6'Z/3@A M?0IB%C.\RCJ
P_\,1:YM?F&?0M(XX!F_UJ8-MG-M_IJ(CY=[Z]-TMVGTU,9GQ._%9/$,+/F8R96$Q
P4>#5'O?46Q]W?6RO+KHT6(V=8C.+W7IH&(B_8[+N&9%=BHF%R@%YC,I?PPYFJ,*V
P/4W$M#9)@?#W.67Y\2;$?$NJV,#1U7E5:CJ8G=A&22I%^CJA@0J7;N4(-5+D+B*'
P%&L3.OR36<\Z.W>%:ZF)$Q+NNEL*X.NT-V$:"FZ^J>RAKH\50GP^?X4MC !*B J;
P-IG#E5VZIP=7B9YN]Q'RI ;[A<!X7H1MNOKN,M 4%S*)"7$^ O)!B&0$AHJ8<XK*
P4DE7EEBXM;I?S:<(30//_ KJG!?BN6#Z)3Y?G9_;F0PBB#T[&V2TQ[D\.]>48 $A
P+$-3.61Q;_D5R)"MI%C;5W:9V $=U4XA@S6P,?.3%MMK"K!IY1V/>A:0SRX.;E0;
P57MY,S;Y]U$Z$&!VM&W7>8S#I^4[S=3@H@1H_H+_XL@G6IN 0)'AUEZ^T;8KKS;%
P=>MOQ2.P4ROZ$G,.G7(%,T-_MS[11\G#!;68X:"8P+H $FI,EIB8=@W#JZP;]B2-
PD'KR?WBX#/CZ<#6[D236UCQ^SS5)R8A-?-?*,1[RDER&H1\:B,;ZO0;/ RX469W8
PBGM1N,3H!+S$ _A_6D\L!2EXY<D]<%6VMKH;M*GDV#M8;:8;YF@6V_%JR;PT#WOX
PEK/?KO(RHS/ *RG$<L=#A!B<#S4]Q@%'&T;%;9HKL;6GY;&_SB5@Q2CKXGII'\]C
PF!'3'!WTR8X\1KI2=!-*A5&X-VOI,4\SK$'XI'5Q-PE>GJ\(&E+^B*;_Y6YO1728
PL6$=VZU$!4ISUKLXAH+9H%2_YV(U,%-)[THZ^HV,5066PD>9XZ3?W4()E);E>8IY
P<DP8O5X-62&9L[TYIFV[PMLY6CN[O?+HA&Z14?0R](W7A.WTZ7AK>\FD'1AIN@B 
P(RVJ@UA.7P&(]L#$,%XF&C_PN-OV_N$URF^BPTM*X7$2./4H&B]UZC6FLX2R+Z.4
P$W'(]>L_39*X.MMZAH?P>TA]VW+0J \X,2& 3W@6'G"H^""8.+L37>A@/6*/+N5"
PD(-W2PDKF^'2,?)>74C&$0&F_^F?8K%[:[MKQBIY<'0,S6P>U6'^H<'0%QJ>NW!Q
P):)LDI9O+%#! 1KE.2$9'P-NL#Z:88N0IPL8X43J,5/LC\N"=\!MD>;0M<1]ZNPF
PW#H"\RCM!<LSB])*@MX&8P]@2MV"%+T5!B\=$) # ?XRV9H0^<;W.PQQD&%@XP I
P(=N1^E0PC;2'E DGV4_ #-O[6-;KF&^YT'>?X/'>LGLP+VXR?$2TJ5J.?H5-(V 0
P/+NO4V--E4.%;A9=;?,_2<&$[;&P*]]V10I4*C#FDLS%!V>405R;[BP*_C+YD>8$
P#_QK =2%=&FAX;WM55JCU7%[*?LR&]L?1@387X]O8<Z<DW'_4;=QB.8H:9"4NU[B
P)Z$'1)";I/Z0\OHFVDY'1&&T0#=@_7@K3;<>+@U^QX<A<=5U];/AX,#CDI_(QWIS
P3&A64<8^P!:P?PN77'<6X97,RF]Z>?)L<)VX\D!-7N\F>?>)2>[;O5"MWFJ'71P\
PD;;VP:WE=/EC:OL&*[X2"8L*[SX(HP:&O:7#WF=/6L;E3]C&957GH4$E^P[N9>+'
PH(LR*W'_1ZONQ33S;>K\I=FPZSXTD'S/]P;FP;X91(V(L2L/6HUF(\N\8YV]_?5P
P57X$;Y@U%<^SE^%N\[=[AHZVY!H<VWPL/NMY5 71^L'/WU>S+H&'' ,9A#(CO0U8
PMCE6WPI>4[+C^4?%//X)T,?1[TE2,=JQ7W^F^^3$I(9_U+ D.2B#(YU'^$;BIJRO
PF]./F*E%">61#:5R6,;[+*@P^9\":;*1--0O4WZ,I.T VES2REQ3FC]U\5\.*%_E
PXVU/[;UQ(KUH8).5L+ HJGXZ4'-M<O:M/.MC-=YO68F.E\N;52*7!-Z0F/XN@F$S
P40N7E"SU\GL98S/28AF4PHI)[HT%C-,;#^P,I[!.M=5:D'82)\.P)!M=5?1!_4I$
PL%PGT2@\5G;D$V\U7 ;C>6Y_.S$:&N-X;5R3KV^31\I^Q50V>AA8A\03#3M84K#V
P3K#FTT@NMV"*FLKWM(,NB)R90 OX\UY94QJ/^!V-O[R&4E=RJ$NB=OJ29B]BZ,S_
PZKEY 9@FF)>DZMAM>FDF/&9RDXR.&/A"V6S@2V%U="^4+$V>N08<QZ%P\F$G]#:3
PN?G.Q!N=MK%AIXX%"&32.KS[$[WE0:S]@4&(?8;3^27#ZEC%Z20J0P:R6)\>#$>Z
P-"A5X9'[2:ULWR,Y\9$&?8MA7Y#I3)9W#/E^U#(>O+P_5^^VR99R^J1+&/TLS=T 
PW6Z/EZ,G"O*6Q@:_<DG&,SXW1 '3^^6Q"+5*R#2P4BSVO+;-9P%+9Z21-"B,<O6O
P1@NX%+G33%<]BH>U7JL@INN$#2%9 <[;&2:1XU6V12GJZ$F)HYAA)S,TQSFK%3M?
P?ZZCC)@ZB9AO0CI_L>R_."GWJXT;^7X6US$L[Y%M@#O2$+B\.NC]5&$>[_210A4?
P?E^^8KU 2CUI5FW;FVM$OR'*AW_IXV9!MF=?O#>)Z:I1^2W;X_XO65@T<;%8Y4+$
PF)F1?IT/_DV7\P#F5#R&1^C7*6\S[CM9>B#5K^X%E4RF'YKE.P8N__LY#8U+$+>*
P %:]&"EBS1D67K1TV;SD5RPI= 5;%543.U(S L%]ZV<L?S?+X2Z 3._IEOJG0I+!
PZ=63@H/&75_\X;*O8?7KVPU7&JXU3(!J)^,Y5T9J%37'MGP+!R6,[U_K6 !0B@"1
PH>!E*< M547V:2U<&(TH+>" 6N'T,W;H1N;')CR>%]LJ1G4$")K*GT1NH>DT:O^2
PK:F/E 'OMR);F^!)=X%:\<RNH5I('4")GL/X8KX C$E#X#HKI,T#I@/M;VAAX>PB
P?I=_UI%6Z^FW<EQ_U0411OWK.^Y6 G^@]#RD3/A]F5Z/!RE. =I24/(L!%QV<;FV
PY!Y:[RA_Y"DMB?4@=::7$%60>XZ7?8A)*L^9&O9<3$.[I$;0S!J4:F&XG%'H_S56
PVM$>J,;0"UI(@3]43*+RN@8GID;!UAK+5RVTFP3-;S#\$'/;6'I_[3I\IC>HF$GU
PQ:00'VX=Z^*:F@6_\CR=.'UQ;3*J+28//7H)Y6>-$O]F 7=5+8"PS)5.V.W,8QF8
P.,K)I^O,6GV'TKLOA!=#5W&=/.#OGO.5C+ -7?"-JC^$>HLT&W#/P'FBPSK1\JU#
P')C@J#';C_G,M^YW*GHI6I_A;2T[ ?'"+SQNQ_11_RX3RA0H*XRQU=+Y._)KI0</
P(/QPDO_'VR>NO%43S'9:'#=\4>E7G@]B\%Q]!*:Y\@PJNJ"V[13ZW%AO!-I?C:&@
P'TBC_1T@1;W(\YTY-G.['[A-_J0*_; Y"&2.\MSJ2UZ'()O";]'D]VQ=7O"&%E\!
P$HQ:[6)]ZW1>-EC[G3G*<D)@ '\0I WL&R!< TLHKB&J>:1,\82C93DD[?3F )*\
P:JKQ,VT$4;$IZ",0D<0&<=/!2PC%3JG'P53'\ /#3,F&1BU\IERI'M+^JX*@HV[9
PHU$5,KC =<QDXWN\107JT]J_#]4 VJ$**C!&8M7JH92*^/,8B\@R5T(AMPW719_)
PBZ@;&Z\-ZP$IT]L>WMNUV(!WBJ:[2=2[)(N6[R/;R3(_Q&3TL- $5_(+E6W&EC*U
PVC]_"^VV\B('+DNYIPD=Z/S%;[F6"*&YL8J,I<]]K.C#'V4T-LH F+F?LY,GH815
P0HI+(#M5V)%CMDYWR4_Z@/! *&3Z_W<,(Q-]QG&B(&[6H%WHC8?.A1=KB24((LL4
P!09&>^RAI&8@RJWHZ[ZE@J;HSJ7<,IF1JP]D0I<@;'?4JKD%;6UN9\<FYU3DWI$O
P>98):9\Z]F2;69I!%'F%5CI?C[Q&.3#NA@)JLAA"W,V9-]61EI4#9Z8 ;+Z-439[
P^4(&^4$333,U_B?"N6)W'EP9%@NRA8-'@A(F=2VM"U^B??!+9C]W)PGPY#)B<55*
P<?-W!V/-<5"WX)7,6T))*VKAD?&R4R%GPI<8_V73"7$(N]C;'N&.WC_6*7"T=8)M
PDHN@^.Q-//?U0% 3.Z.0%D*%$Y"&-1^%T;[:1D&SG(9H;#C,HGT%T3*S?X@5PCT?
PGP!,6@,V36'A-S)A+MZ),8 UO#-OUWA-$"O%I*-5-YK",:I3#[N&) 362T7BT#$O
P:C/C;LRHJX<'#-LCUFO";3\<TBLMTQIFN:'AN'W/&&5R=K8L:3RPOC[-3S;??J ,
P$@V^?W9$%8]+/BJ&*A1^<)YI?4W,2 K#.Z<,J4!J@+?CC_; .-^0?JY6O D GVHN
P!!>'?EYGIXW M&(@"D>6HN;R2FQA;<^9LC1ZXFG'1$A* 'OG\1 Z"^6*"?O 0-?V
P8O&>',&<LGY!@ /Y1%M%9W\"PZ>]Y4KE][?Q[\\&>[]"NDW+N"(#C0 ;:XG/;?V+
PP4WC/$3+3$["!&0U2C]KA=" :^PXJ7 $VM7RG7L?7B(54Y1I )?6PPG @%D?+&.P
PZ%<ZHMYP_K1 !:2GX&!5A@& )SGZ:A_HJ.)]!.^?ET.^:/#.T\1#%3U=E1%;^=_ 
P.OVR])0#B:@L7/J5<SO;UWK*=VL$.B+])0?94DMF*2'"36I^JJJ>O"#,&TL,>C"L
P;CQW@I(PQ1Z'FR/J@UD[%4'%MSN @7HQ'QTX?^W$3D<C^]Z"E(-:2S]MBF;O[*/K
P;#"DNI#I]$F0N:^0P@"Q&7Z!;7 P/T;>*/]9V9A-*DI0<FHZ,DW>WV\1:1P.:M9#
P>2),/"[70!!$4K6QY8TT3TYQ&V$"O"]/,S=J9*)]D%?R\0#KF$,U>P)!=G+.W+!S
PVE4R<<=.%E"H!^6WS@R<PG:0JS=9H:<#Q9NL)@X/GL><GC5D?&5Z9H2\C1'^7JDI
PC6=Y) P-W,7Z4KV!W=;YL8IW5X-5T@\I)B?4KI%JYG9-]*;<]'M*-]Q[P-JKMMB&
PYB82, WJ"?V"3\<G.I )KI\&AR/JI]8UT]<E %F:OLN4RF.E*^I<XSYDG[B UGC&
PD:&5T&0H ('1 UMVKGH:S),453'I\Y[45MF]0\KPFM2:BBFBMCUK5#ST*ITC8Y1A
PYS#0+CL[@GC'\T>422BZA(@;J-/@QU@"C##<E* T(]S]E>%]W[_PO-NNKM#<G=@*
PI6:%IE>Y/I]\5T1+9B)-9Y6K2A$GG&L*H2MF!]F-JGTV-2U9JIO)Z\9,VL'H"%;R
P/2("-FM5_0&3GI,A FU.]K%713P*<A48J-&YG;8JDR%0V?-;3OGX6^%(4T1(@@"^
PGU'C"T7;R1+<@LP/)%>Q_X2;F91 T"U)N7Y)X:@!2<MI)?*I/->>!(!])GC9:)T!
PG+#U6"ICNY1AVVO5RT0=^V(.GA:M1%P57W?.-P4OW;(G<4X/Y%E?52[,[\- ^!63
PZ<%W8H.EWZ\(5I#$REY46W41CMZ+'JG^"1[ P8R72/Y'H"?ZD?4 ?Q*8BC\@+F?9
P#8I5?<336U8[K,+2_U-'@!GB]_QN7,9,W;;OF'Q_P4P27>BSDSC"1A##VMIQ9[C$
P D)*";3%"?XK,V77\)YX$*1_,Y7H'9,J2MPBSA$CSI# R>O33?1Q>Q'Z5_3X4TL<
PRZ4WQI,SCE?K^XO(6^4"YF-80I *%PETG4X$4%L@.?1/\(J"+ C!E&O7U]@<TOXA
PO&Y^A/4B+QI0^QBPBC[2T&C 5KGT:WZP6#9\9"J4\TEQE);*0@0RKBW(_0F#OB:)
PV%^:V>Q)F7[&@@A28JL-_>C/]>15?"XI#N^@;=Q?[>?] \=#4ZC"=LWU[O15 U[1
P**_U0T7^KU(SM1EL0@1.L![:F]2*>FU.S'HSS94;KECS?R\  WLK#1N?5'I'?,.(
P@QKG,-EEIHX@P9X(S1%85X-+&5P>VI%WL/O3=BU">E6"#/6:9V?*7,&K6LHIR7,0
PJ<F23%\OAD]I&T4_@#+# WNB25(J1Q/0DL'L&7>;_23WA&G2BM./I1AI.QR.^0<Q
PHBOI)/5W%4UCG#1M"K_V8VB"Y<H.?(*BTBXM @S-?GAQ1@A28F>X@M,6(S=DGA22
P9Z?"*N[CKULD:@!LG_H \+ !+D"C'P?#1YQ#@^>97,GAKA6F2J*X_(#4?( /\Y"H
PSU?M/Q$*@0&&LS^CWUG)3&2*#J/U^+J.I:"XA.H'\PKLZ9OF5:-/&J3#2#^HI]4<
PXI//[HVG7W<()(!*.FM[+VT!=;&/VDP'=2,-Q;."PLOQ4\X0"T3W&8):&M)W%W4/
P3>0R[*Q@H'9AA=?IQI4#-:'UQ]!>WNXJ;WLT_T?!H6J(!\_H-0B0<U6W$H)5^"PS
P_-4>J[>B^G#,5*$IG.WFY3&B<DWSJP!MW)!EQ+*/\_^BSGYI@O'+UNY6)HW/JL+A
P3';><A4'8LH+ [VO,<$AKS"O1RI'__R<XE7P>)] 29WX% Z/X.4<41A;R<-G:R'Z
PW6TQT#=8P&RAXA'Q:82$XT2UQ:;VZ-:!ASP#TBRSV(E.3P+@#+BV%22!7X43.0@2
PMZ[GD1(Y66B%(?K O*$BOJ0F.V!"*LA_*=0U=N2J%5A!OT]@QT7IN+3 D::C08[Q
PJ7B!Z%,Y>KSX3)@'N+JUU7Z>2D$H6N-3VE.7R-GZQH$+V*_'BH?1H;^:B[6B_&20
P5<_"^00VIXYR\;G;"$Q^C[?(+/*$N)%K^@1,,\TRK/>:OJMS^I)WUBU0?5=;/49#
P>GP48.E$VCTQ5##"X8O(>2 $D)CP!E83YO6S;1HU])0_],FRIKDOSD$5H=-0ZHLO
PR5 4>GP;Z56QV8*::?$*Z_'UEZLRD BI]'$B;X?B?K91F+DJ,[R4'@%TTRZ:#S[&
PTX).D42WU6IGJ^LP;)!FD%CKY[/UO0YF(1R]A7ZVPW+V6&O3 W0A]A;0)H<U0Y*)
POES6<;A)VS!"H4VM:8NI*Q"?I^3HU:9J2^?L^:O3?(],GUMR:BU7 _ 1EL#!#%30
P$.9V0ON41ED'P1'A76T=D2FTAEY5)E.N/((%S\)Q'F>5#P[&U.:<;U_@U6E7^D)#
P^#T0J"BG &X]*HM:3ZX#EHC<_1C&K3BKD]FDZ7UZVP(\C\J\4 &OD%4)G:_U3 SD
P0,,X_Q=#L$!ST;"^(?!P_-3=CSRV%4/+BG-E1_YD;8M]H[G:>_YHRLV]_#"IE%]@
PW1=M^9'6KXRKZR[0IKO)SC8:'^4=$!)"*]$LO5B9I0BSG\ A6'=2*IC[O;:C%1E9
PLV&_O9(01C>SW+P25LNF*R=NUAA.T+ASQRBY1B9LE#ONJQ %(-&#>TCDUG:56)ER
P;HNT@O-PH[S0.^+QS:AK-Q[T0N<9Z2IML99FV5)XQ9T#*Y",\6^3W-LCFDM8L@<C
P(FNO=CO77PSN1^P,58*&YDIZE7!X()##-+2WDQK/QUQ[2O%94NX/??^US[GVAY90
PC%4$N:M.Z&<DO!7G&?A4S!A?"MZBO%$Z-)G)>HS>[N$!1VML@<JL O@R<\3GH^4^
P-'!(22'==@N3$JI)Y;%UOK#:;J]-(%R,Z[)>-DIX-"XEDRCZ X[AE-XWZPTU.:Y*
PS2!C[+O:5T-BT8.V9=\.1+HI_:@ ]5S8K0>6LSF;=;7N"6G;%9 '3QUU^BB6T.!?
PZO1/QU6D0TL0)#2[<QH*I6IG6RYZG(4&8+DH828PL?-Q7OK5-;"IX,NS(^.LO:>E
PD.$O*PW,T>%/ ])6?#!W6-X,+!IT%9R"[M?G_3<,HT83>-UT?^T$ZY*&7=:?^&IQ
PHNO73:YIS3GWO=F^M<IER/C1E.)KA$NP5S=OL*6F:-R^)Y/DD,]OE;WF5P1,N*3T
PJ/&)A<*0P'06=XC^8((I;1G,/'7)6^+RT)'1)7X[[Q9*YTP)SVV$U5.]2Q>:L[[C
PYN!]OO&<OHJ0C*F[M^UMI0?Q5@S3)EJAS>IQTA5V2)\5)^8R8ZH*GUIUHDD5%I,'
PCLK9*&Z[_U#'A50B&$:*:/'X"P\]L<J;=-L*-OT1)AMU55.&7>O+2QV1D?/6X'\G
PLS<B4T1J[H9OMAZE[(Y6?Q([+;%2?\)02)[HPAKWU+&.7S^'2WRZ4E*P!R^I7\UV
P.5X]T\6T]Z=P8 59N/.\6FZXJY=!A3KL7$2*[DO[4U!V772T](18 ,@QZ!WO+6FM
P2L:@09U&]R ^"NCJO6L_MM\7WM;D)WK^7SH-T?7@$W-T9V,#GD.E?'^DRKOK9[\(
P-575HX.]90>%UGKR #OWUQ36Z[/J*/#2*8>T.#4E;^O\5^#PZR0^4CR_)UDK<F(3
P(V &U$&WF.V]\@9_T]FHKTCH(\IA81L3 /LM_(_[^&7Z^A/4<-0L\?_:6UNVD;F8
PK'2G0MCX?L_(M=>D+SG'9TOVV+62U_\:OY>(>=>I(LC7-D)[WD0F_2 /_T0K331?
P,G"ZQ?!+8>.['%7)YH+NW;?D+SYC/)Z>WJ_PQ])K*7QA8-\I,H"?%V'HE0ER*H]M
P,=XW*:G):.9TJU>$,W27@A/VTP>>.O0- PJ,QL[PS[XS/AZ;34%]%DT<7>CQ/16 
P5OCS-CCC03G*>Y]23>\P=70)-X2TP*5#;J-(,18"AAPB.(T=WN;8^72E&EL<0VAW
PU3Z^*W/U=VT S ;2A[$8P<V05'[R?(N2!D#4"\F3DH1P5_/)7])S8'+IDT^F<7-9
P9G>]7=\MG@LZV9P6@L-V520,)2(.CPE2VK.:??UV$+0B47;K$\-U6"7R.U( V!B0
P8NB1C,+>JN(M;G9%N\2;U2"=0MXFO?UXMYG<ZTLZE])M,HM?9[QO9%)72SHR+)81
P2S[Q-Q$]D@20D&RGT71R_&#/.A>XJ5K,>Y/ A:\Z;?_!*L4,SQ9=N99+ER.Q-JW#
PY('LS8/,)6V+"DI,TF7WLS6[1R*AY$A@_9&W*-XZ##G+^[[+4@&;U8%7N'[$\AI?
P%T)Y2DE_/K$W)W %W;)* -\,--MWVV;4#B'HQ$.$&8YX$8\9PGK,<&)L7^+.JAXI
PL,PRAC;XK:=:W!^XGCT!4X<S(0-%7[#UD D4ZE[O?W8[U>>SZ=/78.D%Z%,ZR)%'
P+PD/@_&H)07V[_OZ;")Z5*<U*[ (OUZ(:1C<K(OO.D5:WH2YCSAU_,2'("X[^4>Z
PZ?R8Y,4HW6C*:9Y87B\O@Q,4YN9.^D[78Z>*3*P[%1TK&640P]XD7#90([9W967-
P0/=9#] <87 &3>7,.#E34(B58V%285.3;CMHSYZ+T#DL+,E,L;;7PCX=K\7QSKR#
P^T3DZ"'QIH,\ HHYX!#>O[G\L&O"'RF4 SCI/WL3<IGP6JU;E+/"([.@UIIG17?+
PQZ5#FQ9A/J3Q-&&,=ALQ1:7/O1%]NJ X1'#-GZVSGV/QS7W3(ZD6\GK8WM(4Z0<2
PP+PI#P=9Y\TCF(CF5Y/5.)1>69XJN",UXT_#N/O?*O>SL[ZKZMFY8+#X8R!!;?=<
P:6GS$#DV%M:&29GI?+185QG= ]W.-83')6_,O2A,K_&G']C;@]S67HI WVAH5X!8
PCJ#PE\ W0S84)4467RB2P:LAC3K[*=\]5CC)B+ =R'$I$B25K"_[I1%].1#Z9*Q3
P;37M-$#P6EYA-5=@IL$ZD);H!R 5DLSZ=,BEYQMW8=$9V!XRA.(=W]-<ECPZ >6+
PH>_,CH,ZBW\4B:-&Z=4.[*JAWL^ZY/YEG3KKL*V#0EN:Y:X4YE"I31D,.5G,W"R.
PG->'O)(;K=^$3QCRW^,AO4VMAESW[S]V=J;M6(/JBMRE2=MS?79A]>1;H&@Y\2[L
PQ)8Y@B_4M&APM5VSA9(R'1SZ<*P1Z,KR"J$4K&%;-'/M_?T-!22A/E][?[DY&'28
P_>5*.CEC+^R)WP^4Q2>$(2B.WG3#=O["X#S!R-MWSRQ).9(B42-D7LQ2A/@C9*!N
P@IM,Q2$X)3I2@CINL&?:;\A3S:3W,0A:FHU1_KGI Y[XT:L]AA#G>1FJ^1BR_ -B
P@O[5,<7'FTHC0\?LB& GC5 'XBO\^9^DQ>SNHS'Q#+$UP1V#6N7=W8B''DY-9JG]
PU'/N!:]6F/+>0"$R/RGN%4U!I6^D(.N#GZ5O91H)+PGKD.,G<(+#,W'Z*Q(5821C
PD0Q\1</59LD2-[LKL(40I5T^5VZQ/(P342!Y@,U:W)_U$ ";]@[FM\'KZZ.\> .3
P)1/G)=L(K_3684F6Y_CGC>D#37"F;W-&2.UW4 P.M5ZA(CP'=<,^2=(R_ZS@<W<1
P8Y^_NX9/XG7,6@KJ&((2=)<\UN+L@B+GCDI[!K[5 C'B5%+"39I+96AJ;[;<:#+Q
P<=S6/W%9'X#%5LSE9%!3>/,\;4:N#/=0WAOT1'F$EH:?H 0<42]=&;X3)"KSBI:S
P6$&;RB3VH6'>%S2JZ;VGF)S-I I/@* I" F09E1/:VHC]U*F57;#5@]SA  A(<,"
P_-+>0#"AZ4(X%^;;*FVJ=P;XUL*;G0XR/RIY]7Q-9I4H0E=*.Y7RQ%=+,;$?"_R:
P,8T3+__5<+565R/IWNY#?P3._H$B*+)!XH[&/+^V([TT"IMA6>P/4D6,O<%&V*65
P@_2T/$7Z9!V,N 2%DCP^_;YD;(9]1Y9:HS/F F^RE:3O?6N7S"%$4Z?^LZ+HR>H,
P80GA,D7GYNB:_#2?VC,HX\<$+1(6)/_&(Q9?*@-9=B$X 6><'@/G*QC9L\;/JTN:
PW(EU;"+#;5WLZ9IE,=2_.ZQSJ]YH=>#%J;HV&]O^M^VV"V@HB:JD&>*1!"DU'P$/
PV3SL)OD_[T255_\%3G9):MD#?'ABM#R5)A_='^C>S C;@7+04CLGNQ1]$J>EFD"P
PRQDEY%5[)H!])9WZ@ OR&:F/#?8)7PRF=1]R.X2EJ<]O83TM9I',.*:\UI*59;$2
P'?L'LNMG#MRU#DQB$F>CIGO[CUQ:F*7%X=CQC$CAFJ&E@V4'7I&NEY4Y"V@<G$K8
PUPV>]R$20;A59.,AB#DXZ,_0_*3WIWM O4.]P"&2R^,D""#\*,:T#$%1Z,GH)88.
PCNJ%;,0:89S!!@"!I[Z/7 QL!;)5:--1V)"0*M,\ 3:IC.$)(19!+#M\T67=@*?P
P,"TJHG?I!>;RZRT;GV&W3.PJ<LN-VSB5QO31_^Z-QIQ+8U@J.3J<H$03N*YE99N;
PD28X"52<.]LT\'R7[U3N.Z^3/9:[:>TPD+22Y7ZP/Z. <7[?JIP6LPC1( 5Z2R:3
PL2VZU><(4RG%F\CF5#>9^4F0-T\D^[\_Y<CFB>70G1J.7H^65I010T*1#^_,^N&<
P82[6E& ?-*$KP'O*LL_,4!?\9^J$6+V^?W&@AYL+,2#;4YH&OK9NQV=C%9#I+"JL
P*_0\@W?:07@C)J[I1 &(09@FZYTHRWI&LPQ[M<)*DC&?@ /?OIHUT?/;C0/\50^E
PD3ZLB9W#S)%0!D%]$R5G2]GME7-DKP83S?\UW[^!)^""?_)?&B 9DFKD]9$%!@Z%
PXD)J:%S9Y2)K>^;7?S'2S]@ '[CHS<CM[]16/C2@IX;._@T<*]$?,=T>VZ_I30Z,
P$=+"?A S Z&G^5C>&%ZW]2(]3GDH#QARGAH/X*1%Q2F[P@&<A,>+EX>C(O15;S41
PTO6$)#)W<V'_5P\JN9K%9[/TQX[$AARJC+[:8;9K#GEXPD\ !H-UL=UX#!XK@&@G
P*SG^DR^@R2Z  JD:Z4_CEJ1P)#4J67FL& ;BDXB<$B-OWU<%:"&GE/R?GIY)>FK@
P4PXKKCQ#S+"]=MO4P2:UDKS0W9:+7/F%Y_DB\3WXTL1RB3^N8XL'L28EHZUE<3;6
P^1A72ECIXOGRK&0%>; B3&8Y/R?!3Y+9 R#*(+?7:K(2?+W36_78_ NI@T2^R2!^
PP6X_<PF>"YN)[IUYS:F 43N8X-_+C\.*=9;9<.$>6&RV0:+&V29U:;I0LZ2Q"7XX
P$MJV;#2%P^V!L!G+-)-/_*]Y\Y,_\',/ZF/_R+N\I#*].VAE$N5V,:-J2(^^K(V,
P&S(<"Y?=[(ZUR& 8$%^XCJ=H%1!\"!8XN]'HZ>K)FF@'9.>H^;YB#KOW4AZ!B!2E
P#-E,0L;,^ Y(Z+D&(NMQ@"$=JMBK7+WH!QO7:V5H>DO5A<I&<N*[QI/ W)"C\<+1
P/)_DO-(7;0:7(\1%[:H]'<5^C'B50QI,BG6YK!P$%EIC,4MPR35]##F; L&IXF/5
P_B^D;#WK=//22O: P;"2X OL+YC?_:SZHTO:=7SU?OUKR-@>'Y1[IP*JY%*L,)"4
PO;=R70*D=5&YII("G:Q-[>31@#3#-U\@VF09\90 %/&*2N]<:*SU"\9#Q).M2BD/
P2_(?/7:?)&0TG\#16,IY+&OAV+B"J]@?NJ+!&N(8_2I_<1&G7/],JMMB!#7B1[SI
P@1 OA'3&E8<OA@*K^Y=.MOEYWX;$F?WHQWS2,-P"0VM+2.RL$.";J644?BOIO=JQ
P!T;EIN/9G4\#AX#:<\"Q89&JR<+T5D20 _)"*G_8';$L(/8P2$T;/Y(FI6Q9;!+J
PO"LJEA7P@L#2M*A4@;Y2HL..JC>?+]P(WG]8B74>LU*8: R(79J=9'!@^R?ZTU/E
P,*8I]3D;^G4@9D>70^CP4=':6%G^JYS*8^HT&/0.Y7=:N*)I6@T)G3%.<4CN"RT,
P73@*#JBA@V?:EVS#J-;+R00VO_D'^TJ.RG:#>=IRYCY7\_#-IZ^5[]8U@/(\EW[R
P(;7U)6^]G7G"%XHK/?_L>3_TM[C*YQHYF!UL4:C;<>4 #F:$>K!\]G6.TVDWMB@U
P3U<WT.YL6!?O.P4="K9=8=R\:]7*P)#;#OZZTL(RY-7+-ASEYMR4K*6C4URKX03U
P]P)]6T+G:;SC)E^W5$-DF;UCC"(#R-%7YPR:MMCA/*I=X2B"-:9I9AO!5 5?N']4
PKTRDU%&I:SJ4"RQU=/<-^QY>LY73._\IC$P7J6N,%R.E/Z0.//B#3,2?M)D1P]Q&
P5;%$,@^OC[CIQ;&"@,;,M*@/KHO@$<0B_L[)_?/_G%15TRR8:"I:*]*-"W[2[[F@
P(D$*$$ZJGAOZK[B7/1D:&9.^]>W(VFZT'B\BHYY7B^5B,7ZKP/AZ%WFN:;?)K*_;
PTBOQ_67P-&+5!XH3V!) RW6RZ%M!"7SV"N3 2N$+L-%"TX3?7FT^4UD4SK-NS]2V
P+\@ Q%?U54 J ;Z$9->:] 8MV1/L2R #*/5K?IA\ AD$GF8ML:P[AB&46$\ BDO8
P+F[0X)-T'8.!2Q16C" 3L6%M.-V>2:C[DTE&<UC-SQ8;DCN8T8T>6EY?P'4"DE/7
P)LX-%OV]EO^W'6?>0)6M+.G5AG)!":FX_$VS8:Z+R,X%-%VG 7N*7]?=(: PMODW
PF@H;*D&R4D$!:PA,C#^.?6G^UP%Y($9S$P%%*F_($TP>IX&! *#X7ST 3=A/4XH5
PVJS^0U&/MR6_9UY]X&O:# (8/19T7A^DNDS#*GJ?YD\8'V9\'%Q!49GG((I/'>4I
P\V+I-ZP_>#]GH]0+IC&0PAA,I+']"2<77RBV-_'DA?WYWRKNNU%6[I<?_CV%\3"4
P+?];U\(X+;,<FFP5$$N ?:OA"@6G+,X0!ZTY[FKYS,%U>/T5SJ,SG_I^N6E;C$TK
P@VS%Z;^=0*P]FC^_ J3O2+.CNJ@A?^G4-CV"3=U<Y'9]^O+Z]RB,[5@<D4>"P"I2
PX. 0S(O5*<S$IKKUA&=\ ZWH_R@ OGN<YVAIC4V%0J\Z WR!\8?!?M]@\3_*;:*!
P,U@[RPXI&'#I2\)$^$HAO'Y&D;!C.-V)QUK&PP2@$O5:-G]$H>#;<D62+A6)WLM,
P9P5,)"56]?M59]X^244'&&URB_$2M3 XW!"@NE/"].7Z?RL]2]%$70>>"K3\4SJ]
P3;4%F^\!7AG3&I_DM42:IDB1PAN33P]I\=IXC(N?R/^ 0N0/@1@8>^I*X)W@EG.Q
PI]IL%KU(8\D=G':F1XSBG3"O0GAF%CHS8[D [YU[)NX.$';H>T4/@X%*3HD 42G=
P J?;F_*E0<IHN>*W=:FC;CP37HQ7BVV&C7WD]=<5]M>/!2B] A:PU&$QS5O? $))
PUL/_ @-0#23AJM])!+=/M=Z-!/G!B_. +0&77@K0$9ES#>!29(1_&5=@4ULE$!TE
PX?P^?&J[12AYD3AVV)'7#8#R(NJ%B]AYX+>5KXWI^WQI) 15CCD1LSB6$^+O,PDH
PU D+3.GT!/@/DB!:N;7>>8M*2W:-2.3=O";TN1LVZV!JJNYL-JO4WC(Z4D;.%G9W
P2>+5S$$9*#(\EP&Y5 '/K61P4; +J3?5 %^SE.4P=^[U1,0RG"BNL,T;.-UZ!TXZ
P<3T]N$^^V!]U'.SRO0+ASECG BU6.II@]7:+S9B+(F2W:BI?4 V[6%5'4D$$A@C4
P'813"=;B%Y\= SI"2<E!+B.F0M^H(^8Z2]@(41WP2>R,Q(^:]NB,CYDSC4-E>$)D
P9OA(#OK_C;3(2F"V6891:7,B#I:^_'S=6N;"K'919!7P( 8Z![XB&.I!]/:[1KN0
PA;/4[S0O<H,W! Z!J*=?1TPBE:D:XGE]&GS;"QY3SU\[8@:+\;6T[1[8ZFI(8%.N
PN[RQ#"3 TG%V*^:K$(1&R8\.4*QB%A-"ICX.V&M$Q!L!J[Z>KZZ/<O4HT9X*+[?\
P5#P9]ZGQ-RJ?'O,;R0Q6V8K^?K?]OCSY9EW_;Z4 4.M#2E]_\9B!A\_5(ZI3I6=V
PIK+<=MM@#"S;92YQ\/<P*,,*6&P@:'A%T;**)S/EY,B;RWFZV.V=GK<LB_:]X+9V
PH^(>._%;]YZGIO;JN' P6E (,.I*O"NO\SN+<R/GH,L?"NY.G)L#..G@M)2--,%J
P*=3:0?C40L,:6F!HW&F]$Z1=D!T ,4_V_<G67T@@=*1?-'[#+GSYUG+W3%!%J<4J
P2$OAZO<:5BQK'+?UK@/3]VM=>FF5/R$WU7!5%-:L1%@&Z*2]5S%K*WQ.3LF0].'Q
P[O49-;?Q6]NA77JKB(&#2,7#DBT!8>DWT1%T4H]-MGQ.V[F=>BR\T9-G$O-F/HWB
PA3LV)G::?]3J(83-04=!-$XY ]$C2J; _DE&@ZTA/OWI@RPT#.4*'*2USK4#(-,"
PB(9&"WF:!,E3E!-ILR6 HR^U3+X: G.3A?DBHF(6-GV;KS31N30V5&?7.I*W@?Y@
P";%W(=2^>+9>#MV<',*;](3969=%<^B(*'A>QM'>Q4,\OWP_ATI,,6J ,L(BN#KD
P^171%7]K)5OG,K.;+=YI*,?!PEYRK:]< ?"$AV!']GU20G^I,4CQ+#ZN5MK=2B_-
P_F(A5 P+'"12\+BVH\%V3]ED8Z50&4EL]IL5C^I3(@^W.6?6P,OW I"I]NV.'VBP
P1>(+@X3D-"3((GD4H@;S19&F 5$RZ!6,L6HH%.7,W^A=F(C"".=4'XV \QVST)RF
P*]E\I@JU(/N+BJ :1VNLY%]>VK'X)]JOP0M@<<NGJ$GK*25WH,G835"\M"..5I)J
P9U@1X(@4NW]K&<)BH]C/ZMK\R4\-C[VTM"VJ*+8X; -SA"I( T"0V_IC+^S]CVMQ
PWS".;EO$DF4^=CINW1QP;7S=:9.>Z3-0I$.91YM9*V?$F[[0C2J&OAFIG5!OVY(_
P96SB)AD?1M)>>HF$\P\@7/61@T+J8P>O1K()Z^$[NQ#!D:M/UE,CB\-^ WP$M]_*
P0/I%)#@U#>'7Y-*U,Q'2"&R[.;L_]>+HH&@#(YMT 9/,0F%0Q8*9XP!83/O_U.3X
P0!TO5U/QGM[@Y&T/V^4X1'2=_Y$M_N?Y(+:KE<>^-I:7Q%>RB6336;7C7F$3U/K 
P"+=E^!OPR3EP=33W>=&UTE1+!0Y31:.FJK<R[2UV4Q3M@<^L_X)/]/+>0[<B$X;[
PP(!(RJ1N"I::&98U\] D7@,T5HS?AQKER[*S 8NG$]6S9I2&JX9&H3H[2:-Y8V]O
PM'(&MCRRN,[Z^8Q/>I9I25#C<RYNLU>-D%=O19_K+-+ZFW?::8Y-5T^2ODD%<TT4
PR1QTUW0-NQH8F');Q5"A-A&F*=];W&ZVMD=F^O&RL\I2&ITW^RS-_*13T*XU9,)K
P$A-E4+S92=.=OSG"\ ^O(  X"XJ.FD_"3?<&T8AYSBZ>L46<H__S37#./.)<O2F:
PSJYW,24LZ"E!7,>VX,ZHSU7I(*YPB@^=(?&EDA9I2;6\DXGC>3*YE13NVS8Y@RT&
P^0V<NNDT\-[$D/7!(._8:-CPK?:KN[4://+M7Y(N^ =FDMQQ] [W4'\)R\VG.<^X
PE%EI5EJD@T9'E>-7 1C95UX!-7^=/I %?@H?*'&[TS")>7$O\1L_?VCB%F$US,&K
P/ AS0UEY[WMG9&/2FSP,8]_%,Z\4@!>RF2NSPTT!4D2-DMU/.,X2N/A?$CC8N[PV
P.-VOE^H#,JL_3L%NV@YDS#!Q$NB9'EB=G[W2DS(.6[45D[5WS;O]/-PE1 <ZWZMW
P9B$DHN>"AR_3/L1ZQ3YE7ET)KRWIW_!#&X3NWB+=R?+F G")_F9GYI$!6>OA-55M
P^;74P/7</R)-Q ,LJ.S: #"N,NB0H;L\4O[*<Y-<]F%[B'@8-W]784_A(KX7H1W^
P&T@F<HF*!F[Q%"&O[^V=LV P"%;5H'WPWU2BTPK9<.QK/O?'<^,%L<DO55U0Q:!K
PJK WU:3PXXQ&/<CB:+4["KV,E!!%R @8I2=^T4D6RAT3 S@SU^38-EY(9 #?^R;J
P5W^G[;(F=7>!$*!OW-^$C?(L?F]E2X-L4A?Z(TF\&@$(&_ 97&Z;6%6 #/H8YC=5
PD[$-JM0IW#A")$FUZ=]\P( 6&,Z")0;^W,N>G_+MIOD""<_6*T43%M?G<EL9B_QP
P*M7-;?QA$('G5K"FV"KIO-"..(Y89_"9X13 (D>"0N488=DO17.DDJL[.T!<3*][
PBRLAJJ>:&UW/)IY=,WTLVR!,#=%B9J#?=WO;U)I(19[5 Z3$8I^]XT)F^<[:?U\E
P-XJQ4W1)4X0T]8ZV#CP*IF@$M9FN"-%^Y[!*$1)[K;IFRUX KR@ )ZPPBQ6HWYAC
PT9Y?9L+$1<T&K-(*,E"4I8]?8W]W\%J0X'1[E]7W#:K7;Q0RK<-=$N,%8;L\&/XD
PEUOS:14=)&SXD8=0#DZ,D"/RN,*@.9BZ9 9UY[&5U&"RW(T_P//?L^NZB6\UAOQO
P<I\<EGX(-&G:C7M@(LQ[2Q2YV!Y(BI(U#ZPQQ<,JF O\=MU,:GY RDLX-<*5 H#1
PU!BSU0.K-WD%+ILL3G_?M5'[[8(-<8ZQ1^D#^6+QYQLP=.A,/.6F&X56OZBV,"HG
P_/$JN_*$109()U<*CEA.\FM(7=LFYR)V9@=F<_<I4TI&R4+\$F^E/D,D#Y,3Y*X=
PNC0[7$VKN91(8T;:.X[79;:(#/SG3VP!8BN9AMYA&K1FEOT]GLWI%CFY&+&C^O'E
P"/H\XM84ST+8GRK#>AU(^,H(BET]N YM/OWJ,?GBI^<FM3:&^L(ICUD@TM_*FC/+
P%F"\+84 $CF#GU !*S+Q"XIXE4<"9HG$#H4O_AB*&^=VYE?O6+Z\4+3%\-C" 9)U
P0-I&.G:.(=R]J$3QG;X?VRFOE)F?.<#TDP7R7=-3FE7L^O(3+,_*@D9X-EZ]GL.A
P)A?"]:,BF@ M:0"#_"K.()%8^^R^4(0@_E0IE>#6>G!:/K93_E-8(2+"U8A\!)&,
PW.5UX(9S>CSR<?SXZ>+F%*WDNG_CUVWE.IJ#/:D>LN+1_TYP@ZOB1GLTATE9%FU\
P#Z9 !L%JI5L*%7X"YUCV)J?4=A)@39/Y?KG)SV%\+=<.+SA->["V]7ZJ%_=M0D\5
PJ'&%8I;1L!0\83ME*\4@CM X>6Z^=8J5JKO^\$,PMLR^T-$]CS  A_O)/SBELW,>
P(WK/6>H57Z;'X.1B9D)+3][5A-R4 \)6]#+16$^D^$J\$V, N+XP.KWZWAM]R)T9
PAGYA?!Y0(2+9B2,4HS@*2/V,EW)?#3);.MYI[@[D<);@.*-'_"1G,/:&&3S/2_@5
PSTBSR<3E<I\5FGK(4#ETE-%!F=NM'ZZ6ITL39KZ@81.[X3'1ASW%]'GF(3I2Y@'H
P1@_-%]FUG*O+VY0#G4YOP8WAIBH,EO^V2PQMCS427>VYTNFRG'_[2 GCX8!>+=N;
P#]0 #5E7!Z0#%A&0#7Z5PXH<"/O8$/AL;Q_>I"VC1YTSB(>&?H:KM:5QQ694DX-K
PG6V_YX9I^-=X3>"/3RQ>R4FJR#E]AC^S*Y,PXX]3M%)],]3507MTH,#VA?.$XII@
PPI1RX6H VLJ?$=]CF6\\_OXPH4!+/(Y0I@U'T?0%]7K@)#&ZHLTC=WI"X_;&14Z<
PU; 0Y!-:)6EB/=8?G4*XDS4Z'P$YDJI6,>E/[&:@4<B&.QO$4S2O\[U]LO@L+(R>
PB2$^QV,R&0-@@7[OJ/H:6PMJ6MJ5@"*AHA(;'8LE0QB1QN ;C4P0**R62HVG$) ,
P Q]@'JRZ'SP*&Q8;#T-FQ$0]@L!]X/P,@<I$T7(GDHO1_X2$>DU:2^3';%NM/UA]
PL\JCEZ1U-3Y$EUGK6##LNZ*4@GLXA^4T'-S1X*YO@]3D6A2= >B"_6<CO2!!FXNX
P]=[I=I@\;^MRV@.OP-DG_8T76/C(ZL\=1@T^=,-BZO!M&W\3'.JXQS%Y2;IK]P_:
P[G0_?\(#'&<3_^X+_<,/=W)6P*5_1<O1@[XQE*!5.%Q1XH4U!=%\-:H_)(I=6@CP
PQS^4UW2/%1W,'-B%S!S\?'6Z80.KS4J@6OX0!Q)+;Y>R:\93O\[5[*>>[I: &\O9
P R7B2'_UYS@P#_P6766$07CRA:ZJK9]%C\:X(0>IPQ!>))F>XBE6?/E0+KU3.'&?
P %*34S'U0$9J4$O; ';<63*C'X,U,?)A098<4&K:NE)JJHS^>L\R4X2RQ\^"8,#F
P.0_PSQ_5$J8&YIK0/Z4E(])2DYY5.#$SDN[PG\_@?)Y ZW9^]Q)NSK.LJ7V,XB@'
P2EA]H--SVLLQ[DW?:U<GAT]E\4> A\:3F@T!>:GAU16\A>>3*#I)*_P,;]]6-9?3
PQ6>'H"\.OQ#&A@%,*S?=6?T-I]>P"J+-1 OF$C)=9HB[)B?1A=,K7P]+4?KQK56R
PMLE%S;L"-P!FL?>[+NKX'N+*')+7.]@=C0Y'T)7I0#X L-UO#0HD%LU)N4ET!Q<5
PT\C95#)#]/$JOP2\-KG2I=%W:]F[_T=%3P!\VCT-/32"IB\DPM=A2)ZK76?B.'&\
P?7 +%9\4_CY%:.YU>EY0//%(&<I56MJW3-=!E8PQQ[@>B4*4,/.5*%$/;HQ_;.>Y
P!R/W9XI&RE2M$BBK+76"ZPA!>%^+!<++V!S\A6<?GQ>")J*9^B#EIJBX8L^:!30N
P:H;.5;:4N'W0+E*8T/%-)=A1YW#N.!0I>H2JR-56.J5K::W,FI!L4<NCVU>%=(&(
PP/QI9!57Q0;.K(FFT%E 7$(OA=\I.W"AKY20]P&=R,^?U4+8/&;1!]4( PD>%(7T
PT&PG^4+LCB7?]%Q"JR=HA$HN5W"4L<5?A1D9S2D:6H"&9[O8#SC:78&[5C\"%I>5
P!V58*>HJ:-2[>,_^@=FZQAB?H<V=B?YD!OV5_[M#3;"/N$2N#0'$U?M]J>$AYK K
P7 8TUU.X"5PPB^E&_AKE__8![4FFW#G")G3D@10#P*B)7;C^TN+_WK/ZQ:C'33+V
P/TA#*X1S-''H WX$KY@Z$"G[!26RH4C.T*5S?]"8#(M1'%-&P>*00$IX-8HZE2_O
P+O,3)B!1"-=)J@)X='?)L,P>:M>=1 <WF:-=>.)(S,0K17O.&0B^R<T.=0GT/H>E
P@.> 5MFQ;Y4[F&BKSE^IO1)53=L0"F0%1$J( (3CMGQNP]4+ZS!8)4EE^T*N#*0Q
PXSM.H,2)SF7^W<Z@BRKY37YR?8W-N[$W/_7N7AW:C1H9-1HQL+$^]S((G*X)3HQM
P*<")3!=[3!W;923&)8[-UFH,=JDY5Q#1VF\;Q 0;3KKHRCE6A0L&7P,(SX1*_-]>
P^Z$/,WY(D0^F>LH'ULY5AH>YH/YWFZ;KT&W7T'RKV\[XX!=EZVL?:/&@B=:)'2X_
P@48>S=JZ' ,Z;4F%=T=]3(N@Q/#E$<E;)_UF"AT7Y^&N=C _3#8VE$M#;BBTED#5
PI2++\FFE/)EDX+3O@?YB>,^SM70ZS@AUS\5\4%<H8#%-% S:DDS_N<'%_O+U64CM
PK0MC=T!F+>?A#5B>!6KVP-'TM6N3IL+#3-DD#6LE)<RH4;H8<K05OT")@ZII2=< 
PL3?W$[I!P=%$BV3 MC="'?$Z C]M'T1O,R3DWI+]'KR]5.I,K/F\7=3OMGF@TQWS
PVE-5 J6XY^-4.M_@:ZE@)*,O(YG4W S3)L.V=1A3Y]@ +VIP:F71N(!BULST2J<\
P I[P4[@X0)_*D:VR@+#SPCH/^W=^0M@Q+$HS,^LJ9\O;@Y5K*>4;O& ;D.TVIXBX
P%C7J#HD SQ/??X_GZV]Y"B$!G ^14_.]=^6.5?N]8I;4.;A%>/IQ)-PTR\S\4 #"
P47V:Y7M!SKX4FB0>9H L?B"J#?JT #^.3R9H6[BH%8 EGK7=ZLI#/Z #6%@?ZF^1
PR2>7\HN$2KJN6L#T9R_-J+POO5RMAPAV(F-3AP=I>AEX01N[^I3_] &R,V+S?\/A
P,JJU]1I0]05=T9=#P!/P(O]<62ON8_PPMV?\HU_8*5W?*]@K^D1T_AS38/RA2QE7
P1 G"495%0O'D=4JAI^&%.X,NN;#N\O[H:F)G;2G9RX0>HD:9O88KP4WM&0NF=<[H
P+@$_)^0(=<L?^JQ/[[;]G;]VW$9";Z?@H#;1#]O@L/ V\&2FJ<(S^JK+18##+C9%
P_?RH>U*!D[" S3K_#&,,WDW8=*3=.\_+?CP)3M!9T2Y$NZ7F#D*.YT5'7!!Y/WUC
P#*XI_Y9>W=FCGDRM[L,H4X"I >R/0G:.R:]7\K^7E2TUAC(%(ZS2+T\E)9,&FYQ*
PCULO_=.W;3*^F.3ND.]D25G?O=>6,?:2FC-(O]HMK%O3< 2RE#6T0<U9?8?G14F6
P_MUD1U";-2V0@'%_%U>U\:*O"3#ZKT(+<D3HJ&M\SM:B!96P3%"UN_N<N[;LM\&$
P2@ZG5N>S];A?[36UF(\8K BU]?C&7@!FR02Y%3X8_XZF@)[# >-ET#5;VV?\&+JK
PVKPV/\-IEQ\U25A1WIW[3?F6)'LAH=%I>X<Y.9C9SS0;;4?WO$KUJ95OQMWCWX4I
P!0^4G^A$[5%O/\N.M%Z$PFDIS[F/+2RE+/>"ZMW,*0.;%R7"9L;=UZ8AT9&C=+14
P)+XP&-NRMTTWB?:DG^>@J4)%-ME#6_KO&&RY."C$P*K#E%'=\L F1]6IPJ/?);@V
PD.2% 6(6KRTQ5,7F[L@_ ?&ZC!^/>)V]G "986U\R/0H8#;\?77?K?%4R8&%V&/&
P ZIWVF@Z*N4VA1)'^-!^4@#+B"V?_>_$P#+H)8H*4.A8)?2_=B9P(/S)\$\O2,9;
P:Q<-%KVJ<RQGF=MDR.L]L%CX]G/,]IM=J6KB:6>V@6Q'K^6CQ#9S(O[:#"6CX2Q&
P\"GNG+>K["0X/L-)DL&[(ZD*W3:WJG&#/!E9-KYAZJ19LNUI"SOD)\V;,))![2F'
PQJV&!LYO;#[T+=\L27X DK^+DV24]YI-L3,&YNP]0[7M(B!)*D]K-Z<;T)KQVEL?
PL?5?(%%H?@"6\6?*E?SL3FCZ[<087HM0F P6.;=_&?L8<<2(W+S).N>Q6%7N<Q%H
PAZ408EMQOL)W=>$?-LZ<4B-W/#]&X!@S1F(Y-:QCNL69 ^(1OQU-A)G?)(1\-*4[
P/ 8$2=92DBV<%_MZ_!&]<423ECR3UIFFB8C!.M;D"QL>L\:KOZ9 :@CC(1][M3S7
PTBG>KX_ "VC:,_!N43.7(#D:T%^04Q:;(OY*LE4<T'VC?UR,I"*BH!41A4B?*WW*
P8M'#^38"#P\OVOWBL.X[A 0*A30;F:-6?9$&_^/=?K9Q0J:W9&1<N/I8!)#U1[_E
P 2G?A98,6M67\#N2"O::]-*J" [U#95^X!<[J"^V7F9).((E&0M;PVG;(U?8$0Z;
P0G0M]99[?VH^L-\A*9<CA RI5(7871:)R O9G.^4\=B.-1F>6+S4"8TBH& I91@/
PM&809S>N6YES:S.R02Y<=EDNB+,)EAV<:-X8V*(->_QBW'5SQQIHWB*O-M_=S01B
PKG!3P+X<7H,S786 ;*6HPHE^!/$L<&=/&-N2K9GG,;3*-=[=9)46DO1% [C=#Q>L
P'E!!%S1AU_* IR/.4YL^^:GB)#=Q?P<ZNC][\UE)C>%^' *+.4+?J/Y]+M?>^WB<
PS;S2'@6W4OR>(9OO#Q:H<*D!(PH[ME\<5N[<-^KLXUP72YS^FK1M>6M8>X5GIG5^
PW6(?IC'':F:G2Y7]*6<)H'+IB5G%W9W*C7?/(9W%AAJZ3WY!>#+CQK]:TTJ"(L^C
P =PQ BZ"6R?E<@ORL^4I+<4L(- H$G,XU;F:H-\=?NE*T2.92M*>'0^F8+%H[N84
PPM0Q958%T7,;))X)"PK+L)[R-\.UNTVXRJ%F8$OJD!W;?&",ER_KAQ^6L&(&G44K
P,^/B9$64,XH%%OF@]B\KDD A>\J%ERV'91B2UH4W()01PH*/J :*#6:+X9XV.CT2
PBS5D62I2ADL6C@4*X2$'R$&H@D)$39;,'XOE1;.U=22LSX&'H9=EYM]?TG/U/>O/
P@JX1K3QC=,G1FZ\?6Y7MNQ2R?P7Q%<;4U>)=$BP=\;:YP5W;#62&IQZ!F2?"^_/8
P=/,9M+G!!H(-OLS^R%%Z$)0TV^&&ZOX?MY"H>;?/G7@_8CB3(!8FE$$T?3;N!]6]
PSWVDM"@N221_IZG\0WOMG+6COK,]S!%'[ ?]M][9*5Y)%UX Z-Y^V03D+Z#7](BX
P?\G-=/R7H RIL"0M26W^^TVECQ@^^0@P"-JJJS5)I"'MWU=MIS;);W$%23])B=;G
P9GX<.^19%LW%,H8Z]W;BK)R_;QH95N*V%E\WRR[BF@DRPPC./!R07 T+!79@H_.C
P5I*64_OE5M#*FWCYHC9W-/U$J*2X;WVV>!]U;92#HWB9)-W#-D1 ;@:/O_P2Y01/
PVJ(%7C6PDK'7;KP08-)C']V^E-HODVV\")0OMXU9&.3+8<ROBC$:F&+&$27B)HI4
PN%K8>"6LCK7P%#9Y&LG2RW@UAHRL9C3"*78=J-[%!&-2IOR(M[NN0)9_-3;5L:[!
PX6)\PM\7%ZJS,.L5SN-RA>5Y0&/I3'U_:1S]#NJ,C(F9"JP/#T@3V2A,1L^]X6I5
P_O;4?UW7:!&@,!L2Y@/(?,HT-JX%X]C5?#')(.1/<V4;S/K.]EW?\=YW$-SR+!FJ
P@$](8^PRJ[?4H&;LY;.%=!M'0Q?+[5U(>#1XU?*57U,LIW^F$N5V;?KKSF;Z=('E
P;VF#;E,\DDVJ\V4KC'X>I2U&W?K,47-NZ6J"KM^/>#C8O^@C-_N-09%%["_R[06=
PD,7^>[4KEKMA4_R%]>.C1[)%WVR> UOQXN;';WU[?W.3Y]R8@$D*J6TTRM9+(R,:
P;&?0)I.7(<OCZI<MY2TU(=#8:#=<)VY]^4OE7F-LAN_(="U-<OA!_/=?%Q5Y%S]$
P/QI\:N%J*NFQ5/CX8ELB\B3V&2&003@-41RKHZM3+RY-.9AX@V)2&P&A#' :PL,'
P#7(+66 U0^!U)#*@2_^!GW9WE4!/P-?BD>T0" Y\W /HNIDUU)F%+8Z?P*1')NLZ
P-8J%IN <\KB0AV-K?]A 9H2XU93@X2AQB=->=B@E43H%QOR[EW?]K\$F%]:K\:2T
P?4E*KK(*E%F4XP+Z]S"[5HA.H7P<EB+C.EHCP;O<#TM"O"W%>#@FH('M\'($8I3=
PO W%:W(.TR7EG#,Y\5AON56_P5R6XAV_F62T0*[0K6KVAMWLW%%C*3&-/!_UN#]S
P*@[8AXWEI<[)+# CR5BI0SE9Y%MH\SX82#4E*>KLQ28/M .:0H2-X,'N-C_],&,X
P+L'0<P2U^>-FT];-S*2[8(& Z+:F%H0<FE[2I+LA,I/U&QO^2T/0R+R#GM^B536%
PE+6-U)3?.%\K&^= :J54V&V4IVK$CE+&/I-^WIB66S@IJ]OV!2'U)JND5Y3GE 69
P DEW4UQY112;X.6J+' *%:5"-S)<"P(0.K&99N2HZM#VC>,X=)#_><EAA8II[I*X
PLJ#"S)?_]Y4O! E><@GE=HL"!F=&FRVE_ B]7+&Z*G0"LCF:ZK-68-++ *(?C:J$
P>@PT3MN=Y2*K1&D- &@+Y6P,$2G<;]P;=4Y7(2:X"'@=N#BY>Z$;I_#FCD!]IO<D
PN@7/2F&SC#(VM>X>[M+><?YCTF?A]D1%:(L,30+7"GC;4JVXT_K[J,,R6K,E\D^Q
PGO%*,__.]I:MS7,'MKV_%NK 2PHXG]M,X,Z1R=WY;O'^=CVQ<5D@E."@=S=I0%KQ
P'(&?YPZ@_2S0@5F,54PA!-78###&AE4M,J9VXC#UU<FP56GW]"3,F>2G6!X5 ,#C
PZ5D.:Z*UR;!* </3'HW\K37J5YG-.ZWY[UEDHPY<YYU2WV]'NP6FN<1_S<>LEGS^
PYWAAX)^LX#V 42TT%RX]\C&B3D/H2VLF(3(CS%G<Z8Q,.']TDA@1:/.B1U='1/Q 
PQF?<]YF"%,/MY&VH.GW,T;,]YW#11;S/M $INT/$ZK<GH@49GM%*TL'7'L6\S?,0
P,15=1Z2?6U<S V#"KQPA/R1B0WW?[BRB..A<O)NV)B,I41I'+L<G[X^ZMCW3H0\_
P;;[?.7+UN/Q//\GQ]1#":+HRRVPQ^W)A.]K>P<57+5H,LY.4WB**+_AW\NX#W_ID
P-G7<U\"V1&P.+A0N^Z773O6=]&./5I\+TF@(CM$XYPCH72[91BY2IPI3^( T/[J&
P^RVZ#K82G,(M=OF<4143PO:J%[3>WYPY]38?*\BZX?S;\BJL8:M7,E78-N%L_C-A
P:I'6KVRZP)4E2)2^E1$!A_PTFR83+[O9EP@(G4ST>'GAM!$IC+:>Z>4 G&0'S=.C
P2;Q37S.I4KL15,^5HBA#R&I^'RGVJPWY596 RDU-:A]P=<)3'@KQDU]55-OF*K1)
P,8Y0>;X/HIU,:6@&,WVG(+H[2HO_K[]AF+??VA3R]@&U3+>!KT:?\;B$;R.<NL>X
P1L1A9GW"(2(X*(%>-OJFA.5'L*Q9P<G)YJA \AYL$Y,Q[<H=H1CZ,!?#E9BJ6 W)
P0(CV0D;0_5Q-.QBJ.\/;J&TF5R8?9)&E*U*5$4&RS:5C&K@7<2L)Z3J[-;V:K%>N
PAC<8I3-6XTV:Q0;/Z@U/*336;A^QE11P:1CZF4O#(Z[F1ZC^)X+4%5!RN?A)^(M>
P7NF-28.,6_.MX]NFF:^<#1G/"V>: V;<_>OU!!X.$?[^;%]3<]OB\QG87BN22S31
P->?RDOG]][UIW$LZQM(AK7IE$DIG)>F:H6$&0D JK*67I:"U8S<:QNEY>J,0_%(V
P\"SLUH-/;D04@RWX[;;O6VY&22>3&'KU0V,V] ;$)V KQF>BF#RIJ?%BJT CU>5$
P-6%D][Q4RL'J,!GDC(%S3ZX3(C5?@^OHSMP^<#*F*V49-G>51<J69@&6^AX^O\30
P"]:R*A,TX>#[#@<P&BSEAHR!! 1<9R&7AE+LJKYD,A4N+3M#SI8\\YKX%N8[L]SA
P:/^I_)%A]"46=:D+:^MUA"3P*4OBII5615+G!U;;5&Z,W@_XE)!B=0(F:RG+.>'Q
P<()A]N3EK(^=]FF*C'-/V%V58<A,<7=[/=X\.0\M#:>P:)6,_RGDO-9SQDOUIQ$M
PJ<-N>1<!1F)AWKEI?!$CL=S'B8E';M_5J-E&FP)T'ZX@;W[L$IW*C"2QJ/I=1&PK
P*P8>H=RL7JE,\=$A6[@Q/P2Q3ID:UI7F["XZQDP-B][J&B'(WA^G?RAE(Q^HC;$5
P\QD*QOYGS4$#E92Y.-NV**VF]]0'9^B?ZK@0-0,9W-ZA:X1W*D2,4'-@_QY1%Y*[
PA$*?##>PK@^-Z/DKE:JG6W7Y4. FMA&K3.:9&FQ Y\F7%9DXLVL#/6FBKHJC]@A$
PR>$,X\IN!#Y%:-QD"D@)M7B&Q RV0EF##KQZ-NFE-W JS3B9U7RYNQ*^+JOZS^J<
P:MM^ZCS_4<>EA7_D&.0FWXHKZ@G=#2!W$@*4>1I?+R<AUC^%6,N$F5F&*1W+,FYB
P23-AC]K5 U4QRJ:>SRF6>E309*]8_";OWJ/NAL;6.&;.[/H\+8PF-3HX,;6PCZU2
P=8V4/HA(_,/C?'EA3I0[M4D=J+,'Q UKK8U$TU=[J>0*W)FA#"[-6RO[A+-WGM8E
PAD*TV?(%JPG0_6+B7O/^#/U2:@JRCCL1Z9W#'^-,)F7(80H-8/^ZQ&TVP<L&,0K@
PF\-A,0%KH=4M[=,=0:=CK<786>!(&WTC;PN$!^]XP4'T^<]W0=M;T\)$%3Z73B^6
PO(_=0^[R7_WN^M2R,\,&Y+6"^CU [;DG&=<_#:]H;6-P%5C].^^[VEOZVM_[UC2<
PL>\=Y5Z28\GYCLVD%'B;VP>()SNPH,U*C/"D\;X47<6>3_APL_OU,D74//8J]1J'
P)(0Q[@OL..W;8T;[YXRRP%V2B6SQL63[)AC)/_U+9:'N <P26EC6-;-&\HY$K=W>
P7&:7TY&U:@9/PD48 LU@%.5ND[?Z+!U#2*S]+K$92'4ZW='.VH-BB?UG\%O'P&^G
P9^ :*UYON/,=]0VX!29S_M9;X"W$@X+ NF81+>:W#%$MD,5D5K[E#.A4U%#+L>+E
P*S<A*$R:C=.Z='7JOFW;JOE+#/V6P!V:*+T.H7CYL9\'R/$G,R6: :FG)F-J7'R!
PO\!_:["_4D>+F['\YF(#23:<2V;FMGO?!=&]9\AKAKFF25@/$<=WCZ#,OQ'<2$S,
PVWK#I3?N$G]LU45CSR/*MJH5MOG"VV!"/,#C)[K!K"]SKFR!8^CL^OXYL?5W!E65
P90AZ*BC5Y+,[QT"/30_J';ZO-WBG4]F,&,$G:'*HXED&L<I0O:<WX\@3 VB<PV0$
P=M1;V6A-/4 \M9W\7]Q9Y:$]&3\'$^!9U0',KTH2SQ3<:?5XC)J[VWG%K,59L]0D
PL7I'5N%9>8X'*>RZ!<;"WIJ+9 R,N#46O57;CQN<F9R\S+ZB>R?\40:-0LPY^)*;
PW0OF#@4!<F"CUJEPJH:ITP1\EE 6.]4X=$% F!S2<=W2Q(7%*W0I+]HZQ^N9[3!!
P^XBVEJ.-NG>7JO6P;_M^?ZG0[ML<RZ*3Z TKNNH1 $$G5V6_1UK,\S?W$9%?J<YK
P_O]<'M8U3W.!?T![&E<03F2;J/D ^#T1?OHZ1[>3.SGW]MINDN&!@O$\^^E[WPCB
P")^CK(UP*9\#EH2M8,'/TB.P!7-E*$Q/ [G,4D]89Z8$-^23VY\EV)\?PP2"EC5@
P]K&N?^)O(+\!\_8K<8[:CW58OHU\]-DR)<ZUR_<.HE*:#[-GF$0X?Y'RSW=T\=D)
P1MK*9L&_P:6A)G4?& C2#1J&3*KL8,_$(4''](0+K3]F/M\8@N@JJPJJ\Q+V3HD3
PC?2RK,=$9@E#=W-3%C"!?=5X-3P_$Q&-J%N(_J@-[AHG)4)]\7-1'L;Q05V2R]SX
P]EE%46@>TKI3VV(I_].S8O[9(9W"#+F([1X:S;7-NK-=?;4E;9Y>']L.=VYN&JUD
P.&KV+N#D=?YDDS"!VFM:J2&!R@*B3_#GV&+P@EQJU7P/;I.8P@$KTD]ZI&7=4^)^
P7X0!+.2R)9CE.P<CR,Y\,$S9XSU5Q,MR*A2X6:7JE:K=^#T-L9V-_E&%0+MQ;'9U
P^F* D"O/L)),%Z5H-JNLF_X?0YR4J]K5;FF"-- PAF]O678(7@%-1D>J_']T*Q%2
PUXH<+SG>N8+.7FZ5@)X1TW%M\Z1JK;D%;*:\]EI2<Y4B0="7+3+0I1*%+\KQ2(8]
PY^L/B1L7AL:/_-JC&$ZR2^-U.B-&1%$/1!\)($?=88_EX(1L&)K=$VXG-HX,W,Y&
P/*XM&X@1D/DL?JTE<@@\:2GU]',TI_2%9IRM^6;&!.7E1DWJ0BBOVY35?@:&:/L-
P&_5WZO+*$8Z])2<=%:V.3?0ACT>.#)3$&2;\70Q)3'UX5/E,F^3S(^S'Q@]OW%+X
PN@?C;\\KLZ,(X@L9M^"[M=5G,H%<&Y>4(7;P>UW-B#O)>MQ;-\TP8M@WP9=S!$+<
P6N)ZM2B,%KCW-CF8Z>6.#2 H&,57!:@2^EALP)R68;]3]0$H!U97\8/.^XLMM!K*
PQ3_G<)"'SE<1@Z[0KWC# U)=>B7N@C7\H0$X!%A',=$IYRLFU9T%,O_YX"H^YR#L
P^,4,/-G6()!.@^2/KLF@W?)Q1O_'#Z#[/5:C,?HCF<J#_I;V.JK#B>U$K),?>S$G
P3:M&T\T?ELN6$3G]XW; R_9.KG J<6;39?V(%$!YEU&I!,/Y."2/@?%=7UA:,3*:
P+):.".W\S>25'!^<LMOA-GP+(E?0[+3T8UHD*,#%W4L:NK4&>8EAY@]-3KG]:%=3
P3ZI?VDA4UGZ+C;Y)]J\]SXVA&9?X\B5,G".^@.95P137N#ET,'&Q];]TNMB<'3>Q
P+</_%?410 ZF05ZD&]<G7-!Z,1&^7;_!)GES6YE.*&7E\=:)WE40DN(@KUF1>C2@
PIP;.16?_CTJ1Q+7X;!>.WT\X/E0S!IQ?:Z@\=>&Z-U0?(-BFGASEAZ !1BBPB]V5
PW2X,=[1HX4<Q(\AW3BNKOQB+YBZO1_)8H1M/F(T+]0[2KI2E5'N$J?&)A$;?&D,>
POVWQ =#LHAX^$0GKEY56?7W 9G,8GHV&"!U,]B27WKD7Y>'3[UBE\NIM T>7:"$'
PWY@O'Y<!Q$QR>O&*K*:2Y1@:\:^:"%Z@$6;!Q%4NI[FG.,F A8FLC:Q?F5WN #8@
P&^/H]78&.4@90L*X$PT@A2$<.87SP!)6UUK$@E)$AM!XG/'.P1,?=&Z\1=K?)'H4
P>5OR-(6"K*0XU*\])&AK2'R%%8]J0K6^Y>-'?)#+*#"OG_@LQ;"9#&E3"&NXX0Y 
PU^Y^3-)8>Z#V3%4X+#(6I@I'Q5?G04/EZ3=V'N/;CM+:#*8Q/4LSMD65^.) 7[4F
P%REXH&-<(X1?5B]R6O4>29(J>%8\9[K499KFG*O-<#\,KIR^G'.G_5^]OM,WOG]P
PNB*<2_N6A2,/TETX<C\BL+IG&!>R\!C_X?0/3W]6AJ1QU>T-957!&J<YD-%GFEV\
P(&:H#=HJ/5<UBN,W*GGDHBTW(2AL>GB8_M'@-@:6\6HC#/ '1>Z#J,'T -RE8](,
POCZ1J!FGVMN2J7.2&R1&MGHU^P$N3V&)HDO*N<EQ?N4\=!+X?##[.YJY+S6#NY8)
PFIW+8>^.GQF\Z>,(6'%Z*_""9R=\*\/*;<,/'>W[1G[-6YIZ+[=8C6]^.K""$ET?
P5'@#SMU518[&WC#E3C"*J#X#+#7OYE7=H;ADR5?9_?: ,_ZB>)VASCP)-?N7.4PA
P$#H@5C_']Y 4_>MH?7]3');^UU5WX*!G"'#V\#4]Z"=W%N*4N8B+R$Q7P;XU3"[N
P/GCK3=Q'U#CA-./*8X*Q(N] 9O^]<Z0B^'T+DXQ]QAKGIC FVH<)H8!90O=:B"&Y
PF$W.,1>,*1LU%SX22!6,6*$@!N":2Q@9[*3@G$RETM9GAF&Q.)AH 3WT:&1B-NE0
P0)3LF5#_AM\*;SNEI^-VJQMH/=\R<RB0(<(9 Y+G2H+/++I$KPU4;AR352&P_/AL
PZ]^;51,JV+SB.BQQKE##);M$ZJ=@'T)EDXJ3*Y1(W,_P!MK1@1K34'U\OH/TC4]6
P$-(CX3FM8T<1M#7??T!XLM]JZX]]K3LK>S4,M)W /NV2Y;(@BKFO.CU(*0VT4D#B
P1+/@<"@A60OJ$H\ 1]Z<OV56]P18UA!C:>ZDO$Z]"!7._4YHA\;R ]3):]IO$S3%
P.7BFZ,-DP$2[,'+76.28JAXCF^FH\>F)O@0]DVY7YR'9!-S]!#R\38N6@IE'F^FN
PH8DJ%L="JZ0<U0R$"+[6,E1#+& L* 1!:0(4RNN8Z?'G1X)SWJO8UD9P]KE( #VT
P5T D[+)'6_!^S@-HDS?LVZL'1BZ-4RB\@21N](]7_1RBXICM^>E$\X<;FF&FDZCN
P?I%4>8=[RQ.'@V;#63Q1)_:8N RR()U[ J8FV7W#2KW_GZ_;Y7)&_RL+72D%G!!P
P#GVI2_SR\/VH*['Z'W ]>>E<)+R7;O)64U?$V&=G^!.+X +*S($8(#)/_3\S59X]
P 9_4S;(O(CF$%@!.. 02PN7':=0I#@'6BG(&-;5AS_)LLW[%P6.*Q]55*&)+WT48
P'M 7/HP 5X7LU6]Y3B8-3CW9\!IJZ5.&%W8F*H7Y4&L- 8%[_WSI5&!XR"=%KQ9,
PW;).C;"_>/:WU\65VF@]*F"D?*..^]S$5"?T#_14!(&'$L?<-:-G6S"[,?8-W$(5
P%<NO=PDQC3E7?:8/]3J^F?/'S 01?#&&M@3$N33_,N4%+B>2,!<KK-^'G-CK/,#%
P1B,J]$FSZG-8#(L2E\;G1)XZ<TFEKQVFI2G=)-I?;[NN[^9+Q@E;%A7D0P(M+:VI
P<UTQX/A#WM# 9*L=BJ3)[]OJ:W/ZDZZF(BGLF2PCG%T5B5*M7/3^?D5EJ83<I#E&
PMID+G_U9VFU8^#NVL[^2%-"V)^%;JN-D;C=J'&D\8.J\_OA :F;I_X';X:NQO_S_
P \_<'60T^[MLW\^9BZ_\BT@68Z#JZ/3FRGNT=<#]=O4B^(TTR+^7?]9:2XEOVTP,
P4QH4&#^7W0XY2@^BH!UR]W(YI*+Y_K<%-*VA<++P]$"Q>Q[!78VZ"LL9H-=/"+@+
P_5E%9IN(XKK0^[) D?T^$S="O6O%R'4_9O\B&2D\D#EIJ6DEQ6R)EY%U:FF%M?Z/
P%U6"$#N-EN4+T$ 5"\]B;;P4X6JH7+FY_$.;04_ _(L35&R6V"0 S <$%@P:I^P%
PXETGL31)J@_RQ^S\8"FV@5D9(Z7:AJ)2!UQ2&%R9E['0K>'3'*TY<Z&JNV9Y&Q4$
PYA6B.H9;[;]6JNLR"V,+,?2>KA7O=BA)EAB7C<>;E<^22;@$^6&["4J#%LN\%-J'
P6F_9?S?\("#P!;=QA<9<$\\&;@9OUOA:,U.V2(^\82?A1LZ&Z-(W#+ &UFP:="?]
P1HI*<R.D]YS/@BXF2;")Q^EIBY&K#@<T&(?Z^,Y%P9(*U0X#);NW&IGP(BP^V'_,
P4!*%765\YE>JRH3[O"].D CQ862 CX'\<(4V5HC_.37;XH="4_)!J=;4>T/43TKF
P,RNR@K!%"6T&#&<$E?A%=(9LY_>IKJ!O<"%4ZBJD,JO(]1C$Q+N$![IVR&A2_2*9
PJ!K6'98?5TO NX>CC+@Z2\0:HK66)6UCZ,*4:MDR=F%KB$8C1Z=N*&E.-R%QB1/%
P=F/2!E0:G=0> 4>;$V2NPY9^(#8]"&WUU;K0,AURYL-.:Y#MAK%N\C&ZZ[X3>^\2
P4:,>G$X>CM2^E ;^S(;$$8GJT]T]$%^;,A%W? XE3/$\2RU6G;:U(CE\8JZD?HFH
PD"2-FL=OSB'4C[3[Y(HY*N:*.+KL5!3*[\Z:IY@*Y'%#6L):;\Z\VJ=OE1 J*01^
P%&R^UU8J^,#88&1IN#)"7]^&QMR''=8V7'1F'RIT^QH?\,62F3RV1EA8_W.)-IJ5
PV,6?)'LF0.V6#CHX)! =A%S@\L0-?>27AFW9R44&E<1#OF"6O[A)C^R!Q<J5R%E*
PX)%T*1U'JJ3/1XVN0UY4]_!UF$^P4L!3\S8G?QYY-KS&JI;!FC<[DY_46,'K%5A4
PCQW*22! ) RL8KCTP4<6"8B581,!66GC?3\Q.U34A&A&$02,?9;#(:1W=%C;DB0X
P/JY*SDQ4JJBC6+EZ[WYS)KPDB[7(?UW.WN.J*HVX6%W(,8&&;>I<ZE' BM(C!N/E
PZT/[O(3=*]/L+L:] 'LDO4DB/95"-'_M<5A?='H*]E*N%A)Z[4 ,T/=KCIN67A#F
P/8Y[UH:+)K]S]:DR"%XCHEZ:;^S33ZF^#9(^;JG,N_$?"-L*&J[L0%Z&J/%B[P7H
P45B( U8F[6[^<P1@7UH:GL# B"(0P\&QQ1B_7]2<)[(9P"Z_=%;EOF6H>O-WLVT[
PO69"\J:C2M%+W!J>WJ6H<0V,CBBOI')@@^H\15^-45NB.F"KK2UJ^!K*B:=B*<.T
PM9)%D??#M?GBDXF*L4.#.A@\-GA<K_3/JBOSB T)V19S7S91^0^OS]@0Z3Y>J@EZ
PYS'/%Z'#@W[-Y2$:&U'C:--=5R]4(>=N0J7*4US:>,O*;5B\!%:]-HFPQV':V6O"
P?5Z;3$7XY+FZ8Q<7(N$8F^W5FY#C%5E@GXL%5+#[;:Q8[^$BFQ;3>EY'XAD)T>'B
P^ZHIH$6N?@9H;*,AT6N<3C<@9-#\*3?90MT& D>T."GZ':T1,60Y %4LO+K:LV.Z
P<5@S;XH5>4V)C%X%.* )F#7J(4?#<&9L?KY5G/%D< GJ@1HI-K\BIW.CT9PU:1?$
P<.&<TC)V0M>$_D GPA3>VO0'Z_(W&,97KN UYHYW#5F,M[DV"50]=$4T/2LZQJ0!
P;UES8->]7^GP\4<4[,[8:K=/,HC7;08C>SPV.:=0IX8*SC!9570CNJ52I7V,R^ZF
PGC45N>Q<5;(=ONN:ESP/Y(LN5UMQ6J/P#&40K]O/XD$U3+6[\2\UHA*Z]T?=!HL_
P+VPV"4!313)7K@GKVZ$<:>FF (00E*#Z ,CIELU7Q$Y*"HBG.M(L2SB#.K.G"D@/
PP]*#G:$?8P7[0J8?H/P&T6P>,/2 @;B:[[J^"Q/=P%1UP8QUIZ47WB$;U2Y;?K)R
P1<MTPY-,"('(U'\U%=!W6S>/)ITX2("!-&UB_  C8M)S9:S64CT?K_2]<V$CTS*^
P0-1<[+"F87\AJJ;*!HY9HQ^((HK,ZOXF5IS+.X BBFOL!W2CW4MKK\\$-'[0X \K
PV?N.M&(:.VW"P96 <I788F,X7:%&9*L'^G.C!S_#TW:%SO_I;$@R@<J2I4M$8!W[
PC2EE&,7T3$1XV:2H?% C4(Q=$-"1C$M38N"Z*ND.>+G86I.5J[T4_]W$]ER "!J)
PNJ"*&BWG=A]RX,JH*^>FHNC/&8RY9$(8YI!_1^1_!E&O1S1&FCIG^^,8,\Z4C1'E
PUPO25^%O WDL!OIAHRSYC/K%B*MP3H(U'Z-#49T;&BB&)XD]HRNNM?WU\!ET-S-$
PS4V\E%3J%VU(GP:YQ7[G5>+=(K5(@,X),<()Q6<$Q1@YRDUK]TGI=]"%;/[PKTC#
P(M!=^X_[@R7YV^_-5EDB;F\QIZ"TE/L%5]C>0NWD4VM?3BQ*HI>=!-SMVKRYZKI:
P^(]^HT8=SH+M?G"@^!?M7(9BLAE'-3J]B#7;UM9>24T06??X9-']V@+GBIL4.<GG
P== :!R-3]75?PJ\\?3:@8#6CE*[(MRI<<T>&J#PVGLSH9%B![MXH4X3!5;4(?X6B
PZW_0OL?<H:5$38NDF[*P"$8[]1T6K3"X/O:AA5 </30*7YLV>_FKEW,A<282?!X 
PT N<WU2?SD6VV@8Y$VR$/=/3ZIQP>SY"Z]5]^I3/_1VT@4]>"?I\\DU*', 2SDK+
P22E_1>[-0B%B"PDX:\AY.>$ U"&Z=),02=D5YOO\/\66.91HQ=JQ&:\4>E[-)A%E
PTM9GC0<:GK!T+T(>@<YI!8P1A_FS=<H7"E$PAF*,17)L;#J1=$Z04*;7-UEN+@\!
P6A @B\E]S&'"[)IL'1/Z$1[NCXUMF$,ON1G?8"D^HZ"!-D-99?V/(V'-?X7G,]?+
PK4?A+83W>_%5HJS='7(JQ@D\39C)^XN1S\3M#KKM%H/=.VI6I5$C+.SN+N?Y]9D+
P:H?$(E4T7MCK$CV7L, Y=._R,2J6[2C;JR#T'H73' _2?>_M1)GY%LCI4K(QE7L6
PG!/N:)H__]_+\_X)+X"B$Y[_,R"*?3#>XL?Y:OR*V8%YTH6-ZY][D&U0\MPCKOT?
PY>;$]OPVR#85D9Y%G]?#%=S5WB% P3OU82(J0GH&0:S;2&FCZ(E,B7&1/9!]+C5=
P*<NG=Z 4EV)&3[)):[+HE%3+5V:;;$(1F8L+S<D/1V>F1H62EA,[O<PA-Y5*@SE%
P AED7I*IU[)KO90W.B^ALK<HY_[>W",W5-A(R!XA>8,,N;JSHC/76CD2%0*8W53/
P97A/Z"B@A@22QN4M8J2K>?*0P[Z.Y\PBJM3O]&_ZA-KEK!<,_2?==JCE$2<9H12*
PPA2:_2=WE7.9T_CA%6H"67E)AR,^Q+ZB==S8$%"3-]!^K4=(\J(6)H7R%06H%6.U
PZ0?^84W@&W^3\U,!*6(@\E0UPQ!SL*2+[4?VRV:_'LOG0QCN!=MP$>QXWK9V:NOA
PO<U7D 6RDL+*FXB,_RZ[SX8P,M%D?(C4S,*@,?F<VI'8G[O)I!>W0[PAAN<"?A,\
PYL$%C"5%.!Z(D#"/6.Y7& -BJ$]2ZC)"3Y_R[D^FS8Y@E=K1O1N,KCD#&GAF'MOP
PC/[TDE!"I.5<1YL+47W@+BR2$'1UK+ V=)4_WB%<+S2. @__N@L*N:I&9(6M!59M
PX7X!BYMKZJ UD&:8(NL*I<7]PB[B"/MC416^E\9%,)\HD(7",S8M'%U_(Y>$?"7G
P.%!AQUW\XI=M&^J_WN-U*&!LF-YJ4@NW4AUY(%#N_BO#='"P86[5^6[,D[8ZDTZA
P $0ON@I$YI%A1-\99OHH47Y2.NQ8H="X<+\!;)FUOX.@K(4OAS-O44=YXLF5!YI9
POI6QFN*V*G,BS(QNGY'OPJ<K&(HF'=$UO6@:F66";D&M%-==#EJO>#@8=DE@L\'\
P*#%,LLT/B.[V@P-XY<E>[+#R/0+E45D<2>E@;]_O]Z,/9D2=A:O^;P1COXG GU*!
P&+U1QYR!3P&SH8<SN]L)CM9"RL0'(HRTQX%O".X3/O-,(#M.<S,-3Z/X3)O%NF$X
P7[2O'RTW:?3;Y;&,*?!:1N,+0QV>VI+^</L"9!JVM'EQ7_!\]:7'DYGXA2/$OIV#
P_9 IHZ=_F"D^7CO/7OTJ=6[L'SWU9@[>&':F;/*'G8;VF=PG29KW"F.E\;*\%.TZ
P'H#8F5VTR*V=#D&M,[VA. 3#RO!:%H<@%>U9Q)=ZP)P#<=,@J5??<;! S#99BK J
P5(N!7OG347R\[K-/*B(>K>U%&Z$J?GWKV[C8PS+C8)#''>A%1#\2/9/>=Q) N\75
P74WL:CFX9SQ)U SSG]W& 4;?DU*XN'J5V:G73O&I]XW3@"'A#LF,@SF^0 :@K@3;
P^V#X*Y*"-8>A!^UHH"0&-0,VX@O49 S ?F=87-.UU2EX7V@5*OP)HY,\$M  8V;S
PMR\HO+.EH8/87'?,22<Z0AG%L!6NDO(-B$VA<QS70?U[*UFZO>4578\=4I_ SS=>
PX,)=H$9N&$R0\B5UU[;97B/'ZP%=%@@)35"\(5TI^^R'^'''R#-Q"YU27"!L@\T*
P@RO?I\V\JT0C<N.MV!E@^_0_LF.-X[]ZRQ=B,KIEG1-A=J54VAK$?N10>4*/J R$
PO4FW$B'OJHM.G+?]/36MI2?I[2N%J&C3S(E4W]4US$[9R3$DXTIXJAY487'>>&%(
P8D<S8P!B?_N:T8W[FP+,6SWVK!8U(/1F3TI9]-# EX3!>G.RQ0;+3BT ;ZAB?CQK
PKFFQ#ICJ3M$GZ)4VL*)ALOY+/R21(-#)(.[4ZM34ZUS7C"]]]Q[&A&^.T-9::X9<
P@AU24J#"A2NB^\0W7P,4DJH9.!;HAUVUH_1 ; Q<DB3N$Q"/;<-2V#MW%>&G[VH9
PX]5#7E4A6&"G$=R'3([Y9Y[0]\U[BA+4JKB)%]LNQ0<H>9-N7\:T@/V#1WS@15D2
P#DE_Z"?I1"ZVQ4.@ S"P]4[BO01!J1:^(_#%4Y$5&^J28\?2]_E[Y$!]6L4W[YN^
P0=>_%%:U<!(F[,*[P[J>KJH3)M!"S>Y\SU_[6?.42,2TCD4];1" ?_"_X7K%G$TT
P&S#9\H<2XW.,*F"D.+F9;9JV:.@5D+]I0VP3XM[ LQJU],3W.ZMIE&B,,^HJ2\UP
P%0!#TF3'OP%*>*&Q H\OZ)>6>T6E-ZV1F('NCZ +1WT$P;9P_1VY!'XRI);7\7.H
P@*;!KE?=@ @,_9L+WQ20169KQQW^K9*0J%Z?3+FN_NUE+E<5PH&3#.%<9"\(W6Q4
PY7+H4MJ[2FCA:U8AU'<6(A^=_5/P,VVE%DPB!32PV*KZ:CK8KB) ;:K98X%X*%LT
PWM6$8F@8<= *B(:<"ZH/X2JV\@==HRFK()Q"9O;?+10P1DM=Z--\\[ME*Z9?W#8W
PPH<F*QV3?B(=>U0+R)++?IPIQ:X+<-E>^)=2F)$Q?*4&?L1=;6,$&=]1( X/T??_
P(C(UF?4)T@&*F" 3(G5B;+(O,Y<=,/+]2(!_PQ&.>;/W$S>F<6;2#/9F9D,JH8DB
PFM8?));SY,\#Y=/H-"([,' ="[$^'9:QU^D9Y^/\^?K0D/S4XUPB@%;GG/<DN!0V
P'L?$O'%!M'Z32'2]14+\^4$07.K<8"5VE_2[,T)3[-4\"$K?SS"@[BZ[*U/KCY8"
PGWY6LQP;W+*Y/]+UZG=7;- V52;!PCR"@40I-76C>8T$J_Y>]W[9+%DD#ZV1FK2Z
PF)2XO7GCG@,V%9PD%-IKKTRQ;U#O\CH5P')50189L['(XEU#J7PJ+D@WY)B^XK?S
PF+L:ER2AKT"_LN5A)&U@(*''ZHA:KSS_!J;C/,I/:\>T*9Y8=P=R#M P[-0\("1U
P3+^CD4O-LD7F*IS;Q^>SGN<4JO.Q=="D@6(%W")X+^$\CFNUDZ/C,!3M3B.26W*>
P? XMB/9FW= "2AQM?Y&'9\Q77X8#)PN_QT%V!RK8C6]U1W!/6?V&CCX=1+:@GA.;
PDD>L5ZT(Q22O>FZ5%D'/N#O_I*2E"V0W\6?,3D&60;W5/-D2^)-E.YU1V_-VKMGG
P1OJ>G._JYC#ZJ_O-7&"ELQB0+^Y.1"HPK_G<O?*CIJB.BU_;:U1J,)8_>BMVTJ-B
P>?Y08 +;,1C^=ZCO)0Y2J;,;&JZQ^>S6G\J?KI\K-#ZSNPE^>OMK7"A%VW#6@(*N
PO^V2WNY4T_IIGG*>1K2S$*3ET#05M#&MS"[=FD412@;]GEDA?[>]_9K/-ZUT!"3F
P9SS $+YGU:+_'/Q_W!AUQDL+ RPAX7?,@MY!V1/D1I05F-M.>#1<I?RL[-P R)V1
PLRU 'B^\N X]\NVY5<51R7!N_8"&Y51HD,_9"S#GEO-X+9'A<F##9V"%=6H^D'^8
P?N@$[2?[[5\*4%NM2C-H5SMU>>E#K%RX\7KV+4)1Q9$O&E!EWH3'P8LS9*F6(0^?
PY,G)\ 892/,@5JU,(0:7E4$S[1&R6!L\08\XW8[;^\D&%C**B)FGZM[7"N2R#_X\
PWSJWVN_J)G]/ BZ%O7M(]^U? A;\AJ@NXGAG&RL$CTHV!XW5]KP[KY?(Q=>\FVK:
P,UP)Y1"P&1@P^BA5#<AWFO4^G=)#Q(8(X65._673!EI -B$^XMQ3AQ=]R&17.O/_
P>GFX O0?H)L-N&' 915C%_.QBH753CF\::)VY)H5I62W[&GK;BE+E_H>'@W\),T.
PU#/FX5WAH3E 7'MO6'YC[BZM"XLW=C#!;ZR&!'1DT2'](W6\@3R;SM7U="AB-5/$
P_+"XG],+U#<C TO&0EF2DE%;/K+=7)J\4RY.SR=*L9H*UDTV7:P]W(G<4*?BHUB%
P7MW>.4#!Q/"E3G&CA7CUF,_@4T?@/^O& 6+R62X3QNM*AO*H,5!\A'[ LO+N*3=2
PU3^FS1@ _PZW8E""&'R4&C7?,I4SY0]JX M0W5X-6AM)_#&*Y/Q@#LBJX[[*E,C+
P',O3L*"TDI^?5U%!TYPC++.-G#-\(&9Y+.S%OQC4I_/X?%QZFD)"TX5XT%+\X"AX
P\I>QU.UWM)0:7UO,TYH:@O##GP4<;S%,E&]N]\\?_Y0&W3-_I!5?!2&(" QJ5V_R
PW+:G]50=ZS]$9GPPC5'^T;<.6)D7YV#][[%,@M._^>#-X&^5LT\XE664H4A$6JEO
PZ6&0Y3N/P3\,X01&>U443L>JSMN'X:_S!\:FMB%LZU.D9_D LJ8>]X5TE_4Y)5#@
P76%EZ<,"= K7TDAW<F:?112N?(6 .%P RA"LAK)A@>I;JWEW^?]RTU8550C)"XM&
P)*I:KDH,R\17HY!W0S$2]#+*=N[7@@B8'LGLCP?0R2 1BDUFEEK@Y=B9C8OUKDIB
PD'>J5>/TMI>TI<"I4XB5RUE5A)9#WO\C'Z?MWVU)K5[!5$4@-^/BZUDDXRN'-R4I
P1$FH_"#1B\UL;PQ^,@,)!#6LI9A8\NQG8-Q1$L!ZJ_PTNQ21.JB)*:$NHASYF4T,
P>-M9&WY6 Y/1/C+O0D,1A_*2-VC0>K@5\@AJEE-<"NJ].6+@K<Y%J N!5E4@&NH,
PW8<6]:IL[/,P'Y0!KP%;>1NU(]'&)P=&GU(+1!WGBQ1R>PX.A_$[%<6CF8C#00-T
PC")?2+D4$7C/*G1F?TAP%USRLYS%AX87\/;V 7W6:)2J!MDYX9;>'+12 I-ML+"V
P=KVV?=_4XP2+9E^4L8S'EQ8H+UQP?6A1MT[5W6.Y["*?V9YC&EJRCNJ+ON*Y2:0N
PVNFQ?C0RD<'>%W@1#,L<]-#UO04I*M)&\=+4I9QE2;O#?)E5L;=XL89Y9*Y^7G%T
P?)R7HSHVF380INI& 0V'$&1E$G:P7MOL3DSI5TU@MP(]G[7%P8QLQZH#S(?-.#Q5
P[\][#W5:@0=O<C.@B!['E=G#$W%&!9:L1QM0D$I8U1V*>*0"J68-[T:=6M3*OZC1
PJ438XO!"]AY75RIQ;#(.0^*<;" M=!?"3H!^-C1A[%%<BF$ #Y9PULIU"XR-LCOK
PT]*+Q\U06&NMD+8-.7Q'KB4DER[:HDF=I<K46A'/<VV?W9SZ4&=+?/>),S+6]U"!
P92P?2=]$Y<$H;JMXMZ81>":B4:X3CY7E,&Z$5N^$,+KJ%*-+,!E5O,.5+A<I',RM
PF%!)&K+,L*0U* B?2,C[-MX9Q(TO<OJ*SVU23O2'QQOOXDV6@0QS\M W'Y$??4.G
P7J%G A;5CUJR@ZZ[&/UA*3,&XU>9/\[_F>H[7+^FSUOERLW2-'XC__YNM9_4^N)#
PC#L7(%TV 2T7, ?OVH#0+6E1G4PU>:'XBEC\L!_6)>&]:_DDB@[9SO8@T;2$9.]9
PJN6_:+ZM+[7I8\>)<) 9,]VO/&TCGUSQ.<NC!+2>=R=( 6-VE6/>..BB97=(J.I0
P.6L'IF^)1--4-MT68@]<HQ-,6J"QX491&O#*J*AO*=:F9IH'EF(8RJ.K(G&B0RV;
P1F<W=LAZP$8G, ,K+[9UQA+9,PB#YA=$)J0 P;.3T+MCQ(J_):94.%HWL,:.C@*>
P$GE556\E.'4@Y*T@-F*N:"E+]/9BZ4V&'QV&:Y8.=OEPZ/E*^-_1^Z#]#"5&SS7>
PN<7OY('*\O^[VX1@Q^8CD1PVM%;JXHA+J::R6&QC!*3,_PL[[H3> R;1JL*&$VD&
P4R-\F($QRS3X!4,[D%UL1IL%C0.)7&;4//8984\ ]0Z2$8:-;JVF+H4-W]4.@\E5
P_(<'3&GMZOEW';#M!*03F:H38T9:G[N[NSN9B/L\9PJR Q5WD/!@^NZF3'6'@FM[
P732 Z?L:RN%=T>G%\PB?+OEDN^)%@VV,<H',M] IY4U!'YE' HN(3FE<CM]Y_9%:
P7"9^"\]5F@1>9;U4K02!047,^_E3.4BL+[88LI/$7S=#1EX4:R0'N4U'+X>DT*'?
P:)BZL.N@EW+F7X05;I/N"[L/9?0CJ[MD8)3TJ:,HZD4G!E;,(DV<ZT?YK?>#*$DZ
P3K_C,IU/3!?8*N,>XS%0-4-G_3^^W6Q=OTDOEL\YD=@CQ^%QGMHWQFTDY%W%RB[>
PS2$Z8WK"M1@#LC^$MHCWT-7,\$N<W>+?E=5!$7T>%6Q4W$2XWR"GQ;/?8:U7W+CC
PT[[K!SL!RK<MMR&Q-/YBILS3'N$!R@*A"RDLVQ'B$"D1?.5SL':%3T-Y+PW7 \$]
PM%(_?%']]X,[CY;22QB<OKX1B-LRPY%S1.2P\O&? 5&>^0>P!&[6_K*"=CLJZQNG
P"/N<(#SO[<FKED85_7JF")HW#'H";SZPR=9(C>/R5_ A$O94"[A&@W\$U)>VJHO$
P(Y;:$D #7IQ\5:"CD[.LJ6\?3YX9;*N_+[AJH7X/)EU,[)[40/3,690$Q#@GDQFY
PK%>!RE=*""1S_V2Y&32+@+T]>EG(VK+!?4 6E>LJB[X9WQ+6L  J7U=KB4_GT9>J
P"F^617!WO#2KQ] &\]1/U__BC[2LF3(<Z,>,>42W, OR<440Y4,"-(D'#051EEYM
P:<)%L0TQ_',)'-XG?/YKT/G\C*F3K P$&P+,C\8Z1GY(%QA/>ZDLLE?:?60']&$2
PH/AH 7]O[TL[<6RC[B6L?-9VV4/!AEUJ^.\%8GK'EB+V'6< J8DB4?[YN<RWO^92
P\3+0*^'ZA[N[Z,, S.*KCE6AR)2,G?'O*U+,N":=3$X7,T>3^=6<N3H%V-W)X%>_
P&M5]+[I,#7L2/Y?JDHK#8<:/3>FMU.#"]OI5/S*XAI3-+_.Q*G,TQ 3-:ZA3&('3
P!X5F.KU*E:UW2WO6?E%T7_5M[N1_[.G1['MFBW8]W>Z2L3&AD]IW5'O:S"A"REE@
P<V*Z :(ZX MD+0.O^'!)!8GSL-RVV. G^7$Y=4C*HOF?1'^8M1?TK8Z: 6^^A@]3
PC(I8:1-AA% AUDE&_%0H#Z;22+JEANGG:O?$V<43EY^XO-TLG?_K?'TRC8%(3E";
P*%AIP7^32:-AQ4EF.-Z*[^"2&CY?8N7C]$X?L/3.;K__*-N8V;]B=CT\^OI"R=-%
PK/L;T\-_7^O^//@2%5X;I:\YXM"UXC1<;@T(4H5D0/IY*QYXOX[5S/!_0T\M49$X
PGH?GG^9)ERN6A-E^9L-Z<]Z_:=Q$>L?KL*US(V;,4.&\VC\^ZNTI;,LQ[P%?[X"C
P73NU/QIPSPT9R2I(R6L22E&<#H: EII=![7V2)U %I$OXHKUQ1_+04_Y"KPY>/3(
PJWT52I.HN0D7W4!Q"$#?M#T$ML<_U.WA;/V#'W<NJ+ .3U")Y>5# 8H?._^F2%6#
PR]2IX90$FWJD;".9$6UQBL @V>A8)^<6R"OO9/U:<Y$V8O+&J\J:NJO3](&O*]JH
PFN/*=U274"2-7\ 4)#2!8<XU9P2 ?75)W.:);*7GJ3*-X0*F2F4GA"4H=C_M?FMZ
PM5P5@Y,QM] N+)M.56N@>/0X<V<&D/5)7G-5<=M^MFDAZ.L9BMLP\P ON5@V[?L;
PI4$,$?E:QG26*43@9SLY2_!6+*+IAH2L=4.%_>B,C&LH_Y-B0M8T+VN[R+S31)@0
P!<IT2TS<QQ:LR$4TUC=$^W4UN[J2\T8L^9_#^3F1(#+'=YXGB8*80:(%Q.D=?Z/_
P.6S'>(.W9DKH6N=@7P@80US9SH(Y2LC.+]ILO8"X1IJ@J_<$Y"<$6-8=!1#7L!#_
P!K)=MFJSZR$-+M(0\RX7Q2E+YABRUI-8QV*9&/+QR$OQH]O\J1"78 RGLYK<T+%T
PB7_]"+F$105J&FDNH[M^P6*^M-CR]1Y,ZAF]F,R>'9PE4C2_I$V6)GD!49-_SO\W
PBA_K)J4-8729$/S&9 \[=#K0AQR]1O>@!:*J)V2,WXQD%5_0WKKIDTH--9?L,O,W
P<;]&&EN3EC^D3R708K[8MAJ5P-]0+5/"'LG>^O+ZFBVQ40.;"03B1:6-?#%NT+BA
P[)H*6VC$2P6DYQ]R! 6 @9=> VV#I5C3UKF,.NB6'0MT\\;E??[[^3!0ZY]&@"54
PD"G577R!:T0!AK=H@ WR.Q[#PNP] 05R,%=/]4@Q4S'7];.^WE9H\#BR[1JN$;KV
P<DAC$O?[5V00*-8MC4;+]1(,;*+@8RAL024TW?H![FB01?HEK66C0XQ\E-W"]'!H
P8;U<KTPL2,,"Z'TO9(L FTY8Q4JC\-P\/MW\]]T'&L3CIZ&OBP=7;%66U&5''PK"
PKXXLF3RH&#0S@S_">4,_#FM^5:C?M0(S_CLZSX'G]XG=T%.C:C4-"<K6I3)VQE_]
PP*-9T;(HQ F,NT:FBVG_+G?/@^K62UW28%HNL@C&;5P8,,<+N+4G<N;2M->H!;?G
P%VXUPQ?J?8=2ZXL=TGCH,!N%_+L/Q?AH\&DB4$3*=YG9\"0U@\'TM21YZR.1]A3:
P(AW[IFU9M-5]Y'OWB8J0T#L[,*$I<&CVR*R3(J2#ANOUKT;N<,NCK=+,QJX^#MB:
PC[UB^>&IK)+SNX[?'-<"<L@7> U 3LQ75GE'9#VNZV<^Q3O_B8.S&[!CNNW;ZB$U
PI(MY6E/_*S?_7^E<+G#^U_*R+-<V6=[C\EZSFS3TXYHO.0N[+N#US&8#0*CAW\YD
PX0RRS1NE/9.;^-R3X/;I5YI8"X^\'!\)Z2=%#PX5U+S27\@(4';C'*A55+PER 8A
P%B]!B6\'WTE:B6L@ID\0]-! 7>&-=>H-Y?MM0'PF&<84MB9;\9OQ:*G*:*K:>[LD
P_H$$?V%M0X/W5-1X(Q^I#YE,N:,KV_IAVYYC.%BW(H.3.[4VTS0I@E^'Q B,DH2]
P]C3B> 2#!)^]+6N3<.RR/HX9-FV/6SOS;0;\/DW8('6$0%D]T5D2KJ Z!G?)]U.&
P8Y+F-QW<AM\2&-2?=4ZO6WRP"[DN1A@YG/=%S#>E4"AO!#$4OE8>&!/HO^)O1SMX
P-^QM "1< !_>U$DA92^HDTSC@\N3/\DI >6H/Q%H88G>36\XL=B_3>^RI ,4(#EG
P82]>_BU*'EP6&S8%BK<Y]]DP+!#BN,U-(I>SM?-6&'.:6UN JV[:1W3 Y8*>L)S3
P3IS9JV4F;@I,+E336G3[%,I!4;LE!8H$!)P1PZ'OV#X#^:7''%:@Y5@3*U)QFZK.
PO\'?X-,V@5UO7;ADNFIASF4-9YS[!M,41BS,G_Q!2@ F]\O;BI$SFMSZ%6=:/ZQ:
P[QL<'"W\5R,84W90^-T*6%,'A8;;:.%(H)=3<6B,"R+FJO=QMD@#,0&9<@3/P?+V
PTML6RZ[^ZDBYYNT[)KN:[->\GT!AV8EXCO#;#:\)EU1]T;L93)<2\[/@X'K]+0IV
PNW5&&WGV598%G\9H U(BR8_#Q%.'&CAFG*+-)_S#WG++#PNA:S/7?I-AYH,$]W?O
PQ^$/\JA7FS?5JR/SOJ=A-;H[0N$2?*PW?\>Q%;D)@3R$N=,X;'*F21#Y=WF7";'L
PDL&7P[>X[$U<!.+*(&^"^B>0I_&G4;:"6M]3OE/]*D6BFR&]5TN"(='>)(\#UJG!
P;GQ+KR2CLI0!F!^VX(\JWYO+^6#47XK(?(B.<NNC^-8<YPN<1_MW5^5X)%WY/,N$
PP$&73$!6J0)ODUA@K*.Q%:CH4@M/+DY.@Y-^53;C%:U%;3J%)L=\1'$0KR8.8@14
P&S'*>TOVMA@/Q%O;VC2 0PB[-2>S"@@,'IY1!D4$'YGNI<C(56:''X++:<94*;.A
P1$[BE\N?FIS!DRV%?*A!7$T=R%$/_T%MDT@4E"IR@)M'CZ*<^4S]VF!1/A3+P\:K
PHU?,V>TXV$T (.> XX--RX'DE%;@+\KG:)J5U'K",W8+KIL/2T0X-C-@3XQ"K].'
P75O'7OG:F@/*QZ*Y3L)7&MU5C/$_AM1WSG*3RE%8_J<V+:=^7R\_/-;3U!R49^RL
P$&_ZK8O?,L,RBR.:%Q$(E4%[I6=(Y:JFAT>><"=SFJQ"#W%UYU4[5=E%[=RIECOS
P !6Q!VD4T-5I)[_VF>'Q&I.QZ*-(#&SM#=A[#7<\#]+$V[?2ZWN?S7YZ?H#&,O":
P*0CCK/F/_N3*K* >_+60* ,/+M UD-0W3$:7)%2A;9#1E4)M1HVXTAGI ZQQ+_?5
P01/4>3:IS*PL&T9R?G3- 9TQ&Z^^]<67O)+<+82V+;_=:;P'/MJM/+^MT5QD9\^>
PY. N_=06O99RD@'<X>\'<JQ(?0)&4?V"0R.?C#D?IQ/5V$U<DE>AED]X*,HO,U0T
PTJ[<MFJ[_LNFX2[,(+[-4Y7LI*55PF:(#U"=7&?443:&&/'WOTP&0S4 A*]1>&:\
PV):()07-.@#CA)Y=/BW80[RKBF +2+Y_BY"0J&#_. 0A&5J0?"J(;0>TG;8WG$&X
PGE;E4S 5I%M/@0"(Q3&.HWX)T:83;)(M-YFB5.V&@G1"Y[PUC;D\TD!"LUJ%@D'H
P;8TW]>1:^3[I\'\W1N9Q,90.$=]%=!B61'V:]H J>UD%KEW[1<VYA49J*S&#E*#5
P"I+<)M*I1W4YJ@33YF5]L$=AI^3A*(&I8,7#80CZJS_Q99$#&:>*(5B$Y) ;N?%.
PXV[S%Z;OQK\[FZL7S"4I#[E&.!#"45;$HU0;3N/1<@Q1\*]-TT-+0*G<X<L*KRR8
PEC[C0K\U]9T(77_'^:(/6&B;U(Y'LWP#X=]@9>47N\$'SB+([.PMA7]AG$:C@QA>
PYHC/M1<"LF\XR.A^^'8$P)9DEDH9_7<6L';V@UC@%Z.71[0DBHU$=8,66G-_UBL,
PO&(G:^SJOG3UD:QIJ=_:V3850;5)P<Z='BVLP^[9JS1+-O9T(BP-UP%DDY9VEYVK
P&1/MEUK7DL@LLK1/4WE9^4U1N4V\.9!P-/E!A^R!"[A[N2>.<\K\'?'1'&9C#EXK
PX.-37JL,4)9.,H-5Y8JL$CCN98!-*;$I]C)8\3XE#=-A%,W<$4LSNF-Z[W49D('Z
PT^B@]E,BCGFDD#)S_[,'>;#P-^1HJ2+2X6_-IN<=R(YZ0*=(3MS)J$/,F/2]NV;"
P\@Y803\)V!W9Z=[D7T_[AA$[G\6[)4$)VR))0\DVIX;NC45J[Q2XMN0LFC]V>4W+
PK'_%2D/% ,B/K'&.3WJ61GN/V1KZY:BI/CFV6 ]W<UQJ%D?R@1"D&&76^].4\,+A
P:Z,$TRGG!62I#G\PTH%0^+$9XM4*+7523H36@50EC<+]UPJ7]Z=[XH\<82YR-+&M
PYOEH>NMBI/CQ==' 4QFKJDWJ?BNH8F@/Q*V6[I!3/;SA=Q5DQ=0H3>"CIE&&<#2'
P?8GD7*L+:33Q<T&I2E2 ")%+4I3!V=B* 7%(3X(#=^DC3X97?)K6A2)0:Q.VZI_.
P;P18-OG+T+5EUD*+* VOL+;[-#O,01G4D]7Y8DY?]P#=%Q;4,%XFB?47Q03M$-JJ
P5(OGA= $.>6QX=2W(4-#\[>;PZD.%+QSOJBP1H52#52#+LTV:A^5B&Y0NQP K590
PVNNU)(8!8GV4O$1ZY1>XI+\J^; ?]8,U$<<&&[=01V5N."M@6P+%!HWO?&?1@SRK
PD:PNZWT]V\2<K'GAHYSM*HS/F94I4 O*$5@X_EU.YTQ?=_(%LKU87M8 J^C<ID/E
P^" H$F]O,($V+O-K4,"%[KA+0:&;U"B]PG08,DX6C].L""JMI@F8$0AVO2ESFT6%
P=5814= %V:MY\)>>LH^_C!QGMD]I?#%,#L802O,]4IE@/.ZYGDF?D-:/_DPMNF *
PYD17!%KV9KR 53_.'#*W'I(:(#JP OI1YXX[JQR8:50\R#C5 OFJ_&>%L4?CO:4F
P2^I;Y=-*H)6#3&<7-=2;KR-3A,EC31J!J]8RGF-QN1N\0]R]7$J]'>?8',H5TVK'
P<P-)F-M'KE-@/7\;AON4]N@12/,L^+Y<&&#4":XR&NQK>H ]71U;Z4(B3C-P+XZO
PM)/= _Y8JW[++KQ[3QB/V^=-\I.\T1:&]?)5<Y$OO@$&CGC0:B+E^TJ8G'47VIEZ
P-J*))CD$7\T:7@U7UD[#W;JM.F$8LSUX-!H5I9XSN^G_&F7+]X\VLX2^[K1!$&$F
P)I;9B[J*^\_OJ#'&XR^7>O)[7=  XA1HTN7U[86'0[4NB+TK[[(7=^'?C#]G=#GR
P*(OKZ;*GNHU9>Q&"@*^ZRJ.^7;1A;M&!)6+*\5ALF%5Y/%?3:PL 3DGG+;&G7&KJ
P[E&.PB\T(VBP=KQ(\5*O7 )RE>&/XY5DF44K?^*[(E%+R*UI*@V,_#<*VJ[;^J]@
P8+?MTU]  VDD"YZY28G&"?%?T:*[>Z<'B:+;EBQYSP]G-N=?PPY=!J4@ISI.7Q<F
P_+F?CBFFT_&J'47]IZ[?CGK22]=J9$BGH+$Z,0& PD=LH.\H$?,L"#S?L,':TX+#
PILE-QE[TOX(=5^I'1*DLGT.87, "2-G:U^BK9W6(N>)XRBZ(8+.VUU^K]]27RMU2
P'+0=[#MC5(]U\8+0WD%&80P NK.DYW4_8*0&%>-%:''(1'F^.]W\6 I(F!DK 81.
P*<'J!=*@Z#,3RA IE]<2$3ZNC\/U6-] DF.A90G1%;ZZ&LVH.6NR <U3G<BUI14$
PSZ"JL,T4V#=?$:5].+[B(M8X3SAL<OYV%SGL"P*N4T=O%  )H>U2<\X,'*Y^+%N>
P)" >CI 0[GZZV6#%#JX'U]A+3-[S9O2%QS'X</)P9 !\'GE+CK<7%'=4?G[.%*,;
P&SF&'ID^\BYQIW3ZSCLH/\&^O8>& >D*R[@%>K>%1R QQ2'IY(KP6M%OH#%?.MI[
P0Y?ZHZJDX7/ZN4(:V?C)1$]1R;"6X&/C[[XKNRG(9!YF<D_L*G>M(N$FHLKH\C\#
P[R6"?C2?QD#S6Y75+8LD?7*[.UC! :YU_*-1(I6F4M?*M@,JZF#Z,?LP! !CQW/Y
P1DH5""P1\F7-LYHSM(1.S"P=.BX' (Q!>2%_P^&B:+/$;-6?,)$@A9:]2I$3/XU>
P^'=-O@'6[U*UE=U-&':)>9'AE%>J0!7:#]JS%Q;Y"X(+>Y6J'>R53;<[DBKW(%:S
PQ78690)_X<8\OU-D6;#!3%+1!/5RFY"MCT4)H9M2HB-JD>"L[F"A66A@8*JC*T5S
P&[4ZD"_!J7$,@DA2[/@P().)/4X@"IZ 187ZB_0N@??T1>&1+)8K[-4&>MA@:*2H
PT%#^,W;=\+#1GW:-CTH7*"9.NERE9D>;TMR#OO(:$?Y2?9FMUD4<0LI55Q64L6^&
P5-^#V%<+R+.5\B_+4M>2KX,3U(Z:@-O[[X93V4,28"P2X<\*Q<V/H.5\/*::= X<
P5IXOI'7\X];:P#NUSR +G9FFQ3S,5MB_C&[$=6I*"06^G^9:^^IKP;A$1\.RUM=%
PRS=U*J[GN/;X)$I:2O7E"X[AC;Y"VZ'VQ7N5K70]RK[A SN_E:T%3/J!7^U?ERMX
P# Q#4'Q@^+<7.X"OS2(.&F\*X-Z6K^39Y> @5AXUA>@W:ID3>.E6RMYS]_:736$F
P>AD9<<RH[NP]S_[9G.0EMNTL?R8F4:Y6_>O2D58AU"?>^TS*VI1IH1IB7WB,SE3V
P<6E/M23-1L:['E7 #TX[E*B?DFQHC#WZ[ ;?Z9-.B16.!MIT9925F@L!6E'>UB",
P$JB1P7='!WL<82#5;P9GTD\3H,X3$,_*[!#O<H2*XX2[Z4)5/>]7CV\S'>Q2\ ,(
P_ 5D$\W'IQZ0FZQ!6+R"B)"N*@] L]G$O\XV%KLS N_GB_&"GY5EJ=L1(X7QWM+0
PY&)/&6CGS9M:E7F!0%YLGW1^R;NSS3,([5#D ;Y C+EB/=H9C4^26T$ZOQQLLM]3
P<?6>.,>@:G&$OE";FX<(\Y LV@7K%6H.D_-H<(+L_C8QC'#:IJ&F740K!]+&V74\
P,8Z[^RD@:)%'VMHJ<[45J;V4#[+3<TWE1D)O>RO_4= &3VB,;6]>QUD7HS. 47)C
P7F]T3WS?9XW#@=J&]0XH-AB1CL]+A<.!EYPXTX[2T'=G1R>[@>=5\8A:"-W[5 -#
P699:0\^H#F7V4A+VL_Y$8R-I>,[C*(UNFPCBKA S&:0(#\9SGT/&9>O]8?39,'%+
PL5F\Y97CQ*C,/!P/ TM+X3_*](Z&:_!N31W,:Z'ECO](,@YU>:0H&(JFR$$R+L38
P1S]WJ9GH[<>F?H%9;%DF+^BI4E J(%0?',N:H[6QX,?'MWQD(Q2U2X7U?5\_Q_'Y
PZ_0/,!(M9J2\C]"^!*.,$]YFJ].ZC)1MM*:MOV2#[[#^79HV: U_6>UK\]F0O0<Y
P]J'+ZY6.I?"@95X?P:V9- E.U@P 7+H-TT,XB;-(2<IPWN%HX-F/AA@@($$Q8ONI
PZ=PEN1[ @M9Q6]@7G'B:']Q6H!68@E3UD8Y)?+KQ0#*UNB^K[WQ<G=<##ZM^4: ?
PQUE/0@FD';+ V[GIDF)WDX.$9_14R!0Q@$'%G!GL^A*.\Q[>/3Q5HAM0 @"HBL2B
P'8@TP@O>"Y57C!GP##0PAFPMHT^2J9Z1\3Q]DNBHLK$FM7M0R.5WD,$HX[)=]SZ"
P]Z,PQ]UB^#)T:_JR'A5H.P",!4U4&Y_OZ6KFA8G&NDH0PG/XJ2A9!YUF[$B'AY7(
P#-M%Z&?MF9^1&>^:92-JIC%/#ILF)6749(N;<(\HQ'OQ[5@S)S1/MF.!?)TAZS2&
PC9;-.:LDQNDK(BH^$'Q(;!DV)=++)Q/!"&0VIF<Q O)/4QP1S[Z6?XLBL#J\D7-/
PW(1LM=\O*BUBY9!ZP$ZGO!=I C/\1B\X^\HRBJGQ?<FK4\U'M^!A57^[L\D>[>^J
PHL.BZ#?9O/T!SA?S@P'[IA)C<%N.;$QH%*JGM@QL=@0NKJ-)! TEWGK&#@I!K"=+
P=01O^3U&5FK+_NLQ:_$_6*A?UB^R<3ISS[^7-P#/LK4U*TZK:OKX%H>0]>DS1I"$
PW_^*OX&ZMRG5^H^CAV$'YSL]K?:+:SWM2D7B*:'5B,QC?X^/IP@J4/H]*W185T<H
P:5GMLXG;.VIS\:CLF[& B9S)+=A*CJI$)$=%\4MA9"W65=[5E]-Q1E4SD7,:X#S5
PLIP.AA@ ("3SY@\;G&%2]CKA6YX=@]ZB\[DPM^J16UJ(%:K$NV!P+FEVMV/CX4BN
P@6QEY9A7 IP>%"VK16QP\-%*,1[,E8+"QI&GB18I(7\[OC\4>%"/-*CUG/J[/(T;
P\^JV1;]'D<]+2$72_1PMIGU!^MP7W#3A)4V6Z_F%*LG3B$>9P.PO@1</'X0?3_9%
PU<[Z7:9E\T_A-NTR_E^1Q47%$C3T61:3GF1239>2('UM$+G>\\/WKP7+%RQHWW._
P.K/R8>3+]^04[VQZ,W$EF,DHXC 1F-!]6RN M4I$&70V5_M38NV5*@;G>)^!E)_.
P&R)\=#;D2=H';==6?[]5LB&:SI]JT7D4)(Q]3X+O^0Z(W^E* &E.+= 8O,<G9)=)
P<[K):IOO$'R%:6^QE3TJQI*C7E&8G-LP&TZ!L]T7!_:K!K+\]#"M04?SH3;D/]F]
PYQJ/!&\_E&3ASRM$73WXJ!23P&*<X3O4_XGG>)S3GC>-QT'-TX(D0J0HSQTLAO-;
PZ%%-[+L96RTIY#F^N(1+>B5\6V@AHOE)]__)]E(BG5J\Z!Q]RVE28^0^*W8@LY\%
P,=TP)R?>ZG:-O+VQ>'&5\C70OWRCTSVV0N/\DG]*5:PP1"D^/("I'O3;\OZQMWFC
PTRKK0&Z^LF_IKT 5. F35"=6L44J_V_5VMG5$"TZ7L;3^*Q9O<OH_T4)]FE R,,S
P4WP[I<OI(5Z-=O?:H+N8,,HM.AJ&PZW36/8@KO<5[-*V,>\]YD.'AIH[XBW"Q3(K
P(,#?L6] X9KQ@UXN(1PH'4&-,E](@8VQ6*P+6A>4#F*E/RDWX F36S)B'\G+41M]
PSL'9/>>&N=P":MOX_G]*,%*]=E@.* $%']Q!6 J[)2V";Q(M_@ZW1JQ#'_BI;#L"
PJ_ENWEZ*0[[092MM:F-3>A?EB[:E?,2NG-_H>2&[TCS)VJX17B!'2DW^C)BHB@"W
PA9FAWUGW;?N!_/JYXK=HZ;1/50$I3ZH2-#+L+_##_]P7>.,S' ="W)G*8C,$M*;0
P)]MH6HP[4KF4X8:8$6AC"BT$$QT;%HDD>QY^2"!#3^:&+&R.7 C:)/,>35@!- Y1
PA/$BWB+)S9"LOL'KUE)2,]Q#'<YKS&;-ANP9Y@LE%3>6<$5MROP2I ,AE>N*G-]!
P:;2)(](4MID9: /]GN^17A(MD2<\WA#XGRX4QUD5@1W$^6C,L)>O?/UN'VKTM;*)
PD2N-L+5)7]VF"7AH\[Q^ ZLN7H*WT@X*>!^Q^,BNGVI(7/(W' &DFY0[-1?K!^/'
P]7,X\CA_CT&EI)<EM<N(T[\",O?\R@'.@_[_!7E,D]GD:O08$9JBYV\:J6@4)D22
P/1O6(W#JF2&CCZ3Z_8Z%G&;_3WM/G9)*QZ@H(Y%*;OL#0(G6NQCF+6,;U#I7-/ =
P5:R0V!6F:C/SU^B"R#-'GW([1$QF-B/9AY2J]V8B!GZB5)P/'SRW\Z2"AS,8F\9 
PJ,2G'*/X1OQ]-7P1O>Z;K77J?]D=Z_,!X!WB?+(-Q/LI#][H"['JSZJ/!'^BLFMC
PBID@KSFMV@_NPZYTJ@]DMSCD)\6Q]:GIK^D^^VRG"*_JE,&4,)$GK;L8Z%O@2$& 
P'#5<G$NIM<N\(^2XPWY2QIIMYHB:"C6>PF0-%$+0OU U10(1B0 3.VF][1RI[/^0
P@SU2/MK5U9=J6R7U,EIYVK#+J0C>YG(%A:C6#G 5@F]\_2,I+10=CG>W<Z\C0=KM
PNB"_0VP$)8C0WA2=U3X"J:?5!NJ#48\M)2#8=I9P+<_B B:(5%^T>8AQF1RA(D:U
P)?!#$TL"^M/X*SAV%&6UV\O#BMS:8*GC>D&+]$:"2<5'#*6'PKX[0*Q!ZC?69B]&
P\+[IOB&CU$8][D#,62'8>BUV EOU+=TUF^+6-8AQ]HY0D BCQ/+5_:UMN!FOLV\N
P"BP7Z#-^JLB3[?>CR5@0";FM8G!'1Y=!<#^4):R'E=8^)D>M ,R5(H#6&@&3NU\_
P%O!?IR@*9ECWRK;3%8B!*MOF?K8T<&6<24DIH<8!R[N?":T_7TO[4T@2#:Z$';1.
PVX^,SIB#8A;E*Z]'H7%\W6[G@U@:'"-[R8V=H0;Q60T6A)*T;O!-\ "6N^A=DKT,
PGM !%F;?F_7HPM/;R>4-GH:=*P%%.@'FS+XKHT2_['O&I\"0_VJ>(Z_RKX;B&,54
PO MZ;MS^@U$#N-?7<]''<F3WF1\]*X?>'/K"( TGPJ?QO54.(H7?J7T,!S^Q1VD8
P>91#.S1?JAS--ABU"P#53O3H@=]G#"1FCJ"%0)<&L0-$1ZAP(&.9V B!4CCP;HN7
P,H<%$%#4W&"6X0A%<U#'APU">C*(HXV KJ&PU$%K_"Z_9:^E20?0T8^G7(.Z; $(
P6'GV^**^IU?M)P]R,C>,UM8F*'N5Z8"'_ [DCEN$OE1VU5S_#R.L!^"X,9!Q^T^(
P$$J,0S7+>^L2[\8PYX3H;9KL^;OJ"^)5>L=A<8\%K=$YWM<?B\@"_3DJ)#H[)PD^
P;@Z^1(^^, Q%1 ":O8TB29<4MG*_@86V?85 :?U-8TQR1,N =(@_)E:QB0>+W&1M
PT7W>[S5ED128N0H 8#V&VM:P':Z-1'A%H;D00+-%I/6OU*RN5,@5M%>4@5]1,J'(
P&FKP>IS*U8=>J))L9P78H[I%T\*?T-R2]^<RMR6.RCO%<>D]W69PP>_Y1%X(;A8Z
P)&/\BP@$YQ@07749.G/2=E(]M:TPX6<'H0[6I['?.$[IZ-+#*39)L 5$;C-/3]1!
P#=50?<HS N.6H!,]*A=X]NY <NA7A^D(!W8M -+3,MYX&'9J,T5,\B@0*[XMUR)U
P)B62-# ]ZK2('7\GE*359Z9)K&8J1"-)F9E)4D?["T-,[M9OWXI5!@-4PWK=09A)
P2)O^4P\%9C?:*%KBBYNF06WC+"Y9M=X9RZ4X9*(*;AYJ6I_].S?3:?8IA:*8_1W&
P4&9$GS#G7 ^*#KZ.FW9\<32[L[-ZR?@[>L#P.:3DV#400&(C'N=[V;>^!*ULGP^-
P8#L0%Q6L2U8U"/-!KRS]$*[KAF0W=R,MU.#/'M/-Z6>L'*E54,'E"2&Y+%]1:TH6
PSW"&73,E4[,>#R);UK&R%!^9R]5_J@02.=<TL^PV4";>R.22@365G!&'%FK55!J2
PC&4Y/G4]%FQQM =EM;WLPQ'9<5&&>!4#IQ0^*Y&%?B)V= WWJ%X V,OM1HBGM'^2
P0E]M0HKL]\A!<#-N41*8__X@X0;#&<=1RH#Y">^9[LL@!]E872^30: F0]4 XJ"P
P#LQ=/<>NK*)&EK!=_5QMX)6B>9.H;>.D9VC'29=0"1+@UA>O,:.%T3KE4NP./N;W
PLNL'WR'._R]X@(6*!4WYI @T$W2K\G3/=F,!=DU8/Z6^,N_OF.5>C -R.G^P"WW:
PS$DG"Q(\^;X-%-D7EU\RA2Z98U04N9E_28_STNQ]G'=LG_6#J,I9NIM9+(!4% 1@
P5NB(\;Q?B_580;.SFMXS#P#=#G=!^5>1)M-"O @*&E%7T((LL@' UA/4S>G<HQ,\
P'QN<.HT_[?#0/(&GS=-RLS)(_GA2A(6. _O7Y&+ZN0I=E.LO7::/WNX,XV,P]:6Z
P/=40TOYE?(.?HU<E'W$@AY"OJT(9%55-8#,TWX8PH@9R:_(ALR9QI5>V81NF6=;S
PEX[2/T!!*F;9,RI.0RCB0/*JV 9IX)M#.*RZ'[+P:Z<M/"0_&X(LG,%KACIVH]LL
P6TU$J#Z(E88VLT!WX\_,J:WNU>N6@MSTD.NWN>T86!%,B-SB[](/ DQ@,RTH,7J!
PW_P:AO.L P?F&'RI%IEOE93OKAK]5WH(FA<D*8MZ(TR$D??G/&YT[##GUQ9R$[.*
P5BPH0T3J<>#Z@%H3_\+.S\%A;.<Z-=D3GM_Z#&C:A>A,C4&<S+M3&-5Y5$[!,>H'
P(ORIGBA#4_R>SUT$@/APY9MSO_9ST8_JUJ))J!)[EOK@X?D.WF]'&D7%61FG9O(5
P74'C*"]@EON1.8)B'D6RS$KB@3'>AKQ>TD:= CZ]4+9N@8^.D5I[S4':\M.=L&EU
P:EZG]MZJ77L M1Q[[69=]#$RELTT1G==1F^'?_+'_E_ YN$N/+EH=R5R='53@M^+
P,5U)@3[[-9NF_FAS3?8ZOY->>^M!$F7,KR'_2:I5F.-!/]HA>+GFB_<B9^ES%B]*
P2J-M1Q$_%GS*3\.+PNA'UC(:FH([;A80I]#CE#52"57R"05FJJ(>&T^$3SLJG8+Z
P*<)2YM)Z0AP B%%F0?UUWHZ4%4Q_8^_N^+/2O\.'*1R._]4YBAZY9JW>B93 MR@>
PD!!!C9#0KE2(7,-6S^)STPUO:Z@:!K0/@XZK?Q-^2;]RN =L%4H=[>]^-+4B[\[7
P[G*32^W:\DO#"_ZI#[>&56_@&D=KSGS";.UDF=N&'"_7@JG>"Y0#1>[1R%A1+4R'
PK,@]NL925GO3\T3,&/9O24^ .3XKBJ$IYJA*9@)OE0@79#<Q29CSB-!( F[2R\MT
P+  2%AGKM:@4SC]II+I-4/3]+B PRP>2XV1F[WT"$X8>%K,_^,X;?]P6R:P< 05X
P.]85%"OM[+J0908.(4A+ZF4]3;(+E:\D].O,"@Q-[@)2PJ&_P&/ .TYY+.UE%X<(
P^'=43E9_BJ=W,T&$BYK[<49R CXC@DM51$0H.8WR3EQ@LJRU4FVQG#MP4PH)._YV
P1-/O;YA2VFIPC-H)PE/?+R7!H24.YF*.P_7NDQ=DWHZ)NJV5$!V\ZRS^>$I9/'0Q
P:$."U/X<0CBD8T[+2.[WQW.F?#$O5S."_"I"T;=EW\3]]G-@WIBNN*#7'*XZ0S"+
PG!.<60&79Z(A_3'4<(ASQ\&K='XS+N62*4?1H Z+LQEITX"'@V)L)VJ ]%X_DDM&
P'&=[(FR,3URTLV)'0K8<8NQ%XI#+!@:A:NTD7Y0IPH3_I; 50JHGN!YE>A?FN2Q.
P'7PB@@J35A>B?RTNY'UVXMM/$YW[8<?RY$^V1?++M"@85(P2+@DWPE'%56\U!3@+
PM [B:KUX3,'IO=2XOC^?&+(I=^)4L=&8Z=A*-H(_C&!BW_ON8T4,X;6!8XURF-&2
PW4XJ<5\K:VZ7F&,14EV(:K4F\>WP6.5!J.@K/2ZQJY]LJ:@[(898?9>*'6J=(:2C
POO[/[R_0XR8\#)Y#"BV]1%&](V'ULPV8$3=N?[@5_U#D@7R?75Y0)TM'U>$&^.4#
P&R J:B# +TI'Y*"]+S;S[ 9!#858=J&4B>N3AY8H.C^0$2&=BSP&,J%0I",W[J7,
PKL!$)2?@ B!\;KG[5ZT%38P+">(B*)7$*0#*K],P>__&SP(LSGS[1QBMY&UXNB)W
P0ZVW!QU+A3U_3+JNSC( Z73.[PY-K[:R"AD7VMRLJ:Q83R,P$RT,QQX <J'1VH;,
P"7!"\S]*$'Y/H]O=R%@U3$R(UU[9GN"[J,P*JR.3"1G=WGY6/5/);^PV.?;PB>-*
P'<X@.]T#":]V#R313=ULW3U\C6-9^Z5EX?B>"4J!WIJ&SW?8ZK-,?R\XB-()6W/^
P+9U$'=\?:U'5%UJ&/'/"B2$,1'V@3(I?N9]:UWH) )]L[:P.38//',TW!E -"L0!
P_7^$$9HY0C7-E,>%UD,:R\9%_])*.:7A\+M;LXG4\B/A[V'UL%62=<^[7'S^Y,;M
PZB#"LE5,U4(:G2J&E*F?-8(=B4.5GDU-&$3MJMVN2]&YK$+RGAG?Z/1MKA<MPMGN
PM#CD%]3DL#@M3A+^$ (%0P+-,<+ 5*SI(;(/B)]0C5X<$P=8AA&-U@ODD'IJS7HQ
P#)ZU,E4/)0D(20N] "CLX6K;'>/ X/T68)#^Z;AX^3(X^($][\$#1M3]-$TM27;:
PZ Q,<#RW04BOM]HIQ0/RDD"@MYUM=MS]-'D%.N"R<^"=@N&^S<(X:BI<"C9GN?[+
PS1/NH0IC^*M-P ^T#WCD8#PJ1_54P?*#GA&7>!G.PH;B'T(L5&V>AWX]# ",F>%H
PV($LGT'-V[%#N(S>G=%( 04XS8,=&5UHX0MPRW37M+R;]<%>L+1XLTS"]CBK_K:&
P]Z05/7&>-HB3ZF.WCC) V(_B,X0.T9/*4^YU+]SQG4F)R(^FKE&GGVKWB !7[NEO
P93IO_1K>^(5J)0[WFX3R[BL'^',398XX:.$:@L8O_BKFCU!WDSP3&I_L7A[R7[3W
P]T13\'*V^QQY&7VE=O\R5+F@.$TQBO5JRP!=J$D4MCL$1!QD&MD=],(9B]3&ZKXF
P;OZYZ/BPZ(R7<?T:]B[>Y+)_O2 !;D&60)%N^IK,ZGF37'87QWOV:(6V/.>$>$2'
P5NB>=%I%&7'#:W[0>6?4_M1(EG<"C;;GR,HG)H-Z:57SF$MRS]+?E("JF@VE%'':
P]W1Y?WHPG4N7!WRX_"8<>Q!L,'6*%#";]T0.6%%][%*U)Z;-&\7'_/DG%8:MA/[:
PA,NU<K*23K<2^S09[(C*'5OI>S:GG'EA++1X=PP5GF=VW3/>]@P&R^6PQ.5PU[=J
P15:^P3':; 0[:3Z, 05 LKO5"-W/2++);QMUU&D5FBXP5@>VOM2\!AK9-+6=]LW-
PX%^VA)X@,II/-LTM.+0UY$ OM<"* :+4Z9'6@*VD*H271=A*ENF]RNS\#2J;?)"Y
PV@_.Z%5ARA+7%\7KQ#Q]TDOZ=Y;Q\$,6%U;&>LL$!7(MV'F.QF^A62XX^X6$R67M
PMP3B!+VV$/J>,03H-A@!2]3I.EI+PGY8:/F#Y&-%#<:0&/>16AW3O"L/?ZJOY2^_
P7ZR8O6Q%E(4K^K2RLR^_K$@T&EM2/___;BN'K<T8AISYL3LUKMC6X_%:]Q8<A7VD
PS?7VF[FX\S\LK%)!$%HB C6VFGQ*=8YY59 48VJ)R"VHS#J&?9)-8I?0"PLT$@L7
P*J)1#:U^(01^2MN>>P\6SQ>NO1!!>*>NX.35ZG.Z :\"R] (R-2E->)4.$=;?H+$
P Y+X/&UX5]T3X@@OJ"=Z\I?]C-,5*]LO=YEH]DRL%K5-MT,%;"EVYX8_W:\:/_#X
P%UXYP,S5E0Z39CNJ!*J:@;,.(=NW^9& !:Y =>GZQV*XX?V\KBH]%;"I$F#AD7%5
P'H-&D)$5J(&?+7<82LLF#:#T>]N:0/!@LPW-FF,GZOA4D;G7VV!<HC*3Q9H;-GYJ
P?\5!D#3"W'^TE_@QQ&CAE9\A$C9S!1*FT].JY0K\A M)I5U:K25@$$JCH]D98"D;
PF<$KBBV\.:(75S 6LX]@$6+'H^[C/&@[&A@R/:)]IA]<RP"BYUW6+!\5FO9E?+%#
PJY2"=+"U;\H"#J94?QXLZ9DA!>:I(%&?+,X0O>I14*_YRD0VY6VXB9NZ '-^W54N
P \4#UU"[&'W?0%I_RFF'<_7II,6[=^X?0$_LZ3F<N:4T7/7PHD\$X7BQ1.+*9%$J
PN9(NW3"UO)4ATMR/U[L'!:<JFM*+)Z142\"+ 9W@0WT=':Z=/*W_?5X>^;AK)NRL
P\CY^M9.3G;=W +&'55>_:;$4,GW>LGI]*P;#H?%^(?KY,>UMYVJ=DF"]7&@B]DI[
PJ[&FB$W\7YU3U,P6&:-M%_UJ;,$Q"M+'8N[3IXXG*,!A@]CW>:U=PH:P"[4C"3F^
PZ/+DGM)N90MFAJB]X]M1OEE%!DFT@T6YAZVQQ G^W)X95/W^)YG4%3HK/?Q'ZT([
PJA HJ@XFENKV9KV&;TD4O;" BW8*\.!D?<RJ/0G?B'FD]"NED;(ZTG"2WDI#F8H 
P9+W(&GL_ K/8^M561S07$I8"A!+%'$BR;&Q/J972?$;!C&(F-OB0(6 JK"!M0&WK
PO7@>1,B*^.T#OL<,UNF"0G\D&DJ]&SRC P$Y&2PY<;CYLJJSJ;@['(W$:=P8Q='7
PP]N)\+G01^NKI]7%*BV^CU]UI18V> =:<@>*@-5T02O"!$M)SDNJ>G#=^=)+M55%
P#RI_\2%_/;0N4D?/SIMNA-9S-M(R+!@%@!88\R:M]Q%RKM^N[]D,F4[,Z,:/#'(9
P:;]^[\P%;W,YF3(KF=0'$4#6ZOI(5IK."9@>!%[ :KSV\Y.SBXG,P1S(#Y;98;?/
P=]AX+0%*-11I@SUP.>M-3."*@M?@&9X]2H=*W *(Q:GJJ 4*I(5[$)#B8V]M(-:/
P,$J?58:B;%C*3I!_>0*F'TVP:W66?X0M-4JS'(&C;M+%.DRD9UBU@/89^7 $#G"I
PKK2BEXLX?JK,#K >$6V;F%-_(:&.3I1_[N3Y;;@5\V:GS@H:'91]]\UKK^ 1"H<E
PL-#MM3:+";KIYE--C:77UF+.Z<.,SZZL#83IC>YLL]#:"%8ZGE=>YY7/U#QO.OU<
PF:L\N?.VQ6O! ] K\J=-/O^>,MU:V2O^Y<7_9&?+FIIFXTSI_.(0&H/7D1K]/%J!
P"F1[\0],OWS@*T*;< 3S!8=^E!D/0'1J04#$CX<;#5N[Q@'T0<DF%=P$.AR+$G"0
PLZH(_.TO SLF5%_5)W'%49S)QW/[P!S%T:K?^C3LO=79(W-LO?_ UK?+U@/UAA4"
P4C$' =()#3)C$WC'-4+?0Q^:SB9"$LDR+Q[?\! S3O8B_-%/6*IR-$R;Z!1?5TS(
PM<\38$P*F#X\)+"G"$F<7:=0B5O(,"4VS)$ZD>1RD]@"]2H(=7/]_ZJZFOAL(B$P
P5U@/V-.=\^DY<,$BS#4P8M:N2'&W,=2"H"<A-G%HD+=_Z3$)*+31CMVVN$@X2G;=
PRZ0-H9 RPIQ)Y)%*PLL[1;I;KWJ W<[PGWJG5/(2MERF(/UR@*C!,0..F:DG/M$L
PA0: 2=RF%^49HPFWO6HSX2.T"JFG HCO\JR"'&5$]$/ZLV=K.H7!U\R<9V5QL22'
P;JNP2IE&R49S^R.6OH3_-B%."P7E*@RB(U)8&R/YT"[^]#E;]6&[(H&)>]Y+EZ4O
P=KZC$\U2DVQEQ/^/HLQ/&LIO9,'+I\&'\/-9ZG.TL[BVQD<8$76D0YKYM]&@AZLZ
PPK!&PS.[=Q"_FC:W_MZ]R1!T6DNF/XZ2Z,70;0KY!P,YGG"'U@TS[Y9XHWY?T[5"
P(%S+6 ^ ,BZQQ6IN#!U0HUY+?QASA'4]>IEXT>FW8!W%LS?"8\$!LFM[D000'22)
P_;AJW. 4"6SF2K5,TMGH1?$,_]1Y!V+X@]91,3K2[=,;O]#?,2.9WK"GBSI-9#8:
PG(\[O^27#32L&3'(2N\UFLUR8*FI/6J24JB[/LIC^#0SK06XN']F&B9"NI%W<C!P
P!XC;544'62YW?;-('V7UVT\7EHNC?/,K<+N!TB^@J384&'E+?"7P;"L<>%;"9Z9'
P@^! S-(H+'E[;I,*>CN^E3O^1+D-.L\T'$!CS<-Q73IC[<(.GDM]R@HB-F7A$T:F
P"S6[.;L):>;T";RMG5G<XK<X4JB0_BROM_:8H<8_9,%0K-AW\J5Z;L]>J:]ZV=PJ
PU"$$#Y[NUE(;XO4G@&$<Q+^Q:NB>LMWI4+^0=P$@JCE0/=PD;-PI.L:KB3I%;.1'
P?]*8=][Z@B8*!L&T^V 2/? A76DJ.&CVC&B[=1K#2?&*T]8I@.Q]T??J+E47Q7R]
P*C$I?/V)%M,:2PX9UJYQQHVITS,Q#9[Q4ET[M)BQS](QO$PWOE8M%HSEP^LM2#*4
PU\Y>._ICBI?9/NY,M/-7%>SR"N=["/)7EVQ^;4(;L1<TYL?%E;(MY#1<B#BZ SA_
PW_73HBM7\03VM,^88A8(,ULB@V2-*!J<8P!</BK<LGF%#[:T"C ( 7E1L18'YV1I
PGK\RJ8#DG?D8Q7\+.?B^R/#G.7)\EQ832=:I YL6B_"F"N-9HY7Q0##*@7%,(#JM
PL-I/)4C/F/_]X90'A/68259!]KKQU;>S.AI\RUJ/Q0_KQ"CSO- 0 2#X.M9&@F1>
P8=]4"KOKI!_J&"I%7K[V48OX/;R5N#]^LS!,5S?#)T+C2:A3<XSHZ? ^ 1\PIW@I
P>MZ;!/M_<&\G9;12ED8.S3P[*<3JH!KT.8]0@;1["*I)F+>!N._]5@P.5>HK'"F>
PVES-P==/&5D\"^#+7S$#I,6/K %B='))4CF6P *WRT:'<I\-=Y-?N6*GMHKIFTM.
PVF)EX)\3-D71DU+M).MB0D'ZW@Y89N(B7SLQ.Z/H?8F;4ENL-Z8>7;2T($O9KI.[
PMR.FGZ>G>2[;1 /%$;XEXNKN/0OBBVD3?Z!& ;SEHQ9GX^';'">H5R8@"P/[DN4&
PKX\B3>L6<CJYI/0RFOZ);9X34A>^LX)+WM_3)-\].&,IJ!]EY3"YVY9YHBN:'HPF
P) ]I@*1[2/&'@#FZ>QJO<%I:T$^.8.R/YVQZ!H)B]GR'DJ7*[P,;B8%M)S !Q87C
PHP\%T/H6_QI,KJ\XZNO\<DV;3.":7+=V5X$^$BW^T(Q<^A73R;+$Y"_ \7W/C6L]
PB*101_752DO)+M!;.=)*1>EX)HNDJCG]@U'4#=DY^S*FT;D)V5:^M&@8([]%$6B:
P\35UZD,'5TJ>%:4>V.]-\%,:EH6C%R!C]WL2R3\'8C#)HHX("M9KV(-"&I)VOLX@
P/W=/F$5IOPV*RX^-%Y=(H>>U<+Z]1[,G('V=]1.:[W<3?ZV.7A&-C_=;C9A2PNH$
P+\X?A.4BU?"9%C'JPZDKJ!LS77/"$J(5L2E.;(E*)IU2<2^E"X"ZOAIZWEBM!X/J
PML@F)[^O5Z]@< 20,,8U-92F-QEY::_ #IW+2 OYHD5B*QRY)8R]5*=&H V..<K]
P\A(.?AY7=VU+XB?"B8"9,]-P#@1H)M/=+KIDF8@P(L+EQ;*%]O6C<&"&RQJU4/'2
PYU3RC3H62' >;N\%\B>R 9]5ODI-9EF)5I&584J1ZMOH5R#I2?_=,NUUB ,3U^;V
P68#CQ=G]#).O!@D1SIJ@/S84]45D?YH4_WK1Q(2Q8S,F2EK0@44,L84U4($.4YD*
P-62N9C38NJ ]IM!>Q5;K+6YBT.+)\.M['PW<)L_+IZ[7:FOF%G\=@PQ0']=Y9JBL
P9RL_4?6B)6-. O=K5Q)2%)R=($:W>H*@+! >NL32:MH&EXVJ<SO4DG$V9L.# S>+
PCO]\?[2Y+,]]B>N'GAF_G.:[.BC23*3^=08:96S0;.$==>ARO7R^Z^[N/]*B'A]B
P*OZ^UBYR578I)G()TOVB75C3<4<&I2#DH#;S9-'#I&O-'D[V>FHX>T)A"5HI"1AP
PWJ(#YDC"<\8<GZTLRB&9,"-@%*^"V J?X#O9PVIHK*SV[\!$4BB-,6OQGLQM;CC?
P2]8CKWS[\Q/7":$#ER&?N]/,HWH?;Y,*5 *7IW@;]'(M:3VPW:H'$)OQ&Z"NR,#C
P^'YJ"OOR/.5.A\UIZ1-QO^WM>_7!-.%^K$K+_/7LV\ZEWJIWR\ITSVT"VX7(<T>"
PI>C*T$_Q6RC1_U+7N$T["IG[W"O@;#*, RW&40\1&D'W"E;%[1\HCX_40CY'FT=^
PG0LV](:]!VA8=D'I$'S+"SES#KT*%C'V\H2:/WNI&(+ WM+X(QK[9/AWRFF^2:G(
PY5M"7%2*QN<R,2YW-NS'@F8W#'0^*GK6;\L;.*H2<V<[XEHN*5TN8;L%YI7E&:[;
P?L3MC]$/I4B*->FP"TG(8@D&U5/90++0.(Q_ I/O.JZ+JVFD-6%AI"("2_S'1G)I
P);"=;&9FZ]B+$*?RI&)6]-Y#0WU"LLJ/$F9J?0K[V#M!=9*BS?JZNUAWZ&QDH*;U
PX#UEU@)!2AYGCHTASTH92M+%P\%7%_X?@^/L*4;3^!"LBB"5#&@@W<;X8[A!2:KL
PM>=5[#0CL,851XT]>#U3]"[QF1^>=J2^<9I=X,1E)*/X$PZ$A&[KM#L;H<ZLU1N5
P((]0O=_R '=#2^4Y^-R"*0LYV(S$NMPY%XZ0PL_)Z&9!,,6.\*$2(5L3]6-3]B![
P/4,\!=2\O/RLA%F<5^]DVDEAW_]K!_,<Q\>IR1EP1/:1,;*78YJ/0_"M":N:I^@#
P7(WTC^HXRK+,>H$50KS?RJ1MC$=+/W0M5LK!: O,4/W5S(EZ^.@6)P_9'KT\[1($
P*1.D>(&)C+-N[IGJ<+]#^%6GH&3FH2%TW]/V!-E3+4^:$GLYH_M_6&?8)G:)%)(E
PK\*:;L?PA[)4//Q4#U<O.#_ED(A9;+WUDC?,37CVC!P\>%D\[\0[N@XPQC!AOIFR
P@?8,O-B9F=&[+S/%'J;U42]=W2G $3C>+WVR%C-U8>%\'_/;0T=X.N1$*1:B%O,7
P';;67:<OR$8II7D_EMKI5T$8PGTSB0T0A\_Z.*3;C![&[%E10P]_M#XJ2 !)QF2%
PI>[!THAR+@ED8\>E6?RQ9(!H0I4>>4&UQ+GQ&BI+>WNDF/DV;<*;8\Y\(_1O':7S
PM%4:&,GR+%,H(KFD][]Q[)N[@T,Z6&?)ER(72B7@G@]">F#A'@(.E&\5'D$!])MM
P=AH5Z@.;? OZQ+TUU\AHM;[]!JF\SH' L8[!0HZ>G -^G)3N8-=6_RB4$(2@BZH*
P*^9O6SG=$_QMI_*::S5Q!=<>15BF'" 7N1%64-XS,:-%]MPXM6,3%.,;QQ1@@>0;
PG/01 X[3]:F<THG,FNRW4WUEBDB5KKKU6M!?=(@=KSK=QV^99NQ121TJ)DDSV,I!
P5TM\4\[]90(?M1M0/(R+6ST#!4*0;MF@=6B/'?-3$)0W22;P"A2ZGI]8C((D&?),
PZ3;H.;PPOF+'!,Q?G6V&@KSF/0;39SC.(^_0*O-7V#FP&.\=Z_XPF2YVEC#^XJLM
PCN>X1R$U0-9S!7*[(UPKT52B+\9SX$>0*$H'[T>)SY$*LB"HX/-GB^GP(!AO+P%+
PH:SW6"!U+S<K9LMK*6,L*E!]+/#M2DN"FMI:'M[UM\H424CA#P?\&ED,;*PH0@R"
PO-[%ZM#6,5^<'&KGDY9VS]=X64EY0.1"J1R6$8E;!NI1VEN8/+@N-R>Z(R!)CF]:
PC?\JLL<W;@<XGCI381F91#248CV&Z2K"8?S:?Y/M&U'*U2X'*\C95W@L#W8 C6R%
PW(+(6/A;N>,_9:>UT[%]=H9@:Z5*X*I&7"LA-&S^+H-VT"10H=F@I@A0!,1AWDF/
POM1$UAW%B?H:.3WY!BT% _K._[:_SI&M%IWJT:(M7*"8T"DYE619#ZC'0T5\QL18
PR+,P!>#IP'9*K)80^0M+I0_):\4H/5;'6RWP>(N4=(S,HJ[?6!]3L*ACP' (3D5)
PK++ !D"5?(*,56RON_87XR $N#>*AO[/02UBS0*_"Z0:I(KT2,RP2ZZZE3Q1SKTB
P7?&?\6403VWH&>B+WVJ@D B$!Z[Z(X6=)$YV@AG'-]@TAXV8O3AIQ^TV:U;>/.CI
P-)F#D!_0(8ROK,@ONQ#TSNS2AT..?A<O-G<M"F/KH'2)QN'"GXG (2.I(<5R]["Z
P^+F&.N&"OX<N\[5NXZP):K=9!VNXQE:#.[0_E2$D@X$S'C2)F>:8]"P0]<]*YQCG
PU;%'&S>Y45-?,BD&R.F+:? R@E! ",LWWP98$5O6*ET3H3V(R[SX".P;L1T&:B-=
P,YWE_D1C?EBV<A[?/I^VE .XT#S^5(JP%@7JS_+HO3@CA/ L+01-2!)5H'&WTRG 
PUXNLPZJ-52)M4JT%*V813W&W/:S#X(Q\/=)D@'.]94E008^:AP-#'93)M%(<(A]N
PB47R!<,BZ;EA!R#.1GGPF6A41@Y@!2GR3:F]U\Z+7]*ZCIE<T)3!2"=BTA&CH# &
PN?,[4%Y2C*VV5HP&^ZX,)A:9J4*_406?SU&^JY,)X(>**'/]-37]Z=OMCZ 2AY"#
P&3\K5$M/_%E B^672(6LU$J[C(>]CLCC7M,L*7:OZOSY$BI)-ILW*I<??O_KM,#;
PQ&E+!@1G,$MXK+G516I&C0-@3 5RY0"Y:(QXB2?.IQH;8U@MLF^R"9,>G #BQC@&
PE/NEJYF-]"4="<JHDZ%[#X_\-["6M.T# ,<QKV,HU@CT-NJ74B?@7GE44?[?(<8Z
PFMSXQF$FQ]:4**#;\^-"!!T;JI=Z=Y:C L+*LGJ!H(Q5GP$D:4W&:MV?6!+MV9E0
P7X/,V)_3=CF$?-H. A6%FY?)0X(.I5!HY_Q.[@FUUBJY^<RZ_O;Q$LF@58OXVW-7
PQN[J4B'KSU';ES[*"/XZ/X,VD<Y_-XX#\N!DP;0NS<VU>W!,)!&*!-Q<[_4+*K+8
P 5NMXE66<,Q/*ZSL1G<!C;_-PYT=8FB -$AT6,W/YI<;=5;]KXU"M)KJ[?EWC<@>
P6&&NXKSB*>3'#&8:HJW>AQ>'_&7?H9[FZ,MO6 V3>O8,_#VWQ7A-?+!=\,2SZKQ&
POH;D>9=!JO0=R4Z"_^CT<7ZU2"D^@BYK$P4MYGO/'B*^@]&\< 97PP;&%(XNF#'S
P*!,\85QRUSBWU/0ZI6 O4#4+OCFWIJ;D2_>/ A"G[HO(&=]!>T/V['N'<)UY[2WW
PD#[T)Z;@/LNW/E?H',.#27Z17(#%Z+P /-:>-V5"-=8* !B@D(O/25)NC9; ][WO
PW-& -54SRPDV4 >_&H=8%]=S&QO?PC]247F;O&#;XLD[[OXCOVIIIUSP=3K45RJ,
P]Y>77$)@A$E2H\+:R]XIT(Q[Y4'\*!6AUTQ?_^S$[00-U =D@,M&^;G>6/OE*RP*
PB&"-=A",EBP=BRI3G>B>CJM1SV)!X.Z0H(.SS=86B,G%\0*N/S[DR0_O&9P 6/.)
P%X&\L]5Z?)D7&E0ZZ.251G"RQG-;FN+5_ /D/YGQ9,PE=YCV3<"57!>2RWS055X4
PLZXQK== AB6/35@Q:5K.;WI&>%C)A[;+\<F]N_)G!WF"^!6AXQ8JLL0]A/6I6C'M
P8,_.><HUC--A'G]]N7F:E0RD+YGNHH354@_'"F>8)E2HF!$NZ)4Z6BG)3S?<@(C7
PEU\H]EEZ9&A<Z2FE>^GFS>P 4SY$+/A#JVZPIJZ%KN'.;4- R:)N):QJ<W*$;]HS
P>=AI'6))K^A)F?/Z@Q_<4J4 :)I+^282^7F:354'E_ZXF5\2@^;N&86,AU52RH8?
P><4I-?_T^@CXD['Y= (O;6\->+Z$-A]&2M*:B2TNYW (6<)^F8Z>J-'S$+#EHS3"
P)4'<O3@PQ*?E"-U=!I[O1P+9BL2 T[B@3C#[E[(!^X+@PL%3GKK*%*/4X -@U.^8
P*0^P*N.F_)2TP#0Y7OHK'7<,"+MK\D7PD&.&490JJ-%(;#-#. A=M_+.-&L7PNR2
P]C3CFA!: \AAWXDP&QQ<)/B*:9O#^<'MP/5&'MV"HQ_>OXMC,&7>=*^!%'CY#3%$
P^_,R?:K8.P0]8Z6_/JJY7P,J,903JZ3P1%T>>=2@2.$U8!T'Z4ZC%WT$E08K%Z67
PH.N/0BRR,X3'@^U3M8K(;YN0<88)X*. 3AQGA45// U]LK<[2K^]Z,OYV1[D;[7^
P0/B=J '?QO)\B7K>7$;$9G)Y;8^+08;\06(? 43- "X-$+L@QXB7B3\-KN4 K'/"
PG0%RM]4A*!% Y;ACYU3"X@/8C<%!9XY[YY_(5D3F5@T+I4HLWL'/#.Y"!=&IVO5%
PMNL">TT<M_M!0AODV,J2CN$/3VBL'+4+I3$Z6B[M1 G<ZOL-:U$,Z('+5Y\. <P'
P"XN&;F[P'+][YK].?NB4<BO>;0"NR&_\]^Q)"N^\PS0_3GW!JNA3)]J5!MVQ_F'>
P/5DT$9G2]I_[)0;MK,IH$#N_/.6889.I=021CK42@J%,YWCD/,E77K.+EHHQQ2!N
PJ9+RMQ5*$:Y_MB),T?7IG(Q:/^"CR#.>@A=)D>3]%!RD2(QOF)=P8E#I<('*V&V1
P@(Y_2FS& 1]-JT#"<-7ACU7^Y3O<N&$ ()#<TN@ QP?]X;[Y_Q"O#U\->#(*-[FV
P4EXQC0\+V,<;K]5U94\2C@OKOY]P^>:O-WMLI;J.&NGBE*KKCE-?S+^;2,%93[(/
P=L00V!NR5PJV3W)4S,CPM0F!3@ FF4L@'WO][WW19*)FHO:P?*TK?<%=L;/%NEQ'
P.?]/OLH:+R,TF?AK]?IO^IR8.*D/*8=$)2]KG!,SCXY3ZQ0\Q:;8$)LYW*K,U/Y)
PW2K"9N7["F/I!'GT1RH;P[>];7&HQ.KN6E5<(&\55OK:-J3S$@UG%6SUDJ1LGCU.
P GYS<\F@86_0NN9(#3SWR#^IZ>\\"1__%8TUL&?!!_3W&MN'2N(W1&"^:@R !SXX
P0,#VM&2VBSQTF/@@/A:5'#R./T'V $:*4RVO9O^H13@>$&*9XH[F'Y/.OET/>F&W
P5IO[YJF(I&&7;^[S ;\Q@"-W_B9<4,W!LO9B2-5[-)E.%.+338#$IQ.DD:8'E:?[
PW1'O*,5O--5]DVCY2)V<#"-?\JM;+E;5<JG.:P *YRCX'L+;7R&[<+$?[W9JT(MQ
P<A;B4E1TW8::W=_&3/,(7Y :8UBG^R;D#44H('(YR=HF[,* B6>B*NH%WJ44259F
PY_BDIR+"HKYD*I $;[-V-! AR.^6,[GB_%\Y<N((VU/?R-2&&7I=4(8S,57+>"J?
P_->.Y_E&P%=@S(DT/":52@)VP$32+^5[M5>Y210OTIUEXFA;B2OCP"-Q^L/1/P10
PC="C+=C:;#4^KG>W2=:1Y9-B/R>(G=:.3O4U;;QVP(]W92Z=HS2@(9[_$L5L ,>>
PM^,9OIRFK<M*$W6;ZTC4[ZP%X V+/*\JO9]7PDL*GGIK?0Z[(!&Z"HI'<@)1GVOP
P&*[H+RD<#G8U,W,$-$!]NGPR/G@7W94,>2(.;K2L3LF$*XBO#?%GLZ'S8>EZ* 9P
P33DH$\W&;Z(056,5X=B# !3#(=@9/29PC4NNLO(E'YD0(440G-++MM QED44>M!\
PU*H-&P=YM[WT(5>+2G)C$[IL,!Q*D!$>XGDB#5;X%NM&_2!'W:T5L0?DQ*O/)A+ 
P,^8L:#SSQ)*=W_TY7S>_?N(=P.<V]U#$+/ER.FHK(^2;R4QPE47],U)3CEK#GGG 
PPJ-8@5T'(*\V_-I&E2O+*,,&D8@TF[(9;N:=GL.T1[UI? G^WEUG6[ZY(KXY?W2_
P>1\EYS][%"59TA&>R%DQP290Y%E+0IR4*$'LX^#FIG0^(T+^5/?'>.D4R-%$J6J#
P>W&LE%8$?R*0,*3T\.%C"JKR5F@9SK!\!L$)"4*;,QL1^DL?#L37V% 2Y*[ <S (
P:_IGH6"@7X8?I3E3Q3K>0'!\M9S]\A C.$OSAET+HHCU @1!)@=P%Q./!V,[ <=#
P*#B==TRI)GAN8+<A81VCY.TGH$' HE9G:'ME51X9M/R('?7,'"!S6LQ.GMU4EV]8
P*AWOM9]&%R"4Y=V;XN,WWT+7H4"OU$S>LG:^=?<PPLA_'$X*B4?9=?L>%2OZ["'5
PXC(CYO'BV[#(0GY>F5R4\$]O2[^JGW\$-?3" G!4IABV]H_VZ*IN,_] 0CPF#0S6
P[?6WGV(;$]#N0>%TV9'+X?A_B2.@UN=*H7#@J;'L#4!CF9/'!45AU'!V"4;G+7%C
P] HA\4("S)??!9D1A+*%=A3YI[R&+DK6W4)/$]]Z7$L5*ZC$S'6YXEF\7H,W+@&F
PKT5 )_5)+L62\N<KGL+W-1>0;L1;Y&DI]ONAGF)#Q1;D1@K3A[G73U?YW)/N6=(A
P^$5F:[Y2:H[I:*R\1U],S4SXK<[N=OJT%6:/ZI>!AFPS#W10P)$U=,% (5KDH7YK
P9G!.+C@%W)B E?%$L_CX\D^:75*9.VL<7Y(_8[B#(L(HZ](MC-#DV1&0\/0#%0 B
PJX]%-@H:$KNEK I2H;$>^Z.]$[3IC=YS_8^[/V\\PSL<JZD#5&;(IC]&?N%UL3&>
PRXG:U94^4!CE /R3&/\"1&NUDHB: Y#MC:4YQE&!=%PZI.ZYGE-ES;)>)4!+'T+H
P<\,6R@[[SK.S/R[?[!4 DWZ='C19?_/P5M%4FFK[TH=\68R7J%&*I#<DF(%Y#N&X
P9Y^R6EV9WCRW,A=6[:&TT&'+O5E6%S*R%H.%S01X[3^DS/%>NP.40'(1]GKJ81X8
PEL17'4*]Q(6/;@7_XL;4:<#G1TATE0RW_0^@:X42"2Y@$YL<TC=2/=V#/UL;V99'
P[.E]_@^U:5'O';A2(E GYV%GC]YHS; >$:0[T2 SYJG'[[[7HTJ=31:M ]S*4\6(
P@>LE%N/EA!I]D JA.>^XO^Z+"A5IDH$%XV<!WF$+SH_D8NT1 *<>M*DV/YK(*VF_
P6TC6*87>D/ W1N?QP),"5]1&]:SZJ(CU(B\/NK$@EA_('2D\5+[S[6O!X;@IVD*Z
P)DVK-:<P'\!18$_^>^D86GQ)&WJAHNERHZ62KJDO=.[I!3MJ*>]N2KE5.JZE<D3D
PF2D5-G\QA_JX_O4ZX7<Q2U.%\]]@&0P1(.9ZR&K0*49\SYUW)X7NB5PZ&J$Q&Y86
P]D>PS"(8R$[LER(<XC;<<;L1/( &"G+-=5O4X(I2N/JVQC[H/>LEFX! !"D8%5B<
P;%A#)F/)F0LUG5-BP:'(OM!\G\C'3[R^60(-2@[5T;=[E!IZQ:T_O8:$(X[9]'"9
P,$]&9;9ID*]T2R8JH!.NJT"1*=)D+IS=^YVUBJU[YY6;A55-S*BPZ1=GE)E<2'84
PVO%UN*3NDU-\G7C46 BO!HZ,Q"#PJ*[6=^1,P&>;*T]7/<-"H3=7>E^:"N&PH$V)
P2^-^VTB,X9W@_MUZ'=JR'A2B'ZJ::;7>@ADP35>SYU-)=E+ ]78&78D7DRS4O[C]
P 6P3"4.<0UG2RI1L1K]R\4\T9KYY+4C</VD^+X)6@%4(5C)[\)_DN<"#W22,'DHV
P_X\F/]5)BB=,\[)-8F;S2$N^DT?>5](/*QPN?W9#C4>%C]B('D_%=F_87\*6$G.4
PW!Y !42;O%O67Y==^&*7K0JVY'V9 ,=1D"/L:]8BJ#W@TQ@5K"RY*+M(S;(@/9+9
PD[ZQ$U8& 8JY4*+,?;46YEOV$H:E;[!C2# [2%7PQ;)^Q34+;)Q[RUZFT@?Y7MEH
PW;1O1NFOZ'&]A0]0*BC"\ <V\N8Q8X+:7Q+]C>K9=Y+WF4H$H-Z!NK#^&[536DIS
P>TWI>(B-X=4^ZE<+>,HRVH4@EMK9%_>P^<JM&WDP04EW-K*KV87 !J:$X%G?^#E6
PBP99VC&;N'_8V-3X+UA( 5,$7BG$-O%GB:@>)JTRH%X-FK:__=2&YFJTR:/=T<*4
PVH"5^)9*Y2;$T3]ELOX@!O]6)-TWW#_,B];.;D^O-^[B@BWM'LTU&A7,D7TR:TMU
P(S1]6!'_MBSSO%$I4583_8T@=Z9R 1"Z_NGTOP$)-LHW:](5N=EX!CN0EV!!DML-
P[>*>T8YU\ IC&;Y ;GIQ9SNI[S^A3@PFJILHR-SGA+H^:640"A=WV TFA=P!B2"(
PN5J,2@H>,?)D^IW-A=WAS/Z7!O0&LP% H!9*!N"&3';[&E=G"<P#$SQ=5@YM4#-F
PW.I58L(!E+=DF?;5_]#0;5 #_Q8@+9>6V>TS5O6F5(N%O\V62V1.;<S+ "521)GN
P7@$D"P?KIX<^T8JHM50CTDR[VU="XWALZK6\T(4!YH[/"4Q:"?H$;+"=X+^YR'";
P+MTWBE$>NCQXS\2,%O+^7UWA?W?Y,U0]BM\!U'X@6<!6PDP>NU^++OT?R,QWGJ(E
P:=U>^3(!XIXJ4 5VK[FW;7X\&R/> <V$=P!GVI1&<US-\BQH^6_5*8J;,WR=-<2L
PN[JQ?/F"_4O*&S6]DM)]U0<A\;VW_;E^GQGVY>YR7DQ4Z]U<F*'T/)PE71ZR@U.R
P"VPR#SZ[RM_WF@4,>&&(/L'_2I;= &=#&-T43*_:][PIL:!&O>(-#FI><]QIZ]&O
P*ZBRP/CH*OX+IE<>;SN0.'7Q;3BR<-AD"Z.RJTS$$NX5S !PP(TS8D(JSGZ _9'+
PFA*3@-P-.6W%B P#/F-8AXAG$?13K)0K8<8;]C5]/+^[\+\(RL*\_[,MK!82)>TW
PIH0W#C9R=NQ*6/4HCNEQT8VT:3KU>G8JO\Y)SC*PW-#-7O*$IQ3[#Q*%H9X/!6<(
P\X,Z?FQ;!MN#H>>9<83*PV(@S@Y=+7OI<U8+8$%F&U)^&7!G>A*AS<A/5T$9H4%M
PW!XFU$Q399]E2:3#O;T#YWVH9M'MKO%C923:M)QGLKP")\^&XRK?Q&_(ZD^$*BWE
P-$J.A@;+PK9A'!=DBY%6(<11XGE01@'EWS=(FGPI_2SKI.PMC?I!#3>F""HZY'G<
P:,T8GX=L)D[G\1THT!O*]V@C,?GNE76?? 77C%[.M/:T\@>=SAU0QKF?<PE^/O.J
P\$KMBF@'"'W/"7ZE*Q"Z*5.HN39JDI:F7N LWIU;%'-> $]?2_B<#LZ0K@*VM(/0
P/.QF1TGC8E,&08*XW0$7RT#2W\'\8KH\J0""-M1]9A@L%)#[*-C;)L:VA5.(M/-X
PZYAO$V44H*-#0>L%9,B(2($> Q7O>R\'J7+544SW4.962GUN.\,B'==9UJ%M3*2G
PG2"4UFT9] VPAF>C8Y(%VD<W0L<Z:JKA:^0SQ0Q/%VS;T!<@^Y'J='&6CBEEO)O\
P!P:_!= V$SM."6#1^?)0XLKJSS]\:0?G\N_Q]*4^,"+*;Z[$N #=DMK%Y\$T%FCC
PWA#BPCH%[%)@Y:;;XHB"\DCOXF%.YEO'Y/>#3<.%*R9;@&D7.YU3#5 +T@!K=J'Q
PSX5G<'$Q:U3ZJ3.'%SQE=K*?5>P3J?V-H$?)DCC)U8OY8(^RTXU<Z:>Z^3#6>?-@
P)IP8QUVJ;D$Z\,XOH$2H;LNB\'> VY@&D\>Q45FE^TS16DAXK<)T,SV29@&&$*/V
P^T#H@17FE8XPVABQL=E"ZO&N3,$7T+#/BNI4=G$%7@Y4P"P<'JSA+7U>JKK85JQ8
PO]HZW";N&RV@-7A!!-5L\$0M#BO44=&'_([A&#C4CTG'JO@H&[R468FLI^2+2Q2Y
P*N]<CBQBC9/R*XO"@N-4]_00HH[:$?MRE%4!:+^6DWDO+7ZLPU">I-4DPB]?<^<'
PCOB4J+ G:?NY,>[5W@<<A:*&/X++E+I7!3MP[Z5W+)94A7A,"ALX-*^P=4RC<]$=
PO9H/UGWZSRT/;@E;O5+ ""\1ZFMM641VL7 GP-*DQ4MPD)&!11,Q(.UBZ(QAP8J1
P@!$*1JOR3[%+!XF2<T"%@A>!# *65 !-F-+,6R(,^@%_\,M IAJW_I2)ZW6NJ4D/
PDQ<<$#8<[Y&8F$#318\=X)J1UFA$"OSLGI>MDH@-@O9@;H_("O5/!8SDSR'C@AKU
PFY"6)14>.=B3(___ RJ&(F<#/S855&1T[5$ QHS"Q7U,"!L:^0KAMEZ:.#JAB_:%
PCA(L)U:;;Q'>O+:GW-T[Z"-%QN\\XT>$;EI1;9=M9<FMW$3/GSPKL\N"3(U1+)+%
PS:KLB3,0Z(ITC3+'((8>E-1!<V, =<]@F$4+' J"(R=/I9)C%GC]O'5@@4SHPY&3
PF,9T"HKQ\UR\YD]@CTNE^8+9%WM.F>TSUO001*7+6]O3)JP%N]Y%S_7@93[OW'B[
P!63Z#TLW67T4O-37HT']]<&(?/]H7\R0WKYJF[91QA-3?(#D;U)]+"74M#9)*T][
P^&6-"V7!])OJ5RI:QYAR<%ZB3EZ=;62SL(URZFD $BZX0/(YTT@)U=>UY"Y-I5_=
PK$SEVUU*2[(:*GGITSK8U:TH@,;0X7=[XH<7S^L8/KJBB_/\^VX:+,Q8F8%B\O\6
P'W)@[670,O'_I_H=[IFP05L*<K0=+L'>HE_TK[QVC&BZZSZ]9O^!@I"6Y"BZKKNK
P,S;$K2FO=Y_:@7[I[SQ*ZCLM5=_.A159]#_T5WES#<@YX1UN3B3P;E4_[,(8&YNA
PY8LY3RQ8]3:;JU,X!SDZS[&_E J0D\E8[\;5S\36(0RBT@#B0/N56#C'!;.$?$,^
P59&19[$SN:V CVB?IPV>,*6;%!Q4/'A":/"9H='5^<A^Z6DD\35#L@)I(9V;:H+2
P+#<(%&Q$4GBAKY^9)=9IEFQR#QWZ FJQZ;])O[/?/FB 8DW>(0DC4/>2,&1HCL[=
P,K(/!\]6RLM*JMLG?IC<:Q)FN(CD*A2IO8GZ8]-PS]R[Q)*5R='PBC4,_#[;0KS1
PHM*4G,\L^>5,Z&; Y$!EQ+4=[E.3[?UJ./Y.G>?K0SD:#6]5ESDU4=:E'*[\44-D
PU0A<_P;3;IEZ!C1$X \+]"N^]#?H[%>U0H"X8W"1:N!AE79"1%EMQ3C_^RWN/S*@
P6FIH._'8^?P=\@:5]CHTX-V"R""!VH.](K_OT*X'B1HN 7* =P "=GNDQV0[M?(I
P88?_-1ZUC37_%-U$.$%+4B,@-5R'!_:?BN2_:+)<8!SZBQ LW2!G;PX*WWBSL44[
PYLX7:)'WM+-:!X%, AN\W^E6BGV#'# ,C^DYZBYXT">=/P1Q&+3<B9#>I#(D'1J5
PC4C#=UZV%"#V_19B\)#ZWNKAB(N5O5GYVU]N1Y)\$!&G[ SQE_CRO(6!9 .?2+,<
P'^#W&7;-IR+J 9\ JB042>^?:V@_D?8W3:8W_-/KVC<GCHVMN'XR;EJ9.F^5ZGPF
P>5B2+BEV30OIV7RW9:R9(7HH8WU0QR#"C/>&XN/LSYC W&T+BW>"5-6(.*VYIT^"
P)=5")L579U_,F)2"[%FW#7[G-35<FJ1R:\.T!A%=@(9FE"EO3(?\Y?7EJ@P:G&\5
P]'^7[U.X!?:T+MP[G7[3_I_QXKX/S#4<S M88_A+3Y'/@S(9G31CH9\=M(8[(=K&
PD/PP;&!8H,,(Z%CI<%[19@_PJ'4:,*WM,0K9HU#G]/F-P 9(BE]=I:)IIJ'.[6,7
P;"LLW8CT?:FS99'4X\H!V1/\LK*.]0(CY "HGAL)'7S2TB3 TP61RF:9L6]>QV\@
PQ6PM4O,NQ#@U-UI$_8@YX-#AW=#H!0OR1VT6)E,PBEY\"8<E21]D 3(']XD*)-"]
P;<B[A77J(EJB!PD-8XC%8E)S]A%0>SIDC]2C#V#7AD)<R^%7^%49EI@T/F9SKA;H
P%^_HQK%4!D?E2>H_,R  .H@89#ML+BFO0G[O#17ECV#@;DDQ@!<U.OP,O%8057/R
P]XQC0FUW0F6P&<WNL@XB739W,);+_6/[/DOB!,M/ZA49<<X;)8G:9#O= (I,U!J;
P*I$*8U%TW];.<:^/=*4JV+T.Y=C=O_KKB+97_\]87@%DY(( -EYW$D[?%9JE_ TH
P*$7Y(\'L0PG06>Y+<LXMQE:(V"OA (Q8_0TV[2:GJ5*4-^DSF?+ !%I*XT>%/OJ4
P7&&?B23FND1+PDE#-"NT3!LZI3#,VD$3!V+MU99!H.V 8>>MWPX/&ZA+O,!-E;'<
P+UW9$%@H<H640=U!F;VRM+RTY8UU\6'RHI^U].F!3EY'=M\J4*>-.\BY11=<!Q<D
P@<CW[-P7GSOVY;+TER6>]B2>* <$1W9=WHWRY\ S!INP1NSAT/ZTBM:@5-T7M@VJ
PT\]1KN*NNM>ZG\EF6/B'LNO?]DK#7"A<MF:6"72VGR"#F# <XOUV:B)7F=X0> (5
P/*(-,5>;O8XH&6*(")_BWL%+*8M\6*O1]VH#L"AO3H2^&$Y5DSXFP U4CTS^#"5S
PX/AVMGR!FH&-N">$ZN4C+30V8/L.7*9S-KFG%SYNV#3Z$$%A/$CZ@RAWECVVE/@D
P/9O/8]>_%%/6C[&=WB)1<.2L1'9FLF ??LI@NHXHS#(#.>^;$JD2*G%GU<V4;2AY
P&@#H0DD^K>?56Z';612\C+\8\U-1B_+[\B/7A,[8U3=F4_-%-T7Z2/1#?'MYC_[V
PR]"(*0L#L<\_E$\/X53,3WSXK@2_/D;@<^-E)VFK*G:4\U##55I@F.#T3MOZWTSE
PZL2=[WG9X"D%/\ELME=T+70I.PKLWAC\I<XL]EW/46KX'P7G_3]4Q<)8HDM1?H&"
P"K483S+$YI]*7%?E3)\7IW%QQ7_>&VJ.[@K_W%3VG[3YY^Q9:89F/(X'\%PO\"\=
PL =7Q'TD >))E4J^!(=L-C8*RN24A>.8D!N^? ;W7/[9SFXY[URLW"!9B0VECUD^
PZ.EFS_/B/MW/JM7;K[W-G<9&2VM@/N5?E54\PXFHAHA]^2R^,9:$_G-J[#JP<]^^
P].R(ZEC@QM-O!((\NUZZG)PC5@HZ:D/$\V1 O][D^<#@;/28^[M>H.7)Q_<5!0'G
P_0[RU[>V'+1AJ946.2!PT686F@[BUA0I%_&[8#K9IZR:\WL$1C$T"*GD1<Q>B23O
PP^V\[.;-R3?G:HLT/A.0/-O9Z&GI[&%7C9$E-ULTP?)R-5RIN)XTP#-_!Y%>1%E^
PZ81_+%P +JV8"+.UC^B'G" !H'9Y:/>B]M>]1B-94+7I?R^1BGB'KGT_(W]#?Q-?
PD!L2P?(5IO.INLS7$X<RH%"KV,M8BM736[\KB3/^.A1!OG-J#_TF3)0+T_$%)014
P>2_H09D\9TT*4ZBJEB&F(B#LS@W6]O[,>;,^/--NE2P6/TP\,+XU"M??*9,Q7/)1
P2732Q>RS2/9F@&N%(JKU*^0\[F)ZT-VMS/@+ JL.F5-9C^9@AN5+K4NZ31(:='IO
PXG9%D E5&@H>)6^JM;97)W>>G31!:"Y)QYGKN_;D;^1E=<1%XU9Q3J. 7AA33*N6
P1\930$:X>,>%H45*HO8>_GCV_Z+GGP/P]K!"0SHBO6@W9#=EB%3=:K"R!L3<W""#
POLY%0_143F,JL*WKTD"UCNW,:JBHI@=2?Y)NY@GAT  ?8@I)'TD;^%]U<< /MF?^
P35ANWY<1_=3+:%++5AX/?2;IW(^4?AZL3R4RH1/ CJ'G.7R!H9**\+MX%++TYP6O
PP:]N?WQ5*G(0M7'AJ :]\?GB(,J]"'W5H>E_7 QB,F0GT(U=S)OE4_/N<@8%@]CH
P'E@\/ )NOO5>C1./2TN,^9E85ZFBY<>4T%O$TAOW#_%7E^>[:;7P"J]%J(E5J,.-
PU)WX !B>)?0[*Z53^+AK.?,)W#!B8#K"DAE=N^F5("C]1QP_$",OH01 I?/ ZE<$
P4_?P4D>H-C69.-0!* DG4>/; !HH3D @L5_\9K(XP6[K]C?KKDH,[YSI-]T<3.)X
P8*"RH,=\,2YR9VB+'E.@0V5J/ELA\;YB<>$<P P&[>.<XV.FR-.E5/LM+(U,6()Q
PHZX?)!=_674<$?3^B2FZM856Q+9AO&U[-:(M 8M)_STL'F.6H%NM:P2/C(F[$$ F
P$L^979Z-%3WBJ@!ON-\JA) /!C"[8$&'RP>__)W"/H-V:;MS**?),R'.7!/K^.L-
PL)CG*D"9/3"=+P20H"GKW,;8RQAJF<J+'500Z,0,00<Z13)MM,TDD1_Y43R[*L81
P$;*2RZG\8^PE7H!L!\)@K#\(]+_> >Q-OVEM\)OUG>2Q*.K.K0W(A#"5X3I-0F3V
P/=4LI]"=MMC\')FB.NUPU<1U3<#2@(<698H< :9[C<E?A$3YT"J;X>I2F1QZM.;#
PV[<TGIN;!*Y\U+L [?Z<CG:1_4YF%;_V !.+HW/RSHTV&'UX]E'+<?V;<H'"N3@)
PV!*D4.D$:$@O KDKK4YSJ).$H#_0WYD$!'@MG 568)L[:&L/[MVXLTW]W<LQTNLN
PZ'_$LZB1!LJIQ,,WMR95VT-]G4:RC]?81;+=<%WW4XFD6<X3Y48]( )+#QOWEN?-
P &2C@&=6MNU7TJ"VQ7%/Q;[=LW%N]+MLS>#0-@!/!MN 7 >'W]<\YH6\:8NDF_(3
PB2"/BV=P$Y<Y$7H%@S>[R)ZFP:K]WU4:J&PV&#:5BU_33LEBQ?6H3A@T""F=ONBK
P&;1P(2)S]] =X7,$-!;.F&GO/QJQ#X<%%UF99LXPR4ABK[3$:"QH-.-C0!++3HVX
P92!AA?V$HE^HXL_[7R4!(&U6XT.F]<@&5@H;.(0GB6.9L03A_.<AR/IU(AML[=J+
P+O)F+!7?WK+53:Y7M/9]CE1A<*!;=K@64!LYR8U&%*SCI(6X7UHH;AVRZFQ_L'T"
P214WM)1<IS>Q.MA7F[\+$)Q0/->@/T)&1_>CT/[V-):81W&$=HH3.:3<2B^85I]!
P4]124ZU@3_7&,?\82XF[=6A*J+4)>7?<%#9CG97T1<H<7A!:BMO4&'S;'4@^\_/C
P+Y5\=!X_T+YWL&ZM?VW91]ZT!YZW6,YR5IFPJ?KB<S.2A-:,M 1BC_":-E-8&@<M
P8@N8KS8QUW=-P_U<1J-]!7&.#.O!+%E.00V6MTBIA_+);;+42YA_0L?8_](-*_B8
PE[[47U6,WB3-2T!!CXO:$'Y P9A[*Y6,(DEA$Y@\4D<$%&CK3( _'PPI3, :7XX6
P!ZF!M#([,>NB0_3C3L5\7<8^]&)3O>W6KK1F1&D[6$-B/OE'RG^DV"_+S?T6S*]W
PD"4F_)^2R1H7XGDZ10O0*!Q6R #ZO/ ?TR!ZGITGC&71$'\(FW%[/@3NJEO7K5/6
PXCO2"[]U4JS#VR/Q+MWJ;B6&8J/$&9_K'R\DA=7[KLFI@2(V@*I<KJ1E$S7<1C_=
PT#"D(:'9DX?5#8NR4*^=NX[]XQ8ZG/7[0>?/PX9J(9>XD03Q?<J%8C8FI.U[#1(W
P=WIK37W-*K*.9EVJ%FE@:VT,3INKN#]&5JC1?!*&X[8E.-2\=MUNMYEP 3<D&71=
P(>";ZB;NHZZ;:\(;W!.T?&26"OITH"#+&;- %;R<0FR#JWP!I"DFR_L,^%D+,]U?
P?:\S[Z\5."Q[%&I'DLW65Y33F+GL3:-$,]1?+1]1HMKK1 %87"&75BWZM&<%K"U5
PV$XM,09$^5N@,KE:AO[M$,GT?6FXR$O\B"J**+7SGH,,DA=:.%ZT@O-Q0.G^/>PD
P-V0^E9[MS"+K2\#9']HJ"7/T45XF9W[1.+^,6^F2R#E0GF0\L;<#9WR_:U_6-]-8
P+_%ZFFX#/E)16DL5#R7=LN:)P)+7.C&KJ5ZHEO:%<;;3IN]TEU4M-0-$"+"AX.,0
PA5TMY,8 TI8-P/#9$#4B;.=\>UW&ZQ>@((*PY^=H!""G58C4.4>HHP7Q1#P_F7C>
PC90F?:]=Z^-? -K@9>45,?6MXW>'7-S\TN9F+S_\J0)A),?!%QS0>AIV?+OJW<>B
P<K$:N\HZ0W)3NX1%T];;YE#Q#8.GU2$4IP5RY]7,03&NP,+RW*SS!;X##QG=[P8%
PIF@&"+6J(&4^!7\E3P%UPTPAMB1.&_B_P5=@C6@%[NMTH)7?I^-F7M813AV_\HE]
PY]M#T1R@NMZ*-,JV&G8R6&J'+(T:K6EH)7";?4(CE0" UX=N(*P''OK"I] F\ACL
P(8'KG]\6D'-JSVYI8=LDA1A!9B3+(?L1L_%L)9)]84?'ZVS!QA7%\VXY7S_6&?D.
P;GNE2*?,34WC^S^P&\OOU*@LR^Z8E -BJY89L*&!2&_@I2!\MN]5*OL68$0L.).+
P$O.=PG.W>A?Z9.G>F+>6AOI<2_[3F4I6&ZXL@*17RL]*9_($24)[L\EP7-6*"T'O
P:TOX/V^_/AZ**W8=?U*903\P]BK=]5:^(Q4602@>R4K1,VIUS+P3NK+'-%X$<+^(
PYB06Q#>LHJV3C934_F];9V1JFW=7"V\LQ9.MHP)$AOO(RX2I0K/$Q6FV7M8:88ED
P]5-(6OE/"T$,HZ;84ZS7=3IQMY^A<I5>QY1.:NGLVW"(4/,O&I;NXE"5Y+,SW1L'
P15CC- #V+KY] JHYCA['0=Z7L\>X7)*JL\VQ*D@AI*LR1_Z206 0OHUR0%;,!SSQ
P/*'#FZ6'L_!;-FY<^ V2;#[:CRB)>":LEWS-R&%TBXLX12\/ZU0D"IC<-P\/BJ"%
PWUMOH4XJB(]XFTI3X>15K2I;1EO_J&A&S[^#XQ;'=',B_TGR5\3$IK+X>41-KA@J
P4J9 F8F2Q9P%1Z\DYQ]GW=EDKZF7Q3-%3=SFK6$>O.SB^96$&5=_MP5ZY\/@LMYU
P1L-R_P29 &!#K4G9 S'Y5*VI4.IA6 GGNV551Z0Y"&>\P;9#MY@;,8HD_MC V+:@
PT\-VZ"\#6GC!""\9I8,1^I.K4"Q#[CUS[.&#A#OD]* QD!D]&]:NE<Y=ET?(:++?
P/_7=MPS=XI<"T(HQY^2.'YRMR?N5.LFFLF!A^/W8%G+DCDDQHSUVZ]C0&C-9T!1K
P =+J5;>T^8$T/\&>$4V$/)Z//J#O8X@CQEKO]=N,8IF- O'XB/8*\HVA%6G]0+QE
P5? RH:>GQ<=4Y.WM"2E0#N*C8J<?8H>58[8%<W0TH"YKU@6,H*A92.PX=*&I;;R7
P6&*)9CJ6E7O2ZMO0$$H&KD1$A\_?WF%T&F QA;97"S32?[0A%MU!N$.!Q/'ZF3?T
PHU)I;WI,&"]N_E1;G!M!R+;_!K_\I/6+;^X6:H"0N(<L)3/6=$4=]7,HD(3[R&*)
P9W-=/$P4#^G%.AZ1(VGKJ*\3-DU#=[T\\O]JL3V;=YP=F>@_ GZ^4M[\<!+YV,W<
P=O0,PU7L]2.\8I$V7E@16<SM+P]#()OK[*B'K M[-I(S&5D)GSHLH.:Y@\(T^K+2
PQA.L37# "?1E'"'.&ZK1M\>IB]&M"/7QKG^S "%9D#ZCB2GL^XW_W.'#4<ZJ<;-7
P40IT^XQ.IAV4$XT<!=80$+"QP#>->#0DY4:'ZR!U$I?@M5H8C(AKJ98?KI@;M4DS
P1N-<Y\4Q,"H#14/U)=VN/G%CTX%7]"\XR/H_(ODZE_I(JK+I#%+;1"I(8?4XEW>V
P2OVNFLWS-RRJ@@VAJ#6UCNJ,S_(A^4 XO>9#+J8."QXRS2O1>K!P6QS\CR>"M&=V
P PJ)@/Z$(CQEHKW=JH(=&V0C.!>2PNDRN\7&IAJ WI=,WH^.K[IJ]M*J(B-7K9NQ
PS!MIT*;>2&5<"$<TKXZWB"I;^*(1[NH=D/_CR&I68LNPTXD>:S=C'DWKW@]/#4$P
PQ^RF$D8S_H3-WB#2N<5?N(DX7L+#>H$=[EKNP]:P+0+T7"[+JEOU;(,>B-G]0%D.
PSTK)=SYCV];V0<0SC(3@U&S13GJ'FI#$5H)/E9!:G.E MR(O"_'FVJ.OR61RR/X!
PIZ2;!4J $ON>"Z6UZ  UU*6?M@MPR]:O: A42Y@#M;R9B^O;.RT_DPX-U)N3 A)M
PO :#U G@#;VZN69HS[IXV1!5"IQY2.#4&+$?(;UD0_!N!O'G__F3-+D/EPJF4%##
PF4;W2#$#$QS(7,;4B?K?!T+LD]+D@K3,)/]SN:S30N]^%%M9$E]#_F1C'LQ #:JD
P$:1)G%I/#(_WX.KR>-B(X/P$G/X?4XXH:[!'C>OPP%@-0+0%26 &Y6?YH'Z*S[V_
P0J759U8+BY_Q=MJ""8B;X*SA39/UPY:OMK:?UY</0VDYF)7)@67+GM,/WZ[$]@\A
P78&W?71.V(6TWI=2]2#J^Y0[_DTA;-J:".-;MRN9(PZ[VCJ$ -=C+[^+G^ZLJNF*
P2JSM'[&&OS8X.SG=M]-8$[0*UYY_7T?*.], '.SC2E)C9.X::!GSRW\#;?=RKJ9*
P]ZG? SI["E8/ LT*3R#167Z%1''PB*'2LZ]H *$(6\G#10_QGG# QXDBDHGV%P./
PD1$OO6?[@+X5_JQ6NN-#;GV)Z23G62(9A/TQ]JZ-'A+=QHR0%!)/*:TG! KOL-G8
PH; @1GG3>;<=U<^[\\U0"' TZ3A,$ =?MFFMS]D915]N.W.4P2ZV<A(!T)D_^?U)
P(^Y]D.9%<DJ04@!2!B?;2",=VVYNN>#+O-<I2;^"1+,FW&,69Y89 K7S#1*5:WQ"
P#S-%BU)W;]ONI&\I^-=[!KK95'C(9D_TP#6I8:;Q.;HRG+J84-,9UH(CV<C212H<
P42@*K7F0S$4V"Y!V-#S$X+H^DXQ#HWT'-"Y_F .=C]OZ$191*=NHXZ9GK8BBJE[E
P'V+VQM%=$GCD/I I8Z_>"GX[4-$^[T,)4#"RV(J3*;6UG#Q>HL6737[#JE)YWXIV
PRMR 7Z8#))YZD>J*ZYT $5[CFLT'9K!Q>^%_QJ(L[VH@L M=\3R3Q63!78J&>:A)
PL'Q=U0&\_M+'5!QO1;\,X^(<S>@=;-1_2N1B<^1_3[9O5VKJY\K8> I]XH3T]TW_
P>=X1P7N]\YA;V72F%9IUI4OQ092PN/U\]E%N3CMQ^M(7M^C\?<L6S%:_\X\,ZBX<
P7CA9>['&S^,=@WUPC#KA0S!1(KV4IAD8)0V>[@D&K@R:PJ8J:LK ]^UH#5/&#OE:
P?K3J5&7-7R.Q<I$>_VR\.=A#IZ6\ /X%.Y@^-ED'<,JBID9!B1X>D8$'@O,N*B<7
PML-5-;V[D()K[M3&E]E44U^\'"5#M#^..^8";>E5*)V]P,8B=<^>A903X HK2ENC
P^GUC#H+-,%%_&^+'&=]8WZR/E/1?^UTR>,_>_ T].& &54UV699Y]V[)5/^+9#8H
P[P\[H<K\6!P^J7J;V@-XFX  )9L_9<1)<S;.YXF2(KHNW[0>TZ2T\555R-0K\"G\
PXV-@149K801_QBMBMS^*:CYFBT!:$J#KHC!ZX<@?$2/7*@R(H=7U.KNJTJ!PIJA 
P>4+!4J"-._ YP[51/M+E_^)^:4IR+OES=)*UBPEF*Z"$@=Z\7&0M+8J-_Y *V:3L
PW>H:JVTZ#>OF9A15ZA<PCW_CP?D;GR#KV_ZV43N>5-;)CR4J]7@?VLD-!OV'WC/E
P?1QH;172 >/4&7%FL2!Q5^'4X$N_N(LA\%AMM3L/>+4SFJ,*)7!'Y,:HU;NB#/^?
P?4_"CJ-PROZ8)=B/?LKQ:,/.O08F[<X+P*9I\/X"+I@@2WWCS%?=]4;5B:FC<[VF
P*<;J>7@DJ9_8LZ$P<I2%,#7%CQ<?0(,]]1(I&)ZT<X5?N]OHNE/@![DB<^NC..8H
PLZ5Z+GO6_M\2P(S [V?>,?BA@]4_]_7N -BMT--'"P.K ;\+0V/_,?0^QG0[7EP;
P[2MFOZ F1L<?<;G3_FWA\&(:!TJ+KWGYA[78Q89H[$#3C)6-4M53#W1\@-2ZK?DF
P$T(/I1K[)O>N(WMK<BA.$,$D4RC:PJ,ZPLJH\+=6;FEV-6[/$>YT>I'X><P-0*B"
PZ(5%$VH(A#,-)>(NAESER&HSAQ+A=NRW*.S@X8(P4?T)CB*8K06%RA?=L+7,8SPQ
PUF]?DFBVI:L,X3+-)4:TP/BYF;([H&3M=0W5&+L[$!<)0GK12KKUR:FA_^;&NIFC
PBVZ_81RB>?3LPZXF(H.,A,_#2ZOI#>S%HM:9Y#2Y@A2:#L1GWI#(*2$MJ?[:?E.1
PVE,)>"T]VW[G5'!+"=[I48! &@R6MK9 (N*4%MD?-TM&=)KEWTW@6+F+;9+=&"J'
PRS"&@\;A]2<;R9S"L^0?'R,H+1\F0-I^6Q*]$'%]NRS(Z#626V[+Q='(M9H 1C@K
P*=[A%ITKIJ*+&"Z7D>QWOJJ]M"$*^EFY!KJ\%TTQ10+#13.!G\*5 N51$OLOA)LY
P&\T/E[T/[YW],<RZ,1$G%)Q _/GE:;)!]NR(IA;GC,DU:).)ZG8JMGEW)LM[Q[EY
P?6H#@(3\T^GN"N)M'\<?5RU@TLH4)S3"#0,_D9DCB>!&>FMXHCAD'Z(Q9,/)IF >
P8&M7D_M:H.9 Y%_(Y/FK194C",A0ZOD'DLS7H]3*PR%W(1NDS@!WVELZ$9MTG':@
PZ9[QHEUPV0__<)$*S)5LWFAMC H7T,'FJN*>S<(Z!2LMGI+Q==.O.M*K#7BY%= H
P$&29!%[TZX%JKOT;=3"T(6#6=% IP$2;'D('Y%TPG7;XD ESNH,Y&>+ES$X)-TO]
PD"=8?S68RCOI\#Q..;AX+*EF^&,JK8OH!)5(*WTO:[_BUK$D%L<IR_?!U:Q/'5W3
P3SL*[-RB%\IQ-2)00,Z'S4K+\1!@V!<BT=CPGTM^>R0EG<YXU]O&@M?7EV%':82.
PS--]#[!G2XBZ2R8Z;/<5I[;:1Z^!(,?J [RG^/ ;/#)C!\@=^",0KJ_*P"B"E.A9
P0KW>1.G\Q;T=96*PINT#6N-@\HQ8H7EL;U.P,A9.$(#-96EY65\-U9&"#C;$%T!J
PX4$$U<5RD5I-;(N;+X1<Z$/3X'>)%7<(^D=.MV:BR/QU/_T;93K/S]?D?A[!ER5]
P87E!"X?>? A<W'5$=4A%#0W4VL:6WB(7J],;/-Z(9/P*;C[,$"^^S]LSP3=RL[VN
P*U?^-3S%**AO_SC,1!=QV\,)"1H"Z@K'/%)P3"A%O3RP'RX' "48;USI5LMG;GI^
P2@EZ#]B/\:8G93KQ%TJ5D*Z7)'79->U@@1*,R;B7@27$MQ8:WD_<2&@(4+,$0K#M
P!IW;MIV/WL6@#? /2R7$)!1DL9])QAT)9%P,:]05P;Y20\<!("4'];2]T,,@7Y,<
PE6%Z>^3.,OW/+S]3O\S>VI"WD,;1VDX XDO;O'RR./?+Q+969]WZV9]+ 'R4#)82
P9EP?G=D226 33/81OH=WWLAB7G VN>^OP;(#F7\L.L^-L$?6 :11LDIHZVD[TKWG
P+_GNW8UFI8/L]=RMFP4L'O/2X__+R\M4\-HZ8E(IQ+BD0P9KJ$96ZS&;;Z3\T=;7
P ?G/E$X+WV6YXO>0;6FVVIW[J>Q"W>U Z<ZM*--[<IH-*?8>_M@;NHDCO4)*_%]$
P-L_ EN_MCI)/GY?^#[\:QCXPI I:P=L:EAOMJ$'5%:-U8GW4QU,<+;G9<(G7?XO(
PGZP/%9 D/+IM6ID"*EH4 2Y!WPDY+,@Q!MM024>+E? T?S,.2:1Y&7.)+X]9^TR.
PB)4>^BC!NQ#)WI&-$5B)DPAY,8&["$U\EAL8Y36NOLY,$MID,/V7+PQR]*11T<$N
PWX''?R@^[$*E6.H!VXZD\EX&J??.YAR> FU+DIZDT-<$^A/Q=8P$ B5N2K?0/E?P
PG!#]3<4XV$QTF#E4XQQR7&+HN @Q0J,"TP('*)W\E;PUS$5"D%&VDC32_&[$.#'%
PV!+G4%LEJ427^A$7HLKJ?8@%?7>^O@"_MP3<UK7=[H'2*< 5*V1$18_.7H4G' >C
P;/'T@F,F34#HQ[3:L8F]62"8R1N:+8 B8F']8MVD/>PI4Y0RR(4VV+8-*+I )<?E
P'12>&V/8__5(*Y<ZIQJ,QD*W1][4HD)%.)M@7>O'VVR*D\@/7F[E!W&_PB1[4'Y*
P4<T]+2"2JDU>8R[![ZYXI#ZZ*=LW3BIU\#W>6+^3,"DI70GMMO2P#\TI7X]1M$"%
PKL\:;ZV,#O"#L<($Q6_RY"\=]9T6;<5].\*)Y,!^#U(;/,G9T:2OOMKX\AU:SKQ*
P$^0JWPHA<Q ?.'\"<:] (T](IB<+9?_6:]R#II/K"0/+9$P0]#*Y2#[^:P$WQ$@.
PJP)3J9QMC5F@_@VHJKBJ."1 Z92UU3D6+^.1$[DESRH^8I\I*)A)& ZE,PM?Z0K(
PQ $N_77#%"-S,I%N9R;KPCIQ$J"#?1(_ZL5310_<C0\L+M304;%HDF!QWM!/5[6R
P5<([8.VJ+O3G/CG.E:%&@IO5#MZ_G@_$A"[JRQ3DPTQL-Q/?5M1@N_GW#E;92^NH
P-ZE&"]D)&F4O6EJ2Q4.;Z_B,QPAUWU0$:>Z2EWI/"UCL;!@L4XQ#EG)*_9EF6>O_
P$:$<].:YU#NZ+*.#E@!S#*V,5[#4L^Y9.0G,SPCS?HE<.I-^Y7:&RWAR2M$6&SC3
P'(BJZMMO"@-V(VQ36L7\\KY_,S0_UCYH\BI7MO(,G>#%)WJ6"6,".>RM>F:.-C> 
P:'J9[3GU@T*8U(DW =;LZAC8W!*D#E04[3:9JLE"-]T*Y'FE/T&WGQUN\WG!)*/K
P5,/SL2)?51Z#8Y%1T^2MA=O9G=V?60 TV?>#.N,HZUXR#R")-!*&<6^:CKOU^ U4
P8HDM1\OR)1O=X,PE0N(N"X(^LGPXU<AU;PIVEH4SN:?V0*P2:_)KV("Z!$BJ[!F+
P?P$9GUV/2@I1Q[RSI\Y=+/D,HF=13GH!E,#.]&O)]<HJN0GG;BT 9RG0-8_,I+-W
P3WDVN\NPTM^ELH,5$<-48@RXO^-&SL9Q3V5LQH ^VC7X,T3U1]K'V; :-@<7&$=/
P92:+@Z!-=M 1PG]K &9VQI*8_,P40S$%73 F&G;*IV8IGN]P^L[DQN$H.*IT+Y%2
P8>7CFT9]$MS\WA8BQ*2<IET3F-(+&I^08DU8U HUWHS4\D*_IT*NH&) <?E0\<81
P0/WW'"8:C)YB-G?KP2OEYTG63?*>Q2.<T;O6J=8(<5R#(.AD 0;V-"$X"77$"*0"
PB"BOB!HEM;I1 X_(="%X*LER7S[YX6T+X]6&DRD]U6@!JZ4*\)_2C_&C):!V#\;O
P""O$UAX;U%W\=)\Y'6)H4TP0[7:@RQ6PY,"ZTNDN5*>&.\Z1<6+%HP0R7W "[(:L
PI#P!*CMDUJ"[WRJ7(1G;;Y;BQ[OUUU8H?;(9S--C:NM2Z":9C%@_6$,BK6I:M&P 
PX2ZT$J<HBJE!_%37G%TV\9( !*9G6=)51%"WGU7[IQ=\$!L(]'!<5A!8\,1LW,G4
P6-#VC=H^P=,=;3D%='RJ>X)P?*1B>3ZZ/M"-PVBCBK96HT;#DSM<!5GJ5=66;5!M
P\0]<[3F(7B(K/Z,8AP$)@4^Y[NVUIU$N.EGA6_'D)J=PMGA0["8M9N<CCOK.D&%3
PQJQ"!R4J7Q.Z+4*>OVD^KP.JN=]-L$F4E\-5H[6/T(O_(7B=W@M0H_8?H^WV"EO\
PBTV;F]AF;!XK?K M L9(Z R++A;,A&+^"',=G()LCO=ZLB_F=2RQ3B^+0';ZDV^2
PK<95R_K"F)@ Q^R/8<_&Y9"WLJ]ZWQN1+X_)[P@J=E/D"6$$/1;>%Y#G7C&LZ<RU
PITQR<B0LTL_*B/"^\\\VX<<WPP/56=Q0"_MY9FO9L+YT,ZLZ _F0#PC'B>NR_%*%
PQU.*]!_.P 1UV%W/4"$SJ8.1&3R$&AOY7]!T<,WLV&%IT(D4TEM7EAW1^^UIHIX4
PIR9 /3>A<'L6'J:TS,'<#8WL/2W=R;> RKP!E55L1S[WX/BX\J!%=I^]J/DDYG5-
P/-&*1"#QKX'.PA^"G##[.SQS5;527%@R6$TV1Z_F;J/2/[3>C^V]%ER(ZA\PE]IJ
P*\]2L]04$Y)P7 *M0D0')7TII-H^7B;>KN841*^DL 1C22*+?JS:8G:C*%3!*23,
P'V_8Y@:9C_"\P=ON?899D[(E(#9XP&=(D!&9YEO*!]R(4@0R L)6_RN-T4D&VJ#[
P$\PV8CTN*GU]EQ>M+L6=]I07!?FD^]$U7=CHJ4.R11(_*,CS/4KM!KDO +^(H''_
P/*CALOO'Z9:5AX]"^F)4\/N$O)NR-U">"JP@$X<'.A7?CG3R7?T .@NQ+"SW$ZQ:
P-I&SCM;?)^-B\BJ<5V@D0D#KZ(_R* ]6 "+X$-:ZMWL37/QWR2D@>ZL"B4E:<9$0
PNI[+FP%H6]P K@K_Z17J4SM60;QR"&PLXRFB*DA"ZUTVAC:^#*S+5]3*E__W*=WZ
P<JJ,X(1^UB7LQ"%@AV(8ZD\0\*LBA]('6$36]:&6> &E/4LS,G&>H[X"5L?KC09;
PN:G5W)[]'M/<2$>[Z#"Z/<9O7#*B)3SS=+2P02]68]G@ <U@PA259[K0<>(T5)NT
PW9H^,B\\(KA HI.,L8(B<I(P6I\&1@GZ0 ;]6JG->#(/)/MB$62-NL\X"*)1&HM8
PJZ,:U)(M;R@C=ZJ?*!AW($MA[NRE+*KDB0#BH%E[\SRLFE:Y<=!7MHWYD+_>$OAW
PN&, -'\GX<;9:5]A#ZMHL";XAR^W 1$C<H*41^UZS^I< QCY,?X,\M^?O*!LSA@+
P!6CWLKM*=Y6U_'9\=EF/5  Y<ZZL!2W.$3,W^^X&V9DS:L\6P6IPS[4-[WCU";7%
P]-PXR-S>G6Z>8:>X9#Z:M\0H_$U!C^08HU0@QH=GYVSL D F('AD3[#]$-1X<62A
PUG, >D)'E!MZQ[PV X<H(O@V.RL0K,\:O=F!ODQW.-I09@3A\=ZPJ%4I+<X(G#;B
PA24G0MO$4M$$=7?T U<5DI4:RNZW:P0&65NL7PXAB>NQ^!?M_9Z!!]TL\"%-E^JE
P*>@ 5^UZD"R*5$OW[;:YS-!)[7A_S\N8PQE-S^UP0!)CK?<9?86I.5QF/B0$0E*V
PC\[A%>J4P&>>C,5IY8O2"$ZB%<  ]XJK[<+7\!1-<J9*8JB<V5%H^#+TJNUZSER%
PP6$D=_\&<=VT/%A\XB+)7"9&+6,370!M8B@A#I3DZ0X"N_> U_A"5QQG2IT2K;H,
P."D6OE/8TZW\* KH23II Z?I94JKTF_6H0@G.$4-/8OV*1&L/$DR&F \J]"_<7V 
P/]B)]0,&Y&"TG93J]L&#QJMQ]+W2O%G*&J873+1W_5_KGW;/5P+,!C;# B!F"_2R
P<_WDK-OALP(UG/1]K/!+HM:V '[ 5F#\R<_HJ5I4G4XZ^:"D16MM!9=AJ:F[VH\8
PIW0--(9#A+:>3:6Z7=RKY&OM%ADP\M)^XF-?$S].R&80^O)&^^\$RDMX[XD40Y2#
PE M<NUJQZU7H9A*%/SZ0TNM#4D&7UH&%0H05 Q [/0VCN)26?X+N/+Y!)EWD>QCJ
P5Q1Q"_6+U#*P@$<YX;8G$F\NS]EL@OTJL6CEA53#+F?-TRZPUK*RX*G@MZY)S5?+
P:EFR8J&76!2]_*,87+Q^=W4J&'U(0O =A,O\SZG'M91*U>SSAIR5RS^TD&]MD.B\
P3GC*J0<:J"+*PK?Y1Y[L?PY^^0,(!W8AIA\CBU.XFGD#!4@1E%2J5F^\/G'QMI-#
P$LBF.[RMUAYO.!"4% .UQPZV65@<B:8B-?)$&2X7E+PHM[YEM_%Q;-</(^PO(B,@
P20='UBY<R0Y4&@F0Z 61+(J;JI>2"]Q+&[C[U!M<V['D@3(:/(L(H<=\0KCT6=LF
PS :S7@4#S:M?*!^,30@D&JE2G]-/R=5GSGDAHZ]17) '_3^&E.2T=%!1>68Z+U>O
PLK!%^LNP?[TC?,K(=1-JOD5@+4)I"0<II#']DA0$^EFH\Y/"!+\;\HD(O59 (SFH
PJOJ&)<2^1-!RI '=?V3:OG[2:6GX;7#V@=4U@TX6TTWSQSZ.B1"[(P:SZ7<'N&O$
P9MO'363C,+W+YQHWP6Y.%@KY/?;H/+AU+5U]$O3"O/ZI96$C 30R@GL)\&S.ROB*
PRJ4[<85(-$,7.1UZ(^)%XP,[.B:[E0Q<W/?9',K7Y62PV6>IR;F4!W]-@S9E=+ZV
PG^^X2*HIW,*XID8NN]5+5#UH-5)&N.3Y0\JT7=/.M:G:7:P3&WJ>4>"\6NGX'W,+
P9[4\V6]S 'QLJ;2[3YIU&E^T0HM$1A", ;D\!A7'/%$1)+D"*NK&+P5: 1\WU7')
P'+YGL!XY,-&4Q-'11ZQ]!+1X*W8J4>UOEP'8@@Q3_;K1TRL"X1-%-*T0#(V"*,Q4
P_.>%FZ1UY_=235S)9Q),;2,Q'$D>Q-:V]955%HJ1/-\1_%]T(,:^))(6TV@FT@,)
P[_.6>\#UC0PI1HWF]"K  QDW.A"D^_R&:T'/99#@\RS6D,&+9HOP(CKN@F>[V12N
PCF!)]H=.''NJ <VD(<UEI/4HS!&ARJ$-6=V'2:@]Z <KAM34'9AJQ"76%DUI:\Z0
P?_KLAK-BZ8M-DW0'B)6$8.)$1NKF<J1I(;SZTI(IX\I'.VCCH,GVKKBIAAR$;)W\
PZ[,),G\C9B2PX\T%O*EG80RG7OHQ_D>?8W<%U_W3E^L;_FN(/;[_DA&(EE&0;-O;
PE]R;$20LPL,P(?CMQ%'7_N>\ENZB%RY 'EX*)"EA>4N*/P-J![PN9WG?L-" %>X\
P5L=8F;01MC%^11G+NRCMAP+H&2^1@;XTP[03H@GQZ5[?N,H;8N3X!F$< F^%ONNX
PXP#$PDRO 2"7%\Y/-,!6D/62W9]^O?7KNVG#/Z<$V.F 6.48*+N!E0."_I.V-+_I
P&25 RZT%FYR];$M[&1MAK.:NE'&+6JRLB#&%3EBW4480YH)Q^M,JW!O^XN!<U[ )
P-LY_Y49!#4\P#6-W(X3Z:WSNWNA1X:P%&U]-5&%P(!H[KI[EM\/FZ$^+B&^2=NLH
PN!C@Q,%>$(WZG-:?R.N0Z'@T?'TER H=/9(,P__EA4@'J;>$=F_EY]+@;PA-==?Z
P&:XU6G,64^DX&UK /PYY#B*LQQ^T1WU[H9T0A8MAM.32,R^CPWW*VS]X+9;-&R'2
P[\A-G.4E6F/.INM?RY.6/;)M$1VU^/> 6?EJT*E^(\F476C(;RR=0F8QA 3Y,#X8
PCXM6VN"F!SA=B:/1TH!T1O;-5Z#85 JQZ3N#4QS\/K=TD$H7F+^+UKSG1_TA_:#1
PO%]%Y(<&W<EISB_\5NI.%V\LG)^LD,VN4I=B_).<)GJ9"DAR]6$T!")37W80V1J.
P5=AS-/ZDRTX7*?1>Q\3#1^L)ZYZETY90S40GV7*@N/A[>36&6IO>/YE2!A!(+1!^
PM,"S\7R:%9QSZB^V_]UVNP>,VN"VPB*PJOH9U(*  UX'B8,2<QR::^(@YLP+?UU1
P!XA;FV;S/6Q8<# +X_\0A/V2FE@)/#.!6*ZW,K)9\:G%3,M+N'G;F[$G.87WGF,Z
P=P>H(8^</'L\_*E2)OOKYU0_MAQ3WO8KG+=.VX[6-Z7KK@(Q@=4>T:[RC3/L)TN&
PY0QJ2G-'O?J+(P!?"_!D;D_*<=77C02ZE^H6>#6%'O [XF6Z6?8CKLM^J!A"(#< 
P%YH:Y.#F<,9YDE>TB+&:I(?-SR#58%!S*UN^FE_#'0J0<)#](87*?4<X@:QQZC9D
PWBW_5J!X\[KQ7"#]4 _J_Q9J,^*B5/]14"7'?U-(CN9T3C2"1DA50.C2& @A%LZ>
PZA$^A4E7\Y5[V!4*#KD!Q(9(T&_#:,<AW>W"9^V*RI*C=TR5;*LP"*?0S\(/C8@X
P0SL'ROGFS-.TVV9KH:)9L<'P;"3G"G2A_/BE+FP4G)5<V3VPQ&4YN\*UQ(&#=,R_
P$=6#Z-DVCD6P)ON".;#64RYZQRO2=&-YU50SH!,ADWY* ZO==KY!YUYX&:!/C>,'
P@/Q6R=4;<V]-2F583;?C"-YU4:D+S;;U=NZF!"&0X&#S]T;=AS2)NQ%\5@1T0JW2
PP!HN-@JA)S,%VCF"9O>-->1)^57)R=8*"@8B]CI,!8VB6\\6*[SG"JH>IK)S+@2R
P)D=I9J)V2M&N-\,*M0(Z&ZS_LTL>#K#%+:_XTGK28U)@B2:CH<I]?Y,RK@C8A"Q2
P*>&H]@F5F;_$4&:>F0V3,4X:" (F.,2;N9$3$UB<LPB T.YJP"K\[.VH-%!?5EZ_
P:\6^BKD87<]"/?@)N^5Q0#_"JV<N6\Y5)]&KG7T0G6G2Q@Z"^(%)[+Y,/;F$_)?<
P+G2V7PERU%%^Q\:#0#&FZ<,[@"*C!&Z%YJJ4>!$&>D8)P_.*G2H.LI3EV=A145T!
P=VZJLRJV%H78N>B\C MK17E ?\0.N\(4!<(^%; 3W N2$)J/6K1:*KRU(Q07J"CA
P9)>JH)IYVZB ^:2ZO6NM;AS/*)73DS/8LL@5!D#%Z?V[4:BN8+_2,!_G7^AYBYX(
PSL(ND$D^% &M-J<,-FCJJ14!92WBD?U34K*<=">_XN(15V*7/_;K6M#A!G 71IJ4
P=S"O_4H$&UD=BK4=/]CN4GR6(#(:Q7#?PM+MH\7OAPL4A!-&TZ+"$%=&C(]RW[MH
P/:2'HBLODR0M'\,6!X[A]S#FGG!.RL"R0"_&0:+/W-6'W[%'C']J"!(Y52CM3AS5
PF I.:LQZA@!9>VM7;:,*=ID])TNE6YUE:ER058,E@LI#OU=9H?+>L-F/.1FCI:4D
P/>N(6)NYT,M" %Y0B3X05(U.%Y#N?I6>1XN":2X$X!.8 \CR-G8,Y18 ;=GY?V]1
P]^645:Q7;!.O?3TS0NCFO,XV2;,HJ9:2@'S%RV]G7>'J.$I'T"T7\ZL>$(H.$"@"
PFX)+&<-QHU3M&[*H-(GKI>2':V:.2MDPK<K/(S@QJX_KJV=(M]<;/>GX=KV6XS'H
PMN;+9 ]8$L3=R'/!LWM19WTK$JN&2&;1&?"R4J_NP)'F6JL!XNBS<X,9WBTT 8Y^
PW;Y.K8>^%X7,+8#0L"?\&F^.OQB3?"228A[D+W*[_FL'A%(_R&*C.BCW,IA'M>K]
PMJ7BE*2OA&N03GAR/]Y&S7ZYIYQ<WUV,&DRCO6**?*%D@ T1FDJ1@A^B/K=?9R?G
PH=$5::'USES<EMAT0=R53,.[4U*<N3D!DG 5WENQPGLV#9A<VO5IA04>]&-J%*:\
PCG (2H]XV@1,A_W=&;HRR8)V-!'T1'"WBL]RWS@#0A!<)23EHF<J&//_[(?8I"G 
PR;N<J4:>#0K7GBSD]AK;DQ-C2K=D3-2AKK=N$7Q: ]Q2 W. ;"-P#!(\.9'$^EX#
P\E:U:S5Q=PE2$6IUD*MME>9271]?QFY5X9D!+ATY\61&D_JB_*E[:@R4R$R%BX1W
PE*U^-U_NXA"6=="HHBZ8HE' I02ZMI: K#WOX\M5_7J:3?A$7, S+OP7@,!HBV$4
P>P]8+X>_BC[C!@H471@3P4\SL5P"J@\:DSN-F9%O8]\;$XJ>> QX)A)1Q!@6PUM[
P5V-7[PM?B%TQ'FP*>&I'^B;WP4Y*@26>]*)GSJ " NK7E>?^;$H3Z>-76/>0%2RF
PS)22&(BJ#V(J&;T%*I[\2?]7[R3NC%PNW<D!\)W^:FSG1A&+%R]*Z&<]4'?83Z*Q
PRSR1:>?EC=NG$"E=*.P1+NL[&"6Z[E/:3<(.WIQ'"=)'HS/RWI*2 [RR3IN_G%A)
P",Y@*PF=^,#FJ:L^7BC1*(=G%]B-WO[2J))1SR@&VNMD(S3_;8*KWPT:N1^ETTZ!
PT,]3?T %DXH'X7/7F@#^/ UMSR@E3FP@S$1\ITG4M $<B34 9%_3R<][8< \6,]%
P(!=I#P8")E:]A2U40HR2 6:)7-.KGS:B%P/ I! TH*^/"-.[/EC+UZU0$*-Q#PJ'
PHA3= Q[*2(5\4!+Y#V5F34 3,@HSK+-=2(*DQJ6\$/B_I/B<)U#!\/.OYI1#"(OA
P;!0UZ,?E*'&;TJN/S[>]X?(G\T0GN8&L_28^ D K'QR/_PGW>;4K:56>'.":5BU&
PF3J-=4_-E?D(DCAC9<C]L>D[QG^;9,3JX%-R"_01VH<+ FQNH[/,B:[ME7W?/63N
PDM+SL.ZUGFZ>-*X]<X7/^8*_"+/>(J#G $[<NPMVH2P3Z1F6[*"+UUWVK1,;"QP4
PVLP<Y1\Q> U?=%.&YZ3G\Q*492S,B'3[L9IMCR$NNKWIC!D+GI2Q-)W(S4PF<C7-
PSH0-X(#[U.!,;1QN$@\]GT2<M=9%)3#.IWM1*C/]%Z"NIR KA$.LA968 $R=(S%!
P]/2C1,88F2;[G CJ5QSA%2>*,3D:#0='5CNZRGCJJ>=W]RL[BI0&Q$UO@#</-1E 
PIC/L:\,SJBW-&Y%,M$@/FG*$G:7\HX\ 4H]" 0$<R7QG7:YT&2FK3>+ZJU]Y5)(7
P% (  W ]WCS7+\PJC93D6;1CKU4#*8T*.M,W..XM1<.X0U9A#<["_T"%<(W:#^#=
PUL7!_/W?,/]L#>0F/3;_6A,]S/5WMV\WU^Q2H(6>X#PGSN'K!HH7?$( K"<^?*\N
P$]!B0&^,Y0KY>CS47MDO=7C[B*5ET]?&>"O%58*C('TGP43,-*[]#O]@#B/TF@6 
P5,GT?RR6.Y+.*%FKFB6B")E[W(]E==3I4GMZ_&:5=&_SP:$II$-#9Y65\5X&>S20
PL.M)=G10B>@=I7*]JO$%%PNTCJ"GVZYA_!UVO4T>?CE'I]\6P^'9@?+6<:9"3_RJ
P4HIV?1G'E)?/H!B%/2D *3C 10_[GFQF1CR@@" ;F-]+2;Q1,NY5N!%D]7S=$V$S
PP"%Y\9?[$_& 3;/1.MOJ+ HK?X&V#3%=E2-&.]%^C45*#PK@FL0[<X'U("5*5B@L
PX*C']?'#YU*S)Y:DLXCI@:&FKB+/5\&F:K*J2ZU? !)S:@=B%>I&$2O [X1\3X.X
PS@^O'+-&+$?=JN(@YOWO8LIGB@#+03F8ZJ_.M<(<IU(O@\\4]0XY(ND$LR+6MIC,
P; --=9B)S/[:LP)_-5Y)=?YW++ME;,HU!KX@](N/K<L7KYO.W4$4N"<=<@JQ:ITM
PA&,=UM\E/1D%%'G58?P8]51MU )DL[@ BD,%J(& WR4[YB? 2F8*QXZ(YK@^-0TO
P#?_=+X@,3!WY*W.CHB^'>F,!H!O6^%/TWLSG!\5J-!NHAK&I1*F-VX! CAU4V08Y
P^*_Q)NH^B.1@U$'@E3<TG:NEV]FC-W22S-VCJX'(NEA$[R<>&KQGC^*[I9[]DGI]
P&,E>%:@)M&L*"M#\\5=1)82.?MB3X'530\OD)&JO6%?YD>]B<CQ\)C00,*O^G)M]
P!Y@LR 20/>8$'^$E&N+5DG][X[+I[;4]#"0V1K4?D44OZUJ[[+3'>(?Q-".?$)DP
P*#GS* 0@*/VA-,/$12R8C6!_(7K%A:JTP4.K^5W'V-(/CO7%/>09Q\GXULA!"FEO
P1!Q? QW*$SR$1."9ON0_%/=IRQBI3GO/M)4]JO.C AG,Z9^E9?0TM#6=]R^F,LO<
P.TFT24^7H#_1]F+N="X]E1U>5\L-;TW\S[#"K(J]BY<AW9W\6,+-?19R;#0&0*>1
P %DW_O604DS-=DH&&U*V+2OO/J$/H*O?_R=5/X7![%KV9WG#-0#3/@\@POVL @>M
PW!$JF-'R['C+IUPZF9NK=HF^Q_I$_P, Y?2&]"# :#ZGAAQ!X^JPEL4LA@TK *"L
PSLAU14S!=A3/^QJS7BS!4H?SKA#Q$5Z%EVPLJ@\Q4GA<!V^1/JE045A1T[@"(N;8
P^3/QL<5:)?[ Y:J0<VU$V[D\WVVX4GL3&*G?I871_$-T:VL5C)DX*ES".:#.Y4D1
PJU "+1</&ID+ KQ.#HW9V6D>J<ZT][J!Q),^BJQ_O%H_Z^,I$PH;AIBR]7_U6@'@
PSHWFW?;L#SP_E7"/(>B>;5.5V\$PBXV0>V?1+^-LJ!'J<."K:* .4=)8P>#5TW5W
PE4]^$F["]OG*=LG=K[#:UPD>6&$]V"I*QO  8-/@%;5$P;>;X7IGEQJ/UD4J&_::
P1_>YI>QH+1$Z\Y=GF3P84_JW+\^'O>M'T6V1G:Y=C 4&,+E8G+0V> #WPK9J:4DQ
P/Y!NG<)@D(#?RMF##ZBXO*#J7:UWLKYXJRJK@67@OM8E56"1@,K2G,V[0]CA&Z"2
PV$W12#<6O$J-&[*]58;597Y_7>^69LJVBNV\4_4Z(8&'3QO)$!!6>*_<[_N@[3^9
P"KAIK<:7S<F2G+!I(#:S5A7A-P.OC;X@[VM&240BB2GFD1UQO2?+S]<V&"\* F&.
P?)7 L'BC6G89E.0W[F4]+(V&&4("3S@X=#.KBHZ]+5?T5=]VA+IJ'!\Q#6;1E/PH
P6J(L/-I.)8HTPZ=PX,]2\V7L>R;>I#64_FO*B?$(]'A<P^!][;6R(U%O3XOK82TK
P>D.81A!4G@%QC[@"_4<V:9!-;MVOIYT2-.K%3A[-X5?MK3;P>;4+G ;N^ Z/PAR]
PF'[D/42Q*D'_V@S*Y3J LW5?):7'AZ/E^/7&JB\01O8CU,+<VA+RNTBDW?J9V_* 
P=1H36DPD2UY4+,D&*U7ZA?K65[V#XC\KDM1PO6C9,PVA')[.'[M8^U+!E6]@'2P?
P$9@QD'60]XA6]UWG\9H68A4<RULWN&A9^?23O)&MP .N>)BX3OZ%&+,6W"(3-WL/
P?N6I1UJN(WC399'[:B*Z7?M<KO/=+"28D(64!%H="IL&GGT=5O^%D>9E_^#.\$X_
P#1&*]XLPH4AL0'],16R*.3J,+MKPI+@T<&=P>:LU/JI%%QOY0IL=E^9G6BB&BV+<
P$O/&.J+@F+S=&=I9X]A<5&:)8A^&%SP5C+I#H?(]7)/+@"L9V(+D(./2*Y)>V<-Y
P2EK=TKRR:.)5T4#-AO8!S1UEA+?P<:-"V$KEJ&:PJ:]Y="(6Z0_$>D,#:-.-=(V-
P6GYV;&QQS"7[?4K:/+2#_&M'\QVZYI#88K=?M.W*Y>E+<VL@3V;P\:ZZU:'B["V_
PR@?@.585A@;N?Q=39<HSR?N.UK18*DM9SXD17W6*A-JCRD>G,WI#EB76<LP']=R'
PSZS2PCN\1HSWK^N.TOS>DVX7S.E/%&)&WO+A=KH=._?E-'V1_+^0>%9Z)'.9="\.
PC?2IQ=>'+_!6%*7=C5*9D!U4CFUQ-'PX>[N:EOZ!<..0R!9:G&WD6Y@[V/Z5+OWA
P88\[T^>+%&2X'A.2L.-E+A)E%J:I;;*J+]W'YQC*DZM S^18=@)QN5*#.NA@B&&]
P# U=[&$!?7-*5AJ^0D*QH,VCY O*PUE5R0?=R:&NL:;8<C\.QD;0RQM@SL%YR # 
P&$#PR$_9V8SMN;;KU"8[>]\?MU/J0=LR9*OU3!&#I-O(=Y#YM7.#H!C^]6LIJ6E&
P1J*/J-8R0/=F5@7&;!"Q"+&B?GP\[_S+U1=HXB$/Y^0]!EVI7V6Z/J9_3@4+,*NN
PD:90C@S<LBP%FQ2"@E7J8.76W?Y>ERU'/2LU:;O#OPRP$,C1B#8*)7>1ZB%G44=_
PGVD*,6J$P#4<P(WA+?O@0&<_R&T_:K3"XC<+E6,'J*59NMP0$,N(A%6YPGGND_E.
PU^S"]1YHL:W@6A<(%^M1KFVT_ZO5G7R+(W"'9;^E!R-M_7-VC(,'7-4^DM7G]QD.
P<V2)0FT.GC^CE+^Y155712%=&17O>BWVNQ"/(R:1/7FV+".6[S)>F:1W=WPA!X<%
PTGX8-*Z)I\,0#X)TIM,#^%"@$SDJNL*8QFSH,8 %#6!LX<2N<4\/=]RAF/C?7]SU
P:EI4^EP:71M90%G9X4M6B=1MXV\39XM.1 N\\T!LBII&-*6^QPV3<V!GCKSKQ::U
P+5C+T' <5C"(=G_SFE6%5P:$@NVB11I:T;$KBCUW9EX@I!]D)Z'\% QT&T]S*29'
P*R5C4H4K02>-<2[I*<+?#<:%WA#OQHV?)Y]X&-?!/*(;,]]BX2W_F&"Y)TU4+%[<
P#4)GIN^KB-5QZ6I<^)74OF'Y*K4V5ZK6*&6<96T-AJQEZV*:NZNE^]=#/,?AGE>J
P%_9TZ0H\$\EQEZ9!"Y;?Y$SO^#F02GAE8\)A2M\I;\AH7OI5DC3IL+;S6$7#]JN%
P[T>[Z:Y<;+#F(\P1C%2>9>,L!$LN=B8L+*&N4H^WCG.? ]+N?Z ^DB'\6K-P<H4 
P 7;@V4J\0@?A2E/.3'75':,G]1H,1;U?6^?K^#S@CK'*.=2^#'+-8A]#S\RU&>D%
PZ QMEKR5Q1IT6*[XUF./3G AV,$GA[0B4!U+*9P\FL[@7G]-AX,9[L3^.R*@B"JX
PYQ:T?9/0JS3H;9E[C'-G7*'( "MH]M/PGDC>;7AT*0E7S<;$@DN\?%5X%X<!HS=T
P],H%!2%G\;%&>)[$7-!9%O2KS=)FM_MI:<@XP?Y%9 E_ 01!83N[\<BY=T-$3].,
P<[7YJ],]"AK'6F%LDG O[ZD)B@ )<X\E;K0XFCO/<ZY7-_FR,P?OQ&Q*P@WS1Q\T
P \#!#^?)S&J.*,8_^F@3N#TS_2'GKM2FU,@F8B_6=O^38V@MJP<Z8]VO=0;>PAZ'
P6C;1N(7B+*_$+A#>TA%('GZ<#P1Y<:=?KH25+EDJ^=1,3+4]F#<F.& Y7E:/P[I7
P!F10)<,V^AXH7IYI:4*_-,QW >Z(#/=Z%%:V/*5+:*"><Z$0H(&O/:P?IHY! +"S
PV=VQ@2"VBWBGH:1I>U%>@]/[RA=#6K55T6+:<=)5+%Y<R5?R0T5!^<IW7-BW[IYZ
P$:,E US?MG6/ROS<P%*&-KVYE ''S7U&SGRE'FNQ/(ALT'L-QFLV"3+1U.WR'^+@
P0E^&UV*$05O)=*1IM:T\)9@A:UE+6\#P@2+H_0D//A9; %I<!Q3PH%,U[ 31'5 \
P&=D J4B"1V[V)>--;3$<H4% 0_2+=")MQM&=C;PUO2F7L)=&V&F8/$M>&;FMOME<
P(.CKZ![PZ\>6D33A9P\K3Z7E.+"SUZXH5E 4*\"Q';@/QUO,@@/X-ZW_Y>.*YBK-
PP%52.5,GCZ9M>9&>N,W#2[[32K,"8%N,,H\(=<S(O-YI0BT+: V,E81;32UX2/0G
P0L+^3)<PFA3)3S@PX@Z5"A9 SR<;3P%X+,FW&0X^,JL'?JMJT,MV=J[^%[7]%+?8
P:Z_I2;NNC9)4B;Z2;X1Q;9O7AX;DGY&^I4 EM_B2P\17QZX+>8B'SW&IX$^RQ=-3
P=YVBNO\P%EZ;:3W.$DR:@EHJV=5J[;R7]=F+TF#<.2<@=DLAX5"!5H!;@?]F["O8
PAHVGK[>U;'Q_H VV58[H'J0K[^W.>WB!PG,-L(*<#GL_13>ZVT%<Y4*C 1=8^0/)
PR 2".CGTB>OAB1#"#^# ZJ ESG\C.G]$0"M*8O9P.#A\6*Y;:T_S<SK(&,P&U<TV
P=H\^^P[I(<!^:V3-^FV4QL."L9IU9X7\DP Z1M&.UVCVW$+OZJOD&?29<L+U9)U)
PA]4>%?G0FO@42Z?8<1,^BPMXDG@93OS;GH"4KYZ/N>NPWHQFK%$M_V25-%.]?63B
PJE+EJKU6ITZ[TA=ZXB\ 8L6AR6R=],<?P66$0F&'<,ZK-@Q3%1, YL_8-FG&(7+'
P)C02WL 3!DG[G-CR=/0 ;4^PEI$BT",16R.1X%P9W0N^$)0!VNP@%IB%C"]%P-7)
PL-6ORREPE?)X^/_,D<P2YZ?2L3Q)F&Q<-$W7_(V_V"#W\T,6U(Z3G[K3BZ@.UQ^2
PKLV-V./=(+<-V"=A3U4QK"HT@FK,KRM:)!4Y*]-MT_(9W/TRPE(M'8#^V$Q!T]W\
P\!)K6W:XXL$?@N9OKGC(X)>_6+G7N%KN__6 G&<_98QQGGWA$K$C<'#<NN3^QOYM
P+51S[*1$Z^Y$(VA=DV:L9;=(G4%#ZP<"2'^+-DD')<\2,^_SL%T8__O6N-R-L.<B
PNDQXU*RKNJV3SI?*3IPVA%HW'Q:V923W'[.---^","__=0 M%0V\E2S=,*MF04#U
P@!^-OZ'=O+,;O]!G+[G0)&WC?;=)^ID_B*;4K)-@O@TQ/G/X"O4@=E5F:O #MX\+
P^"C%WYO!8808M:QR62]\%_D\@AY(1)PH1=*,S.]9X(-2T%1AO-/U:<%Q=+C+W..I
PWEYNSF'U14&.HS$&\B\+?X<3\E1L.:,5/"!(49A);[<D@<#F] [("4I-+:)">EE=
P9;.I\&/[%[+S*9+D3WTJ?\  J>K[7QF9S+\L &ECY!W'\;C;EX&@20<,C7Q&@SSW
PY4L^F\A)@;S),X)\]X?/%8;=U=:#8$58.SNHP!#()#YK!X^7+NWKU?L)=?N!VF#3
P#7OR08*U_*$9S?(DX_J\WJ'2&U*SBYH-2F"2LKWUZBT&MM\$"<1B]WSC@"F\]%,8
P6<^?>$(ET!PQ1B*5^)*"!N9\2W=#20MVX@ 5C,=&<+<BEI4!GUC[L6.Y-#"5@C?Y
P?YKDM,.W3?O*M$'V9(I[+ZDN!8IT2F&-%KO.&RA29:I&>&TYQ--GJ:"4TFP'P?X?
P-LWTS3M!^'G.8/!F).M("1N(N-/$5<.-BZ++I5N8U<K:_RERJ=Y!(OW(([VVB=QE
PK]6B?-3F AKY\^[#UX56U">IICC-8".0_C"/F/_%%K[@3:0!+A73/,>I#*HYM/2#
P*^DHG0M.VU%M\04.'HRG !;_O$J2Y%UI$0<P^J[1?6?_+6(M*!KA62QK;$=L^79]
P9ITGD<([:V][:/&.O7PQ%CE8'FAW:F[Y>Z4ZF!?/XO$CLCD!SA' #/[WUQW9LKM+
P5HYIARQ;,QRF8<U,O<!W[KJ,R#:K__<*D561R))/(6H&MO2UN+&.F8[:^XT0=F%0
P!C6_;%:\E3UFG3ND#SI!!X'JX&MGWN[G#I][!OMQW$.,'?EZ'PO'JXH%9+&4Y+4S
P8,L%O7 ?BMS>.&QXLVJN&/*/E:$07E+)SX%F?,Y=+//=YH<!<O>2WUT7#PT=&/*7
P&PAXB=**,(228491$X17(91$>4"3^=[T9J:![72O@#"<P60TL$=MD<K-YM3PX)10
P_@42BF/>Z[_^U9@=TU<VT&;OHKWAUVB;NP+V*?M/H-;ZH&/+YRAP_59)L2NVT/C.
P]#5V_TRR%8]3"7%OZ1F)H\9R8?CC;^90BQE5>-$"NJ^ 40!";R\IIQL.(*CAP!R9
P )6N-\=Q)$,PR)0#V<?9XY!\@ [BS^D:SXIZ,Z<MU1$ASBI%;^&WJ!*0*[N"J'X=
P6 6BM5:J5]QXH]\Y#4/2L]IOVFT"T%I+OF/662*JIVS.=ZDKK]AX^(!,%#Z=(&A-
P-I8YIMQL*F0<C.MPL3+J/)L@_ _I9#AI6)\1I@[)#5%X=,+Z:(C9<RN@\X+M*%<Y
POE;Q8PI41ZMQ3?H 7$O1J%8ZC080)K/]"_F5."(F:TH3*:Q56:C"U<J;348"KYIP
P[;#9][+XD'M#6SM"W>R @6:=#RIP]N;8$A(L2MWE%'228^R:?!++Z\R2(6U$KFR$
P"& +G3;"Z83TP=GWI@'@90-:-6DB&;>&Z)Y<5@V97)W,'X7"5LJ#(F3UE'\.3@NL
PBY8]1BI?\/Z<V=0SDMFMLU;1B:=;;M[ A4A Y1U9;M<RI/IHF^)#XK;N"0Z%,P9W
P;X!"]IGPTWMC[9H<O4PS N9*\8^N.G76;6Q1A,PRQ=\?'#.XM^RE;0 2[P+ZE O!
PT$7:M5+/^  ?/S8 $(V$+T$LN >Q(?.;D?C*[B'G),AZS0/1A!YWKG@#(Q[W8F@F
P;HH>5.)QU9H4Q_XZ[J;DA-Z@L5$S9\_HM.'7=$Y,#$UKK.B3BP9( C?/_0XO6/U.
PN!Q].+=%"U=VU8U W_IIR4[%;FW3*6HRGV!:'!5<C;OQJB??1(?.DF/6CM$5FM@^
PWM[(8HZI\>_\ *#8^)"4GH>PYGGE2J&QH]3"I+9A-\Q/!5JKA@X)Q.-.49$^S@P4
P<CW3&7ASGY*X0T5Z\46G_.3FHL$'FDAX LX/^/?6?DP7<#?*%>A.YM1?_W)EBW*Y
P3H1XJ^2,,=+&SK=^W_J<LS@6XE24X=[OW[,=E>4]JR@C.W! ;Y'X^28T--LM%BR#
PFCZWF)C/!M)0TS#HLZ*D<),<DNWE3^O0B"]+<4)NJK3L, VN"3Q[V:7#5)W99MHG
P!U<SDSCV3@ RMKCZS@'5]@=3@=QY>IC,+7FMAYD8US)<TJ$I(0/<31.(N, P1\&%
P .<C=Y''L^\<<I<PN![T@K/+C7:*/X$U'1M? FH07F?:W 05OLK'PG$!'9$[QD"L
P8/CPCY\#J!N[04<B45?ZI2I#$:AI'SD^Y<H%<ASMJ+RB:2G*+1*L\\.<[0>I&]2?
PV#SM$YI3 "%M+>0KS+$EY9!1H_YHF!_M/5;$80(^3I5T#Q,@W%VGE9?D8C/GU%UW
P7/MD_:WRPT5\T1:1QS=R4FD(Y>K/*C?7W;HVO1)._R8'5OC-N4YG1/K>I:'0AXYP
P^*=$+]I4RYGOP@NG[_#;&\-8POVGGEQ%OFGZY!-.8HK&*DI,AI4][]SP>6[+M134
P&^OER-H=J@&AZ;2U(W],HL-'<G[,L*VDVDVJH%9,%LDYQR@2$3-><'J-8-K?@@:D
PFOZ4'^XH)550 T].,_478+1GUE&YN=6'/98#GES#EA&8T?7NZXDL>RK0;-K>]G'<
PD05I=F"LQR$KX:"D9"=!JOQ&[$X67PD-I#3J[!SV#W1[.^7/(K]LC@!#]W$=]EP1
P6$GJ'3"OJ#Z ,O[P2DYE@4""3D>SB)D0[K1V/^CV&F\YBPE?3EH_(-1IF6Z8O"W!
PDS[2SWB[3NF68%R@ AGU^T\YL45G%#VQTY@(.-""[MPH1Z%;F%Z;%ZJ#T=S7WM%I
PD8$1$FV8.HUB1"CO0N/HJO>NUFL@"&.::0A*&I 9F":E[9GEQG8K;0FT?:L17L;-
P;W_3(FH[4,1SYX%6B!S1S,NQ@"I[HTRZJ9'*]:E#.IOHLV3G*RY/)V]FQ\\1"#V-
PY-W (,D7EK^6FH(](8>J9_SV6%$K=W*Z$M@P,4V+B8048-U,- %V?#1CWZ/D+#]C
P4XLJ.,%%FC_2[RMRG.\>D0H;6X%C="_"IER5;9RH?F22[6XM'X,'(5=KXZCV0][]
P(,?7;WYFW*!$T.EI9+!XZI,ZZJ\T<WN$*VJ'"X[D'?Z,N\=]8X,@O*IDO5$_TFH*
PD3&OYSP^3O/&K,RMEWNQ5(G-D#8DL"ICW98UZ:8J8NNKK^B1925(.V*^"'PYAZBT
PZ0]\M_HW:*&P\V!!C7X ;B(ONMB7OP?8]R+29!1FM6;VV/FL+LO$"KIY0A1[-IK6
PS!A$Z;-0$_];2TOJF-; (Y0$3RJFA&47\QZ($%$#7LA+T\=C &2AKO6+?IRM&=L2
P=D".<?-WKN_99_&R-FOFL6/:'*V/XJN L81R@^\9!& '6J.(?X;6:689HM)9>H5%
P)L;K6LN0NG: L6U^PRB[1_XH?E?^2?ZX]2>#AD7Y:[AA7^RQ-]H6'_8.>B8N#V+,
PO?/XO,P=@( P?.%+_!U10<6Q),).S+H2L^I"+#[>10R.#Z.AZZC2!_5YR@SP&>H,
P;XL6(3].),(,FF8L>:]H**M-J2'T-^PBY1KO7 PF-3/I'Z]N4LK>Q=/4[)_*8#:F
PBM,\LA_6FU[ H1"3)*XR-!]>>D.:7A02F?)$9\DI+B:;P^%H+JR]95N[YTRVQ@WC
P7@L>6,-&="]. *KZ6<8:! 2X/=1>G9YUJ0Z\J,:)ZWFW%-$(>?./M$$- D8ADU9)
PT3#40M">NA&+68UW==!OPR96+C%N<R)A1J9Y>.?Z!W$)?_VX!^*QB[L??A08%7"Y
P%!PHL9+G<CA),Z(/?"X7%.S<%@)9(U?651LY*1(=%\CKRW@G))=<C]6/\;X,:O_9
P]-J]J'@7;VV$(O*[+'( >"1SCG]%Z$Q-D3 NHL8&%:UKY!7W"!MH4Z*N?QN&PE(^
P/S:#%:+N*X?BDJ5%7N3][K!W7)O@?N8D_E+61-S&VSK:1H;C'D#6N]4XD7<^_JQ5
P-?6ULWI7@]=MJ7-^VLDN!IA#"D![95Y5?ANHL-M309CM @B+'7.O8-.8;4LLL]$.
PLUS&87\_>I=+S-AQ&"TF&B</S8$&]88^<'O6&"'8#(%*)L39#2NUGO[A(Y[]F?L)
P&?@:&0Z^X_I?V2L8(2O@<\QR27^[3"'MHPKC!.S]0NLN+/6^M+@J6B("KUO&DEJ=
P2Y",+@BP>LL65%%2&T"@Y_KK'QV_WQA]/\W2 [_G07+KX09F4:M$*I@W)TO\LTQ0
PJOX647EV&'3(!T.K($[\.D4UG=3]E73+C*VF+HM"&^?AH-[4S(T@6HVL#7^;'P3Y
P0,_8%.6/:N9CC.JA2YBMY3N9\\(O6$ON\L+9-N_)@5F?4P\S7I6VBBVE2\+4,):6
P>0)$.'^@?@4]2?0H\$X-"+Q.DISDY:MHEPX6_X>ZS"T>\)?IGDX+H1%_6G,[Y:L9
P<BTI!S-\5"S*N?;'IK)7WE^A@ $?_1"+2[,Y?N2@>$X!FOLBP,-AUB;D^NL=K3F^
PPFD<W5,O2<EC&Q"N6XE89&=OTK/*!(M5.*!L]Q^;[S"]ZE6O%J,$W[%988GHX@2W
P<'+;/PV8$!55H(X]V!1IK1DX#)N(B^3?-;< 2C&)&0VC!I6'[R C!G.!__V FONA
PGTG$1\GHKW(;X=0(GKTIF2F42$4PP#X5NJ]@:JV_F>N1XQ?3/8_C_+/.3G;Y\( C
P"H=CEDN<>@H44T5;+WRJN!85LG_\2J6)UQ$18+Y=\05]@_!%!TQHJZ$,AYDZ6DJ&
PN694 =0]#/-I 8@)P<[3A-Q8F_?:SE90Z'K#Z'"&%,^1*6\R!V@VV2O$-71I3XAH
PF"U65K]FS,[<,DYP/84S+H!=U\0B"KDKA^-%5%L+J2VF)<SJ208S,>2/D$[)O9Q>
PB C)_Y T=)'CI\+HQL)QQ7^K9AY\%M-SQ45U0G?2DJ;7!1G-6Q;7" /O"%:NX$0Z
P*!%W]6G*^%-Y&QD*'Y]H5@'C3K)WK ,E;Q: E/^IVT=7CD^.6NS]Q7'V,'O?H%9 
PK&#7@B.L6#9@\S^3^B-&_VW=)G$Q@TW]O+KARTW$YR25W]5R\I8%#\@A&K:B1_8/
PL6_[5U^M9+%WOICI:'&E+M&RE_+;"(V=*2.36D+B;^/!+5F':6B^= PA SL#:6GZ
PAU:(MN83:L[Y*^A-:(\"H]8HA82U(I!'H78X)DXSLTO_?W.X]*CD$5-I#H>WW6_@
PM:;!*^Q'\W/12@_?J*EDO7!:E11D@T9>V%RI#J_M8!.GR+7P\AM14JQA-I!$' D6
PM'>BOU9G!>E1G].S&]4/'N@-5:P,5:^"8<!B!!77"*+RET!&3E\*P:-")_0$B[ S
P83\-O-I-DFUU:J,E1]TX0W8;J%%;-%D_YDN._S.7<2XAX/C%[SZ-Z=/%T!*A26[*
PJU-F*XP;T\ 0;;-X5:45@M- >7*/DE*J$6M;6I2"7 _<,#LB?F8SL7"<U=:7H:C(
P@!G6.;L(.(U]S7$M.L!:B+.%6524W[KZ><-!G1PK8VU^J_A!N5T>^=_EX(U9"&?.
P9OK[?3L2>LLBEC;VU&(+SKNW%0^-*QLX*9J$SS!]OEU-'J0:&B6/?>F9ZD95H^^1
PY$5JO27X^8C DT>]AN/:M3B&U39IGM',U.561"*_EFCJ[A*RDU,YQHO(W0VP,UXZ
PWR+#ZT$6@WKD*2N5EL02-(N4KP39 9(V931\M.Q5PH@4;$+"3JY7B.D(DVOVL9Z>
P; 0.CO]D+)"TS_QG5K ]QX_PU'H@)TBC/PV]; ?K!=/"&3L8.NL^8O3-;R[79U/ 
P'R\.=@@6S85.FN8">I/KIHFSV7%%:,X6H$,172YJF;DC5BXL&=>I!6;I1#VY)XXJ
PVK[.2@A/2X^OQZ!P=]->#T/TKN#+C.[8B[RS7UA$H_ TQ??J>YF7-B1+AY#X"T=E
PRR'M"T?T^[3QC;O2E@Z&,U+[P;U=P67=!6Y4:M=U1YS^HH]IO[:\#39+!\%(KJ0]
PRFX-=U?UTJ9N=VZ%D[RN]3Y=_&S4WG.I>$,: _7[6"3*UU;> #.6R]QET_CK('UA
PC:\^,K@OL;* )6>%P'TF65\8<S/TU(9_G!7E1(CT@-#L8WY\*BCTRK@$@H!@@ID?
PD?+)I4K:R)H(@_RXTW7;GN67_5;/4V."'YUCV=+^E8TW_TQ"$7C)@TSM-F&1VO8;
P1\R]Z5]=\RQ28F0*AD!04(J=V,6D[$8BHPAFGF\,.YFY-%CD&E!.L:ZFDZY?[.+A
P+U[HL^H=>PWEE$A@DX^-L0MDCY:%[:.E)S4K(.0$AQ>^#4=8RZ<'=0JMY7\^/'A*
P0%(D:_;T0YWA$U[?#Y;&L)DIOV1S_A-]^^UXU'YD3\<4,>V8&K;)G6P2&< \9B9,
PM+C"')%_NX_+XX-M+<!F10QTL+-?0/9'"I8XN3MT%.GG/C XI6J1KT'* ]C#+;R_
P8[9) V-5+I'8Y)A.2+(*?S?I^,S?5>:YVLM2YGX?<S/@=/9(O PPH_.AG=-+"I"#
P50HXHMW-U5Q3!G)"=W,*KA>U("51/ Z=B!?';<FOZI[1D*XZ9/'*:F0I#VTY!.4C
P"MJF[+#M'A+\;H?XJZN,\157!VCS('@B7DQB=,HK3!:#8X\MG\9VT9_SOM4LHC8\
P%XTQ[SD!*>D"W[IBX5=UUU6!I;V8?YZV&7XI9YGE1OYY!=*[+QLO:DIE)@H$K#7&
P4/VL@4;4:1T=,'QG^ EY+&GEB0-CZ%?(98FW-_=6-["T?DG8-_[!<DAXR4?(1+=@
P_<):8UWB@UMK'\A=!%W!!WG$.31^Y@;U=B>?Z@E*6D?7@3[(48]MW7Z(:*0+N_!:
PXPURER5&Y1S,@R,D <P^'R!\*_OK/A@YQKT\1U4$0[<I0R;N)H%AV^;?GCZ"KHT^
P<;TG)LKQ9#OU02,V>27G@K4#0IWF4H-2QMJ"TT# Y,O1@,@::3;U?P+M)X[ .(%U
PM-N[Z"4&2<<U_$>+0IB@Z750E/UUBTS:YYR'P"X+13YTL6CPZ -Y>@";'1UB/[4K
P#<#]A23MWR@T\]-K,<V\\<G>UEU(UF'"&@ " ,S66A@0Z!#M#T097,?'%/VX"WUN
PC3:+<K<L J@Y-]6K'AXM<\RR61B:V0[;!Y^G\5V4FL5/OOQ.?8VMO4C8.]<F:P__
P"EC]%PRV#>M+LV\*9FY(7M*;#;&YR+,8!2 8>UE+H+4!2C^(R8 TLLH$U0ZG:]<P
P4Q-=S7[:,1*JGTNM&MO[6\=!]W(TGZXDA9XV]O3E(QVFE(9FW6N=@6O?[A7]A(GB
P3TOK2LIRQW[XO^W6JBM:M*L:F[G<\!TW<N (#)9=$7^Q /\AO<6ZKVLE;T8$C#.[
PMU/3Q)66=9!>C]%"R9E5'^C0+?MP7$5#A?[C,EF':@B,B*A?>+,9&&H"L6WKSY1N
P4;IAM5NC;%EK<=9*49"! QMD'Y09D.>%1LL@#L(7L8M K!5,(!P$</F8H38YUY*9
P LP5YL%W59Y*XER6VS% /L4,5=-PD(K=?#V>6MZ6($H@8-B)W&SE*4%[%LWJ%-L3
PN8%9PK=SAZ3JL%$U*AGR>,5@Q-I5QF!3AY$#%K6??/^"02?N=MMA!XH!!S>GK?SW
P^^AU!+N;N1D_8>&8>+U:R"/(#6,\39-<*/(GIN\",TC1!W+/B_*"3,#CU+(C:>Y*
P;=)+Y3HW E6%BNLUNI%%(75K95%HO5T0;S%=8Y\,$?"R-JL%V_<;:@1U+>$]PT]I
POUH==GX*@H[.O+"L)(9KW<D3,]ZE/GG(1%S_E-NJCI?XM&/1 ];H<^(%5Q-,(W_N
P(F1A_1SPR%%_>));&Z!2D0T#KJ4'K/E7&?-L%!90FG7K86AEVO&UMT#63]>ZM=\G
P@1XL?L>8D<<GH)()ZDSX/YH 96%W7&@): -R9-ON+'E8-#G>RKU;A)1CD*))JE_D
P6F*QY&?"KMM[GU;EP#0V3VI-8 _K!EG#;QI$@G83%0JZB6)Y]@6UE.W#_EG0YX.H
PF;_^R+Q16/J11)QTCFJ!KB>O+X<8)0LPZJF6 8_1%U>!1AK0KM:&@7[!]VHM/YKT
P=70A^*?.RDNA8K?9HCE"3130&,??KA8<$V2U]_U(@!?M0!FQ.&#&[3RUL^+T%GPF
P===2C@#94] H;+U)+>RWN?*@B^"F?C7VF&5YRT-'V!2JQ.#E\\L#YKX97HE$$X4:
PZS-108-Z.;PT"4(+OUH8K33J\)ERM2PDL$-8/56!XN:F._AN2 @$!"F[?I&$$5>G
PF3."M5JQ3'!/&M[R6@:N/>9R  !;-$+WFE+*,)EAP/C-<+C%U5P]*%HH56%N:;"3
P2B4P%=(:/K(S6/$E?DR1\17#)JO(J;@TK9]N,%_H O!^CSWUOTT5THK"B;IC=RD(
P?<='[KA_IXR2E^AVSCEH[K&V]RN"^=EK ;;TJ#;.]U'H=!C^#!: )AD/$TCR$,'3
PK!PQD2K%<4:_$2^U'B#6'B:;A/C)7C31972'C^6PZATN!G6:588/ K[A4O_ND)_<
PL K"U!Y&7+KJ._!0 ./)(Q()6%$96=#P2(_RU)W=A;TQ#FR!"3469,EX;OM6JF"J
P9+)D=5YWI?RDBL[@[,'QW/D2SRLT%0'>_M+[_=Y)T=8A^GPEF+WXB*-\+(1:?=.-
P7P/*^)GS#\+)W''X5]F]B7IL;#R"8D(7J!D1R-"*!4_D _+ ?V+BF!SF!^BL(PZW
P\1EH2YH!'X >)9M-0L><HS#[V>=T"/@+[^Y>6&3NMAX/+LVO\2^#J4PY'>UXHO59
P+5Z#LKV0\MNMRZ0AUIA[)J]4K< 3Y@[I?7PZM6=CFT75!+L;"R+[$17IO)^D4UJ\
P2J?X; ^FJA$DY" G'KX43>FL8_E]UB/)<\Z[6??7^+ M/0T\=A?8Q[V:H5_J0W\H
P[PT'W^*^T"A>'=5WP7J. ,S4>U8#RHB:-W4H( :1"T??N^6@:3_\LYX7+'K_3J/6
P%[/(-Q!NXPY^&0F.(:3A8Q:\6-Q,VI%"ZP#O2B-FL:;+W=S@%G&&L&QK%OOB45Z=
P8?(/*) AW>%K'\G,Q;Z]_7X)/6OET\@;MQO;BPF."["0B=<6CY,TNBQXIV M9[%.
PF#EV=U@C:^)1B.5:+WN(& GR@/NA,)\2;%0TL)9:<VSW*!LMUOX;,Q[Q0OZ(-;J0
P0<2+AN714ER;E6:HYS_G<OB0Y;-X0XOWHZM/HK+BX81_\ )S9I6N:P"*+O/&2$DS
PS[&0)R:<$^NDR9PM&9=Z(W_IF$M29(01/[!<O"633PPNO1!(ZA(*:<AB&PMC:_I1
PHM'EZ79_.X2N"9,4WK-PWLL.>V<W"+;]@. @QM+)>#[Y3CV=IB4S5+C@^*Y =9V"
P=S+7)82=B.-#$*+HQUA*',T#_Q>#V6VTESZ6RPO_\G_(O'10<RNN5WM-+JV6/!S=
P\CGR*7@YC_\S80.C%"T12"U6%$-T(N'A60N@/=@:=$".UM$;K)E->(<<F.^.S]9'
P"TH!G&D=61OZ9V\7Y%!O5>__,6V1?4,,%[ZHER9/-74LN3%#&HTK6:=/;GW*1D)3
PM3"6S.8&/:7'/6.^W%1 W-T>X0L+;=LBAA$;14CJ.TMUVZ@;DA?-7[&ON,RV/0;8
PE-OUB[=>-ZV]*5V*J8\==2=GICS>##=+$TG:2=V8&IQ6-2J=?<B0Z=F:JF$QOT^S
P+06:!DWA9R&4&O\.=D*%]%TDRN&KQA/5C#EVOCS#%7YRV3,,Y3J5"-&;VZU[NV!3
P3F8Z1+3634.H4!&(*^0T(%+O+#WAJ-0FH4P?^CHZ4"3.,3_;Y+R?+>=']BL:'W"=
P4Y#"8I7S*0_)X3AJQL4&[+BR9"6)BY839[]7-FL\H]__Z8'5_CY2% ]'.AEE8L@K
P1(R^KODT$R_LD#<3M^W\+$40Q@$C[LF;0>"HB7,N\U_,G$ XBXM<-S QAKVVEHD#
P^SDD$EC>\Z?VV,J_9505&[A0B/:[$L[#C]4YO8&#J[QYB0#!MPBV/H<_W 3/  )(
P8;N9=O_*=9?*LEZ#\LDBG5A!7]+\=)KMG8XPHJ'-ZS+]F259P<^_Q?QN-']>_8R<
P(&HR;E&NI?Y>X1E2:5XFC^ :5_?;,4@#26T"Y7@4GR' .75EFSZ(L\TA(5(@4;?7
PC%@W%QS<2VV8D2$=3-L.$"-@J6$4M.27G#%?+AOV-6S2(Y:NRS'=^;A9(B_SV/+&
PKAAA4RAY8H@!W_(1%,IXZ.K.CV9@F ST<;J=7QJE:3TC-Y?)P+X-D,9&.+Y=MS8(
P&4.567USP'1)NOQ0MME_PVTFEA25P'=X@)K!]#)0W NQ<?U&,V<+L/RWD#FWW]M$
PQD[ML[L23Q+"ZWV70&5%)4>;I4P O"S6W>92LMI;>E8[#.IB601]*:EH!S5 _P!$
PJJ7C.MHE!(&"/UPD^^).:K,3AV#,QX#4U,^2^>EV@8\P#V)'-\,!&]A"<(]'@3;,
P@GYF\ 4[1K"'ITGTU.&D_^ZR8&M(F,8YA$H<2!RH3*Y8!9%,,O_%<I8@&.H!;E2Z
P?@=R.8L^<58\PED9#%0#X:7&0Y'NYN'"'LTT!56S0;J2AR/ $Z7$B0O1:7GQ3B*.
PYRT"F2FUYFC6V3% ZT:[KA9)^J"D^NU?5K\=+=?BG.00=\LHT.N@L..C6[(ND&\>
P25@0UMC2^!_J+V#=1L9N]:5NA5<FG+S9TU63TTZ])+!@*YR4F;#8L>R#/.)]HD#:
P=]/%3XF3\14K<%KK$:(<:O01&MB "=BN\;/RJK3.ID^\-R_]5@W7Z=3 >9#VGBZ]
P1Z*\F.3%NSV]8\6&Y4,._RX8AEX=L7EQ(Z(K1U.XSDC8FE_Y.:/,Z+!PUQAP? ^5
P@NH0O-I-_G(&8,)+B,?LE,M\0!5(UG'9B50Q%G2/]UR&:>YSI[-C4M>6]::B*9@8
PUCW9/X@0[B",K\_Z7=I4D7[DN=Z.EHW5%)&'RG5!!;K*WF,8EOPVW^X;;?\SW\RC
P@"]P:,"6:6?:8)R[B:J[Y:V/]RAS7BR@**6T5PSE3#28*==WRM*M3*5?VO*SJ57\
P\XP^LK-B"S982OS/!F3T#42WIHQ$Y^YF#C/'CX2Z@NI=N?&$\/;&>]HSS+@5^;7 
PWU@XP';5,;S?4Q/?_O2Q6W)?':8CJET^#2.-'O^3 .Z^9WR<?YZK[FP?BG#,J0\I
PA H-RY0 K,Z%*E&F>;/$QYH)Y4?_GIVVSG,6JANDDI#;ZH>YP=B(,0_O-T+*@XD&
PN>]#(WRDB9X&'V-K\OEKJC.;RI?>VY'_K[YNXPV)))GP3_ZTZA&]W9>K(K$CQXSQ
P4R;>>\GT>\XM#M'+*P@^H7B!^2EW$IPXJ?&0J9=9Q,B=,^:?229\3BF;]>7"QJK*
P;OHV!T&X4<%,X42G<<^:+?2M-)5N>]WN_-Y&V)IFAYKJU]%=8$V09A=:.,>H41J3
PH%20@QZ82$M&H75?HJIC184X/UO9['-D#,F:>([.]3$(O>(9<'YL8TQP[WZZXMM3
P1F<#/S,N[5$P_V$NVHAE+.E';V^]19">$\5_!#KMC)/*ED##2L,9'9,0DDD,'&CS
P%]4L6";#^)SE=58ZDNRU1(QC3O-O\8T+DDQ"_G90N%<#9&FR&S0:GDVCW;P3F*0Z
P-J-FZ+#2]_@$G@[]F$S1:].FV'B=YPWCD8:< Y64A]Y-+LG&!I^%>FJ1>9+^/9R"
P_@YM^-P5V0EF&+I@=0UI:6P'ZW7YQR=OR(YV7@.$ %J\,E 0@BJQ%8OV'2_M[0UV
P,'R@N)A[%^F@W:8H$<I*A8?RV\H\+_8H=>HS;N7L&X:(9"A_-Q]!I07;%P(VAW+G
P8M#OY5FF*0V =#7E(?UN*9$P3;OI+\5:$%6=@3BT=+&7A$NC<YX@LTW<O+D:7E@/
P[V-71DV+^\9[['?/VY@>DDI+,?''D>"\/SA$QWVO*L@I6FY04!M>"95SQG#CTM1A
PS8J#] \3I:("^V-@ RJ+&2=,SO(W+3'SUI%5TBGVDIXZ&B';>FK*#&M%[<1,.NC6
P3[W Q/U7JR)<+I)=CJA(3QRJMV<[EG#QO:KK1V, 5)+[V;%&\IHM,QB/-"L5GN9O
PH$\7^0A=Q!"LH]?C1N<DUL"#9%@B+#JC(^)B F)>]%+;%$-78RKNX,EY5_\S!\BW
PO&7KSJ:48]-PN7=PW[=D \K$H1VIZN,F]URB;">PI"$-A?7$;@ZX/[-6)OX%NOY;
PJA/J*-=8.&@>/)4H0'Y.&+M['2[XA>>CXBHO1?@7A$MD^EPC=N#KQ[QDGJF>QLKY
P(),Y"9GPG2E#A3K>&_O_+NK7?,@)9N8P'FZX[QBMN!Z4H<$?.*)O6D5*C(T68WQ\
P$TF]AOV[V\/6QT1EXP16.:U%PRJ2;1PJXW*H!,Q;^/Y_+H?(C^C.Q^%E^,D2_3>I
P,(PKU9968=#0HE"<^G;?&:[)0'$ +!#/+B.196FK\:6!"N*1'[I,QZ+NTF3R),P2
PJW>_\I,=-J#ESE/M[]Y_=7^6S'[6$7SXU;I.J7P'W]\G.&)2QCXCLI[5-Y<^6YSR
PQ>!"K)@O^CH,3R*B+M62,B//U_;WP">D#(#8X8YE[>6F[))"]25K![F=U_&Q=D9L
PL@!%[T#QS<CS6KPQL68T\[TP8*^IEOFCL2%=;[E\5N]Y8*/5TV)<]U!P*\HC%;%M
PV#1*4S%3E13^(DE]+S2=!6+69DOG[B"KJF5OV'DKA-]3XXL";V.VF'B14$E?E!SR
PG U_.PWU7"1^0X)ZFBYEE;KTI)2,XI3F5P.$2-^D2VH8$7__V^]IM)\)+U/LSINT
P\3<1_K#?)(.<5:UN\/UT4EOK@-4<XUS8%F[!:V>7M9^GDR,)&!^MV!AG\9^Q*EE(
P*2XOS\BBYQ6Z%],-G/*! AX?3>&CO4Z3\P5OT]QNG3(IK?EAS($ 3TV A3AA>&;K
P4F7"W7-C$JP5]Y^@Q@P:8/>_/90JCK^VQSSL-SUW'3M.2VYIL".,OY@]N=@M-_I'
P)IN#+NQ1=O=QSU5_OD7W]0 MY:R B(K,>J87Y6T;A@C=D\]G+B^XZM1MJ B0)F%-
PA ]=J#=\#E<7N.9R(:0YEK2I@N\3[8]:HE'^<T1^UM%J&>IDE*N%Z+[S[--L)B)I
PR4QA0\#HT7J-G.$)6/UGG<=J$7?FQR<@CL:#TK$XGN%,[ 97.S-6L'"HU87LJM_G
PBM-?E4&4P?&8P!.&SP7SF_GYUJFW[BW.X4:= 3G8*:)W:P._1Y$Y1@.I1)TU8%"W
P3K\[G+''$5P5K2_GW6B")/A8:-6TPS&[@*8S_2S="/:\0?=99A)N[[HB,1LD693C
P&S\>]947Z[!?R%Z<-)%2.RBJI,A-A92/!Q5*TH:_EZWM3%P.D)9#X,AJ3O+)W"T3
P&S7Z6R7,]"&'1[%ODEQI.BX=!;J7!*V<^WDBEW9?D9"200*U_@W+;&BGLL0'_$Y%
P3N5+Y$"P>91+,OM>"'_,%_ 75RPZV^XA^NNM/$4?H(1P%I/4WT)\9YEJ;5(T/MD+
P0*H:RM0::N.;+4]^T7R[Y?VUBSF)1734 %4,<-_OY*RE/:V:3=F(7L.($8R.A"25
PEXJG"(GHD6>IB V>1?PR?R@1Q2]I.[-?^1.0R0X\VGBP!\*ZFICECGN@EWJ-;<M3
P>& -+)/R8<7B%ROD2IW1R$?_FA%&,9GP;?"IU[!:,8=<.*%RD6G6@0JPX!+21_6!
P$["(O=8' M>B"APN\&@KXRS%8OK('V[4-IT:0&':P*C5H%Q%>ZC"H\1V9^=/5-.-
P34AU75096;G&^M2>U;0@M!Z%LQ;OAG3-3P"1BGJNJ':4JLXP+A$1 ZN6<D*2[ OX
P=C\E/.U*Q $" "$!J,B3HI_<9/*@^H_/;+GFT, T%!KPIH*0*F  ,F_-.P<5(LZ)
P3D:8C\W?9 8G6+5[6BB7IM@[*D*:(KK,X#!; ;KW+S1GN9,-)EH([_V 5^;]A'^]
P'&?1<!\;!R0 -[A9S]?G<V.P4OO=U8O&_N+$.QWGXZ;#4*HP8[UY.B\W% 3@ATML
PP]JTZ8$ZFB IS?=!8;&_SW=%GT%D4TRP^! B8XLR&.I]:\)T_#_&<?Z7"59YR7H#
P!/,TB3LE?)Y6GQ-M _=)%DK,[N7&LQM#4'$PE36^#$F@-!\[]U-52(0 N-&*VJU%
P"8CT?4#4_%#P&(6GP015-W:.,AV*98>EKT*83/0!3GU6E9=F'". ;!==H<[,:;.&
P@WO(+/LXNQT 8=JJ7DYYN<S#0OBK#JZL1%N3L1>A9M!7Y<7.9\4(X$4!V]<2+7%3
P1-_!\8QCRRIM<H8<HA5:Z[$(X(//B ! R5&XCANM8]_XY;V<ODL"NXM4>2.9XY?-
P*#4\8#(O@6Z+A9!=1U'\8K*80Z@<ZF=L'S?)4V.>$J#)XR+*6+<YFN]9"Q0.D8QS
P3.'NS!A"H(S4.8T_LO6)RRC^%;L(%<TXN-H#&O$;8#GPMS#[<J35XC0(>H,C%8_N
P.([2VMO)%XNX*1\05<G[ 71+HD;4R?B_&G[0!@);;CJ>,)>'((&_*FCJ\G"1=;C7
PL*!V';HN9QSG#MHM\HTX'9HZ:75"TDU'+<,V\:UF4G;TJGYR@J%V--/])FQ6)T@;
P+?'3U =^S.),SQ2"FVI22"6WT.4BW ?$GO!;ECWVY8$(//R@':B7:J4(KW<^(KV/
PE8(;\EZT+:40.-#4&@)\%7AX^UP-)7'\ G)7&-AVNV8R_(&+SV3YCJ;?PG%BA !6
P8T54@*;5,#_0V517&OPD+C(*(V@/"5^)ZHU,2^@O\'S#=9ZRSB'%XI!-;+CF:&MP
PK@=QPA#^V4Y/.!JIF=KL L*]N3'O@3R>;)==&E\(8Y_NL3D;3]X:V\L6%XL2K+ +
PKX5!:TY8&KY@0,;.H;MHF8.3&?HO")Q+S'8$@=RE::.7K]*+DXOC3-!^DFSIL0AW
PWI8\,8\T3),*J_?U"W>A?IVSH@1 34@[BEX1^[=8ZG1P=_2G[<#FT;0FU% :I;K 
PFHYGZB$_::H?A:$$V&P\+._<TFT98LU(^JX%?SJ[D,?1+J4IFCGYA28\_?$Q[%/P
P Y+OFJZ<F&J0H56GN6]\3D^YH5S60T[(+G-]XPR<W U;&/NP[) 0]-G3WGV4,L-C
POX'_NI:3.K[2_0^'H5XER5VQ?>BUE:"2%3]SRA'UJBZDIY!CL;09=21JFUY7JX"2
P!;*7-(%9D_6H+.9<LF>K=_BTF^*8&;AT_7RL,R^M[CG3#5K@*))&$#1(:YL.@I@$
P3^T\/OC;,I8F\*4.\>0-<OY_4?H-T=C.0]7*!3AD>KK0&H5'N-_/'MU(IX[4^,; 
P5Z;!A/ 2I<3EVC1>+/-T0LD)DC5<R981XCAZ V(H >6S53DP1G N TE'-D@;:A&T
PNL#A$0(3JT!T9>')01*8P>%7S&IV<YG'VRG"   >>F92OW]9'TZ:'S1.I@[[3@>=
P!&821J(/35!9KMKZ$\B*_J9TW9SY.5%[9?@QP*@X!V4*OKY7[0]ZGI2DTAHY,E5X
P/40AN1N 36+YT,2>-6#I+K_1$2Z<I+_QW5\?2M+=[I6CLR@AO*C.0ZG)\I'PR706
P>5R,%/H!='%B6]70S&WC'.BG=U9YE"$;/F!O0;D,%69^0;0*)X8N]*(/MZ2#*WQM
P\*<D-NM7V@3%.$#!G+[D(IZ2=Y2A)UOM@F*#3R<J95/,Y'O4FVL[+(4.-K.Y9+6X
PU50CQHK_WHR^8_!K0G]W/U\?)T7A$]-2>D)Z*)L \ A#(M)[G"6S*\,UQZ(@8(CE
P48;-'"13'=6]JU\XJ&)Y9@>(<>X B >T4G\XH#<=&"^-P [4B<+TK^%IXA%@95S(
P$LW!I7#5Y54/VZ4\M%!(:P>W'#'HIVY5 9Z0]WUNM0VH]8>_I ^#9^P+^>0ZG\XZ
P7DZ]XF<DEL6>38ZP#/S$V,G.*9YR.?,SY[GY<IT_*<2T8@]K6]-XT8.S_QZ\$\UA
P1*;FR!M6R ]"R*;P&-R"X_)RZ*3?Z3KSBR!^J04-E?K@I&T"]E23L@OSRTL\CB$@
P-8R4ID^82GV7"B:Y'L#W7A)P"#;+$<9D![R5X./Z\6N&2%-]O-AM(X<H06W@!MQR
P.Q2A;Y&)82P^FM?LT,0"AD$8 D[B(E*Y#%8KOH$>NLFN0S^_!4 4 8]\]+@C;/!4
P[=)43*N65NWC;:A3TE%=9X(E/A%<H+<VJ=*DYE@]V0@$_!5RZAHYB/Y$?<Y/S[(G
P_V9M',E\<C",KGXFZ![ 565B==C-";Y(GLP>M)Z+Q?XSK'L^JVM8RQGK]@VX6FDT
PD=1F(^,9^:OW,]NL!O5JWV2E6A>.JU&^ ?N\P<LG FE=*8D8CWK:RO<C50Q^/B=*
P7J-<S3K/'DW?;9Y@GER9$5%%ZQHQ!R=[-YGX1?9M$^;0<$]M')LR C6[B *)&);1
P /I BKQ5N(O+XWG^:4A+6AC"TX W*/4I '=J+1TFTD6EPJ,ZV$D%?LW ;-DUBQ<2
PCY>O346=XG)&)\YFG3)SMZ3*8Z9[2K4#4DOFP,/M]OXJ@DN?A\WV9,RG'%E-NE)_
PMJ!JS=IS&I^AT'Y??-JY_X=,6\R\U?&]<W9"]B=ND8$95,/6+90/*C5TB(GBF1[K
PK6N[,5= 9LO*W"ZU+>7B76FB5?M- J-^,U<)"=/#P<]]]>L9ER&@YN"!QTZY/>H-
P8S]L\6E(7B!-E:.U4H:!WV.G[V=R<B!=K8;80@%>U:HJ<_JA%ROJMCEVIGD$ 3P=
P9[*S;-4]\N^:MQ;I/!:R5%QIDJN$ AEG(;-?O!ECI>7*4.[WQEEOA)L=RNBO4UJ@
PJFFQC*:?I0*L;6[I!:<I!F0UIBH=HD"__X5:(*'7Y=UZ33Q'X^V$D5_VKDY$G-='
PFG_>-1=+G<UNXLAS:O2G0X#5;>LW): \+4E04G UBZ$[[599?Y!O \V'C'9E)*),
PK$X G"S%S-S#0,DBC)[/)DX.&C3;2)8T&=Y1.UT=/O8)<"P\F<"6-^I4D+EQEAND
P\@N.P0!A<Z2C:)RY3FA_HEMI4]]73P4>*(_JIFIZV Y)Q9!FY?7:7&52P>6IB= 8
P8)E==Q RL-Z.SP!P+2=LN B^<O[SR]75V%UX(P9)PC'F[)%.Y6E:FL,8UQPV:'>_
PQ1CMQC0P6V>6$)ZVSML"CMFR1EZ-Y?P9WJG&4,V@F_N^77!8@K57_VYT;E_/TM?0
P(PS]+1BT5'&-LF-A8PQ</U>E.5JSGGA\1*ECA>1<U^HL#:A8%D"]:D7S')(YZ[KH
PH$&%=\IY[B:$]J*DTQOF1E -WSN:P='JK&PZLFX^/!?DW6C/BG3&(ESMN:"+/BVI
P-X%\G:Y_RD0*KZRI\?^,;.&%6WX?4A\;(;^5[!I7_A&\5E-:M @\F,)!!XOY0>PW
PF?,.L [W%%^]I.IQ:'T^.(W8*)IM%*7 T?J6!RY[!:)(X"1VCT_Q6*/AW")8R"&O
PR3CY4UPI971->I/_#@D&#^8<O*UJ]/JLW!V^=H\+H_2%UW3 PU4_+:4<7C"%_\X&
P.6Y6P/<*RE-_-VI./IVUR/%"+YR'D .O'K05*B)DTC1@.;:)+[AI'7]N&88J?I%S
P%*.>\,FB/OV(^,U]'+QD!<[.?D0,51VE,_T2QY]&^JAT.TB5IZY"+6W#&JNAVHLQ
PL+=.G\BSA'TQWZ<*SC,XXS TG_P3R@97TD:WD) "-#R6\"RK*QYBK@KRO(RXK .L
PV98WJ5G[Q"-R36M"YXT>F*[2O10$E(9'IR')A*L)S ]F%>8A5(@B#VU+3Z8M1I))
PZC\Q_QM >WGCZ$H>!(^=]LOZA@7=Y;S[76U WFK?HCD,%#+*.M;(Z\Q>"H'#I2TI
PG&DS%N2!J(<6+I--(><@L0O&QM,8*U.S!+.C5D._YE4&_K@.=/0.Y=A8*W"8^<7!
PMR S.QZ,FJ-9K@CUH8A]^^-,IV4)NE)*BJ@6"". 4H)@ST"R?P$(!\QTK8R<V?JH
P-;I(=%J<%:XCW[D;(-(WC--/3.?,>J*$8A@7O2!$6]'^6*E^!;;YO,3TYB/TQ]F%
P8$=#<R0W@@*TV&XK)377J/ERP>N##I'G_5_XPC,$_F1<H2&6H<2@\)ZUFZXAI#F:
P+7XWE,%[4?S2!K(;,?PFC<R,\27VZ@,< !66T'5&<;)>,/#OHJ;%."T86?.#Q?+9
P8_K1!Q-UU'7\6B"/S*8\>UB.G>(>GY0A$G]=FN(M,;9^))7NRP^,594)*6;M<STY
P"$WT*S6962&,[=:++@'&>6;@J"Z<(\"&*K]&'\UW41OZW+&Q:DBNH2RH,G]3(>[M
P-$^F0(%HX) H;=TXTYAA6 %_+3[8=.K@R$$B@!H@*Y8BJ/GG3B3_GY[JU@F7V0]\
P@)* 9,Q'G3B?%.]?R;U:*_:H;C/8A.SI)<V>KFU?^[K4'_2P_5*CO0$G-6E901,H
PSSWK+5%W(G4'>IDWL/-=YLFEBXYPLGT18(K@Q5RR1;U>GDY)-K2/;\V.@SN9L>QL
P8(X*]!-Z:"3V*I6\Q;1[.JUY<G1L!JHT9:.:=-2J.NBZFKC=(BM".WSU7D[OUV@+
P1!*71!8F*N-#="\>H<=8)RF]KCLUC*%%_NZ9CLQC'6MB]:<@P";?^=F]J^$\&*4E
P?5DAI7T"R83PWZ4P')B;>-9=T;\U?%G$PT-3),0.057ZYOF,*)3( O>,^RGI$HW&
P8 7NU&E3"6I$L=/*GUT5]:%^[#,\LRNLFZ3$KW3]!V>[K1=&1#08!HF662<[5.78
PQ)#B>UT-6-_XD18\,PAK:>NM>47/$(0&VBS+4)L8$?/TI !%>"%<>.:7BB*@#P2&
P1[V8I@A]\Z9MD<^Z[!ZLK0S9D^B:NBZC,!+@1T,Y=!AO6 CB)EIY#Y$H$.WI$4SM
P:"^EE 652&[<)JE9>T\C,N=6/YVY0@6%0LQJ\$*14@//%CVU!)^OT!X^8(0)2T8'
P8)?2FS1!?,3"M> HC'QRP/A-[GHZA\?5!#/>\UM02^\3VU('E51<?0XY@;QF4VS6
P1@[XV/%PC7KJH/30MR/,X2%^+D.MV$E27SM9DP(]^&"M;#FW7@,BIURW7'Y ?)-T
PNV@+WXNA9=2W*HBF'^AE;GO$*&@=&MGOG#<8T!(L8!:FCG,H#F8Z0]AS!:64/,".
PI @CL%*&C=*#*143MD#FC T'],WWOP8PJRP#VG"(\$H0RW:@>/ %69>NC&'^*ZTA
PX>&^\ECS IG#DZL'C"_\1].6V,@PB'W@WJAOVM$Y).(T^NW?IKG-3N<CAO\WZOP&
P^, O [! WH*286#0G/<+Q>P4FC?1R$4=$4],/!EUCZ-C9EWOUILNSHRM<U!KM53%
P,*(L*5#](AN.;5C-)Z. A0KK^[_80F.WFIW ORXZ0,&OI!N:?E#I-+#PQ/"85D>>
P#L#>0I]*K8:5"I1TV1SWDHQR$Q&K;@**^>27*=Q+U5]I=1O?P8C-M4WKLI,!>WNA
P"SO"[S+J.K0_AOB"I^/K\C%LKK80=:X\NICJ:<K:RD0+55>L^CC;<VM31RD@LUO@
P)W3M2-"6R^WXLGK[O(AR81$*KRP$+4Z>187&T)L?\FT\;M!O-)8MOL\U/U<?:K=9
PRT%5Z&;T[CH#GPL9(#*XB/14"QK=_%EQU/J=D8^]$O!P"AS*:M=O^7)5618^47!S
PG?'A)#3U#C1[Z?L6EWAL _MJL3<7VRU(%.U%V":KO!;"R:R&^?IU+6;22O0EX$[Y
P3%?:V@(OTVO=&Y*[YE1:=[C\R8'(/^'R/,S+'ILMP)WF.[EHFQWEHK$B]42?0JZD
P[2Y&60Y^IC9#^69,7;_#PR0G_X\Y=#KJTB[L4/:+=4IZPS2(03<]MUZYI$+^/SKR
PF1/_[&97%K4A[(>%NAGY<[*!*X=E0,;V$3_RO&!2/61/@K1C\PA3)>71'"9R9)4'
PL.Y6Y!7'^O'9\)?^.TN$C='+9NM NWY+T_YMDM1S:NKR9_'^KPA$A[">5JABS$[Y
P"79DSS@+VKYXL Y^5)/3I 64M\=#A9:C1;LDVUREV(Z-E9Z6D'Q"#Q?(40JL$K;)
P2J63.JZ'J*6(/1KG-,W/@V 6X@#^"0$(:\>MFM* <,#AJ&"JF,>4(46"D/778F,?
PNM?Y'J*?__UG*<A&7OE86 "14]5P/S&V/M?=Y*,QV( Z,W+V)Z'J]C72IJM[1V/R
P@*2^$$VG>8C$ZZ'YX\$67FI?Y%"&8P[:!/JN>@6ER+1%A!&_TVK073!D:Y8?9O7>
P89T1-=K?_C4(7YY,-:[(>;W"[[-=ZKUITLA2EI7G:H#4VFQ_ZK"@RUGK$P$*#M@0
P\T;<8)0"(Y%BO#HM-<'6:)".2X .Q%9(?Q0L+L3)F$YA%JS1TIK9(NH+'*)&06C<
PFPQ%7XM6O4KJRU ^!300S'R"M.S:Z#$-[E K#*8,J1B128E?N3GV3NGXH!\[H;3M
PE]*B2DC6?@@<O>_-TNL12:$(/DQ I1B8;N%K^^)#7\%D/U)?E/85(&$_0$C!8WP\
P@;PA=LJ(RK012X#W?R3Z*ZU'[8^KIVD*?)/._+_H*;4UY4<GRQNX<HOO#I/&42LE
P8JWX=<YVY@-_4#E@;'ARW,?&V1K;[O<%+=TQ*RD[X QK$1LU,=**EPY<VL$C;2C5
PPVJCY>,G>V^^J;$^G@-?_8&$Y&"?GO/&( =-0BD#C4E.4EY3>%D/Y)HK%M#FLSB?
P@%F4O.* G99:_;$ M22^'<7"TRH?3,%A#-"YTFQHN]VDY:.NT%@OF0-T^&6G)Y;K
PHG&"ERD]4<DT)O_7"^ 1S=K#N0YB3/WS$&CB9.7Z!.L>MQUA5UB-_6?JV$!EB;*9
PN^52VA.WQ -NG ^\R>VVYNP!PW=IVU#KC(VB]Q*S<*8KZ\G9P[H5X;'TDQ0@\6:W
PFB4/A/RBU^E?>)U$]=B<O/.1/#V3@X@<.TW0M24=CS%?))-=(?. 9$$;8YV"PFK\
P6U72YS$)6/DUF2( MUP/? E?Y8,P*$<&;/W8Z 1R1$=30:.9@;AX'CLL87U*8ZPO
PYMI0T2)PKR\7-8A,#Y)Z(R;"2"[84[=X;#A10.;]&BV^F_(-1/F&QYF^QP 0_O6D
PJ,J^4WSDLZ]L_B3V\?MHH@H*9LYO6J^=-AW/0.3FB?TGZ5:-%KT-!T)9G.JP-'=5
P7SWUUWJR5)%XZI/O[,3X .-I*=-_?55<'Q/(_1&MX>R'B+%7V3M+M&,^NJ5S[P* 
PVVI1%"U"MS J<HNR<;G?GDZN[;+WVLU]%)EM@VNJJPVER1.DU+N2KBK*=FC@)MEK
PL%:#D(?_T<&K);V23D3F9@$23-3!%"\?C23Z;5I0RG1E"_TNE[T3BM++10\2DF6X
P3L!K /]%*  8)E<[WNN/1.A] (K(O1#*[:8C9:O%FZ*WH3+F]YGZ>?9)_NL%XG[=
PP472!CV?&^3/_57V8GP/VG-'MJ=UON$GZ?\G#4T5U'-%GILBN[\%GS<^#-W795CP
PF#1\Z2M$:!H!B]W9XPEZ0BR%.P[>5>5*V>)3,S5J'YFFL\99FU5OED3 WRY6<\;H
P_2,%1IL&JW*#<I=U7,[_VF]$DCX'$HS<QZV//.II1!Y'0G6BJKKQZ)\ \L=^"\DJ
P7DFQE<1U5UE!QIFN00NOD<DYK-KPD=&"VYCE+S/]!9DX[_L0XCFW0O'$W5%(\Z49
P[.-AP R<6&IT].,A:+,6B^ZJ-,8M;=LSKD7^?TA*'<A&RA7L4KK\U+^[Y/LI"OEN
P>V)>=JU-$@UA6]6OLY@I?[W+,4$K4?6QZ_,<@VAK^:3.G(NS<@L2CC1XU?3=3;ML
PL<::Z.A"\#630L5SHDLMMKZ+.5"K\F<?+H2M*=1?YGMYA6[= V.-:/Z^;B3T_10+
P3N<S?X1TC/313 PP0Y(JU'9 *R@BV_W&G-457IKBK6E)@(0"P*:=-[+-8GW!72[G
PAMHPP_:]9<#P']3\B8A7Q.W2I.[="W@'9(RCFH9#K6#3LM'^1ZR1VJ2B?!QFYS=F
P='XIRHXZSY9&S  EC30D2RQC,()=OG\[U;XU](S##9L-H?"$5UI5V3@9!&*./ZE?
P?-GNC6..KQ'/OW&_0 PG;+VH79#<T)T=<A=9E717Z(H/]C:Y@75;QI+UV=[LP2P@
PHZ'WB_\X]>PG5M[7-$DAD@8!B=JE8LODF)$Q^I[6Q$LS>,W<**QO.A86.D4.Z"M+
PCOC*5+@^K2+;#R<Q8"ZAV&ZK[(E<5>4IW+>_F2-TGJU>\PET;4R#D]LI&5?"$3&P
PO8.1;"*U-O,GK_^LFEWN3'.4,U.9(.5#6)$L@=(70D"M'N'X?VF'=AQZT-$PI^W_
PDUPHD*.(=<TO6MC;LJK(IK>5SK6QBZAH-GF":5:TW A-VFW[WR -N$$(QH0(%^.9
P"7D+!>\5W"UOL1OQD!WX"1EPRAXQR:N"F*]0#5#]QP\O)$%55_$Z3"F\*K-2\\01
PK>18>1*=5@9MSE[+JS!:0C .?:XEV:Q6^BZC/.\5")7?FH]/9S3=H94GLQVY!F;"
P'7O&OT4N_[D,A=Q$ D=4KB_T,];1*"@ B3//8XB01-:.I__4-1!&&<N*1N<Y8JKM
PSD0(EJ1M7@-R@TQ@".K:[DT0&. R0!!M6:7[+J:3!!!EH$;49F[ 9>>2M ZO,)1$
P*V0L[H&Y^.[=82(:BEK\(5U%9OF?TBR!0E/7E7$+U$WS\VV[7QY)Y!?$NVQ98KF'
PYB0@ &BDFOF"C=95HU"_PXYBZ]/OV2('HDD3'0IP8,W3>>>F2_$:,#?*]=-VFGR^
PRTP[B [C,F/&CI2A_A+0J-.)&E*5\LH5GD\6A+TC)L^%C*E])O;A??.U<:XHNX1.
P+#=4W%ZW7&/@)]5;&6ZN5?-Q+.WKS!2JPG1=&&]OH P0,A,<.(%-A:KTKXDUYCW?
PCE=[SOR;\B1$2@@UTQT4OH*Z$^(R8!!A?%X*&='7 4Z8MM\$M'5GTY^4C7T_8B7-
P89N+#5D]PJ@)16/U>IQH-?,H]TYYPRW$"Y!<G)Y_[!JRO]SDH$,9;P)>V[VPV("8
PC@<)TXH"]WPD']L)THKVDP"H9YY ,#PP>VXB&*:>@CB%>@R:A/R0_3&]H@%L:B+"
P4[H4Z%V3AB.Y+'Q+;T!;V5@G@O5.("9^=!HF<CY$]]&K+PR%\*,#Q,JLE2BMJI4.
P%HEG#_=AGS\WH:@].Z5/$GP!_2 YICFP<')%@7(=>PL)RVEC*_VN7+TLU,,,D%ZT
P,?%RDN_G./N='^U)M)1)QH=;UQR0!L%CM]!"&G< 9U2?+5M^HS,!DS*TW?61VG_!
PK_8_&XM>-/VM!-I6TAI,++20IGJH4'ON6?2/DBD0&"OAO?L!#$&S-/7EVS=(H#-=
PN$"2[J&5D1JQ4,>_V$B+\DEJ5T:L$J>!J[JNR)#H8_I4PS2]4E8\;5MIN8"!OQ*P
P6?0LYP\6S:%IH,)+]G-^LH/$)!_II8IL-2SH114OK2F$"EP.@-27#Q%U8^85Z;!0
P)7W*+-1VNN4\#=ZE[,J5AN%J@-,'4C\!>$V:-G8Y+D/9H8"AE^V]SD#.L^2V5<X;
P"\97:5X'F[V;+#HB"N A#'(#QO>7X)H5*!PATQD9XE-M[-G8)9K%J NA00MJ7R0'
P^O:U4"@$%R*H"EEC(-\NH$+JTH(;^C2/M_6GA/@P64 ,)Y"C@12&HO\:?9QAZ\'*
P$A<>%9T'*K76ASM2M=;90["H30\>/;B_@#IR\90,;AHJSS3"1.ELM?9*:L:3I@O2
PV,Y9^U$Q9S_^TS&R(FC3Z<-^YHPRH>R7'*2[]3&'X;),#/+294T/6\_$J+9Q"O:@
P[5_;A,@'OS H)]FE ?+OQ=GO[.WL#N5=#Z\,JX)T*WR5/0P?5I!B@)HF4"DVEG;:
P8J@E4!)>E?TQH+9!D__R+BI,?=I'1CL"#/.ZW0M1)%O[VWVRV_W!:FVB'6GT*&9>
P2,%NX;GI<VZ8)5C4,@Z]N<<1GHJ_1Y:)*\-A\/&G$1(C_0S22/J-51H6-'O3+$Q(
PF# ,(7E(X>T/KC.+] ]=U(Z4GA41=A/8;3Y'>4KTGGZN*!B%&C["=3NQ<HS.S8UF
PO)M?:*?IW,\3(M@@2SGB2D<M8:71"CF8:$R5*/0"U!DV%B ^WJ&V7:'Z7JZC:VP5
P':=TOASL:JCDJ LV3YA '9)2:]_(!$OHCT9N+@>7:?"%ZA R7=\D9K5+97XZB%N.
P:WGN,V8X;.XM&_,.AG,Y*PD0,GN3U _J_W.6YK4GA#KM/E(V,55KR.)0QY17T0JW
PGW94I L:>/2Q1<D.Q3)NH;C#<3#PT_71'@]1]PSD9"-RIH8@';)QI2?8Z>Z#.]8.
P6$/=^'09(,2K*%"7\G.MP3PJQW]FAB&_^F!'H7RN2A63_&/U+&!1]O'DQ5R/IU=8
P-W2P@B6_8MYH+GC83[AA8/MLCEA:&SW></9DUZ_D- 49K^/= $5'!1O+SEECM6M7
PKD$Z.&%]P^Y(OP>O#18W$U6H\'D#MN^YII-BOKI2XLON_5QX)+ZNWF20$R)!%4&8
PHHBS.O+?H*%.>%LLQL8"OUIL_+NOP)B0"EH#^<"R$N;(UI!^'<H26.0$FQ0L7CNJ
P]L#N"=_)SX@Z)2V<WT0WZF[%?M,+I!-4Z8:ZCT@*$/?S7[!F2P1!>$+]$LJEZ,UZ
P\3T,^"NV&D"9$TG5,9,\VRR,UJCX4B2W;;_TYD^K/S@FU7AXBUJCPJP)?]36TRKD
PQ-\+#JV^%QDC.BY^!@<&@OQO*"5%00SH"2@3=G[58KHUF$>@5UFBW_IB1G&SNQ\,
P3\\?LZ1ZQL1'G. 9E;)Q^S-GU]>N02O)^"-O)>ZB^TQ3 TM5?2PM745Q.^3>?Y+<
P<&8WD-8CZ"U9TZ*?8[)JU1)XW5RI4.5=FDH?06ZJIS#E:+=AMGA:F2"6[75V*FXJ
P&96$OQ0'AG7$"%U"MDJA'CJTXJ7O![2N+!]7]+F\61:I1DX<4CG^2#3/BH(QZ89$
P=8]77#4RRX#&7OV=7O9(N"0\C)'52.K9EEFH#]A\^6;C8B8:V2Y8^C$&*M4-"K-%
PT ['_(I._%%(EZ4#[Q5S^V%P1TRR_FL69KV #W7C-3"!2K@#;& @N;DEVI6630C*
PJIC;.@E,0A<9*JA::Y*)XTF*WI]!F)A_AV$@:UC^#1^) )KQ7?WSV-4@W&9WO\M^
PBC;ZKFIZ0UOX45.>0C$#D$'*>E38\^\A4WB#\94\YL\/3"U8O0H'('X%M&(L-MM&
PI9D[U9?>S30L51:+1+8=FL!''O40\MQ!0$C\B#JV'HY'O;'@/B#0,9W$L32=6'J'
PF7E\*SBF"Z(9(-%E?X3#"_>;]TW747[BFRP:=.IE>O3)L'$_5MS]3NT(B7#R!_63
P13R$RV&UOE/2/=GARC[EA<#S18WK2)INN.WYN+6#KAUL8:([)!C?-F*-09=5U>#2
P-B,(-%QISOXY@2W5V^9?7U+"0%&K?JF4ELF!9O>N%-%3W#R$E]=MH]15"#UL=:_)
P0*I6$D-"*1.$^RMLYR]-6[59LE1"!"-C,46H76$M+-/8TZJ/=2;[@MZY;C13T14>
P]=W\ZY?2X&CKP#2X3.5&5'F*HE,/D<@]Z;0Z!%?X&TCN0O$;!3E5.61<D\COF)5)
PCB(N<1._H^] \EL;J32^RX"8)$YA)'Y9J@.7OH$NCP%0/!!;J>?/#(9&IL[YV [;
P"]OPJ"HP4)\NQ1L$:*;.@T9,^W168V0%X[Q-C1^/$?9+AJ\660S=MY+:#FP"MW-L
P>,X\6$!?[S39FNMU3?_B,H!WX_E@:Y<!*>=YTLD CWD=6XHRQ# C_@M=!^TJT:]&
P:6V" OC\[M$H?ZB6'-"<M<DB1H,U:;7*>+Q,^]TMI1[_;TS2Z+:D?)(2!;5PF:SY
P.:LS%A$E4V1Z-V5R=!\**WU8OU!GH=V$+&@A]/7'L "5W7N@D[R](O-EC%AL8N1Z
PV<[5!>,ZAT:I#A,CT]%E,3PYA:;^4,+8K$4AT^+4L8&RC!*?;2FBJ.G^\.T$G\+:
P9R*M)H5$8B"<;(&.77"L_R_D8]2=40'6C9WOKB02>1%IE9=TJ9>H_$@/[\?;/E9N
P]M(#X-%A10%K>1.W$8"98'AF[M\6SB%,4MT&>G<?]R^Z0/:BT>F =!&\KH'[&4JV
PJTZ,2B5..(]=2P4GM_,!Y&]-XWI'B\#E]%:9RU-/W,$-9GD,^S@'!+DIU[V"3Z=Z
P=\5_J11OQ<&0&'1GVF0_3F8I\:69Z![O&Q/'O/A5EG;<<C[T01,:E!&15#XBI ->
P6SAJV'@IE8@X:@]F[] K.?JQ^#2?)WT66DG,=R1G;\'&ZF"+JV1A .^W^+UL 5IQ
PJ;N,LQ*P%G#7V)^YF_=].=Q)[;#. +"#:5/9(36RWP@C5A:NY@C4VCW0"H'XIE3L
PPIG)>"6X7##!:)X:UV,8]I8FA[Q6(;G&#J2""?XU,+@1T'("$FZXL'OIHQTBX$FA
P)5H["!ZN-5/IVIFJ<,S_W&_IHF369/Q8>AH%CRF^K,@+Q52;IW7#/U[_*LNH2P/-
PA$>=[KYC;=<>_F\@J\5HM/OH^NF/D@UZ[VV#[)3$6-JC+$9Q?7. NWC[X4-'MYN)
P*T1]/.C]NFR#/R5)]R9C]]13,*/X'X@Y%(U;)1IWIQTS<Z'XB_1!]DCE7[;'4,#.
P=U6S8W;$S>B[ KRONZ12L++Y;<Y']X!]^9PDYXR.BD6DD/,,*6H01$LTL:(30L2Q
P)BZ^JR3>=8P7.66U.OA0L>E>-PWMX/O=FN"Y"M[%WBP'<>#5PF0'Q79[&#6JY.MX
PM#P$=V&L:>PWNTL?QF2#!6MEE-7-$D19>F_%6#/BDV6KKM1^O(K/QP(V'Y5")+S:
P=4D556XZAW&P\*I[N72J'QD=TRR-%B8?1(UYG,6);/CF9:UNXD^(7+Y10](Q,\,_
P'6#+EC!U M+Z[5PZD,\8,2<N)PPP?G21$>M /^27 9H0$##+7^V8!!Z0ERT!JHZ:
P9"0<B>RS<Y<[(6];_MO[(& _WJ)I7+8!#I@)DA$Y%%A^[,\#=D0^J6W5I7M4<C L
P"K PXF44/ZX.01:GIU&5:MPH8\E)4%24/]QYE&D2(+;-]V'T.@A=NM1)4W,X^/,J
P:#]/P7I)+O+:U"0?8>N6SM)'"ME#4R[F=?,\8IQAC%<GB7R/-\N*%E-M<'TZU*$<
PV5S=,/)9(>B*@8W?&BOXZYM(N@*8,R9:35<WCJ@A9\V54^N?BJZVG%O@K7S1:F[\
PS[%61A@AFL+BMBFKOTO,,B_Q19D+/.1D7II9,D"C7^+W^K/C8,HN&PA2V:LFC7#@
P:/3IJLI'OPJ-6DEH/F&3@QI*"-)A-,V8.A%.^LO8+SUNJ>;VBVH&"]TAP\NO!*YX
POSQL-7C&DZ&V\PZ35.9!"$60R&7)1^J$=_<2#O\''I2Y ,#><6.98"GGUQ2=9*AE
P+=1I174>0!FML%)/K:#]_$4%(P?U$^C11#$RV9AD1J==E \:24BS-F#S@- "!SCW
P3TO*XJV=AR.[?Q%9M];8V.1"NA!N^!48SU&C+VT@[A4M:H3CL4*ICV"\5AG$$0!,
PCK+SGP-W[ (P.V;)*N"-4R@%$J[6'L2K &H^PCBBZO:;L!%[ML91'BEBN.7-#G%]
P-^Y(P(<<K9.?,/E$;B*U:I2K/AM\U$PLTS3>D<01S+K7='7%8/Q.:JW1%@ANW&H2
P1H. W2!OR\8-4M:CB&'.MU;A=E79IUUB8!G?J0\WM##M=DLN_#1D]U'=,$>03AD4
PZ)+L7L6#IZ%.PD.:U7<G3-<%#4I6]@'!0=NU<T<U#I[D;*&, \<M$4\O>G,]M-T%
P)1"X@]QB. J\(WR1$N<GI020R8[8%+F*+QP$Z"+R6H=/'%[W55<R.\($BE]"JY-N
P+WA0;FQW7%//P6:_FK54V],PM\7S 4^=2T;Z)O>PBF.)1\FD^ E^!$@/).)N;,U3
P<%YF"#P>Q]_<>Q$<S,1SI=DA.]\8<+'J;&0UZ1^6TJV*?Q-;YH2CN3*ZOILSK\$*
P+\H!L<F$U[$#$@KJ-QH[FA>^2;<WC:$&>&N>C/3.EAA!Y+E30,X%LL5-RSHMR@ I
P1V%LR<R]AZZOVJ)D)JJ>;3@\OR2MCZ'\,XI41F\0K/NA=XT:\'7OL_Y1AYF%5WL"
P[HEHTDY6W9;.GB ?>E^G+^\D3EN(E9 !_*-C3B,+#Q67@G2^Z.@PM(%?-D\$E_KN
P@#ZQY'B3&SP7=-U8+ <-:.$-'?><S($=\3:'$"5ENC_D6 -8JD8MJ6I+XO>D_WHV
P]8WK)?Z@IR2_(523!IT_0IW$IHC_FADU)+>'.=QVWA>H-*A:(EUIBB^^_!U.?]Q)
P:;;OCB/U4'VSHQ?<:F2-B#'6AV:W>P@B*,^^@.X<;L-#C;J-QC/7DO"N;6]C2;,!
P 7 464YP(.QA;AN6'\OBBW8%O%?,X1AK<^P?OVG$.7N$@-(!;2>AS; (B<>C-(RZ
P#>Y':BL?.GQ(_IXK8+V$>**'OA@K[B2CLO=6'Y#0@/'JA<.[ORI6]"\(92F4EU> 
PN?;>A2_[_6H N9??EK$P*]'Z2BZ\*(#!T>.F_I"X_;=>NF59GG4#X?BF8+/9#,)Y
P9T\NEG-@NZLZ;5_T2)+HF3=M!R/#<>"SN.U7L/@0(#!TATVB)N0-BYZ.)+)4I4[ 
PRH\> ?4K+#1E):1?$Z7%=S?:'AB)5CQ[$+B$]$K"_"O=W=<U\^MEJ)\_B4=:J&6A
PC61]'*&[4VI10U8,%'*AQO=D=D+K[2!-34_VV+I>^.$9O7&DR?EGA;-G)@1X^EU2
P5,;K08C,(+^=<+_SUK07X?&[L<[B94JTG'RE(RAOI%6,"ZZ"23&>]<^N\J=KG1H3
PK\!L&Q$H=O(4JR/VQ]-WMXZ1W_U'FDP1^,YOR"R4*@W.Y>U^9&]Q_8E8!ZN&4CX3
P%@PC$#@4**TLU-7#X]I%[E)"J 3F(DG-'P1B\?;[GSNQ^X-@(7Q!N,:S"HV@YU#2
P+F>ZZ>9_U#@QE;8E1!/2/+$( DB9U;1O_0R8</\!:]V7A6(($IL'!DB8"=YM6B[(
PJ@Z8G\WE@R;85S&>_&D-9VGEU)4,JC3* !_A^7BZJJ G^DAWG,EUM\?!4SU+J<CZ
P+$ODSYQ@U12B[>=5V4/]^>*K>4VVJO[4*^%76[!,8)8>C!J*S&8YFT<'#W0Z+3]I
P,AD?)Y1/%")(,_/AG#5R"5]] ( 0Y)6!9O7M',S[Z'(Y+733MA<(A7A_#.@0_>0W
PCCHE>S0XAK\SW.+%DR_@9D ]+9"QF&(FNZ\5++,L$TA=)8Y\98XC\F8CC) C34/K
P%*0!Z:9.)06W:Z><7A2+L>4;_E_%7(QT# /,Q9%26MD$#WZ+%2NL16 !$N[3"($;
P])VNZ/F@M2RA8W=&;LN?XDL+<^S<.J]4)]M-,3W#@.I.-.I %P-9)TN_(@ACEYXQ
PR"P ,Y:8WRK'T]+O35+$5B4UI57T!\G& NVZ2S9DA?$44T7ADM)]IS!2)*I;0^9T
P,/4#8.+(OD'3"D#PJH>\N@%AZDMG>'-!U#K"J>B7S(?X?.ST+7P^)$5<$LQM+?+P
PNOC[#'A;L^12+Q\@T*\%1:P<AQY?][\+F96 EGY5+R^3[]>/0VI799AF5TGE]N=L
PI,EQ4FO*':!7X?O=:^T<X\HO ?I&_L;$"Z_S>UIN2:\?<I).ESCU+]XH\;KH2<3H
PN(_5"'-)+ X+E7D8YCSG,B\96KT#QSTBW0VJ!4A+;W<-2*M0%\A<XG_0;EBR0YZB
PZ8<ECTI=04*=B=!7,S_SW.G>Q.NLM']=0$]0*'&*Z<T'MO; #6!C';B<"["_*@UF
P1;U;6S9PTE7XW?7OT.P&SD:.]&2_G\.)BF,4_TW[%JAL:F<X!.AF\M3.E[%BYF>V
P_-B2JK?(9OR3=2;C<ZL+8QU/3,Z#"UR&4:QLVV=J%6;EGI4NN>W.%A?KW!Y^GQ35
P<1V^"^K)?".K9G1(8C8VMS6-U1WY9DFS]>UUX3H=H#9LGU 0ZS?VT#M I8\&X\7A
PZ0FER6D]Q>IJ4@6=\&A9)&N&;[JHY)5?Z'*F=5\]W]OZ436?('.=FZK@Q428 W/B
PF'XWWY!-61:FUD4,3A$*+/,)AV^JHZYJ^P+$YP)=FDH<D:=Z!X]8"'MU_[6O(+=;
P]:B)QS\PKH*R@TAS5P4"2?F=/]V%,("DFV*!Y=[]#EZJ-&*$"1ZPS]"(>8-HEX[W
P.2%DU5-;E</[D.4K"I--+B:H:H^^\I"V;L@6P_(T;'M&!^I68((&$46\N29_= ?J
P^"]Q*G1M7HOGH\09CJ(ZM(A85[<_O'OI ,(>ZC76G:R&V>$93!XWVLY6=ZN 6B5)
PBZ Z'(.N3)XH>\3B^HWP$^*<3+N-ZI(+HSBW5@:%-7F%8PJE0EDE0&YD1F:OMI=K
P$JLFL=HS6311-TI%BY0ZN%#Z_"-UZ#*)CLP*>#=OT7^XXBI.-?L6%[2E]J[]2EU7
PR]H="[NXH%<BS34\G>R>@E/$'-.$_#&R<7GYQ1_W3N=>XTAY_T $@<^=2;'I+.;+
PP&J;N=1!>#Z,Z@-MCH)_=ILZT19'H \J]K)+X[5([2GTG"JI*DU02;8!5E>VH[E"
P9+L8(DDE1)F-,K)MQU:LNH1_LF;^SV3)>/'DSY.1;$+O(-+:R0]VG,?-0#094A.L
PV,7G:,SD";-G\?%4=9%F%9Y\7/"Q85&?;=KB8=1EI! :N)0^'/). 'C^NQ:AJS';
P@$PI7YZLZ[D;NPR1Y@?DQP^B&=VHG8;?L@H?42,#&>*3!./P>CIP_@W)5-G^',"P
PG[Q;WU&0&IN'Z1<)*^!+'I)C&)T'Y[@%H18[S-3T+4G#)N,GO'@%DDJ:.FA06PTP
P?.T!&)*V.JV)DZ?J(T.WU8UK(6#?;@=&^$GQ@KXM@ER8@[X$Z)OB3"=GS10C;5@(
PWZ=2F/!Z:/<G(0!WF4Z 5VLDS2^#\VVR^67+5R*BVVC9R_#/7QV)\<1GA4*,CUG5
PN;%1EX4#BCGB2QEW400G-\0+7W"7%'OJ0MV8C)<V?C1H>C<HAR4^OCA!^>%VD-GS
PI$"P=?7@BX IZGR&'^?.5*2>F=TW&5_,971L-<N*52$O'>[CIU]0AT*9Y9MO9W$T
P.>]\APF#\"VP[0K?%R4FB5\<=1N0E8_=Z!>']="_7 ZBYG-P+215'+]W4'9@6.'B
P+L>GV(^JG8V73<'1RT&V>O8C%RA(SO8<Z\X/D!E=A[B7#J,\K&).%VPJ- )E*O:E
PO>.?4RY&1N;5MZ"C>FGG/1T1-:[B,H95++5+O+"=>H)N^2>F#R((H%L_U%NF^3S+
P_MW]=?.VF"I?35U]\"M3@,J))Y<]S:>"?[/=(,UZ=+W8D?$;$&R\;_YT.712\6"B
PECH34#\<I-)4%N!RKCG=\[J7Y6[S9B$[YTC[#1^9<FQXJ!ZKM2^8NI\!_91N@L6[
PP;#W32$03G99)\MK=X!"[)"^,C#GWO?Q!;/@K!8!GLS++\BYQQO1YS.[TSQV> 2/
P@7LWD5-OHVG$&#=H9N*T.-5L&Y@)AQ&,<0!R78CRY;"'V3:&3H@Z5A<7<S^.(,:9
P_VE3RP$:C\A98'.EK&&W!F53VUR(Z5B?XFD%T=&.PE*O?MK;1.Z$1_F*U7UA[OR[
PA>7HBO)J=CRYH[RZ!94@QDSK[/?>N#*2A.-_O2+U(I"DAE=6--"_]L6,<"H]U "U
P)F V;V[?GB"&DD^Y1:-1^@"@OE\1,-=5SM1W$#4.\U["P7D'=C%QPC.7\4'18[%E
P5)VK*3RVXG2 QE.B/@X;GZKI-^NWE*8/H!1A^&(MP%^[DHT#WU+ZN]S5J1+&K0BS
PPV%RTY8<^-Q 1O5VW^9+1\I+9'V[#=]E(< DO?'%PYM^I@]P-G[WX$_U&\Z'"U>W
P48K+4.E)AEZB2!JV!\-Y:)=VP?._C2A]EXVW:9BPUKE%Z.IF,N*X*\7P$E6>=M:]
P^J[C2H6HG ^-SQS_85I]?*!W0IM%J'&,QDUW?-FGI,.C7GVNO/?^($X3NZYC/M;R
PLK05M9\J;'^/=/OZ'VZXB2%#!V_Q)K3)?0&\(E8>B_SEE4.-;HJ\\7<M1A0U&_0&
P2AZX)RT/+,7$Q[P<E2:ZR8*.B+.3O1&&ERDMF\$1!EM"^</D4S+RE,*2972A5PS!
PP<>3(.GH#W*(9\YUS]_765?-N''OW'GQ? @(;9TSE9"^[?M!*=\$47R9X]KWC33M
PX9OMH(+'MF=4O95I0$1X7."WIX+V"")GH)([]NCXD9;UJW<6Z6)PO<!D\>Q)A'W3
P,?IPT6ILKM>=QN_U"7AGPG='>)IRQKQ5%(UFO@1LB.ALM_C&Z5..2:RBS\)0XRCT
P[QOIQK$A%4U L]9.,/L 51;W3%AYR8+68<I(7P, 28DOHA<^YN$1OB,P)*!$\FMW
PO[7$A.\M6O;8BYZ#_M9#]GOMZGUB#V?H=3CD\5UHSOPQA0&VS: \35ZP9B0N2X@)
P>>W3PY JETFA)?4QUR(_4QTHO=ZO!K.-VS(\D-&__"+U5QYA_IWE30S 4M)*]*DM
P+OA/NOJ"KN7Q_X6+IHSOCBS"[P:O'1Z/:Y-R.S#"=YW'F$4.",NTW8'?NKJ,4V7N
PUNU.2(W[83/L<=%AV!@]VB6)RN.("GH4Z$0HL5M!6(T><24F[R/<I[]$$9>QO*.K
PBM?*@%KBW4ZEPR.5G(4@;%8%$\-Q]U-&5K6;T':6Z4U!>G2UY^N@-D_O>[&5&V%K
P0BSFJAFB=J'B6NA&FNN5BJ] .G@.?'M]<SGV&^@9J(A\D"#IWS^"]$)8#U+U@A@+
P=JFAKQDI_$E$ILOVU$CQ'BA%/L"CKL[USDCJUS^)WEZ(UMD%JX)FIT\#&]!O9UJL
PDF7V6\P6_?<H^9G\-AK_,.$K:!!/_(J18JXW.@_I_7XI(H7<*$0'8"M%<[,9,I2,
P.@ )"<H.I;_(P-[/DG@BW*#B@CAM=^=(OQZO<LM_AVXE-_04]J#/DB?.OL/)QS)+
P[[KHTI]F_LA!S92C\=MMXK]4EVP)]/#X"E>FB\@) BF&^JP,10;1*%+QK,":_PYE
PT2\U91,K[-[<]OA[B\R)?)_]P S;!2,"@.7$HIK)L"$8-=LB7 ^MEM058#HOF_>_
PO<M:,AMU0LKEY7^C]OW;H[?@90$MYZB<;EU K[Z><CZ:S")6A:YI_H%+"',?2MJK
PL$!$?7#1@7A@QBFK,PC8%VO?>>]P?(00'%&\DIC)2.+4J:U1S*O_6%*-))+ RH<-
P:O/#S(\%%YG;$637[_Z:^JCU9'CK</?27E[&",J*]T@B_40.\:KM>+H6A/>QM^<X
P>-J,>Y^#7UQT;@1:KX-[,SQZ.0@"WSWQDEH:\"^0DB\(PR9:"RL'XPG&@<Y7?W#+
PWCI,K!"L?@5')+8_W1HTMW=*O.')R\V6JWEV9^]/V?:<@$M 99BHUXYT*&D;IRQ4
P$I2:<O%E#..<&+3JWFF]&,7=8?HU_[0=Q&\*R*EBS5^7 S'82@39W\MQ%76H_911
P .Q;.>5P2YU+"O V>\@^_Q<92DM>7#2$D1D!5[9^JH+SY.#S71\UPQ*5YD;:&Y7:
PV5< GH48B\D,)) ]JLD^!2+V\0(G@*Y^*YL6-1Y(32##ROY53T^0F(7@1&>2G@Q_
P>->E3_C^?[B 9GAS^HST8^Z2HO]!N+5MG>]RW$<"\P>,CL4[D(31-TY>:N-@-%R6
P9VBX.U] L/(*& 11]2@\J(D>AU.C((&ZY?WB:<!4;%"&/PSH9ZLK@_1=:E-4!MC>
PUB+A,97Y^<^?@%'"/,'K<9#LE]<: [\WIGR^G="UFX@Q+KX)/\BB6*Y1C=L:O7LH
P?E;/* X>[4H3/12.25%&@DX_8Y1#R'!5C>A:&4"?+IN30&H7;0;_+)MU6'6$1Z?<
P+0]4T-X4E3,N$RRS"*";'W2&_T).)B2SY] ,3(XIQY6ZF>VS:>8 7Y]WE27;)],'
PK->E '?VU22OE$ <B5ZOO>8<TYFB+R6*I>2= ,!MJ^2A-QK(\GA-F:$:E+M.7,9Z
P:-;I;N:F-J@/+U\TAR1K]E_I+>^(35'1)(9N,?P[J[1AJ-0QF1'YNQ9(CGAW"(X=
P'BD)P24)S1BL;XO_)YV(H-"3W(RU4RM)YW3R[4(AG,]F%.WW8'V-$W;'"82>.GB$
PP.^HC&BF<R!8_/_9\)8[]U._^O$%:-1RX<]_I;*%R4?60/(4S*V>"AV!RC+B9H<1
PVSS9HI4.Y$U[CD37O0+/G=PN:YL8^]K8U,G#.4$5;%$Y^&W/H874PA23"090G'=]
P2U&XV.^"VB5ZQ,N,PQN2&TZ 6W6:(1A!$D@H:SG15L. XUT7"(W-;%YN5/%>M6M.
PS*6K#MQB^MS*>JY.%9A).U"(%>15E<],MHI.H_ZFK&P_9J+-K]A$ ,?(*Q@(H:QJ
PMV:!'O!DFGBOGWXG&46Z#[7HZZ$U>8S;/Q1!]07O5N.[KKS&15+Q$+ZVNLP#AG\<
P$\W:Y&H=#N[6RAQ8L@5_YRVK_8U.G*^+@ZMQ_1Y]\% ](H.^NK^L1->OVTXA!PW=
PCXR:09]:5FDVWBW)D'U@P%\V34Y6<<NJ6Q=U,$+*T"%DAA;MB:6D+I5FN^^R)QX!
P8.&'4BY.VZOU_AN>3E41=>&TRD0QE+,EL_@R9LUXKG9OPM<G(F ]VM\'J%VIC@N^
PORIX<@4LB!8F27<%.4PY"R3Z#+_\XJB@T@TH7]%'B\#ZF_P?5N/]@'HX7G[JA)\$
PK<,7W&21730#JT,-(TH\DF"C&4:RTR?!I9!KQ2%@0C)-K*2U*\:0@%R3;V4Z[UHV
PLW2B_AP:S%\DO,3!2'G%S%*4/51BN*5@N )='!SBP;T;BBX)_2[-:,8G;J"G8*SP
P @$"$]=[<==&HTI#!.9+O$7#K</1L#S.SBN_?9B"]LH9?N+DX!^7;P#NZI#M#)_9
PFF&X-UTV!31$*1,.<K/'-'Q,R:1:L><*1T^,:I7=O.=)SPZT52)^C^$9:[N,2"FW
P@%P/+F5Q+@S_# W8=B((G(%H4W<SQ_BIU+BJGA/P,$ZTGO6Z+?]K'11Z>.OOIJMI
PABJ5K:0(7I!8,:3E+C[:63O@P5U6.-9XD^!$?9]8E.<]J[Y'FZ6'VZ=.OR"I#H,]
P<2]_:)1Y1MIMO* Z[37R]I<.Q(X# !M\>SYVI;Q:0>F=/6=B >#C=/+9K(VL2?84
PR5.=:L^9'5"@21B.=V-5(<U2@Y&'<A.!CMP*JCM&B LJ_1F1*J>;2$%0^L:4&;J9
PTE%BXX+NWAI=P.7Y;ZI2[@FS;]OXCOV&[N@I2GN&J0Y.PVFQXVFE09L7<>G<CU)&
PG+8V6Q==D$B+94"DT).!L8C8CP:G*RP!<(?H"R+Q?B1IBQT(&XIS5F&%OS=F=M0K
P.L()T,8J BYLC]@(YK],I+V&@Z$V<3T*G1U68_&XYEJI,Y@?.PV)X)&,XQ6BT:NU
P<M(N1[=N!ADN)K&79^&]F)3I)!%;%6KU;,:40P.Y5S'V7V53UQSE2Z]ON,EUSY)%
P-RN+: &[2[0XO ;D-1QK )^%2<("+;<RA1 O,)Y >NI*$4$U820-70'CIR5G\<82
P8<B,W1BAO' TT5,F 9V==1_<HI9D'C6UM0W:("+!9AO/4AEZEJY6LO4V_2D:HILF
P&[K1CU.+R4QTI"8SI&?8>^BL*FHIXL5).'AL%BP_4=?5^DW4' !(XUQ/^V9GC"#'
PJ_6_( 4\<N^;:P;*NEC>M0OP3ZROG!.R.\>/O;%"RU3\>V.16_S^:N>=Q)0+N2Q5
P0VQ#W.RF+)#2W/MTJRF%Q&,<O(6,[$A8B0QBZO)'LDH[6$@!+B@?,84CP0B4JQ@,
PWJ7^57N9E>FKB#;=P\**#9SO<3E?[_[:L7/$[^-O&L[4OFJ5#(Q.\0WR_PCL#7'G
PLI\@H_O-7+=ME 5;E,NKR.;A:O4L<PW2W^*+5",=_?\I#%, \-@5QPJ-1#,UAA[5
P G#.P@(=11@/E&GG?&?5G& 6+/-5YU,(:Y "N"B<:2*N6K28U519P*.XLHL)#VAS
P=H %I=A8L+7$)^OD??R(HF.UY#\Z8E6._L/$?:;5Y4(XFWD\B/G\QAM)AK<%[,::
P#W69MKC"Q!D6;KXJWH]78RQC.?."=%$O5G6JH7-LR"/1D;L(MCE2&4C/; TZ%.NI
P^HR[D1;L&38\2YP1R4<B]!7W]A;.YKR,<@M,D3GV2]H^E7M1Z\--"=6,+%VU*03V
P#M#9Y.31A/0%"NW)#&3>%Y_((P%T$H#X,1I+#;H5F/6^HBBFAQT@82+S!)=7\[9@
P3*'+JW%>%?L(S+87[&&'FXVJ:H<0I. W?4[PVS4A.N3DUSS,49B=VJ1]X):L=L*O
P7BX#O"1N!,BI@]KCM1DX*,P3R17(6).(@-(!7JJ<FR!HNUSBL@<X0ZNHCO?MO-Q&
P'$2I?KUYUR@6J[]7?#[;KD0,:9%%<>ARD5HC701PTHL]* Y)/&-KU-5XFZ])(QO5
PI_L9A3O/%GFSFC;^0+W]N9)=-;CV-I33QA@V$T&DTMYT8V73;FDLR_"KMJ(%O^+"
P@.8[6LUZD-HOH(Z)$3<Y%Z^9IS:W3OH@ ER3M2(B6'Q^H?''@I;EN1L?&*)H_0C@
PCDW/@B2J)M(IH2VHM48N*<X\9WDG"LS%CIGG%UV&)QDW^NY#(HF_KNKJR(@:O[_I
P$F37ZPL8;1/6_Q9&XU6L'X@P<;]Y:#G/*M\.C#7-.K2F>.O?E+KW>8*14$B2:'RL
PJ7?T]<433=OX.2+$]/38=205!V- .\HQ4I!7SY.25NR*%JT1CH_(S@F3R4M3KW35
P5GDGY\XH.I7SSBA.1JP7W,,08EK/ V<+H>ZR<K9=)(+,[&Q6*;5]3^-ST<OO0KHZ
P>ARR$2^\T=5LI$79&-D,@TKD<CU2N0+,&6A+B_;MB#O(4]P%7P:^WGQW**V61E<Y
P8"/ C=Q/>G:<P;@=C+G' ]) 0ZO(]/-*<XA#VMWIA3@?MFVR#ES;[7%FE+H"9RV&
P&<ST[?U,^A.KUKGL=G7'FL-1$ 0'$EI+)E@E:S/BS_7)&7&IR+5%X$,0YUMX>F*N
P9")HI=,;^9H:C/8"BV!->3VXT,$;Q;6CO H<2+ <H2JM8(0LJ!-1X"M\$"&"54+<
PE52)3ONO^W:-\A]G&^D$B+^("NM3.GDILG$O)PTL@[#I'GRUI__4T92>)-9S'RN3
PO6[9;?'P5I^YVUI&QT9TNTN=I\'+ZC_ 05ZC\/2*"$B&4=CH5,^F":',=G$T;P[-
PV"+4CK5[L_MY3\'/3MDMB*WLIK7\UY<"A?H($+T3&F3D1<1(%M9:"IVH$W7'98DH
P?W5>22LIM\$?4Q4;;ML<D5\*X(,,76#9 >2!]Y(D57'7+/31[M&L_A11PPAN/X$G
PZ"-[+%.1<VQUJN A8#_9;?ZY[V9Q\N_SQ:JJ/2*'\G?> U'*(_2T3+7,Q/>9O;F2
PE6I21;"M'F:5EI#KOQR"I@/_!1U3?&F*0&&W+;Y[FN3IU5T@\8>=F _C%+C%KT'8
P*BC F_A1>DAW]GV=E[L#S#7JQ@GUS/AK!>&*>BF0,PL6:LA;P!#IJY0$TIPZP>1V
P4>MX[Z3..C<L=ZZ7O04/.2E&9W2MO@FY#;P\B;3OUTZE.&V*<<"4_)1\O)739<N,
P_9I/.E!^OPQ#HH>9?.TA@)I-]T)](@U[_A0? #:"*%!\<:1010,$4=I5!K:L-6[H
PYT4((K]83H+(\I(\VF8B(YP[^X]DYJ!-[*PM[@1\2562\*=OM_.S>R<Q@PFUKA_=
PIWGSA+[\D/(NE?821+XRY]L0;G_:)2I=9,N$#(: 'EE&A%^5)0 3K/B)1N^IZV+L
P>MY ^2ZU"HD)_-V#P:5VA:/C6;P?S)"BF6OES"FX_ C_$W/FJEMV\@H54\?C(56\
PHZ;KU'O'"DZ;^>=+T+"<%7<<0B*X6&V:VHJR0A8#RT@D8/.U)+5!1Q81E*AQ8>0/
PC/0D3;$HZ#:"S1\[N=* 2WI0_EA54'8'D <B^EH_]=$206/?@/)0[_YB-)D"2ZKL
P6\X9B21?12GGZ!&[V%TGX<#PDLPZ&2:=?FLI8GO?:SEMEGLWY<V,8/D*GX0AE^!:
P(\]DJ:.OG\^?47+VF9>-P\32,UV)/PM?'?L&5$4W<WDP7,C171C\!+_31>DMNIA%
PC=]3Z28]3^!C\>?X2#JZ_%WI"O,V. &H-ZXN!48O]?>(RAA_1C5J;T2?^"5%1)NP
PR>?=_+)5M]J<;<#D\H7]'4701'3[U/5830W#.3-K6CK\4W$\F XWH##3(B:,R3DL
P:[;T.?GGEP!6DY:M<J8(H84;,W/EP1W1K6DP^B7XB0, F\1;V#<&Q0<YES T#-5.
P.[H/\F<[X.F#,5,NP=3I=VG0\8>(:5!%]#/^,"8BV8M#1#%6&'S*PE+D24JK(QQ3
P$UXI[%AZA@Y-\%NM$@;\;69Z3(TZ8OUIGQ4:FL>%(Y'C@PV1JP.V]2U-]HT)4L+F
P&P::S+!0NQN&5^!Y<\7-%[/"'F>I^>!H.DE_B#Z> HVSIM#(^\?G7I'::NK*6%5I
P!*:F' M'Q?L>T 3*4\M)"QI<_!%W?^<@]-0RVX$OP?ZT1-7&' H?C[>\.[<J#Z,*
P$T!W-B2\Q*A\[UB]..JE^M"H#>&I"J/!AG0+13B,W_LK3BT7?U H_UKJ<44MY\CX
P,@Z4)T1VZ;P;E& DQ=[>W%B6(9?Z0KNO!!G"ME0#B#JBWGEN8,Q[71\T5FP9 F,&
PF:0YY]F:]W5>7!DZ7_5Y82M>UR>=VO(<T1+7A-3L@8 ''0]295GTGQ4/W0ZT;,-(
P7SO2%<H<QUH$E?+U(Z2'X)&3B$!8DM+T_W$CX$%,4(D5*1B2(4WB7SB</6!'PUUO
PTLC" (IVI;$KD=1CLAA?[; F%"?/^S1E@; 0FT\I0F2VJ817$#R7"?*I(S+&S>T=
P8]"SPLY)9 3SDX>4!-#@/:*S[[0:AGIW\1IN(SUO.*3  O7RFU,G[W>@*)DB0!WE
P"T&A/N9F@Q&_JE#63<CS_"%#F^8\#:_(\2S>1^J,XMRO>&.3&KG)>SI)(_;MPD<J
P3,!N:3:5:6BCXB8ZK3Q0939TD4)LGD.C< #8A8 T6LS$#[K':WP2XH6U4YI6JB#O
P7B04D6N(3V&'2"3;9V?@MH%;%G*#Z-B?,@=V+MZSNG.Y(2I"S2GP>8*'SWSMGY$J
P4+/AM2-9M#U_I7K[@W5:;.CTDQ$5Q><P]A-<.C&4P(JM>3V.# 7( %&+B3^E 6HD
PE^3-@:WS;N'6F3D&L2/+FFO2C.H G0+FZDGK-!HHKXIS-\'L@1Y#RY[7>[";I5/%
PX4F!AD#%69I2GGS-\?]BY'6^0AAS!*TG"6-P,9+*.C&5E5JBP(SN<H,]Z]"!(K'P
PSO05Y6R!S&>WZJZ0%IXV:PC!W-(XRD'W^Y(@XK7ADT=$%H#'?(.1U4^I=L#BMB=H
PHIYR<BH7^>\*JZV+@%0$CV#2AW @ XBP59,0MA!1%;<D=J5U'S6T&3MR9)%P?_EU
P6PHYP]4*Y,FHU3IV<@S0Q/ 8@"&-%EM8*",2?H+A-*:R?R5>X.!=ADT 4I>M"NMS
PJVT?=)!L@J]:V'XO9CSS'N+>6(1YT+T>+I54HWSJ67YOF^>BY^DIFFKO640,>H*C
PJ:!&FE(Z@LAY.8E8FO?,3F+;J QLX^KZ4;#Y)UJ[8;19H+O]*;>DWEELQD'DX^$6
P#5JD?!.J'9>RI%P"YN.9^1< P5T9N1O<^U_$#7[^%2GHQ<OI7SDCR(7Y])"V@Z 3
P?# 47R4 ?R?PL*\82YFM$5 G@+3E+NOL&$E6"QZ8WXYPPJR_9"CR@N;VH4JOM"?H
P6TX49+C@@"$03"*+J[^_G5R=N$DWSJ6.VN>T#C"_2((K&135K93.U;6"B>1N+F8L
P",!2.63?Q4S+ZF4[[@0.<W98U,U8HPK)][]1S&/Q.#8!4>.0?\ _/PT'U 2PPAO,
P?WXNH)^Z0)=9C5Q>SVUN!GR28GAOQS?&(N[.!U2:#*0^!9+>1<T]:N$YT4C4:5#7
P(^VLNP!?Y2CO E*VG'=18';R)A.:'O^]J3SA$G@3L'M6CB&ZGCS\>%[Y-D9=);I'
PC\Y1("%Z][])[-\K,-HK"TP\:ZQ.>;L.#@!^K'=RZ0HYEA1OK]+8E_<FM2<_Q3+$
PR[VU8-/!O"@(-F\BR8*=V7\85-]T;;K'HVI$KNC]L*HXD^94!@S^WDBE0\,8ZQ*6
PVF2 4FV0AR7%&8W(VQRW3R5">^.OD.1NFVC2E,@'>I1KL;N-Z'4#&=IFVVMCWE7?
PT>: #[SU&IIV+8^ H188*V_-PDX_W]O(Z"EF4H=4%E*9>G$XUSV#]] IY:$N*R/L
P_4P<Z?ND_ 3W5IU$L\G!Z@D:7\!!0QWD/&W?<"I&ZAX=@;2[P/8UKQ\?.A(/4Q'(
P5L!#CG[*XK:U4Y.B$;+VHLI/]<A1JA^V196('\W>K"LS\MWJQ/!X G7ZG6G&R+YV
P Z)7*&LQ&?8U7)F@#A[LN"M&L^J-/F\U"ZC5]67,R4))S[EH\@9$XXLU;Y(44@^2
PHH2Y 45=@I?";,T,3I2_,+8DPK@E-=O6'_LC"-62S%]W685\M]"+M'-CN=.=89Q"
P]&(#A!6<9Y!VAV_7=3NHVGDY],.)^O+=$ BT,%K J)EK*.+^6(R:I L["Z@,Y7-Q
P%6*"LY6D1^6'5'KS-T)1DZ%1AV+.9-EJ^T$TU:1XE="0D#!\VK>GR!Y,6?*6W?OG
PP] #_5[$QQVL8P]+ORC%A9L/HHQAW4(H8>D4%%Z,">BJBC@H% [@,?DX ,9ZGP 3
P^ZSV_TE[3%2>\?(MC"M6I9.$:Q36.H]U/NMP_K@&@^ H6W0)Z [SA8CC+M<F%!H[
P2BF=@C!2<]30>19"@J1V6!BZUZ61D-U8)Q5A?F9LA)V$L&!@YW8A_Z6+H>0^'XO 
P+S @II!;%2#*L6&'=1O%Z'R'DIT^N:=S$P7/C"ND7#HX.9Z'*JA$/SZ5-<WN?T<M
P+5X;7_&S42O.%WPYIZK\1M,'$A,[(ULMYC2Z3]EWIJ3YT-<_#Y8K6,KSD+A=DY:^
P$*D? 40@_4G)'=L;DL\)\"@UQ3//([P ]#0KMFHICM7>DKZR'E /?4RDI<PV=LPN
P[TU!FP!9]=EP-7GW_H0(J<WVB][2& N?M<6#G\%M1ZSMJX9O+';>);"ZR7A07@Y+
P-HG_5CN$^0S9C]H^<C,TH AO!J ]H+Z-EZP2Z3:B^O_6ZZ!!8*7E_-</,:>VZ@@*
P:]=%1VPTKTN,R+V"[RXZU1!T]UXHDFZ_B;61,/21H*W3A;15&M NKVZ 06ZH*E0_
P6@<X5[?6/7CX&=O?9W!C*_L>KQ[E]R:UKB*ZS$/4Q?6UM7_@&I2KD3;QZU9EIGAB
PV3[NF@$?ZE*2CV6>O[A4P_I_'H]OJ0)K_<97Z=[$<F-T;:MMPD\+U8"=1($N?GH6
P9"+$< Y,((BO]R&N,N*$3QT L,5K9,J8%!&R()%P5G9I8Z[1[WKXQAU-#(->*T9^
P80XO-=(Y@M&@8(P9+$:[_DF==H':4[E!WEK%1[CT#YJ2U#<"7T2T=FI^MRV%8*BZ
P:M,VP2H8XRU;8E$2>+!F9-:\5 0+^,A-<L,<A 4O)$NH]4K8/Z*9_V"[+L!2%5BG
PV.[0RNMM#9F0K'@81>'CU$\:<T,EZ"%NW%<7/?%?G(@?9;+F.;6!FCZX[!3;4:*D
P$J([+A8&O;']3::ET#"/W3\8M;I<M5F56^.//Z.2MS'W A-ID^L2MM6"ERQ*8S]J
P_O?W:4P,<IW9;0"_>I3<V]^V#W)3_<$$S[2C6J_\X#+)APXN ^\Z@9JX81'Y!#U9
P&GY^%>__# X>M[1L5D1)#*DS.)^_= 9,Z:)&EAO4_B[KJ1GGG6/R9[@G8!?%-]OI
P (OU8?E6XBXE >?.^/1\K&M]9'D,#GN-;&FIGY[1_.UEF#RU=ZDLW%*B7*!3T5#"
PO'.^^<CGJ%;OT,RQ;!N#H[5'F+Y/+1[B2.%-%V8&:BQ)% CKT3OZC#E&+1L4(K5$
P)'D]C^)X$>X-90N<V*[6'/-;+^D\U'N@7VL[_ *?6LY7\G^?7"2Y4'X/.;0\].P 
P+KB^UH2J/4D0+\ >'**1F_I@A^:\M_72?31(G,8M+MQL#DB6Z"U(?K_FW2'>GIL@
P344AB[")K:M*ADV<$I@O?SJ.-W5>,;$0Y@".(6O?IF7PB2[</\$C8I((3Q=[_4\=
PY,R/5T[&.?FON"T^NWF,;0N%AT3(L;^1O.8]@>&\CVTWE:CGRJ*DYVCH"CP=SF"M
P9B4!D*W)GM(/XHW+.B]:T.CES(EX5'@BT%...U;*+BCTV%S?*5+(A3)0'H8*PON,
P>;*X!H/2M 1@G_2E<IM0QEAG-EWS;S5@NM_\?&!QW?EQ]QUW/=Z'W"_O-PI_SC1Q
P[%(D")6BTF<1YT(T_"EV*VV7PG$*\#H8#CKU)2?SO69Z92\/8?'@I\1\F&5+%#<5
PD,(<0W*$&<*B/2+'CB6NKBE4@QL3(J;Y:$.JEPZ]^+#+IF]6&A+R49$N>;Z7L]=2
P$N97XP'J](%4S%885)$%+KIM'GERZ:^N&4K/$]50^SK_H]$9 S]LVO&7^)BJ,\"$
PU] 2EQT.4FWUEWA)"HQ@D;5R*J\5X=<4P#@'S>4*]AVORZCI1%&NP8Q%]GHWZI?.
PT(8$0:9!]^R/I?9*)Y Z/J"T\^U;8L-G\6)^O -I";0J <![M1K=",/"Q_(#9TOK
P?.B"&D[?(E.O"L'&"3*Q>^<",HR:#L BH;87)+F:)%@*?G*<-9")"LXFDKPLNTH0
PHF?355BE,BIITY7IF&IE!R)TLS!D"2?61N]5L'Y]5B2\NR<8<J$*]H]%:4](''^X
P'8IVO=M2Z@G@-$/&SP3S8&XZ#0Z;$,/8*F.,,O;,U)B[A@^,3BJ]@)YYB,A<!LDE
PK2T-X!YK "S9(W_$@&@)5P^AJY(^JQ;/CLK$FTE9VV=$A9XOC;@>3K1./S35RU/O
P!]Y+;DJ1^<D-ZBI,\G:.*_S@?8!'1^_/*3T_Q&X/CLL4ECU!'\V'P@\$37\.'^>9
PEXJYYK"]-H]Q$X:$ZCIC;XM+7/YD9>LV1<ZT9A\GJKBT XUM:=!L^IQTHPXP%P+9
PNO(40!OF9%RUSL836D5]$2A,LD"3Y!=GT]EHN3NGESK2T(?;[U+$G$%\CHUFU# >
PXA9BXOF:'J7%XC,A"+TA%SM.H[@^)<>\0A).\8NTMU%]DJ9X>5<X1 77+9-JKP)N
P5Q5WI0C&S,JC&OLQ);0W+Y0)T31O%VN<#CGD$9*"C';ZI_X\FG@C Y)]D8R90@D9
PP<51$G#;,;C2I]'\K$C!1K_ED?7*,&(=K3]19L]I=%>SN=DPD>_UQ<6Q9?B-!G=K
P>POT$(&94T<*I)MQ#1A0PN @;(>X8=&;W8UJ\IXMMWL^&C>78"+JX:BJ[$[BL<40
P>HNY-+TS@H5")?S])#E0&L'#3_*YZ[A!<.?!ZTE[&! '_"H2DD&X9C]4H+-HH$;]
PO\PT,YL,,6[U7IDF */C\\(0MM?3'A<PAA"A$#&,1Q9-,$&.S!I0:\FU36!WMC6A
P4KFY]P$5.E3WE%F!94DR7XPTW)A+. _E]?"V]7L:/HW87"NQC"Q]P[-05^%YH*O=
P9S+$QQ6Q*[-(-6D8HZ<#R#PAXVJ2RFFA%J11CC96/O0JS1)<'!"B^Z0*?<NK!^M7
P2<^A-A?_>1E1^Y!-OXXPX8WP*+.?]H&X0S^%+]W-K2<<OER O:T#9_Q(EQA(?VH 
P8?<*'V9)CMAA<<"[@2;C^JJ[K.T/,&L"\XD3[^L$(.MZI^3RD:+,76YMZ!B>;@)"
P4\'U+Y+W:E5#=%A[U+GX\[4+'&MSOE=K0 QG$P>_4\_?E80_J&'COZ)HY1VKY)OK
PS?=\6!1ML(MS-GPV>;>&EM)WX:$N(* S5A[DX%-0VS3LO.6VM)$F/:":O$[$(:+!
PJ%C7RSS=O]-F-[QI'SJ?T.4Y/N,_**$?).WSKR-D;CT,D]SKKUMJ=WB.("W:G%"6
P'A)Q?"\8IVA".KA$"?M[=7XU(UB4DH72NW >IDP6$T<<!ER#%>7W^"GQ%)VBGIBG
P]>ERZL-5]NVSJK8PRL+O.9*^=3VTE)D*.R"JS'(@I*0Q==#"KMP64XK0?6.5Y:HS
P8"!%O=]P.HAE+$-G,#UD;+=I;Q6'<@O%I<EPMN3]U&DP68.\_V3YV#1;SZY,?@>W
PB[^OL #./RK%M2T*T1QV3#N\#-RY EVO>GU 8J(<8^,N"(0+$V(B<VX,C[)Q.@H6
PN[X)"ZK6+H34@"I(RY/P#P1I-\)',<FNAE Q:UN,_'B)0QW223NBQW_NKQ8_IXVV
P_2.["$K#N3%7HY74NJUW[]X@+BJ+G"<&5_B#DF0"#Y">9\2N9<JPY[E26]F<W9ZD
P$B^=^*UEE+C$.X1LQK\M0H^]F-7PX))257P-?_4YH8$+(=,V2ADFP1:Z:<'W#RX$
P;P2)_BQY"3\E8_%^:=N#.-7T(?!Q%G]B]P@PP_ZR=<Q8GLMQN\QNQ)ME_IYA1%=^
PWZ/WE*99ALV)/QJ/_MG_SE6Y&=!"XN8O_;W\:]T!KY=\+*L@98S7A(>OA!A&/081
PS<RH4%6F_ZR2'" IV!K7R$K?6IZ;']I!=D8,/HTM2["^G\?=4":[7XR?MON80TY[
PH_2%815-ZPYKG B#ER@;E8+H(4]S*$FTQO\_>*1V'FP-"_,CO!(8]O=80PM<7S(J
PR*?/X_CY"NO31,*PH(A^D$UE^&Q;IDZ/TDS)F4ML):XQ$E9\$! EX^=UX'TX(RG)
PN)1BN0>K4Y)T.Q;9W459L /[K]/XQL]*VH^R&AI+L"GY_,Q6K2(F$7D._K?POC4G
PAD:K\#*-WL8JI,PI"Y\9 :H4AU(*/R3=GS?Y09L7I8#O>$K7&/T_C%OSQ7,.)+6S
P$OGR5(E5J/2Z[#656+I^"_N+#Z;I&QZFRX258,YVK')H9 W?D-@B[#TASYQ-2NV0
PYRX#UL5)V_2I#XA@>-L<<)P*?'\(SGE?33?S@)A2(*;Z><W/*7"C!'(HO+,DU^E*
P+M6$'K/E^\U=G0D1#T/;E[(=L!//W4+1 $FM.F>&\9 ,O>$HJ4@K?@JII6Y[N 5.
P/%G$)G$CX/K_D"9P)/5,*/X4:B\,AX8S([018,CA7.PB&8]GTT6<WW-YX]\?9X&6
PA9@Y3V+/O"PV;:DJ,1?]_>VTE7RJ^M5G,EL'E4B?A5='K<NAZ#*#5ESO'W0@3CIG
P2BVUGJG:-,&Q_5B9YKZ8;CX)%A':*!5P<0LHC'?N ITROHZ/-$I/PS'TJS_'H,E;
PN7>D2G8*QT@P08_$P\J[^RDF:H(A8RVP@O_++VLB3<JUW@=>678UVPS1D$KTI9N^
P8;DZZU(/'X-+JC_WUB.%8,%#0HJD]6#Z*SDS!8FWA#GBT!(=08R2U'<5U\YD<#!C
PP%$58&4TP+ J;3DP 3 PK@@O6C[(@87MSDG&V[4>36F@P+9KH/[$[B$:;LA=IO9B
P#ONV[^7&QA.L)1^8!E5<\T]:LX46/@'T*VNQ;W5N/L6X85-^W(9/!?+\294<]UP$
PD#\&PWF>KCB#5C3UDKE85/4L(<$KBN<(PX)J BI>L3X,^WY/LTNAD!/=T!38=9]6
PP[N1D]).I<ZX/T%9#U6C<.GLB*(O0=KYV_G^D)^F8!W]Z><G#"(PC[CV)<:*O-D;
P5#!2]O"1^HW\4SR)4]S ?Y4),P"INV5(MA_/">D"VO?,K5FT=5VY7L5+TC1_OJOL
PE.I%3 U=M(B.ORM!/9]=M*$_G/3Z+1_[T",8=#N+@ <!B6'+JRRB7'TM/9V$1!U@
P'^[92D-.$_5@N$$/FT'\Q%EA[TW8YB>G6 RJ5_FC7@]* =6K)K";G?;'LSAPF-N.
P'HD;C#58BP&7&7QQZR:IIB@K?B@['RD0;L\Y^H'M,,$R$83)TM*&";1 GH=DO(['
P=;X7+9'/EX?6]J7-$EWV#0H"W$2T7>S@+LL;>%_4+!<BX:0L>+1.HBF[P,6<%O8%
PK/_D' O73>;%GY1 &U379VR\SE5N/S,SC3'&M_MG/]?-VD%O0[ZR1/!SOVM<_=U[
PC^1M_[/2+$KTF0>M\@[B9Q$="V$U_OP-%+6IAS+9])?1(I\ML_K@AM8)@Y/PU M 
P@ O$86/%/.%GU$Q,<\@E!<G9 48)20EZJL<UQ-HDQRE.:+XX]EGR1#Y:AX"<F A 
PT=7=NRIP<3;SK'0<4NQ*,;D<8C=%AXC/-W6+W1Q\Y&2\C:Q#4]SHM4MW*]([K<J4
PDRKXF:'AICB,7?X<<[X4?'DJ>AJ\N0=P7>UR64G:)X>GP,PRS7KIBXWNKX.X>DZ!
PAKU[R5E:CJ50P<S4"&Z. <3.HE0+9+(I6!:8<:L&ZBELG9VU@S&,-4?9'78Y%ON8
P)4434P$37A'_GR6YO=_2 ;2LK8;AM>N%R73^SO$B^-]/2$CIY.+O['<-%DK-!0.?
PY14GW)?XM1F1"GT" 6Y0.PK4'#DT^06.,X;&9YC'M*O.T;D.'/ ?KI+VVFJU:RF]
PV>BOZA\B[&ZF;EH47B1OU"C=U;/RS+B_]GZ"JMI%,C7Z>(G_^ ($1[E:=+<HP2(6
P?[H'CE]E$Q*2Q$_"FF&TK+\*0.A"..T;:W.S 6Q.JD]7VUOPY1N&00^N*C L)ZJR
P<N VX)/>0'XF]0K-1JH&[J4<O6GFF+E=C3%EW+&@1*DWKW()M?'1TY/.Z405=ULL
PJ#;B>@EA^YN@\CGG#(*@8]PX<6.!/O(&+JZ*R% <,F&BU7))05I)NOT\PCUE8=SV
P=U*:I(4-0%N;52(#S!.N2E@Q;33Z'8I:QN8%9_N"B0FG<_:5AFU)=SAK-BDXD"AW
P7JL/:+L[IDZ:+02:[L]XT9VGG3]=1-*_ZPZ=X1 69*^6W=(&0 .>LS?**_!Y[<^@
PB^N_;S=H>F1:S-8ON?2>YG5NZ&K'*J.18^VZ#ZL45UJFGI'GFLK1P>RZ;EJ-'>JD
PV$B22VY@43UJ>^W#46: UL8:<BBE/$)1?*R@=[T4_R&.E$<7N#;7: ? J1".\LJC
P5::G/W58=<YW/H?03XZ]52R(RR284U0^%,[_5(%1@VJ:R0(I0]4HR&#CJN5%O<@"
P1X'[66<<1@D4=R$[K^Z$.QZK!97C&TB"DI[W!?)7[UT;OQ^E/CR/N2:_3N?)UR+%
P'(.VZ1>_W*P]9\RS=K=Q/ &>UO0@FO./+<A?'2"/Y]ZE7.UHV"Y60),YQKK \(79
PL]%KH[@>CHUZ[7;6 &X\>[.-QU_2>0UOTS6OX*X"QURW7=SXDB,0#RC!!MP3_/IX
P*D*N<XVC I)L4-H;N_G.'0@D/TJP<V ==H6\]$9:E _Z8BU*YWWZZ&+T3A/Q(6L8
PT4D;OIXQUI'-((]U4SQ*;:N@!H!:;2*7+2CLTX=Y-KF:YLQRK;G[9Q]AR[IO6J1!
P!>-6RYDQX-&*673A.A79AU-N5HZ%VA$8G@S]]*M]"<SCC*,OVLO7*S@ZT\'-!C(Y
PLCP8US$BP#I-KPI4R.D=PJWW#T018@D(&CPS)N-Z[M[VA##.."[:I&=&:GGKK)K.
PJ]3%]G*H3+.]PDFXHLY"*V95W#GY1IY@.W%I75PW46>W& & <XNI A2B0XX;1)E1
P^B1B@KD69/FT4"7W+5A#*(X2&(-+QH(N Y%)0K$L:J'2[72O-OB:ZQ';_W!A>3*H
P?S4,$,P0R;$:#NFIRXYDP/VJ&7(+&GN<#;#PT4"! MF%A'K?X2:C^&(OA[I:<Q*P
P6/BA#Q$XI]62*E*PEK"3]$.=-,AJX@R''VZ=(61D+BCJ:5+7+AI)L1]0S.CW A#B
P-\]0T"4R*2@BY-)*%T&4M78JJR&)34A6,-GC;V :;VO;:Q0 X:.CK 1W;R1 3_.G
P/+Z4/F+,,*) ]^J?!M:!3XT>>5(4,U3'0R,[&E:Y&*,%-/@WEC3>BYX*P8@Z-;*S
P+@5@&2Q>_)O_B3/PE=E*>_D5JG%(RDW)X]9KJ I7-X&)^ZR4VX0QYOC]]9J3R!P!
PV6-E@MFG9B>W$/%.W9.N>JMM=.7]14[DA9V]05LOCU-T%&08'_P\V=?$YGZ5#MUK
P\,D[N8W")8X19J%8!+1WT^C80]:,(&)A=WTCT062U#=@7+AO(O@M'>$:I/O29:?]
P^H8Z#,?/.,EQFV%@U(_2#O7VX$D;NWK7E$F&09SMK]+E/N,O/1AZ/BVFS"'E3)OL
P/0RFJOI2O4O[GY!G9O:QB7KJ(2R/;HY_REL6?+GV / \*Z=(5?PO<0E3&@/@E"%T
P0=*XKWI/NL0\_$7\B0EW3G"<)?8+"=@>7>O]G*\VJTH3#ZI8^9O"2DAQ(SF?SC]B
P+!3.@2%[\V5+;9]&'B730((.KJKAB&_<#$P:^%!CW.!>#3&>&&+N^^LQJO&U=7OL
PG8CEKAM'D!$#=Z%$+9H&%2PEC_(C]@4</5-\J>@W)DCFU3KT=__0C!6/!CM%P5DN
PH7N:X#ONN$=XD]:W[ B'_A5=]AXA3%-C7-!_IIFR>!B8DIFG4/V/-CB)D,)V?<DT
PO';:WP++HX)?,<5-*UEJ:UZR"\BAZW2O(=U52%HCNDD'TA\!?($4WG*QP[B^#+ZC
PQMEPSB6A+G?'W@FEXF [>7E.6X7*D=DX&&X4AH5)J76=/LOE:(#!@'=#*)5=1K9R
PJJ2QIU36V?PF(TCWNT 4=;Y%BHBYCT)##DV,-D80DP'I[SG#(#>6F\VAJ8<A[(KD
P<K*T^FZ/(G\QPS::NZ1)!=B1Q6XV6_6>+"75/0Z0 C&_>5_;"6"9P28J\#+Z(0>$
P@(!..!)=YW[SEV(L"A5E%]X)N#:4$,A%F=G,KEF[@+K^59EZ:5#"MW;DJ92IEN^Q
PK8&H/LF.WP#7)4$303UZ 4W.4K]3.$,'UEE"660DO75#9'?HE[?N-81I(MI9_/&W
PL/LQ)CSW"EW%*^ ;QW]:2(=V+K4Y5 JX1%V:8SJR\ZHYJQR)-$NU55:.T,"'*7YT
PX-PI1>N+<"^I82MAXRYYS1R:?F;2? >*]3 &G?[AWSW2JQ:=,D)13B!WU#:!Y2OY
P.V,:WQWBW9#0=F,"#TZ-6T+[XJ9,5B5N[LB" :Q.+Y$HGEIIT\VC*>;]>+3K9YO+
PL@2NY8%8.JX)-U3.E?_=C;B3LOV[S2GA%8"(]:DU9,WI:TE,CJX&D3L="K>>3;P"
P?K6.V:+!X1VOS),45\H<G"+M826O_5 6:Q?E1[V8+>T+]8M*&-KH937[1*(MX.J]
PZ!3-RLOESR=C,J40&4TWDM+S<:<RCL4MCRWK9IVVS:,MB$^$+!='@"]YO:BC!UB3
P/Z!4)Y$+.-CFXQZ+;FA&Y];5[A+IGZKQ,)SN^#2\1*5,#*.(@O#4 >@A[4X>(%IJ
P(\].23QN$=,8LPT7(?E&?PPL&9.F:")&AN27R"E8"92W?Y9XH 0O/2.BVW18OJWD
P4@Z9D5@LZ2#Z*#/SK'RNTWN'+_*KU +IE#>>B+,Q*4I\^Y/8!_,C[ 9AAA<(WIQB
P]8$AFMWX\*]NXC1C> 8RO4Q3CW>@Y18&2T]YMT:-J'L4PF4S_L,U*(&L,9"?-,<Y
P!H /*LR7T'C*MBM>]?M7W1GTW=<\3D<%(5GI-\\ZN>YQ8.309A'5S%"R*44K6.IY
PLJ-VF6[N].Y$_A%P4,X_5V*7E(*GL^G;@ULAF(.-R_M>'?9M](WTL2W(]:H_XE&A
P%GASE^J9_X&E6L%^"J,.%0F^/]5CK"UC:HX<@U/^13(%F!=S5\$S^EA,:8<4S=2T
P&;\N,"ZPNH@0@J:-9 I-.G>?,9PD3!\4;'#%6Z\AKM:28&%!]/!4TMS75JDP%7#^
P)Q,RW;WM!W(]>_7\<NV.X;)L954L\@[[WOYJ"".N&GBJE9;)4_[=]A/M;)H%1;P6
P"=OOY=__".90+%%J+/^SH]S2 %\U$4-ZG@\F4:[ @=JFLT2U,9"6-AA&FA9O-5=3
PA39K _MN8(H63$8ABIV65.M+D9SF(#0!19XASYL7+>JIM 2D4[4\:1U<6Y%@<H,C
P?3W9@^GIT-H^U;-:Q:,W[H>,%\1"?O/\A\]-,4?@ HK2]@+LEVRL[VTH&-"&66\=
P%5[NT7B#Y<FQ0II[L!W[,'N+7[<3^-FN.-,%SV'_'6"T@V(X>E).8[1Y]&&DLWC"
PUG'<3?N!3PF"C)9F]T^(G@HVSO;WDJH4GF0P<.\'#B_  67RT .1 /)I].];IP\B
PV7T*W]XJ<47X".]F\(7MP6W7*+;HGD?&<7CH*IXD5(3LL2214S4]8RP.7NZ.^+/=
PYB3USR@:K%:(3EHR)S**O@NLYQ8F%O7 QR89WO0"]&-<."=&#M/E":39%[N(A&'/
P!H?'G.IFPK89BN1DX1KY,6X\(MA18"PTMYDL:@7,HR4FN%+,; ICI0;:K<S*F:* 
P6^<":@0N!: )DQXK^#]A(,5#['$CMRHK E8H]2,.<YT)^N%)##>O@(HI'\<Y*3W5
P;6/CFM2BZYVUYQ'OS]@!LR]O7ZJ7X4A)TE'N]0WNOM"8<8 K6*]0 *J%K+* IFK 
P][L*'!:JI$=X\?%U$K&+:L8-1'[?!/_1LYB%WX$,]K..+U<""%<)/ZG-4T-=VBMH
PYLM^[H/S-5_\GU8X^)2U4%7VIA7GPF:$%[_=R O!WQ?>L+1*EO&/GX]F3-_]$3XM
P+OENHE)#_1$B:><Q7;YQGO]ZGYEO8!:TROK^5(TDDB#1AUG3&3'\@->"R0>(P1CA
PY<%[.O$),Q[Y@.\+,"<V5SRD$ #4>\@BER?<"R;:2NSDKV>W5N*+'K]I0TY8'1;6
P'!KQ;O,7,NS_1FG%1U>MWYY0AGQNU29C%6C95VP W-@0(63CQ<+EU[%[LSE\EM4)
PB$FS*F%^];6./.J<4E10(@$B+L]]&6P.Y7WV6A!EW><",%(TLITKHM_+F!PTD.]&
P",\L8.GT\QD#%2::U6K<W;*4M4-5/DM4(,?C3G>6-_N)VQ<B.3 P"A)8G3&C?!5J
P\66&@8;&0FKDVC 1IA?9^(%KPKZ;@!:'UC>-Y_S& =&?Q75!5.M^?CC^2'>S2:J^
P89DNA9>W:^.F#0P-FD_;E@H$_.?06P7-*AD*8XTN2+F68R]^0B,3D^+,PK=1W?Z/
P_8U&/&/L=J!APLTE.H;F<Y.N(=W8<MKUQYG9/%?!GZ)I.]$*[R'D'/M7@&#VO>XY
P&MDQ*!F^Y7U&QB:)OI#&#>M#^)-\_.-7.;&;K\ [V,BS\8('DS%M05K%84SB*>RX
PL(] BOCP%^*-24#$(W<BNL.LY'[!1O#3HZ9693CAMR9*]]CNT>Z:N@U"9)B,3 C_
P=XNR?>:D*Q\5=KCLR6<X-H2A)E)DCO7<5AN]6O@8>KY&'F%>CPJ,QVL/.H=>]UO&
PWT01.^TQG/(<)DHK]9WC!5$VV]DK:$WSWXLZZ,QL,A/):2K=9UW9<0Z9C>3*DK'X
P)]A7E:G-TFB%SOYLKC@[K:BV,HIK)501[M%O['BPP99ZA:^TEZ8/Q[K?1,XI*GM7
PZOB(K9X%K.4_MGL<->]4RG);!2USDWZS@=#72@V9./&TA;:.<$H,UOVV-K?TM<)Z
P)'U/R?#FCOKB2UZ3H-9N>Z,=:7Y?5!Y8IR)A*:;;V:Z 9RN#?VH$'SY[@\)PA(PS
P:GH;\].Y#4O$[H6T 4.("HW/T )'CT2&84:UWJT)+H2+5FK?3B\GYOSR$_&]YOC*
P#J'-1CN;^P'3=C7(S;\8= GO%).-XUCQ4%2:)U4"-,/#P]H?#PZXP;[""S]Q"(UY
P+79^_6AFTL#K!K^Z>,2(;EV3%JI6S4JLRH6V:#:I7@.(M.K.(6H_G87(6 #R-"@K
PRJ&,W38=<RYHU:;(EN@6$K#5A"+TM#GD,9^ZEDL= 3_\2UKR<E>S+FR665=!YI=E
PA9./^OOR#0-2?3G\HE.'!@(6#P:Z3#"F\XD\HTQ40$$V#KA<AME(15N^\/L_&1<E
P\GA.KT/736Y*L:^ 5[8Y3/FCF0"K[@PK9??XYZ '*-TZL@A9"XK[W5T#,AB99<YS
P$TG;__IWP&]%K77)UVC%MNQ0[&>GX]J+&5C3V<_.-,\T1TOO\CZ11UM\BEPCW!N\
PCGG1B]L#'Z9O[D%?>,DFEWH5PS>FPKQP9O=>5C1["Y9O&L3K9JEOK.K$H/A!3F;R
P$UKH8JJ.<JG5;K*\+PD$L#9BD%>VS'J7,8G3B>4P)M*A)O RWW#:VH;$BZ3G</U/
PP>^1"-QU52(W(6K3@]:$.=9>C4*YM(QP4\O"IG7S/$8)13@-9#'8,"4V)4FFH*\S
P@V-ZS7BR&UX^^O'BI.ORUZ]HZ'^_$*?/K-(L):(40@TQB,YL3Y1JY+DB"JT+_ /Z
P@X4.QJ^ SU480PKBQ'#O42$7WMR>]!4Y,LCGL.[X1SC)VT#L'!CK/FU?'N;UG-_@
PJ2;3_[8?TB0Q9_IQ>)V[RV:C"YJ;A;4F/!#'OAL8*:[Z=GAK'/Y1W@A5@R;[7*.O
PGO)<! @)CCOZ10JV/=$6W<2@8TOU=G+%R:A#,OHE=%91J1E7WV^VA[2^JT1.B'%-
P+HO\?N_*ZGJ:+,?:.WL747,-DN5-/6SQ,N1-JG;0C<Z@:2YA18Y3B/<#4K3<PP*8
P(@KERRJI%S*J@\#>XP/.CY@6/\=.9A/$YG*T_YAB\<@%Z4L >5*W/OI%9IB_?%G+
PYV@."FTEF4B:PD*!!;A GF1%6-0]+AK-INHZ(PC\E8H;#XZC<1M43NDY-MI=0:00
P? ;4ZQ*ME%&]U;KS<CH!;UR4]RCK;"Q>U<87\T_&L@#*0L%JV!%2^H0NB9GT-8#R
PI,_ WS/#6>TZA$Z;UF',=NP-56/, T4L^-8NXA[(AM^\A9UHSJ['K]L2% D%/*'\
PO/B&&&PR"5+[T9YGE!$#\?25'(CA.^;8+_/:U4JB7I.8=":H1L(E6-.^P\58!;T(
P5@0E# /1-4)E$\V=K@JF\/>#FV@WI"MK 7[<-O-Z;RB5\E-^?V]C(\@4KXF,S]9?
PB6U&'5:2<1$;C$Q[UN3XR"C'8+?NN8"(4XL4/C1L-->6I1K:(:DH:NSOQVNM##Y#
PZ64$Z?Z@D?H/VR-([%9G3GK)\G2N^/RA'95IS,_G%NA?-]LP+'B*RIKA.IY:L4RW
PM6KTLG;>M3>]\WBLS!P6)+2XDI&J8XTR \;[;*O.B]3=ATUO;U4>ZIAMU-E1T#:E
PMHQNB.6&\T[3B<365/%5DB@6^B[Q@>DMC\7MX69]<T!6H(3Q&I&XMY-'4ARI-^XK
P@XUIR..Y<%I/XPR"'9$&A[N)?8PG[G0&0OT/Y'U0%A:MK;37LRBF1LTW*X]T:H64
P\(>"HRK2,(79")K'#AK%BV@TY7\W*%N*9<M>9=_:O()*?;3Q-/J^HI-BV8G%-#PD
P79G/E'\3LUQ#]OJF"L [<0RKLNMI#H03:"XMK*^7WN]VZ9C*!CE_!^1 JH=K#/BI
P\=Q7('B%#-C0FAP?[2,'M;:C >O\%Z@,"-JB6;8-3C"\Z;UM^ E/8-<FT!Q*78A&
PV.T/H!9X^(DUX5(MP8BY(C!4.2?Z1!6D",+D;>=@ 59,(KR_00%#8?BJ)47)?\3-
P@-A(.S)OA1A+$!*F.GN-Q/JVL[U9'>L>^@LA_=DBD^_)'%P6"\!;K\V"('MLA_PV
P^UK>_37N9\9<IBM7;B*R%U':;1P%PQJ;MF8&J(. =@X67(B]<(^#FK/Z@OGE4S]#
P::4$5!O+PZV.JS]K]E-F*YP^ON2GX5+VG/@ 3I\%A%NN.B+-T6(^^B)BDK\T>JUU
PS*Q"L1<<[H'_;$NXZLO2+>XOM3*!"/P3Z(1"S2O?UXU-,,DGO]D14B!5>D1?3]+^
P?GCW,W^LD.F_2AI0HCX[Y$?AOA8P93@0UTC[S=1X8)@.^;<:VE:Q-LD';I]GFT\#
PN;B<3_[Z8ASU^XB3(RJ)']6IWK$O\_LN>I*@:O4-_DFVJXP"J_]"@,1Y1<%HUULE
P$RW8FY)1%B&([97E9T-<J!?X*[1GWZX6J6?ETEIYY+XW2"$KYS(<X7H!/V?V-2!M
P[\][)[P N;US:'H1\[K^=M%#UJ:V)*T7.6:K9D1B,>\*8D5"[+JJB8L,*$Q:O1",
P^7>6M&2IHIR%G%-.0?M)I=H!7OVTK 5?PD\+"M]5K'1E0HVW<H"<8]&M6#0/0!X^
PS4;H9S%W-BZ"<RX+5F/AKX3ZA3Q?A"+F)^7+[IDF/Y503/-*KN)5#[:7HP.8+$8?
P<KM.:GN]G24+RS+((-^ZG 25  II?C*1*OYX0KYY9MT=6O[Y;1%03O$2;E"A!RL[
P^,3WJ8/FJ3Z<Y4Z>+6I6XV@9O##?]0NHV\H-C,D03OW;AV>YZLVK;M3?6]//# MX
PEB-Y(MHRUNI'5R !&R8/,Q<*-GQPM#K&)/%#8T0/BI_Y5&YU1E;&C2!5VL=%"%[]
P4T=_K/I"+"OMK*F7I]I!2Y%*FT6^7@#.FK80Z81"!U=KLFJY$SH3P#@DRS%SX*1_
P/ &L-,'QA-G5USE,@/U,<[GQ:W/(4$*!;>_IQ5[O>WS0K-C+6<)PIHX-$;T@8[T2
PD:C*QZ?=-ESW<3U3$_A$K4 '; 859'@]A-K3S0&<]8O"M.J$'(P?Y%$#E_V1=@(S
P3!OB#A3UCW H#X[!(U8T+G^ZL]35[/8M/IJI*U6*#P!HIS-Z7*<.X\(5?![9A@*K
PLDV+J;(]J)V11'D5D%.>Q?X2]Z>]3];#?N\TJS9F$QT:3.Z)%3'2P$'51&#8SRIL
PPJZ2U N,YZORVL1*3K[&OX(]29I*=W766^DC9COJ8=,A<!?U.>=2YY\E[&<K1I\&
PS<K?Y7(R.$_NR?^$ZAK<?CYTVQ-MQNR!'-WU\XS> VT99^F._"[ALE7(C>0F'V7M
PQG)- Y$<-S@KV-8B&60[\D]+)X^ZH)$AMSP^R?=J)PZQRB36Y*/.G!K]1:S^ 6[2
P/$163Z%IB)4AJ^KM30=;ZHM7\$-,7F)JA3)MQ)F]';5STABH5G$5AP!R>E,#7,TM
P[#&G*YTG?$6I9$&BD6E&LZ,I3)./M"GH/-=40-93(>?;JR*G=D*]F!+[G[TUE5B$
P9*!9^6^2/V@!YW\7+@E1N6K:G)E92!B[U[PAZS\!2Y[AIMDW\><H/[WM=730/9*+
PI.0J5"/9HA^[V?@.*UM6@(87KBOSJL4,0[I7,,EYBS1Z3>UM@$0=4B**>H!8FF%B
PMRBAC67=%EP8\^IUQFV3Y*ZH+2YUCRY4F.N?2&S'9DD.)!O+. UJLN$3G:2E&BU&
P(GWY]*YI<RWMD43U=2_ETK[K]>.'H)T'(EOS W^?=H&44%)X;KL8TC(]/JR#!28"
P]G(^\"R3+AH%Q$<:E"7U$"CSR!QGD32P>SH&*9\#Z%^<VK72S^91X7#6MXVN!%<8
P?(JW@Y9H718!Q<JL*U'(T-#V,_'0MMG,^%Z\!'*.&Y,\DE_<Y6(#R-B>P#YXSI()
P\1P^O#F"0]#J.YNT: \@H2\=NB*WR6M6BY#DCLO=QJG+GW;HB+),@QCW/6VX2:M/
P%I^UA']90,!HB&K*/K0.SIW-8E.[&VZ@M,5D=MM;YN&[!))^)DK*\:NSUH59W2W9
PA+>[RKCW_2M60H+$O(^I%<IS7FB\58:ZZOO2Q@]/(D5ZY]SC&1FOANU]-8L"$L>S
PO06E\.BTV1B-RE?X/3[UGO8A>A7$[-T@5&PX6-A"^0__I>R8I7]QOTKD:Q!'0EPA
PC)#%1M9=34K QH/ZQ-B@%NLGJ$A"'DC/+_.$A^BW>ZQ3KF!H![JP\FWW2BU&H"[6
P?.TZ#_W,J3Z^BB@:<XYD$UZU@)>JWX%/.5P@;Q6*QJ)V4?HE]ZQ>-]B!E??O#O\9
P=Z@_=RER$Y9^5(T3VZ0?RU@-JREC%O4_[X?2NW:9YE4-[.EBW[\=6,(/'K:2ZIJ(
P:/.AAFLF*T]87)\$9.C3Z\=O-\T,\_\/@O%+828V:KJ4=9M.N7]:*; :3P^H$WXS
PMA(QRLR]1/Y)OQ+:OT)A'VR^J8O"(Z4[ 4D/8;-QHW<Q[2G.<TV#>HATJ%3M-F&C
PELH.IIWUD;:R0L#/FRZKRAC%QX"I#$+KL,5]2ZWG1#H[JGT .-K.F='5PWU)4;?(
P,_9#?"D82J@M<N#^E_5^Z&J]PI:*M>VB6((Y\BJP3S2@0=S"Q?B=1H:I>:FEDP\3
P^WX)S0L+45W(2V_%NBJQ_NB0;PV\T&C3ZLM5'Q6N"@&)U=I'D,;#H B8_8-I;P77
POWV<0 E.M-UUH<TVK126"E$M8]&AV:&NDVS@4S$.0T3/&^M&3T\05^M&6;HI@ ,4
P;E_PC7?XQY'R 1!)F8,"N:S>B09V_8"!/T 4)L!)E 9,[!T+'W2ZFI@UX$-5!4HB
P;5G?K0/(A1<02& ( @:O%:Q]A<ME_'\Y=(D<"'!6F+OC ;,^FB/(L/GD[0YG:LSF
PA>1I[]\E 10)]>16YGDUVVIC5PHRJ0^BYR[2Q?&W,8&];[.]!!CNC^-LI?[;9T.^
P?J=$[44 &8E4\1QXHP>(X%T2 5N^,A-Q<>U[30#-"A"XWO8FSD!D*#H.Y0.@NU#G
P!R"!.6]</<()3_7$G/#R5(L<]A]WR1&OBM?LY:#NX^>8^S65K,C?=C?,8N3J[EN!
P\?NBBKP6=!8M#-Z>2,C*C'K"R^RM]H O98@LG!TD6/!U%:Y?#EAB8NGT,IB!KY,)
P(UH+O*W@R?34O9I)-C^@H)#=3(LJV\'CB1'"_<%AJ-KGW,P2CJ'+%H3MEY4<.B2\
P6UW:VS(&KK)L,"CE\<,;QEI-@[SHLBGZ&__VM*!WSR%S%G[.OUX-<K>)MDF#)H-B
P&B,5L_9/H0Y@OTWIF8NM@CM+?Z8";@T'NWT)]ZAP;R.P'+N)5;K7U:D6GRRL^&W&
PX9>V"L= @"<.N3W6M3X !C9EZ[\?"LL1HF<"Y;X8P,5>.-YFI@)SV]#15-JDS$$K
P9VF@6QY^=1C>[&H?U/T-:6>R&09)I=:,1['S)DX);>6!?\#0,:4?@U&OA3'G^!LS
P81>RC_:T0L.!3;LRG>W]1QO1P!RD,0=#[\W__D."\/J\I;A4#1=^04T2.W#.[O!G
P*98Q'K]OR85;2B)=J9TN:!<-9Z"\R/3[I4'$ZYR9G[T\<_J]5?(-G@6>9#6:GNAG
P,N%]S=&Y,B(@#XHO%9@6V1@?B3_V6DL1@V2$J:Z_'F[X62OM@Y!ENVV7K=$6GD*X
P]=DO&1DUS-K\4HU(MWI.WR#.I(W%'V[:" (@1A_&Z@_H<1^G(N[J[Z,:@4B!2<E0
P,F6;]CUREMQ?C@%B2^F0%:FZ\)NJEZ(# D*G_2+44QEUG1:(IG^#/=)F["%I?B? 
PO'<M(P[^ZOHEA :(NF&NM]!G5-T=GSOIN<XBP:_MWC_N?5H+F>_PT$K?+WU=L9$G
P<^)_X$T<W*!!,S&,QZV0_\M3!U.90Q;$NXJR6.%^LBO))H7/ZJX6+IQ/ABM9\3X/
P$+&+8D9)N=J']F%N&2]7.@7YZ:()%$BG,6-7DT@B7 YGX*%YGBGPE,/YXF=]NP$ 
P^ZSY_L<K]J[&EOHSHR*=9=)&V(>\!NO4R<JD>\46LS@/Q-[M*22>?[OP,CF)) 0P
PTF0)SP*I"9($B+#<.[JQ/O-%+'SLWLJJH\0 ZO3<EATZ2LSJQ8 BI^N:"3^X@0EL
P%J=B+$J#)]4I'-Y^BUZL\I+*GD9Q@![X5"]#&O'*3OG8)T.*P:P\1TW1M(3<=T <
P#S+GVX!I#T=1]GBY]M:+1K"!.\DLZ,H(':[=P_86OZ=^GGVM #' \-TPYD!!C9N<
PQ1!G:+A>$QME/+W"P\D[>N0,?V1A=H(@*5)NH[((<_N;;N2HMR9Y$=3, GR0(-&:
P:D5&KY31"6@Q],,RD7'I/(JB"H]7<[CE/> ;LX0*).H]8$O=4'@A2V47IWL\Y\FQ
P?KWCR\3(=:[13NFUFU\9)SB59Y7PZ5#P\2X8LXOV0<73H%:A?>EO 7CXSS0X[4@+
P\S!06481MV:TC9)4NP0.0Z5?B1-2#?0^9]])/3]I7[,@;,I8/W+R;KDTXM-=-=]'
P511A$O%<(N-]MS11)FX."#M:DAE*'-ROO26UF/LJ1!Q"079&N!WO@G=[44JZZP)#
P6+E=R;QD-KUEQ*/;OJ=54OB>W]C_"MSYX"@DAR^PJ&D$R=@H5TE&)B-C1E=ZNTKJ
PY)8.(EA+!5N0'^/=Q AA8WAAC'J, 08Z!9+H.T>P4_"+:1,*,B3HI0L?9X-;( [)
PM=/P;B9XY(M5O?C"EY\*W,[[J%C?BZRFEE \1C<\@C]X\HUA;.E]QJ+" L,2'BB\
P"RV+CHM=%+IH6,:YO:BE0932L<$&$F!>V-LV]TU3>:++A2^ A*U,OO$KF0#D9FZ-
PQX =9X++-55B!G1X.NNGOO*82+_%NKBI I&4[9;6P%V1_]DJVTI%&&7QF^&7[/2X
P=T((7Z"@S-M@NC'D!F_+0^R^6KQ@^83[+:FLI(G?'RRG5="!6'U!4AUW.?1B'XE+
P_> .3: "C=:4Q_^IZ!2]BW6+Q FA<UL>)Q/J:S^34Y.%C<$[E@92NF7S77@8WLL@
PWXW*$_>\]$</\.NZWAXTL'C71JP'=AH;<!LBSIKMI9OGA8<7%H=DL3C(5@G;&KU!
P ^GO8X%Q/#^Q#+X5;RROJX17JZ&T];<W/3Q: /M25*;J_S"-8;S.T*"MGD2-*2EL
PGQ?%JJ"4:$Z6RY(%),R M'/BMQ;#9=FT]2]U[1V<&9<E_69B_FY(A^H5U:X=T]E6
PO1A(:;>4MPU<KB[3G,'U@2S19?G7&<\=U[=.GYK'UBZ)+ ZE>73I3)2)_@)>)O\,
PA3TT#90!H6;Y93?WQ6]1THC6;91T2IE/S,QPG&OVIK-CGR7K>,:VE7H7 WYPW0)1
PS$V.IT1V@_9Q(.V4T@_H5X.+TKAERO3 </ [MD]ZDBS91@[IBNEAUT2XI&5%^==X
P)H%8\3G'0CYK?USRPC5>@S?VA:+!P0-8_IUND3S,!MX\"BYMXB>9?!W58S=!A/".
P;: L>4$VHCAY0]EZ6M@%SG8:J&S)1=I#J5]2IN&UT\)@ ;Z4,7@X/D1)-7VW#$B;
POAJN:MDU L_VT4?EZV<F ,&TY7^OX&*/K^+5#;RYG3HHK>NC@%P,P#8)#S+^Q"?=
PU4Z7_^7!$=M_8/29+$<?8/,%Y!09B*7B8M2_$5Q#B)HX>C<OIA]R<Q[Z/H)&+?Z>
P'M%"# 9Z<LQX[(''?-5"+*[$M:F(?2L%&*"UM7_WL#^,N&C1;-G7\0L%56LTYR]*
P6? #E QHDGO3)>'^@EK-C/<J#>5'L9X'_,!Q^N=(F(:WH3_%Z.MDS"&>LLB+4NW?
P9U*EJ(6Z#,4(1XY;E2*+;++88'ZT!1*7%3*%?TLR'G7-7]3,RX()$Q2D\@SJY2 \
P6&BVR)GUV(EWPO]R;1I/,<1E1*,DI2B0#G0.\698C*PP ZZ!&_B'YXNT70[^NL>V
PWZ(S+G$8MD1Y%MQ+%M<7(- *_^T=OC:D#.B*7!O,3!]B^@8RY@KDBKC%.08+NR58
PEO5K/].[EEW_/#SS'/+T%#0H9'3"S^I@DWULB3FFFJ+%=29.R72#-FK:*&T.S9D[
P^I=2\6KB-^X>,L.G,XC.D))DU1IT-FXR+=D0&+^4DVQFC\J?"_$ADZ>P79[!&/9M
PO/-_4]V;)N2<=XR:M_.ZKF0-"3/4D%?2D8B(H3UPU:.5H+V$('43-[U9BR.H@E.8
PD[RH:Q?_!$/X7*S0Y+,0TDL"3.:B'XM[#K!:[8J8=%V.[[4-T#Z41!H&SJTQ;&80
P>Q&L1TD.&0WNX#-NF7IGHJCF'5;YI[F5B)3OSX-'WR7=/MI%LW!/AH2&C M*_6F>
P &L0TQI1/(,.=<X?*9K3DB@<BH"=H7%.67*Y)W3W9X:+-W?-\7PZ<S_C?!5V>!^)
P<[-QT:0\K(NNZ"N_BLEZ<AR?Q?_(2U?4I#%8Y%W*K,9-N($R\EJPKS;&PP5M"A55
PWASE%8"UJ "=3MUEO#9?1.XB/?SR%EA0+(^3GKI\\['9J(H<Z56-]^OO6'K(\UCP
P*'WM((W*.MT#_;_ENNDK*IA+:9S_$U&G1L+E)FNI&-,E-WMJ^?S /WM$[_"3$S]=
P^V^21ZV3$Y YM78-RW<9B1 L4*?0+8^Z=C^>7UG?W"O?%O-X'-4FXV!8EB@B[OU]
P)9_2Z\BD,3AO/?H(W-N*P=GS@BVFUS1TR1Q_TU:>H_(X024=R-A,V]):%^!B7I:E
P=?*#SU.H^\2-\AY^@E#>"+AT,>G&VHYI],"DTJ;J>V)HA:F0LCFAY+U#FR/3[_+H
PB&@BX"HE4*]FZ'L/@2>*DMLY67D?/2UQ!.MA<S4R]1.[LM$3_+6F92I;QSX\+970
P9[=Q"7K5^P)&4D$ VWH2DL+,68!SP42C?$&3!MMZ!3W5]ZAEH:#-J9<\4EKIUN1 
P,JDM7I5XLG3'CSU2..)*L,2'EL"S7MIM'CVNB\XW005*(:M"O6^<1(SHBR?[5$!S
P&$BCN_JI?(;KJO'$GPD;)C-&75=LA8C9[]VQ'>_T:\!*9R/); COPS<I),Y8#@-'
PV%O98X)>U X;RHZ]6"1;&-/)+LR:Q4\_!/F;3HG8\A >X/N&Y7-C14)12H<&FUN;
PDX*;-!P%C!72XGH4&XHE;,8UBENJXP<Q/X""XA[M3(#/O"! >&VC[@7HH&_W1UE\
P^'Q7O1I+>(M!]CJ_>Q/V29D B4!H%G>&%SI\Y6SY1EBHWIT^C95 I3KQ;>&S.8(P
P$M#:]N\!=N=/NF?@FPAW&VL5!BDBRJ%3^:,HO:A8;AOYK\H?+2<CPK@T[@B]% ;O
PIWK3QT ^)];=2/0B?:R=522 ="2<45Q_DI#?Z_$#@V/2\AL(*:\,=R'@"#HZ.PK*
P/Z2#'D)^"7.58E#C2B"1HU*.&5W50SV)SR>-FL+:]!$/K.#JV8V[;P[!>HN*EJ5\
P MW\(L$@L$&K305=RS23G>]J4*7?&J@>T;MJ C_\<ZIJ* OD1!F:E<@1EVS\C/57
PLIX6CLC]4"N9<OW&S./Z(;##0';5$/,[*'HB@T?GB),"T)7F1%E/_+;80E=YNH#'
P??ZJ"+K3T-2O7;=,WHMU=!I;A(C%H&EZ]Y&8Q;03Y.2KATNLAFBSV#SR%#WTTRC 
P@55.F\- !5/(1<I.5OY*,RIXAP2PD;S4,K[VTT&JT9LTA^_D;/I(J,(W1 B_]% 1
PX3CH[K//AM(2[Z]0%*1XBPASV1(0'AB-+7\N&"!SR;%D]FX(G^'WV@2PH/]F)ZN.
P._9%(Y2K#6!%HHI<P7W>E_OHW$O\K0<J;5+*Q6<MAMF^NM'H< <*,"YP+*.7V2E1
P1?-+HHVV7BS_(P" SL8UV*0UU$<Q;Q:GR/2Z[LA9KH;]PV"$*2CSTF9OSRX\=5DO
P\+(OP1^:;A2"&$!<,ZGKQHU6R=0UH]9:V9/^5PPI7IJC1&C)-.-R!KOP6;>>C0A+
P"EMUF85#>59>D$VR;\.9JH3EO#"DW<G$04YO:XHWJ40H'O&<$^B,7HYI9(KKE>ZB
P^(P[1/L3Y&WYM7RQ7+2@=<#H 0G0=MS;+_YHX"YQ\MJ1WM6I#7B!B_0_C%+IP^,2
P\Y/EZ?V/ 6Q$;8)QU5[JR%O]T8)P>H+!%7(<N--U$<1A99Y]< 9H,(.#7)%>DV,V
P",!='J6F5"7_I59PQXTZ]).\C9T/-7&X1%O;CW(Z]PB&5"O#X+ )U,OM B<Z U"^
P^5X4!G?JU.R8LZ&X&SE[+3)T8(V^W09_THXW =1A2"UA.0O_HMNIJGM%]#@_W<;6
P?5F]N_+'V2ISX7,.WD'$>'2L QM DGS?WP>.=X.VUF,FG3GKE3\KI2)#FSO[OZ>E
PZ+T%!ZSOI B+F4P):L68SN:G[(E!)QSVL.!AUW#1,:)*;,&5KP@FX=]G/V>#KS9U
P6Q\3/(U<RTA+?A%+\7Z;[^<<Q#0RZ'"&DW,9X?PAOU\Y5_?43,9*RFBW0]Y3,YF[
P=4;J89+>.)V9!%ZK[J_?5,K>&V\TE#Z=E)7!BNN0S4;(8IFHV]F+Z_K)%HG0$O<4
P@QT^ GSB$%Y]/O"%'0FE6.Z:IPM[#EZ/8>9QKS:=N(FX:+JWI)]K^,E/\=SF:*XW
PB9QV])"2"&K=KLN>#*[6'R?(9YFIJJVBD<%&1Q"$GA(M?[ A=(U!Q$<;1-NMGU]V
P7BW+$T3U/B,N*[E&V,8^O=&X>:IK<TAX-1KP!,V9AF:G>ZJ>;["^&"R^?K-3"R_N
P&''DZO5(>LAN$3ARJ2-(H\>22>O5DVPKC6\W)VP*1P.%N.)IH([/Q^OT.@)*U\/)
P272O:ES/B']7KUKS_W6-Q/8@%H)1"YT%=NTAI>[."02JXEDTJC:O6X:*<KP5#_K6
PW5& I8 ,]BZ:7O$I/E_FBW]MQK4J^.^J:[/_0];VOVL6]K8#//??;J<E59M/(.(7
PK?6FG4%KS02  5'E<(O0>9K_  [/*5<E^"]>CF)1TLM3O/-A;&/L_X>K.;:I>-D"
P.1QY 7IU)R:+R,M/ /2$V=]5/C$.</<!]B[?67^@EJO6*JCJ>_^$X+#(E$+[&O=]
P,"E*+Z+9ZRVD+39+JTRC1CZR#GBL/VAJ_J3OP"ATY:I6".\5CPSDN9V-R+E)247.
P,4,+:7;+^0AI7F#YT^+]YNI[6$(I+WTQB7RZE)P=B!E\\_[YVC5Y7-FHEW/(%<(5
P1=2&M)=>'^\XIGJ^[TY:G-J-Q/M**4S2JE8F&QB%(^/KCEC>ZAC1O*PR#P!'2? H
P@%XW6# G89%ZX1Z I.$A[U?@)U\='0O%5AUHNW-GY$'GF=)BKTF?#0W,R,F<IX0.
P6PKZ8&TV<' TIN9QH\2#.!+SA1$$?2 C*XW3V3RZT+X.6G<R:%Q1*M<KR#7C[G@H
P71,H?<U!LH1EMW_0,A9:06/HNA_:<W,:Z WT6J'OL>M\,3E<N$34NFS,=[]%MY&$
P23/>W=4&,"B0M,KJ>NQPIU[)"RJA_DU(R@*V2_,?CCJ.K"$=(ZR?9/:E"SN<XEZO
P2&060$^!;.A-C+#_ (@+8Z(AIRUJ+2ZDW%Z+4F-//[F,3>DL ,(T#\W,SS(1\G 9
P]I%T,ET_3_H5;_)5>U@Q<ME]L9MV.3!I0GV:OGW+5JO88#75%J_Q'-) LBR\KIR;
P#C;8%^I,E=YQ"](6+N:-Y"IL.%_&4]UGN@L-$>L-KEYPMJP,D"0G/C1-0*3^U;VT
P!*ZS&CV;70>ZS;3?0-"EEFZ6RZDV$5_8 >_$?EH3\'/M?W="Q\ODCQUB(!+HSUIO
PUQ?XJ(M&0GC,-E4^H-16K:%W-SNA7E>\1(QV+?D3V&J-1:#E)TT"]"8XY5J4>O+D
P30O/RCS3^5)C:9>\_JR:,G6O=*,^0UJ_WN7,-VAC4WNMK!<D705$'T#1Q<-DG:CR
P+@K6-<K0L674LOR\BUH%S>?TI1.35-QVT;E>9@;CSH^>[4"3@4IA0FJ4EM\'IW#S
P8TX%+?2>6T;JY .C2P]TG.91GO99S'R.W]1S_[GQ71"?$E8 ,8FZ<4_^6ZX-IFZ)
PZDY=;O/Z>8 68B =(+4E>_OE.N7UI_U'_+V-H(%GG75OHA#7868V<@BA-96=%*P&
P@'V&F2-(]@K_6?W7R-YG 46$I0W:BHN90+]*TP6O,804.:*9*:=#)#;D21D'-\##
P&B-* _@<E,RE!<A@IS.ZF[&-OZ^ECR'>H!IWAN4'Z>>:M$+=7899 0<T#%D7SORQ
P8!P "F0@J?I F$B_ E!(6<N^SF2-8D3 T2P"3MIZ\ 1<IXJ:%HM:Z$/JSOO&9OBN
PG(RGUN7*W&L5KCCQ.<IN<$!\W78/!-OGM7<=OQ]DCHT[W+U/S!)%@48=^>8B6#L'
P??O%(_@FOY/ /BRA!VKY9=5PK9D<@KO>B%+-RJ1R3DGAO!3+=/]WRBO!D%S=(0N>
P,3 %Z4+^6J9.HG_)Y&6R0D;\R(#L^_63JP2/YD6UM0+@'#K>V9J /Y6"1FVT$(XG
PL E5$Z=R)S^%"@!,7 ^A-R.WY_RXT3U*H%U18,25_M D'A&$T6?_@KK#>MS.^BL#
PL<R\1KC45D) !(JSX9. 7>@!$WV _%:C 716$\9),#V(!5H#\'E2+$YI/;/34M>K
PP.X/6->C"+ 5.*5"#*@++E>P@X5QKV^=_WHS UBM#@:6MF/DTR^"\O(2QWP_<3&+
PG]"R+P"S2X!PN!J6A6"Q\>*>NP&516?P*EPIY ;TKGO5Z^C/6MDT?980DK:INE2 
P*+1K<J.5R_\2$)UHF67H D I@^X"->T?A>1A+55-')XRXM=:1S%?\WG+$M*R8%LT
PBJR(QW*R&.5,0!"-L"<4,0$9-BSXO"6R3*8S>#1'4%&IF#6I#/N>]&K&;8FZAFG;
PN4&>VL# G)4OB<<0\$3HC>!:2*L\#)H!8Z$T#\6[SK#'X1FL=J 33ZR2D4XKZ$%+
P)W-.DM1V@UOR&1EC:(2<OYV,0>2PIG\ ?N):$X2ZI7N-B2AS)Z75#0F1?+5A,4 K
PZ6C %/)%&%)#76ZX.,B#^U8HK2Q_0&,B7WKFZR@C\0GZ9^6$)$(-.VD,\'"HC/)Q
PZFDW+ O']KY-<B5Q$O6<)G8&A/!'3BU.^:XDEA^#+<+MGT6-)?(\F4F=<'$#T0'4
P@NG>Y5F!@$95PE?Y"O Q+(WNH4<[;-&#@\(TOB=D9&F1/AQNV:JF FC5YH)5!ARF
P+MH84A>.E]&G\+$;/=S%WVW'[NWM+"K6T@;,R*2R\F+'*VJZY>TU6X!="15-M657
PK=^J?1KLF]<'X8Z(8]<6]R'VVP84'C7=F68).Z#NE,%=?^ETD@7">L6)/+8)(H@ 
PVLQ)#U;AF6131#60F!?9P3-A$G ;TJV>,U9'D_V.A&'&D@II%C3%%O*GL8JM-$L2
P-@LVF+F\>^Z)&3[M>HA$V4; <F:Q$_"_'<^'0CEE9)WZ;DM=A3G*HC=RM\=N&"G>
P6(SW5!Z"H".P0KD[&O&@QB@+B\@M)JA2"1J4[Y2X6P&@Q8?YG)NA(6:WUG:US1O(
PYB[-]!,_KPG)N%H,&*L5 8R<M9S&D7\=G%0]!LZ<]@*6DT:(5?V* +/PE1'"R%JZ
P.?%3R$-SWZQT7\@ZY55-%,VU6Q<M3[]^>)7RPQ/Y29M-1\5B?)P#69)PK^0HTK-#
P)(N;\(9KK)\5F831DL8O;[T#)R34U"PJ[*P2(I C#$6__1@*%Q)5X[Z42\V>*XDV
P *@*->A?WQ_IRTJ+BP%B#9S9Q#C7:QS_9#0][$-S$9@\XZ&X5W/W#Z7J;MW[F^0/
P<SV??(./E4+J@M68B.M4!O01M]!EZ/RJ)OJ<^OJR0PT:4$8TCQL-&^V02696CX;#
P/H @&-6G_Z+D']4V"=*QC0"NX6:5I,:OCCM=1HB7L[;8TH"?.]2<7'T,#<3T=("3
PG8-^6S*YP!NFSS@X+*+0OM:CQ$+_E"MRCO<=#IZ*[M5R3#Y6PL$2?9WJR$TQ?/U0
PD%#"/( +6,B D_GR[@ZUXB$X6(QM'2Q>;)4XD-TW<)J28NTM;0<O ;:7B'G!:+C#
PHUJJFK?HR2$VGM/NTYZVF>*0Y(I(%ID^2=@$$(Y5N^Z#8YLN7H(@Q-0HL7_$VNK$
P=XR;\?[%OT\>$2B$1A'PY;[6R\<*$P4WN>=E666U1%*4NBNX]Y>2LJ-:J3!+:O#@
P.F!;^TV1=5L\E?>C.*#^*(1-%4,%Y UV5$57\%<)MVD.$<F=\2Z$;LG64OPXDF7(
PQS5,A="J/#OPW>J'JUC?18?P&R6&AJCJ4N=C63=,$6TD38;=BM*WU[7YQDR&N%L*
P#:5\&[/_ _>PQN&9:&NX,=_&-=/.6'Z0L>7G=!>> VL'26!(+++NE3 FPZQ,5U'5
P&-&\+0+9,FE\+2I+U)@:B.M1@Y:04GP)\)@\[F#!4:: ,MRTK'1*QZ&=2T:C5]:J
P>IZJ^C_$@;:INU?*]I;T+QH6LG*KEGP6IN6[OC)3<.VII]$.G#I6X3?'H1].(+@%
PVO,H/;;/> >Q#+":E$]B IP9-UNHZ_AG]]XMA>>6[G08ZG/528WG>2*W</5)Q@9E
PM$N>P/:EF#D#X_[-Q',Z4A#/$]69:TT'^H;B: T3S%PFC13,%^K9HZ'B O6Z$!A4
P<7C(@:!TU,BD]3F3'JQ%%.\P-("NOG*()?^;(SD.HPO>8]H(O& D3_5MTJTT48I)
P%?EGD*YR:O[KR$R9W*]G-9A(?574<#/=54@->?%*B(0%U?),HN!BRY#^8E,Q5!/8
P&LJK;ON^?*$=5Z$V%AN#@Y! /QQMC.NT$.[VGL_1PE4982Q-G7Z$U@WDZALBO>B)
PQ!E^*2ZIV#=-HP&?/7L9-CO@E?C\MR^E4K_'ZAVJ2Z^6ZJ#I4$#$J@NO42N'RH!>
P":-#K6J=E9X=@48F=R[]8M.R+'"PSI/O*H]P.I*@ *67NP<. .6;F 9J#>:D7:'N
P>[A6X"G11-2>W((7=KCZ1&TN1;U>7:W0V5>((.8AF@*T@Y7,8?4M@XP)OKGQW*\G
P&%2_J)R5$R)(4X#)PY@X37D9!;* ^]Q?'2O:MM3VG^6::L[7;&MZ("D#.E2-51[%
PXL^)PVESY@O28Y?VMG="&'X;$$^2TE*SX@4]@$/5]?:GFZ;;V8*_U4YG9A%&6V4;
P)IB$]@+:+SE'*@5Q%+(<^T2 FOTQL9F2.C=,ZM::V":-XL]G\-2C=[O@W[A&H\_Q
P"4U6*61[K*%U0,%9N\EKX(+?ZXX0@IL.\@'*PX:/&K,W$:\L/L>XR1KDT+\?/865
POK4$_O\9E(T#U*X>J=:8LU@[1',:2+Q,.).,6<,2)!6\9Z&?&JU\*GMNQ=99J7W 
P+/3T;-QJGTUW.17@(AIK&X62U,V75E,#[+>+MCFKU=;P90WEV][ZHH1=B+IMN].L
P!(NU.$.Q*MW8WQGCF<4,?!QE'K(=A,MQA-,5_@L%U/V"QZ;=]<>\\10*"HG*V_R#
PKQHG?LOW.Z\[M<BB5YR_'O\ (P"$_C[ &ZECQNQ;*H-E@CE!Z1CD"O40_8WUZG#8
P2IG@S-D26S^9(YHB1.6Q^*[$KRE.W_INC/<_F79'&YRF(U1+YE@!TM*QZU*<+B#)
P"W0-A3FE1\Z46YE^^*..@MT&ZM[ &E8,]!*_G"Q2]DNK),7MXYS/%=ZB&$B 8[8T
P]ODSI]Y*J'6GJWH@8JM,T=D[5)&STC94$QX.V8V4)[._&P)]9RRP.K@U!"WW@$<T
P'UNHX)1Z,: 7-S U=6I(T9CZHK-82@C[(Q1[I0'=NOR4HU"+I6&X%GXZCO_C8EKF
P]L7 8B/#X94#C*"+Q<23P)N]14_]SEC#]J$,5G)APLGD'GT+=.M<!H5WRI@S\"0?
PQX':6.R2;$,_)R\OT&".41#;%<YOTTX??NAM=2CSPIDFSBV3B9C-7GJTW;V1WE-O
P]+7/87BDY%@.UCY0-U3 )Q'):$JA]V&H9^ZB;QP#%D8UN%=!OH]S9=:<^W \;M;9
P'OT+C$4DP@#%"IZ>VRN:!6B>VD-F:X&2_&TX"#=9'G<6R8-XDX%J-$^8<E(8K??2
PB[OJWR--JUQ>\AJ63JV0MJH*AW^)VYNH6FTQMC0R?HQ7AX!P]*[7I-'"[%'#,HAD
PZRBK#6)GZJ9C_\XCP*)*5?]F*H4%FP2;9[6?<?7/S/&K H2BOWPG40*M,[:&L-?/
PVV-\$M5D)6G?7;Y-R,O] K9@9JNE,!Z(0AZJXX8+KK$ RS\PES6AD0CP<9LNWK-4
PK<O57]"I$P#BBSV,WS@Y;\V-+]5>[[WJ6*(*CO,@!8'UH!<>=01@_ RFE#>\ZF5D
PIBU8=RP&#;0#[FH_Y,Y E^EG_"[?^:PNBP[U^PH8B-0S^JXAT>O=];I+CR$K"&0E
PH;9R!:99X8@ D(%8)]8:AD8C'8S,MO;3_7;7$J](QQ7)C<AK488S*_5^/M!Y WF^
P^A#_8R,I2BO;WQAR3OI>+;X0@+NX:03.]Y.6LD@+J *##HOBQUOS"\[*5IP;=-?Y
PL#J:GIXK)P94 F"M+*7PY+V D^#G$M+RZ;V).5IMPS"^G_0**]'8+J(7S# /K(8=
P6,8,ZE,I/$!M-(:-@HI:VN2M.+-0EH#98HB<N;9>%F_M>2&!<D@2\AMLNKR"F77K
PXAQ:/%.AJDEJ"B7RL1AM6V*78W4,Q'+XC3?/K6M]T,1DX_AHFWCE$U4!%8Z/WO8K
PS"0RO!39HV=^W1H4<NE7)F_*_A9P$Z*I3MG,H.2W0BCN/9_!DRSYP G DP.0"48S
P.NJO?F]QYWF/R*.B,NB(D7)O#7U3B#O.U$WF+"#J!IF*ET1@Q>"/,V:U>PP=HO-]
P()<V+8D"T4:Y R(FB(G;<#=DJH\02CM!R*]W/#<Q.GMJ4++!&MN D;A"4DRO-ECE
P\[3H!T2$YYL<Y,$C#60.TIPI4$6(60P@1/"=4/5P3;Z8/(Y[[&KR+ B^82B$+B'G
PK^.Q;N;VBEF&5%Z^L9M7D=+RC^[4=;2@OP=+RU\2$.,-;79+01NY':/=GNG/6)LI
P8A/;ILQ8M^_U_"@KDF[;W9Y"H-JA=Q2CU8OJMD_W(E[6YZ"N$2S:]=@*S#?-P@6I
P;$#RI!')[,!]<B6IR8VJE >UY%9[(V=\N( W->/*W]Y37AB9$V-=TQSXX,AMO(WJ
P%PV>RUJ@@*9?N*KW4N.0OB_%EY$7O(3:UKM<(PJELO#!+W8M/ RF2]\+M>(0DTT]
PGLHA+]'9XF="B[F9L!S_MRW=*IP-L3#%\USR3%8_6':L IR6:[/314B;0IR:5Y4E
P&!=#NOJ8/&%\,CS\ T)\>R?:'<!&"RE\LUW,?5TX8>,*_H>!Q&M>@Y_UPTM<T1N2
P]##9[Q8&5GI7UD !,3B!PFVB]?VX(W,C8-@208_I!I_*4Y7ZT:.=SX+8<6!72PS(
PSO4ZOY%!;51TZO[2(FM+JC]IGG==A%2[L_>A[1-4BB"G,8G;(3-_.K4' !.2#S<O
P['9/+C"KG"*J*DY$^9]>^J&/\*G39[AF.C&B4?#S;/10F+A]D(I7JYDFE]:Q\19I
P//F"%(F_KNW4W=\EFF=6-7W#TPY$KM_S% +Z6*0CD5I Y:SE4?4,=#H/1H!JMAFS
P8=WCEF>)W?CYEAU^\3S9J[0J,<D+KX&)E\7'1+J;_&=TY]F^Q)@KOUW3[8[!F\%.
P<QM=$A5GP)*X9VW )-,E>KOS]:V$9YM63)-SZ]#:U] ^CMRS_02P48F#;F+ :7L'
P:Z :-?$1ZL%91DL+.4H3.D1[&"03&L=%/UU%]E,QXJ0,7R@J\N<SO'.8"CKX^+)[
P\G/E(8H(#%"WM!EN#F]FC_'Z_"W<Z"1^R%P*_6H916L0SN:23EGN])%029<R2]1/
PJ@[U;?>9KJ/OV<#YW18:E3)+ZD;:;WW'=+ ^9C,?<(VU^:T02DJE)S*C^I@&)V^0
P;_+YC$@:]<VJ#24;&3F=,="D@)\26/YPA0Z*AK;#6RBVN-_0RG!TXXXW#9KZ<?W3
P&BI&GF.B:+,!% C&Q0R'[J5=,H?;/;T(-1I?#70< <6C-1:#:\U$*)NCQ(1HMJ%+
P[<)+(3,W+Y-/\JC#3[W-;8-FNO[-D54KAQYM&*0GUD1"N?7 ="N]^'59SI98!P8]
P7'3?T'.+#'LZOF_-Q88)041 TK6]5:(<9&1(R9&+Q8>\>6X#T=$X+9(.41<\-K[=
P3I8N]"-(TNX_%M55BY6<B!^./*Q>VF5\U5?Y4E"5KW7PCO%9IW3'LI;4\L^/W\E@
P*YBEG@0&:W!KI@-P'6_/D3 _4B) (6<:LAU89(#AQEUQ^"TAP=,CLAFWR4:/ #17
P!"Z%*+LLKAJ;0XI_LE>\8.\0%>YXO?\7^JPG  N]5BCG\AT\B_.2&23'))+Z6[E<
P$>.S=ZC!J4+U]A\YE\G4EQ@CT+A:,#G'!58S0!BXC5@L& GM DV2NV 5S;PC\U=&
PAV'_3XR53FWZXL /:>:!-JS)FAE 7C35*X_$$D:>#KVFFY4_U=_#7G&GYL/@P=UX
P_WCZSI58]I\@BP$N@'^W3/3? \X26:-7,I!T_-V#@ \&6G<W/E1V=:P9]?AP'ZCY
P&TP\340-EKHCI07*I6$.+RE11K[P(CBD8CTT4MFR>%&]I.)Q-ABOF'7W"9@:QAN7
P+$?V^=:+$)Z'LS3SRD^JIVE*<>#[!P&+-S25D'J@08@*B)QNQ;^)'2&3[=_1+SCJ
P[AKW-Z&F=%$_RR%?H&8^ W];RIASXA WY>$/MN7UXL.<.075!<I%0P)%XA]';WG>
P[/,ESF!!-VRSR_<#P'1F<[9M1F0A3,(H,K-8&)X-MKM.RD"&<O&1 QLK-I]KD\W)
P%AJ"I!_.^:N/:-#4"V<[DQ2'D[.EA6X,LDV7K8K)0-%7V/]D#N)L@M>.L3X-K"&*
PF,47(126[C)=]EVI,*VL6(-G=I?B7@ZD@_,2M"!RZ47AF''&AH&E[R"I-TY"ETW4
P.T&G1<L:,R^_.Y+.&_Q4PS_Z]1YKY8DTB)1Q'*V.OJ \7>^:CY9'J$>S+]UP//2N
P?UR,K7STXI3F4HDK(1G?O14#*,7# 5%K O-UR'KA1G81O[U'S)L2OV9]DXR_H&QJ
P*NH2"*W,'G('IDUVVW3PC_5,H\>>4DCE5\X_VMC?S4'40S%SY9&_TW.*!8"Z 6DD
P:@PXW$Y8PU6+\N*:R?(\Y!WB')N/="47==GDQ5HI!=YF\'DLO]N=]JU8UK!O=/C7
P%I1=9;9>8NY./Z[IXT>UNV4F3,K/KR>ZALKJ)00U%VM$D+!33\Z8853I/$X'FF! 
P'W_2'N.PM654<T@[&3F8X6%JX+;;$(-S%PN+&:0Q5+/ZFFEZKIW*EJ^=';\A0RVN
PRE!=69$$*\4;F^+N D"0ZE5V"Y#;)[R<[W%1*5#D7.G4]FEE &$R?)DKQ$W/1[[;
PJ216]$*]+0LWP=M9W[V7H&7@EZU_ZM]%XMQ0Q:@%L/F1.@]6UK>@6,'X,%H"WMB0
P/%(1\5SO86W9O(Q37)&SH;\UQ*X?W2N$TQF4EUYVG)]'V7E:DSH&>W?Q%\:#.BH,
P:\$%@AASRVY-CTJ6AGL%@V7/Y3'5\(78!!6!-TRVEZ6W<49UB7]RP#$P%%Q!BM'X
P4[M$ 2/B!T:(I4I4T#0-<" =D#YZ&0,?/5=DF6!A_,?WUGZ9&=U]0^,"S,PL;7GY
PC-IMSZ0:0UZ*60RM,>BN]J+F$S,L,UG 6YJ>#JG/O81)TEZBP6!/$#6;3X9 /]@C
PN[US92O73--U<T;M&_2#K28B&A;=?0-*)UBQI[C!RR^A^M\]I7HBR_3KN^ :/;@"
P8TMBT$@BGD&-!9*"A$G$UE1(N]+#HU']E!\LOC<KP5S#KI4>$_V>G,P<@$B .I;&
P,[5PL:MYRPS&^HMK:=+*" JS52AA?+L:_^K4LM_"7$@.Z  ;])T?F^"5!;*$NY+V
P,9[^V*R5$.':=[(F5(>3S[#'1"(SKVUB=_Q\&FZ@+?L2YFO.D 2O-S4[I7)P35E4
PI> EY0<*+]"'OZJ+OQ>P>>(S2=G;!2?WQFLX$35;R!LEK#U>!.^)4N-_*R!L4Z1K
PQ5_*:4NLUFV+1ZAJ5PB&R0NB-=[K>+/JS(:Z%6HD7YGD?9=($'7&SQ)4&VXHK!, 
P'P$X49PVD>@O[28.ZY;BA.+$GJGJ8L(,&8@9EOYZAIY- G_%F-G>MHMT-7>E,M1 
PZSH1R(\TK:!LRP\L4SQ B+_TX8=C6JTYR82!>Z*N=OYO;FQ^/+9+.*YZVN4B$U8T
PMY<J$:W*(KH*=)MT &>C#A>A%,RH:?9*I_+RE5:Q!!Q"K6]@,O0J,)Q?CS@IOT+H
P3W.GE'BO!E))()V-ZX)W/)F[G4O].ZXJC1ULD1? .<Z46G>KS0U?$>QLTJJ=2.R<
P<#6*0T'AC<C=WZ<$'#M+ONO0CE(;(:)<QP(;IS4RZ%AC,E6MY8\Y1:2.F[&Q"G,Y
P'*1BD43%8_-\5?B"S%AUZ^3%&!@1TN$:HAURMP 9YF;^HT<J<BY\WV3.'4E,*J& 
PW%YR9/)5B/G!$I^-2Q@J9@89<&H6Z:]2?+E1HR&*[H>59Y=Y7U&7#YS,>$S/I]FM
PP$":8(. Q0$*1=HIRDGEGZ*'QP3,5+5X;6(2S?(UX5'P60.6J\4DV[L\["-+.#)N
PV=;;363+?+3#01E$ES"@.P.HFG5J-KG%3E<.#M^X8B"M*)%!N9-L"/;-+'0.*/*?
P0X:*E1R1([&4W#)YFRW_/H7HPQ/7E^129O"T&>AU'H4W6^KK9'[=4_8_1QE9LC7Y
P[+.K2XD>]0N84]R9R!",VQZ6SOKUCT(11W@1:A-_3VTS$U\3^M!B6LHW&^J+ /18
P+1G^47I?B-,6CD3_BI2M.=:TF@O1-BI*N\G$B#9U!P=!E0>!I\;/ UP6AZDAX"(<
PHD1Y&K/. HW/)V&.S>SLGT! 38MA=Q.E1,\2YP'BQ3#WUTSY=$#)#_:BRYX\=D_K
PQD&:_\C?Z9.E6ER<^,<>ONFTI>Y*CUJ9H[*G!1 3@+E(8+>]JWU7(L2R*?$6KZX2
PR0;<E-$[APTH=H#*F..TN\H9-5!NS!MHEOMQU>]MB/Z;U*DE@5>3F^>-L/@,0AY!
P/[]A(FWIE*,B=T1)FF]6^8K87RAIKQ7?T3&-S)RQM0JWD*>KM0QEMO7!A/$?'FYL
P5$KM:Q5CUS5EB*J3IRP&NP!>CG^O"IQJZ%0,[M$(J&-LCN?<S&9.%$+Z#R].XV*\
PCA_]+I<1^((H^XU$2VU_G*)G-<>4:W8ZZ4;YL:1 P+_C(ON0L? ,ELEB^Z9$3=,D
PX>'Y68E$R[;)BYU3R;YS27,'Z_-N5QYW^CP'^FSIBGL<EH=P4,/WQ"OU[.&(@LU2
PC*;51N_GTO6X8Y8_V<4JN\=ZS4\7++6 C+*@/NMFWBYL[PB)0;BHQSB[95FQO/?>
P[5_%>^B2&7&IZ]LK.YY5H-G]I12T%A)[=)KO7E7F]HP)C*81JIW7^I]W+'A[O27W
PLKP4.W6X6>B^RBUHH%0E[T'M^+T\MSB5.1&FLC>[*?6].OJ.5A65G\FFK)"!%(4F
P:!PR'8AD^86$TS[".2B1K@\EN*RO"7<BVP1$IH>]J]5D[ST_B ([0 ",IS,1'AK"
PI?J=W]56FI1=-%ZRVMZ%]3/=;^V,-)^WN3GPM*%A@QA&S@*CD]M[%45"F(ESPFOL
P:>J>-,.8I)]48O6TUH,*^P>4[VQRTTDK'& ?0,?BSUF$R"UR+<O)-/0:;9\M>X4+
P>M?L&)F)5,_\E>>MV'_<'[L4,S%[N!>ME.8]0.;ICWRKK3E1%, DXT2IGT;< %U?
P&X[CQ(B")=JT2UB,-7#X3@+;LO+9QN-\-J$C12V ZL1P1WBO3))A*GW36@.#:VV]
PI<35_E%71#4[X[%=77J"8Y1?OJ]!?Q%!<H569NQ*DO>\/_4]H_-]\X%S%1-[7W2C
PS5JWZQ\K<4PGTUYK 'IY?+D1+OBTM"C2#>@F=O!(,=?>]PBFU1;EL$W4"FZ2,>G.
PR6W6LC%1NG1Z1Z/6@54T6]Z0L1[E+M:= /)ZQ%@>C1JN*@5_OV>I&)7..C_6FU67
PO=76H::K7Y"XL9J6(>6"<'ST>=ZT#J4)B4D6KUONU0"6/0N6U>TGTP9/GIZ +,X'
P]#TM'M"N9YK^L,9AHRJ51>U74O3! G/@+)B5)Q'+>B$+BX_908G&J%TT*#>0:$.,
P ,7YN0R7C \AM,<_Z]@:%ZEEMK'2^%YD ^K_>^.TP"Z%13JOW(Z1QYX+Z[<-ZF-E
P A?QGL&'>M$F*@WJ:'^>BXV0.-7S]*F;MX=7S,0"L^)5*5'7"]2YPHL19R_N:$^/
PYY=.59>M.8&F]6"SZU8G)O=PY:;5K\I_CG26NUL#,3(<TZ\A.[G73-<?:W%6]E? 
P=$-M(OX*%^<L!L(L@=R$F>;#X5&O>3-V$!T2X_8HB)LE#0E5R"C5RHI4WYH!<8'L
PF>,<*V["D-CZE644'<4I'K,TTO[X!L7F+Y#AMM67::Y4>9NUVU!CE$]OI7/MSIO;
P>J0YC@EB@_WJU*(*$%GOK8\;_$!035]V8*/4S"\6Q.KX;739GP\OY>!L6A5<QP08
PW2>)QB@"T;?7TOQ,T/O$#(,Q>RS;\*4T;(D3'Z'XP3(6]*4WAF.Z0&P4*9C@=98N
P)9T H(%V7'X7J\K!F3U$_$,R3"GC)+?#W4!CT>C5G.@8.R4WNI52!\6VT&@_E@IA
PBYUS(U&=JLUX>]!:R3=CI>MO\ MO.XL)1Z5Q6;X$W=8G#(DY3OW+JNMM]4.,%%@Y
PLK\RQVN5P*PV0;Y^YHA43P'I( &K(;: @S1PEB1<(-L+(;;[AK:?)1@#1(4BL($8
P! *C?"31*L;T^2?HTD%_V*I)>?WZ 'GTMM0P,(%"%#NO>5%U+N->J&@< Z>RQXIJ
PL%E,64,(VI='YP&J[CTD,1G2.!&(36W[-V(5-EOEH!<>+XBSQJ3Z-=[+9Y.VDC?W
P]!'M/[);&2QZE4V9T,#&H,71-/V6>%'\?A>_8V.OY2>O(">9>JDH7![:(9%;.D*A
PN(;;J!^#/!H 1!%M!+,&1_'JH\FX7F"/LQ6>F,TT=X>5<5(H>D]G@_Z:G*.+$)\C
PJ3F(V3?^M;W@]L6I")8C=V?$L8Q,1J<UBK$$HH'K>0@(A$S103#S-S1@G=XD^B=E
PI?:8@9/T'PAQ$_\MV!U6XEUK7U*&9TXF0LS'O>ZY_-H[WSS)2PFL F<:OY0=4GLL
P5Y,**)W0%Q^+\Z,3H$*$%RJ^@PKHP["P"G#+HL/D80N>6XOZ8*$?B!6H,@EBI#@K
P7C$\<;\WX;5CC93N!/*P*$DGK5Y(!,S-QZ(H<GGE(FB1(?0^6U9ME_F',JC2ZWY^
P\-9[9\"'O93TS6VL1C$42WNQX:YS/(BB-4F/X'6)7KVNYC'_4J$Y&%>V8&.] C):
PRP&&((6N*>7Z;\3>TS8C-I=#5;KQA;5;"=0QIGZ5];)<\LW6&KTZD"(?T!Q!I)T+
PF5 A).G0%;IM.FYD*;)9-$V$B$D<QEB0D?H'S,0MIC/DE<54^_FW'PK-"K!6T]O&
P!@AN)/H3.!NFO:LU8XTPD YR4.1''R[QVXMD'K^ZHA&=53C7FO0PRZ'WP'<*E>Q8
P-'ABA,9VG'2Z=Q .+$Q3C6H^DOJ_0)K1_BD<WQ_.=4/24J[A,XS2<K( 78_):-+H
P</>>I#CC0<9?B65PDEF#FT@ +N>V[_ML5^G@NJ-4(ND/9 4K\MK&8D'83/^3&M2$
P%4+Y7G@C  O7W^MQ#0ALGU+Y^BKRXL!D?K./Z^K*Y#JFSP4@_=+S":/AGM_!8+*D
P7/.M_WD@J*Z$:O+:Y[,?L3X^X%TM*^>+G\A,ZX6="P.-.F5CRZ_/OK(*'T5%]O8?
P)*9T"5HR*"LNR-SS=K*G:<[1.2" 62T":31KCJP!+N9GF)%'>@'QBAT;0H6EUH6*
P8TTR'--W(*N+SJTTUPU9@15CQ@S)-N5%#4"2F+&_FU+7R01K?RIRDG 69M_.SD/(
PML$T#&-)W3E%?3X8C/24QP6P3QZG,G52*S1F+J-F#V6K2YT/0-X_Z9\X?32BUIJ>
PR#S?'TL I--@R#)(EEJ7#I.EA'#O=\XG-3:D=(JF8R^^%N=JXI ?XQ+^I=;;9#-P
PZE_P8M$[N#K+$%^W*HS7?DWU\P:?Q%]5,.RXLMJ0-LDCX%DJ2/X+-!0 -3%)<)$)
P*:$H=W=)4Y4YR.^^2\'#2N'W)!8XQBR;@L180F;!%?JE2')'ZTG&_+G-EY[]2>DH
P6\,!T?(KK5ZD:W>,XF_!BZCZ >+)VRE5I8!$>/\0$(3*3;+RT;_U4=N-ZL>COU3=
P\F31[L$C2E0O9(!R.#WYKWK\;P8+U?=NH0LI_>FGG\D4@0K*ATUA>*G)F^%$J2&&
PIA3P#U;U)#-1H<)D$B0FDWW&U.UF=-C.#_C>>MJ121'OT"IF#6;XFS5:.;GYB)3)
PC1T'6UV*=#4?(F03V!E>CEN9_TQ'A40+!CF8YBBZXG^+K7+^!<6>+&$'_K1[W>I0
P9O:D#2-=WP""OW);<.W^-9O)ID2TF"RM:E5SSI>XJNDI&[7<*1[N J\M(VU2DQ9:
P" ^""_Z;]C]F1_O:K#C4;TRQVVX 1Q"'-LQMHEM_[VBEYJ4IA!-D+804P5VKGNY=
P"2>KQ[W,#KL 49B\W.%&SX6;WXA\RHO# A^1E1:5ZD$)+;Q\P><[H<=R)H[T$+W?
PZAH&D=K 5A,,YHZ5C=P2F?JC< GZ1BR\WT,3CD%[RV7;YK90(3ZEBQ[!7Y[GJU+(
P,*1ZFBKP/KJMFE9)<LV%[,!_TNV]&HA,ZEZ/4X)4)Z<8*N)USZC8!WGNSQ_UL7EQ
P^E[GW4$*JHF^Y_PHWW6'D(IIT%;ETR]<40AANO*X9-EN[$;K3N\/,FLRQ%>K H<+
PI&RE)>4?1EQ0V O-(3*FCL(>+D''!%YCC'(F@W'  ME7+E(F"9T<J\)A@/N90BI$
PA@#H!VD5LKU13"A?K<T#KV:;?NIS[OGU3E2]M^@L/$I338E/%/U)\G10+!NAT(Q!
P@(AHMP!VLWU";;4/2;EB=!BZ0Q>DH(N@.CS%O&HW 99+"+!E\@P&\K\9S,S^.HV+
P;X]7(Q_S',]??VZR4\0Q'F)TD8SYN'PIS ']Z#,LOY7E'\!-DFS(0>;FS\.R)YB*
PV,J'LIL^23^$V@>SK%GW]R9S1*-C.!OQOJ [+SE+8Z;VI]]@!OZ8S7Q.GOX[A!",
PFKD%#I(0OVC"K0F]K4I IQKQ42.?0]VY"O#"2HJ>D+\<VPEU5-P(UFE5D]#.SP)7
P^,49G)N#27RQ$RTI>K8K9W@-J%+73-,N[*-&)[)O1 #^@DC)'J#342Q3E'=M+P8/
PO60VP<7!S\D-<#;.K"  Q@=;1TYP'R?#:RT(B[I!/2:UY&;^USCZ!>!?!0\^]T*Z
P+OZYUO85&YORK/3HMUY9J92>Y(6KBN0^XU#)\F_ZUGE&TG+2H]A)36(HPV0;5B)M
PS.5E[-.4!)U>A<'ZYWDU@8B:UGIT=[Y!GMW=<3I6U1&<+"^IUT9G6^0K\,]-V^_7
P)#(C"NI"YXG?SIE(S\'9^CJ-3-DJ5FXBOYKDI):PG.9K=V(Z?Z?&<;0:([==&3G1
PSB8)[9Q$$(X#]]O[9JC1S OW3Y$-R\$GV,H\MMAXV/Q2.RR*I?6JHKN^Q/A,2QX.
PS)7S!A1 "SP/?0U*M+?-@33WX 0N<*+LK*,BS=Z5G!2Q3IJ[5TV!J9'JE)J'$GN'
P'^0[F)Z6^>]$!/PY''2JW9 =;AVO;U8Y"=WMG>+B4OR-:]XRAEG))N])NPXQ<]&4
P^]F?AY-V4.BQ2>F,AZR>L#XVP\5?,NT#>CY.DI3CATX(2#.\5ZC&-_I=.D0X;\]3
PT"<*BL=UAW#OB*F]R VW-^V,K"_B4J47W7>Y5JY![VC;^=]A6N*0#B70I*M9OP[ 
POQ@BS_5;&5A^_4Z,0)DH&$1^J1M;P)I^,!K0$U/8@?ZSQE1[.Y#Q>(]*Q1>NCM<_
PCY=O8QUD<*B'V=&[G1U*H4:^< N'M?&8I5Y+7L$Z2=!?@0=J2BNZ&N;QC^<)IKX/
P^K.!C E'^DSR9X7T"W[T");/B)Z;W/;%_+IMZZTIB]-EYW(\B/Y$FS> X]%V2\=<
PT8,/L]"Z=-)6&5N!!.0,W3Y7582-0)5U=I9&^;?>C<W%(8U?=DI<"_VU)T%@(6]5
P#BL"_?WZ?VWOG2-JO+<M/T1HASY]4_0<F^Z]6/-59@LY07K/;<2BZ7[V1Y#P5OZ)
P\?-7N.DM\;.<?HM%B;#[E@:_U#T247W870K(N(W"BIH8ZZ(?,0(^A2E'&N\ 1U_\
PR"$WG112_ M1=JKK=LD<(Z>LE"BJ6*T'&B;)WSEGF(Y%W.[.&<1G-[H@W0;>N=L>
P=9,45<A;#6[.D'D7OMX7U+W%9CZJ:9JQ%A?SY&; -J)O;8SKG;#HWOO$'S3E*:$L
P\K1=1YS;J"_T1EC7PU.G_.24?L2S0;?"%&[#+9V/Z"8K4RE ^90EI#KFS3 ZZRE]
PK[$>]055'^C7"."L.FON4&G0UA@;$G,(N((A+^*9A9"ZM)9X_=&O7D8I"C?!5;H.
PQI=W2&P64H:[P-C9<PF%=W05K.AS]T=<,=%.#DD4423NJ)P&M,&OMBO6<NW,%>5"
PP_K.R^F3]33Y=YZXX4"6EOB?B[CLJJR")K!4GZ5!(YSWY,(H\2!B7A ;AY!.XQE4
P3*K']5""G@T7)HGGTVZ@ZE&\$<!0W:/:^'TWT)_[2\0+7-<M9@7?DM/R6N9$Y_U?
P!YU)7:4L"#H/@Q_-HX1I.<1G3.D+YK"]>H6@A4AO=R[73(Y"T8861B.9[4-F\.+]
P&WTH2:2:;"3-,>[%-^:%H+#=%7_=;.#:ZSFIKE72D![_^V:,1M9<A-[QM7_,S#/!
P4VN7+%; YUIH\FU\6T?7.+RU.AN=D$:NHC'J1PNZD%V+2]6E(? HWRV*'2_[*#B?
P-.B_CQF96V*Q7T L ^S@S>HG"#*5(@5!:"Y\HP1!5A^^33T@1N+")Q?9_\L=B]WP
PBE-:H+[S[Y@>TD[0DR06M?LA((K.-1S%99=]Q;HG[@N0:,,2J=:-LMU_"</EQ^>P
PE[FQSFZ9J'2C?<ODJXVOP.W# ]KW='737K3I@-7-O&7'HE DV"HK0.S"KP?2U\$A
P'<K0'6%H"^D^!F+C;*V_0C\_RX#HVRGRL8_Z14Q9P<5'U H9#5GW]PO%)<!]CZ"V
P&>#,^!9L6?8+>R=;22QK\Z.H63$4+J.YYR54=*_22-]G&^X]EJ3V78[*K=:(PRQC
PH&8% E/ 6W-Y!_^A!<WSA2%Q8SZ'RTO7"@ZM9M*7Z$<;^CF<?NX)[9498 <.R2:M
P /<@A-5W0/TI.&:CN3$J_78%N4S=U&P,>2+Y%!H8])4PKFDNU5@&[M!!&?I57G@D
P;^Z.F'Y](0NH=#F,=Q+C\EZL-^\[>#75WK%<-\2F)\D@S.-(]#IJ!18+QE%;;OI<
P6+\UL.<Z$WF+_.HZ$C*"QP/5?0#[GR79@ET\IE&8#W:K&H>?'O/0F 0I>!EU9MGK
P5*>]XU/_@"'MI_/?#1K!(LK(.-IJO-,BL9T.LJGB1LRD&PZ81^"L:L'4RDD=/%&\
PWY15Z#3>L8#&? RXF#H,UE/PY*1.MK"Y[N'.:T_0K#4TUJ#[6Y\T0X\-=3'BES@F
P C 6QM7/*#:M/3@ ;^F -NQ[]T1M;;0"<[#H6-<#N)8/*X#C66B7U&0[/7;I_%?%
P0&9T"1H'!QTWA6L9078D4YMFC!>_D5ACGE)V2S?YK'C[94VU(=[L[!TB!_[5/?"G
P! ]!GSX#TK7]WM'/YGDAB>)UZ^G-C[5!B79,OHPI1<2G1AK:N;GP,G:RC',V0357
P4E%Y.H<>DQTW],D!1&WSMQZ$YP,O($C8R1ONT44+YN">_'"N^11VP>;]V:IX/7OW
PXCNWD32Z'/)R?/O+<2E#TGV^C+DKBT<.A2X3?]!]UM-B2CL,L.&6(^_Z5Q83P13/
P4?@Y^HO3B;%->4R]CM+E=CTQ-IV\FQE7P%-RW8"KC(E?+$V-!.S]$9EW8@5GSPB-
P7#.II7G:!6[FS/;(6O)1"WT/@J)H!D !2RP\/J580#*WDLM\;&CII->L"P9RW_NB
P4@"I$Z<*CY])AS21E<2.?7JKXHSC=LY%9A5LT2=)_P:_R'OU!!MFNIL./A!&G%C8
P,E<5S5/U&F#N_SJI&%17[+2/4ARE=;=9FP4HH/ME)#%"Q8R $-VLQ6FS(%YKD\/ 
P#\*4HZ\VK=,+$6.4GS8QS=X6@6=PQC&GN(MSG5MCRG.[C-=\OW"[__<* B5KPMT7
P:/V]MG_G]AN:N$ A#Y>YC1Z C54+L"COB-6/TXZA,1=SP=[VD7*L^_K8-[*QNB31
P=Q@$N4XB%>P<1[W)QHK0D??6R\=;4P)-,U&DAIR#:&#O&9;7L<#9AC!0W!B'A'K1
P%%:\9:Z M?J_O\LE!I(PR&)0(.U4>.<NGDSY@@ !P&QG.#TH75*:,4I8MD-#0G12
P:(9OFZ@__:K(3]X[MV=:!Y+Y]&-<)T,TEEVA <867<:+>Q&0ZM7H,1W>*9ZF_IH7
P1UJE@4">W+^T(P>%1C2,&121S'Q+;=9E/&:7/$<V[[SG =LFO;Q7:ACDPW!$_]B#
P066$U48$)NN0T!-$?O*S"NN*#;]0;?WX%7C)TR=U_&QG,-H?GCE1<#D$J@=)GBS2
PO;/#2?L2'46^B[#EYN\BOYR7<@(+>"\CVX[T_?F&A<7-=H&MQ02BKEIO)+'#P41*
PZ&_NS[-,RNM>PH2U\Y)F&^ 2AM80:^/#.%[GDMQ92=1*,$%067NUX(1RO.KI?:C2
PNUX,L!#/]-^9 A*;[@%J,GA%VILNM/_P>F]_]FHRLP7HBY(!L<F:8B2<LYO"0KB8
P:)3^HGWP9)FJG0C&]ECX.W/E$ALV\7++B:PJQK[5N$7;XJQ/B&5)E<@H#,7B HJ>
P U<:0^ 'CR0<6<6R#LK$O3Y 0V+/=0ES*/J=Y"=)(1X25%:ZCON-%2^'5M[?77;.
P_M;L:B[PX2A-JU%5?:WC?  G0B +.BAV:.3V;UMLCH59]).5B*&)02Q[W=8#0Q78
P/G#7&I+OVE3R+"A_WE2^;4S(T2EAEK4TMWG!HSK.PK\EUDT:%"1763RGJ49_/U0_
PXB*:?%R*5BLJ1$4MM[CJ>3F\EV8[L?N$ K"IC_:5W%FV/849=[5LGY'<;0L-EJ2*
PE+FT0;4Y58/8;^("O;7WJY/.CC>$BQ; UDN$#'7P]_.HO&0= ]1_  FHOH@CH8[4
PBTI<WUD/88TC)PKZBE;!'RT"R6\^#CR 4G<%@+W+ZA!%23=V#3T^Q7\&1"AOM=R9
P<7.0%M\E73/IXACHF-6I19ID;"A3XT$V?A3J^9KT;#7@B0<&A>+@1@LJ+_0.PZ1]
PJI=@3LZI6_!ED[A*X)A$Z7%8"MEU.-6W$>-VQY5EFR&43%I71Y?/IFJX>>&9 7<*
PS0?&Y%$7PZH >4WFEPAC*I^_(.KP6E31U%O(J7 KHL,D/65-^^,ZO:Z/ZIG*XV$J
P7\::\Y?OUE'N(W BP;@"I"&-#<Z.. U[VK -#88-+&B6D9R@&Y;6+^E^'P]@4[;,
P*W.)1![OMVAX*1BJ1UF%7"=Y?J9>SK(69.NPWV&@R^CRAT8JU(DFN3>?KXN8C0O)
P*<TN_]3O;B:FZO(VU7J?:<54*8OSY0!8IB2)HNQ67V26=Y(ZV+A1;<WP'%#=I2A2
PD0'\*C-W.CG)]+H;0.V*S>XP;G(*T(@#D.VML>G22-\\M"0IO]YYD7='2*# /1]Y
P.1II.K0T6LF\ 92#<?!A(?U+],BKE-U*R"TEO'0D9?\+%VF;F7*5G0[NF-? ZHL6
P=%\U/!9Y,\4RB^QT2*I.Q+  ,Y;@5<5@T&OL"1<J[=K85:FG>XPV.@4WL8%@U>LL
PK0EV0-K[2SVF6[(3=!KD.M7UQI&//,1FH*/X-W>ER>'+4!E6ZXMU)6:[3U!5RSHN
P]-Y@X(Q*00',U(@XOR(>OGF9" >13RS)-2I+4L,D\GPNY.L32T&*(4"/BCM%+>JC
P_-A"MK=S2#.8K#S]P_1#J1-Q+2PJ+\^BRJ/W7$BB6V!DL<X[L/ 9P+AX$LRZX&?@
PQ,P_*EG;]%A987L4*0@GCC]*15] \6F\!/K:A.O4"3S:CGZ;[3\OPA$3R\2.RT61
PB0?073MD \SR&0VDUXH.VQ-CE\,<[3Z$T)G$F1."C0+D2RMM'XTC&6/)1/@FKT6%
P/@QTV0ZE!SV9BL;F-Y,D;YSEK66V1C_5QV1P!)%H3"HK!"P.#^?F$-T14W8!W^CX
P0'@)5+VE]B!P]*"_%$./V40_*K]T^3RU72A__*T1!L_2CF=A0?K>QNQS]\AZX[D>
PR#K4M/]XLHF0Z9O356_?P._LG9]6-'?79("W&TW]*H%K+Z+9_3:5]!#=MJ<^E1U4
PUS\GS0"64$LK@P52[=)27'=7C!QNHXKLX3Y:<\)I-JY)]UZK+TB)XU["_(EOO(;X
P^2$/,#U=D**-XQO45_O[YCZ"645AZ<(SQWYQ3#FGR)B$R*'ZN+<.*.T'[8*7,SM7
PKP2IT<84M&(E/\JF^ZX94.P!O\]])16%%DR+X:KK"32ZO*4XV3<1WPQ<^3['BP8U
PMCDAJ+D7BM/>E"4!JH$IN7 40"065Q@2/5-^3^LU]5#6 _T.9XY\I1@T@G5.X3Q9
P/$&%IY7$XKG>'UK$6%GF5L5@3G/-:&</X?C)",K^](>7P:VS&8GP4'=,6&_ "]"4
PX_>O2CYOEZ&(=;;O4XHI-M++N)$"'%47:A?A$OB94 Y9%530$Q0*(# 37%V2=>*8
P',!5HD(Y+UL%9TFEC&Q&Z7,MO,XJV2D<$&#1NMFY(N9HO9_8!B)8[J[D)\IN=::D
P#U2M0X@U*JKUVF_QX1CTOSAE(Q[)':@SUN'FP#U@+VZ1%]< Q+;S@M(X30G/8=3B
P0CPW,2;KF>^E,OB;CQ%=4DLJV8"3M6W0D#/_H!^NH6*<PD^MJ=-FC\(2AO-3\0T_
P.!IW?#.XM(W]+C#UYGBQ8O65N:WTHAN/#0I34H:]58: MSXH!P +IRR+>YCE@+I 
PJ=_.XXC#4<9R\4BUO4&%/^A,;I^T"=3 ,8MG"@"#UBG0-*9TOGR'O;]!["SGQO71
P\Q%69_4A^:$C6-K5L:-.&_Y7 .3;T^P-+-4=>4$;T(/;TK .)R9*9V+OM@>6&(&5
P17%O8=CA6'70=CLDV4OSC#J^57K!#1EE&O,^2T"[Z+<2-U#  _A853AGK5XBG$*K
PY.K[^=+Q$6Z6-&U^L&L/^G?]2/[Y'9,#\55"7!:XR,RR67LHB-@O;6=2S9G1(U<H
PCLN#,O2"ZL<359/_!_U^1K?(IOBU X48$5^$MN7ZRCSQI3>T^3DJOBY^\9  (NWS
PY(1Z@W:90NR[2#Z(X?EO5K8C"V?V%.2(UN"[,J)/7V5FS_)TR'Z:-)62W?*17D=^
P[M>KM]LBC A=]OL%7[U3D("M>Z+-/9\R%92(S2**>U18P^Q:M9$72!ZYP]XGO4AA
PF[K =_IF*B\Y9-;4]_ >WL&O3@W+;X>.GO$?S1\1F$=5?B=RT[Q7U^N$"0<3J;BY
PIF+(A***I(+*&D[Q&YJI)]TB12*:)(-I)$1]6N_&-(?^@?4T@P/MZ/($06U5D3PI
PNDNT:Z'#XF"0(,_ZU]Z1__+' F11?H5&)"D2YL%7-XUK>XTD1]%\ST_<0$^[Q,!X
PVY+';,!6+P-1!YT1)4 ^: 1:8JO1K( ]CFE1_CG)%U>CA]L:]@[=7/'W2RV:7V/E
P=D-8.0!)PQUQ,JB8[I82SCIP:^3OMR*T:9TJB(3#?SG,[W)<"P@FYA_R03)[1(".
PBZ"GD,0K]J-&ZP)K^LOO3X3FX!K-L+A*@9:.U>-4=,*?1X$IK>._V!9>8"W M>1*
P[;=1"*/\EL!C@-"'^#/Z>>(B0&Y9C::1U&/5<8EF^Z._+X+C233% :Y;=/>()0-V
P"WH^!D&)*@R]TQS>.R5=?%!EY'O#9#(Y<+CP& P7^+)H=<N?CR8PE"20RJ05.&)I
POQH^XZ-VAGHALA8/[K8G)D7HQ)$5FEFPROP 6%.[<,KH=?'@6"WRJ&AI[:\\XG,X
P*][H.KPU:&5PN49/6>Z!"*\;4TO-(;JAK.-6-NLT  WQ2S0PBV<V/2,G7\"//%[_
P)GG]=$F'IIP.86,LUQ1"(%+B.&1X@)#))(!_1KA(MZ("\Q"L,_1(%P[1WO+RM_5]
PS*TSHPC-M\A5)!10D>[(\8V\==Y@S$[M*ULJ96*4__3:24$ETC^&$!R@/:JJQXXE
P4?8',&OO%.,E:5,D[1DWJBS/"V"?\XH5-,*L,XNEBQ;^%RU^=YW+=H'U74_@TB'Y
P Z$I>00U7./*[\DKR=X^L@RR7J^O<+G;9P^X7,QTD6C:G,U2VQZ(.48C!L('"*+K
P_$!:]*1&[_OI8C]![S3M:!)3Y^1P)8(W$@L/-=$Q *1R+S)9VWJ,I0U (M"$D?Z5
P$.N!N1?H!-PN*Z:>0A\8'S I47($4'>P1UGLOF%]3_\9<\585TG5:A.U?A *X\,)
PI11)+JY)U,>U6S857SA6VKI5N4M:3LL"LC4_*=' $+$QL35ILOM.BN?VPW%9:)ZH
PO7U-PU=;@9RT0<:)020"^9%*^A%'2+32Q'C[,8F615.D9S?#(>4WI\O/#YX:V> @
P3E^2[3I:I$^Y((EH!*_@TGY<1DZ'F>QWVZJBO.(LXR-TI:<TH"+ G)3)NP]+6#[%
P;ATV"9B^#2%#-,GP[0,"0!!=Y T[QH#- U'LD*/;3WMVZ'GI:4"OHU(E!BK'?5[P
PY%VP[DWYP0(DV3_'-WZ(EO.F_1YJEX@+V^KX:]T-ALT#+3T(?O.\D#7+X,\@6C/(
P<@:JL48!TZJ$2:MQT;J#V2IHVE&6$YH"V>JGXVA=)/G0C['[J"=!757FB_Y[OC%B
PWJF7HN>W?;<CF6\9)V8!^L_&:("'O\B_I $"IIL[-']/Z\//QS)SCB)&->/?N$-O
P^N!1R'<<1I;1%' ,?@,9C&%6ZVK0EGV64.MKA2YYE8_4YL=\2GB0D^_M%N^9+'E&
P!0I<&9)7;,2M5%,<&[-HDAIAP?UD@!B<>?4L'?Z2:9D*,*(J* W<39 9=MO6G?GK
P%<5H[OD1B:OA"MZ2I 7X9S?,['[\!>%E:BQ,L5/:2"8#TL(;T$(WY'.]IVZF923#
P$Z:LJ7MM'1^<RW<:\IG$5SQQ"4BV)3$G9X3M%@:K)UUQ6A,?EQ1&=&'.$, JJ'-F
PD;.P7O4Y&.DE('',%%013NW[T&U)>P].R#?P<S[AVY$]7NZHZI+   JS"2W9N(_)
P"/W@OS'RI>UG>S@@./13?F#K8.YA-*'8!VWUOKN634@V!N!BZXS/0L6DA2LA"^/&
PCW,3R\);SN<!1<ZC5H)L95)4C\);\A:%Y$L*G_9%6(V>Y(4G9'OE?.3Y 8M"">3)
P(7\L2J1#_!!312,0L:/GA1R)\WY89@76)4"/'2]7@ZO,K-XN7[IY/]0N_@0M;=(@
PO_3LH<*)6NAMR92-S:KB;Z_=8.AM+2G9:5M[N_&(5M)*YN % 3PV:ZX&LR9*0+&J
PO3-EGU+6@M6V"KHB74KK=8!)#,'N&25*MG=6_EVHL%Z1#=VFB"WPUZV$S]&KPYUW
PP3O8/BX/P+RL37XC_'?5CSA]?Q.37^4G%K)""H]BC0UWCEK,(95BU_BD6W%+:NE 
PMU XO <AL$:XM;7D>7HT(\C\LV7-SN4:XWHL:G:UOY*@OOB0JWE_^#B-5CN</3NT
P)VNS$_""%[R)]+]MW8OZ4GD%0P%/-L)MJ/;7LN@/:@_KU"P.#& R'5^*4REWJ@U/
PV;54F6[K6H)/+U96\-QS)!>UBXBGA1U))YGV7YHJCT]NP()@^J#5F0SO\9[!V?->
P.Q/D7=8Q=E]G"#IYQ+Z/*=^*\MR8X4'5XQ0]82@_O]<18R+!/,"BW>4D)Z8J;=O!
P>7ORWU J(=C5-ZB+-V"V J5[Y^1NK;SAP4^L,T'J<E+68)(RL<)AC]Y[05)LU\%Z
P150U/]P8,7J(:0]BUH7FS4E)I22AB!7YCH&&$B#'(=B07&F/%K*J5W'(DR1B;\SE
P8J(S-ZO88#4SL'70L_?T<< Z?' ?:@KV]3<[B8UAVJB$Z[62F>B 3[W$C8-<A[$=
PX M*Z'O23_ .$7 G.1Z."V>\D7P)@+,/+QDY59/8,<%F<_JH[E(0>#QIDN]3B9,D
P6&#8?$5@+"H,4+.X R,=.^!DQY'R9_3WX4AXCJH)%"J\9*RI)MIWF(N2#P8\[BQ7
P-Z#42=TW"(HX\&;$@#'A2(OK3X7LGD>C!JF3NQC^-[3M5%#$,H5OU4'6\@0??#$-
P$'Q&%>P+YR4S*S:M7';RR!"U#2&MC4!SPYK"G2TN[)N(X,^X2O3W@FC$]Y[YXV1?
PWE-\H[>;K]>&V+F:SI;17K.&D+J0#\_P1$2^T]_>%[CD(E/<-.U9;I5V7OX6>!HZ
P&G18_U%B+0:N^+3.^&$QBO5+TDJ^T.[NI+(DMIIF6ZY#%U*>E"T?L?^.U\A:6"?J
PD)7M^C6B#NN.C+-;R/J,QUC[F+!LG,T1K+L,5SMW:!*<KKG#)1'SW41H:QT41]^K
PB"]SE>]HS3ZAI=[6B/6,F,=1MYA .,X!C7^?=BS4J3RHJ!EGP_^7>.0U\FKSV2]\
P@Z0IH[Z9MJXIE$/I +!!/SL?[,C[3C\,G=5Q3B=U=%,*I$J[4<1@IZD5!O$.)W>3
P$XZ"'S,4\,49M3JC.6/*UO!#8%+"5XJ4D8?2[<7G,.28>PAN"U>"+(8W=+=%Z3QL
PQ3RI[++O5!4\*I+4"Y6^G24/RP>URG@'A/0[Z:4/Z*O;BNL8DAX^ND9:^HE%+B-[
P B-B%5P)YGV93,5?//BVWOW@%"TO?\(=",7E] $JHI",I6 [@@:OCUO;_]18MBJN
PJ;N&3^OT*L"6."=+Q04@%\]>GM+WX:<C#.HD#'\27+R4>+>&!!>V?M&(*])!NYTF
P@7?#T4^K&?9/>[?1?N#W)QCDS[C3VZ*<<;?V&]5,E@7@O<)2&7*FY03C[-44_7Y.
P$47LV7!M3UOS.SVH1?)(6M3ONB\/=;F@[+IYN0715!6(*=B3:7;=LYRVH"J;8%<Q
PAUAC<*#3C%7$.!W^H@2NO4=O*<ZD[&!*04LLU_@U,@RYFRH-"\TM9$,+$=TJ&HF&
PUGYD>F ]6#G\O8I5-&>87)U4&XB]KNN06ZR^2.J:N1VC,S#BCHJZ7$Y[;'\H'(NI
PY2G8M=HAV7]-,&[QS&$MWX?,O;VAWEL2W?TF<+(W&@^C251QK9U19OG<ERZ\EBG9
P!5DSN[[B=G->$DYM34M[=7+'VSUM&$[Z#V'K\_1RZ9P"R?PE5EF)W2P# ZGV.QQ0
PT^.1*2[ETW /W"-]<W=-N?E$_2K^)=,KC]PMBK$59 92X7EB9%]BW@UO6PG:U3$+
P@? 1WN 'YN!O".EI<D!<"26+OCI1,A\M5# "=/\MC5D!#'K AU3?NU"#.7.]/YM7
P" G_'-)W6W1[?%AU8L))P"HKA,!092OXT.-"6E7["+[G,CCKQY:TTLI_M/S$?:>5
P( V*=B9 Q.C-D/O8,:O8UJ"J+L<Y)IF6]CI!5D49VKK]FQ<7UB1Q47/GMFXADJB>
PW/"<Y#BY;JU-WFU;GT.V)NQE5V6?3Y$0W3]!L;03M<9;D/ZQ_VP6IVS:31.)@B@H
PY8EP5',310T[))(/]J''/PJR_[=4:1&ZI?=1[.5EFB]@[[GE6T@A%E'=K$#6\+W 
P[?VP2J)J94=HKD+:C>G!I"$01@#$9);R$_![IN&-BKW1U#=]Y2 C7N*D#(,@T6\I
P37-(?<<.TI@M-MB-VTT!P Y LV9>.\;0-E=,$0:NH>I []DY^',5*Y:3"VK=_QN!
P$AX^N[^W6=Q(\+K>WBCIW(G.3;G)^)311G1Y,8<">\B*7P8/.DR;E-4 K?M]M-%E
PMQCHVG[-&F>%KO;_;5D75:$LW7+27?M!<BDUZV$5(SWY9'$( (>3#:7'5[0P0,N$
PZ>?\ .F$> Z2=^L4P6/Y?TN+;!S1:0>[XB'M[ &6[ *YN["#;\9RN+X#8Q4B5NG*
PY(C[753,G25.J'F\F5!T@^]"^]'YP5/[[T;O8?7+9[?MOI<JVJD_DQ%"$]TU6E.#
PF']#H;[H/!0FI\=Y-P9CO5M.NI :%.%8V$< *?WC)94QT?SF/WC8EK7]#!HE3?",
PMKAHN]^AY)IFHF(6GT+PR?%(>TTMJ@NIT%IAZ0M(=-!-ML/W:ESBY><RN#<F$@O@
P.-M4!/5UO;<WOUO]K!PZM[%#9O;6-CJCE'VE5T0>+R34T(*M%!1QN^EH:^QR#>@@
PIW(+Y7,OD%<*K=+$OL">&5ES*\S90MRJ[6,S>XPN:<<;,>\-'\+1]XMQ0HNI!,%Y
POS/K>^[<=C?2R6R3H2749_5W7 O^A2YNHSP:39M<.G4.D^>. VRT)22M?V%$V(F/
P+?%-D^]_T<\1]>'#'PT2VV<MB3(]QP"G"J6O^F2;8"NS-^ ZAVK]I!%-IJ0H70+ 
P ;^MYQP*_^GZX/),KGG<=9O)]QTCFES5YHDS]CD+_RDHQZW;Z4-3'==7S=RHFD5I
PCGQ0*' 1FS#2Y2GD@+"R&=2LA(GR"BVO2+H,BSBE!;UZ=ZJ*9W,I03I[\;.M/Q E
P//U"SX-X@MF;*%I3K5^*!>V"@;K)M"Q\C(%(](-?Z92D8_M#&S0L&$I$Q<#2\L+X
PC<%086BW<3Q[)R33S#SS?>F<C\Y)K!KQGJ&>$O>#^8;O19=GDD)X0^JS($XIH/TL
PX1+D>7RD^4-,:JR+X@54Q=]SN_;_ XJ'5.0O;P$(;QO/PY7B_LQT+OXHWJI[!#1$
P5H_\W1R K;_9D?#BFHT2W-&5Y\.JX+1TX P3O_4OKV?FI/+)&B:^3_<*Q,?KCY[$
PHN:<+"\!0#LU,AN:O8-[7ME>65_>Y05T^W.IP+ELJUAJFH_^J]@@[2]A+@,Y7O!W
P_K%E%) 5$:@3--NJ=\5_CT.[<@X]IT_@LI:$*'(+=NIG@LF#^B+\S)U]_YJFG*!9
PQ^IV[G8_SWT=59JU>R1HU<EJ6-.+S=;UY?@O?< KBMFR+&IX$I&!I#J(P-I+2K),
PBU8'0#72]!X? IF>(HTMUJOLTZ#2C>E8(K:G:F+EYF4Y<L.UK-<P!]-QL_C_4%.+
PL>9CQ^# ]C+E7%3:U<]JJG?4286V"+(2ZG%;&WV[T;HT$J_4JZ_+X089]NOK#O2Z
PBMH]*#0YS/&.  V!F<K!"">[FSQ5G]*U\CG<>?'_<;F7?XE263GYC<?LM5("5$I6
PBQ9*+"8BSJDF+1:_O3V 4*5$"[X"42VX=$O_P"!3#03"!SZH8$X[?@I&R6]D4 ]3
P66B5T1=X!?B>!EZE>SY.O*?1 !4D?S>^4[HQY7RU=V;H9L&DQ1R\E)++XB_::UGO
P%IM. BZ[W&1N6B/F\'"3*39S@H*-'U'2U"HD7APF*MT",<KB=[$P?DKD/[9?[<K*
PU :T:10F6^HI#25XY"#!CZN=/0$'ER^#&Q$MC7+M(H/T./G>H);[] R3^*>KBW^\
P!=C# QH(+!.>'.U'S?PW81!?)>RG:8<O8D+ZCY6G+;@W0<E*-/5WC(T]MEAUAEP&
PRA1V=,:4S490<F@H_9D/?0RLP>8-DY1H3QY]W3"PK2>+N=.FK+^?GK[JUJ_\2$B;
P8,.,XJQF\T&W\1D2DM!93)5?"5($UOYZ[YD6= M629..8D]]>H'%[@VEVW&6YETL
PT?%&IR3*#:[TR7]I;J0,F1]TS-=HN<-X/A'*13MT8-9'^/609GHI[>ZU:/V-V+G8
P20)(92,D'''^26&N3E1"%/>F*HVE8X\I:5B/6+-8E$*->$LY6\%ZGZ-T;+9#2M!_
PIYG(:7B7AJ,"?'$2("3"D-,6_>EV:J =MYHQ*C/M&^I,Z6CUE.Y&&5]S9TEX6-J'
P'E=97%+$KS^3FM[-'[J/6=^6!!$4 T1UB4,R(PUE06SA:I>_&FH);A!-= =P@Y!M
P0P-W#W)BLE+;J"SOAE]PXE)HT@)M)KB2^6'.?T>I2B;J9S,XEA7.ILE+CM#3=A=>
PV<X BB2^+MIWLT^+#N,3QOM"G2!0>SR8[D\8]5> +[0:ST00!A=6NGM>K-*LB6GK
P825IQ-<2T)-#FZP74>5#DN6K36$XSZRPUOL@^T;_6,%LF+TAK=1Z9I*C#E5C(--7
P$0N%P1T+C0W';I&(4$CD$'POPX/U<TMOD;\&]X_)MXT=0ET1JNQAOAV3/W=48J[%
P/#=[^, EH -S]$@.4V=>TC5975CR1C0B8T.&!<IYEP/P:SN>WW43YY[L&&4^[L73
PE9"YI8GT+X:Y,G[CQ(NO1Q\)L?R.YG]G])OG-@$9TI6%*4J(+I\(E6&]+\IZI+$ 
P@&\^D>)08#YR%X!-$Q,XN].R#C1'T$I1_\T<RZD:+V)^9,W-D;XZ2ACZW X-.^ V
PA!H6?7KR-T@#IS&;9<@"",U#&.34RTTVD>;OKG*8;Y\ 2KEL[B&B_>.:B(PN^)D=
P+G%<LDGVTLP)%YY8CUTA@(MA5YF5]B!/J)MH(;8W"8$^YP//\H>>TH:58\)><]0A
P>]!KU!X3JQ;&$N[X ,@<_>&<\YU,_TB!@*Y?XI?FW7J:__W6;L>2E6II'\8M41$1
P@FD8P)?H-_RO#89$B9/VD)90QRWE (#V-ITX?BK)!?+@D\3 [>JLR/^4W/<4>2PN
P.8#9/J=U?$C&A<>!%:TQ'F@%]U?K_EYLAR"7FAV@A/^=;M SFD:OO_[:Z\_<DO\2
P',\I [#KV^D!?/3FX@B%4D*86^F9V.##6V*A-04H'\VWG?+L9UM[_:1CXPQ(%_&0
P&+2-YEYLN[9;]+&5&V1G42K]=PP+,*RI[ZJPNSPGOZR(VL)PN+=Y"G4<@@C7]4[8
P@YB,!(&(9"34T_;.<)\]U^ KU6&@WL,D%S )D!!@1!M\&:,S#FOCJM/=#,#:Q[MZ
P#OK_?@PE*0SINM%"^:GCR\:&I'A"KW[KMTRB;)5U[=F2V_>WS:-CXX#GXB9-5C\D
PH0OQAT?4;C.+S?2[5/#JPP*G,99C^+C/GX=;KQ881#A'ZYE.%&VI@T;YJS\*5IR2
P+'PZE8+HU)*^!)HYO@OC,ASH)=!8<P$?"H,KCR5^]JE7/M7C-> XAV,!9/:4%0;N
P-K4QJ8-\*>((JFT^L<%!%B/;Q'=SI3R49A>'7Q<@.E6:3Q<1J:#H@RL!4@T[/3H+
P5,(R>H^$6R1M%"6.F[$.U3ROMNO:#XH@9I'U<*._1('C+91)>6C)UGZIM[V:5A X
P3(%6H&:)M2$DWL@M9WG16SD%:A044 [@Z-_Y\@H M="\].:T-62#ASYQ^C'@[W]R
PMS17>I>J"D[=+N1-"7RD55S&&CE&IA]&9FX#1JGH,[P_8K*W4L9(<AXMPQ=(D4J0
PGUZC1B_9Z]Q)R)$@IW[:;--9,B(7W5A_#C8CPQY6;HDUXU$W(NPU87=J&'WF*J\>
PV9RPQT S5Q5F7#9T^%G1B*3XS;&:2>Z@L-!1BI'ARZ/@R8>H[LRJ.>&A1::[BOGF
P(C@&LFH*I_<UL*%*"=K[,"*W4KGW/+#)+?4<Q,(BO KH/JH$JVB=GC/GQ9(!J^9R
PM7X=JZ3B N051 JOCX7;VUVM"O]:)D(EN0[R'*\"]E26&T(X6HS3]FVG:3YKE1M(
P;15#_I'YO)<4@G62R)MY=J+DR2 '$HL*@B4EOCK.>[]X:QO>J#HTG,A1#M'FH$[ 
PJDIC>GO"* 4I._@&R,>=+V9YPC] [MQXSS-C;%JSP-CN'?P=/!-E#6Z/E#<(035I
P?B/N6X'IIG/D=$SW6U[GEGC%@I/W"Z1PKF;5I@$$I1=9-;DZ0UN1E([\LK]03]P!
P"FNT/DYQ^@3!GHMEE8\Y9\!-@.@#P:U5,>&J]+!Y%P/0^&F=G7 F6OLM$?9:TZ$D
P'8 6>/:3^\:/4ZD9CDZ&DB9YREK0.N8<Q14-=_\!4%CJSQ@V,*!GPB\:6MB7\_53
P"5K4-V=\;ISTR#NR5Q^/B.SNOSRX (@-BO7:JEBZ+9@X_SS"8^S-E'N.P+.C_!;X
PTDRW3O;QXE&MXH$KHU@[@K <(4==](5N9X50@E7.%8_R'YZ%0OO6Y2$T9OFZX&(=
P<8AQ\5Y2_X!#E^J#I@&-XC)>NC[87_NOD?'@470,_C@E1DO=S!_L&O:M\):+ XNZ
PX1=/+P)+X@$TPJ4!21\\]?K$V@&;/(#ZG0_/J4!A523= 3FN* G\I([;&)B+W(=\
P6VEZVK#]A]1)LVX+*MWU'L+)0<T-R:\8%S3I)$1)/7=$!FVUY^0*'B/6+>HH!=?K
P%1:H3X,!WM/RF]BA<C:-,SE+^WS?],=SA$[G=&Y A980U1;QHUC9#9Y;R=]SW? Z
P_&>=3W\"VJTI<Z-.I Z:7MXF<3),\"?[2%JA%<>N*.@J>?EB9"2(N*IGYZK?GK!F
P.Y7)$!ZB7H&%2J(8@W7^AR=:2X]-8[O\?#0&RQ=KW7P\$VTO@0P+?M*GZ%4K0KW1
P47N9.*D<CJSR<Z\H^(WL$+7@Z@(U_J)D?G^42#P8R\.>\Z2Y[C+Y.6U)4EF/$K(*
P1OHLPD* #\SO@<0D_]Y2OU!<=B-TH^Z"AQ&B,;HM'R"8D=G3QG:((8H+MID%AV"*
P89J-=1OD_4LK/-4![/LXI2G"GR"%'[:+DMDK"#_W!CY:+E*E^E4XU $%K"UO*T0E
P7Y<FT<$!#6ZP>U\<S+URCV25=6^(+H@L7[F)-W&Q!(SZW@W)Z)>090*?9P]#0BY+
PRIQ%0,I'2-DN'=[JPO#92L<H6NXI]M#?->B#]7/1XH\Y89WM ][5YZB(DIJ:+O\ 
P_>YVO&E9HC#0I] -IJ9;^>Q][/WF/>Y/ +9LWGY-,+$,6P4KY"&(7!M9 YOO!H;M
PY9C5"=59YZ;VW'C]&FB)LYNJ/ U<J@U5>P'5,.E<4)#".,/=-?&VIX@ .)8MBFDQ
P_)>N IP7A4S>?;?\(]K_S"&"__0?]WNQ']%D-3G'CM-S7WE><X3QX;NK]6+M@.;+
P4\%N>_0#[WZO"JJ& XH.5KJ+6[ TZJ8?.C\"I$HN"Y'>0*[D$<\8^;W9 (SOV;]*
P11O$4S_;!;$1/L0HO.5Z#ZZHDW/]S(1S>N<ZVAHN56^'AGW7<OI1CD7,9S)"(]N\
PH&*JPAE%QNS'"Q[9I-QCSBR&SY1SVT<AF:UJPFA]N1($-T3L3M _/!S>$WS;OC!2
PQ,=ER^)K>XIUG>P$L)U],SVA=V<>$-=8]AK@X:XR"4\5I&7 G['U%*DF_AA9"@=*
PJ*_-C&.3<VRVAA:-8+"*72"D*_Z;-T'5^<?D7/H+JNL@"<#.^4CMXS_(C:;"K;NM
P_$>Y\38+@MQ9 TQ5/FDR838BS>2CSO>K])9Z$8I:A;9V&Z$D1&J>&%S0+R&9(P+D
P)K'$">OFLOS5A;*.&"=5)@7;KRLOIW[__)!0957!$L9O2MU0(P?X;$7?\M]>Z 73
PM7$((6Z6F#N("#S:JT0A U_<PA_VOKX]1_;.#)57?\=#5*M1A*M;;X;Z$37X2'[D
PX_9-C'--;E=SUU1\#;25L\0%NHYO8J"5XK\.$RNU->NB8PR"'U*&,1AJ7_OBFTK"
P6H:=[K1H,R1'O[4&!-L=/ZBMLCRJBL=07Q9C/T8 E?;H_X]H3TB+ O(&7"9WUM&Y
P85QX])5[BEAU@O?S MJ-RX_$A-=K]%^=_;OIRPL,'1C%N]@K!=E+?3 V0V, EE:)
PX4?W]:D,DLUYCU@5IE6B)#[BROQ<<4 A#*XZ#&53CUJEH,V;DZG@J6* W+K&V-,H
P$/;.G>WO%[G[1*LVO%5Q*C.)3-R5GK5:,6)JC#$^S]1+=,G[F+/X&6?HQ0^(7*NT
PIO>*QD2L>.MI">0C>"1JYE6*QO-X!<[<NJXOZN)-SYL3(;B6AG:#E(X_8X;2;I[9
PPBD&L67Y\;<Z<HUK$M]FOTU<M%$!K??HB^&,X/7*3F##?R;L:=LCN?9J!2[Y8Q N
P(3[ YSQME.XZI$F"$]GT*AIMMO8$/R58X\GV*)]_1H\+J1=.NUFD@D:Z!WN;NST+
P2ZBQ+.#7F)^!),)G6Y^XL9A".AS!(H'QO":0-^1-9)M\<4:\$7BB+"'YXA:Y2W:9
P?Z(G1#D?E%0\NUVN8LWKM!K^YU3MIVI0Q0>UH,[6]?PI6MULS\E:,//^@Y]5J^2'
PVOW&/<Q&I5D,#WB27%X:=V[M"8-;'>*GT=$"),TI[*P4SFTV4A:2U?:&_LW#G )9
P]^Z!O%U>W@7^O)%BUH,'(4*M,AGA+T2IRQX_1.M/BS;Y[OL#]\0M83B@!>G<^R(H
P1E?GD,A"($VC):A9S G5^]ML638Z7YIO+#N-"+IEHA$MQLY)5IV<=+$!"[2\9>TO
P6Y]-XJ1FCH,G/CHTTFU];FK\=<&URM2%KWZY9E'&4P_NLX=2Q,-.18NU &GIFS),
PUS\%8Y217O#PD"$JAZ\[H&/*\I3#*@DA#=0,S<"Z0U#+Q'SC*#:YY/4VM_X\66I=
P6;H&IEA!/E@"W_;F9I/3/0 '36L0;^,Z/_RH@KIIZ[J9R4+.1Q1%)2@-@4+BZ ]P
P@C0 (<^3:@H=^N"G(S*M^@07!E5>/DF6($8(:]G(*BNJ50 4Z'2?5?+ >21WX>2W
PN.6M'RX',"^>FE.@!*2WK:D_&#5KM0O! <6!3)]^^@4U*8;^GQ_GW%."F3KZC0[9
P-\4$1C^+AG+2IG*P?D;7TU25[+9/TKQE7^('\=3K[G4CB8K2JSM&X6=W7R(\4)Z'
PLG<&PA3W;>40!]K1=*S- 'B2!X&?63N$X-FAX>LZ":,2^NC^8"8>8]-XGS#5N.+:
PCIN9<%@1'J#9-&)']?7-LJ0P_%Z7T8$W<K001FHX7CRR8AD<._(&\S.0UNI5(![!
PBM]Z7#&7=]/EX-<II;J6>T.A%NP@[W*IHDR?2\]6?:9K[%)C86XBN*]A#&62>&CF
P4ROVQHCF366 WYJ9O@ LQTPM7P@9^C3;TWW"K.E5H"A/ 8 *8&^O],=NUA1<O+R:
PI?TQ<4+/JUX?I4IC), 0CT@IPJ*PF;>;[">-XKCPZ8*ZPQ4%7U&^S-%TJS2EJ7'H
P2OVLI[>-UL8G\0)F:;Y9IH&56D/>,D%MGHP/</TY1HIV[)Y'0T #LIOT](F25HH>
P43O"+2H5#AAI60!@V$(T)RE8/68"1D&N9&V7V?%0P3N  #A(EG)VT=6<F[O 'IA,
P!*_SD\%!*S3?E=GJ3[;R41SD8#5LZ4JL&$XT$5HBYNG&XDN8Z/J!U8L/ _5)EX6Z
PC"A&U<P@>;"!@4^,SH3[OK\QXS4>3%+N_CKIQ05%I"V.7GIO1 Q.OMI]R)#E+\;8
PUW-F<ZT?:(:81Z$,ZX_(5IC(4ZP?#YB$SLN5**1P-X+FZL8*G[!1ZW6,;1VU<("G
P*!.L:1DPP[78CHEC/&P?N,^.LU]3/_J&D\]J8'&HA=[NFC-E<FR?Y@R.0$DL.@L_
PAE"@P$;-_1W"X3ON'1U^$#6&0UE:5-'_%L< @OH7HIP--?FUCTBYR[101A-'CUJ9
P >O+/R;N@+:*BD5/^'2C:8=(6-/=R(#;W0D 15\2VV!6>DVW86G\MU65ZT; !:9S
P*(7&=<1\9OIC)Z8K</04N')UM$?6%OKE#S2$MBR[W_/6?!,QMP!)(,$\LD9F)=Z;
P4((ZU?LC$0;KJ/E_&J,;JS'5+\VC6!]V).J6T>'?ID'%?QDS3$^'7W)(5%%HJ,AV
P#;E;+NAP"7N]=KM],&;D7K;\;&-D2"RI!1!W&"JMJ!<H1U!YEZ7IX5YT/4;SGTIW
PQJ4X*DD\E_(:*Q]P  8TC^O1D'L+(?IE&9MQS/^P;#":0U([MY7"<L3*)B-%6>0#
P^+[@BD_X!6:-8.37,>?6A94*^83V]@4P%&2@N<)SOSM5EA;JJJ=>'V_U01-6]C\H
P (-B-P"*.(+F[QX0T==IC;!%P3!^>;$#AJUIY,?H"4?(XYXB^/TJRYTE_K*(AJ;8
P Q=$,$O@U-B&#'^ETOX\9_7[<QD='VE@3%,?&* ^WD24;G2)%X58@'WS4)5&,,PA
P&J3S>:5\YQZR MAB.M/^H[W[U'L9<J>(:#),3,7K9X)(Y(R!7D$?O/$/Q&I0P&+0
PY1\''EA/J9.[V.L.[M(S 8X7X) 362NH:]1\V^(7R]#&'PE2CSB6DD4($0VQ/;)W
PU\+ .NH#G S>A;Z7O=I?I+*>#G:NC_-4&#+V8LG_#D9>MK8[L(%RC:G0\JAYER:I
P_'):-OMKB;N:]XJ!]YE)6AZ4,^:)I08_M50SV<F.B;+_4\ 3J#6>E^!7QA*;?1Q_
PM5AB+B/Z26+?+@P:"-UA39=%VU.%@.7N*>&2]@+\&E>%K]XVIC-[MID\'DIG/9!A
P&Q*#RE\DC;:Q\+EIZB9R %W"R_@\C*GBAGBXLA9I.5$R/=L3PC!P\93K\#6Z@,Z7
PT\YE]RSX[.0[#:5@X;/C-?) YA$"]8J&"13^I&,3W^I\&$C@[\KQ_+/P\BS%-BR(
P<0RM2/@XLYM50RSZ-#/$%]I\$QIMJJ_^2S;W'P84RI:-IN@Y>^B:D"9S84\"KR\-
P9LC6 Z^1AVL+(E&V>)37$46FXS8BL?D ^'?M.\F<ZX'\K>Z\_X)PC3OQQ$@4Q:6G
PO@,S77VG:!ZTO%5M/-9?_%H5JJ^WC_\'OOQ=:_.=KO?^-?]>DNG]D\B!IZ%_:5_K
P0=+>JZ5T$IS8@A U(%12ST>!T]CH,%PBX%%K7+_.YQ(XKH%2&<]83;ELG[<1[:7(
P*7!"BV3[/Y:EMRYN9F<8(U'H0T,GI97&_*L]5LYEF).5@,K'F1G?O/G/RDBR$ "<
PH>DIS7+P IRB%NYKB&UXTFDNFBZ(HS)"C8 B#[FYD7OWRV6%>87M)=#M<_,N;[\'
P,\J  _^_Q ]57ZM<(LTNBZ2';VLP.6-^1^QRLJT/&A)4NS>3?#ML8'P=,I\4B7PH
P"N;NX3; I*03+#B>C$021%^3@66(U0F<<D)1K?=M&$:D(:VI+59HK66:\#TS[I4D
PY8DZ,+EP.'F">D_1%ES!@NP):VA24]"BKH05=T$M0M SOM62Z2@C-\%8[<R;\W%+
PBO 9@@(\__/N<2(3&W"7Z/X>(K67]3IZ>X'\&YX 4=.3=+5""AFD7:(.[7]'B>C\
P!EO1&\!EG(RN)OUR!6M6GQX/MQQ*3:\V1)_U^G^>#;)"GZ&<OG\*-I&=_YZ[OWCM
P@\<$@GLHOPK@T!8'+\S,_IL>M4Z\(N"RRKV>./V)5[K?/K5ZC==DPL&*^#"4,EY7
PHSH:R!2Y?_^WBF,!V<^E9!D_^^#3:S,Z%O'%Y[I6!FKSO/[:QJ5034/">_[@[H,7
P,A)9(-&_DT6VHKO*[X!^>2FX3_NG<MU/&[X<TXQ%3>K>Z\<QG8KMW>FSF-IX%5,&
P::)C(RZI\>SMWYU61XY:R5;?]=_YB2Z=+ZPNWL<EJIR7$P ?7(OFT'3GSQ;,UNNA
PSW#DG^#-%Y@N-+:X.?[$'=:WQ7%T8'<L,GLR0'R<9K.K@2^5RVET+MX\*J#B*ZQJ
P^X(^NH%("(J'UBM-!39'&GXY"O.;Z (]NJKN?F0<WYP> -YVBEEAV6B /EZ"EOS4
PR[#M /C:W^R'TFG%>C)KOR.RN9U%9O>&:$$N/@[EA#$L 80-\XF=BX]X#$BIKQOK
P.32"@;H2_<,M,:6N[UBU)Y% 6,WIW-QLPN=IVLGPR^(2*T4M/V>!V@&HB49TZX%J
PR%BDN:,\RNCHAY5V+LB+X[I7FQ(A;^E;5\LKY)B.A1AGO,@?3A=2/K6RT1W2_H#1
P:G^/-X(! 0@,A4IN2E]#G=<K> 5USN;_&=Z""!2SS+I"!8ET7\U*1P=L=J$2H2-K
P?3[?R!JZ.L>P&3=Q&W7)'#";!ME=]L8,B_:DBS--$L2.AB7ZX:C;->RY,>+*.H7V
PSL,!Y:>KN()S9"L!M)W%G>NC##W&@T'/NT>O/V/6B;3RLGN3".^/#%9%Q$B^+_7^
P\R1];Z#W*]6!%OP@P&DRJ[%!"@'YTL*^C+9=\!!]D[84N\4L8\[^)H&G<.P<AJE8
P8\MA H>C+2_4'GF@RGBH(-^<8;_.]^R#+>]L(]6B[IK)+F&[[W6@<GY%%"J7?H<^
P\20YAKJ!,2_[.@[F\#A>^PGO%@EP8%)S J8SA&P42J3L_#@O?!_"+.A'67A)?$@9
P2Y?^W1X?9;$FOL25VC2>#<LV&(^)\7J3=@T8>W9)1$98!BFJ(LZ%G0QL@2PT,U3/
P:;<>M,G+0A.J>$#T4#C@$QD<Q]"Y;_#\@3RC7IA*Z^BG/XE 0+$!CDWBAU537>\$
PZ2@ZUJGDQTE!+[URK8D6HI)H1YP@?[1*('<;<@"ML6*D>@N-!-B7QEH1E<WA053O
PPH !-0PW5LT5_<GT\*#V#SE50$%\*[OV6X!JE<'C+_SNM+0-_#[OEC 0Q71Y97$?
P^FXM&L39L*<G<^?VLT7U-1X_;;B"6Q(MW;O "6/ZQ6,Y2G06 &%'Q-Y R_^9>',N
P#>$";T+KTM"[43UV9<!,KCV&,(#D;"\HIU\.G7LV;.OH).  _9 W:#.\QK$AY[R;
P21YNRLIZ <[7#: &CB31I)YX76_0X)UA\8HIT9Z%TF\!9&,(OAQA]BX F/@>AZGQ
PRVY];YUK">969^G6MGD]. 0&)Z)',@T4'"C7_YK)XZW@]C'!TBP2C?+W-\=/,W<I
PE,09W@9,7=V0Q<8*-A[X6^B?)A$"0OA'B*NKQ\\CP3\!@1Z:UZ?+9*N\5.F^\%<R
P)!I:XQYOK5# <1:US9E7;$GBE!O,R=BMSZ5?8XJS!&?F+5;Q=C&O/N/DR&T:W>UC
P/<&9>0UQ_@_4]!*(L0J"Y.%2'?VKD?9XUK6=),.M1D"%8B2#Q:A:36[Q7C#FEQKY
PN,/0R<Y\\0U]E=I%NBH,M!#D_BG:,IA_J)CJU!:VL-=[/.O%7&<#3ME*,.+RA Y8
P3@W"F'=S_>Z*O7DBNG)*,P-X?W$8D@VM^V&YBK&CF\:>9WJZ@0=-X5D!6FPC 'V)
PUM#0GHV)I;ZOD.75X(.>;NI-D0$;T:[$5.\-8UF4=0_%%;*%C,"TS5O,Q/L! .%\
P]5,75!/88V"VI,8?$/;.GK4S;-=,R"F33%JBSGA^4J*"FWCQ,[?4+&YB) ;ZO3CT
P#SKTM:'@)\*'.'@OH%<7I>^XUDYBT#D&9CVUHV_75 \:)^H$NDQQ2'N(. V*8J,B
P8A-D:4<QQKC@-/+/]DVF:0%I?JVI>IQ3 )<8$)5DI=.S@1.Z+8ME=V!/7$V3ZV@"
P#\39:@$#W7<E_KZ/''VM/I<]6N/1TST^,!P/P=W<+2]FJ>R8S>!<A>^0*4C^6)48
PH]?.5JA=S_2,_B#;8=P(>A*U*>KFCB^:]-4FJ'BB.<SUD_DM+R0FS?<Y8I'Q8.\V
P"F+^UAT136]]::9L4SNK5U4$>H)>!( !];2<$&W/CFB?,R="$FV6!S]*2S;H$7ZI
PMC%X-*G'XL&@7Z^&,IY-2^N&3[^!+S"IJ%+NX7MSLRBD&TJ;7>3T( "!%4>FT%:X
PI^I\P#$'%DL+IDH49#?+R"DJS)0J9ICKMQ2$=W4<Q=%CYW3.U1\_0QY\>1PWI5_Q
PXV/&WR@ZSNJ#1Y>[.*MW%@_\>1;2"V2[ZDW(@I-Y.$E+LB0](-DOIY.#P@%0M\)0
P],@BP[7'1_*SDRU]EIZ\1+ULP84E@Y&G,_/\%P^*S#= AQ..8T]\<Y^J&OU$+H/#
P4O],:IT,S/K:6\:0SDFIY<_XK&4>]R8="T:[4"$H?_MXOV)&2Z$^S !=&58;)A-J
P3S9P H::*!M#H9%86UD(D$9_-.T^SX(8])+/O<YH^7=3AC2;B%HXY<>V]HI52T)*
P -;?-*AXX/%] "H(34!4/JDJ6U >V;=V,_B%17<U#13O3C=-H(Q.)7-K:%#T41A_
P;UJ?KL:_]I+WNHH&9-UKM//-'X)5PAXPEEO0@U#O*HR&?3SB!&<F.B(K5GE(\"TE
PS&=/M) !6>H74@=B@PO3<&L&O/]=*QZFUX3C> _5\11+>M [XV-3OE[(YD2':4M6
PVTC+4MXB"1L1:B5D>3''$W8<W_F\)(D3*!+J7TRZ6KOQ=--48JI65@&RHXIQ=L%%
P*W_8M!N'2H'W.!/NC,.)>E"!V2XT1(:S*#WCHW>X&S9#F[!DOR<EXI_!9Q/VT#G!
PHFT27+6A'!B:JJN6XX#R6_VW]\EL%@Q8D-UFXEF+A!)9IQ^K"TI-O@S8]*WC1#,$
PP+)L)!T!;OALPZCOTT9<K9J&]8,4L#7 2W1ODP^8;X: "_I\_2"!@@$,NU %5)X7
PJ6W>P0?$K+ZS/JAYFEFJ?\>(ECJU."5(G'1/I\,>(:-5G<N>-NN@:UAGQ[@#TE7I
P]%K)H/!T-#K"B-= F/7GRQJ+IEVBX88/4BDI"@^4'-D$&V\9USTX]'S+F^=]?I_S
P7Z"X@N[%I.Q,%#N8'^0GU1:B)S#1MW )Y^O9S/O+5%;38N!TN]XA,ANMYJ:V7_&0
PSB<7#7C,;JI59&&B W!WF9QU,K* HP;2X<1_C]Z!;93;>D0\AJK7A/0>=[BB5TP\
P,Q-SL6RU)+X"N<]5G;=\/,>J]#MH$5B/MRXONU."VP#M]V)U6S!#? ,K;R\3WIBA
PX1&A&=RB<L7C<?+<.M!FPK3YRKG]1%[K)+?_E#,N&&Y/5EA=\4H#O7JDAU3^\;ZJ
P *K8%=K'^M?1)1]9*Z,E,$6D'4^+^_C,"8"4EHJ6X0MY40!8)S-WOY=K/0UTI('W
P:&L4!H%::NGDSI&]E;V+X$_67Z]5+3X(9\,2]OCZIN/Z-&,$P@9K9UBY]S"6*!,4
P0Q&X![PVX%;OW7T12)!,J>,O++A=Y%PD])U02EH+JDD#\7/"2!0ZK\.J--$I3!&I
P+DO5/U:R.+X8%+C7),<(U LYY'JH#=ASD+6:G$<=,39I4WV.YX'.:+%NA@>W#\\-
PD<Y#X6BO!-W)Y&X!9 S40\;5-9L$B%.CD'VAH7!)CO[VI7[."YW6>K$VWAG!4D;!
PN0-\H3$K(L*;**?KLJV8BH&^O+LFK:Z'0%YY&!!I-VX:*6]&$BR)*U.FFZZQV@7Q
PX=&(@Z^9Y3\MLR!HG;<ZSI<*/^0=%[\/SQX1&7%,QPM=IU-)^,>UG1F:PO/75^4;
PE]#8":EA67I(7RW;9]XF$2'N.NS8[$+/69'S=ZYMLN&BGU[79S1@.S7VL3KULTZ1
P_!A+;*;G!-MK&EB'LE&L40TTU1*GS(S\6P>7.U"VPJ&A6!1 :J%)6"#61;0,H;$M
P"4 WJ+(HT\9\HR=!!_.U9G?(_-"@@$G"@$ #!!PH#P<]C@@-N.ZQ<'6&.4^(R65=
P*HC$#ETC;9-$[^%,[U4WXTKN0^S8 ,L1C67B:)#36WM-\P]H48CQXW>MQ34DP=5-
P.9IK^[TVD $X0N1@CY)Z$V+MDC<Z'4KK7^4/D[2]'BNKG.AW%T8M+(3;H;EB?TI6
P@MF$QG0Z*G?0WCC[A"]@(.R3D['XU.)O]ULEJ;&4(S?8[K#969<!@;?O1 &4X/,%
PD#W:Q?1X0-*OF8&00>M*4\38N&7EW#0J'M17]".3D-F45_$6#]WC!'*&^T,*,=O_
PEBP<[7_DA#CB[G9=]_<X@$':ZT["SOS13&FAKMU3?2.SR.]1V^/<IZ>[M)7GX&&Y
P++SK,(%O>>J^79*#,44$"HIT)LPD3=$&'\+8_D4NX05?;FUTD! ;&IN6Y> 7;U7F
P%$DF]L9N4/&=]) LJ&>WZZ>#N*X&HD !Z9<\_7'E9\,8>3U;@7P'75C<;?9>W>:D
P=#L"/<2SC%Z87'&<Z.%_QI45D315E'(]=[H.S]80T,:<$I/&^W^\0 !\]N(" -S.
P9D3R?4WK</F,=HX*0&F$XMK+O<WV/,G2@66L%<JNU(9'4E_G>6#F0E:.;BY9LUMC
P+T%U,F>65!M$V36J'3&WG&F$;QV5#AS$.*^BV&;2P9PBG29JJZN YNW, 1LRE6IT
P5&L:=@5"4KZ':-JV\B(2Y3,OM:.?G1[;6-;"EXYBS75(W\K(YIUOT?DS\?T9G0@_
PIYTIEU//.R,*;X51=J:K(^(E0==H\16:?H1QP6UWJ3E$:RH9,I@AOIZQ;7GBEN$Z
P;[C[<UAD4!!"X' @ZCP$?M2S;/NP:25BF:\0!KD;->Z@'JKB19XY)@\?! (F%X/1
P4P,XFK)U9T(M#.$(.'%055! E]R')742";NZ_E.,3BC@GU,G'48N6['5NK2K7N!-
P.N8"KA\BPA.52$!8.7TFB:$Z0R.N9.%C+OXM2G2I!,]K376^.C ^8H!FJ=V8=+7$
P2(F11UV)@2NN)\UQ,[#8\>7>=Q7,0![]=516IZ,JHF?(;H"JRQ4I12"Y)C9+D"T[
P4H*9/V:7*8[9-.V&QCZ].<JP8S9:7^C]D>/Q1V7?":O/.KHC3+JZ7#Y^;D.+!:^R
P*;9[E$3 &LCG/D.O-ZD[&-@__4YVDQD@P$S6[6J^*X_O;;OD9UVQYUFZGS19T?]:
P&DL;]NJ1L7=BC?X6NM<,(=M:LQ""Z-C:YN(Q#(AI4F&JJF JJ@3I]-HT)K=/8.WS
P 7T(#8XM?=T(/T 4OQ78QX1_,&V!!:_MR4/#BY/S/FJ>RA'ZE\3^DS?&^M]FJ >4
P[P$FN)@&V?MJO<..![UK\P.K.Q[JV_9,3V;$0]Y.+R!AS*A]^L86;&O8T_Y'K%D(
PSH9>=TITQBJ&Z"+R62H2%[H0?U)IT4#T#O;=X5(CJ&]CZ)FK%T6516O_8::B64J$
P0SI )_2EYA6WK1MJ<5-9+H<8?MJ9S>@'.$K=Y+#Z&K!SI$R\KFTCI]M1]UGWOM:*
PVF 7??/R[Y9!=%Q6CQ%:]Z9WSQYS<J4BTJ8-!^AKY^K.)*FC?X)/=(,QJ>CH$48U
P3D(!XDWV-5"!I7W391N!P4 E #+U6A.3870O\SMCV+$A-_%I!!D4J8&38H*K ST(
P1._[&]B_K$#P8-.R1AW2#86+SI,QX)S'KC,VR&P4OE*EOK.Q\:4NQ]4@F34E\F'1
P,:-DL:\.7O.[\2WMB"\PCP;&[$JGS9EN]U'ZL\G6OXI!5;?P *T)X8_F(]1MF)$J
PWT9OS8)[NK0J=P0>]Y:F+J?5Y*$>Y9T8P4KI?"T,Z".'4K_%3JO3$,., (Q:<CV!
P/P$1 &X0J5=1M6U($P+GTO!D5\10O<I%^Z X:MPGQ$KV7^?V38'$H>)G+&M:\P?U
P>8!JW^TCS;\RMSTE0;54'!4QRR'9;&SB#2"N<OD<9MJ.0%1"?KZ[MK'V7'ZS?Z'0
PWCOETT=EX0'46_ZH]_CM0YOTV;%-V,%#HV^BO!](_F?D2>L324MQC&LI5/U"ODQ=
P9(\CQCE^^;87*FQC[4C]=!:[F0.*MPRW4B0Q6LOW3%N4,V!N/>QQ3+8G;&'6HD<7
P0X9Y3EZ\&<;NZM(AZK%/_83R7:]->(141CY&@0M;/6@24*+!YW#V)) =R\#T%C)&
P,WLAH&^!ZC+J[GI_%O,B.%'L@!.0>"D?A2,!^Q[K-3/BY=J.%_RUE!O)[6EYP7SV
P;PI?MK.<<+)<MT/(3E/.)__/]VB.K!'\(%N,Q(SF0]BKPSI<S4",(_4GI&JK U+7
P]+55(30VN,, YTJF[0*C;DH>)/D;&;(V"WQ(!*[,X1RW&__BS*'%8$'A)9)1^6$[
PN;AU:E>W/]#+,:V<]C_PA][]L7MX?R,F727H"(:'KD<-'7V;7=9'P&#)[X5/U 9T
PED*;VF?)&D.8J;&)$:,)VR-"IJ2,0GKU^O%<]LL^UZO$'P\28LR=^-8S.7G!JS)S
P2AN\YGY%URE@;VXQ;Y9X4()AX4Z+S!J)0[I+3Q9W@8="<[R#P,I%(V#++:ZS1:Z_
PHT*LJP7TN2CIE@&@M_:*!S][,;50U5+)IRSB:_O/^J8M2)H1L(KXMBN<=1W03<SC
P=R_215F\*2![R)(:JID2A>NX[!DY0&O,K[B+/C,S4C=;P@YJ"N:XK<;''_0LS):Z
P&/_\&BFK1#X?*MZVJH"9G$#M1311.L<[)!#R)<E,1(_^!;)/\XJEN'Z/"M4.FU0V
P>O.2P#3-&1DE$3N.T*V<; "0(+HQ)WF?+7GV;&_/H@G4*7>=(4H<[KJE.AB^V8M(
P(@'\D9*GYJ) *,6[<,Q-/]1>[]6ALEY\VN@,R3'[Y,;-_]#1S3"NBOA$4HZUV&UR
PQR]#TN^1-+C<%YHQ;ZUC,B<,P]6K'O?4\4 4T1A>,V?+B.</Y3ZLDKF!/X5)9E*'
P;=$W7L-A$PS0;!A3&Z%OFD/2K;]*R!5SS4^HW'C3[F!5+DJ*FW1U0>)K\^LX1T,Z
P-N+U1<D6:'ZO< =^,3D)?XO,CD#F0Y[OW4J"MCG*C OB4O 1-) 7S,D8XN3OLXX<
P'!:A5Q-GT-)]11W)E+4LH1'@KWB;&]!LR*?W+#]]K@2$$2VB,\ZHS?J%RHA_%LHT
P% 0O22R=F=^S^GQQ(.,OXO>;&EZ&%<KH'N]2S>89SI=Z9FYT2>TB_VN@+CPZ%":W
P#&NA$5BO0!&U.#5YE+UFY]T#_;7_P;W /V]+J33+!B@P<G/NLWT4_R;0P&BDYC?/
PT"TK(U!,HD98ZC$=5Y%6#(148$N;RL'+@SVPM0.1!S5#4/-+6/^^L<958^J77_- 
PGR ! (GIP@W[$ ^6BNJH5I0G32R-=#"P*TO2^6ESI\INT7W57'B@C\?V?3:,8)/Q
PIA:QL823LMN)C[?^H#U&"'H./JR5ET%2\W2BUFD,30<&P\/%6XY);XN6_1"L^T%D
P9H6YRC=>KCUX!2+R:H3GMG1=IB88 %"T:U,>LB0NN@&WI]6[4X<<J 4=TIQ+Y?G.
PCE*>8-+Q8./^];F3QFJ&O&</A&I<?$QW4L$OY/L YV/&:Z6;@TZX2O/IQU\&:L;U
P7&TWW\XZE6(39JN_F'LW]_^9B!=#X?O\.9@^JGVSVL]XF']Z5[@AL%K_*EW%F]^'
P,=?Q.GQAII"WCR$.#X!^,,"6'D\/4Q QL,B[1,I[6\LD\&W[S4HX$J:7ZA,%V ),
PXF+$L/]W2QFCCYU0([NW5I>;'RP0L;%<W (TB7]25#)Z36[OW1=G>8K0=V29$YE#
PK12>2Y@6=VKHO P!Z?V"?/+6=-/"V;=+(<K,IT?L&#(168AU4;XFC.-A&1M9C #3
P-TQ'.]B<\QXWD8IMCBPN]D&1W:-NS_,*(K7/[^6R&_\<?^ X%CW"O7_IN>#M_E<3
P(21A)OP(<4_S'+GJH 8M\LY2RNB?.]">O_I*(&;6@VKF(I$0O"LDC^!EX[N7H U/
P/)L.^I_\X_+$=QP,)#'R-)W3 H/)U7 ?THMX:3U.FPP>DIY"[E12@17534J( Q\(
P,RI-+&N"]27?+WD0W[=@?^C"VD[5]QZ$6UUR.T0,[K#ZU=R;'85\@GUK[8:_-S==
PM$P[5E\8]4KT+6+_2#%LL;QH&[%B7L. KE"# 6PNEK4-UL(T[X;O1>8_^*2AS@^^
PC00>FEC8R#*)VQK2(;P2__R3BI;NLQ9@K7O+>?+1#+PU#HF1*7Z7,A62CNH<7Q#$
P.D :E30R.4?=3?34U!MKP>-!FS/+E99\?F#Y.!3+$*Q\5K -2-\*&G58^3U!P3A-
PNR"7,(8F@#: I!AI0MQ2,(@?TRH'#-!T[E!B<*88$X40:WCB^BQ.?P<427,Y'M"E
P]B,?)X_3?X4]9E9^P[O%<XO3>CM.#_)D]C#T@K-*0<-!:WB>N>O@C',,R11/J4T0
P(/?>6P)\(.5XE98^B3?/)(+<:&:+3\SP&BK^L$S1]L>YVXXGJ\/!)Q$<*TQ9+BRH
P45/T4AA.[8GMS\TQS4'DF$TD7>T@P_&3D8<BK-_5KRA\ %Y@/CMN78$CXEI$NKH2
PIH0<53].OW< E5320-];6+$RSE1A)S=2&K4%4CAZNOFJ8_HVY;\=FNP,XA&EU K5
P45N3*F=K#SMJ!2$U$E7X_G_86DZ^U(0Q<'YB<3(QX''=^F1_?"(YH#W;J+W&>"CP
P6'#6+QKO+&^=O-V2@^3T[&'6LBI:LNHY3V0*2M>Q^MY[W2!++2L#TI:FQ5OX.X^&
P1Y5AJ[]N$YEMT1)V=]JY6-"G\U43NCI.LQ#QC>5X&X6[RQ^E*\LU!R#9ZD[1U0-#
PY)*-QIU*U$:TGJTQXNJI@Q4&%JA%@4AW*\=5P\FJT2N'<OJF)6Y QD/ZL&&U[.-#
P4$P41FKXO91'7LY=]F31^0W)3.4V;KC^S-(DS(P1])1>['NA+)\ :<:J7F_C(R0*
P$Z#]FD!:>S07+==$T?A8)=3'-V4U\ZJU?KGE>+(R;C7^%QG<GH(E7?!TE+>V0Y/5
P:Q/=>,=N5*<VM:49]-*NE/NW&AV!?C'^"FTAYFW65^N_!D>D<8R"I-I9_!.Q-<FH
PQ-J4*AZ$ZITJ3]-WA&0VL6B63AZA\\-)CF&U@X],<DM6J9&UJ]4[K"H.0B5(DD9Y
P=1HEXS@5^=#K)OY@=S6/0. =<B(;)$"RBPIV#H?;OJ9.^T#<H .5$AU-6354\WW.
PVO:KNY%X L=Y8NN%UJ[@@T+U]966FMW('Z.T*%:7G(L1B#.1)$9WF70?7N5SXJ:6
PQ?.R\X7PVA*FLUV :'MEJ_/.0A>KNI)=2/<R@6K-64]G1Q'[64=O'CN!R$K:O.$C
P+:"+-P!N,4S"S.=3]D TL,7"VI]:D+>.\<3 J5M;]6H)5# 01J]_22VJOMH1R1.Y
PL94;?4IUL<)<.!=0J;[62.=P'X7,.\$QB&E5G=&49O!>RT8TGO'OYS+1(&H;7/)?
P-2E5Y1EO\]3O[7I!8!?,A%]+%DX/V0T8J#$]7).I_U2G &R!#(U4N6%L4"."-DQ+
P;?1O X8B9=!-R'SW;@"WT3P5;6$#*[JYJN4%FN[O9E;LW' E=Z5D)3NI:F\^!H^?
P2I"KWY-SE:WAB,+#QU*+?=B5PR#)Z>RX^ +@*;2P);CUS]K2,($:@6^[]*F1BJZ*
PVO-UQ4""Y\2;@X7O.W>:W'<(O#EQ$2_H#V@E M>GFEG,G!BD6H*S"M5N*:1=;!->
PU$6T]X1:SK,'3LY,!<2Y=V8[=7DJX"=YXS#95ZHA%^5AR2 D7ZH%9P*IF#0 G_CP
PMV64.W?.%L\-VWC>J"6V?,(08JH\E@.ZCC0 8:PMINDOMHB3F(4IRZ)P+U ^#D/*
PT"Y1<6? 5 J1#H=.:Q:>ET!J%X/?Y:(WF^"R5"-N)R/UKI1OFS >AT<NI?"[?09=
P,1I@K05B&Y&H"-ZCZOD?@)Y,OV+WIOGSEZU]QS)B9XO-A,I<_7*Y)BB-A1:&+@*L
P9=.9I:O-^.CBD&LFL?: L3ZI" 821.?]MB??X8]<+TU%7UW=!8>E#M#8*+MA"FYV
P?=GK^,@:$J,@]2?(0GOB07#_=$_?*>K;9](L9]BCAY]#KE" ;T_EDD>CMW&2Z@)W
PZ(+]!EK\"@W:_00E =[*=I1> '3<]*V=U@@HS/3JFSA[FE@"5&<?</&FQT@DNN.7
P5^T_)IQ;:>:#WP%;1V\FN$[#SUF<'\6=3MKD;OH_*R%X%E;Q^;88)H?3PP8[.!K%
P8''_A!\YF_L"S!_%"7045,_V\L+\%_^S ,E"KYF#\H7Q2I\F^2YZ114^F''AR?;2
PBZ/YA_+Q^B<#8M%[6R/MW(5UBI!)<*5;\J$!Y=O.4D@!Y44!C4-+!_LY#-O?;0SY
PA$PD0-X/BTZT<-UNW.;#GM$]Q33@Q]^D7&D=?GRRHXG3[YTI)UTB@+ER8%6=P=J!
P KB:WXW[ [C_6;U',! /\6%IJTU2:]W5I,Z@B?]OKQS21?LD<*U2= 8:)EHH6F>]
P;J0H42U$02Q5,)D8@T1RX\"K9!HDIL$?&-#,>-F6<;P?&T(4ER!\)&T'JG%JF BE
P>?W!>'7'B?LS\FM.S8O*O6TW:*L)X5)IC)5-#&=(F/5+=8?HGXC1Z)OT?^2[Z)M_
PL*WZHF(.KJANBY,ZHNOPSV<.Q&3>T4<(5@&:^@)I28TUE)QFY8U4L]"8@#Z:$I]C
PL<8TP_A_$#8^Q/MYAK6?6)M$@('@F#YQ[P<S/[>G#REQ\9)%5Y$.*[W7SO?P$(-%
PI!V<;T)=6*JL'R^87YA$LD]^;.4\U:<N" A# 91/I\?H>HXY568@9=="!1!D]L*@
P1%N]PZ+L9PP#(S:XHZ 8=C$MVB@*_' M]V555W<K^!*G=4*;B@BE]01Z+RVG$21(
P+ZO#,D%3MLJA<C<.+#F=RN07=^4Y0BG^MIGEYH#(%-9CGNEPH0HK'>59H#H*\[)&
PV:#.!\,M^(H5$\5>QED,RDA'^;I]+ R:5!<L# ! B^,[%+Y%P!".IA-V:IE]U+B9
PAN#RCM(<4UPC*!>5V7$OES!-72VF#(K2W-RN]2$)UQSSV\ZCVQ5._MZ&&GKY4(05
P84S"1"A:-T VYH[%)S?,T[<V"G??,#H3.\X+2:IR0U5I7*DL5HQ5LT4EUB*VA%RZ
P,!=?O7XX)=2MNI^LC6LPUPNKH/[EPGH@>A>N"\R7#P4<=W*-(.6$9XF@Y$7H^U(-
P5*R70+X=O\>> SRPXJUBKB@0.^RZ+F9[R[!NNA4Q5-+$< + XU:]!7C9;_KU(P>&
P1MNNV7)]69%RQVV$7=9+.;WADK\D__I?SR#1I^_?)#ZN3Z:)I\3RN)"HM)0]Q2?U
P+>+E.@IBO0@3EG.<RB(<*+;$-2^K;$RYXN48UL,Y50@DE;01 T E)VG7P^/\%W(2
PONET#WT!ABB=1H ='Q^ <5:LH5FV)LVQLT"+43ID>/UF6Z\)_G?*L#Z*+E[9S<?6
PK4I:)')#<Z\.\5K?CHC:VW5Z?7QP[9>G_6.4F'Z+4:S1*H"-4W+"[[\* =8G.&#X
PIKK)*_(0A8Y*LV<&08H:RFUA+&IG>Z0?-),%NJZE*^X0QC*_ A.9\*\<PF_VH1#]
PJD\"Y"02UQ]#44FZ@BB[]E&_R/[2IJ*,E@M*G#8"2=VLJU- O=H2.4AI$*0L2K,J
P9W!5'/TT+5@XXH+"WU.CQF@>R45D_1@]F8K:TJZ7Y;EU?5LPVA_L%'&;Q$9YH(?H
PW^^2YP40'.9*BQ\ E#=TOUU?O8,Q1IR^-^Y_$9%U%3C8K5[_?PG^N!) 0>S[XO?=
PGL:$U\-YNO#@1YZJD-UCB70YIU6C=MD/U#2=;,5GC! Z8.?MT0G_@+MG.@<M@QG#
PD1\KV:.(.(K("K$1:#*L)?6D)8C/5YEU00:- !/H<.%&F*6+>K>X+PL,P=?>(7SV
PGF'F8C$[JK]ROT\;*FGT18#,$?YU.\0!C*'W->8^Y\_Q/*AUA2D2*/$/R,]X-*!U
P[DS'KNBYLO]4GG2*7#WJ/Q;9<:0BN-<OII$+ .13J;M6K6-,]J':[)4"(O&8 YS>
P,EJZO'.<+<CV^NR4&:S= 0&W2BH7+!&J9L[&3%I>%[AH[C%'=A6UI(<\\8'Z55YU
POMG6E=Z ^X*[[,$Y.L0C/FK,-VA/"+N#%!&MXX 3U-M@':<K:#\_\TWD[ZNW(LY:
PTA J]6'VO=3'.TGGVF:_6;#G=N3 6D+WB/LB:2Z$<S;_@(_( I2C-4V^LK_PU':!
P#KS1&L!XQ]+/",.4+ 4&'1I<_L)>+9+=40()RNEF'-ZJ[JT/!)0U L8?F5E:3<8J
PYP5.?3.=$O*64E07:@1+5Z;9!@KA&@0-;_*NTFG29B1?(@NGJK/BD+O%>@=MVS\/
PFZZOLLK$6E;R^[;=.],$"Q!_IR]8N'YA9Z*%X>AFPI7)DS3@?LNI%-37ML(;L=&A
P:JA>T1SQEJ+B@WAJA7Z<[<8E<:QI/CX!H^1B G.RIF8UZG"L/(Z://-I](D/C7(-
PN(\ 2?/W'*"U@YZ[C!WD?'-W&.]W0W>8-2B2&$4+1(=&[M@Q)"VZT\>2A"!O/S0%
PF&;^0OI90_CP_U7YW8=(6KWVR)4+8[\"@Q+SNXMA^'_@1L+2F3<VN1+:D922H /L
P]9O?.2J"DP^$6IPW0YR'^ZXP/KU97[YA6V EGK5*F'Z3JVM!$].H'0\B$Z.J=D84
P/LV$QH",=."KYU7%$BAQ@ZAMVZ,_@3/U<.=18U"$!<9%\/DL.B =/NZ"ON"$3O[)
PENAP]N__Z'.W6W5#7GY!0>KYL3G^7&DDMW7MTR#/Y&-C&- 7J4=K%Y&76)(A*H/ 
PD8#]^!CP]66?Q&_^+:!B^ <>3-1M^U,\\ "*-: 155T&WL >MV>B2[(A[Q3V]*= 
P)26%'Y=TQH@<5S80M0PH&2&2U(%-8)\PYG:0GF+5B)XYF"\WBZ"390%R-W8]-,<:
PO+,TM\B\7 XU:#_KW@2@;O@<@5I9MN ?DI^<<^0_*;;S3/.,GV8/&N+:V/_C4B:*
PTKFL]%3SHBM6KI.C>6>17>):;3^-HQ&=]VP_1LZ'.B/!,:#V^P$GE#*<9DQI'R_C
P8,.KD^H,(8[]@3S$G[&:$_A?&964[R$,#M*CT]4$IW#?Y(8[YC=X\4)^Z-'"B)P:
P;VZ)T^Y#.2*KO<1ZQ@ RU$,41"YK& 525(#T?B6LSVQ%(V[OZ=3S'(T5A>Y;HTSP
PE6$!.N>#/(9>1IG<,7#PS.[Z9XGYRE^J#,TAAXWU)IMX1?EZ$_>EY"[;?[RJ?^6<
P\!Q4Y&4U1HA8VING%]LB*C<+Q5'3H]?*\MZOH@H_4V[Q/;EHX5F2>OYS-^25*PMW
PJO5.'J3][7,T ECNP]$1+?!G=0^;[I>!<L6!J>D"MUAV3>T0Z$#<B=%:_69FE3L-
PTD2'3O9!F^%=$X=^9P8!T/3V]DF23"#H'U)]*YH6; )IZNF:!.=:D.NUFF9^AQ&I
PD%X3V%K,-Z#?R*5%#^B2^72$O ')T'?VC/C]CF];R[TWQEB-"->*WD89 Q\\X4LL
P/IM1";MC'!$+@>N2=P?;U;*(J^F?OEYH&6?(FM4'$C15U'E<8U"O/,TY ;/9KEZ9
P>AF["30RD_N1!AJ1-0W@>Z]$DO%N?1M6O9#6WWDR(::BQNGNSPR+(&+%%D_+MY:3
PSJ<@P!5XZ3%BH*A_Z;N;7)P5[P6K+<9*1S]@$]4N*7M.3-36^]FIQU,NJ9IW=F4%
PW?<_B[I! )CS,_/+N>-?#,%^/]$BY]#XANS6EXVCQ_V2C,9?.HB5)/(@V$MK#[C1
P&(B !U(J*]IUMP-%G%699R^#Z=D(2BV8>FH=XX0O"Q"!??AVOC(\&:C4.X33>)X"
P+''N4>Q+'V\/KUQ79\>Q31/$Y8,(V++]W0:1@6R"87YG%J:^<IO@Q6B!0&6)_0"!
PRS,EDIC#TYW[AENDMQ&D]RFX<C2S9?%A#9QR^7W5B@&)7Y^%[!=Y]/YKW>]0A<]-
P/U7'0WBDI=5$.++^,>U]042[V\7FG:L57NVPH)([R9Y2?X-M6G_%6FT@R-;()</^
P6[IM_93Q2=#S'%I$Z)UBG8J_,;3;]EQ <:(E.F6K5M@,F"G3+X^5]GT.?&I5^H&R
P.=D=SHP92EEAVY,(@Z;F79^H38AQDZ1NJB\AO!%VJG-7ZV2\4IWG!S.+[\M%TJT.
P;WTF"8(K4]C8F<9QY2M'+H].?H!OO..+^#VK.KWW9H0G_HY-'FY$8J6W@]9!#4 L
PZ1:%.=3P&!=S(6?*2N&22IZ KJ,[@9\SH 'Q."4[1S*7O?9_WNWL]<GEI>ITR(J8
P1Z*F?7MXRYB)Y6<[30+EE;'IP*3-=ZAM(*01?WWOP(Z@$&"?ZA>[\">S0],&ZH_%
P])1PS>=<,0?2J&+-SNG<-Z1(O^<G9YFBCK>4NDZC4=J%T'5+G:A#H?8:MZ\>$D1@
P>'&5MZA*/O2_<\DKY:X=R]WUV'PHWY@2=?@J3Y%THPD[L .A,],B:;49/RP[_1+0
PKB5^JQ%)),3<!1^?)M'<'>==O1G#_+;H\0&9.U:I@U+IEI$8%DLM7GK%PS\^HM5A
PEC$K LE-$3PWFX->NH#B:8JPXRN55):R1I7-NS@JR7&'%:O#LCQ9-A 0\_?#589\
PZR,;KWZ:,P.?K'Z 'DTO=H)#;'W>S#H'$PVNHPK9D9,IKO<E0J%/F&Q_[DZT896L
PR4VNN4$[I487*[3.]K'"P32==K-EF-;_\>&*YK(0MN?^/ZY#O8/BW824DN2F%&<=
P#Q,XZE026R@( $@3:V8>S6*M)2*G5K ICAJ2!")5#TT+W7<=J(M*VDKWDI[DEA8"
P([73A)9-V7")N;>SM"&#$"H_/,G\L\WCT9B$)>P[SBP40"M1):\,E:PQ)"&#X\7F
P<@P#5P8ZZVA@(!C62!X\&9%&.DEYW-/N<R>C&[JOJD%?"(/0[5>Y=4>J[59VDE9A
P;_(1#? L1BG70+#&?6R::9\@6& RL*-CT(B$T4T78WF?4^3W*^'T\2E(&H*'399/
PXE?++P9ADZ >!"QDZE)2%#\MP,O$V^=G7%C%!=3\IQ)#KT_%0Q..P9,.GQ9?A :T
P_/;@)"3WZ8'S1&UR-('K0_8;D?:W/]GFX_V%5__-L^]34D_*^44+.[BMV>K?LH0_
P3C0P[H=R5/ZZA0E9$ &_7F:L.X!WF%_^G5)% _VM0K;=!YZ,QDU!U'W][B&"KDH:
PTEXB!K'[[C,3E4+!J"+S?G,2?*% ZN]E\W?R_G>#(89ZJT 2=1JG_=.MJ<]EQ<Y.
P8.ZA+.UQC1(6.Z'^P*V#,^'WO&GE+9PO5APM,4@74.V1.UG)%$DF8@$^5/]YE+!A
P+6Z[CRS_EY4,JMV<KNBM3<K1<#T+9I^NFT,ARQ5P<[O\39 H&3TS D<MT7.-8<EW
PN&?-T.^.7 (.Q4\LM@L[JM;@',*@?7\F$V*?,O@C\C/-Y^Y13$ NQYYY_ A_;<I"
P !:Y)N_3CX#V6IJKCXR=A\'UQH4Z&;U62^'T!]%]AOQ8@[!MZ;HUU"$#CL;:NDJF
P?'JOC.1ND 1(94D[FI8.%,'GO4BA]&=GG&V+/6J[*>AW4.R1B#0- W.[AC_A+-X0
P 6L 68U\/DNZL[$3)S>9$FQI<Z8+9#U:55E@)8(9#=YP$J<+AG  'W:^?TEDL$Q\
P1Y=)RO]*+2K9@%N82N9S<H+;);Z$DSP3 ._I8A(AJJ<,:)3>W/>K*V[<0RC)> ,K
PN$9YGS5(K@JMT35QVHL*F@LAH:VZ[Q]7 ?]N#US]6)]=3Z,WQ?S2OWG,%O[VEN2B
PN&B)'[I*B;- 9H-ZV:[@LK%4)[9/8/%@)8D_8,D>'5T:&<S9K[I8 X;_%,\SW_8X
P9B'ZDGR4.=LTS%\CT+Y[P[J[SR@Z1<F1GZ<7=CD1$SX_X+811B:-4M5X_(LZ]?>Q
PZ@9CSWF6[HD*A-1*54A0*]],&L56@IBOW%POF68W5=!J-NN-P1V[>2*% [ ? 1U>
P1FJ]C_K]^RF.*B+HU^+>S'.7ZO?"5T*@B4O!K?DG7_=HX5D-Y]R^=>$T2-.V#O+S
P]6V']$JM:$$$@ 1\&BW704 K@PV\ &^TN]_<A+Y7 DR0MU_1I/84W-+)+*71L9 J
PLHP7/$U;<39\I&WJB1M\Z$$[=J7_/08G!N? =,-@UMZ$_(KRHVJ[WPQO/=#F^-(&
PK\]424'Y7KJ8:L&O0BU3O\TKUQ;5PU]M4U$^DK,Y!SG9J '>HW=R;@T$]DP$LPC)
P;B!_BY8!&2W5,7M!B$C[$/I6=#8Y0Z!IN\V,9@+EE2?N@#JR66_=IA@&6,_SC1GA
P>,#3!7ITD?,9(6J85;QZ$(RF7*;QVUK>A:RU-/<T@)J+;DG(/P%3#X03[W%&1*+>
P0\[QAU&JHA-T5Y<P(AP$]=M"PQCZ=+Y_IEB[P$&"41J1G"!.<2>NBWY5QSA<<Q^O
PRV*7-4W;6.R)T5 ;%[02O-E'X'-;447C5B>)9DW=>233OC1SJ+0'%&S[LVCBW-ZP
P6+=>^:R+R#B%04><3KVO]MRH9C[9#BU$SY<!]T\^<8?0K:H3#?LN2 P].H:+MX1E
PR5>@V.4<57>:TQI:RY^G\862^H1EP:C7E.7H7NFX)!D67&U71\#O.4U:IW#"DO%1
P%NMG0=$E]0*^&7[,89[2DHO-I]![54I"15J];+19;6SD[-1 :KE\SP$OLNPC$O*U
P>J(,GD/X5>CS+;:%!'@?WVC=V5".Q[JK^Q+PEQGXB:BB3GX'>=*51M[AP>$U7U/[
P!<\"(:GK6,4N8C2Q5"A!/5G?&[L2GF&2CTPB3R?%&;B9QK+?JTPAL-["&=T+'IE_
PX&4W7"IC62^>& #YO;*P'^_G)P]]=,:>W\00-$J*AAY5ZF\!Q./*EYO,=4%+^Y[:
P^AQ[\MTCR4(]UL?L]T>] =&&#VK>O(4=2M% SR!H9-YJ,HK777@C!#Y]X\VT3'4O
PYLH[NJT@>KGO=P;<=?<?PR0K99T_63\,<CXUK'H6CJDX'AWEER&<H\^O/1K(E7[9
PENT_ZM:T1@TJPJJ/5@.57\B&$V8FDLD<$(U)!]'[[T&[YA>R N>W.T5S^/O/>_K_
PEGH52P?C R&&4!KB>QD@%J+A4!67^(5I.Q).RW.@%!PB#:K R8C$&.#QAA"ISNF#
P8:!E:(@L).>$34U0*3VG]6AZX%+X>TD_J3HEV_&7O,J'-"@M3;@46&9]3$H&R?AE
P54P;RGSE*D2DUM4I;8\[-'M.^81MW(*23SEQ9%GFMSN?P2T.[)+'OJ+3]?0$M$ZD
P6*1^.&GA?0GRYC(5!K,5N';YK3*L+N< G.61+H61G!XD :(TP659L$N F__XFN/9
P7O#J_"%U"VC9MM\G=O8B@K];L;J.]/*@P#P8F5]7H.WM)N&N">LP48#)['(M3.2)
PEN(8%*QY8O2EB5Z6.=Z+JD%\8S\7">J.7"9EY*<)TSF<7?ZJ:Q&S%XHBFYX) 9GB
PGC<I,_%0%S#]@T,PFG1;-<A9X&66N=TQI_$/WB0A.U.?Z!;'$&48IO@U^?OS.88!
P2KK]U38C2=H +8Z*R&52-I:1';.?R:KYF)?O$JL3A&^1?I[9VQM+/?"[WY8-ZR<I
P8ZD/BPJ/*LTZ<)89!4X&31=/\AAK%H%RXW1,XMUK@:UCKQ K?K"DBF*SCJ1[$BDC
P:ESH-TE>B_R/Q453(H3?G/\=?7.:,HK  GJ.T'[;\V7.OFK%$;N!WB]D0873K%$-
PJ?'?%339Z<E8-6D8(D3D&9+AALY*FDRMB]EP!(&0(=Y",D@J6=^WD85$F$B6#R7-
P9!&=O[ =0B\FW;+Z./C@#+<4TVJR%XJT83,,5GX6WN_D32R>X2"P!0CFICEPW@M8
P\Y/7"G]"F24G->,U2(V)H@DVQ'F\K52^(MJ%:YXJ4?9#Q#EO?H+FCZQ7MDXY'C]?
PLNK$I(FP>E<%IMGQB1#&=MHV/!Y'@WZ!-XF\8^H.9W/5_R)-V0CPL!+0<N;TMGMU
PS8^&P.-'#75ZOHA^?$L>$,8Q=,P%;8"+NK,2&-W7Y>]]-R,6+/"T"V46*>SZ$X2!
PJJ#PWQKG6B,7*NOKA)DS0MUT>7N0*LYDM$-J%A^S:G#3Y:"P<AV9UZ#>3]COY"J;
PUY1,3+8YX &ZY?,OAA=#L^&(K(2K274Y^G,\IUO!CW']<.'RD(L8->&22:E(^W]Y
P!N44$Z'UE>+OBFY7F%4?K R5^M"]=34(XT;(A1=$8_0^--52PCS-47-4P;P+BPLC
P<RMH9 (M;-@Y83JI*5CD *JDS+*(9/[M,%TE@5M.#59U:B;L1> 4XNUY'Q4AZ=7T
P5"S<;4=9!1Y[,B&QU]AB^.KUVM2=Y8AZN+WV%CJ?U=KU8A9N\E!U,%"03QF/:?JP
P?FGG&[?*, V/1EBO:UW5AV\JYM!9%61>S'.A>3*XY*, 4H=7-Q8Z=FEW2S*D#T(.
P1TG5H( O!=HU'_<9(LK)^[SJTQGF_X0%6#0HN*FA4_U-J.&A1J"N/(0=?'1\;D*D
P8CH_ 1_4]FCW"A?S$RC3$U3G8P#IOI$1<77UJU ]AA$@AC*F>Z-IN^X^ ZFP:$05
P<I(1RD^(S#&"OAM(2UXPU+]YY,:Y1GD$<*T]O=3C=UD&_6VN/;HX.0+L2$[2T&=R
P^!5<D<DP:RA^ 0ZO6@V1.) =D*2/;/_WG#*RN8C%+$@GF' @)QE_3S*PJ)-KH4+D
P\J2!IUGNYW'X@L1+S:24K\E)W?6B1$3%S'E7V<'-RN6 YGQL^9_HM?<7G58986X=
PQU1,*=ET1J1$X@?.<VE]WE[M9GAGOOC52H0NF_@X8ZR1*V>>(/M 2"S,9_B,/(],
P9K.FCIG<EO79[LFJSYX8NLE>=*)GJM/P91_Z<_\1KR$9*-*)I.NR7"#*%:>5):<&
PG;+>4>NK[AOK]S*BY<^BMA:Q^IB>/J"HA9BB9JLY^WSH*Y_]4<(N<#3.'[*&C$ZL
P\E;L.R!+LQBHAV)[+A=:$H$SPP-HCH :XOVSON.0M[KV,9(?VMD?/#?/20M^JYJM
P*QN"&!A(CB5[/49Z2WM7-%ZK'-XS37/JRB-2^M.T^QWA1:<H,U:3]:.4?)6CF2H(
P/"M&',,] (O\WB8TP$O6'N0W_4:^M97-<1="]_J\@"9RZ' E)K=N#Q-N$$R*R9K0
PQ^T=O5)K'=OZ$^N_#]SC8SO#*P6O^<!:^W$TUK;!;<F?_=[[+H<GTU6D],H\C77W
P8W-)'OK)+I209>T!HQ(>?[/]$X>FUV)G7ZE6ZEG$40YWDL6ND7;5_L*5<Q;-)Y_R
P7+#B1*DR6M/JG!QL-&/VM>7'Q6264@+A8 BN<[*2"WL-Z1VVP W0:/@EH,]ZHZMU
PTBJ4S:&"%MQ@@".M.\UZ!)%:G$LSJV_6*D=)/K*KWBT]H&V]"_QZZO:J-PKVUN/W
PWC5\!0^L^N2\XP,X"'OS$,L2X5O!Q.)%J@Z]U?B*;T*X2_ .8&0TXU^7Q5?A[;[D
P( IZL6?Y,90ZMI5N#7A-$NT,Y<%B@6N!XY@*[KQI#)33H).'P=ML;AR:)J(2U:S(
PVO=(^#;+,\=0KMNHLO 'UH%%N/F  6J:2GEGR@;&;);7BC;)DD6AW.U: #F4QY)!
P'K=OAV S$W4\W$D.$67%UE2/2.X-5+DQ8K>!\S"->3,P*?N:$//9.TTV'KPL4S[5
PYLB#*/.&U;6/K 5MJ_L.QV*9L^";#'Z" U\9S)40FL-N)II:0OE3.)*_&Q-P/S%"
PJX%U,G\1%$G2OG^3G!8B:-:G0R3E+SN-O'#PV-]- TP-/JP@X&UR?8]^2U9-O1'!
P.E'NI@*HOWWC*^'@'KAQQ* 9R]UY?<Y<;"RQ<>&2P-FG"TI<&IRO<PBTI@T7<[*0
P&O(H64_2+^(T24QN$Z#RJ&9G. (YJN!R/A_ALDTO;:""8])&KN]:M@T?CJ'DQ=2=
PIC7CH L;7N7"NW_$4/H.CA_1%G&,UZ9SNIU>1K#O?_4M I7UM@[*Z6>,[2DFG!1\
P(,97SEC+A S9NZA+)@R[C$/B@$5Y#HD*31Y?[W9$@MV9$,4ZD?T!4N=2R:F+K*T/
PE?&B',<<9'G18@>R?=Q/+?!_R+8&J<6BBXTCIER!(^TYMLN5XG+$#\-@)*ROG:=S
P__#2.NIC+I_TO<HK:3]?ZT2P@C^MEY=O4Y>WY:YJG>U!*U"_OW1CHW3+0^G^<\'=
PS>+(U**+QW]CN3M_X;TX(M2#)"GL:[%)">-_9)40:L2$2FU@95/C%Y=^U8E>O]$W
P]Z.>'CVZ#BRG 08-Y<R\(^=ZD8W!.ETC+C/&(6I@XE6/%;B'ZY<.\ ?4+GHP+6$*
PM6]K?)_NEDPA=SQV&9*HK A3TL>W2Z& UZK! $LVZR)[^9H]UIRQ_P4>AWQ''QLL
P?/+&<O]&]+C+)NLAU"O);'*7[-SV+Y<P3 >*>;4.&MJ!)/.MWW2W[N'IE1X1KS*U
P/\PLO$&PR.BEW7DB>=Z</DQMGNG^L>OG/@B/E3Z3^)1=(M'!5S1UY@>U%JYJCT!#
P8O8[*2*ZY3 3C27_EJ?"Q,;?+;+V\/1\MO0B38\\;WON#)[+?/(9!E+LR/^R$S;Y
PPQX*<&_PCV6VZ1W8I=:\A:?H7]/LJPUQ(9_L.>[-'U1_7[E5\ZD*J3[)K4T SWC,
PO%@A^O@!EBR*\5[.O4NU61NI&M_BQ9$E25RQ^^ CN5\.#&M)Z_2$0Q_;'\>Q9_CV
P*_.VJ1I#QWG2,4\>!>"[D FM8VP6+JF@2$C!D*2OKX&;HZ^9TB,^S3;0, )0-1)]
P!P$-*K+.-!G(8\VT#,'0IH.\CK9$LF.7Z@-J3D[;(_0@3NT/&X$R=3*!1,#^1J4;
PA"[5 \[N(\-?(M^SH,U/N;]6_>:$)B $(0(:RSOTZA)P->P=(N+JP 5F3Z9-IV98
PQ^IQ?=Q47-8237TO.3:4K3HK%W>Y^U@I+T47TQN%(1\7>/'%P?^\K*I5SB6A24T,
P8++F7LA081UR"6(28\"G"3L<(>Q"3/<0 7F^( (D\9;G.-2+K<A]OOK\"#(3I-RH
PCX9C("P-P-M820CD="$?5C_1SO%PBE "-,#W*$98&;0.HZR2,S,IG#J8A!,3$GUU
PD08EF3B']0@3]>O^5,MP1LDRDS7  D7T<$W(5=5]:VJ-5UBA?378X_#_W\,F/+#^
P[?#,QAC_IB#KU*71LO5L/U>\%':?^F4V2XI-0+\ X^\L<3>1;O7F>BQI48"Q]+WX
P #T,M)\K[T]7 F*:&N@WWF]N \B+140B%R-6UY$98Z<[C%\TIFG6S^U='(1;:("/
PY0736U/..BD.G,_ZL]KI<N$8Z=5U'AA(PR=6F2?NI@C\<YHMDBIXO00(BWB%20!N
P/KJ?Y_E#D ,6?(/_APU[O [.1\<W:XT$>/M6&X&7:!W(3Z%H2A)7'8P?6>1%3O!<
PL:&Y"!4](5741UD3 <%A/VQ?CDTE%33U?&FL+M,^-7.KLB-AK:#L("IQI*M%Z0G$
PZSX<U.SINLR]ZAJ[&!K&/=1OR\08^^/UI[(RNFOA?*DYJ[2@XG*:?T7,Q6R!<#/9
P(EQN)C0@4Q[YCMZ@OC%W=EX[H8N;@D7W.*@B\&E>Z]HZ4I-^!NA\ 9Q0*V6B;$]Q
P</-5GCI*0,3#G#@^/\FF,B$00*3N(RH#\HS R919HCP4 04:1.CEBQH9[EFJ/IH%
P4LJV2'=GIEKP'YH:5AD-4D16$UM)TH14(BBF,:DS[R3U7V0:<@D7X6XZV:C^\B[?
P8-7"84C/>AP-=GX=D;X$O1RXGI24BB>T=$GP RKZ:!MU.Q]^73.7\E7M-V7 K?(Q
PH<SQ-O% G1KF%0,48BP_J_3D*A_2GA[00^9/LF0MH_YFZI5X9E25@B_#1 2[_Y%0
P[A FCF5V$J-#MMUY1MN=XZHYN_)QHL@&[\'I^DTH\B^R&@QC,OQT9=>^Y*B14/J!
P$^C0NQIM7V<)#H JIB Y VK'*^YR]9L:] V:2^2B.FX*ZWV3W]F/ #E_O0G]P2^S
PV@U!=2H8W#_ ;?['9B%M"#K.R[ZF\\0BU@PQ =.?8,2.T^W<U'1O+_,?@L,K0>.5
P/68%2O>,UU+8VH<2<. ,EA6UV^'/NN'3QFF<MK"RV349>[*]<Z!;'.;A9XXM]JYR
PT,1]'X\@]F75$H_,L!VF6[ KY*%FT9J78OO 4RKG@^U&@0M[M=?Y^ZXNQ]7D4[[A
PK!U63,7J?W5[$> \4??&TE)E*/$Z:"U-*=ID]0]#5#\O V09"L$":L8"&) =^BCO
P*8PU.-.P,DG-\L']_W]-.YCMA4R9BV!'$[!B"(T8FTG?X;WF$A7LV%\02F(Y241Q
PK''N9VX,EIT/(\,TW6O1?*B+?)535V?8V52$PNEI2IQ=O?E0"OFW04U8NNJO/D%U
PTCA?Q26F7I4/9KI7Q*X7$\-!,WT)8"-@ DZQ7CF'4$9WD*@.<WE07>Z!KX&)[ZV8
P.*A&1W(\(,9RDLH@FN<L-XI9,!=1KDY)^2O'EFSKJ-8[NX49170$#A;-='WCTGBQ
P5DO[#CQ">?6HRI=1H;.;=+[@R3S6,E@1S6+]:#;PNQCC"RE0"FK6\-0,U8G@JU9I
P#V!K^ZE[<1[X+F%]&;(+H-YYF0F ,9& ([T_#L*V2+2GZY424H_%(\G BFFE.J*;
PKO$D2&:2TTMX%NMX6K&^@%H1L+SJ/PX2#UU5B;1=6C(F33,M#N$$"-LKJB$0P-[>
PIH8>U[D&!$TN!G>A%WC1H8^+Q>UJXZY$FKW@;<XFO!A1K@5KVU3P^"Y_%B*6CR'C
P;Y;G[")KI\YG8WX2=6?-GGJA,VTS,2C X(X$((1#3-]/DI0-/PW1A+%E#$_SCNC9
P"5,*V5I2R16^I</ N,4I (0& 6N-? )(:TE2QL1?,;6V!1E;^YM,$"#2%").N#6T
P@KZ! ;$QG+._(M2CJFJT)"TR95QN,T."=4ANVO8F-G)F!#D!W!D&O[),,]$5*\!-
PC$S?@K >5@XA*T9-:^ E4OH:L7/F)B8WLV0JGL^U.7BEPAJ"_,0JX/(5UC?S[_?"
PG1= %;=GW-LZ"72'KN"Z+*K6:I@!*R@ZX$P9%-2)MPFL,4P$V'C(>5U6]GY!:T\Z
PF^H ][P8+C34EV;%U F;/(>%=#<2(;&'-*M4A8+U:6=Q+YQA<X4WFIO%>R%]Y_^[
PYKZ0B!EC%1,D<]7X[.LT>K-?LH95.LF83.BP @1290#)[-7VCNZX?0X#&' ?1^,9
P>?*%66*%JV0*H(!RV_/YS>K#F)*X.2VW>5^!7! TD&/&OX44)E39V4RCL?MRG["=
PW!!'=GY<+_#P9:[* WE-LQ EO:?@=B"$.*+Q@2'?=7=??ZC/?YV]="=-:BTDE52Y
POS9HT=BC+S$):W7H'P=9S+G>S0_T54<%XF73,8+[MH]>![B;AJ\MMV'Y)Z:/ZYU.
P>&!V*\_+=L^"9P?=HXB6"_B S@R/VP6%7"C=_=$JIUJ<:$,M1X3KL\&OGKQ:6_?:
PAQ@SR=[ <][<>C15%OKDQHG HXPKE^/+"D.' )-*4.$LF,''7Q'81>%$QQ_MR1[I
P%;'$ +?>R0R#D/(Q0D80*DCDSKZ^,G7W0-*+%W25P N&J'@GK_N-;^!@,*V[2/C=
P$2,M_@2HR*."C[) &1[<[0J]/;3*%W=R]PFT+[[__4Q5*FAJKFG5* +=V)(,7]6$
P1DD;.!-#Q9TS:T8^5\-I<-_&.FJ9%V9#R<^.1]TU H\W\_;G,3(8$'B6HBQ[EAL%
PC/7.*HQ))U?<TR;%6.<6IC2%/G;2VN74-'7ER'TTK@("^\^CN-F87418R#C:4GR8
PBTM:HJ^6)K OSNV6*%UKCB4A?(#6G5*9N;I!1B\(A<?5NG>(^'DDJ2-'S?=X(+FS
P#AB0O8ZO\ZE,8^RO2W:Z2P!O1/V.V4QMALA'J+R#PGS@0A!V2YYW3]<JKB]!X+F:
PH33MZ6M)%YRR]$U8ZH:J,Q]FLK.?P-F, 6?H7&L8-?6?)4)&MIU#PD7O\)_U*S)P
PL2_,D\,+T-Z:)ZE(?T0L"IC_NIQLM\8\1Q$C2UO'"ZK%Y= ^B29A=7(XQCLC3O1J
P"^$D7,6<O ;'\I1$@92XDQ77/'GKUF%]4U&5T, 9=&&PSV,"$'':&W+#E>"NQT&U
P&(F5YJLIQCZ2!</\Z;_N^_;S4B@ADP03<!3%%M_HFV+($:5P(](/Q?$+#V2\4(P#
PW>5<SVAL3\*5@KHTVF<M;/UX;*(#PITS\8,^3,CLL>@NY0+/?!XIY4OY/% ?=5G-
P=,\*8S9C#02<=X"]\G0'7T=II!R/4X<M84U\D#G6QX]IZLM$*4[>XUCP->*&P)03
PGJ/$.RV>T.<W'JS\J\)>WL:_<J.]R(T@ YOW71;3T4I,C*W+P>.WB5!H]A#BQ'%,
P21E:ANS[U%EZ<&1EWVRX% ;:\6:@@@5GUF/9=.V5CR\\>%RHDV![J$T.0&MZW%;*
POS>K<(XO=(E%9/JOJOCX;\3]V2T-R7_&J>O/F00WWSV!>2N,V)\\%AQ-L!S4CN).
P1V;+;%H9IV3BX8Q+6VM<Y0"/J@TJU[5$7ZYZS!@JU:1MCVUEV J%($^0E6XPEIK:
P7@4)>^75RA7]]3FUMNQ\-/FGPF&/CJ9V@PV]*D4$>>P7+E]R@4W^:^#TN<>M8L?M
P;3N6G9]L*MS> O+*CHLM*$[@P)0?#$ $W[1!"!B/.HB&4&_ G]+,,[2OL:53+QQ_
P\7A\J0J>I.RB,9FTY*"535MV;LI27ZPIJZ.*_9'O9P(X_HG7"O^?9^9L@_PD= 9S
P,6Z(-3N"EF96'<&S*!A9"4HH'LNI"\,C@,B;5D)A9?"'VA6I8?4+M<JV<4&LVK.,
PO7#,UT*DT7.,Z ;NXR"!(:SS?XP3O>6X]9;CAF=8&5VN:8^D;9T0FXT_6XR6B8TV
P6/JYY? ')6P"X'']9S71P<[!D( )?+'(I!L9H$!8VK8@50SX=]$>4(<<(+=(E++[
P$[TYX5@E:)]9IY:)DBSH<AW;&X*6?,0]:"N]XGF["H/;2V6?Y+4(.IC;-2;RI1S8
P/D^][[_W1CE99T,R-8"A3$^0^."S9X8-MJPS658)TV][(\JVR''*PV;&+%%I+WLJ
PK/9_)O3V6[.LLV"28O"1M_Z3+EC:+>;P%:M \06N??:ES;[ST/;+ W<X0#@E3@+*
PO!IYAJ(O^M8X_O,G#-IFN]A:K?P&.RB/G-;+@<NQE0/V*6V)EWF_#!$'I+($<&D&
P&%6\RMKJMC^SM_AZ\(QHR*08L76(Y\X+88;3MDOG(_AA8#@V]$5*\>"\>HS0L =R
PG,UQG5DY8BI78KZY7OL,G\C!K-I([5QDA9V8-W]A7;5X&?&'"N"0>?NOG8SW8CL 
P2NS[U(,S_"O1FLU%C8S8B.:IDMWK;656%Y<;E\20X# 8\#J*VXJGSF^=K;@B8J+Z
P&XFC74AL7,*G%V!DH4TV8"3V'2VQ#V8<L?BSKP\I,IWT,:MW]5 J&4XJ@34.=!VG
P.DL%ZW@,=D37]N&V(3>LIQM!;3'H53\$Y8H%>S-JO01"0J<4(Y'E=6H&./#=LOYQ
P[PFS=VS?1*5OM0BS_[,]&1/ ";+-:ELO-*YMBRP^5%#DOX?];;;@0T4_E9'6=2%M
P$PP+##)D%&8C.BXK_E1TVHD0#W?>#U77]H1U"1GU%R$<MZ*0"5KN2"!F$842 9V8
PUQ_2T"E;<H:Y@I)+Q;PX*-Q)\9K_LNN#SJ9PG7 \9O)#$(FDU$/HL78<']L'HCPR
PF_MF BM;]+N&@R!]$IG.HM:"+@B1OLS8QO \?7+,Y@N)&>DU3/@B*NR^X!AR+S9=
P=LO)NE@)<5[.#/(1OW'- A=#A ((JR?,UEI5I1.)7V_['\X?$.L?%ZN__7Q;V/I8
PX-8ZRF@4_CG0XF'0WC%KX5%R\Z6Y5"?K#F@Z'I&"V77?E\S<8&+9V35]_Y^@Y:&Q
P1\IOX#IBG@B2$8RJ_#(<]O>\#=MATUP:-I,/3_!,E%(,*095J<T2&.9U3. &Q2"2
P7C.D=M!W[4DWB]BXI@SYE[@<+(/Y]&)3([,&'549Z]_(ZR%?T,SH@IECL!00F*/?
P/"S2];7RU3*EDWB KZGQS<Y]VOOW7H5%Z:B.=!MK&P1NMD&/TU8L/\.$$.'AL#L[
PMC'E-2U",;FK!WQ*-,'&0UUT/2-K LHZ[$!SZ]W 77?@:@I6F!(T. *9V'4?#EV5
P\IDP8 $(AT1*[H7YA;\Q]7[DJG/A&]=0E>7SL2!<!*22U>S)%S"I(<U"BIN8VR59
PCV)5N$9+#D8TF6BP ;__JCM3^$PSV9:HE6OR*)Y:,Y:Z]T4LY<@CE)DG.7'#=FZ.
P,&8Y+F"@U1:8W1<#[&C%>.E]P7R.6A$SH(X-3RS]/R=;ZBP%%S#Z)'..7E\\1(W8
PD+*B%^:S5F9>>H;C!R@G"5/1E?XDDV@L^-G(3Q,( 3?\UGVJ"Y3R[<>.!VP-QB6&
PT,.[3[($/*%I)A[_)R28*@QY@,:Q9&Z,6[05PMPN1UY^[$DK6+,TU>T&&FAQ84M:
P\P\JO>-WV_C3$J6R>*/4R"%W3[UP\ ^\]JYRS9>+T0%,AUF/&7S>8!MPPP3MJ.I=
PTJ<F8#W(;QP%J]>,]^-7D$-%#$DE1J&AVVF045>5-7A2;#L;F4Q6%FH-V6GA"YY/
PQC<RX&X>56M7:$B&&3YK?FL><</N#KJ/&P@EJT0,'-\A@C=@R&'JP*QWS;E]=\-[
PFZ 6:EWSB_:25LZ.\45T+N],W1>V,QQU&SH&B:U;0J=M1O;.KX?##5]H(!ME+<*9
P)B/A\EN35[KUG);*,YYZ90Y3;._MS2YAC@6$BG_%G:F,%UA""0KC(/-W\!\L@KX&
P9P3C[_6MD0>0-]3':*421#EK.OS,W>4_YO(:""PCTY+(TKCH?XL47:)S7QO<@5$J
P(KPYS8*"'*3Z1 8,X.0,=$5MP]?:@^4]H*_W>_FV.CG9GI<4N%_5N_B[/_1W*-H:
P3BTZ#8#WZR "B)RX>.Q820T+S?N<BPYZQ;0D.X[A"T!XP5^?A'UWFIP>)4,[-,(W
P>O+8X%:^2"P^99ULLB&;KKTBY?:@FL7(8E*&%JL,.@L%L59;..KC.$T)5AOG]F\I
P,0H'DP-(%0\+#"P7#5FR^ABJ<:V*;A48Q3=6 2!51S$!J.;,B[II;ZPE+=:G\9I5
P?:ZLAR8,KO\V+N;!R$C?5:?L-80\V<% +(?Y2SR5+C12EE=(+TTSX-*EZU+L1RWK
P$2<:;,":]O'_U:O8-;X$,$@YG-5W*4RCOP'<J$KMA 4DU6PG.<,$811D*,AX!',$
PN'0P+M*C1+K8QOGA,, ;J$T2%[U:MTEQ,RVSO\":==V.1S6VUI$!-C\:PM^,=)<_
P@R+4+!R&)@:#%YTN8FYYM?JC<>Q*P/,5U3J:EXG:@5[4X.R=2N73,GA?_KZ-9[+)
PCF3I2W$.MJF:S/5SR=TS]HF#[4@'UXEMC'.9DG(Z"E>(U/I_<+A;NR>)\R=MHP94
PZ?H&C*)NN2\==;VI9@!3SY!H)N$L&L?722GC98P038_OR41GEV"0#P_''8"2K8[Y
P1Z^]*N?O<1!G-'*8-G6/DBEBIU5:7B$IG*Q#6&U[1;&5V!D-H/[);;K4&%*2MRK,
PU>U]PA,@[WLR/'(HSB/W>W9C>:KM(BZCQBUXP6ACH4UA#;N>/ !FEB,]\;5KP*T4
P_IC3Z+B=0,$NXY0FX&F**J93.@.ZW>0K2#R##Z$'(-!P(H_YG?LY/MW@= &8F/LG
P6G/,M3;>DG63D'=B[6HL>5K<[A5A')M_^C_EG]Z=C+AX5;OH>4 UMY2ZV3R[E([R
PD#H=5W7Q-.7)&GRN,<Y<.P>LND5?5+7JR? :X*E"CKP.V'-CB=N>CX-\IDUZWJY>
P9W[HN/U,<%)VE[6Q=+IRA4P<_#AC60N$HO. 1?0B5E@BP+H)19@!K&Z1BX+ @%[Y
PU9X27L;A'!79C=<KOVF8(%WO^>PW"!IVS*1P\NG%CA-@N=\K02](KZ.A3)X>804R
P%4E*<OOB+W;H>Z-Y!V"V(<[?E@OOJTF=_$O-N2&--Z)2JXL%V=46;#R-<_[U!PLB
PAC8B/WBYY]"3JB&D8!($82 FP^3=\[KZL06^:MEZ@-;L(Q7W:7YUE>XI$J4'<_EL
P2F6E6VZ _U.SGR?R^*REC0DH'0$.UD%H)\5P5";0\66[?AL$)UQ(NG0(W-XUK]^G
P$\I3XM0%RQ[-=(K&;"<QX,>*O04^LCLRC?-3R>H5-U]KEWQ'86S/X#>ROF ^A ,K
P_&*:WI8W(AJY+NRLA.]'!;TM6Y8C5_;*W[8/P!.PSKK]WV5$Z\738TW;B?25K0!$
PT,19R9GOV-/H2'(AH 7S;'+>5Q4%=]V0 O6Q'D$Z5'[*N]Y^&"7A 80B)A2NK]\$
P-+(B/ (AK+$KY)'VB2;V)"Y$B+]'<9H8NY+@X]5(OCG!/,?E>X&E$5?ED^LT.9]N
P%)_<P!4I<Z^^!MN)"TU[]&GNI7^0LD"Z4E1PAHF9QXQ9%PN:;H1MM/]*<>HOV/Y"
P1ZO0VW:^"@]^,YX[HCJ=?_O,8:E]SOY@/7J>[ /8#&-@T>=_ C+2N&<E(L!L*AK2
PH78#G/$QGODBF<[41F+4ZR-+UL#^-H8C6D\7Z!CYVD<:[A\SFAH6AI("^LWHWW7;
PS@9*H55(.B%Z", HC8FLK7!RM\]R8@,O]Y?]5C_!4;+%#MM8N&@NL6'%4/+K9GSA
P$=3Z9L76'6ZK*(PB5#[)*G\&(Q;BU3/6.D[?:.:U#H ME_>3DQ2"A2][M+.Z2M3"
PK>,DPNTG/MTJ#ZT?A+JH<&P]GN QW2R^>$'8^FB40%6?E?#254[M&IQ_+,PN>^"_
PPG7E:J$#WI\:3TW^4B8*-YR-E[<PC!Q$2Q4>.#_ ,$<5?5#Q <Y74%Y#1==Z92\3
P&\L[J3X$/=?1N?T\[I"SDSB*/OCQZE0*Q:?._>&[4I*4L#)2)HZ3P_*D;<ZUNSP.
P K<-"L5*C+L -F4K2I5<R]S);^ U@1RMP9)WNG?K(AN(8&]A&[KPI5,RO42Y7?_B
P(;0D[DG%5 / =!'5 %R5?*2GG*TE/X&R[_'JZIDJOK_'GLESHJ<F%G[XD;:;XRKX
PV?%#6(Y2\K-8["B'O'T3(9.E< 5HD PR+R_[>CYNY7\1P]8F#VXG^XWT#8;>:DN!
P'"!C5_,?9E3.45J&>GE[>>M]*H@GD]V9CA9LPV_."O/LL0VC[D#ID.TAI1R!U[. 
PP19YBHVH"G]#8%M/BT1&.',IR2R*K;7O'D@C EE(%'>ND=@@-#$*N%&7-NWP\UP%
P"TLQZ5\Z0VG6X^\W+MD:S?RR*EC6"O^Y8S^I86X_"E'()1N="P]OU+)CI23P;1,!
PULLEG^(YO;K!X@POR68 ?\HUU!)I<^XL\.OCM3==8<=HU+NMGE;6O@2,F(]X+[]S
P5D$]QS0_4;05O$>!5:/1F"[BU0524<]4<>'.Q\\7[EX/-^I$,1^9D EV"R\+,_0<
PQKR"&N/=R<M _$]G.5SNV7:'3!M.ZX>E1_;K*WP:T(G2LDCZ^3<1!!1R>@)6#J4Y
PGRR&V%55V*N^6Q19+E4&27+@CIQBQPOAML.N:Q;ULJ;;@@-C^6F1UE'QQAWMZ$)^
P?ED$=/#9]M_Q[5FB2CS3KQ..[H;$2'XMH[#Q'FQUYS419@I)R%)2\;B0>H(3QHM<
P?QH]0+A;ZR_9'?HJ8ZMV/+VE!!C:S^6$(B(PWJ):+T(<2H&D3Y;);X#LB^0&KQRS
P_EYY$UEV5(.)U4IW4!TXS-=6.<_*J[%>Q1OOM5*+Q M&GJQ?0/)E<BTZ+G.+<=K,
P]][$0C] 9*$F$"'?)MV9Q)3< ^N9&"93^M#(69 =MQ&^=?V;E99<A'XK_PN3]R34
PZ$W;9P9>E0ZG>H2K?+0LA6$:5GYX9^!=4N'9LH=/7?E/MCB84C6C7<LPS5;)%^F>
P)7+0>'<FM:=?[><9=[>U.#JN;/DP/D(B^1EH_)0PE)=N%A7:O&/7EVJ6 "I(Y9E7
P",;YL_256(:$.:#8>$RF'PR79[#?CUYQ4QH6=7Z)LX&(6'(PNRI-H$XL>7XD59\O
P-B:?93\(N^@" E\T/!U[#FSU?NF[80>'.(0[J@)30#D>!W!W,5D$NOJ(N_6 7BO:
P34/Y6NBSZ$(4)(_15VFS"CL9_$<W5'_2J<E)$4F4@Y7OH,3=)ZNYZ;\+BH)*66H4
P8M>W0('=I(YR3)G[YY@Y]A#WY%02D,@XVS7,U2@VNSNU%)S(40I*_X6_<K5SI+;6
PL-%:R ;%NX7!3K/?R?O> 3F>W!@5D@' ;3\WVK[3.;J@#=>@\,CZ;+)8DXX^@HWW
P73\N%(T&R:9CQR^@V"EUPPD1M29=O8P]I/(5M4GU;8QX2%V? A7B);#T-5F$605%
P5]W^LNSW:;RS(X\3_2DFD*PIF[>_\9B<BGU=)U>BP]?*%O\",Q5B)FO&"#?.:.@6
PAW;!NL*#]4IM&MA&UH,;P6/>B\;[@+E(2@ALK&W6K<PP1'I,#GSNZ?R2'\0%H_.!
PD)CR11OS0N<[" 93"R5<TQA-XEAD119E\V5+C Z%X];;3@X#L"KHK^>6V<Z_$HF*
P]G]'TU5I?0;S']/WX=I_%DB:WJ$#T'MS+!7FK!@\!XN9GO'1VAG2,YRT]?M,0)*_
P3>P2?&5 :#<24X,8?SBJ7E,S)?>TW)-4F^NKK^DLUU6D^%83:# 9?L?VO5T]]!QB
PK%N8F4B8.&J,/8J_CG)C^=M:^I[INSR<O9UJQ!$T?=]G6;K)74-_Z_ M9"F8?A]9
PJ'= I#9>")VC+ 2XR+P;*9<2+[6;_3UGZK41]3\68.-];+)RA&7W/6I<DILE-BO;
PW&Z;S"O0GHA58%0#:_SL]&4*BD'544J+27=I$-ZX0M\E%:R452MU&SA5.ZQ.,MAP
P)NOJ^5'KI\4,ZH+Y,">S71_G@2^^PAR,+6]22]?2R!CMHHZ!857$7G!2Y'$779;I
PN9,9^RSH^?WC7-',SS D7NKB7HI$QA,I2N;L8/M *Y1GM8^H<>0P;9*U,0IRY4RH
P/1FI.5]B3ZA25\J16,3<W"[R;EK4J!UL)!3JF]+=+JZ SA'M.9.^A=6IBHE[CFH!
PT.#;B3+:]M)2'^9>$F@DW#UQU*:G^Q3F_$NAM1OG0UE'[+BG3^<3'DS11$,VIYLH
P&@Z%<N$5^D)>)=? !,<WA76-3MR@OQAU O'9.ZJX-DIQG.[>;H\7_;W\HRCE2:Y9
P!K+A.\5.18:H/4X70XRYH=%AYD*$>=<3YBB*%1L6^!?[R*JX8NM,[3E;/1^<>$<K
P)&"IR:LY%9P=Q)6DNG@9.N2G@ZF:.TQ5 #:@9+8AM7//U\D:0^"5Z"HCV<+HF+S(
PN2ASN,O+>/B1M!%^?^>$L$[<OBA<V9BIIT ^A8>#R8S_0LZAH87CXG8DV,QP^7 F
P[/&AH#55)GE8?P$Y&5"8='J'!G6^,,X1Y@(]C@MEIE/*Z%)L!WYDZ]TV"O3HBB%>
PC7,NKT#9HGWN<ZZE&\4MTFI]E=NU&MQ9UH;; BMI)>)&47E&N<IMC,, F&J&SA)'
P2Q9V$HC9[=9]6F9KEB5Z*R/GI966/3]B($Y!:-SB SY8W<RL2?K^5DJ]&CS7W0NY
P(P"A&Y86'B%YM;WS1]A]NY8)P@5$P7B@M+?PFB\H"$I.@K[#4]5$,XY1&^0LJSF>
P"O]S6?^*8[KT8-7054/9%?B=4$*:F$;C)WR2;6I=L/GD?VR@57!J1[[O\SR=S/;8
PUVWQ4> 6$RNX[ !VY(/&DUM ]8@!WS$;3YKT[7 YIDMX_DY'/=Y-A!AOPR=0[%RL
P)3">)JD-K!4I3FL[>:]U]NW3^PN<;7USF<-C,;2Q-D]]9B+O426%":==K^MQD]5G
PT-JY$!DKDI=8<IRBSPC>#:^+B:\+] 9<PM?S_X!8 %.BV'T0+OH/-GI[*0P9_G,4
P'J=K,<G84X[,9+),\3\>,ED-2QEH9NHV2!+ZTT5#YRJ&#5P];=[NM:5I,RL05CJ?
P.(0.?)T=Y@H27G%_I1[FDU3L7.@K."+$9USK!1PS;/),:>7HXE\2>KR"'5M&R*3,
PJ9">K8J6!4E:&C;*E1-Z3;(:6@@Z2;^ :IGXS)0>CM'FHB;N^_N<!JF )#2VBFRN
PL0X,0C- S)CW"%O^](&7"J#D7(#<.:>+^U>U68(HW!7D:<@CPF9P<CR5CY#;UC8L
POZ=:, F*X-0O0%\SCF+T$UJLZ#T=+*7D#2D8:RN(^)2(LM9@\OL7"=GE'GB1QYT=
P5#('!41F$%B==L=>VMA  FP24QU9^UR,K!X_R3?\]PB:>LLREX2<J-]]* IRN9JN
PRMU4-^(OK)JY"2Y6>S0TM+A\%2Y("P3D9,YCF2G"6U*'0YY[=F62VMR+T>V%(Z_7
P6'([A&8/ %@^K?$\%]_&C?&AE K8.W QK>PB96P/5 WV%BEXJ'3VB<,$GHJ84>O3
P,!8=M:>!5[*3FF6+EK6&OK>BHNH>EL7!.1;\]P>*6Z<(4W$C:SA#%5K D>L!%@!?
P-%^MF6!<9!6N;&1-.+ =>7=7#<8"/-R@$E#8I7][*:*&#E U0"0\&L286YEK-7-$
P*/GSCA"5+1LOH?B6+EOL^_CZV\J!&DL-L1/X^GC$V$*98$!,4,B9&1&D-WD(#I7G
PW(M)HUU'9N:;_D5CO?P(A1@Z34!L.*JWCL=8$:=<Z*F$0OR[!C9V+^<4E"^,$J(@
P*IIT*WI35RV0)H#_D$-*#25&[_Z"J#X *D*?N8HZ&4__^>O<%>)?,/1@_^JGKO.J
P@R1-_P>6X CI]@]0Y(_B\D7/+7[&-OYC_'?)-4,TRJVXF[K=(F]6:DQ4MMD^(FR.
P!S8:F87#%>(KR]?1<-;\]SP2$\A4L%(;(?FISV['HGRB/9[783A-\4?'98\Q7"/W
P6 #PFW##DI216<> KEYR\"W]GC8AC?TH#J/VI)VG*VCUQ:4[I;/[O"/5^E$% :MF
PS3_85>'%%<6[0_BVQA*N\1#O44NR*U&4.;E<&>ZCU1H%[_O,88.7*=@@$]"_9'R]
PWP]ZI]=4(_DNLP6RM2\J.,G5A*@C',AINFUMGN]+$,>#^Q62D7KHB-8SX"4X,IB^
PKQD:,XWJX_VJ>'I;HM1WX]U5$>@R:OAV)T)O&C 1%G::;7Z^K!YP+]4SC4@845DW
P%38=+*C5M5_A0F@D1N"4>TPCM=%- $:/1P\-CU'F"\PHMEAD481@9J2S+^\84PYF
P9H2O2>I'=8#,M(:T[LT&R/SPB:R+<L5FHC'[CC=E;V]G-@"@@AGM+@,<P+6SZL&.
P*E:W!#U@^)(,!_P6AY:+')\EMU3(I=^<*MGI1K^]34GP\G,O#PQ3++Q'QA&\V4O\
P^/[&\YF^.R!\('V<0J#+'Z0:-E46N#3/L7S^@:Y$+QB-CYI9 _@2)VU>%QBJ>9^S
P2^=K3ZAX8=EJVE*L]8)R@ H[DMJ+[.Z:%I3H];P:\() 6/25)B"?HN2\JF!)Y3CK
PJ5*M(BI9JTB4%U2R[W1$2%.JXVVZ<L>Q((QC:5: ,&QGTS_7'+LPBBA16<9;WJ$E
PF.L7SZ$"5(!*B)' .).(I2:G )4MX!;[P[,4<X>A#L"MHN55-30''RU .(22G98#
PO)N"6D+[VDO9V1C"RS%;?T'8JTPC=41#G>2EG!ZAT,]NARJN<DKO0GY5T( 0A_* 
PM(YUN68\2OL+-',.-*>T@+J0MGBJJX?!I.%7_#>+]C$9*YA>1>2P2U:-W&U!CD!Y
P/XM-0GI,G1I:<)-) M$?3#(A*"W89Y:OJ+B;>.>3DX0YH%JG_: -QBRECBH"O_(^
P3;KAX&A8LNB1"A%0 _[X7=.QEWCP)XVY3?W(V'W?C+/@+0H)^#X+9I1C!DB^$[7R
P)0[SL((1Q E)B15))PI.$]>@L-QZ=\P$=;H+V@BY0!XY8SITR[9+'R=>#CVM.5I<
PYKL8IV8F:?,#DWR_1.)V3%K47\!NX[0K^6&H]]'=4R1KTJHXQ:#26.US<_<>F+2D
PRUV6ZCPV]:.&!39APM>8^+>1(X)I_*640=C9RQS6E/?4&P^B8O8_SLB=&("V[I"F
PWRE[G#ABJ4+]9WH%4])46A(& ,RXJ/ZE)2#NPEH[-S5L>3'X]R97,H;RZ5FHK+57
PLM0!U_ (\RF&V XQW+Y=D^^5>.NP]ZC M=Q(3L5$)J/14LR)[1RA54BM[#B6GLM8
P:F9.PY;KR1.8=]@5%UC-Q:_=QW:\.VYG2N\+O_>FO0X[;Y&?LH$@KL0A% H5AT,@
PJ6($V7R'X;RK"H_[AGI;BU6WL7TYT9K*.'H-"VZ@IH_WJO28M' \!S W#C/*2XMY
PM"VUZ1"25U(68% 8[[?A8:+<,]9YW4PUH78#%_?'LC%PE&#ZM,AZ8RL4I6+Q"J6Z
P\G74^\VHBP,M_<(^[]LD)GI(IDJ;"_3&^XF)KH;]K\*>6R0*G1M"*R*'>S':%/YX
P29 .-JH344",5]1<:J_970SHJX-OOM?U<")*[2;6GIBI7=']AXIP'='EN"9J2'A#
P-C:V9W&T/"W-8 U/C'/TB99+D9G[YUR&^O 6F^5#GY1279&:8E96-Z]$QSC_W'AM
P)82H:+_GY1_ =;/XQ#L(>9/:7<GN\ ._YF<#',;YZ+?-$5#07K[_Q1>"/?ZU:]QR
P)UT_Q?B^*69.$D<_W>DC/5MN;*%K("HP=?Q0'456EZG^:_E7E28FS*ZO5AE)>N5&
PC(9I 6AF&/(8JMVK"W/W*\B6YA(PO2'W-SYG?H;X -E_UOHURV]OY(+\I7K9TONX
P]!!DG/T<O_L5U:_T-Z<[[Z!R#N"&WT+GVB93%QC*T$.&3V 3&(M\,7*-'7%*@,X_
PB-&M@RA?=CS96?/*:UO.M/H TY&J<]:=YKO-O,Z+.32;KV2+](',ID^@LJ:F5V4J
PM7FV7]];?Z3>Z#WVQW //&ZF(<<G;#8U72*;.7<<NYY7@)W17IF]5$ X6%<OG1Z"
P"OSMQ&L)]54W$Z1$DBK^[[KF8GAY8[9Q"3?7Y?4J< C)N5V)W>^UW&4]E NFV>Y;
PC% \7<1 *1I99Q[%D+T>RK)L#M([;%@U4H>>G/ZJ^2F^!]*'%$[0)D:3KLS&9M0 
P_LG*(^9X('MJ>D4@7-U2P^(FODW V7 A]U=40=;P"%3A0=</WN@GDC46?,N8)[Y'
PM3PG+=\ISIS@%^+\M/[3J[S6"&_R34;BYYTA!-&! ?\^_UN]\H*M5'!IKF%UK;PT
PG#=*[R+I$QI IB&K\M91UY;Y2Q_U:<S%=)H;09'1.//="E2R\K1T"F *Y>FH=3$Q
PK7C(KQ^TZ5.H $7RSFJ%><\K_X-+YFNF:6R>'[AIF6B!>82%@C:O%H'ALO[Y(12]
P@A3MV%0;3$OM:YE:[B=41NK*OT^@<\C!(2XK'GDCN[856$=+G]RNT<?29>)15RN4
P"H'71*F\W04)OF96Z-U@?_9*;BMG4.7]Y)0=!',+(G8JV'7 2WZO5WI2@\ NN:2/
P$TH<U61PJQ*O"8;,T;^X1&O6,G^S_$*T$M5P\IX%<$I;"3+Y T.N74^YY<+45F.X
P\+,L'FUH2_%IFSRT&I#>W5<ZLT!1Y(\4YK@%2Y.;9BJ_V"-]JN'+O'&%>& 7K1=5
PO2X!8CQ+6.>&0R1#N(3_GT]U;)CBP'I./, <"Y]SS+_+^4UOB%9%;,PIUM#UH3D&
PJF@+$;$.Y$)X];8/:M>0.Q![I.:,3.$UNY9(QI?@]P>":[^EQ!6)?=_9?RSD" /Z
P-/Y.:[$&_'@P%K!@/E#/-H /Q4_%^1+G.207X2Q=]2:#+HQB)MH[L_<NY_5_##19
P2E854(+FTN7BV#1I+K#3;9;Z.HJ:0'E-UTD3"FZ*EMLH4H%M_FQ15:^W"NKEB1=J
PO&+GB6S,(R\A=4Y53ID=Z6<TS2%RK^VWRCB&S+2)W DE0TUI.8/:1;@,R9.$%&+'
PG&3CK4+@CE5WJ0,F X; .::P2UAA.-PH4[A*H37E><4$JL:H'62XC_B@\67_U)N6
P.U@H5+Z"PV6QZ_5$)C1)0:.%!>E'H"3#C!M8>J= O2VWP/B"MW4A*;5W/)':)(9!
P4=EE!;/O@RLL>8UY4NH\#RFHE5#CG*#6E*B(.;(15X)OV$L;H]913H458@^1T0(J
P]-@R^O;W$?WCWWY^2#U5F#FB7"1UFJ;#2M]*<Y<M.K9G1_ZL6+3/R-3TT$/1,O97
P4<_[=\3*?^$H=(6:G(F$["6B['T3@(;$RLPWNGR)A[_>H)*A^EPF343+OE9QR23;
PM&LAQ03UW_7"0E)/W:<L[8H1!<X-Z%%X&.6R-^Z)/R%[DG=WO3-Q/#_47T0W7=/U
PI/ETQW%?'?2 B&&P'OK>!HH1YI]FP_,. D<!JA:ISRO46&0YR'V)RP[_Q31($\T-
P<@-35'6==9IB"X/E<K :.@M$I_*-]>B+E8WU\.-(EO>F6)&0[??E" '63&>0?PM0
P,Z1\.!!UCJAQF49Z^6- 6.L@;8NQ:@G<@8Q<(1?T4>H:\LL>649=IE=;=) ^/Y1<
PXV[\9)@J=JXMK6Y5;5;->K$<!*6-9@R.BT0A_ZTY2WA3NW<:/UH;UPJ0>,AUW%%Y
PD()-I93'&5#;W]1#-JF0L$>)/'*HZ9-WU9JI;G&9D&4_H:Y#4& 6T^G2)&#H6L5A
P:K=]4W1LFGO]>SA&].MV/$L#:NA54*"*^%1DB*0(O!=K&G)@UPYQ(;[J)MR=EI@G
PX/R'76/X=O<4PA]N8MAF$113,QPM'@!5\:P-/Q^I"*RB12214QO,D7',*T><@<<M
P=RHNN31"0."N=6EZUVR[/>GN0J^S!,/^_L$-%)-4*;2-UTZ[[@JA2+T+7';E>[/3
P7Z,H'#*I+NVPD1]QT)VK71G$UHQ+VAIJ#2TNOM/5=[\B<S-UR\-U=%2\+<8)R-71
PFG7)/_J5C,17$-N8:-.Y#?$N7ON*B\2[@PM9*4+OWBK,=@*=7^:Q^37=G@+D[:9D
PM^AC2D_B'NRH,H2EJN;8,N1Z"]F\#,-,RVVTI_8-J/^KSE;T5K(*'"FV][[+O=/V
P4NQ\M KF<XS(_& !(1"N?0:0ZJ]0$']K%3:"?)6^>1^15-UUJ*2S8AW29/)DU]8N
PT73J/9[L(Y=BW92^#G6W?KNG\37,W\%H8.-HS6.1B::*OAGX6]-BR:S-];)-N;F,
P)G%>(BB%RZY47JG_P#'QZ/,"T,C)D!35\5*#JJU\^MLIBVZ]^&T1G8)&<>" H&XV
P?)/BV.[ 1D"PV 3#3/VF##;GUIS1Q_'('_J8 ;^#2[,S[0]U7&2J=8' ["22 C&&
P<D!DP><L>\5%R<&&Z*2M=^(3KU[@O]4D+M>8 ;$O,N^?:#LRRV"%37\B;#TH^39Y
P:0C#QPU<TQI9\#E*425L)=B%?4L8L1['[B=_V[FDSRW,AW^,YP,&__U!@VVD#/DD
PRWO14@/:<^A>Z,?=W]B:7Y%2BI\:;)\&O_B:#^E19(7A59KZT:AG N"(55[X::[S
POAZXL+H'QT'O1;0RE$IT!I$1Z!^>%) SE%NUS0S^R=Q\*\P;76_TU+8BY^'Y)\%6
PLK!YVM3'.'"6-XY_IF!U5T0FZK+X'[Y(7L%^W&S&4^SP-3&JNBK1"6P7^C9BKRII
PE7<!(MRT^0:[W312S?8CK 'Y'OBH-/E].*,T^D'>DQS8#<I2\B\RQ6^#G6\K1$L-
P*JM[>"H+U%)W)XNX? RL_>B)Q_A?O_8;#9Y_5&CX#!WLQA%"N,;Q1M;$N\=<=5/9
P8E4X&_,DJ0;^!W]OC+MEY*=K@H_$S,M[FH.HMF[96BE**>)H:S:EIXY0=)^7+W+F
P3$'&Z7W4(,WV#,O<*4=$46#S1W)_)--VE5-(2+:-?M7T8U(E^U]*^@O!!+K$X+:0
P)DK7&/X:_EQ%'$/<F-9G.?:<+D,<1_%9<#B-WRLV3[D<Z4[M&B_Q_%QG\88D;1>J
PC;+/JWA2($+V6QET2XE-!YZ._>*DI -I-O80T>=8>][]TCKJAQ [X8TYB10AOBA$
P291RZNF?( &20%^TR^Z-P[D"-\3*PA*M636HB]\/MYOGQ\"J:?;]B@T(")K_5I5D
PZ$DP7L7/&")**I_1B(XW;'- \8KM^_2Q@?C(V,Z;)@C;T'QDC((%B;%TZV2H-G,$
P^/K"X^RQM:0]XYKG^TE(SN'':XT:(Q]2:R6]*P%G??&K/G;:I11UWGS<,\WXS-T@
P& 9GL_(^T#M^>61,75<)N,(M<V&2A=( <;B0T#17C+Q995*!\M,4@*1FK-Q<:1_S
PTP2 MOI83>@2(,*D\MC&L=,.@B C+HGC-ZG,1\BM/+N1>:@8P9:LW7.M2#K-,@)Q
PR4;/[L"TXCR5<?;^;D+5J6U '28<L6&;$G@2 ]H,1--LR,[[L;(_Z^.A!Q;V9NC3
P?C)4=E(F%B8OU3>)XC>TUKKTOLU*P<88&0OMZ2/8XT_9AK*2/M[P?F-OWVO[K?+Z
P^!4D<@]+\=5\^T346R)E76J^'XS'MW-R(XG<T?TFC'<4:$PM'37^,DLPE*<KD<@#
P7>#D/;F>F4#(H.82G._EH]L\; O$#3X;@Z%_#1CVX'>/4<_4;DN8LW 0@V#^T<A_
P*</E%=?"NL0.'_0$!8MCW# /FV'WNKH4<$C$(Y:=]6A.'P?'E&"Q.TZZ?G;O:+=*
PF(QDJJ7J$%'(KK$$\^5?JOBV?-1)S#5_R%?\P)&P 35<QMTG0N*0:-;,+6)^W:T$
PXC'T6YU+Y2HS.DX6/2(2N LN]MTB<OIU4F=O8VJ0ATG<I3S9::P00R@8M)X#ML;H
PS&_QZT>B$H66JT458UOKS0GW,T =*9&4@-(M4YI)Z:VN+2.9B+W.8YR^0X:;#C)1
P%*:V$'\207.+VR?;$;,IIM)6_BB/CD%0&G&R(41IEL O#-P+)R"PRL<-O5@* Z,;
P;5<.V2T)>WD[1+QF@97FH+./S=S+VFYZAU!IDS'X1I>P4W!VQ] XDFOZWBE#=G:N
P$F 8^:FZ%I+K_H;[G] FY,URNI\+,AC_-:D,CI%7F@JM$-3W;(PSSHIK9.(AVA!,
P,EAZNU"#CF2HS+L:7^ QY!F>FD]) XIS.RA-": /1AP-Y(]_1I((;'6=^(I516VK
PF$80%>?Z,^)((\M7JFE;OM'?W*?B=>4SP2B30<R+=:K6FS2^!#BSB.+X+ 6U0YXE
P?:KE.>><DV\+$AHLC.( %P8WVZC%RT3XY+=4'$WX/A6 +RGLE[:<=[>F,B"S*6O6
P-9NK5!PG-0$XCI%+S(V1-K!.W(@*5MT^BU]7RR/AA/FN"NAU5=JV#0KDL6K>T8D0
P6P[#&!9(V-*?J!6QOR"B^NHX(;CU%BF%E_%=+M&HQ[CFLT-8>6^[0 -,+#P=,I5 
P20MFU).S]:2:V*Y)X]Z(V1(-+Y"O;;BJ.XR8F/^\>]8X\=!30?$ASFW+JPC9-0:%
P<D:\ L<J0'PP+CC.%\P+X)DRT\N]=B>?1MMC]F3'UD*\\7J;72MJ/;N84*%\\E*;
P<<,YQ.Y^8^6.-$C=#!]3S=M[2^YO:DQ59,6&S3R+%.*;B$XUN -MA9H*C]],1H<9
P*US@)76$+OV/,<Q.P"=41 0DG_>!O%% 5%7,<H$ZN)!F/%?B5V]U,+6M5>$)N[0_
PDM ANY-^RF2W'I_)0W+N-8$T=(MAU>7D0;4ZUPGSCTP#.S&F6U#DZ GAS?@32\L 
P$VGY7':@YJ-50]GJ,)!JZRT/;H JY$7+W]YYQ<YX)H,C+=&M!)LK>#>+VSC*L1?)
PC!W@&IY=WT<]]<"[.TQ;D^96XC RI4S9<G=FVHH5S>OGLD5?"W<S5$]?5/OJ<M8J
P/)$_J.$9B%XOKZP(1MR$^@K,#*M:%1HNLS9',:="-CG\'!XLF52O,0F:A)]'2;^5
PYQUEV1.JZ?Z3RAH-<>3JZV8-F=NV_-+4^@_-0U>Z").<N_8R_W62+:98B^IMEH4C
P <3EUX?=90L?!<0]_QG9]43\@HI&US\;G6XSGGR294>,<"AWM# :E3&QRS.8=]B5
P_C]Q_A4N?_LH80A'G])Z8(6\JYT75H,9T[?;.F)0"AB<?P%[X,Z^>;/!1HCL]],O
PU0#Q9VL]J869QOB"L]*#%8&W5HW2_A(#WG.E@F\$RS@?%P'6RQT7DLJ0K01KXX>D
PG['8/N1=2$H$'?-J*E)^ 1]C5Y:F@KL#UPAK47/(?M,O*(4N]ZU:HEA@Q'<PMJ&W
PMRJ]V^)WQ#O0ILQ_"8+;]<Y9%4FC'HI5ZRH[I:;U;<NV#= (@\('T?.@BNBQ7(:Y
P;D4PJHL@IM:)](%R$0#TRJ=H_H^/_%]>%UA5TQ.TXQ!_)O6=B23G*Q^L"K)3SR^:
P#$_^8\&& NP[5E!7"EW!?RNKHX'S! +0-G2TD?.M]+W#FXBF.]A;A[/E=27RNYPF
P>/^U,O&:>&W.4I V:GQJ!BSZ*R6V-025RCZ#BWC3SHZJ3#9ZQBEXZCP.X#;/X7\%
P0X2'/4AN,ILY+1Q%[R[D9X*:1"S7H6X!EGUMRA[."G<4^9VD3 W20RJW^)6E$,#I
PD[ ]$WAF9NBRX@L;RG+MDZ:Z1!Z3E54KZMS),T!2*XW/]58PL4T!O'I0:LCY0=UQ
PQ+Q@-5HK5R_5)YPENI\??=/^,^9RQ)[H #$)6TB$9:SWF[@EYOL/L27ZB^Y>N%3K
P<Z8F #:7YK*<7D9[_Y M>_&<2%2+CEEXFB3TA+F_P)>G\5N(*K'*,GG(; IN(HO?
P?4G:(IAZ=)))65*!#BU)&Z#87M@>@ A*1T?:44V "RR'6JDDT8$HG<[<'[L9DG4\
P5AN:)"0"-<4(JTHN=)VO/6$C]:B&&Y"LQ+[25"8TX8;B#RN;RZN\NF!O%KN HR,R
PON(]0@X,0C!G65RW<W'SW9JC5ZP=F5)V P3"G)PZM"<@+#_^LK(:,=@C=_-3-D.&
P@->(LH-H4 \,XVUI%">_5:C QT:!0(8XJK*^Z-KWR7B*@S,_37ZO\!-<?D@69(XP
PT$(!,VJI?&%*JD=5UJ?!O#ITNUP613FG0&2E"7]&2/A&!\&%J9<L,%C\"M!&4.^O
P+EZH[(2I1]6QNG991F1=UJ)<XDW<G;>"/]8,]O6YLFQ"5!'TE0"C9A6N!?8"V[Z:
P2;@EU]OZ3-1HO^_>*),P[2[W%K:4V_:I.-&<\L.P#]<_I(&J=$<DCOP0SKN/5$P/
P\['3X<!@'0ZN)"43,N[]UI&(&Y3P0'\PN9G.'6023T$;8H0;.KGT4MDMX0[($Q\&
PB7SF.I"<%*>_-R(30SSOS?T8<]*N?TM@KI\K(9B#%.ID-DY=9N/\0*=''7BG6.&S
PE/S]&JI?NH>U+I_7(:JF2P1&4O?,GMPO*M71\AP(C_W/> H7SIDU'VS:;A>E-$X=
PT&LQ\5NUWB=3_\%WMS+$Q-XGERZG1<B4).M1I+9_9".Q^*;\?26VY,?G3SVQ##K;
P-L2_?*GM8,$V"BSGA2_919,S&N.U1@PT2'4:K&"'ORDF!XO%[<U'8+(%^D:ZZF.J
P"99WBWUIP*^.N27B0!(GV ,<#2'U.4%\]I#0;6T3["*X%7D\4,$4-MPL]D@=)?K.
PD.,RKA.6-,K'83X]^4,6('&6OC+R]/TQ/Q9J-G@!SIY-/J-',]?BIV'*MLQY/:*&
PF9O\YZ+4_YSD_\5"91<K22/EH$ Y>F;\KN,N:)T>B0( :%*H=+%#/: )-3GH>Z @
PRG0=&4*Y6[\JK&Z?19%\'Q=5TYINW]YV&QMNOR \<5D,(_H5F=DM.B4X'7\VKC1A
P,;76H\=0]PTH_+_9EG+7OJ@<=2HWHY86_:0?(3KPHM6I"]U 4[L#&=?2.>]\PUM_
PA6U?<NXZ2W083Y5QB(HE@*JA4"7+_&OW1MO(V8O=:O8L9M*&IFE&B+NDE5E[QO9M
P_"?E"R^R?7::&8 W3Z36I.B(?1*#>.Y.+.0UK6\^)I%#47Q"!A_'$+8OFU.*'JJU
P>2+[4-!N\4Q,6L\O9TO*"-<0L/U45,IGWX)Z ]]_<DG+^++>9R!RG12^FUL(2Q&'
P3?$/8F<TPMI*$&I2K;%:WM.W,RI)Q# I.7K!]V:/'W58HIGC;HB*'&0 ""NW5"@.
PUY"/&3J&/F7\9NJG<7++7<3R>8D=3'<A$X#J;DS!4JO\ME>[($5T+(R&6"Y$/8%W
PQ=+3_G]QJ&O+=.,P%!YQW3-LJ(.P#.48)DH::&F!3(FNZ1E?-NS&8&2$@;GIB<VM
P\6!1DS JYY)X]U?^*L\Y%T%H+0ZA9%+):% >$=A_;QS1 ^AS;1Y*>$'R@+W@,L3!
P:/7)(Q^3=IW4QEEY7+VE4VK:PKU!U3@$%]4M028\_.D.1S$TOQOB1:NY#U[!:7B,
PA3+N/V]9_Z7W:=7.TJ+PIR6-;:?24@%SG=3 GO6H''.A(U8012OM;_;]V)<UX<HN
P*:Q>0\M0)$';)67;+F?7YC#_<T%Z,_ND"C7&Y,=7GF/Q9!", [W'].Y7?!/4_-VS
PT1DCT"\F)<#&9A=WSR,N!CG2VW:XU@4=[VHK>JF!FNNA[#UY!(*=*+V(<-BB/FU]
P]ET1C,CW^YE5S)PM:YX/'((K#." 4G"GPE'A8!VDJ4#27&$&EK ]^#@?"<5'D/1'
P/)Q9I_^3@6XSSV[6ML]Z<*)3 Y<C*0;PC#_%9IY;*B4/.XHEE^2Q[5>XI;Y$$FQS
P*,S6/KPENEB=Q)OY/,A;N+$1+HC\;NH4''+"@W,3:=+6,8]UJS?WC-;RBH#YKE[R
P/.P2UVHSIHY!L?UBRG$E:3,9QH,/5^3KBIE&H-QBC#:=9&#(F@\M>DX$_=(5"S_7
P0]'9=MZ9$6>AG2;#?65VN8!.10W_JV*5D'C;.*@1/J%E'[IP<Y'6^MGR^3M!!P9;
P]>)TBD5OVR[Q3XX6KZ)KPI@4W>>:F[3^+BF'D>%)@5BRR^#;U35.0B>?U 4;KY5W
P1YF.'*:)KIYY7CWB1J"2U8-GRJ-TU 1UZ!XW6S+_WKX&M\Y"L.:WP)51]1<,M[5H
P,N:PI3BDO#'[BEPR:3;5"?/\[#*$JS<8US=/(IFUW)+4B!P9RW"A. $@,TL>[Q$6
PNBE<6$8"0\4F/8Y1L[_ZKGGDMO9B$05>N=2T8$3?*MWI*N@AW>T,N(Q#RGK0D1@O
P1IUF?JKGKY3+K1O8I?_6O[6+A[("(Q70765LX-;TX^]_0?MAO,WN I155-SG_W(@
P7[JI1Z$R3H.Q@.>0 PP2A2Y_\8\S48Y6-ZMA= !BZ.*\,8MFX6>2+(.O1@HW?6U-
PLP9W1M!_Q\]#"M@4JD_>A5&R/>!19Y^XDN+DZQJ;%\?BF;+-)P<)2PB87DSA$L6Z
PFI>)+A'P&[I&(U5@ BC&JD(?-;HIR'+)$.CPT);F9*>G\I0SNAG,;7#FIEQQ* \+
P&6H3MI&MB$WC\UY 4^"D_ 0VXXI^^49E)'!1<@K81=$?*+_>O .!M_"%*QQ!0;2_
P6J4S7^0]DA:D'2?9&L"H9X;H8RB&0_D LU2[IXGE<CRRI!1'21B&\]EU='2TIA^9
P%GTV/*J9*)3ZA[.)K%G2*5>WJI&AK83 %UJK!6J14.<4G&7K9QR^"L>YAU0P7WXU
PPE#F6VSX73NKTDMOW$;JT\.:@&^@OVQL-+9Z=&R9X:5]5_CLCU>J*3+5C*.2.XO\
P]>/;R ?][ES4']@CO^T$8"XS<\PJTQ</(Y@4-Y3CT8TS/PJ8LE[):?1=GDVFK2XS
PS@>"^W4!01L>RSD0X2)05<=S5*[&\?'%!FJT9!6Y'M$,OSXA6S3\0)WU+@'6!'_>
PQ T95<'2R7,0YPYMDO%+&^"N+@W_P=7GC3VL;;TV]8U!63P9;HU!BX0H@&N!"L:!
P+;8"Y=4F@CP@M-0/X@#^K\SUYUQO;@R*,)N(!VS3L!?3D^\P%6*R,G3J'5\6K/[*
PD1RSBTP*5?J>B1^J $ 4<=8P+4$HP/'@.$BF7&+DJH'[&D+1@1&0-M3&@: JXC_=
PC?U'N(<&_DM8(\;#!^VP2X^1] ,\OF-&A7Y)=C<OIW]JF5ZY+-CF@O&67I0,9U.:
P"@CD(:HX>PQ.+(P"0$;MMZ5&9P/\MI1N,I%PT2X!NQZH(%4P7&AG>#C$49\7D7@G
POOP,;D"L?/@/H?6 F]M$8A/>3V9T>Y"J2I5R>L=D6K4=:"PH G2K C-3X]="/)22
P\/<>@D T7Q@R'(XB#['A\QZR$E_]]C^8S^BRAMXUI.%:'QO&*U\-("Z\^\Z(>9]$
P[(Z:U]GPB(]<]7*@!*?^@6FY]J!Q_NR6_*)=?&#^HDAM1+0NXQU]/E6</-9 _97M
PD#X>F,E?(3#6X.NK8X>BO1MF989OFIR9I'U>0E$#K(,DY*5JPD2A>H;-VEYU=3>-
P;1R1\VQH!BF!)WNQIWDZE1KH*\Z?D<&(\[M&STD ]@L@P:/MANHD(?,ZFE)V#MWV
PI*,\N<I"9@!%U N59@?@"H8FQ+%+O^K/XUF\X_0.(45P@"$J*Y-Q;R%<R\]73WK7
P+M,4F$CX.WD!Q-2N4D+X^ A;2E_"5P(ACAX@N8)KH#%R+?E_>2>@Y21VX=%Q8O!)
P2:R0.S138NQ;G>$'5C&N? JC"^_QL6#/F".4'OI_V^D9O^$<G=<0-$0I^SU]42[V
P=!H;4LL[T<,;.#6NOW\AB+GGZR12N&\'0:FZJBF[0S@4:U@PGA8X%0)D(LBD 1>,
P/J_&HQHY@]R^(JA7FH_^T2X^]N9\YLPN_ T#YM3RQ6?N)'.K@TV$0U#7LPJJO^06
PP*U0>? %R82,?CML5<D4$..Y@H>$' 11*"\ 1+C(?/91J9V.JKYLZ=(1/%0>L*= 
P<87R*T^_($V=.Y<@R![90"L\1:K!H!$.2%*2*W$M3T7W>"TMX=&:Y;.ALT3S[9S>
P["+I-O(QUA(6^9@ Q<[70$K5+W0GHWV\Z6'*AN51!W4ITUU-V_V[&P$4!T# ]%GW
P;G7M GE*\GWE7HZ_AE8>Q2G$)A9 VFC4K_M6=OGCH-+_ 'A&U[,*\"DMUULS)&D3
P4(XH+] QR><6J/I+0FP5=W*PU8P#_6+W@T#J-HERDNSM:CSX2,Q^@VX+%#>)'OCF
P776E5K^#7.Q)<^NAT5N%RX]#I4NW:+3N-_P*%!,U,Y%48[@>$F%VZZ#\ @IE[9B!
P\K)^QWJ=I3$*#<>BF]J$T32V3EWI%"8 31'X?"+9+-;!-)L\#[IOGJ(J9\+>OO+R
P&#6L\X=]IAU*&H1)@QA[@<GW6*H?-"56<=+XN1D'MGX])<DFQCTKWK/B]GH;#$-0
P\0?Q% @XV(FEUV>'!= [=)!5X1$^(F""RE")GD*Y,J701OQIAQ<%7>0]>^QXJ6O&
P/Q?QW;-^Z_D1IW1A[-EVY%ZK5>KK6_>T%\19O3I%<B #R_IVI2Q&(<&Z'_K_7B+?
PTKFRQX0U2TF>Z&M[5AFXCGB?HAR W9@L!DE) %!)CQ/O7?ZSIV*#&KXO>J+4+6IT
P6%4[[-HL$ZIW.5HMQTEU(K(YBEE$O::?[,X]9 =J0(Y4>Z@4<" 7E:IQ0/U&1?$J
P5_G:8<:R.=,*%RD?A+OU"Y/?(SM ;B^9BN::[;Q7&[5ZQR,IYQL.YY=&SM4UM!?3
P/SI1IRQL"":YK-D-,VE&?&MRZ;E/I)<P#0ZQU^!T7JJCE?RPZ!HO>-%8L*E&K+9.
P2ZD 1YG>,N*[6D^-F0Q4NC($B)-$ Q9B8Y_K,5'JTL@6(;UI[\51>\41C-.@K\-T
PA\Q,3?F%[@5**THGRME(#$)YR'S4%WE2B*BHQ,OS=5SCI69IQ$D@"I 4_1'/$,IM
P!"%CXU%R9Q/57^>!NXJ$&8X-HA$_(;75TJQ7/$,SYCRQ4NO8JY0[XK[[$1+.2L5<
PB>&7L"E4RR'"AB=&GW]D^'[AEQ1'PP/HE-$/9'-WQ(FFVO:+*U43"1\M"(SUM#*$
P_:CK.B[R.\4: 2A8!3ZDPJC:M829KM)!&OF(&2Y14*'W.3"RUD^67.^U1H@6#Y0F
PR8R(.@I"M@7"G361Q[\ODN66MJIVSCAJ!W22]7?STG-_0"W/#S)?%+B9Y7N2CP]J
PK])R<K* =]C5!+)WQ+P* 8W\NR,P+QDT2UC9@^.\>^D7#"<O$VB=C0&N\)>3RLLP
P@&WPIAHH(.J <_K_.$(B+C:L1X9C)U[XRZA,/@.07=%><.C9CM RO(DR22)E(1RD
PN'.#)PR8<!E[X[AO!F L 8T8F-;EU]NM1FI;9NJT1H1^$2C7)**]3QAU,4B&2]$T
PR-4*5@OWM0/FR.<LG_$Z>V,+:4STQS91D86''-R;H6T%'"Q#_-XZ-T.?S-/F-Y&'
P"ZQ**+SM 0-%EAC"='<-+TMA'-/IK>+*.NY%!EFBK?)'O2;"K:1HF?DAMKEH(^;O
P%"5$A#8G0/LA'EIZ+RS]#M;%7C.:?#@1QLNS]^BOSDXJ6G$G!8")*[,KRY[,H:$X
PB:J=[RLQ17E;O3 @E0H8Z;T4;6^BGKEQET90\8Z@+17U>=W&6@L?>&A$W';7C2+R
PVX3@G5F=  S[U:[JR2J,(RZI.J$RJ3F_=:&@'F=!S!*07^^GEY;:29HUHX7) "^(
P!Q3 %_!;20%-JFU[+12D[1V^HW6''9#/_\ 2>(HQ2>9:@V+5<A#7F^L+DHTEJT8_
PF"=ML-5K*/9H:7U1R.Q=,H-AA6>*/*/*,'L A*'(H?-'Q:S8>+OIQ^,0#;J,AQMN
PU7]FU=X)RP6.P\350.>J-$K\LJ9 -VY8XZZ 4IFSX"3)JOR8%(I,W]V,&$ERK*+1
P:5J'6:/+5 [O6\U1BL@(UWLB=Z*IS#@W[J\@UM^62<-3V=_1:C?RKZR[6-QK/Y5W
P\SE8;]CAG7.K:_B/</[*$Y"++3X]-1"YX>"^FN5.]0__AYV8,8WRU@8"+AQ)TCG:
P]]R8ZF@L*<85@Q@V!$>&2+)T0W=7;Q-1; LE'XM2J_A.1K7AYT9N^N<#IQYE%(8,
PV2\LP.Z2L*M[<8X/]H%9.?0TQ7 +_@Y#:.J(=!C+FU,JHH/50^^ ODQC8HW/D%2Y
P4FI"9]K[H-XM[1#A2&'Y+!8+Y)]04?#U"D ^F=.L]]HQ>7D>DNAM3D?F6^@M:+LA
P5NJ*PLQ[F]>"_^U=9H9)OT2O).(&]OZ&=]0Q_Y8["E6^(&NB:J4FJ%6+))LUY3F.
P^2<<B_@'Y6P"KE.VZG0,MA(8=&,W;Q:$^)+MBRN\.-#%%_ WG5:)M1#AN3TW#V K
P@U>PBC.,B=4^96E#^LB!,K(CJN@VN.Y?8(5LXZ=M[<21'1[^N\C73"!#AT=#2^_4
P$8':.X!WNQJ6S8U_?GZ^"A>\*T]2/F[6/!G\MLJI4X2 :LM4#.MV^-#*!@UCM+=0
P=#VBE;-X&]HKB_+7CE-T1VL<K=+1[:!M713JR+XCE0G3"*9-\#N;"1;7=-6R90L'
P>SA3S[<R=B$WS0]V*/8RRD9&%6]M/,(ZA.+IT12U-P&_H&:#7428M-A,HVXY1?SZ
PUP4I*;^^+NDTCZ5!G$6JAD:P3W9FB $]ZA)_\I!.6\BH%^& F=G*IB42\:>R/2\P
P[/3N(ZG$S_N=)9.E/IRFA9%=7";=+R,:(,Y\&KYWSC3T\'A-YFCLT*T><'HVFEM(
P20U")/QX-6CK?PH^,:?)9_7#N,A19()5+A7MQO03_"X6L(?^ ;9NPRI$(KS64QF#
P<DG.TM2?__6>YUZJ'Y J61QK"LDICC/! $S-HKDV>P4?\,!I 69Q&;D0Q0=>96XK
PL__8TC5WPR[\]D4'+!YJ/KQ99K0?ZYD'](6  4< I!16O"SX/[F6MZ0V_C+@"L&,
PX\E+OL4#<E<8FE"TO(Q,@UFQJ)U/+TC_&3#PJI"OO*$,V- "U!(#DSAA17<5*^D]
PPE]Q"SV28V@FEEG$9Q5R5HC!U^/8C9P'-1EC(%E\!(E7.4>(I>J)[C17J>N7X'8L
PGL\R%]Q48WB=W5H1)B6JF/,C-%>%':,AQG3^A+DMT5IPS:Q6-Z'QHRR0P^BF4&S 
P&[!PYR51@M@X@S3<G$6U<G,@<((U9\H84FLR&@W52H* N/<ZC3^.YR>ZB$Y\'3Q'
PFYMN*D0,1"&9K<#?SY-921DNJ&_G!@!!G+PILXR(9DQM'FWM"6B9&FVKNP0N\RA 
P![C?7#;;CNQ0@ZFND=IG&?JKFH=[(+[-S%*_3,MJ*G.LJ<SKE2I.\; OZ='H  3X
PD2>VV4R@(VK-"87C<OUN+YN81[=+(5O7-*#L-J1K^H6"; DDTTM*Q!)"WB'VC,9^
PN]T4:'L2TGMA^<J=H.R>XJ*=C=S#VI,%%-\)P/NR^]$@FH*9MS4 !_EWD-DH21]S
PEKJ/KLS<RR\@2ERS?_4M][CK2BZ9CUAXQ0 G1C3>!J!^WHZB/R-'LG6BONN+L@PS
P2!1Z>RNOAD3GO^+!G!@0*!H.*NT_K&CS"!G!_2*GI"<O[S)[^#Y>[69(E(!J>-/(
PMCTG-G.3B :J,ZS5RT<W/4=DEL@]"%O6VTD-3U =WD%M]S8ZD&JFZ"Q\$C*>"W%V
P92ITX-.@V,RU0D$4]GD25\31Z;VR?YNU.]P';'<P%97@Y)!<H"06':9QA+4!=%X_
P/G_K?A(V5 >20NRGL@YV;",5C8O!J+<U3FOVQ6RJ8^$P6_D')C?UE%F3Y8&H$S+I
P&'_9BL19LV&^'5E+*EJHVO\E6%\6,&KB)0_LHX\>RFNK<G%>VLQZPVE9Y <7P-P*
P[:GHVBK[V"?0XMS(1Y PXHOS@6PC;Z=XIBH5SXYT8I9$R<GE%<0;=?=1@([TRI<T
P-KS,XQ=XL@R0Z8GPCUK_6S>2;\.,B8#\=5OY] O!)<$_:N2D-:<OHU^1!HKZ+KV<
P]<TY\!K5C5L8/)JP-%Q]35U5+X;1N,P7$B#4:=[&:ZJ,&'U#KM5GC.^M#B, IU)X
PI5TK[T!2_^-=OD,K2I-1/@L\H5SJ2S)O;ZZ8A@7X?'HX&\4 %XUTRDP.#>UJ:S9(
PH[H78_@>11Z_<1D@EJ6AIW>/)=7QZ(5.GB;8>11L! /03^D! <^2,62[!$@O:B#Z
P>,B/-RB)FPC:T=F<PL@(:0O966<=')JL'WDW19G<R+7XV:R$=]3TOS'MM+6>SM/_
P3N4LL_K7ZAE(FO)MH[Y#MW]=4-?_ELS;T@%\6<PODP:FR/H5(PA:ACY^-OO/E+! 
PA:D#GE9*8V.]J\I69WB&.W _TO&GLT:?GU.[]>A1J<$BP"^Q$0S7J:#T,:(S.H!P
P< WC+='6US>N-Q2?N/(56ABRC[#1"CB)2)])P58C(M!J.4P#$L8KYWGZ=":*@C,B
PH_H".>NT[)Z :FR,;B ADOLR(L;HL*X?*:]VU:72 WD6+<]D<!A5-*J64(A#=Y(<
PD[I=BHQC1RNZP<@:;S4#[58^^N8"07R7'HV4U8))I!3\VZ ^-T93Y/+=(Q,K4@Z=
P$  [4'@WGJWEF"FPWZMXVSHZ2@%L0(@W&2)Y9A==,RC@=;CL_AXHN\)YQU*_=9>K
PBBI+,U)B6CHLGEG@^SW[;B\>1$M6T[=5#-$T8$-;\<AM3E'OF)^1+V<JP,*C_YQD
PMTDQ1M]VZ4@$B ONWX$,KJV(<?X.XY0)'#P;*Y9<GICW6D!KO6,#]EDNXOJ $VYQ
PN(28./$5</I[<8>D?I^B;9D$\W/94HD%@FQ+W)^]G\QD()<@.4"%K>BB\N:PQ[6<
PFO<R=>1>3R&'P=B+\MK2P2#65 PJP6992%@]X!95L6.)I*%ZV+K+'\P*9N'Y.8C>
PR?<<M7_*QHXEW]:2_#%'__H36H6S8JX=.?F3 AY5*G.2Y1@XO3=-X&NVXO".6L;R
P&CIZ',9X 3+<1E\!HQ:VH&NZ_K&8]_>^<!]Z#^=BZBX>Z71?6:O.]2_/P;9H!FP)
PMAQ6+R\FN.QN??-I%AIVJI8+ *N3](YG?-04K^8,Z&-'@Y?"+/6HD^X5#5'&/_UA
P43F-+IKY0A89LJI2$ G/VD '=9IX*[)$BSJ#D'@+H@64XYKD@J*K52[,@9?O7"9(
PG]"^*8)<;B+^Y;E5SU*M9QG!Y?,H'ZR4S8Z";@^"4OW^FY[M//?S+%$$U/J"XH/.
P^+JFY?^[[>ZNNM0/'$_TM+1&6U+K] ;B[>EAMSV*$&E@H1TB5!Y YZB.?4*YDTNE
PY?-O$GA^@Y*G;*)32-_L-KI4\B>.*=$XU*9Z*A7L3%N(;WU^X(;/:H,^RA[6O&TR
P;6_Z[YTOJ%W7%D'HR586W6<L#OYVC,9[X=;<W&:GGFCW$2J[M 2_'&G,L+THQ%;^
P,(+<OU/B?%7"C]09%JF'IM65X[%R4F=J;HGI3Z D-%)%M7P<H_-FX/[N-0HS/?CW
PH'Q%@O;D7ATD9D(<C>+OYX9B(TU+02*@PIZ5,[ QM1J2UOE315P^KR CZ!->Z6H 
PKLP?;TI($#KS$\MR)\>J6=Z!M"VWW]<3NR)1165I"9XZ9N"7<BYO,O6HE6.2J7>D
P?ZF-3GV"LOA:4TNK\!L&!R]*015H>X5?*_O66@;J,7E[$!4+;@P$F\/+RG]1 A[B
P,<SX,F>Y&*-''4\M#T(_E;]M%IK.^J%6:BHV]K"LA]=#8V+D>KZJKL[GXV(D 83V
P=M "\3YBJK#6F%Z5ZZBZ9?/M%6>[1!5.@?ADG6%^7.7&)VU6RITV&T\55E_>9\!N
P6][W/T@G(CZP-(Q,*UERRY4IWR\HN,N_8[2+$-4:='$0===]Q[M75F^-0P$:C;)L
P))&OORFN%8^].&JA/7BI&@F&(N>X><0MAYI0F]RHN5'=I:<2(.]VY@6;!M3AJTI3
P\\C-[R%B#-[>OF;I6)!YKN>+]8=V!$ZRFOP[.".5[L\^!0I\-]@UFOG+T0E!J-?.
PYK-[$P(,*@[C9 ,*UM&"EB9-ON.8SD9'&:=Q[T#N!P]$!O_K)6^C]0DGQ)NTR-HN
PW L=R&O(<P'#]K<Q2T@;]:+"DJ@5[QR&)MG/3"L5ZM9GY&';/8WS<PC>1>:\!XNX
PA;C$22T!(K>R*DMJ!.N)448Q*F)62SGRMM'E]_L/3\)[)]]&R=;Z=M2O]^O'1G<7
P/3?G+0?9W^";9<A+;JJ()L7=@2WJH"O.W6,)QM8>\H"O%H%2@@0]FV!U\;?TQ"&J
P_ZICV+/FP;C].378BCLP4"W_]";NPO!>C><.0NROI^>W(6(G%C37EZ)0>* 7M(!-
P?[L:+-U6#M8=9QUX%!*BP)E2AN;)ERC%@=(G=2N4>?]GGK/FKE-O<-3\+MT'>8C,
P08$MF(K+9-08/, 'G,G%&SUR(OG-D'%O!TF@#J-R3DX7REC.>J:_V&[-:H)Y\($Z
P>%")?1STE;!I9PDX23]4W"GE/W3&PK3T-0NWYF.VX2,MLJ>VM[T.-RMH9%I+ +'L
PT$'[E:<Z?:'V\OWDVHZZTR/(13UUFL/MNU9.ULCC$I>J0=YCC^6Z=>Z$A;/<OR?M
PZ A^G(\UZ%VK)MKZ ]%@_H8#OKVS:#H.GVWCJ4AL]8D=*7@.S?&WI(6/ '8!51/_
PM[P)W(SMBQ7]8>8WR@N\HRC#U.4>E52LX7-I4"33@XD\66H7=OL?B?QC0>?PA6R^
P0 X#R%E(X7:RKC$!)/@QOT+GH\R7F:5&^2!U+D?G0,[_0FZQ[Z")13^(!;99H,\E
P&-QSZ^%.J?3<IUJ6A>76"@.V(LVP.@JH1OPO89)=* 15XIOVC?_E4( 2 ?*>-GT?
P:W6GPLT1F<U7S)S6;HAD@]\T9S)R>GW."GY+>5Y"D'F3J@^&.1B8!K$5DM,?=8X7
PN@(.F[%(&^+5:H1%1(WU$Z=C6CH@F2Z%@K7''T#;LP6+D9/E.KSA2-X4H>J-:O5E
P>&/U!?J5^,@D)4%O>H0Y'9;W$\%W[*=T@K1I&HN7^$<%Y G^-X@<EN4L)G'A9<7I
P:CZ9WLE+?[I%4O-E 3(#57CD?LEE@!R2+LZR6!Q$D4#1K@1M7JIJ H^V4P (\%AZ
PXCC1,DHV+5<ZG(@VR1*C&Q")IGQ=MM8FX89,99E3-?]6ZOJ?Y5P^]TBS6!D(3K6I
PIQ$D#4J&]Q);H;. -- )+!N&NVZHOKJFN4#B#9E*4D8F?SW4K?#R*5:IETK>8J:H
P$]/8/+SKL<$5?\=Q@) ^^[L/Y1MR/23$S+O[Y0+CHT.Q!=NM.7E/.T[OW\M'-#\7
P:LB"WTU<S332*8-:;G\Q2) ^I#\\GF@<SV"5.QBQX8@TG&DQ(<GT.]>NJ<;R<%[*
PGY5^IR7DU,,?,<'(I G4;'>3<IGNZ\_G:/_;W7%P(R>?<J+UF4.F;5A*&L*]J::!
P"+_S2364>S'CP0&.JB%:_U(K40^RZPTYGK/DS7.MB=]W?$%\G9D.8I9#KKO Z'++
P2KQ8R!"E9$@9.2%A?B141JHQ3WAQ\Q+WVQ7SF6M]*9HKM-E8_#2J%W;LH^08+JE>
P:%K&&],GIX[6-MR9()=E<4-RKM#]WL:7U\ONOE-X&5TU]S6*]A&.&;WM-8OCZ^Q4
P9=J%93D1>!OC($+-(+9N ?QUH9Y<4VQ)%6C F<0M_0A@/JMS@Q=QW\/9MQ(Q+I;Q
P5,;H F3;P].,!L*+M=P#!J3H@@%WLWZD.!G5GP10.4HN'^@2<<LDO;U'LL#+RD]]
PR",'.TFK-WK"'["(_V"REHT$A4_AF+:7]IZZ*8FM57"8V&Q5@&FM?LXU#H,:,K@^
P"D8D! _8:Q.? K*@? O*^WM0.\8J3$G$^^.6%X1'6""\ZM%2_KC,/;I/\SMD^I*4
PX[-J>* V_0!<EU>_3:ZE[1D%*[D7&=]'NH]PQYQ0SXWON&/.M*3R,<O&]XG/"@<2
PZ:<X3O55EG?R5AO2; &C, ;?:QW:"P%+@%_.J)>E4=M-!4GC?EXT,*W\OC&,-M#S
PX W7O)J>J[3)0];PQ?,(MCFV*A[)?2CUD;XS[^K?N=@ %.4 +!_7\OQJI_7IFT>"
PR:%N9/D2Y7WDWG-$8QCL ,#C>@:0]$CNPZZ\RKF:> Q2!W2=*,\*]GH7$!$IDP^B
P+GM@F;1A/+]UI(]>WJR4@3US]LJ9<:UK-FC(!>UF G_#'4V%LLGQ C:>:1&?03>8
PHH4 ?+\^^@CSYL 6)('.,7T*[E:M]X+G7:FS!!N,YB3TK$:1R% [5MR4%J9]=722
PC,/T$QPXPKE6ZV4H*O_K6YDB/\/&1._Z7LK%/"32.<I&[1XO-OJ8F"K:8CHR<B ;
PH-15,FF/61TJSM5CK=GT/V3=)#@!C;&>NL!_+^;3\+J%4R2:T0U4L6ZS6V\!*\GJ
PFD.OD"LK5(<P,06/WK>&B=/5 0^PC6_F%'8\$I55$D?5 Q3^/;[8D:/K@^.UZUE4
P^G!4-O6HE0C@-EK<G?8$)LF291Q FCD?[53!P=PE=T]R?0[.(PH$1?I5\K1L=M:[
P\7H5^(#-\4<_FDOP@>0P8)P[XJXVAR6YL&4BJ.>/U,EH&TZ#NC3=VKFT8K$_F_T6
P6 K >*9&FE3QI<( 89@8$,T0/76GEO2O#N3OF4+/8:DLTA2 YA.1-O,&*7V7R'8^
P$_X8U'012H0^,[K]9IZ'.6_"6$J)3?52.'H2=)U-:J]Y&04:A'@3O8NZC=U>SU(_
PU\S38ZYC!.I*YJUX%?\))%G?LCWF^^\Q.O=$;O#WO[6/?VY\6QWK1 \PPUUQOP&^
P#O7LWFO_WW_C)(A6EYWW_<;-8!X8^6PY$R)LBF'-(I7<H/):(\CJK^@%*E#A#A%/
P2>B/%].!6._=89J8_A%:0F=?$ !.U(M/2 Z(D@5)7_O3:R="@:I<5W]1Y;67<>7W
P/=>(5*^=;,M+<<6_>ND%\F@L5M<21]:A&S^5,0M6)/L6&!Z%6'ZBBXOOZOGRSTG^
P6E@YRK'KEW.[&49OWH/\6B\35Q$76$^43=Q5;;-&>FVDW)/I90PI%1;XEB.%YFCJ
PU%VW-U? 1$N110PM#8S%A."R6,F_XM"43BK)FX%W[KA!-SNAKD,=_3*%FB$>F2M3
P^+>6"4+D:WZ T)HQ9KWDYZQ/$#N#TMISVCO2[\&+]S';NYE7=)B&JHXW;E;T,6&=
P0]"OHCN\&$G%I7IAZ$B!1<A*^R.[/E3RL<&*1V1[[1 A-27G&/*H*['7H.WOBYOA
P-GD-_B!ZAQ&;^U2U3 :$^JN19,(:FK9^]=IW]XHXV\R4E <JI=A4B[-Q0E]9V+#L
P?-UBRW8OTQY<_2V2>^&SN!$4<[TSR3AG"_!, -&$@WH/.76^9CNTVOIBJEY(>EZA
PQ]=ZL'S@62*9K#V"3[?4MK@\ ]A8T(MW#^P32*N@]SZ6$&^6\TAK!"9WFYHS,P6H
P1ZM/#/LZLD1P>XKD7,P#&]R6 ,Q?&NP\ 5I)G4405U3XZY R0Z;OLYF7,& [;;>J
P V59G(2I)G JZ87-"_*RGVH^M[V!I9KLSQ8:L=>56FT$F8^-V<R>JB0=I.J+]+ @
PE^\&',A<,N:/6@9.UA8MM0@H\4NC\K7&/GD-%8'DP0G#S6/NZ^*EB')N6?D6T.N]
P^E&'D\UBYT18UM4813+_88_3I4C<10<GF^%AK=-%F.]>.U&3]"-+EE?:@P@F5\*H
P#;VG7K987:V 858=7$2<[0<9H?ZF1.N_N6C]C51EI<QJ:8^]65W.X:WJ!,%*)8A5
PF2F3AH@YX7YD]I3E;.#2S)*U1UB1FWLCI*M/BEP"N*?Y"-+48.$64:KL)/_Y4I$,
PQZI,B@BB+?YJ9M;FD6ZEH$,X(#)6Y)(3:S=*\0-ZPK\F\9<IC:_4N+'=5#CEL$OS
PCP#GP].NN-V4'O3#"<*7""F*OC;V[T.^AKOEIEQUYH?M?+*[1)*CN!IX<5/ITRW;
PFP*[^<)9O:)=FYF7;@6XL(8@\3.8D4*L.-&X\A'RN^O88RT/,>I,=DN19FSIP@&<
P^XPY:>A-M>C 6'.[]L-+_<%0XN!=T:$SHFB>D"<Q.41''S4!YX]/?7_,08!$XG6@
PZULL@Q"<,7Q5H-5X/XGXG@X<*1_DCR4Z$H-E(\,)SJ@]'W(VO+4*UAX5VZ.3*>CJ
P>![C+0 72HUUZ=\=$XL)[F02:U5 RO329+FEPE7.CE>J3B Q$"M^$C5F-R59B"4K
PT<DNX)E!=WDQH'V)-JH1)]@K9TTI,LLBY-PW=OCV1*@1*N[(L/H$1JV_BJ)1TEIU
P&+W/+]HQO",?R@%E\S[0%)* 51USK*Q8M:Q^ *],;1ZGHF+=V$[KVPE\23$'O0PN
PC4R(4X:_H59<^V'I> SE0Y(=PDP6HG!M4""]3AF35!V2.;I/LZVYAFR^(DB^<KKW
P(BK?SQK$:>(3+T# />XKL'9[]0R:^(WD^A3#8<#?:SE/'WG&8V: H"WUS?B"4-^-
P_I?D4F14=>);\@^Y^MM\_I1>JTA2MG]Z(&"#($49<@T'0,/PW#X; PPO-%6"0T: 
P3#"0+(($!XG0+H(QD%S?_?TZU3VQ<7OOBZ*L:*'DC!_]+D-&6^SQMS['&#>P- :U
PO[R%6D3;\OKC.Z+3,SH:=D?*2U7?IRDY(D[D,$T<9U8C!KPFPX1_%7Q]NXSXM; %
P?4T/V67(NLQAJUV4D_2W&CV7@.UIQ+&L&*M;;EV%*2>[_>(I>@IZT9M/'8@'WGT^
P 23:'6<ISD47(6/4E:U?"/&R%M"HGA<+'15QN"M(55=E\33Z*2Y+28MQDS6Q*C+M
PNR0@M6H%ESJ0HEDNIQ=4!K*[/9W*\'"7@ 9N_HU$FF0M;] SAM7Q/#S,CQ;#'K(9
PE.-C"SAQ5F6M% ,8T_C$>,;)1?=#A<</,*L3:T60%H_]EDOE=\S0(0-#0THS_1J.
P]$_,LOSDIN]?KX"\RDF^*D8/'\)=3DS:=Q@;G?3'6.G."PI!Q75M\HBD6W(MC8+B
P=@@YVORBE3,/,?:Z3GJ3@9N@6DEOH^).MA]1M@7@^"'<'[$O3@][!6C\O]$$I1G 
PH*C"OY78F)<_+J^YW5+-"8AY1B]0SS[ K2/A[608L93;J44Z8/3KR3IS<^)O,B"[
PY68=LFUGJK>\N1]?/ 4SK.Y!UX%5KC_?L-TF[T-N=EL,AZ"Q4Q^\Q55A  \K>[*Z
P.6F*PZ"QK&(E95C>D7R>49&%2?\8W3WW,ANI55NZP_;K./50OT3\5$%=*UL)A16"
PP66^?3Y>/2;"<A)Z@!]W:FT":\6 J0CDBV\(YYEQ&F!Q(D&'!4VU F=;E0()=6QW
P_T5A,KBR;F5>.H7=.^SH^;7GI!(=Q1OU&(IIF$BU=4<S""W\#GV0OS:3-$A:&BJP
PB/,\((V7CP$W"T)TC;?.$D1A-))*"4XP*?;EZ)*F)?P/%3A#Q= =)\9N.,YB_I=.
P54$]V]+)-YQBH)2@4_)8;6H;XKS.0-;$$J3EQ9)&^ X[ SS\ <CI)%R\3'T2SM1D
PA%#M- UP=3Y8A(Q:X.SH@R9=",EU"Z#! F ULR^R:$+6_;28CC/PICE^]NP3AV;R
P.KYQ/JEQO4'R@I)@QET(1#-I@MOPA(%90T+P-T" Q_ESN9W$,V@9F$XEM183H89D
PZH.@#_[60.A^@-=11.UKYU%08=*Y,UER*)?\:X[9#P!5,1L,DW"K[\$?Y(.'S(A 
PYXU2;1RQ1(=SZ2P)KX.N\[J!NPA\NA"HW*3>/750W;EIQX/W.AGP#*BQ!(;HR04,
PHOYV=6Y9_B!:TN,>[K)3% <^$$/U_3W2X1.T1_<2SP^99<!LE=^O7))^]K0/I@[G
P@>%>/#SQ_%0Y2DA<F&AP=VGT^[M1( :'C&PC W3+:@V? 6[WX1?),CWSD=TISR@-
PG'?[3Z<7F \8,T[+ YP_0_36 /[CU'TW)JBZ'"+R+MYP4M4K0#[P(9L[W*3W'6C8
PP4 ZOG]US$'(*WAK03^&O8*F42!)/='<^[C9 TJSR&Y8>#)/U<MA,T.PJFKO[Z*Q
P:MA28Z< "%9]M6B3090$1&;SGF'U='R%#09DF=\E7.J$/LC!,.%Q'ZQ;M_T'L%^#
P;2%@:6^"#07X?^M]&EU&6)<_!LPZP3\2+HS@J9:^OB/>N@RMDPD-SZB5<%VXDC6'
P>I=076],5QJVJ\;]&I!C)LQP>#M@Z\^%CJL/8!?6B@^ )'<4%0FD0Y-43&A,6<D]
PM%Y4!Y5(0,D[:0C$?X\>7/7OFLRT/^@KF1<&,U>^9:+,."YY_!+-WC)3<FH"/&Y3
PU!IQUFJM)ZSOZ%*2%1UR*T'=1:_.JPY_G7JH?N,BH?H'*E+!65HR96.HR!1[U2-3
PZ+="RYKY%&- 4"I%:G>?!!Z\"DOS2YPOA&R)PH4O+M0[!V?@WP@[Z9S5-6C=KH\M
P$X!>Q;.<K*W?JF5V \\1=<O%C'/"0Q>?H>JE0HT\EXP%X!/C:%?9B1NIGU><R&:<
PT#3JV(FEDNJ^_"<DIJ+'_)[]FN!->?;L1[M]K30)$B@XM.X<=5=L#L+N&"Z8$JGT
P;TQ[+MY'Z9,(LAJ^; ]JZ8,>[8L>BJV_3=2;#M0YB,O7ZCG\O8=@:\ZT1BAA@(LX
PB"W0D\]><%QH@B UD.*+QF!=%H+T^@G/\\FMXCDX>DO=P M;;H?^!U>HU#F:.';I
P(@;<YJ< Q=YQ[O+Y*$!EAB\Y+.MC"3$O$>;=Z>@@,B438KW1(^$5.?."]@0$5Q$N
P05@?@6@^:8[C>BJ17>UP#8-:0=GIRDI(R) @$%_S%2_ 3C5<Y#E@[X$[AEG27K!0
PT;X"V*N&&DB#P,S,B;[!#/WS\>7?WS;4"1D\>2KW/YL:)F+I%PE[!"1]: -:P ],
PI&+U9(Q[BLX?>5[SZM,Z6AQ"'.";Q=/6T&H'QJ_3I@R]X3%_M-BSM'Q"5H;4BLMF
PD7D"6%W \[^+LL%DR92]G^6(N<]8<)PU(U#8'NV6+I=??*0NXS!-].L'#^/C%IMY
P>)D.O<;R>?K,_]JC]$LBT1'G*WQSUN=EIN<K/+4L&DVJU7-[!]/[WRIX=U+E$XIG
PI:[X1^AM-HNCS=OG30Q63R4N+U_# EMAW?B0UOV.B%&TC.WC_U$N"S$-=5';*TI4
PO^TB]'-FN,<5]@3F]AW#('C?_S8,'^];WLH:J9A1>%>L*VL4]1-%1ZK.[4C'>':)
PP8$G62[7CB)\QW=247;?D*<SMM\\AY!R&P.Y;$K3,1DNJH@\9&.H6.I!><'V:(M)
P6$1KUS1IX!';QJ&/2SC)N$&D%R/V%&?\2KO(%9QPK3J.OI/Z?(SY;";N:G,NU2#H
P\"BHAZRWWV=MKKFJKV]-./M?7J? "*8AI8^NQUB671["?3%7A/=UMHB#[R@FJ6\U
P0(@%?Q=[@%_;8^&NSN!8F?I5^4[NEUJ6].!5MYV8,L4Z[*TEDE]X"A?Z]IUPB.+_
PDSW]T?507)01Z#W59_-BDCLO8!/+$<'^H,93]_YA(#[Q'\9^9I<JAU2"_,4R9P1X
PRHNN!%C;J9#X0AI  L6K[._=_;P8:[O#H]TDRNT#ZS%]%6-QD@9CQ.J3M%OC >\A
P X2]53AYKG2#"F+$:ZZQ9+_7$LEG>4F=X+,M6&Q>U*O! D. 3]B,*0)<I.51ZR+O
P1,,K=#;I<^>56FWR/Z08=_7H6SB->.<N+*SDVT8+-&O1X'Q*2:Y) 93V[=JC]G_>
P@!C38U/IB4#GTFIG7;F"OS13+I,/".(NZ/B*5($J1<Z=@E30ZNXMB)M!N<0<>(QF
P7>K0Q+0SMJ 6!LA876U<0.EKMLK%R?KKA87&MFA/5<81?[B'NB+A^9+5VB+GQ70@
PWVY_4;PVX5%+I]S<35<^ZRL3,#_J07>M:-8DYHVTL39<3CJT&_^WP^,*/%"_V;7H
PXN4HS-E97QU1\6.V19S+P#)ZUWP0HA_*%T7KXZNR'>7;%Z+$?K&OZ4S=OV7-QYD"
PQV#2FU^\T>37@UOBO$Y.-7GKYJOFR70T@<H$0:@24L3!0_57Y[KZ#\.I=*&79CK(
P2,LY%SB1:AQHL%@TJ0_,=9TSG3<D*4+PG\7P/W3(@.L.<QZXR[4Q_D0H:WIOG@"D
P+ZZO<DBXICY FQ8%J^^6GVM^ 4PES+$ 0E>L5H\O'ES6(( K702T 6W<,@Y!JG;)
P[=IO-$;"WOS'U@IV+FT;),Q=,G-HB_)C.[]R"$9GE5Z='NHEM)C),<<-IRZ[&(EO
P@:PH_7U(+9$4**+=$OS?Z$7_. &%37]*ZCP^1F*TSPI+;J.R3%1?6QB%8\%U$J"9
P09MFR)[8_SG4EPU!-,VOELJ_*@'O>;['ZE>-FQ8!S3Z@;!JC7%]TG$2_93 3/YUN
P,#L8G-6BK\DU__ ,-NG;]L9:>K*9BG/:@:1H"*&_6<#_'S^\!CEB8,"Z"T[C2Q;P
PR[&&P'Y#62T'_[BGZA)$QS(PBAX:>/+!MJ =3JW7EW:7"+@MO*$Z/<: )<&1Q7SJ
P\G'=[,\I+6YDQVFF(*DST;(5;A(^7X%VE%#2"P?[V*GROS,[1A_IP$D/ V_\#1$#
PUM/AOU\N3ZS)77 DX^X=O?^1,)(7"_HOXZ6]"_<P)"_,\=P^L-\6 O0H!#<+::H^
PU _+#T@<X3=%\>5 P!??C+M/E=GFGM(NA6^2O&:YRN*$:^$;\?WR5R8>.-WVC5!?
PJI;%H/!WX_^->[Z2SLSUQ\=P1'] W6A@!U-J&G!G'V5,)\:;(9(K>":*&(/S'9B6
P@'H .-_:&$..MXY7T2CZPK5$ZTDZ,+C#2M5!O4$FJ-N^LF,@3=TQ$21"3C1:7R'(
PC4TQ_(M4&*H9!<7]F)LB@3S\,"Q^SYVP_FEVUBNLNX) .Y\;_)!CRO%)\]^3C@"W
P,C6W;8OUY0KG4G:5<8\^:F,)ONRSIMSP?#*]UV6SF09QI539@.-(5IE/2WRQ?0&,
PV@S/@?LNK/Y)KJ)=K[G'I1\HM^F(39$C$^-<M@]]38^J?=F7&'!!%+\RT<=%F6A5
P:\*HMO1**+^VL-^W,,' K)XKE3_>$:'NC_D:P+OCB97;DH=!Y6RL9$0BR+\-;$6?
PT"5O3LQAP<#51,+<?2JT<":Z<<%ATSCGAE(<$LW.$(T]LD<X2-8LS4E!0MVITEO>
P9."]_H5K!9)62/=IREY"#U>=DYS. HZS7D0"7KV?I#0TM::L3B6E?Z47L.?=NQQ/
PK>]7T[L00O0<A]6SL'PDB-0:3D?K<?1]#D/@R\^?:0OHI HI8ICFV?C<Y]PT.I"&
PM6:-8H0LD_#P%_$10/A5/&^MRE<,7LVLEW]B1[,_)JKGPO52[A&@&H"2J2 +)'7<
PALPUU%N3-@.J:DBP+,%G,:OA3Z'+S)16L.!EYS*__[*'YFO]'ZQJ:B9K[?5+<&5Z
P<9\3X%[VKT3B'%.%^?Y?;8V'<-;_4GYWEB^@782AD!Y+U5P.6CJ$5/=*])"X"!B*
P%1+(@672C'%E+<KZ+D#2S?A';"1/>HVBV3HM\6T=2FFBIR(),-B-_X#IJ^BJRZ/S
P/D9N^I3B7C]/U9#,\U43\SJN4=LF2$83 D6;JJY=,B-G)]X4I1+ P$?I@U&>[@L*
P-"$!Y(+D_HAAEXEV>'$%1M.\QG:G]93NBYKQP^),2M'6CN#9ZI+]DDKE,[(TYYPQ
PNB6=S(C=1QRE9B]T/=>0/UJ''Q'<IPI*BM*VAQX2YR&+30O ,\Q[$8NA@L8<!LU(
PY&KR&HS75FFB1)(K\YS)"K'\WT/Q4#>D/*X6%9B<K^?U/]5*1]M'153'T_R%)^/<
P\BP1)XN:BDTHNQEUK= K'+<VS3&L9H%SFXW,;$W\1FNO**:9#OVH%-*EIM.0A+.N
P?%T'-%&3&R0B,?D)R7T]N,@HT?UK$^O>ZB9P&^CBPC2I2H_ Y8_R?O)7SMYSNN'E
PS?.2YXSZ4:A/')G)1:M.>B:8*@):NL_T@WEO!8XV%EZ/'O4FP3?O+$2+F?H 061X
P9B$<9[K<5F@QQ*N1Y(;U)9NB:XDS8W1?I,$!,'OD(L/;=/X<4<@&__>44!6;V:Z-
P?:ZN$VN7O^G*0E.IY8Q]H;=P9WQ3L0#S1>5\\R"3L->(*R\(N<7VCE2*?(]HK\>E
P]!-D*:-W<72=/\*'6VQKB.]]G](F7Q,0B" *<3+S04\W)L.=E),SR, 5R*7:?@@*
PO&_3[/&,[S^LG0@?\2#0]W^>N,2LGE_V/G%>E_AF=A^\X04)<3EG9C;K3T;ZSXHP
P&;^CPU)#?@Q4B.QNVP\228DR$P"CG!P\K;N8T=71;#&$C,A3?NW^PK.2"S&!'6I4
PZ= X%9D'*0+/[])M2!BW3!_IUO-EAQK"=IJ8.B&;L:N!VDZ;]L#-ADPO5-03,A@R
PS7P0W\:DTEMN2)CMY^N0@*?G:#8JXFJJ00?/V1#AKD&GWN$7Y&EG)C,JI8SX<-7&
P)\*;L*6D'7M&IDL"B^"ME7,O_&^95Q,3/];D]]U_L?18=<")RT]_T0_Q@%%XB^!/
PD<^S)2O?J"AN:PGK@,4GVR<WC0B%H78RZ*#SP$%'%T<O[V\]K3^9A6=8\B7#UC-/
P$1%XZ-A#,IDX@95404]*7D=S^7$LI&>6 R_"Q,.*NHB@5N.SDSF:U==Q?\/]<+3/
PWGQTX.L^2TA7_)%]XQ3['39Y/G<N36* /:AE'BU<G@2OV*R HB>*!GI(J5<W:P7.
P(1&G"G7&">+KR4ST,MFE&DE0A@]U(;7PMP? 2*05Y![CJ]>1(<X!*LZI/FW_/!7V
P?7?%P))_+G"88?5S?K"T2@;S0)G7+5J(X':'8D5*)J[>OQ2X918B-]^F3.6]54C 
PA;JM_>B?I_#''(K5,R 4,'%_04!41ONT&UL]>+3%_8-D]6BXI*TRO*ARM_";?29L
PX1/E?_UQ#.QDYH*BH^C.\EC7JG?\J75_=8E'BAK7L\P3PS1AWZ4<HQD#^RO9FHM3
P%+%L&D0E>M8U9+[:6@#FGY$!:/LU[=LA(_W_XH<YQ8#XC1;$*+DR]P'[0^54O>J)
P=4!,P&1GN?I3 O+>57R\'V>V*.1M=*OQ42.N#_X4.Y0DG)8/DO1"V<!PQ[_"J,]T
P=T%;+RHPQK+V'7Y"NBBF^\Z'GWT(\ZR5#0?R2K;21F]#1X3.JW+8ZY10][?D-O(C
PY< YD81A4,_RJ@>!&$F? :5H25^=2T_0]'QI\J^TP2D@7II8%_U+*CGZ]33ORH3#
P1?E9_L52\ULX.$H'/^+"OV4,:#/ M(UU=FSH\#I,)Y<;I:(_]#T$XY9)-/#R;(A&
PLOW!E5.7*U;,C^Y[6=,'TE+9PUY>6; ZK4,QL+CQUIJH Y.+:4M?  QH#K%CNO$E
PSZ-;YFY:K[8^1!50TX9K='JN"""DV2W5U\%4>/4N&GX9R&N:0)AS7.]^:7/='-V?
PHHM@&BT6.DUT M@2V34B<VUE)=]D/?X]SI\GW&#FWK)#H[ID*Y0YV,@-W5M,!X&?
P< ;*N6$_!*=6AX^^QT-'E-[^=4;2(1:"!0+NJAG@.2)]\H&S[S=BJ^5,$[OWMAGQ
P,=>L63EO3HA'X,6ZWGX]L*2K]LWLW1XX10+@JG4YA0"[LR)Q27 Y9;8"_]7WQ@UQ
PVBPJ\A7]59W.,!&8:]*1NAL.X=N$R J3B@1.V!1G(U@3CT^I/WW19$&@3!C NH'H
P$2RI>JMJK=@*?9)1!!][Q-7B- 'AIA:)I^J!)51(_?KN,O^V^8\XU8+CZ;ZU 3XE
P*H$3X-\].BF4!8X?/X33C+B,M('32G*;OULK?.)\4&0HVR7:MWIX#8Y;8S].:55"
PU E<G=$??@*9R\C,04-332](-^)29W</1P%),;PMO27Z$<U7IPO?I\RA1X&M":1O
PW?0H,$Y6;P8X"1]"*XUF-867)K27MU@WW[R@V<>?1'9YR8>[C\#RK6V#EBK]?$M/
P$+>5(!Y435)GPO,(6#O(MTM:I)1"?-5_'>"0Q"O"R,C>1+3,@4@M<SP-.6JO0N:G
P7D:R-A3/)DK!EX<(3ZQ/>B>23#I18J2*T)Q]H5:&ASQ/A16VZ"$=O9MWN/</#WT[
PH)?XF@-N":7 _MD)GF[>%303^GJ^S7S*X1J^&+KYXMHHZ\7C]1XL;]3E@.?J9@<4
P?M#XL5/:"BUN+3W<+A$%DA,N4C+0!1#09TAMEN;68'2]KDQJ!].H#$$K<21ED'17
P1NK-8/^;%JD*'CV8+K^OG#4"RLT5I%7RV+G,ZS+2P]<L"T%4;#EKC)[N^O9O^A'=
P$IQ[2H1NYK1Q<>WJ_QZ)8&'4[&#?AEW="1!QW;;.R?WT/BLRQUL(M1STVD;)-0OI
P\"X1H<1W(5S?_ %/6*#N14FQH+O*<&.L20]Y)G1)XD\]UNQLMJ^O^1V);:0)%3[6
P!!?-? (:P7;Z"P0DFV.E:KJGLM(K2^X'N6!&3\JX,C!1U(LQ3V8O4G55&B5AU7T-
P:E5)4[QK_)KCF&\Z0T/%:>K40AH=A2  X\FCT[:/0ZVXTF_>TG39UY@#ED(=\/=T
PR''0MY?(#C>FDMY@BT1./9A,:IK  #6$'CD/4F7V5$D#H.O8(*PG<XUS7CEP1*\3
P\91@3-(7P=V5ZY8G%5G#-F=ID@>,6CBS:J(/!/-UB6A%_2(Y-6;+NI.Q&@^YX3GL
P<^^@#-BGD>/Y+ Z JLH:X?,JQ<B!5?F32,#C%DSX$R\2(MU:_K:[PH1J@A]#QW@$
P)ODJ;L&UMO9)^/^*"MR$*KP*J['W#@ _0;J<;^I&?)-^7Y7L[MYWA, 7/S:(H7&R
P9T-VDJ*^:J6!+"KA V!32IG;4,DL[BIWHG"LP_FZ_Z&!Z0VDW!=SY4D(0G!PE#=8
P02#[3MR;D;5["")5:[A 8D0DL)GT_R1=J!_#R<6R"*IG_)IKUXII7*N74#E-*O.#
PP!H2BF2S HT.^+/#LU1M*4-3$5J$),W<_"B>Y-!'4B3S1_] H=%J"^1\T@+/[@3X
P0ON%Q)8K6($;G R/DLP-DD,1DA33&5N(R"[MK(B5C7DM,0Y,SLR7HX\@@CCJT'JO
P]6V]-Q(UOZ,@459"*)M9R"BOTN?[2R#2A[MA(35*]@+3"_<2=;A-BX0>;GAM(Y'L
PPFL*Y*18>0 O"/C)+OM88P$7$HW6\Q,)\'0ETB*WSMH+;X# S.[R+=+F@=7SWO( 
PO!ZQ;5 90H8EZUS8NP7;(]AD1A\4RFMDMLRF_180RD:SELD>)PI/E.%,3=X8O[4)
P8J:ZIL?^U@XZ&9C*IO@D7C2>GQ>;BZQI;[1(V%SS FBS,%-9T!V.R9U"[-L3'\<6
PJ0)P.$RM>+TJE@"$E>I)4+K<(W4&SI)^FK:]<(%76=RM?GL7$6H@)MQ DI8Q@I7R
P,".UCT8Q-P\D"TG=Y@)Q;;S-8'X\"PO@2<)A\T]AMRHB<<%53%OAQCS6BWMVQ,J5
PRC@(ZNZWI]+':?B8F <GB+H2TVG$4YQSN0C<?N8JO_.UO/1*8>B2&G#J8&8:.N)4
PVPL\Q/>EJ+=)%C>C_1![.O%*L\<AIVS.T,>2N;!=$__XU;[Q=<]YV$KU_X'MG_(;
PC^1#0J&60+5'J=NPA]M&]P- ^;;H*4A,(+:ZU"<G-93V':^L5$SWEO"*)<6ND!!!
P'O8&1\@@ECQT20PYO:8&LN%Q'/GCBK#]<$Y"F5;,QE1A0<@]A?'CED40] U%V1T,
P8H8XPI)V7B]&>A0H7;JXA:R]IRZGWXS'6+Q=CA#;P4CW&2R26_T(5E>+T&%P*ZAW
PN84Z=9S,O;&KPLI@HU> H+@%!V+$XZR8L3GJC!EF34>*:/N]L20I'Q]43V6IE2 6
P*:?_&_\YS_+=\=^ @97(Z3G5&"37FWCTN,K!IQ4Y"C2%<PGSG&<^;X6QO/8\4RVQ
PTD?7-MI B!<1%)4)%S%-<N7J-H .GQ+X &&)"])-Q-%=$'E%<0G1WDDKYR!'2KP(
PV9@Z)DUETI!I?Y="2 N_'G7A["R0/4R_>3\=;+RO>+>3_CB-RY3;[APGH #F3-H3
P<E8;I!PU;>!E%5 O-?V'NM%!.+ZX:S(?^/:IE3-22W&4$6H=P5C$]C!/$IL!'IFD
P!H.?4L^]!M+Q!WFY.V^#M]S[;*0O& P""ZO.!09H\&YQ+:Z^.[S$^PJ[M);O[6B+
PZDENI%0Y=BLM88N"IBHS.%A4L6U2->9>4*_*I _.\ I\9'"%KO0;2'O<^EXWS'K[
P'3ESUCV#]I#*X8^A)M >T;@>3&HW7P)G76PN9L7!:NQ0N/HLS0=D6U:0]D\=?M\O
PL/4;U+'!\$XN*,9\HK0^ZO3#"B>D45(0:B.B94.=Q4.?7SH6]8JT_G6@W6'(<V22
PX=8X_PUW>>.H3&PEY\H/OBPS3@3_-:26\>+CH[ 1B318^)/@[?R,Q#<05QW+QGAX
P&3X)&9YOZ+_,LFQ#L"!TGLSAQ38CY/F(,R-P'073);V8',M,7700=?%0C<U<^WS=
P7FA0E34O.V6<EEHOZJR'3P#.M1&70@,KYF9LHD",4/?B3+L-;HF;^[?V @^*.H;_
P9A4:HDNUQ6Q6N1J(W4]BRC*XH.6F6D1='FA6WTWJ[C_Q=3JT9.PO4$U*D#8%VY3G
P(%V00_)Y,0:'L-ZA+!%&UZ8I<[+)@+:!2>[$B55-(/%L^8OFP#$!,)'C'$D(>=_3
P_8(76KA^<Z#ZGA[#."D[\^;B4BCJ_<FR2/*V'(+MM7"OXR%L?6F]G.? 3.$;DUO)
P/I3URZ?Y"%A&O=)$_?3S3F#74L,5<U<7,/L#;!_HLZ\8TSLTL2%O_Z,T0*R.UDJ6
P1H7> ;^^WL4G[>S1,$%&:#FQ9ZU)+L*KGM<VV)6XH&T /H$ 7N$&=VO:.1+]FM,R
PN!(;<#MB1CT?Z%LH(Q_JRPSOH+D00BK1B"Y;IFT;W,F [-5J$P1V9;_G!EEH^/1X
P,8*,"#([F^S_G[T#,-F4#!F+40WJ/?<I#%T?VQL"#!0)ON:''1A//EM8>:]_JS;H
PD3%>M=@HPA6:0!(]*199R&JDP#.C++Q6$IEN>:%P7,FWM)-3YD.C!XX:>R/?*=4I
P5?R\CT8JQOMH/7KSI#F#I"/KP;Z*IZ9C&/N><I.QDX^4)*F=I1FV#B_M9B"0,!7R
P>YF#TK%,VMHW<XMYZ"+-'&42C9<'LLB0.B5V'K)T%&U5,).:(C6:@?*VR_)]Q($,
P C6$Q-B@\A=S1[[%6C@ V$S@3@F=9\4XKX\6+GS^AE[?<POW]DN*?>*&O^HELZJ?
P/2/.#M2\W1H2,(#U&<O,ER>X'"04K8=V=>TM^SOFQA"3'5WW UWNA<_<=JYP4$L;
P8S*!B[HM1BK]P#$1G#O7HJ(/%9A&%L=F6Z>4^F=-8T.3> DPD"<Q*!^MF"A@+<HM
P.@!GC9V#?]2 _)G8IS@/88\N9T?:K<N$?5MLKQD3D?,0W3VDQH=H,4J4T!B 8("1
PA-*SR9Z;O4==VX!N#;&KO[5D!-BL&4,6#'5S&NST?2 '?&B+I<$C@W*ABA^IYUR>
P1@Z!=Y6+--V>LW+_7OR/JP$DE,G:<\,=Y9/EY*I89;=;(^5T!5_SBA2=>/WQ*]1U
P"][B23;N-)T"F/][8S6H$0;=I22L!"^.G<&BLBD9D$>WN\A<%?2J:6"9GN2ZHC%9
PM71>XQ=).&RQLU\UE+7M(KEVE)&J\,&.7*=^G_R7(55 .!SQ;_CD.L852#9&H?>4
P J8[F%GG=$L@@NV%,-K,@.?&B0SS0 ]&2!Y>ON^Y3"&;1A@L+S_?;$Y)L!CD Y0"
PL?[4^"-:Q<ER5M3UB#M@#PC!,<.*P.3Z9=I*<B=?6[L+#EM.I3=E?PFI  3F3*P@
P>.4CH58B,QB:U<T4YY UBW ,HFO0'LA W*E)TS\A?H'OAFDO%(&5P#]\U&43::L<
P3:$\N'@69/$[0RV\.LWHQ2W&HUSP]E.2R0//)51 9.5(CYC<.J$?5Q1]C@?+CB$:
PKPGD45L9!#EF[,54V*I <VN-^! <C!8_PL54#$V7H2/85,=#/!3$#0OBN:C?DCGX
P=.]DKB7)X^!L>VOU?6#\3,/=7S A.EYB%DHF2;[:L2(RH)\'9YE,E<_S:B';L\X0
P*2&^/OQ*:9?\[_7BU&S\6Y.XG?77_84=&<*:0\" GH7Q3X!5A)GQT#FTJ7LH J?D
P-+F,6_@;7 7[/RI5^ A9$*FU=?O(KJ!_Q 4!?<]B[W.)DX3'[T?-28=4XD\'LJW@
P#DGM1O0^]BH]R@VMFR;9MKH WC=%0PX$1Z6_7<Y/#R6)8%FWKPN"08V'W7%MZ1>-
P+B<(38U'H.?$>U>%+2DQL&J86#(H94""F3=)RY\8Z)#';] LB!I*AF?K@H4JD?! 
PX 55)B./K$>T;PP:RX#E0>VP1E,7GLJ(N[G-.\MT#CR7));S<K;FUF^?.W"A"$.4
P%L?:6+89J^]GMA=]TBM2>JN#9.RIWX#(><</!YL;G7Z>-'VGL4ON%2*1^4-,\([Q
P8+\E]LN\;BBPY'G)<GKP/SIW<%>?9>G?=B^=PSB)2=^Z=X=]D,L2B,YAK6Z94WXT
PZ?Z4@HC6:Z#QO@/J>DDV3:C42"EF#.R=IP1,9K?J5N 6W;PP#!3;^7)W,E<MH=H+
P,XN9H<.HIVX$N:V"(AIGGOYRRXG6[(B5UNV6H#?.<IELG2EZ'&(3%2P].$,J6'9C
P1NIB,&"4OZ'UXFXKP1R7M*038G8=NZ? K>!X:@T4F"V?CGFK,\^UV?-#-5XQ)R(%
P;(XO$NG <*\37J "IVA8X"N4.;BU-& :BEW]:I4Z_\C8NUVR?2' LG&O_[,RAJ*P
P[FK]0^S_AG0%[ZHD&]ER8YDH^D0Q:NITH38C)6 OZ_YJ[S4'7?(G72T[$UD%[M;,
P^7S(@3FBAIDYRLG(2!T/80*"]45UVL'9YJU6%1^F!,OF-N)+0 "X<U$K KN&$J1(
PU;D#8;+B]V(E8$#+B2#OJJ>$C31,DGR3M4;(L@(YB;$DIFZ^6MB,7 W_'\.. -0W
P1WG)Q,.P=Y;V(7__.,/B"_[\$_'IN%<A\9D8I&KJKDMINMO,-:@Z+5SOV:RM$_/T
P,MTXO9_G(Y?:I..^NL,4OA1-# <-KFW'T1'D<,7,\I$_:>![C4)\'U&M6O4G R[?
PGG6<S(Y]VARK!Y:$ 58S7'*%=Y;ZB9,S^UN'"B70FB(G*2%I6Z%Z.S3.#_E+HO!H
P.6;\FS3T>ZN0G@3FHR>\X!2^[_T- &=+VW\Z7F<S]VA\4*CA%#TNX_GM%61!M?-)
P;?C>0[KG94]$.)_022]=4@6"7$_LY%5V?M#@-:14060]FO5U6E60*"@#G9"$_)A:
P;@4F'\D3O]7QY5DC7N9PC=+AYHW$/F,*W2TBX4EI"!OWS[KOA5W:FY5X?>+O(9W9
P.1QB/3ZZGSHC]H0=Z1"NG#7W=+E%<*W&,Y#5PC&^)BO962EB_PJ!0<PZ#GZ(7-IA
P#RA/WAQNFO0NQG\ST,4GE01<+MD(OX?"%"N!R76J9Z1,+B09RMI&B9U8G7ASC\=!
P^Q5:$I4N-#PR0FR;F9.5OSBZN-K5MW=4;%/I#D][7F!L]";>L" E3/K)4WND_ZRT
P2VY$P8:PUJ;2<<>Q%C7WFW\@B!OW*%AMS(!4-%28E"ZE]J?VOA$6##R#SE@&4?!K
PM\OPJ9T9!$L"H6.?#G>@X@5B#AI$L>-YP)29C=QG+1 XYC\K=W&'87@S!\/2"YB.
P%WE-?R>5)1,2X3MI'IRF7 _E)><5+%F<'("*R5YC/LF^4&$^.#JX;L Y1Y#!_X6J
PZ-9\Y,X;WRL)MH=.^Y9S6WI= "(.()6N3<W4_QN;FGA"DDOO243"*IRT9\>!E@R'
PC["7LR'#DM0'[9 ,8R2*-&G7687RO70E5D)^H OCRUZQ\'ZC(=9@HT ,GR T3].M
P-*7-M265CWV7WW3%W0'=@7+0QJ2Y%X\UN$RVDH://!H&@U4N/9W$-6,$GM0R>]>=
P1H1\IW[> $^=RU.RUU3_W;;L*JL0]549CU,G:UZ'G^$D:)(9K)2&(HA90%:;FS62
P+]*[*NACV[.(L-54BTV*/ RFR2!M</V3>G[3(.:MUS?P5^N"JVE!LW0NB@"5VU E
PO&[L_C#FQG&G9$Q5Y)E \_[[=*!.DE]=ENP@$8J8'$!0JY%*$!71Y J+UL2,/K!G
PX'I))^6UY>)A:L-?1O/K5:IO-"09-%!>/U6>0*-V2?Z!C(Q))S=32?0&+M5.&DKZ
P^O$>S=_\><%)8K;'_Z[%?(A'U-U,4:XP2MW\UT0S9+7$HH1M1]@4.-&?;D^[FI+9
P%J!L2^7['!L&"B\S:PC-\R1VV3!B?/1>P6^GY2DF,&3)"1_W$&F2QPCPY:]H5^,'
PO8\GX2I5(DJ=II[6H"Q=WR\^8">A^:JN<'.=A7<<7'I1['ZZ4DYOWL/=KF.X'HJ+
P8('P,X6J0#L1Y=,3TAM8D)S*#:)8=) T-58%;?ZW>)/8SCE(P&<*?*-S%'TX5BBA
PP&:45*=VSM4X^+75+.;,25+$8U@ JKZL2-VC4"G@R7#MLF8:=&F95SB:R]S301/:
P!A)-%UQ-JCM^6 "&8G;B]!&WU/JM-'TE SQ\8?18 _/?'A"] 36:%*2\..]SM2*9
P;=PZK["D<'-#Z]MEF:%A(WO BNEH!0]V\/B,5:0A!U35OL.&2!5I7(R(P 7,GWUD
P'%QY6G=\)FT,QU8*S#S8^_0 Y?>HO&@=Z99!J$O)^1JBU%BFA^F7O\J9FU]\OI7;
PL9C$$ZXZ&HO"\KP"U,[KH1:D#' KLEJ2S\/4=,^DMNQ>#XZ-_)_+GWHK6L=(ZF2,
P4,,LH1& M.'<T%)%.>&1,5>5_VESGV,517I8F:YCQ+1UW7%)R!K>TX!Z<DWL(%H7
P^C()+=)(3'_&SQ2_NK>EJR<Z21?Z;Y?*>GBUZ_(%NHJ7+,TZ!'C "D/._"S6U\)6
PUV3>48-&B(V)$1 .#4FP'$>5$JV"?+YY'\R7$V1O&TYR>G[*4,/@#EO+8X00R:8]
P6Y[L)W0MA7[L7:0C$J2G(K$N[>FKRG6+B8D26-?P7Q\/.F,?Z%$5='G/OZ'G!^3=
PP_=A<6A]*"4_PRTQG-ZP61+9NGI2$O+?EW+\UY;,G^UR1H(>.2J?_>X]_RP./39*
PZQ+#/+U05BPY*+2("1.T4[ 6.8M41.%S(!&&%W^'^3T>XBX5(.Q%?WNT_\=><<3D
PCK MHAM,T?JMCSS2340''L/:>>XXK<7^<Q.?[G4::>@--J$Q5G6&*;'[T)1#-_T/
P41<$M^NWJ!Y5J13H(Z@^*+ ;U(][J]-KY4Q62D0F@#0-QQD)(F@UAUGC$SFS/GGV
P96Q!N4O/HF3^^=]0N>.)7JL&1L3D2N]X5B/SBK*(2&]#P?M2I44#Y=]1=C@N6<%0
PBZ#CZG O- S:6[959?YY;?N7N*N2XJK\WGQQ(LY6GYJ>5?GZ_+"5;P_K5NAF>>9Z
P\+V=-RWYU2R"/Q&9]3HPQZ/U) V+ZX_ZN+MNF,<1KUV2.=1<SV[IY2S7^"FA,417
PXH>0%!Z6YWVFUE+GAL#6>SL["[Z!#9YG&.'4BL8U[@NFU=5&2R@X5\5["]=0<C6.
P=IZ#'&4;M8*C+*G>A*:6E%/O0+J&L?A(IIBDKPO2ID]"'Y=IJ&/K^D5Y4ZJP.@$T
PW [W81?::_GJU\&9L6%U4-N36\LQ\G]'5;SS),=("Q*=;0RXP_XL/@$N04?-X!;9
PAF&@D0NY\0Y[%^-#Z8B85P5J/8%G@S/_G2QVHKAIQ+LFO\A$>3\H=#4]O4M;(:1P
P$!8-SG!%P-W3%(ZHZ%R+>20S.%7@$)PJ='",=-]\8%Z^73,5K]6+9XKKT&7MQE9K
P7#XLH#BQ)5-S2<?&,&1-ZOO+6ODH3>-+<(')2C$#D5YKY,<2JS]]C-U3QI/L0?Y@
PI"VJ4W*!,OW1*4A87^D@5M:\-[FXE[!W%(U;@/M;0Y8) QV6+])!$#NFR<^J1*&-
PB#2<=53?O\$((Y+YB\=%VJ?EU3!4#.946 A-B5Q7Y:SKB-'4FTJ?>?\3K"*=%X&,
PJ96"IIWKH*5_TDD2_&.D";F\&;O"L<71%$&#X+#J7-!E0Z@!1E2.]UDU$,-IPQQ 
PK+Q:P.J!Z:USZG:$;?^)PQI__.%3V]MUZ_/2+;J.QQBMOEO9KB+V=(ZW]'6:2E."
PA7)L2F;2*NGX@UC&;0G;WI3'"$B5(73:.3?%[!$)"F/1&LJ@*9C_E;"2PZC%^R]?
P5+H-59/PC*VTTJ BGX.VQS^?T[<6+1"&Z#Q2+3KS]1=3 DTVSDS]OU)]9X\#/G(T
P IQR'F66I%2'\**%MI,WDK%EBA-VCF^7"=!#"2XJQ=3R%I:,^Y\1!M0YY'- 7Y2*
P;<LC(F3!/?>P5=CN=*K)4.,N*S5#GXUV]VO=]?G/^3!CHV<]^RO'#$!0&?&5(0=G
P.7A!"AR#9IKZ@JIKNZ24J6W[T[!MU8;'I<L"H' '!@Y(#0TA6E-M*[\$P$F>0NC 
PFV 0A>S*-4JVITV(&W\']E=LT<"J-6!.0_JO^+GD+M&;5-GPCQ!3V2U*3(._V[6?
PP@3;(XS->"$O[+!I?8<01I\C$%SJ\K?J8>>PM[+)F(:5\+X(ES5#RL;3AGR\;EI%
P'=MF]PGU??=!1+3E&TTQ*8R"T4^59F*;/5[8F_((1G.T-GQOT#+(+^ZB/^J(^/3%
P*7;_FUUZ!1[,&]YXQ7 J4(!*ZXP" (<\/AJUKMC_3C\!WZVV.6^"!Y)4"G=L.-N)
P[X?A.7SROKW$W=H@Q5(IKR:,W/_RW<XA&NSH:%Q7$9;W&]VW1;YL%V"Y(4GI6\1=
P,0Z67>-PHU+^'%:5>[V#-\ESS$H"YBINUWPBD*88A\/.4*OO-R #DWH@2ZQ'F7KJ
P1SG=!XKZO$[!NXRR;9"%[Z7O(5O$O3TUT/?C#I.EA<G%ZY_XM'!AU*.[[Q,%1HLH
P#:IVYLN4LKTHJE)2066P*X ML+^\+:F1W!K!>2SI?ODM=G.C6: ?3OQVX=#YE] '
P-[LRA++EG@9W\V2(X3)7/?;D,.);(?4C^CL6@4SEW[4B@^TGY],,<\2?Z?K$(^F9
P+QGF5FB,<=!>_8VC!7*8G:B+/T%5-A&H'!VLH]@29WJ_*@)FN+DI978F+R?.= JD
P<:)R;TY7#2]:Q>=^^@4^G99 X13CB6\/-KII*]>G#.A*"''<]S6[BN03#U&DV-QU
PY^WQ?-$T0X&P\"CR"D-^ZH<V,(Z5[_I%VZD!XV>VR,1C8G6$G6YE\3I'NR @1G#;
P&3-D/ZX.B;/DAR6=%PS(B.S9Q>;B&;4Y![ $8"^%^UW-1.?9"3<F\=M*Z& #"_19
PI/PG:&=-+.": U^*@M'V1. ('=!8<&/J[0.<H?X@O[WG/8D:UK2DKI"@_+Z=!:PH
P3*<VF"'XWL('P@;-.MFA6,C)3M\44>84\A2'']<D6IP'H&'J\:^G!D@$T4$RHIS6
PZ /XMB(\"MQYH%]Z^N!&[XFW($@/Z]XYW#:V8C.<3\]7A<Y21F>$A/!QM]DR8.)5
P_^AU^"X\7W. )/[/E4? 0J@1LW:%8OF1.RXLR2$O(#8!5IK?[_,J31BIQ;9%I87 
PV5D\4J!?";X!F+=*8X^.;% _9,RV42Y6WG]&MCR>3=5WX_F^^E5#5?3-3\R[7)6/
P=+6;?/R^+L-%%PT2X/QH%FGN0:<DZ4)M,Z4M^S.C<*L:4+"3XX6O8$7?U)FA+<.Y
PNS0M0=QX722OASOC,]@"T'EQ50 ++5FW^.CO@0;QI?X)H(H;6=&X) (CO/BN*=<Z
PWUK=J$"L^%IKU!@=I=U:*&"':7W% U4C3QS'(WX=%I;58RO8[**4"6."TITK5E4B
P=NR"87;)$[2<KDE5LPVWAR[<-W/"[M9D1K^^,#@,?=;[IF<N'C6GR?=EZ-4(T$U?
P0@X "QZVM._PSR'!.$\>^ 63+<G"V))-$Q?$J00!EU"=M+6/I]_EDD#BX*O)[K. 
PA5]F]"91YYB],,VQH^:NLY3OP5XFLR=04FL[Y<(.D=8HNS9B>KJY\@9\?(>"T>8R
P'7 4?#\-3J93C!RBG6^4/!RHP2(GT3Y6(KD"^?$SB_P8 !NNW)"?=PVGV-6YL+OK
PD:AAPX=LGP'9D4?>Q,$G2ODSI/=6&@Y0*I?&XR+.13/#N4<XC]O-M.Q_-RW>W<WU
P7CN%"/-U:9<9HKWV91V7 FG>-"5WPB;O_%YGADY@7<X JP8][T(XSI=MNC121[SQ
P$^F7*KTN3(Q<YTUXB)*@C2OT,S-Q@%?YV%5QSNR XU/[(F??:'H.6MVK*&*G-C93
P"PY@NEJ!0^11ATA[6,I.4_<T4B6FS5DT9Z.:@\F(:^JY(RG"2WMW#.B=@Q>  CLQ
P.MI:1!T9I>(_HYG<*>ZBTB%41;)WT'EIR(^(\C2_*>-?/0].(;+,$WE&=%%[-CH-
P.#/PQ.88XV-[;XX ;U,M?.J(#C[9NI.K=+F<O\\;./^^BG<&9U*Z]9&J)*!'"'F*
P@>[7\88[-$Z,XGS*5!&_)FHL+NT2/CQ'3BD$&$43)1D9%P08(W!KB[L]?_8C0A=8
PE/$,8!ZHB]L"EEXF<RWG<:O?I [MBT"E^7=:;EFGO;B+N1O>A[NLZ[SEO\1S_H2D
P@GT&G91<_'D$D-1[K4MD1F@6O$A ?8\5TOO"=X6C:RJB--'WUD^?EG(W>H8BN@+P
P#N_MG6P=&ZW=I9MI(RH?M:,Z[KC!;$Y"_EZ@64!TY.  YWL4!/LX^(NEH<;%6E\Q
P]B?&ZXE]/>$(Q9F?2XK\.G3+9#.KB=,EYVA1DMZMO@E*">^9U.;@=3;91[]4R84?
PG3M=N+:F/LR^&+>DU<#-S9?1NJ@]K?%A#3=-\@BL<X;WYJR[4$CQC3#<7V!C9XX@
PRL.#:F5"1Y=K>R76&83;<">NV0.[!=$PD*;O3L)E!+5HJ9WB1?;./0_"$#^HC823
PN0B9&4-)!Q\@-1OC^ELH_$AVM><]"B"^7SDIC@P9%)DM,MYCT#ZMQM<!+VGX-BLW
P>:.:;.?"4Y#J3W#4M8TWB-?73?8^H^\7>L($2^;_+]<$9A_59AW$CF =5-E/D#<'
P*K&?Y/F4*+?WSISH,Z6D8:.J):$7?*7$#:E\]T(1R?+ 25BVW,[,DX7U.2U%E:YU
PU5D^H3(I;%>^-UP20[C8<@T U87V9E'$)7VA'-Y&CHTJDZ@>Y2D@,+:,3*FY)YQ1
PM*_IM7Y=;J-<3:;?,O[ZK#D]_DY&0XZ1(^0F5^:2E$6+:LN7I<R_?Y76?.\E[9M^
PJY<Q(%',63#]1O!,*;['5?;I@;T]_ZC#].4:8<:.(""]M02@;^6  P:9/Y$7MX!K
P8DS")020)[(VW1?\X!!H&FY2]J&O_6N=!4%.P")"C[^IJG[$U@BZ][JMIFFS[S@G
P;29Z5N;1R*GT(:K(2-L/<RZ<M.E>?+@DW2MSNI'J2.E9:C<3/ K^*%K_Q->\^4>E
P#-7P7@4S':FE%BGJ&1=L87C,W-^)W3JZ'?:3,A$UYV%!<9O1YHIV,T%UGM [<.51
PO;2/Y5?$:O4(>>"1I@>J70+_>!/E!R9+8!^2772F92+^**@/,0:V!3V'*BM6@T&'
PQ8F<#G$,&0SF$3^+B#T NPI"1UNFO R%(2QMPI:D'*%98X3-9A:T:T)EJ23!>%ZM
P"UVR>_J[(X Y?:VANB'HYV"56AZF(A_[-$ ),JT/(!Y/$\05X=N\(?0D#!@616#N
P"YX6$T&5P,&<>%6L72>[Y6$VWOGT8S/3GZ1K<*E3J/F<A4HS^0)3Z0MMJED 5L-W
P6^O/XJ/4G 4^4IH,2>2[<MT<UC;TL54;1^B+)HW4,6_C&2AQKGM6RE;3E0V&@;E&
P([SJTV"2=SS;UA/P9*Z#\" 8(N%W,+:HP*.R3=:4'C8@*GT2[X6OEJ2F@5W0;*>4
P'5ZN0GEMH9UZSB_)5R1Q;?@H327& %!L?9$EOJW66V5'3WZ9@/AA0AQ$E_$>Q_S)
PZ,>D9,!XV>Q-]AQ8WS*4Y6P=<ZAN3OP-7G@0>OJEU!JANMXCHOB[WG'^N?VF&ZYF
PU#5/7:I5:O(^%RN6^*N2CBE)\'/M%T,0ZOT9A6NF4&^%S)5AGD#U&7I(-MV9&D7=
PUXH;DP!CQ%>0^/^($:@BX=U[O(:4WA5#Y$YI,C5!5U;J!<6+V"U_NL6^CD\9->0/
P[\F 5H^D%)%0=L;W '#/+/@23$]GB(AHU"56=UOZONF5FC+B)WLU%U:SM93&V^!C
P<M''^V90WC!720GISNY%U^)ZFI;6B8)PS.H2"-"*"YB.H19S>=S@ZC0<=-(S%[3;
P0*=>[5D.7WZNCA_Y]?$FL9G=OUQJ^_#0-N) /45_\(2(S_X'PD>MK]HQ=)0)A<2.
P%F+>&H$=BY6NR<QT[U='<R9:4?6F]BM'Q>#X/4K89AK%#S%,NGMF'_HQVKC?JLF^
PTC81]*H'0LRSQ?,*Z!N_-(1G.Y@6'>]TCT8"+7*ZIGG^EK3G7M$P&E#03\2[MS96
PL:RG12U.QZCH-WS:L@I,6PF6=&A^RN3WH;:1]%< GO47NDT \15P@&;@.B@UE1Q/
P)NR(=5U4@0)91187<<C"5H>H-R_*SS8P0+VRS9!3<^/+\W:MB!U?7\D]4S%']E,&
P.TM#J$5CE@*H8QD+RF2=HBI,]",[I",)A#2LY,V^*X]O'60Y^=I#:*"7O2!4M* *
P4?Z'L'@CB!\VO=G/1XMJK()'<VU_6!:SW&2S=S$-1U:F4,282[9FCY=+707%<.[O
PT.C)+TDSPE#RDQ"1@C;_VP#6"[*?SIPZ0D@^',+&&A+2Z(P=4Q/EU3 %1P8&\V4M
P%P'<KZ"F@Y+7NF>'J?(U2\^C:P.O"0RSQM?T%>'OF>\LL!QPRVM.C56+_QN!A5[U
P@,-8J@)1]*2+>\=E"S[0MCC(KC1+C$^9N?)/. I O<YVY ]@:MNM<ARH+\AX"43Z
P&VWB? '=\%:A,2C:]]"F;I1[;'_#TY5"/YS[&] 1X3/@-%DNET(?H29R8[\015'"
PK&D"\_9C=H45D3>?JW1S:MQ,H,&\3*"&5(^2B77&LK,D6;"[B'KF1'WU4_B&3ITG
P0?P3/G 9_-XU7<G(1>NQGJ-&16(GXC,R&Q2&H''B(M_!:')!V!>J;1@9\%U63^][
PV0W 8NM7QI\L%5TR:-2L#U/TV$FVA]$&.<-C5QO<"/RHX#+@I"^\B@P^K/)/7CIU
PZC^/L>*T5SG/&LU'HP?AG9!X*>VEWE5P*5?:5_BV@"3I^TO[1M=L$+4\H]V,)QS$
P"P*#0P7_=Q<,BOZ\96RWV;SP&C*(>/@J,7/<E2JYROM!7;>Z^0DXTOCKQY()C^0?
P$$?D'.7@L[$;5(;XV"@#4W#NI4^ H;O*-;Z16$5:JE*]CLW\N[DELY/^3BW9H?R$
P"BBPA!"0;32;OO*U1XYSK&&X288>7%\-2",20;>HM];A_P62]?P*M@BZK@6'WJK1
PI(C0BL(_KHO9G>5FE?SN2N==/&+I8X&IQ/4PG[*=L5YE!;\]@3\\]G >FZ1%@*0#
PRQK&7^.I&"[\Y&*<<W=R3[7+VIX>,*./PGO&3(Q0\."W^/X3XYI)I=N'#'W]\]("
P\K$6],VD]WF/*A15FY*>1F5 'Q>:FR!01OY8PK"V\P7DO\R:PE5Q2H31AGG9)< G
PN#17!FG.P99=J)1)%7H/"66D\KH=[1B5@."1J8Z7_>C%^AV;M=PS4'8U9D8M;UJJ
PW&]A'U_WA=@*D2R3'3$+LUF,B&-2S1RM$5;&WJI&!$RSTMC]'VXMA@_9X03_R? 8
PGNQN3\)?1LV$S]]T\>+6UD97<,2]_/GN_9#[/%Y'D>>H2!L ,%*CZV;7I\1<_.7*
P)CRP,:UBW=(Q@ GVN#1^UFK0:0# %L2IB_=Z9#5!/:$>?<HY/JMA'6L?:DHVI/?7
P@"!ED_SS]/5]]F57RZ34$U2Y=&RVCD'BB9QZE:!]8IRH>")R..GGY(_&3*1=),WK
P9J)!=%\V23PY:Y/K.O778A?'&LMC7*#%?-_L,[0/; 4@-WU!A5Y!,"\ZADXJ_&B#
P58P_N#5N(<:?+@]>1XP%77FH I!EOH]_/O0RB4Z8%-KPP:ZRB<JJT&U.^<;%&Q:;
P4E0N9^&,IAQ7%52)L@==3WY7D\LMBM)9F<XF#Z?TB:)B'ZW&&,U2A[3A\]EQYBY3
P#Q[BDI1-J_\ RW&70D83-)$N@T>QHNX.H,:G5D60;UO+1N3+:ILVO18 EXF9@.?Y
P:FZ6\58O-2'ZMSA)I]1'VH*(!+\W_,FKU'$0+'WPRU,O\T*?S"LYF\B)/E9 )>M0
P/=GCP_W*BQX5J3X?3#C<=4OJ3"X..E;CAB=?O:S^1W%GK"1O]I(/'<[OH<8^W,I=
PJB0ODV?)" WK=)4</KVS,RZ+U6%Q?^Z5F:&@_-PGXZ+I_5'(\+<>Q 2>5\EX):B(
P4_[T-45H$GA[#8(W6O<N[53GQ^4U*L:-"]30B$;S4L@2"P;)1.'A#T)T/[95Z-G6
P<]<L(+L(H$>"Q-!,L=##7Q#W2S/5B'.']LL%[*2-VM*;^.D6_<B,3&U.S%NF'P;T
PV=D50'HSE?%=J/LMT\!.#"D<2\3O";"1_2_SIUB$Q=JB4F^^R5F1@F]@Y".EH'TR
P,[9%&X?;\[;>"/*@YU6 T3PKHD_C5_B8+K%E#79+:V#/)].=5;[\2UE$E2?B7N.S
P-ENS2X*W,#3U-JX4-&#;4DQPRC6-DYZV#!40_SQ+G)/N7&*,'.O>8-L593P_V@*^
P(JTT':4.@S@"N/F69S,H*^_8&)E10@$6"BH<1]Q=XYBMXKY L@9+CCNO^N^%-]3)
PK0A O.NJ24*W0\@?3!Z=2*=[XZP9E'2LO1/W-8,\>,4*Q$?#".!C"P%<,X7>D[5#
PP0UG2NC@67\[<U!'IC2['H;.3B--UBC% ,-C71F!'B&94GTQ45/%,L[LJMTI=>^[
P_@> .=2-\(RCWVUD;<::GOC62K-&GS7*/=E396A*8K<T(YX6*\T5P11)HPY=:<$U
P,M(^J'L? O>(5AP1N+[M14VR&Q?QNA.ZP >)U^S%FDZ&BWDV4=6RA5\W?$"X?&-)
PT2Z^P6+NBW!% "C3.$8X-IK_XQ4-TE:8JJD/A!F(V+=L_'6-X_W<%S1SR<;\?4H.
P/&*]79,:?RRX=?UC,E[2,EZW_,0,9O\).X[Q7#1V)G/$#O?F'BUN%EA^GXH7$4ZG
P+N%D?"R3)XP0GA09% __6N!F2>FV"^RS1-"UICX^FTT&_V+53K(,S5U057W4#D%'
P_B7)UY593K0["N?M*Z_3LET4>U_'C7V(0Q<*;AE_-SY\<7OVT5(/\ZFU],:"_4(L
PVK6E72>F$>TG#<1$L(M$<2CHKQDHF,$XCHL[5U#'@&?N*#6C3 3/0CNV >#'-FJ:
P/Z7O]_F^9QCO>F8_;2,O7%,&8S&2_0 (>+XU#(\E)@A80D:_;J&H-T&#@:$"MJZ)
P&](*!U O"#/ &UM;6FM:%G//RY/C # (JQF55-SX=RRR0GR4\98Z7\":)]J89\BI
PE3 ?""[M$*UU\G?86\MN_9;Y]7#6V@N*F^9*H9?DN.?*&Q<&0HXMCX):>/,6P!;O
P&XE/%<$G<C&RQ(@'4=_JD2I0>.H8>!80WV&115A)5W=D:/ OK5:K!'%HO)IF;U<$
PCN,WI>4.(.N "[B])Z@U3ZG\(6WRTZ[3J%Z.PKM(JZWC)2 BQ!<%,E<^AJ)$9TGQ
P\IT[^3,'/C7Z;U)&EBY\^>O5XLUB>L(124_&O?HTW<I _;[C)T@X)Q%D\Z7JKJQ=
P%UY\.ZO&H [N3%IA;[O>JZ8^EL"N:+50V[]",AW8(!AWD4X$5IH\J7JG%<GVS,+5
PLS\'580E3AF4?UXN 4FQXNIL_6D"2^7G'A^A :\#3!M]IFI/I] ?(IT?6K8J59I=
P/K+5/63X55'\!.<>MWE("-A.</E==UR[2KA.IDWJO%<_L4%@.G3@],:///S6A:1M
P2*ZJ8)7C),3>42N,)\B!IX1ABOU*6O\SKT5O7%TLC;Y*Z>>&24L4C[AB=575)I<O
P+$&;EL$E^!V*/K#OGF"':P")_(<VR>.6#8RZ,ZC#,\TRN./<,AX;Z& @/S"8/N'6
PF,KE_<KA-]T=K4QX>"O "1ZS1!LN^-RJ(\+N=FQI^FG:@2('+J+**FIL1!M8Q;O)
PT*TC-"I3MBCT0"NF 0-@Q/]O(LAOX4_<&_\&GT:5YJ7V* P'-?A[I*NAT:"L*@D*
PT'C$\,BR:1V"$BO?7AR%NM #>8]P53I5S<NS A%14T/6,H3</[8_S8.#H!8W"]UE
PQU0VNWE3L!/LCXD(O8YR.7L8FC,H[EB>6[1@!EE^=T/:(JG;6DEHKM(Q&M,H4U$(
P52Q^C0G17"XW!KX"'/<K!2@TU,B_Q_PU3+0@+?#!Q4>H+C0&_CO?"U''&EW5=XF_
P%*8;WV8PNW>T&TV<8]2;+_4NY8T->=^U/;QS*I]0GHCI<E VGLJ%W%O'8)SPF4W]
P4Q'L4XR[IDMYSC@:^5Z L.28O\AOLV<E=V^S%_%4:9Y_[THB2_";O %#)TZC_7,3
P/JQ)>>GIW*:,K3JP']MOR4;*<G]3!5W(@4+8[85NW8";8KZ^2YV#%S-;'5:2EH>W
PR*PLR&:X^[N@<2CTC+D0.[+5E=OJ+<7?4+^NR:/0;PF!%U_REUKX13,:F.&XN4^H
PQ")0\D&'!%#QE9>\5H>-+\P8)CY0\'L9>NRN7.51R P%9?"*A152[G9A,]+5S$V1
P)/GF!.VCTD)0 /%^<XD?#TP9YC<ZMI^PI"C3[H&U.F_=L3B8&E=L@6. *V?#PX 6
P,#N[ML<#RV95X@=B@(R@&F=4ZIK)4.4F+0?X7!>%=]Y;]EWNQ8O#B.0UTE<T$4-!
P>:^C9I,.M)^R'RVTT\E%D$;3?$,6P6/-P$'%J0[AIR?HV=\\>7+-Y1&#PSLH/$9,
P?QH-R$!K-!JK^NAC0%2-@Y:"MO.TK8TD:9;',*)20)BB_\ #EH+/A/%-&><>9(SC
P 7(CYZNP^+TB?NI(5.(TP^!CHK> FW<<&B/!VWV*KV.CN7T'L@5KSG,?->)1NPF_
PP-RY@]2,0N*K7%/_<5]N%3%>"6RZS\C."445R=D.3YL2P=9RSQ=#5!,G7\)RIX$G
PPT%!4+RG NF <VS:T$W'EFH4\69=%'-GO50%DW_Y_V/^:DOPB7""QF3$#*J$@I%=
P<!!R,R&X;/:JM%6QY-_RT(\XS\I:8DP-IAGP32O "!# )Z83#2/Z?:QH^,[0]K< 
P+.)R#Y]#);A*__''UVZVSF.C#K8U=:2+,JLDK"B"PYZWOA$D!9[Y82,&:L8U/('0
P*/Q@PHZE-T*MN\[4"UP+!<A;\1X"OFY G%E?O\V8M1%8\&/4[T!R\BKK64FD407$
P<U*9L.6"S_A0=A4"0VA]KH!78ICQ]Z> 1I?"?3<]M3[#,QY:B!&2A>%!LI1D_^G@
P/D5^(0>#ZS=]J%W&]$SK;,GZ?$IUFX[OQ E*:R>X[KWO]?;78[+'2"%&R/,MVWCL
PNKDK:NH*.N;F,!QZ0V3Y+3M3K,*Y1RJR[ _NE7UHO!Q^;6Q+'P%F;7ZX5Z8<4'-<
P2= #C$]JDI"0F&?#72> 8,*HZ?L3VN >VHF!#0M'#44[,):HDZC1.O'"F\=50HIG
PXVHS-Q9YC0]!K;U3+KBL_^CH^<IHU)*).)\B9ZQ%JQ/G"B'KBY?31?<NN"D*>*:)
PFQ_35%+:!S?."K3BRCR4D,99:=K0I1D'>;_;"^2S$I<P?!_BH=(:"PU829 M=+'0
P02T\G'[:-5"2+52_:VAY;"2R'Y% '-;R7<S\4_! 9MU U/Z0&4_:[9(5*"  #O&-
P%+S^(12!3G<%E^$9RT9R3J2:%Z]'<IX9++4>!;BLT.%: 7,(I%%4_[DX)!T6FRAU
PPWPZ3_=I2=GT?SYN6Z*.M+BB A] 5@\.8PX+*@J[\WZ&PP9<6:6-?T]:/7V./&E;
P%>)'E3SBXL##AI\PVW]-!BO*81K^HA6G+/5<TBL9UCA.S2E>L+/11A4O,/OE#99X
P(5Q!<F$;62K'-6\C4LA,^G0_CO)DZ858[>"O# T4H2?!#!5;VS\:>OK$0^S\'X;@
P=)%8B^"9_TE],!M^0NC,$=T4DP'YGX/HE_C_*PG<G2"0ZNW)C<T%459BM55E51S'
PRI;K@*)PV:* #^(NN,LO1_]V2\<E+.%!5X^Q$O9(JDW1\X84;OE\"@J6%Q>IKQ<*
PU &S%UG*L"DJ56T#<%6U9E@".\$DC (=B76>/A]><XD:]9<M\#U+%L.UV2@8T+2(
PC9T<*\(M<E;#5;8J"ZZCN_(?? R'VO3R9(W]4)&74>$0Y-:Z#_9%3PHW*#>J.P%F
P+>IML"@3*\., CL>=Y!?8G?P_5!X'J5HQ=!>MP?3$<*I*+:)J-G?](T/D_C'^D5P
PF"W.;_R?EW(V3J,\?D0FMP.%_,#$H%U[@51Z3:9VEV_#3K?"M&L,+KM.RY7/,VZ?
P<N$4/6N&2MATTA@UK^+JVA)(KNP@>";#>AU2PO(W^1P/("&'=4,NJ6(5?] ^W6E<
P.03_=:U2KBAV^?"T0& 35>@0R:1^)"$T$K"WIRO/^Q,OW[$T:5>O([>K:^,9B@@V
P3Q1!@:&'!SFGX!+H+(?K9#&+0;.]!DNY"/OPRV6)Z$NL$&@C>XOWS2;64_&:6L"$
P^8C- C;B9'[<XV5.[4[<-8@L/ZL>8T!OYS4;Z5LKP=36*Y< )J77;"^B#>Z&_,&\
P3[ GG]AK$3+ HM]_^?!'[/674G=E*(VHE#&QU[^404KY\?KOSO')R92]UH]S_AO"
P +/U>V:(ORY_9 \S$$DIB +JY\;M# SB3\W53;EXVG1!$)4%D*I0!#S<Q@(HJ2I$
P1OG(LU:W6K0 Y+3^KA,16@0T*=D4GSC\L5Q2WS>(G""NEU&H !Y3I(Q7XPV-K>(#
P="YL?Y/7^:PS<"1#\J<1W"3W>ZR.2_>N@V71VO-WC)Q;*2# U&8U00_^R]-&SN(5
PN52Q'*ERW(#[@X^@RHME5TUJQ)L8SZ".TCR0P$-N@!_]4A?D8SGF0DB%10B23'WJ
P_#H@M87PK+-A&^:N#,J[E_25-\+2R#_RF#L,-H1^%1PH)4YL-.ED& @I+=[*0#X3
PA$]F,I7??'ANE_V&9Y]UPCB\S.B*\7O--V!PN*I@ERP4LW'AV(T92:ZEK@K(/PF!
P"CJ@RAC#T6P9;\5]^7<1K+-0^64V/@-KM,.F(JB_E76W 1S:; %;\HXWNA>&>C&/
P"7%3WY6$>VV(,*]&&,]F3X%^E%>/F6O*/@DI1&LHEZ&.&BUH4B,'T)0OE"%3C+1[
P_B]?'<0S+O)=._[I'! A W%2]<53O^16Z74SB8<W;E)WS&7)<LX6;Z3-@C+2U=NL
PZD]);$Q'G._W[]N/2="=S:HRSXEPX>'+ ?TBEF254>P$I">9H^]S,+]7GEF)#YA_
PG;.ME999;=4IJ7!B];S]FHW+&]ZN4K6X^>LW=NE:^ <6!T"94K.EI\U)#TL#_A?D
P;(G=^L%=ZVE>W!>];3-;T%37Q): QI3DO)(G"<]4?5Z)Q.>U+@"7OI([N"K9]#1)
P:3W=VZ1@F=GFN7S08+.EK 3P1 L+44^%DYV9G,1T9M38(V<F0$PXN'.XY-NT0 AP
PNM[#[$O(\BFUHEKPYF -F">K5LPS0BW7HHP6L.%?2_60YNM*_+YIL5)07DN,HN-2
PIE_>KO;T6;UI**]%(KH;D#[[W/8>!?_\)7?_NHYFPJ=_J&'^I/FO1>=)VG$KD3OD
P 2K.P^;X4WU^"KR9DR^410+A)C\KHFS!\OW5XN /)&H?^92H+S(@(+-D1QIE0$\'
P6X[EWO8U8DDB1KR8-?,8#2 =D$BQY=NJ7[P1:IZB&/H0"=?)1/LI+73U,J_=#NL=
PHS=>,J'.9EUUXVD,XA(=RAOY[]U!UGO3&\M*V'4 D",4P4('G3ZF6>VHDJ<KD]!"
PK;P<J,B\ $?3YBAF .=J'ON-.GR@F,-T?-+.XJV;>=((PM*K ?MK"YHOKHM1E+SQ
PD8R+\U4NWAOJ_1TU-H]%5$*<1>U\[R=+H!=X\"?[MR&[Z#^P8TY8_!ZLU+IIZ>YR
P&T9/U4$&(8E-EWI?HN13N, \3Y(F$_3O -WIF)^VJ.+&U8EB(D$'TI)+T=UKFRGH
P_5(4:/9O=[=Q?YA<*I--CK2'0VJ?+1^K))[!(]I+A5B>/G01?B4"+63[>K60/S--
PA3:590S/),"4QEJ"?\(IP3IWZ1-95=\EG?D@R6_+AD7*<F+2-Q)R+%50! V?GF]?
PDG&3JP8LK?"\LZ@78#'+FSY7BBG';?+)PTPVE&IIKG;#- "%]1=%$!FQ!7;PWYSV
P,HY\^&"8F3.[UY *D<N6N2_/=V_\%$\5S-44#H8130H&:)!M7^>3,=*9<[F?'M.7
PL06."Z?5S]T+=[EZ757/K,PN:A_4OAT;K?K&YT?LN?S^6!VU-@=&N]RH%>OAMG*/
P5=@**07^^FX1D)K269P<@^P4<A6&(@H5%^X!)2%@*\X4AQPL=78PF,0($?.N*%/P
P?X)=,F!>A^)@^,;]D:=P0J%K4*V<MEO8@X,C.L=@Y)[F9F3JU;?TZQGM=$?=0GR>
P5,I J,^X4+=ZXP;E#K7QOV=%?OTFV'B51=-# DDCGCC\'V^.!6*^@3"</9K[Y(JK
PB"B&(0RA#;'=1H3?W)XYV2>$[Y#\9R/%TK02@I5M@^Q/_>]1>D3RH "4FK'95-PC
PSI!/?*^JE66,FA*U6"*0%K0;;"/YAC[Q4PRN$Y\!WCN,C)U8@>6]^J$.X"5@U^0L
P/:)I<_'V3Z1XMT[ J9#OH37[I>ZOW:'6,IXOS%GYDI\O_<XH5.Q32.&&Y6+UT!,W
P>?5+1R[FM QCJ_)NGOY*.T0"XC3V-+M6+G'N!494YM$8\7O^+OA#]*9*.$565S95
P8=LE%CG5=T/=H\_4/#EGM*9,X/AEAZDK06M5V1]S06@^8T'MZR*C1T5;Z4'*NB%W
P5 2VO=60!* !/J"T66)#F>O'D]2I&)KB6XT,D@DVK:%33F08U,X+[;80*\_D=*IX
P<E"P49P:,"MZ)A'SV*BV9OFV=+>[K"\WC_\7F/@RIL T3W(A)V$(ZK1-D_0RR03D
PE^BF0XV=?,+^KV776>#\<'J$7TIG*:.NB<5NW,G;4*7P1WR9K6X89'RRPJOH0&).
P .:(M3AZ@IG/^1\.J#.GV")],=F-,M:677$X=5LBBKM&0%CS" L=_<[NW*O[^NN:
P,JM??]I_M["4S3Y"O$174/&-;6T_PV)UI11E*?/42)+[!YHUR(9!_(X32YX:!^M3
P2W=E#&L 45\!*"+)9[=HU'ZB&D%@.5& ')],Q3/46#C1%U/P2*2W7!J5H@<ZU(YM
PB92.B/  0IC.XIA?X.;^ND:;QE3LZT-[:0(U5*7XB&^02FX7_I-?Y^)"^?LDQ9(;
P=:6.FD<SF'3J]%CX&CE.XQ#B@M1JS%*>%XEF)Q#N;[[4?V.TB+!5+)C$F#';Q$>\
PTT%3[BL,5$;E4]J>)L9=X7(8N7V:X3+\Y],F?4UNCW;!LBB9'UJ6-T;CC;S&,][F
PS<$V1DEEDH '+K,/",,AX$!/*"Y"-G7="//5^;IIOC$GKVW:RIFA8[_\U>1&&#?:
PZ&NNZSU^W_^*56I$D3.NKL=%:-T("@8GM;5*!U<I_LJY3/ERV8XIECTNDO)[&:LS
P.D$>!B6'*63$BG>_B8*WSM!$E?V3?(>;B) 9CR"D&H$\/V,ITAZ$+=U*P-/(ZS9S
P.$5!3^X1=D E(H;I8,7FF6MA\!_+2-W2N/49UR8O[C-W \^S!JE\F"7E%563.X)4
PWJR11W;C BRUDG25M[478#IZ[^*FGX5 TU75'!&A#^.\!=MX2 PK.1T:32*.!I'^
P7W>Q[XU4?\_[",L8N<@=";X!?8J"=13(Q;N!!"(O>Y4(7N=[P*@6J4NC$!LMV/,$
PRW6JEZ<=7QJZ$\6$_;BAF55O6\ASD_R1E45<$Y,-C1'/!"[!GHDP0P^X/MS8BYG\
PYOFG^!M5[5(7OPM=^'=$(1/\JRD7M5*Q\#8ZQS3/11O$X://[C"+=^S2A8O+YT+"
P(2DV2'S3F2Y.R.SKB>^U!%C/P</N-9.W:Y.CH\NWE[!)10$!&X-%'@'^NK'KT']X
PR^9)4%ALA6<X*8)](MHJL@;SZ(EY&\ C1XR?]I-<>1STCD28FQ"M^YC9128>5_2X
P>:8&=_W$$XOBGF $XE3;OYX$\14J^?AB[KNYQ )&\#F?HHLRAN%"JFIV;(=I/*/Z
PW)(-A3=3&<)-R]=:"KF'1")F3L0RST%-*(I],0T8OUD#1JB#>1W)W]N?C%BGG,1\
P4/5TV>.W>GBIQ]M28>D!8#RT6)<:F5B=)1+"II2I(/S6,(2@7605<NA?,L\ZLGS*
PZM09<O6@S&U_%]ZQQQ^R)2> 0F:;\;1#@MO(H?C\RQ8.1T9F\"U7I&$J?"#!$<OI
PE31.BTR0M"W OUHLV9'=$L8BI&=QM[ *@AQ[1^>8R>71#PP"X^1L/]XA8UUF)<"K
PPAWME!I'!3=*JH6V$)0B6GW]%I!YS"B^0'PVY0MFVGXAX@T=RL8=9\04(H]N(U-4
PD8<U.3@YG//R"$L5HW4Z#&N4S>\<C[US3R>(;"8[RCH3^FN(EJ)>/M\) .B/R#(\
P!VA"FFL@H0.4QP0SO]RX")PP1 )^>2)Y+56/_/W*(*;?YV>L=H!DG%RPJWQVNJ?#
P:YV..1V8UX-1*Q!A3ES!!>=G^;_X^.67AY<.!Y6JQK?M^#L^O%GO>GRT0_M%55&)
POB]S/!: Y@0DJCL;=DO;RWR:]@T[B;QJ\\%HUER[,+DW1HL/%TV_(C.2F!^X9Z9#
PIK/?[-WFL$O [B_E/+W2M#++D4OOR0U),4"KXN-&R*8ID%S4\"B?)13")Y^H]%N6
P^0D"[O-^R=_255V6$)(V/B=1OC9^F4I:5GI@ZY&P5RFJ,@NL^>%_R>V7PK?G1W"S
P(ND7H0E"7;N3Z1F[%!JA<AT)\C'\\^'&^G66TQOF !NT9W](EW21 "#JTKJY,9H(
P6PK;_9P?8JYP6[.ERM?HP1NT>F.@8ZZ*9T#[8ZPY-)6N+V+=DT+0:.19)&XF1DQ-
P!"ZVI<#</R-/7$2T3.<G*@]Y&KBP2PX6R/TG28?<QND-:!K1#V7AQM2$WX06&)G.
PO5,7XBML18:31A;I"5Z:#WPD(LZ=V-0MJW2 (X=%&@:6LE^FWK<<-P447^FC#]VQ
PQE-SUG*B9PG*H--O+Z&L'52"WT^1HQ^F@-VA'=KNP,X1;7E[\.44NR==E5W-P(=*
P[[:7Z!I:2ZSI(QF5@-B5#8*U56O<2V# %Q]P!F8&K>-7.!0M!X-1X-CFYW='5;Z%
PQFI,Y$W<XUT-]DP*I'!N4^IL$_U[)PAI(H$UC*;HL#X50P/#$TO?EU&5."E*+Z57
P=PL\ASY<<:0M67*;^XZ07[)4YNVM#*PX341!; ^TJ1+#'PWJR\XPGL!VA*J0_8_U
PU,VS/UP*+K3504<CL^98Q8,VKV?8]D;S$>098=9>OSPQ_R37T0C-<VM\.R1Z91IH
PY4GZ5'SN;'X-M%W:8NV577NR^_Q:UF(]BWBRDKO72X%5/X8 OO" 1396CQN6P<S%
P>OXME=)K)_/_P@OF]#Y.*F+E!EUM=*$%Q55( <HQ2B5,!5-3.K;EA3!(06N-[B@@
P<H,=;(D5EKS=RV3"<+!>6*3+[23?N,I4@\H[VDUER#N)FDQ\C[S3/31W'Q$,L),7
P* 3,:M3^T &FG'LR@^Q!'OMH7@4*TNWXDHW^*?V!2-8S:;N_(+PMMG"U'<&!@.H7
PU0C)0/($[_X<XYSY&0Z_U!(/R>ZTBZ1U@M(OS,3 1(?!T49SUD!)O%NOB1[S%)KS
P'\'4$@LY</JHWL%A./6JD+<V7B[254JJU;M3C(Y>/,Z-]WYACMJF@NCVW;,JN(;:
P*'<[H%@8KS$<$/9J?"J&YVF)<N12(2W?'/A'F,J590-AV2 'D_A5<<[,17(+NX+V
P<,9Y,\!(4-M:U1M("H\5N[,-7@$<^AFW+'W4PX<K7[I5GL@#R;*13[2'5,J7#75"
P(>  1P()SK C+L\,Q2UUH^!HA_#6#$?2+'0JA6E.$=]DS#43_5XA7[C(15PUF5?1
P3$/ ;=BVP1A>6E^([A%F'M2@RT"Q<EVZZ>Z^YB_!:2C2DM4AK!1TZ@6J^.,C)J+9
PRR=Q]TA\0%G*L$1[!:!!0OJM-HN,*@(J]PG$PR6*VPSO;E-U9F/TX#R==(I1\!^V
PY=)X_)W@B#V ZV"DT=R7=L="OE*31E@WVAK.7R0TQEJUMSHLE>[U*DI SO52$>/W
P0&IO;9Q#H,KC#:&.7@+WZ'AK\,H 2N7YW]_O[=%,G7GQ8_+R<RMJ(K=CG6&ZJF<"
P$;R*O+8+XE+I1<LK!N%;$RU =/@>HZ W6Y<U.*GS)G[63?L+X[V7%7M/ :S8C;1@
P.&P77ZV0P\^JH\@3]P"\M@YPTYMWI(ST%UP]PD)<MMATBE+(I;.6Z([=I8?U)Y**
PGK31'$#[0^IU8MVP$H4M6&A:XMB'L+T[KU2?S.]@&"31,KD[J>F@5EFZ8G_J.%K[
P1+I&3@H$^5=1UHQ\XB'L"[-D*.".6+Z;4RSXLV //M#W3S\@@BWS^;&N.Y_ ZB_W
P.1BC.);_&2+^;$Y]?Z^8P:E# 6738"NFW&\L+=5LY).89*#)&W3>9W='_!=+?L#"
P?6,)/1V,E-Z4@+@C"ML!?V(]_,Y@KQ$'=H[C$,O.';]Q<):9\GA:J.?9B__5)],[
PXGS]_:I@@LB7=V2!M+UZ*!W6+S1K:7V2(<=@.83W.WJ&O<.^H>8!KJ2H!ARY@>1H
P4]I'0!C&8Y@=[8/VQ,/*K#D7#[8,TGN[C[NBS#3?;+=JYQ97WHM?9@#\A^IU<,K7
PNR($RH#VG_O!!PMH84:OAZ<\A=1S48)+A1M _,-:/+*P'JRMNF8V^&3DTJG:M"V 
PAX=@JJ[GZ8=U($;''HX$& 'YP"/;)I'2%V6=X)"KZ%620DC/F>K8\EA,!/6Y3A]L
PAQRB(7QUR!I*B0;=+[>)P_6P) #Q++*Y;E-9C//30?#(1)R/CB2GOCYG:9IF_5)V
PV>='V^X^VV9'%5GU>$==T#_?T&?XAKCNM22>8C7?>-JQW54CG<?D=8GI01:^BO$)
PM*_A >LS/AXB3Q*FE1-7J*JO*PC&6 BP ZN3*,D<HXLF;%X8#%(?\X8"3S@I*2VP
PT,_6GGY=B,O/UY70:( KZ)H;Z_GVP+X=1J'KSF-MLEN11A:6WZL6=R3SG.P$U__P
P#""0].*3W+B,'8A $BYQ6,59'5RX).5D)$%(&6+7%B[]$CJZ[P65*9+2%)4Q]UFG
PR'441969'6;K[6E:ASO_S@8OFC6Q[KCS4U6J!6FOA"-;V7V-0P*Q72H%6"-X;.[1
P\W=2K 9!> WW-BJKXP/8DM$-("LD%SE#*_2<Y56%Y^?7)Q(F5:<[PLWBUZ#K> K,
P&XE:72JH81PJ*/=2:\(PBW5:<@2+$8%9 AG[^1*U6FGA)/I[D)+G*^66\9[E3;E&
P@&?3OH)@U5-K;[@B<3K@T39,1R^[-4&P,9XZBJO\]]'O@C)Y!=D]Q?:P,)NFB!8#
P2:4*MBRPL!+-366N9M7O+)3_FN/MU5^U]8*FZ.D[:.YVY[__GYR$?Z"@YTL_0+38
P[<F,".^$9#?R[)JI$X^ML*& SXDX7Z,B*,463A3U5>6.K2.6NIK/MW[^8@G4\X_9
PY4 +(B=>$)Y4&7R0:H4H)N/*Y$4U$2A8<OA%0B>,ZJ#E65M>!A(6<S8#$7OE+!%.
P.Y_XJ"%?*O7:<?[9Y1\@ZTX:^1Z&R?K5C?GMW0::,Z^<?Y0'2AB$!VOSQE:]QJ.+
P8V?ITYU$^"7?.E ?%;])6?9_'(8G09#;N6B5].^YTTCU"*5XJ/]@U#O/3.FT";I3
P0>0LY1)A2 DIP?.HIW#LHS ,3:,)V\8I? :ELG9K'1ZVE ;7&*R___\$1!_TRY/1
P"T:_7DY?D(+1'^_9]6PI*T%A9S,WU.Y57N!TJ=?'2@$UHM3*L>S#O"&]?Z$9"N[W
PCWYH1[XOB0-@;TM-;#NW#X>2.PDC#-82$1<G*"NDIL_)_BED7B3.+Z3T6L&M_5+P
P9'_DG22M#V_RR]4'KX94=6@A%N>>[A'>M!7(SV'H$OBV+V(Z;YQQXV/I[9$GH08I
P0,Z?ML@T?)FH>;-@IO D760&6+,0HE*O/!'I,7"?8_1**'-_Z"]3CY G-K]'%JY6
PVW@*.MR*,"8'@?)DDKJ'+\9;4HC"&#]'0QNICV^KU82_@)"(RWKP-CZM+K7"%RB'
P%-,0,E[@;F8;NGLWT9[(_ ^+ M_Y!'!D,$])HZT<H9 B<F^&X0\=(XD$" AM6<Z#
PJL8U!HGDA6,9@4'K=%8R<]7X1ACS($LZ*!I.JS3LZ88 !HJUU'6![#T;]8$=J+P_
P&S'FLR^5E/K95K#A[EEIUZVT '&%1S#C%N G[7<^KLSC'@(%H#?69Z2,!DS4N>/>
P$CXT=^^VF^[[XLR,J8'-#:*9=9PV7Z;+VY<>Z3VJN.UE&=YNB1R4L187DC9G;"6\
PN$:%BB"'N>"HZK<7JX<K\'N]S^"@_$I$G3R1L-Z.VXS.@LE D$LTR1^MR?C97>30
PA0LH7^V)QP?;P\PSV'>E&HPA]^9,ECV@,U8Z]LR<KH\#M9UKU8.T_HA]]LB<->VB
PSV^>*MP8A_-RIQ?%JY6?0'"QJX41D)"[,HV) 4&OI85I[X-5QBM)D@K+MH-;=B5V
P;:,SI"ACV4=K9,J^@((1BL',A>-WV4(Q] 7:UH$@>A5:IUXUG*_]VIOZ)627(E_0
PK80N+ 7AS!;%56)YM0*4#QH!1X)0*T'Z7VYLS681 +*;(!58&\^%"+>[L6:_V>!6
PWVZS5,FWV@'S.G33@&-E>T+Y3S,&SW_59K./<R)+;!/AWB'CG13+OO9V12L&=3,O
P]8(STV%0M6CP)'TO0@>5XH%Y>]!'/[UF5PNM(^C"VD-KU2_!%BG'HA"!$UKK=P%'
P@B;0ND:\=02"ZC&"?8S;.UN:H=1R'>[\,4R)^\C3DXRFSC:!/JDZ?1CDO93]6FW^
P:33_6/L2D=^1F\H1P)%1Z1\Z1+9^:#34%DZA\.0ZGV6% +B MS.YI!D4>!JP/!8-
POK'V.Z"/OYU!^5$5D1N5*Q%_0T]PWX ;JC+4(,"\JNL,8 G=.9>5WW()PUO48Y_!
PNP8!#\:5P6H&K9)\6D3C1ZC;B# G1VU1V%',85O+#EJ"B,Q^XQRX'".[F,# /Y7U
P:DUTG7[I<\U!Q!J*QN36THESBR0WB\%5:FH0?MPI0WQ2/D!(GE]7]U$=YU.DBLQL
P\,="6ZA*-;D9]UL9EZI1SGJWY2L4P=1K#<YOXAS;(1#[GFZX#\R[9!V#F&1:BI\K
P\_NIR2<L&X\Q.L6 3C4P?]=2&#7]R:U2B#P1 /LE1WSK)E.%FC[]&A 3847;Z(SG
PIJMOE$DI.%4KG;_)*=5\C/H.(<HK_!M0DLVO\V/C=]V# DF%U##**S9AV.W,%+H0
PWAMZ.INWEQ\?\8,7#$,K'17&S0_*CG *!,[%LU"[,C8_C64O7B'\ZP7XQMN(;43 
P-<7TUBF ,Q-%;/;+54ZC?C<(.8YPKXK>;C7"X!/"#N\H.YTX\WULB0[?:U6J#[V<
P4*K8V!Q(FCVYOL<>.P\]34(=4[1GKK[?R#YSO%\-MDM^V7DLUN6=J)YR29.B6]*[
PF<]W]SU<)I!98).M4AHKI?Q49LC7H!C^,+"75%!_9$:_CH2'I<I3:JAC1A0_=DE3
P-!=\JAJVPP N"3N,,N":#G:=GZ.+X#0+\GO9Z<)3>%/$YR[44CFQHS [SN<5JK<X
P#!NN9Y(D4+1C PD*3,A$K9_LDFE.=-3+N(R8[<+)ZJ&C:_0&+7D'6#_B"A!S/3'S
PN:QV%;0=5!W ]8 2[A%3_O2<Q&%S=0E,--XB]UFW4NE\E].GD^13G*D5*B<MO:+U
P!%-0.!.'G>2-CTSGA36!^BY8NS@;6ITWW^Y?/LS?:3'WS#QSB82,C_HHOEUFYY;Z
P@W +$>1GP>8>ZSO(UOP3;&;Y_\K>AQ>!I5:B>0X,#'G RD&RN0X">D_&%J #@<"/
PQ]+F:1<V.,-;C %N9GL'HA0 JW#+I5_4\/"8HR7Z&'S33ILP55F";5-.P/JH-8[3
PT1*+'^ZG1"GZQ[2FY]'8,1\4D?!1H &3NP#T=1*8<E/2(@+.@T7)C/=+,<68CR;H
PXH!R7FR>Z/,'!X< ^$W>E2,L:L'ME);)4B=87!T@9M@9'AUU*O)U1U%;'[F>S#[>
PTMNI*9)^:1C]_&JY)Z GAG>!='!\A ;[,5$'PGM_%5L&AGL%SEH!+<_R-3&(3T9A
P[-B"F<F*;?YT Q?WX".N_SV"-&0<]]2N3)XQ/'2KGB>=/(75Q\_UW!(]%U_]:3ZQ
PXS+46:J5V:BC[N3?O")MB.G@F/J$,,EU4G4"R8]U+C@P; 3,-[.SA"?5S*OF>Y+Z
P4[1^,3MHZ$?'WPQA4-DOD- 5A9][L"<X-1A))7*$O.S\G0@>U"#-=]?JO9N-A!Y<
PP/XZZQ)E20Q">+\P3!(IZ'L>V*/K&S1^A5(A=!/R02GW;WY #UK@JT;6RF3T(*>?
P1)0&20,C 5V_?[+1QF4;,<WEEM1<G5XD*.4UB#6:^_/L3<!^8IYX-RI2B^[[QDC5
PMI@F6#BZE#LG!$K(($R+$YJW';F&W9=C^7C7G*39/J^]+,Q6_,EP[CDL+3(@IUZ[
PUDW>7M?$ ;U@'0W<Z\K>+Z'HH(I9,@8[I*^#$OJ,T'AP\UK=G(/K'[X'A@$)\V-+
P4K!EN8#92II&.N2ULH9RS%2^93T#^WS^^U^1LT6K-OI]'A1^BS)B'.NK.XX;. /-
P)=V;H/8L7&-XPLZA]Y3)/EJ8P(T_^#(G^@7W92/>:X;E&#%@8[G]/"0,IQ^^,* :
P?J_U*\M:'^$S45"5_23!T]](-PZ?*H5:6/,!P&VJ@S D,<P:'FM L'WZ>:)G4&,J
PVXYO[#F?'T0+P0>D_&'=_SAM[FU>_;__FI>/(GO,3Y.;4.1PKM$JL\[;, B+8LJ$
P0F)'#Q2(@>]]P7X- . U@'Q\&=]WLP_C7S*"^M<O$C5YT.UYG^&=)4:@=1S4I!OJ
P;M.4M$_R-[UL;C1JAEH5H+Y<JM.D1X2H%X51%E+9T!K*FDGUZ)8[P#44C$H@KQ4V
P=F<?! B(.N_#A[PYELWT0"F5#[$.0*(DSB<K6HSZG[G_"!H!(L@ZFW*VFCS4+CCT
PS$1KSX2;01!+"!? LRGV#V_P7=Y_>2)Y&Q%BLA^3/,QO@309!K!!N\(%$:8L4%YN
PT*)[EK4%[L4##I8/AZK:VI;EXFM&,!S5")VA#=P4]1=E.#'"U2A$8 @0FVGYCC5U
P24*IG_SK3A;SZ\YK@&;Y.0>IZ%LXQZ4*W\B+]1.J?9K62A>!Q]<)SO43$R?MLDC_
P*(EVSYI7#NP+RS-VUJI*^9#!4&DJ4:Y6-M_DN*[,KT:[UN6R]%/4CP+D Y%2%A49
PYBK+[H\Z1<N'#CW\CKHM22; 1MO7L-9F)IFO<CK+(E"8JU;,FV*SY%Z<00DF_[^Y
PBJNJL8*^@.YKR$]U]'A+LVO>TVD&H$96?Z!"#8(6<B![6%[]!::_)!15/YGBSWH+
POK2LY-]RQ!*JESW<=Q=N"F1!'KS26"*X,WC'O*#*L\<1055B<60SHU4YIG':6515
PQI/R?7K_+>^7E,H>*Z^(DFD6%QU9$SE/++^9J2-KJ69OKEY<PS.$LY@=YXK_8?A;
P+="#!#9[[9!<H,^VL6-1^:XF2\#_B8G4W$UD1C+C="I.]V;%U?(GC**L>*ZX5'>I
P9$MGV"C+===UP(V<5B$.+$PC>XZBDV/^L%'\1-T&+WELYH,T&0KD#,@X[QD_@[>N
PE> V' _J\+2"NR8NIT#39Y__\["2("('_@E,]([_38LO\I4<C2_23_B,'%G2K' $
P1M*IC#IJNP99T*%:HF$EN! ^.B2$98?J_:!9T]#!L>W@ =BJ0!K!<720:LDSC=N"
PCK:SQ+GKFFU%V U>[D^S"F*D7:J4=XI?N>G@*?Z2RQDS%SRQ(\=FU&LBK+PP0:'P
PV21VL?QJXZRG6#OI8.VA&")BW;@D<"?M,G( =W#RUBC,3"W:"\%JF+T%+"(+1;N$
P/&PD4)ZXF]7GJ1_Q'P5D695X?4)"^YG8L*$6>8!Y?<@J9"M<ZN</OH(">=D.*%N]
PM4@A'>7+!A'YS6A): N^7[N_3-SIY<DGGH':XD+V$B^*6$JN^OU4GG^_'=\5UB]*
PD\?.]/C=JXRG^@Z+0$.6UY6R0I5"X%+;-3@"F<:JMM5W J-%O,']#--NTY0.]<$B
PXOY;YF*2+&OMU3*M;_9]< ;9'L0'_:L;;LX6,VI;*0-(GT",A[Z5%#1HEMJ38";A
PE=L&DF 1\S;<[F,3-)NM]H?EEG<')M_AR>-1*X<.!1]29]1]C>C?_0N-L+7[!TEL
PQ;1FC^&/^:N&H"- 6;G8L]_<R(5'&0(DD&T-7 .X531@3QSHF(.MTI[IP9@)>)7&
PE\W7'B2U$'3-[L7.(RQ1BS)A]<K%R_8?#:%,H&K=X8O*"QN/7RP<2UK3O*9"J*&@
P<=T[+A!\Z 'FE>E.6>*AZ0'-M[G5SSL$ST>5!^O5\<#L#?4H B><-GI8-9[.OE^H
P)F%P3"J>&(,OW$VU,"^!3RM($5:G%S/<$G40EP<"3/!<&'R1, RJO\F:^^UNZ0^<
PI1:!6#N<L#RV,'I-X <!*\JW"D4%=?%JU)5_(KFPV_A_QY&ZR\6UQ%PNP,5Y.3Q-
PFO)-/!^T54K"Q&3</794=K^#BFJ;3O:<6&O>7TP_HV?X>P #$V: 'J8X#[\)L0:4
P<4F:%ZJ5AX,![58^!>.X\I&\*0O@3I/P;2@$Z#R/W+1TS<0[]KBX9 'MI@4,[ FK
PSW03=X6N&=.?0;RWBX"%:C>/BD4D".OJ(E/>TQXXJK9JM.?Q!,Y JXM*W*"LZ(9<
P3D\*9=HP_BG#2OZY&58!1=_ <$Z.;1+: ]_+%<)X/^ 1-,  ?68MDLH!OUF_.M5N
P,9=$BQ ^U "Y+[*UE2_?M8Z3\YMY39(^=8\C.=;4+X*Y!K*&,C>[X[R#@&DQ2C0*
P&%F],+L4 6-;-')[N\&QJF&7R _(GNV#GPOQJ2#(#-1@\\7(%]';=V,IUDW*^A !
PC-69J=\V-.:P.Z:(\79'QTG/+%)</QIW0V6[B&]S5WL(-5D>T8Z%\=19H9+>'R5(
P('K8>:!?G7A +0.9\>NNON-K*ZT%HR\OH2T6/0*:VMR,3@Q ,3:<?5@=T]2IM;>.
PK%1J<Z:O?[N/="H/=F#+CQRI6YJQ@Y>,S MZ/A3V;[-8'@"=>]'^W79>A0&S"H>%
P?X. ?G)QH$#@A]13OA$J"WUVHL[,G>J]AF]:7]V!U"[I*T^"E:GJXM]S-6<2+[8I
P%M@W(C[.KB+X/.HV@MB!8XF-[E,@V2V"H$++DQS3<E"BZ R@91,@:?RM\/&[_ F[
P2V8XSVF*GLBCLPYG]_5?K!I*=/[VO6)%@.BH3L9J M<-*<56<@<_)UK 4U#[&ID&
P%\G#<YQX0#]Z>2*&R)^/A3+=@GEZ'T:G!O%DTN/!6FR8.-<2-,;W8ZI(>8>Q/=?.
PM[\)PD13-LY!AV6:O297#06O9,BDF:GJT?>2+5H,>0J#X![/"RW1*0E.*LZ6XWKX
P7><Z?]T$RZA?C5P-G8A(A./%RZ_5O,009VZK[%VNM_IH*-#46+!O1OJ>1$E4X+H:
P<$04R!=[/AF0<MVFG-Q49#(.A%]\:ZR560)[4_+4X[_\^ B$#%YF_5^X@J)BDHT 
P8,ZY &FIK<D6Y1QK1<+:/?(3_Q88WLH/'K^SVMU__H@,342<S8Z8$NV?EPVY4>OT
PU<F$_BOU%_D:S7FPQD>P>GCQ9)N?E)CGP=^6\YF]T7DAI54K5OOE8CDO^_^>QJT\
P+5%>$?PA8B%R=PM_5Z@=>=K+,M5>+*L M1PC]R5E<2[2"RBJ,]83A7R>6;[Y1#[9
PV%FP?!N\54C%-<8A$F]-7=*A9X<V#,U@+RDT0Q9OJ)SNL+)L"U32^8%D0N>U[M6_
P ^P50[B4ZFOS]$;VPM>H2\Q:0VB=N[N5AC+#M"*A:"[^]5_@ @VT/@WM[>WJY*'W
P,,PN*>TS_%+$ZPYJ[MR(*\*-39)@31-%@T1<TJU,APP_U.HJ%O"-IFCBCP6K6%(G
PD]WLQ64U]L)-;=+*\F\UZ;?C3V_ !Y5>OO<?QP.;ET;&?&L#PK8_[9R2H #FQV8^
P$J1HM@//1D=X<'7V*!7\M9-"./7D/6;!TX(P<2^-J_V6MF5:GC.5Q/U4CWU;SA5E
P!_FC?$;T.:1QMEV L 0B%J>E3 /C@R1/S_8L?*!X*Z],$0#./@!ZJG3X MYO@ HB
PZ=9^\&2P8M2/8"F5UT90,L!I^#2=?6VJD6Z=9YM\U!$D++_>1IG!KJWM"_I'GZ,I
PP^=;K'#^%8MG#.A&EB!2FWV[(ZMZBQN7RE </H,FZ"$!N$]"7Q^(U0C"V$[$A%^Y
P-MG<RX0OP_9_%PIX 7MIM^810#@$@*]QGY?=UD0[)$HHL^%U\]3<W"#<=NR XO8"
PG1M.!7@=JSE!HA\(N@ 7\SI^8 M')YYF1UBB7B%\L<1SNXQA>)RAL'1?(P\)-'Q$
P,RTE=K+7L(ER)K\BS$G^6R'0\*T)*+/;(T]YU<^LXLH8.\X"%M[G&VQ<Z?V796Y"
P$36)98FJ/*I3&:VP,=4CT[+,(HLB+#]/+=,C2<\*$>"2+N5G17OE,A.'0:W[SNA&
PPBLT1#BBP11$DZ?  'P-R?*D_EJQ@DIQBJGS_DC"*G6_/.US"+_")%\*/X&>:9["
PU9>/P^^H^>H8X*??<6L,3K9I<27G:DCZC@@N*5.[FH*,Z14N=&#Y83O+\$=WQ)E/
P 6">L2+(.R#1?5#/5X#?<LPDXB?R00@PE/0.A]Q63IE^KE=?,N86;N&'7L-H\,=C
P'YN;'@W]@:&6)J.?Q!1+_S9XE%1>0=\;.07 0(J;&^-+JJ+J"?\ LM.+V8G95_ 2
PJJRP<X"<QNAGSAP?M[D"L6;:$(J+;S35W&3Z)MB5&[LAG79H$H)4T+S<EH*PR](D
PB7I*ESOXA%7*V51]6@@X/?,I:CVM941VG#$ (X77P+@C.JD;8KJ6,?A%* AYHNE*
P2;-+;^>DJ&J$!G)D;$4#H3M]=(S: -?[X);5O(!K,5(MKK_8ZW+!1'<,H_Q*BA27
PV^N_OR<G=,I+XOSZB#UZK?.;"0ZVM>,)E=2L6U#5ZQ/'@7DJB]5$KHX;QW@584:\
PG]^H,LO&[!A198&PWATT^KF&]D" -9[$8>:Y2SCA?)[UX:']+/M4IV8G3<D*./"S
P]YSR+"4'XH* 43(.<P6FW\*W[4E.W%8-=AM1UE9LK_V\\*KZ)FNV+GHUWH1O86+\
PA(I#$+&F5&!Q%!TMR^!+M4$,N\&B2 BN(!DO1/7!KU;A7J#9F,7BV(9SMXTQ)A2P
PIH^W6DR>]G&AOX.D]_0C^QF04<!>]9:N2,O+5(&'V(H]V)()%G(L6_W-MPYB%U\5
P5Z4)TZ;CZ&*L76A5&EY8SNNU%FF7=_]H>E[IAM-0)VR8<5M.S00TWBDVM =K1A=D
PH/N2C4YE/<N?.V,ILR&<EXK;J[0=.216+#NB$"HIEH1O!-A#L#0V1S7@.1+H\NKZ
P$;9'F?*Y.0L)O&V.ZD]2G8X!AI;@V/ :)3UC,S,L+Y_Q[$FSTY0P'+W !V-M.G' 
P[;\6=3LT#9I,#$;K_Z @#"T=*-9_6UQXK24F!TKYJCH3IPE5>AWCY%KZ?2,,>B64
P?Y"MO@VWX".HAI=>X8:A=0/0U-DE"CAY'P0HGT4HY!<OI_'?'_&1R4#LI?H?'"I]
PM9093]X,-S8;D0_CW9O=_.^3%,O&C^1+7>I]V"1ES5O;,:B/?X[*8RY&H!6WPC78
P$;,"1NH[..GN#$MB\'M*+2<W09WHK1;E&456)T54>._9 NX\@"0<7+. 3XC;#H#)
P3(H,?GZ-*6F6\?^V;L'(61?56,JC:)M-AU0Q0/9V,U)-=>\(LOO,JP UK6Q/X.W:
PZN6>M?:-LJ0$XWO30^N]>B3GOH<T1>9_O(XW]R'GDXY8H*RD=#XMT8I]#.SGB]K>
P)-;"OSK8\:SP?QR 2&2#8&RF(D- JR! **/JH 9V35' .5M23=>F-ZZ4A@8(G):5
PZ GPL2D%.;O\ 7-^768#0'2E1\'2P84*^7I<^LO))\RS(1@W(0Y>8QTYH7X<E6=2
P[6JT *,,6[.L8GKF:=X;?-9OC!- -ZLAI8BLE9T)M:VL0S-KL+W)&Y0BR;HL2[3'
P6N0,B"!$N2Q!<8H%MG+A=8U2_K<SB(8,Z+Z%[0G^L(D;@ [DTZJ&F':/]]X_^C['
P":?D!OJ>MB$-$4K#7I7B#:73WWA]DJZ5AW_(DG9$]=U@WJ!UE3]6.Y?8DJG'ZI+Q
P;<#G242QYBL>C3Z.__5+)GT30_7L',9'??TF+-2F(1@3TY(R,7OW;G9>@FO,_QC-
PADH>3T2I=PUVVAV<49W?4@!7.FB(H,37K0PJW>QXVG;L5# !\&*QST;-[TT&E0DT
P[#_:ES!C^IRZ.*/_SPCS]UC^A_GH'=ZVWC5YI?L.<485G&E:>^OBI'=W&]TVN?Z_
PA#1I[F]M;@=0ZF/[9ETV#R_>GQE#IT>;P^8=:M_U_",G=R NBZ9$"]RSHIFSWH'&
P@$6ZK$J)]=-F0T9)05F5S1&\<G7,V=KVHGW/W)_?IW9[Z!+4T_DDGBLC*M,C4+:?
PJS$4-V;E*9)1H-)WUMY;DLC5"+1^FC\257*$7DE5GDZ2JR3IHU$$_F3. /]EI:,%
P"C+'X;"[ 1JLE2MI?!3)CXAA?C96O@H&Y<$8??8K.O=-E,,Z?F\T&\$LQE7D$!;8
PWD]9 '^Z<DW >IO!'4)JC.7*S*.!L5(IGV=3^EJ"@11X:>96K#.R:0V D$5VQ8U,
PPT):AY#:TAOT&KQ4ZFUJ=8%@C"^R-*6B+(SDWL50$>V:SX>Q X-@#2!O1S)CR\!U
PO?J=PM&<09Q9OGLZ[V28-R/?R1&%O]>15<]*2KC[QC5B 3\38WJW-4)3TA:=;K>5
PJ:&LG[&&XM"I%5PL,*I<O!_]94_Z)IDK.XNCWDL@G:7X>O!-'LW)A:X2N8%DBG0#
P]]!W\MVOI*\E*]U 0K2:XLD2U9?E>FZ@+<+-$:_>*IJ" ;6#';%*6HQG(0:98V@U
P;L)B@\=*G17*:R'J8)_790XYKY(Y5)C<,YKKQ<TJ0VF'6<.$\_# B3[L'*:N UZ[
PO#8FZW0GO)8M;UJMGBL$&Z>A_Y9_^*$R;T]Q HNG8+%4)VK(%$TV+M6IOJT%-B!"
PA"[ZUL1YZY;S.?ES7@LZ%K0CH)2#UX_@"[37W'(/]\63MLS^OLI%GI9BAO?LJ)[U
P7+),13E&/-=KCT^W&,OT%(*4T$:7DV0FH QY+T^G>!BQ!^EJ.C X2(BNN?+:XN/;
PW!? 2F0$<_,[=+G+R/9QH'E3%5LB@UC5:&GX;U97L7Z]7/J8.4>RE\@#@BZF-"/^
PJ.Q6=7,Z(!XO*ZC[I#P>QR:VT: @47D%:R6/B(^*<K2\ %5^G0N<P?7L52:-6LJ(
P!.^"RHR#9U7,P0D[V%T2\+('T/,I180G$)0(?$3 RP%9)O*EA@5\JH*$DROA) RP
P/*^'=X@'PGH'?$\FN-&P17 UR\4G(J893@V.B\Q\TL[X ICY>P#<<5G[BE<%!6C7
PS(VZQ0$DL-47!3PB)AN_YL/&Y2!.>QE\:+9TGC>T+*VVA@9LRSH7=1A%.=P?L@VC
PG$!JKW@3YH"P["LB7F%A"\[&U,7./L!\U"FGI?S\G'R!*HA=? M]":7^]C<@.[ ]
P:9OZ,-%[P'8L5]>O ^8\K&(>!M_<V+-S?T')UNK3;2;+OOPE<:0(0Z.CL,X'1!]Q
PK'\4NV9.5'9MGB*JFD2&G>I7(PMG&%H'JT=XB>Y3VNS/TBC[;Q9]K-_;=8^D\"V[
P5TA0<D@E[QVS[PSTK2*:(47)SZ%3=A6M,%$!&VE0/,1%,=P/AZ>K=D3WE.Q_?2CC
P?1IFN653>$W*J";%N GH0D@(CC8B%KN]W.MDTQVK5N8K^]TO5^]APB>!Y$1+#0_%
PWEYZ_]3>\T!3('D'UZ ?+_V-"=%&W+$''%*%>L#5LM46"R[;)(FY!W,'4-S\)D%W
PW@T@O<ZRUP=;1\KT)@G??SOZZ&V?1' +.C-?C1R7JXP N:G) FGYA[;5[&0BT9D'
PD]>RY>./<7_M#GGE1]"^2T36QRMP+T!0&\:B3F^H%,RYYUL-Z*<L4!)",N$@DQ6-
P]]]-W\VP(V/?\=K6$_N_0 F2*^^^@+>+,B<LB7"8K/R^D_K \CK=%UE>AY?7-'AX
PI$!#$CK5LRMCM2%O#%)4;3$VG%P E?+ \_7E(*F_]\4R/7R &AD;)1^M][M8TTX4
P(E*V1"7[8!@L9^VH]] ?A]9]!):_7K' OU'&G2G@J=HFDVUQYS-I,MCR?&%T)A5<
PS9:]-D)=6L/'GMP9.Z5YR:*1SUDQ\HUI8KH9YC9UESR5D,YH,[/PI^!"\J1@/M9X
P)/GH]Y;IE$TT(@3>E3.<<HY).NF=6-4V^M19H$5AS D%'7!E8J%1X?$VLY7XVQ5R
P]@<"UONDW::?:!\4,:*H>4T@]L=2XJ$*]%J<E:2!5R_)FA9Q!OJCM"Y'WEJ.)8YN
P>BJ4#OZNM&Y,8/-OL7*+$8?9,X/>K/MFMW,G.1ZHRJW[0U3AE;/8=QZ6IG+M7SAB
PB89A[2[0=X\/2"]B9M@0S-I6@F!W7M,MIU!HGNK\%+"+K]]&#9)'D38=\UZ!\HO'
P/$J@L)Z&SP,L'*:TR<#IK$UVCHDOX%:O#1MGM;&3!"1X=]U#K-F.UL6(MCE#M 9+
P[LTF%<(#A_X==86,$U/KGLP4FP\6T%W4=:@\SU&SK, [G, 69H(YWN?5,5[K@W1H
P,[.P _-8OR+--R,(-M"Z,[DR(7_N&#M@&YZS"M_VE?*Z/,7<[QSV9'4&BN8,PT=+
P/*F6<UM2TG)4SU5VDYHS>/%\'Z=PCJ3"_VO,9I@H^ &YJU'R;EPJH9=0\MTX2R%'
PN'(4I) D^V!7'%4(?O1'6&COZ;:",V_J82QVC#Z[2_>,AM2Z%XE69O-*0LIT.9(\
P81J74#)H=P3%Z@$>$@QU?C649A*VY1ZL;?=;F%^*YP-;A-.*)]<R#6LH*<\;C#H=
PF!&KI,CZY8%Q&FDN/5-#^X8?*9],3\&)B,T0Q @VP!Y:B]^B-E R,B_V^VZ:XSFJ
P[@DE*E!)F"3Y1,,#Q>*P^HTTM/LU_/DB#-8P,RT6G"E4NWM)GKKNKO\TKE/3(K*<
P^&,%*9B?];5M]EH]DJSQQ77Z#GKEKJR.='&C>E7V4!9J26M9]^HISC[O%ZHJ6J 7
P.O?#";C1>/T_4/$WA%I:PF_5_$\A4N :ZS":<6#CIH\6KSED%G20LA<I*ZDI."V\
PGZN,1DVSB%IT'I\K5O[F-WW^3'OKNR$=N'Z-S-53J!/.GKK5AY\ICDX$N>V]Q^V?
PB\CI3U,V+D+3!W\6L^X+3JF).^P)!. A$I2SM'17IE:$.D;7U9(I%PRJD&!Q&V[T
PU-D)+!F&_=3>,E41@9$ON=9+Z-D&A,.YE):Z$<-1^#O:>9D6X<?(Y@LWV+GD_/.2
P*>U-ME;QGPC78&,=+TI<+8S+[V9,:*69NG VVG(97H3S^S.-O@F[:1)"DI<34VC9
PC:@RN@- ,YW2@/CG'NK<Y5  [E1@LL<IR[#S^[AJ,Z/=Y'WS7DUJ,*#ELV:NUM-'
P3Z$QN7<_>!MS&B!.96).;J5L<@*BF8G])0%6(@OA4B%*,\MXZ0DC(^SPXQ(,$Y4"
POHKV"478:9H=L.'23CKDRS(>C>PMG"+$RM(F]B:5^4C6>N;?UN4W.BN)DP7?^.#?
P6%1E*7K7N@VQP$C;>S"VFG?J#YEFNE?:? ; (Q<$'NF;>Q>J8IVAU;2;?1FKU12L
PL;3,.F2T"T%SB[(\F_<2V*)+CP%9ETBV.[/%36*[&@5['+9QI TE +]X"5H,B-\E
P*%2DL.LCU3D7_?B#SV7^K_N1DS)X#?&6/1(&ERN^7/T_!I)9%&KJ(JGSRZ;9ZPD!
P"I!B++%9 I"</0V4S6Z](O0^EX"<O3-O#$S3$JP[&"9 1+MJ<WX7,DIV*TV!K;<J
PH3H$!D97;2GK%&8V"7Y-0P/TB*^OO+[LXIF>HY#\KY_5+'(U]!]:AK;O-A;^N9*J
P/FZFT;_DI_@B ^"3_<%@V^^T24]U4BDP+J&!ROP03A"EV! 24"FYN=LC6C,6VC>'
P >D#>*1HTC1'0(%W%S=;<FV0G<$7T+ZZ$4HR6\/<%; J 6GLF8R*^_25?%>2 $F9
PJ/S[S0ZR-H#JP6F27-V6? A?GO]GZW$DTD\SF#T(LAQ8PA3<J5H$J"2,]#UO#7%,
PM(:M%8>:?$5^")'4 OK'''S3=EZ@+]CQK>$IS2$"(L\^Y$E<&M'%UM*F38#+HH:S
P;JA6L<#%=M 6ZZ".UB"[WA+8P+XPUW1H7Q5D%6BMQ+NK_W\0':2<-;$?E\IW)UJY
P;(Z=X]I4(1LA(["0UZU>?ZD8QMZ1V?HSEB,\.]%QT#[3UJ"SMJ_21,Q(#TP_-G<8
PGO.1&0L_;%M&&[%M$:BXL <3>2^B)5,^#,%M""6>M3CS-<776G6P>#XKKQ40\^ %
PJ/F&,U<\K(I'@*:MG:58EARZ:>WS]&PZ'QAB/UUM:+"L_Y=LDSOBVI9EB*-S9J"S
P$:Y)L!!C3\^TFA>4M7JNF !JR-C0T$=.^UL#H+.$*3><%BV5:VXOZE!ECP;9U3*U
PIT$ @/I%%5'\YG%)^M[TV 9Y>>:;NASR(7[T3B<SW-],LFB>-8S7B])4Z69^#@5R
P;IYH!:/VYLMPC9;";@8G/K6-;H6,C;93S%K<.-)&V%$PDF0 %W=G"= '\)0?!1&Y
P-R5$7/FU1)BZD->\\TFZ/1#%L1XDH].6@M8 ^:+LXDM7PN6AN-EC=3(R?$6?9)XC
PT1H,8^ NDB@,S@<1_'%KYFQY*L13T6\I^9LT)^2#KJRIG+)N7<1-J!(<?0UO73XC
P=I7A8OWCB2J])_ECWC'?/>/2'3UY!?3\61-^0%1%+6R]1F_(FT>+35/;K0N+@)!V
P?=;MF/176+Q?%M,#]6YLU%DDE[+NC)UTV@FE(L$N;_3VO8.YHDL&0PC=R9([Y#D8
PX4:Q>BLT XB8<Z--MB(;I_A /V?^EWU/]0MKNRX%DAOJA963<;>^%;BNU?L[ 56:
P\U>HMJZE,P.9UU6:F#&!;U7F1\*B0:/+VEZ(+ TB$W;H.?8T%<_H!)+U ?]9Z8/F
PKM*B.08.!/"6^P)# V A^D.0_1T.N%HP">7:PD3GJO6]&Q=/@_.<L_B-U^> H>&!
P?\KV C<?&W00N]S:-@[*L?#Q"K*  K,*$980]4>+K'!_$ KBCYWPA8+)+CT)^8WI
PF@UQ+I56D1Z?0ZUWX/ :.F&6/8WVU*)IZR*:RD/^\OV/#K]J,Z;LT8B]UT<J"#[Q
PL[;LJOUWLGHIA4U8@[-R!N.L]=3>^W0X/U]*PETP@FR^EE4?L=&6%>LA9.XEA-=Z
PF4T]!/H>Y]@P00VMFT_\1F8QKNW=.F%U3==L>,%7GFUJR+\W"ENPWKU#R+Z#/K_(
P-[*NI45(4.9/ +E7-MB4Q&Z/]K3[JG9V(%+ 92@34]E9+0>QA^WB3W6#>7VGG:D8
P6,Q0Y#;P>&C7IW1>O0NYDN+Y""A1A3!-] ](ZNR4X3+Q@"I.-K1#ZKE$I;L@W2FD
P2%KM,V&7= 7 &(]C0 4_Y=D*$!T=!8Z<?Q\0?N-U3*$C M\,(LTMWL\=ESA4I";6
P=*?$=I58Q<K;0A)Y=;;IRB6 E?X/;^Q_GQ7Y1NY<R0YT#)5SZ;9VVCDUK@?MP__=
PN<1=DX9/G.P/1)+E0S$^C C22/4[EB.0L/J2%YX,G7\R4 C"6$1XBVC(,..[<<.+
P!B:ECECLTF)+1:6WF.DS#M]KUKBG=A#ZZZBNPSU!3@Z $EF^; ;?59&3P6\'G4&X
PQO=UT;':$U&UI&AV8[9DX7BR?:G# YG$='%5^MNZ)5PW=14@KR+-MSNI]L2YL>-L
P#@&*=#FF[>^!=)?%9U8RS;7VT?O?-!G69;^F5\2)7(WD:Q=@]2:2_41W+"Y +T^R
PPM@7I.Z6=++.$3O(EO]>LT5(9;"]1Y1,L@FA/P+1=AC6FMM5$@7*QNB',U,-="*K
PM!EOUG!*C9SF=VN["\F_G8T>?^HL(BI-#*F/WHF$J;\G9(O1WZ8[F(4]2/)BSFHP
P,9SUS3$&,NX<>?$\U2D&8!KN!N=6L),;P@7*#?EQ(:U=WC2QES#,FOK[@(3J@SPT
PK49]E)TY74.9YN6->BAJX\^@AYU)\]D^O/>=GTVT7S78H'^22C<G*ZR1G,I#TCHW
PJF# ]24Z)3<QE+TOAX+R?S&6JR% 0\<![KEE'?K>5J-E\! ?!OI^.02^3_-1 13]
P3Z;SS-:3^HJ0BY6[TK[83_0,+L<]U1\UU#H_JFY5:D(JUF##'<@GUD30N#?/4;.P
P$$)S@G8PQP<8*3Z%-L ",_" H(_MH2RG5>?$Y_$N2FAQUEH+3B_8^2G<F^\$:#T:
P_FU/9$%Z]!VCF;\*U;R8\ F0XY@H=]KV@G[N>BM.PGK1JG4G5UQA#94=9=\..;[A
P @0?Y: :#8A"QBR8&&6>OQ;V,A.:+Z!I]_8?]I_GGR?1D%B?8 ^9086LP>#K4 JU
P57NB. 7VA6PD&K_2;Y5QL59?[RU,*W.!*IM2929]0:9SC[?XDBQ?Q7UCEIFF_EC-
P2-QED6'L^S.M@;>3,6C+'_0P'_5=*E=L0\RR_3(>I,0Y#:SX[1I@ZCI>LUS@X3)^
P+6,D IU@A>C18USW0GK9A5EJ^.C><)'3ZRXO*6>HBRA5Z D @2K+&^)^S,EY1S))
PH(?X_'=XM'"O-TUCZ(QJW2=>31#ZT4U-(+$5F=]Y$^MHM;&*CPIBIQL1\_'@X NE
PL=4E9KOC$/X<<)TSE"EI/EMI^LWL/\LTM+S7++?K(31@YX7%"B9A1*Q-K0#J9?#1
P[\BHON5\JU<P6SGYG9OKJ+$4RQ&;R0AZT9?OAHB<PO4=XM$%;W<^:*@;6R\NI04U
PV79]0&*,>IT\<C3O-=Z\B^KL>9]QDO!S(IO%I#R[,'%WS4 3V#41UA9IX&LN);P 
P.&,**EJA7V&P5K1Z.2<#!$UOEJ)?A"P.6GML138_O-$()T_QL)<(C;,<'0*A\J#F
P,)=" R"(C$'A;;P ,,6V370ZJ7FU>98Q5FN,A^*\/J^03M;"80L.[(TFCL#C@"?Y
PNF>#Z>3.)C+],?['1T!D-<P5+-W6JZ@?H1VA4#00ZD&$^G,7\TLWN"DS0<N?'.8$
PQ&'WK&NZOOE*O8VHFKAG7L"Z@8@;;Y8?KG )R*B8*NVOLZ[D#+)".*= N?M$3]CY
PRW_"]I/0:@,RTXG=E:N_N6J6G>F?A(? FVM#!@7']L_W\N4OPFY!W96DESH6+]R8
PJGC]F%HYSTKP4)F%[2T2-EJ[I[&JFQ2+4;G)P:U81+1JQ+ISW+.,3IU(:ZFQ;DBN
P@LLN48%O[<I<'"M30U<M+I+CY,ZN)>DKC:#IA G!78/KP&M:.MW?M9/.H)IRB/T"
PE.%HI_96%^8-KK^B_7!SRS>O$G]N4><BMEF-+3OOK7P-RJ&,UW[^P3"2(BP(%YM.
PVQ4<3=HEE:<6AJ535BN\+.&Z=:?OJ$5RG'J^+?CDS7&_U6 NW)!F%CKQ^" ^N0(8
PTS( LLO8AY25 IT\'S$T#>KP_^IT,[!I J&W=;X, ^XODM4Q='=#ZN=:_?$^;-3Z
P2X\A'S?PI?:E'4GXY2%RHG!(ELI/QA1!);P'S+TFS3QEEXH&Y]\"0B((+3\R60+"
P3D99[O4E[H62MOF=SNS R7>*S3\%\WFB?UP)Q(^FO"13/+=U^"S=L4^3"*)JS5%W
PR+UM)1P91LJDN&1@K7+M2S7I]?:0_-.(<""+C,P;!UPINX?>F?RY ?308RI,NVGD
P9=0#A*,M9+)%<N"Z C,X/"1:V; ZS2WT3HJ#W1W],#81P"N U,9,"[PKSG\9D:S4
P:4EWNE=1NCW0I23[(\ LP**F"%?-56?^T;?TD[:.GZH[1R]'\R@[;0FT>V'R")9^
PW)F>>EGN)N#QX\=Q[L_#Z62*VHG&=);_TO"QIOY3 J^"H)$T]BQ)_ISELE)'IS2 
P%Q/##?)EZRP6"50.Z'4YRN3X87V_8S$D0Z8@:(2@)2J2^PXR+&8 )5_+"%S?,7XB
P7J+_M2AQ1Y4@1JU) UVWR%](-8/,I4(9 ;N-F0!99!B9\2VN_9PM4]^SA-GX"P&(
P"\_KG';M1)Y]2WR"LZ=L"#!J\0;SXKF56HI,(I=,7:W-#L(OU!-O_K:>Q<UH]#RR
P[R%N^S4#T\XAEI&'4 OKJ>\?IA8^[  XYXVM:H^<[JTJ!*29NS(D'_S.9GHC+="V
P[83=KY;K,,PU8'.\HTD*_ TOF!$5-)*OE:@]6TS'9Y*3))+!9<J$6]76[R-&EW@"
PT2"OGU.OJ3[7;A65FG$<;2'C6@02$! W=<WZPXD4_0]"Y 9!A"Z%:JT[3=;]=\T5
P%K(,NFRCZJ^ZO=9E0Z.\549 /5>R4G]8HF."OOMN]NB^C2,\9^3XEQ?'IF0^H[.$
PSDL=2J*/7T'L+&-FV--RSHTYV)SZC&MT_^7SU"V7)\@OIHJ6=X.4)J?DIPS)TUVM
P]U]^\BR^5[]?EGFKRI_4E<(+NSM0H F>+!Q7=C__]/I/W:%VP/H4WA!%LGU/7=OQ
P;ZY' B"T $.RVRX4"W4*>6*\!Y7YJPG\$K\E*G?C]+Z 6ED _= V8Z*ON>?FLRFU
P:'&,YOGMF5ND/?*OFLDVQ7%)N'>F?:OS@&7K=M7DUQ*\1L+$GJ'@F]%C4S?LDP[_
PX)T*9PS.S1?:GWM=4,:T60!U(.?NUU,^]%:C%["6V9M"7V.!0.XHQ->_]D+L@HNB
P@M-.2+!^'B?:\!B7$]%A01ERUTNB!!/L]7:>+);7'5!8\1^QK"J.-9@#_"\<K$1;
P+)X6O':&X)_.I?ZIN*$L]9.>2 _3\QM;X[%%)M,)LOL4I_;]?0S.M'=]_#5E.(V<
PBYU53JA-/_6\0O55T4/=[.QANT^:3&'I7#V%22:L^XZ27+ AP)%F+G(\AA/BTA"F
PF)QH,3L4*P-52ARVK<RLM^I>Y-O@Y9GVFRVLMR:(!#SN4B U%2(Z=YC=H FO94?A
PM":Q=B%*#\7M$=/8X84 5Y7.QY)B@\>>WLO<,#UG&"F:[ROO"[F?Z=53>'3<7)4%
P\341,4.[P_0%@]2J&G@D@)V=URNR@61[E%+-#".4A<GQ3=*WU+.?@1C;<,AJ*W2M
P(Y-WYYB8,Z7!O4NAM\%0;W-K(/1]R5"*+I9'[0O,0R17HUV<&*[%5A"LPGD?5_T"
P?$KJ*KOHJXB/&I^3?V+UYC :;PBCKVE'>Z7@/+-5VWS"WLW,KG(1Q^+@L**_7"04
P_8&[WA2]%NHE8E['$1'T;4MQD+]\L TIJYI\2#I>GZXEE;A,_!*<*[<R_M/;2CJ&
P*%K-V%1<>MW!SHIA%=AB=BZ"%I_*&5JM'><MP'3.[>#2E02IP];#*>SU#FI#G(-B
PQ=0'=C:3%P9VAO@=C/(BH*.A85NJ#6&C''X?%PL!ON+%@D(NTO\KP7[P@PA]!(A>
PN@4Q")DB4[H:(FJG9HJ#@(A3#NR%'+*&8-";X;%.I#5'#?8-;V#NV8Z\-:3G? "(
P<5HA<PU*4;/G]!*\#MW&"UM0;,:0]7RA RSF1S^W@(2VPG/CBT"!_CJY-7\;\,*_
PB2%F/7_SG"A>BX/@RG:3J%3T15MC;DQU;Q)TQESQ;9WU#Z'Q$>YF->NP*XK1O949
P(L[4=RG.,C//9>K  0]^)K/ =U"L3CAUD>"I06E[%TG8+.-R-ZWHR-(OEH0>(+HV
PE,54A+/VX2;HF>47!DO<AO$V)&B Y%,=/30&+]7 \B:6C"<<M!5@3IY3>!SX:T)$
P_G]:Q<ZG.#?6WL,Y-1O'%;G$JV-)A*-G!\><W?'7L[>Y+V59ML#\*4I(WZ0XPF]A
P]0<P248=1"?X".W"^%J84BZ3\L_NH]*:)S2+C("VY<J(.L4'=-QO;5K%@G!YZ=74
P<ADO99PMZI:LG).HF3NV;N[^+<?0AP6F$S&W#S/<G1]ND]7QJ;GMMO,I6W-GV_Q'
PS3_4)C8U* CIPTU:TV2X+;@]&:53/E@F<#=-8S>;7VSW(ECJK>2_UGH4W[???B*_
P6+PS28NEQI/U+(O8LR:M@ F Q5(&GKZREH%K/9;4PS376:!5N41Z:0#++D%05OHN
P>CW9]PP]:J5XTW\6%Q&YV8L-S5"04G 4FL3='#%-//TL'S&>M:RPE7%3SG5O!64R
PW;^C1F>KVCK1F)F8<6)B"MA1M!3K?8C!#>2I,,]D0OH]BE'=5B]C3:,UP';2@['V
P(Q@D7T/F26,Z,2NP)KSZN&V@O+ 8(N!:CV*I()KX5UE\GMM:WJIV-6JL\&OC=73G
PY@*VY2^/PBSJSKVMB6AW8*7A%V;, 5(\X/@M><_9W#XEW[I]'^%_<DH^_ZCO/)[E
P46R!V=;W(@3'ARD:$\@)]8<'Z.WAI6O?]S)'M0RI=+?3/F &B7YWP#-V$,ULQ5<K
P03V\$AL9QW55+%KY.LN_;QI\E9 NG[<BV]!SLX79\7%GR;^:#[[C:48OA[5ZIF-7
P])2%&R*"SJ7#()N0LL2W)Q#@P8B<V1/"AB._M!#*OGX^RWK,01L)420C4><-_7CA
PG EPK_T2XQX;/FWB*$Z/?Q:41.R9K?#"F+!\"=TNH#/$/=\4^[,@!3%>&N6EQ[@4
P':$Z:RUGHO4M-*ITD$YIPMUZ T=U$<8'IKX%5GS-D$?&K^D\&6,4*9[E/NS7JF!C
PP^- )S>^.G].) T ^UO4UHUM>ST[/]A?Z,*K_:Z4<2LEN<SB0FZP@%SI?SZQ6Y64
PL "5=0V[P+@WO9U+6FW9JE1"NGNXXMPZ'Q7MZ:Q-OM .!J'+7M>I.*Z=,/XE'JYL
PO\6HE,])U,7=&."ZM@;,HF.O1GX089J5,Q&8PIZ%IXM//\2&?'I,#DS0,HWU1T@Z
PHJ<)@B)CM0!EJ/."W!&E<B='*;E4*QW%VIR7@U. 1&SDHHM!?*\3Z'*R_?^!^EF,
P[\+UU6J.VEX"U37SLRY7,Z;LY(RTV?LO4@<QT)>.2@4-@#/;UOPFI>'%9W?%J(F!
PU0A=$*'>%Z5A.--.'^B;]Q5O,X?1.C[B4,) /*M?,P!QJTT3]W^U+W-;]2K]CITW
PNB[$]MSV6,N26%MTID?@AYC<T[]/;$ MGW=,(D*T"MVSW[TW3L+29 QRT:B\=H&Y
P$[@Z5T;[R1@9H0X $Y.2I,/W3G[K/&F9MG25J'P0)8MX\GL2'7UB5'%>9@:Q#Y^O
PPC2H4@!K_C5POE%Q'\PD\)%_!HL8YT[^'P1*'QK+-U!-_[IF!^;X#^*!3*!UB:DI
P/4$335SM7QVLR-C[+0/\4]1LSPM#.R/O,, X%H&K90%9.RX7FCG!BR79("1T/^ 0
P9UI[I#2])=GN5/Y?^B=,ROEVCUQ3BM&=E\LW258F6"3KN8J5HS2\P8G'8R8ZRN@?
P+D'>Y82S:B#F*T*)NJG*RS+WM,96'^FR7B<>:F2J#4"OTD.KLL>Q4(AFY3'U3+ J
P.IX<#'@32(Q:/F9G\T5,X@AD/:YH1J+LQS**<\DPE61Q!> ]P0UE>/F_4D7'ZP5(
P\(A02XU8>Q$+AC*K;7^O* R6G1\$[HK0^U1OCNKAG57>P,TZFB3SC%PSN/<4:4!6
P^%K#M# 'N Z-O^VO=*.OM4Y06#+QD_C-?^=2MO:,E'E;IO_#24@.7NS'CU8-C@R<
PB4/*$K9KO4IK^Y!V,VK[,X_#.,QY,LT!^1$+[W+>O=_'O.HE-5QAM[*.=3.P59+2
P13\8TPI47>.9>_1C#&DA?H1MUB6V(O"!0=$^(:"LP8NOSXAHP>^7AN%RFSQT[JL'
P)7/!X=9W%)ABBBRPL&0+QP4_7Z!2XDV*XQ] A<CLY\Q+!)SGC%I:2S#I)"PPID/O
P'M*H:5(WF?#(;OG&A5\:,K<\[S 6GS5QJSUJ1H_'5FNAWQ,&FAA^VRI][VU!0E\?
P7'I$A6>G7[TCA>B>MH%,([X%13 B0#CO /!Y%@<3Q1+HVF+P, 5-?1W0]#98Z2\<
P5^3ZT;4'.! >8IK$QC#?<,M85!)V AKKFCZ[Q% RFQ-6 LNHJ-VNP5O!^!:\26 ;
P_@R\W\ZH&-*1#HBDX-9?U/I2Q?[P_+0VN^1Q%5\:_Y(;9@.89DJXY/AZ;MA[WBMY
P $4T]-<G7II2XL"O5G^8\V&;47K4O-KXUN!.Q\+KWS'=>Y>%R\9K?0"*5A.WK^SK
P4)#6:?1$RU-XHR[E,8EM*Q-[>9_B7:Q#*C(,3)JR^]P)9VU24^3=9)?ZP'67Z,DS
P.H/E]-#[MPPY<[S*2DO#!'(&)<IZ@@>T" C9K;Q)1F1OXX"/B)CW]M7:LZ!WY*0P
PO%]5R4)-.1OK>%KC1DK($FE8T%<2+HW(?B =>W:C/\8D!#SYMXKNO$J'U3AL4VD_
PBKW2"^?.5EP)'.J!*9;)N(W//G%C2R!M1G6Q6R<5V?T3(0'R/FXR6O0U&*EF/W&7
P2E\@V1EEDK5Q+PVQ[_M!!\P=_'R>EY5.;"NN;'XI5K2-?,TP$\GM.E^O% -AR:DG
P3<BV&O'*V3+?W9.?O]H=9ZBO7:UG-C@OVK"+' 4&##M\# K?Z:C"(>7(3HO+:G<I
P\H#68&,S8))10+DC:$9-"+=!!$#ZTS^W6-%)1Q2X!'R0?Z_ZB4;@5SHWE4"K,3<G
P<O2T".I\.S.R364W^(36=A7RFX22?%\\5PK]^D5=SXB3ZM<9LT,4)4J $''I#\E,
PN2.U:I0<^BC[8H<H\!?[=92\7(Q,!!>< N6"5)$71.82FF]^+[HYBC!6!XM*4.<M
P.I7+9H-S@/"/J*=HKG=.I!P'/M_S_O#"2%E*99537I2ED8V&:U9U%2X57W=BJ&U2
P^;FEQNU\\Z2::1/]\CUVTW+=DS#<"/P/NZM%=>"9XRL[WJ(U;R#,.,K\>60AN(80
PI9M"-^AA[)*-VK$UCS*AUD._<K3D"Q8N6'0JS%V8+-&/-HQF<&#ZRAW7@0GEN65,
PXI8)D>(9DP@%EED&4*BON5PG((^N12#5W\9Z3_U;$+1: !&4+% 8CDS^(XZO7+U>
P1=:C<I$_?H;FU51/Y>PXKHWP+C%J*:C-NJZ#DIT>(XKCG8$A&15TG'OM@(45)/T"
P8;\8P22N\(Q5SA0O?=\^]IZAPWJ;^=<+T;,L\$#.S97P<$.J[S+_)F&Y5#N+-H32
P+3I3US;]SFH8Q#*,UZE4\Z/$G]$=YBFR2]X*B%5\QJ/B81(:CP0"W*?-&SO&&62S
PO'&2P?5S3(R.7FPE/EL8[9]J6,2N]@@2]-X?:Q]WTJ0!];W[$3;*UA#8=-'*=O75
P)\IP EBA#8HK)H1I7%>WR@1R"0+3T.AZ^97>D[7JRD8U_>.N(^ [''@0U:F_Y_Y 
PV+:+HTX88MAYPQ'$-RTN*50DJR /:L6%Z$CP]+6"[-#HBO+*9]GB13_=,<$7M PK
PT4G@53WW!(P2,P]FODACME$$_>"/1C@W)]! S36PV(D7530VY?L33R.%CQ+O#>ES
PM/^,[19VEO(D.'@DGEA577 OG?1PR7NIWC!3GP"2"?R O!?%"QM,@%MIPU6K9/<$
P'4\^3^*6G7ZQKTK%OIB/[U T^YO8ZO,CG3;8CY.D@6=,K^\F\BNBB@BO^E](EN%.
P?-CKT1.4N%.&BO$96ZS-2$!4G$^ +C#E;-^;%K0/>&\M\7K8!OY^&6F,\]!CBHJD
PO+%JC11"P@BK[EGSF($'%?&?4T\6,*8D3!1O!:ST4]H:@_^V0"#II'0Y6V?%C^<-
P?V&Q7>) D1N9G5$S^#\7,J9\WPEB.O"-3TISJ5,0H*'W(JK%T$*W]I?7,TQR<'2\
P.ZX?(INXF*8GF[^,Q:1CO>?7($#=*= 42U+M)/]/I]W4Q%E4(M);^)*?/3D:5\1[
PB _<Y&='-!$:HJW=CD) 20UFZ9,KZ9]9IB")BA*0W@)>_*>W+P)@(#;=\' $424G
PVB.Y;ESI?*C!EL",$#/+]?C0U1],RR.NT!6,*1&(X4Y B0>9&V+]:8>.YQ^C6<KC
P0HJ _'V^][+MFH^\6 Z7.%Q9DB:"?287562]UG+CKTB&KYH W^B5,?G0B+3D@+;V
P (=T5)G7^:X6:* 1 I;GT,&Q['H&T*Y&;[:N3=@87E8K[N:X3I>LOK3ML0(8_MX!
P:)SO$8ZS.E0C)7GYPHO0Z!*&P4Z^'?IOL-/  RI^P1J=]8S:.;VNA1^1P=2D\C1I
P)989/#B0JDYE/*".6V;I@)9M#Y+0P)1*TW>,NS*"KDDP*AI5RY8 /&*^M.K"\1O8
P4^3Q7;"47_2J\E!C&5PC3:QQZY3YGJBS:G4?2,[N^HM51<!<9V3R4=*;2I]CNE@\
P1?MP5T*".$^T.9(#'DVSG S A1QE&%GE7-0:B5#ZWP_M@X\S('6*[E0&]([-\:X@
P3"*D,N*NLGO%VS,H>&8'@T/MHT@'$R.A?4UV,6"S1BE!RYA\\4?0!#E8MK'?#58%
PB=7(*YAJ@O&5L2#I5G=M?D&[H?:2C>')3IGR]$ZE@>@PDCF,5*Q_)KH,)>-;TS+)
PUZ/KJ,.N@/)B>UZ>7$C\O)3SLS!B4T&^>0-%*H&)KP$3L,(>Y[,%=\T=:C<@*P;<
P82\) ?4:>!&55)\S3NT3+_#NAL!!->(<%Y_61P=5DG<E ^ZO&!<-E??L2'ZJ44G"
P:$PE%RK3]-+-H Q:GDBUP QPSR!IBA<U4Z66C%0/1%O> >4%BS< \0[E7;!V#87V
P@ZI4$YY:]E31^R$/,+ 7G%B+R1=,VDA4^_!%$2?]*D/,M&J> FR@Y-A'7^(@RV^C
P-\-62KTPIK:_@Y!HI87E<9"Q8%]#G8G,]M<M5C8!MU1A:<F_L[IE?R&#B!Q1X  K
PASG+[+[>#>XZ2<I->>ZX_=GD?$^ZG^7-K+[]O\YQ;HR$-!/!=M3X_7](IZW;CBCC
PBCL]\X9V:JOF"1&'C#.%D 4VC>.N:W-C,Y+SW(C4]@Q'1\Q&>M PY1$+ZKZ6,8A_
P&P)BX>P-TDZ)K6;TD5J\IIU"6GG*J(K\%&;86TS+?6? 9^5Q,4HRR_D(<RRXQL(>
P4T>WG2;,^R["-G&^HP%+!WE-\=R'KN#Y:&0&=%=6GKEX?/2Z'![HNPLTZ^<=?9I4
P8CN>/[?\N^*S4!4/[_5&_ORZ4QL#^_H<^F?EYS]MB=Z#&V/]B^8 #H'D&6-BG%5Q
P>(DD1:-$SG)W=[#)OAZ;IE[^-J]6)[">Z![NK8P^]E)=&^VZ.L]YR<X%#]K@K9YD
P=3&-YOIV&DAS)4+G53&R,N &Q)0>:,IO@ "Q<@$YT- 'W]UO!)TCALWJIF0PGGH[
PG2QI<"^F))V*0<Z&QY!FY"5_*K"5C1Y*$Z+5H/C)"SI:8#)%LGPV?6<E>DB2WD9!
PF4$Z)1D"+:/&#<1"TUY2$?^LY/0]G/CX/Q[Y(7]=FV?F5X:I.Q:5_11X1#_H6,=(
P;6ASR\GGO7UPN+R4'<"P7=G(%'.<T8F2C]VOAR1#VG$EV;0R>58(B320LJNU17M-
P[0;<_BKA1!.EZ>P"IW7F%7HT%[&T\GMQ!3, Z^/\64BR.$H7IZB-0;#*1GD3.;Y^
P,WSZ] ^@)B446OI8KP6^/7TC>LA_IS@)"-->X_PH(A!BSS.9-)$!G^V)D<-UX8@G
P,- IZKS-0I-YJ*YLSK.JP"L8)PKL@EXOC[M<:$>"R&:AT'2?@<(^;$"1T&8K#!_#
P#J#_QXV;M$;B=3C+:VR+:[1E4),H:D:YLLT@LYP=&*+FS:2='"F)^X)HAQ9^^3=+
P#A5S5C7$!&F\Y U*C58Z.D7(-@T(;:KNF6M8B>LAOW535Q=";B45R>_M[,G=S3(K
PU+C03C%!9^W"$=V/TE&)35O^O>'.NKT(I S_!4B^^PG=QE("N[](A#JSPGVK&AO5
PW:'*1<7K%OM5,5>E^?.ZOFH@\UUYVSV#5(\&Y2&-0"VAQCQ:@Q31IIP6(2"B(E1A
P7#!S*Z06C6/])HHNC,EEQ)K(IGW,Q6\FT?- ;W#1D[YPI#KZXA<^"S%@FB\T05)S
PYK1U>M@V65HXA$H#(^N#!WY&\UN,IVS+/UV4#S^G5MMV07<+*NK;KF230<GAPSQ]
P8EQ,6YPPKBZ81@=<X=0 ?X$E^&:Z]8:B&1U? G :X%ND*2N<]<90W/@!N810NEGD
P-G!+8C I=Q8C.->U5CFZ#*8;':*]K!JXT=*X/4\NW]F=7X<M[?$2,EBG+Q/637IP
P,??E@$ VC@^TIOB+#I?K9,!L2U<S*EF#V% 1%^X3]\$LU6+W7?#E[J2,S%M(12"*
PG=3.)=.&TE0SV:XM=H_U&T(54*[53N>:3^-D$,K8\"_8F*(.!AE246! 34W:S0%M
P]JCK4!/I9'CD+6660;GNB#=G#T<2_AN-^"P=OQ6?;CGY62J,Z['KGF(5.ZD5X9IG
P)R;!ZHDB$%*R,6^M*D1,@F6K-%"<$E?@EN8LDWUIV((H7CAQX:D/I64P\2\IKLYX
PZS9WQ-NS,U?P\=?1+6K#ZBK?4LMQO46R[Y8( =U%"\3%.E[YZE(CU3B'D5:-#M0=
PM(\&Y(&A NLS-#>T@=<Y^N.P]'945:VHK-O,I_-&/ V>[O#T:KKR/=\'>ERW5=O<
P8_<!A4=9@FJ'B=;^Y+ROA=F"#."T0*K)]:GML;#4FZE0]6!\!P\MIGBU$9D<^>>D
PX1FLB.Z9;U3RR M4-NF9ZFV/:ESNBQG.Z6F$%_L^S/=B@Q/GHPX&[^I914XG2Z+#
PEWA[+A-?WQ,BK\Y\B9K[!241SL#IY$M003#.ACW-!;'Y*1X.77[F6W)<<^H8JHH&
P4BU+,_4&4AC&(*'KF;1ZG6'J6WW9\C]H:HT#B>!MR9*.P1<W&U"/O48F,.3_JA_?
P8=*M0'#@FR*17(YR+*/']"@C?$*HV@.+2E4,:D7'-8A0=2E ) )2R#IE?W<W:.>=
P2-M,Z>AHD.KF]Z_@/@S5Z_L?(5_Z@O-@4\%#)+%SQHNQV_%2>4G?IUPEY5HN<@8E
PVO(46]411"!!7YOYE#:)NC>C-1E^1]<6KA+U"G^+8 J)QB60:/(<'P&(@^]025]7
P\;+U I2_"X3MZ1HWKZ@D0E2\8 C^!I+':JVLNXM>C\82"A$9,"C2#%2J&98%J@PR
P38^X;0)7-1LG%/?4SU>Q%J)[<3*U#!/2EK-W[H^XZ97M *AWP"C GP4PTG"^2IJ]
P;G[T^]MD)5=MB-?QS S-F4WA\[]C_2&%<)'4E!!.]%2,N9'I%JS3"<MM8KO'VCWL
PDL7DW!$U2:QFF_HB^/478D??[_Z'IB0UULY#C!B)'VJT0!@M77BJ[H)N(Y3$Q#@ 
PV)229V#XU]T:4,VK3Y6: IFDJ<_T717/XO,H3Y[4Q:*ZV.(%J_?+2AU%EAL!P!7B
P98_A-3G&V)E@GCGW_\GSF]U0Q;PV(<9>XDQ<+;W/R<#.VO[EZ^.$0C6GQ:SMA5):
P8A^W@+D@O\V&,7,W8&P0!L;T4VAHL([E"$"=![^0A7.U#<@@?0 ?.B@[<)?J\U1G
PA)3*G((@0)]N;WR8O9A2F0AV_);KH-0O*BZN;)P/*-=EP:7LL;J&'=>MT:]Q0ZJ=
PEQ8%X*:THZ*-PGN@<_W]5-H-H36F71H>6L*'LB&%\W\(K7V;)"+5*G0M+CZ?_!!<
PX$-29J&/FHZ^250%@\MU<_-^65^$VE#<<8M$/X-0%20^)F$$B@SH%^R0GVQ2]CGE
P2TW+'EMSPK\3_((UO>FHG3@!G#K#L=%#K/?KQ?O9/)4G,'6M&& K6-D<@1=/MJ5M
P/^@O.PXX!ZY/#V0!PN+PR,^+F_TN=:94#<SM1?Z$8&6+"[.+0 (4;JU]E<6PCKS<
P>\GF8;UI$[NQQE5F16H3YGRM&_FUO(2XKLME1E?]1PS45MZ@,<99=Z3QZE7>"*W*
PR5# \73764M6BCF?27K:<L][35-T3]$/+:A3-Q_RERRYCQQ]=+[,6W\ I+3BOC%\
PR+Q7!+?2 JZ)N8W%NSV]80B1$YI8U^XTQ8% A $#@AMTYK)KU4#\FV?W'+%@)%X8
PC'DLN[ \EJV^,DP:>H4N<_;>)-(&MA@,[^X-01YG0MZ'_'FZU1T1+*X@!"O]=ZNS
P8U!OED+ YZ^(?%]YA2;9'0;HDHV$8;3*)1^D;JG="+WH#Z9A0IZB,85Q@3K[<5EK
P*9YT09$PB]VJEZZ:EL*S[+)%#XJ",A&!5Q94H#Y?*_IM8 P8^ZA4O6EG,6503)"S
P'H S.(OG'Z^JFN,<C@E"<;7X1A^?0\Z#92>IPCCK*E"GZ&N[:\0WA3#D$S0Q_$@E
P^<&E+5QE*8^*P]76N72C]0$[S)RE/V';@([5UN@)P7%#PT?<U7;V?@#X!1-/;W;*
PLEI$V:B$8O/9+,S+TGGO:TDT<# D&KT'%29>"F;$8'8J[QM\$%SKPV1M7+(.K\8"
P%_]PEN9/U"6OX,UAA\A;[SL2A13;EV_-<(N#?"A$*S7BZYZ1CP8H<-U A=U&GKFN
P&@'6=YYJ>?0680&2682ZO:.P;<QNT_9A:F+P2H[KC2O,X].RD1MMW,A":"",X[CD
P\]N1+ \BE@WY) RPY2IU2!3M<=(Z3&G14R1@^Y=I2QP"&M.\7YT9*](?<U#-CXLF
P3.?$[8P5B,"']KWON_$]Q[S4E9IP32>VU0JW."B /Z(Q'*U<"NP3J=4.[<U#'"I,
P=D =4K@*NPGSS?"2/)C Y9/!"?W= .Z._"$*LA=^<3KXVX9DUI;9@0>2S_.@U5J 
PD(F_/_CTL:^U&];S^*_&NRPPQZ<?R"#7S1#DY\J7BG#I*I#TP0K&WGG%/;H@N4A_
PE"7IZ =NN#8;R<2Z(T"N9^K&;:F,XV=Q!#6TN'=9RFH8;HW[=KE/%_P)4#]F.AGE
PW,_WN=U3(PL^:OU[*\C\*J=-9[D$TF[' @+"O/W>C>+IB[>B(:;GA%==/%9H\U4J
PNJ\C_I&P&,P;L-#5<+]+[_D+-'5J-AO0CVCN#.OT6H!>]9&5%$E!W-HKHFZWM#)\
P;YDB>K4D$FQ B$V"]@3Y99E"_8:B5TQ,Z@/W"*/L;5EEC]NLL J]V&C/+*"J,6]_
PLKHG MV6'I6J:J<#K34[";!D)@ $].FN"@89D'?(.@DI+T7)EUQH5>; V_-7B%0X
P_E7UJ^%"5DM":>_Q=<OW-+P@4GE['RX;%!1^KRX1E7M XKV@^Y,ZHGM5J*2.?II4
P6MMW9E:H"=;*L7T?QT;&#"ZM(/7N#L=;J YA]*%G'X]S=ZLB,8PS,<WH$+<9H<=*
P])N K5TF:) 5\MEIU;$M\XO((EI73^GDM=XZRPU6M&V-*&%FR=O-!D3;*!D'@3R:
P"J$TWX)SURA$@4*27.2V16K<AA>)YGM$\T:LBR!UQ??#W%(5)NO@1>73S-?)KF+H
P^YLG/$]%:X%KZZ=="38SRX7BAHVH]E+F&HN;_*;-5#OGBY,8A@AMY)U/MW?Y:=]Y
PNOBSH4T>X>I#T3/$1@ :SXZ,UNV+I,!Y$NW;6I0:NK_<>X'^KNV@KS2K59!^8O,0
PN:CB]<$:2J):2)=A+PL BX=+S%F86H%[I4+_UW^T:?8=T/J*^0+_D&F?(U)O T)S
P0SD@N;XT_%@IYPT[TKP6879"%@%S4!M'%>E6@,SN-QJ5O)<KOC?';.;EY5[[BT*C
P,%*P[-S'Q1O&MSVAR__@UU MM\U11Y2UQKC:]#'2^64%/)Y?X.P)UO;NGZ?< DLU
P:ZQK!5>'"O4GNY^F[#A3"S%:PN""\ K!U;.FV1J!$ RU4C2?0^D6)=!2]3G42U5'
PW$]%63JK?.4W1!U0Q/335XVB5/W\JFD$M1F8<\E@O52;@6I*+/D]%CYNH-XS,(9.
PM!JHS.5CA>O: +-+D$J,14-YC45W+78)#8Z-PB5KF$J)ULRA)$C.25WFOK,V!&3U
PLDYX]F$W]GTK6/7BG;.?%E)Q]S5)+0,KKR7S'E-98%#;#*V*_SZ\MU19DEH_Z*M9
P[_+.7\;1.&V#1[.L'4;",<1H&2IGI*6K:)"R$/1Q"UU/" MKHJ/[B7("7OMF[6)I
P0G]8P'_^ -H%W-(GX5K!;_9J<+]UGO)<P+)G--6H^SV?^;\0UBAP"Q>R_G(N%*U8
P_2TF8^.1O$%NV)LR,L5OJBRTS@!$'K^F"L%PG)B[%.3AG.J\U^*B9"?>B5<+@>3A
P94!5R?XX1('9LU6HWP>)0V0]X9N2/8T,7NAJ>,IPV08/5NKV))^=AMHG3SQ]F.%8
P"X_O14_M)Y/)ZM9.>-SINL@-)Q=JL.9?HYS?2*R;WE<^S0_3W3;D_]0->'*(E@Z9
P1<O>-8#4D57J^8935_(<B?JSDX>W\B6!MUZ?@*_NYZW"@4EA7&%)V&5HR405JXK?
PRM5RWR\Y>K7V2Y]8D#6Z-V_J,.M.:2[$.F"E*@IUOTS(J,*2KT'S$H+8^."OJ=?_
P]/+3#2EJ\"[E30]Z\^-T]<^V#K_'*1&:%C@6!*84<?3>\YG#Y()_'@3XI#5-&]47
PK%1^M3WVX-S*/LI"H<HT7M/]0*<$E_#FJG>=9P,VUP8O-)BS<+RG7X@88Z=_/"^J
PO%$AYUP@'K*&0=53%_IH'Q_MJ,SSYG*CK'J.ZY(/[SH]UREKL,)\,JWR5+GBS(K>
PL=4NR11PM;V )T@X"(=VLM$"/WDQR!UFE9\,Y)0!=N.PNUZR?L!-30MZ'AP50GP]
P>5V#0E?V_'Z+Q\$9F@;%#V^[RPPZ '*J^7?,=#1SHNF#LI@@:Y))T'/6W'<.UL(*
P7+*2[JT]:[8'O)]2*2LXX>5X^G\I.4"U!_:<BH$HBC/VF6YU:J]BKU5)A08/2!9"
P[/P'B(JX0P\E$80;6S6X(B[5-QP70P$T,X=X:=[B?\6HA;=QWW4=1_(NS,$4A^H@
PIN<^66=NAD4L0&L=3#%UHAZZX.RQQ^Q2_BY.^F!.Q44AQUABZ+HFSS8H!^3CS2:L
P5?0RC"I'$?K"C"C&WUJ 22W7M:?QM;/?=E.,9B&AJ@ZS ,I2F#FRPK_#NUVS3V_<
P7YB7P<[??@S11/P0_KC,XIL8D^'E]GSPWJ[;@4)VS:/+.5^QDP0O!=\%.221XT?E
P+H#7G5"K$ F$?SEA@-AGT0>4Q!/ZQB[7\6ZBC7IAB;Z!:7^L]<X'-2CCI3Q$2A1G
P2%3!(D NUCG%NHD]TI%?)<:7.>RSF47H<\LU %%5XY?;LW=R\>2R[YO-:#_#MY:C
P)2T&\C$73:APG@"9*IO9?%SZM+ L")G7J6OSS1;;,63 "D@.*GK'A)+$9D+Y@KL 
PGJ86'?WZEE0*CDZ)J\RN;=KR$ADXX!KTI_: !'E2C^R@Y*HPBQR.%16D>NQ@QAM>
PY_-!]+SDE'HZ@*5AE2@8][QZ(+ HB:!(?-GYONRJ!_8O(D>=X22]?,WG+GY+<KV9
PXF](BQ?=\&,BWK\N>X"HFK;FBRXZ1AA+62!SF^,.)&$-MJ$^*I$>&%(-Q@22FUNV
P$1:;87']-M)97>NQH_X>[J*?"V+7CDK4H(S<TA_;<1#E^)YG,]P85YEF3I'5^YJ(
P \HCI9 BYPSG'/Z8B:X$(>DX!!ZIR&+^1&:UHB+1L@H,]0K:P>8AZ(2OT>\=OH<T
P6(:%0]K/)FPR)Y&[E4L7Z>8$0>T8WGV(6V',1K=*1-X>K#[TF/-VA^I%H$V78S8#
PX5(5('DCW-G><6*V\8Q_%_?4>%".AGR!X.$YXS>@03?[#Y6^4=HYL:)11;TYN6_O
P[Y8G8);(MLMM>@8H$VY+9PX:I2AEX1A7[Y]!3F*KJ-[C);.6Q69SHQ\501[ _V-<
PFYVKIR6N)/3?H: JTM6EKRL4J3EJ ^$UTA4G]ZI9R)\(?M5^"*X)/'1"N/#L(]!;
P1MNRX'/H^]:5*<!AJ>LV/O%<N_+U@ZHQP4#J=&?7LQ45#LV6#,X@$NIJ%0T5(*XY
P:'\HIZXU4+YIZ)9^D&!F0R?9B#1YA]*^]$TTMKPJ^6Z#K]F=%KJ-.F$'YD4#/@"R
PI-]I=.J@XO31W9L&+Q),/+):J3^*FRVT.6,J8&>_8&X10)52)O4)>((=)D9G,7[?
P2M4R"-HZQ7.HGE8"']-Q!M%%W"CRC]?$26+Z ;N11A<G$;Z=U4/YE53 KS&@RD.U
PT.%OTEHZ/W'C&1/=I:?J!;#YNK.:)J4,TTX5?L0W_&(D*3=TKE:Z];5)D2525/<(
P0YLM?$GT@%C%VJ(^>-[P .A$LT)* 3?]#U*G28@2-P#CZ&]]/F6PVF_O?$VM@):N
PWY\COF6V(,_4]RD^;G[(V^;V-V,H_>5P=EK(_OXM7\2?4\=SZ;'\0)S)3JQ>@4MD
PSUWY4R2I^@@-V?02#DY@AGV6\9[:2EWL]H81W_[0:31KL%*TT>ZX74A'RB@]U&Z-
PXWMJ3J!M+<DQH,=]2O/98'0! []Y=8=;M>TGJQVN,;'_F:*5PWGE3E+4[*JG:0N.
PK$?)V870I*O&:C;*R!ZIE)&F($B#N,3_GJ^#G)-D[$0[ @#=JB2[(_4\0MXK=TL^
P'D)M7J8*-/2-1[KG7[ZG&'VZ=407O&D71R;DJ3RC<E*(WUBC,:E()+'\JFF0AARS
PN%=.[LW=90/E4AMO_<E&E%[O[[^#1CZ92QU#&4=Z4QGG]CW800TZI7$+7$EZZLM%
PQ2&G@5E C'GD?<MV+!,&V]U&RN:JL9>J,0O'NK(SM2^W>UFH1LDUH/.PM!J$2\:[
PP/)0[@B*;3+ ?>$+ <__K!J;?KR<@_Y?94+5-<^/30<DC\?*$D4ZG8M550,P^OQ<
P[!:?&$JW$-"KW</@ZV7GQ]$7S4]2QN&NL++O#J1>)X?=*-<7FARAKQIW>+]#&VPY
PF)?*JT,&,52@:H/EWP#,A(=T -4S;HO61""F;\IN1:'EI[6P"$$G#$]P\EIY)Q =
PPL+;#MQ"D5&<YX<E#.*6TULH/<<4.E44,>UT,**_V?-1,;0C5@B?RZMG-%2X;%1U
P!9I=,D%''E[Y]X=&1H0B0T7I:UU HO)M8E4G==,/'3X\N%OZP;7&L0\SNO^'8M#9
PWA8(B!$;+NQJY<P )OX5SUS*1.4<J**#N*>5020L]VELSYK_BD(-7N3_VQ?PDXGL
PA+0/I7F6_HE V1.NGR1>XDHQUT)+V#H@!"$@#$N9I"K=_?!;(0&:+Y>O$I/2HI5*
P]]##C;N+]Z)(6W6O#&X%CJ<#P^:8*/2YU/:7G,F>[ZGQS])B^FKO[2RRNAP66@F/
PZB&U;JEK28O(;]@71]!M\V<N5\--]R DQ/V$*^CI-@41N-)$14/VJ(HQCY$6RPP,
PX)MELR62H?&1CRKN"(F,(IWV<Q)P&B,,H<(2\+I4M]D7O6,.BT-^*#/DAJQ%+:SL
PVOOV\,=U7RKX/$LU654YR22-'*;ZN(I,&B/08C. !Z\@$I&N,@?@.<')H$MW.Y&D
P/4(P&457'J'L;GS\>H<1,#[%">1;T(<'8#&"FDV0NTM.R59+ D($-[_CPH3O".\$
P0EO*&OJA:JWRKJOH./32NXOCX$0W6;#'4[4":F.:ACMJ9$4KUD7%;QUEP!HYM5VJ
P=$W8^Q>H_8RQ>:3/E=GPD=A&8@".Z.3E'N>A"8AVUSIXM>\&G+T&.[!HVM9.8SL@
P7U9TU*K <^NN)AQHH)*X-@CU=WIL9Z/B( SO /UE1>>HAU9/.M\[4R%=.<;7.ZSZ
P,9TNL2P>*5, #1Q-!EO8(8M.$(7D:5="?AA.0"G,#I]6P0:V_>U+0Q?&JL2G2TY_
P0(.MVOWA-(E>74-WLA1- O&W+3";J^_4HH80+%+ \RRR;I.Q"61[<&+U%P3%&@K]
P0IUK63CXK[,8Y*5<GO._I7R^SO+L93GE(%U096I.H[L.'G-\@[:93T0-4=/&+PPL
PHUK:M+YMC+4-55'/4>K("3<9'JZLWR7)>J!/BN9JH)Q.P):RGTFY,.,]BY/P0\- 
POBVCG\L>Q<UBQZ>"*_?G9PQ4WNA\LA*SKJ/'8ZJ5.60Q;T.Z"Z/UQ7DP79$097V]
PLQ19*UXT.62PC*QI7-=:#U0&WR@'#3P(<F_<CW=\%NZ-:353)IKW+;SN@<$ACU<J
PA,5;'"4("<(XCGOF<!6:-@8U3I)E-$G(1RWH'^\L[=*Q+%>_+,]"%(.S(,\W3FL$
P+:*;%@ Y^=(<_6)OM>#NON@$TS+Q-6;6HM"[S300V6\7;\G+KN $5U@$UV>P4K(F
P$,$;FQ-^V>8=C?5'V!OB],>RM@@@X+X-B%H+9)3"+*O4A3<Z(\2%G^!<&GL,M1!N
P"J93@,5;>$[2OS[F9C;TE%3((6G&FUX%>CSSJ^>\*MA;2EB@L/ UW%J;-C!\0>,C
P_#*L>?6?1O?!=K;8@'B!1^B3!#BU';1[2*;.^I'='TE&D@G8K_?2<GS4AP94D ET
P+>4G+01GJ6B&>$S^5Y1CN)0"8!!?KS@ZG<K;]G"F%F4@7NRR8B#=AO )$QQ?Z3V!
P\<><GZJJH^1U(]E7$],T*#0*QT^-S$PJ,4O -=<_?*<V9M);D/@4VIF>[YI"9=4B
P\)O+"GJ]2/^+AW_]A$^''1O?VL1-_HFS?Y:=%]7QG)9)#H<9.1>D[(9HHJ.9GCQW
P6=!*TA#<+8^V)1%!O,.V8SN\1%(@60S*9Q4O<\7L(=)5UT(JR*RR 0EB=*BRB'Y"
PU;>A)7_3HUP"@!KY8I<K/_L*N<!-:@MVN4F,(ZD(9QSLY_KTC5'T2E(Z@2&].3Y:
P.0"Q"SV"3*N'"!V(>ZP&1&^RF>T#ZU%F>9]"(H?*G^Q$MKO;+#JNK/RP 9>%U(7J
P>Y,&^V V#?V[!%F5=SJ2RI]!!;*I!@B3LCM(X/KF<UX=_8Z!A?C>(PB=L4;ANA= 
PLYH:PYBRY6I*2\>4JI1P[ ^9=D+W[^;V'[)5FFV4SYE@#WE]+6TD_:\:U*S2)ZW]
P(@6FZ0*(P?)Q(4I;.N%#G*K"><.0Z+4%A$L[:JO/DN X)1%>J']G]@[;B9CH+Q+,
PRJRGGK\DS("9YI0[?V- (/DAIR,J$F]3TYN&/"K4Z!\O'*;Y44$2C:6AI)O0;?Y]
P?["S^6 &S"&.^)Y=E[<VAX/:%-K-6LT"[GXPOSHC(O!1Z)B$WH5%'%UWTFY1)]0X
P[+E '$3G@=\8N4D*1GA;E6/MH"X%VGQ>WH[?LIO?3T!/0 'JU'A"%:G -[FNUKLR
PJU=?I"*C<J%TNI\'%/;IZ4QFDM]LA*DDTH7*OAIL2Z7=0K>E8)L^#]5L(T9O':U%
P2ZY*2?9M#?2MH!ZK/G\#O5B7!.=^;,L.\X&7U:[OH;)6W]9H-6X"IAC=H;@C7Y1I
P40H)A9YR>N#MQX:+X#,\>C&U87(J@-$?^R"H\VKKLLHOSA/K?J]66>Q/$?;:G,:7
PT?T6%+CZ$O3* Y:-!,"EU3_;<WQY%S-"?N\3WG6QEGU2;0I"I&\R\.8E)^A&Y:N$
PA@+_K@CL R&YKV$<I,.)M%+/W.3/'O%&+01%O+K'A!YMB:+6>V"OO&X&'LQ F#2:
P$8"A]3XF.@%8JQ[C/?%L5L6#XQ;$/ZB^3EN"]Z/,#%KADW[SF*X1Q(BK@$72#.%S
P5]PZN7T+<IR/%>@,+GRZBV'3C),TB(4,7WG7?9$LK:H_*JC9UZF,,L2!^A8E*N--
P5Z&??7,4=H$TC=;W1V#M6Z<8$.L9\.[SF@Z+L8E4-O#]MSCK]43'5)2C&,2W)<<>
P;(!<TM!C%53_Z:3EKP:M7??2F(D$, =HT6@>]\4)9+8BK(/N(G.;O HZAX2;K.T>
P0O%&(ECX&%/($$0%Y57"3TP8[Z?[_?"X'%0Z8W'6FZ:T_?WVH#.NR'$1\YFAA56X
P'^/6-YK>,JTP2$4JC4,3&$V3F^NA(O<9YZA/(#2W*.IT.];+A0&M DR35['I3$NH
P#7R*.7OIU9,_G*_;RYEU<;%OZ?Z#&!UJ%VF<V50J(7@L(GO2#Q^OT!IJ@ET$E3X)
P,N>C7E%=7GF0W(&:.#U+=TJ:/ZPSE@2S:H)@95<\M[6C N?Q)!URQ*-);KM8(F+!
PO>! Q3<[0:1N<[FG%C4"=!Z>0-]DZB:$$O_H)DM-U33EM\$8W.^.;@/#%/US11( 
PMTO5+"6+(\OS&8%5.EBFTHI?6J#:_=0<R1TI!P1Y&5(8Q?P.ES08_D!/#ZV?;CJ@
P(=']H(>P"8Z#=\)"^'LS/'^?R&B2]/!M9S++CE?EN6DZ3]F3Y.$V=&JE@N>8,"*U
PI'LA6BQ%;:<%/',(["_4UEC>?(E]S$2!(@*36E-W/!A6V0"#U;D/RBR5.8MLP9H/
PZ*FI+2G$UPG>(PY-65$116%&%8H.0[)@(4-L\2;,B9#!0HB013J03QENR^/J3H#Q
P:/-=9>-58-7"!@?.5>32(UE"3TU84NND 4]Z=LY6=G$ ;*H)[O2"-]-:VN/1KI20
P;[^9:UH?WQ%B>WG#XL'KB2M%:ZEEPE*I(OBRAT@*I^.:4-VO/,AM2YC+S,?W@C?4
P8U7KNF0LF)IM?#/;-Y-BSG[&=3JEIMFDYH\UD;<738 )N4%9 P8(9#0\5%73AI $
P_N)'0_ >."J9%U#X)_:=%7L*/6Y$5MH9#F$J[C']*]?:HH3<.S>/D##AW+L)1^8>
P& W7];XU<J%(0:4JA%1/,--L>"MJ^9$0,E95?IA? =C3SH5;.G4FXN>UP!D$Z5S8
PY8SM(=%\.NC4I_APY[5/-3#VVKV_[U\N35E3)5#%%1QW9X9U 3T?%R<!T09^.1C#
PO*O:>7+.JY&L%Z7WM2GKN%[%0IS(&QU[2?!&;B NQJH(>0I.&P^YZ+VC2[: W=&/
POB_!)C*]OLHRW'D03*_!Y9O$V*894E93- J,HAT>2+Q;X)GL>:E$.:O_]U>E:+=4
P'3"^+5@'IG?SXEG \7CCQ"3D.+:3>DX&891Z7O8+ DP19(#)1&?T&]UOA64@2YI3
PCE0DA@&#8NQ1:Q4#0IY1>8R9^ 62+ ^CF7]Q'6H+6E+6#T^7M(/I$1QZWUSY'BRL
P0^UAKJYYC@;^=2[E>7Y.7OQ=E)'ZI =I\M"JY]RU>!:51%*YZH,@)ZSOP8"9SX=]
P3RN#GAP474AX=\WROT:RXA (0'L!)LI7&$VV7Q(3/]N(^0I8<Y@0X+:W"*LYP'A'
PM#IYQ_\&5$6.:;F&2*:B[(2'_OULBY*?<X^B"R9Q&HX# 6;2[?CV) 2<!*@(.B6X
P=B=QD77[=+0_,$)M[T,./$(%]78'K!V@I-?R;]X$?]7#B E-A56448:>O="NV_6U
PT*^W&6*14)+Z]5I'F,PS<=MI#4>9O:&>"W+O><4'R)TTRJE.W1\0,5/&\Z97(T07
PV4T/C!ABL[7/J\%>CT&% N9AA.'@@!D'\_F+.UV+VE'[SCLNOQ)VUS9XO-<_E#66
PQ=4V$'9M!!J+PC,OMX]GC,)/<._U_W:18VF1-4!TVM25+2]<PAX;D'#V0QEX((DX
P./''_&@67>.&8B\;]4[]K=-)=7]?!VC(9W(!1$(W-$:5V43^BO::_@>A.Z&^/8(_
P=^6*X@%6'AS2\?Z-725ME^F0.85<,HG#-Y%$LCQ_M]IQOVCW'UVW!B#<6Y#IP3I[
P7?+*JC_H!/L/1PK%E3_3QO.(:9>#2CX@@H7S-5@>D_KV1J@.6(2FL);Y;+N?]%8A
P,:%V6)".YV4^[?OH!@XE/\="&P;*1TAG%, K .G_5IH-KMAR<([^!>X%+_4;,>HJ
P,37;RVR/G#=JN1=58^S!V^>;E0ZO8 #$\MME/NA;Z?IY[%%?HWB*901F:"("3C:M
PH'YB)+G^,GQ5Z11LC"NV7#5W#5_,6\0<%H-PH17X?<D%!73O &7/R#:]?:B?3M\T
PM<<%"M_ZRRQIH;S-P7\'UM$^BVXEU"M-PI<=;HS8R?"C*1%RG3>3$W+A8(S7C![A
PA]Y7E8.- IKTI[1,5KZV*20EBIO_W-3/Y(!?%0PQ_]7FT[4\AA)<I)XB^];7,.N0
PS8;@2)A>6Y"BX56*>QZ_$4]_PVKUOB+R+[D@FW+QZ9 $!+S7?9P4"?$RWGI2:'BE
P?\!<X)GZ=M\;L@3JVE;2;]< SM0&%WS_YHW5DLINS$2%*%L^RK4^.<'T7#>LM\:,
P.#YY:\M15."IXQ+!YK0A$K7UXIHD[T52I752_W5W8'/>++N4!X!E:<94V-!B9'5D
PL!71GH$1J'QO$Y6!/'+(,JQZ.PE""S"Y"J@+0YALFURT.1\4[0UZ79$[TVO@:2YD
P\!MRPR^(6M/^R:C>4<J\,[TF]_$8)E:'RZX6=LFN"*Y-,87IO^-W?00K)H&-SR"F
PK+)*SH,H^<'2.T*N6DK<=(*^9)33+?I0U_3R=$PAD^1T96\>8!BO_?8^G63V^3&'
PLRXR,"Y8QD[1%6D*3^T38[(TFG?TH8-RQX-:;2@ K%N[0;T$_*^J)^QGE4DI..&+
P\(V%1!0Q!?M:2V>#2<C@E U?)[_![/M9XH^ 5IM^+L(T-;9E/>LT8.-3-GL:X]8 
P/9R=L>NBK]'1.S\*P.1(G'ZHDI30RLQ?>WE!-SO2)@.952J ?X%P-<->.<SQ7UY/
P$S,WV[;['/><'Q?Y@W'1;6D%?;I4 K)]+@9,9=^H?G _7QX(.H<^@!5 Q4="-KK0
P(J?)YZW19DH9#,;ML#\$C*9;SM.JJ$W<U7N%_UT6G\GQ(<^A,XA<-S]!Q,:/=H6M
PL4UFL7'[H9I".Y;OSZX[C4A*$T&KP**.GDWKTQY"*!EGY#NI;]D[BEU 3!U1O (4
P8M]6!$<==CAF4#<:DY[)4C3$KE\Z44NP#\FM(B\KD'S&%5.6OX3KT>NE@GV:0S%?
P[1\H!)..@D#)P15A!>))U#I!GCV+:ALI3?)5\B+9$TDNJ5</B7,#P3BIM@?_;^M2
P'>&>$*["@F?V@&!5;!D4G(FQ=BK$E1UG9<XC:V@- ?=FC']!;,+^-.?J:H_%>)'8
PT\H;FR'9&6N2C^H"F$O!O[G4[,'<=N/V)BTZHXE-FU"+O0S@=IMCK<B-_'K1O/.5
PD^5&#ZF]"-,Z&L\M!L^Q.B&QVHX^VD0_,"L\+8TBW#X [,L@'7GFE5>$HL@.CRRK
PR9OP4<UQGUCX* P&X^'+RG1J7?=F-O_ZIA\Y+0=]=61;Y5$ F&D(LJ/NHA(4()W6
P;2MB0WBRF(ZK/>HEABX-?SVCMX<!=B+[&K!L['B$=+HJ1#,NS92/I8#,@*;QF]J-
P"TQG9US^6 +PM["+7K*[8[T99VEF'?U' B*HFZ[T/$FYJ'9%48EB4,$KV+FKDAY.
P.2*,^!JGHT%4S$!TL,?E!2D&:C%[Q)\"W&U[ 3YGOO'F6# ^#/FD&DH?PUWM>.& 
P%$_2NU8?QD\*=IHL)^OK/:G [: !7+S/H#/R8ZCTY93'> 8TZN$&]^5\%ZO6&G"H
PT8NKN%FI$^6AB;(?+;[L44&X+?ZF]UT$T_(HHQGG'6!&4D@MR*.^'NYJ=J)C82B;
P5-676FO=L55RX!+)87,'/%$'^'JD*#Y=\+HYE*LYYHCF^1\L>DQZD3'2%+%"P)$B
PWG6,7F_PTK,\@5'&#>)-RF QO*.G<(DRZS0UG#+H=[_]/F (OD6WQI@NM:A[.#(A
PXK06[(!-=_+EEGE:7G*9B6;,63(^+%&4X$LW Q,,S'9^QH6\M)YVA:H64""GW"/P
PY91T_'33DKG&T<WZF0Q\)%1\-/1WH7XZ4YFIV8^=<$LEQ1H5-84M(1OM]SZ0#?0M
PE,M$TI" >^[D,]>COG?2N5C;UNW4H.X&P@.CTPB .!(T[W-D#L"66@JA:*?]!R]T
P4;>F(O@W@Q>JDBJ:<3=M =2PF\BX$3IL I[5G1&!Q4Z6]&^<S) V9^X%^2;YT*W#
P>^0K][>N]K08UV4:!,;?5A5 '&);%[TAO]IL(8;X(0[B"QXW(B*?1\5T)GVHDJ%C
PIS^P_5;H268E?"?KX>!K8=0Y.Q 3>0!\@SNTV ,7Y<0&F?)^'Y"<E/EJIT*_9+6F
P]!-E5Q+S:U^5$J;Y<W4ER+M99CGA%4]2)E,Q@U6[%GLH,KJEB0Y37MC4^0ASIM[/
PV&;MW3+.%'765-*%W @ZLK@'(X-02U4R<7!UB&'U!FS7K!MU;7=IJ5:;:- 6K(?C
P*"._KXC"]_Z81SGY-_GVA?(A;.1]QTV(!3]4]M7X8SF<E,%M+9SY/(I)U^&9'#H;
P>N@8ILR!YL&JJEXWNXIBH@=S)Q+L%*MA_JFFJ"=$)XVP7(-O/E^N:/'U&/T:( FM
PV^COD($Z$*R-24WDG*U^<>Y0W<;B>L;1A$<D^^+&>%YA6D"38%Y+4PT1K"Z(0/TI
PH?#M]MB'H[(.'(I+B$<UF]0U29AA\P:,:9E *VD%8(W5N16)27HD?V;+0)/_$'7Q
P5I9K@UJ6I\VEB"RVI2(TNE_BKIKIKU@>SRG1I"?25JUTA(L+4.6._D?6H!](,AYK
PD ?O#&S09'[:10[2(4=3$-W:G6UQ7R<R"UIIF=(H$ ^-:!_ZS[?HBHT)R-IN.H#J
P>_D^> E4#'&QH/7.? 2<7?I8P=39%N7"K!K+*J(!@PY]?"C@4D!</F71H0)'YNJ\
P2;'.'JN^\NM=.(%7TU/V8$A$WAWX0X9@@7\&K]/^+U0%Q3:M/LIIAAE&PM-M!%DW
PB?H)F%9ID<Q9!!!3@HQ -/R+%9.D<C5L=[]M/4O5!':SA.__5FT.6Z<#&!,@>WW,
PQ4Z[ALW965,G??2PSO9_S@S\N?>#HELK?XHU@!QS78C&PT'/$F%**T%,+2K85/@:
POS0]%IGF9KCHDX7DLSDW/KDZ(V^9#T&U=X:/FSWG1R\);1O?7>E+NTQB5C9'=36;
P5H]1[0]%J2)M=[_O^2P9GB?4U\8^O,\+];Y-#K-N4#V\;].G-JVL-.H5J!Q@@+IB
P8CC9/F-Z;3#2MZ=RP2Z!RVPY6X]2:&YT7<@,MV?XKAL/QP+\2MW+ V2T"#WGV\O(
PC[8#/PJVLW,L_Y!PS>,4Y"LU]/EPI-3B )-$"+3?D#5NE95AM-G/_Z-Y4Q& ?Z;?
PQ5&=,57*/F&4/.R8O*9R3I8?L@L4,&GQM[AX)!(<9+2."WLN3> >2VT,\FU.[DY9
PL4$,E5<>]S8R>@>W3B-&64XH>(DJ8).VHCN31FES!<&YI4-A[D: _S#^G"#98G4.
P!9+LDAO#5F;OV']A>5U7'-T143P6_T0%'_221M[+KXA3:OG4%.W;57[X)'Y0'Y13
P)=P3ZRWUFBV_^)W)8P[!0K$ D.9EX5.>7Q=))T-;V=[/(58UPI*9 DV_LVAAB=^-
P,UL.S@N>NJGOCS *K%&L^:)WA;RZ,9M:K1=U?N&WJ[,(1LJG8GA8;O/0%$0.W]WY
P22Q?.*-$)3#XPX8&F"OJ3JDJZC)=Q)\.DTT*^CR)18QWCGUX33+PZ/S@=?#Z=,6[
P"8KW2W^86Z#&:Y2S !-B(0/2/%V5M.>C7E+%C>("H/3=+UQG\B"\8>D2YN%Q:^5D
P?205%PEZ$'*&,(5$0@P<\X/^$7*54GIC#RO2X4!J$9J3BMR2M)!12BGS/$!,/V20
P6SL>&4*&X@BE,=#)W _[BX*.=<.@+X,S-)K CMM3JV@;';:?)X>XZ2H:OKJ+X_[6
PE%_A6UH%]RP5K:\P*WG+9@OM,/FL-/Y+.6YOHB)F X6^D/$E2F#XL3UZ-;HBV74^
P!]T4W9I0]K@]Z'D)U/*87_-ZS03J"/4BGP(1@3]_^R1=\JHY4U1;)Q5U?)YG@F@Q
PHT(61HZS@;AO+,".+:M(;+>Y4B8?(4!5_I.P)/+=^//8T%L\&,P88_,A.-!F1>LT
PI",?_MMHRA_U8<]#S4T%1.RX3(4ZRR*#-I2%7(ZVL3G"01OV>T+IJLTT.LQ)05E<
PM. ENI/B41@-[,Q?S-0_VB_'.UL7,P#H2VK[O2R!CQH7Y!@>UHK2KX6$8L+B.!?Q
P1"<SO%;(YHN!^-_#M,ASCE9&R61CX86/+)8/;A''.#X32ZY&/ZP?BI"L%D+$'!WF
P9Y09)7NO"_T_+;%_?&+4AQ4N_19/?CN#FN.7W(K_.=7#8)MYAEIW&JE\B<)HQ N$
P+DANI:@3'RTVZK$PU[.Y&_PR$L'_R)ZK"T&,,=M(H!5JN:*>D TOG=JIU+2NI[KN
P\OZFBZ3;+":8G9=T#VQ$G#IJ.-K;>"LYK$UT(0A1V+C;(L 78W>]/\I2N'NN,)OA
P:2?(/"\6!X;,RU;RN0@8>B#IH@3!E^VLV#C6,7%D.+P3[H(!',_E;5/TXC-/NXEC
P;&F;6.(.LO,.\$GBTZZ\60J*1"I#CC?747>"H1!%-)_V".1;A.EK.^I8-ED_]Y^!
PF&MY#EA \5M3ISZS:$VV 6@*J0OG\X]G<QNK3=J)=6F5_,CTAEZ4 0Q,V:#%3Q(:
P?;L]W"Y$7",VO7[I8='X8LO-UB6TN(Y,#H22O.]V\S"$ML]'-I<4K)RVPU(O3+*2
P3^+*I <Y@277I8G(V\! >TQH-EP-Y+,PQ_/P2A L,)6V.J2):V,&2EH(1QUOFR 2
P (M: RD^-AGRO!8#]NO_U#T0N>F@KQ<@02YVQ86=3$*]%"$3/,[]Z>98GE9L17I:
PT VP\WQFS(S;.^ZK08?"H38808[C1;DE=A6.^1B!6R?3C:= [!920G!\\,F."_(Z
PXB20GY4XD(I)1G;8,Q1<L 2,XLU5</4#?>Z?U>-RW86MIHHI29QW7_PJIJXZABN2
PVRP-7:2=.TRYI S%(O$-->H\/8?HZM;M3F<ZCR*Q,>3>Q*QDTKOOD2B"PT'X/^.M
P4NZHP[MDY'Z8(^2H#H);OF=_Y.4/I4;*C-17W[M*] ,*# 39YB0J'AAL;N6T._01
PZ$J- ;JK>X9314[&,:M"!O/K?JU+?;S[9&.G\_WOPI55!O3"\E="91"G_@S(S1ES
P:9EW]0$ $=*TC/;" Y"D]FZZE&/>"GS=1H.<N9B5Y0J ZB:8E>W)L6^S.?EEV4FM
P?5>AXVB?>Y]U9^B"63]4[;2L93"ZQ170W&<6YL =]K-O@V?SAECAI6TH5"=?EYD6
P;!*-_W0YW]6JRO2/8L-%VDR2Q!VVNK,&P9#6,F55V;S>$UIAP/3'DIF^-TZ#6P-E
P6$ ;FAY-'/135(::N-JTB)9,?-K)-84]!)\FX+E$ZY2;?>>%J"F9XW&4?;D(FUI?
PO(K2X5]9_6_14)#!H9-G0B%=E^W03T:(.R3B:09?<QTI+U!LZ%$PO4%/K!MS@KT-
P+>U=2/^U;.(F3 8X%7_?L>4[VE"KO=LC;IU716$G1O/G)JRLO0V3CHGVBB7A5V/]
PSQ#*@K>$9XR_S4O%LRDRCIS.#>(2YKU9W9T^>Q"C+TE//^%I!1.*W%_9KKQD-?9B
P&0N%B7]%-,6/RZIN20N5BIZF<$M ZZ_E&E"5^"+ ZXGZ&TS1^PVY.UX2X5W301GA
P<"^=DZVDH7B?/#CS>=&)RA(]*%HE:X7H^NL@H1O'K. _2 B=9O=3QQ^ U43Q;(Y"
P<1:']A>Z>GDN!"-K#]=$1%':&_LOE\/9N@7%D]1"!8YP<Z=<XY^RM_7TTI8'#L@K
P%[)<F&1)C!Z(<%EX10$?]3X#'D)4\&9,B)AF2Z!N1KQQFC'I:9]V3KK RH:K!.[3
P\!J*3 SE< M(:D_O >*UQK190RG8?]\,-,7N5!!KXQ5_O?G]SL<TR/>N55V%/>L"
PH22&,_<Q3.=?)S'1Q*)[FX_'3D]V**6'8]/]"V6A'N.3;DK%^7-B+$3Z*?,ZTOE,
PL,;[YN&Z+MLVU(K+^8F@UH \S$X;F^VCN^@XB@356TS"LZ;,(E6+;A^VIN'C&F?V
P=W>2J+K++13J8^'S>K<43#+!#)IUN7.2NMW T,IHH"! A?!%GA>OYC=LJ/;YCCS$
PQB5<U;YB5@8.S[_[,JR+[ >06B)=")L^'>=^W)P-X%]U6KUV8R3!I&FSPZ@A#8WT
PMN6_-9%90#UPS0:AI"HSPOJ=<*D1.+<V;T!^$766J2,&1RH5M[V:8R3R[Y6935G?
PLK$K\U75<_!28FMS:A;+.RF;:%2.XBHNW@D,CYYTVWOWF1?_-&ZT BO-O.'5ZM-W
P_N8<QT6)64L'4C/K)!AN1+9_$V57O G+G\"0N5II8T?\5I$8@$N[0 U3!A3,#,1:
P3[R88Q%\ B,>8Y-V]DJ>7@0K8N.1B# ^/^864QWQH^@EJH=4M0"2B([J5B ?]%U^
P%0^+J".[5\^Z=(]7V-?;$3S_FZ7^:!8[OPJ0Z*<1E6-GI'Z0IK%#K /2":5%%W>W
PH&@IEP+,OR78YZ)7!;LQ,;'X9.\UZ'S8J=."'VH$N&AO^1/L0_,8\)@&9Q^U$Y;P
PK+/8PT-"!N1HON@0XXW_@W,L,6M]Q(*.;>_<8($!L=.E"D@@L*D2E65/88G#("01
PV?5$EOU++OEL^!M_)TW**FW_Z!<W7W@UQ_G,C#91/?\5:WX+-M.!.BU].<5;)D*A
P:O*3E<,$X8V7)QHEX^+*)HO&-$HP= .7<93@U5ZUS]]^V%U?(+)XDI:8B7_"@-VT
P+I[I3UR5<UF-4"THDHP1:DPF3#0PA13\[!?P#JJ1,,\)%64=24G:X=,ZG9K(V%)_
P"OR]58WI_%L\!5A#)%3C'3-W ?=@H158J&N^7'*_C^QQB?#K..K)+T+!OV:VM&SV
P)P<H!+:W<L87E<RS]67(>]4[9TOSN-=*@C]M,/!RV_8;;D]<T\P5_^Q3J^XUJ^F,
PCVG::W81_/0[/O$K#.$<IS95R_D >ZUC4.AD;ARF<&$8[\'G=OGCO\P9^J\AT=V@
PQ6T]H$[O#Y:LNB,-62'N^C'D?(V[V;]ET%@XS[*71@\)6VSO,6V@)OL> .'>HV4<
P)RG)-6[[!=6* N.:9?!!^*]=B<.K>R.H9@M&0!%K HJB, 5/=9Z+AW'KGHCH[:.3
P'=Q.2E_BI&3G/]EI8MQ[&RF_.O=6T\V@))(Q3UZED.:>]0@ _P#TI?*4/09&S"<D
PWF[ <G;[6P:!K22D]O<BT;Z;<3K \KQVU. [O2S(-7L'M]V4DS:>+B&+B>ASCGZS
PX-]U0*]B>WU2:\^VEX>IYQ58D$C3(NV#77F1X6_M\[E^?\7>2,5)KI<:*:T*; T6
P'3!%'+9O]O]W\3=AHA:KUBA3SG;-+ZSFL0Z&9BE#:/)56%_J<K]1_R_%2Z3J5>.*
PW']P!?I0B)9<ZX@O#U&Z'$'_H9<4# 0R;%ET?9TN0)IOQ"L$,(E+V'K[H"X<<W^6
PC[H0[D3PG4EDZ9FWI1/RF10-QB]Q;96H9OQG7&^$37OF\#.M%.&H1!B^F3^&Q?H(
PIP,KIWP/H::AT8D5,GB^F.XN4^SXA5Q4G,SE5]YHS; <HM_DSPU:'2Z95C4U6!3;
P]$ZU%TDI\R#-F4KUX3?B0?1BFTXM!YSB0U0?^;/9*64F0C9G/\U'O?^9F_O#QQ<J
P:T$R]CU_VLTNP&;0OJ>#,*]%/;B>K!5^C@DJM,ES5N#IFK=E=#RVV[W9PD!<C4OS
P^[5CWM=*;(QF!6@<4I;&'765FT)=B3C,-F%]R>3G%N. CQZ'''DEM1Z2UH"&/+MP
PC#L1[Y[&+.]5I_XSG))J R1_+"+@]0K%!]%M:9,J4 2MRV'@B\:BC8DYX)Q/BC+^
PI-@.<U"!_@MKGI&@.(BDWIEVH@[J73\.:@!AG3F&$/FIC6O"/&7O.><BOQLWF _\
PQ&$Q[JF3 "V0+'<ZDR0\JY$V[V<V/1,O6H&KEF:AA=Z'S2_Z;J&B$\%M(O=#P@6"
PZJ7SN.37HSQG%H\?Y,51CH(IQ+%NX2B'?X?U=?WDDY]TMN P-3JX:H3G6*9S[OG2
P%2V6@2QK#0^9>N\5YD_I57: ;MFD^H2K0D99 $N,.J2DY!\R1UP+@!2,]9L";]SU
PR2(QMVZ!C: \!U#D>R.)O$<!*S<1%_! MHA7]OF@J$$\P<&V&G2NT)]7<B;W&Z7@
P_U_^:G F?J22;4^95+<98%QR9ORGO236?H3_%MGA&-];T,3B_Z_Q[R)+O73T,3)[
PR))P[G" D2Y7M=J2;O8T@[,>M"*O_5,(6GT*E^W\]5)P22G[PLB3*2!S%T3QCE!U
PH2(J3@R91-!JF 9 RM'WCN450.[IA5'G'S'\DES-.Y,Z^M;6!4^IBK24,4[Y357[
P?@QE4",6L@R P3B7Q_YH=T.ODLU\>Q_MR*Y5@TJQ0)O=%QG^]!%E70Z> 'I??IH6
P)LF3UD4S.H)=WDJEQ.H).>5/U=ZA6X&U+2J5/#E8U)@D,RS@,(E(J]PE8'_$NVH6
P=>D">,=,Q<%I!%=7:GI)A1:V4=+KU_NT]#A(<XI@S-D]7_$>Q"$D-(ZN6_L[:WLK
P03/5P)8@FY2DK&<&NXQU4B(*X[E['37DU&2,-V+GGQ3W_R$#92RL8XU$%XC6G-PQ
P#5,IH9W)HRV9Z=F?L5(W//M>IRAK3 =0YK7E!6,$1ED&*RU)3@6YT_.U-]SE8)+E
P&>)#5Q7U^H: W6&O)48%6%B<D4]L5QG./_R'*>3HZ26GOV^('UD%T9S =,K@=":;
P'?X*\M]E!BJN('-7M(X#UGO(-W^2X;WYJ#D6@L4=[:&=1.YPW>$)OX^.*>4F)UK/
P*^U/PC[(:(.E?:0#BC8-[#GS8\COIJW?'W\1]'-F 2?]Y9=Q,5UMJ 3EM)Y4Q:S'
P?Y!2O+*57N01SM8$6_SY(,-LB0(>5%5I+I-5Y_PK*^I7-G.$OR TX1Y3K44,Q89_
P<P,(9#U8F:![_ M1OJ93)&_#3V>]"['C4;];@##A&6/[DS+;H50K7&X'B"S>5%9>
PFLJY%C>I?4PT[RJ&+VS/\$)M]1+#4VN9XS3E(V 2;6F@@$E3.5H*GKUPLS0,_M6%
P QK21&ID"% /-4<*W[>3#P.PI:P8GVXTX,_2K-Y<DD)AUW,"U).D(S$D&FY/98()
P&OU,G"AD6*,'D/*S[@H*7&DPF6+:W%#X$>:X_%^T+(N"=!#+IJ(2\;-"V7#EH,HF
P]IG.$J(80!>PD1XV+>[D[HB!3Q05<SEX1KDI^%0_QG7]96EYY)<"$D!>J+Q5>5YD
PX?IY 5C< C,P,+/=I&G&UV*EPXFA:-$> -2F,3:>PS_M"%9?.R/S >4!!\%O*T)&
P3P7*&1<S3@B2K71_63B*>1M2R@9<>NMIDGN"AAHXZ'XL<LF4="/GO^C=^-@8T8V 
PI=/R>3+H;<</O?K:AEH U^'@8<D%?S6,:TN.@B:D9@H*"DYU2ZG+<"!?R6[P[_UN
P9%B+0?O=]@RU:YZ;Y^L.Z>%<AXT2&_M^_+M2*Z^!1;1-T<ZD/31XI@BD(G.<LWK7
PMW%@]%^H]U->$_+CRXG>6E>$@6@Y1$N^/,1]%OO2/.;+53&MN.>W73*][U,?8@J9
P]I;4D=+\^O XVG?N_NT#31?X[X1PTY2,1ICJ+^7.>$F J-2'IL%XZUO\=XX%JV9P
P-C9IR+,;,6,RAFW];QGR'^)G+<4UG[W;]I])*RQ/G!):3H4RDT'HC>77:" 5:K48
PAUG4>2TK>%G@?*GN)L^&"HQ_CF3XW^SB"?TN#)::NFJR!#0A<)W)=A!X'W7'6&_O
P+F_2S2%?/AQ=&Q6B4RX9I('.$9O*7__#UI!8DW6&3:50#"J8'AB_(MDV'0H6*='H
P.%>[08S0MK;56N!NT!%%,T;:4[0"&:<\_;1IC1A!.;S+[S2GCKX+]9H*V4;W$  R
PTD"=B*[&6,,-*YP!G-(_O=;T9&>_(^U]";%<ADQT.9.\:L41)=%'K7- 9SM#DH+?
PCWX+8!8E!WDB<*3<^*[;(I[L1WI:@2,_> QG;;48O:F2;08(7F/BXB[Q.[4>P89B
PE,=_B-X.89/^2H3B>CGM1!O9^2C6N[V-T3I@4<LX;J@\0C^TNPII4V3'/W@L.,TL
P,9/_&F;1G.ZD[X.17GQT"TYYKC'VET&I'DQZ[1X3-<T]#D -(-?H9+"+Q6#R$/G\
PKKX1HS./L(OU=&ADQ/ GSQX;J$"O#U+A3X6,_'Q0N'Z*EVH2^<O,4H2_C5:B;<\)
P"1VD,D[/.F/V">, !X1IY#W_$8%*7Y9=XL\OU1O\O<3-?^$VJ>"<0H5V#!1T$6YE
P*!-+<>] ^-SK>3 U+D8:$'[7H:E%+V6'!J,<>?3UG73J9W; "KZN-7?F$], ^K7,
PXD 8HSU;@X%.HICU.5 *.][=M!_<WK=V?V)+=\C>VKX?OTHH]7PW>N&"2PBB*"#"
P97PD.MBBB(YW00(#Z73YYD_VSOP?E5!<"N[=T!71PM;(*XMCP:R.[2F?QY0.H-J^
P4EP8]M3IUG236LJM3"4NFDD179PI+V-(.K L& /=8VLQXJP\B\>-_SZFE%U49D-7
P-P]'APR"(DB^D-!9V5QL=<B'#A;@9-]IEMPRZQU.J":=FP4=49?UTWAJ']I>5(GF
P_L"78?'X!O\)X35.Y=VDT5KRT,.\5C#BP98B;T+7 -RLST)$!Q_7C$H/*F?5V+]=
P3(+*!%GM7:;%\)F=B5SY&J:#^&.S=RLA@%Z7P*N%@ENG?6^MAH@9(_\?G;RZ0NU0
PH],@78 JX0W &Q$SJ"5H,N,1-%M3MF\,#6%AW07=T8*.[U,'>B8+;F0_J:"T]U(T
P2J5<E2'+<F,8)(,<TH"08;8:6Q\ZTA:_0+;@CM6^),DA$,9&ZV6X?$[L@Z:4M\W7
PRQZGQX)!)3I3=+A+ICUP3;S <MF_(D[^$F7RMA*E 5@E(T4C>6<<<E#4Z\XH99D9
P?@R[DA_4\?;YZM]85[M=$CY^VL-9;@)V*>5Z-RS4%C)'06R^:%T?&;R=L#L?&)^Q
P=> P*W_3YT<8V>14=NK:9S:MS7)6B"!SW*L*-+@4WQ_%'HJJGI@H"U8KH3 UR,U.
PN4:+78RM@'R^#*MX_6KK-_F"2BJ/$?JCK&(M4\[DA1CUW(*9/$DJ'^^!=7T^"0;T
PG@%\Q^80S%!5)\!CP87+!"%RU@@WTAWW$V4W>NCV$[U.M9F0-0W20P^E1FRGI66O
PTI VY_9 ]$3A!W9&]SU%R+R\)#Z@[.*.K'.B66_C3J<ZRS)XVZG@)K^91D^*Z*0+
PJVKN.7/@2HS,(.M)QN8*W/1D/HMGJ^1(M7DSN57DV\ 9]^]ML]X%DT=O&OQ,5I]_
PR0F<WRNK#8C(UTOI]Q&K:,IM8?9$Q1 ,0M>)!>U1&XT@*GSZ9M>&]ZM*US?%=F \
PTGCU]_P]4,!:"-&Q:780 ]Y+%33))MP<)8K5OA0F13^$W>%&<W9 O1BL:S@R\P\E
PPY4.XW/.(3]DP939KH@KK1G8&3%8G7F*O1"P$GG5 ^@T8=0I3T,[F9E9^QTI K^1
P]7N%AIQ/IV+417MT@UU^+;XA'Q253.E!J?.49O\]Z.E=H"K;Y[^'>J*RJ>U_8)*U
PPW7/M* 409\;)$!T8A4TBU.Y&K>(@-JK<6HX '!57L(A2P#]8;4,)76-3.18D[@%
P.N&Y^\KC'6,TYW:O#"%NM_JNM09+XA%QK?'*)@F*[XI%? &.%(R+"@/T ((2R^B=
PE[+5T\2V5HWH[L+^QNQD.&+$GZCV*3U4+0O"?&:MY+B#3"'3*G[14+K[Y-_BOH?N
P3RZGOJH2][1?JLX$Z(E60Y^2+8MIL]S8%RPWXNS7=TY$%S<E6H>>NW?.8S&GT#F 
P@&:ITJ[N#0J;VN76!I2]P!)QPZFSVZ/R<2K!X7"M?100(PW[7L%(S& MKB](@DO.
PHL<[2=]E7\ONDC^,07GN0Y8?Y4?.M$1S ,S 5AA_*/M('VW$MI>J Y=?TK[N14IG
P(8Y  @QDDB+A=E0)6>7-V0M@2^H6NH=U4UR!W)H[8W[A]K97RB&7[_+?\+7)&77E
PH$-Y$TBC*F3/(A.@IBQP" <11O@ZFPR@X2&(5/[G#J/#Q9,D_'G!TWADI8BL33$N
P,W G[8(]/_-QZ&SR>VKWFZ:<C7C.0R/;FWA=EGW#ZK=:H/[Y@NS8_RXY:2M?GGQO
POA*KO<QW+P 9*<>P;IQJXZC J,AN_ZE#$767U,#IV85OH"$_FMELG 'N5:1H8Q2W
P8XU9Z$_^T]].B][Q%@+=9/E:UNS&$J]PW?)[;Q+Q?O8YV$[U%M6WWR\KKQI/+L5P
P[0*?ZK:+>[_D,,MT>- 1];&]C$QSEVW>3)BMPY;D=Z5>9^CK0-5?6[_F]4PL<T\V
PRMNF@GX.FGJ\L-2]$&2L5+6'6G;'Q<VN0,B<SRKIM #RVF)'WT@RJ[/*K[T'RKY)
P+_%<19QBZG&C2!D#).$!7W=\?1\ZZ!RT!)V_.3Q,4@\O_.G!_"2 PC2B9*A4(5N>
P'&MO?/'C?4&B(CAC-?/O(UG!^?-4P2DKV7E=E?IB>"9KRO2A=S8AVPC.URA6MKN!
P_LN<4].0.2WSN3@4*^T;>7RE+K R0O39*'P1F/;&;QA236@Q>H?0%S_Q;[G?/TJ9
PK&\^@>4D_E>O#(C2Q1=\2]=J2XU"*-_\S0*<]FGT+GMW:32\9RF!/[@N8.#M!%+'
PGWQ)X/U +RP?)2^W3;5NX^:Q;SLB''8(.<7R#W-IM\2S0&4"C.6F.-NH_[?H7E 5
PR1?HTK/XW^Y\76',R720#[^<XTB0>C&\5F)P)E9EO88IX$=!M%\_@]6M@2I*H=,,
P 1CH&<J( S=5WK3]U%&\ZTA$D;(T\D3927WJ>_E?%+:",(49/[)\XR\2#C<%B69,
PP^^LX5+?G2%\L/X-P?PSXP\MY>GKEQB???5Q.0OB>"AY[6F?;R^T8UTN&F.^6K2=
P$UNJ'<E/S8CDO<WT'P*$CWX5_RZH)CRML/3@);(WK6 $" DXDE4Y2\S>Z_NG5TU+
PK7V*]/T-N*Y<IDA?C0%>5!C56]#6LO*$PIGT<@5Z'RER+_J#2=]-#M8ML<":<Y:/
PM+3?(UNU&[\G9JBU3!WKUXI]FTG>?0X/G"]'ISN8L#E[-WX/AT[!977P'XR_V>)#
PM.B@Q!([%$>FL>'B=&!R7R=O)D6M1UP!G,A^*ZTP?POZ:5?F;@S4B8G%#_X9 ND\
PFC.,5VQ+$0X0=G5PJC@4374;@?O6+?!8N*[Y([T[R,Z7:C7IK4(F7U4SD?L.7$%0
P 1FPW\9IL7?EB7T/#=W0>'20)_C?7(1F(V&^+US(*N\S 0T?W5D[ZG"/>,D\=#HN
P ,I:'L':4BL4NXTQ0<<&!<\.JZO(K^0/Z5:0J/<_"_TH'V'_KM\E)RYFPK4%0ZM]
PYLG27.!BKDM6Y0>&#+W@,\## L'48./*F^):RMRB$@<PUD.E^E1IYTG29 B?"62/
P,\<(PJ'"V9>;2D_MZ;BQPQ=Y[+>[B.SY!E26^[_U>JA=WKUR?;B?3E*'T%*N,G+?
P'/T:YC&QL-3E]09H<UIY<E(XS,F$".(B]&(RCC%7+\Y%E\H8^]%O"].H6)P7: P]
PX9)OLM E-+[FA T @T*3+"70Q6?\3H=Q[IO.%G2-M\(F^5F-X$YS4U.0-.3P^G_!
P.)YGH%?NXP600/G'F>,OIOHR@^_ R/^YG%G36,H@2MT2>X':+-!#BY2(TW&&\[5M
PGM^C>"!>Y$F\C=SL'5[S-WRW<JLN]?:8"-\U&'E-KN [<DY3#MTQ-#\)[4L@6^4/
P 1GHB$%QS'C]*S2M*U:-I)UQJPH=D+E'G9/=F%$P6B!*LP P\YXSN^49.?._(2F?
PG48J;DQ!.6VNI,Q8_ 0L1HD&5[*Z"O'/'0^N*'<QB'PA967VDO7V"-F[7K!*XY9]
PE';1A=M/R=[P7+UQE2*>6;&G;[> ^]J>@<*\^U) (6V[O^J_1-<C:@@L01J;4P;7
PG@@W2J\"N:_A?617FDF/[KE634P4ON##WG*@3/I3A;: _921K&5I2^ =G>!1:%]F
P$:*[II;,_2K2+W3JT'U'8I(9::7W >79ZV/[WFJ?*Y_Z8$L$[K:R=OQOM2]*:$8J
P2;;:M2.F@,+"TF+16BGX;HZ<%\0?0SZ6='?X =L;)=:[+YIZGY)"-&]>X! NFY>%
P@*K""6:?5YC+Y _\RJ8X!9&$7.Q2*2,)M $5PN53AWL(A&L,K8=4.D.*J14!MKL]
PDMB4'U%;\;&(OCV&^,6/K5X(0(:Q!HTQ)X5X(1J'";S8D(:\]VA;7RI)0YJ3BXD@
P@G-O1NTW?_P6,]&K4OR([*O4&<?XN"+MAZR%5S^T4Y/)_'-;\ZQ*'.3;)6L:TV\5
P4W2_:7EM?!15,'MO0/VLG)=B1+2FOXG2FIU0\9VL4E1>2%!L"<&W/8!;*C\H!>FC
P-6+0V)*;$B'G_0JFR>$4PC%;^+54J>5Z34BC^SR< VL?"NO,0>>4',_EG%P=B&]F
PQ7S0>MMH(M:#Z,LO-(R6,VO(NN76U'BQ>F%/5 9[Y5&HW#V:"!6Q%(@XO.NAU!T/
PQ.1$,NH/H^!-L7,A? =3!@768$**]R&0H3IZ3O5WO&#W-O021@@Y*ON9YB>8O6B:
PC#@3:/[_/O;3@!/CVC:(<?+8TT!OTM4/[E5_@>,IVKYF[[230N1)JU?T<7S'K112
P:.S=EL-!9S__A<D]??/9W W\<Y$/% ,>S:,-^6HT#<K<*EU?! )\)""[=L,ACQ/$
PV;*;:UZD%D)FIM".#24G!"/VJ+[U#'MT<C!&*92;)5$LGZ1!8FVVAD6\# #7-FW-
PO&N^OSTSH"/BU ;-;H7)],FNZ;6>7_*04JT79R7@Q5C75(<.X*-22Z [47#GX2(Q
PI>_S2P$"^3S*#>&Z5-'TN](=I2K4N2!JHP[TWVB8]P*7E]'S:J'5=Y8JWS_VB28Z
PX?J6L=:F\Z/:ZS8*M1)(.0X*\JP5UY)V1F;NW # SW76.F0(.2O[_2]5_C[M.R(C
P-%O[I\_4E]OS8CBLYZV:V-\C43VJV/J;>T%GFYV_W69*?K1L(R:ZD;1,:../2 LA
PWA;X"]&NGG#0H]O<MDG%TR))?7:4;(]WU?3@@9:/;0.8K<H*Z$7I$$[BBU_(P(;K
POEV<C50:9GA/'%":"\V]7#4]X%=^X,Z6/]P:"SDQQD6X\!6F>#B+6S##R#=2+QM4
P&LG%Y3(>$N#F3OV9 ,T]G>PR[&UXXEF@$/,'G3_*^DO*'N@[Z:<;_)2=_?)Y%7EM
P?%"Y$KD#"D\>@GF\J:<]*(700_H\'=._UXS&PTXYKFH@%FV,59/B:"_ &P:Z(>GJ
PY\7O1%*F4-)9#3]@5\ZQ[]"Y A:S[M?*=:P?6[*P"6+)RZ0"1FDRP7;!)KKYD*UG
PJ7E/_;PN&/\;%D]DQ]"#LU'NB'U>Q#91SS!..\J)>"K"FS9Y;B1<M[1+F$+3R.JQ
PBL=]6)51QI/GYDK=9Y#_F%*S!P)IL-8X'<1ON%DE!B^IF,X])DP; >V-X*F]WP54
PN"PH44")C5+U,\)#G/+?CA"LA0_OXN+PVL<B:IA'(SQ5%X$==4U>F/:)D4S&Q_7;
PZ6:-SFX44 (O>)7ANR4"AC3WZ,34Q$G:OG)N@@Q899(A7O5&-B1BJR&)J/R&I"\K
P;1"ZU97.MAQ"BV9C!#S(89)Q_XDY4C8#&K3AL?4LD=]$3:6$=#TQU$?8^#VGP<)G
P>Y@")3.@RV)\%6P9=']9/%A KW/#%::>G#%3:EOBUD<P"MB(=5I?*OV!E+X+_9LV
PXA-#%F'T =%U7^170!P3B._Z+$NCI6T@!:8V_VA](E!CK05BEK_LY)7>;),[J*S/
P L$$, .=343VTMF"2.CH93M0_S@1<6NT69#'F?Q ,<MH,\#E-&"B)$D$YS@Y>9W-
P0;R@*@&+G5+="C2T0^WK-&49>.44K&R8CXAL0R8*#FLO=]V>#KTVWB@:(D6EJ4N"
P$VSAH*166>"@LF.M'[Y\@J1]^]L.XEG<TRQ@WAU"3+_C-$^'H">3I![Y&4$*;6%K
PVE@[7=N(JM19WU/S%!A+[);4AJL/CB78*MB!?*V11Q2V ER8UN]_I84B=^YL<8 3
P2W_%[S2OJ&%%J(W^J,C=N>=M+I[:EDR$9P>7,V%:>O5C.M]@Z7> :1/8\"]CF'.R
PQ;&&-V1S"(8SI<O[7/'7L9J@5WY9GO=M/>R&K]8&*GQ9?K#ES_95YL:EEP&2T?5&
PL'QJ47*LK331=P1S(GZ!??M$/\'.)L'JQ$7!G.@:]T)UTH8&T![$S9 W#RS Z(D7
PV)0LU68()3D%\R_#3(^^KC:;(-)_V=:04)2<&&JP5L=ZV,.<?0ZZU!%A@=C]J#_]
P+/VN)4IO<_4@9FX63!9CK9%H8>6CR2?QV/1P_L<T;"#K""34>V0.T&EO1[(^?>T'
PS*E%0S!5D0TP"RB= Y/+,J>9M;<;!R?<T_Y00:F": WVBGS^CW9W1?7$KI=HA@(\
PENX";L:-^6 OXB\80BB+GI&R))"I>B5&0"CD3N<372'# 83T^K0<V&CC.>QS8K:6
PO!5#\8.:.6W<FB*33( ^@._?70$32GRVI56OA#:@WY?P1A+7X/]/S5FQ95LQ?*)K
P&^HA6M8HVPVG#[QWQ8YT6W;-)[H@YW2*?X^W_(!BLR&A@"(J%FEA$UP=;RX_.V]9
PS@*3,$<^6ZTGM/EX"^1A=)[BU"&(SS*1ERGFH- .QA#W9FNBSM0FTXQC#XA??51V
P##[^7(US:6<?.PB*X><G7BI7LRZII:G75P._&3+0[PH/;B9E$YTG2H_$-R##SK,Q
P>)0Y:JJ1)=Y,X8$B^[B-*Z#*0!1C)Q9.?EW_O2J=KI2*0:>@S+9?+'/L-N/E/C<$
PSRCA-;H!7"PU8W^H\4:5K;U#0)#C=([Y>_\CM3]X=^H5A-*YAVE9*J+%Q"C.K9IG
P;/O&Z=4"-! +CZJ_>ZA%E6CQW85'*EX78J/LBE*QWF=F*9O!&%;2'+MAC[]ZAJU2
P!#H0Y7T7=E15VSM4\R/XL&6+HYK!5HZ_JJIQ7>#%,T\)6*"66?E0(;Z[=TUY@JT:
P.H>)NTZB"K:?F8UPFQ$/9&54W<3'BO%2\#7U;EUHD(M<B(, 1&72]%@J4ZGO;N5O
P2*@@-)%;$KDE+S&I>?0@E;,6?B!#&I> _"1N_@:0BW-6\/$L48RS_0A--"L'I&<(
P2-_;G=XYLDV\W!LMX T)KN7PJ_A.O+B7[?2^:R%B*<5)+EWU_/7\D-T.5 F"NL?=
PT3(^YLPH<]W]F'8C_;_T*%PAB&1-*L;#-8YP,T$G<PG%O8)>L=F=>"HN#0\]UG#:
POQZ_.A*AEADY,SA5,-[E?]MGW5N_55ZWZ#,9LH;E"Q'CS*&SA(L ME<S?C*!<T Z
PK)->!%;NPZ^,,57:GYMC0$\+SHMAG5>\S@[B+C+(NM$93=M)\#CW(1N!W&*XSDZZ
P"Q(X6K/B<)'YKWE#'/815P/8/JXT!.)N S.1QDQ.8-]Y7BB!ZPFI$1\"*F;R9=5/
PPS6,N#,IL*"X/6U=(.&P3"ND.1L(M99A/@&+[%?2<7O,2V8@WF)=\%6)O@E, *-]
P2IP<TH_(;9Z@VR(NQ3P*B7Z$TKJW&4-NFDT^?[- CC<VLKH@#^&1YL6Y$TB;PU/L
PZ<H-C^RT$7Z/'&_;$HW+PGGD.:" $%:6\J"!V;%#(>0ZA;5.CI&C".!3%N\(^).W
P1,/J]!/%B4F]Z0'S799Z28'X]1#\+76= #_1IQM(=="L==78Q/4U;8TR3PP[3SC"
PGIQJ.67I, ([,=H@NO0A!_9F<552"A+KF0:_:^P?=TG6KF9O5)&@D-TXHS+%!'\N
PU&&T5_98%+;7D$.P('=N@VO["<E9)Z6;\0K<^IFA"QZ#(/U3"UDZJ.B;-W;*>.EK
P54L@=&#/:D36,R.$Y!&7/(^7V5NCR@-%7QT8NZ$Z)UH SF]7,8\)\_&7E>O7^,75
P;1DO)C_C_:@- _OQ_@X]!$"4+B5!<*%AS]S$MN)4'[^^W4AX^D/+X=>/!%\X=A-1
P% D'MM\E)9"Q^;[_Y*; )!LU:+.%*X+P0IGM)MJ\Q;I*Z'*BQ./$-<!,$WS-WPHR
PX%333")1AVCT!.WS.U_PQ4'TPT]D8&RZD)6VK,@D%Y@>2$T9 I?^ZDTZS>Z251@:
P&';\MZ8!-#Y,O4<A$V%$_;XV:0P^PK':(1#6=]E%=<@%'>S]D!,2>'1(=O3XL*2C
P=;2>/L^1Q0K[?6SMBZ8-@^<T*_28)1YL9!^G8L0)>,;;F6=5@!TME[>XPFR98N>>
P!W2<X?X5GGA2B.P)0F#=QB[;X@4<3;4U;50RQ1":64R$ 9_I)>.8SJJ^QP3:6U])
P+MEIQS]:NV&,0M,HAQB[S?2LGYT'M8&Y23FGE2 BC![N8.@-3UDVI'>3\50@ZE.L
P4:PGO+$A_2%F'P-!H+%H>-5.7B3KT974B.M'D&)3^I*>SM-"[\I,UX])A'<3+RA5
P'IH89CE$#SSMT4_=0#SLZP'+%++N^)S@A,]]&BK7*L'@?W^"\4!20'4(0ND!%WDF
PHB%D6CW3B(K.Y/@9Y#6"%C]]/\FE7183LH>2'T*P)$!PT*S?DG_F= R-*0D1+P!J
P[:?%UV;$8.],H6,<AFVVGOS;S_IC#(/FH4@3!?W=A P.9N5RFS= Q!Q<IKMOZ)"/
PEB>XJ%2?VV7&:F\U!0S8K"G%F6*V/NQR\])@OT6B):0I/^3$,MJHYM54L(H=XLD+
P,Y4M8R_9,T++I8?;"L2>A',B$D#3>CL@ZVXL>S02H*^PT4&A#=7#Y]1B%HPI&H#Z
P'EMV GVUGTP; I%6F'0ESW,+IV;6"-U:NS.&Q,(1G?];=B+W2%J,A':&P35^:@[U
P]KIGZ6*TE$45S'C@GT@_;QV0,OU3%M2J1<X*UYI_7-E]?@WD_A^Z^2"&8BWX%A":
P^_LJ.M4*E$?PH1,617FW?@1"W?A3F$QW]NU1!2^G1])TX/G5X7F(3O\MWDV>(LD$
P+9RNQ1(3'68OC!NLF<!4-RW;;/?FKL]C]5=<?(>@]79&3<BU] @Y_-L(+6OQ&"/O
P03X#GJ1.>YF]RLCL 4T = ?8[]2QV+*]<,[4J30R(3,RQWL?/H"Z0W2VG.:(&>R=
P&19UHO#V-"U!7LO,S1U&%]L\]E(I8,ET0Y_NYGFDC2"2/?ZY:Q4(B\13R*IW6<S*
P!'*(6$.96;2Z6DG7E,IC-U8Y4[I9+ -/=0##0PW^-L0G+G1U::V<7?Y2P4=[(X&&
P@TD]8OO-C _UP;N:+"*[62K3!"8U52VX%>J9-;5 .6U6QZ\SHZ32J.3L579$4,+G
PSITS:,*@"JQM;F(YN)(WR>X#M)2CQ+%9A3PK[<,Q%X%_@ \"QN2_56[&NA%KD0+5
P%;L0;90,*+]4[7["-G(#(@&Z*CB5T5U6HZ,/Q\EK(]I$CPBQTBW?Y'7;>GX5 P6;
P-LPP^,[FGNLJ1H;,*7NB=05RVYB9P]/%O]1,W72 TN&4Z3FF(77O#:X 3LT4@ GG
PY 4':4\-CYUP&(=FSA*<A1I84- Q>*B^NAA@2NW*P+C&BCP:3:!:4WQW218()._F
P+-6U(SF/TA(7 CR]!3CUN[OY6N;%IW>-ZM?1-_*!V9@*MMYU<:UZ+<<K)#O9^)>R
P\,Z: %E"SFF[TE#*A$_ZH[<@-?HJ-V7N04%^E-W?MJIQ=VDV#I.#G2%ND@M<J"Q9
P_F3TG:$$3*.]&C T0&X91CXR &L*D?O#D0D=HX9D2#\9]-8.R,,:F)G]N*K5G*D.
P"U\UR]]M[Z>!,EUF/@A270^=-7]#8JF),X5X[!FJ62\=])?@M8\E=H2<P\I4,AKC
P<>FHQ@>C/!JN'VL8&0JC:!M]8,#+-L[+(4]^0UNMT> [LG%WEZHL[>*@%.@AO9+4
P)5N(CB1V[6TA9AOJN0)E:=#62OZ69^T\679G=J-^LKX<N"T1#N73ZJMTWF;CW7H7
P>'F(J*5'GQZ"';C2PHE+234R'2I^N1K/2G35%Q[G,!;C/L&>4Q$(K*M2SPB]:?%'
P[MG3*3'XPB  /#!)*U,\M9B98/"_L3X!J1/HR^N/8XSARSWX[)R_*M[[[O8GGL#0
P.I;FR^/C[3"= ^@3@UI9ODVM4&T ]@.UXJ)_'&)T730#F2V.?NX(1$TJ=@@I2>-E
PP_Y;ND0N8::P_:8(@D R9G_W0W5/Z*&%J*<&PCCP/UQ:D'\XISE%/\*45(E!V?',
PC+U?#!"* O=AYRUM>]^@TVHL6^V#)C55Q*%^(U3*Z5@1U_6K3%Q6K$M)<@N*SP*_
PLL^BIG.I>>A.O["=0] =IJZ3&.&.5(J/_-$4^&(09.8E("Y"&!W-RQDHGT]%N<RF
PBGPDE'7#IT<:\PT'U.%"I^NF0WO=8<%S]D,*9?]6,NM>I,R\B1_I"OK-.=_YHK(B
P_^P0(;%:VB_JN35*6:,BWJ_#\^V)O?@DPLRP80$+Z<""F>?-LD 17GN^27,7-'T'
PQ/^[V0X/AF>QQYD4>T<0A0'/6S@H&,0=*2K))L/X''&_OL_;;"VLM-#T&VS90[!.
PEU;V6](O@*GCS/2.;SUH_9]B<^F_IKA,Y6SO[Z)KVZ$PWXEG1 VZRVRYK&%!CG&^
P2/O1MEL+/;<+#!&>(+.\$U,&F<>BR!"D$O[.KZ4D3&9_*CP;5?DR7 U)?WS^E3=>
PKHG(LFUTTJ9KD4J5!JI0XH-N1:N#0@F[ Y&S7JU3K7LH<V%2ZK<;AF9Z$YW#NQ13
PTTQ0M$E' U]&?P]VI=V6/7R=9^>IN\2@+_DOA>CLQSI-"Y*WT_O)6X(]7;.V5O^,
PNM* U"%8T&BTPX:3-%<AI@;P%&("<[$JN!<)FB)4\TLE[ 63,Q]"*&LN/HRV/ ":
PT5OO$MC=G;LJ2@PE-%1?] UN1>$;^0A@I51?H=-W"I2JX.  4CX11_O%!NM8JER"
P>DTVJD/EN4OZA!C=3LB[;?H:,0KS^AQ[U7,+&3O>%.7FD1P=4<'S\:R=FV:JYXH_
P^GO"W8F-R!UK#D7FJR\1742^)OP'0Q#K"_ 7G>10AV:[%&GX&3BOLT9;<F1P^ -#
PD,?C+3+X,0+?G"Q-]7AYYT8NOQ3+5;T%NTSUOA/#7U%GG*%(J%DB$$YOHH=CKIYJ
PH2C+,W<Y%^2EI,(I#P7ZSQPR2FOND56Q<:I@L>9/ALS,2@[CZ.2)%CW),T7F*QMT
PVO(FQ"[EKF+IMHLE)X_S%T)&'*<)D?B'9\JTI>^90CA2B]T::NW8.J9[U1.P6JK@
P#W$U=0-3T+8RR*'^)^>?!]3+O1H#F0E.BG<2J)DT=[F4TLH?KVT6N&MT0XO@+D*$
PDY3L#2"I;#F<3!0"B?5BD!G,+-BN"#Y3%P44F/_(>CW*^*"-:]<'J Z!!S@"H7=?
PQ%=_-C9]-DC*S=JA;<_[4<$5D4=)ZRYCF<80.5#NY)J\0'%V+"Z.-RFN,+%OAF!<
P&'1GWXGL6V M).V]+!\0WJ_I42@[QP,[4\JX/%0H2(Z;:(R@9%%VK02K&&81!_@;
P3T^C($LB%0"Y_^^._'M:&-77PAP@]+&:D$ULU%V7-QH=P( N/Y*J6V>DUI>J)<FX
PU@V_CL7\O 7V.T*-Z".RK#G]V<^+2,S "<SCVNK!/UU2*&83=0R[+P/(8>:?P9/1
PK*J_O/%<RD T<T&)R4>[V,\8GMNVR)-\%O$IJ./YK&]LYDW1B0.EMBN8]=!&=371
P)^BQP?0Y^JA#-S;N34CH']+@+"4W8S2Y-3\L*KN#^16#H-MR2I+3&>Z%I26)CE\(
P]#H@4EZ<V)\RJL"-2\=7&A6H I.Y=JU-UH_*WJ/]%[_I+Q>(I9XL$\3>[1C7#QI:
P$ *DNANB,)34'QW(UT4[ZG*(Z1VL?<Z$)]8#Z *R\<]I#>#.#GA-+#>A[VJNQ)!*
P8W<P0738^3I^AXPFS>9A6K&O:34#I?%,1ET67XGO0P\GQ@:8XAH7Y\]=2F!&,(:.
P<^.E,3XN**R@VM5OF]_2Q WJ"?X3OGY-$=>WN<[U=[ZQH6C;)"_RY:FG0Y.B:Q3M
P)?A4YF*3YP/0K$G'0:!:>61/TVMH_ !]"E0H^*2B,!H (=H17^?DQTIP61ZES'Z>
PY&J[=)O<(H#YG]6SU15NX9E%9!D%(5P8DO;SL3."#*-G4I1+WT[&)6]SO(6$[!K\
PUW$RH)\F:4 RQAVC=Q>O$VZYX&FORHG6N<QLR;)?Z-QVI]*0ES7AXUU_6K>.\XK[
PD!:"I:T5?1(V@T(G W;_I)H#A(.]_,(_J+;G$^^6Z-$CPO&^)K#NA\?BRM<::SN6
P\^=>KY++?X5^#%#VTQ J91Z_SV08AI@,B_VK?[V/!0ZK.E$+-'^QUJ33B51OSS-)
P=D8P3'3S:5&!I\MN#IE<T58W.*.4/U5O+)Q^#WO,\2<SXY3<P[ ?<GV?F^%>7;R<
PI6,3[X-/#_K_I18^\4>TZ<%?(820G>H3!AOL,^Q;[_N@W"L8==ZQ DYO"XT=KQ_<
P'?=5?V8;S!RQQOHDK(LM+:ICZ0V%OYDMP=US:V@7\8_03:B@63J].9CON3J8!;%&
P,EU)OCEZD\X;3#$2U,7'7,^W4<GP-9)49#0.=(-JG20MO#:--_5PD"2Q^:48T+2G
PX[V"O::6SQME+* #2@SI;8RNO%VOTL#/J=0KE2XU<CS&2?5B,#]N*57FC%@.MV8^
PK;KWX,K*&CZ@-"D6;<2NK8M<O7K):]U:Z'7,8\ IR WH#_Y5;XKG*9@/)4'D*EOD
PM'"JO<,\A-8.80JX>D7/R;[>*%,HYW,?H!2_9YDC2[:EV_=1XX6(P5_( 97H5CCI
P(8@+-2GWI:-2[J=>&Y\=^&Y[#"JM[8U.!J77>RN,WY#\11CT(%QO'T8^R; 10\G&
PJ:*6JD_SZ_0F.E64F+NY*6.3+D@0#AO30SU&*>&,TCI-^J=6A*4B:\&Z#4G(42EG
PH7"QU)(,VTGX83[^ZZ, '4./UW89]A# 18\\,CM81<K%X.WBAXP6>GQ*WGW];_(%
PVNX+,6C8UG2/=>:=DK:0 Z7WC>$-4K_Y+&MQK]2'.9A47C"]E_[(B7X8\6.O.$6U
P3:P&)[=^^+@7]CJO.2(&TQ4]/,#<SB>4QUN4D?*F7^A<WP<"\9L/T_QI*?4/Z5-*
PND&<'KU@/+/WB[/)4%.#C3+DS@*Q)+"X;YVH+/9!DV-OE?!U_\3IW*/BA$DH X@9
P5ZOIWNFTDY-<QAXPB?IMK+I6OMH=E)?H[KMH+N^ T?R[P<-F1QWHY\KI\PDS,)J9
PVKI10BL<DDY*IP)+2-,GU-?A8CJ3 %LREDCQ'#1D*])18J;9I"PW(G-?X"==\=:S
PC5?>\)Q!N#A.CDP#MO1RI0?$J%:,R44>YI$3;QTNC[%&!H_.'+" FSR4G!C<UJ^Y
P.>WNET0@21L*0W^EF+2CK2@)5*VW[="=7I?A5H$)J/O!VQ<:A2>,0-:XSQP4Q>,O
PF=+U%-!K3IMBC?IV</0IO>\1E?)66K^JO3DL*0H0%9&B_+.DMF!5_2VMY4^G7:78
PZ-M:@)@JI-BW\P(NS#(^8/&FG[.NE5'+S%,Z09+D/H+UK=E)M'ZZ3B=#;M35,L:,
P #K_AW96Z3WH&4!VETTX)0RJL!>\/.?5H3I_GQAJ*7]VD[#?2@+!_K1J@"CP')\C
P?H<L,0;@[%BR]KA=5-3HT;^IBO?+W3EQ4P_Y.+BNFH9NA4>R;T@,.ONB#9?JO8J;
PSPC?B2G!J#8%GI2KN22)7RQ6E=H"SL9+S(I!1\8FUIY,!,!,BJ4OO,2^[C:U/"\L
PT"/V$_+L^3E0/L!V<Y/XS 9[B33$CISBYW3:<,^7L(I5)( 1Z(YCQ,/Q$R^M!=81
P;RC$()V*+_=JO<;7K;X1BF6EE^J<$G;>XR/933DY2E/&:FL$30':(C@/R_5X2KF.
P/SJYXMMH1@):X$7$6E*'R)=U%R;3.7P6!R,?&F$,AL==O-;M,^5_UKI;BP#@.Z$,
PJ4(*2=M;J7W0!6B9=0P;E&&]?1:%Q".B'X*<?8:AF4/XI ]9BN5J*>4JO8$WW"1<
PD+%S[2Y*LJ!I7,?Z9B%E;]71T0G.\E/+-;"+EZ;%WA-H?1Q'G&3P(O;Z3=+QBY7/
P DE$\'J@J"%4TP,YG@=3RL3_G56.GFTR%QN*8Y!YO1DF UP3VRACATT^J#5QA$*'
P:.\LV04!J!0.S#XXFILB"F!4_\#F#W;$$J2SP]&/&8XUA(HA6;*KGJ[.YV!!A3<.
PE!'LU%$:$UQ:F)Y5-O23S@R!H/R3@E@8&V#&"Y9)PWOLKVJ\*!5QZ6?Q&T.GDICD
P3]Y4>N\@_;I41-/;ANATHL\&V_<\**^VO"U"<U)>ZN&U=413$49?B3:INO,\\!8)
P(SZ,()"<K6@ 7C-AK4RF:Q)40OYE-76S=8>8=7?<*^1SC(/!M7@2L!JZ$ER722R;
PBLOXW[F@X941&@5^]>3I<TM\F?Q0X\ZD<H_AVJK*S;<]@B1:=#>$ 72H4=@P>QOU
P=-;H1*(AB'8>"<OH8,Q5:;=G=E3<Y;%8/8NJ'7.UW4M S'#Y[Q2SJWHI/::DZ.&Y
PCX%%T0\2&KDD.&J2>HP&=IZA^)F+M_-8V$-VW+9NDHY:T]_7001=9]ZN&>U27(TI
PS Q%0>]JB/IE&2%+ EJL]';*:N3L!U V0PVY;:]KQ;"P)=LGB[+O]%+G+X?4R#P5
PXV;E=&_GI"B&O2H]Y" "3IEN1V2!U, .:&GK?)FC^L1!>AE)U( 5>I( 3&-.-8GJ
P>A1P.T<\(TE4 WAJ)/J&THI:;^4,$\Y0 6@U8&\L=KV//X[KIT.HKJ@OK-M7E$C<
PXER')]3PTUDS"8-\;*[J82U8/D58!S#_>OB?G/(R'Y/]K)IDF*<O,MK[RPM:JRC.
PHKEP2S 6^#/8S+$YOC,JSO07>@"*\%-IEB1B%+,3C9^LJD_M'9\A#7.B\*3M\]<Z
P-7: >NMO\.T)@^?721YVYE"S3JY?7\MN!O%9EB46!,8=96!5I6FA1Z5@S/9L0W?:
PTYC,M<)%RT; 5@4=)B.EBTGRE3%L\SC2]5J+0!56S3:8RV<VJ79T!$9.F^KF%/2\
PS,%B#;.KBE/[:V5:3";FRR]'S<SCQ&>K/D^:0JUB[IU9?^)_G@:R1 -%,L",#^E.
PKFJOEB4P7D%F/" ;.*US2#,. \_^"7WNYN!4;@\B$9'%\T%\CIWDQ &G&IP<^5D,
PJYYG3,A$<KT[>&.V05@B>#LW#0=[+7;UX?ETX,JO4&$!1*QH@5>!".@/#X9-L:75
PT(VO=$PLJ!L9P!T2]+%)V.PSD%?SV$QD;)XQ%8]TXS:LPFON-R'@67;!0&/[+F1<
P'!KM]T+8> ?N;-.F,$]U!OCOLP?-CA576D111(4$#BE)]JNA%1VF,T5?V5+OO%JB
P]]1^6G5(68-V&<46'(SB+<T,#1GV0"6%#10"-?P"1J#JG:.A1XOPN-'7*(0VD=R-
P'40Z>3=3"=;OM\E*?#F8N7L*I ;0.5\ &&'%%B(_"##YWPG2WN^S3>)C9' L;AO=
PP*E4T6Q7D7]FE,E5QG ]O,1<C;];]$I&[Y(O=@2MZFSF\6"NMP_@54P;H_B'SGBF
P@(J@Q*8F%4EAHJ*X8LI]L&XD[9RW7,3 ;MG6BI_%1QU+TL$0=.:KZ6+2#CN>]J]-
P111ZM#+55Y1#?F?)&A*@F,PQI-M:T;.E5'?3)R!]EZGP#2SLK%M!>Z\IL>7A'!36
P1)9T*F>&(8$2R+<D3L-^?53:=,F^Q5^,1YWX4D!G.B9RDX)#1!2N5]1J:3W)=;&,
P-ON2/M/2TBAB#Q<.BK\!V:L0?DR875K;NJ^1"9@N8N1Q,"(4#-6KL[K>0Y_IG*(,
PO;1"(8:^3 /3NS%O';@TI0+'V_P*R >YKZ4?H1T278#3IL\H(:'S/5S5=JH/<P?U
P%[J M)Z@ID['K$5=H(NJ,!KTO_6Z-'7.;2!T6N8'K[]7,$S9"2TKJ/RZ6"V+(_D-
PM3GEQ'OK*]RDY(Y+)M)1M_?KZ6EXZNJU.5U%U2#OU!+FWV,43*J)N&4*5@[7'@3K
P6GQZ")5O"$G_/)>X'[]CJ@R$7NWFG_#R2\_*9/7WC)9DB'NADW*(,T<-I0KQ!U>V
P:(YU[!U=^J2OQZY'^5[&,?V50'EJDO_5 SN*^/_DR437"]DK-NU4V95W9W:0)A =
PMA,_X(0MO5(NA'GE\19JSD-.?%<)<'6/TXHSANPB!W-&'M]CIVD53F/+Z(W\1[_-
P.9)E?S79)3@*J62?^Y^;(T-HT1"KLN<[;N08,#DQ1BC'(N%."L3A'.)LF<%I;^W3
P,Z]D\G>F .(D?H6='PD'HFL9W%XM/I4=F]UG:TD:R\\P:_,2>.H[L)Y*$0H$9+%V
PBI'NDY>?D]-_F?UEYN8F_JD5,-MEV3/U NZ W%BW='SQ!QCT<9QL70#R5Q@PN\&;
P5)!VJ:=^F;@OUY#&FQ_GXCY=MI8\LXQ+7M*ZAU'/MO4RX#T]) @?)8%*,NXUR6XF
P%->9U-9#D^>+']E+>K=)*2>1  X <UXX:Y#S\F#=0W0#6B=75Z4Z<9J,3+(^K95@
PD$G&;C:9DBXA8_"+7=]_19#6^CJE82+PN+67>!>!X;6#:G:WXIT JI*0KD2FFUAU
PQ@5#MMCG:>NJ&,4]&&N SE.NP.V3Z^;KSK=[1#'*/'C=PKZ&/L;(7.(.]KEI-/<S
PQPM0:F5/NVK>JSKEKC/Z!7,9#D&04CISL17IJZVV \Z9QD 5"DKDK^O6%/2- ] S
P/C(KW!>SUP]GZ0SHXK4(()U.D9S-TKG/Q/Q#J"U$N'?U]K+@,DR@6S5R3D]E1P=M
P_)7P []X=VV78E#U'B0BHD7)QNO$BGR?]E.P3?X>H\?1?]F;4V3I<A-3XV5C.XC\
PIH(MS@/)/#0N7%Q <Z4IKC9HA%>N, G\S*6G^A("J43Z8E)*D<(!3MZM2HE3ES^,
PB-5(8!WSX ZZ5'074$)$H0(?.(K"=_HKJ*KDEO]ML*!^L023Z1P'NVH^2,":B?D\
PW-^EV_:56"T/TC#(@;R.?O,;"\XZ##+ &C-\ S-C0S# UJC<K6Z+V1+$DNGW4CN:
PVLFSN@%^5HB6?2WW$KY3O7+BXBO66\__(7^E3  4Y!3< FB0,^)G)H"57FW0 R*[
PO$=^3[V16;WA=&F"3[W=,T"8!!?(@;"UU^*57U2@<IGW3U\:5%TJ?%@.ME%G0F5N
P#Z$D AS-(HKB9 S3_+$)7]GZT$1VOM(JS_'S<S[__ DYSFCZ(Q17*FV4R#UMAN^^
P=!SM)C)RJM>7L9GH0ZTEVSHD%(4R6GS3T9B:08Z15P:S$9^WDAU3A'4\4KM8<+&[
PH(G]RE\P%@I*JOG=X[Q7.O$"\::3IA+0'<,&LPR%H,(,L]\UO)F'&SV]V>/)80\4
P5BD"I,[>;XW5<FOB1N,YSH?GT048L7OQ@4FM'JF5[M7R)A54Y-W-\4U($438%8]<
PXLR/F/QM;AY"7[:<Z9H23S8=ZK_H@0K))UIYD/<S=%"' #]0W7SO%E0O>Q@M& _X
P@G\9%0*\71^@R#4=\C*6M ^<%;D.WN+L[E^WZ-/)0DS]4(C9*"*&MJ<<8:-#. ;7
PQ'&4[O8$.11X%G^734?IPE;$)=M+**;S9%ABZ\[W @/'G1ME9-XZ0$"@,TO[$2]H
PC'E>*!E">S,%E&;X_H.S?'TLO5S9B+:T3DQ_W?@7DM,VMMV 6RS1H5+=MFNGNXJ<
PD9JNE?@=?K'Y[6L:LSD8-C)R$" B(VB$3'6#G\X8ZSVR%FRZ<I2>_8R^33@B'-A7
PX::UP2()&8-?T\*8F2SOR"JTJ:K$N_U8DT!8%8%L.&SD+0"NRJI/K4,7*]E5#2^$
PC4?Z_/F,Z])-#P\_A)9[&=WQ+W9-@]W=3QMEBO9@Y;.4^KWYG"$Z_*UK_/4WVVU/
PVU/^+-IDK?O2BT;.53MBE70,5LR#MU+*<CY\>0!=H-[Y@--A4#$P/8O3QB03]\B,
PMNF.37*].QY:=2L?$#?KFXUW,:'+LOD*HN3&K_GH^S%1+ELC!H!+XIHX4WMV)"YL
PUBG@MG?W[K4C^8U]6W;>]/,4;C.O*,KAXKT"UQ9F\"E[[+?I6_345=1+:XX%E,F[
PBA5;XFP2E0?,EQ&<*:_(VK?"'?(G8;.I8/2&E3A,:DMXFPDEN'^R125"BXLSA S[
P %L 9:EG@VH?LJI">-M#0:8TD7@T':("A^<P\3C)Y9N"J4^.B2/<M>,8FEF7WWJR
P]BS<>WEK/R@W^()Q'X^;,LBG=^9_60'NCC  <K<)HNE=RDL@/'"HJBEOZ^-/6ANR
PGT,:6)_OO\WZ/2F_1RA9]*S(7@C>,R(YH)-NLBH21: :U62:4R:*F-D9I57Z)K@M
P/A\M6$ ')KO+V:^-G/"+;I3SW./;.[I6$5R[&W-[%!Y1562\AP>55;!:#1NXV*_+
P&[$3._U$"6@$E)F9=3"#\OP56*7M4&)[B284R^^QB-WPY1.]"U_N@2!$+0KK U'8
P9B _NUJHB2="N>P)2+^9EJU!)NVZ4GB@!/:2"E/^.6E6'=Q,!^T4EKG4'*+:<,8>
P7BD!QHTP=U7B3$\;\EC C23JKG8['!?3_NCW,K_'P\S,EC-9Q/7FA[ V4YS)NOV_
PO:F]K)DI%MY+)M>V_!05:)#=4?;W+ D$YL%Z:ZBB>;IUQ,@-)^:J+Z ]:TY@E&=Y
P+0;ZD3?T)_,;J %CGZO-R<@L)ME'4D/W2/\+$:!G*Y<KKC@WY2+9L@V<EMC^G-3I
P:9&CKKGO8=TKE;#$8%).J;QO]Y9.0(A$L_[!@-LWS;K<Z33OOFK#4YBU<^^N+),V
P4?2<UH+7.F0.I%"PJRGC'#VA7_#)-U ^_<_<O?B2/8,J8$@-D0/UY9S#Y^7_)=\'
P;#8R52:%TK*HH07\ E&8HVKRA!P</C,T,HT+G1^/Y?8/^\]D#GY(/ B^,0.8BART
PQIZ>OVN3J+F<SF23<0+1>JO^9@GSJNK41@U4$*_>UOXTZ!<'DIZ4\[X%SD/J'0A 
P,T/Q\9O313GE95':GZD<QJC$(@EC6O3.N&SPJ><&1(3"6F*-7H<//,4\ 88RP6-9
P9$N%EKPGL\G19G9HUG>RF,U,:BARB+.'4KX@^?D(>J1)ATB>(R6^F]^Q5U31NN&+
PE[L(ZA:;PGXV$?&7O^%1T+AF?R)W0\ @&T20HB0\ #VO7I>/:$CWH,3;8K]_Z<ID
P<D7XCZJ#Y)KYU61@L3]-_L#K1"E9>0L#D]P?0WIRO@3NXJ$3>RP:98;:YF+WR(ZD
P=: 7,#:0QZ<T6N8^C'L_@'1+7.I.!*14WXL4ZH8(Q0WDKTP,1F8S6N#>(93Y@-3"
PF.N XEL7I G)4I*&2^&0HV<5@T8>PS3,^MR@Y:-DSB>9&E H.E] KK!J-=@P6F$S
PRI0; "X6;6!SB:_9AV)"XU_N@/J!FX>V1YUFACCK=J_5P;?&!WYC"#K7NT"94A!N
PRY%QX#@(3>V=&XV0)GRQS6$/1T(C:_$0")6M)]!BIVM)0NGV.AJ<;\+GQ1 F6,3 
P5XVZ;7Q:[WC_!8!<7L'K(C]>P-+C'RZT4AK C%+00<*@Z45OK1IAL-AMYOQ ,R)@
P[(8!5/DZ#K>\>F\4;\<\^URXP$U5D5LRQ#<J8NP7T-(?EV&]BU29F34UVH\N0XRF
PF@:%*.10W0'C8'@Y3?6[4H88EF!8HMEH$2:D:QO/#/).TZ72I+;VX)Z +Q=N=N2_
PTX>*6<NMM0N!XP_X!#8]!/4OYSB/<OSZ/9>2@K60266:)M*"]\YS.H,1,C&;6GEF
PR+"CIS[MAC<>W]>1&#3K$$?MHWM\&4IS-L[AT$ )\I?M#.]FH>L_^3QX,?D7+X2V
P#'RU%I'W!AQ^:K@:N,3]"D(H.6%M$B2_7L\V3H(9<4Q0?.K8\NY3E>.P7Y0PDIRV
P"E#VC]%XS=I.'MOQ2DY6@DFMMA4S-*TVQ\6+*8:^Y[T7']TLXRU1'D8 LU PO4!!
PK/Q.'$ &RT;CE33:AX ,*Y*)!"(8=*9<WY)8&TPO<4:I>!6(;%@89_4) )Q9\LBX
P&G)8$ZXK/2X-5%F\9+,RM(QE8L1+00/<HU!4UWM^$.E>AQE0 =C.QE>FZ3I&L6-'
P3<W#5H>* >W%>N0GJ?W2I16%2L(F.N_0E,Z$[W^9TZW]=56-8_5[I_D*;@E=/P)G
P2]S5-]: .ZYWF._(<QXUT-%^IBEEF9ZHL[#G4V26H@.S^9OGHSHW&F#'_+PW^HCW
P3*YO<N\<YB"'DNE=,K;*@Q&\V]^7JL9X?\W'.G<*W=SPL\#_OE3S!$=KT:5^CKI#
P Q>2G \&OE(=; XTV,-I>+L6?3@RJKL6/D0A,G=N)5'V)@7\BLDB7CI.34.0.^1B
P41'^CU]S]QDV6P;'"M9^5,P$=M56_J,%.B)DPOUW,&"$Y5TR$I .<PP>=M#U[E1N
PH:\9]W6#8;#0.--JCZ#[I\QV9K:&0TW!YV_K1*R=]I (#?#&P^NT=FZ^/1+"S!,K
P+]WA/[ZDY7IP7-LIDUW4XN/9!\%)7V#&$T#["T24J4T,,#7+ @SNF?8LU&)4UFI-
PQMM">XE+NV!K4*F(7V9(#56@W-0+?G%L%'BOM*)YCV3-2.W1^FEA+:?=OC4R^7!C
P47X.=UX14 _N9KA,Y;UXH:V7@KMM]_/@D%P5S^TS2GX]"_^5&K<>SS#BI2&%)L')
PDZF-)A%FG,Y!LW_(_VE7D)+*;(8"E&.8*,+)(E=9.FXXO.E#'53X?0X R/-RR[0"
P$49U<?.\!F"$_%@V+1U3!V EMQG4;2-?;X[<Q&FF'0,X936[.?QBH5<\\<-JU:N#
PV86P)[,ATC2([97JY$X94@\UXGZ/O.-\)^M$<VZG_M:37L:;L#?L&@Z W$'9;&#B
PP2Y(/V^'7D1)="<#Q:Z$'R9&8.>.7B/T56U=AO_,[B5FVM'/K0#,@Q6]FYJ';FHW
P!4_U0AN*@M5_#A'W[H5LM ;==SJ<_)&""4/ J4M.:H">&&_.:,/3KZQS,K7_ /")
P6,,OO^J>F+-L% B$Z)[VPP[6WESW4NB$-WO,)0>T-N1CO2O2^QQOD.W# +[C5(%(
P/A&#%0(@<=G'@0%F(48B[<MS\]28?/LBS=?\YRH?)4^B=YX[7PD*IO/>[/HH<N[3
PI([,,RW8)09J9CZQ+)&Z(PNI(VO/M"\@V=7KV_8D7S:E4O$1MM"B<]#&'&_L"!8E
PJDTT%VFA:KQ!J8X$GEA^1S547BC9Z^\KD5UG^U>-3]<NA9LYB5U5?@AE:"7PU8&7
P_ILT,8 WBC\GZX*'27K8X^Q9HO(I!+MPA2*.)&\/"L,K6E1D%@]]XL6FW_%V7'E]
P>9$,Q%;OZ>8<0#XX+D\&YN\C=0I:@N1W"B\3BD1GXYW,$5^(G/O4PPN2/4OM>E3V
P$+=;;%+"]O>!)<3+T^7NT0!CDR,@D>: =@Z>PD&R8)[O0R^S_;,IL!DE+;_3L7V_
PSZ7!>FE<E!)0"P1W@@C9KI-K+C,#KC36_UMD)6^MU[C=DD!;0?3S-)@U3M4TI'^,
PV!NS=>),Q]3L]01AY?>LTN)H @78+>Q]OGGPYO[L!))OQHWJ,Y57GP,HSU,6=+K]
P>'+<QB\ \1&_/+E);:_$P^UO"?+R*EF:4B>[,RQR[C$!P3:-C!L/B=B!UK-YO::C
P-,MBI@ %GZ?'\$")"W=(AFAR>1%>H-:7'F&/"TU'0H&K5\[VEC:9<"X8M_  \AWV
PRG?0P$L8DA";& O/P5'MDP"241>R2^3@+U>5#KO:^'4BG\J#$CCEXG=I]B,0#+?;
P@51CE^>,:DUKGX"9RX-I>!B6CTJ#SGSW;+MD_J_0Q/*HBX-N';M<E?0$?:DY(X57
P$C]$QDU^1EM$:9>QU;" 2;81.R&[5.&!V @6MA0E9BIH=[KX0'L6N$JXVEXS@$ZM
P2@#T\];8C,9NUB9R<T)YL4Q&IP4.8%99 SPO/.AE=M?Z-KD0)&A_B8".E+!S'6ZG
P>2,CC0X9:/A$;8WC3D*S(#\)*(''!;8#X[( HJPXH<7JZ!;-T71W,MM@_YLK[5BM
P7PF='7QZ_A'/9\#!S+QVHN&<XG3'=<SQORE=NEVYW_ ]M:/_E0D)(FB&;3P)3LX2
P#R^M6@ASX(#L&).#&#TFB5LZD1E>$JE510W:C:CT95PRGL[%167 !3T- $/J\5W$
PM5,R_A /ABA,9IU_  7@$%>;*.!$#7DJ>SB4:ZN=#5 #O10O*]QQ\/J0GH'6'O1=
P#PR [XK*Y<2+MRWP0F$7?AI?ZXN"[VCIXQ^J$'@E<*XO6IK";:*S] ].9USC^&XM
PQU@UX0%"1"TS)26[<]C%(_!>- S151/.+ON$]G_']XO.(TM0H$ K=JJ0DFI3Z5--
P^QF"1+2E'U!F_T %44V5KS<M'#+-P:G"5(MU+Y$J3H9'@WW>#8^[!XWA)+*H<V2.
P@_U-2,RVS'C?/18/'X!*(T9]=D7O/-XL"R]R,T5CQV5#KB4^7T/QQ?AMRQ?U +LP
P)]L**:5#N(B3[P4"P48@<P2JXK:_3"RS+;-"):D19W'=OSGYRH1 F9_)7V0IMRG9
P-@ 6C/KW/\IHH5Z1<D0)'DZB#,&NK?[!*R X_$[P;AM(#%V-XH1*YWX\&6=U61Z/
P9HVL:OC9!UB,6 $$0C1H?<(U^G.GIQ+2R\C(-FZVU7LAPIB[JT')DC<<$YH.< :Y
PQ*3CUB*NYMFL4<L:JN->,HF"7J5]''"D"5ZU6,MLA5' >@?R:PVYJMCDT[@'7V)1
PI,.3G'#Z:]KZ+@10PJ>(DU=BQ98NN9M^,[_B.[ JTP DW3#8)8\+R!&5(HA1(U+,
P#<W?'(,#_=QZWJ>-DQOWX+?MNQ;GV\>]"_+:( 8]9,X)521?Y=!$@>SZ.@7F$J= 
PN8/76/GW61!>)'HW/W*&NWR;:9H0M;(>JI@;.U\59*[E[I*4SS )S:'(*)XI+.=9
PQ[B=XQW;/J(CAVP72&%=O/.:IN#7-U,#YA&WXSA@><*Q@F0 <45G6!+ R6N>#!R$
PI<V\#_B^_LK>G25R\&'VS',R)+ZF1(ZLV,0;W749=S\&>?2MI=G*KO1 #=2QANV<
PKOD38D.WW\C_8TSAI*=B6T= MWT-0$YE4[:;?BO_$5>CX^>=I_MPX=%"G&VTP*.6
P[[54_=TPX0A1?25-'=B36=1V@-GNUM%KKM:M(TMI=L07'H,W1.KW6D-@PG8)(4YU
P+4!:>$] 10V[8 -&FD.BQ]0NFL;O:*@@Q@IR,2AE-A<=E>9I8#VCJ>=&9>[F*RZ0
PB<D9!DR;Z$K2%%J1Q&ME?M3=;]-1>G5 V48%8L=#\F2?W@BP:@>/7)5/?0WC1Y+?
PWXG_<2$2"?X6>1 7#U-73R<Z\1OV(/MQV!0/X5]#JSYAR_&H<Q$N+41Q4OJ[W+%F
PJ[6'_,XT5U-7JHG#*U&-&M>@Q?N1&<T-I2V\;<U:<\Y]*"%"X1BK#]W2TW=68%$@
P5JI$#"%_N]D>@DXX,9W=0)3:W%6"FF'ZY"*_4W)"MK/7R1?0KT.ZF!0*F&D04P,9
PXX"#1K9B]^Z2*;^NL^X>&]&XB-T]ZC%Y'P9<FSAM G]SE-@%J3O3Z5B9##&Q:9$C
P/%DL0PGOQ27:LLQ20?/?6F-'?\)4H+6[1J(<.6GBO>*,\V\><,^&XK/=0N,0S]D>
PPS!W"(QH(G!SYNKC?#?!Y!V<>'1]!,43JOW+Y2!#Y!FN^4SF+Z^;DHC@(2/0.TR&
P#Z3E[.KULG&MG/1G<7!;[LD4WT"T78:Y2G9<C))\F*^-+SQ(F:]-*O'-=A?4^4[$
P"NNID.!K_&ZL7X=@7Z50.!%8%U\]X24;X;<BH//Z%@??=WHHK^O M&=47HFR9=;K
PW;XH(W-^VT>!Y)RO2GK^#_.0RJYKL/2"2=S7TS8J",3_R<T):7X\#1@_>!6FX#I9
P^#O-/[(:4<P):QSS!1@LY!.H9^O]ZW1,OM6Z!\1DR=P, LXU PV89$ZTG2^C6]*N
P%$+R^>QK$5P.69]+]56-8%%[R1KF>S1',V3+Y7M%>,J#=_Z;1]:0Y .*[\-;$WD%
P R2%JZSF57AR>8?$8QSM4?^/!R((L84(ZR#@<-MT1SA];K9AGY&X+N:-H#-)Y4BG
PM%&Y]%6O51XBA25>(ODD(% _$#ZHG"Z>#BP=Q:BRR>4:8^>''1->;'VO<&V9$0V/
P<;I^F#8N]K)U>1#VC&/,3B-W+Y: &5M8+K^G*!X4!U&2#^PH=$>86&1]5Q#A23W;
P-9OJ^6([J"1H#J+5+0!MO$N7G^LJGIE"GN>@XO9[$11 @(9>6?#MNH3@Y6K@"X%\
PZVWJ[+G8Y[M1D?N6'S68SC.GY(C;?J>[1$K/)<JC/ %9*+M=,YV1?E7Z81SDCXO.
P")66.VZ]VO;<Y/Q2[:ET*X[8EKO=8Z]V. DPB?]DM]E*D%NIQ?2#YIV\NY7T:LEB
PG?<NY*DO&1(&=KX:6ZYF>@#.?]+W?).+K>,(P)<]Q?4_XX"%\@VMKP*_-H2;=?4E
P@Q"+OK@?U[J\8/W$5KS9CNHKJ R2TJU:O<&/*VX327J=D?3U./+'#-AP*4G8;3/-
PAS#'89#*UE!\&+X3VP'*[>BQ,OX]RHMN1A[5FX"F?$A:$ /+G^Q@1IN_EY-F*+,=
PG5?TO6)[+_J[2#7%&0=V[X@%.(1#IX1\V1621(LT:3%*R3$5VP31-L-?%_IQW[K1
P;(?/LQ7G?MVK$UW&L4TUIRAQID"X9PG/G =)@[.@@H_&^$F80$?:WF7.@*PFXB6O
PD,"\K#]5E8<[E8.O]H,SRH(]5[(CE5 N\#([N<VZ'R]JF84,#:Z)FH^?9?(<%W](
P#K'!7WO9[?18=6DGHX@XW5%V;R^=Z;]3YB6O"1D' /G,9$!C+ S(9/"NP*&,($/)
P*D3Q1-&I#']H_S!!X:MA&KL][M-6^C#H[QSEM5=0OH<G]0"_D449_GOUF$. XHUT
P5@-*^.EZ1(FGDYPYQ>G=N<I+@L$C-P'WIG.\>,9Y$7+$ NQY:"GM%0YTMWL9]6X[
P# MR**3*B[VL!4#D$=9P&WD8:+55:!6>8<D>AR%#G%@$\JQ"@;3^$G+C&\^.^NN\
PI;WHY[8JVSX,-I?N>.DVE+CW.'/Z I,CAI*Z;>CH%O1S[48X6'EU2>Z,UF$3'&ZW
P=@UN(3+0[5"F3O$6'J-V/SYIJFU&$\P[VV7@\ _\!FB-9GP73=UZ%<I:9^EW'OK>
P(_#T//1YSHWL'(QQ*WJ[!"U=#'T!(]5]4$"!XO_2K\EQ3?V5B0=[O'^$ZDNPU=^@
POKIVSWA7"_YX@85V /D_RZ]38P 8$28 @GLI_K': C/M VKQQJF(S2]R*](&G!_E
PGYE%0!S@<<!E_K5:E #657O:TOIXEA1&#H%CX)=P]EH'D2Z8]$L+91#^\?_L M(,
P/"X<A/GGF,*':C_>$F%*,$+@/(7KX&9EE!<=A,E17@$QX.H3<:BY>0LY=]_+;0HA
PJPI$S!'QM T%QH&,6!348<F23S(+6(XU^R$;/W6FR/$-,&^DIR$3S[E]/U+W,4\O
POJH#%>"4^P*OH.?'>#G0E :WGZ07:2A\!7Y&&*P)0/RA=SU(-!,F$J,\Z>.O>\X8
P(>HW>$M9/]<:$..POW-"[ $NC,R49&YGNVIBF!)<+]V\6&]$>""/2+]%,,$&K?00
PS@/>=AO4)\HGK=N_#9'BRIY+(7.\[WX@I/&%V1=;OE6QW5X032^>[H5P92TACY;4
P;O( $ ,[T;_LNYP=I \Z@.$(X(Z)*43K2F6=3BG^>=@O@B?+W-'.7SDS'"U4L;2S
PM! >PFG-J- B^6V*B X&=G*AH%(P[9!+;J_7^$@;4/[7-4>NER-KX9/TSVPWK%T4
PLUOL^C=**D=!X8%G/(5!ZSU,BU3AX6(@[P@YS%)N&<IAS-9#+S"F6$W,[Q)9"MVL
PGX\6I [.[;]HS+#4Z>&-N[3$$HC3V_!)]GP]8%N)C_RB0+ -DV.H_V(\1JS41 E(
PFC365=_3C#,>C>HA1'-]K3A0/=5L<5EP%2<W,@SED*Z./LI'">8M.9.O/W8S^ TQ
P%KBVF) )ASZI/!&OQ<P]=&H]GQ3?I@ *%U9$(9<:(%V%BV_.)DJ7QE,*C:C](=XK
PTBS# +_^>3T0U/[&WM .#*@& L=-[5M!'UDNXC,L[O\KI<% 2TKZ1)PS91.98"-#
P)[.Z4TG(Z-C9_@;PN>1R:OJC[0XGN!7W2!Y72Z,#^96BY_6VL*NY==P=YF\/RLJS
P'_(K2NN#Y(FDQO7-2[@4OI931_'5+D_+"W'7^(!KPQ39(MON-$BQ?L8K]/)PGTD5
P=Q_,>E&FY13$4OYNB"F#AM)F?BV_6*F9<:=>O;!_\5?=&BYW?Z;-'H4+KF/ 3QYD
PM%]\\5WNM&#5 .>K&M-E;0;/?,H ^JF!1DYF/7R\!T0 <4L'L\Z&C[_@6X.8!CR"
PR-.!Q6T!$1@&4[.^A8QC]&D8A(FK1*OQM.#)4H:T]*BM-CJ!*OLHEU 5:E* \4@Z
P(RM O-[:^U7<M)_N8P7L#%G ;.2/'2%E,2.45&Q6O_N-<1_#I#&W0@]5!Y,^.:MZ
PVEL$3UL W$_RNI<4:#/ ;EC0L'YE]HN@36>1_[^BA:0"L 3$,S3+89B&8 ;7^*TF
P/1?84F8R(GP,EK5:LU)8K>$ ,+)*[;;U#R)@:\7,IX2G?#A8CWTQ!-R:NA]F6II.
P+' 6M 'N[M[3MRHWOV%G+N#VH/G1@;T,XFH52W"MF_S.OXAI?KC 6Y$(Y8]63Q9_
P$W&U<K?O4&LL-0X3=.@!R%'% UEJC7'N3M>M4L;(I7*IU,A*$K4I?]?T#:?BKX$O
PM4.%OS8353K>K[9N ^O!ED4YIRQ93TXZQ6&?16G*N/J87\&WJIWA?V&O)'Q8\L1@
PUPE(CKVS^%FME"25#,L+F,W3/?%TJ4PEC <NQ9P@!?^N%N%?N? ,Z%>5IL6>R+,O
P7,&]Q9&[.4_$CB5JX#!I=0SZ/E(0G!KLE0Z;"><%CTD>*):*<[N\0@_(.['%4\U@
P9SP?]P]!B+989WX^O@I%+:<VVV&;D#A0USH)1%XH@1#)AI<K-*[!\G;;1<1)5>'W
PGR<Y=&TA%?,^&1:R)-(Q:P;!84=RJ.FY.(OD::R2*4H\/8:3>6/Q4DHD;-Q=8CDY
PEW0ONNU+]=G29UON(9-E>W")<N!"OX_*UI M_365@VFX:_#UXS+A/!G\!*-:;>/=
P2$B^<*12?5IAE8S_K0J<7;WU;TC]-?DI54K6?O.<A9Q':XCN\.KRRCDYTY^FF"DC
P=THW,V_,EI3VKJ.8>KC<+A_= -S7&C.FJ6I:8)K"*(T?L^:>'68>GX["C[I(--\0
PPD?WQ]2]!Y4XW(&)ND7CV"-O4F=@X*@V]]P"QHY&#(EH0YG.KVE6U,9=FJN9=S-F
P6.N1D7\Y.[PV6T!\V!;=#-* LB#U(!L,C"B A)Y6$/QIAI^*KHNIN?>#:P %9_8M
P# R%Y#4MT0RC6JWTDR?GNT.AZV?-#THYTHST+H39%1I<)Q<)Y>YIOP3D 7#,A((5
P(?P;G8=,D7U+R<OM"&XM?A!@O3G[/L#WS5-9 ?"(?%,#J+#:O2?Y#K.Y@K7?\WY-
P!.F]]6)P#O/&7.>Q7?!*T[00'N,^&G]SG.N-($(1B1F([7\4^S7I7BBZIEGL"89#
PV"E<U*)%'EC.\'%])#[<FY\EXKD#A[P7;'7#]O[2X11<2_XZM0)Y?!QZ80(D$XJB
PCP7/0()7B0O5_[ ,5]47_A:AF?7BY!3Z!X&W)K:679;6J-^:W@3]^\>M28XQ@X7W
PKSN;O@LHRDN*)$ZQ3"J4;,:V9I=L&T!(TW </2YQ\$)%MI$I;?262F)9HIL!4)S]
P>8]\+[5T#YHF&41.E-![LRIJ6]#1$?(ZBQU<7ZY61]@.^%SHBH5P[!JFR2":*8XG
P#ID)")U/XG?\[PW@A@5 Q^GL7479Z04UL,6SS:/-MN93(LYM[(GZA!'$I0S8(V5?
P  ?8SQ;,I1$>LI8^TN)(A.AP^;05.IY,3G+=C3W.X!C243SG045O-OE .2+RU4V6
P"7S0?:9ME=._&'H_)4=A[?R!IBPAW[ G_TJB:N%5D"RLV]E>H-/>S]&;O-LAX >#
PIQR:,PNY?S>M[$E["QU[-HKTRQPM)];H,0</$AX)(=UX<4,1)+ 1U]/@I'LJ]KC9
P.'OV&O7H=ZN"%:7+M_RB5VN HV8D.JO#& -+),G@'4*NK77"Y0:DL%:\PYBZ&-D7
P,--J[Y*:_>]C'O_4X-C+;_M![_)<8.;PTZN<7/0M_':X;&['X]5X7*C8?PJJZ:._
P09&2P?T9LKT&/[/#C.33IR$_>2>MH O/]Z5=R9X!Y.G L B$C'KH+VQ+@6_']*&N
P7]+DB3EOE;CH;PSJT$;B@@FZMOM%=S4CHTR:I9A+;#Z'B\<2#[\,7%P_K=^..S,&
P'2J %/(_'&G=,+<D'>]">[5<ZWBRN"@$3I$<C4SB<RJSMT7^3,X6OJAPD4F*\;QS
PC=(LOA8V6&)VL6I+-!>ACAR2ST_,X=L_F@/I[8!UJAR('BD6I@4D_=I.7B<L#6=D
P74+B#MD9%[L&F%1'CH"-+F7,H1:%AZ[?^7IRM9BZ*RJUXM"A"/D-'2,7H<+J@'4Q
PSX/O'DZRFH ?)Y\_GA8Q6_(13'/T8)$H6KP9G9H*[MA1<<;<9G5'!L9&1K$/PO;?
P()5:H+PWNWA;CN>^-$7K*;&M7L6F@C\)TBYCS,;'U3+S@'30@NI#J1C9YH5=T!Z'
P@M\F9>?X^[=%M+8"1"CUW6QD3##''- WXP=-<,8MFA@_@2[8Z!D[R>@SZ#WV:\O'
P%TL8KYS!$<0ZFH6? J-OS*H:MOON5GF:MAA/DH9C8JS?%<>.XXWJE:%@>VS3N+W%
PJXUO".-AH.> P%-%7M $K90WP -<_G&EX"QJ#.T25'F=KW MD7'-N,VY*^X;@2]Y
P!HSZ[;Q-RE=9JH/7N!6^(0>FO@A@*]W3)C33DBL3F+>8P%G-%A%5O31@I'P:;:9;
PQ..Q7%(JDR D]P#-HW;'@)><3\3(06'-895XQBF(83$\?BQ-80YPX"_SJ(C72WO]
P.)?^574:A;WVTE-9J XAFN!,94XP/2R^\A*(F_/9R1E*0Z&+[3 ?'$(XIU59JA %
P=GYE2_H24HE+_4+S[CS2MN\A:(0XX.:H([G\@:+Z^S@S;[J[2*)W^A5HF*H]W(=,
P^S#:4.%M9?2+\/P>>84 O1I7.BOFLTX[7*[-HI6 [0<CQ'B4U4I3 /\%X%T4"#!0
P+Z6P9/#^:[:4;3?J<T47"9F_G)$P&C7Y]^FC($R'M;!KA>1)+;!]F!G C%&C60+W
P'4J476\S :^>_C@/4-W3I='O0^?5W<'D1&)-HKDVU=L<@",?V(PR*M]BFK!:J!()
P$\1PK7(PCVTHH"GB%[DW##:A/4RF/=YM4E0%M1MPH'R 6SCI"DF47MN-W.OK6A<F
PDK7MNRU=QH\-LJ;-JUE6ZFN+"!RU9RR,?H"/E,]POMPP9(IFL4*REZ9;GWT0]IYQ
PX!(+/F-GDW5;$>HLE<@7][1"*Z..FB#@C9!R]IL987MJ3L,[W0?/?7](H<,XJ+:=
PS$B:,AA%F"9F 8I"9O_R=Y"HVK\EL!Y+9QL6[IL\_9<MVHA9V<6919OGSPN,_=HG
P)3PIG.()](\@O6A\0FMOMAGJN8R9]M:4 PJ</7BP>O7')T55@*)OJ^N",^CCZ9?-
P2TSFSV9"3 %:C -])[MBOW%1*P2F9]\6@A=6[DN''7,)Z"/>#D$3O#-M$RD 958!
P.)9OK/131ZB^IZ(024AD0H1D08?3AA9E%X2"WC)5*IJKH6O#DM E0#Z5V79"NB_D
P=760LTZ7<C(VEZC'D+ _L8.<Z^]O#\Z1>%'^003#M.!,%4.)!:'RFZ1%8L2S?GCP
PN@CZ'#;=+"]YT[5R05/(<PCXR?/;R)&1(Y"^.JB-6-K RW)=!G?8K%R,)RT^<)+$
P$B6-J_L&/+C[LW8T3:($>5C[;<@[A-';#-0<L R'P<QFJ7WM0>Z9UC/[]UW'DJ^K
POP]7@QVE=7QKLS/$2\@YS\L(=MPF "<-LG<;5*D"\)OW0R[1V W1Y9;DZCS06!N?
P^5/O)541C/VJ)#)>6P^[#Z82TBAX2(=83LG$3#52ASBUM_)*/JX8XH0Y9(8%^]ZD
P,J2PSO\'$=Y 2ON+.EF@LLM-R/I_-F5V0*&K1 ]^20\,H6:\+*E;7BX#?SUVRSWL
P3*4QOCT2$0P&B[_S?1T>>^%&@6N:#%E%*%QX]L[,K^FFRJLXY1,.URJ0F#;SV6T[
PCO$YIJQS_.\ ]>ELKPIQRHG%^46SCKJ$#X4/&CG&A@'UJLHI'UZZRNJQ$@*OE3F/
PF&#$IK$4S@Y*C..(S&96V'ZB:@J=4=M++'4)A+\%G*%'?1PGK#5*=IX6")G*VQHI
PK5_^25X\(O*':2I"J^# Y(ZZ%9]*1&6HNM>"6:R8\P!['N>@@?I?W]<HWKEF@NQK
PEZZVMC5N>,I(BN=4\-9N"0R\<I\GU1DSL:](H68VPN!%?E [:CAUH3" EGJI+A3Q
PMR5SA3V/R_@D&6D<R4F#!,A3/-VZG,0D):."@+[BVJV'3(LLP8QW0!08$+R%%)Y_
P6:OB3N "#+ E)*A 4]#<@88HA=[_TF0@UKB^Q7M(-GS]"40IOJ[6GR^30F8;%I%1
PV@-4VI;S3><:FQ)7O*4 ^B'BHJ=$0R*\F,"8!* F3%7O:XT 0.L/7#41G@HD+DF]
P0QM6/QE#R'_'%2%68XI!?/GX"4QA2&BJ;!?_65QRBH?5:UL9L$;^(> 9%KD2^^;+
P/EQ>W@4_R0/R+,(V.$BJZ?^.W=/OB'E(J>*Y)J$>OLL,:>*\I)3@%8F^IC#X\#]F
P' Q03]NV?RZG<QG.^6_]%E3J  -R<[JY[H3X'?&KWQRO4A-O/*JI8&?&Z;^9$N:U
P3(=R4C.$*9T.4>^X[+4L3SP$;L,L\"6EY=7(&U ,9XBP7=?4RXTR33-027AB5=)M
P<S-_C?Y6*'<XZ)K\3 #*]O-[_GH[E>OUBFF'6BU9Q%/MZ%DU205E]IW#<[BKG $P
PQ1\MM7&&3082[3FD!N%!TI?^CG$\0NJ'&;-<E-=[H9J2ZZUADE[_Z944Y>^H8DEI
P00\,_<3#+RN3JSJH%@D@.PTRE\4]IZ./%$V\@8@&N&*TI@MVF6_)'VB-SY'4QEZ%
PR<""9"6I[P$YT)NOX#M3!4')K23=PW-83.&KL5*E<:B*K?W>9Y3T" H/ ;B)[<WF
PN!>I]CVCF04K#@&B =Z+> QZ%EYN,,9)^PN;/8 7TQ$F$[W7YE=U0Y%K[M<]@1:]
PPLUO'TJ\9^/J-34'3;QL*:PU.+Z8:P,ZI_>^&]_V=C33YJC(64JK*&U"(P[ET$+H
P$GJ$J*P)_H97$Y?[@IT] 2Q,]U,S>$^3ME\MMJN);(C6"KVHVBSG5*EI.AVKSKTC
P7EA/>8TDMYVN>O.7T?0(&L%8-$XS*R@5DH/L"-5!.304U2$EAK:KZ!C-;UEY?#8<
P S6+Z/X:.#*V?(>?7&BSVD>?KLRWCY7>M_A=^B2GF44<M"*&CN3A<%OS<,:$\PD:
P35/X_P<M@8@@Z1'TI8?^5>+\#15^<?RA$<D2DRE$$_H ?!9U4*W[4?F"14WV_Q>U
PIL_+1W(9[/Z<#TWT:%K&CLG!>?B2,Y^#M3 M?TC^H8[W52+((;VSCD_,YE%/\#\ 
P5=5>C<S-[;X7K4XJM8SC1M!EATEF?"S]]2P:ON5I<2)H&X6M[T@>W7CC:E:2XVQW
PB50EU'8>6^H]&UA_4&9=;0H>EJY .;Z)&OCG$[1X:';&717Z^!1^P@DJ_\R\W.W<
PR^G.N< $4,#5[,?81T_9GPD)@A!K_N-\$<K+FWKTY!:6*74>&(T\)9MU4R4HDT=:
PIP\/GX<H&^O@4C!X<^4$6A #<*3,+I0YRC2\QE17-TKF OHKDA8KS)G\S>D5\<AE
P4712#6H M:"#$;"_IEE,F7F3(4>%XO>%9(<8 4692#[M\&$3C6.:JI5WSI?65%M-
P$XO4Y!<D,')&P^R%0'8\8(N>K<2GJQ&&*>C*7SE.2S<E2NROE8-:Y%NZ48%4*N2D
P@B4$W<;MXG#!RD\]%<'9V@SV\(P6X5]OA+)PJB-A(Z$XK''V8* QG/?*6T,&V;[G
P3"ML6U(+\]9!;>_[2NT;^ALHYX\SFV5I%4\I;'C4N8J5\#A<13[8^H%-'"^+$F5L
P@TK2,L4M1?FA;J3S<7VI)@@< S>WM+D;*J!W8F/%H]5W%A+V5;1OMW1)C).%TTN]
PZ$>U.(@UB*W7[*!B0JJD@S@S9GNGC"HRCD2W-NPSQU'N=*]"-O52;0M09T+8F@)8
P:VN7V&QU; E"T64Q"3B5B9[]@;F3\V4Q]:@3H2;I3VNVV,&"-/?@)-7X?2^U>0[:
PKG?G_*/Y9OBPT>_.PP('?,;#V&R+1@/#W^RX)^O^PMF,-'F8JP/[*7+.A=?,&T-3
PFF+272HPF9E:!!34#V^EL3_JXZB-M2$+PQ 0ZB!%P'^H%;B 8-E0Y$-:C+>4NE)-
P<"Y VZSVT]\5(\C#U8PG' 2"@0,V!8P-WY;^4LF?WT=3J\]#"(DNVNN6GFBN(D''
P4]MYM9(;M ?4D+RN7P+@H.0A@7=0V,["= +W!J3FU6.,ZJ]J 9=)7X2', JI7;]"
P<,8LL!'>;"<(9!M;/,YQPM*-_NF>P'TQOU[]#;/#MP;"BLP-,X%TO]Q?>K^D./6<
P-0;2^42Y&)X'_< 0_F<!T*-"XSR691;$AWW0*%5<7:8JZ2RO14D&F M1P,5JS3G#
P>!B_2E.R[4"]-T"MBHT$!+>ABPH$/Z"M8.S?8#D47\XMI'@TJ4:+-E4')2R0*+>:
PDZ:E-PC90I#- )@".+U'J@5UZB'EZY5DKRVJD^N#';KX-N%J'[I-]#+6H7!9@1MS
PPFA0\^TV:(&_6I$RJ<^ ?A0@@Q."JCG;U36*EB+*"_^TR,.ZA?EQ]#YG)A"A6):\
P.%;P/=9%,7(%?^#*Z^>"GBD3V\Z#U9]T]"B@L[[,CAJQ11ZIR9!4C]5/$6F+$H"E
P1RC7EOXZ7Y36BM+SCTRV;RR43@C^"J;QO1K,\?S+,>99"C($_8K 'IC+ S4MAN=K
PVI82.=4F7>L!'ITH\9=%]ZZGGKT/.;G(SB3\[<&G2:&2[_G7-D6W)FG]1FKSC*!W
PBA !>MA/+P[Y%.02>I!>)%^FQL.4Z74,EX%Y&B0=G\;0Z,\S;) 0G>686+O>=[8Q
PC*56;)6-E-,WIU:T K%DYIA[C%F)3RHZ%5LF4V^,E?J)!<+$?D/U#7Y4N7GT)$R,
P!UY1Q%!";JS*CR3QY6)!\NY(LTD/Y7XHB$4JZ XTH60+89"DO[!;&0VO>0H6P7ZZ
P6.(EUHHD7N$2-[*N2M-)BRJ )&Y$Y33\V[.9X\C0^N60-G@5]4]W=X3JMITT%<9K
P?$TFG,-95D/_\&/KN&/BP1WV\*$KX ^]]*$[:T&[UTQU-6LF>2;L2I)^RU8+ABX(
PCN>+BBPCXP>)OB*:QU@8KOWK>DB.-T<P@,3FR+(W\ETA93VRDQ!974VTY#\,3^'C
P]R6"IS.@CEG1)![@V5U#&4UHS;E%F<^0'7Z20;MJIU3!S,?O>^J#XF58N)QG'ALB
PF[=U&'JR"<4Z.9@4T!/D>J":<.F_1*QJR)F'-#RRPPKA^>KXAT!;:[ 5*8HP%A%>
P=1K@G#(V@E8CZ^GNAM4D7PP/]K'QF]B,&-FW<A%D1D@=I$K-PD%<J(^F#67UD&\L
PL']] I+0-:,8259>&.[#J:Y&#VFB!BYRI?1<>O=HIZ@7Y'&-\SEY]7EJ2HM>!YK0
P P?.VY$!F E/9D>47"R?XBU0VNKX5X^4N1G!G<YC]#.5P(77;NX7\([%2_4GY!Q(
PKTRU!MU#BW-02 ;&I!7=9SC%NK;+$!94Y"+=$2?^8[6G\&EK=>]RFJ%.3CI)RRUR
PWVLR_#I7 69ET B>QX3IGKCO!.9%"0!D%\0O/.TGQ0/>W!STV82!:I]A-L:EX)ML
P-NK;\E87FBUW85;L18D\ ,.:I#=O,FG9;>&A&/Q.+-Z[02M*<S-M:S[N/E!98 :.
P=BLX?CZ*/H281[5GT=\R%%A/R/FQ'#A-80K/!A7,>!G(8?EL.!-&QP2-]B:7^#"'
P#3&AR)UI;YI>&5F:Y7&"TI+3A* X_"0+GB76,]-7JYPD@=)66[L#5MA2KL!F5U:O
P4O,J3PO_Q6'^R)]4C .\&8I<&JIXH$;!FF.=6BJQ!:QFZ4;8:]U0GVG$XF=[[!6*
PT/&Z\#$95TA,84ZAD6:EXTULM%ZUH&MWIPQ6@LX=G"9&>DQF=+Q<1KO%+@A8=\_]
PDOJ8_8%)IYT5XM=&*8;:D5M=80!0C,AWT_.<NGG8K90E$G7:A3N%Q/S?"5Z-=9XF
P>@+9.*[IV2E$.C7"E-GT-V^1J2O]_F49:3H>O+7V80IV$4:[X^I[.N9J?B:N_Q>.
P>T?104ABIY)X3=+PZ.!.>EDYU;61L^[NTJ?/##E1V^\;*E4F0M8B2*HF  4^C&5 
P%J0EJL8/>L-LBD^Q>3L.>K0Z*5ANBE/SOAUGA9%96I-R'W!XX[/JV)O(>#Z(@CL;
P6>H_?_*#D6&_]=C_R(^A!=_K-J52_GM?"'8RLNN+?'U8:=">9P5N:)=5Z6NV(Y@_
PN][94V/])!"RCKY4GIIFTT=I+[C*^57"W0KC_#VWDWCTR<4[Q$+C'DO]UV]XJZKI
P#42!?RF-%,8.>_D8B ,#0+%J=DL#9$0&RUB/5#9#ZL\SG.WU3^\<[UAZ;YV\,O*=
P_[ /S<2PI_IJ@<;T+>,(R\1"3I51Y&.&?+[+()L F6[M* $]7+"B4M0QR_>M1GGP
P]W4+;9[49-/JN.KA4!^D$]?/[!>8T"ZH%J90#]M<KE2'3K#UWH:R.V/J0N!/>M;<
PYC$/->U(N]>:HE)_06]R&(T9]=\&*GP _@85>67'TTF 6>"95B\H#0V_V8T3MJM7
PKB_XP*7VS#2X8Y]&D1!%*Y'8KF^[?X.FY!+2^[,6F:?J"3U)]JKR#S&@0U"O%(&2
P,O$DB2@^+.DHXXQ8Y6V"KF9AYSV4/YZF=0DJ%+@5IXE#+)!%R+WTF#]&I9$N@A5K
P^3R:*SCGYBJ;Z5H2J>?0O2;I/)B99M?NH<H^?B]!.ZM_7.W"_&[S+6! Q" 2UTER
PS(SE+6[]BYT&K%MVNF]9,*VX%V:[P>LOY!IP&'$$\L/BT Z(75RD)?W$)2,O>*BO
P!.K>$$N&$'F3<LLX+D5)1_,Z$+WX&+?I;W#=N6%HW,4'*ZCSVW<*)3)[_56&:JBG
P?D_I545C%^6K 9]:&GV)>?2?V4>IS@W6 \UE6D4EJA<"^T@FB1#E/$2SH+5H&H*P
P Y*PH!#29I>ZT8*M*;+?$J!\, \<LPAQ"/\N_-JG2 ,?1L1C_>?;M.>4GR34T-S]
PP?Q.6Y'78_ [<58\@&31J,X33K))4P]P$N<VGE_G>73#(O^G_[/V13H@2!'VR):K
P^(4HA&UE6C!1_[H<986M;ON@W"^@_<"MW:&)J##>;LYJ[2)DI +M<^;DOR:F(3#:
P&WUB9;:![,4;%FWRHKQ?$KM.9I2+Y.]GO@D&S[;WI_)\EP-!"K'-_!? 0U!(0JA*
P:U:)($4-U<4?4!BA4@U.KZJ!G55DH8#9HI9\97YE:>TIV&X%KIIKN'=WTCB_]-:;
P4N@'[Y<KYOZI)_R9[%6-F>:GPK'T/5*IJH-%RYZV3T%@3.#.W-29QX*A-KZ%3RP.
PGMC;HB#;F"&W:7XA8T-JA!*XFH\BN^$19/*^6U=+U+"&Z98_!V3A#_<!3+6;CZ^=
P ]#B.D7^5>O&<![4AX4F>+W(,<1+I_[GK8I;%!MZGUYAM3L("^K&:I*^O7+TC"K2
P#<V&$R7\ *+:7]:0RRJN12%,DA)K=F]YN<!^N\N/VRKM=)MHIZFUZ'$#BRO2_E;-
P7 E(4AAXCM.:-JE;(='DQW^T0K9&Z"E%H#;\4]X&68'POU/T6?R<B2[F6G3BR<&$
PHQB0!3R'@OHN%1,VQ1'Q32 57<U:&Y^>F<MR  4M\9R#W(!0#\X:KJ5<FA-+ ;:Z
P46P:KAT* D*?RT_\[:1.IYVO-[/;L+$7^/6'9,OBO3;;0P$DQ!=59GB/Q#:WH'&O
PKEXRV6F^=S D69<Z&V81E[H(K :%*%KV]F9)/!F6PP#UF'7I3/*G=#%" 0/<>!>J
P!>9V_W;Z8+AA]:I>-U"X![BGT-BTZ):18C&LMPL@@D<Y4EEG9$N/DS[A5;L%JAXK
PB:5^6:*3)C %RP.T(P/>/]+BMKH:1=9AYGH<LAB;\?)X!9%8^!PO[TH2.XC#)\/8
PU##JSU*:]HB]YWKUTXE;PP,T6Q!C'R3E], 0Q;8564.=ZC+1:AW^,B4]HPT?^P8*
PSR9>@F 4 *+9<5N,F0USIK^(%"SK+<7AV9URF\I1T0J[RWBK-Z:-!F$8F.51JO:^
P@-/T,E;!WOY(,/6NW";Y6P7C ;H QJ[/'-G%6WHTQS^-71S+7@'1$X#38A,Q%UID
P?KR&J:3_IB<:^BQ&_P"W;=0K.&K<>\+R^G'C$*>2I8 U0N]@K#P]74<.(N"VMCQ3
P)3F)T=4%F0HEYPLOX%AWC_4SM8:3BQ/1.]SZ\P.6M6]6,P5QEM]5C<:4I<!J2JJ?
PI((E=.@G'4F\V##7 MN%*XF@W<$DK3P*^ZDFC1 9".^>#I+N)W@T;DR_HLBM/_95
P2D0^&[G^CO3-1@M#Y(/*7L4*#+4'F6[T";]M%#ZJ,ABM5B&\+#06.U6$<-N$#$'9
PM.%21:S]U=#N*_Z!2#&G+&6 ;N25?0'L8?@!>KRZ,)\C]8D*3/JK0=QGM;@RO\QX
PK\5W^D4YZX;Y\7!W26P"V_6[/*NTZ %;BH-%KZQG1(2WV5D@D0/Z;Y-\WX'Y4P^1
P7<9/BH<96-Z^:===9Z/7B;?ZY&.DR2@"-&36&Z#:+>.NG",*B$?O?9TB968I8P$9
PE0XF>'W#41:AK?W=3+>-L0[WM$\6;UQ<8*'F]7_MZZWML]8953=]BD9B(W%)2RN3
P@V!G=-!><^<H#618T=\4,F]S4[(TJ$KF.IQRL!]^-=>K\6:-FC7I6N5 R1@>J"Y[
P='0MOJXY*7-ELA<]TR<!)98OO^;Z7JWL PS4>'D#+UZ6H1]8>W?>LX1_QB4OC\)Z
P$^3),D*AI!S0JD[\KL'<I2+L_U8\([IN(#6??1HM1F$#..BML_$12O56[_'K@3;@
P$95X@W%53W>?HN)50X-YQ&0=-+,84#\; P^8_!18=%LT/"\&YF_7F>;4<KDAL1OM
PWL(.HC7?#%S,Q2H&6'9ONORA$-RS4R;7#+\AJX+J+XF96ZH'7J1IB&9-PJ$SK7RS
PB/PB&38G!/(:EWZ?VHK1T)3^:5/:;Y0/CB^,3_O) A\E+Q6<LMG]%.60M?#-,:I&
PH2JV4GS>XD@AZ7N2%+)R$LT(.ZKQ&*&#$?GD.&B:7R\JSYKA;L%7C]J-K5FBQY-)
PE<9H2)#U5["*<C$-?^QV2$I*RB_6*E6MP;G!K.C \+SK_95U<BBO^2270B%KH!>;
PTOA/S9U)HPW*LB-:@V&67T+5+HC^-)+'PJSQA$(1O@T?4!__P9@9&<C2](:@ND,=
P/O/J?"-'L5M/U H'7U66%D&<@0T6T1$[I"H!2#SU!S5'LZZ/!>&P6 0KH0N3JFT&
PRGA5_5Q'OW=._;KA# A+WTHVUW_T$0W?<"\?SHBZ9+\G"#!ZJ]!*I0EN ./0Y>D@
P:UKP;1@=J7Y%A@8RK5Q@&V+DTOQ5HA[*ER\J0O)T\0*4^H"^",)VL;93U_394M!/
PI3F!,UF6<('9K$ OHBO=*@XFY4)S*KFY3+7&F_NCJ[SXS\[]0&R#!8F6ZT&._N]#
PU-GFY8<- ?8S_IPF>G9[U"\WE!P*/2Q<;6T_#;0*);;/Y[JD8H"5,]_VC0R$*J-P
P)GTJ9U=T7E_UJ:31LZ,-<19*Q?^Z.5_+UO+X'WQ3$ Z=L#GX81%Z)(WHPLUQ!J*#
P, EA)Z6<\^/Z%;8K_,%7.E X<'0UW^F,:?!(ZFJ!&QD.0[@(_*+&55V*S#=?UQ@H
P(&0Q.$/=T/:AY+*.7-[3!(J+0P3+ZUJO5N2;8M"^?XY;4[''"A*O)NT6I8:C@[AS
PPI%BZ9*Y5X0@,8GO^S)V%H \W.YTTP1S,P8)F86$>DKGF IUU$"4!B)$G45UZ5=4
PL;A)NW+T<=(W!44R1L>/)%G"OKD=Q%6/H&IOQ>B^G8)3,Z[#M;1.(:S?'L$S*)!Y
P&VE$A)C.PK/LX[K;*7**,I*+M_B,8M_9ZRZL"]J-Z2D,(K!)@?!ZQ+VR(GJ(7-%2
PD#%N!_ZM$$GT3KA10]C1;@7*P'+PH9WM(TJ2,6'&U>IV@S]DX0TC'UGS&:-(4+"5
P^9ZW<R0RKBF;0[*T.I-UMKWZ(Z5,@^][4G+>LC/<W(N2DE4C2LZ*F;'<3_1SQ0GV
P#_DD)&5D6%K4$D7XW&?O,V J^AA>FKK /[@?V%S*R>27E90IFY;8@7:AOY N>"%K
P$0EW<3+?8T>&VYU=N5)L$3-V[[_I0/5"R -K<''25R_^V5X[R*.VJ,+>OKQ=XL:J
PB^) \X.]YI,*09MVX5@4<>R^' LT2^0>OJJHNN<T;\X,..XRW@ ?F\VV"V"=L)G-
PM0\XFJM[ ILT5>0Q?I^"9*P+KZ,OQ<6>+,,XNM'/Y98(!WRUX:W'LGJM\4QY.Y]@
P-=D?BTN''OCG*D)U3WRT[([7( X&A\^UG1)\_//]&C_.9UH\>A:$_SRUB\#S]2?6
P2!*UUGQN1-7T755\6:XQE1CG)'][/KH##I<#0=XD/"EV5=27XPPYVG"ZZD+GYLO0
P=XBO0Z%A9L4)FGRC@G%L3G[MV(4.H.T08-%/_AM9O&=+45E5=<.!H=<! BW5B7U6
P>F<#*60&>C ;(KQKSK'775F1"!ZI,4"(^#]'4K)^F-1&YQ#=)TF!Y?EPX\8F< 'U
PLIYLZ>CM4F57/7 X7G%F840"'&JB](I'VI6,J^NS1GC'FTC\^DN4QO)&8&Q/4[.A
PIKQG-F6C%#293FZM7^8QPX[Y'* 'DG!:9F2M"U]R;G\1KP*5ZV# Y*Q\ ,'3^YH*
P$1)E,:Z^:PS>3[2>F9",2/:>T0VL=/(:6#"SR@VV4Q*NPX9X=E;V&0<%3FM0T,N&
P7R=#=5FQM<\&3'[/T8UQ6D)C+F4'T--Z,8QA$"N0EXRGCPSZLB!&G1!TFPCM:&;9
P=;=GF1L >?G %<:F6-W>N\3"[3MC(FO+;8QAU0[JG526'*D7H4I:WCLCXKW8Y'S?
PS= *&7S7.6<J!W6E,5NL-ZU\I,.F=[$WO2IM$.\;2-I] V/2?+XFL%;9C9MB^).4
P\FZK%;AGS:<Y"QZRK&.<F0?$?L4.TA"D<4.Q8ILOQ^+XRUK?(VA<@5SKG6<UOC0A
P;P5//*Y\(X>+":%^GG;!F>)OYPQQ==-GD&.+7F!TOA\F*@V7GZ&[QN2!)+/MQERE
PGD28&P2[O!ML80M'*\_B/H7Y/63KW ['AC0$LC% LO_:O9T)#$F_)OD1W/X&CT7N
PSN'T8=U$)TT2//GE G$;:W<6UT,73@6)4]Q=0?>/IKEIR"U"\S=G=\?X@K6+B/7L
PF;1*H"H!(JSC:!C!@+1;TY9\GP481NMK\SAN]14C+:%.1?G.+S%1L_& 6@ 0-B#A
PMB!!ZTH;@K)8 ].7.E7+J\58I89:B,8_JU11E0RVMT,9=2A")2HZP4;=HF43LDX4
P;[SXZ2Q0]U*XE,6:"Q9"W]>NCZM'<W'=G8[^QZ\]*J;1J8KQA-E,Q.=I52%3H*-T
PBHFM^LU,+TR1OJK_"S\=;=OA.\ :Q9RM],Z.XV-VA9^5X,=&J_TV[4B[:U2[JF\$
P P1/@+? ?;1R["LLF![=YB^F16\ TPF3ZBF\LPY0O-_2BNXS=R^Z[K- >^&YRCL5
PS0.$$(0*\[^-3[5?GOYN.;, 0[<49\G^W3^T=XW;2G0QB>"5D7$7V=+_#8KW(VR&
P$OC(PT^U#OHVS$$%K^['S%/-PJU1\RT';@7#DZ"J/XL:[OAKR7Y/6%S/D*X,TQ^;
P _\[AQDJ31-4'@!D"$/$C1BP167/2JF;V5:SN9?H1@XW^E)< >HD#[?#&YV>9/JO
P58C\#_Z<L\:,GU"A-H51G>/"0+'QB.?V(_Q:UA\7S'$2X%LW%444\J8VDKA80 E(
P!/444FMNG+(4HM,&'''1 &'J>Z(/&IX!%K.C]7?W!$"71"AH. 3)7-<V0 FAU;L,
PXB EP!RQ3@5K"-BLU?UL3&'_8]V=,3K]IT"1^I-!CF7)X1/^B<G9]SV"(2]'[Q5>
P9!Y+4R-*!O0I^ DJ0:"V5-,E.H :D- :, '0=)]6XRZ23ALL 6+A#^\PYI9<7\=1
P B4\M3"#1ZD)IJ5W )[O?$]B2<0S>E3%IDO4U\L1FG]>X[H6LC8+@/^&7='V;P$B
P)EJVZM:0%-_-*.&D&+Q[>YD@=3CZICT&V39:$G1[H#&A2TQ)2635P.A5C78<<*$W
P[;BS0\ _#=/,9>M0[; 8:2*V@E9D:77C@*8(1<?/KS[7>F86D/Z(T3;JJZ1M5Z?F
P(5E4;PWIDW4PQ)C,-?H!53O?<'!['*SG%U*6BEVA^L<#CC%POA[83BF-Q!/>>D1!
PHMB-#"&],,'4WUWK  ^_#8;_J(7A'B9X4.L4!10-4E#7?4KT7T;*T?L3)\BF0MXM
PY%1UT7VR"'N5RNO.U:+HC_OY.TSI&7ILMDBVJ2><?D2"70>W):H-P26Z*_';OT:*
PVK)=J_YT)Y1NW>:<AW%_^_BCZ#GH9YS1Z-%LCEKVIX_A-.JZ*+Q H_]0>.IF;>5(
P35#3J@3J+LWYR<UNCI93&-I>4C41L+) <R$]H$YITJ0)=N!'Z0842X79WD5%0<I@
PJZ/_'X%1VOBGP@IAS2C\BXF=?*/WW#1_3E TJ/AL\YY['CXX2,![',:W$W$,9C>4
P>7BAKKD_&=M.!XXDRU/ /@8H"UY$E63J2,^I'JF;9)Y].IRH"Z"+/,D3-5_!WW2<
PP\Y(O$?Z!'BR19E^%SQQ3,54Z\0TFVC4-(?#.(@]>+AF3R9016]? \E_-E X &WL
PEBXOH6.)T!5C<D=TJ>SJ<K:V;*F@]JSC^_V_2"Q%T]"ENDT0+;Z&8L>%1<Y%$PRT
PRK96]M8:<QOL ]HU?!2(D &+B#=L"?GHG.AQW?CX3U<M73Z&! JC]'!6#B:1R@*[
P&4]0%FR/]]8_X0C'&_,+"G>]G?:WTNPG+%4TC0]F8 R5:7O?=0(DR,?6; *"S\@4
P#:+2A[-C206>GFG)"R.&PD5W6]&XO:6I[L'F'V9FD:3J('TS5-MRT439N_:*)!*L
P?X2Z!2C<$4XFN<?CU=??5-B1RQR"(G0>B1I#-7#5=D^BK6C2.G2_SZ?]E?;*SZ;6
P0ZNV'^R>;A_T $*5?:WOM*C&*_94]$ HK5DM?9H[!V !1%W!J514D WE#W)X:?[L
P <<SR?AO5@G*,4>\9,D);9RAGOO2+C=N??0'U9P]R!I0J;>Q]7:XV,34#DXC^7M+
P@BMG)<C 6DVC[9L/9XW,4-83(;WW<X?RAY'YCH]>Y%1[-H<'EHRXH&+T9GF<X7M]
P\B/?)B2$T?CHM@!3M^4I.PZ1L_X[Z^^$9':"<OT%@*"I3P/;O.3<F.>J]UINA&7'
PYK0=K-]#<ARI&FO5Z1C-)LP,LVV(TTY'YYF^3<\2A8:LQCE:T<2JD&YZI6X"=?KS
P 8"S.,PC[JDZPX:E :1=RPR^)1O0TAD[@5L"<%LT986B'R:+E*NX,:5W-HB-@*Q;
PI(^1VE&K6<[81J;=PUDE".KLF6-13 *"IHH[33[2!N.8,P&6F$#'_!\J?.TQ1!%A
PN5\MQY@G9F&8VAQRDO$/I0[B*"CK:DC9J.X'(4TC ]!,<V@>IP(KAFU?T<\C'!!#
PB<1M1NO*<7.[;AZ?3^GMED] ZX^;F]ZR;_SZ)U"+"M\Y_T8?/R44!P;J^E=L8.1A
P\.C=W6I[#MX&\/@3L_1_#396>88QX^ZQ&1<@=1W)U8W)O/-R9D,6Q$RW[!6MFWUH
P%62\5TD0X&AOEGF%PFXXTN%FF3@J?\- ^[.+5"UV;.=HQ[H?*YCC+__&D,Y\'Q92
P\616CR3GS)F+/1/@J4G+3%1=)*9_'.\+7-+O E5E$)5^;L SLD1A;/(4'I["JFWG
P VP=RFE=5MDCOI.6K5#B^@S%W2Z:))>I&ZK,",RCEE7=>KG[7%,8FH[NL.#S*@ 4
PSF2PA+6]H$3);.WT9-0J=P1D#YD^)Z5E[);#Z590?S]QN!Z=8KP[0*LN%.Z D*0!
P6ZI9H>9#XHJ3RF(99>UD:+4PKUZ[=^Z?]5Q<$G8YN:[YP#PJBW0!  [%25J30^60
P;+)$@3]BXH]K_P;2R"T,OK.AC!G1+MM=O%Q@R8F;P9NX=71:P0JB$-:K9\W#=]\6
P4\5+W7..#NO=B3YW8VXBDVHE:Z.67JGGLD40M,\NXP\\@XA*[5_+C.&#I ?TJ8%I
PN4'@!:^6"BU&]Q\4OA%:S,2F@IQ\8F$0(UQ-DKZI8J2,L)M#0 (Y65\7![EZ4T9J
P"!J(2ZV>@U41Q4+#X5+M,7L@\VE/T7<LG=[2>$7O!:/%.4)H1R4;I1'083/&8\ZR
P4889E$<8(=37AO8DRYF2.W7T,!/DS0[/-.\A2@N_FBF#2N>9JMR3ZC<PGI^W]$T3
P=@<_O=3.'RQZX'^Y?%.-!J$&36G0? 8<H50 TJ\G_;^7G6[BY5#7B44B59<#!I@ 
P6/J:%F[$INB44&H)E9AARG DTIA\2#;S!%B^XK6767ZH*"ZU;K$F?/$)HB]/SE$.
P_>,*%XM6<56(@CKAS=/\VWSL=D47C9;&.%PGO?Y(*GBNJS&O/J$^X\")&;QNRQ&<
PY5;9[''\YSMY:&_A\,^FK#W&/H/PR;WBT9= DJ=6L!A9.4@D<&IP[9"JNW_NP:;9
P,N7&!2;?I)$8" ',V5)I-*FZ[Z+"R[W[U=I:3MF]$Z_B<.Q/>+R2.$--.'[UF.P7
P7'8%5^Y4T/W]CCK8:3[C"YXGAU; 1[;ZMM:L3&W8.%JAOYDOI@GB/5IA)5C>9OSH
PD[?KJWK R [W#/\I\;J ]B*C5E54$H##LDTWQXJ++7Y4-.N3?4RE4//&,@\R['$[
PVWT<MS22(STTQ1A579J@LK)_P;V2R9#X:[_8P\):] 6W;KHD1%@[&HQ(W*J*BFN-
PS(M5YTX\_2]8&:P.XQ$A?RMMS-G>@M,+^Q>&5=P 3_'WQ"TK=P&[."X;7D  _C&>
P-F(7'X(D)WJ8'@<0^65&%/ID)9'. )B!:2NE@L&YK&-N2KUS+^B8LS;E#C<P<?L)
P8,W@7\_<T,JV.>B"X\_4E)WX^T.F9B3>WMX1230/FDR",,T/#3AI(KF"#:KV(6(Y
P; ODAUGGM&AJ1,&:27NAN&. _AI$*V])^-5GD@V@9"XQXA(D@T2*W8 &(U@J"4.W
P9N*7(_X]QAV29'</>.DD:BJ$,;14LU_[ZS?%A%AGY<XJ3Q&< DI%C"*]-BK?E:+Q
P+3#H0UWMED9T<=_?Y9.K:LK7FF2E3F?&VO]:2_$') GL:X4?-/B7+0!\]'..^CO9
P76&1K>O_SR#"B6L*^&'7(.L;9J&\U:,=(YHC)]*K$ #U(W8X28$UGC6DI0;;Z'V-
P*@&]FY>0X1!EI.:TM-(GI'=-7UNO,08P0_CF6.LA'$MP(*;[+P]<LT D]Q4D'X)Z
P MA>4'AC9Y==RT"(+S<V3[@_TB3&OP*04R5E<LQT%..*Z^1E54C*92YH]GN!*YH(
P39"*D[#CAR#@:I6-J(S0$MQHE?@^)H'?20N.L6<6'^JQ9ZEAO#=0!EZH4ZH(DB#7
PG4:%_O,R2'^=W'2JOO_S"H97?-K3/MBT -R"<'9=1T_YH Q!>O"'CQ5Z<A?RK;8R
PG[(],JY=^3IT1LYCZ;GOVO">D9[C@/F8OUZ$DBZ?E"V1=-$<RT(G.V#K#^S\NMY\
P$%'46;VXB^9)W>1F 9*-E89^O6<HZ2!O8: -!3/T,ISS>\98\"(^5SI40YT8*:3W
P(^FG]KFNL:?3DL45"-?4_CM=EOV!-VM3>=_<!F =CD*I+MFO5JN^T_EYW;6WS(6D
PPYI9YKO1J2 D*\WV7H\[C*!/V0NQX]W?(V/Q>O;10%2_]3US@L@&1?AR=+[9PN>2
P&JSKJQ(!64Z;&Z H#WA&6[$Y,2_ZZVKK>4[W-J,VLN#&![SJ3=;<'7>^>G*71W'9
P&3+6(RT@B[::09<@IAKU)=H)&W&-?&U(9;>>VPYAL\75_=B6V=F'TSZA-Z%+K=VS
PFZTC"ZHF%ZQ5"FU'F::'T<O/ <J!;NQ]^4^AD:GZ/WH[DM0=VPPGVTJY)[', ;.!
P.[N0X8[3SI7CI6PI(A$B#Q<\M5M&1D897V3-&4_V5U0 \_<6U<J4G<\;%"-<<B\)
P<XY;<)ZN2,3FL9,B9C?ZF!"GSD_>@YV$Q(,*K<F?IK>K?O/KY^)1F^$[*L'!(X7U
P):D8\157<27+T(0:F87J]7Q(#?(+.$0*FYN+B)R*Z745=T!,[>K5'8.LL.#-%,#B
P2O_>(# .I4&BC!VQ)$[.1[-G;'Q28K#9.,5.@C4&L)G&\-.KD<$'*(WE'E,3M-*<
PDXAR3CX$/O]29K_U Q0+ZT72<S1Y@46=KNF83N*6?HP&8/+0W$6)5'XKTT?DV$.G
P')1GZGAZ_+FD5)F*7G"$)-HY3T]DL'!"H?+=L?:,[U>2.J VDW^-<>'"Z"@4_M^\
P4.SE%+*N%DS*CS]M49 DW6(6CTWBY)9%\,6VUC>,[LT+5?]G0H6[E=_M\$_(O!]@
P?84M? .SU U4*Y85]?,>'EL?4]WMPZS -_14#+T<H:6?KH3+:(@S%P!-ZH^\P <J
PCW1[=^<2EJU[DK6AL4">W0A,'R@+.D^F_E6.6*=4O)7?E4T)E71YOA8:6.JC3D/F
PM8#+3?HOV?-%HY6:V.4UV9_IS+H&R$W]HD[^<_&+VZ%7@3RK0[0<DP;:V^!7DR$H
PN'I-GW;CO GIX+RX[9/H2M[U3294/[@9!*-R)^:O8^&BAEK?C\.%EV*=%!$7%XO@
P]78+YP7#H2PG+RV*Z(SEFQH]3I0"1$1?\S!5*G"WILO$^EN*9ARG'WLW:A;HKDC_
P?U[DR8"!*K80)!F/HB_K48H3W/WN2C"S[NI@D)F-"PB4QG[Z,&Z_VB]A)>:]/<0X
PKT+^=<KEJ*P#R:G6S[(-O2PTK%,S=]WN5KV!T=5T)'GZM(H,?FEJR=(T 9Q"4Y8T
P;$A>!A=K=<,F%SE:(OE0F<7SE*+XNF9Y]V U(.;'1YVF<=R/.8>>65U15!JF^[I]
P;HXC<.(C'XO!DY:LD -S$3_75W=HKDTD4=X@XI+:P#%9#"G\S$@&FK;//=%5_'O]
PJBGA!@JG$7D4,7RR4*4C*7V[JQ"N,EVW-X,A/P4'GK'D=K9^9;"K"N"I]DJ91]JS
PT'@4@U9+?2D:POPB[!PKBDIL<G;'HYKI9+\32[)LP"@DS(4;7"6VIQV]9=9>CS !
PO\/9!JHT<0B#?@"L05<.HC8>L;^K?= V;.K73?F7J<>_NZ3R#."2("2[>WE*!,7 
P=]#.S49PO).4J%I?/0)_:;2Z,GUKF@ERG+):!:]M9!\8Y KV:JB>,TNA9<WMQ!=W
PQ%>OM'QN^*^A=WV_QMPGCOS+/'=;E[$EL:G+PS'[CX_,:G_YFE-!19""@@G'5QO<
P4A;J3Z-'I\D9X,#,S[">H][*EY4A!5KZ8Y5I(&5B/\'4J>-*+06^ SDEC//X"38W
P^[G<).P;/<Q07WV/?.QXQ,IL(*B>:!;%?</4K+C42?O!7SQ.WZ59[#,INC$+DQ*[
PF2#3V9 D9<@AU(XP]XB$.LW6T:@-D34/&_YK4A8^[11?4N;A-)I1&FIO5IFSF^I3
P!\']VE9L!88%&HL T?-K0P]TS(3?!YPP(;B(?,A/OL5#)FO6#+!@15N,%[]0_+OW
P5E(#Z>(#Z\=_]JPVX ,#1J)E6>XBR'=$RVU.XNHT.8CH [9C 1(/>C*. W^&4_#Y
P@V-)5*<K/&><_'T0G&1X.2?(55N;@U?I@H?@2L84^X^H=KR"Y0)QKRV(PNI$V)O;
PI=19I8G';4$?5]5HK+5;/];1BDQ H<]#Y$VU/YGPU>,98$'DE:W^%W&:416$_[6X
P@(4@CS;YZ FJK^;L>86W4SR-&GJ15U+(9OMJ!T=3&9_S@2,'9..[X-^6OOG)GCUO
P_&EGATI$LQV;'HS68\<!B!-2KM?VW=, 65 C3F\?:>.3H&&?)*QYB)GI7YS2EHQ[
PU*+(6,".[RR])_ *YX@R,9?:BX?W+702G"_A*]^]_[+ H-^O F3V)L^.:&'OA!LZ
P+4E]W(6EX6I>EN2]O);2./39F@X*CAQI;&!T\.X8J3BB#<@/+C/SC,RW('V,*HSX
P&>OD'7_MGBYU1$.C'&4<[?4HE<,<3EW6)?+M%JC4O!#LWDVU-66"M\<FJ/3C@Y_B
PK4]$N0P_C^@+TM.^\"W,^\075M0;QKA./KR7G-#7<9M A6SSRS%^'W10Q&F$=T0[
PEA_#Y]>>ZR[4TYYQW 0EMYEW5OP)^LBV[!'Y #R0-183]XOTWQHS@H,Y:^,F!7$J
P(!\VU9V8*7OIK]]!<TDZ$!-@!I4X7Q!GZ8Y:/( --K.<(Y_1E_QC,8_,,O;III0!
P(5>*/[E6A-76I?O-AK089&5#A/CTR 0W?,?^,E@A-:: T,3&Q-M!-"P(L70D$\VU
P>_5O"@GG/%$7/D:GV'O@42<Q*  \33(OD&YY27X6=NA?*:_<X0F3CZP"K=Y*UCR0
PX"U]?)6Q-T?&6F1D3K/&CPW>5HT#+RCV//<,DR6-F$_KB?]I?IB)KVDZP-"T+9VR
PP(<5XS."TCW;(GV1T'X!<6E7;9NY:#3,<^;+5282,JU%.FDN:8V-?A%\H$2#FYYR
P25W72/#L+ Q[+@-4]ER1*BP$@=,;G&*V,_R[%!_Q<A%>)+RB,V_%DJ;]X!ZO[B&]
PK><#!Z2CCZ@4MO<_O@3-TPG5@&:8ZI$"JXR\ !07SA?2IB,%><:GU+KWL*SGF(#W
PV#/*\KXL4&HZR@8DBXAE6";PAD>U(O0S2)BV!O1Z8W["S%^RC!7ZJ?/'ZV(18O*"
P[*]VTS!V5Y=DP-#%<?HM4'5&"EJZOSV8 C'KT4CE^]B._;LN.*L",JY"_J.,DB;@
P8;BCD_?S2N]C09YM;!<P.I,6VU%#6<0)C^/8S.T269_:RP&<@0Z!;LA'HE?:.?N,
P=7E]?L/X$44J0@"T>F7\#&\G:_*%/C%K[O8$@/ >(**:DKEX:\"I^9=Z38,.I&1^
P6U5EJTMZ1D#IS']EU^#.J*N1)CV>P!EE?6P>/C/[-T:99??XM@O[&>BFC 9X+4OG
PCL@=+CFT5;2=57?5*YO.',@\R@NT14@ "<P_I-1E)FJB=2J>!2!M&JVIZ*>*E&F+
P(#<&G:U\$?V*=F/0DN1)IZE'@R4URY,4=%[6H8$ R1ER+ULAF5TW*_J8NUWD$8^1
PI+L6GS&C$E/?B(9W=O2B>T#ACN@3Q1PD[RKL3.5>92?'I/&X->43?VWM ZH?3B1E
P@#;Y]P"1D@86\RHG8Z)-S.7=D+>6<&RE\9.WTX7QMKC46FL>)N1["[N(#+<SFVYR
P.6U@AI[_#T!<QV!$5907IPK<\B,2L:-^K*0+X)X60YU7G'20R0!O')!P.XFX,R!!
P/_2688+$#5*]1:'4MGCTKY56N'N[)1"[]'TE*$=8:EGZ:L@;]<:9E_YVU!F6.1[%
PPPG&1)W%X.[&^@3#1Z_7A99!*3J[W$RCB7;A6+I'LVBPZ)M5\66=FD>\!R4R*\Z]
P>@>TJ&C3B^^AK4#O-O7.Q$M14WE! I:HHNX\6ZN/9<6R ;%-I$@&%%2^"0KJNQ&!
PW_9::_.JZ5JM^52%\U"!C5 I_I5A0:V-)IJRM\ S(%NSZ,;W(!E;NW#5A$2N)1B-
P5V]\0^I6TN17JS53VC)KLWA4JD]4#2W+I8QW4U88DGZ9]_R?UM8">"$L6^:ST7Q3
P5YN2,[Z^1R=^;PS)\F:/9^;(.D\O47O](@[^_D[4')[!.RV#^W.0\*$GI!\!(Y2?
P8QV3ZZ,4I)2, &>?>%8J?_6"F[49]^^6-=JS**<ZW85&WSS5\CT[&]@V44QZ!XYR
P2?Y,P+5^#+64C_+B$9[[@,V&+9_0$GP><QRZ._^]'V=-1-JM9[*2N/(:;5,@,%S/
PC EIGF_XU&MRCMKC^83.I^9<9<%RI WO+6LP^""E #&0Z#D8X]D73)W&FM$*Y,XJ
P"*AD!5MU/Z%!:+_,A6 6&KV:$*S',/;./9&-2E%!_AMAZ)XQ$H)-?ML%Y2B^1Y,+
P#OK\,99M9HDZ2\2([=(ZU]I@7SKO+A6@0_WNM>3T^27.N8#.["53[&FMKSI3FR,Y
P9_U\#[LA^=A!W2,PBR\ET\)$$%G%L8ZG4XSD 5;OT<[WI8@3_^J5_>KW\B(^E#K*
PK*OE;LK KJCS@UVO(A]BZS//3&*T695J5*\%+U>!*5IR8)&9RN< _7X93PMV?YZ#
P?:?K;3H+N\_:]-Q61#78#J#M2__I9\ 6%#DGR)9\CN6*8-UIQ@NTNL!GOX%=Y5=C
PFN-: *8>!1#"9 /XH<F7EI^V6"]]IW'Q>'!60A%U$AB+DD*H&V7,]=_;V2< SH8Z
P*/^1C+52::J*'68GJ 2=&E:,9'U*-S2@Y1VK51#***CBT]ZC4K<9^06*!>'#%_ML
P0800":W5<+-;5U]1$<T:!QJN71LK"P,P09M>)4 $11Q!&-Q FB*%OV\[>K97@G84
PHY[S<:UIC:TETWQUOL3@OHM0KJ2_MA]OG.BB@>#*>./)J]K3IUZ3=N/'5WS%Y9TQ
P23M#V&#(![726Z2:_RF@K;/F4&K:&OA[B#+&:'".FZ1F1P&9XB@&'&1\3*#E=D],
P;+'3Y;.12EP2;]Z:)/:S#QL7B[R40R=6_8BK["'M"@M?'SH6,]ZWC_EZ8:B?.F9G
P]S5D6/"HM:@]/^)1%6;3>>>WCX:?]7Q>5)A7:@I^OMG"QC<G*>\3((ND/]3 CK51
P&9M5@;S%8" #^HZP_W%0-T'KE==G1[^GQV)"AC*S[.IF<_G=D.>-A+EJ@#=#P8;<
P2E)!:<2,XN;#R,BK-X."SWW&,^#_]-U+A6>NRZU94=O$)]I@QKZ"\TJ089-5O8H"
P?$?TL$'@U^?EX;;OCDY96O4-W2E@ST?)8*20OFZQ$9:\IE9 S"SRB9-GXGDT.;PX
PXE$]0HXQQ+*RU2[V)TR//7$J6]")IRPA#;5V\=79LMR-4%T#"V9/Y)F\SY/"VK<T
PGF>2F_D1?6)./F[=D: UQ?Z@ZF H;:BU>K5W+=AE/)R" @JZX;8=,:0X=U!&259 
P4[:B3CW3?9AA ,#3REKLM$&T>;.KOBW&]1MND?2T1XY"T-.ZQ#4?,:M7.81)K-G(
P A8AK+G^GU8FVB@=MQ8J<]M$O>)AI)43$'<?2TR<53Y 6$C3!7795>HC'!M[/V?6
PHIM,6]&%VO+,R2 _/6OUO[U-*222$\Y'S5;(^!LZK*-R7&^O>-^#7C%AC>.G?.L9
P2&#RDU09;1;> -)M4%]1BXCGDH]971#O.&0TUTIY@QGBGA#&[1-:7B]BIZG7%Y=W
PV7<C0ZT2%S%"!C"E)3ZNP C4N$>T;+!PS(0SP3"G9&H.!K1:P4 $JXAO4\K#!-C2
P!D:E.4LZ+_7&;M&FA>49B_>0J<[9%B//M\(D[,066ERS1FW/$AH]B;YT#RY+0=L6
P.C$Z%.CHND9O)@8&"F?MY77VB5DQ%P",X:*$W[1/.E+>Y$%G0\ ;!3X;PI+&[!&=
P0Y H'BX"J?;*T-V\W@4:%+@4*>E2#D]H+\D"/KN]E#5S#*M<-FF$WDX>;ZV:@9[A
PR*9^<.#[@N^&]Q.*8/(BF)V5@4G_\/QIKN %:^X()D23]@"<C8Z./38._CWO":P<
P'>1_RESB^*1\G;B..]'_$HV8H\Z?(PV(K9-A1M62O8L L&8 Q*Z]4!1]V3H,,L]:
PUU3UFN/+GS!M\1ZVF9<\-B 0"\@LR4>(6!!WO;#T.;/E"OWY%[Z/%'[SE52U_>%K
P+N3#']+RQ+6.<;:W\<%<(IMW$QW\."?60IE88[WSMK<6LP]!JI/F9NU0'MLXQHO?
PZT6@;4Q#?R3,E8SEME6Y%\\,B/$Y?@79/51&:K,[='8RNXT4:(&*XI2Y]G1O3?EL
P,KO]\88-3%FMK.EQL;9EWDI!"S.SRU4+?397]H."EY[C"R'5P1 I=O4]:,+#N])$
P.QVZM;D@5QWYWA;+W!"]M/H,UG%)(\5QN(? 33J-D1R!UVX!=Y#SJ$W#3J2"C02J
P1M+%N'+FB:A_]78\.%GCO3;^[\M[02'?=Z2%MN),VBJ/L/A"[_3Y(/C^\=.>[!I0
P>B#P&[=YMUS%2<*<X.&Z+S<.*?7=^M A@!C.OGA^L?Q26QB: >22>K23#D=#6:W>
PWB$6&O]E.$W:@ONT[OV"D'& Q1'>FK^N>))(_][7Q&-7U&_2QHH$ 2AUDANDGF<6
PK*")])^.7OU\F5-O':!@G=U-=IWN-!T@(/J\&XU)$(8L,>7)-8POJ42VB5JNXM].
PE>E3D@EJ*9&ZX3SZ0T@:L6HR X-Y/<['6?"YW)0$+FR#<VI4;&UZ.V)R6R&FUW4I
P>B-OC'%=A'QU*;1C7T:Q8:=Y-'T^J_%>&*B&G9ZP0"<%'R*R$^HTC>WJ0\)D\*T3
P8%ONS+?WCG6V95!:FJ=,>#S@YA3=(I@E1V%\1;GQ6GPO+J-$TM/ ^2IC(CWETN*T
P6CC^0]XA^P8"J4P8CD;)U]RHPJ_#1DND'I&:VLQ.MFD'4A\7WJKI"OUUZAO1BZ_E
PT8\+">HHX#(W=P1QW['0U$VPM]3KV.GHJ#OWUI NWKA=+,KF7GEAY.91YK8,_T"3
P9Z32<C)7Z@ ?G7GMXJ9?(Y\D4FDPR]YIA\?L"FJK&::Q3^E4:U1&UCRH."K]$%C*
PT ,@[L;JQ8QHG,50F?.#S+PC\KK?DT!Q>I+-5/76D,'2:5I[>;HIK1RSMO&ZU/";
P,8*;0UMKK3M4WZ5(L3@"V38%^O9I)K[C4_H>K!^F>[-!&2E+E_</+A( P/;I\(V+
PTVHX KF-P92O[WF"(*+:&%)0,SC^M^K/'G'F8$X(FTKT44$KTU%?A6?2)M^.=5 Q
P(-*]=EQV<<$T@2;&B5*+=$!_&AG=HG,IOT=*%0!4"$;!C][14L-)MY,'X.WL=R4>
PU#DOV9^W;) ;.'**]S//JQF-6ME:VNWO3\CL]17K[]<2!5@7F'8-PYLMRXL&RBPI
PGOK<V=?BC@3\$OE54Y!Z3/Q61/FKREK./3-ZG;R%ZBO3E?IQ]B6KL:I0WB4_6P!#
P6K>K%V%S[%@,;ON'[(ZR%1XY*<9Q*K"&;U%^$FB#0AR9-\7(US8@P] S!:/YU"GG
PFQQ=V]CCU7^K\6],EYJ);I-OD2/M(E=**@:AC0VW:1O4Y2]F5/6$_;K#U]HAQ%4 
PR,E#_L9H!7L%)%8-RXU$J"S^-/'=@%AY3&OO*D\0K;2PCN(]C9]P]F6IEZ+,W%PD
P/\[(689_S48]<&]X#J[=H@T5FY>_FQ6:@]S1Y73)/<+*;=K<=;T$T7TP4\]IB2O3
PB/4/%Q0<=@4G8;[,Q,-LU"ISE=S6XF^(Y9"I/4A=IZXNY2$*G9N9\V5Z^!077HGP
P7/U@T?6FW>G3HM-!.LTZNROE2HY^9Z%[,]AZOP'K7?D//14 *03TOK0J9PT&/I< 
P\0B@>_TLU;WG!C(T/K^GY#OU'6T%G3#P"66 P :[C;9>3F54^3WB. G'H$GI\3JB
P?]UA'M7]L4JZ\;_/$:;F\GES>^<M[8?.#I=C?P,N-<?>./KC9X0)3S\.)5]GDS3L
PZ_1G.D[@"TR*A-U[&@[?%\811^LBG7X\9#8(;$\#0-Y'=ZD*VM2UB:UHL7QM;$1E
PP.:PLP7[3OPRUG$\O\R'QY@4**#6TXN,\G O:K49RC_+]E*^C81_("O7M*V<(/S'
P;D'ESF7E92I7\Q,"R"A=#LM-RF7$?Y[+.]E?CO%K;67\Z%N<,=).CTW4Y1H(6 8L
P+&<:8V$A0F2H(/\GAQ=\'XIN23-02N9Z1$>F?\,V8B/.E=L?[>9.NA,.NA&6(G),
P8GE"'L;%X?$WEB^69HR0\4;2R<DJP$F.BMEUB9(?OA2:0'NU9=80!5YPZ&1/ +P$
PFJR0-D /J'"*]_@*YME.WT!MG0L+2(M&:X;C"$@4#D?$JUB%L7(V)S U:R""LI/5
P?Z*)5\+::HQ-430Q^-=(J7SL)2L=0;D"C^%%Q;UHX\<389Y0\>V5$$UM$Y?*:.*B
PIPY]I?1DC.XGIC;5QF[NOZ:E;F23=\MQIAV%>;2(5%?DKV,^]9DJ+V](8GZL.(9B
P&XJQ.KN#!7 'J)XAY."_2,'01 *F)ES(QKBGXK-S5O3-#DA8VQ%:C,'E2MU$1<VT
P[YF*O-C4I-]_3XF,?7/"C^ ,+ACX;W'U6WKO3:3+ZC-,MF(W3+.J=O=/I659J22J
PTXJS'5T[$52L.T@)B-]$R4%11^+5^/(9^RBUL!.:TL_;7?J,S6$?'YCDA6 .6.[U
PXW+8U.FVE(%DJF1%WF5>HW5QX3X3?/.UMQ?T1Q#VYF\X]/K[AV%FGYL;@6''%U#3
PLD'/7T)V9?;AAY0@_A]79:=PXO_MZ#B^E76!POEO<:-OZCGT@S*8\&SW#<8W?;@@
PCN=2'" 2J/+>_XJ) &PX%"$.Z]UX$ 5V!YF-%BA9)3=A;_II3,R^0]*H-,C98WE"
P5J P]SOSH 4G%J_F\J+"/XH*I0<HC@B F4@[[0>-(#+:?!KIS[2P?]!\V( ^O)%M
PT!)E_S[NC$?]UR$A(5NHEW$R)<!P44%*.S)]48EX@+G@8^MU[9AAKTB.<,*A,1WF
P5WK+**8M6Y"!,RY(11 VCETV]?W6J;72Y]UQ+H*::D/:W8^9URK2LQE=$D"IK79C
PJE(>B/4.&_1:C(G<.(HT K[.H>"D]:U7Y7W#6!>N>(9S-KR/8Q\.!=.HM$D%  NT
PPGT.'*YI<F5A3_S>Q.L3/=&.OKB(/C]IPY]85AI.I0); >ORPY_;^YX\+<OM'BZJ
P-J>.-OK> 8NW/Y0\_'9+]@_O=R7?ABJ?$,X5JC*SRW(V4L7_N =0)$LL*@S@!$MN
PI[APAF0!],6<Q89O-J4;OK0YR.(65U&GE7:X!^M1H;.NZ0_^KA,V?]F$&Q)TPIZ<
PPQ5("<K>+[0KI#:ZECI>9N38+M%)#U,FR?EMZ//)M-.]>/I@!,P" Z!/$MOZJR]=
PKP>1.!"^ 985>BNU@]!#$$6JV,\43^L3@MM4LL)%==X.8"G=_W;S/'7.%1V%%0+#
P3H1BMY_@3JXEGP<!G!'GFHBHB\1- G=P3XNFR>I>TQ\I2[P0:)FO_4 _=GZG0ZUN
P*)]^"%B5_GD ;C6(9W/K(N)/SF]C]5]+'A?_-$@;XU;!!&X;CIWJ1I&SBKXLZ=38
P'!^\L:!$/EUW&6?R_#J'/Q2(H*A5JUSKKH[F=+GGL.6%:NU;33&,1CV%+W4F\I!$
PN'029$Y>^)Y:M%_6XK;2(8C)O!K<':?E<[6WEPI1W0H^9#;9 94.&E4,]X<*5$&D
PZ-OFZ3&98IG,J<P*@F3:B.HQH\8[MI+G[JD!'(@0R7B'GWY0_A>#HUT<:- D@'UW
P98= 6*C2#*:Z+;<UY"YJO;O)#Q4G5'',>W=EY[.8(M.-X3@)"KN%-'Q@,C%Y4K]G
PZ80.%#4PH>&LY<H8^M=.AN78\9QV,.E>RC$^5G<[TNB9^I4EGM]\@S3;FQVP&*@C
P% W=?1=,,A$&W^.AMBI)#= &M#3LETJ44Z7&T;T; _">LRC=&AH_X89\"QX@V7<Z
P3*QUP2C0R/(!9R4WX7OX)3X^RL1BVL]R&)+O=TP\,]+W!GB)6-6]_^ZSWE2<ZM:/
P$+[L0T>/PCI\VH1$&*1 ]?\ ]LS5<R\FKW[YH'9(JP7*NU VJ^T!D.S7BBW1SC(I
PM)S8I?;90D&:Q1;:E9:%=)6EIGEU'47]YU/&@*968HO8)%S*T6+D7IHC7^>,9YU_
P/H?8J +/S)70 UR+3Q3(6QJ*Z2S*2=[1&T-U) S90J"PA/[,3M$-Z+1F7224>1GU
P8&/MXW;GP6]B9F%H01HBA(TY#>0_4>5[)<M2NW/SCOSK8W=&X:%1[UE@G9O\DS@M
P]+1=KQ6G"]!@'O/S5L-DJX"G_@O#P?SM_._4/Q 8S7YA3K-2JV,+8&=2+:X.H#!]
PQ2/$B7\7-GGB9N<H:N(1-()I0:&K/9VW3?(\+Z8@*S3=%M7/*Z$7_F0,LW?F.8BD
PU;6G85OSBYV\^13(Z.SK\&P#Y6(=,KTDQ.,+M3C@3@2/D@"INM#'?:2Z.,59*N,D
PVABTFZ!^W]WDAZOVBU#R!O*J:7^=M5-V8\%3[<S])KA"!]980P36;YODW\^O%K'W
P)CVVX#IBK@[W,3D%BU94PNOXUM0?[]]E<57V'.Y) _UT_;($=_A%_I31:.*63+>&
PNY?<P23SP<.08N9J[O[UP.^NPWZV8./4J'??&I;A,Q(R!Q;7FZ],7 NI/;M(5,:\
PI^JU+EL<]1LFE<N_G1FCNN.B58L<(T21/6T>VU@2\SS!>/=;(WZ+.=>^D>UZ@WEV
PK L0(0L@-4/]0-EINDR M4;%K5>SJD715>H^UHN%3U9I_BC(*9+VH! UW1>[_#NU
P@#OXS4QOV_-Z&WZJI&\68F?#25<SJ?$EPCB1ZDUX^WGR&%BYYL75@Q[3\:W8ZY#2
P.^V%?3O,;J%HC/J&>Z+# 8U,QL(.>VQYN(DL#HMK-7YG ]N(4;"0RQ^V'V9L=LAR
P%LX,)79 !P '4H'$='W<5)S.K6-6>:$##>ED+8JW15?^/+38S_7T?>:HX5B8)Q3@
P4_3;0*\B.:CJ07&B-+IVB2'M3OK9F"_7;Y#8UV>1J5BZ4NK[00EOMCVZF;;8JVU0
P7;L10:/=TQ+">)-O.V?RQ%F"]8O(^_59<%6VLE==.Q'-HGN"PJ^S]%RF\\Y+M884
PX3)N[C(6.X8^61^BK<(+W12GG:E?A5IWN+T=D5RQ=>MZZF)OIB\"*UVB9GR$NS5*
P[A;*]%"46Z/R!XAC&&FF49>Q5SZ#>T/BKQ7"F.@E^N4-[<]?+G2#D?^:PHN;H"0(
P._[A_Z4"RP>59ML Z>U<TW3HWMA7'E2 "K2VMKM1W%?]NY&$CW>'$U-_V=,:4(8;
P$\QM=J766<IQ;E*LF_HQS]C]1T>9*NO38DU:2E*^HAY#-"8N YKGJ..Y--[ F*<#
P66C YE&^B:TKGDQ3?IO_:,EV'WSEX D;3)0+AP74*R6XJ_2_(AF$R=JJJ;LSFZ3<
PJ#H+ =('=_Q,1-H5(J"("##N"#D1Z,T!FSGF[2];545P Z>%S<4'G*AC$U=4426X
P# ]-I(RW44((3I^2*+Y,-M<AX/L_!!@' %0@806&5F2<1J^0A1TP$2=3O]'B)[SU
P"HV_,/-7.]V"@>J4_G3K.\*Q5CC JA:!$'^X\W/&%Y'=/[68TR_/[0S3<\>S93%#
P*TPKY\N&524*A/%//_UPXNKQOK6'@&7$DOU<@>,YZ \YIMPF<1E!,"=-]W?IGO:)
P,Z-3G=4]O'WC35'DP#?.B5O>_U4"$;1Y8CTE8/,@RGJXL=QY%+B'*8-<L;GTU*9?
P0E.N":"[3Q)OH_R)E<@TI?$AEH'DQMITQ6M3%^(7:,=;NVJ,R[@G&_;0@MN2,_*V
PA4=R?ZX76G,NFZ>CC:]15Y 8$XP'Q.\>3+%9WG#F<?,!$<@*LAZ.+=45\=:;;6>/
PVIL:QD$2]>BVV:$]G,YC0P(03P^,YJC-UU<]:\&U-=Q%*ME H A=59<*?*N?*733
P3 6(W4A8BJRF_'#-\?Q<A:0'OS2!CQ,&]D*>:]K/0K6_6F5G$B]!AZVSL<OU XC:
P>P,-0=?A/?H7BU$-^7G<-JC!U*3)49,!)J$-JI?1)$V67X;HQ_";/N+U4=G[C/X)
P]M3 @AK+(\Q),"XP+,&0X9)Q@-OJL%IW$(5[@-&=OV?"!.%'R^*QH<^G:D-M.BF&
P:+)\2+SC8E))$J 3=>U8_))!V$-?+YI*7#J/E,3I,T_HQ*@)N8N$>_T>=!M2W&2 
PCM<U/WG7^$9&>8G_/Y2@HNLT:O+Y^9MQ9]&*3S]L8%G%/'P66"3=NF.)O^0V_CC&
P&5S:(&Y=,U40<!9T++2H1!"E5CI32TU4 8^F\[H=MM(3')X=X+#8N=TQO[N@]EL/
P.B<R@Q&4TRT1>[0Q7),A*T5@SF?;LG_.\#O5U5-@US_Y)/AME(-AS3:"K^D1;N%W
PIP6Z;)*1#^I=9!R*Y EQ'*);.X.FO<+A"QWCBA\</;A<1?F K+\I:-OMSA_\XIC0
P%?GT<[TC2;ETY/:ZE#&W^##_IS-G(8V64H4.RZ@_LT'OHJ,8'T+_BDM8@);RRJT?
PF9.OI,,^_#DEVN.PE?(J-PJL^*MY.!J<+[W3(%CF8O._GZNZED/COF6RE-AE+T5]
P*SW&X2+D4]<VHG_D3+_9\%MQ4AO)M0(]OYM>]4F2#LW6V*23;%XGVY6K>FSZL[+ 
P4<[.W)&(H1$'<WD8:IK]GX.$3V1@EQ#&R3D:V_'0U 301]2^B@_),UV[Q3&^YRUF
PG/4$M) 8_@L!S:OAS*/N\_PC2=(!RQ>B8G)O0XFL!X7ZU]C_MMH0A A<FR[PN<!)
PRZA@;V$KTL-H#)@OI,DGX2'[J.S/9&TS/>>D8RL?9KN(CZW1/M*"%F?-6._LQZ<M
P.%!Y\TJF+:1B :*D7J=H;VH@ )9>-G)% [CS85_H.[^GAU1,N_J6A8Y% U#'US\>
PW4*$>_1,:T5R3(3@$0^PJUV<_J><KOM!3 FJ7-T/]^FV:,2?PJ'/[G9O3:JSO*E9
P0[ZGION_$_A&0WX:]KN^-$Y5^3#JR<U.U!:51P=E&O\<?B?7(_V&0,/E^<+>:$V4
PV?3[%,T<^V',OGLGKW0! !!"L2)M5C-3UF3G7F5M.(+UF7&!%A8%.K#G:  >0"P;
P0%J;1+GD5GA[LQ/^]Z'Y<(#5XNGZ5YUJ'-E6'4RPDNTMKST)UXEH;AI'4T#91V:.
PX'E8?&2]-\Z?9%("ME;%YL.,F*?]<9GN\/OF\T_6DH?\;-^;M!V>/9I(GMNO+/@+
PJ11LQL$_0N)$G&$L1:R$OR5D+SKH4Q^MP\0)"16>BOO>)I%;F3"TV7$*TS++8,(]
P]/0*R[23ASWL SAU.-OJ78%-8:VFMT.3%<,P>;,64E#+1:QOJI=!,3%7*D, 1Y I
PZ A6N)) 2S)+N"C!7[I+<8#'5OM&7,Y$"[4W@H"=XN>@?!0ALOBX?Z4YUIW13>U]
PA!EMKGA7/')Q\L4RO!ZE2$>;N@Z(FY/EZ\18B$-9.*0CEPV/-4T=ULO&2/" 3MT7
P_:_8A/!&=0HLY\V5@!/8Y^I.O/4#%DNPE7O*!&BR)4HRE@56$*Q#&0DTTUNB;%S0
P<U-NVS $Q:K$&3R7V=\:Z;/)[M(X2Q6,5%2TPH@__F(A/.$K2808*[G17Y#CEV7<
PI2U<Z+17^YO8.,;6>@V-GQI@Q&5YJ=['S_F;DMR&-F VOTH1TA[*N41T8%;VX!=X
P0*>]U"YZ=K8]I'RSZJZ:TQOWIUD=(^'5%!PJP;$TH1>Q#N.->8!ENYEW-C? ?!R^
PU((%2=T/PZ6M58!LKT;BV[5/(F2'Q8%E)?D^<GPA^586 &9Z\DJ?%;:/_Q.;; N_
PK0+*[-ID?.U=!FI;W@4^'> 91/I)/GEER\ 6X576^^0T<33.T'%J6X19>-.P/+C7
P\! B:->?F$4EA0S:$?L10U2 B'402:)+:Q5E[CI=?6SJZ&YFSA/VQ@R/(R.,ZA"8
P?,C2[;=LJS&R'? 8WSL7H9/1,HG.UK,[8%J6?\'LS1QI01)+@<*#MUDC=@"RKL;2
P=Z?88BPOD:6>^-JW.33:@071GF=I;XY!PJ")CH(I"B)(^/5NEL=1&MSM\D)1ACK%
P<4\]S!6- G;35?J']6';G1P&L&2L8TQUZ"9DO0Y<* W V,G\07F ']V_V3KC03>W
P>N20^><G[;#&L_X\Y/2F[=>)/A8C8F_U%- 3C$" V7K1VXX4!9$H3(!HNI&NI?4 
P;F=0H*AE>Q.OH"_?F3+4KWDH+U'[2$6UT4@%-#ZYQA YLV1NRN^WT2J YD/R$,E!
PKM&T3E\*^YS6>Q?!IVW2;_HW:0G#,_ORE,;/_6,W*/IF4+TOC9])ZKH_@,*CM?M2
P>,WO[U;KDNCFGJTX8(^9"])TQWQQ;SKIC+8@ KF3^D<A+B6!'0UI'T=2"22[M". 
PAKMS,TF]L>-<%D856>?#=16YZ12>#2R!;!.+#_[<<X52."_TS5P:%#@!'X^$Q"8N
PP;]'+,T0VZ.(YH\"0C*B4)^117@ @\@$2OSF=P.H516ZRJKO"[":HS8S_H;W*"*_
P9X.)8'8E 3*MLZ""5 H8&)<+B.8=,-B*J=#S39 =TLA=^5*?%>$!B+</O!H4H61G
P>JY=Z?PV8\/15@%(U B-)D%GESYE #)E/(@'59+BX_V_HP&VZ3L7JPA&].1\?APK
PTODU*\'2'S0 '2XPQ8R%RY=*<?AD5=+R77ZAA'??O1B=@<2PR<!Z3(5B'PV9#%M+
PM.$QUI9;0R%GZEW@ES3C&S_PQDU%@.78](K!9?DFYY)!5:\".7CV/J^@E:*\T0I$
P9$JU_G!:)QDI7UF--B.FN99:'<C>=V%*WX#$G\A#:>G.5),;_F=&@(I3CJ$BE[M[
PB2*-CY6'403!.[V(6_2#(GN-OQTG>JGTP^CC<#7S2A@EW%7=EL>@,Z:N,'<:(?K)
PV+.0/VLH4=,K-6XP=*\*7S1;&=]9RK(_W-SQ<Y82@9]7K(>IU4TW@=3A\%5P WTT
P D52Z=T6?*NXL<K\Q!S^]+&S3=*%/55;384Z3O*.PM!!U$#5YMQ2??@Z(O[6'MP"
PF/??B#Q,]GSI2E?AZ1%BZN=V;-J\CX7.K<%F;O>-K&$?VCDQ0>DWXV.?.E)F1D!C
P22$?ZL%9^WO^I']^KM?9]XH?B$!<K9D# 8FBLZ&54V[;L["VVR^+"#+RF<SV9:<1
P,9*"2S;XJO>@IMG1%)Z\0AGY$);/M0B1!T".C'@F0[[8:AZ+X=Q)3K+;+G[:G/XO
P7(9$19])?,U:G*46ME&18+76T*J\"E?5<!T!KROW*AVDN34R=IKW)>M<;/%A& RY
P"]SC*M6;>J;4O8QWOKG^U)0X:#)6@(=C3-2/FYJ'K2]1-4T^6A3A&7?Q^ZA!-E:\
PW>_?%DNR+4;:(HT_L:9UWBTBT]90R34QMM]C&G;C("2E0'C,++,!ZIF--6IJ%AJ$
PD/CN[/89K5,F:-#]9A5  Z3;J=6A;(>285< 7X:=?A%U Y;9R%S3WQ:ND74@7+!)
PM@N?-]M(0<5![O%</<0>CW$8@MNM-J1]W(UGZ=C0J:AKCSFJJMG/#16IJ!24IF2V
P/5\>1<TM-CYR$K,$-D4O7>8Z8C@]XS^5-OJG?XMPJ\?%OB(.%]'R#9"L>L7(A1&9
P\./WXFQ#&=$\R/I6SF(WMFXDM.ZS6N+"W_D%W=7$J)F)LP['U["O:3+U[(A?QG/&
PT"O[:W0*1GPP](=2-*VZ#RKHGTVVGW'KT3OO\FUH,Z0:64$! 5VPH.K4L2F.W9RW
P\_8PEB'F_4$NB;@-F]O[4-F'?U,P7!3*9^+4P3^.4E=O%U._$'=VD)5*>)1N]X'-
P'N)0"*!A&'$G4%C==?.)YT5ZK0]CL?&J5/)EJ/&<>.3(XEX9=7N[EX9F]!X<YPWA
P2U[RC3%9#%%1K(3N!OU.,B/Z7JEM3,*L$C.?ZV%W_Q:$H+$J_)RU\EZ"@8W,E:QB
PV'O>R3A*"-.?$^VX//KG>8BNA9[-Z:CCQANN9SKAZ@"3FG>R+V;!LG)2-<]::@;2
PZ6!_9U-_VN#YK=FTPCD5[QLNP&GD[_#-[S.KD;;C)L[1H(QOM@=GI()3P<1*H\'R
PEN?)%JG8,<LB=IEJDA,,WD4RX9MS&XP$0X&9*<@?<M;P"/+-17M>#;=5@694=N/'
P$.B&'3<S"]^Q"!O7.X\=^N-Z;Q*Q=@:%86I\3H2H431V/:=D!E&\G[+T%/9'EH[8
PR<^OB\3!D;,G##!9$DAX2XKO$*J;BKT3Q#'6]ST5XF:?;@TEY@R.RE$1XT^,1QZC
PBJNH2^.\14C-H^7/\X^9A$[ 6'/DDLG-1%!2C"JE$EU;I%5!M"9T=6?QC[F^Q"?&
P&, W.SOS6J(]OM/1X#5'I=#B@<9;3\PF.@-9*6/J7Y4^M Q;_4,"F@)0LGI=\QF+
PCP@_/(DO<Q'F +@.:W/+&A^C?T??L^ZOHB'9:DOPI"I(6 D"O$7^X4*FI;<SWS)9
P%.GX^D"B&X*MG'N>2[]]16ZN@SRLXZV._+%5073:ZF#M+MKXXQ/NA!CI^$5(Z%RT
P+I<0L!LM\XCF-Y2(!1>)@A+U\8268P@"LUB#?_7JG>A<@9 B8FH#]7[-UT@WU@P;
PSYI\-T!8(/)8C*,6E@>L+>_G/@%94T"V!@.(O/'E5ZI_G#4=I]CI_:J#NTW/]5:>
P;:7K9&O@"D)M<[P^3T23\INP8QB'EK@A32Y?8R._6>+*CKTO?AD_41/L7SZXD,_3
PC] 'NB=N1ZKV=AL0EYZ%ZT/;_5&55J24VL8@;M"ZI.D ,<\-6%MW?:_%H#TAWV*,
P8HP%:7P#&@CY-/=M_'@5#,UKMLKTQ:YBCB!QLFQG1FI,J6EZMK3F;WIB<=YXH#Z0
P(ND_/:>T:':IWUH"^GUP->] !T-ID3FD>Y\L8 '25I5-K0HQF$YB[54+46N^%S(]
P9L0[VFOL]L5RDGAL0T]; @>^;)]I2H_+L(HP%]H6$7A0 1RGA6Q*F'K^$.&&<-?E
P8!VH#1T?895L7++,.Z=:&/7ON_R)ES QME#DWAKK!3YX9O ?*LH_A0I?MYMPBX%!
PG-W'WDJ4V/] =H7ES>L/2,)4B=A@//I=[T9\0QR3L%4=;(-\O*:C<H9&]3UJA)PP
PRK<H>T.@T8?0) -U>E4@H<>;*<K0=#,^V,>+J=CL!Z;-);?J7D)#;R[!H'N10&<7
P,I1R!#W1<X6<DL:X223[X#TQBO+W#:-=)(?UU1/ZOO V[M,5]3GG0E >_%_>" W+
PKV92N",!+5JQ@Z3.&&T^@4J?=C'P GC%_I2HS]R,"AVC&^>S?[0I2&9N97VNU6(\
P;1;@]$QK$4]W4NNM?2 W./R6E]5ARC2**P0BU/U_#:J\HL604_(^[]T\]=.CU^23
P>OV'J;B7?NWQ%/B8WP>%.IU^B3:*;^O&3WL?/_JLWP\=^%A.N](?/Y]0K4)@?Q)T
P8<$RP4FV;ZR^>/IMR<6GU:R2:4NI*H+M0.19=?'<+V!02+5I269(LFP3F>W<5^!@
P<0V6Q]U."^A6X1%TPE #!A6E<9:50$JURS%UO%WK*51>%^_)X<1P&LQ-=&FE/JHI
PMDF;:"4ZG,Z(KHY1S&,?7%24NIP$7#B3Z4(:#>;_+[F]]M.UV;DAP17.Z>V7')**
PT,//**='8J(I12'0U58/-*%1_BRB0WP;9@N-!!#V+[^ZHLYJGBI(,3!V3>JWB#&L
P2@+EUI>M&Q<UI)K]%/QAPE-W=! .F%'V J/+.@"W;B=#RQ_S*KJX13<MOQGQ$<S>
PF;SW<':TY!HH!64>A%(JUZB CK\M?:1T?5FWA-E$4L,RFZZQGZX=6+;)LI8!>=$1
P5;J=5? 6N'R)?!J:YG>M",<FUY,4!C1-4%IY;5]ORI="%TP.+;PO#[, 9ZR&/QJ)
P_=HIZQ3Z[XB(H%:=I^E96S)YQM1=-4JO)KJYB1BSG_OSA])#MFJ,7F1_!]82MW8D
PCYS=,R?L!VA42>?U"'7-H^'GE;!_J 'U%E$;UIH#9629#X=B^YBSAQ=>9Q9G;/)A
P5B-R@)5AG4JZHXMYN]/ Y&_%,UFD\/.]EK2Y9!CLZ;0)0-6K#(B/;N^'/[G>P@[U
P.IGT'XV1>:08;7Z"@LM=;GTJD(I2&?6+]$Q('GJM6#2_O66A$5QJ$$N=?+0IREY 
P+V?D,!T9B*P<Q[=T1;LU=@P[7^0%#G  L0^J+B_E>IF4U*K3!ZV>!1\O_K;')NG[
P&F,T.?YZ8<>D;:UEVII-U,$LPRYW:'^X0^O&;KW0!QK0@'V#VW+??![)X;IDH=ST
PI<%1N#W?P&?,O-^9)^A'J0T1BOLV)MK94K;_#B78F-Z[16+L=X;;ES_?[IFMO*)B
PJ]0ARO^<,RD-^4NM31N\I2U.P\%&D/!Q7RUA9/-(E,SM5A^.: C\B(NFQ'S2Y6CY
PCIHX:L<J^V<J&9F[F\3560.T"NT4'X(2V7'YSBD47^/J885FY%R'O9A4&[\IB;>X
P/$$?1$G/AIZ 2W_EDXFP>.,!)XM<L!DEB4<**N?5[S\UU2H0T''<[1ACT'\A/N5:
PDH:'N2,=O?VC6 "DN*Y%G)I%?I1_.?HI1FX]N;]/OD(K61QMFKL\"*%@\_@?Q^J8
PB F>&G_*O[/9885$^0F>O '\@2Z$JO(EE5Y2 8%Y>PJG*M1&$X:P@0R)9)'30GU-
PTHQE.7^/8LOH()6.)!DV-MJ_.H753.5J/![W E>,]"2M:95TI4^-M/>4]9<RTM:M
P9:[DMO-.V5 52 PBF4[0@WQ'&ZC<@7K\S))8Q:Q!C#>_&ER^YKW,NP>$Z;9H$5!3
P:\&*[E'2V-//+29Q+.Q7F//W+R&99OX"B3M/.U63+3IL_6 D/J8>9%#RZM*2472A
P_&JBMU8M^;9/X@T\S&D#N.XR8^P=_=#%,T(\KI?]#6U0$J#H'0?HR$8[T%<D$SMO
PLO]%@WP$/B&L"2"BT4EF^<0)8G4CBKN-U)QA2>BZP0)W$@%8\)ZB8;OM$;HX 9M=
P$"AK3C6Q1B@$-/J&I*,X?B>RR775Z_A#9ZA2<#54LS3,T6]?5&^VYY]NMU!J25@6
P#H35@2]U(?#B%&.+9U&N57ZG>OR$H]O_-ZP!R%^(/<P)5<"#CY]]H'V@6->Q7 DU
P*$ZNNW;CT9WJ7$72(44R*  &/78*C%@QP!]4['1I\_$3FG$&#M!@U!#2J=)(/)W(
P>%OWQD7\->WM\1FF=O6N:! W:^^ ';VS6*Q..K'YAZ9VG]:=SQ>6EE)!=Y;L'DED
PPMVHO^6Q3:@>U6?C?3! +BXKG%YZ]S0HE1?M:;W%<L:,**G?M8/>;Y0YNJM>4,),
PE@? X7&)!1,B^MVW^=Y"1DC+ARDGV+:005;\Y![^GL=ECK7JAF2H&>F@:T=K-)F$
P[HHMBX\")TX T7P6=1UJ8_OBR0'%O>CED_P?S)]65J$\BG" =_LSEY=CZLX]$<Q0
PN'EO$)*38<E0\2M6+@WN"M[XJ+LU[-*EF(Z.B;JQ[')N,14(E6'_9$^J^RFDB[5S
PIHBH:#8;%\),N0\1T:<$O+33WXJWN3^^FP*'%BG=@ R6HLMX"*LS6SNM77<^YX@2
P#KM2)$7D2TPS,([WH--[(?1G0^]8?70&@W1P6!^>7$$-0BCE15 *<YFWTI9]S2RZ
P@G%I,/'C+H!!I=CBP9,BKR7FV'XSF2T<&?/A.1]LHO;0HJ.)3U#8.M"<X^B S9O_
P/L+_]CA@;)5Q;9KVWK71202]EGXVG359>D@\O2"SG][PBAN]F@?+Z2.\58S?+6<3
P_8BKA=C7DFQR@P/YF@8$^+$XSO\^<5"7;,/FVWZ&U_Q&NT>B:O[DS,B4'KW#9EIX
P>M^0"0JUP\DMZY'$?!(7%!/>?[I>2%'ORQ"O'+=I7V/B.7JGX$T*_)N1F/%IK26;
P/AMW=*%=$WEJ'QJ# @,ROF+*7*V,Z9?HV'1:G=$.E*%H"8KVBS*VX3C7?"=>V$G=
P\!VLJ,_U\[FJE,=$-:T%+<R+?U93!,9</D. *@&$FB&V:\ 6Y-D<MYHC'Z-.L?&-
PBV!VXVFYQF'Y$D""NF'@,;>.8&";1 'L)6)F2@<")$N/R0V_R27B#X5RQ -XN[!+
PJT<UP=)%*\=Y0.JRM-TP702 L>JA""<NCV_R), M5L;8,<]B@4OK;;Q>J%X9_<5;
P1HL&%C3W;LG=O"*T3KG?+G6U<_>I,K_-&I3L%7S7[28>I">=S?\E2W4ARUTQ>CAT
P9."R^;P$M,P\^0Y*\]3Z[$UM>9.#-P%GR*:H+J?7*L:=:Q<&JVF>(KOS<4HN>?#8
PV->1$]WNYGWH/WL#1Z*VK2,#O&NA*V'Z>TF-Y##UZYW<15WO.U):&:4]U?WRJI&O
PK>%;*[+2UKYJFZ!]RE8WD*G>W__@M():HD.*@J=7JRR7 67]%$ 5-9 =ZXSX8(ZB
P5=K('9IOCW\YAJ O[5FB)ZM74DF$P#:7T: \-W)]D?6*6N*XA8ZZM30H0)N1(>\A
P]U1&!Q-9:6!CV6RP@P4D_E:GBWJ@@D@_4 YHHS/%A7%2LC@I2>MF?A'K:OH)G(@"
P,.!H->[NT6&"2QM&;E&HCOAN#0P4S=J%K9LO/XF.<;'^ O5]=NZ#U)L5P(L5:*G^
P+5GY,]S08GN=]M!018'1CK$,=LO#^KH:-!4+J7 .05_7A#QU2@ S)?56J8DJ0^XZ
P#PU2H\9T=( GL P(F^O:NA-DTK%!*^L]!AXZ Z#TQHWGRE:O<C1Y*ON%![!X@,?I
P[EK?X$G64^'(V@9&JJX!>73% 0@8KN&W7&_@NP BCO</9Y:]NRG?>V@& GU'Y#N3
P.54#+5%-/C_<_, 5"TGG%LV$,_$#+$\I.HY]3]%:SQ==77_NT54DJXP>V* ,N )O
PNI\R+-#0XR5R4Z2*[YXIO[=/+'G&RJ\R9 G_TD3UO'O,*KHQMOQG"PJE4Q?IIO)\
P6,Q)LL9-.FE]<K].S!PDPY.\-=[XJ_&\B#KUZQQ627\U *P2>36'95V9HPE^03XG
P@X;C2?/0^Z>6X:8"P9MUVE_RS/JT4UZ8S1ZCI8B2'=+8IK*Z\)U5+3-F[#9%[6S@
PHA>#C-F1S'G3LEI@:C74I]_DZ5YJI&TL)$TTNL9HDP@V9NV[LG9Y^X]9AT1D8-7F
P"5&0=K>L'WQ81%TN2RZI1HJ\A#R/56_?F*/63533=NA[7&ZX63)B_"'5QA>$Z243
PXL#*_-*<WW-#4WH26N@?;/!LOFJL*].%V5P]6E\?I0>*J!)]N=<>>]Z7)DK9(3S/
P=,I%@$$A76J>WH41CY&C,PD*9:J[3!_8?-ZMY2[1?6D,$70>K/=J ^7/N+%ECY-.
P?U5$<&?()\IO64O/H@8?L"1IC>D!W!_J5F4J%IB$\(55WMKCB.)4*R!EO*T,LANT
PF,NP%&:G"(=E'3'-/-<"8P,365SFU+J"40=M*1ECJ$Z, >TG;.=L3R\[0M-7+W/J
P\#GU?C/WLH=^97([:P&]#2U X/%#[?NM+R_%U39$9WI/T4O$A)ICA,D68>)M9/'(
PN@DB.@A_5#*M+Y/Q'#/C@MMQ,06NOA8O!2-I&S61NN-2LG38]GY5KSAXIE8\2Z,'
PD5PM=>QH!1^O.%DH5@F19X-AQ6SYY46'\:6BW(J>UZW+K^3B/ ;6LH;(9S;EBU<B
P 7CSE_\:KSF>^ ^:_&^4NH< $]^;?!E!!HAL4JE=N,R(==L6G7AS[8,,HDH<:8(T
P"/PV1-8*&QV"GN*<2+HE=>2R(P%O:>1KG;3KAV$ZL8$U7$\@0%%186(EI9.R!Q$Y
P# V2:Q2K$PU(H/,CC,A(:&O?LGX%KVA>'DFM*51J&I("^U>.W?7 =>,M)T5;$-'J
P1EY)S5BX2T*MIEYY!/)E(0)ZJ!"_>O\BI/:>B+OFU?M3$\&9O]RCJ0]9255UD;EF
P''987<QDVTU^[ED;!$N.^L>R)&9/ PJ]3V6+PW-SKERCW>4?X8*PM;\UZQ!\NLC)
P%.4TH&;8@OL#,9:;!V$ _Z^#<8P'Q<EZ!WF.#2D& 06%$C)2M_S+V)_C:\MM<]58
P4OX *DD&Q717;DIX9B-(A@GL$9'9#S&ETG)<!&<L%'KDP=#&N+8GE.FACG8R\+YN
PL\C#!(Q&YFT$-<-J-K$*1[F,3=D7/:XZUBCWVS?X^*LR:,JZPU<UJ+8NRBZ7I?CI
P%L%BR_W6Y;1-6O6&Y:WY2M[-Z+:+&W-MD3)%)B -1G MRWB'$7/,U4ASKCX';X&"
P/VE.P ^J1MQ\Q/W<CI3GL3U-K^ WULHH&NK1+ND=Z<F)_XI_;;&=8Q;)4%+K)A\>
PAR\ALC+YHCZ<WMH?,S70@M(5TB/LH,RID=CC46XY#P3T905X8K1228+'U'>7#5$K
P\IAV<"^!&W;3[.Z-U::.,-)1M?T$9[*X:7V32S.(<!O=&Z3XY-7KH^.:'1\3Y=_;
PN;I)-Q1RX':3G\_F&($?TZ3)RW7RS-")S"N-;@X=3]BREIJ:ZU!Q1_1$2:JNZC% 
P5P1#>B3;9X82%>J ?\JK#EN?$P"2]35I>?D\2D$@8[%'_1&#,/AF?[FLQ'-.X@EI
P$ 5_-S!)L1ACPB-J(!^A/-E9<\UBBL+;\XXY[='4WV<<LS[Y:Q#=9F/9.6Q1CI%H
PKMK2L<"P5<3)"ENCC"9DA4UJL8\Q\/+N(M?<7*9)N#=$,R^&(\72H[]LJ('>H<SD
P,H!KR"V7]8?/,$WK[+0Z#$CR$%&F#;M/* 3I1!F8M(::"[=E7;*AYJX\1"\:]V:]
P #VMEE;3?>WCWVKD[2I!W>AS\U=7E\9X7P\>:(#(9Z@7=,R0;#$E:#:4-9]:9@72
PI1![:XO,$O)F:@DZ&DVPO*(5MI_XL32Q';X3-0M<I\)$?<ILY3-J@=W8D68;?K@'
P0K\<%.0V/=%\O+0K>[.GAO[CR^):5*O";IKEGRG:^,KRM9ZU+3 MZ/LHQPT>8B/(
P[;4U1GS;FA!2&&0M75[#"B;\P3#4LI;H=,3^::"Q?L,G.N"!E!*M\URU4%MN$K/T
P^!/ST2E@>2DM.+HW6"HG6QCZXR#H-CM?.>W31 K12+/E&ZY/"><G7SZC1PUI']/;
P.EVP\_HOI-6V>PQ8+>U8\JA3FE=\D/[53^H3\@OG4'":B*:[G?GZ\. I^3$>-"0B
PK:5$Q%G)BDNS/AG%2.+@>ZT:H78_+/HRT/A(C5:MH37I9-,-SQ_EMEY5-13&\MYU
P3C$\;SYW"%T18CH*8["]ZNMATY5H![H>;CQER!4R07^X1.GIJ1)L+/D.M/O;%CH#
P$SHTC'VY7C&:$">BC5V\+0)CA:;XNT8MQ$MN9$G,S+9]>@A#<6@_V8;^(F'9)!.V
PZ%</.7CQ*#M!WJ%MF]G;^'G+!3WTZ-XC#5., ^)]@&@$FVF&>--P>UND8:K>3G\<
PM,8(D4)39R2^DZ:^^_TWDC'N#G1^':+40N3,]:W6:TW&B&8F!=YC]-%==@M_*.#Q
PG6IZY9E9SR3M2:R6*HNEUH$RU[#WZJKN6 X,25%'!!#(R2*HSO7P^870=$ZS/D6:
P!_IK?<7HLE?X*F=<DDNW7K5O602^9F3$JC7$YM5<!@':29_[%]J[=U/*%,N0/J-6
P6TU PD%=_.'T^;=HWW;G2>"P%=&7!C8U;HE]^<<BL8S0)?=',=>JY-$7AG8T/1(U
PX)FBH8%6^>/*H'8>L=".1E<IT^55Z$(>[]$H%4D\*P(\J/P2OM-4W/";&D*I?C:Y
P-,=/GJJH!(HD$0JCVEJ#F /=9W;#IN896RGUS9!= 'VR:65C\/'5BDB"O3,\CQ+N
P@119[EO"$S*^Z IX!EQ]@5U(M^&YC%=&@Q*+17_=8,\,??;N.RM; +9.Z)P'//7I
P1W6^?W>@U.T5M2Y,#4@9CUA^SN/DE82/"B*X#&2]VSR:4Q7?)@?9#4:RB?BI!COX
PWL! #6BH\A7K^WI2FJ?P>A8LEZE<_XZK3\D@*JIS(&)I?E[.6[ASPM!]>JE<\#YQ
P"6;LL Q?8F]:6G[8'AH7PL0#$09W49H+X;> ;\E6K RN NI )@H4QG*'1@8<M UT
P,0H-=Q/7/!<J] 6N2%5+\J6)@0E6:V4.YXVUZWE3>&AT8F+*O-K@?=H(Y^E$!Y%\
P[69\E6Q9/SW3:PSS0*J'H/^BQBM^C]U&'7M89E[$5#OD#OAZ*,6.TP0S;ZX@M#Y2
PK7M'Q)8[)IJPH7)HK>H\VPQW_-<DA%!SZT!^Q5Z>F6K>1HA85 =VNV5#:_!&KNIB
PX+QY#W<E(B@[2E#R_HAYTF>,4Q](]]E;8$?['UL&)>"T0EO(6QF6I"A<ME0V+(?Y
P]M 5$Q[Q 0KA=AY!&@2?$QF\U2T\':F"4W[9$Y=^K;53OZ"19(&A% /R/\)<@>@C
PW$SDMMFV#0XC)RGM9IC"CL?^4X5I@+T!J@,TW V1B)8SPN7NZ[K%5N6J2?>=MG5Q
P=[5[13F\)BEU?S_N\SMJ*>S17U+B_[8<L\I_96-L"'TY2\W(EY>@_;+:FQM./>D7
PV9C?ZO 8@3ZTWEUNGU#(R?\(^L]:J$<OZ**/RM@P77@.S".XUH17?@@6G781<=Y1
P=5:#S4D%VIJ_5HP43RP[B0E$!B\\(H<*F(5M5T8?20Z$[[1=;]AGH(6<DDMQPA@%
P'\@ZTVK5?CU-0R22VQ7X<ZVV3Z_Q50F(FXX^).#;8T2+'9G\OC,2;&AGG[W<HCFF
P?EV$LX75Y2[YN'-IELOV3> 1/S7RT@]VC2@1.T+,7H<B4R6D?*:AL90X2?'H+]V?
P8G4,P'>G=X5L0[+/V7)L=16_!XYTK<9]>R_9.98\6\,6R\6)V"'!5KJX(9(2WUG?
PC,E440S(*&UC>)+Q1N1/,Y/_D#X!J1ZU,?JXPZF9WA=P,V+WIMBF.83D=$PQ5)/(
P_A[9Q4E'M&AFMC!3V?/?0I'DS9*)5$*24L+(%O%%H&"EP*82,",99!?UYOA"AR?9
P)Z3UPQ65]\FX%)L6JG06]!O')R5OJ*/VDH"&R-J&DOV*;'&KO)PVI =*K++J[2FZ
P7+J9QG%W^,!;I? #D@Q%)(E[=]+?<<S[7=>PZC5ROIKH*>^@'[14O""-S)("CX+A
P??VA!RZRB28JGCR6U6CWT7*<R1HN&H^<3OV^7A&:QF_#F#341QWQ#:/WH$;GX@"6
PSVV[VE!T^ZO(6U]W&\_,0;+WOUT9FFRXYXZHO5U*NLE,[IZ9WXOZH-[%RY7=LI'#
PDBDC@%N/Q<L<JV]ASDQA]:XS' KWHV,\Y)3-J-+BD$F=IILR?_D));2CBN#8FNK@
PTX !:DKBP:S[]<6=</'PK/0&#A?51 J7O")RNRA(_PHCDKEDJ=+:P=G";EC7>8^ 
PB6,@SXM*:>6D7&OO3#O\#:-0$B#%(9.CB7$IW"*N*8PK_O3)T;Q.'YVR+'LPM$GS
P.LI<,.!LM'EB9AB8Q0;P$VOI-^Y!0=M(H%K"G!H%*U$1!-QM SJJE\40;.C^<E@N
P]^SR1:0F2"05QL(Q/$U7 DG9*$Z)0QS\ 1[QM5@J?YO];$5Q_3C^8MSH@(S2GX"+
PB$ #ZH25'1B8:RM5X:J]AXY1A-!RRR^9M Y_QL;=MI-VG5J=?"KJR2ZQU(>):M.5
P$E\*"Y!"WL+8WVPNOLD!R,AH4JS5)QBN^WBYTZ[(*HRO9@?,V<=!. MMZT>,]QJ:
P>I_#2^?6[-6TGP2]=Y5P\H5!I+Y9IAP_)5.@-<5V"\5""Y0<,U.SO"4 F=(O:'Y(
P,Q6-<O%'%DFLOG,@+ ]H)4Z"2+5<!Z$7])>T(=[=M 61WKI<VJ]F 1;'I-+?;X!+
P>S8-A%KE]/?9< 8$#O0!TN-ZJPWQV&;,32O<0U;/@U!PT&';DE8WQ%17"0/=7\$\
P(6>:JS 7RV%:LXLN8BD </B<.[:UWZ_H1@^BRW<W<9%YV_D/]MV"S^C=W#2E:_5*
P^CCD(EQ9!P#"9F0G?AQ!D,'=R,@"C+!<4A7!'_4(STIJ5SSQQ6;269D?7QA42)M5
P(:K8F!SSP\MY@Y _'BNU;'IZT@$>@N'NJY7;7H3CF.' 3_6<$<CA.R6&T\P_4!DF
PUILZ9W3:#R*A[+S)3!:&$I9K-UO%/1TK7MV__P**'A./X5) UIEGWV7F6C0].YT]
P]9+:<=G?[+W)9B]Y1N0FF D;"N<OZ2;=86PW UR-?RR2YD"4^;J07XI*N/:VH04*
P(M#<"]%$C^=%<)7D+'3N &:-)G 1<821Y>+Q^'<30[$"N#7AK?(PR"7&C]DBYY^=
PKL4QH?5_8Z-F]AH'TG%C">4CJ&\[K4M+3?GL[%M#Q:4A;[R>J^<DZ7>&:!$5Q1ON
PSOF[X0@$-;3>:$;\"LASU?YU1WRP4*M94X7'^?PQ+U2_1V)?R!.MU'J3S?L&O\>5
P9,JT]HM:HR%*9W5Q]47K(SY2%LEK&'NEIKC\=;IRF!!MLT:W@/F3G3<[XZ]26(5L
PL;B$',57"8"X/808<OM[)8G4OV(1 XYG[HQ@QQKQ7T)XM%SVQM<TAT.>6*?Q15;@
P&08FG')+Y7!D76R%E9I"D$1 PY'FMG1(QN='$:R0WIH*BGS;1R^]9Y'_':[61+C!
P4%5>-_[].^"Q@TT04^IZ7(*4#DZU:;$V-EM_H@EMJ?S\WU6>RUTFS1G(P;'S7+D"
P;U^BKE<.8C\;+,A[K0-K&VZ@\WPZ'4"1976J6"5#N-O5_'<V+_1;(->>1J=Y&/=-
P2EO4=@.WF=?N#WI"-Y ($H*YH/\1'(U38C O!']"U%"_S*9-!N13)EITMJ)C]')-
PS&O$I+<-.,6/<25;<"*@<ZOL?;^'W19I1\]H!'&H-PC^?H;[QZG=_>LG!-XSI7Y6
P*:HX+!L.(-]&> W"A M(EDB3'@=SOIBN7PH@?^"6_NM>4>1,6KPSY14R38]9W&R.
P#;;!\+EDMH0JSV VYZ6[56TU7!S1G'SQ.]YZ1[@!J GXV@<=)2(\+D]4SG(!8T1U
PB$FVT(8!7HWSW&8]U?"(S(U$%B-&@AK9 2U;&9.I_)IL'R(&1F74]OZY,#X?\RSP
P*0"$X$$%^NQ6/YNX1W>,,HEV6EA,N 271:W[M,)M/M2.SHT/HL:F1W'CF[T9]N'!
P?FI\Z0KKG2OP<B ,N""0!IZ&[9R[CE7I/XKX@/?;VWS"J(,Y3KQ@I]LI+;_<9BV#
P^Q?S,32M5S3B9C-'G2F<.>LS@,V&<=4^*BDR^"EZ(=FZ?6DH^&E3Z&/8!"A3EM]'
PLW>)%=QM3*&4 EL,R :_UQ1'^OF5W<NK HAN:@-E1QT#*29CBC7)H[R:VVSU.Y\4
PH\M?'+"J5R%J=T,)ZGX)"KXRT3N<#RGN88QBQ9K:LWJ2$XVCC);#ZW()D4R(I_<U
P\F0#S729/\;AMW%6.A&05-/W%")V1M3 8E)(RU>"J@"&W#RZTC,8+4!JR;2O67M"
PE51,\-S>V,7^>->C.JY*TE?.&.-ZYCYY(D/=U;Z8IG*S%P84G\(L,L^)'?!9KLT]
P"P+L;5,"22LDEQ\)&3@GL@GZ<_1XIRS]_>K;0B/1V^LXK^C^BPOP-9T\""NL$B (
PC0@7*IC_F]AFGFPCGTR/<VDKR(=0Z"$Y;$YNSZ.AX@NX+'IU2[,F<<!6E\P2XF2V
PT?!2X+M1@;(RNE0+Z4WD'LVD5HUM/GO/_X,PH(SW)QNXDO)TG6:2S12CF%(X:=8N
P$=".FGM+@FE;82@L.^"?V%QWBEM6.N3()D4--9O.NDJ<O 2&,,#Y/##$$%Z1BN%%
P%Y74H*0.C?#F@+Z$+6JLDK (0?*M1(F4.0XQC/7)K=(2#K/+^!Z4I6\KX1,%"WUQ
PU_Z]!X$+9@[&VVU+H/M?=Z$B^\ ]][2,*QZ+=H.'Z3TKKP_.D,:QMD6HY#E.567/
P!+[^[+FDZ!(W+0Y+%1>25.X?\8" 2,IU*5@PQD'KW,C<5)#))]%5&I$J-[>%IA(M
P;UL--NC,L&,8(I%"!5J=64Q Q>]N(;U5NUEE%T7;=:QI:.;X[ECVYVN62';CXC[H
PC>@2 T#U G<-FZ=1F<;GZ58*6=4PW Z+&&&H=G23#?><B$85D1+BPIB%SIA@QOG'
PW#Y0MZS>@Q=UU>G\Q0:45=\RC&XD'X3C+*3T3#Z"6MFG@5?RJX$U"$OWR5_6Q;P[
P]O.YLCU"H;DT3BRXEHNF@?9):K2QO+^GT_LH3<+UQ3@F7X/\)'<)X59('KE'XP1K
PQG(T'5?/O$($!!>PX&M!QBHQ+B5"&#SS?6)ABE*T3*'5Z>'W"%\T(^ZBTZK,X*.)
PE$7]S.]9U&UZM8UQ1MV0%2'DFPE<O$Q6A.B4\96,14%'WR@#J$H15=X.8#2X<L._
P7=#3*-Y HVQ/P*W\RPN&!(5Q:=$^(-(Q:EW82Q\P\L\*^W1WDVH*&3<ET56T8(ZE
P]Y;11[7=GIX65H8ZOK.[X&J;W+>=7!#E9GFI+# @Z[>;50&Z9D$%)$-A4&"7@$+3
P(#N!.*<-&BUYLQ.60?K9#<6L/R'[%@+G#Z@/.U*:,E <#/VZ/G4UQN<ENL4I(".@
PJ)]8FX'C:")(.V$'$>:C0?R<:5_=__G#_+,4D?/+2\H _E:M"X ^*"-M(/*K^)!A
POQK-*IY&DHM1. .KZCXZ(@D;OEI>,0LNFE&!3)]6=>,9D;?V4-!B=M8RJ,I5<G^E
PFWR;XY2,8@/SXB\KA[$;WUKS[T$>I24<AP2Y-(V8Z'\Z:B+ZDOAO%?&6Q5?=?1PY
P2G50QB.)3?/T3\].H2D.63&0,LJ"?0G\CC[#=D*N>%O@%/ YDB257@#WU",)9L!!
PH9JG@S)N&KX]=^,\?:S#;98ZP@J-+5B"'\UT\!ZU(QJ^?7CK%M-;285<!A%QC9PP
PS:FPA"Z":24Q(NTXJ#\SQD2VB9<:%"QQ3Y&('T!!H7*];_R-'QGS 0<^S)'CIB$/
P10=W8M]9 C&BI%[>J@F H>ZD'V-RE1SFN0>UBNP/M7[AV0[API>3XFB;0T 5)_0:
P.1K>ECV$M;%"3[#H.^O<=NN1(5;N7$S:3A4Q)E]74Y[3@^^^C_!+CT+[,B"AZ,"*
PC0F\.@X5NC$HOMSX/C1S 6CCED'<H110D5O8+-E@'S*K$IP9]2^=9P7:N?>##.8;
P7J"2Q@R; $]AP&=LTAO5=QC^\8BA&/R"Q5FI<U6'8#M(G">;YQMR1^)H?^4JJ%8!
P L,!Q*77L(M@"LTVUN BM4#<K,F6@5G^< ?OC]&4_K.P/:?/XMV]@"J^%)-:OY%]
P6;+N:G=0+@LZWQG(K=C*(2.I6S+>D_?0!VU718?YA;CHY]M2A!=5$%O\]6I#?/3G
P+,NI:H%<?U#EI1A_H[7<NNNB?PGL"\SM@;068%[2SL:[><MYH<B(:\5K?Z W>XV6
P,-D6[(U2D53DNZ_SNO@V=/_FY-W)QEC]B*IKOBS.Y$$I#*36IK\@\_)1VW>[/ <$
PPZ33E'>V./V$I^SZ+ QK,?94*S =OJN-IQ(JXL.%8H:2$"CI<5?A0BVML)Z68!W%
PC9I0W$&X?07#JE,=((-<&37H.$(% KBM;5(08;:VH]=9MKI"_3FV/4&G=4HF3$Z>
P._P)0W/9DYM'9Y\!JDT/LGM"922=E-3-+50<(5<'UQONH,]_#?_6WYY5..M4^N"&
PQ*M>-K$I!BXZ=,9!!172_%V'::7T#TO!:"C7];;FO-1T'CV=( 62E[3;/%=]&YA?
P%7H"5NO;^72(H\/0U['GVHXPYXX5%MD"^LM]/G'B V? ,^T*P*0$K+@T0G.=0LS;
P2::HCP0&TF3W(D,E:FG)SPCRH4&5/ Y(1@N\_^.),"RR6>LAZ8X5*^).>./WO[R#
PBP+P-'IAB1U&^#I]S!G_NB,3IHNIN%>@!%(M9ILHIEVME3Q\M+,^<PU6WF4?AQ2S
P\S[R]?53AEF<F(BDJD35M!:3_D=N2A$RS7;MBG(%%E@29^L0D9NX&[&,AEB3_Z!I
PG\_X_>:@C*Q-"VFYCJS7="%K4G,21!S\DOK7>3,U1U%X:IE9CBS%JM?LA-AFD_ZP
P#\@9#YWF6^UL=ODJQ2FFN8J<JTW+O"VC.QF?(M+!PWUM=\ 9?O(;^:5X#SHX%3B]
PE7E]E?8SH15:L2<W7QQLJA 5!Z%.=)Z ]D28JDBS\0$EJ_A4UP87[6[<!IV=Y]9]
P$8GCSX#@2(@IJ)O3Z\<1*Z1H+1HPKZIL_N=*,G_3>E,]QC-2>+JDG@[" L*&0-[3
P 5+K4FBV<40K:A'-OQ1K"H_C9]\8%F73HBUK!@'ZTNISG;2@V1!57?'?7XK?&P<S
P)&\-(\X'7VR"^[=9Z*PN.EW(EDS,]1'C^\VCW7U K*_))F=*45_Y @$I<!$6F.>1
P&JY-FX\+L@@H-H736H9Q(M XXEZ$N<.;Z?BA0^83/>0H2,S&9K"[A5L/3FMU^;%;
P50H6>HZK(5&/HBB61M?Y+V"Q/EX*4OTLCKA%+R([OW)?.['#"M3# OY=1 4L]3Y:
PCZKL#,LYQHK&U' K1<;5ZKGP,LL18VN,:-4;-E>!J6S#E1Z"F]^3^I<44S7?RN]F
P9$8-"$-?9 YV[$;+\^RK+-T*?E:,/>=9]5:NQSZ5'"\X]=V(&3-KERV<N@M^9^]"
P;)Y\)*I)IM<N9!S:4_C+>ME.PKY""G94;" 19YY'H:=9 ^V+A7AAK_1WIWJ!)C8$
PVN'T-A6OC_".A)&/'SN)I* 264-?@YA9PT[ZW:]WHYR:RT[B*WJ9R\ WQ4G@"77.
P^A>G,>R<E5M<R$;^I+O#EMZ\'SMH/-/V 5K%I"E[]+]+B+54ZED4/ML>-0/K7IWJ
PCS=JPRY[*LF O:@3)7G1%(#XKI4=X+-?=3\]-J[1,Q?Q+"-%#+IP_]K!/PD3'YZ-
PX-F>6P-)Z> /F=]FR0V:7^>U4=#(Z;VJ.1=KA EI<@E6%.<7<9#^6)EF@KO<3P@E
PJIH453L3._93[8G,@RI*M*,@0N@]9G<]IJR5!Q3$_KXI.%ZLDC%N/.8ON]?>E?QD
PQZ+]0.$*_]UT(!VNW[X?=7L'P51N_) "MI36K7*[TI8S/O]FH+KBV(@DZ@I/;T[K
PW*K?-Z\1Z'(2,^).)Z=Q:@X,6BDB*@#$]B@:1$*W>[74T'JS#%0\VZH<&7WU!-><
PZ@JK%NO"C,)/:H,\*AWY+)I= 7R[[Q8G+(R=(NL1"]S%<SE;$&J=\8>L]%9-JYK!
P&CU=9A#)SB<OQ-:KA&SC@X>LXO<D<(<L4Q5(+5&)W *A(EXZ0YEQHDB=8N/8>NHU
PE,KMM]_B-_$::)'.U4A^UJ14^H 'XO3C;#2JE)+"0@&>$9M-T[2;R0CNK'%\9QWM
P+32OQR)0C&L\MJEWO)E7&-D D8?FW LGF\6<"KSK7R0.F->-]$7"0++U<Q.4@2F.
P?5S3QX=+!9#@DC%G<BF6!LGO5$T9"@LSS1K.X]P]?AG(\V8MZ?MJRB'A[;\M&V?W
P/X<S<L<)YZP@V9!!!,-,?[&PA'2>7-Y_#9WD4'1-*:H2%Z^;8@SL K_>Y!V6(:C6
PFA#U;1:Q;06,+AO%DPJ(QR##0/,3JX ?UB/>H<E<X"3DXJ;X"BX9W $V3AZAZA4\
P[97^V+*L15\TF]9O9! 1&_,NU"+4CB;S[2GX]_';%@[V0MS%9^P79KB>;ETW$J.O
P%"L%SC8(1AV?POYJ $=]U*GK-)KL[?L7FYI-;GRIL#($1XZ'H">?\+SE:*P=8,,:
PUUV7%_MHDL72AE*3<'S,F,3!C464?U$Q4P@C!A@+V%("MXRLU+[X=#D?#'2[WE(U
PL=T6,;>EP/:>WU/9-9'2N5?"/X4_5#R=,C*OIO>+:S;1_PY!=/<&[#_\E>GU6.B,
P2+WB /D>; PU5LO^N9 /%LJKY05PO9^=P2#)9^MTUYT4=J!N :SY;?I!A$>^%OIJ
P$_/G+3'PPR6D(5T(#@A($$'L\!)$!PD8- @61[3GIR#>O"S].1M0D:!$Z*P2_4WP
PRE@<YYCZ'I$_J-#+XKLKG:!NIU 1=OI#@)DK21YV]FXXI3D9B\98-U=_!E5[]*$E
PYC7Z\X[^R+<WKSZF^,ZHP?O?!\$$EI*+-26^ZXH?Z8PLJ*Q"F GP#(9EUU'&!>WM
P]$S?WZD"XF(R0L)>N/Y4Q[D5@+J:$9EQH(+P$@U2_EX<%^TJ2(6*IP!+2*'Y]8[#
P)RA]&O%_-W@IZV/"CC*G6A R- &(-BYM0@TQ*H!DR+AH1Z9F2*J#VZ3* *W:9R[2
PUP6A.O%(1@;\(8L+3F^,R6Z?63O9@D:.EMV7X=CW1"%K++H3LKV[ (FC?9*Q& 0#
P3>N6$@+%.^ UW,B@%19$Y\Z'L$%PK)$+9ILEC[OU79%/83:&'$C<[T3>_-8^/8,O
P4#"02XQ=%SRSJ:H,J#4P)\N3QA&VN<=GG59F+^IOFC!SEF22R+@]9+<]QQ P]EYT
P*-49"X8H88%\E4^:?U6=9KV_>_Y>X9AJP^Q=)C3YIK971&34*[/6>L_=&?V W=X-
PN<IGB@UUT/!U%"1\3)_@/LI!3RIKV3LN($\N9!>X3D6P:&I*T(H;9]TU&=='H'JU
PF)P1G;)!<88/Z*2D66 '^=>E[]-)<W2@?!YD*/:/8MC%HV:4!$UIO[)W6AU0MJ7M
P[9MF<*T7I8,.\K0ZN_R$ US0^\OKWI3CZCN39Y&JLE.7:F3$U."?[G8(,M03#W=Q
P?2\FQ"%WE'SR!'*;RL<J^P\?85=.4\DQ+ -=*<N]"6,M-<M#JF7D=QOAO9JW!TAO
PJL@$065J^R6V;=E6GT&MQ;N4137W[K@@$AU^!BX5K1TZ3IW+=U_J]6I\MIS]%<7@
PO':MCW"=^* K>QLJPDPM;+!_1?,KLD,9RNP.F3K(Z.  VB([N&"FMM!A8ZMJ,EF0
P=!)WV+;N,,$LJ-@A(OHF;/H?4UMO$UFOC[%04&OY-BAZ=[4WV4$1 /+9'OP2GRG 
PZMR;$N3 'F&@*I_][."M#$/(>,D!F)DM8B3'*&$!^AI@@L\83X;216:AT'&%%ZF"
P3%#O;)D0,,<*V@^#!#74@-OW-I/Y" :?V[64I;T>OBGQ3/#O3?</5=6KS\3%_?T5
P6?SUG>HTULW?VZ=439"XT(?(6$93BJA,0<5XY=.8SDGDS=,B,RH>B$N<!!Y4K()^
P2L!'9U1\')S3Q9Y0;1ZUIM8Q) M"G8U.)K_$3Y.^:>68ANVGC2/CVX52X6B.'$B7
PJCRIO#DHQ[PQI9=KW/J'%>-0T9$V<BX*K?0081;\'67G(D.J1<7M3Q*A@?@0A0&,
PS>@Y#4UBJ2G"A:VH#%P=P$;3J+8IIF&GQKRP]>KU+$&PC*'2EO^;<9LJR.=;=O@T
P9MPU'76B,\":(AEBU$@1MZD)([*G]LK&R1F3I'T[1:Z<; NKU,DZ.IX!=+S67@F6
P_N%G"TC2X%&5(O_!$0&?KAUL-X.Z5/B_/NJ%M)!1WZ0RF%=Y(@-DB-CP710A-3" 
P,Z2-5!I.J6X_"FV_T9.U4!#$U^3K1.MURC/\N2MU'*R*DJH8LXET&"=H5.J*G= @
P24Y_\^PSJ#1>K!(-Q8EF6HAM )=ID!CO,&@H8D5>LE?H6(*U/:TFM,)2]9D:4\"L
P8!1MMLG<G3^#WVD'N99(&O%PX"G3\%,00'^EG_I%,MOILRZ <@*!* ?/2P#K3GU 
PU['A>QZO6?=(XOT-?;*B#>GLB!'UTVG^?"8WZ2Y)[K=&HF5C8AX.P ;YL:24M/6T
PIKX7 8NKOIE_YWCU;:P7,:$O=*X)L9. I7!U*[\*D'W4W*?0&<2!,2?_'0T.Q[R.
P?0_AV];@PYMY%)F=571+M,;%:-8TO;,XMJ$5)N,X9XWKYZ(3-P3/^.C-Y'D&I?8V
PJJM%*&R"UY7T53:>I';FUO:'8Y0;JKUJGI,>E9WVOAF6$L/BGD#(UJD)D/=UVZ\)
P'8^F0T8S"K6SV=2X_KYL T!$&&#$,0V R-P@=@B.R!29Z$"2_DS[9WX=81)=.>1+
P&$?<)Q>0=08*A(?PP#RGDD_)MT<B:SW ;=/KKG"((P9J#CN,[2+^E(08!I7%/28*
P.7,V6&TYR.88Z(1E6IYI^=]Y3,!EG5;O !>9.0**-H1\TMFC_P) @YRHJ*QA,0QE
P'F6]M1.,ND%P0KE(UD7@PP#!C8BYGQ7<4OY MM#7G-FH*=@'_)LMA3P2F^+HO&.F
PV8SB]:%MQQ#4AG4I&"*M2$^/\;A<Q1_V8[Q$L(#=*NY<C3-YU>\M5FLF 1M=3ND:
P#/R]]FB>UK2 R-<T;W8W=[[50OS#2R;NU7+!=!JDRV71OK=W$O!&,\<"\YOZX15U
P9W*+U6A^\*[K1B6=_+?:;:BY?PZ(\><V*8P[\C:ET0<VNPTT%F5#5+&?6DH5/<#!
P<M<9[29A 4*PF]P^ J-4N*(RU[ +D72?SP%BBZ76"Q/<C30'>5?ZG6_OPTIJ/A1[
P_[^Q.E9_\WX,N0SXGB@)'8+%A='9(M)4!'!$>7VA0/3P)[7O0*8/(4/PB5V2"6E?
PK8LB?6(5QS;].[UR+I:4IFYCH)]!X8OET;()PO(?ZLT_K>QLO,8'^U/#KK05B,A/
P$SM:'VCF"6%W61//I7W=^.]&6&J6@TS447KH;%O.90V_-]_U_?7CW-^WR>&DTQ$1
P$8Z\U(Q68\V;_0!$'JGCYLT.DS:'$UM]_>9SZ#0*-U Q4:I7#F(/+G>]2Q/;TV,=
PCY$26MRMT>S6_#NP#TKVI8"0, $U8)H2BH4.%XH=$[=PA6K."6!C >P.JD.-@8RB
PQ'R[$KEA(G.63H'8.1@K VIX^M0+0&7H(VT(>G3@_UV#;R19KTDF0>.V7?V#EE*/
PDF#L!3+ VL=C RK)6R67U#!Y##4<@CQE[>*E14#X,!X0\ J>QC5Z4I+9',#7>T/"
PU&#5MR$.!U2STZ;GT!0GU"I"DY-#-*/'J4Q?X !/2!&7'WOP2O;#"&IN?Y#F:EZ1
P;P1RH![MJ=L9^=3"6BD(5%QW?G]A7RN]H;R86A/PL()2D]T$\[!)<O91)<OB&K;J
P2A2G#IX4OIUBXJ_Y."GPO]&BSF#WF#E/=[E]VM,&&^3I,EU(< )HPQ)F0;;@X).<
PNLQ35WE#]",.8@V>4NQ\.*=>V!@J<5"GB^W/\9E[C:?EHKS&.8DZU@6HF,A54#E\
PPSP%V?,G!N!E'7K<^2%:5G,+P21!7I>3:A<YCF"K)2#L0@PQ/DW_]7L.09;.XLS=
PST3RN2T"A_8W,YUFUI>D"82<N^9EN"G>T<SR8]0L)#NNPHFG!9>&$#^C=U39[0Z[
P<?*70Q6EUZ)"149FI(#YY@IXOW-(7M$5B9@#)6@<<(X(1)KO;9"4WYPAP;(/KIO@
PI)JF^<2^8JPC8:B"VT08JQYS596'I,=:2?'/6#7NAK??=\-POB(_M#6&;DV:A.WD
P!HU2\2'L<UR?]Q_.T6%^*E8]3QJA(-'O==K(E-B8<F(L?#3>II!#PE; *UY\J&)L
PL-/\1%1 )5)4MBE 5%K;<-(-(%8>:Q?8;7FO8?Z]2>4OPW14()'@CRZX? XMDV8'
P-[&(LIT%TK>+BCK5W4[<Y!0[=@K$M0Q6*3A1VX.\-H4!@J*EY?N31'#2/3ZC(-F?
P1B9"SQ&QY9*)94@;M8AO X7B/Y[:+VA^:SRF:4+0/02%BQ;RD.?[HJB^SF8#@5"0
PVZ:T5&CM@>B R&6M=E!B-NTPYO!*B4/C[0D5E3I./80G&=I$:1EHAW9$-$8;QK"M
PCAVU33L+''R^+NRI,4=!G'J14_X_Z B R#G.VR%P0FBDD*I8%!2BMV($8E'7QDP 
P*29,T+*09&$WC&UM0D3XXAL1?%.%Z=.SY6CP=Q5#P]6=IZBI=+#@<,IE^V8[-S32
POC2@IQ?PFUBP4HD@6'^F0T8)7S6&S!BTSHY?<=J[13^'#V]#>(VF \4)?7\KD\2S
P0[U'DV_D![#F^RR=O%\%^3\O=4**\C+;[#&"@D_^F[B#D(>NC34VNT\=I7 ;J!>%
PI@B^O.^U +^_9 !6GG4+.?X$N47=DX8=2HH<U:D<"OKE&RQA=O"S3LFD1YJF9HAE
P+N)W6G>7V_0M-S74.(CF>_GUSS3PPLJ^W; 9[2]H GFY0:8*)8JEE%ZW=UJ4?M.%
P\4V0#*0(:Y6CZW)'FHT:*/_Q,NOQF"FZ:YO=.P/FYB27$><(RB2E8 (F.O6")*"O
PIS$"Q-[-(D.WWH?J2'_)B.2N"L,.MY;,<TKV;4BQ_Y!2VHLS](K(:D:50]V;^/R?
PI;O^37ZUGZ)(,D]%J[*L$>A^E[1CA2'7SO&,&D3. 8H=?#06^S;T^PSM3KU[!@E#
P14R$1QKO6"8O#=N(P[K060]MO75.<:BKNZB_B2P^?1%AOR1XM!7EISX E5^\!>I_
PE U)_<S1LP1 $Z?]..K753R%KLBP$:8C1VI'H981\5@7 Z.J"%F\CIQW*/<ML:=-
P35B-F''W'I@45_ZKE9<DKL)*6X(IFJ_VWU<8CN6P4N3 #:9+E&X!TGC2WSFL^W_R
P5H(8>6.9L7Q [3M-.@DWXK)A,E8BTHHR5TPXU<\$M/7U#ED'?X5?%^JWXTQ)?[#1
PAVPV!87UX,&R VL/U->"K8AA_2VJ?B58IMOZS(8I8]5,S<$=_9PVB! YL]:4NOP\
PEP54R"<YS&?WVC,QM&V>N;Y!%0$8O/E==(*AX 6>C&!$#NNR=P=T6I^^^BI\/*E[
PKBDS^%*WU]'GCRD%$2,NN]R\YP!!%?=V9C$Z0:C=&7/_UGF+:2;HC6B"75"8K,AM
PN=XW'1:\5B;E*:*I</V+N/8/=@(I-\B#<AQ/V\3__(Q4#F9-H EK:.H)XP,5,^!!
P$S"2B48S"][T[19K))C@[?G@Y6=B8X0S=U\)*AT,/A-PG(70@6H;C\>!> O]N-AJ
PEGY;4%UK$J,@P'R7@7+NP=%^OOGF.O3WR.YH]C8OW4XPXUQ4[?"KW'^DKNSG>BD1
PNB\WG]U:I>%,(&59,;:,]7Y@Z1D"7^)?X+VN"!'3;CRS\[+(T2OE=CNG2M][SXM<
P*1Y*0(9C"8LR0H!$)7A9(X$0ESL41$K?_PS ^Z@VP=H&)SCORY/0+%R@$8NYZ<]6
P,UH]<+X==]K?D8.D<Q$A;NZ/7L* &(SN=IIAN7G! $6:O]G75R8VF;(JK[/2L:/D
P#I>T1[V+4*97-B@[1+065O!#Q[I0@-"5?V!F44BS>FW[H0;@[VNIFDT-7D _9AUI
PZ]J8[A^WJ;.:W^JB:DT/R+/7=U.W1":\NT2H[<X1>_Z*U-HHOE#-RY>E:DY4OU))
P'!1O653*)793TN- Q+$ R5F=A:17";-J6%(->W[5 SRS/=4T%HB#W;P/&.:;(K&F
PNWO3H@D%ZY-?M[9)*W H*!V#P0P1W[C<:JNU2KY?&P7L<607);*5%<6[GV.U5M0<
PC/#*O+0HU"X+W%8DE8PW=CI8Y6RN'(^=MM>]Y7L#04U3<7L[?AWT] G5-9^>*HT\
P%!#(XN\J\XR'-H;$1Q8*=?@[.U]6Q$TK\V_2(JOLVB/Y]C3J:'H6+GQ$Z;\8SR_'
PK6>U^;:Q4I6^B93N2J17 =JP#QK0U@BM]2P&*F"4T(&.B=R7?(U&>KQ[AZ(Y24#+
P(LV-,;]JG (8V:82J=>: )"<KFAOB,TNU*L%V?-+#)+/.\= A6+0T=6%7JU@5%= 
PG (9AT4+@Y">8%<$74^&'3DLSR.HT-<8'0/)(-FT& ]29Q"ZAG!J[$4.LBA$1,]6
PD4:V"+\I,4;!*<N'%Y,(!KTV^IP6H1G#LL7&IRJJ4D/NFRU 5!E6[O%J9\['][\;
P8"(*+OD!#@MYW'A;+HIC%/N *Z 28=;J>3C(LM\-LV&MJ_QR_]*$'&4$%1*1)/Q<
P15,/%K&L 29E;1('ECV/_PXN?7">*J6>L $&(@/ 5#YH5OJF'I4K.2)8DET6'*0E
PE5A:CE((/.X*L /"\UU8[TG>U6?&W\<Q*YSA"&GN!Z$B). VY8F,:A"VHS]-#_EX
P'"+B=,D%0^/0:3DR6Y )VH(5K(/CW0%S1#^?)6J>J02F%[,JH8RD]O3(2UI^APVU
PKD+L/@@P:VG0Q7(RT$W2_,8RE!&> 8U[92ME'H%LQOJ* Z)TZN\8-]# ^A0FKR"C
PO/P$MR);W_!];!7?/:\S*.U6/QO#=-'!'D&I;S%:#8XKYV9TG(:?+N*ZML,X!/GK
PT9VU+"HX8>'"^-0($.@A5RE/M#JY>2_Y/,"\N]?($..1+U<1LFYWZ69[%IO]U "Y
PWAXC.!O,*I>K;_!8"^@98=3_8R38.I2E\D"4)11,$3/ 6F"=C#ODRM;%SMN(<LAX
P@V+Y6!T41?CYBRD?@6A5  LUKHA+EB!H4[E30L2&^K;&%98-VP>?9(F#FU_S%=/F
P'D NPN1$D&0V2B5FMDNCE3UL6(\&HY_Y68^J(M2^6)XLCSCT1ZVL*+@"+B?<4#/7
P_?$,?O^577$E18#A.\[(^/$&;'L'PY'.0-\DP"(5_ULX ,B1_,8*,",K9>1>K4"Z
PPH'#%^$+WFL,G'H-]#M1I;3UCWMT(?K.]: [7BH'<T=@==66?(8([3(>X&UEU[?K
PS$!D9 [2T(R0VXY)Q]]MVV-0432POG+?LV5%F![$I2 DO\I_[9_-D)I#(!A:Y:QT
P0%.K.T-G*EC'@'&1^L66S N,1,*3=H TH6XC*)Q$984(,AQ=4T2$:DDT\-&F!ILT
PR=:^QASY5;YD#4J46[VCT\#TXHW\51S0(3ME]"GY4X9[AL1N/1=A@:K;L=\[O0F&
PG?C9?:<U^S7RA)O,<#K%/#HZYA*X0XW<245B,$_EPZ[6UO:\X\,.;V!"ME^4H"*?
PWHJ%PS%<^WLK#VN<J!C>;U)T%V:@=&)S< 63?'M[$^K%"0/7&^H =[L+Y&=4*B&W
PT<)W"Z4"A/$5:TYQ?90+UTW>$*WZ\Q?]\3N..TDNADC&#1O!0SGRW>([T)#&;E]@
P J1M@&Y8(%X,^/+5$&Q:8NKLC!NCEJ]75/2#)!8E63:7Y-R "(2H.T:W]KZ&1^A0
P[;+^*8IKEY1)K_K >SMS\1.OYQQMR;R3P30>88CD?V(/SL^7DTU0S"RFKX\THMA<
PMTM4=?BLBU_Y^Z+H0=<^MHY;N;3NF<3PLR6GP?73DLU^X:ZJ4Q'4A0%.>I$B30B3
PL=$6LBTZ.0/"7H&K&4*/PHGQN@]+U3(BC1^]:[6U[0R(I_-A:9H]SYHQV+-6W?$<
P*A>XF9B6F3^>VN 17;Q.1N 3SF O\KD+YW=Z(0)W1TD.PIJT0_9"394H&MMJA_&O
P3QEU'1:L!4,HFD+[GUW)OR2XI++LAPYBNR7Z.^L]'04Q?;FV_TUCA6&8.<RL@&)4
PYE$'2:E*?QE]VND\S_O7'."#JSC<.*UIL&"G"[^5?<O<$((B-5R4B"U 352\$/Y=
P7(2&_@JQN5/86-!SE]AIW&I%2_1]Q/PL53=&M-O'2WR!]!NB@D8F*NRDL@6+F.>L
P)Z1-!_CT)FLO R$G7:R.(.: 9"N4N10?,9X%_@^5D7#4#G)K)''0^WV(_YM)&"86
PVQ*,M$IUF,9UP/VFU$V<Y <6DKK"F<.E)OUN*7P#30ROH2/^DSH!H>L)4(S EY)%
PC7(.8O'&^*0CAG()11?]7Q,1:&>%6J*:=37*((?O-J*O'0+BI&L]T5]3_ 96S+*H
P^IM(/RO?%CZM#Y_.61Q L"J^&M^9OC\>?J,_^W@BYK5+GSOK:M<6D5&2Q0>%1<GD
PYH%<A!:% Y.)[B^^%F]9O:!E46WZ>=2 VJ:6CB2ERR"N((8]@. ;J& <U2#=S4=/
P1?0>?D,!W?E=FN\&78:[;2(\/'QD$_KU=AE#<E%,Q<![FF2L*_S'=IL2^D?</G@!
P\:K*PLUJXY,S>6TR]!ULXV('TAX'03,]B3+Q5=N<YB*C' M85% 2S/S'+(B/OF*M
P!FX^ M -9F@4L>FIKQV9BX(.2EAC);K8D.'$]2#/QMI[^SH6VTN&UL4;DN\I;X[[
P:L#L\@?>H;L*?I$@K/9<7SE'>1FNDZX$:)-V1/>@?<9M4GP?@6OVD@H:KEY69@%U
PWL+3+^L?EK#ESQ=?%B.O8\&NHJJZ/&%^YNKUYC$P=G-3P4 W59YJJ*+V.FWRWH:O
P'.Y(9IG& BL(@ E?"V6<9<?/'??2/0TOP#M6]$69Z'$[_J%FA1FC^%,MOE\B$!:W
PQ-OJ>B\O.**BVZ&4/N0G$>_1H?!%1,9&+?GJDNU#6,4.9KTJZ@U])SID7! 1Q3YY
P-YOIN8/&,KALM7'T-V6/PQIH8D#A>0NN;.X81M)?R 2-H)G\33:IB*+1OFGJWO"Y
P&0G$E.8\M]17T+<]'=O"KREY/5\5\=V EE&NN6?_O6?:P^2YVV+U4*@Y,>7J(%B>
P[A%^B#MZH,K!.@W55KWABC#K_C171NTIH[BM*B;LGB'0>=1+3:7/&H,*3]2@.[T)
PN"I7[Z0_]DRW1WW0@&273RC;]*</^VZFZ/8_L+1'0:<:IHU@5#8ZGV0'Q 3CV*:]
P[LB8O_HE,ISO0O02=P?AGKBYZ+4@\P@\'^G9FTYM(H9(_!1SY?T?QJ"*J\G"B9)Z
PFH/[7G,]Q6&-&!?FO-M/_8"/T2RU%+(]1,T%4GP8>&7C@PO:TCXBF!E6J1A@93W&
P2-G!3F-^6/+<B"%7!CNMRT3P36GI2LYVP&'18L#U,1G4#GFY$.<9CYPHRNXM" 06
PB"9Y>\(012B49_16<.VX]@Z\P[*AK=WJE977?=]@M%6@8&N1SDHV01TXUGW,/R(%
P(3,J<KFA%K@6@U?0[XF_SVH#9[DKFRC@-Q@"<:N+1584Z68RJD((( R0KJ4;SBHP
PL,&."7.4FQT4V-ZVPUYMNFIJ=;<F_. 6WV4NKIWI)_BHZ3@Z^J1J9P-6+7'[E,3I
P$BJWL9W$&"Y&&%&/)4TOKN9@8C9I=RW TX<@N6&,@MP'C2NH)U,"!9^:O LK%;Q7
P9' JBEE&F2Y?]%5&.A>K'+"QEY^TM4E GBW=Q%B0C]?YX/*-AF?X .EQ9-SC72IJ
P52^>$!N4G_Q\_C]<S<</E4KS_NI#LK96.*@OG)RX^=5J/!):J-O7,7?GHJ E*YR$
P:IWGYTQ$5$6QB#92"JE[L@A.AB.%JY"MQGX)# 77MMBW50%W%C_#GT42'.$W0SQ7
PCNPF8,S?*I7Z?;;N+?[AL!VO0?54'CG&8QW-I2!-ZFC=!,^\<FFC'6N&=Q+A$E3W
P[G7'J1S.O'XC5%]$+\9OS_,F^I*927^*#.T!2/M=5W28X$K--7+BD9P$#LA0#);*
PE#AX)?*T64_ ?5[O"?/(GQEX'!\ZIY1;TCK$)K@RG-N&[L+#4P91A[IE&</"Y\3&
P[% TI5C3$-I$AK=T9PK:!:-4?Y  5O5$9#WR)B;^K;!E,N$$RZJ;*&H8/[V/][WJ
P=6&2<S2V>V-P"4LY=V,GU,&.9;25AF-S7C&EO3M"4^>S-K>(@8:,F,[^0(3%;,2<
PJ\FE!>_-(_X6TG@TK=ALV!*9WM$H*5@GMN[UG]N\"J30L&$BAI[FIF<35E,5VZQA
P+=P504T&1)TSB66@(D]OHC?OLQ1-T;U<<].YWDRYJ"]JRH-=-(*1'@%LQZT:_%K?
P8D*_>BS,(X3ZB:)V/M30,<^2:&?T;USVGO;(1=.=+&(-"MP],OTV)0$AI0\?3OI 
P*<MC)75!3L+:O=H=YQQ ;;=@J?/NC#A@Y80+/N-[3<IID#$U;0IE][J.,PB)@QWJ
P%SX:"J&(G*F,)4":/6K'P&2M71DQ%;WA<(^I@/+JKY7\G46)K,<9!0%KG:Y2)@]Q
P>A:FORM;C;U8!7FKG%K?*9P)6Y%W@M[+7U<QON4*4Y9R2*CATD4@X(3_6$S _Y2B
PY%FG8QQF9;=CCIOA4.NF02 Q21;.0P39D9QQ5@#4_8B*9V6MBKI&6U&6G_6A4:[=
P:3&)6N*(&MW.RPAB5OP*BT3M/CM3-1<$^51",&)L"\4KGQ&1-]<=33YTVM5DIX13
P1]P<XJS#B9V_*;6H?0.V&28,N<9RCP^R^]'D!R)PZ^33(8@?H/GR:D25[ "\Y]_R
P=FJRMCK^-=/T/-<V.IZ1NT*RV?!GZ47!%/GUEV4UM^0,;)_%<I691B.6(S7P *KX
P5G.G-<+G7,!J"6_HU:CKPFSQ5EG%E,+Q&]#ZYTE<T@O*;PY;;ZT2_E2725YW>CLK
P\!,BNOOT=Z1I"Q6KYN=&&,(B1/H+&XD*5R;N".;\:S=0MJ],AH7'*4J6..IBQ^LM
PO-3>;6G0M#$0ZEL9D?#?:*+B\6 WGD!O#+,EXH,C$?,WV5Q98?2;\XLR6?M6V646
P/?DS]!%1AH8+P> &:*KTY4I%BF/(_Q3DL'T<6UJ;!B4,U6*"K-[#-BE+3*O4&Y5S
P,2.?D>+G01X%94X.(2XI0=NQ)<2DU:TL.SJGL7$#AL+8Y+FMI=Z_HC-&(*)*F)P/
P1.-7STQSAFR;H*3^%73UK-FTG-9S#VY#.FL*P 29+5K&H:P4?&K*:9CS!^Q:?9M6
PIY[7M(WZS \2#Z):P#8)5&)H?_7@+$>7KP8.A/5)N0-.3TY%_58(7C:P9;\AKD93
PR5I3DJZ&(_#S([ ^CP&FC&X6!]7=:Y,$*IJDZ(XDMC,T54MSZ?'MH5G/[+VZTD8&
P,_@BX ,23_3M;^DA?#)/\HV(D5W*A:H;KG!S"FV:@V55PV1M@X?+>;]&37$^UKAN
PO'WPR6>%X7F3>67;\U.-)(L!VB5\&H*)^#6.R%$ZD!]F8FPS<9A>^F;-AV&D!#F[
P*P^9#:K0-J6+\BV]]LRLRE69*5\N5NTMC>[]4U6=4()NF-8*4%44GDW:1G;JO" T
P^JL\3>_[]2LIQ#1)I7G];'EEM-RY>D%4YBR!"=6!ZD9R)DV#-75[&/R;!43ER?BT
P]3X3I$;&D?2:SHR:'8G&FFREHJ8VYX!M;R$YT]U8/.IK^$&G\T9R$P8%9U>YIZV8
P.W[PP794<N*B_.D(0XT?H:V9>@#/\S\FYID-Z8J0RZ$O^U,KE'_F#'<02[UVT%5;
P)8KKC $S$UV(/O::)EV)EK]9F1Z1L.U?_G4XGGP3=A:@_.B@[:KN\2.EA8,!]V]4
P*/O1-=5[?H]M8A&QM;K'>9*L-#F4/0(!GH5?7XC2;HDY%Z?VWNH<A\QHE7R+8G1D
PJ+JNV@S\DLI04[@Q_N F#"#FK3*#3VP/D]4PQO,5KN ]?\K!%+G<@1]=/GEW3B+C
P:YYBQH3F=\O=+/I2\__)"7O6JI0?7;N<S1+P ?P^&1O:LAIAATX2?9&!B:"%-]%U
P@'T=]4A%)H$_Z-K]K!0RV?$D+- .L8(F<=%_ZJ@)#C$A_I>'OPYCE%Z2'U15[(])
PAI)%.#OZ26&4-TE!E3%_V,W N/477X:UH4:\ Q5"7?4XITUZV39REY!:.*<PL8_K
PZV!AUA+.&"%%XI3A&F-"0T1 ZIEC/,I $F77'6<'MJ/BY4#AQ#S9[2UW 9PP@NR#
PI,WR_:<*=3'A8JV>&R0@=TW-I_A#\XH9V7&H \ \,O'L-#T0*J:I\<::-0:>J,Z\
POIA.ITG HJ^Z1\,DR_SHIV<.[VOW)E)[-BD.="C/[-GR*F&L%$$Z9M/X71T@P>4 
PI==C,B9/KW?-^AX]1W]\5I!+(<- 3Y8[F(/F7^0T^DV1*3@3[;5:*N;EC357I6Y,
PMRS-;[)4;>]Q^@3P^EBM%5F[=WM*>D!]9[3I&G?7&S*/RQHP^3L3Q_ -_=9NK%D^
PQ(5B23OY7U_Z??J/9&-^@?$:S\Y''$FR#YJ.(CSA;$?U):U%TW/,:&<&=?$Z(.F)
PE-=6Y:/3$T?R'GZZ<Q,A8<&F?R4TV)HX0,R $,^G]3_=)B.AIN5\J54$M4Y:?GI1
PF 57]?7[K=]^N]Z6/AM*3SD]&387 %'34&YR.,&R'X$OB@C-AJX+2!#@W1KCF;4<
P>6A;UD4#*<0FR+)6/M-4BW;A@5N* 0"3=2L]0X)@OZ7@*9!@$0D*F^:(9PLPR5[9
P"Y10OFU <APQ9A(AI'O.')-+\);7JPP*7\DW2A X$7V;SNQN--'#L-=()1N#[^=4
P<A[]-%1Z]:>!<8AY$I78=^TKR YGAG'GG$]!L>F@5L[J,?+WG7>,OZ %EV-S.9TY
P"6@;<LD!?&YL%E2_0+E'V"@/;AP[5AI$^H?=7?<4G<$JU'1B83,BTED&[#R3Y=!]
P)4X]4!']","^39X3"C<U5OF-Y*RC^*[:E-^.":%^&YZ:"]WRD256394;TDOS0).F
P7MVZ> ,\8=B?.?V6!2DW-I9MCX_(X)H_E:XN15*R-G9_D&!4+BB=UX1VNJ++Q\G[
PUD5RF:J@IAF9?O2PI:]PHVE+W &@$O-L5[[Z$"X8D,P8+%.10+RA&XKDD^^ C+8M
P?!EXGCI=><A[5(>%\DLX%^+/GG=8%80\9-C*Z_;FZF9MQR$GH>Z8%C;U:H]Y,]UJ
P#52[6QPSZ3\]*.[KK2>7?)N%VU@N:V:12 *LK3:&:?"&R%(T>G[?A=0D2]:@Q7*.
P4"5?>5*6";^/IDPC)HR.E5T"F>BLYD=O@\5+LCYLRTUHESZ $I^F8'MT_3.R#I!W
P$^*UJE6 /Y->Q5N?XL&+JR\<$5 US2OM>\/)3I9('J=18DE:2& 7CP'FJI$OZ)$W
PJE#JPS^%ZJ6%73 T#S9 1J-2\BT'A8-[4B[P:#N-GDPG;:G"R069^4,TO.86/NQV
PYIASRR,U0%>F=\',@C6>3=^^3):4C]QX9V9IYA#[[^\70<,L0,HV[X8<P C_L!U?
P78_AQTGYICAF!DICFADU_]_QN<Z=C;/G-+$D5DNWYO#F;?#F5T[0YB5_W]PRXMHX
P)/^D.I!YL&SOO81S!N3NI1,$KJ'>'"<R_=2MH2L,GN:$8!F\A7XZ"K=&%V]9DS3*
PR;[H=J[9,8KPG'$4*9:6</3?D^=EYM,<?-#JLU;@_XK_QGH5[3U5&"D#-M0_66V7
P>'O8U[*=/SH_GC2QSH]3ES$B76PD6V+GM'-GU7D" ]'@=]@SI^FTZH%_ -B\))O]
PWU5[\]27._MOSU?0 [;FBG+88%&PP)'9:F<.P]_LYV974S<G28.-*KO\Z(B&ECKA
PJOCL^ *7DJWH=JSE_U;]Z487X+>-X:TM@6A!@UKTF=&]HYBKB/+(BV>AWD<2:]PK
P6Q44GV?5^!-;TZ>C,HS *5$!0+/57K_2G,A8C[*_/B44H-S'#4N[Q*P8@W]#-TWB
PE_[#4IF-_9DS$PNQ0^$U$_@1Q0]:@R/4SAA4S'<>7FBU@^81TNDWIV.*/Z$1%_FE
P(/6'XO@7KI[W<U)K%$BCA8-%4'78_G(K":')CIQG3R7?JBYVG@W -)FC4"V0][8S
PB#2P,!>Q'EUPCB5:)A)OCOADO_%)5X+Z<N7KC/@IM20\K]FDHUQ;PF9'@.5C%.QD
PH<_=/!"4 HB:P[5NZ4H<7VVNN5T7?%[*$NLA)J"V8E]UP#,^/C+^)+L6B<,,B6%'
PQHW$8]>\_J7U:?=%[0\CZ,2:7 PA-E&SOEYY 4=J\F>:<=9>GZK+"VNU4!G\[XD5
P*O=9;%M9X:!* 6KP@7X&*E#T&_<QHG"%/QYB,*VJS.>H$$IL&XWQ=JK%'PW<F=*7
P(T&[^3@T>[[YW%+/+LG8J!BIYIA(4()DZ2!VJ#UL1'4Q?O/R-W#7$])>,&M5;Y0B
P#$@J717]<)$G!MN]ND;MJ,+M,20Y98!58 >;PM<@B/N0L\NQ)X!9#TA>*!-)I\ZZ
P*0B?065,1SU&NB1E,AO0NC#4%9W.3VU_C#1/[F$D27?OL7@('6O2X)"A91()SBWH
P@[K/BY(58ZDGKO)634T.M3C]]DV>Y6IWT%Q;^<^U1_89'-S[VNCT3'[2/E#>-VZJ
P+ VA[-H<KMPJP%A_54B:M-ECH^TR/_-+  7?#Y?RV-%>]4\9MX&V_94,O-UFE 6O
PF]?*!<&K,*2<P(2H?7RY+HECV_++>DA/5W5GG,3I&CCRM4T5:*QW!-%UJZ=G1M=<
P NUM@2CVM7=P'XP1AY+E-V2,T]@M/<F@051.+ES$YLSBR=M57*HMD5%-X=2%5BG8
PF+/J,^J2W;G2K_V(K ++E:?%7L4 P@9(C=*^:>E40J&FG$,_L"!*5[U'2"<MQ,G:
P]X9X\=<*!@X('5"$MW.6;PF '/G*4#^HN^B]@Q@XBZI\J.]H2V9',/]9QF02;;#U
P9&3FYQC*N9=I1K!.M@AKD%T,6ER]FLC?]=?_-;>9@CM^9RFT5A$TQ#$-B(AOKGLA
P!]B;=C'1$I1LZ8P@BM)FM<R7H@*AXI'I_*T87X\.#?=Z?,X-+[-%9L%7U'ZIE$L5
PC")P:VA5?'<,3P<UX#U#C)F%.-,CT,@T8>U!NB/N?8&(T&6)&-CKR#D64-6<&U&#
P)L^5_MO(XZ[3:FJI7L)$4P93I(AKN/;:)[W>SE3M38@(W,1X-"6BZ5<@1MFE/8:E
P6S@O^2Z_OJ2?!\=>8E"<3R&WK89E0)A U/QO@;F?ZE;;W'"-VM4)4/O54]B/$7/\
P, OC2X^DYY0MD1A#': *L;G8U?$\27]V[?2:753*FH=LE867GC^9L)'3S74VQ,K_
PFINKRC"\Q= :":,2!P(,/6FMB)2439PES<;A7#\#W W.UI(IPR-Q)\QB#1Q&!N\\
P@\J6_-DFF@RT$D+:WN8/].>62(LX&6TCN.FI..:/\5PU6@:(8O*[H[Y@)B.DNYI'
P!'OP/IK6P$U*A2?A1YLI8[/Y(F'*YV6,_[%0(#!+6XU :U4* </>SF8E<L;C65-"
P\$3#$2 ]5RO_R"U!AD !ZZ-]A1H*P*>J53FY4'!&Y!79NV/B]37)0A8_]?M@WNG8
PT2W(OEG(FHF8VF\_:PG7*'E0QB1?YB  2G-  %%^]M/F]ZWQ]3<I/;T\OOGH&,Z]
P4SW@2KE@RHY&!*B_G)OO&.G98O97I G9TT+H65)B:J&C"H?ER4Q)3;2M#FRDZX$#
PYY/;GH3!6-W'TGDKE++))+W^4](98:F0JYJ6T;.MX5\VXU%#L+N[LN9X"=P]Y* V
P=D$H/'/Y@0+QWA^@S*U:+@LCE.';<"A+\2SR'4&8E7 $T "& )8C>4A>;NMML=M_
P\7XIKL(FR)_.<R6*]X5KO-DF!ABN[O!.78WOHQ0T'$6^V=AB$<B1;_3U9P\HO!SH
PGEW>6H.>>EJ;LY0[%50R\_J\'#NABL=: %\T*)UTVH6I=&B(5-F JP;BVUQ QD>\
P@1JRM@J 2AS*E(/+@H/MU9*C^@./PN&V<A1)!!M_OY0,M0@$(MBY(Q"!$E\_PB@8
P2@4P]?I2"T**B>B[KR P#?/OGTH;ZA#RY+Q",.%ZX$;6#NY&K5[978CYH()JNSJ<
P?PEEBUES-M,O(+*2"[IX&L7M+8KW77XT?^0+AQNICM_,W7J(R_&8ZRSR<#;EN3D4
P4H/ ;"'H]M>V53 ^!N\^XA;> '5I%6^"*SMT9]T=S'O-2),$SE9?EP0_4]YP-!M8
PZD XUB,KVN1#X=V3HBK)C+D):9KX9N*A*#BLIK[%7Y86"7!.CER\%Q!%Y71A)2#[
P\Z3;CEOQXCGJ\^B7<#>=$'L[SW+-.E_0]:1G()AM$B&#AL#YTRJB>(HA<ZU<0[Y%
P1A,1,!NKO,B=W&,0"ZGNP,M4F6P"U((+W (2C.ZW^FIP9*IR,A5HO.#:&Q>7_RTN
P]8NGR=5!"%2-'0+"HNH'>_@V?%B_P1UET>X(4#(8>)\F=!,5SB1\88XJQ'!'!W9#
P!['QX1;45YH=Q+!3K/^#O-GU5@(7757C\E;4$6.X<;,N!2<V&X2WK90)+Q0^[I.E
PG)2()H-B0::G7+-7:J#/7T$5^^/+*M^\+.(Z"0S4SD'.\4-K''.H(7A:9 (W'GH:
P3^?_9?NZ#N7J?,S>-YEN<VOT7YJ^!W'/@NH\N>0)#+ZSI:$,)=[V0>CXFDZ]/GV<
P/*DG=-;V6T'0<L8)XG+UUN''805U71JOQ5.48&1/77G/! ^5M^'YUTI4)Q/_@S5"
P32<DW4&ERC3N+=1$<4> I1$B:,33Z@[$D$,<%1RE([JYP]A@==07-8DOJ-[#J=3J
PU\<9Z9"LZ!1D4!,9(5LN0QQX4[YL9U+Q^)ED=%QFL:[I)MG25D]/4/PU17L<;[#A
P<2FHN;1 -[WH)5#+,I")/T+R'S%ZD/[_04WN;<^X("D1:KV<TV*=I@E*-J;(J^WO
P@Z+322@J=+A,M5\M,YZB\/&$Q/_JOCZ,KJ\;2U#WNW-56(1&(GIJ[Y6VU!M93)Y/
P:+/]WUFYISUF":&Z7,'U8"PB-6Q5[H9]IQPBH[0R#Q$ )ODEPV(-A:<YN:LCZ;>;
P^RB*K<RRT&K#_%_-SF5K47481_[.P2KA7!TX!=KY<0"ED7;<_3CF?IO#N6%9F6+:
PX:P9QLSD<RT!'*>FR);U+'.-&9\A$VG3A?:ZW0%D=3=0$)U+YSN)M DDVQY86/IM
P+?G;8<,C5#N$I=),N6#4)9U134E.+(Y*.T7!HG\33-+/\@2SO3DY'\??]U!UY4W7
P^48LWH#X-;AN[XJMSD[ACBKZ8W^O T-7=C9K_[+#=S<>/V]E^$S[1'-^MP19/<;_
P#D1#Q46>S@OU-9\S/= D^W/F8I-X<T,K&M2DAP;6#9D/TBMCMJC^DF99.-] &B -
P)QD!HOP\>\E:!5KA2%4$5]V^D2'S=<.R/-!PW>AMCW/[%V;6'?Y\4X)*:$B_CU0_
PZK^:RFS^J_5\^#EVQ,.^NJ!AKQ+,QTHB;TV_:>4':AA3:I7<CM#Y%LP*TCN*25]C
P+I LECJN?HDRHL]<*R\JU07IGC=1'85FK68?[,41G3_$!'OA=-4U>?M[AQ8];CPH
P4C>Z.7J$1%J<5A]W3W."E/]D6\I^@^?G8+4(>I4&EY)=38;)+C/ #YK9)I3@"Z?,
PAQG>.S*_M1 A'G);3[8^U78H"^A=DI'4A1;$+Y)J#!%.4SIM):':7JFWBG2.OC0 
P^M):,B0%^OR(*,_+-9$KSDY%&&P&$-PO:N)M),\QOPC)=G<J+N[O;9E,%;ZR>D@.
P8@*S)>[2 _2%#"A)R?/*EWO#'9'5^B.-$5E@[%[[T411P.@%\,TN@!-H@IS)]/(1
P'0&M*>EE(:(Q$JI$B[37^QHT E*W=: K@P73"[R:TZ?BL8)ND"<WT%11*BT$<U0O
PG&0O+@F^LU%<"S1!^<DH(6*'=.+SD*81+//ME_\'*\,K-$4:)LZ$RLSP57E&!H,I
PQGA^G[+2W*F'WWU<BKRO3CQ?<2GI]:"\/QA3VM&AG<8?)H]$4&\O;N-:&I#45##P
P/S?GZ*H$R:2W.HW((\@'8UCM3=%Y=BZ^AI)=<TV*5+\ 5@F#%005X[<Q(:Y&O? ,
P+6J]'0P_ET.8\P K8=2&\E2 U70\&0]2QS][5NZMC&MQI"G$-.V,M=M5=Q5;-["&
P27 ..G!WC(!74JH"T+9S7E]CNOMA[+Q&%V#B-?4;^.=J9*W_SU_M-*M#40$1#<(Y
P;)+)+J.6>Z3'.FK%=Z48G7 8I%L!3XK2E[9]-63]EQ6N_+\[O17/Y^<0./(6DZB>
P'9$$+V!>#N!F)9+JSJ2,IZF5OTJ4_F;>!-[ RH'UOK)/4!.EY@MP )_*O2BZ*6!@
P X5-/>MT%0@Y'Z3K'E'-2'NN3\WNYXH9;7YB(QI?=-2VWW)O1P[W2$):I;EY%>J*
PSA3/[46]E\CSC:\J"Q[&"4;YA>D@@17(B[,%LOI@(;<S=!@)\!++CW;9UKP&!_BA
P=(H"HF\>"1Z?E83A[HI#&55".S)Z> G56OM0 7'Q!0?+OL;J7'%-SG\:NQ4'>G?^
P&GZNRNB?PK0MD  ER=2FE]H4GABP<R/UI; 7]K,23J5WUDL;=O";__]1:QWV^SR=
P.C-'7"GY9SL173D4ZX]*EQ #Z"?QB8'N81('E>E3XS<*.IWRIZPTV8A=9\;7JMAW
PM&V0#\9DO/9G&%;RNA#D/)V%)' @*6;5\E+ZFZ=92S44)QU>!@U>V0/RSR.SS8!.
PV92W#BA0'YH$ IBLJX7)YG_(U:V9Q]6R]']%[1%6FJD]6U S#$OW2:(")S-&)D0T
P(M.)R5G)\*CIGPM48^@?[0CS&<D:K@+M;7$$./_:JI\[*1)5 ZMD('ATC("_!1K(
P!PVLK4@Q)VK,/&SRI(^W>\WWTS*@3/+\,,I,"MK[A?ZZ5186DFA@W&.>KXS>DHS 
PF4@%-C[\<26+(P!:4$8.[@L&CP<J-(#Z[S=5#O&T+X+A?P#+&TGMBG,(9@^VHIHQ
PDS3.8$RCGK[]$-$5*_HO !I,N4O?$\Y1_H[RBJ=5G]7ZB@_]N<=M5<KIC!VY36.C
PNM\\[(G>[QI/02PG[@>=A)6L&M01CM)\>^H]9E)!1>J) ]RF[BS#E;A@YL G?8F=
P%0X%^RL1Q!?O-'XGQEQ?E*1\JVPW,0>_,095SI.!P]:$5,-LH-;8K1L(P7@VRFG&
PV(-0X]'/75*+L1 Z@QSXJWV9(=WBQ"1R<$LIJFB:MIT8))-!'((9:_IDFQJ_5OU)
PJ@;I+3=T?L$_ "5EJE#Y1%YB0V!2[4\:N^LT&,B-EL<"Y L"/=%49(/<@O=50,1G
PN'PJ*.2)JN)CNS&Y]D9PMSSO3$Q!1E+(R*["1!7+H6]%!?O^A#^3"(J3):+:M)T>
P< :0#<9E^M"9!?8EO.<]L+2W6MRO/+*1=GI2S8EDHBA<GF!Q<<(L0868TZY=.[Z7
P]]/Y'5L^%I-N[7W:5D@B?]Z+RAA4HO9)CC2TE&8 VV>K/( A,!^]7Y+R:(MGMS_K
P^GE[-B\:P=3L1MS^?OZ1;\5\<E!^NO<.G+08+4QUUF->,<2R@N%NB51K)_FI FL>
PSP'C4NX7'LNG4(M*,]] QA6D?S_WAO2TSOJFLH9,8J;I;]52"XF-II[E"_I!.3/]
P8L2X1E1#5X^#1AUS4\C02BJ$7=[/-1YYQMZ*-J&W*WXMNRR:GL:8-3<W0E:WD_F7
P-4^L[XFP&3678K&)A[Y!\-56]1+9 $\/F28T+I7=6,/^V?T$D,<R36$0]G;"Y0Q>
P%EGX M0)A@5S&V1G!XXATA2)I_Z*Z<R#&4HJ<0&8:/4.<Z7733,U=)H\6YRP QKI
PM<4>A;#P\W/,SX2ZD%2;P7P]%NB=.@BM85<5R1L69!&,G[(8JC^.^LWOK1_Z<A<#
P#S+5/[5+@^#_\U$%R;U6H<I3,"S%;U"JQY7'NSV?0^4?W/VVM3R-WFD&\<0VK5;I
P@L]C JHIKUCD]DL;ZT,V)NTZ:$__"%ZHH2C+-G5/!W7DV-"@0]%M8_>X]C3#LI-@
P\]?<APWX^AU$?;?G1^K$G4G?;'3O<,C]%&L*S0COJ/&EB<=G)DI =&XE8RN05)"F
PQ%HC)+&2,7\ ^:LRE_@*O *:K_:>;;<)*I?"J@,?S=0WD=5@:= 5"'<1PEQC561(
P3^8D7_A_2JCZ]HQ2&FQIVLD*\"VTT>K7CTQDM4S+%M#$2/^Z["'VW&3*/<5+HD$)
PY?89IWK(.UAOT#'R_#UWP1'7FG\'*3'WE8:FELT%PZ*TY_1I25V6>+G .?&#'KE5
P.%?R9SEI3:8172HSY$#NS[#*N-%7=A).8C39[_?1BO:YY9DOGU]&#??8P!(1'N;I
P#\5X:7\(O)^T;FIZ?" GB!QVG3=*47EG550+/H%AWNZ%U;%.?G&#&XP]8XAU?+W>
PHZ0G%_#M6$NU^!=E_[7@.[!#.S*V<GG3_V5XZJ$.;5.AM'C&,&[)#;%^'- W=4I9
P1T,6G6]R-QZ'"TY#),21R2L/U<F =U\E*J5.[TABT9H5$>]%71A59BY"@']]:+WL
PH F(KP;C*2NJ:1GW)H>\%[&E7AZJ TZY,Q8A)2C0P@"TAIP F5*M8^S93)G>Z?@O
PSW&H;VS6(L](N54A+KZ8RB/F^+^2F D!WL!O)(,>:+%-R#_/1'<ZN6&4_JM)4-T>
P0P<?QY K%.A@U5/)7$RWT%0+A$S8DO,>WTT72Z=B==TF'Y"\)X#!1YHVS-:/U\3P
P+,'D 7/]G-TT&I1$A>CT@57K,Q2*6J LSEWB513(<M<"F9#]VE\WHM)3&'<0>S9(
PGHHEH.%MX]B(PA(C589 BZ_CJR[,:3P],>)*C%,9T\ 8-OH%[$7B/->!N!1%DB]C
P/14S>RM]<DF :(Z\ AN_,LUC$:A.RSV"YCJT4W,:;D%[GJE@)C9^YC7[B5^SF&E?
P?$0U91*:M.:23R/B3AO.5U^%L,$+Q=M_P=GB;]KI^USVRPU?5?[503('&Q;W=^.0
P8BLA^_'B7>,=\=_AFL-N)H5TBN&PIP'[!I6TJD.\C<%>=$(\N$"*_RDI@6&;M:ZZ
P_&Y?$U4&6/5<GX9\]D(H9YM"=\L= SY1><]\EDUNR=*IA$;%<$@)_@=Y)W-RB+>]
PWJ=YN Q=P]>"++MC-%Z9MH3&BU3HRG=VVS;8C M[$R7T'6&\<7/6US!3P"V%;^*A
P6XBY=ZD5^9 ^TW&[WQHRQ5Y+\O!Y_X[O/?8]B[@A%].E#DJM=L297Q4W0T4$]MM9
P7CY*%[UY^&(WT;8.^E!>DR#'70?G]TE2#S\N%0A(RWU%[-5W;]5@_6BUPGGIRE2-
PW\/%ZU*R%X) 8[<R)PRB4@PK8"B^:4ZW)[&";ZK$VJ)K&:,+7S2E''(V<LX0C9CA
POM-RWEQL>',)'8R"P8(V_@720"1<G$%BMYO=RR\I4/F27RAQ_A(YC;'1(0:F1N%Q
P$)E<3$XW8FKOZ["C;$ZXE+QO##63Q^8I>Z/KCIX\?T>H)@2(K^")/-<PS?AEHXI>
PO'CC&1Q+G%>2D]FS6*GO^P(X;\JU<X.QLX\_S.%X T[7=M_82JZIBU\CE#Z@"4[T
P?@&%;)%6>%&/YGMEN&FK0X+4 H 6I*AY:DE3!3LF>\T^R(ME!VDN!9+6>$>K3"[M
PL8JWF-$2AM6AT(F"$V+;10]B_G?& '-PQOO*O_GX<U>> )N_4T&[FIQ\F@->1"HW
PB]P!,0YY:!V5GTYE53(Z+0TM(VA3[^*C.-& <2L[,B&*>(,NO8U<* E'+8 =CW'-
PKP.!KN/I)=V8=L4>%53B?!)]*RSK;QA-4SQ"BU4GBY@?S^X/U_ET76 #*N0(-8Y$
PMZ9>,*A;4\LB>^[/@+E;1$(**&UD)5]"D 'X13%_/VB*#(A03S_.$6MW:+CFHX^/
P])JE+&JQAY<WSW9HZ,[/IS2G[!I20WDZ&G%33D N::#*$PXH*FQ9AD&KH2NCCDS%
P[?_Y2C*^D[-B*VU8$$.PEEXJ) _=TQ.";1*IOZ0-#\!8Z.1F/=O"R]T+P3/QN'+F
P\^ZZL/\W2AO8QO3H-J4%1LDFWO&HS1!E#M>+.'S!9^^3'W=K!JD*0NC1KXXP%!JL
P"02A>9G')MB9R2\S\-H-'W^EK^>V=ZD7'OC:KH0IV\^RP=Q?/:ICTIF4[SCC3HE&
P*L#I'XM5T9N$>8R6>:X]6R0F>!KU+G5-%O$Q6=30._1+VLNY=W;JC!,B1M+-F)>C
P>* !"7,,9P0K#S.K]12BO[9D6IVYXR9^8HS$U]+(2U(J0.M4+^W8C/,E9$%5#M?6
PNL8#%Y,?X569.JB.X5 [K7BL$\0W59[_A/[9ZL@*X-7GY<K")ST8A@E\%K' 04V&
PAX*,ZQ2UE^E38)YV;E-C1F\4VUTJO!A1QDOZN[0QD'F]H5QG)NRO62@&%L#5QL>!
P10B@=42K.[ 8IG!F^+3;0LN,RF$<H$R?^I.U0/N]=YL7. RT4N(\)-)V-.;0LOPQ
PB1X.^43 S#!RH<>?WU3;@\HK'81O!=T]0AZ?_0JG9('(4<$!G!/'<\?.F]QIM_0@
P7GN%GG1#L.JSRYZ@8926B\1S%PO1IYU*3J(AR!TCY?48)N:R141KBI!F=<O*4E'-
PJJ/->Q /1D6;34]V'-$32ZXPW6O)3TY2W@D!#8;T8]4[=UAK^1TAF_"Y&N]>ATKK
P(+M-\LU_?\ZNL2D--40=8V3A^N4XQ$+:PN-XO:Q18>RRY[PJ",XS HVE39V9E PJ
PTH\H#1Y5UA/^S=$RVLSN7(?09D>:/1WM+CKD!1QMP-,P@.82@[4^6;R,AN20"GT.
P@\A[N-4UD E+0'WJ\TTD5U)W&@O58^..%UFOO*@D L#&<M\E^Q7VEJP3\"M ^^P3
PW#[Y/%P*OO0Z^;\=Y7T\K!>I.J!K!^_(C+,US[K32FGZ!0%N6R@"'2K!IT-DRX4U
PVP#2;=^8\$>CL-S" =>&;%B1,I3%#\^TDXO#&*,%^E-Q\UUBK>\$T,AF&%3Y6KR+
P"% F\MPA !1>@3/)LB*QY)Y6XC][N"^E3ASYHZF6KVC22[XPBYG%JYBLE?*18$OA
P!1R(76T9T+G^?"]];OI_>0R0IJ_*0" ]4RX41%$[G4N<BIY)HNBY52^=@Y1D0ODQ
P7-9D2[@,\Y+>",0Q 0$I?7P3$D E-#V9LV"98^S2C*B/RT,%/MT>40[_<!;KW\K:
P]\UB76NHG/T7!XRVFA[L8?4LN?;62C801H9J6?S TY:(BQLO(MYND2+A$;X,<-%/
P.;&2<SZGR+%$M"P:AXC.BU0CHN>>+95\MZQKH[K%C7::?32$>N_$0M]A].OG!<^A
PE8Q]%#1[]CE09>.K7N;BUC&==AN]&9!+<I,]!&H0;<1^NJL:(LG)J @7O1<$S;/>
PU%FJ-2 ^;H!Q @.MGTPE\O8\&*9E$"#RJBCK,V;%D+8KOMDX0BW @X9/=08[8&FZ
P@F@1\58<9O0/8^^KFH%,F*PU]\@N[&<:^XR+4IR_=HD.GJKED $(\AV#U1)Z2$9/
PA:PD+B93VJ[L,MKH7P&(*?-74"E95GPH$JO4UDPLRU>D,E@G\KIBA0K)/,4266PR
PZUE!:4Z%3XG=4ETTI9SE2#=K&QPK&5*2MEO!A+U9UK98D*'GR]" 6V''\&@:46[P
P%?X/H7@:C !!)U[W+;#ABL35:N9$D3EE.VRKH[6[EAKI5.1[_C_957"\,1<Y=B;B
PAZ:(AYHPY\@"!Q-D&CS6&ID"EFL6),!4[(!I&]L;/IIH_=F#GH V7"R:QQ-4_S-Y
PMGBPKWJKSKNSU^;8I#\9VA^HE$)L3HQY*%T=<5/.,;A1RC;#^FP5=N=>OW.HZA^-
PKY2=/,G_8W(- 3[2JN)%+LF,H)#90#,Q-.VC+8<2&3)HPZ3B7K0S@'K':A],$.@$
P?1YL@7 9Z42+&D2;.(OU%^//9SL@6B=_-6E^,BIBNFFEUZCA&9-$O1J/6,M(=5AQ
PL;XK>,BH5PBY-,6-&3NXZ+%T.#@XYJYY*=1"TK[_8A1HODU[:X=;C3PJ2K&H4#7$
P"6=\*$0?.[-.O>NB*@42+]VO$8@/)FIDV^Q?]<- L<VAFB3+,=&QZI3*9+=8P$=P
PYET[H3'?6_R6UW<50&.TJXJXVYQ;1 ]ZUBVJSZR%Y]A)-4-T\/J:-W/XG46QYZH"
P%!A=,OSA"1MX_S?*;C]F*0#O>SH;+=9(*H66:<_?EY1EH.M-R&0IMZF>?!PN8^RW
P9X?N?CFSE;9KY#DB#</?D:"Q^-45V7)<LV,R4;U0!X>E_*:UQ X\1 :[?-\MU&#]
P"-YP&2T'VW,RF-D&FSR1<G;"9NZ[I0.]<S/+L*A<WY(1S;6V16K+^)5AKDJ#A=I=
PBP="-5#1,,EPJ%9-%P<NRIMQQ6-)13EX]A5FAC\4L&QQ68_R\@@^^BMA+)-\=!87
P%EV+Y4?+5T$\C?TLSO96I>%E"]T_=(]BYE9E%-P+Q*BG(2.8!"I^H,/;&=C;QU*9
PR=TG6G(SM *Y>%LW=VL JT"+#FN<2USGYG.1?[Z(2M9G=(55 T7IGJQ'2AX\.3 3
P+. XG*\('*G-3S0-N=@O8BW1BWSX2%S9U! 59@0/G 0R\%D;DC"2GH*+:=\-I?+.
P36VQP4)S<&MP]<U-#,[%F"_CK5%0QD*BX8[!H*2$W0QQM]R\F\2.JY364 W#T+2W
P(PL],[L#4?",-7#(8M]\O$TL>]\6J^1<W,W6KAY@8\[3W5UJ,?<RDEA@MX[E#T>Y
PN5]?\*+<*_$\WXP45_W(DZ4%7 E'-HI*6P4^C1A[V!$%9#;O@^DQ1)Q#1IX8N\(Y
PE!(XQ8/YFLHO^J;WRG"U[U9U%<R2?]L@!%+8Q&)[D:.[1D6RQC]^I".632-W1P3@
P_]5VI?9ONX%B**M2.A3H-K 9 AM(M^?LZ>:>L6*26\<*%5G^BE.$5A!8?ZE4#@,R
P0K8@&! (SX2/?H4-T.4@HYYG@41)8K\M1(5/[.I)*=F TNT_XBF9TN9'"GF69@ G
P>5][J]_1..F$OKWS]GTQ;\ZBJ((>1 F04THS9DJI>E")G3 W0IU.0/R6B@M&*PEN
P;.@T9)@U+_&?SDL #^HG!Y!L&@.Q2_Y.9C=6%GP'4U/WBHR/71+SCET[*X%QI/!M
PE8=)7-\.L<W,X3GFJ5N6X384<YVS/U5# ? W1E3BO\]I\> YN8XOE$G.>3PPGY0@
P?N@^;HVB'>ZG_05R%.?'L+GX.22<)0->1* 6]^P".&_'.K#4ER KJ0WMBR%O4NVS
POS2,>5J*Y'I\>^Y^+IE%U6H_ -L=<+2;^ZC"GSF?R#B:5%ND'1YAT)6\(^ZX&-E"
PMV4AX Y0,=>0B4ZS9^L20BTU=<IF 2982WT[5OZ#RC8IIX&F0O.XYPN8MT8/->TM
P[B?M1N<J77W?2'"D;U.W7J7SHKZBWY&/1]X<@C$(VZ=?%3,_>6![0+O=;[I_?ZCR
PJ$]AL?+[R.5%CBZ9D5=&U 0]L@[33$(K.&(G>D,ZI-WO>81R]=T]5N7X3YW[#B,$
PVC1@.D[126L<8&H?CJKMLQ-PI3T:/G/-3/FH7!H,GKCC6:!D78W]ETRE1P%L(= T
PQ0;WN )Y9,I.;;/IPT8G-,'RN< ]N7?-10,?\:3!%T"D[1MVT39Z45HZHB/J,P=M
P'=8M?MHJ*HI._W+@56-Y3R+&46QN4&FDD0#IB<'85T<6I0U]+V/P6'*?_EW[J,:2
P.0MHI[0D1W**[D]4\?X :)1*%,?+:0W8%YE(^OOK5BH!WSVEG:=1&/._3UY"7L?W
P2+6H#)_%9@.$%_?<6C S,47DR]-W1;1: 3D>GT"\-DT6'1[<$I<VPN>K.J9P88FP
PT>+&D%6MA+U[P;GNJ'*P,CQP%Z3W948]P*GJ4(T<?==*GML.Z[,XXT74SV(KKV3@
P-56Y<D4QN;44*V5S*D>(6Y[[ZT]_\N$BL'N4SZ^GO4"Y6^00#WI[7!<'9:CF97-4
PT0N7K?NN<2=9,)PQ53TN# Y32B46Q\BB_UA8>^ELEM"S'DM_Y4Q54@#_[2ML '11
PRJ5'@L'1R9:F6<4<32(<%AOWCWJ=D1W;L2?U"4TDT4^2.D_Y>,)89!P@[8LCCN'.
PJ8>S&&-1<(C-E6T?>+YZBB9*F:]FP7HCR]IB^I@R8]I>(]PQ&4_CW&G634*PV5N7
PS\;IU.A+*MWZ8 1^9M(39*V5=L,]1ZAIFM9M[@>5#AD!06A8O 15$G=!>A)NJ(J)
P24UEICKR]@< 6N+IC[^:/7 #H&E_@($'_9I%@F4)D!"D_>M_?,#6N+(HI-RO;X\S
P87"@J6=2:VY[Q1LI7?.5[L&=>T+%-):JG<)>"?O]*>)#[UC>#A-[#%$^GF;UF #7
PN809>VY9"-"74_;?ZLQ'&-/!'H1U6LV%U>4S@<,F*=MP+)DFA-.\\!IR_[.&1O'L
P2)+84$P@\L0#,K1F'%&$N*KM3>GK*O8"3^ZF=2DH!12@P1#B(TW,AFO5&N>_?Q0<
P[*UA1&B>+<"L%L45&P$_O7#IO-E==GP;B'?UN0[C!C)QAA8\,@3'JZ!UK)I$VGQG
P[93)Y1Q4N7B[<5N+XK,$0[Z&ZR#OSF5%9S.7Q(2NGQWS%&*7X^AAOOT+;N.(H0Q$
PP(CY3-.2S>FE==X/&Y8#;5Q<G-5:I03MTY*K@A-CW]DI/*X]6H8],/NS(Z8PJ:5(
PXKP&)CQ>(^7=+^)8ZCZC*#X1 14&_/?1/-GNQ(R]F5=6&Y:CAAF\-:1W^R^Q%X8;
PA3&4$LBP)!.SH16SL=+'ULN,-B[15G29T<8[==:7&V4F8F+=V9Z@0SSM>8'+K ^^
P+6\K'@@Y"?C>1MLO0C)/T2"3SS8!%/W\>D8[2"K_9(L[\99.!S29#@]A/0XVZJ_%
P.!&KUN]1M!DQ+S;$@EAZM1UQ0XMQ$7J03I:0I)$0 'PV58'UVHJB%QWG4?T:?H=.
PN5K1[N=?>6$Z2GQ!D,5)Z-HBB:DI"H;.^)#IGGP5\(Z/#1.WU65I$#.<$:$:YUR$
P"Y0S]GY]5KI'][W'6V-83T83PJ;3U7!_T1Y@OJ35<5W[%KT,R1U:5NZJ]!C)ZMP7
P"'7D]PKA\7K1H+G9PEB%[6?#2B^,:_5A7\1OJJ)&9)&556(+)"52O1&G7&3_->S3
PPT8W5:>N0G/W5Z #O1TSC8-Y]*P"5'#0-NFW6K='9$35"@+->(8:Z<G@N(U7J.2N
P)IEO98'A%MXLT@ZTVL+8()3F@XK;1=#,Q*L$AFUXC9_K+#HB7:&M_#*$P)T>_!5I
PE_9(.0*B2>/X"][!#*(7.&W>*I?[ ?:D8U^W&7>\<N(,T"B1L'34S\O+Y6S*]9Z 
PL<@6BPNL[SZ_=\"M3B1H=?_OR4K>1&#@>5_.18J9E<$LUJMAQ!B_,ZTHTV4QX_$T
P6/"GB&.=T:!RB5.N&3C5>#]. X(+RJXH=(4:'-J2=M?(K@?RX#Y48X3M,?W,7BX8
P.>,!:D@S?#;0YC+!4:4N'4RSKTXK]!__SAMFGQL/H[;3.[/-[=42H>CSRXZO _V.
P-;ED?^+Z2I3@;0[&.^_4*3EI >K]1LC\&Z?_"&-7F7'F\ZY*!&TG9C@_![IS<G!2
P"]R>,)F@B*3+]#%C:Y<_=Z6KD[(&,68B[S'6-!G?V*KUJ7['*>S6X7-7\OH0&C^Y
PQ"XS(6)=)S[-6Z^YI&[Z#J;F/8[?M7$:<\2I@LWKL+@8*"1L\TZA1553(K&'ODA$
PMH&K[:!SDD%^;/55*\G^2W-; ;Z%)%E;KN'_4WXG_ZA#R"@_EV;-C,5+2W>?DH<S
PZ6@Q??K"O^L(R\-7#:0@UE6Y3]:,S$&A1)(,65I6I7U]6U<.X=!IF>2S+\</G!>;
P/<[B_*"N;MS)XMD^V.(%^@NB+1PF^".)9Q/4WZ(YD\1,*:[//UXD;\T,,QOAE>-L
P0V\S0\'<NUSPQ5T&_",#L0.2BQZLMS#)>1\"ZETH$<"&Y9=F_1^$0P&08-/G\7V6
P<T#H&LHC23NLZP#R4 2@I!$KC8Q/#/2H;#0J@"R2E_;.PI838%/T[=<ZMDW>+HEH
P_H/N#: ]@-%1=;GTST[*MQR'+D67>OX@$VFEA2QOPBHY1@#EV(N6.$/=7!=26E?3
PSRMU,:6UM&H=" <WSG;8S@4^6$6/NM]>IA=72KH%^=#@J6^'L+[X"L[KJ8KIM$[P
P8EJU7GB4PP,*0)[?-NU<8!@U* -E@E[PA_.NILPS%^A%Y_54-F.JA%PDL0Z7\:6M
P$N>(JECE,1ZJ5/_J%U*+S"U"V0!V[,N.*6R&M%<2 4A46_65IT;RH:7HF^1;8$"@
P617P@K6MZ(O_5I7W*7H@2OUNK(P3WDPBNHW1SDE%)N>G T0"QZP@'*PU@78<W91&
PFTVX-WNGJ!<TIDFIYY=W837B@,(ROGT5JUND)DH$;XV>9S?I':!S\+>[1"4T+-=G
PJM%/=(%=JS5JQ;X>G*X56X-OFBM.5&E$5N;5!*5P_N-F..]=?8SIJ:2N53'G#<'?
P6+,[.O5=7>LB=(%'PQOK?AK)WJP4]2&.24&VH/PE)'I5(AN5L_Z9RT!KU=T]W;_@
PH?*[GYZS/:$P#)>A$O5:F'V\5AG2_O_2LD0VTO(T&&C6*U#[-[%N#QFW6-@E/V>1
P<8GYR.W"(3(WN:M1P['^8*=[*B"A@4/U),T/E^0+==6_4R:*V?J>.7+<56H/6+6Z
PL3A 7#A@AD<<3B4<?%3G(&#[WC*U5?L3F=FPN6I&NP!A[YR1H%D$(\N<)9_-WR+V
PPV)C?3!RB7,_B>MGY](JWJ([J46E7/G_KRW(!79>#_BVGH_'RQRDMQ;,+H2Q1% 2
PH9M@)%];Y"?:9RJZ;#I2LTY3.)$JP2N1RL4=,<M>7AA#&,O@)?"<&!T7*Q3.WF04
P/M'%A&<55J#9Q*'"%W?LEY]S(&BW]WJ$T24 ]->Y]<&TF7E %50LC71R*GR21;DW
PO<FIO'WC1H%]+!P-+7'/F+50,_YM:P)H0029:5L]F::!E,]??__2VO?*, WT'TUW
P0,A6"D_VP$O(T87<_HX%<&[_#^Y^LX4IL#LK92*^R^N"(IFPJGC/W'&A+FIXW/>_
PZP2?\@$>C?S /:-G 7^D-H_L/(W4<4%PBS3:4P/ OE4H=QLE7##7+^Y=Q+%9(_6D
P7=PIX?.GT(Y9I;]LX[#3'KI.C>)(#E%[GI1F;Z7$,,T,NZ%;/7F0'=D&EM!6/0"I
PQ\4^=\_Q=AQ$:>)]*>LM.!\0UFND[@I84PA6(F/G(>P1!^6EE8T.[FH.+K-2='. 
P_XHQN0_O55F51U%Q.&:D)&;-*AW5-R)G@P;D6H@U-8%+0GZ!LIG:22+WG0\J2>&T
P9I5K?J ;S*28/'J@TY-D9XQH_#ZL?SI&/+=/=B,B4CQ\D'++@?$W$4P0$>CN6\HW
PZ.ANN::$&#<5A&7%TBA&+Y;+>KU:3JY7J[3V9M:0 60^4?PR]ZWH(/0<:DOZ<A2.
P7H0_L*OZ\"6?%R)Z#LY_UB4AV+4X@,=XR7,%W<Z 7#0V#?Z_-*38YLDV-;S?GAP1
P,5/D%V->.7MNCPP3AP7?[S%2EFGW_&<N 7FKF^O"^-%1Y=[J3<?'7QPR. RTH^?/
P\=X-P;=RV#M?T^7"9DQ/$";R.,B59$N(E%.?Y/-KPO'(%/!8-75DS>ZCW1[9ZL2D
PQ66E6A]30HXA#!&;(<7YD"C3^>MGC5*I?2)"[)U+H\/:5.ZQ1/8B2,$<<[HLQ'CG
PQU:W&9$)OX 6TV[F(!4GCV8JC43G4U[S'G#Z-HB+R77"/]^#5B-L;87(!ZG*&5 ]
P/SB?OM!W&FFB" % -NZF !'') OWQ;[E:$O5&[09E'K51_<O2VZLYA!=26&\L;#)
PK(>7(WIJCWHI1W][UP&<;C*G15@KQ%>ME+U?%]F=ECRD^2/H,QKQHVV_L^+5D3_X
P*6^V=(<=?&X/$_G=16/@2[3B<2BEU58#&WX9O(8B<+75P'X9,=[6%JD6!THKI7=@
P(1DZH*?-4VEPEW.L!SX_Q#\<X0]>_MUD>I(>7%1FD PC[29;D#.6U[(ZO8E!8JNK
P_70@!U#B#!3+)C"5!3K&RN]YDH;3LIEJQK J&2: -ZQ2ON3^Y(=BF=@(MV\W@">S
PK+[<M:[5B)KKLKF(\\V5PGT*YGCZ$TDOZR&%^8N$?:ELU&(49'$K'YVK-B?ZG@G"
P0+B$8.[5Y^ ,9_2 Q#NBH942I)4E=%Z1NKL+]LM:N5BF( VQ/293V^T)USZ2.WA+
P>3_W>V6$['[K9)Q\F-1F +HZ'R3J3\\,&<>47"?E/\K4>S#H6$Q]^WPES=Z*PIJ;
PS14#\:4 YKY@X(OO)ZP6T+YTL/TG&,3XB@2@@_;//GY85"HD]\XM?X#<V][GO=?(
PT2C5U)')7@!9$LM"-C\LU>C)4P"U)"*%]J8&93A8'AO\?ACNP/G7NIDII,4.-D[9
PE3%@VTF]>Z2XLU@$=O:F?U^UL$920IXP"":V_:$:JX&S8KR1"%CNL:IW\G5B6T/K
PYX[J0^EB52-@BL#%;"MZB2W6@78O <(:GM%K;-_$_AUE7N9,O8_GZR/AGI'#@/E:
P,5E_Y]V 4\:WN@#.26,IXG2K_K(@AZ1(8H @"!S2C,0=>.>^G>LA?S">=N?*;/Z3
P9>]1$N99Z[]4_3&;Q/Q979KJ1"-\-A40B.>K\D*/^/=B,<I.@_,ZR1';JO+.5:$G
PA](";8("HC^,%0F7[V.!,HTY1)1YJ ?\9ROS2=%U]?%&:3]6%K_F? <5W,T_>K!G
P.4>+__+F%BV'GM/&!*KQJ$GVDN+:[+K,P8G@K$?^QQ"&=JX^"R<^3*]*Q09P"9>N
P;2__WKMTUUA@P'D%A>B89,H:"D]*V-4O&0*RS?0_$[>5AJM #E'3P8S>_;,0*_1F
P-K(/>$88\@A%L+[>T1QK<'8</H<O)O??$!P'SVN"ZY'4_$@N9\>OZ?&E^[\G 56@
P*+>ACHK@+W!A37G7$A1+=HQ$E#2W_/R>5&\#K9"='\R.;HVNL53UER@!%WV$W;?D
P0%NJGOF[=Y*1@"&G@WB?R]Y?L?)5\/9!]8A9_-!T&&:*D,12=5;1'+Y2R^(<$!-&
PSX*+%B;$^S]TXXDXHSR=*/WY@0-A6T!KNSU#&>^6.:ML'Z'E=$"H5;H]!/4'",PW
P;'!8TW30E$5*S6^^1WT#+IGK$"O@#Z<K'0)4BJ]839W^$^";LJX;2_"-+B,8:WUA
PJUH['"(LP5GB9D>$4YYRL@6C31LN73;4!%)[ =3'FW!-;Q_ D.4NH%95S'V,['^X
P^Y<W0M\3>ETR#A1Q!<@/1^A>&!FPGP:RN+JUOK.54A0LKOI(?'3-Y7':Y_#8ACI5
PC_SNO=FU-2KGS'+S5C 37C\)UJ%,I;D[$238U,,5ZICL*W.QLGZB\M.VP\5R=P:>
PI%.MJYY*027_<$C,V[O-:>'V:@PB011GC_^H Y&P-[!*,MT_B_.$!&O) 3TA9W"B
P07_-J 6FDP7C Z3O;EK*&>E60/XJV**84OYTW>L,MOPSN=RQQ4%O'3M>.Z!9Q'\1
P51SPT)%>25VUB8 2\M20O6UW[HG/3.[@*IVGRL;-1@/ N32>86QT$--;$4C']O<A
PM<4_F,[/+(V FM!2?1(1,[.#_/MEV%B8R9+O'P5;<">-'-N\CDPO^F9A;H&+.[AR
PL8$WN6J7C\1%%%[6FSSH^C 3H28$USP =).B+@H4M!90^2_&=T.T*7=0^[9:8C^K
P;IH#,D@ SP_G0%VY$VC?GT\R8NZ%'D^#=AM.@$BB'"&^YL'4&Y: <RB+9GW[/WVM
PS0BCK=A9M@$&8AZX9##5*RYL=,Y8X/]M,*)+,_*/>X &]'I9OSN.4=JRQ:ZRQC?X
P[+>B\WIJ;_8 'J?HT$Y' 9+? C7Z$.^P(+B8.&J>@>-)=;[&=>Y&W&3J\G("_YAC
PZTX;G48=QS2D\EBGA)RBE(X+35-4::M4DC78N!QW#OS*^H'OEYA7$828;\"#-PYT
PA5^KM$'>J\^-QL@OJO!NPGA@%$*SH\FDB"5%#7B > "#$VD#E+%DH-)1EWLO&6!O
PZ(8F:XI4=%TQ$*<0N%?.M'% );5>!-0[I^H)BXRNYBHV/&'$V;E]!>MZ?$[DZTTE
P7)2>L2H[*(;&]-M:#7B4Q_)=%/Y\W1HS:&B@KI*T)O$*GU >W.J'<F^6(@&7N'2G
P1OB]&F%)XEK@G;^%<=!+CU1X-XANA"\?P1=O.??-.4^?J<U/YC<( $NV+_+MSC87
P'-JY>\-C(Z8" +3$542X_&2VQVX?W%R)WV^(]Y#CX6T9[H@0SD(!%<;L %Z_IE3<
P<6)$#9P>EF"4Z'A( DQ"3D9D)5>A?>]P<^QDT!0VP&)M@\GWX4CAX87_-&EU :?O
PIA!4I%-^W_.8EQ)UN$$,_--'\4@L49%S )I9;$/B1L@'58]M[/D,2QQ_H1B]S 3A
P0W=0\LXX:GN45>KB?</=%?B81RWR]$@\=#&\ZX_LOI3$!S$-,3^I@0#:=-.713F]
P,A+Y4[Y9-.$42.+9,?O2'HIYC2C!R8A;+<+>2"3*Z'!(D8GYLU@%XD]YR@$T6X]O
P)+-R91PWDP>?M#UA[?CS=F= 4@Z E<&L7P?$C[4L9ND>/2>N9^U\P=3#+0AED'U8
PE//X)022]UBV6!<XPJH Z/%P(Z]NI^I)>L@!@_>)?"_D!7\C!M&,4V%KV^[$T(?,
P,482F*F'AJ"=4"*B7AHLS;B"1_T!;LX8H,;28*YL>QG.RN"AOJC"7":NIPB:L"L9
P@0;7ZQN"LAMPJ "+9H06*'@$*<FZ3AXQ8))!5.T%Z+XCN>&GSZ6]=$D\PUG8CF*@
P\J^5CR3+9OH_V@IM7\M=<5P>2(:%!>;K*XR;$#0!'V)S"VXD9+-#(.=T0A'UP9RX
P=B4CGR^0$$>A1\7JM#ZQ2KT/_FC0D(Z!Z=0J"+WIH$J[X!6\2E9&.^.[A6[%18JJ
PO+T1#-AH21%1E/\=Q#O-6OYZO4V%E5J:V2Y @,<6 5)+YR,)I*3?38C<'HM^R$D(
PB4K*NBF1&&IY5CSL+/N9CD=ELGUN<<LXO$ZV&A^E"WG-_?#+9-CWI>)M_,V[WZZL
P)2!/LN',C#%"_=0BU[$'7$*>@K[2>.SB*X:^ 28:F<)ZP9Z: ;KN;/PS_P&XERKL
PU';^?(C@3*QB]&. ;'(75J-4](S3I0?'OIAUY+Q1TP1W@=K.%55Q:H75^ *6UB2A
PM<-0*.K&=CVUG3L(>,DG#W"IP\(THD/\N/BFB&G0ZX\F7&S+4E<_.#PXJ0OG0/"[
PJY<0EBKL,;!]SV7M_YBA>ER @N''NNXM]H4<2C:$^)9=+IG'#O;(I=0%'S&LJK<)
P IPXET$:1F0\7!L0N\,!X ;.)=(-B$F3=*ZZ^:KAOGE85?"ZXVQ_@GYTZ(YU!=GY
P$]9+-4>D8<^'PU]2C";N26 ^\/VW-QX=[3R-I-L1HJ)OWT(52 5'[8JO+Y=:PQ$G
P43M*;T(7?*5;$N/PXV.BZAG,VT>-\C?F%%5U":%YK<MMZJ=:55*!&2B"Y#I:93_B
P 6KKWS3LB/M/#[UB@KZ&%VAU0* @QX=+ZYC2'_E4NI(T "2I^AI(QM3!Z'S3R/J!
P;0"_"$F)7?V!2@[+DT,: 4 ?76'DRJ467]HLQB]GV2^MW]KF"L'N3#@!T$KR"N@(
PF.;M*MH!Q49OS%,YH6-H/UGJCU8_P$!W1U9[U><S9%"[J-Y2@KN_)R+$(*-L7[@3
PY#C3C!L%@:2.OLCMCO)4L\< EXBZ/JD_AW]\B$L678U87E^U?(>82V;![RDS$.@$
P98P2W_/['_63A7JJP'NR/^J(S.)&$=6B'DW@G!F*B"LKB:-G<@*E338K=Y4"([[_
PS/JX9]JG._]QIP=87MG:7\=#@;WT#$,K37Z/R22WV/==(2!;+7V&IY>,@4.VCJ98
P.'M> 5O%ZME8D]N$;)3QEIF"3S!%U[J_:29*Z04I!Y]G*N_]5[,<]=P01R]:D^M]
P"0-'WW,E'847RP]?HY^]#**(7VSG&8W(25:<OX\+!_(D)#1V&S92F?A3M!@GX]:'
P<K*R:W)\F^QOW$0AT0Z_9=:C=":>T'@BHC?T'$@5"!45PG6R"X:;>) !:2$/<-T)
PK[;(1;,ZOE)[*X<$,?%^]N!#F-J)EA%L*87>11'),7W7=Z%B#,HYDY+ OM2&'4'\
P6A+2JWVNOO"/+QGW/3(^B^=(W!)3?F:(NG9].*?\I$ >(9$<IKJ^*P/,1B-KVT[D
P7YTFXH7),?!_6*<>%TD)65'Z#=_#EZFO%^$3+Y5^HX:T)8":&Z.]_!II>IRDEU]1
PP_DI+XOTB$)4(REC9"*3+YMK<UK7E[)^H.T\,+8$C\&JL85G\,!W?J/E1OH4^,9]
P*6O1(V$S4*?9GQ>_'G5+B^9(L2@-G[PD<@(YV-!VCU99QR6I)D\ZJM;,X(Y9E>DJ
PLEX=%$MC]S07JP'^3Z/QU'%*3//9"XMM!F@)USTHH?BUM&]L^D925!=VUE^AG?6E
P/2FG."/.\[Z2\IM/M] RA/"1T9</K?[==*DGWNV)Z#=I(* G4*[@F&BTYVO=]OX-
P4RB"!A)SX@<>3-<'$6HM-AJMU;A3/H^+#T4+P'"X +Y?EE,S-N8]HE5>W#V<!8@9
PE Q>/3O&!DTL8$5\D2H=1= "QT9_1DZ5$932,ITJ],-.K\4\T;%2<?47QP-_6^-$
P3P;6W QKC7J1.ZWUDX,0OS2HV$"7'SNO=^PFF\&0>I<#UT)X]_#/%?90(L_R\J)W
PA36/=[F3"ZI7-4IB?> R? ^S*=]>2K$/-U%6E9!P_29=@%JW<VM8*2U>:K60_IWJ
PKK8"_/RZ8FYI]XWG,41PV:$S,.=;3$UNI;1I^1Z*M-4GU%#MU_"M?;0IV?2MB&2$
P"+<$H%(H*'C[^J @8S"<#<S!AGO=D0WT_!7EU0@):ZIO]OKP],;X%,_ E= R25DV
PJ.S]W2E%<_,='/\[U\GGW!#V2?GJ^BC1TC\.!:-/XFWC,+.464538/\/^(,!8YR4
P&,6P,#EJ+K >W;@(JPI?YPI7C(LHDL!N -&B"85&S0X#P4,[*#+CLUHN,68+&0D"
PFC\I.WVZ#LS=GH2X^TOQ^>AHOD()%XA 5'*G]!M]RLS!Z:3R&7""3.7/'']=G,2V
PH)]O'H>TJ=B19-M \$0F#>A_EWIF.H$)O_PF1MMEY/O)?412=ZH9NUI"AC+J2*#,
P?_69/LKY4L.*6774L8*) ]((!LNT3.CV^[8O(JNTTE7YOL_\A!/8M><:N+3YY7%Q
P@0)^Q&<,W=O2O$,]MN6K(79]=77#J8[EU2,W,<5"#BT4:G6^4J2^5A3]:<R2:..6
PB0=HSL$],8CM3+ZN2QG!=L>2[[YWZB8&)_6H7[P\^<]K#:@IP\X>>Z/6)P*I@'R6
P9#S)0"S0'./W8K(;W*]=LYI<<=2NY"W&J170.-.C&!YV@O4)D])K<#K'8/;:$NSD
PUJ:TI@)_!9=_>W?G:%.FQ#W6=<,ZB49 ]4 RQ]X,7$QN8S&ORI<Z47LY\HB0M/S]
P:#8$\--E>ID-O2=+[>..Z3M,CH#7H2#R2+#.'ESF-C"OEASG^IL(-/9U]709KT9)
PXUB2=H>>)8>!9V9:/>I=_.D&>497UI_#+PTV=4YKY6Q[1H Z/T 8'1:&:?5F:>'Y
P4;,J&Z<,@[&;)&\;DP:)3<=PV]UWI5TP7SP.CEMZ,._ B0/.3?7I :O/_; K3PG4
PXPJ=L>_4,=YU^J^-7:42QYA(73478>H4'CK&+[5@.#0$%,@Y(??](%$K;0?+(FUG
PB<I_B/?4C=0STL#N^9K"\X2Z&^/H?++X,5&'><52,\BDZ40 ;AD#0OS*"'(^K-4#
PAEU,V/%B\#YFAR>%YT'4A$X:=UGT99][3J_OTWV,:]&/H V*YRL:\Y,=X5P8Z^+8
P6TUATX27P.0MB2F3K-4==77$V8!6U\?%*+#"^'#=?<"*<AC-W6FZYJB0,&1Z4/@)
P.?5E6R#9X4N!#*:E_ED^ <)P+5CX*+ZVF_LH:.YU9]U<.ZKI3=3B#P;(,"Y(^Z,2
P5O=EMUVV4PXTA/E1L-?R6NEKZ5KBA9F>XE:U?CEY&X'Q[RR>*/7T9\^9KV&"5$EU
P68Z,&NJUM)GG?FD?Y0!R)F"9E\YNH2EK<>U/J&#*@]79B@%F81+8-#\$&X3W<GQ>
PVXP^:$O'KNG6CHT< $L>Y^A+0LZRFO9 E992R,>R(OJ:Q(U1&J2?+5*P' MZ#.A'
P1/$3Q+&%2'1NER]P:*@["@&];Y:F:3W0XG8..X.JB4*:YGX]>=-_?[A<8\ [A&OJ
PJHTTK% JP9PP3%X$6TUBZ<QVPYG0EM).#N;212?UM=02D%C-%,RCU#E+Z">V4(,Z
PSF;&;8V:U8TD=>T6#3D"FT=B 84_;AY<!FR@.5\J[<]\].7 !K7G_5Y2K+E"3]F:
PVEZXR&.KFBD#* R-/UCP)=@W\FINS\L^)VQ:4WX=7B2]*[A(-11TF-UGSX-FPXF<
P(HG#=>M$5@+DJ>0-#ABG?449_+C56"L!<O2X%C#*%D>'+Z\9@XV05PMZ4YQL )N;
P=,[[;#H[D9_,*+"RWBE_*M7]C$*!E5'J?\80#O(%8"IW-\;-2@4RM"OB52XO4^0#
P'-%8W"LO9G'_*(E\"]-7W7\H5QU V1U"R=A5LQ[43=>SI'B&'QY8%D@IVK::#53-
PX-ZQP=E.'!<.;SV?O6-O\_+(SL^6JGENQN-,=Z-/12AP_?]ICK)R@\X*$!86/.'U
P,[J^4D-"QO1.S7^1;Y;I>;L[.*I'A&&<AQO7%*1TU)-++?Y&J0]:&MG' +ZE45JC
P+."\K&;OX5+X/#KCTY5]PMJ(?'X<*"QFP9.!0,AW5;%IZW(*Y78^ /5 NH'_NW[1
PYCA0A).*$O;UO]1R2D\5;/4E:N5??)SWF96@M_0&]&<JY!4J-C&YK$2,_6-</DZ8
P"#<D?2*GV"K\JEIB :W90_H)S=R+Q,:QWG8F]#61\8S8(B,O]NOL'=+CXGIN[IJ$
P=MZKKR.KN0*?B$*6B[K\\ ]Q-CEI6UA^"PJO01)S3R]4H%$?R]:BA_'*3^U^5J=W
PY??DD=968&=Y_Y\$AZAB-/P\E?W:,/FE1[>NT#XDZG&/WT OZIUX(23B()>Z>\G2
P14!94P+LNNM:/)B7G\]?6"'IXIM5:YP(KMX@"0$J9 JK^PB"T)H.:0&"PQ+#)@T>
P=C9&G>]5QM!OBM\L'^(<LI$HE3<#K1&JSL)CU0&SR 5(VI#];![FE7)N!T@@:S3,
PV$U>Y1"'$3[O^;!I1L8_DZA)UG?70H?_ZULXL061LF2J"J)BB=R.8T=1L2_=F4L;
PHN2'(5AX/Y!N0SXA;U3D_JIXX3U"OP<.N!<H\/3"!'SB'B)=:A'MPJ\FR)4C)^04
P:%%9S*1=HA^J:"_/G8,!)NW^_&,,G:A)?J-#.Y<?2LVS$:59-8G5@V1I;'C'P>4.
P7MT3TA"H6Z@N_IT"Y(.9/![23)P. I4C0"=A!TWF0(XTKK_ZPWM@GL]@6\_%75TP
P@T%JG[C<GQ^W]B0$>ZMQW-R*T]5\VT0\"I1#2?/N!V;O 4J)ML/A/96J8SZP<F7E
PXT]JS9G_]R!0E6RC[P!5FW6U;E1Y!PG'G,M7\Q[E!N#FQ4S1R&B>:KS'TG>\'I4@
P<4XDC#:/&5]>4,S6K2=3;9=N>S4\=0L0Q!4)M,'[]TKM1[F40JM+!(0@+P0X_FDC
P-'^$G%A7GA,U1(;'KMFM^BU&:2#'COBAAP0]3!#<'_#N+V2OM1"N5+T%X#E$FN<'
P!#Z1+CZBQRK&>LL,<+'TGQ^/O[EA$*^P>KIG8HN#=V&#5&=G')WS<[%D_1!)8(]:
P']<=MNXAOW>KC&@ZW'KU]5%^]HP]&*V?+O;1^9)VP2([^XK/0J4J9LL2.SA])U>#
PH2IO$TR@PLR6*=HL:][T#VF30A/&EE=!A]1KAY^!Z=U#UKF(TM',[<IA-KQ&1Y!P
P#X0H[$WM-GOC7OI5PZ\+I4@JQ(;XTC;Y ^?X9.V%13$+K_H)%F" _X16Y.I%A5/>
P!I [H8UFVKBSM':3H(#806Z27];EO4"B=@L?RFW(:>S2GK@8Q4; ,><\3_SPUI%D
P")<##Y]XK8_BE]=F+I]@7M?<)J@1Y)M9Y#TQZ:E)HS\T$UTGKC;M*ON(2.F74=(Q
P<6XEM)Z__H7R&7:=(>2_8W9M&VEE4I4P0JWL58^[9 18$6*J9Z4BS+W^B0];XDUC
P,A>\I?_#0 3SG/+K9N>VJHS@I%YH8)FM1P*IT%%]\-]6HVY%J/K3PW@#DKY(3]/#
PE7VN3A0\VA$LLDQDP>?91A Q9\FYKKUS1&<D'NGB(IEZ@?LJ9O[RL?*HC LY )DI
PDOI;:#@0;#ELM55ZC[AL6)@7Q^(!>J?OY5-KI+C/&V2[4T[5D'T8J(;'<6IX4B:[
P#B9)J2WD=WH3<,>#6P=.".$7]QE1LU/_LHI]-&_DUS?P_%[CJ66F+Z\6H];77:#/
P=7M+;FN^70:^*[7*#;1EOOUFL6N?8$VXWFQN;2JW%ZVG$9GVMEH==-X<L35CM_WV
P&>&+94( =!%6UR+)R#+!N4H-L0N\3:/)%YO+ XN@"4L@K1*-1X33#74M2<),@ML-
P]N#4<&5/![FDU]4W@2:!*I!0?.9F/%)]<(JB.<7PTW[G]!7B&A-CI8> '+F%DFOL
PDR,U1B/A$>2@9&L175.&J;GKB*&M0W/.C\K#?9VV"Z%I53D &F?3.WF%"R4>^60-
P(F7>QZALFL/'J?N+QOJ>2TZ>2ZH[^Q*7,MT0GJ+Q+"-J,JF6:G>A*'F*V> *V4!'
P,J4%Y]-%GEG-+D:5"OG,OM4,/#(E&2SV[JNBZ/>-.EL;E-2BLP4YEJ\(V);>"(2D
P+2MLA2J[F.0ID:<D_UJ9H^.9N+NX-9?".Y[N?S?N98OAMI@22.^">-GI5'\572+H
PO[FKR?0YXU%R@4Z;EUVPV87=-1VIFD0]D(W!;?3ABK'&^4=:24JSGH74^3UVB=W!
PGZJECU PB$.+ G2@L??5WDO0S<ZF8XE5R@/^&OZR)4L>4]X_!GTJ_V9Y'WWUM?M]
P\&14;^9]Y#416M#87Q9XG+[?GUZ"$617NB#T_<%%H@EJ_.M1D5+Q]G>.0VJQZO8Y
PRG.U2841$T+^TBUQ&"<!D&>67/3Q!^#Y>9XE6M7Q?=_Z9C%$X.^[FA?]7)\+PT;K
PKW+D(%A% WOHSA="PS=&#05H!';?3)=R7[UR!R\*+J%<J?T8MMUR@AW=R@H.Q,B4
PQ>>1&.D8.B/\1'O='^'_[@BD8%]PV9H]KF(#67QLX=L'99\W@D7 [-I0X<)MX2=A
PL+7_O6YMMQ)]RU6P_MTPJ!]CS]_+1AN<'N/59I5N6<;!%19K=5-9"[RFR6^M2J+T
PL@,$Z::DSU A30GM:U(<#+H2A:V\=/PY/N8X],^9B>2!*B[Z$L[;V^C'E0%:<DS9
PG7]/$L#UUOAJ3Q2SO>(:?;>EJ8CM-8./:0JE?/U<U]^J8[F#"+V(NQ6BO3:*N#/L
PV:U2;Y-I_U0;?!4KR\>Z'R;EZ:?^2IUAMX!:MD;3-9@6-!=]S FLFB1IVA*-RC+L
PJ()8LB8'"E+FW .VEOAFUFR'$L:5T&$,2%IF? /]%ZJ,Y"WF&,XE5#,;9=-J\R9M
PAON.1[LXQ%2+MK?+C-ZM,<5;S'5%G15B2.5++O&'U9EJJ<W[>\X4E<.6M/]6Z8> 
P?'<($'A:1XB] /WVL#?/(:TZ>Y )L;]!MV*]N_NMF/!MF_7@HVZ<"2H [GJ2.7*C
P*]@;(FHR#,,MF*C^_3U#]Z+&];,S ]K/>F>Y.W,+P,L )ZAQ )-BKZ8$":^^E3%F
PZ>,)XYIYJ"Q>688V"67UYGU$^X7,.9)P=+/,!M[8M"C"-?><M4/,G6RA$Z<&5:HZ
P4CSB2GJ7&Z6[F:4HXP'&]X%+CZA0,R4B>V=LWL]CJ@W76DDE1[_I)9D$$O6X[)^[
P,ZM-Z[C!903;)/_#5)*@/$;(<&ZJ'\8'#5OX>)\]U"N%&\5]:8+(KW):/,\SBD$B
PI]/8F+%SB;-[NVN XA'O]4WIJ2-D'"1;Z]8=ZLM,>^R=1=>-$#;#[E;7AI#ZU75O
P4K=>'7'W9,P/#@.NC" [\+_>^>75=4CW]Z\W+264S#D#.8VU6:?Q_L,P%17_6C9#
P>!Q<3IV$KB6N^T@0R6K<WGT\A<U9;(JS4*9 M<2RXC:Z$B8P-HBJ"4-;BP?^:::I
P15__;C:0C0M3*7*%1A34\EQ=9L@XH:P]2RI0I4[[!=YE EL8BD\TZRY^I4I'$6GP
PU_G^G/?41RU%(:WH+-A2>B>"P%"58ADJ,GK*)NHOH:,\H9PZ\^%)WI&@8,9$_+L5
P:?_6XLO3]&U>% @!H;TK"#8.=]#5"BL-?31'.RAE4M1F7H?BKD#RG\Y E4BPY0)%
PJ5PC;3T"MJ*#$3A?NW7=0O\R:;V_AP&-IK*^[E)57F]FRO5[L,G@(Y]__Y"9D*&2
P'ID+;OUA\Q:=9"R">.$99IHSV\I0KODEPJ.]P/C+LUC"FKD$ST<UD,>_2MW+*&['
PW+'>9ZJ4 +\M0?<N1E;H[<[*Z6@H.131,Z>4VXV6J+?W(&(.[7^4[\*UQA1<M2Z*
PO*,V.B2$J)"TJICI9OFM(IG MN+&#CO^?:DF(^E1FJ?A4KKNC0/(/_Z90PTAYW*E
P$1O!922OF"!4*[(>2 [2U)$"+&O!,!D5XZ&ESLI6S""\-)M^V8<LL)[(I+OSI^]4
PDB4Q?-@YY5P(6%'B*D4[H[.W=@VF:FI4:+MMGP-$IZ859DB6GB=KAQ_*3!!#"KM6
P]3Y]_/[^A%7[6!QI@?^Y_%ZC_2#-7@EBU/.#I=&>L*^)?;-C+H/'SBUMGF4H[:,,
P_@UW75-35!U!<KKOAH17OKI+91(512H*D_2.IV<S*TH"!A"6#V:L<D![2(RTGN<S
P-WI9G%-=?:4U)H-<G*!6@, )8@)] 820D!&D##DVWO 9 )J9AJBX)]M/J"SAZLEY
P&]#*NM/L+6(BGI\0":QT#,QYR(:;5=$BH8O3IQH6[E"=&DOZ?,.-M0..."IIBR2=
P#G)WF:UT-3_[_ENF90NG<J6&^&>;'%R3*X[:LFT 4ZK"!\5T]AMT8^CL4L&&'5XZ
P3.%M1DJ-E1FW60%4^9^++5*V>F_TG)W&CJEU Y_<++V6PR[W96*ON0!-O!CW>3Z"
P"(^G;5L;P ?<I2UF/F=12_BK'X11#[MB=>RI1+)[F\+H9P90E2V4A=2>-)'Q"?V(
PN;](6LBE,Q=6YJU5U%&;F$$E.4S3KCT?OBV]WQ:UT#'KM;)3H/:LLR&'%F U169D
P7I;!/[6]B8X1*YS,4DO"_U*WK#\,7(NY3+40'/8?&?Z@G! \0OA+$=M8WACA:+U,
P]K1KQJ'V(4!Y/0=T@[VA+#1>NP1:&4B0]M(G>>CUEJK:W%O6W"V8F4>G-#<XZ<(&
P4A?FP]*C&GOF#ALV2.PR/:1W4=9CA]N [U>L%GR-']__OA@!T%-D#I9P@4R1)#\ 
PJA5O((4^^T13?$P14T"1+%FCW)5\]2]LN&K&Q]#?RVZI?^;K(N^ DBJ)X'R;#+V8
P^3%D8.+D\3@3<':TR9P/2E-3O,2+3'N/3-34+U<(]:YP=73KY95!!CNOD$BN476,
PE<?\<&P'%I5KH(MA7ANMM,*0TA]]XB7DKW=SB2!^AQ.&"^GBYR1]VUZA)$#%!.$I
PUM'G>+*]5?P%\D_H>NF7Y\5$#[UJ]%C;X>Y53@K68:#MLTUB_FG];VXC=/%HY^*+
PG.>CJB1IW6"DTO=H)DX\%?!1Y$QJ^) 7&!S\M)>-I.\HBP9LFU5%("Y+Y-+-R'4T
P;+T+LJT(>6$<G8-QW &CO*=':QT#EI$[87764GGS!)S0:6T1JRC-3/4R['LILYQ9
P#P]N$+Y_;7Q3CJ@Q[]P$*W#.L/K\MHN3DOOQ[PF R+H)%L5\(5Q<E$2>+*@\&)>;
P482L_AKZ3(/AGPD?BWG;>F02DB<;2@A=4WTO39<?0GF6N%IPQ9C*DO>KA;]3]G#2
P"WY_]%E'F%IVF[<Q1&X<7,C1W+N90MZ-7HGA(GG0>IPII4-\3D'!'69=Y[Q/==/Q
PA-9K<ZA+()J'?5[*6NQ"4%+3+6A[42%A^9CIL'$8] 7IBINNV9@ZL*]=B13[.&!6
POP!$<_JJ##Q"7>)P5LE88I13>RK06+I6G9%@)&<@CE[%:1@<+2*X0:&&%OO\< :;
P1DN6S$,36H_S5[.DO%<US^A9&75V#AIUR&>2L35"0%;=TBU+] _34]:O [E_WG:U
P\F*=#"'0(Y [_37Q6?@R<A+.YV_H9J<9PQ8<!M-16!,.VQWJ_<:%A5+_AAY)MV E
P0LUT>0/:M24\ ,JJ5#TQP6X\ F]ENZE7=[U202M0;! Q_9-!*P;1Z&C<J$<UIY9Q
P9;NF=$7#\G&S?"*T/A)I5PUR\,R$$MQU[Z%T(ZI(3QEOK5^10Q+!M35$U-V"%] K
P-0R7@EHJM]I0J%&]GEBH7+G%+.+/,F,/GIINN8S2/GKWWB:IK"@*O*A=:M(LFNI$
P"2W;^/#$O1_H:VK1(Q?0$IX#5&[U$\R1MX=-LULMUH%?X@UE&^0LF?A+G&@U*Q@6
PY(F(B3R<U^3,CXL]*D7VJ/+N-'28(X#>R FEW##H2]$]N2^<H,)D(OT,R;*K6<:,
P+I2Z/ U&T#1JY67^L'=QHBVE)B/I/1*TS=[S&*I=B19M*A4\?<;"B3P7EB$[80MA
P?;&YV%70Y7)#2C 5IN8@F)E6)HF0W>8B=_D+>38O?KHEZ6CW>.Q[24$/8!B.;.9B
P*F31['FY7@]4OVR?KB0_1-$L+'KQ9N!N61#/#SS1((V;4EL6,O7.0^=6(+E9%O;_
P$^2H<S&!5I= KG  ]C8NC4Y1PI)G%_5P 185$0OK\,W$:Q/ RMO MJ?=DTX)"O+K
PHA.A'OJ\;E].9AKF_'$!8#[%V(F) (>P]'H@/3)]\Q9BDIS?^0.C7X,(K BW+MIL
PA.#HVH HI(QC4:^O$"E(LGC1<2=A9!>I(IU_ RY8@V/H8U4&ORZ<>3NQ_3JAB87$
PMO>C\AT<'D\")F[$3&8%XRC<F4M'6R0+(GXZR2,3,$>'$X?\:^KFK!5_>!-T->2M
PQ.N81P"XVS!JDE)U#CS_=U"B</XIT=RGH+LE4VS7.YW(1*66GZ.$E8*?_(C4FH*1
P<+?#F4CW4[).09^>,_4#M;MPW-*OP6JP0WX1VOH&A\#=F0#2FP:(UD#Y2^ABJN$4
P]>H8%1JLV(8F1T7%WR$7QX$)\J>4G</.*F>NPI1$PZZ7Z6=].  =55B\774LC#G_
P!=<JNT&B<%D?<UQ8,W&.'$"#1E/7IC%B62.J-D!5]3H&F6G3S*Q$=  H;$8!>?!+
PC\,M\4 NRSCUP4H2OID_8^KR@VQWE[T )4:W/D;?!5'%')%O>*I'"?@ZG[/4,6RV
PLK"W,OTD35PE:#9LNN_/T_B#)NJ2^G4A'CL/W[-CAB&6GPB@@Q^',M@R^R'I%V\W
P;)K_AM"86C.8[%-DA[89!I,NB?3-6D(E!KB5'O(KD(OK]!$EW-,SHZA*E#-O2W_Y
PG(ED/38NE?XUI#8-8Y)6C;-66AY6QCC)3-MA]C\-(HQ^B0#4^X%C73^^ N9VW4<%
P?B1=N?YF1N\_!SDEV718@ZDRB 2:6L;[W*$4,'=SZR#R4$C=Z8XR?Z9G#\(0&.,U
P944G]T4FFM,64\J)D)FR\-ZJBX$4P'OD0(3M63OXD?)[[NL/=^\:=![Y2M.C([$I
P:DZJ(8LWMML:I3_+!<B[NC]*[WXP8D#P*GX*2M^)^-').E/GN&QW/GR1N3 :BG\V
P#RT0YCB=J(Q\RYC7\MZTU96N$XP/P+=O8[EW.EC+J#"<-G-(W"",:/?EIM998I76
PX8O&@![J>!&#]%.C4591*KZRX06Y)S5;3HR!6D 2\ Z07^%FA]V 5"C+CC Z^5('
PD>'_M#>ET4]/M<FVS+:FKHH'5_0VTS+FD>^"G#M*NC5"N_>D+9#QYX/HZZPYKXR_
PD/-$^7[LN>E//Y'MGF4B/4L_NMVT<WP"#+?7$B6_XO@_6TA3+T#G^UI#W=$?:'D+
P[AQO:$(6,0Q?SP"_J5;1C_SW\GDT+VOZT5LU@+C';C==-3?:G,CR&O_$B/$<V,0 
PY&P1P P%4/*P__\R71>@62JDT6%Q<6&;=JR<EP,5?;?,)V4&X^0B-./^$&$,=_Q0
PV83QLIDK7T$#D5$&B'"G-U]=HX3%VJ;U^+I+WWBPK@)W[0G98%N,6-/XO7#>JQO;
PE@1KG8#A3R$63^/WQM/4R#H!TN!MP;67/P&BQFV&D)3N)E>3A5AXB?&G]=&]9^1!
P%ULY2K,0*IY3VHKY.UCC3!!NJSGIF^[Z 9Z%!P- 4?(1CCOE_5_L=QIH*PTS?>%_
PEY ?#%%XO;6[ZO(83S[I%803FC"F?:05L/)5DBIU)4WU;G/#]G!L< W,%R]X@C:K
P&:Y/^5X>A.;#HKV7UUJ,(-NB8$11/W-U&Y.T:(D'N->;27_!HW2&^M,Y1HUT\S6(
PCD0V>74"%QYE._+B.WB[(X3[S+&W<FB:U;:&NO_FS_;JO "]\..#>^6W&V6?B<?R
P;&DC LEJI[P*M__M\P&0"$D<PD2$&"#>P/)&Z96TH<2SI 6-WCPYS QB0GF.R1??
P[3,_Z5,^&8T /N[(_XXOIM"0:[EN8NL1#XE>)=U'4$*6WL-O=K TO]KX@C?MTBMV
P<!^AL>INL#R^@&IXDJ  UU SJQK8X6UGQY-A3QU&/4DL!1G3O8 ]3O5J:\[T^I"O
P/,RZ1,W4JLQZHZ[=5WX%@@\YO%KJJK0WW;B%Z=WPY@9?5I,9?5/B949<H5V+>O[F
P]@F->4M^.:B[(2M6O&D@U9^;9./AR*9UG5/CDUC3=<-3^V@+!;VHQN#3S[PLI40]
PPIV5^(%-0,1<J[FTR&+ :HY=V&]R\B4!RM,"A?$,@@0)" IJN)J)=0S$#Q TDIG9
PO"X?Z[6H!;/@3!Y)"!5DCG07/*=(W&7M_=O9% Y0[J1WJJY*Z"7VO_DWYJP9F7)T
PNB7UX&3-%^NQ&I3N=^)K.>UF4RK81<Z(\]O:*#9U.HJ^-[XM+=[W%$WKJ?)FF _/
P=U!/BQL*,;]ZT<F\2/\/ J#01&.6K+NPT.$$W-O6"K?IQA%&K&,NIRCB3F1;9L^>
P[8U,5N8V+&F3 7\YWC#99FF3E?A!"?X-:R 7*RF0[1D>+>;#/\L;/.5/WK'-.WHJ
P(D0E6H"!SUIVA+MI("3\]L19.DOVS=[S*.7 >%EZ"Q0)>3Z9[A, 2N2T^)8LD9-A
PB /+FXX[57G[0M&R)?[#) 6W4.5C,YAP!@J/WU'!>J4-9IHTL5]H\^_.C]-E9&@I
PN2O"L(N2/A\YU79%68A4D&S]7-*^!K:I4V&)!D3$[:=^*.*&T]8\X*]?7/ZQPUS>
PFFV9(:9^2Y"/.#ET=>)F9_^S->KLKM%.-0^T.6Y8/,D3VE;"@RB_7:P@-+C 4!(%
PQH I=2^XO57$[LTN\_2X&=#H$3\((EW.JWS0:(I<4*9%"F'0+GR-UWR@:[)PZ]VZ
P@B6Z4490*&!./4.L*G:ISJA]+W?"<0:CNW2E-V-YLFW$/,?'BL-5W#*<XM[W&!.H
PZP=S5_2Z:8AMU"E4*,Y=/YA.<'IQV?5/:].;@X]WE\.XT/MRUA,V08"6U#EG0KFG
PD<C,# =QZ7NE])@\8-DRE=D DIYS3$H"<!0;$%]=788F\8E""]?GK?Y= [/7IP3Y
P?DG>W;) 2!6X*_<7L1L3D ZX-<&%L?" $Q[FD$9EU<U6JQ,]&P2V.^_DOCY#+3[[
P.?!XN*N8L>P@SI518-T./.\4DDLC<1T:1!'5,RT2)@CG)RW/4P%6$)N=T(\*%]XE
P\1\&K&P54?'* D):@:N]%7.3)?$I&,E,N$I^VA*R)^0'3A?])#_[G6MJ(BL4"Q^Z
PFJ/]&:M=XG):8^GW4 \,UN47$88U;R^"GQH&ZK^E9PJEJ8', )S$B*P^&D]*'07)
P4351[GP?9/#;S35MY>WQ02@E("Y:='^]]=4/&^#7J;]9:-6 $5F_-(]*;=^PX0C+
P\@\6F=V1]^QS6+=L+58W[H-*77#E:R%,4 C-BCN*GFEA!PF\ 8=5@S_+';9,/<4*
P#=:H -Y&$)RJ-\;D_.UJ9ME@D.5)3[TW@@BYKKTS*"<^ -_P<=&'.$2'0'=&!K& 
PFZ;2G4XM5._!)'6INL!$L]E#BLZ?(3FO1[I2":JU*I:I&9HHC^H!VG/U2L75$P/L
P6K(":I/GS%)?KBNIP@5TMY<-D2[FQ-SI,RG<\W*1 3T).T>QN I\M(K$RHNLBP?=
PUF,W5+$5Q%W!-XJ2<Z,=QP0?%*@9T"U3E63Q+^7=7J-1H4^'K **(D48Q7T35.=(
P1Y^7X\J4'Q,UAMY9<>=NQBP=F@8T]E#!I:&BMMJ.%"+7*O4!CQN%1>KII<]:K_\/
PWS0[=H=*WUOD[Q.HKR8MLU<@N1@Q+NUBE6&>F(U KPRB<#^'A_9[3@"KURU.A2NK
PC;>:;K28! Y#7<8ZCKXN)**C1+OSHF*(J ^C]'%HQ3_.&?ZYY"D41VKE4*$D/_#3
P\;(Y *-Z1-@C(1B)E*,G:MVY7V68$K='2SC7.6Z!%*UWH@V;$:9_DT:.-%M<)%^-
PLFWH8=&EKMQ;B+KW,,#-9GG* ;FBG56;4;]O@,&Q76B VZ1:&"&;;H*+*QAL0715
P=_6\-*X_,#<J$@_IAJX[51JKDZU>P+! 5=-CYR9B%3T?N0 +V(D@[/^E=6TH.:0^
P]*+PI1^Q!^*W6#T7Q:'<Z0ER#GPW6;8K"N%5[LM:X9:"M;>Z-ZQUR,2'+B@(I?RR
P)QUHFAG5)N-KI\^9Z4,8#.&&)HP6<V@9E;-6/JJ0=&%$>ED7_1B-M"ZDB59EMG-&
P0Z!:N15&HXA0EM?,I#63-K2C8A.+)!":SF"!%5/,G_!?RV[#+UW3Z)L/?@&7L#!7
PEB59>D";BX1#HFJG8H2:@.EM')UQ9Y'?7?5< \2R6T@8]]CA:_9&-OW2^I,TY.!(
P+?\7?:.>3PZUG!D,Z.V"R_IC<'7FA:\2.: -( .<>PRMGU9['75O/L:RVX#=4(AN
PG),+O=QR5TO0L&Z;I3S_TO#/2AT5-++KDI("<!)6U$?>BEQ 9]3?I[/W+ [YSBG%
P'SW(!^Z^6V%_MEN#- T=W44+^N >023D15N&*ZH+I#.-@\N.[;CLCFR.#^G9:)/*
PSFO^&HZB_0!8XJX:TME5U_$+#M AMI\]8\)!X>8Y!QH_C:R#IARW)J_XO%$HBLZ9
PSCN^N7"AH.N$*+B)V'M4 O;+/'(8@VV3,6UF.C].!]/"R81FS8[VI[=X+2UK9D,%
P>+X77^4]"P&]CIRWG:[0C\L24*#^I7$5,P&(D>A7'$SYK8!JS:(EOFYY/<82<_I=
P?_=RWAT5F-8JQ[CNV46/SBFY8.T:O7UV.7K&!1Z&ON_,@&-SKG#)C9% 5>W?;GXL
PL$)#NJ<NI_<*+.M,X[^> XW'6)_S%_;X9=2AR%@<F'3V^=: R.TF.I&6D4#OU.!-
P4MWD=#DLY.QVOOA%L]+9,2VSE IL82*=O-^6S)A8G^O1IPZ>FH#0XDEU/_"Q#,]J
P@Q3N42YU:"W7BA?&W8M-X=LS''U$V :3HT&'Z;AYZ'%]93,5W9.S-$BXKU65'T_^
PHKLTM/Q6DTM)..VU(.U0^'9/3&CWZ6'RMQMF.2#$Z%1E4VZJ5V4-ALK>IK<(Z0C"
P%%@8*KPO6J>I*B.3&XZ$: <)_FE@XGJRPD,C&TSEZL1G3;TK.VDE@'K?X)ZY U7<
PO%J^U?]TIT@>VS7&X-'P?',C]C>GW?W':-;5-6$3\<M5U""_U?.)^8GB/]?(>^4@
PQ2IL?#*)W$^0D1I7%^ZJ5'9S(_)XU_SEES,"BXTE[3_CZBHJB\M_]+__Y%\JUILT
P4&4"SN>-) ;E'8(+XJ3A;<OS[->UE>>ZIF$>\EFV)=]^J<!T&.!2/)<#E*WRQN&1
PAD\(>UAV5,1\UDDRS"$H49!3#>V&\THTY8E+/_8].$T@9+,9HJ8526_-@.O#4Q(B
PF!.D )[K[6,1V(R#* 'ON28I,PXSX"LR%T;*P]+%'R'Q96Y]$^5DXR3,$ZQ):Y94
P"'S^6F[F\6=779'&_GKZ'+P<1\9,U%A%V01X.4M9-"N;W.4]I,>1J S?WN7_6OI'
P#7!E5?4>)!3T2CI.GFSTZW3)4J8MW%Y&0B-P$6[-%>?!+. S/SE9]_6JB0,3]/A)
PM(#<)#.K:A<1C.R8NST+7RUWYI$Y"-\"VGP^X^<*@$^6UO?'O\O#33!]CXTP#A5.
P'(;<5ZP@D/7LX')E1BQ41>QVH2*V1@V*>&P\[=7FKM//YSNU[X"T"1(]_ NTJV*G
P9R+IQ7WP#,-OH>$T3,6T4ZD6QFLT6FX$,"3Y[>_<60_CXX]\B>5/)]EKT(.#FOKM
PU6TBNG);_Q F,/.]F8>0^T2?-=R^ B6DE5_$@2"66HDY1N%.L&"L/B6@?8-@5(GG
P%:&J^Y)?B/8\ [?VLH9GVB;[4C@5G66>A=YY6%^-D.Z*84FZ\/,Y4]77]H [/2H*
P"I8>,B*$-@I8M@'NO=)V*V)[OS9!;3>"CT%WQ@R(?[,^_)X9;?75^$;)X@F7B!YP
P<*,Y^QVXD+[+@3=S1"W$W-&20I0G$YHCXF.!7=1&_?:SO>,7&$52W\M+8S7U@U,'
P1JAHVML1"F=S:T1-3D).P23ECZK*S-T.R.L>S=CT,#/V=9/HW<*4&[ \#*AGP-Y9
PI#IH&0T+\_:DH;QTV$P/1D/X=]6(,_2',3;4+)LDDF*<%^] @J!0S]+LBA+.\BS>
PQA,A$>30QZ4F,G@ >4]C'#Z5AC@TIKVI][[1!UEM%H/3L<]C9DB8H&_&3!TZ[1#H
PH@3 F_J<'8 AR:3 KAW'$<M#ZX1@#ZUOSF0;?<2#[MEX-,0Q=I/+*:PF,TC*;XC-
P9"^DC=":G_UU6*=8XI'V)G4IU>&R,8IOB6 ^H&MU]AD5[>/$/[J(\:H ?@^84-GJ
PYD4]'GY5,(\M(W*<"./,,<I:/"8O\8./ *9&*Q)9R<GM_,[N4O@00C5!!C$[?&D_
P]&EYD'&2AWTWU(0/YJ@[$C@DI&.*BWM6.@? R7ULR?VB5;ODUT9\G5$(-8:I.&ES
PTA>/(B%]9Y>ZXO6],9'*08"%:.?CQ9O[1"WGS)+4"8;U(KF==Z^K,3R+/_RO;QW0
P8ALX6V!)-$X7R&3=6D,LB<+.@<J+7585S>._J[%*^%?XOH==MDTJGW)PD\=!3Y1%
P4,XE&C=)S>E6!J%SFA<6\/%5QC09EP_5>;QMVJJ5X3C,_V29?\$.54O(WPJB@B"5
PG]9]D+;=$;9U0N<'5W[A*RY,A?Q'F\7R\9)=+$EK?]0N_/ABG?9[ G3BE5W[-AJ<
PI,\J+1MR,9KQ,V.J+'8J"#C_,J>BO\:FAEI-1M\5\5+@=V1:UEJ,<HS7NP7;+F<P
P7T"R($;D)M;".0=)-;2LVR^H6MO@=5^2RIEP.GH+C(NL6KVC467!+9#GH52%+SH[
PI?>_)$V;0M@1_D$N*ZH#5RRGL&MX(#@AG@!_.V2!Z]!'RII:_-] $K=O.](B(EQ7
PAH)/RY/@XI_9?L?VW.K>I-AA)YXK0C'<LG8V+YBPT'J3]6NW>-39)^CA"9W2C\/$
PD1GCET%9>>+;R_-_]_<, 1_5CB@ "@E/2GO93:HYBTT3<.+U+;Y1F?RMJ>#ZB!LD
PWTMWYD*"(*]X76KB#TM]+SDF;T.C;..E/*1R6(+[YF6:G!P0;\HQ] )8%2N,\EG"
P.BQ6.IOCF-&ZWJJJZ^5?]!J/N=ID5G-(CC3QYGESIOM%_I[*A0,)^;/BZ'5IE!R!
PSDI#2A;T&-%$,/O!/9=O&T(L.9J_)X(!PCL&+-\YC5J@5E-2J<?I*%0G?0I&CHZ/
P'&%JNSLH;0#1(I0F=9(F^S27M6263MZ-Z5FD3%2COK;AK7,HX)]>Y&O4M"![Y%8R
P72:)[XZ/%%;JW]6-5W[/45>WJ[^8>_W#AXG38J7]7%BE4T?@E+>/^?_M= _#Q7IZ
P?Y\$UIWKW\J7"*G"U1217HK.5@0 :JQA30I:V.5?#XF9E'^B38:92TVOY\T[7<'&
P3(?E^M]J@A3W!!'H3?%*4;53! @U#&3[<=EUB%4")ZT 8LT#6.%\/_Q=X&:(8@S)
PU(AK&_< 1OU5#]3$T0+96):0^M^^5SGLH=2Q)/U>DXS$S*$S=4\*ON&5Y_*ZDD"F
P#'8YX,[!@5VO'[O?'!/[[,5=NVOY>^'?JRN\(>A^S+71FE-17]5@UM>S.G3$C$'Q
P*-76"[QKJG]RZ'5A$'JY^[QW\/ 6"5[C-9Q7_N[+"*W.I8L!&/MU%4G/%@,_U#T_
P#4$K(7A]R U!(;Z R9(Z./^H_R?=UR+>Y)_J6+S%,F]A50-8A@B1N^M1S=^*A!P;
P]8Y;D51^9W8X@6+#^=3<IS"HUHB.Z$U3/RL8_$,+!YHIW?.Q=P#SV^M&H:EN9-<_
P>C(7B"=<_I!?RE/K%9 A@21&O03[A-[\JQSO+0$CULM37X]H N5@U]@ME0^@$0VY
PW^C%]1/POM2I;%;WCT2Y"B4Q^CJZ+M!9HF:E<X*?H65^$G@IC'9"+FHDLBV;=^Z5
PO@UG@3G86:]39#7V&8E[.QN;N/ZR3T5RH$L_6%Y(VTF8/QWS6T/,V=V> "\A\5.W
P1J)@DG:EN3TH+Z<W"J=\IVBQQ>A:2>6_6-()3HR50S[5I^Y#BRG.H<9,0>%>1E>C
P$/9O-,#SCF"I&0.0L,+A 4(;5S&SVL:B7@^&YM6G>AZ K M8,W[L\.A\Y;-7?,9 
PJCI#XW7T_XRQ\*.K4@GE&95JU>!F3&CQMT/J,R,*VA]JUJ* O>7$>D61*2_Y$>':
P1M&3HL[%M\4IR;QN6VO=&.SCAU+O'0/I$B/&A*V@PT)RYI#?7D[.D3';TBR0N$W"
P0+&[V*B?LG2^6W#OY&:62:F%8B/V_YZ@_KC^N,(*Q/DG&:1'7,NTP>A!</]F4!8K
PC@%GSC=10Q0\Y4DS_!V^-A\:3!?OM1=,W+O9">[UA"^GJL:QF$R'7,$!:?837$> 
PD&)X)#6PQ:"C.SPPP+XZYD3R@KG"&3B/5DT^E8JLY38DRE]BV<$?7_N&PXA"^P6_
PU&N4(7"=KR)_:_8@K^LA+"]AV0W&Z'ULY-N:Q^XQ(;C]\-/(0*MK&-IMT?#2H3S(
PTC;!#U(!#-AIWN#F@58>#W;&9)8KZ_\!/_*KE<D%[KF?3AN7EITN,*9,PL]UYWS:
P#P/*.G$G3CUN7E""R<YYQI/4P?&#;:&P1]Y&Z_\9;?X"9&E7I*7T<IB+4X^L]>\_
PN]L807<B]8:8'KJGQ9]M38#P#]5J.@ M'F=2/M0<[K/JD(1H0E!/VK2X!#R9583F
P"$"/X @MH>CAW?U;ML<V/<VZ[-4F CZ(7,#G3;MA_G C@S! !FNG\7B9MH2SV"S3
P-O@ZR4+6M746[6'WN;%9N?Z=D]ZYMAB>CJTKH5NXHO:J+N'(YB]1_#.9:^FXG!7!
PT3'U+W^N8VJ5B5[F=R:CW;IW^0#!XMX>DB!>,CE2BAX77YP./$+5 C+P*U)?8)YL
PJS&13Y1#C4/XA_'&1LO?M'XRE5H*C3.;Q83+,%Z!H^C*.L:#:;/+#[R),+FV'INT
P]BHPCH_)=#8;G,!0EO )U'%[[8'B8A6B%#Z10[0E8[B;6+4]_<LE__N$\ID%^\6Y
P\4:)(']40G;2^UN,\!83',]ZQ!=98K&L?538RKEP">JQW-"!VEC#S+(FJ33KW)@#
PQVZ/\;G?TN6ZMGOSF0E=CFH0B)E'T[EYI^% W4<,)X*;X2\;HO?@W.;GY?&)7079
P^[F9Y9<X7*P# %0[NN/G %7O$3=E;6F:_  OPW3T+FG7.DP0:I@!"I34E;.XX::0
P.R4;*B;&']Z^E19K1?H]F@YVD+*+@;#Q?DYVCH)>;;[Z+*%-TH;ZL$:E-B#TH!Q*
P,KIO'>;F"7=KF-?NJ_=4U<[K^+BJ6M:O L 0*B$\R5#7'LJB(@K%L3@97G9F!Q]$
P_/#E\@9'A7%U2/.ZCM0+K@4Z *?P)8P+I EO ,*9LYBY-A9/N;LYM?2YHD EM$ .
P*RZ^B$G1[Y1\R\:84<9C+-#73C ,(*H0'\F)76'5,HZ@-AF8EU^$CZ>;BU)2-C*W
PT[YZ(H<:X=07_O$.(FHMK/0U+.8;&9X0T :4E<^9B\:+TQ;>M<4O255EKUX.S(>,
PGW;X3I_PTD10ST\07,E=YBS\.(+-7(7CX4 *EQ(F<)AI12)IBRZG^Z(;3^Q<\R;G
P+\X-I9/MA)Q/&8X_[ZZJPKO0'HQJ3<:4!OXM$V[\L"G, XU:MN&OG;0I]!ND;"<5
P$Y7NT O5Q-WW8S"*!_$[D(O;17;,\@@!R+;.X$)2Z]"]CUAY:$+:29\J+.E1C3(3
P!&8ZRK]<2"6<H^7J\770/$.IB;R9X]F[3L9^)><(O\3REP<UC>KJIPXCY-%OC1G[
PBE0&*H0N.Z.6!&F[&_$-WQFV%C&(-W\2K+NHN<I:?W C"VH4E<I.;^!WHY?8]3_:
PMCF !C![C9"@?B4Q3VR<V+K221XKK#PEOVPV@9ZN]@7'\)*<X#)(O%;=C _>Y8,'
PV,O0('?QEE2<*]5?Y\1K0720(=!<*7500/_]15+-D8WR1.)\/JB:$1EUH8]_(>D\
P@B,>SHTU'(O14/P/,L+$&\W=GJ%OGW:D>&^(^;V?8.8?[1F%)5^7<3L-A99(^5@:
P/MCXDZ*2*$F"T*U$IF%2I!J4;I>F'/W>A;Z#X7+>9QFXU>#/3Z0> .7HDP7K]J/T
PPV %=L!_"XF5*SR&]G-1AGF*!YT%"\*[Z_2MTB%0=%?V_\?(T,QOO7IPYT)G R$I
PP[\7:DJXCHYS D>=X:"_V5QTB@R!]-VVQ@Q%7-[.]@ERI:O>.;0&R<&(L0'^%EDC
P$1EE#K^^:,(2 L0:Q)^2"/.)TCEOL[,$UDHO:</Z\/J"A#S5M<YD:*9=+$V#5_$4
P0-&.@EN38<PO=(N-?69-<I6KPLX&BFWU.4E^,18&?J0K&XNG\QTBIXXR__9DXTDF
P.C.T0^J$:?LLB7()>!^ DHM<23\@^"UJ3- _ZMCQ6>RYJ*<R4PQEM_U-G!B@'BOD
P@LR#O@.O#9 N:K.(F_-VRVYFN1#22HN2ZCMXRHG1<;WX^E-0>D(IEV=^)!H!-UBY
PX<WS@[!Q6>JIFRP2A"@O+&PD22PHO=]+*A'G+^FBL7S6MJ^R!L4K'@XD]N?8!?I0
P%QESL00$<@*WX[10=7,\37^&'8/)&S(B02K3?&%KQA(,=I/9S6)82)"'I<',.+[8
P6=+ )CFR6G[8,&(,SENEJ)ONZD%"1<MGU9D??A-5N:C0S"A.F\E9*QIV)7<R3P$W
P$SR0NLHX0-]X>Z\/A P!&30C@P^=-!V3@JN^/L*/VFY%T/D_KNZ$E-R6A0MWH?C9
PI;! 8D$ZK6;^X(O(] ZH$)[$Q9:Y8[ZCEY;1T6V5%<T59(F-?5-TA!0'V_F<A9D(
P-CM<"A"TD&'QM@^*7X*9VY@LF#L. R!->Q*F0VAG4"J#=-A_(./8SWU>YX4]/:TE
PIWV-ED&@8 <R6=MY1&LK8B[\O3,^J57Y/]5A&PB9ZCJ0F[#C%W!"TD6-C_\E72P$
P4!\(QA+ZY$YJH,'YM,N01%73+:]D[ .+=6_U' @] D=W,Y>@0@7E:O-S&@,GPMI*
PM4L)V]#H.,(N>U:G/E.["WSY&NR+?BXN'&E0KE#DV(9!Y852/5K9B=W2>>3@A3?8
P(T6CZSG[RO2]ZY CM^V3%4=P =NLL/,SZ2 XP1/@Z[IZH)1_HM$QAK&4T-=.XEIT
PXR%LR\Q?I7"A=;F)[U521L9_+N^B%:<@L7A=VR4#O?SGK%/,O2F.LZ]WFTEZD"6@
P\D&R\!M0&+H3)_E4?NE&?TW*F.W2?[11[B7O CS2TXS]CESM+^=U_O^V$?*.?0.6
PYH#?EL4#^41GR![ED5M:85:XV%(I?3"M[\-"SP%]L*3?:9  5GB58#)V^GFJTGHX
P;,9O*KRG[ #R+ XYN>T7<0=M"$L:ISDE!E>3&ARHT>L-^#_:>FL%^F24@E]YFR$K
P<V2BGQ00%F9J5)J)3C=N[XN"C?H95W!@3]=^W/9LO4?*:P!J"@5!YX>88>E= +<<
P*YEKV\SN HXN844S#-V(#,LSW?VV'Y'U6+^646F+^EM:L7_!&@^-QY::Q:[.#D*X
P3LXZ,"?Q%< [83=2]J ?'E-<5F;C8.0"0OZ.=)^)]ZB$4)^D55S)E*JUX.H[3K<,
P>,!=72C?-0C]& $L3EM=AN%EK,5%UB;CD,19K-J%O)7'GE,,.S=\L*^@,7-=V1*;
PHQK^G83T;FX7 ]:]W0<IQ*L2_<PO\CMWOMC EN%4-]P=Z,\P6/'N=Z.#J@20&HYY
PCH:9]:)/XTLB#+<THZD"AJ8\2,]$T-,S+D])Z(/HB$%8%*)AK ;:PF.Q-<JG<VA5
P!4[SY(N4=H]5W]4&L$0\=YCNO'*IB%@N DQQ&&#7^#K@CTQ./0P?EFF*8V< >T/"
PY7' -G9:3Q])W#]X$)0\$[3K^(S6R3)[3?$, I4[^^VN);_K@QJ;]WYAT03J,5J[
PS%(UA+*L)&P[B5VDBT=F-NJ&3V[IQ!3^ W4%-+M*#:/7[UY;$ N+5L> ^ =BT!UP
P<YF4A,V)%+"$I+H1 MJ=I&A;&E,-.=?,!Y*[@T82P\4,!+-XWU+)39//#M5C,FG$
P[55=ERB$#'OUO-0AB[9B,DG?+Z@D+D>38>CR,=ZF"0;0F?8)6&"VHZ*"XC@&>89O
P+7 ^]<Z:W7A@L%$T?#)_W)'&70'/38Q6H\B2M7^/DKNP[NP!">A<63;)K1 /MG/3
PC'_Q?R^#2KMN2\3AYGZ[<.#0@ C7F[6- ;JJ?O0^CEGP;>L@*>26DMZ*61F4Q4B5
PF_H2G<2O-WK[X0-@1R")8'YXGL\[97=G!TSC1!QA[I4O NDP@NTPPV?A\I\]*.<@
PD-H[A4@?H>P((Z84Q$':0;A/JWZ059&KF0R(I1 _Q&C@Y)&]<K1H6HUUUVI!N0>(
P&C-<281B%FRG6H%UP5]YLGBY4IO5W7[H--[Y..0-W"#CJW@:E!1PR1*(98727D*K
P.\$)N;0@C?-]VD)9632NT E*4W6XU.1%E?GM=;1-CT@9QE8OX&[,*((SYV=-W0<Q
PL]Q;%?NB2>Y1S6 1?A!IX]64$;[=;E[!L]*\P1=FKJLEI6F*P4WQJG<PM.=:O?Y#
PMAPE@LB5S+4A2!&ROPDP$1BAKD@!)OMP5#[H:PO1VI +77,$I8\BTC%227RMK[2*
P-$YY<.6-MPG@,8[)/U?/+ _EV-#VL(^O(D+QG"9)_A6/F&-2)$9()A("]V($^JU&
P^]S'64]Y6&C^V24!=JEK[X%F NA8XX;!AP*-K,^T794X V%8$.$^_&JJ4G$[(C9<
P2_E3UE#+7QPL"H' A&>F.LUL1QG9%I9T+$+I8?G]Y8UFS3A U67 GJ%/G[_N!IT)
P>\.[7J)J4A'9'00&_U\VL9>DG+CO< AN2T<6Y&KC]P?".]?,G+)+?SBT,D&'C/?P
PHQ#M*X/>AB'#8#$8LA6^GE40SX=,/"30S1L@G,S=.RT(^T->0EM4*D.+)U="Z!A$
P/U@6 2)W8>*T2'=F,=W3XK6$]FI"8PT9D>1&=@6EOBMF\9@.E7JQZ5[QYN P$N7K
P@&D=#MND>AG>SFZ\!*)VH"=DN YM&]B"8V&>2]LN&B3Z *'5%5,M5<R6?S8OKD;(
PY, $X? "$<QLN+A"<085I$W$*?83'5"FQV3 ),54,4NTDNW?1('."X.[P$@R6J:$
P-S0A!S&RL\ -,:?5THP++OP5L%#Z10C%Q4$!1GYV">0!R%O%MIL3Q3/T6_96WG+S
PFR5&8\OY$8GAB0(1 MIL>/O3+($449QA(KMJ[*3TJ1B-=]C77C=8LUU1HL6/M=H'
PN61J )-Q'O_HI=30:YT/%<XNY)1M;>R]0;XX8FE!6A5;[7S76O/WOI)%,T C\/7E
P6EQY=]9/T S\IQ[6:':L*_-@8'.+W#HDRDWP'XM<8\KKNF2W_DF7M+N0QEO9'AP\
PQW0<UBQ>\K/J>.6&N83[C/B[=.@<Y@"I78U(9?<6#X%6Z7!1$XKRGK>M--AJ?M$:
P)C/BM_KWA4U^T$27C+O3T H+!+C%GP[=OD!Z /#1958HMV@05VY"I/$;#NLYJ0R$
P;*1#P'_\E"'W7C<=)VY0>D?#[2%%2W0TIF[%0=?>4<[T/;C/)RH:[R8!NA6N95//
PT0*S.2N@"2?5B'BEL4.)X]\2(K:!B=CG_L,)Q2#^KS$Z !0$I54](".8$.87319X
PG!IC0Y.GJ>!"27KWZI5BU-N#I&OO;O%1Z2-D!VMDB(QMD\P85YEL3<OXX NIJ$&[
P">G)$]*S8AUQF>[^6+>5/NB%W:,T24UQPPJF\3I50OV%,C>%6X&GOZ4S!SXUL)-'
P]YP[LEO$>3)3SR?"/F:+.BMEW1>2NU^G"7Q_\:ST,492.7(9+?35'6RP>6GLQWT*
P)$QJ_W.G50Y.;=1W_O3IY +-4]U,2"9Z^(A&^/1&F\^0I78+GQ!1<#0,3*,S9!B-
P-PTYGT6JTUM'0N$8$T_37Y2LDL\[*CP03K=.ZZESTB8X<C<74D::HRIYB#OCG/<>
P_+VB-=56]K@;'7D'OE@+0 AD29ICS K]6.X02Y[#\ _P*[LDT*'XPUW(]>J:G&PH
PH/C%-/#SPI1FV'*RVB(E.WK<[8-P-Q1ZH:S+0ZJL*DXKO8O6F'#[[*R.@K,<$S74
POUNH'%\E,VGM=C1Q$"GK6\,./6%P*^HAA@Y01?#_FB^P\K;C'NA8>+R30NF@T.+6
P$2";@/<->]W"DS0F1'%4G$D>;2!/@);M<+%LBQF<BO8.>#60"6*2I.K8ZM(9^X"9
P8O/ !E%[%:2Z!(K.H\.M]X?]93.9"W&?>IGWR\JDH.W<9ZRY--U#QFP+NOP5&8#Y
PV,+V';/E*I2Y]D?SZIMY,21OA^K]%@%:Z 0>:L2B1F!*1\**2)9 S<0L*@Y,RQ"5
P&J]ML%^[5GT_HHE3[7HCZAWL'R9UE.:SLC\6#%.ZB!Z\N"(]M: QRC%02W$RHN1=
P_>U*+[LGR ;A>AJ0NX)T<$O)K"IB(_S_C/EL19/FZ=^")3L9UMNFG5< >.:5!6*U
P64H7=-TY/X[M=&6O&$."%HHT)9M):H &V6%YT**R3XV.4VC2-5;C7PR8R08&<.?0
P6IE:^C/AZ=++B?=9< Q<)?X\-[\O]1[<QI%!K;C6KHX&V)W-1R6^B0G#*+5* ;J(
P^F)J(8WF+<V M.4K<Q [!C7+>)H[1[K+UAS_ ]VSHP/ F8"?(/D_"M:5N3SPW\%C
POO'AW,;_&?H#_]!U='U6;*<9JW/%65!Z1XXYW,Z7DCV:B*MH92&+9*J5V2$2M.'@
PN#/:-BM,[[-"AQ#:/UZ32(XY$\V-^.9OA^Z*LLG T&@C=ET69N.S4;\BJK(!0XTK
P6*G&D'YWYO,8R/]CD^*-[^9OQZ)AWY["%YIM2%",.'<WU_J,H]'5=[%W=D\7WVGR
PM6W/8L78?,,D*??D2T'I![Y80!.R"BW7N=A9U;3I\*0<"L3TK;J%P$@+BDLZW46$
P.7K?_?OSJ_8D=M@'3#$.SAKK1]OS<KAA8#GT-%;%99+A>8#66_""Q;T^43@-D>N%
P9MO(NFKIO''2)ID^\ @#(N/$:_;W7,2'^LJUJC!3/'9F#CLM!9W(:0:L5\:2"R#7
PNB>+]RF)\[&J[U*WDE,@F<:'5J W]WH)Y!X"!Y+-45=Z(_[,EH0*R(W0E?E?KJ1!
P*5PNR-O)S+^TMB=%@-%93-K3CS*-_P'. $>*\;)NN.-BJ7=.<XIS\!G6NUU_,\@H
P)-5H0KBOZ9^-\[2+HG _I"); !B46QXJ7?;Y4V(&LD(](H['ET#I:M *AR@,5K.G
PD5%-$T@NTJF3%O#P WT*Z%^VT( =23K@X6=MK_D@JVL[+Q/2I 0\<333%QH[&RA]
PM^5<55/E;T7MAY WVN1G,-5KHEGL#E%7Q.,0)QB+P9R8$DS ,P%]R6=R^(8 JI@9
PD3 5I.VQ=O\?'GUE)MF9^3_+N7_^N).LAM]G^+%D&F54#U56\%2S8U9$PMY8\3GN
P]\G>#$N1@F@_^:;X*;HTVW'YA?TO(0S/+1!N0,63@Y KZY<M5>HA=P>OHJV=!NKK
PY/@3ZQ3;#0?18%569KKD[-E19<;^%H! 0TU8.BRA&""S'4]NO@I=$Z/^]'*GE>3+
PU"-+(HV;'+C#)@0_!7P1\G,EJE#^,R$/FZ/C.]O]]5%@#9(H?E62]P2VV!T9XH9:
PY@CC7QOQ3L?M:7-R(*"RAF(JJU,?Q<'R\%]OCQ%7+3OWCGP9VS:%/ET#3RIR:)!-
PY@PER., F_<@:_;F&,#T-\$N.#O/6\8(N<5?]TFSZ5B01WQ6;*%4[$$F1".HJ7- 
PM$UCWG3%ACB>-@*[(-8#8IVIOB%!+SCEV(5)7MULO8C.-"79]7:U\>S-S)V8>Z4K
P/KEI%NX2<+?%1C'*/"/E:JR4?X[@>SD6QQ/S-#))N[YMW&Y%#B':TPGLFY*_8H8*
PQ,3.U<+ZP:U)1TN\EY/>OE["CH\R@W(W="<B.>1=.EI_C.=&]<LWKIPU_>:7ZF:6
P;4R8[>M38BHC%:Y\\>,)L=;0_M18&&/W?ISK5&T+8MM_*Q2UNRIWGB91F9M"SLI*
PT\;0&<S.0,!8&&Z@X_TM VB8+.<>$IP'A_]H#V63?/#G'>H@B8G48_0YO$5L]:] 
P@TNA.0, ACBUB,]B.3*"9==$(,V;^,''$>!G_M6#!^GR7_B)-7F+95E>???MS##&
P$:-BT,:GF9F:D4#CEL&!G_0QBGDB64)1JWL/[=H/U =(\RW]I>#[MBFH]]EY.)OU
P[B[*G@=DLT$[@'ZK>M//!IQL;MK)AG5LF7CGFC[Y8YR!^/(#OY/O@\O\L&L;,RHW
P:QX"I^-O<!Z4@'_A@>O4='WD9T;Z2%(N2DT.#M>,=9=H?/P*]N@B#S)D"U7FCAO/
PCF&?%E_(WQ/<ZC8L]3-.O8@XIHJAMGDX=.?D  .("DCMF)3;F/>.%U!8R16APT[*
PEPBYMJ]04NBVI:J [%2+>)V1_.B:I^@H#HU[/$SNK[H(2"3%=]%OF7P8;F),])#*
PD#WM^>#0]Q4?XK92$?<S:FG\^SPX\TP%>9-QB(YV"_CLK*7:T6-MGB]U:5.8 98[
P%:R&\I[VE0!@N>![!WFTN"5@A@^5ACI6.$7#:_C3W:M%E'>>1% =L$6J![((OSRE
PR^C( \YS:Z4B3S^4BR.G]2P/Y^20#IGN\XB&$[3K9/Z,5@E^Y!B6&QE$(VZA" 6O
P>.6$N@3V7*DV>F[FTP+C! +,?TLJM%4>>./3,^ALBR4&:*SX2'UXY9$SZ.1X1?Q9
PH>8R8.DRM."0E*1NZ:&I<J9>FJ(];Y^SV[$^PCQ/2I[2C>@U-1QK&%@KF6U%"M"3
PZ6U3F='9ML$]@*202D.F#QDM,_-68GHGY"Z$DFC*.#PCP/Q7#-ZS@NV3DL@:#Y&\
PE/+*5T!440M)'OHK^L;@I+?^=Z<!=5+8.RTG-VBO&A<$ ""JF;B[J$W#IT(F1+2#
POR#;:'QW_V7K<@^O8KS<I5 LJ956K:*N^WHLJJ]5PT]5KV==!T_XZF[@S1YS9NZ(
P"]0 3>UXES&E]VSGZ9CA3X(<"/\*520 0L0>(,,IP$MYN6!XVAQ_MPA#=&<+N;\.
P:;=%^H253)([Y +0M!Z=[#*4+\1G>TR'7T I^6P2!$%)+JQ!8.7<_=:F357R/T1_
PG9?;Y#+^N/AS"!FC">@Z0^<=#6(=ZY2DK)XW<N1A"Q'.2"*X6^AX?.R(]L>KC9Y/
P.YDG$,8K:)%'_FIOPQ@NLM<$.&+JOIA0MQT"\]O/4L[+57;W+#%O*Q6J \G.#9N?
PNK*F0$)[ 3H[M_;IJ0Y$9EYY]C\C/^25=.S!-..C_Z)T?S#59Y1Y@%$'6LM8 ;BA
PVXG5DT3[4:VH$+O+D!YQ@6ODV *PB\WV5@O5.<VGOLJE65SB<:'/ OU+-W/F1:P_
P2R20UO7M-"ZX$QW6'AT9$!/?,45N*T09G!)K,E@;IPLQ&57L2200?9W9GFZ %7^L
P^"&LD2<!1H@4W1"?I[0RIBVS/>0'#I))6LZ]XM$WEP&=QO\-LK#>BB4)5^6)582X
P^F=?>[ O[P?Y'5/9\8I;)?,*LSSO4EZ^P4.FR@8"^TIG+S=.=_0P;P]YTI/AI'19
P(_9[69J#$268#Y5$+?)VS=)/4K=]K#?A5.V;37).H"&TA/)S?&GX;+]F@M9--\_?
P;</ZSIN47W6*K9!WUNNUY+/6KS0QW30B1"XS<08Y%3_8HV=400WU"XC#E@#;[O5:
P! T/,U%] 6\9/:KD'E@ZU[M5IU24169W,$5;K%\D7#/CQ82X7WYKNU).I;I6U(;Y
PJOQU#5J5'R7?4 >RS[W7<POAA5]2.-68=M>#+"WC)0PFX6)\T%ZS$L2%O1TVMVK&
PWUYA5!*]=\MF0!X(1 7=40$4<GQ+8 :Y\O 51Q#2:1L_N"(7TKN3 1NI-<=Y@UR%
PZ:\<^5I@<"V$QQ@ !W_Y)5AR(HUC97 +H7B7$VCC<LQI*ONK^*/)7Y6;D! :OE4@
PNG\D<QK)Q(33'Z56"-X<F,;TY=RS5D4W'I.+Z-#(08VA#"CAY$LJ0$!U-LO@3Q3.
PDHBT4B8)>EV/4J+V?9ZMUTD'BOR/)EQF14*(GO0LK4DB!(RZ\CA3%?_OO([;&T#T
P[":=:5*N;E-;BB]HM9 [YO,B9!+5 MH8 C&YB6MHQ8[3N@)^;69HF)G"#1-@O ?V
P6BLF09XA#WY>:'<?M2R]1K7&!)=[R=%@KWMFBU<CJ=!LDBHQ,1C%?JI9!L#9DWJ3
PO*?#06 W6!FW\Y>0KNV,M^9E7$@Q<J>7:V/M[#[XE>L8IC9FWQCBA#Q!=VO+!31@
P:W/O:7S][_9'!M_^9$A7.T_*DJ0_G:*Q@.R=^1Q&9IMA:<8D\+!1LD_('$3BI4\;
P=UUM(+\#W5>J(0UV1)QML+] !Z$(.5Z[MC3VJ_XXH8[6"!'$R%.6I.*PAW+ 5O8E
PD'P62J[:(5DHO$82A;D0D%S0)A>\065*7^!A+##@GHCJGD]>@'+%<5%)3*@7N*T;
PS1A4Q6^@*(#%7WZ>T:E]-LT)>[LUU(]=^&L+E2_P3Y*!W2*,9B LU PH6\1Y"Y2P
P$.KC$!A2^J6.0N3',$P(;J)NGLT\_JS!DG*X9I.[IO*\Y 9>Q1T0!IU"&FJU@%E!
PT!OK]%"S0H"5E&R4@'TN58[I/=_J;N+3!<#;X&OG)N\E68-)C0&<2:RAAYANGD%!
P]]C+T2>(53I1'QY\LS^D+/%'KQ'FBWGS; H2=V^]@\E(PJ]"J*?"M7_!X.-S2<PO
PE3P&&$8I?5_'74=GH-4_.G*>SYZ:1T?UD7@C_#P8V*K5)>B;R\=0P0'C$IJK X?-
PZD#>9JN$"B?0#S=NY^C*H[7Z>F<^__W&)X6KUW?[M@M?_AJ-8^S8<)B@/*>C>-^,
PL>Q5N'>I-9\5GX"_&>22A<+7]-#(-\V#J\@.&\B\C!B.QELMWRF,?R"U!DM..JB-
P?[=I[0MV& M:5/5N839\RF=R32_H1$N:Z24270LEQ'?1NVOHR",XA7@2]T67'P8J
P_--%7$T*#,'A)Q$>F,O ;H?09Y'(+()M.-OZ_98P?Q29PNNO(V8=0PFB1N!A?Y9(
PY50J6DY;1A, OL""7.%<JD ,1=?@14XW4I,@&,TR$99_2@;6VH-5N%Y7B:WVISP.
P*F1(59MS+H3A$O7\@"=;FA0F>B>&8S8ZW/%NFPF"W71\AEQNR0-N\@5N%,-"WW\Y
PP#V.^5[(O*J=Y,.RQPY_I)6S<\]UZ6A]'*V^<1N(EAN%O-#J*YXWTL;#1U_8&O"/
P&%_%1M)<RUK2NJ*^5CH'Y!P7W9 H%L)E=\\$@Y6&#B;0F)S6\G:.7V:0*PY1XHLR
P(9GOV=ZG3?-JPV:V7-U2)2^*ZTT#,K;Z2ZXHS J.)=D%[C.8UWH$.JM_>,14)H)?
P: 4#8R;T-AZKBN\KWW93^6I03DS1+-MAH2LN!3^_V)[ $UWJ#$HAA/(?P;RZ2QUR
PP[R948A$=[H>./""%]4)P+DJTD3:LE+'1CP/[G?SBJ+$MM/@C@C:P_B'\_Z2J7 P
PL50HDL'V]P#^M\![<#2^E;$D(@31R4 K3Q.?^>[7U''$*DG^U:V$1JJ?D>**'#,S
PIQM)ALU$.40(4C#MRL#?T<U2AF,""D2=X_:JF#HH9E\GV5VSA0\1@S?\(1C(1@RW
P+LC^4VW\["64C<D7[F#O(3-V0CW/"D69SHAA70X[IN.UZ9J1DW$1?1+SK*RA4EH>
P/TF-+EL?ZQ1B]);4TY2]C"5"'4HI9'6]-E4R]J]1)K+Z,BQ+U3JPI9MC;XO(X=[A
P9E&'QU]/S"Y2)XI9;!OA&6N)>A+W"0J4J/B-;"+-R5@?/A,-RY/*9*%DM"[2^@(7
P3)1&P!*YP'C-1J-:JFW R4 N!F68NE%MX_-#KRT/</:FK"J*OGI?WD+MB_,U-#9$
PCU;K406FRFVLJ U,^U9(%W;)$NE!Z()/@WP?A(E6M?;V@8E*!*7"WF^*-/QO7=L^
P^QB-C>_.N1H2,MR0 ?JSDZR=\S@V&= #62[\B)C92PCOD 6!!F1?H@90,YJI5KE"
PY:)0A35@H=*' Y/6C68/TO&VP(<8UF1$O/O1]H*KJY:6WN?W33G#>%C-YJK<TI;"
P%?"U,W@;2']))/V>-IVB]4$--CWLGY"-AB<<MQGHY^72&F"5T'VIRW?1:E213):;
P<$ZHY!Y:R^4B2S:76(MJ@,OQK 5PS:CK"VX)[ 7RW$9O76XWWG<MJ24,*CF(B74*
PH=;C4F4DOFE2IVVM6:IUGVK("&#*';C:/\ZY'XHJ&!-H&#+HPN*XT_GZWX)9[:1+
PQRXX\2.U;<'Y:A:J\T0!>&:$E;6M['%04IP&0;\/TY$FAI2PM# <I("H33LBH3@6
PA=512@L]%.\A.!%)XK7AIZ5OK7._*HZ)7ZBZY%7&@8J.IB "/RS=R6P]V*M?JYY3
P(,#A?O]=1\7759$%*()%F5XI)UCW\NL<RO2)]R6U$Z1>+N_/+3Z0=9"0IES&)#W<
PI"=BJ8%D0?J1_\LC[;%YOYCT$DX R4#O#XKEVYB4RCI'O ]C[,@!555-_7 ^<N)"
P@Q&[5^*KAM36%5#L4[_+YG=F*%:"!D(I ?43QBK5^#:P_Y<\\YYP#@_!3TEC+UCL
PB>CG_03HYYH&.]UJ(6Y.CIH>F;X$X_;M7*S6G2\7OX*:5Q]]P<N[^<6&BL;B!/UP
PB)Q4*W558$A3#.02$3DN64/Q\JTB#%YA/DM;1$W]\TG4<%CU_172-1F8*/%RAX"T
P)#4L(\,]<8Z"5^/<?E0I'.SZ/N5=F09#UD3,TDV^XJ%T+T^RS _G[RLKJ#,"N!T2
P-M"Y\@L;6PC*O(Z;OR BZ$&/BJ<9D/2Q)W]^LO+=>0F UQB:4HV?Z\I\6^B0 +6C
P V \/YYXI=5!$H<_U(LH@T@:!#M,ND*N9Q-$?1E0]1<9<"?YYN(<./JE?GLS3;#=
P*FLJHWUL\DXXT-,(9^DQZ-Z?T2R551?.W[PEWY9\:UO50 4< 9=(<SM?<4PQ*EZ9
P2X8#@5R,O"K31=%[O"FP(M>L!23DJ-?ZS7)?HS'7XQ4^B:?B<N%UZ?[[ 15Y6F?X
P?UNPLDFI:6P>\LHX[<5B-0J>2H3.S*LZ4.R X8[I3-SF'C<:!,Q1V+/[E\EZ^@Y?
PI];.N3;]$#OS*UEAD.^%[->7T-%YX__BF&HISTA8XI<-\@Z+[P'2+=Z[B3/ZO;%W
PL^[#8V=^EZT-*;"0J!H/-#BJRJG&8C9,^>0Y.[AX@M"'!)UMF 0/8W1BV&63)F]_
PIF/_$0W^*50&R83,MU%R.S.#,=)@KC](62!PDY3IJD*QGP"<ZG3XG?B\\I4\X!WX
P-/!#0(AZB&$H(!%8/-HK0^/EW5V@V/ <7?L7+J'XL7+./_>A4W^72A <_4,O4/"4
P[7^3CX'*3W?/;ZRGM:K@E"8XM"*%V.E%\XWA+*NGN4:H)5JL#=2IV7\#+U"+\]!:
PKA[F$M2;A?Y;;7M@]3?#YRF+%.;T8,VEB&UML((8^PL*'LT\W2.B)9+5&[[E5??>
P39<V0\[] $%)JE3<ZI5ZM70>:S=7H"E-9)/8@W*.XIUY+)PX@2'\72M**IZWV-E?
PR-2,J>K1"TP[D(EID'2T1=_!^?P6&MV>48;L6>.DJRA=+1-RHF96I6%0,=,!@#(9
PB5M?XY.B>W5%>D3D19F'^)M,HW(<[WV0F^;-X-V_G.++*X[8[X"G6K&^<O=(.T)7
PEF:EA):58[8R63:EY+?)DI>T5QV=6H04 ;J0\S*GP$SS H-+.SYI5>5*E>)AE4X;
PMIR,$D[7) "J[CB!&/[-D1RI=,'?,[[^<2?;VT%0:%OA.AT2\?7 ;K&2FA](.L-X
P-EZ3>X$@Z<@.4Q5(#L ,H!?"$8%[/%GFYQU^X\I\[A17HF E[B<3__E5VHN'641W
P *DWL6%6DV5YZ#+%R,UD%]GU+=20,/3^*B=A>].Z":Y^NW7H5!$D@E;DEM\C57Q,
P[KRW<6RY'=7UNVY-5U:-<'&\HD0AQ<WKYW+R&XL/P73?.E)7(3(<O>.8E_R&?B[Q
PIW<U)JU:IG;HOU<2"\ZPI!AOI/X+;NBLEDJ08.WA//\A>R3F!EG>23NY!\HE;(^M
P2W''R3;N&8IQ)ZGO7Q':"4420-'-H(&OZ"_ O%;%R0H@JF?U'0M/D%!(X6RA<3;P
PG(K1AM!!:C6RKELO*0NL"T:"+\$<2>\4"Z0YCNL6K,_/D^.7%B\Y\J5%!WL^KYVZ
PS$9TQ4Q[2SS:'2N>_ KP8R=B0S%V,:K/A*;# VE@)X!R=&?I WVP^3K1 6AA$RXX
PG>@5&70"V$P77U$,DY>I+AX !4&Z 5"3N+C^.X+( >HB3.YP=Z>#Q5N$ [YL^#F*
P2V/*5 C1P]MQ"5.Q(99GO;ALP18>IUSW2ZE% /U_]TC&#6@'];4,0]Y7*?;.*8Y2
PC[CT%G-H.NN[]70N&X" N:MU[387 GR*"G@POR%$<G:.E^@.[V6#H$9\F$AZY8Q'
PI"QZNS//I0@@AV.W0B9W9\45YKEN[!,Z;QMA%Z^,NNZ+K3$ZDAH7=4Z:O.V=5?7K
P6&D#:,RPKL ]&6_>&U3Z>! -Q_VLVBY2Y+%53JO*1@Q?/FB#O<[A%[XB;;\%5I+"
P;OB)0K)VW<%#H[M]U@3F[B-,?F)<,3'5N+\,M;CTC3T_"2@/-M-K3RFWVN>+]$5T
P4%UR-U8G(Z\8M>5VWA=A;#&%MN.)OS&P]ZS<.@"N*LO"[C$EZ.I7<K3RI"J>4X]:
PV>L6*)^ 29'BB:X,R@\K8PMVV)'>LTE"WKCMXZO*RK&\8FRB&2\Z&CDA(HU169UX
P!'MB&D1CZ-<BE"8[> @MS<B/A8EI)CN+6^-U8J> -)1G%)&HV8WJ3"P;FNX,\FV 
P$Z)OQ/5,/49#/@C"UD5*;.8K8I,V-2,AMN.TY@G^?Y%$?VGJ("Z#B7O'?!7(*+5]
P JK4AG#;M,&'\<^7=U'9L_O"NJBLJ19Z"'^/F'I=[T3$.&&37/,-X'&@4D8FEY&_
P,JPW^0:$[G""84RYY*Z^=[=;75WG/89MBBX#3@W56MR4/'QBRM;FIE#@'?P]?CZ)
P>&Q%#O&?U:05_*^?L$@UM7_/ '=ZIW=<T5<'Y+<N(V:QH\RK+(\7/RA9H/MOOL!?
PX1FN6MH.,?%FE(5@ ]>1PA6<:0.'$]*)A7=)8I;\(U(1K..F#)&0 ^>>2D>J^<\-
PF,0]%06,O.%IIY0>LF:R-0$O+VRL97Z9#K0M25HH'UI+J/^FNXJT0S0K .N]@K+1
P$6UC: SOV&ZPV"D4/NFF. ,A!I/8YU#X'#3&G>2Q,EVQ1PBD"@Z("->!$$CM(B?7
P'%/W]D?2G:V'!/U[=8Q R[KJ$"=1N2!"IS3LP$ 5]*A016365?S>40.[[_2EALO:
P7JETRY#$BAAL[OP.P6"1DCJMH&;RSUX&#HX@39I''CUO94M^[?^09IMX_XKXY,B7
PVFC3E$K,,]OJ7N=U)&(6H]SJCCR#J\KUO=9G%5@U*&_50NEQ'.O?*8IPX)+]-]W)
P<-AQ,49S?=J,.$4]S>[\;,PE^!&FD]A[_,7#3IK)_]2]6R.LO C''W=(!\P4XT#K
P6(E>@]P'+6R_?50<2P?G)), WI2D]-XOWSA^G8;7'H\Q'.^,&6'6#^DWLT$)VB3X
P'8O26(:_BW+=]J$=DW29;T!F:F!O9^:D71_P2#Z[;C"528=08$8CN/(^[_9K>?@@
P9UL6V=M<U(IENZ9_3FR'4OU\X-U?%KM3-C+$'T)@B$ 73AKZN5%2=T,PFABIF&U=
P4D]'%%[)/;\QPQ^O$)@,2@,G[I5,N 79#T)G]&XD="C'6% @8T]=:W8;)6[P]']]
P8GQ+3"TX(2U:I3[-,,X+*'@;C>'@T4G)\17ZEXD.24U\*SD?[+#4I.6A"G_2!M:6
PKM6&NQ$F#\&+^/ K(UYI'%(-I*G ZB/6MWK;"TYESY["(7]1(S]]ENVUE2>@>C.Q
P%$X]O]'(>1;+KSB[:CG3^2179D\;0PPW535"8O;4IS+TB7LQMQ02=3ZL>BV3DG,T
PD=][>C4GL/2I:%07]APN[+4TWT.'(EAOCZW)#2"'D\AVJ$1$;/F0I<Y6+6J^>G/M
PU"2AT+?98?Q!P)J'YD-<5)SJ]CR7N=5,3/.(AP@[>Y=B4_E>%2P,8V+66&#<_LB7
PU<O_+#6]@=\DJL<8WED[M84K*$K$=X2+XY+%]_[F3$:VZ],OG["9+?#D,#)YBC;$
PWY^.9>'&Q[DH<U7 ";.M]7M."8>!=+70P#HP;).I0(X55=_/KTC2M$_< T[DU74T
PR. E-<,!?.CDHXN;@4V3I)!W+.#)LK^6TO)(ML8U^=D6\K"F(6")3F@-L..& P^L
P7$D(2GQ 'L#)<@0C8U4PL/K82",P0KFK\?3S('=-<%Q\'O[^%NV>HA[@+_YEW*U>
P\E^*7OE)I,3>(%@RRAXE)&$^WC]<P;WTE;\'8.!V'_34YAC4.%-L3J&Y0"^Z(O(4
PD@GS8L<6VVG8YI'F]?.@PKS6N%0GX,R\KB.2D6U_NAYO"% YA)$.>T!^$(LSQ;5/
P]5QU3Z$Z8TR^+BE;QOEQ6D)1Z4 @+[X@<$>WVWY;3E8CH35C)[N@G-U#,T89^P^^
P;:$6 UG]3(!4)I@R+E85[=$6'(D8@R;&TTHHZ//C'<ACA?ROJ_YYJ;0T]_HU95'L
P//A#TJ/>Y>8)]]3YSC,JV"H+RK 2H?^,*G3?R>6F:M5E%OW9K-5DH)FV%5!V+6YV
PT#("8F'77P*X9[.?'!H=1HT&LEDYZ'OKTQ\1"SGB=")G T4[< 0_M X6W^*9 'Z!
PUWK\G[;Y5#WXQ1:L3\$(H+G!ZVBZOXY=5\#[&<=Q$BA)A'H@QEC7$1E8<+E'.Q!]
PZTA;J0ZL3)'X\("KV-GXD*ZJVQ<B4R&=KVS0%K X>Q3OY=&_%@\7"N.CG?EKG<SN
PUQ'1A=8K"-KOM"OTJ2]KE)YZ"!V(C 692H8Y-F ,L.GIBR+0.!2[.9;9 L;@P)"K
P3GWDP"?<% "YJ!BMU7NZT?/>*CHEXL>Y^Y>TPYNCX'>X,BK(CDA'<DPMU%_-DWT?
P4*LY.W<IK!-=96$84A;?'W)38**[/IFW.E1/%?I+#DUOP@?N4M8&DGU7,K"%<T)>
P0N\V@/;4<X%)2?\[!1CSN#S&56^?>N21-XG\63&[^599M-T)1-P,W]SL2P<RZ$8^
PQP.#<NG;;*]Y 8?>*_I(0H\/4L>H"C-!ZB427^G1L]?:#%O<:.VO<->/)OEM%UN<
PM 2BWI>\?W>U [>9MI(37.$AE([Q/IT#XF":/<1F?LK;IG HYF$/2D'7/[.2'_PW
P[]LCQRI<7S1%" 3%7**9*/2V*+AD4UDD47XOD-TI<2U]&S4&6GFS6,J@>-9X[!^5
P0<::+/D6DV1^;B\<,QES4&3W'%2L\K.II:G9_4NO^_:!C&GOJBCKS\UM)\L&( ,(
P>"? 9-E?\6:0EQ$/K&FTJ>"A*E<AB/]<F09+2A[R=5NU,(G<#D;/-!4#E><M-2><
P93Z_I8*_%2'IEVF<L[!W1G%_<D=HN2'UG ])],@WU$NI? %L@ &8.OUH-+I!4K5.
PV+:O\U!;G#V?N0N"D6=X%&HILX,!C!E;]$!T1K!ZB[Y5X&F_#E]<E$+UWY.%?6R(
PH'97WX*<"5@'8RBRS9+L2L>N/!^KD.(E[T17VZ!XTW6Z*<+&##2'2I_Y[[XW2*4U
P@\CV/80S]HZAB(ZX7Y#3X/I@@M,Z1T(TI/G<)!4Y)3FO\B\?#)VC)].^ GHP2V\U
P87(H6=4<7-LY#5#J\@^+/QU3] 5@\;"/"'P>9/+5X_V1ZS3>0YW!:"IP>^D>$IM-
PN!K!*))X$D^]RYFTQB/M3)>-#6'ME?%[FB+*BP;1P[U-]N:XQ+&+HN@?_M7L9X!N
PH.K /_[O0VLX'%2SJF@0-)"4F,4V_=!.[SV!-0JF"E M^[<V%+L9L6$T&&V46SHT
PIY2^"R@1-@QT_Q:,&JL5.#9)HBR-FFI(VAH>I*-[EKN?%]2CX8WL826?A JN%F]G
P"@57LDZQ-R!73.BMQ%1OU1STE79,<Z(5^;POP/<L;DFYT^6\?*_A97HY>N=5QF)8
P&YYF4DR$^A0-/H;@[*RS>8IB#XG %U0@@'_O:[$QM:.YC8:JPF>_]!AHJ0&@'/,;
PSA@T_S?&&[\+:24@U2S,"3U(N5#02;#MCCNI*Q#*& 483CPT%?X[S53FRF,\3#D&
PC'92?C#I4K!%YJAF^MR5NM@(3X.>HKG.KP=M8O+*A7$C/72V-M_3@#.>.2X6T*'K
P5N<&AB7N!)SW$51T9C634B^)S/A3;>EXDZ6;_V;/J4#V6KUB/96N4O\279D:3X5%
PP\D!N1I]6\KX4GP";"N><:D341#16=]\Y8>>^VJ7EK<SB!#C&)?BZ)<8?_IE-''A
P\+*VU6(SW_K]BWA/(,RC/GFL2QUP]W1B1S[#S[>_F25X]<\_+=@"RQ0LVJ;)I0CG
P!=]=D<V1NHWUC'ZNQ22D?-NED@5Z:UK2XM##1YU17:FISC4V2R-U+-$C-HKR?2F^
P6PX4@@ \7>,O6.W_[.L\R:3^YV#0B8[XR^'I;B(9%L]G@]8##N;)HC/7W,N_8E=#
PPP$O"LZ/BT8$F]/OE8PVL%'?/38%3<'.61TFK6FZX1&!.NJ;(R_[873W.GG1%:"M
PR[?7>5&JQ7=-A,2H)E!2%&>D=:VR>P(X=\L!24LB-&] "/SP?4U23@0JR<UR[5&(
P?Z SB%D0,YCB)I<(YJ;+E'B &)&X+Y8:PY]?[5%Q![[?N-=(;!-1)ZR]?G7#E_F;
PU#> 2-N,V6%E(JX!$(SHGB^NHV,BX+&-SPL ?/)0X-T2"5@P,H;POU/X6D7'F#*"
PWI,'PX0'K8?,3_88#-YO/5G!07HYH8#%KIWB: R\%>;Y\!AMXC)Q]AZW=5?:%F_8
P#Y[?@YGKR?K(4<NZ3MU)2>'=S'X?BDS74N!YCK5Y0J5:?^3)?\"B:\N(6TMJT9O<
PV8 ;52.CFMO4&*<P=2E@S"^PF!!$-8#L.W&^@SWG^Z V+J9X6[87W:6@8V0S0N+U
P%1I:6S.@">S93QQ^OV:',%.#RM:X93A?>7Y@BL2&;#"A6/!" 8[GYV')1D(:J+P?
P$U6M&5U<:5V,-(C6$9NH,A3!UY3\5/4V_!K,KY,)VKV9+FP5'X$Q_6@?T^5R3$K]
P :BF"\D52?#;A3XKL9"FCO)$ID^]D!A%K.+8'QEV?B=[0 SD]NAI"NFE+\ZSDB=X
PPE\!0$^"?ZB,D&CSJ?_G^MJ9%"D:!M$=5%EZQ7L=2M;[^I)'Y//2J'"P:8][8-.&
PPPA^@H!P=2A'Q7CK A=BNU$B7K=>O#:;H>V0LB^]LL] 5F"&,8GEC.KHM1IH?,)P
PH^GOKV6L^@AXN&$:2+YOR0)>7#7)?CSF*4RBATN=.(XP0Q^E[SR@6 E.X@B&EO+G
P<I;0,=CK?))1/S5H+H5IN0!R\#2&\OU=_'="0IQ$[T8QE/YL>\,#V<>8S2*UO%C3
P*IQ\^\78ZH!"0AYW:3J1B:<"7,%H'%]Y>5)6C16.E%B2'O*,,.;-KK;Y5NEC#TH_
PV/@>.?(*O^$K/D3;B,A^.6\.8]';8#\S;TN?HG'1Q=@%+B)"ZJM-"$N1]U&R2$&7
PW=9*@S7J(FLH8HBD-/_OYFK\<2%A,+^;&_((R<GW0_[_J4>U"?TT1:7$9LP5[CZ4
P,A%4X) ,AMY0@'#=G%A*\Q)>2\8ZT>)"1_(N>YC98$V?_:536_-OB6'^F2?U%%$2
P!\>J(W4G/[FQZ&AH\A,9B"\15\IUM=2;%_(%<TPD%X$-D,XQT^SF?\?8[C41PESL
P[_8WCPSO:\=HQ-35 S+ EHE5GHRJ_E08,NF*%?(GOR[>ZHRHD<M$@OF#@)@4GV:Q
P1[\53CG'QLX"L5H59,$2#P-+M=U]*@I0&' DNEM C_-UN<;6'&T(0U-M4T<,ZV [
PS\XQVY>@^8*0T$;+5!XZ6ZY%S5<0_JEP^=G!P3R\7V@(VDDF16'XGXW2!8&PRMEA
P>)WBILD#<EB%>(OU?_=LT?4;3F"P$J#T=72R#EZ,,>0F0+G@>52O)O?>QDX=FT13
PMRI07AYU/G:W+$3+>NOM^0NT5/FO+8%.6KKO$/4("[7+!(-_77VX1$5; KGDA+2D
PR_5R6A;@Q%,V2X@9C)[M]M.D]A\A.@_$R*2S M/@?G[N"1N1NO61X#TIBK>J%9J[
PCSK'A)-)8)4'N :.[0MUC$PH*$*:]0"#V/[NA(1)P/D("LT!QOU_9:09'N7H!TO(
PD[ VQ"Q3'>CP3UH\].E;FI)_<Z:."+'3'MC@04+L1TI; I5^P(T$*[+"CB;MT5MO
P.8FGL'#U!FBF(,YS5X8L7[L:$0>M,J%:](<:5K8N4_RT:QLA9&1ZARYQ=%#CRS%L
P%L*:_O8JVELA=C/;LJJ1@9<$K%LE /[U+M2$AAN&*8R?7:&*^[U(>.$Q=*BXR;73
P<)Q[T]:4:,TC5]D^/\W%&LXL#L)Y@*L]5>U?F0PU/W!V@ J+,C L2=_")B9].X:Q
P9I#1!+NML#POUUDZ$;\-GP>$3LH#M(@*6RH68&8.\KF>3,?2L0C5^$E&/)Q84T,+
PS1U(Q4D$0Y,V+*.%N*%A316ANEU>T<__UQU9 8:X>!5= FU-EKF_9TD%/:74EDG%
P0_ Y!V-[.]FW.ZTA;-OBC.;,[1L/+7(9UD=E!N'Q39U100=)B7FE^QV&&?[G6GEH
P8HY!]F7P22492DPRX0HYD_Z282%B(%.4BNL:.\=/N=$/1=Q)8N\,>N]9X!=9)M!I
P W)\V_]U4<0$N:6!>-8V+?%=[I36H_"0C-$+^PGCEYI;:"L>_..<\91[4O%8VF]%
P]JK7T\3&4.622^&$%RK/.7"2*I^SH#H)GF!02X)G/X30C6]"8T*<.H68?S8G'FU?
PQ"/S QV-P,H9VR61QUOO)Z>ES=3@SJT6>EC=HDAQP?7TM6<,>P";=Z.FA]$^T">(
P+EE5"Y]'H+Z .P.UA_E^0NY0-(+U\??@ZK,*[_S?J.GHOGY ?*AT$K9BEBG"X_#=
PD?N,'7Y\EG#*FUQ;+/^O0^8@,029;V"V)*O0-L/,34F-A,Y>!E)>LP:X__@DJ@@X
P!%%F_':R*O@A;JMZ3C>7%K'C!F2>L<YOV=:"_*2&;+R'#]".)+6-YRT2C+SDA!Y%
PL[?[D>]JCS\^VWJ*1QW"?; C[^\_R,XVC!+-6G*;T&EE,.])LZVMZMT_Y74S/FQ:
P3MS%\)OF5#L@Y"_=P-VI[Z,8Y6G'"#28F'=M,(O?X@-2ZU<ZXBA F,.Q/\VWRT8@
PWX0'WX191>>.ZZ1:>8RK?^-@-7?D.Y'FK]=E096%I4,A-*O-?.G-QXFN/ 7C CT2
P:^3.*<JEN,U:8?H-R">#@#V!7_RLWD]CD.&2NV.F6SY?Z3DCO.:6'L60N&3E(J4T
P*IW;6/6^G*(5/[M(Z QR85ZUN=$&[8A\ZES^H7%YIF9,RF2003D9$[0JG%;KZPU_
PX9D((Z'_U]+>0.H@J-I9\N]3W"2__LL5\><3O1_FE\&3P/[1H^(PF^5N#@QT?'##
P>'3R3/S"13\@S*+&J99E(6V=_V^7GEVKITS_6/=#._\O8L2'WWV)FP&\6OOYH 7#
P3_:4:*(IL<^+#A0 B%C$,6@W3**;LI+GI=(BL ?H/^$M1\ -_T/.^V0/+<1Z>_&<
P!M+;QLL-IQ@IADF!\+M$Z1A?H2U DW71$'!)0 E?,!3-EU%S.(P'<UC?+JZ%3O@^
P#7JS,C\0@$M0%7:XC8 E%M"NE>9F3S3]>&HU-P/T &C @6:,^>!6,)G<,+Y_W[/<
P]AM^1:4ID$LZ><-OWM=F^!,QS)C#R<8MKQ_. E&Q7;&^%58[IPB%H;SZJ]NT#;R(
P^.;*L,+NJ<$;]TW^IZ:5#V?R!?^<![0A%_\Z?$]W7H$B\7_F&:?^'-7QQQ-*T=!Z
PF!J*SDE1MOPB)5-:8Y]86N MH4X TAX=>0\),M+B*[7ZMQCEJK18 7PL"K,%5JS2
P2Y02>:PJZV%UT$+OY^9J6"[/>&ZCE*N)VILPQO.935C\6J/J=E"?G"[M%*B*WV>[
P"ZMNPL_B<TR+=;?C*8%Z8D;@>17U(O>:C!.MY=QR;SU5-7BB,1Q)4[ZM1A;%117)
P\K*62?!VS32/4<""'6@_AHM6<TW<M#GMY<6O\RWG02<6,CLKA)?) C,C^]XFDSQ+
P&O[*[@F#DNEL0:J[!O_ TA2*]:OIR.=BV)D*6AN\IHL5JBA.CAB 1K%8\O'SA#V+
P4+Q0/Y'JEQT@]&J]8JVK_&,D A@>-_?-OTD"\H&4[HS.?Z/GWDB^?'BM)F=:F+22
P?O,W02'3-L?@3\..7\%[^HAHH!<);Q5C/H%88@S&#$LS8"!3-9[K)/34G%N+#U/M
PJ^^&<F?)%H/Z%I,*B?JT$6HTZ;>YQS+*G68C\ ^-9-A]DQ@7KLWKB9Q%CFJ3E_;W
P\MUR55C4:G5@>-,Y#.-%0>+KL:U3!\P@UR")7@_'\,,^4^(6)^,9O\L]7V-YXM*P
PY1@O1[+1PAW_MDY[)+O$&6EXU[ONN#O 3:U!K7-(G6!F WN>9"/&O;:X+K(6U?Z<
P&RW.E @<R4.J>O@J^,9YY\"4IR=-['3?OT>'DO<75LVBHGLG F?;LB,3WJ:]0K2_
P?VHEO&K,1OYNBU 810I"U>@/+.WS1,E%S"9FYQ![,^>EQE H'V!A!.QSIF79]61L
PG>(!C^Y+22\VB:/'"JDKLPWSN6@,="#U("FCBC9C;&6_4TUP)/RHJ[21Q??RFQD)
P<)8?\.\&ZMA++51E$^:C6[HDY*4/>6$/7UE^%&CW7J_R$U<B(%E&/[.H!N)L.H0U
P[=2)8#UM.-1 ".VZT-_V,"^<!](BLY'Z$6BX>H(.&7;S,6(!T"(^!QN2??+# A6N
P( ,;0#S^?[VT;"*0P>G!  =]0-W:FNZ^537+V A;J?[O>F254Y<2=R)SU )T<0( 
P-ZQ=5"QKSEJERY@_^EE8/43RODH""=29-<N\PT4" /M(WQ8*)0,$KI+YKW>V"@;L
PJ*\OL"G;U.@\3:T[OS5(M<5AKF'C!D6?'$621N+IE[N H<!:+=0R0_[QC.J2X/)D
PY.*J\9+08B8S!OI$]>987@_9C905IU&^K6\'Z#.8TBU#X!-@TQ/D1@CX[)N%R@=E
P%9J'A!C4A/(^+L;=7>1.M-25&D&%UR[,$T%*LN]=O$$0V\QSI)QINB3(('(@$9=4
PG11!#+2B]]D0*?<I0W C6&76&);G/6YA.#'Y"QJX^39#&]QOL[JA#Q(JK\L@H:4+
PB?"0,Y._GMQ*>DH++-M'+KD!VXU*A7UV.B#^LPB&N_($E,LH-A,F?XJ^H.D1 C("
P@#Y3OCRQ<4MHQ"6G'+-0D<EL:'?=&R^/S-Q*U1I/-YQ:9VR0O3X04.HE_1P1!K(=
PJM/^5Y>\9U1(/_5[?^X=PU5;'T^><8 D!#8G!T?3Q1?UK,T-WP+B,ZW@P89W&1XU
P;/>402Z\XEOL$^3Q?*< (5#(;Z@545#V9^=P(UA2>Y-F+*5(=BN$UL;LM"*:RDMV
P4BU7BXD1ZES/*FZ*[8;#E!3<$1Q>^Z16:#B5%:A@PHL<ASO).]SEF:.J9!'S4C4T
PN:*)XVX^H3@/]?Z%Q=FC]^7,;?6I1X_DK-B+6BF]<TB[(ZDJG.ZA!Z8GZL-?+Y"E
P5.KI0F)5H;$^J6"69P^8BDI"-60K/_$R5C+0V12:D YD4VA$6"1?7KDK71@"[Z3^
P@F6)?6P(CH EYRR!G&,/_\:C3 *- /)O()M>\CP2(.-R3.- /K8B-/ ;\"_'TCKO
PFWOKH@3P@J29E)\@S&$YGD,9<#LY+Z61L01*-F"IVO8:;;TT.7A(>"S)]RIRYNBT
PNR'+2:]/(_[9O2H'O"L14DW:G7%L%MV>0CF>5AH<+> W;KC!!]\@DWFA^#?5 *E:
P\O=\B0-^7.FY:RZO\^R<..@I7[A+IT2:K3#/>J@?_#CJ7;B:<%F;Q2OB)-[GHW \
PA36S_V-OZW+C0*3-PDC\9WFW@#76&]I6ZN2FN6CU*.)>^2D_M":! %<S/,E0?3&%
P/MT?'83\.NSCU0D;T @O%D8&_Y: *=*=*.A%IZ62>0O_2#2:]/A^L1LH@+RL'B(/
P+RVUL26VEM<=F5VB=E)W- B&G[K&PQ05:(;Y37I"Z>VL22#</IS$,J>1HW*]+!B!
P1#[GQ#/SR;L.AE-Y?'ZY@'H0GG0[N%) P2ZR::'T?]@7J!@:;'_EVI^_ES<YG>I(
PRO&1KR1E6J(ZK>2Q_$M%ANCN"D(]$9#M=K)@&0B8(9V2BDS -0>SM(*A;X9'%(SR
PAIK5L!4J*E6?1 X29N$V36]\8WE-G%[J0\#R3\-%<*MH<N_DA+<O.ER_55\MR+6)
PFRU\@>,'U*%9$S1-N=4ATRY^L4BG>4<*C0;]LY,R%U +70#F=;C;2PLTP=G![P[O
PDV>]#SAK!B&[CF?P$[(Z7%_:6)WNT$^X-DK+_4GP+!R;XH/K(YLZ2GBW"+U[]H4Y
PA;Z(Y +I$ID&(A_Z#(^"$69N=Y>GO#3=&0(+T9RPS5VJKQYD_6B-F9AFP&R)X@/V
P<R!.=W I^EQAX./DE#9(J&4@U%9!.7#P6@RD#I/RVLXQ154UQ\K(LN;E0SBX,-=A
PG.7R%0N]H''XGCUF4L8]P0^QYW)&4N1ZV+ZZCX#I./OZ.\9-'N<\MT>-RD7 &9:0
P4DG<TV+./E3D+*'/5<$LW\%R;2<O]96?IJ%X'56KQ^CG >N>^7CUM[0C"A)8!/V_
P;#NTGU/34.8LJ!&>1(+VLA9>SM4%\7*%=.:,H=R:SG5M4V8BI=)I[D8H;^"FLGL#
PU76!;H-DPB;)_@?/L&$JWG[S9?[:L8BQ.#BO8ZK\,Q LZ3;"=Z^UC0JKK]9\D5Y(
P6DHV52QRN4<&AV\^*2D?\K%WI\H:+#H7LUC"A/]C!AL:]<A>>>@U]T XT+2)FRXH
PM9-TRW."M=Y#CNK)/1># X4[C\:GO@H'$Z*GIAJ7<#JZE&<LPN3.%!(=;N4G'@PH
P!OK99)Q" ;<II8E=Y7 GO>.$788FOMC2I<_=L",)5SZ?+TY@O<I3(WWG"V9!+KI.
P54]3QR;;EL#%>K&S?*W\?$%XJSFS>0*ON:2JE9Q#02X)TK0 $7E3Q,K[EF9/RT2R
P;63@U?&-_-<CTF.5F_NZUG=D#94./D)/$TC 'BI;%C2K?>I<9[OEZ39-)CJ3.^I,
PBZ\CQRTQV7X^*QLPCZ%+>YX_ E!DR8@JR8&IJJQ6PIBJR&,!XPTAX,=4V+?Z9%3G
P*CT]&N/&[*QR^ZN<6</3&"(@2Y:COU,NT<'4_9%"1*$1KJ&H(.[?]]/9CW(Z-5UW
PZ#Z/DB?WB"3YFP-^(?7OVG"4],^RERY4'^B&$91V!,(SB?^</.0PCF7T^#Q,B3W^
P4SSID1T+^E!];W%+QM/>I6.FD:E1B6A:9R?')<2?]3^!_Y%"DP3$SH088ERO>0I3
PASMYTLFE(_UQM++QX3 (_Q;1U^P[-G2@G[P4H)Z:4Q-*51D&>Z$H:C.M%@1L7BWG
P<X G)L8$DU4L9N9%K 7C&UF":Q:FJ@45C@&@W0]3;,RB@#X'(O/UW%S-L4'@:??%
P,LOCS9!T0\A?T7F>;(* Y;G<Q0!#C"T=V"3BS==B=G&5/2!4-A;#V(UKU7Y]Q7^[
P,*7-OI*YS3 9E_O-3.N3I*G0Z68=["A<8NX)FF%?/&0$MI%'-N!1A;&+^@@126%A
P0GYF APMB#(*Y])C\@+;OZ=H7F[G*)TL"70NU\9V/55T!-M?&U!6$PI@Z;5#H$/$
P4^"L_"4N"06;47 /)W0 $W\?PA?=<TXG6DB*V;-.15OD_GN1+4TP1;5=T)UB '2P
P522'OAP2><(Q_3H_O[<*GL/M0Y QP&WYA/8#XVCT* Z/V6646G\] O SDK12@<7K
P%,GGG'4)SLF,'XUN@J]LEVX.V<0+2!EB$[(4_O*M=V( AL7(*P8[;B2^-JTT'^$=
PBS*K2@"AS^>AD"HOLU#T5(H'BC>[DI*1_-BE'\'1**LI,MWP>?=))\A*#[--F_71
PI4LM(=],:,V*;$:=]%/4S%4$XY=;&%[6\ K\4\M&6 L701I9$R![[K)]OK/3\0JW
P1CL&(5.*SYZ7GP9"(I/) V$"0!7R]BJ3/MK)X!$R G/=B8)I4R3U7^.''R:CG5N?
PB]/O^G$R$ (9.38VD8M+MR[]Z$6?N<Y^$W"/V@3IU#_=$NH@9@OH;=1$#\0<WED;
PJC]5<VF,'4/DWIHL))00H@%#-U(KKV"V6<EL/L>]<O;1VU%!V-YEA5?0QIT4]/+=
P3OSY+<+'HDZ/1-KWI,!^]8V'ZS(&6/YR_-&_C]#7PRB571M<2M4M4*$@_89=:R/<
PAOA+\1:IA_7GN9UFYJ%;7!Y8Y%QG!=C'ND9G/:/_++?;P-'7<8LQG0F8$-^R2#)>
P4YE$]VN:;D,SC"DG!5>5/HIV#/%2MA)CD@621-15"P8E_QMGUP!3,M%.**U$'8:2
PW[-PRU> .[LS9U#,\*@XN<(%W%YF44H+$8_)#-OMQ.FX=!?C-?772](W?[B++[CK
PM\4M&]>65LG57T?LR_:%!EF@[R+0%+"HS"^&>PQ.-==G,>+5GJQ&L;@T5.=5%)S0
P?IBU6XO'CX$).D0_B)I:D!X+$#!")J-P@BVNW?9A+WU=LQ_9[U,I-O#8VWGBUI@"
P+</S1#@RBQ/&""L0#HH9?]0H4"ZG6-COY#2+=/,/R[6W'%.&UF2-1T(CE[6;4D;Q
PE>IL)YAJ\$PDE$>)'L],L7P.EL UZ3C#8HN? !FX6XQ2HHG6V#;,T.ZXW#(LLSE!
PIMG,=A&FC-#:Q)^L%=T$?O'A(\C95:X=N\(FQ&S$78H1T^T%779R*=7GRSKT6S"'
PK2N_:U]Z_^$88L6UK_*'A?WZB_']0H%1J\U>(3$@ VK(L.3N[8"]-X*R6#YK\D#<
P<ZO2T#2?"2.FF*]Q*G^Z0'MCIM!&@._TH< BQ%5-#W>4\O7B[>4;/Q_>U&UL>HS_
P'6W#A3_O!I <5)HO)D$H)0B'B,W7K(I8 "W5H%&.0G2X^-G!:MXT^0WK]FU'/*;'
P[Q:1%L+OXOL7_"7+OMH@7/>7NY;G9Q(KI4EVL;] @4>M;&I2&$&/3 9#Y:XVX'JI
P6.29_.KOL#-BFWC="<%8^N1?F3HTL(>=Z@7(\OPYT9RE<4E60(]:%E7C:W21AG!Z
PQVI\[E9OQZ@6W<I#O8F,+D>4!?SM ![X/CP^AX7H;$K]UE>!!X%GLM/<WXW(# AC
P<VG0 MK61>\_Z ;PBH04R- TC#/L: K8*MN%;"B1=,R/#&N.!R]M_A82M)\");F;
P+$^7EI*(3,*A3\!\ERU)\C/KI%=-;[F39H+ !%L:;=0W 62<.RYEU/O]N!8*9A53
PG9#.87PP>S*Z6E<]M@GS\1E_@%9R=R(#[2L ^5>&KG&FV3NREG8+*\MK_KE<CE&_
P&$ZPZAM^(DM*U::[!>20[3(#:]_]Y4,&S;>17 $ITHC9S*GYE&2D@J((*!8-=^OR
P?+)M"^(I'5W\4JX#0H7_PJ=D]3+XKK]_3B036+&B7"P-+0^)X.4'>AJ3__5T]F)!
PZ(#;PD8#CR.C"?4ZX]YQN(J*8+*P%AT+?ZAKJ-VM/O'\<'GX,ER9VYQ1&&,FE2;C
PSZD%D)B15R]OV[N$WF->'^%MRXP8O,<RB-?,F/YZZO53K0?I#RN<*F,Z ^JCQ)1<
PH,B8J<9.HFMDJY;C9:8R]X&,P"##*>9FC+&/IG;=EXZ;7OEM/NN'EE33L5:C.V#F
P#[:IXIX5YL>3:GE7]% '_LSI,YA>70;CE%=P/.="!Q9[B'*EHHA'WLL0#GINH>WP
P >%"L)+\H-QS.609AY)5NS'+^ Y]*=VHJSW0PW+K91JRCRU4/1H>UL]O5V,G;IA&
PY)HO4$!6@Z'I,/85"C.!3AS*4SG8^,JY,>%HJZ.0]ZHN!9I9S(4/!BOD+9B3U^&5
P435#V)U<-%A%]]+C^Z]A+P#Y;AWGQ/1;I\HG<Y?,^G)-#IN#C?!PU"P_.@:B[ 08
PP;IN!R(00F=*M&!BY"\$K^*]TI;^,,&0G9TV $+Y@[6CX[N#@+W=,($/3/*" O,J
PNEZ-J/ M: +<R.G?[8I@$0!T-^6)/QY%1E*K@?;TXG)=+#T#;_6;A][LEM:TGR9+
P,59;@^UE>8?)1/"7'5;/.*E=7>/ZXX'7+>O=,)]X;'@![HG(MYM;R/Y#9/%W:R0:
PQ,$%\Z;UYI!DVF;N=OX:%ICCOF572SQFKAR'*ZC.=?CF!XE<L96CW.<^0/P P<IR
PGIW&P @2-G2OT]LMKH]'1]&'J*&XJMQ9^8W^7%"*>]GR#VGX^TK L_PH.Z1L(95&
P4/6OB;'?<G:GCR_-1Y,C]V \)8F\P".=HD?H?9AW'C,K6RS0[LTYKT(0*!(DXU>5
PE'[1K8Y_JH87@#ALP9O 6Y+G]PN0[4HL/^E\'*"](1I>X[0UOJ/1%&/>77?<G>AT
P3C2XGZ#GZ]!'E5I1'K@ZDP$!.PM0(!5VR)O'H15O_*3*=\G!#3G?;*#)79,%)>WH
PWN+)&T/%M@S8!'\9SA@<?W7(CV!I$K:\H39W=BT7GYQ#;8LE]A+7&<OD1Y:ADIY<
PS_"L/O&WO6K8'(2:F7RTV:%TRY@-M1NJMT+$)*A10*Z!R!10(U]&SY#'_)D@(8UH
P74#ZLG5E%!%[[V$[Y]SZB>J%>*L5SE9OE%87DOP\(H2K4V!UQTW&RN@/D%7#AXU_
PON0A2%A'<'9_(1LR[>$^T *(!EMH/8>BYW"3E?IUI(E5)[R_GHE,E[!0V+/^E)$?
PEQC-K>S)C%;L(@BC@ICRT+53@L9$I^9Q-'6@33*1&F/<H!KWF<HY7XD:UTZ!OL5 
P/XY=/67;LVQ'.G5V4/\M\^G(],GF]0X?[(7_?4/)XP=MK^O$ )&<'9MH-!KEN%,/
P_"4V]KXY,_54/3G$F\V<VG>X<7+I;7%]R#/5'<^QU/:( *-NJ>XW>G?M$S4C0DE<
PT*8M]H?+?TD3>/Q/)^:'<M7M$I- 9%A)G U'D0Y9^1_'5=0:H:E?<\\P:Z3AAIAN
PN%-:ZH29T;*Y&\@(Y'[S),_&*%X_%K%B(OT$E^1+(Q.3N!)VNN0=PX]</4&PV*.&
PL-9S7Z_=Z-6@W<EUP_8R/IK>XM\VC&#^I(06+[EAY<@Q<=7D#/)_!F5?$N!B,0[(
P3N^.\G1M&\>-7IM?$>=2)8<J?2:HF Y2H/PFCM1TQ+%^+/ZV--$D&F;<!&,N7$>]
PUM$EX:B+"V*\/:PKM:>LZA@B#')I@&QE("*5465^$A VX-%^WL_;XRR0N/<2 \+.
P<\[+(QD/?<0+M(,D<ZVGG4<7?WWOZDFI\RRH<\RD)#5L1P'OUD[A8TJWZ@A;QC!S
PX[+EK(B'3S^64@?I=O-IR)"^) 2\,4C#/G;&0;6T>)WX!-GYNK(N ]]XKUVC&!J:
PU[#O4OY)>/I!/+^W$-8LJ#F7Q_UH<6VYAH4K>M>",6_K/FFE7+<"\"22G<109'/W
PG9BD:ZP3$LZB8^]8Z-<$(AAJJ7WVT+)S#ORE$SX\D?M .L>?WQ3Q&Z'$2U0./4";
P<WN?#24D3WL[D"55'X22=R]EXO.*B V.;:CR=S$3X89%PP4UH^D(\ D,03;;4O#7
PXL750^KX,*F^NF\C")JY9XC@06#>$:<B26& G=.I?J+*;KB<^14VC\EGV17U:;[5
P5:JZ>EKV6"^8I8U15&)6<%!V68$E@HL.D &!":S,SF/21B)H7G ["?$/$XG0+3)#
P^A2=8W N?^:)@(H$396SA!*+2;1$?]%^BJ?,2VL?6@?02>'ZE*FBAS!FKTN7IVGA
P &^V3=O_1W."XU[M7/6?H5$*:A%!Z_>ADPA<KUKY:TS][7CT)?.8#W0Y0N4(]"E+
P%'2R 2DYEB2'.X>NV/]H(U@ N!JW7W+D.H;2 3*:&&V@R.H13\[[I E)C4C-T5#N
P"8<Q1GO&();1."V)2V1@9-SM7/O?>U(K[86>!V-T^3QFZ(CTW'_V*Z*OZCGU15PJ
P1@5IJIB/#-Z+U.1C?W@3KMQM?S0</MTT#95L-(Z]PIW:8-SGZ14AJ?@]/&>6)X%0
PW_6N98CQGYYRB9("2*R@,>8H07Q9]0UE ![ZD=4!<A:KY@@@1EW:X55^W]S-.ZO)
PO,YH,T7+$P=KM;WM=MXV@0.1/Y24H307#P]0)US*F6N@NH.&1T+PQA',!M@E6^73
PWKZR6U8:P^TS>4]HHCL$Z(X07"2"+^&?-<E-8P[X>=:K#YZ?\',5L(MR3[;U=J.1
P5UL4/9 2T+E^I"_<$\$E1:2[LF[ XVO*9TKB!640B/A];C=F&@BD>ET.J10%K:I6
P3_%@-_'Z=S '#"><.)O<P,A;//B(6YI=BFH366* W*@+OD4*VVC<IO:XYD_\M"P0
P#CK( H0V:(F-XF 65=_"?-JORZ>MW\R2.Q6L!YV@4>>X?/-#3Q)P196Y,AZS)*>L
P*ZPTB:TS8:REUS4Y54E> &9\[=K_!;X0[VJ26T_'WS@C)'YX"VEU@#H@*/:?<O,!
PJ!#H66+\YL"?I $-?:O!?P2&6^2Q,C5P@M8 5"-"<D_Q;2TJ2_;WJ01?!?(L^4WV
P2NT/5=YT-/[<<C/E!J\ S'[B9G]"M_=S(=ICI^W95;_%0R!/%*Z4T]*T%^IWEH_M
PAW_SDF*07>FS)GY]RRUQ2KN09>0*0//0)!.M[V"*^.1)A^B+ 'VK.,_0HN\/FCOQ
PA, .0T*K)@P45?C-AIV'D9+/8XZ3D92,!XKCM5U*9S@?;E(\,ANNM,YD?/BNL9#G
P7NU%OXP\'."7PPSQYO;)U;/#;/I(T":G$8H=0%MAO,Y8HJ6FE8. %K5_YQU%;7:F
POT<X_DA(#(JX8?>R[\*3!]'%-2!N#1AU78/DXPBH55?Y0;R4VLTU,?0IRP!RA4#1
PF%KQV.B58+2B2N@.)I9[SAWK8GO[\QB;\F1(.B=E/=%ATC^9<[$[R+\84-+N8>L2
PD ]M C:([B0NC5T<5A=31N9>E?W2R+,1T4!O62I-&B!GZ8=T2.>J#LK B@;\==M0
P%>^-99GOUB8IX.U6SG9MPEQ>Y>.0W150Y*L?BK]3G,!?VC63K(R6S-DS#)\H!O6C
P%9>H,GI::$?85AN<M)1D@X(7 5//YG;9,UG/1.OK%NOJ3UJS7)1&-Z2+H1*4K=C 
PH:QV5FK9#;N+;[BP?EP;PFW=A0%ST4:Z7\4,^;_C#;4XC#A#34\T3B2#(CG )?V5
P;3=!"$]GH0M)38>OZ^H&(&=& $&4D:X6SG/45<]CT=S&-AH8S;L9H*WU8]TAX0&A
P<MFG\3Q"@16T&NF*)'=OSK,KG;#V(371!0$!]5S:$<S_ZD4P_4M"ND0?YH_*[2QA
P^)]-3 )F^B:U]-WNR\CY343"2A@>DU@K,VS7- 'F-$D24,KM)O,9TB_!XM3-S 00
P_^X8K,#-C"7[;7ZY*X>V+< X<=HS;EWP,^Q2N";0?3JN7L+WODBN !B7GE+Q<4S1
P/^'Y-L0F.D(UJON!; T.B3F.L[*6P/FDD14YRCU@@ZH1H-_,$$,J%+OX("QG,-7$
P1AYL' 6Y:[*T&:;ZPLM/&7[Z9?74ZX%XQFUJWQ!U>MSA6\HW!>VM- -D>UMW9=V&
P%VO5%/H'M(HZTN/OJGOS>%<LJQ- M+_\+,<5,X;<+S3@!]PD6B29\HFL'(4^;0_E
PSFF)6MJ2Q*K>13%E.)73F-W _>UF$ZT*INI<J5#1 4KIH3_8\)/+5B/W0.<.0810
PT:U^XA4&9[0/].&,P=1>H4MB*5YIT &#Z=Q_F^<WU#[*P\,OXNQDS8CX*B%KQR[*
P RHT@((*_15O")-[L\Y.,YX\#@7(Z$8O3FDH#5F$])P2J164JK[#]AV=H_<13W;Y
PN=G(JX*=_M(NI:(\.75:51&^]@*D6RX$A8BXR')UWT?.-0:/0YRG;)8B_(#0"F7^
PL)4'7K\V*@*LBRU%94"N]J) A=(R5O=X'QWF*;/E)KROSS)DF/93T%:AO==2JEYJ
P[)UNVH2$)OLQDSBYVB1^;J"^1H4WD$TNZ<&ZR2@V.F[H)NK ^Z+Z6(C'M'R,$6?A
PE(N-4+O.+P4]%;R'L;YLKHW7CGZO=4VJ5T3 Q<T?-NQ?H#5>Q&EF1)1@N@QEN&)6
PGK6;[!@BDGCAQQH D8WKS]<6)SL27JT"<7OJ70S^S8I!Y<P,Y1UQ]NE)FN =+ 7Y
P@$T7Y#)@CA94SKO/+*:]X>@5:Y>23XOAR'D!BD6%M+-,"AV-[TZ*/9/M(%S9K+EC
P_B)!>DEEH1I13.[ECK&,422<]($P3:%;@\BRWFK0Z^%[4F]_OOAASVKA35'"N1(-
P0ZU,Q8=NCK?J;V@0V=GF2#!W37OW>TO@3@^[C"NX3D*Y?K5)A;>V#7&WU,SJF;!3
P1L",+O7PLQK30(V5LY 4H^UL,+53ZA,Q4!,-\SO68-9*Y+]G*.?#[N[_;O1 BS''
P,U7:L DM EO28:N,R"97G.ZU75S#SB=:5;R:!A$-]N#]2EL.].7>NWS7M= XX27%
PF.#FUKFPHPHE9T$$!^6<TF<-85' ?=@1\Z/P8!5F$6A$,!\?Z%LHL7-9$UD5ATU4
PG<=R).;:&RNR'H9%;Y(M@VRZIMA(H!^(1@X>T^.<Y134E(ED]+FUT4[GDZ8Z69OS
PQ6H]M9FLU>!'(NEK+6?UW>,\4QT_C+W'Y0]=%QXVO#)+\3'4MI?+88-]Q'U&[_XJ
PLHW *Z3S,D9+VY3-BA5/*/(T@W@6&9>=S9H5#%-_5B!#-#AXV'64W'FDT*/LS@@9
PVMF/S>Y$G+.7X\(3/DK(OLLN(M=CLV)AU% ':ZQ#$%%EP+#5'K@1NBR)7I!@W5QN
PGY!=3B5F(2X\U:"  ^(2>J-YBCAW9C]7+[2J!^E+5AV*$7Y@AW0;@0U16*AJ,G8R
POB!UG?,[&EXU,H[JO*Y4CZ5PF&U'Y8M&@USTX0 (MYUO2R1[+?4_ESGF#HXTST*'
PEH^]732P>S["KZ(H@D$FW890628M0%QXP@&Y!N/G[F:M?*3FD";\@!="X9H08]E 
P:9O2TF2P^V_SN;! MO5=RRZFL1,<9=VDAYL@:IL-Q<<4U>M1DVZ^(GP>@'/_S*_>
P#[QZP/@X&=H)PDVI@%_/^)"$H%U9*5/!J4(L+0]"!R=GWC)]KJF3*-Z$2JQARL2$
PZ )118G=HW?*1_@+*-)&.X54+O?\[X'E)!4E;D[)9!;ZZ2)[)UK<M".'^=.Z?9'M
PT #Y*^GG= _?P?F@53O^E/5T>_*T,\=G'TS\ZJWK%>+()'R$UO+IX"*V442I8C E
PQI#D(#J*SSV]78H@5]^UYO@*E9RM+$/ XMS$[D (QX H+[B'$SE0G^ :':"9ZYL"
P154'S>S>\_W._'58GLR[A)F24F_ >^/H>O;()!]2H:'"J<$Z_ [35X\TLZ0'8 3U
P+-,YBSM8J@N-?8/UC[WWFI/R8GXC 3+0.T$163F]X4X)UZ,0P)N$BJ3Z?%H@4_=8
PD73$#B&2I0%XN85/MI&[A,;+PCN*#(=S-*D"/:?;(<XU/&Q7 \+XD-[\GG3PH#?F
P$KI-JKA?7@WDX>_4RE9-FO7?>N#1^@8$>:T#<$DLEE7G3H[./0\-VF-%4=*':Y$ 
PF1>0*M?GOJL_!<^,F?[&?DP<*1=ZO_-N,J\SC-++7)5@9D*V>%KHP=<S"9""-/.P
P>5XA%_3 &D;)*G0?ED1 V^8MO)(F,68%K26RS^1+UF&U^Q#78R?AZZ%_LH, S-:4
P+MQ%D78(_WRUK8PE-=H8!5_B,WVHQQJVB)0/19K3'GM05@+_!+VL^>FV7N''59AB
P9AP]IX9$Z[YK9BIGYH#62"I H9_YY73?H<!DZ:V5/&"GH"Z 5>0F+NMI[+T TJW]
PQBTWI'D!=L%D&^9PYSG7WCZL*V?* 1R!!J#O$3;*IP-#5MK1#$KC:+];"4J0R+=9
P]7*=Q,,+88=NGI&)\R6;&/P6;J^$\/8GM686&43C$@)FOT]4;O#Y^[CSQ2V6SJ#^
P<'F2D@*Y!7C_])J5-)#!6V%!>ZG+"O_2'&"T?BGV91]/?.OC=((!^!R7TBG.UAO0
P@+-D\KX3;LF-5K;<WY[>5M4F@H;X]->Q CF9L4L&716D9X#Q_G*]!-B;"_ O.\\0
P!7$I:(L,UXA-Z-/+ROHK%Y94X$UDKM3<ID"63<(*#\=TQ,I3CES4!PR6G.W8$N("
P5N/L/"'G5X!9]'T\L;YU'!D,?V5#JQE?9%Q<)D@$.L!K)HL7%+&"K *0JQ8F,_4:
PV/N9T7A*-;+G^QH>F2[ZG"FE'[F&M<=5WJ8.0H!FS#G^%Z"'+(CR&^'YFM9KG9[3
P)':$7Y5F2XP>30GC\PZ8G;3 .<N'/% =5A6WZU,)!<@D;."%UG%_'A_,'_4GF'$S
P(ZT[!JNG\94CGWCGR#JAI"^'<-V5%[B,7&/P5_<%6PQQEBV79G[+8/AU+KTC<*?\
P!8]Q#++X 4BPL4G0$II]1JV)7<>)EVW"FV%A/S<:G;-KA@7^H%6-_M,Z/:GU#\5.
P@>=EW\K,'29I^)LPZC-S6'J )US[_KCG^G8<0ZZ'S)[=__P^'>Q56]=QE BN7RYI
P(%M]:<H,M/5@^D1$SERYAG^+%#U>@A7;U-*^YDKL)C0K4=U5:6(*-G:+_0+PBN*#
P2R!Q2QN9U;AD5)]:4>#U!:S*TJ_D#K]4),2J&>2F6.^JBS,MUR##,0N?E#!C*I?#
PSGU0NE@GS8=[]LE#;FYTV_/@0DZ]8!SZAH7I=&M7UI\-4(%-;:$]?4KSR2+V\V>7
P72G$3>**?89(X$1/TL<%M$]"4(5EFSIL)G[FPE''"1*"E;MZ/L:>COJV\%@6?&?%
P^;TYEEJCUZ5>-RPD/" *L4%V*(LT KG_Y'.D,#4 :HE9I #1L&N^]PUM7_].-&%F
PH^-W7(\>VG4TE3/(SHWLWDY^[4A@M&U,AL"^WD(1+6D1.7?+<L4&B?7')W#038PK
P?A<'3/*J@CF/0U"=M]GI5O/9Q0\>7?/GWIK&.E;Y)$*Q9=NI$!1T;K!X(4H">&"V
P<HF7,R]=![A"J]G'<V^?ZLOIHD%CSLL]D\&]0!56%I"5F(L++14*,-&C-:!=IE8S
PQDF5@GFK/F@Z/ILL;.0!I\FCMT?$5GRA(E3.@KH$&*7Z#=A';^M7A3-F,;WQDG[E
P&4A7Z-00W)^HA* VX&5\:T!;RW@PDMR-36Q:29>B#!#_VP,0H%*##6+JR_-LNU%G
PD+=/AI?LE_N.<)[2&2F!O0"[?2XM/4\J_.PM\11C*94W Y.:LAX$O%S94@%9UOU4
P_D[Z+$ _\GL5$)1Y1\KEV2!;P#SH?SOAP8PEE*\!,*,S3Y$B]<2Q6!PHHJWT&36.
P!]!1'@@Z^I @0%=W*2^#N:%/:=<^$C&11&F[YBSZLK]]EJ 5]AUDG9KZN^@'/J5H
P59SHBZF.X9A<+NNY+\T-RZ<5V3-08A!:!E=XP=NXS8VDD"(L\K.'!BC'U&H*-G"W
PQ;5\+GS,8T""BFT"!?_L'ZM+ :6ZW\%SH!?"N_*UU1:S,=20@(DN7>PG1ED)F8((
PD(_8G:#^0HCS5Q9]/X7?8]E=8J:K_L.9\EI2.*M TGROYX :CFI<@QT"[$J\%T[\
P8A^T>7DC%,$I6C#=QD!)"#-SL [&7B\"6C!M$V31&LVXAC+']M9R)3,-4U*JQ8[7
P1MJO4K9#WD3)@\Y1B^/I)<OG=*.P0,Z9,SKI4B Q N2!JZ4F&"G&S&MI7Q?665 "
P$\\U9VB2$&:-9$OWM5R1;B];M?@JC]W7!?O&77?@7X[&8P]P@#NP-\.;+HM+&-_2
P_T24^;"81%'%KIX26+85B3:3!9+@%Z] %"'Q!W'LHCR\<O [6(HYOFAK!SR1<[P3
PE% VG3"ZF4XFQ $^$!^JPD$;/ #/XRH=-X5@1 *'O45H1W-(/(9OU,N@CGG8Q$EE
PQ2)ZJAAD"*<U)^TE(QC.=E;OU!MP-ON'S:Z4T&&CP7G9^+*H#"4NWO?W^*!9W0>:
P6<BL3R4.'$R<C*SQX$G="/A"+P=]?L0QH@+4[IB&^1Y=MK*$8AX]D"DP/5S?<SO]
P2CK9.Q%6,W]B._.2$RU)_8 #Z#BZ.,RTXI$J!ATPE,#IE=<+,LK_N9?^,K\0I5,0
PGO"!2S?&#[4\*[25=L7EP(6P+AQR"UI["@,HT]BR\@%JI =_OE]-TZ5+9.;)4R[M
P^UJ>*]U?UZGQ>]'F0!=O+N)0H8:TGN..#:KDJ0P7D^L]8 ?284E WWU!K0IB4VD:
PSRSW/Q6_;KJ8@]@,.E+KR!(O>_W4F(BL\2#-Y-"YV)';:;#@92B%EOE$>*SX2%I#
PACBY:BGHC$23$5_L>1OQTO;A/L]A@XFZV:L%B76Q:_R^!#RPUY#8,FW*A7E8E-N8
PQ4E[23H)4Q+N:W^L<P9$)0[WT9'H@$2]9M?2C[:$]+[%> KR)49W5HD8\6<9O6<,
P^;2?!<:X6]6)5G9M]J3TQ]+;$2N/?1I$%Q%=U83V@4SRK]<?&TJ_2LX"#AO]-8FC
PC%\[WE4+PWL.#Y2,P,)8]GC88>+@K6H@*1^#Y.M^ /6Y]U=^.;M]S5D4S:$=.56"
P'5L(??F[6, =?.N^40QFD/Q/!AED9P:3P0+ZQ";6DM"JZU%W\TY4QS6Q8)=.*(J=
P^(X',-_K 8[F'O+)0@*G]0I_S@5]?&</(1)G*BO<6)L^Q;\!EAX[.6(6JZD"HRU\
PVP5T*6Q7W:)H_OL52876R245$@[H>::P7;TJ8K:X99CE<!D< P?;3OZ$UU_^R##$
P*^E8>1=-<P+)1&V-[,Z4SV(IH+HG[; NM38P>&1+05S"S^[ST*_R,%TR-#F'X/1+
PLSF8FK2$I$XNA'?9M>,2BM=(;8Z?>,R(== ;J67%QA_#M8;1ONXY#BZHLQ1M\2H#
P"@QN&A$2P#4'PYFR9UC)^+K&&,B7$"C53W#ILU$K"GMPJN2X^&AJV/G\VT($-=OK
P&&QV+MO>J"WI.QUB-S7DQ9+N5\D3.C5K'!H+86ARH6OG'WS7ZPL>SCSM9C(;^ F7
P]W!F$:4?Y_@"-&U(S$--C JJ9@HV+MU>ZFI_:APVM:G"7_,ID*?+9#:$+J13#T>-
PU$>G88YP[XHLA_K>33*Q,."*R\FDM1R5IL&W<7:'_8$.1/2E:9]0=1A7ON!>K[M"
P/!?K+;OM;R$1'1]#]\(1W2WTOLIN[K_L/KBY>%GSTB70#)&B1Z&WF9:7909?@5N8
PN;&/2AK,[<N!B5KFN(S:]?_G&<R*H=532@M&O;M-.0/S#HH]]Z)-$:S8&]Y,]+(T
PPFU;%%(,;I(9@S3"?)D[766FW%3.F.*"O\7'0BPR X)7?U<S""IZDR:^3F"TZ%4#
PA[(LV*_#7E:$$HOBU51(J5ZGK19"Z_CU;UF/P-"0P%M:G7;T?LR8R\8"V%*-P'_ 
P.QF'CW\061D3#T(!>^QS\52*Y;L7<(HRM=:O%&<CB%7($\+J8Z 9,DYO_>))7R!"
PP;T[M[Q_?"B3GJ-&.VUE<@IPUT8?'YM+H87?$.M)B"7I(J\R0^)O"9;!&D0>W4"R
P9]L#=E!*RL6,N/>5S>G7$ZNK)P,@E24L";WLSA9JX?LF(%)E6@UE;/H,WL)*%-HS
P"J:6L]]A>>M4H"Y^&E>6HC/="B0>V>YM Q2#_M1:(8]@#2S.Z^!FQ$>_HJ<CL:O@
PH]DO31^X!F\<=B @^Q7<(9[JE>'B_0EG%BXJ/=(G6Y^=M4H!7*V^0YU=R^=:IM/G
P1I"<;9$![?9YVI6LI337H("@X2_X&4 A\@[L#FZ*.-  4&RL!TJ<)NY$R%S>#T2=
P>&ARR[=>H$4:K]S[JTXY['G,TDN7RFJ(^-R K&,15KF'B\!_I+% W;G-N_<V^!G!
P!K:IH'EBP[&R,OW-QJ9T$_2>BUAZ,ER#T\0C(X+*9@&.J8S1@B=O,G@H6AA1217V
PSYUZG\?T9O_<IE/8ZK#Q7/V$8WQ'.9\$YH1;B21OO1NDRZ?6U>3\2FHW]!1W*UW/
P/,6V8WV"=;:-55BN-?8KWDAS2\T-$;E^^=*S@^/.$=JP"A!ZJQ/M"[V7BFDWCC=Q
P_,]>3LV3?WSRHM1<PIZ6O]89K@B#'O,"YEG9WW]=K"94,&%[>-H[=0(;D$!?Q5T&
P,$M+W="RJY!-I^2/'".>HHAQ:"OYR5;E&WT\>8E^%UD"*_A(]U5SV<V4,!0_<Z\\
P%"7 35T/TGZ>GI^SWP"@JFWV8(P%,E-YRS>P&S.U:F<GD6W.JB0;2+KC5LA!5#.L
PT1M6JZP%T-[F=CKBN@<.//:).XX VVA%$'31';N5U[S^A.W+QR][ZW1GF3:66[KB
P)]L <(N",/*N?CIN!QPV836*UOBP%%B)#J9E[%:_12AH$(RP3&\C^^%YLKUQ/WWT
PT*/@^:7"J?P'Z>A1WD,$)DD9DGY&CAZ&O 'K7M<5N1_%1]&S#*U=R9ZX)S(GW<4K
P7_G*^9RV\++>&C&366UKL A5\VD1<+1;6J?L@KC#]Q>/*$BX ;I<2KEBJW*S,W0)
P9[8*@X9/J#02)9?F^":"?6 4=3MPOAAIZH,<M77D"S@^-WN][$C9,#E3< 0>(Z_)
PS1PTTC\SK-(/$!G:R-1!^?WQ.4-FB=W>^[XTSIBUXML;IKER?L@W.P5OJ)U<>V=N
PE]:-%3E=HP-V!DYVUP8LT-CFQ9>LW!"Z_'B)OO<</4FCKR4>%4 3M*&6GSL,*^,0
PB8E0NYG@ #5UA4W,,V\&";,C5X6GA+5!+ !#%Z]"[3U8V,+TWR2QZZ]Z4[KBJ><D
PN,T3Q%L;H$$48A-6'R,XPQ>"F^D*(_M4'>:*%\FZL>J2C7TDVRRF3-CW.\!L;<)I
P7-HM^?A3_G"E&M32UUR7 0EB^ RD,.IOKR!_;D>=3PSJ\+[@I^S2+XX^(_ J<KEI
PM$J#L U[@S-=3^FD8HTI"/+3&:[G@0_F7%;Y*52?G3M>,JHRJR#[*MJU;XZO\^6^
PIZK%<BPNS+6)"1KR:R?AFTT@E3 O;A?AQ#RB3M;B;8<&Y&8DB+!$GA*J^A,V=PVV
PE>MI8/%^XPW1_ETQI04N#4].;U=B$')CG]FBH#N RH<XW,Q#9@,K70CFR"A-4\K#
PSHX_S%@G4^[QT+&>J.LM";7)\4@N3] 84Y$LC)YJ7GK;6T#2<ACI:?DY>4<'EUL-
PIJ:DKYWAZ)!-3/8/+]_M6M6.7R^$7 50.O)SUF\.;TK3_)69S7=/B"L/\^G_*YFN
P8U:5I7+8%WC&D)DEN^A4 4(];L[5HU<B0<D$[G,HFB6=\,=:<8*[T!U0TZQ5TM&6
PCE-<(3L *4>]%-M0F'B5KI'9%^@'+ J1V>_>\@7Q")/R)W#=H^&DE3X=ANF0-$UP
PY^+/0C&],$V;;^;_FWG[J51M@C'0==7_6"1])712M=(G$$YIO^R<NVFW^JC07H '
PZGK_"O13JAC:PRP I%_BS!\339D.Z9]9_O9>L%(@/QX74VC=)#P0QGYOB*Y8QIN%
P/HX-BUGB46"\PQT" [85I5?OFP8-: $DI.NTO(DG3#.K.BW=#*KN EY:"5L04/NE
PNBX8&4U'9Q:/!$2:M7KGO,G?0Q&[ARZL:RLA< M8EQ,,DC:I)BPK\G*P0TN4.#H*
P>S,E^HF>>NU1OT_EU.]$-Q,1JH.?\ VPD.#065_@Q&]/F*3OZ#X?>N[:$P/3N 0B
P/&N0-UA9'.!;X3/&U7GU;\U+G\1ZT!^X@EU6V!,(57T[ZUM3$(Z^?^1U#$*\]?NF
PR*PG:Q(J=_-M%AP_, JDCW.WN+FKR_*E5+/3KY)PE&\I%:;7PF.>U9 J >GM<BG;
P\%E[#%*Z3^1&8P2/7/)Z(.CUQ):O3'LOFYS 6M[A/^7J$:,=/1AY3H*4"JAS1@.%
P$J+/V81]/!?;'??6PKJ1+0,X9&IC'/GOR(Q8( "?[??\Q]+(J@+J\A]D.\I.Y#)S
P/5R1UUL2HBW80\Z*N FNZR0OWGSII.M[P+->@!>M>-_&8[B;748Z4FHKB)2;:TT!
PL#PYTK<^MT:HQ#6%/D,%).(&%.>#/-!HCY==G<&>30WZ%:I-[7EC$93?18^(*\AO
P[#HV)"Y3OD ZS<)>^/(TTO=E9?;(:2?D,C&0KHYB=[JQ.N.&J_GSIJZW\]'OQ"5Y
P*A>LOXX27U0=W<)IZRIPIT4PE_O)!I<)2#-CI2U"@B<.4*]_33\5S42KY8'.E:V&
PE?J07W2;LB^O.4 "-@J?MZ;/\=%[_C!%:]AZK\PAO) RS%F51;WJ79FN8M&0" RJ
P?SX;P'B-/*U<E='0.'O8JB-X_%G*8]QH7'V$ D77=370K/A\\/\BL.%*^O1&K6!!
PZR)_Y%8F8+8?.P9N^\I*W?(W&>=-:Q6*]80YMTV$U ,;C'XGA];EIO)'*E8,51*1
PH1#'M*68TZ1P84/[>Y18%CD_C_R:($/M-W9_EX>DBZFOUGVHFB<W(5*X$8#]@+N+
PW\?8PE#.S1RM$>[#9LV'# Q"I7+\_)Y2,:/^;94>==R'B$WPHO^R(Y(:.7R:JC*T
P7']-B4M6+0\8;6_M.28W=_$Z.FY!L):0 "VU5.UY)9:,!*0O1ZB$YRJ'X!7%D]2(
PNHTIP-PE :ZZBA;?G,8.84M+ F7WP8/0,Y,WE6)K)RBA%=XVA[W\$\*LIY\T%&[T
PQZZWW?,-H)F &92,,R'_7)%10U825AG+[+-.<?C5ST+C7X0?/?F%CMP)T?1->_G.
P-!6[$37DQ]2#F,-W+%P+BA>"VH,)M,/&.I(8B9J2TJ2@Y_1M0WDWGNB7\?>'I[ O
P?/.&Y/Y?:3)J7:\+7W2^DUU#2E'A_G#+7O+)7E>K#:8Z>!-W=)*M*!AIY)N^D^ R
P?K4/C[6_GS=)E&BQYDC3* :N7JN;D_-G]WMULLJQGWK+L4AWF,N$+UP:KJ<88]TA
P?(\**P5P(?GH-6FM2)[[5IV^979-(;^F5NK?7A\=YNL1$-NH-"$9#%K", P@HX5J
P+91?F0GO."1&>VT!=SUNU=#%7?>7NM-CX=5YI+T6.]6<,@/][9^V:;L;CN,SF^%>
P2,]E9.0(BTK#]LQF;H0W=1(P@9$]Y2%-(N<G4_T;BLY>4@6%U*/X,L[@AKK;.^47
P(W7^*X9IA6-)(MITA3^!UTM+C+O5UH' K-QZ@'L[L1?/;N+]=ID!ZR.;KMW,\, N
PL15HN<?Q'R^B5ZW"$\9^'#QCTH]"RH96$K&EGZ$;.&$E)[!FT:X4/718[Z;>BBJ'
P1"\;=.H7OR$Y/G$0PKE;E=4&P(OTQ]2OW1)=7F2C'5;$('ARBPF=$Z7Q'6\"UMJ:
P#UD?J=E0A"6KTDT_MV?,W/S(D07+ZUR6:3)#+>+-6N>T96NO/<W'Y.F;;EK,FF?4
P?P89S?DQH-K8OG-*_+>YB"6C,52_:4(R((?(\&A!+W'04B)5NI6=0P>BP6:W^(^+
P+PS>G]*N:S6Q/8NPOC;N'^[SOIJB06U.U#\<Q[/R\'!B?;T]1",)(( 9UUOP0S\F
P_[G&_6W6V7>E6)W@B52HH%TV3J%QQT>$G"'X$HZ]T]UYL#=/AP/^*AVE(2*U]*6<
P_I'G,C8Q[\TLD/@:_3N&E[4"MUNX8D69$$V,13JL!=]:.0FA&$R';N_Z5@;[84RX
PM_S(F# ;?&]J8C*5?% \+5DCYBD!(VJ7Y4,L7E3HSD,Z7"W\,*^'=97N1Q$)1-C1
P[9F<.0Y,>A'$2^:H%1>5I4&)T[HR]/DBG'KBEI.[A3U8-\Y1C0'H+V[EU<CT/GKW
P1'6$U]^^EU^#!YGH:"0@$IR(M++843J0)YZF#_,2-S7D:R9FM!2&SZ2SE^]?D^LP
P*NKC&NGUV+ML2W=*AYS]1<^LX2K):*EA9?M2#F3[4.4OBOHP%0->!R$\#)/!>AVV
P!7J3^QGO6I6B_Z]Z>Q3YQA<Z[V$#[Z8^_=8T]4/5MNPXP ]F,*YW#R.^Y"J_)>].
P69GLOWG2S8]M?_GKT,ZOSS.(DQKVL0(GXFLQ]>+,IA4CVCS78 #]I)XX5>LRV;:Z
P;YG$T-8><AUL&!:W<-![V*W_-)_)$=)+I_W4P\L[_HK:!QX#K?.949M5?]W3YBH!
P*.+.)1F+:<:_ -S5IZ2KPJ</(?2A7A=5LV,5V SVZ_!VL?!CXYT+B7FW!/A>_PFH
P2HH.*'$6]321]]\),5KLM)RP.F. @"NUQP^6;_/*WT8UN^)T/_YM%PU8=C.)$,J4
P.@Q 8?:K&!<[FI<"5/D5B=1^ZB<M:J40T]@A ^A@#8U!TY[V+>Q5-!5G(EF6X3];
PH!CA(.S(;C'=R>#^#,N?M"(Y!-DTH3ANUS$MF9H1JIBWM$ _CNV2MBQ;?-/O]H$#
P8K@C?U1)ZWDH)I.IC4O-[!,@4 OU((YJ0;@J![0Y5,^[OT?:PBO,!B$=Q;*6[\PM
PO1KTN)$'Z!K][OS3^=;8N2G*,W-9%CBB@!F'%L"JA1CON=-<-BV"OGTM&RRY,HN5
P>H<Z$XV-U#G+]TDJF*9.VOX"0G6A]_E2T2Q1%NR47,#ZLM^G9>=]G2E=8GH*]967
PISWWJTVV_U"MQ0Y6,'+LS%GV3(EFNR-82=(B:L\0*QB?=&4HH,9%>O56*F^YIPCX
P(H%X_ N>U0BD8<VB>S:'5,U&0K;!P'_+[Z/*9_XUA_5('FFWLUK//6Y7I^<U10I$
P(E\@CVXT/L88\6+0NE>Q' 9P-^=!4K,6D;%ZB44NKLQ?4'O _VF*96!I8@G@UZ"T
P]R0GOW6><:^),P]'$!,0X>EG'GK,[E4+(FP.!V7)V.8W]DT0TLOT0_OT7[:^N_8.
PS%_2+9<8-QPK19BC&R":4MJO]Z!R+@RB_+?1H16@_>TXNI_:_M"/Z]3$-Z1%COS%
P4"RF]/TE\FN1E^,K_W>0W)=1!"<#3):N8-Z/XV/F5[I=QSA=@R56PH>/@$!C4]V,
PMMI4WMWAD!_7"\H#I]\>@, 1=H%\Z5](50;R:B5;OBWTE@P1I=XP>CP)MH"UES89
P+# +JQL9LF%0C</;HV@%N5J:Z.\D9R<@3=C0-EBC,S4BUXXWF"X H9\)9/G+!F&#
PEH*%]]^"/??5PZB.VQ(4ZQ&C>$/H?L+&;48H\LAV"QR. 5'NPK,LZS5;[2=BL$H7
P^8MVI:)?]/6(K27^C^O9F(+/!(F#RK/EVM!O7Y'&H3?XNVUWYT.0@Q=/6XS@S83I
PF"C3QVDGR^8+''#4'F;.P<_KVW.#/S6%*(E62_71>-H""L'XMD=)$(/_@73Z9MYF
P6O+C1R 08]RI1OET;3FD2,QH#MK*'TG0.ZJW;;]2Q:3,H<>Q51]+4"PFRZ;VQ/;X
P*2"W7/9K%$J45N[9^0%J8OJHH=J6K+/,/4*V?PO]#Q,\P-I!7I[E<AE2/VE:7YM:
P1MZ)@:M+^P]MR-17H]^ [I*IG[3@@P'J<#;KQ)::+'@NC'-L JO'8-_L@P23*U^E
PP)"8.%.0.X&RW/%0=/, 9T&Y(P]9&/X@ORHI'OY>O)BPM'(R9)./N%I#4JHC.=J<
P'=."__RF66?[<HU-#'U8K8 =S8NTL?58JY^0HO7X?:7F1C<P\0PX4I%"$!\T5VQ,
PRVMMO(JQ*7W;E]I67?3([W8O@V<67AP*Y72<Z5IK[FHV>M)NA>^5\."60.:C2!K5
PB$G$8L!8T!J+SQC<TEI#XE9_F4=GZ+G9=0(!RIU=+3 &D24_E! 9]AEBVA-T2&=[
P\W-EW0 [RNGUN]4"<10;H^KS[^U3D[Y+?,-".#EI9U_ "U'L1S8X<ES^ U5<'BKO
PS'V#-+9.ZSU*@^$@O3!KD?#Y!5[9T96XS:W\B&A=#KAGY@'@X\6\.JEM39\2;\7B
P8*J!T&8Z_Q^=,[E2E.K#\#CC6"O0FY>D488JU7.Z)N;$MOGM!2!UF]][AVY7;! Q
P.;Q=P/[[9W3%=[2:)GHR&-@M7TQG.\P?+$MJRQ$/4W8^D$5B18Q$8AU_;*T"B>FL
PYE[;___*.&5,?_96H6=//C;<T^4!#=\JIL<P,@/APULZ3&A$>%J1,FN_+\.$!^&W
P>3:_8GD' %!?GG]M 32N8,8OUO*93^-/D8Z1CX0DG/VIER'<XZTQUEE@D#C\J+8.
PV1R:"? *E>:Q\I8"=T]L7PW2"9<6Y9"R53<)V#':GLN]0(=>82V8JH51.I2FZ2E<
P7*3N7CVP2QC!4E"GDK.3RRY+\;L[6>5>?R=B]IP41_<P0RQ';05A38.>*DO7R&2<
PDB1#UBJCL>PU.PZ3"QYO\@&1IA[P 'ZN9EX0$T\ !G_#2;^/1"A(&>>5A>N-.C+T
P<9UB=RBG,A&.].,I:#?F%347%*) ;2;H^R39,5>V!>E."['PU$VFVN#G&2;$O\H5
P+*&_5,0I38:S3[19VN!NXTA*CU-K"+B;UD"$C#@2,Y:=H,CO)?TDU/F0EB<S+C%B
P;;*B]E'L68]\?_W.07PC[2*-.QPZ4&KAY1^?5> +$SH.$V<65!I@?R9'1N *("W6
PS'=(6T6R4!:9/2ZX)FS;7#O-A7?"43\@X*=*;RM&"WCJ :$.+SMTQ[?IFU^'0:\#
P\+SW:E^L8O7W)24IFA2GHC]D%#(K%N_,X!M_L,AG8J,.$[X&F^AQ+BD:ABJ#S-Q^
P3,*I6FEI2_)-,^I]U0C[07,8#3A@01!K8+8@WIR0KM0KP \PMS#,Y8Q?R+ P1MYF
PX3OP6C*)G9'I'B[(0JZ.]*SI+^7RIP.!]XPHO%_*P&E8\]+)W64XF 0WS3R8<A^,
P@]K>%P74<^_>PGPL*K!1@>0.WHE4NS 5Z8KR^EE8?;TD[0.,E%?6%?&<-Z5W :)"
P1'9!BD&!D51_SX1XG"EQE5/4K'=YA:A<@.NV^J:@=:6%3R%:I<\YPCJW9IR]'>."
PWFI&H.]2\)<Y@6+;K(_7&:JI@BO6=9Y3E3*S_PF5X*.06+2M?8^#1K#22%#<=3S#
P-YY-(S= \2Z6"'(9^(H0VUU20FQNB-!"M;EEYH8'7J&+J443!'*A($S28(K/;I]9
PS<"KN)-Y\^.MH@5P?.'1P/G/LN"Q/7C(@3'/_,*GHCT+CJW_;B='+=RF3PL3DTMB
P0,+["Z,(/?*K=?.-&>5]L8J^G)R7A/M G(DV0<Q6]YD]47^2^&C1&(,A])(#(<BL
PX ?F=4!)X[ 2\:^D3GQ2A28#'XUIZWP76SO1\QI_C:=XK Z#@>6>F9F[>E_IRTD%
PRMW3]OG*0<KK4!@]XVO#2INQ.YDRC.*ZSI072)O*57N5_W]84(3<!D5?K&+/4QK*
P\JBF<_05'0\#MYD-N806W/FQ[.2'A=R9A^6''Q_3U,[; *" 1O38D"9OLU"):$YH
P&S\BRUK%=IL&<*;B[U/7@HMMS1F18QUO#*U)%IK'VRY70\FJXI?D( /U-6>)N!_W
PRO]NAVY)&3=\>EDIA&Q@Y&>E;^- [?.W^_+=?JB"79YCMT=]X_T/,_@LY\94QKSL
P+VX%"",==5]1V,>TU$@[PHI8'F<2>+3U5QZZ[?E^W2W%1-(K^\3HRMZ^N&WBUHNK
P&B_](@RG4[9-#*%J,>,:5OF@QAQ]L/.@MZ\S82QS,]^$X?=8(A>6_3-5/BZCDN2(
P=EW8>Z;LW7/A?H"^]!%IGL +V51"A^-#2E!!4R:ZVQ_#5%,:LT'2A/*6Q^ =D,H"
PR_C'BE8L7P!M!2NTZ/XO"@5(>%&.34DC^3QO:?I]Q4\;[?@G$:*RT$107@5I?;2/
PGJ75E.W7&#5[]X3MK%P!Y VC;;4WV#5?CFC#D(JA)J;V;GNJU*&[H%HW#$^&W6ST
P\V>*TV>Q?#G+P%/$4:55/!]<=R &3&YY;AI- E*AC!:R398L'0C\:K45+?S4=*#O
P]*'_H)AX32)H.,(OX*3<VW@2=5>;'IB*'089>14P#R>=-,*%HC(0D5X289$,]]38
PU[0C%V%C4OW0&S'3??-KGN?)^YM]>35O[(/727QO4)BH(/0)S&_%VT&U3C4*C7E&
P0(;1M0ZWDY8MQ>6#!7T:E_!VL4C%"7F2KJ9 J"!4&@;;>FR2O7A<BVFOOQH0Q5]7
PL*Y53&MC%P[]#4F&\;$B$>-LE_K6?B]NW\ 6GNV_I"BI5_1B#)?UET%*VO[O3=!]
P-_W'ME>GVHI<*GZ8;I655FIXSPU[R&,=O-0-!:#DZ@\*BLKPSQ,:[*W1&B+G_]LC
P_>1@'OG/1G)&L^$B:!+',6LKC)\_RJ^V#Q[CH#!1B[I%YES<V0&YJ&/ZO*UC@]]5
PQM2>F05_80 (-R#^\<<DYU7C!"1R!/0:\<K\RO9]3]X+O:/0&!H14Y\M4A5'\>D"
P^;Z#%% F09N?!T7YCB/;_88&1MA8KO4\0%G*MY1EHJR7#),"7/()E9_WP3$D_?M*
P;VZVN:1:L:]07!P!8OTJ'Z(97-Z6K]*$$R-"+-4%03W'=<>XBHE>K9MM"\F<;DX4
P'L[3D@.,"7.]Z$A[]A83Y#E</77S$3Y3.Y0)#;P  *\@^6KAKZMBG9SGY*JORPRG
P@F6BH/'\'^BYK<.@JI$&3M06%^!-5N$+(: ;D49Z83[W.F$L#FXZ>S*L4OM,KK3I
P8*19@W3;R4*=CB5L]EG9&0]HL^0_F:?32_%$:N'.NL8U[>TU#0*W0L++CDVUN^I,
PV@B**#&<>[7D$=NLC# TA4_;B:JUQ7D=+BV*4UEEGP> =;0KO:M7<^3140F(G1.'
P0LLR!CU6NP _8".[U8FIZ;UG^HB:=<L*I.^UF]*;P!,IEZ1E/@!X2S2_!>,VN5LF
P"/ZL#OLR89#=$DK](8X,1](&:NJ\9E>)%"&=>@@GK=TBG>F[MH\4R;W).19WHYVL
P=57X%D5+I)!3^0.LR<B0&#>0KOB28J0M7! N?RZUL_O?WBB(3 KX-J+:@]5T7+J?
PT';6V5MY5Q]= I %V"^%K$ISRIX/L*K#_;NDDL1A !/=K-CP[%F39C7A/,1"'E]O
P?F/]1FJ[L3'*+O@&_]^J?FCN0<IX_%<ZGPB,E6#)H8G0)7"B]]-#23I.@+"FSX3X
PLA_)B3 :"Q.4:>EV8?9:+2 A=+=XY5U,<[T@?>K8 ?DYF@?>/Y3X-N4J/?1>2AG4
P?$MFT%8'Y>7+"O($=HJ&NJMXY[5J%]V^F]F4#(M\_U7DVY4V+38E<:UPY-J;Y;ZJ
PX5:J3&T=+4D^QQ)R$'7]KX?570"A\TS@YP\Y(/\VP70,V-RZNZQU,UW>8O=3:K'A
P7A[:\]BT(WFAB61O":?0X/U.^X,U'U#*UR3*U.NMA:T7*MXQYV.Z5:$8%LF$%;]Q
P(HMS1 32<KE 71!544 :L5>\:_]^;9-D'"% [K.NBC.;6X?1I0X-OA%Q]$8E! @/
P]/)-2R@P@]X!4^2,/'VR6>ZG86SBG#WA_ UIMV"(D"+;C>?N/^0<,D4-V].SMK >
P[<QP5]ZW21U+PL#YRX__V,<,=&*08Z%9F)P53;37T9JP!+^\+!ZGK"#B#SR/##9-
POUJQ[<K;W__(/N2G.';?_7:R 2?'C1<(XEQELER_3\BAWU=6,AD)=]Q@$,/CYG06
P.+D0E;!>3#$Q,R#T3&/DF[^(;BW3N75WCE.6:A5&4MC4@Z@H?163:?91H.F"Z9/+
PU%;%]))8&2%SO<=-(NFIA;8.A8_TB_=+!^@=2\.31_1\D.P>)0^")7T$'\2>KTP7
P,/UV)37%78+^_O_&*YU_K-^FD?TUK)QEN$1431BFX$=A7^0J.B]Q0D6N4Z*X*I=%
P:F-.9>V\:85 %^FU;9P 3^%2*0[:'3EE>1*!BF@()/2A(ZL5.,>2QVB*=VO03D# 
P-+]U/;(]*?8@"B>#FR%B!;\?CO0)%YN<-:"@W(ITA472L$D:WC]XBG0ZWUCOI)VC
P9#Z\D7%%"*UWP"T2'P0I)$._G@_*MYX@$@% !&)+BVO% K8<"$_%MWJ$B4,C*%6H
P)V%6!;\@HEE>XY\9/) ;TOF/?;LQ:8)[4YC5GI$-KG8-^;Y.T&;<[VYQMO%3E">]
PN9NGT@"X(VT;(7*KTDHRC![O.2:Z4V 1'BJ];^_]F SWR?OD.^O.7K2VT6ZTX/GN
P59M_NW'N?%FBBDM8S6\@NE%%$8R;9EUX/O]@@MLD!70%5 LB2D@X!T_"?RY<H-48
PE 7:N9)C+RW'4$&<6/HZC&=1?#6UL]F\>9I9/6Z(5DH^5 3W5B9^5=L-W^HGW$BL
PDN>%?.DB_N?;MF3WM*I#RV!6"UCU^LP+J;$@_+&:9)VA^7K:LF-H!N%(V]T _&76
P/BV*B V%0T*[UNCWJ8^<_,HGH12-I"4;8 TT3FA2F-<9U#QM/UE JRV7F5X%[;_Z
P)S%6Q6^O3.-:-W?T"*!<>9JYH,W:D+#:%_RZI4_H4,]+(8=';K%^E[@S%<!+^BLP
PI$:$@X'>L[<0/].ZS"GJARN72+^6V\2?,T?2_*8]%^UOG3]ZG*9-E<4'\$N0@Y> 
P&VIA&L(R;W%'BY7)+$A+&B=EUAWAK 77KP4=3K4X:0^>@$31E9MU^P_;GVX]E:[?
P$U-D$$K2(<Y3VT-LN\!&W:2Q&F)^,LJ+!:@CR#05J;^%AUHS:/V):)D13)J[I+_?
PI.Q"Z6.V8Z$$)<$?9VSPX"YN0MO5L?P*Q4NP_XWQW*4+-G[@ ;(TB],4MFC1^6-^
P@^T#/U\-+D^)EV=&V<32N< C:B_&FL)6602"=C/72%5YPVKKKBV><03E]+U<5+/;
P9J,=A'^0PFF]G?5I5>Y;B+V>,#212ATI%X!,.I%-O]B)TP^M[T.@J*P4H@AZ0'LE
PDR=9QD5K$4>&D$[0CB+&X'57P> F%!HV>M-]+9G9Y_DQ>U9W6N"9RA!;"?9^P\U'
PW%-/MGAI&07R#%/).QF"W1E [P4$F4W#1M+>E]A>@]RT),XH>A% ASAM:@BXC&QD
P316N+SO0+!:X&*7_S(2E/.*,,VLA;9M]<./"$! O!@+%=UNC)+ZW@NZK20#RQ\P,
PC :S _8E$C&@ 3&<Z5?E*=+2H;S[=25_8$<8Z^7K/7O&7B96J][!T:3_*8=#-\?"
PF<[P3_M.Z"R^%?^F\T<\T1MQ)W [2:J.V#G/(<<OBPP*U-3)4>9S I1AYRT>.+R7
P""4*V8F1;/U6X8PGL1NZT"0CHQQ0+'[+M2Z]NTHP#39-%*R>]I,(:%@M"3:&:,<N
PL)Q'7[9.7,X<XEN#!>0$;+ )C>N+[5DLC@RHH5V!'E/38OW@31^?8W,O/P!)=[1H
PR3W6@2'X"^7B,\PY5'*OU7J7^ND34&!&X=[;&,630F'SUTF:4W_/VKH;U\[ K@9L
PO#5B/6_7-W]WY=27Q5*G)19 5LLO?O]X5S57&,QKV;SP[)P['3%8:+YE;"7,P?"&
PJV@=*A@DMI*&7C!9>@G>;+7 AE&UR \YN/<'T&T<>P-5%RU=ES%U;DKU;ML17;%1
P)NFFVB Z8Z3H6!D&KO [32+@0M$BT?$"%R/SV,:;C[?FL]P'L57(60%"S.3]D5O4
P%)R2[9^T7&^/)JJ,L6O()[>=6K^4@2"Y"E[LYT0VW\2%&,!N;NC<0%E5#I3=4%;G
PN5G6B;HJ5J%10[A,A;C;ZJ7=4_^DQKX=[J@MIN?9'-L6'3_]H3$UH:'6X[R(7%8H
P)8#78C]"PO/&&ELMO#RV8NXLC_K&1\8PC^E=)2U&64_6&\R//@=Q56I&KN7(_'P*
P!;D^,D,78016^S^93^SN+UL:0.%P<\P!2JN1[*Z2-$MD&2I^W6E.*<>_%#$-O4S=
PV7/<1)KU-^.2@%.?.)NU*1,/ T>+O+V,OLPYNA=]*->(3]HWT^(8-O_:8 C/.;#V
P!:TZ^3Y^>L:G);.14@3.WE<D*]C^6/H;.;!)R6<!2G[[4IS =(#3#K#?FK4* (.&
P^R1R/E=08!)R3Q 4I>N'52.<.$=:(9JC=7/X^5QR6P#/Q6H5P)N'QJ *6^XY=KU@
PN&NM*6)TNZ=I:@L5UJ"JB[;#L3UWY2][\LT#^V6,"%R@N ]/[ABDC-PCZ8WJPS5O
P+EZY'%^]%+<\HR_]II=!$%)(N*B3SHB<6G#H6-;U\!GLVY52_N0V.OZ46<-_3;8Y
P2YP:@%RJ__*&!=6A*5LVM#9_6V"45F!M:S)$8I3OK">CQY*QW 77^4Z9+K9'0CN:
PL^V8C*AKZ@,?3[UB(^BN@W V6&K,,$#K&(9YYCG#!G2.%T0*YIM_X02P_!UZ<X,/
PRHHWL*WC>.QL/-;#SF#SD:-':_&QGRFO,#1=JZ*)F;F0YA7X%U\@P+^;^&2DE7B;
PF>H!/;)8@#' &V/83S RI>@'54WS*XPUVF-[0>VTC<#R -CNXU*!?7>,AFL$@]?*
PU3K ?.6ULS,PD;%N[.O(%&2RY+["'T20@;4D$ESV >(T?R_ =@'SO>9,FF!IQV\=
PM_5-PM9F6V%24^RL2NE1HD+&. 9N]Z*OZ++J"^6+:5EQ8YJL!ZV>5.UXU?%3XPLO
P.13(+  NM7-C$<;R$1'N4>@K5C6AKTN#1!^(" F4<ZEN? ;4GZXVN-)LAP:E5GUT
P.2%WG5[JE<@BB1\9I@=\ :KYB6&.[XMXB^SR1D3,EGW9A(CF.!Q7PJ%]Q]!CAR=Y
P-O\\BWCV"CGX+XZ7'H'P3;MA9"G)*?7B/U/I%AST['J/]O?=:),#]C\I-S%&^=[R
P:KO,HO=.@)R1=C@IQIM+H>3#$AD?(9-OX#JVV9D)81-0B*2$N3FK)G2[]NY,C( 0
P2IN5Z[L.D>N>TE\YR@8WZ! 1K1Y69(@(Z0I'DFIFI%!$[T]*RO5\"Z(A%S0@YR(W
P/6\9(.SG7H>8HIW!HN&_O;*(QNDI=S.NJKB?37?"=D@9LIZ547Z0[:O=K!;A:S)V
PQ7/CM!]JQU6A\]%]<(5&KUK"5"',OK*^T?VQ3 ;K6V$O4 .9N NA5VZI80_9S(:Z
PH3];B[ Z^O#NF,LL^V)<53A,X"KL==\8W!P#KQZ,25_D<+:/6&J^UYS2($?O*47S
P_$GTP1WKL=['BK&^G9)0>\7@DU -'T]8WZ2)8(EVA\]TT#0BTM@.2L#6J*<D*RDK
P7Q\2 )\9G3!>5+BP$JOFE6)/%%94V[DS@.F%OAR+CTE!WA?.\%IFLVNHN/ H;)S)
PD/3IGX$.1UVURZB-NW16E*_CA+-59M;V?:XC04R:)Y%S_)+$H2N.<']V*E/36FA5
PTS28AV'9G-)D!613(2 $J%\Y:!>>_C'@G%JM/P34S1(R=64N@L=4<L7XE56>(RY-
P.=3A(*L?PZT3T2V:78MW+H=Y4-+\OX;T=*K@0U"B=>FTP?7?^I9)4=E!8<T*0SGQ
P7FJS?5.<_/9"?94+P/EW;".RI^X2QTZ4 ]&5.@$\:[:VV9F-MJ'@:^=L(B\7.2DF
P^@3E2D$]D5CPI:W\-Z\+:*4-1SKZ8Y+.@M%LO\R*S'AC!29HQYR'C_L"_D6(,2#/
PJ\I@+\T& C[S_[9)79YG>]HY727^&T'+]DH(:2%1^;P?3);W6%.)=IW>5\NSDC\C
PT^A ?1%PO5QY3NW![V]GI:@X+#ZL0JC$@)&\D3/V'"@?/]&0^*\B7R+Z(0[!Z99?
PBU<"?1@7^NC]^RM.I^(<]1)(_2MW7Z*4D-'R12+748:VV+DI"'MU;I]M24WREH1 
PQ J[']?+S=N7<XD,2.B3WL54'UIQ7Q2_\Z66E5WDZF;Q,1'D8,:,_94YM]7"%IVF
P"L\KHB7-6G8YXWHU7(_*\JL]$M >,279N!0>2&!&2LE:7JD"^O*\R'PP53?7I.O.
P9&C+H=,VQ_8MWGIA*C.;6.].;\_G SW294##W]'#M-1[91#GK_P[WP>+8 ]0;QTX
P I9\UG]E:9FZ^"$&(#&JJY*8TBUCR947O;GF4&T?  F..&,R<UV%(]B?P4H%W>[$
P%@DJ=G@S.<[JY:U],79+#ELV9MH]\@V*89#TW;6(3M6A1LM[=+#D&;KLFVS2E". 
PLY;4!DCZ'(ZO@=?#W*&3&IE6-IU:"30,_>M&O[S<Z*!1VIO""F(G#$B]S?S)@..3
PMD\-,QQZ-I8I64=OIG*W!C_DK2R\.6J_3L.U<7_2A+9MQ&34L,7=)A',S&[(#:V#
PMU*F:_HCD7:AJR^H:4WKUTL?/EJ*OCC38.T2>K."7H63)$+G>[C#'.U?S%HO>N54
P$B)MS1[CZ] L!RF^LD@A=< UNYP$.$FMRBC':1Z+RQVF5P('?7',D:)+GYP0N<Z-
P_55:6I:'RYP^_-I[S#L>U0S6I822$<0T[%=8V(F]T09/0^;*)%!P6 U.#)F"V"FA
P/!\BW,Y7)(G/ZFPI+ZO"*A$!K[.C.H4LNW7]8-73#^FS[VPL$VU\?WH\#*!GDNI:
PA8;MSC5R"7X(D91XBLX:>+PA,^,=G1,DWE)*R\C!1O"0"\'H5Y3($>+-R-.:>S@C
P3_RU.+P)>[H3?7FV;J_Q*%\2-89%P;*IZT7.R"K>T.S[!BP3=5GZP(V UCW;6#WV
P[-*(EJE^*.3PP4@D(';BL)F)%C#\I.*EA>T4M5GZG0@ >B;-^9HM(@LVU%+-!PY?
PD9[Z)U3M]_!ITR &BP)(?62DAY>TR4R[<L:06%K3GUO8F%],:0T88.WH*]WUWGRA
PMH90DD=9GV)^I+L2A(5[3N:)KFB,L6F^KD*5[I\7L-,R]NSV1#^J!B+*F=YVPLR<
P:<L&!.6XGV":&Q^\H?A"K'F/5B-1F\;I/Y?P'&3?=@S)Y'63BU" )V-519UXZ'''
PMJ)@>!;25\@C-KBA+NPCRW5+FW$QC81IEQ'QPT.<\$B3%P8].(!^6*UX\Z;GY(#>
P7PLN#JA7 SW>5HI!KG*8>FV_Z\P1P88.%NG33-(^2$HH#[0[H?M$;S0$E0]00R1D
P_TJ!WCA_?RFU+%DATU0"#ZS'AAX&2J1U.H!A%R>E/=QUTZY'N^SPXH*WQTV;E>,]
PU'UTP-::>6\KP)! 0>W'7;!S"(-]I=A:R(.GZ\%FZ@9LQ]:\\VX+YH]<#Z:PQU?=
PDFQ2#P//QPCT;?S&/2[P8[N5(RXC<OVTCV5@&UW *B"'D=AJ#4OYWBYO62>=4L')
P[@D\4D$Z[46DORKU;RQ;]6HUJGY@C)YG>1R,H95USX61-77NCIGK<M?\V!JC<FDN
P5".K;5^XW"?_N!/$0XI/DHG9&7>4CGUU*1!E,0!F#K30<\6@K@F;KYSAA3:IFKJ1
P:3L(#N@7H2B^/DAH;TLRQ!G_ _2L,5<*QM]QUSLW&2@%M;VA'WTRDVDU1[;Z)N5+
P0M_"$T"U<FFZ29)"R3O4;I?QE(J 8M8Y+@/YEJ2:\X:9N0\5P!-[<CT&(-ZKD>PP
PJO63#6/VNGIO3Y1\OJ&1P5ZAG04N"#D-@R[R/$U8[[[EB")XT3HS5.,U[#V8_2\[
PJY&]#[*"SU0[)U $TY,B:&S[42"9.[HOO/[+ID(L?HK;+&41843'W D82K#J2-FD
P@0$FPS?R]'+"H?UF4>XB<^D?I6N#A^@;UNM/PZ9/>*W4+QEF$2,3T'6 /^P<%@!"
PW]@='@,KY5'VQ32ZQ*R1=ML8?;JMLA/&*LE[3FC$G%UVD\V8,H(GMS)>NR*DR56N
P /1G/[EN65Q!C=SRD!*OQ3$96E0,5,%OH=XLW1F"2T+K"@OZG^+C,RF1PA.DSJR!
PR0Z&NSX:%;OWVWX47>/,&!?S% 5'YL3?9[\G5YD(!,!\LF[B$GOR]Z8P#(AJ4;?W
P=V_8[KC)GAEP?TP-1K'18):3!S<:$.* RB8R?UURY>X/7;E#2U0G\+IBC&A5=*!W
PT,XPE\1KYW[I,MG#4_G'>$YBD5]>H%_N6CI20OOY::[0OO!5]XYWW,/3B=00WZDZ
PC&N602V:TSM$F^5'T^C7"QO9ILIJKVXKR["9&L\5**KH5E35_00?LBN;GLU-J*'J
PFD[H03O&T<IN,"ZG#AJ9AO( AQ><8K^_2KZ:, 2>MTDGN2*E"5 "^CK7?AWM#9?I
P"FBKY<@"]\+)\YZ9>IEUT 02!M*AHY]("Y33A*$@5BRO*HQP8B_VI4]?TN96<I#T
PIM8Q(6T>OX]E'QUM3PZ,Y@<,4XQRIA@,CJRJ6!<4<:9I*$H$?1NANL7>7S'FT7<Y
P BBZ]5J,H= [?TWV$&C[-[T3W[S2ID EW)8T/';/;K436G4RL^0Z&KV\'N2.?$,L
POO+VMC=CEG7S%Z7G\+&1%F5[+]],M7,]N>0_*%# =,^F)D>/G5=:T:B?*+I=F9&F
PA_&+1SU#2U[:K,S"4#H'MB$3>5TW8ZXFZU5O6*U>:NX+I#Z:7,A0[(T!V4& W'73
PF*:76.2B8?=-(=MP]M^FN0>7HZ4FTC"+JO(PX=TW#!"4Y5_?RG4%Q-9Z=I%P%;F;
P\S"H9?0U3BAT'AX#-H6$S!YK.3)^QN),LA.^QOZ2R)7DK>F2O)I6;P\?[/G2S_*1
P:I0X+23 87 0RQ;>?V3:T"]7_Z^4;I2:OSJ!UK/].]8Y%6*;?@ ^8'T/L]PO##-1
PSJ"-1B!KB8 /#]A-5-?[JQ4D3$EG5X^VFSG'W_D5 MBNF U6\5)*$JJ\[>H8N&.'
PC3_+G8@U$KTE[>]\'7ZB\^:Y7WBO+"AFQV/>$S=^ "4=CHT*LZ?03L/=> 8 47D+
PK]"']%B3"]D$+.*0HF8,%NJU'\GA=,OOO$U+&[+$Q(1T9W:--]ZO)L 7UCC\]XK3
P8SRH8QX*+FZ664F[4S&@KQWT<%N()!X%2L%6<P88_K?]0W*N!W\^GS(,_";>BMT0
PHK5@.)4P$M%<IIWS0Q1-/_&.?X^)!:;%J_4N*>K;GGA.NZP-^-A5PS&5B I6//]8
PAA@V92N"HN5ZQIW=?32W0N0\>!*@7=0A"CB;_WB%KN#*5RDG?X^FGL34)I#/N>*D
P$  ;P@[ELQ<40<XMY+9F]C&^Z8.-1IPRK<N48=)N<2(-\W[)?8CBE#7^'XC:O_,:
P8 X"1''XUUU>YY]U>!B-C$Q-H.\)1]@PKQ'A4,1=ADS<-$!+%5'1%Z0M5"_L)E8?
P:5>9XO,-Q"-#5WLO ^)UN-[)#3^C#@3JE8XU,(G .O>QGZS$E:E$JMG=%!WH,C@5
POB)+ZYL9+E2K;YTEY8 _11O4DYTKQ*G7L'=PD[-:J<B7-MG;66D>^<QGZY^BGBIB
PR4R(GCDIHX2&UYC.YV_9:T+OL06,=>$X9 W#9R>*],5=,>?,0#LF]2YG3KC5&GG%
P',-1ZG!M5.6L[K"1W*;3%\#(M\5@5I#.U5I*@[D]XB37NF->@V7D8W 6V31*3/[-
P)@_LT$-KBJ1K =$\BZE"KV,FKQQ2WS%T"LHJ),QE5]FHB)G:H X>V<%CT64S:8+:
P2IPU^4KE\L_ D$0^0('2#3%R5Y"<#F"5+ASV)FJKJF3.6O>D !TK@"FOD!T]A;_)
PS3UFAZ[VHZDU7*DR".05T_XA<S@537N?\ _;?(V35D!P*IY'EA61RX03X+:S71$R
P2MOC#@1!-I"@,[!=)WQ0O+?W%X=:KF@&+H+/]3:')RNA_@6*Z?"*_^(*@,. A-%%
PI.:.DU-8(0)+9EIS*L\I*S</N(2,5C ^" RPV%L%U*[;H^24;,>G:4,/R9D[3-FH
PK^[+9PG5:V&,1:#K?EI7_7["4#43+ F(@5\D](';0"7KM DXH6:AJ?$0FR[_G28\
PG-42I'69JT]^BF]@]XH'*?@#(7ZEMQP?<4I0>%CB3U@\@--EOZHF_%$MR-X<-*Y<
PEKH&(YFSHD?A@ P3MB9B"_C=7>Q"'R.0<]L17Z&ZGZ6A*&9@9[X??)B[^$+WK#GK
P;&@,P F!HCO[:5LCCP4" L#)]@NT&O40LV/L_$K76>1WYHU6@A]IU*1W/Z#&TQH+
P )=Z8;.Q\T*,N.IE!X&[Y48X<*#?41C ])<E%7YU%5[S/;.%W3'3"&AMT%A,_[ Y
P\#3<?;>:"<#>8X:BEIK[4)(_P[=73XL%E,M4)./=%!$.,)Y3[$Q,6E7"E[1\]*I0
P#WX@+ZA(0R%*=+814R\V,NR)(#QS9E>#_I[KF:I]3_:W\MNC"@HCB4ZCOMDS+M?I
PJY"]WLEQQ]"=+VQ?(SZ&\WI.@NPN"L)<,*>3T0GHIL7-@:@2.^Y?BZ?.T1])KGV<
PMM2LW3D/HZ,I:-J2>REI^X\1[E]>A8R'.0\D75$@D)1;V,"\MM*R+GC7T+^/P-#[
PO5-'OO]@7<(_,;] 2E/8Y3^209:; M^TL_*T)A"$D\1WW.>J:)IZ#5[/L@@Q6WI!
P"75<(1%5K1<EQ.//?'I,C:2_B[_H(&%6T]2V['TG3)F/377@NO,/4GX9K*[H>YZ4
P8S"\-.+!;@LBU9</#=5#__\P&FRU;[/I*VXMS 0>/C187W0+FZZ#?2IC/C_;'=N7
PP^<H5H\DN8S".<88"HHY2+B <8T?G.C(\&U*@[E-=A,:KY+Q9F))BYS3YCD@2X4>
P[R5]!)UC/MSUZXYEM[HSDKLK0U; JXV>FB@@"9)!%>/8VB:^5;U"06!1.:#*N9:1
PNFHR_!I35H<C5+VG<XNUZ[AD$YRH38G0I0=C<3<U/T01:A1:LZS14X;G]QFXP^X?
P10RX)AF8%"8T5-DZ?8)TL)FQ_@MP%&?UAX&D[N9TN!QW4B,2W?.\@N,F"]"Q]Y-F
PC;PN3AER*FW]9P8#X\R1Y0ZDC;C48H-%F*Q3DAI3/?^X[!<GO.D?L'"[L$>@UZQ+
P] ;V;?&#9]9YZ]E:#"2-^ MD]0F'VT;0=]2O(WZP&B@TS&?31<>.2;02'R8[T>?&
P.77Z7GVONU>JJ+)F#=:=^.7=E)$8(U45DVT!,_$&G<H"$JLL;C],7!'_*8PP'KL2
P<-WMOPO/"#6N!XASZ3<./ME]">M#4Q%GD"82&BKLP5X[\@_4"7&4C/%G333"T!?$
PIMC<J^J CTA K.R0UI'/<5M=9KH6\WIC-(_=Y_L]X'1"R,TO*6$'I4ZBWU[,:H__
PT=9@U;< V:96-CM0FO8[4,-S&(!<9:+M#@ *ZE8#9FT5F!9\[UF-UR05UB06-NYR
P6>@5LYJHV#P.:7UQ\YO7/B437/Y^#/=67:TG ] Z0(X4!/!P'V[SAAXO2K.X?ISJ
PH.ITG5=/+  $[BH8W$=]99HB)+G\MHV$[<.Z_Q#M@I3&Y=F#T@QJ(86XA>?P<8]S
P(2)XE'@DL+F=_[0$6D?P [OVS].&H72BK-0#S3;HDI$"PC:^$D/G57F*$G+[<_P;
P9,%LF/&@<R#;'CL9+KU9++? F]H,(8C7^KK(R 4]+ FF&&L<YSHUPY[!EX.>"6QR
PR34@,.+!.2_];]%%/6[82$'-S#!Z9WN:R,VK82)/(E\&%3BUD# :+(VK#8NQ+/9T
P$KY8#^'+-CUU*S[98::#M>>HGB?&H_=!4=;=9-K6!\^M9T8VR ."=7"*B!N$<#,!
PD'P8+-\M9) GE+7#E%PDL=MW2I#]S%\KD4;#I:!QM.E3U%M!V#PB1WLJE2%\>#-O
P2'Z!^5(9LZ,P>./2'YXWY<%':+LJ^0_)H+3#OZF'+3.$[<,=3=.B$HC-VITD!=&U
P<L@2JK?<R,]32[*.+4B3:L].[W2EOIH4GF;B:Z?_Q$G1 %UX[5S\=YGR2??JKG@8
PY=&=/[_1_A*WQ3MQ_TW2D&9M&G1>^$+7GG1Q?PD'="$=4R=GK'3^E"6NAQ0T%J19
PDI0[J'%]<Q4,X>Q,2C%BOQEZ+!:K&2VW-'N&C2#47L%><BG!Y.A-UUN^\G,<Z??U
P2E"4 $+]0M5[.S52>"/K[*2;/M9*"7S&8ER8?94#M+?K%#[K@&+^]8^T,5?0R"@_
PA,I9G79.WBRSVY4A_>7 <9O\6'P<W*0+GZ-J&A9YVH=GIS>XUZ*V1G;)X<^.E($B
P[.\53.MP! )AXQ3I_W*2+$16-VM[057TXN**HS N$/MK*P.$18 @%AS="&'Z<B>2
PP7'&7W']>6HD/M.\YA*WK;"@E(HF\#QF%+84+98L%.3H]IURF)>"B=B#H2S">B<Z
PE?+1,TNX6S,Q+L+2!+IA_;:W,Y5.F)<)T>,C$[Q-"$2P=#99I)R#A[I75>^C&.DM
PT:0CQ8X@LUPJA/21DR/TB95!6C9^\4(8YFJ/G0;[C[L3)Z(;OF$-0$%"C^,6ADJ=
PO[+;_#PL,\1IO$1.R/?7[J9#V:WX>5&+W#$-YE0C ZV=UB_<30F\K*MEFG$1NA0O
P_UIJ=2WYE>C]DOP7EZY;K#U,PF@V^D=M"JYC4]C?G5S*2ZR??]A$UYGK3N'KI(.:
P_%+\C+_417MJ[B@P.MTI4.[.-0P91T;>&_(,MYU5JPP(+$.5KRNG]J33R/[(7<_#
P,D. +:R<FPZ78*FO-9B(YG0H57,/_Q0$@>:N?_/7]R-;&*BKA7VJ"?&PFT.'22TJ
P+M\C8Q)*&[>/\MNL(1W,Q0=U*02^EOM6LSJR-B\G]0WFE)"YE8A0"2KL%^8FQP.4
P/*8X1FI,4/&C],JTH50H8X/ZS:L_*YD:P'B-2Y*6I2/(=,SE?D"W[6#%N'_%%7\G
P^OU1HD^%-*S@*9<%R84(8*7/=FAE?(K>J%7H-_@CA(S3VVP0I >S?0.*MFIQFG:7
P#AQC 7*48OB9,'X .TQ+V5!(Y+A5VS],!@Y"<A3842F4/B+B&_UU9%^M5X^D@P72
PQ5Z]*#[*4];!5Y]%@J:1KHD<SWW*?HVD(/O,+,';I#5'3NHW3ZH8OVND#3]BY2[S
P[^"N6F]HV4[WN?:F#ZZ_;:._AKO;P35%+\TJ!L7N'A)LB8%0I>FB4I;_OPY_293G
P^EX_OX""]+#?N813S:8)@'%!F]4IB]M(IX&3L96-5X.X%"5*DB=Q+KT-MFO$EU1I
P@]><I+&_JG'G]6W[+LF>&_J^K.GLY@<9DOILGCW;-,)$@)R]<>NMX,(WY:%6<1)[
PUZG>KZSJFH[Q8<[Q:3E.>R"*EH%D3%%9R(^[8=]Q\U2-XRNB%%J6'HOTETAPFN*W
PIV+?N-G)4B,<:\U%MOV^X96NHD:;-^B80V!JW\)6+HT_-=SS9,SP'&M]C-Y\.$B>
PO7)"Z'CLH2SMK(45>;.I= <A*1X._M[6,1T7>.H"?!%.8?4'RDW^0_WP6)/T^G"I
PF"-G6PV@>_OH:8MN.SG\:=TAM59CGY7X1'WM%_.,EW,[MN<=#^BTX9[SD<'8/;\_
PX.%+"21^P!W6"_+NI.Y(Z5&URA+#="R7Y^TQ5*(_1.9RN"VA:Q\65^R,G$M8 C*>
P *-Y4VH ^$;IPK:B/MPZV0^OEQ<"'_.Z@O.O0HT?4:TGE#<U/>Z)414] 4]1:P8C
PVL3E$MJ<,OG0^OUD--AV>,;?NZ&Z.=;X%+M=6U5NEWW'5N6VS^O]_3(;1 .8*TA&
PLQSI$&+7/52C_>F="#W4!1^EALQJ53$+>D3@V/&VO3":7+:P>#T3X"I'Y=#4.$G0
P[9XB+_&YBUCY>TW;238Q6>@X7FN!0MS<:"8PS2[3/6-72\AS\]#5>_B,'EV948VJ
P[V4MP:]U(DOE+?VZI7; [8<O;Q\>CB>4]=Y7BZFJALT<_GM.(^OJ<8X9*(CXXFK]
PC)FR0XDH2G;*-!3?*\41$8 8%;H'G>$S9GBL)&ZKG]O)!J)DMD65PL*!375 6@$.
P6K%"9A1%$PWG>+*RD%,7AA$Y-#B16]/_]?6)9#*\GI'9T[3=E._9=BAM7PUE,&0+
P60G(ZZ#KNP^_\2/7C;0R]>5VX5I_U/S9H58W4$ED4<?0-6^([B"V<;^]!?YX#> I
PN&Y3Z-DEE!7JWL55N\2YY5'"C[&^T<H=!C]<%!TF!R_31@U<%2@$$W(\FA(1*'E*
P^=GS5L0Y(C0OY9&="O[CFO@C*L3$?J=/.I)0(T#K*NF'H#O&6%"@3K>)-4MDTV7*
PZB+T"3^C!R!":)5>F/(R>%3YP"%GC+4R^G))4)Q!)3!E#I:=^# U$A>"V:Y4R"]!
P=>PF[G.?8:$ 'Y?=7_/T 9.?X!48>(Q5;8HI@-P**<=!<^\.>[AQ@5WKWPL\ CZ<
PH_#MG,.1/U!$&O8RJWDD"0'89E2H,PM3S';[@T#G8)J=-]Y?XH=\+,Z#OQ(S(]*Q
P_,8!NH:#!;F52/T+6%])\-.E8Q?TB"4,YV[>9FW>(;9$2PT6Y )4W/VESNQNELD@
P[0RQ;\--*_(Y2[33+X\\[X4WY9'Q+Q\19^,=Y> /MDL'"_1D0(HS#H-13GG)'+*^
P@/\.)Y]29%K^H*6OQ!-'O&C])YH%#EE+N3"^=VNL04JS3>5R3T!_&[R<)L9U%3"W
PG=;7(F!%>%_T O*X;Z+G,!+78@M*FO-RR,%6_UK90B4#M*9UQN[S#L,A,7J"([^6
P*3=9#Y69OO+A$X@X@R91\"Y@TG)A(I:K,>N._B?$?0H_%W;?8!UH'BP5-AT2Y;>0
PZX2C!2HUKWL>J*H#[#M-/;Z$NZ1NZ9* PN1$@C$'!%\5I9N_!T%]K56^ __V::_;
P_T'J+2]97H%DAWM,6)S>:PV$]-C-[K$>6BNI,17V(VPP50 WZ-B"&F>-0D_RN7R$
PYR3LIG<6%R!M,RHE3&#Q9*5-G?G=<"1PM0OZ=#&G[:^H>NX!_8$4;WV]E3EF:O*5
PDH4.Q+K99]/=FKB[BS"LY=HLE(8XN*Z%6,OLLI<(Q"+7Q)C"C[;R]1(V)H]K^!4O
P&7YW6]'\)NM<CTB"D3AVN:7SEJ3X%S?$%TNY9 !,PIH>&@4&=C#\#8!I0V#B;S<Z
P1KL7"D,CXY'G_EI&\%JG!OO=+WWZBYJL[RB:&[^#97G#=;(1Y7Q=/<OX1Z26;B#R
PBU+.XQ18'P=8*4+"EQ2O5R[G^O+7'P*\D-4V@K['>^8T6R&!@^)F=0M^$OSZ *.W
PT#XYXS"R71F@V)</A.0M[I15M"5QK',!U4-TJ(OAB>S.J7LI!E\8R7(N&T@O/+J?
P6]?2U$NQ\,C\']ISQG)X0"%*Y3_JL@+4?]:?J]P)G/SB/7M[T3-HS8:1"-1.\2^#
P X_> 9B?CJ4C&P8#87P].!VD3WV^/"[U04S9%>N01"WX/>W.U+NAC.Y6'?JC]R^)
P2&W'>]--Y%#.#^F$<HJ]J(6(#A(5K_Q9-1EHTVHN%OTX4>_E._&J0NU:07F)WLNB
P!7(]R _#14!B;!P[0I?UBK$X_VQQC3B/:!TX9 4OY@\P1->P]?TE>J]TN_>ETQI<
P16.]+ M09'NS<O:PE=EN(?A9PK A@4BD=P\QNP)<S;8GXELD\TK,D.6J"W8@OJSL
P0__@QNB,5K*Q5N4Q3HD/L7^/S!IER8'I\&6L\CF'B5LQ?1P*+BSORW7S-$^@Q()N
P3'7'UJW:?@78)N4FX4<0;>F)C#=!=D&1R(7LG-YX,*EZ:59I,U?0NK+<(C!1C27S
P@(@I#W7(<W&ZGD QVZ(ZD/J:RS73*XAS ,0^I\]I%&QXID[0T>*U>BO4G*]$W#CB
P-.I,<A]:CY=RS#\XKSYJGQ#7.FI6$U;D%Z-]@M&1IJA1T.7Y>=)).""1PA4<[=_*
P..=Z=T4SO!+3(8?C.+_X [5$Q.7$\G1GGS)($6<.D<DAH2>T<!B)^P</1_O"RK!W
PLKV:@<'2#S^GMK^6#EZ@4B"-'?_D[DY&L5]Q%-T/MZH</4!)"2Q!*Y2DH/4> N2N
PFQE<PKSF(:+$_Q:DW1VP7[78]35(J1EYPZLW]4M"]EES,SK,[:$B4J1F[U<:C6AS
P6'N=I6R0Y P5.R$] BR*QQ#'#YUUR^ABD#]V$FYP\TA7<!00B:/R#]RYG[8C[D[U
P]!.GV,&LT+A,K/P*%@O@Y>OPO:&*^<7^>AS5UM(7?V3%H,T*<E,<V.JA;Y/4C^#-
PLX?T51%VF3\;;MWC#X+I:"UA>NR6,]9K+;:$35IXDLY+82D1>N]8CAQK3P_ F)U>
PGK%MYC-\NF*"M810\%+L):Z8]?V@;Q;CO/^J\#\F:PTN\Y>;UR[BI,B".Z>XWI!<
PN;?@N@&B)'98N@SH1RR'TF@GXUC<9-SZ''#U2879\X?H3@^"=S93UJYMQ&M_"?_R
PFJR9T[3ZZWJV68D*O^)@M-5R!*T2?&(QM]Y5[>3;EYZ+FS':$XI73Z+SB??)XS&W
P)\?7C*0YNG4?+QG:9'$WTI0Z*(U$Z<X3Y#NDX1\G:F)S?"L: '<W$.4&CPWA%2L>
P!<V2;4KR0H'P>Z=].7A(R+\_U*%?%V^NE^//0C:RRF#YW0]6)O.K8W _$FX),,_N
P N.JK)TW.(Z#51"^%=Q#:MUH0Y[+!(-O+;-" SW^+D7J ?%/3L7PW*IAAC:TY_X6
PH !G$CLQ.V0!I$F4+&@V$4% "_O]<&1S;2:UXU2K6HO,/4Z@@((7B1(Q_JV@(Z;)
P_\OI,A*RB>GNNOG)%SZ,2B^P/#^6Z,$1J A3_T?% ,SD.M)II;7$!35I5P[$DOZN
P%<+DFQPP6F7 NVY"6C@.,YF!OP4&J*S_D</CR5P5%<S\!8J10F^-XY(:IW^ZPI0?
PL6BKWE4*O=6>CT5,A>5%R"">1+G\#$S3%<S4J/(R>21A<V=2H>Y\9@U>MS[#\7:G
PY&""Z-P*Q:[A[UI5MQKS0_V$0AY#DEMPB_!=%@",V!MVT MDIT,:[NQ)HWSWPF_<
P!G$,-(]*@D4:JHA!C6)G\6Y=]4M$KWC6O+IPVIA63\!L?7J!J##)%;7/Y>B2K>U+
P+DFS(J!^#KD6E0&GEFS(<'(K?,F^O3U"J!)&W(79^1"[XK#BI&Q>/\,F00?$^/1 
PP2P-+Q76>*+007_Z@<T_MG1^!_1!/N\P>-ZEJX9%3)$Q!R;U-X[DW4'?6ZN= ":3
P.VUJC 0E+?,6"V&KAJ]Q*[M3XYH9KPS==FGLB%Y^G3480$5=#T6HN@#I;,BL$:7:
P]-_#*GJ;V)UA($BH88+94V7&AF;7C4//'O[<N7E<N,[K]\NR,J39V6W&4EQ._$0T
P#:9.="RI,QBQ27[5D.AH3;_03Z*@:"FK*&!*D:RGF387<[[?)9>/2U:EGU"!*6[,
PL)'[H,J=3H!G=#&#;^"_X/'B1K*>B$?9GG528(L\GFF[I6M 23X[(WK.%:N1+60N
P&+M!&U8U)K$;EL8HJQ6K?0XLXFETP:Z-S8377\,]7T[95 0>CV#JU4]C<..Q6\FX
P"4ZWI$O4"TY):;MOZ])26@HM)_&:2+N5XC.-Z+VDD[^1E=U"/F[X.K%=G=B@_79 
P%MM+0:I;%B=RRX9RLD[B&+:K/_7)I \!YJGVV[$$R I_],H3-?\.H-EX-$O.D^S#
PY'W [9VJ.L_L4J#J2<[Y5(@9U70"1$1!&RWMMX+8)MH/H7,E;)MTWYN&O@K8TA_!
PC63"^Q#O^B&<(*X>+X< !@<#%4KO^I\,B)0(^DY@?XYW5!@"ID],'8>/RDBD.FI<
PF),EDS,.:UX V&3(-+JW8 ]*+!.B_[M/I4-+[051S_KFZU!UJ. M6BRJ!^'5>HH<
P_JXL/Q/J]SG./T\< A@[K]N3LBH#YU2 XK>';/','2 5%HY3BQW^")DNH )A_?MT
P+1%Q! 9,U<;KDIFWS)1"(=C?)JDG3;Q' *VV[R+CMRW*M\[L\WCDPVA!*O[A1R?(
P'%7?:PXI"UVK;M"$6?#3<#03.W]O/QU)N5)*W)A0.51G#*HC]D/_#\] !.5U:G=.
P!LT;S E.^<W\HOE*A5Y[%[J9T$*D3-]?@*>&@ZQ4+? !LR.>5< 1,KGHV3_'MQ90
PKC3S@L([E#"+(,X^EV^QI\NV4@/T.%W5C_]K52-$-)=O'"@7FQT"LI3?;9T"0!LV
P-Z6T1@N61Y@+Z,US@]]79+\VP./JDL-7A?X *5MY79&$.,R$Q&!C59S\@)(?R)! 
P+'J59>P2(2[/8F]I?'NMD572D6T9C4O.HQCE?FGX=?/@JDRRX%C@TVJ,%S@7H&I0
PH\KH/EM-M+P6<M"GFCWQLCIF:DKU#LOTEF7UI_@-'>)$\613E_/UV<O/GWW#RQ 4
P<A*]\T[O\88R\ZOT.=!?B6XHWLD?6+6[! ,KWN]T%W@M_V.C7I8C3@:..AIARW0(
P<LSBZS=CS&P$9VKG[$KLY;[9VB<K.7H2SK \$<]9_?D87.35K"5M](ME7MN&V.(#
PM:4'7YC;.%>#XZG#SUC^#] TJU=B9U@/L.NS_E[>>Y" EEC@3X8JOO*'7>^=^EK(
P(L\='_JI+8F7TM:L=AAZ$58![ !P)=ZP:Z7.]^R)!/NIFWX_I@3P_0-K;W6D#-@!
P3E)/3>I^CJNTC05(BN8%C6KAM,@:RB_R48,P8[*.S%_IBWGMPIE?6-I"0X+[B(00
P]/,&D)%*0MU."V*:YA_'QZ^--9,'Z*P"<:L6X:R[;O7W+RJH'%[!4U8HX.;^>)_$
PI^(1($SZR>OL5&/W@L5N*T01NAN2^1<(JW+PXV1_#3G5@0P=!"" VK@_D,]C*%@Y
P>>)F8D82]VG8;Q@Z0!C_.-=W!#$66<H]_*0/-"#D@OBO;!975.1TH-([.T^.[92D
P(-K-)0HD"C_(Z0 JB4'5S2"F4^]3BTA$__NCV#E2D#@1^?!4Z8A;$,O^O6DJ3\W/
P82_L8)>!<A4>MQQ"XJ5JO$\J54YW$_MXR/68V)PM)B-H'Z_"4C37K4 5GHF?7+9T
POF)T;N@[L[A-4%P7+><G1N+.,[ )S=J\I_M=&F(_-[@_0_XCVS4$](3TDFJ-F[)F
P6T77V?18\57-[4KE(7O<7?*/\<P0?Q=:L6I@ %[1O:V$X!=77@@7<U&J8P8]*E:6
P 4WU:!%D_"<+QPB[,8>@5*9%Q@EWQ,$O4IOJ"56[V3/8:A\6V-+"8_CIM0D8*P>,
P;Q?')C\Q(9<UO(:.5"-SM( _-D/E!9*6M<[1DU"5"$+,NF\.[U>2G6G(ITA& F<_
P".AL)GYKQ@>,DH];%-[4%R.Q*>@G3E$4^87J^S(@>T>J;JKW(LTU3G"E .M[3@7+
P)8GR'0C,/B-#2RSM+U?XHUO A[N]HJL;?>R$U/ V6.@3K;XDBR[(R%SXMTX2VNC5
P&U-B*7OD"2^GJ8ONR8"FR(P@>T4PWV6!')NNK;-?4:DY0?\.'=>',)'C%K#[9QTS
P-S+QZ[(QI^[.BU])!MG\E(F1/4_E"54AW^A3U3@/5ZWKRZ9EZRSH6['2$V'HQV_/
P62B,/O.2A_P-)J#.XSMB 7]A5,;.P#V 2WV9NIP^TB;L'A;\R!("UT\81BM.1^+%
P:@I>W!N@ZGJ(3D0VSWYPV3>=J:E,?D*(R4.M)C_8JX=%$+YK%-7=$3W@/KK=9,Z]
PB8&B@[M7[R7=M%=M7S'J?LV*U5B+<6.!C=D.>T.79[W[H<2@)QR,'0I:SQ6R31&R
PLHYU/I0%I*C_Z5NR7HR%OYNILA/S"SYQ)\I=]NEE#+Q;ENQ;6SKP&(+&#[XJ-4-V
P*AD?K_:^**;XAV?<J%'7K^3#+XFA"6;74P^2,TPP] @&X"HJ=X2\0CRJJ'3ZQ&G!
PZ3NXE"0WY 0U=FF[(_PB;ZQ, N9W2Z?/4<ZMU(WI^+_:ITHGWQI(9?!>)Z^&@V_G
PQ--DT^/CQ0GJFOSAV3N6 7\@E6:W+C$(-Q<,1X_>_"!!FN4T-V1]>]%?[I[.]LE/
P1ZEUX6#'0,0%FQ6ZPR\MS<-RJTRNUAI, __6/VT4M:.&5F^R!WN/-S8=$"D7F&K\
PY4/*R+HW"O'[WG2/)T9F[7VM6#;/]?GY^GU>T5-4?\X:!84P6/)TBP6%XKF>ET&N
PQAA=)U8@D9%+EW;_&.ZZ@5NS-O>TK#%@KHK'X.;)4X3[H.25Z7-+)1Z4SC>N"155
P-FJ14 D*  CQ/:"/B%[YHG$)>-Q#<FCBKC"$TUO7Q&_=%%6^* HW#A18%TZT/AQ_
P8BOFL*8'&<K.!D<K&H&I,0,)(@P%Z;\>)2)!V$:VGI+NVQG Q5*%*?3W5;)*8XO.
P#?!%:;,*8Q+6GAJI%87#IA<*1VX0->U?5V^4Z3@1 DO2-*L##%EV"5E5WP<9E]+L
P;2;2W-XEA<D@EN)1300<2RRP%?<H5AC39M_3MF;PH#H57?P(@0"77#XP*TAHP,PP
P,0W?:=9 ;]RGA8F4'W)'=R,QRR =8[K]O=)4MZXO@2HHV-2?' ^&@ O+YW#LH97A
PN5?X=$ND_'9KQ$^)S)L8=XB\(;QE7V&D?:;WO"8)Y?2-\[]G_%H!4&-0("--"<W0
P"HYE4 /0!.CC[RD;R9I)1-Q:/?JX=PBX0; MC!(,51@=_M8!G*5F9H5],8]_P6CS
PWHO?X>_Y/=8(B-\6XM&3';^)'.]ZJ<A[L]4!B=Y5>TR/\O[YT+R-^I!@Q,+.*6V$
P@1$*>ZX/PNL#?,S\8$10I14[CR.T!8VB(I[X=9TB]PZ"%LVY&=+,YGS[L?^N6WU8
P"?!%GS[W9E\LW64((#';DB"TO"@!O14II\M-WQ!$Z<WG7294U_(!FB@?"Y.B>K9F
PY A>RS_=2&SG6F$9L;:=T/N?"')^E9<>B.Y#7-+UMK%I5/Q3Y\\K$E5*;83!1,IS
PSKA(0I_]6DSPE^^:":Z*#H!6++H0)9*\^;3C/,=[70.2,J"4B;_]5<B22D5("A2V
PPW_?MCCR_2Y6S&DT?<"#KDM%9]?M^N/')$$[9;%9+D?[Z=L#PVW#L(7N3R3]<3.5
P_=!'Q3K*H(E4+/RKB_\_AI.'E3Z:&J3YAEH0S3-\3]P -7P4BA^H+X_WK/V*^8+7
PQ0H*(2Q9$2%L-0@B6W))_E6.Q'N\L4[=W61Z%L22*N#Q*']CD4X4 EN&;$94P/FK
P<USUO'P ""W)P[-LRCN [#""Y5'C%A]&O;\)/T6C411O=3:@-N 0AK"T@+8Y#QL?
PSZD[G\..1I+*UK$"O[S#><=8P$VSPAM!J5T2^\A$\#O@ 2:XV893K^91&*&()W<T
PNRA9A:EOFOK[6G^4F",.0@D]QI))80..!]MP8*BY6Z&$K/=O2QL91M^/^@-1&)E+
PI@58M3AW.O[[ )P.+$JTM*JB,GIY\+""RLEZ^J.6V3FS3FU,S1FD72U?8M]!X%;H
P7Z=0:G1/A'7@.)R#/"OX<V<^C&YEO6C6@(=;$RZJJ/L;3_O3FY>!9\DN 7W/!*5I
P?=F 2[C[YQ-0_MHMD"32R$+4/QYWJ*2\H4O#\60JPAP1BNF%P:B@&#QLC]2',9UZ
P35/QR"2.1X>H9B,&Y[&T'6=_&SANP7X43]O>G-"+5"AI#,$#U=?]SYPGO'<O<"YB
P1F$V)3/Q2$1X^#PX_J;2G&D)<6AEQYH<$HN(0_E@_%&E7NLL=#!+.:T#[[HE!RU8
P='2$I8:ITI (%_J_R9+C!P]J2>SKP.:I&_\<A14 (<?+"9VY^\'UICRR-UZ];(ND
P?^;TDT[L:%S%#4A9B+5XG']R;6,0H'^0U-1_*CZZ?<"G!D@/.*;<I#>RL^\!CPQG
P7$N90XW4H5Q<LU@3OEMO]I1R2*OI%$I37$TVS4N&6NMT-D2=V++-:&604!_-Z];X
PF+V>@J2).J6</*]M)7LN=6HTJ?:X42Q;0*]U?8<A-Q"2!<+D3M4CT=OGW%<G:#/ 
P1IRFA?#C80;X$TE@J.+#N $D 5Y8,\F3-XRL&LM_+EB#[N=(8LZ5C?>#>;)(:43H
P7R 2!3^'"<")^"J'C6+)Z5QJM0_!X_UD6WV9(^C9I_S-VC1+I3;U2;X]GZN9/D\L
P-\ MV3S@.6&#_<Z5YH\RI,#;Q3N#W2@*S,V/.1^Y[_S0HTVU5"T?*X$,-FB!@G+0
PHF1PO?(M&TP-SU&%1?3QM)H;(Y"4-_15\Q"X!NXA!_&_H38.YN!H$;'+4\/0L7N)
PPTWTG9.BC#?427XX+4#B2A;MA<]>HBN6A3ZHG3IK\#2C#^5H<-F?$I(A@CE"@>-H
PSP.(S]P8 J1,*)E$K@H11#>;CJCJ%SX7TR>REK]A!.U:8P.1KED.?K%=M3@/]KX\
P_3)K#=0?B4B"9G.^.Q\[/4&:BU77/PA2)-$1K^\  EOR9Y^>8W6C53K80-3)#H>]
P6OH:[3X\(H\- 2=B'LN9ZO#1I)F(!K-6A"=P?7$XQ>M>M#2OOO73Z@N:Q?068L_#
P64FY&=;_W:U($QMC)A%(P5F?@L7DH/MIJNU0RN5<^R[(-"+D"F]II\S!(%_-':.9
PM4]HF!KHO<_CFD/\!?X@V=I0&6(:2L4Z%.#$MM@X8("N]:^ZS2[:=B-/W^N]XA'_
P01^5G7!='03B])#877%3LJ9^?X4RO^^I1^^<M>LC'I\]:9QEQ*:C#Y ]BE!/PM<L
P3URV5'"4[]S(J5$CT2P<K'X?AO@R0+"TS$/Y-#3\0J&'X3PX:E ]JM@$(*ZG;C\Q
P8_4?$01)AG8;B=B!TI'=FO3ZV T5>F'DQ.LXVGB!V5I&SO$#=GBF45AD/5[46IP>
P:[3M?ID5CS(@ 21!)R*2)TA,@M#5()4ZM).CMDI%DCNK?E(#_(]O* ,@;_80<;7+
P&CSN5R)?@%E"F2'F7;V -?B]JPOD'MN/^<_?B-/*&-8A;O%0L *-%[M 8%O;%H -
P+MDV_W&IL6?HAM=Y''XHCH"51);*GN/F4@'9!BXWW!VXQ^-O[ZODU=YZ,C?K 5LR
PWH)&VO/(*DGQ=WEY!+2O)4%=U1DMPN?,+V[@[R_,>G@K#DF]W 8I3C91@"IGY$=7
PSU;R5J^#X1!KIP>P 0#V&.2D=N1\)#* #PI:"TD11'3V_D#J-"5\<4"24B) ]$VK
P5/>M]>7VHG+8GID'Z-G)XSM("N[#DS# (!*NT1[#'Z%N.O9I>]*Z5L%)\P;YP@_9
P !M+P(_F%>,-P 6V/1OX%R1*[;X\P(7(WOF*,*WB!N#8[7,1>W[\^# V?MX$K7&]
P"OQDLA=_>DO3/TE"G3<D@P,.L%O*B)P?;.TTP4:4,1 3.9(JPX*)GL"ZM0(<34 G
PGR-F6^;KQ'%.9Q72#U\9=#RF66:*$4=H\F(SU]-O:\7L9T1U\NJ4Z3]9]>>,>ONY
PH@01&8\:&,;EN*Y;ELB,WH'KNG;^R%*8(^B+Z9M PH1;<*V*8R#L+HTWX&ESP_\9
PW25]$X)B+E.,_86JB])9ADM N)D2^YB!O+;LT2B2"7<M N;"!C/K*YZ6MG4!#GLY
PT(R=-C/YL!:4;=O=!+"^_<+KT)=><_+IO%B7\[+6(WP6R4<OB2M?$V(DOV(3MP5^
P*_;)V,P\7-I7X=,$H(0#G"_^IZF-'8M8KV L:U'P7>GN_6=49$9YB]PTNHGP82* 
PE MG^D,M#"Q$J=^P& VIN\<(T^_[5E4.8 .?U&G2!9.1'62="LJ:/'3HJ9F"C3]"
P"KQZK=:5;7=-89G*&LAY\>I!;*53G8S#0OF117="FK1XY!/E[=20_$MDHZ(>NY8L
PM]L8YYS..L+UU"9TC1A05,(ZTL++/N+P!5YB_0=<:"=;_D.BGT1(\(QIR7?1ERU?
P=KYE#0^4I:2GQ4_B[1/4]LH5H\<2CE=[H'"&HL6 *&77(0;YL/]6R&:. ?%V5KKG
PVE1;#.@0A;B.HIOGE]44#S&^5OR-8HB+)MQ\/#E=2Y)7:I^RM2'Z^TT27W2]3LR#
PB2%N, S0.@OMXC%$F2EE='"/KQW#W^\%^C_N3F5Z" U(%9!4K-^!^MA/[XZR=3U^
P$A[ZCK1)<SDFX/;R?6!L;=C3)&B7</',[RJQ?2Q+8>__R5R(90Z+AV:#8K<2-FK&
P]![9%F\-?Z!K);2\#*:?3D4:;8R)/V;Y2O>2&*!F"[$3C:,&<VCP$X%D>B-(7R\+
P4:)4D,?0IL!KC0#WO(3Z S:PBO7-3IZD?FRMS4ZS0!IW9 HOSWD!4P]0HXFI6/Q:
P"9T-O1K6@-O^/5%_"4HM)?J'*;4^G<D_I.S%Z)3Z+\:7^O(C9-[S=DL#O"J]5A3/
P:>)%W^F:_*..TRUIC5Z<D1S,^<@ON$64/XH=69#D60W9ZD-"!)RM=.Z8!0P1TKN8
PNTM?V:&N;.Z;*.JN%XO4)**"%/+HQU>[80WJCS%0D !0GC=>J.M-[;NJ$S,FG.O*
P-7IPV1]@TAM\LX7]Y\MJD5!(:J_"I<YE+X'Y/^?$S9 JQ;'6+@'-[CF*#@=;F_"_
PDLK 056B:'H&!WN*(MJFQ:-A$W.U92TG4;-R'I'JJK3C!XOQ-P5WGG7U]%U7OP+U
P NDF[(R<]9/DQ*4&@L1+6DJ51'9RCG[:5>#1+/F#*)^>PA;[IS]7XE0<"T0: ':/
P8C2C!(SB0QOS9I/EHWXA [=V'@<*BI.@."$2^HT<PT!R@^J ER$;&Y?MGO(HZ&.Z
PS2&G:=42.T&Z&CR H;HV/W.5\341 'C]=KK[>[VJ+"T$RM@VU?+TE<634E0]SF/V
PZ_@3QH2F\/4'@Z9L-4>NK4I<SWD20JZ^R#HS+B:!HG^$OW@B*89T,O052=&CU"L;
PVXVML=:V,>&9BK/H;"#-"];)G4#;G9C>?]UO5NN V,;0,(RAAGK$7_9,HD?&;4^-
PK)A=JB#'2#ZE$FF/TE9/?V61.%@V(PN1)?&\*TUC&S>A;1)>,T[%+5'#GL='9#C8
P@%%([?\EE.!<Q_9>04+SHT;<VWC@+V?JZ)C5\W8@-;F0)K=('?;Z&-^%%V1(;GHA
PLPTT$B4\>\9QBX:@\_&7.?CP/_Y?=@8P#.1^VQ%^'#88 T_J%M4MO3.6_^-] XLL
P&X<X;QUT-XW8D6-?"\Y2]VO\A-EUHP6%M@2]U\[>N-1(+B>^(7:3PS#!V J']OGG
PZ.0%\IO<ZHA? ^/ <YA8)V,!T1;+$/ KNV[WOOU2:2JIS<FN[4Z0W.TH"YBJ0(J?
PEW#6+Y[N]TICT6A:?:V; 6X]%2.4,AW VX<S@9RYD XSP:AR1;;[=\'F5GWB/$@!
PKVGC/M_NP%B3NI=6;>!DQ[!!4I*(*H18'<)..9M;=2>/'HE>4&R78L F-TOMMLET
P>H85?3S]6-FD\>@9 4LB%8*YMC0\^2*1/3M1HW],-Q-@6$TKOR_@<9S&(L!_'1DP
PE\8$^Q58/0Z^+E2=4<P&R6S8W<Z[0QTU>HBQK"^!E@X;?[T$BGBR=]BS@/RK7*[J
P+]?3^0/C=]7=E/KF0%%Z^4P,8.7\:W8@RH:O.Q)9EQ7!NA]>G+F.+@TAR-M#JB\.
PMU*018'L$PRDU9GE\7*]M#UHJ5F1++&(2G#BY;:7Y[=K^:!:ZJ?E^<U.&4*28#+W
PBKYGX1;C$&(2FSXN(7X4=[Z@C'L\48.._D$S*UWGNUJ;X)S\6^!-X>!R.;J08/R[
P*RH3GA0-NYDZ:9:"H';PP5J3#E=Z>7<^6ZO3KA9R.E_";ZAIJ>H<#RBW@+C5<$QR
P_,K:,KX(,$.PBS+HAYI$0=+#UN"H<!?)B@V^!IO9K.+O +$3NJ95'+1CL;[[?T-A
P[K>M!JA=TY7VA\4YA@ELJF(.'Q"F1B!'TQ9WFS(R+Z IMCCO@K/_::ZTL/7V#]OK
PD/&OKOVY]JTAU7G1O.*!5 T)YYL()36U0IIPN@= XR,-$-1DU]A.W/HNO3U)!0^:
P-I^(*'"5I;W,NB:FIH9PT_'%@A.1]VL/D:I<=Z)C1+*UL"M.DDEE>789==$LGOYT
P+;<-KL-9#&^0CTD+QJ)@2@A)IF/8IC-*0'&J;O>; +1LNMDOB [4Z4R8P1O(N^'+
P)\Q6LF_=!,\'(\9.W'2_B8,E*SJ9AAWJ<8^DF6Z*A7F$U@>VU9I(BD6+.?HG'A$@
PUT<U6CX??6\-QFJ&/$J]-KP^9-U\38TOO.#C3F]F,TSRMNE.Z'NGY%H[:YWVI^P&
P]07?V%%[(P4&J\)[_!\O01QY0 "UN9_'F5R"8#T,!?N3:T@*65W'?LWLMPR;'3?L
PJ13H<_/G?;Y1*;YMD*K-(WQO82@'-0?TX?*.R"M15L@,R=?>^ R>8$)M &>=)%"[
P0'E--(R:N\ERNHK\E'3O?-2Z+!74"DB#"N-%,%,S8!DYE='=[9VLP+>(#/A:4*UQ
PWG-.7<]<B#B8+!6+5FDE'#7JG"21(+ZQ*/L PE$C$KT!:1/@U^2CY;)^@LRG5'1N
P1BG0JY>4JH;%8)_-'K3#L7H#2BME86-B'F\ =0LSQRE:V'9H48V<@9[!^*SJZLCS
PEN<Q-;<(-!YI+]M0EV=43WC[A%=240@RVA(2+&5PR#P"4F %PFYW][FHCV*;5<#/
P_*PV9(XI:B /<B%%KJ7TI6=%7#>CL<H,@[O\T(3)'ZVJ8@MRY7[*$\'49MC]Y:L@
P+YV&,K;&UL)OO)#EI_+E[>>VP?<C#<'6[PLB2#=T##?;MQA(Y.G6WAV'5-Z3E]8!
PRVZ ^F1EAVL(ZNX< JR5+TK>E^Y30EMU0P+!1*^P?("RA[4!0:)? 6C,:)K[=,(:
P/STL-*R<Z!SYY@SBPG/>_QJ>EG<:UYYO/1CJ:H^,:OJ,@E]//D,9O?!&YK6=4A1A
P3B:'RUI]QB1.4&L=M+('W IBQ'VA"_7/9%B]0WI RDCJ3@64(6\+NR(S1&,IZ%]Q
P!J:H4]>WC[.R9OW_TU5G8&&EC>P3.E*_^J6^HI_VKR10/1T8DV,ZGD8TUYEG+K2V
PSI0I.7A 3A3:XEX!K^<O&8P5+!&KILX :V+V<+R/C0.=OI@P^(:D=^53+D%V>(D<
P>WHD&\U1ANH'BJ=B?ET;@QH^:TSM2#ZE)0V/<5#$NALR0%\CS;D59U!)[<0'_8TV
PZ1\VPT[)<^R>!0U(:['B"/<-]=O$QBJ*T_>6062.UFA*;A5OER@)LU#17.26 ;^J
PEAU T55&;;K4_5@_,.&[<M\QR.F<J"1IW5![NMV%O],,R +:P@<Y5*P>^];W4S,O
PHX?']H#UX_S^K[9C/<^16Z%Q'YM-:"$RFY 659>)OH+8V=#?Q.,<'(B>F?LHLL7$
PZF$=:L(ICYTJ@6)S1NVETD[4]E$A>DJ.?F5ZF>2VO!IO(,.\%[7OK5\(+9\8*O7-
PDA_'*2)(4?DYJ7Q%GU'UY]1^[-*0WDVR9]V)<L(C%SF#VU7">2HLIQ2A>61^G/+5
PKXH_CF#!KFA[#"P^7,]B]:.: *\0$,3B_XA;>I<!-]MB$D1,F4YL'L%X&)XJGM?A
PDA@[ G-&C;M5%6QP:&3(]&NF=.F[[0:]>S4DJXSSN0V>;?6S4!M#;YK7>MZB"-2B
PMI$YRW1WD X_J8V'_!=W\/I792W%M?1N.8ZAM$V33LIOR*5J]!7J0(_[L EMF A.
P6K_0SJJZXD/MR@^,/.C J,F];B'>=%9Q+8J_<_;9*5E(\]][2'V&)J6--E<,=\3[
PL6'O9($XTH4B@LQY@2[?F<&J(/W%;>4N+IUPPQYSQ8/;Y.,0,%N]#</WOZ[),ZL4
P55M>FUPL4:AQ*JT%@R"!,[%'!NP0FK6Z+QOU$A*IR9=A5:?*O*[_A<S!S=?L$B;!
P5IE+!Y./EUN4#BHV$;1<9<_;O&Q(^-Q3448AU>F@E[LO(I85KL:'6MA>09O=ZF;7
PA;_P<93%M495.7('OKCY!D2 ZKG A%9Q/:[V)F<@PMF'>=0IFZZJ*>'0O^8'0)('
P&.QHZ:6>4%4BB;(0L]\8D?F4/,&>=_A_^78O4<O,IU:??O%.Q]6_\!<$3VT1+P(H
P]PAR2.&H590='<H FMC/+FG43RRPVOXP'S&G=](B?+*495---Z[R&A+-^O$NUX+9
P82+PVGOKJ)Z/^H*N#<$47E_R1CRKZ,?_AQX]^CG5Z^$K,T,GDX' LC:%45\3JA]P
PO,.O$EBLKIY%7<G3S-1,IB?\Y%EB1T7E_!>V#@&K>%S=NC4YQ=K1V@)9J0P1K 6G
P00NJ2D30_ZUSKR+80/P((R)4YP*/UO3<A?W4<,C'U\:G1HL..4*O4[T1#02[IHR)
PI7]DD^=H8*%U=[!&HTWXPGZY?K9FC'P,X9)!<S#OFB@2PA_M'P5G,\(+\%"Q_0U/
PWLSZ'B* .Y56(T+X)4'LM#@=L@ "8&5<^Y-WBCSWU,_B/G;[O-XY5'1$!UZ]GZF=
PN30])GC>Y_79K@) 3/P2(:X.L!=:43HTN)H>Q[&29PEB"L4.M[E*KTEJL"/(8#OH
PH89*M*1UM=O^G==D;.[<82-P2O=V69I',OCW<,KN;O_4PK&6\CT@5 :FZ*O"0OLR
PY/%+FN#P=6W=39:JD%5"E*QF:JXL(.&2!S:.HTP8=PV,TSQ _72^ZMSG?M@: A/A
PP48"KM/RO5Y3J<):L*OX?5P1_!]8>"SL@F51,D]YK$ZFZ5L<?9M+^PZBTCB4,V_Q
P?"Y(% ?TG''4/"[%UYPGQ;>?<WHB7$L'?V( =H-%54W=GZ3!P8P1"&#@CX6;3E,+
PF.8(1;^$V$I$7S[Q0JU<6">*?,F5)@%=!Z@+O-"0*8UBOXY'(W-VN4.2L6^9G")?
P:P08I!:6O;)MDU;.5YXJ1(P-XCD 8$$XJ""$'*3>WNZ_I=SV?#\]@0*J/O4;32;.
P>M%\=I=^9!N&&E\Y%3>$O&&D!,:?S$AXP)=]Q80>'8;CP^#4QJ8.!<^#'"$NWYM%
PO5:%A!*HWV[ZF]?BS+[DN-H[#^R491I^- WE&R!74A'P:W%SO U.8.HJPW.Y2'!;
PI-;Q0AM.57>OZ(QV$DJ(Y#:9E%HV*T'".,TD_<K")B@>)FKJ^'>_G0CBN8^"Y[V=
P=NYY(EM?BT%HL]3C$=G6HS6K-S" V7?&1=_C(''&):92CXQ'L1@YT.&OG>9$G44H
P*11(!^?2Z;8"!&M ]1FI7[<.AM0?RZJU.1+JK>&W;2X43>7IZ5GO[( HZ7CY,SQV
P JJ<CSK2IIQ-3(JN,KB)JK?3\G$9R,> '/JZ8U=)H\=?RZ[B.;W5)^.C>\TTR_/Q
P$4;$GJ/F_J">IS@C EC?T-"8+B,B0M&*#J??*D_F5E\WEPXFQ^^7WK>B+*ZS58+H
PWH"C@CX@YP_>B49_@K='7'"0P.O!2OVVZ,N\3.6N8HMH5.4AIQ<I9E"8"3K(/;Y^
P>F :[NAU9>/7!T""+LYLU#.F1R%;Y/EC)2BG%,8?#L/,06[Z@@.,KW6I[% FHB.C
P<<*GN^[$KFK\PJ\" %];%J.$<GN?F(4;-7X1/E<XIE>%IZ7E\\'_5'^OQ,8P*&$4
P)B(6QQBPD4<TF*Y2]I6=YZO" ^VT^-VB_G=W^X4. )P>-5<:H^^5#L@Z\_S_IS30
P@N,QG\'V,AA3\^S69-Y-Q&6GU+3R$%=2QY1)CFX<NGY]_J#_=6D:9S?1HL88 'L\
P&YR'>HPE?PMG!;Z(Q^1*X0@E8[9VAU5]"_5$[<IHI1I2K1YZ/V?O*CQ3R@EO =*:
PJBXLZ=,)$IF#N QZTN,\* J-8Q)H@43,#TT =$A#P'(ZH:A+]!22.^IJX+X26XFQ
P["W*_\12JMJ.:^BVX1<)\2[!/B8039K0;GRX>UJ.]C2W3"T#_ &6RKLZ&OP-&>_9
P3*4RN\[T1#BP](!!_P;4Q0;M(2NX.QDT!NJH@:8PFK'E*K1,,0I; ]S6,-F8X2&X
P&E$BR(KQU0&KU#D-#:_ITFT>B>]W1+FI&=D3P9CA:M?!B+CQ\FSCG4DU2S)ZI:T"
P!_@9V?(\N%R4V0!*E) 00&AH)G@*\X'MOM6)TS>2[^(?9"/'<13 @5!*CK39&AVV
PV:]1M6DQK3V5"(W1?BK+4YXRO/'C6D8'SZD$HX,((.V2C_D38>[6(252KC"EUL+/
P3O3)4).XAY!WC+[K99+5*M>8E;9A)@$57J;#$L'0XE:KPB55,H;$77"&N+B:8.]9
P%\1:(&3W4EO8/3L_)5[<Z*#PX^_^O*YR[Y(?@)7?E$!U>Z *%N,;8>LM]RG?0[5O
P74I?U*0%<J.:O3/5AT,Y1YT@8&G#_C<C%JB!3?V6>2K:0<B/XBU' R]K63&J4[H5
P903;C8T^^%K]+'O'R@-B)#]4; $ 8P?\[\;PY*T6TMIJOE8:W;UEIB?&3:J6-([=
PATCHU%!^P-2Z.3:YR)G7)?'WHC\9Z7I:=T&?T^L94Z780/'F=!,[5X5GBQL16LYB
P03V3"O9F;=E0D(!L@S9ZTJ9^)54(*3^4U5WA+(HP/]QWFAPR.[]Y:"08KEYH4XS[
P:>T(:J\@T3N$;LH=92?@7LV&:U.!LH](OPG)_\SM0A\7%MUHD.1(7M ;H/D[C?EL
P)/DY(I7X><WYY$51:E;.LEA(AK/F"G?$V,S T7 %1;ST]--36T<6]L ="%7XR+@L
P!RY%WH'A=C)S%DL*-3QR1T^0GP2U.+1WLY()NO94=8PH17&M<K[3$!11,NX +U2+
PJ JI0R2KYVDE:A&8^.:U[U/$YL%PBR1N$X$57 .]TE>B -BC?WJZ/=E45EB+DO&Q
PF^X2KM+F2/G''&VA/^W-V<L],4C!@I\3$$$!SG+J,!9R(A';K7MG?U%35#)5,R4V
PO)9+B>$)0[]Y*HRH@(4Z]*4U$U^ES.&@'X?2^%O#8?_).OBY3.W,EZDFQO<D7HD'
PEH"5!T[$;>/L6P*+"PB$=[3&9E==4N+HAE%0EWROFZ^I0?VSW8@*>_D(13=B14-F
PF[IX/8$VJ/NWPE3)T5GRE.+WWWO;PAV1(OU3DU8>5#R Q*<K;$"3WLHX7JST+N';
P+2'6<Z'!;4CYV7*+%4].J<9EOF$%OAG\+RCQ^:XD9Y%W(O-#X6Z62@HL#)13:-@T
PH7@&F'*-(",IZO4=)E59N<?WX]IMC?*W?SL \=-!/K')=A.9$W)ZB._7][70,S@-
P39!#]02==C4PNC/"O#&HI# N-S2_80[>^R/2!E0H6R,A,/2?C;[RM(Y^ZPM4?/?/
PK>U =#( 6S?XC@ZZYDH;]I=T+T,6D$3'^7KDU0S/DP,<0WT%L!G+KZ0$NKV_9/]2
PHA!LP;$8UP I!6"ZWY >$V(!(K1OA^ _.JHU'XU+I((18I[75EDF[NY2@I G43!7
PX([VY=D6](,Q,QZ##/6H& ]N6X71BB$<8[,'Q1J!EA[1%XS_<RC%QP9:/#RK(C&@
P>=%$O4.6Q.'2A;.Z<T?)3.QYL_CG2TI&5\'3/NW0F:=H5&X%Q$POY4IA61?5P'I7
P?D5J);TVY]A#V"Q^G5G_HZ."A.4#$V'D64@HGY0SN[,CT<6K=)HTK33)Y_='HRZ5
P? IQ;D8)$%U<"S+?NB5,YW4^PY( 7.4,?$SEV];$^Y(A]JJ)J)3_VPEQJFBX<:TX
P.Z7HA0'SG(6:^]2#._]X"N][S#;G]RB[BL'#_;"/\"M&[EO'1G_V=PN=9:!.P>&&
P544UV7LGF7#'%35T5)008B0\+S9"C :6>(:EJK'-'6,)/J\,M_2C TU_*';AJ8; 
P;-/OA=AAGMRLV2;;58X7XQ>EP#[28/^P:I^ B^74[XN>('IYZ-M%2NFKVM+"!/UP
PRODN$-HJ :'9LF*B;^)HMHG.7"Y) ?9(+BT6T2&B)Y)34):QX[GX;,U2 *8#(AR=
PS^TDSS"34IA!(9Q"C\*E@GE5_)2E-@BDPE-#A[E';B%V S.JY,NBW :#!M3?L-;&
P</"C-J;,+Q=S9MC.!--J-ZU)&V5W -@93)\R<4Z4&16[\OFA4]G.#IH#OG" L__[
PN!C:--/ZJ[:"M#4;8D5V*:;3<>G.LPPNG=>G\HQR"1H_2TQUS^G@T*F%6PWQ H\'
PT.)R0AL(*P5:ABTY?,T$"'OJ_=Q\J^,#DPZ^T^JNZ6B_XCRI7YO!X&H#';K>1T/;
P#24H,4M%\Z:HXO_J7.:XO4M[ZB$1G>9QZ$&+G4=BQ!:NX)<FLHMNAN09Y2@FM'60
P;.5AC <N_Z:<X1' X@8[8>.SBDE#?7A?>9[@8#3)WY>?;#X&-8]0ZK=[G!^RLN0&
P9FG;OV<,:-MQMB#KTMJTAKY+UTDG:PN?T!O#3!2 ?9=TPA&7P3\X1R/L0JWB4.B^
P-E+CF^H6B678S!BK"OAVC*BM:D"HT;*-+@1>A738$918.=WP;RE@?CCP[ZEV3-KS
PF3"1T)Q+J$*5-WA-AS73@C:+JS/*T_RY[O%-/;P2VCS'Q8(4KCTB;,U;".+]=>FK
P7*J%FR#HZO(=PHMV2+)3A(1H#\GT633A^,6A=B_+Y@%R8['L)G)Q,2:<6<&_U,X9
PYE=7Z^89Z2=J%V!*ZPA &$T7LN6J'& [WN-ET<*J);@KHQ+"U1;AZP(8($$/55'E
P6LV'.HB.'N&Y*%SSX"6HG5JT@@5M&9J-$HH^,<MB2T53&KD;:O"8;,*GU6,/6'Q%
P^X^*U FSXDKH:K!$5H9694#^[$L8\-$TB]!]'#[]86WO]U.%88MIX5'ZVF;-P8%0
P?J7U*BP5I[UPU;Z)XL6A-0+1TE!-9],D7!_D%YI^9W8T1%L?VIW*5L!%B0A>_#""
P<Z5BY_B;%=3?&H^)811B!:T5A5':51*G:[EY+M!XN4@-(09IDVQ@G_HF,X4F?Y2Z
PH1XYS)&]\S,9B-)RD@%JT*2U)K^"J(+0W&(D;2D+5;;=MK9)'P8TR<6? *?D;Z\ 
PD<GI+I1[]Q-G+,;/:,#BY%F'0&7A_4WU-";H2+[;:<0OBW^;#',B'37$,]P82]'+
P&;F@3_-;M?J\]<7W4NG'<3DU_JN\YR@J5_G1=W3R!I8\!Z.U%I6\CV;'058W;5<)
PXC1:$]G"^S3_'0E"B=+ID$6 =YG.48V)*F[ V_+"I)SQHV2]B44993S<IB>JPF>[
P]5S'DE>_[G:ZG0>3K0IXG][;9=/Y!@6U$GI[]=D<+PO?,!]!JXGJ6]K_TK2*:9I=
P:48JX4Y_P!<UPR"*2IP8<CMHJNM[AB^L@PW=$.]SABDH2G#!H3PR?TA8O$<(MOS?
P5.EX!67@*OW'43^2J?E>(\^UK JN.)3J^X-6Q&UFU3$6B+P/W?=H+1\0$,BB:WCA
P!J.B-#<_K09>W"FG8EC>V\43J[\?R3_8Z%&6Z$K9"AW07%P_&=',PJ!FNQ(FI=&V
P'".$V(RDR7*I-+W\QZ_I:WP JLUSY)UPOB@$J>?DKS==JN<TAQHJG([.OE6'6+G0
P+V>3GVA&(]5=>\REX,D83]'M.]%<PD)%/4!!".%4TZ]C#-EXIOI)_C+Y(7*VT!8X
PO*C^>=\B.:5V*H,(L43@#%SE5PX!9G2'BCCW&,J#YK7)X[6UF]T.['CZ:!R6I 0C
PS)J'BD+DG,D&3&V!SL2WXBA<^D*-/ZTJY_N59?YQ#G:,K:V2!TCN1G<&&'G3)_?Z
P'IYP&"H .BI^.AK:]'[X1_*2Q@RY4,*;7.3_Y?F;<95;JMYKV:S85]GZKLN69&K$
P8@_LJ@F+N!! ,ZJT#YV4%[P:?GGPC(VI[?0S_V]ZBR4\19R@*!$6Z1HO<IT'NWH2
PN_TNA%2Q,A6&C)8?,U2+/BM_NA;ITAK]UABC"/2^33\[<ES3H@<7_"X6= 63R"L)
PZ3'@J;7S(N1'SHK*?_S!7]H5X(W/ 9/V&%)'$QTJ;:Y2OE:@&V*W4\QC<QIAVS/^
P-%RNPJGXZP:]' /\Y4_.S1O<N*5T<J%NGK1UINC7CII)?=US?(.:8[9E:<,N+E0&
PD_G#V>$\9"7>H?ZJW%N^FYRA=U85H;]]RN-<\CK6+J6* TX1!-;N YK0A^77ZKHC
P7^%J3[(*TIA.-%-8=_-^B1./FP0ST'3I ;IUSU>G>$@A+>BJ0'A:T3"4Z .NC2RV
PK?67'6S=+I\G/BGN6HI_I&IOK.T9$4#:BKB SF#>&=5BB>RN'[1_6W:]>4D3Z<V3
P(I $QW0 F.;/GS\^9*$9A+RB"Y\I=6C#<."Z/0PT&U87=\\/-<^D]'+DMJG]CBEC
P[VFB+*-7.YLD[3!:K(HE[\+*^\=<^"'AALI1J?A)78WV.?RQ5.3&/@+NQKT\PU90
P?_NP%TEBW[?75TIT7GF*8IW?1;4=&J#<RPHQG^',VV=P?KF,1BR0\M/IK^(5?(Q6
PHA,3+N.M'8!Y%>*+#&-#FYOZ^C6/E2OZ?,G8DUGDE-'^EL$$K$JFQ40D)JZNYKC]
P_*BY!3=UF.RET9POP7;V-%[3+2D(2U1P12QJ[H\M#(J0[IGJQ9TR=C2C2:A<%= ]
P9?BU0P;!OXI)L_>6"4M1>0$(T+9 60@*T=V+@XP]6%'PQSD>'<][8 .F60#T4?]^
P85W?H)L!G N30ZLS;_[\PL?)QJ*-2@9!5^%1?1?P*F*OF[M;;0@GW'@(HZMXK5TX
PGF 4LF&II>885W 79D$0T<;4"Q0-##*WB2U1B%$QA867Z\*E*RGQ\EO@ W3%,OS@
P(&3M<=42069 .L^O1V5&?=%AZ9;X*K"*I^9$E#9"BZ+FD,5H6- /W@8A"SR-,YDT
P4/S66IJ_4S(/<[1.03=@ 12UCL84K3 POC(X9G-/1(M;EE?FX5=;E(JC&ONVE W@
P$!]K5_T6GX[>"CKM,)J@FP,@^\./R0+*Q#QH '^HO;I1#_$'7CDMX'<FHW00F"2S
P&!KWNW97_3$Q^  E&V3-"G5RCTU[-J2X Y7/U@-. >W2E#4500ZI(K0>I9+3(JS(
P]9W.%;*MH0F&1[EN/]O)<Z"'H\MM*WLF%?K/%^V(R=D]6/7ZF);\P]H<7=H>;M(2
PX$L'[3$M#8!V_)2ZNMA\$C[&< 79W#S7A50R9&M01!>6'C&S9@)J*$"B/TC.\B]@
PIAU/\J6>3*T^-LG/);N7C1@GXY-*J!55^Y?BZ2O=-[SG_K6Q;G <D3E-GCLB#SJ)
P>7\B5VAG5M<YXY=-T018S6OQXL*"G[]9!+&TIRB) 2)YU9=2/.^HN>"V:P$3@(=K
P)K,A9DLG)].*.<K<M!E/OQBA1B@291 F@(7D[ %Z+E\JE>O-ML PBR>?JG+\I7_F
PT_QD+J)59N)1/>"7)9<!H[VQ1XFI?OX0CS !/V3@9=@<//^L%EWJGBN"IPI0O-@R
PSIQ5 82\LM4\V%2HN%L+=JEA .9ZKZ:$!G\G:0X1!%Q;7('<6S-*NO4$;^#>OW?Z
P_(5B4XV?8[?-]E$D!M2T#RKDGDE9K;O>$HY_[*2!\)@:U;C(\#1+44[2ZS:.DW_E
P3)9I'!R"RF,,*YV;#-^BRE/7.D#11Y*?7>L5Q86"%O$]#Y*88L;D\AEQ/'\%&TC3
PHFJ\U1SY$L%]3K@#C^+(L%[E3X_R135BL*'N"DI%V\* (O&;W7EN6+T8V]U7PR2-
P2:\.H>8=?$.TN9;&,B(Y.%^/R5/#>B1#_>KSJ#Q;33,54T%_EY3/U7DQ@C3@F[[D
PQQ=O5B<ODWPED-S8L6V>QC0J(M-6ZD9I9<U<\^*$.-:CXO]."39_9^IM:DX3CJH?
PIJ9K A*!<N&Z-J_9!Y+S@09#<2K''C&'%!UO2_!;8Y1BI;?ZKP"726)[/NT.?E\H
P3#,(A'"#[?SD;>/FYP\BN$S,OJ[2)Y"%5TXEY(K1;_T *7U%R3+KE,JW()E7W]8.
P/=_U?/D1$?7]2Y4P0'=OKHO/R*-DQV!MU+(2A5P\39\$)R(=$T?">,YN^U%CU!6W
P^T2)[_.E9Z3:HW!+@R%)G5BY76RD'9K=>EE:,FQEH1*4;/X+?OO\LA@3$TL!\_0K
PQ(J@Q-8\^ -#AU.!U,"8#4R";?AS['[ZZLM6Q*'NSV4NI-=P8(7#Z!3+O^YMYS<8
P<:DS1VU;C3 =!1ER'QL_/=*2&(5 \HW+-ZQGVHTYPT_(@207]Z?ZT9\%-;5,$U,:
PUN ).'^S;N 7A!Q4BV>_I/P;B='$-K;#<B0Y]*_#>,:<QYLR7<0X_V;(CL\$U9);
PUT6M%]'I37F?L.)^R0QW-V'?6<>%'WT[!WU'4JNT_D38,?2R/M1KY4U"B@#:Q!]K
PG>C*7A2Q2U4[F:YV4,7'RR?. YO5 U.]_X:\]R3OVX75MKW,:Q^Q7@?QNB-E9+4&
PHGN_6TA@%LL&/:T)5T.'Z/>DL+FFT?8,RK+5R!0*N0ES\L:ONW/*OH')T2?84R_A
PAM+#F ;Q;%XN9(5J#I*N"P9(&^FWIH,0W0\L''P/5U,8"0/>+/(@R$8):.O"Z#8F
PU_);IM*7449B9F7?!OV#OZ= (/G=$2RQ48.D\1:[HIED)TXQZ:]OYH/UEY/#A#3)
P""=YS(P$[H! !\'8%G'0?;L5TV&K<U]/N#;KCB<"WA8*C[CUQ#ZX7-?M9?0[E 2F
P]E.O70?]5);;<__ .#SU3'_"(BX9(GOU_"H'FI/;[$$6+.57MLJZ%)/V/>4-SJX!
P&R !F_#N:6'CMVW&(]YK3'%766H5(*?:H:VTTIG@*?FO#P(T%PQ6*6TCM]T-LZTS
P.#U='G.+-:,(4-U0JT&./L=T.<'K_M@)4LXG/]Y^ASY8!Q^;;A/)_E&O2QO0C6]=
P\@V2EK0Y+\\P"(ZD!7"==F\\[O6-BEE2T>49LM?@>3]:F*5'<\U&MNS"#(@G#55V
PX$4E6@K3FAHF^T&F+!^,IU8%%: L+MK"<S1O8=-IMS89<7Y37*LCUH<LZ9\_LE J
P-?;@<85![@8JY7=N<C+)UE3 CKE"+Q(Y#)$(>L18^G'?!B3$%[<S*"T;/]4T$TR=
P=<1V*\?(N!?  )'&UP[1\/J4-@ 21BHX_-+TK,"=$HW(,RZPNJD$)<6BV3>%W64Y
P*CWM6$QZ<R8&]3&6<O#$G6@+R;)&\V.>V <C<')><F&J@ALHD@:!]/LTEL3*-+XW
P.Y\E?_T^40.$L66*BR]8$F#@Y,B:\=P2RED6N_4X!X: SSI-  :!/<(E[_P\ 5;T
P56;J#GA*IS8.O\=S2H7R7OQF]V^4A2[5&N'V]]B+WGS-\)?\V"S!0_W:DZB&XMR[
P!,/[4&X>&*I:^GV=IL@);DP<4A*-QI8OTP=U[CDQA](%5R%CD?&*=5W=U=9] YM4
PJ#:_<K5:Q@'@!)9/RL] 0>+N!@T>.Y]5NH.:&,HXSAL"*\:1RC823*6YQ)LR\!\P
P*),$5W\CE]:[2QLDTO^$CB?9![S30M""0U7N)<L+%+TO,C*D/-N-.>S$V ;[J.X5
PZH^>(T97UE[D=(YU4@#3]+UA_H^^V2-4EAVX=EO;Q)QZ8LK^G/I"[&QXP0/_W2R.
PC7G :B/];CO_!)MCY[IPC456&YAS(8>I_"DZ\TGY^Z;XB:/@T-F,,X74 L%[P08.
P%]!A._/L"::_IT?I4%G7+/FZ 04\BE2&3>TP!!F&(B WH=O+FE]-U'9&;$/=LRVU
P?.U$H)OIA@ZRG[6.<"G?YV!FC&3M)#6W$=J//E!#,XSW*[TD[E*$46>9.X?8Z,_/
P,SC9.=62G4W[&:,GE('@WLS]N56K+XZ*GQV^A8\[N@\3RR&"T$=['7,3EWS/#0;U
P ^RPPH7#W85W9I*R:0:JVFP9C<[Y=FWWD!4,GK=<&X==<$9KMWY-<,I[)0PQ%D>A
PO;Y*F-EB/&DIOB[M%(E9411BVO+">^@>[F3$B&*VPSG99>GK*1!L_6W6MF^I-2] 
PG;N,<D[9J"^ZBHJ=#<4RBY1L_K>Z)JB O+(*2: &LFH[MZ<(\@5ZVN(5E_[UH73:
PX-V) IR.TPYY"9 _&1K;/@#X0KT3C$=N8 9I-I]DE>C^F<@7-)##'4.,* [2I/G,
PPXPQ\%A,L])ICC"V,NL1\&GR\K!>Z0RMS8N31<Z BL_]6N#(4R46M(WUK;X\_TOJ
P>6IGZDPH$=:@@TF@#>=I7#53PKV_<&][\3X(D)\$/T"K?]GS4/6'!:G!,^Y^^](B
P@$-N. ^N8^U'5I?8&SDKUXQQGU3L6JC?D^<AA);<05.BV1#YR,-JH!U-31%P$+&9
P/&48IA4?>/P9OG((V'OA"IJ&Z#Z QKEE2W&[G$V<OSV-T;<W@!0-T*+-">\7SG:7
PUYTR1;-A1/;R?^ADF#Z]7:^H6CBV%,6-0<_<4[G-[?+?E(QB1G"%;F^_/H81'!D^
PMHJ-1RN_]5R2FE7RA5".JHPJN>#RCR(]*7."U4AHYI<H (34_/$3H@ VK-H6+]_.
P(>?QMKF M>Z)B\FQ,_OPM(!5CQJ\0^.LL->_IOOH*(TJ/M\80TP*@T,5_-,"NZ'8
P__':3MN0OWMDR%V9VRK/_'>"3J746Q.FAX:=R6@>3GIU]6_U=^56/4JA&)"ITT%;
PELW#HOOU0P4-SNK:21FE/EN%1DS]B&.K\<+2G2.MV$8R@[,S/1L_%91SAO_CS3W'
P&3:ONSK'V=UBI'26)Y97(+:+A8S6MEAN6:N^U:_+UUOE"FUL6&D+>12A1[G$+'D_
PCF?1!T)C[G+&S74US<[(N5LQ.,).L18#M5\P,G\R"EN<8:8V/H4P:X)K.TC??;=A
PJ5H[A$RLY?E2HH:UL&3,>6T5^ID'HQ$^OV]X:J7;G25XD%V6R%#QZ0:"L+5,B+; 
PD--[L6V#^!5YSC.(N2XF9DV5]#PGGW3%)N)+$G[2*D?SJM-GUQ5[O*S^A2^EP6]*
PMM)00!:GR3[T"T)C-M'7*I#A9[XFDH4)9&&*B%GXW!B]M=!PG#W)/YLFQ@"Y=N1Z
PQ%1 P^?65U1;/93%5O93'A<S,,&[@!Z8:)AG%5=0S!!JUB/71[F%P4%^4CO&US!4
PGC8U_']^TR+@@GP'NQTO/'X_+A-)'9 3.T?D]\D]=#MC%HRR?O&>]PYIE3872LRC
PM>L!YEDJ!0B/P8(<R-E'_6_+>Q'N)!IM2:O*FKJF41C*2XX?^;9'NC4:C:&$8KDC
PI)E"BO6LH"-[PBJG&>#_C>\;WP%6F,5!%T#ZG[@>!NRJ7K8(YV1L)2QM<51I9@J#
P,9-@#8+4O2$X5(+H)U>QY]?)J)ADBH!F3_HL BL>K<P'3(RXX6Q<N])SFU9Z17)I
P4@CW8":%AD#;T;6"BFUR[X,M) RDZA_!"@"PK[_9V>-6EL>K."5\IY\I02!AZ\?I
PMP" L;EK^Q,"9KYC]"<B])?1B#1VV7>J>,1+],?C6R=,XOP7L#<-1*<9NI>#P%9:
P4P'D-H,S-D:&O(6@'>\JD>($:ZV$>BYJ+MFT8,T?7=-$Q*+$^<Y( K#)Y8B4 <_"
P2G+"'P1[)&H!WV2 G_ +.1-,[W="6F:LM X^S/=,@ZOAVGZ7I<V"36 &-B4R4_,E
POR]6'27-*0N]Y6+4"C^!JO @VV2TF@/8RU0.%Q^<C0&Q( ,94.]__HOYR0L"@%25
P.C9=#B0)$Q;#C&\]LP! 4(YO(&V D$E4*38Y4Q#-1CP4,0/!T\!6SKZ,$'3$E_Q+
PZZ"U)^F*R#Q-R]_3F9+I7]*QRL]L3'>G07.*A;N&PYJ6K-P4B11NI;PZ[W?'3''3
PUY/T,Z YU[5!TM7%.R<U1GAGU[5X;PS??$7@L=F)9-T:E^C"X8O1UR\^H++& <S8
P#&_T0APT4EL1<ED+=7DS74JSB^T*KF:M#*VC(8M6JYB*XM-:QC1)0/N1&Y0M'C/8
P:Y\;V"1C0GPJ\GUB>J>58O!;1"F?C!=G2)N?NGB(P,9"RJ7P?.7Y=XNT%&'*3NE0
P)8O/I#9"9_9H?+"^GA),QQ_%92NEZKO!)"?P!P2W^2KPC37(F-Q$G"-]*UR$=_L?
P0!/Z?NX))%/LB3&6<_>&*KKU7SEN5E8V\J\)R78X=S%O(GI_BK&LX(365T@\1IVV
PA#:H6#]#I<'I^,)(]6+E/HJKAO(V0\.<,G?S6U8M' )!]Q%.>/M\QB@4XFT^L&SN
P\J\BT^S%A&06;P;_S?I>MMAQ++U+OZ(JZOG@AR-#E%D!=05;(S?^PZ"=#BKP16*!
P9-I41>B@[TC2=R/KW#?.&62(9!\2D=2'*. L&H 6MO*0<K(IY@%+MT("8@V._5$5
P!W,%WDLWN,P9]%!6Q.*#^[I*P&?>N>_)4VWCM^2YH%=\#CFECG!N!TU Z&43D@^?
P5J>@1GU)Q-2UO6A,'R54;\W#HE%DTS#I)(X5GEA)^CF4>OB>O&!I#X1/H0_-.]T\
P1ZRMSQ.10,H4!!N]A>6P3[%$;7H + __Q;L!MQ]>6@XAX&55BEKZ+#.<U<D$6X'J
PC>(;5AH_BL(LZ(!T.Q608!K>L!(X*\_6ZIMOC"0($JX[4PP_>KI0L9#M]S*S$-CU
P)O$\7P#$ (!'6A>@Z0?JJ%!DPHA=^;YG-VYV2_=]<K,$\Q+$6SBE=MQ-:-,%6HHY
P9[;7(=.N5UG-D7!AD))Q#V.S''&3ITN.X([K9W0XW^9Z/R9+O2(&K)[D3+DM(K:7
PF_NB0@V?K]4-77HB0C%^>LQ/F;M:49_'W*,T'<H#>?8Z7,I 0@SGN,-HNS^X22 O
PT^;:M?HG!UHT(</<=NLYW^_J=IU_NV4HD&LO#U/LVJ<Q4&J0#J#X_0R<U!N9?Q 0
P@Y&]?!&9/T3Y8\M7-)9-$WG TZUL*N32L?W8T%0MC';-0,ER/]._]M6Z))E'BJ5I
P9_FR6<NPQY@)*'XR!^9)UL"8P^QTQ&_4'%M<K8Y;/7S*V%I>X:V W6__87'"779 
P/A:EMJWI@1K(92@U%A8.P6T5<B9E4Y"V(J6_I8V^/?2C:N_OC "]3AJ!3L;&Y([[
PD:(80K$[Q,[]PGM;(T20/L('WG[^5XTO;NV]&P("]OZ1T$1E( "!O9HDV%G*8;%D
P,@E Q01QL.9V0_%F[D>)B[I:OBWK74D1.-4HV0.:Y+@K"1*_KYP*^,$/&FUN9>18
PQWA6H8'.K\9![)N@5.26Q#L/;.76.%N(H8F<[[K94K @&1>K1+66$K  A?SU*UYP
PR?ZF.CY*M[B;/1%FRUZ3!@H7MH6WO(O+XT+Q'O#HH;Z$"L0$DB/=5B1A.'\W<^S!
P^S/L(U3@G9F:%8]R0J1.!J,2?4\= /;D)T?G>G7XSN#S>20&K"E$;#AKV*$,&KX^
P2%NUJX@W<8IZWY1$W\M1?K71G(/7Z;.MBV5TJIY[XH #AF'IA/N9$NU^M*$<D6/A
P&0Q%^Y5%SBCY.L=UW1\1E^QD)%%T#)8TMS*ZLVS'J_TJ*HLD(UFSVCS0!HC9]HD(
P[FQFM7$)Y;B@K3W__D*^:(X7 KT68&**N7!U%W\ ++H%*4#@H3Y*0(<9700<:TW,
P+PT@^FF[Z==,55U<>+/@MRH=\MNX"B<,-[7NL<-$E?6RZ\B?DHQ7WWB&XDA)?D5I
P85 9]V*1"#^#*.Z8&JJ)0)7L%A &Y!.AP16,/ZA@X^!S$P0"U\[_/G<1)S9?"N<*
P]>R>K@2+C6=X:;"#^F*U:/J'YIA5P5-H[5TY/R>V%6C5T,K_67+D.*5=,K9L7F64
PZ/!\RZY"J@\=]NB$,1TX1V(+WP01?V[Q>H.VLI*+*(&DW[K,H,M*24NZ,^;'\6;O
PJ?OUN\7A^1>#3"$"F21^:'#NUER, ZY=??3*L[#978,I.,A_;BN+3[02?@G9"I%&
P[F 6=/*5L"['^-9$<YBV%Z&$"Y:W4N4Q+7)Z]"7T#M#(\!,J^%5=%)2+E>X#?3('
PLEM^]\FU?C03""'XIS3BVT)%&^7F$6V9YSW747\T5,T;%5MJTIB(7-SUQZLUV/?;
P[4458WRI_*$\INZ_UBKIB)]Q1#:X%60TWZRT7^70?+@T^XOLY0E?OWPQ3,'&<=+!
P()S8QXN<#I<IQC7(VB^4RGAJ!?$TZ@^^SSR;4Q'POY8_&HP#SVV49 !V>SAM#Y-)
PZ2EF#OV.YZMO&M*2^0:AZ$6;ES@;'P?P$S(=R^LWY'OK,OL)QS(+WEDL4-Z%[D;?
P4X L7=<_Y_,C<=;S4'@$!H.TGJL5'X)T-[.?KZ71$RBM/UZ6B4XI^I H[8+]Q18D
PK9"C!62])O#.P9N9N$)B!X7J"]L@NN\E[JZ4^6=G4(YDXD0,)S=>47P-3R.(%Y],
P51,-CC@%5^/(V#1KRMA:NG^YKPFD.2S4?O?FRJ4)GV;(88K2<066TFQGTYAD=Q0&
PFJ;<L28^PZ^:+WJNM#LZKIZ_?1CHT)43<J=446D 4'@IBJ%:UCHG72TXQ>J%1V:]
PA:Y-_@X" XJJE77A?E'Y=3,(Y.^<,=Y>UA+>[_2S';#63IC;NNWP@H#=G!'J)&07
P=R+VK]ZJ%4[ZAG.OELR&IN+-*A](9ALE3AUG1%47["RCL<I8$K&4K8#I)T&':AA3
P7;ZCKM3A!).X83:%M6[>M?2E[+LO+(%JX#'/QTIOEE-ID^>A(('/9C!J(",&(&ST
P:")EYWD"4T4FWRM=F#2X;,<:0X9\^:/E)I^]@&=ZGB0B %5R,_L0HDRHMJF1I?L'
P[[U&R)0CCS3=AR*N''*X\>E*LP9E3]EGC+M,'YB<RB69>@ TGA,P:(O@]X]7K HT
P/A<&7-?%W@&63-6(%3/'O"$6+9B'F*1CK@6U-%-;#UW%J!5\W-5>$C'S4=)QF:<M
PAH/I2BY+U>3#XZ;HQ"45!;&XOP('4!F<B+<E?P>)51/GLA@".KI!T<;@C;FQ H>M
PT;M;:G6-]LDI/"JJ=K"BD6SZC^MT%5[P;EWIHDYY&4;)(,(:=\DEMZS><1[^R=MF
P(N-"R5>#+IE/>R"#_^J#[9< 5K^P</"?#F7[=_'<!M4+OY\;GQAO.U!(0_7Z2\Z6
P;7:!3Z(Y>T^(PDH\=\O#4C&^%GCFLVJ[J^.TU>TIXR9EA1YX&AP%XSX$8)YGH,$]
PZ8(F*]/4XU*.P6;/'6A.Q! 8/:X$),!&;JJWYZG$*\]XZ)N<$>D@8ML;#"&9BI%Y
P+5319.%QG?]Z"<GXJ678CG(P(&$<,,J^M,.543>QTZX114VSW13*M9& M%JP.DEN
PR<.(R HF,Q'@"VU"765'%\=\-.S?@D!47;+<\#)Y;)D=KC(2^# M3$CN-H<\3GSY
P'A!I3$M(G+;D;/]A;'E%%'.G)4E@<49@YGX+FTQQ'T) :(2D9PXQ;;<:REPPMX<(
P1T#;>G(TY%@KY (S>HA@<Q7I.RHQ@C]+94@3+6D'S[K=: #S_:]^(%ZM_['_LE78
PKXI;14W]1$[G%_1X#3(Q1UNJ$AS^OB^D?68=Z[2=0?TW#$(>O?A7;Y\?/MU-;FG$
P4:H8-%8::V8.GTBC#CB H$)6JD G%;1=OB-+TV\#,3N7<F7"?>] ]K F0272*83J
PJQ@B'@1I5-64J&(I;R[0J_%HN[#5.;=E0[S_+E9-,[L#'1TC@\VPN5AMNID"CG>!
P"%$D]@[IL&U&:"6M9"<U"8>F@04(_S.G /D,N0FE SD]1_J+F"T.VETR72L'*U^<
P79W?Q6K#[R?RSM<62DRH8"M*UQ";\ZE!RQ3]V>UG0S$MQ8&3$:0= FPV4$-$ JX%
P<RCK=&@F2HEH?*M85L(%]N_> "FQ,G-Z'Q1F.F)2S\(G? ,FNHCKVUNN*H]9I2?)
P ;OA;O"R7YI>=9W/H1(/Z-E$YRE_Z!8- <[)Q^*(+V0P*J4^!OX9R:&8ZJMA0$1(
P6>7.?:\6J8+RX-(&AO@S[0J;&A3*QX/?;<UC";L +LJJY$*JA980-65@;H79ME@4
P@=DB,4Z<7"!FKWI[RS(]%%ZG.CS"F7!DWYY*2$18@<$;G5]Q=VKF2OL1  ,+!;N*
P5GO"ZY:OJ'QPJ+FF9X6>06-D[@2,&?I \@G=$5I\&F)8]/=E!LR148%8PQJ#_A4A
PW9VFI=QM<N/0^N,=?2CU@&$OT .#1?N3W<_6C5%;/H=P\)_P!<&S#(U[HU+QF!)6
P-D9+*43+7(:XRBW?$2O\H,-&M4U0M#\H!'9JZN1OJ"'2@8Y>V?2)3:_?E. RR9?P
P/H?:G">4?F?.@8!T=W(--W2]\*C!G;@>@E"BAX8!T5#2].&6_K)^V^# SR%F/0_,
PDG^O%JE9WQA)&K5=W23U &WP38D'1 PLB)JTPM/_J/1F+D3M%$/A,)T%RQ_<G@Z7
PY(B:(Z/!-$.X4"D*](;JY>I\?DI"V_(8&B)C#(I6JE1GPV,K5"]3=<BJ*-3;&PXB
P+F@V[;4!0],.]'+,?U"X++2 B16>IHP(7:YF6;L\=H0_6/&!B;^Y WAK4,IY<U/K
PL/$0D\6_",8$=8,*@3=+0#<R+1_K780X5$#U'5M^TPD=IB,,04W=X JO<N0/W.CK
PQ8O\&&JE[>8E1()J^ $$HBH+241%BE*'IN2@ER2. ]GB9>ITGAD M3\9%0SASK5+
PW_U06Z#_]'HUA=0!8-"IN8OB%2-8'6)]#&6N^PR1$XIJ./#1!22JBRD;(H@83C:F
PB!^QH@:M)CMU%[GN>&]ZJ K^.4+E=&PJQ[1CXY<= (X>P1EL0\];NFR#HM@8^W.S
PD2+3H7B>9]; 8@YU3'9K3-=^(-4<7IQ!F:(WZ0<'+$-$1U/S;VF)10T2O%A!;RTB
PX=G\V_ :(Q\ N1)':&9_99OB-XCN"16*%2*M<NE</ZIQ)0%1"0XFUN+\!:;\<NCZ
P3'\,-;FNSA2"&97][3 *,-Q.N+Y2$R0^!_<7L,8Q.,O8]>0TOR0V&1HO !4\CBV>
P:6[M]V;NILFA5<LHK>%H]ZX+:U_6GC-@:V )]RP\QAC6?EVP^R7*7>$D3$_L+12A
P=(LEIP#=@)?V)=)J>JBHHN%FK6FUD,]_._KY2.7UX7FJ//T5LN;\G]9E'.FK_XM4
P54#$5LLKTPKJQ=9^609."G#\/.PI_PC\#8BE_?FA6]'O;1CB> K50L;R#,A<U\=_
PN\,D?TZCG*EV#J7*R^^MJ/S]E#\(]#TD%V5IX[:A+(@FB!)XY]<G!K^2$55J<W@6
P8D?4W>TF4DZGM5\  K*9_69I+QI7K*:M=D6G,)J.BFO!BZ?'.S94A;N5L!"Q)<'/
P)NT4BY-FC[%-2@=)]=G(;+.@Z(O5D,M[;3RYS8HK1?#Y#>0A%[+$(#JP-6%0<!AU
P1Y=M>L@WII!1<&GG(Y9B21Q1%K.XR9%J<,^\]#@&JYL>W"E+!:(V[YZ<S1;TP6#6
P=\9C YFVG*N[&EQJ@-H:6[$(Z8V0%=$5YW%C2AG7#9@>)IL,X=$ -<"=%&RW406O
P/DQ:^$Y_=%M1L938E!=!VR'!H/FDQEOBI\K#:6M.<:)L=%NT2%AO1HV$,GB9$YA<
PK?^Q-1[U;<J0"O/<\N@1,F#B]Z6%XD4PC6^^5J.BCBI>]=!/D3B^-"+D1Q'I2>7@
PO%J.W_)^!?J2H[69A0WZ5C^V)M% 1[ UOM2GY&7WX$Y77GWWZC'O]_ZI+CY(W1N;
PKM,*@A3SO,R% X37E#M)-2T-P9L"BV;=AR^S3Y!-V9NSFECM#.P>Z4,P949(6!&4
PU;;"*E*2%^"2R>X :5<J\Y[I@T^W:=3AA,LK.U".*D7LGA4;%&OG@L%Y.7ZS8WG_
PZ-=9W-;0#+'05G[+B7ELYX?(MH1K(=;*6K0]+((VD&XNN"J-67#?<_WY+]KN!?"A
P,G[M2G.0GQ?>:0(\-_V;=;J?(I7QQ\LXW'ZG^R.=_D,I:L]YM/$/"'PI9W4#=C:3
PI0V,>UB^&76HZ!,WP-%:(MB_OY*]/9('05!0>+Y-8WQEH"C$-5DZ"TZ1J[M7  [R
P';0!^+-WRA[+TNYXOCG?&\55D8FL!&Z]R?B76Q854([XP4VH]+FP<CW35,'+MGK^
P#]EGNTY'>@Q7OYZYH3>!&R17-,>LF:)6?R,A@T7;8"!NF.@<)$6__P^ ZL/WL1-+
PVZAM7R'(BCY7HA+M]@Y<(0O;)C<AQ!-B(A&$6F[*-Z6EM>C<Y#U)@(12>J/@>"^O
P:LE+;RAK13N]UMB;>ONBE*6RA#WN,) ]_>RCX+'OZ8+"*GA%F<C-P9KA(,U8B,$:
PZC@BR'(2E0I*Z"ES8PZ2[F.19E052<C=3(Y*X_K3?<H<F5Y+5;)WL%*?"+"X2<TA
PIF^?&;/48X"7"O*4^Y7#A%$BY9[KAG>!>Y/E4&-9]0]%P)<4CJ' => %JUP2-4U5
PK>S[J5A !6IY7B,(%7(=\5@L@;I^#U-B+^Z?"64LSSLV(3I-IO:"6$DDW**=K,[;
P_IB>-QU1\)L-C*4Z3"'/1:0%)H,S,@^1JH,'/N:M@L(N<0R GRHL("W(S+>=/JL7
P@2:/7IV*J;D2911"R"\+C'&YE<=F7"Y>66-2Z^U #/<;&=VZ* ^%QV1(I]<TFXR#
P1\#,-_'HB5MTR'J8G)3(\D ,:L:KN@TX* "X@])B'&JH/W6'\"8DE.I33SVH/@GN
P\2JR_F>^\/Z@W[UL$@/RU7%:X5O&6RG/[/&I8HL-@/#'S2Z2%O^52:^GMD8G2/T4
PATZVTJ.XL;44!U],HR(IWOIXJ^^"4NF/X1]\H9$'2?C&.0LDKR(HYCB-3DYDY9[<
P3ZRQ?GB2%>8> 7MM(%99HB:?*XMG95".PYF0^Z R#>8MW$,/W#M),2GFAI+0[RQ'
PC).EKFE)*HW6L!;[>6872Z4L;%%CQ].9OBF],8ANIT FD+Z^Q"8P!R$^QE/>PYEY
P5!!=!4SSZ;%ZIT.7650LF(*L\D)\8WNG$=)W)Z^H!NVU5@V=E+H)4EI#517S6@US
PU2D/V)12=>;V0I>_%>XK5;"L]#?W*]N-LM&8-@=4J" S.'TH#=.$R.)MXZDL $=V
P2?^]#[Q!N/@(NIGQ35<'/C1Y@LRB<_@G\]+3DT_C6>'%'D8P:E_5#*8]TS^H+FH]
P;A++!^,T=(44,3(A?%L3@6LV4L16VA#';-E\*+86&\R;!.B*Z"?FV (WP+_?22Q#
PJ @V#6[H\Y%*<"FEYR#+5H7,=CJL%9D=8:)K,?Q=BYI[W:<SN==)AB&0;<9%.D@K
P#D+-FXB>DS$-1G./\&[SOG[ '8]S5(#"\"M+;(A=GM*-;\_IS]QU(SE(_*F";#Y*
PF1X;D1;ACBW%<[H279Z)22/'GT"IY>6Q"T8O"MEQM0#5_6^;'LS:+;VR?B%ACEB(
P5\'3_7'@^SO02!\QH1\$:Y'*DP[!4#B.X=6.*Z,E_.C2B:>MT.3SX@$!>H^*P'9+
PG<ZJ#UK@8/QB\7LSDC!)E06V?Q%; QH#OR\E\&ME$B4P0T[MOMKMK&EAH.A*88Z1
P>!VK]#XN3./01&-/NEH8<+YO'$(M#.R+:$Z AD_IXS1+UD>W,V2]KE[M*%K:J]-;
P9M49)GMTEBR.)E.]J4^V>4M!A0O2X^\' \HB_[0.$F[)XX%ZLO:[S)0O+M6Y^;>5
PJC&<<CE_AHQ&$LRPE:)$(J<154W!Y5+_<G )LC"=[VN!A56!>^3HC(MNZ,D-P88_
PW,_;V*&;XR@A@3*WYQ:#JFYWH/;!2*QR?9I=^-,I>/G7)ZAU42M!G^6C; NXL-9J
PXJPJ"1FF+7(04DB'SAMN-"Y?0;4H>X$B%21L8YN]\B0'"W.P!GV0C^?Y.G0SH?5W
PW XNASWASWX679G&9YEDXXW='UT=ZR)4H_YZZK1P(R+T(YN?^%0<IG[[?-6X.@M8
P.V1%/](M$O[WE#6%K9@@8Y^GO_$GT&])K=L^[!-@_I3DUVR= =ZRU_ENN;#U06BW
P>2E(?K0O(IBBV,W_H:;/>Q471H6V?89(LB\ 1]0,L])M-5/A0  /;F_SKV:CF>\&
P[[&J.F8L.;N*(PX)!'-]/2S[B.<UEETXDXE9K&=:YF;L/89^.Z&#?AIUN&0 #FQU
PASJ.UPPN@\,[?/73/CV*K99WBG,]]<]#GGTP$$;Q^]_:]_:J)VH5$/:(K:- 0 32
P>76D$&5*HB4%;_RE\ZDM!^G99H$;.QV=OG>Z#\T^L?6<O^H/C) HKSJ1_QS=BXK 
PU,YE7=0X4'W1TB%05@!=C\XA^74^-A-87@Y.GY/Q]H?KI?$_*.F^8NY8WEDW\DE0
P"7P!-XT5$(M\25HWS;$>SB2*F'1E8N\I>XE!A90X4PL[X1PF&^OF2QS4Q79R"WSZ
PS39'HMOYJC?W<OXKJEVM>'C-2"RGBJI&C\ 1@BYT3%X2<JO"G_*-DP40*BG0GJ>!
P_GO$;;18Y7?C&VG<=4/^LTH&EW%<UOLGL('/#;;76;6X*S]0*C<3IRNS_,<)!HZ#
PX4 *I>\LV$H!R>E.,>KLE\0:E?=KCW)  ?$ C4R.]$E/3)Z>H9\YTZUW'%D9JK'*
PJ);_1LTTA??'X<=PB+G3 Q7Z\([H1?,VC^.Q>%L1^9+Z8'S_\-:2U86KX662BN:^
PHVH2Y64?A&<W%7(EO%_M7WK$OU)O\QFB2\-7+_E[EZ9^=OF29@(K'3+F"#)AWU+%
P3R2GUPEE5D$JX="$9$*^>N&KYP))8E6;$'CH3 \G@0MI>**0FS'\74+&*)7OSBBL
PK%M*#/!6?#4G'FIG6DW.^D"&XW8P6LC>G0@R\=#;T04*'BDK^^\8J!O17(U80$/E
PL/[@/]+EC\^SBUW XV\\L&$G=]GZVHP9,A<)]D7+"IO5_$Q";E7&)NIG-"&:CCOE
P0_I9T2SSTNL4,X@1>DX1BNEX,&O0<&QL@@V.TGK%M]JX2,;_ C,\ZU9Y>JA*4))#
PTQHL224-"BSDRHC>6&(S*2+BV>?&8 (KNH!06:R$1?BS[Q<59 *B(F&%NBET[R)"
P"9\>L295$#Q)<S7TZ^-H?S@RK##(>9Q<EV .7\\+^ZAY9PK24<A&B"M$KOMBA7>_
P]-AOY<-,YYI9V&(*../"@Q)Q%'+QPZ^J!>[GI>&K4K1GG:!,Z]]D@5&QKZ,VB>? 
P1D?:JV'D9-F6+UG6YC]GQ(#52S$__1.JO!S6OJY4",[V5^[(ZZ0:/+>%U-*EE$_H
PR1XBRZ2RY"'T:V),!&:AU. &_4BE*G?>0HR2M:E:J[CSBS<F0R/2U:?GM8'B8(O^
PK'7Q('T,Y,2_Z7F7)N)[M05,,%!]+NYY_NFCM;,(8+1%GH].(LB\W!(I@8?8CKA>
P<2@HL2#G7XR^ RDM?)S4>VU?IU+O#3!70>?RKJYQ=R8RTY9%R6UOV;^B;T6&+;3%
PD.U 9.L+TOS$O 7O$_MFM+6=/O8YI.S'-7)T9VR!?&\(_"H_IL+Y1X00QI2CG ^E
P(BH9R1W>O)$:['JG4:6S\[]*_A6*Y"]$$63F.!1S4"=^D0L?Q4/!Z5%+2!L>X"$*
P[:\2N@>P((2,YS6K'!"CNO+>F]BQFF?>TDA[$A8JMP>Q.FBEV3H_!Q)A?WSZ5Q=V
P$'\LA>65B8326IE)=712W:RTP#9P8J82:$T^8^'<P6-N:M1ST-KZX\;AA@]XW#4:
P^[0EU_T(8N(9(R/>2\?]4/TL<BI$2BOR$-/^D.^J$5<7?6<EHU;V'3#THE^*92:)
P9RQQV&<B SI>QL'3&K@ZP[N:_'.I(A[VH5.O59;%+ME]+L&[4?S1QSVO<5Y?R600
P\62:>.FRGL4)SDG1'?D Q+R'1P'C(=^$'CL5_R[9'=<U2W^K]2H^_:5PBP0V&TH=
PO027'/5A[U-WC<1<Y:;:H52H[K?S3[^X/>V?*D1LQ1R@)%:UXW2!8T5(+1*NL3\ 
PK;#Y2.+RY!F46]+^6Z^@,L$W#1$_74@BLRNMXDA M(;2P&J?2?2K069COZ/(L^ .
P2JA16WV-LH>CRE2HK[2Z-5ME46WN8TJB%O05Q(%TL&KJK6:BQX+.Y9(K.T<(&^PH
PTX615)S=?!SNF06,N]N^\:]@41UJ-#(*C0%L$.\\:V3+,0.]AK=P?AO"D]5RP,^B
PUV*8?RV!3MN,TC6.J&KKO!V-QI#OZLII3B(.E$"D2FN4)KL6)Q,$H\+]_!\M;@[5
P6<L\[>":-)B')'1%(2GV-'PN%#,A$AAQJR/'G9J3?I7U@6\!0@_&"+5U7*=4?98]
P(?FG"1;:G&$RM2?T\?UE>RO]!HU%R=#09GYA+XJ@#-:(0TN,N/9*7(B75, <CZ)D
P6SB_)PW"*:?9M3_IIG\NH,,VI]O_N)#T0-^B(:!Z^/6"=M\<C0W<9X+8D>S[=Y:N
P7F<]K29%K=@'-\R%A@R37XP/6]L7J+%72O-0GYU/7(Q_/WVNN0A00R!I5X7]71#K
PV9&W)?435PLVS N#+T\8&57N7??*Z.7![85&E_W;5@]K-3(BK4^3JGEL ]1TW!T*
PI06?1E,BK:JI[E,35RD>Z&<Z:^E3\T=Z6/95'$H&GM:ID5A-W]3=:)/!UIK*MVUM
P,]UBT5[=@_:TVGJ\U(W!2MIGP5;O_&C3]%SJ6 L![M%W(YOJVLG0E@RAZ?'U&,Z#
P1X[\!KN'G*EY2;EYW*)$^@A'._E+/X=YP!"[G"!/649N'1;@X<H0IR$ZK*];(<E*
P97LIM^Y<1N-?,PZ''5[O($E";3?+M0NU%$F3D>_;?"'D]/J!.E/\KH+X(6+">Z!=
P]5T='E;1:. NP22;,#O82DA$8>G3/@JLK:&V/5\.<1'"PR!_SSV P5B)WU( IH<@
PS.?^H.QVM==,GY(Z#+L<T-XS54$USYQ;T9%0BT!V]'5@W@T#2X@95+U"_62KCKDY
PI>$''<>6_[O/*#B/V68ES8E__:<2^W2J;D%V\< +O4U&%L"(9<*,I>VL-:/IOXF)
PK G#^FD97DCN7FS#:$QJSXA+BG"2']$[JNFQ;>V[ZI^FZ=.WOFG!'I8G;-;@CY?;
PZ.>12NZ>Z)F*F44W\7Q)Q]A:CJ^I@3"P?0<1@_.GO'904OT+^%JPK[:M&]JO"?9H
P\'1G47&ZQR:QG]%9\R]]2B3=V3M-4H6BH&C"(-S(33$7K=Q3OIJF<[7=8(R%:5!;
P[$5:Z<"'_19:7*.4JN!DI3MLP?IRJZ+](N1)_622E0\90;LT8*7)1'SNT_D)ZFGO
PJ$J;=/'89V^5E3.TZ^I@-KK SB_].XKK>J]H<^4_A>$6WB150%UZK4>3DF'>RSH3
P,]UL]4>6&N<-&YA29.U?)5C\R-]B0DFR)W E"[-K1EJM[?"6K22BAW;9:Z;)V<2N
PT=M6*UVJQ2)F&*0 X:1RF?O%+YOTF+I,87-C4?KPFC5FGMNDT_;A-@46\VI?[\-^
PV/#0PM7L_! $A>LEN[C07N4ZRYC%2?Z=_I[(RU?)C#B:IZZBE81SR++ZD&K.4@#C
P5B3S$>N^S2#*M7S<N='_]L"P6T]M?Z^1Q_ ":.-9_'?CZRIKM!/[R<AZTC2H'Q"^
PRA^G$YXU,#2OX.1OZNG@,QP(M.!9U.%.X>S?'-K_P_A3@L; %T2;.FV9D((\HX%A
P7XRN*?U: M-=9"D]P*K&T7 X],<8;#]Z&!^X"1>P-]RW1N]CK>9>0\J@NC/5\[3-
P)J4G0]J-&I>_9VCHFRB[0)L1FKY/ /)?:=$112)&$@D#OSJNJ&%5"7K!&6$P$:/%
PP >UE3PO]4)M90VX8A,POCB\M.7(O6\3'/26?B=ELY/TM+J)1OG':@SG.)>OT.EN
PN9#$\@H0!7"A17B45,]*D_!0I1B1:&6B\Q+<\*CT%K^RX4WL2KQA)<8&DT\!D-)F
P0^%'367,-/=G. Y->]$:STM$?NO:Y/[ &\EQ@L;@M!90(XAJZB(A11^M3L1=4K':
PZ1G(]T"*+P#S-G,3QT39Y6B!8NQ'[%I9:/,I ?X/]6"ZP?&I'+F$NHU7*4-UVC3B
P-U]0Z^-DVJX=3MCA"_Q'_O9DY-KK#P^"<HY2]_#[7@]#=,%$#CY89+T0E$2Z6=;K
P0"PZOPD0(=XN$'_NK(<** &Y'E(P3IJG]>U^4SG1.D]P&$5:H^-F:CI$_[)=<HI$
P"'400[L<7@ )]T#[.P)1R]^UN'=Y+2U L71]N(:(&U1-<#06,S9G)@1*)ATR$M(1
P[)W$Z^\FBJ._)!@UG"/[S'@8%6 #YJPEAI0X-9,.XW)^PIO.EN=\ $10(@D"+Y>E
P(7CN8D8-[EO'QQU5;D15!XKM(S31L%/:**B9]HTEU4Q3/!K[DCNAU\XF4Z'^5>D8
P5?[$6=PYC29'4%^UK(XU R%L4UCD+E5!]R#LHR/ 6;/?KMPV2(+FIF_\+DZ.^$%0
PD047R]F';#],D\$ /[L%65\%;<<6AKV+4F1&+3+6137H==R6B5^">.4U%V-KKR&(
P\(XA!TK4Y>HDEUX1*1XDT1![_I\D6+<(DF5I>%KT!C*_IWRWO;$LZ/VV=QR6%=*A
P:<JLWZT\G2'-QQZNV.]3*#[;?=4J0[>U"\#?I&W^&17IE37#DZJD%F4CO=V'M)Y]
P1HSJQ/DNE;Z#*3I8NT$1ZM^I=ZZRT:<PH#7K))DHG$\2;R+LHT6(FH;#HDZ2M"R)
PX.A1XK!,ELS8D9J4?&,,!(QWPT^.&2P1-X@'HA*(?S;N4$06(>=(+A\]R,R=,@8^
P%*HYEDZ7<[V:.J CGJ^](@+MTF1+D?O@H%"BC!7HW:Y'\"1$"9A@%_(]]I^]ZN#(
P 75-_/D<OTZ%OK-9-?*GBP$B\"'"AV@+&D&40U#G4<=/9,5W$,2]!HP"X$KUND[(
P$8I[RK(M_'0,;0*8[Z/$FO4J;.']DAET^!/LDW!076]VA=Q7+ WYPZ[>%CT3B!]]
P_XT\@N8+?UI/U6*-']C[I#B5_E)Q+YDUW.JK9C^7,TU]>!KKZ08)'H='#FSFV-"#
PVS_T0J#K5]G2)1^ (0#CTG4B!DDL[08.RJXKY)(+5.>=J?97' #UY!5<F$M;=[=/
P'^12/@0(G<J M'\PKH%:'O"'ZH22FA)K;SL/+A<V8U@D^*+?/Y'I$=6EP[3Z85F$
PR=W3_YKIRS#$6N#"Q%ZIZB%A[.+N"#<?3T"0A ?8P*0^Z;6%6%8M]=?>;M7QP$!*
PQ#WCFMV5*.90 =V3JH)2CMM/ >$.8OT]AR(8&'8$4C' +(1?"XU79"5.:DBAV$BZ
PR+5>9CYJ:)P1CFDSK 3M!;[UGM8\9S;IY;%PSPQG>V7(O<,N,@HTJ */EC/OSA/F
P()J.3]GBO1*;KN-!'A&VTKL76<$X(M%E21XQ,M_;@-+'V =GH940MB#G(0>/HK^V
PR 7#F8/ZP]T>1^7;]-07D>'A,WH#A:E*N/)03UIKCW72?B7IBG&^]/I%4Z''40_(
P'I;R0C0>^G-XRRV_*X#@2B#SO0B4X]RJ?7,Q)[>2-C:&(:9:$S^XSTJF2,^N%T\+
PR_8'ESBPM[&D?[,E$_B>FY,H#A9MAQ6]H!85.Q5,3:+6+&K3=*S4]X7A3\F/",I>
PI9PPRBJG,N>;L)S9_8LS8$Y/LCAXM=Q738>-4>;CP=>7@V<<!\)GT?MF&I@)YF9>
P%[<%.B948;<[?9UC3L88I *WH<-G7GMSBX?D^]XH^I.CEZFE(KAN-'5>-(+[K?OT
PNU:7K\/= >L" _Y^3T"=<EF=?]'I,]Z2TWD'Z(+8?5$7ZMM^#%(37EC:)UQYU,V*
PJ9TS05NRA4PAACFYLH%&B\DB[&K1:1?1W5AUBT 6JW)H.0,T&R0+<,!GYO?XLWY&
PY]EDY5?%1W :['%_1V&Z_#QI0R"C L87&Y\5U9AT')=Q4T2%ZK8;2M\(DDTIP5OV
PRT^S4J'RV__8FGB0;@-;8]QC<XK0E"XVL[H;_J@HY/L=]W7-.>OCU_/2!:XAWG])
P5>B >HWY%S%IT-WN6/:TD>$^.MY'8 #PS*!O\7E'4.7<6M<&(W/UJW*K;\XE3V%%
P>!=EDKX>;O^IWD5E2@\!>UC1+WDJ(2!MG"'U@QN/F(S;:8AP,U>,5S)P/JR^P*OF
P1X'F38P\BO1_IZHO8=S\'YHB(7&NH;,)2LSRLD9J+$%0.&XBNQ&&^-?\Q"Y1(.' 
P8LQPZ MG<H\!B-T\<G(Z5S#;\_10?'$Y!GI:>>Y<L?_[+A;,;A&+[6?!%;/3_;MC
P-WASG%8;:K[@T$3L[!:9>6S4.'DO,U?(TF9;TGBN(FX(&RY@:'T-5<<^;]61S&'F
P]33G_U_1AE]N*&*9]1NX@+=;C@-1-@6MC165 ICI"ZN\A".?4N%C(3"EN*R.@[K/
P;[+PE &UG)$]<P=_V^PW^HMX1A<\D&C/)):3V"\,$_WG:8.QV[?,9E#J@*I&5UW]
P[-#3A*_2?=W< ;J "B8+]+1@2[4PM):OF#/1J,^SCSV(I"F-,0V(1Z"I GDTJW"T
P"8W+)K#T=NW1(-#&,L1JQ[6 TTR7$IUMOE:T *R6MZB0@7U\A=!8W9U&J"Q@F'_V
P5JO:^X3J";8?#31%/4)#-$V\>V$<888^T./69KKU5V"Y$'>VN\<]!1G=&,SGA/ ?
P^'B[F^?3MR,_PQ_>$&1UJ^)H!D4D<(K7XKW2OJD*3)B[LY:N?,06*5!94'GG80*W
PFYM0W8M. ALB8A\7481-:%C*"Q3@E4!V^I_+3?$R^"T+)S(.2O[U]T:VRC&0"H7%
P-5L,[JR'>OM5J;X4Z]\,B> 9?)JRF*^A257;1,&VUR>V5C=?X36&U\D1ET@HVSOI
PE?XK-*400)(H+9HQI9KL_4S95B*.?1I.XU)89N2>^ST(H2"P3<9+'0DY':).%$. 
PIS^,/1E)NU3NJ+NW0MKX*-40.W:CAD.D,D3L+5O/W@O+G<IP/;A.:E\JANRS\;,P
P XI(&6O1_[W@EG-9<T N;O;Y[^P&R4O%JX>6[^FJ[,^FS2(]$]F2EQ)+BB(J_$!M
P O;*3UG]D+@-]O%LOE[D'<4R6=3SIP>N?>+(ROB(N S[:ZOX:?Y*7OVV-&T%A3UT
P U:XP-2_ -N,I9B!NF4GNH1S_I;1O8OU4K8Q\D[YZFUD0WK $IDQ#L3)()(XP$IL
P\8%&-K_E'Y3N%M5\XG:0N9W1_NI.Q]Y,^P:8Y:,1,JI$PJN<<7BYV#,!I%4]BQY[
PM$E,E_1OX&N/&=9%_JYN+I),'[FJWIF5AW+#OXZ^"Z<#%V4,,FEZTWY._75@;6U 
PT2+=*I*D0 HV 91?/$UP4)/[VC\-L )"N'"]YY(1C[EO^4\IFB%#L6B;T0PQ.=,0
P7&2)D[90#'--:Q :+8OSOM':"PYN9"X8U:'$8QRM9+._X35E>8G(3G^+)/^7%>!\
P(K9TWH&V@CJI6J'8F?^HXTNU;^? Q7L1X8?_._>PFE*$!]?K'%2@YF#IWIA=*#K 
P13CY380;)U_:*<6!=ALU!IU/SK!-\UKMAQ9-ST0.2ZZ>U]03L+7/WP4"& \]0 @W
P"#VJZ10%=BQ4O1QG(ZNXLDXL355I0?2TO<ZC#/2L&G9V[^17A]GS91W[!?HH.)51
P4M2>&Z[%"DWU1([R0UQMF_C0[RR*I!787?(::WE4MD[7.3M)7$W?/W2M2\Q]TV;0
P?=IY_#O:.!IAX?,2-#LN- "ALKUK;,P4KAT6#=R0+(-+958RSF="1WI+L,2BS4&@
PRN=3\1?_9B=:>F%_7.1269>C*QLAN)V?0XW8G=ES44T=N'YTYC8*][1CP,W)DQ[R
P^UOMI6K$CR#A-;/_FK08ZWO+FOC/7;P2Z]QW1>.J:HW0]7)_*H$'X&X0[?\Y;T:+
P"1VRA%M]@A[)O<@N#NS<-Y1],&\O%+[?+&N*;'[X9Y25QWXB?L,368<C</O2%&ML
P@E.VZNNU+]];@R\>.\5-F)A>OWS'J E=3Y]^ICLVT0GS"UUGXA?8!0VHA-DO:-GZ
P; Z[DZ&_E^_78Q0XJ( =74*)NM'4R@H8B#G3KET]H;)FV/SYS^HK5M4:;?R%J*.U
P<_25Z<_HIN_$K,NY&44.UPRA84L^%E^27-$EN'X70G,*&E@X7W3:4"H8?QJP)5T^
P#O*>#D8'%<(72XD=EJN $'@4H\1NS)(PQ]X[E5I3BTPJ/V&G0EG!T.M&=0\SF68W
PZ6S,,2D0/M8.;[2XOZ2L8]F#1&P=U]/4,,?EF,FL=7:\]!TW#:M?.L"?RFYGGP#;
P*R6Q!'V/:R):$??[Q%R>T7:GLT*@M*7P7LX7Y$_^\TKV!H?^<2*S1L4$=P0II_Z*
P9A=FU5@*JF1PAM(-W:(%7Y4K]JSK6<074W+_;[P 6LC9;E]YP:3'F]17()VRE7 !
PZ2V]T"4)V:E7Z[J/3#8$?00E%RR7U6@V_Y"&51KCJT ]2[4G<HH+K+,4[=P(SJ3U
PL:+&/0*GDH_V0%K+.PK'0#GD^U_TW"WA/)^L]\6X9%/)%>S+\L;WZ1K$>W&C)':&
P\MW@'NU*X,O]S#A_0(<FMCA5>#_46?)R16-\&S LZL_8O,425*A#'#BA>!2M3TL^
P.=/WQ^09=2)-5,IG'T?L--=/-'@PMS"@7ZW-,ZH[:C]>7K>Y'"Q&>3L>D/%D '@H
PS81,F@@X68 6R<5C5]M4Z)DA0'>G8D5S-M*RX5S;GBY6!5AYJO'JU;:OF()%54E&
P%RE/>%[1[<!;"O,5M_%E?"T;64+\I\$DA7BHNFFNR_7QN6;Q?XI6'KM('?("C>N"
P;O5W8Z9A,/=K'+:5*9*N8$?M9;?V]+;6BO+/>;7B43#WW?<-$&OM@K-1]-/W[4R?
P!%H1).3:!UEYCD^X)MKOK92(,B!8+NBOQ244R+)1)3S'R]\EGW^Y&UXA_\:0'N2T
P/@ZKVKUY=3@E>>U$#6J&S.,8"P,DXW1Z<N]'SJXR.XW@"@2OMT3Z;W'5@;]95K>O
PH\.C"=..S=P0(JL>^"AY7LI CR[ )JY3&4YDL)<^QLO6L=2]LY&>?/Q)BKSRG6QI
PXA44)%_CL .+YC9EP=GMIJ1I4<?.2O:$]_-7S*AR4;B$B4]"\I=@D^[^6#@CRW_R
P)S5UV3<\1_0-CV.>?>G]](.4!99OC]#DU?DQ0WJV9D5&KWEC/SKP>,CP+PD:3VVH
PWQ> 0 %>H;'\4GQH127BKA[36VE/LO<,.FZV=@'NXZ+S?&!*CNS+ ^SKC-(S(3=-
P9?2+L8"O159U=#2M@L; ?#Q3F!-%B %Q+?@>4;)D<QVA[-E)OS2EM@&7*I@#WFK7
PR^TMX:6<:E!^QF^"_P8^:2D7JT<MZQII]]BGTH1U)Y+8N&S2XRN8>6%I7[_3ICJT
P:LT+#U:S3DL309K ?WI7Q]]GB<CO!+"GB) ;]D8%Y-)B-A(,28,5EFQ<NR1$4E.E
PR_X*^H<2)^.50-GT^7W:CM)9WF^$^.V!PX1E]UX$Y,YIT_E(:7Z'(^'6U=BAF;&*
P!R);K<4X>*<.B9ON22CH&T?ES2B7ZR?L&KR30,:_U#DJU".(#S/Q%"CY2N;'QF_N
P7_\(!L_0,I$)\&%RA\;K(#1XF%-$+:PFV+&Y>H%8>CVT*,#.*6["5,GI;)@A(&UJ
PH<JX-EJ!N'0I$<D.:-%KA!Q]^8:2;0.*2E#&F/JP]>)1+3NL5>IJ6)BL%?E4/'+9
P3J69M'=DXE/AB&TWIOCD$L112(=K#\IN5:@1C!VNN>SD+"$AI"/K;FUO/&^OM,ZG
P2T<GJ=/G2[LQC4A[&YES,?;W=1DP#F,([37M)("H_:,O8ZHO0)DR8KA-DN&'2>R>
P=^[JA4ICC?+"&Z(,$2Q'?VZP.@T=5Q6>L7^I/ZD%;&KO#GJ]6M[)5@ &Z(X_M9BW
P*0)R\@U"OD:+S+?!]+#EJ![W@VU/2\SS !?!SM35;9QU5$^='YAU'% 6?M;\// 5
P^&S-%\ 7O)]3)/[R#B;N)FF22L_D$V4= SKO\;:<>9B#6"-,-<2MI6;^\!>D,.3=
P^G%$6>:AED0RO)-+3;352Y+/[E3>V>\R0PCIA5V-U&::F(O2+"9L''BLY9L:IO=@
PS". ZY/R/6P"\21ZZ8=++AE7?59'( ?>L1OY3!!MWGK/B,[JMN&-U*/=-87K23X6
PX+L$=,19A4I>+K4$9YXAQ!E@DN[YI E;YR/8W7H0!ZNBD&YF(_:P."FZ*+3!"$7C
P\ P=80T[7#IR$V0/"C5TT216:]W%&N>>#H+JP%].0YED"!/DZRVU[@S>3]11Q2SE
PWL3.N6$-U!GI#B/"TWW1IH8;2H;S[3F)<*YRRV\LH4;*J4=9JH/K [6 C23$R7>%
PT>PETJAG3?(%:')M6NCHIKWO%4%@*8A">=MPO+VBA8J:J5*KI!\K!A"$ZV C/WN?
P/#S(96F5JO+[A6:F7<"32%IO=A1;'USG2ZUN>8KK0/WC,I<D,IS6B<"YMZNYHZIF
P%#J*G3@MXC2YK?^4P9W^=9I8M[?&/Y7K,]MI'#F0SJV[6H(@/V!&7)'SY[HH%!<3
PEG.[!7^<FZK+86K0G:G0+T'1Y.*S[Y0@I]M@7G4R1_7M!:-M\1SY.*9M1$5B$7BN
PV)SE,,5P&CG%_ W?(KI1V_$0WX-EPM2-)E-F*S<:VFX\^\^.;@N.D$NLT0/ K%[@
P>6YS;[QPUPH1I#H/6^\^40N/L1KV5#JFOR<_K&](C(KE4.YMY_4J200[*O!%XE<>
P]5%OT%HGA.&8%)$45J*;UM26B02SXUC+$:?0$1FC1E_)_XA0>)!H:&WLG::R9XZ#
P*G;WZ&-.:70?YN5S=SD:*XN8^P<C_(#6V>.I5I_DOQ*Y^D0V2W9%L\\2I>$-V'@G
P]"P=EF)3_>#9_\7<G@8\+N#@^<M@3)"B9IHS%3^HS;%$Q/B:YK=:5%G851I["!9N
P'VSK.DX!&?I=?J-Q";6R01<X7KV@:4(9X6)D_TAJ8*2PO/=Z!OO.YQE<.XVZ^8 E
PNFS,U&SJY:R4[3P_5 7SK9JC:\?I#T)5E7QX63EQ;@$>X@_&)L#9[5GWB19YIN"C
P@%)PKP(6%'^?9J0E8D"7@:&^KSP_?4/IP-NF,9ST5A7!8_0F(?+ >K1]P;^P5&C)
P@JU"B+!/_/+K0Z7EKFR=CC0< OYWX"/IS=ZB;M)*2[=GDZ>*E[43]]%(";"E2G+>
PU1Y]"G8?)SS@(<Z%ONK!AWP^36B$, ?5K"=Y'W[L&ZLEKI75F7Z>/!&+V;]BW$ J
P.I&!)O]O>LX89P"9\S<IXO<#6S .3"9"&HJZQ[@01W[Q3>3;;A&4]_K3XOBXT;QK
P-E?*WQ?9GEB_[H3IC\$N;\B2=>VV.OQ@Q"H!)%^](-QS"YVDEHM'AC!SQ!+X9AD8
P3TEX'TJ!G7N?+^0DM!04L)AL83W=_=-1%=[Q_:@BX =.(_JDF*!@%!^NE^YVW88:
PM<BR<MC$>\M" =#PF[#WNP.W<_RQ-^Y"\WSR7:K3AR73-,@L8V!=,3C<)E.4.[QA
PQ-<T4&*ZZHO/K<;\=!C0(+RAXKL L8+%>9S&5;8XI7<^T^UX2T^U?3MD=AJ;X;V"
PJZ&-U'D)00<H,1 6 %J@\"'[6(S=UJ)9S?O?L(=;I>2A_-S&/B97>%M;=((HL[TJ
P<I?SV3F;S.@B:_NAORJ)]REQW:+;.TLP#*_9E/5,$8-JIN9^UZ#,GP$P_3-5QZ8=
PWO;+)7/$S7X9=N%IB?28]_N0=;2'/JD\HY75X8BM,0:MOYS)/D<<]E"T!NZ&^9'@
P=L;C7WCUN$,C(U= %KC,AG.-AIBQOT#=SOF"BM-_8QS(+?MU?@ 3%+]^P>?LCTQI
P2B+'7M],[WG=!=&@$-:5I.'1;/GA]6HOA>H=70( S .R$H;%NS+E_0/\179!I'V,
P[V:'GN,@/)0@O&0]/M1G+CTE:,##Y#HG7F2K3OO([60)\FSD+S#"NX _:#77M0.V
P&7(C@$"%[6\W%D3>>>[CFI5VJ3YPG$]]XEY3@56'W3QOQ:VBPXWIZ-,P<C@:8G%G
PHB8^_-# )R@\!,'-L7"Q@YD5Z.X54EJ^+1& V@V)\-]_$B8I*^5-!1IVRVCT PZ3
PW]SD5ZYOX(UPCX83K^=2ESP@<IFU7KI.<I/)GM=V-/LGH<-3DB)G^V?G23V#FF)4
PVU]XW#(#7F,POW7++BMGYF0SK)[;CO^=Z,2ZQTZX^B^=V7E\FE1S"F7Y9PYV!!6Q
P0#%,=&Y;VK:QZ'A1?3^ORS2G$?T&O4,<OS1;,$22B$:A7DV_@G=U2B?<M)W_!$O!
PU(N3 H;A^E6'.[,<V!$M^@EDA"FPTNPJ!5*Y%&Q[B:9&<=/)@M7S<T/P:!_(E?0\
PDJ^^:%S9Q!&UE[-F=R+,HNT;D:@07XLIDID=?CXO56Z8!RQ4<;#+I*HR'HF--P*K
P\<;YM9&L&\-=Q;>3:;K=1%?V0,P%"PAX&IIFNP%>#=IWE3B26$T]0./U +C322NR
PCJ%F#Q4A-.\I?+!NRX8[D0C6UXMUG4S]CW?+>.*H3_Z X=IP+--I\M.1V.+*IBT:
P-O<?V@5TQ'LQ=TJ1_)Z/?(()\WU@)+XQUI\:3/> 6N/ 3RDENU874VKC<FUQO35J
PA(I[O)8%/"WC;/#Y^B[O1V)<\J4G1WG*1N56$-:=*7B9&9&9Y%SD5O7;<N'8_Y5W
P>Z1 <9O@UFXE!E[!;5_MHS92^R&($!90J_L9@?2[V^Z!&@^L#/9[.ZOJQ6&(M';L
P?9BZP-=(@/B%/P\4.DTH//19!:R)<HW"F8T?;)E@(N21"WV/QWF7KO3OPXH($:])
P:[,R+(8(3: *LQF..+^5P,,S-@E-S'<RXP6MVLWQO_-GXI@=O(KS\G%JO-AE9NM#
P<X'"Q_L.^0F%F]+>F)<HL5,EN7?C&IR8E=PI]>3.$84"$ \'=(\CL_/7P%Z)-UQ,
P-,EC%='72LN=BR2:I';9W>O8;&]?AW'W>LD7^H3Y"%",9UN-OU]HLQVIBOQA.<BX
P$UZ5A3F<Y2M/$X8)Y?-]4K(PAU0!*]^$^MS^]1G<\OMI)Y@'Z+[$4#?%X5#2<_<2
PA+O BW.^\J"@N/8S?Y]DK<WC!)H,7#02HL')H6(&X 7?<V\;TMSH#^BG[@TQ>N$_
P.TROU2FW)1CE$52"BQRXAWA]D<L^"-XK^1$3'7O(#>X7G8BP7BAR[Z:%!A)K$KGB
PS5=R[1Y.DU9+^ 5INM1XIH"%)91I]6K- Y1>/D\,E$<KG# UO;5CG_1[9.*3(Z4\
PDN4;^D()SU@ZILY4:'OVPGPD+"91*+FG*[SA +(<TXY*\CYC0*/TQFC"J+ZUXPPQ
PL=T.71,6/RG"QL<1R:\??[4J-KXES 4.\$,LC(BI(;DCYZ/P.B2WJ>@9Y3X\I-2F
P<*70F+,,=NJPVL5:VL'JF^K[H*6%.>V!?^9$'<_)9,'1A4@NF@%LP#R3/V%2G1'Z
PV'V.1^72=T(K$@$F'9;M(S 1:8""+W2,9/6>/'#B>]3>U! +&+%TRRWE%5W>Q<I:
PY 74,?IR#)&Z_5QIG1FKWA$4B5ZW(Y,!4)XA9E:1'/0H\XC$WSV2CY-Q)+7HKOO1
PCS<\9/.+07(M?^;^>#V[>C+XNS(3#H2:N&GEX<:53= 9/3>Y^)*]N$]IBD<-JW.R
P\_I('A+2+7FP^N=22*G<G!JINQV;2PB[(<,Q$"<#]!)B:R@J7.KQP ,4^Q7@&*;T
P,&$^!$*L;\-++3R7(\^PS267:S9$&2,RIV\-2"(R>\<I'<W#M;)"/>DWT:\('T@C
P$F\CDJ-;G,!P91K%P._(U6(6KSNSH:ONWZOM7IFC35:R?**\ZIMH<;Y_SO?C>?V8
PJSY ZP(&9@,9=+7V9,>W/6FE0KDBVD^'$("811>W.U^ .6[_^IJ#@]74XQ+^MO]8
P#=AZC9Z_&BJGEFL4:;G,A=VD:JF5M8UXP9U-!'M3IE!.]HH)N$_#@S#<3^Y)DCE9
P_ UIP;U>6I4-J"63@<A$*+-<*!==!MY2=2(_WT850(@7J^^G/WQ7M1^F*<5484UQ
P^R(X)MKN=T=E*NHXW48U4U,PE^U:F_V^+_^-#0UN+GMO MQ&?H"3S,B6AG'9'"93
P]U&]S[+ZSY>#&@J1.VI?.G6>'CPF6F3LP?!/(U-H"PD6P)]+:_4G(6+?X)>:<D<<
PGQQ3YC*^A&&G$7Y,0 ^&"^V[U:(9BZ1^<RW8XRD]LNO%[;=ECA'F6BQRI=D/(? F
P91&;828AQ;7C95]2&\#1YN*.%0MJ# 7;2Q4HY,Y4U X:%N7I"2SF[XUN-E[O4XKP
PCZ^K)9X&DP0S\-BA#3ED2VB>-9TMKKL5-G8,S,</[]X4YZCY;79L0^XT)I-2=%=6
P[3GCABSS7,;[Z_/7%'0N6:D)K<]^$WMQU+.EA&/M^][='$20 UY@?1;D(C:=AL)H
PI$@1*V-1AG\L@FU>K\H385\DS[?%<>[6%&6U2F._=M '3VB^26:)QD"42=>F\3[.
P> C28@'N.DB9+%_D%7_A.VZZ#JP\[Y#0KAXIRV:4S_BS-S^#"#VU<7*TTE?Y+@O.
P&OW4&EHAIW"LT;"<S%7G7-S+V@K8$T-G!5Z#E /#!</?"PX>!_FLTTCSS$Q3))JF
P5.205WD* 898@Z-*]HSC^EJA3NVJ-NW@9^.;U>76$7=:_8L9:31)AWCF9%"7 %OY
PVWY ].'HNV:1;&E"-.L#*ZM% N'CVH!UPG)/^W-H;X FNE[9!N>L;J3\'' DL?,K
P:4(RY&Q,Q/GA+IL1_H!Z"@H ,H ;3P"5^M#&=-M R('+(_^EQBFT$NIC'W<QC"*,
PX^L)J%3;[[QLT@B_I1\/@&Z\'>H;ZDJ-)RFN9(1)X(6#-Y%!WL+P:=FBCJ*_CP(A
P5 @=0:5 16@GD'R8,%I_.CO<"?YH>-8]NA )0-N143_GEN_^<IP2W[T%0\IH@8<U
P2T"E>QJP"S,)_>?"Q%+MXUCB:7237YJ0YKAX]U]KMW>P34#^]MC0+-LI@\FX3Z$\
PP#^KUWJ,A6?T[K!S*PI]X'+X>M]'&R' OB-L,9,?'G:KM 7GUKX7X124U7Y,FDPS
POD+TC\WZ;?Q;&H1U7 "\I R[R7#VS3BCQW+!M9VAUVE?Y.IVQ 5?C5L+^F[&$1W<
P,[=0B+79'%[1I*L\$V2.^M:\1N9WF1)7=Z\J25;PVW7Q:_Q)-V\LIP#Y:R:=&=8^
PE)<<[A+L5+#(/K^'H1+)I5V[CK3%^,8I2. #B#&)!"SS,W"Z5[M"]1PN%;1_-X]J
P" S^,R(9'PHF<O1Y ^:^03/^N&?^N$V:3N+)E82M/[J]1!A26)Q6*6.2Z]:% P>6
P'YK:EVAJ/X:I7.AJUN^F?XR-&AL92>D<Y:$-$,&2N/R1S+T&4SW(V[W/=C$=>NZA
PGUM'1,)1ES<"&H=GJR'X@;YLWLTE2@+7_$,K%%X_=>+/F[[;""Y.R/!H(?V.B%?I
PC(D<;SI&RAQV-$R9'3SULU84GG.B>7<-1PL&_%%$BUK_/!L\2,0JWP@;6MUKDU-W
PG('3#I <39(SD<<UDC+SN,O_/6\ W+=9!0(I<)>0Y?<^U-,B6R596:0HA1@7/;&#
PUR6:I[*)-PVYW(YO"B4F#A-&7 H-\A*F50!<JUB=H\M9X-U\FQ4?&?<IZ# FEC[2
POL$:0A!@D%LQ?C06U)U&HS[BII$#:F1!-[B^\L*&N]/Y6$3785_4[J.0])UR-1?3
P R]4+2T$7U9[0\N"W<?-@Y73"=W*T#UZD,G/LO"$>*?_%1-*T\93W6YP(.4J K2B
PS#@8\.F?869<X*BD$J77T,6%,/"Z.TV9XM#PTA9>R<+WQKFM((B^+%%C*QH.:=)?
P_.RCGY97N*HZ49B<.Z_Y$[P!X//I<%,Y2F12E47WYKDEQ5]Q(6 &_,HJ&+Y*;E\?
PO6Z)_$T<-KQ8()?<*PN*F?R-[WW,@!RHW=L%3!TT:)J02IMK&HUMH]YGQ36"K_V0
PY# G=5(3H?.FW=3Q,$W3\;:=E9<@P?T;4T99_#\\C\L(PH#T5!!1^A/)L-ZZS61 
P< M78NT]RZK4L$5W(I]EY)HYTQ8,-C&MQ+%J1JF&WX["2\!/*S8$XDF[LN/ )M@K
P$5]&KQ2B#:U#7&I'D*ZIPTYH,)F)VAHD$ *0XL(MN;$:E%L9> 5+,!)JF&#MI5/U
PD[%"$77NL+?F!+([I$]L[ 3IL4N:]U<MWL:T.'OW$249<0;,D3UTMCKM\"]N$B<B
P=SQ)/X("@W][8-EHP*XR3FVHY"EG4$P[(35TH0_)OM&^OD#,$ % XA+@';TOVV\3
PBK^N6@2UZFTG8'@090][O:(BY,56 &0Z(_N<?H_X-5G__/>O4*.T*:3A".Q898N6
P11;):1>O0"VUHVN7:MC3[FV5+O GTB<>9\*OK201]LPG60-/')$8:8]5=-@Q/?Y*
P@'[#W61'UB;YKT3Z $&AI>^/7S9N&;0YP^Y+$>6FV#7W+Y+%&U803X&&UK3=Q""-
PJ<#'B /T#+ !\?P08'8%(DTWC!(7*5K*0FB85:RY1;)4[T[C6*""  +O#"_5@79E
PO-PW\?YL5,'*WG:=Y/L9"YW*9UG561G8[/A'73)<3L,!(WM,4.MGQO)L2+[C2]B\
P!?G RI^">8_B<'?Z5J>]F,PMW1?IFDX8J6L?7*UGYX/1C6NZ_7GK=>Y3]APFJGZC
PS&T:9)Z7EP<+<@H)%<^<E^# $C8L7OKGV.!0?&B8(WCA.Z-E>@94'+#JRT2ZVYG!
P#B[1R ] ZU\C/*3Z.&C2Z$@VPAIB+:[("+\1G_6IZI-T'[T*)-4&S].45MPPX.Z*
P[I2<]A8=W__RVH"\S+-_]S-CE(!&?]!!/9]S,*;GX2Z??TI78Y)W&6[)E?C:N2UF
PY*<N^HN/(_CJZ?(*Q:Q<?U%\'Q2YM"94AYAK27SH=OO6<Y\]WE::CK_<VO8W$\4X
P393PNE2(UXC!Z**95C>F@%@^G/$-984A9?=A\C@TD/M>XY PY#QA(;'QZI!KHD;%
PB Q*JB]\\$LK5Q0<\51,\>.YU;S0@Y/2CA@:=.:.V4LJDP#./I!_KN]ET15L8Y2G
PAQR?M !$PVBVP B/<!(,]1?!>$Z?&#;.+[K&"VI&.Y$26O5KH'/4?_>^-W)_$KOY
P3C*NG-DJJTEVM.I"2;O*I>J$[>)6XKFF;2 KD46$4FT15$0^Y(D#YZ(03C-S*BS%
PX[>FZ>Z4$X2CP*XV<YMO@2LVNF_#3(NR<,MZ-TE'00LM.%5ZEGKH>"^*,V"/;*E4
PW+DH#'J_1>E?@$>"4=XYY?++R1[8J=2BYEV0Q1JKI3TO]_$S,$RNCZ?!LL):+Z,I
PX=G99^*$D8W,Q[KPVM#O"'J31VK+NI3I.+XKYQ?@07]ZH7M@1W28="E8"Y&JXU'+
P'?S*:#=@Q%K,UFZY<&,I'@\+T!58=_:\T,"9!_][JO@9CQKY5Q((RL0#V&MD1ETP
P''_=_J%+8+YOMYZY?QWM>C29^U5 *)*9M]U_62DS2+&<*'@LG>P)VU;YCVKE7XYN
P)L2]W.F' \@7?IPR84F <$]P@H=U:[E(O/TD,Z87+\:C^"GNL\(=K6N1^G?*/OE 
PNN=(@"9X0#J4YAX.N?%0? !;H/Q.E=<&C+I."U)AC&B^M)EH$6C6X)TGG1PEV#+W
P7,A# 35?!JX-2'/$)F=7*N C76K>U>R 7I^:\RJ4.X[#T,Z-)-8<P1!'KK[DK1BD
P@G :.G@MTS;'!XF>'W9+1_HU-;0"4S83'0IMODS:-[EQ .,4_PX:+ICC[P,I*%R-
P&@5/F(53,=TQ5+33W38-FS8GM\\0L&[U2'N%]07!H340K%S:T4VO3_\:DV:(>D_@
PJ2:3S\>"WV8<.]G\N8VBE2F[#?P-.R=.,EXX/11  7GX1/O7!S2WM!7G(UA__G18
PN3YKEKDH:(U9V"N +^].9^\\X^PG%^4I]9JRI['#3$WN8F)N:5>W9X,K\[VK)D,R
P8A=ZSX<M/_YO(Q$%I$(G1W4 41B'9==EDYTUKP"4[8LNM+IOBP-"9N'73^J3JVP9
P ?\T!FH!(&-)IH(Y!"C>XA ""Q&S89U0$ZA2NO$H$XPXFFD=76$GA.TUURI^*N0;
PD)^.:7>OLT+DB\)K/,X][QDY(RAX?NT3KGJSG;GV\."M@C4K4]FA>%'':*']L?N-
P2Y7>$_Q')E&P6BP2ZJ&73D>/+:@S&D;N=]B%![5ML@<:.@\'<8<GAK68:#YPO<5J
P$N@UZ&+ )YUW8J9K;D\2PWB$<G$T<0@B/&#96D.;9!>G37,&P;P;[Y*7ZX],#H-"
P/=V1=*/["!+V0B\D#O.$H'0.^CC=!?UMEQ\=R$AJ1^HA,?/D7!/.*J(R_2)62[,4
PGW[AH.;=1YI!>9IX ,"UB@9VV;;T!,!Y!V@N[+'QGQI)@&)V1;$23S*JZA?9$ICR
PQT7>< R[;X&4L*546&WG/#)B7FL4ENT^L[!\A4IC7L5TZ92/$&EE%R&2XTI!FE8'
PXUUV4K6OHN,,/@^6-Q2B1T4 \#*7NUE@XUVX#9,L 8T!2?%>XB>0PT'/,8@(GS'B
P'3C*_YE(\V*GMWS/AA-OQ?4TFNI:5LJ&FM3$R58=0%0?'A>H\_:0S2@I'3WR&)7(
PK/JRZ$>F-AZUV%EU5Z=[PLX?T^?CQ/SZR[-;>C*H"+WU;@MGI201"#A5&\H@1>H;
P\$)H[]"!:0_>M;M!2V <VJL% TG-]WZ/E'D4V&7V["ZW=D5A#9:6M.+ITDHR2]>+
P\!NPW<WX1OB\>A>1Y&F@8;K<2;NR@R7%9*V<$8.B@-YY@.N\[NAL-6X23DM7_)!*
P#F*D<DCEW8!$T7:H  D0%]S5S,2ZP;^.@KH%EPXY=_*'?!_=SIQQOA5ZEHF18R.U
PUY74\553RJ%G/V0)&>="NO7D!O CI4M@"4DT:VZ40L58"8"[SXVKB9:C>%<P3[^&
P99<..Y[4V^*\@*0[U7Y[Z]808][$8OWK;,<.Q)'@LT2LVW<$7I/1F"#$]TY'R!3 
P>1 C&:&AI;F')25%5;A,Y#;&G([M.!434_"7WU7#L)SHP6=.*-$C7S(SFU(A;#?4
PRI^FN(U 1%,^"2*U&L\PKIBL6/S<H1:08PB%V?G2?B;6^P;9K[=,#2$5&4#E=]VO
P[%UV311IHD[8QV#>'JTNU'WY=I&DEDB.!TJ\9FT*!6/QP-NHX1THN4%%#DUF?HU-
PI<3/ #"4+78WKY/]'^$+@P!AP>;0URO%I^I@V,?NS)ZJ(2*":#^=?Q-(_-8'SZI4
P.=M!L2**S/QR_SZN'.)<J^TK+8,1OP/TGT[,--.R_DP.SU@$M*2;DK/S81DX)9,N
PS8M+)?9 4,6$!C!O%5Q1HL?LS-%%G(%,9D+,))DHD^SP>J=1=%V4C9@V[&2C15G<
P+,>1SOW_&76@*!V,.TFOG[:I/R$*IQ>=AADW;6.&J[#J=[J=:0A/<0L3ZYE 3L3Z
P17P)(9*:/QO*Y%TJ]&!>)NYF-NMG5 !?=*!QU5>O7QPEP HK][_0RHQ%(*[42+%6
PI+GS*,AG>(4THR]S'Y]Q&!165JYY5["9V9BB8JVU)D_&QNLHR,\_$<6_@3:"8@#^
P&*<>3:RI2L)G+7E/["FK2\;\9!'R5,<>%MU@J^<!(PYL3"I_T6>U,X_^BZ!S5'VP
P!?2XEQ=;P8\&:@T*1!T?+$^W[Z9!NZ]'DDO @>\"&;F[$T 4C><5)=GPM#43K/.X
P9*A-N0=D,=<==ECM^ /%/3E/)8DD$WX#%/#@&V^C;U!;UYFZ)IH^?"<@2FM>M#*^
P.%Z7Q*>=[$#QTJJIH@B/N7!<"XG#&"$C[3RV_6Z#@M1XGW>\-_J'C(9E;M7>6X,T
P![R8Y+THITL8V#2"77>G6:,[2PM>3M;N@YH *X2MV.3"D&@,%T-LM9CGHPC%WB%\
P. (:S[>3%':RVLA7&CV^A.4#>LP4N'@R#[4( ;V3,-Q$45%ZS+DZ&W<X-S!N4- ?
P1\G%.SV4'%_"#U.33XPZXT3L$;<B0S-*. 'K**5QS,;K3BP%80%V4!ZBI_<D2W*K
P<5%ZQ:P8^X#T'7U(59[MBMY:UO;4[B Y&+X=3<S[K 0FO!<X.$ %LN"V_'?E%\)G
P>&>(_S9^)'H[O#DVUPLZ;6/GQ/34K9DK&F^C*,[LYG],7,J^=+T3TQ%7!85..[?O
P[B>9YW&K2MY;7*H#LAS]>EQ2^84;?-WS]HRP7/L&ZA<3E_>&@A(]BG1EZ7#:#L3M
P1*UWU2OO?;VN0)A]1A98C'\;^^.)9%HP=6;1F!9OT*+8;.R%;-E)[S5[(H#_U[>0
P>3HI/.FL/V&K@ KH:"9F3QR.",UF(_FN6OT/863_U&C);_$H>%$ -R:'2O> O.CH
PMS=?+/:ZR@"ZJ'PJ\!4*$$4[I9)0=H*[*<K]MU$>2R?VB-@=>$3,\D(\M>6!-2&"
PAAGD%_TJ;X?!:6#K:&#;DD@,R%=#4M%(?M9"+QHQ2_1,!X29WZ^\9;CWWPO1O %W
P+-@N/2<>6 )ER)QT"*EXFTSUJZ8V$[?4(S51EWHCUA!1Q>WWHD*@V=)M (#"873I
PX,OMNC;;[KWY52NG26'R F ]F4+$)A40W2].3L]Y'M4KV? !O"2FXR909C7OU'US
PX'&V1G!62)F\5V]>P2S]O*1B(^]62;.P>\_DYR4UGK=3V= U 9(THZ\[Y!(+52@8
P^S]#L<)03U35)Z;@%9=_>ZC%$0_;HI>N#]3@2HT"H_A5;EP2NSC?_UL1LW#  &&J
P?S !A^NJ<5)&O74=G$Y=(3 7Z]Y5>[9&4$45XC"P^E^/H:AT*(OA^:>U4<9;-[4G
P';V:T;/N]4";5+A=.W#P(8@FW.F;FC>>SGHO6] X0T"T\YK^@OE5GF8(;S!^+$M>
P)9QSI+KTJF?$G)(3[HD!L-W.A3$UY7F[SIK UNB*-[&/Z4HG1_F<64DV*O1X>2(.
PICAK'5F^^=(YW%AZO^6A:T9 YN/?;"8+\::* B+CTM.)W:&GGE^D?I:8EM12H'P*
P:LQA)TR_U5(*'I7PM:6.'ZY197F*2E_<3%^W\7E59# Q+X  :.R2%=E8%VGUYM#C
P$7<W%(+HYZZZ;>!]FV%DQT![5?*"-)(E 'VI:JYDU$"S808/Z#/HN5DHA'BZ@)#&
P=B7_H6UF3<4<R,^++F@E??%PS-9&"KKV-C53123JCGHRT014]-,(.Z[W&#T/;YY1
PGB)]P-"-^>VZ;HQ3,*T1/DS4'B_O"/YUJONR!C> R3@:"TR\T&*Z$EB$?%[!(%KN
P2M8<"/N^*,\G>6_'3]>3%AC^C4#)-R(I-QS7WVZ@QJFKJKO:[B+0I.)BR-55[ DR
P0/58U=M1JW?PH'R: X*&*@CCC&W(Q&ZXCHF]"]_P!_1P&3_C91EDIPG1Z,XJ6>WV
P,/V,M2#.V112$DM22YQ"(P#_3_T*ZHB#8^2MXTB\O[R_=YC8*XC$?JY='13Q!= '
P._]G3+X6&O$9N6-V0;GD#  +YY)@@(R"!@W-@JQP!'D/!O4 ,MII%!1^DV']$F,N
P@OT&8AQ20 ^A:_*WDBSW<D92J;E0/2;OV\VMJ5'*XV?H;K2SKEBQB'!DW80Q0HY^
P"L?=N$-U&0 A^#?V@!L#R8FW8=M7'I?9X2!(-#X9#(F_V,VF?N3U;KI*:X7,NEU:
P&QQ?[=/SBV$N%/\^MW[6H<2;&H"G@=D'T!T!3^),H<<SDWUNV6YW9AD<::3[6(]\
P)=".G"0_5R K7C!^X <H=B)U'N8HW9I:H!:Q_H>@9(OS69)AX^+;@2ED*#&8#3EM
P[F8&LZ+E_S+FE[7"A9=I\S2V-^ANT$;2HY^CX"Q560NTJ?P=^G,Q^#!EL[N0@>3?
PVD[ -Z12#;',-N,BVQUE"&6_*A>[&3>D0J>>F-;OLR%*CME4!J#.B8$HDS">\<QD
P'K_>D8J29ZEE.[:I5C/P[E]<_BUR\AC(8B=)7 Z* VMM'SJEZ+[."J?Z7(U-O:_\
PM^A:_[_;S]FUE'Q1C\IWRX+.L?XT5,4[CZLS341-!+&/^1,5LRZVH<MTU ;QI98S
PNV.\:;B,U\WKG*;J\;U0^,Z:TLYDK'B\7[4B:*3E@1*(]O:05GP(00OS?A(:TI?:
P@$C)/[+TYATALK5<70N-%T!<),S%C2*K0A.\5)M9A]&=?1!]#>$4!]Y@^:0-RU*M
P+0VSP[N-"L'(RGRK?1+^96VT(B?25G%SG+(A;&'*FD0EV^WGP,319;JVP:(H5)!I
P/4IQ(SX#(JF$S/@+S9EM%!N-:8V>;Z,(CQ_[CI;Q6T>%>S0**[,3C(7W>;W</,)9
P%7J1]=I')#_3I[WGK?GWG^N0EPWCA\M*05XHY)[8DHA_5Z>/C<]($9$6$ED<:R$>
P>#JEY6T;H5F39$%^%1STJZH,C=8)$KY[*>I0_P82GZT\KEX-!3S[=H-P7LKR7WJ 
P)UYH].7!WCAU<5*B"U*9!#H!8&@YZ%-KN:Q34=Z.)//\F&EC!EDL!W>2$:Q**HJ2
PJT+':Y5B[5!?>_%)0Z[3?,Z2\,K^-??52*BUZ;>[I>*15?RL7W>C.,CG*UF;G1K5
PIXHL<T30"9@[1/@512S/C.L,-(]HW*FWE?J7,(.42)KI>!'RCZME&AI^21PEA ZX
P/==F66JVPHT$3]=2%.D"P9))UEJ_@33SSYL=)O%<20""V!WHGT(A'#9?<^177HW[
PXS"!'?-4QGX*:5G5%]]GK;4OP("ZPREFF6KWU:ZB;$X&G3S74RP*%]DX>-M%?$ V
P7M8MXRU:OB)FWB&2'\P,E*/AM)7 *>?4Q@MT'/W-CO6CHQ*.FO]U)_^9\@/ JB6.
P 7K40 /ES7S\'(?O@Q";O8!\Q(0U20866^X *Q*N+9< X F],^\'),B/Y2)\GCE@
P"V<GC]Q/.75<(0(10EDPN75/I/3K3.?!C[W?NG15SOZ:#W\KSG@1Y<:VJ"Q"$<B>
P[M?-;6ZSBEV^TL.&ZL7T0\"X4HC:>:$8N4G9)S@:4#*G[ 3EV?@B@\=T64H.R7Y3
P:/&A050@*GS@TO$[$Z?WP@RGQ.F'DQPJQN6;A@=YI[[_0TUDL$?L?BK26CZO^7M=
PLDL1!:AO9VNA8*!Y]^4>:O7(SEWNJZ^&E%)628OA!#(-F9<#31[$3]LGZ*CC!G"-
PG763>H8'#&E(0OK/1&E%<3Z](NUHBT<-#:Z++F[=R;@H 0YA*8*JU)+C"!NL'_BW
PH[^).-= Y.GIUFL3^HG8T+E;QKL+^ 45<S.J4(#YD?;L!]@H/SOP#,@<TZ1,-A:&
PV?;],*[,5G7YE!KZ$';60\K_U"),]A9R!)O:6"'Q1F CWW&J)[BK6(50W4+2>!(Z
P$?^%IA<RP,!"YQ?"Z.-:)"/C]S31V,]'P2UC?L4QSOF'P*7V-Y85 7NP&Y@J0&36
PCB3Q[5L<?9C@BTQ4S,&WJ6]]7LFD6/A31D[$LR+[9CMNT?($2WUJPREOFZHTGKP 
PGW&:!&"F2)Y:KA(H5G5U2&+EE^"FS+K, 8[=W_;ZA[6_T$'8N^:(,)I?O(2[2/'X
P1VG Q)_'.>9JVB!<BD.++^5H9%';:\:0<@?@^5/L2.5V+I"W6\)86I+H>#_"%_!S
PE>CNGOG'Q11T#.IWM<E@-A E*&K*S@1>!KEPZ<WG_!\_-]*^S#$T/V3FR,I.E3$=
P?VO^S!A5:W2^GJ<6/,C>GB<X'!>-\LZ5!#TAFX-2ARN'\!>5-B3?HZ(LP:^QP&D0
P/&897,3T+#X;$!I.4HCA4E/7M'6WD#$2>/Q+A=,LJP,<?%L4V(-#0=;72^N % IO
PDM?LUH!LSGJ9:0,.D8H]616X@ II;>.7Z5099L?O,3*-R!% !:8^HH!^:+KI/UBW
P+ED@K@(FC-M@W=@Q_BB[=D0R#WPJ<XX>I5"KLFHR\Z#RUQU%#*-N<L$Q*&QT>D O
PW[[;_Q@1F$CLHV6M>^:/@)WKR<P1E'^4Y["*K%U9P@5ZWYU@1'F+T48+"S*));;D
P189*$R^V3?9+]"BQE\&&9_*'6U"QX!)Z3(L[*H_)?PWO5)%SY[TU]I)&WR^D:6;F
PD]!YDTPH-TBU7741V9H[I%K)QM.)!HBPZ\2 \^#QKG8@YO!6$)^$-\GYWMHHK*&[
P]_"=BAH*PT%U<V<-&'[^W%<)DT4-L(*YK,(/*T0]Y\ETFOM K<D8P"!N^4U>_S?J
PM#!:FS9PM'O/I[K*D8XP3HA?P+UB,:'M&XLK)&O[=Y>@TH!^S]TQA-A:A:^/)!FI
PN,+43<! 'J9'Y:4I"RW ,W%6#O\Q9RYY32TO_BIL@^D"*8J,N%U0!)=A& N=4/QE
P%Y?-9J846->K0,F@.(U"$XQGW50) A$=$9QOKU<5Q4$)!890H(/%Q=<LE/MILMB,
PB@/KQJ+-S,8I;%YXS@W>FMR:.>T))</K,/=:+* (%V5E2U7AKKTC&R18(?<89B?T
P4\FA<;AN&Q-C\'<RLWX44[SB^Y2KKSULBO@VIS#VS9HHCX)SV'/\)+K?:5'7]J1R
PS?>;MQ$0=39DLK6Q1$*FZ+X15%:<Y!CST_DSAN<AO4=4>]@FJZ.(YUJ36Y2:3?@0
PSW 4'Z_@3'VQ-5?=,1.S=_:]?& ^#/EV@:HIT_<VXN^<6*Q(C?E%D$O'^9O!RJ+:
P&0:OL*\<FOF1:"$,V.FEJ)23;0LUA@US,"\Y\TKLVS5[598[]9F3_J,('-#*6Q4[
P')3 4-<(H:6B^\BZNJSPW5SC.WK7RBB=(=3W0%^95 9)U]%>"A\6DQ8"*1R[\0?L
P>6H"8YBN]33IRF+6X0S:IGG;>K&=2-WH""_>]!53/_)'ADKEX&N>N!@\J32^5%5&
PTE3;4@8IBZ<J@YH>2_E L\(L7">U@R=0,"@TTU_1BN$)05,P%1!0 *)ZT.D2<(*V
PC9IR&V*NVM]&(I'E)T@6J'H@G*X!JB36QML!T'65V7+Y&=]=;G0NP9P;DY)@NIF#
PA8KA0;CLE(^-"OU8G*8%M(UWOCJ=C>)2@K9YR5++MC=9%?@='U-+&'6^%.?:U.F2
PRW\JRR(*%_?>_)*^.^IJ_63E52S]_$P9B=G0$/"5/J0TMT>K6#AJ4VKGC%*"J/J?
PJWB#'TV^EEQFUS+-W4G69QZ@V$&Q3R"3L;X)ZZ#[8PT!SR\$X>5CV9G+!+(XC5[]
PR6< LD7*KX3I]0_/8#H9%%XBB007*V3:^WGAT$XDT^.!56LOZ,8F%X3# ^KI/I)5
P.^D^>PI#U8Q72[SS/U*8H!XO24+,'.2I[M  "NVAB:5;IR3MX<,VNC^XV)T;])CJ
P4JP?=,H;LO2@1:.?/=.*%T[::<.<+?" 0X^0XA40'H9'DRKJ](I0-Z5$%5YBJ/1O
PSVW_]S9:B:RY([PY\?'\*BPZIRIN%1YXOIVGOB16.N&.N_2IZJ<F)GPG ROXRG '
PH&B\5B&S0TMB&UW7,Y@JI_BQ59R=#X/KA/$F)!%I+!L)O: V RV'^Z>SO0L)?)\S
P)W9\M6%2A_H2S@)M$A Y/:UAXF8X;[*[SU^XYTU[?[:EH;Z.]S8O7\I HGKY^4?L
P' !T9Q_NDRHB_!?S:GQ0IBXDGO!?G.I9GV#IGL8T04U;A<Z1YL_"3!A(A,GTBLA^
PAL&^_B%D-F>QTPTH$)>;;57I'2=+PS/ZU+"_^FE\MA<=YH-XR0-J?C<*5!/L;&,H
P*2)1F0>()[*J5._@@,AY6*+7^=&I<%T/_,";ZR9K]A>4E*,/:F\;2[0<MFH0C$/F
P6#;OCHQZ2O^$K6&7ZI1TA8^U.F4N2L^V[M:RP,G)8HL;5+0,YD8IWA$LB5; ]J69
P#79_FSQ#SALJZU$<XEILDVQ\Z,C3R%:"R7[^[&4JH%)*5B302L@!A/,D02'E=S( 
P8;T?L(VC$8;@&!3/O6AJRN9;R7_+2R!F^[@Y+[M7.F,"*>U/E$UO;:W!NVI2YHTD
P%DOSW7?<1 X]L)GR2,.YYR%S3>[Z<^4$;8U1JI-J &\:XJ!T(!:U2J08*K2WL@&U
P+W)J74FK&)V$$"K,ZWRD8TM-R;^W'E/=RVE4N, L@6W=B8+2>@*N<=4-:Z$]^*)4
PGOIU  :EO,>");,>U.:Y^00I--ZDASA[V102U$MA/-\LF+K1EMW.XEC<C))0W=%+
P3&2NQ<0/K$79JWRLDW_A/+&*:E!\QRQV&,9.-3%=M7(15/I06\<28(F^9H[=Z6')
PA:1VB+FZXGQ29UKBSMBUW\'BD@TEREY>N"X-QBHU#%AW5,@2-/>U_,<9/$*,%01P
P'DU-%;-=2,(0_";Q=&*"V_\)B@-"^ 0#'3'$_/U_3;]P*WU-.= PP)] )A@/'62+
P*4I.(/$S.*IU7CC6IGJM<Z(;N) #"28BK%WTXP0A9# 2S%'*_, \N+Q-CXJ<JB7!
P)A\GY!*H^ H%^AV)S10*FOCRF*@V#"\"]^;S #KG8K>2QE@%UM\2P)5)GSKM>>&%
P1YAS_D)%2DGY*S*R>$: D$;Z HN9*2F+=4]V?F )OV)SG%Z=$M67 PND@O4(EARK
P,:<CB8P')C.M&QT7&B[_?/;CP()_):'V@]M\\N'?S# W&#89;UXT2K^4AH"5W/C@
POH-3P$\-B/]"2\HR4PT(:6(_*;:6NHK[B-(%Z_R8\]VZM3O'O3W":.8+IZ71'-7E
PQDV@1%F<6^T.A83_RZ[;<_ I*KC5LS"TC?3YZ#GQS*;W5]U,O'C8W/\-8'A3,E4/
P-_XU/BG%AT2^==5U%JI7A(FC133>+F]R'J6CC7?90E8$!B:XI]&%N6/[!Y\AH0G*
PB:ZZWY1X[-<&I##MMJ#C8#KV)V8"0A."(6%07)@PZ-5^;)]SYE' O$XP.N4/IZN3
POR#E[]=HU_W;'PVWV'<J/1TBK71AA;_-UNH2+R&\NAU\4BN+%S1BY+B6_9LXUJ:!
PJ^?0P23I7B.\N287RK#5+B54-^73:I]E/&<ZR;/&;&_86[WSY$,FJI5$Q &4@HJY
P^H&C76;\E:,8M)W*CQLMJP69+>$U%/>@XD=1E?6*39P>K']]""PO$S!7QL<R3B@K
P?%#"F!0J9MT1MM)O)ZC^=:YWS%B%?^VWQ4Z/_, )TJ;MVXW6K.&"N(%@JOJ>/#/4
P++:E*W_G@K R#T]!!:PBP(TD&0;KY9&=2$F,S*P3:H^@M]L&P+N=D=1V'/ /0D$)
PPR)ID):%2]\S/A[<!JXI%YO#0.>'6=D#) #-JQ/\?1CY'6?CEQP?9MVS:3-#_J(C
PF\63_!Q(A7($-!IXT<>/@DBB_5KKW)"2S*S,=]=7'%DB0&$6(=O(FNPU,.JMPG:8
P'*"^S&]I5%F@4H\NB< 25L=Y0]'CUV>A$YWW9']Y+AI(QRVG>F38=TZ&S_0>%X[@
P@*Y;;'\/:2INYA9"\HU_58GMZ3/IX!LG^X@A@+R',<=F/3:+[R)<5.$ /A'=@] 6
P@&VK*9FG2="ER403S1GNLAD_V'+B9BW$>+) (/]"CA0[Z19$6)&_XN<_HF9;L.I+
P/MB>PGR<%H__#* N<!_+=892*T4!+KZ');I?7^JR].N6O!%%A U$B@=)C.K08B2U
PRA)H.T6R9?_ ]A%V,B@HPJ=K0!7HW[Z+$Y$JXXZ7_2?Q[+JX B+QR#XC0)T"V&X(
P0M- 1[2T3T;P*Q(]!CB,*='5[[MLERDEM(WCW^?PK>X$:%(CD6DT<X&]J"U'_CWT
PKGDE1#@XA;81G#<N5;VK6(("=XA_<!G!C$R5589Q@$IZK1.,U]D'?-]\G8@>\XBE
PA(QP_K++!=G6'L8$YQQ.FLJPB2[41+13;$*7RFGX :'DA[3X; K!\F)#WBO3/TVM
P47B3>=1'V;6AM,]1.:YX8ESE)/M=3Z7@ TN%ZCX#^\X#M5H$6I\URR,>ZO'3FC,N
P!5+:3W2$-$S RIF]P, $@2 IV0TP#1< 0,M));3\P1]5>?2[:S<_Z/,"85]?,8Q3
PZQS=N#\V[5IW^L"O34K:N!^%J7:\&A3ORI)EX(*%6X"=C(/,G?XZPJ''_>6[+R6:
P&#WB+P5V5*(J<D2?=JRH^I66%=>=@O>!2H9D.H45$AU&8Y$C-G$PRJWZXSJ?$[CY
P;\;^Z,P(:X;(>PLE2E& 57E&V%K"AHF\(30S;F-7[<2E#3 Z([<,RII^NZ7\P@OT
PJH- U7Z8-:Y9];IXP&12Z]VTJ!J"XC-A8R! 9V:!%DZ)%:K K30\1ZIF+GBE-?NA
P"N%@<NB\<C1UA GF&'0,JQ<?:U6^!LZ&(/:>QQ22FP0S4-)-U#PK#PE)(RRW([[1
PS\BMSF1V LSPN#DPVL2FIS0D ,6D9Q1U#@G"B"PG*Z.\*,+0B($^SM_]+@B/S+4E
PP.]E;TVFH8/F&&TU]1!_-=LR@E0F7XP09SAA_V8TK"N3]2-PXF0JLU/^TPYG*HZB
PJR3BS234*&N#LE34ZA!K>JE/(<A4TF,"$BX:R]ER^N]1K]+NX6R:0T;Y(,?SM867
P/4)N?CECEHSL1=<I8N.Y4EU3GX/6N$6>=]\<L'0#,P/&G46_V<=(L6_.B)ALWT24
P^K,OZ?T%P2"E>X?@J-X]_ XSX;Y/2RYBZ]5+J#>\H:!GE3-(3M+ (OH5O8QO<0-4
P/"H]6451XAO!8%SDM'.)'WHR$")<*\_E A=E??Q#N#!@K*_WS1AK*;N(4C9':BDF
PW&'7I^JYXL0-?;T-K'XG<X$$?LDNZ#<4%6PW(-;OLAWI+2=A'TL:UV:3CU!6IT)=
PH^N\*EMIFE>X<A-7W0G3V\]_W/LLXL1HSW^_U"YFJ=Y]J5T!XL'K17W#)"3G1]RL
P*1'V 1?[=5%'D5; (9#3X7ZX,=IN,UCN8"%(2I61(L6C%,CC6G0"MM#J,PV<_?L4
P/4OV^DF1IDD,\]J#X@I!,04U?*?<0F12G 6Y\(01QC[YT!T'YK8Q=?KI0820N#%O
PY "L+]2-E:N3 (T')RRD:I-Y.Z0))*]928)]:ZD(5TIZK]\M_%](5AKK=OM3V10^
PW?H=EI_]RZD17252(?Y-JTP>#4V3&;<)5OK_>!I^R,/\/0G'VO^6E57=<!;B6?WG
P,!:H9]KB2VH1'7B3P4?J:/L;X0^%UD?#&%]$QHN:+F#@'=MELH9-)_>#H>@RC=K3
PQ['&"]R^BLG@_?W#:47+2_4(FDLOQXE0.@U*1ASG:H)=W6,5)(UA9@0NJI"JGXD7
PD6_^1MS#!ZKG-=0.P386.NZTBJ ,ZYMINVU=.[H<0, *;65COXI+BB SPU01.#3$
P5Z JFL^-&]R3%OCY%<&EOP]=&"$UN+E;& P<A<U_Q)6M/,7%)>G96HMQ$YG+XU4*
P@.*E @'_ ?,4^GD)((:X>0,*\FVQZ5 P0U IU9HNEY:3<86$/](9D02?5S?C1,:9
P[LN 6N2^$[LEO%,I%,+5'1>2%KH#T972IK#/W@ VLJ39EZ%!1[S<R5,X3+'X,\CO
P&X[$J?\SC>@3^7O<#<](]9G8A64^:=EQ/FO"1^1.$E%"9=P5\(M+C=F?T:TA:_F@
P!$ZM ,^WB H$MF)/'+@3_' %MRU[,;:LC*S4HUN2KULD>C:YRS0SN(8SS;A,,L<E
P=SY-EG;>DF3K A[!]4UO:"(*;UN@;_(3(_7:V19AL[F=VF: 2J6$5G"N>Y:D5F&3
PXG[^5/[:ZUF7Z.#-*Y=W[5=55B$KZ-U.SWKQBV'IAT*KQ^N(A,A)?^9IC4EJO'#'
P&WH,VQ/5S>Y5+48E=#,'*5R\X#'#(?C(,,#AA=DVL.2J"SX?:K:-GZ3(.3]R3#J%
P>C<?0DVV3!K/L3;8V20%!Z)*ZS3H#8R3*29HK5^.%-_7Y#Z]<EK90&5U&\=\ 5E.
P&_(E6UOPV^2O9D76<<^C(!M-RXF(9-46:&2G=__030VIW)\U-VO*6Z!QJ'/N.EVC
PDM:H&A5RM0_>#]AY15#]0=+!/\8,FE;7&*AEEE$.Q(L>!4<\O)>*K*I?T\)?+8LU
P;<0,=">O"_MOD=6(!LV[I\6=OGNK^/0GG*@C6X3LJC2!9Y>I9 NFOB13XE^MUY67
P,N= "PUP:,^:9.'BUMUBZBJEY*><0K3HC>YF<*H!=D%6!@/*)QO^N$QZ8T0;&-2\
P"+)A AE^.G/PTZM2FX_14&; "=KR=!3$A,\4+;[/L'$3]LR;Z7 DVA#1GJ,Z9"<W
P28C+D5Y/>9/[/? (;Y[M<BC[X_V+_L9W7R]ULMDUKDGI2GW8WU6O1BG];3\6HVP+
P4!*>R-/O.Y*.QL.&U:D\ZQ-'0AU-I%0_-Y?HZ-#F[Z&!V82R-9]/6M<MG9I"Q4_.
PLS4DJG7>"].L9[VS>[K,@:XK( N4'R9>FSW.<\:,\_<S3OF  L8W29:1R-FZ?_@'
PNNWSGL_QLK%6?9>-394]21'1],EJMT8?EM&C]-)N**\>>+0WK4KTSF2WY#[BQ.YR
P_*R^/UL?]0'\';'"P]'SLRF"ZSO(D(QT#8<N)T!E:*&3A(OLMN144;_H-JFYN)>=
PW=\3V8V[0%@IP(_+;Y66DA-UL-B)H^M?:%\N'R3EFSYM.!"%P_;ZDJT 0D',[U<[
PZV1WA].N4B#6#0>'"^V/0B<N0"\K7UU=:Z[YF]EGZ_,',[2O=4^B'%Q>!^[M0&2)
PE@6JBH!@Z/OZ#;&%O@<3)^ R:9(6E$4#?<(Q]NN5;P+KS2(,\M4NI"1X6= 5%V[Q
P6I7),]_H<:? WG-FS2\&Y&PL924QF1I_N#AI\BO7.9\TY\Y6$I9!FZ)A! %BJ4=[
P&N5[5%^\D/FQYQ\3K=G7<)56J+X$9*D(?V].EPD6&*?!0C]/LM[A"IJ7KEL*G^U6
P,D,N=W(JU_NCU$>Z%[*H6BOR7K5[8J6\3; :%9J\7?"8?<Z!S7 (PE1W:A&RKRI<
PS/2EI%RL!3M@.5D.?#&!Z>$7#');+$H^\Z<ES9?Y\>L2S]^>?3?O%%JI?FV;>+FE
P<KI)6F_BTV1X4VH_O;J0AS\!ER<]"7%^PE/M#]BFM7T+\2>UW<+Y-2!F#,V56W$?
PNE'A7YL?IL:8#<'*PN M8XQ?<QB!( 97@XIA%Y0+-<)7B8_0EMHTB]*B=04_/T1R
P=)28G5U0D?T@X(<ZQIA/4M5D5.$]3[&Q@]$1W9JM'W M7:3;A.J/A"F?IMJJ#%*2
P?^&>9;IK3#M(7\M57LIP30RSPJ\:I)7V[/K_#A+'*,^#_4OV]W=S]HFY1-LE[$:#
PX=]QSM9T=R,NN?]^-OO_.CR(U:),6EI#A*5<^M8S3:]S9S^Q%8 R;!Y<YL.!?OC1
P.5V5%I%^TC5L%L8PF)=E'^9M&#O^4,MBI;/TB[/79/@<XE$W^86.D\T8_<MD'J/F
P&G#;Y/;O<;T;\3T$"!-R*L8F_BG.8/^':/6;5G,7Q(%X2<J+YF37R+%5:IQJXN>.
PIA@4$D:L(V78G[1[4:!IN>*33&XOD\.5JL"XP;#_NI+5YT(O;4A9OF&N-N4Y?IY\
PB-1:5H#1$W;X;-?P,!B$#!$U^UR0PL,L@F?*$B^!V!R*_ *V+%RYVF/X3)VHFP7X
P7YV-FS]X)<<3"L4>JM)TZV^H*2D_4TY<X4'GLE(UNL_* BKKM7VY=7BN]M@L+R%Z
P8K)V4X=U@]]+.77H7M@7'MXC$@=H9OPZ\XTUHM*G:WR2?8^#->)-P;W?R0Q?:.:R
P=<//#*-([NR6]*]D^FB?Q9Z.5AU_Z!@#R$'TS'@Z^(<"B<5E783K:.C/.N6EV6N.
P-"QR.<CUY!:C1N/K#9ZYINNH.X-G4$9 X/6?M96XGF5VV=CF7@![W-/@.5N_!27V
PYC22'MXE>@9L$XMK\H4P:Y><1&O+6CQLK,0KYH= !=$E2^I$8[.">T0O\;;NY5N?
PSAQY]=VQ>Q!D75X/^47XQ]-&Z1755G04"Z688K[EG#"9EC4@#CP 8U&N$M+:B*B\
PO Q[SU>QWXOL-#97@DP$I19)? I8A)7<@XI5"1C62UEQ#E]_&M7?!BW/'6H"C).U
PF'(,\$P5&;(06,'%I._MTUY&M"P82H51RZYC'[7$I*6#\B<("&QJ<1^]'\!F-"=L
P&#X.MX4.9_-9#J>V"]TC$BL*+CFN2;$LD1R^$K\4(LJIGL33!Z9VL_HYQ^;W28*=
PYOR48[;E4,GZ:T-=?52,_;;Q;50+U\5"46#SH@QG^Y/3?U(!X454GDT\Z>Y*F!:3
P!9+*([L_-SD]+0VT]'JU$M!'JG[I/H:8SM0\3ZX-',!/QI29?J$/,\V/?\A?#2.I
PIV\DW#%K/41(--9^)ZXIERJOFVT%?I1>N387GZ>A!?4YPBLUF#7[^,!B+F4L08(S
PC<*$J&\^Q3S6:@C,=F^G\,N#VWU9O(F8KUEAO'HF5:#S(HL$U ]@RJ"_>_$WP.S:
PQ/*/4'>NP%P9/=G$S<WPAU % 1\6QT2#I3JY>7837T]K2(0Z4=?CZ8C?E&QC>.#'
P1DIBMI#=14R<1BTC)WD$]-)3;&#1!</F?OYR@ @'F$2CM+"F,-="622#-#U-64K/
P*[:N(!>#^PQR<1V'%P#5]G/V'-W!1#6A34$ X(\QND".!_R+]NN1INNF;3+WE$;G
PL<!R5P4FC MR$W=LLZ7GKBV8Y&H<:KPXY/-VC.:HP79,R!PF/CJ9;L<XJ3^=N&/?
P!-IDTF0V\+R%2O4WGS&@ )X9MF\PTQ+Q-2![8W&G*7IN>G*3C=]2:D&5S/#?_175
P>J[ST@PQ/%BGVUTP3+?1L(]S]16QRI>=I:&&;.KYO"_A<'<\ABHZA#S<HG+2/*42
P6>> @Y2CA-7ZF]11/V4(K8+7_Q"-";+AVPEO&> %%%A]8AFNQ"20SO_A68UW:/3]
P<5Q^NJQXU=)9F5B'B&0K./QN^8/Z)^Z7"#NC"#A9-4>PO;6O=?D*"A1C24)?L10#
PP?SWX)_C&>&]I+;.'XM)JAR1,5WS44X)^[Q7A:3L,^Z\XLLMP31".'<<X!Y'LG(+
PU.X+340EJSY7"-C=EH1E/1!>JFAKUA&,R/[,MN](;KCIS?E9X7@:,XIG7$!"TX82
P]69N_^2,BL4!/:]19&ET9DN4/P\1#2E^>H)BC #3H5+.(S1&[FVU7B;&=JV$M\M+
P6X@S801<HVH)Y&/TX2\2Z+]_4L)>0#-KX3C??/].BUKS *&1T:CME?RQ7="L$Y0]
PY;(-H .>90SM89_$HLM(+28/0ZW*49;FP;:H!9>_'*A:O,3?]R$L^H9L#T[O9[IE
P@-SZ2=_UQ(^HN:$.\ MBY2-X$*9MQ1'@:M"+2[2Q>,^<=#2#?INB=O' M(GWK'='
PZ(Z#+D]Y7Y(#L8H$4<'D2Y0J(D4%@:PV A0VYM$0H$7/7%-0L:+:G><#*[ %-=;#
P_B]7);8ZIUI,C8GUHLV*L1HFK@$2$Y'FA+J.L<V6/=CJM!R@@#IX#$?97C9@2/0R
P1]E_IQ^P>DVJMPQN*A<_8G%\^%?^LIG+/:7IG<Y!F,OCJ7,LY00<B^]7\F68UHH"
PJ[[Z>)XOXX,=U2P/^ WB]Q-$G@TR"+$>4,$*UH*0K*EV9OP6.FR2LS;__=],Q2AN
P.ZFO99 I7;5S>R[9?TK?$[V%,(:#CM3PRI&< ^;S9S1832H;\ [4QJ6O1N+-G]^L
PK9-4@!W<#3.IWL<T:24**QFG,1*F$Q*O9N&?94BK[T2EA7K_)0[>A,IF5:2NGI>Q
P'/=U)B\P7 HX;K/$$>!H]4QP%"]:CSBB2'A\B2D")V*XI*]B0@;RL4:YI8;)]/U@
PH-E&G2.$&5;6XS!4?GC,6LJ=;2N[RMSL6OC"X0@,TWC);V&$J7R[=3M7V4 BFGC3
PW"IY:Q-7J5V,,8*D&>'_.Z#QBN>YH>,;2*1,S6)M=@ WQ<SD;=7'C@DT!\!VSB&<
PD>2BAU18_?_ZWY7W(TXT^9:&H@WW8A920LAH%!95*$I15QW:SRR!-@&/NL3E-4(%
P4^^S9_$?*]W#\JC*,4R')!*]KL$P\5Q/1691^7^*6=+X1JX,&&HE=>5K 9KQ_*:<
PX1E#J%-!#F8(E5GLQJK_K+]RZQ*IB7<QL0<1T8&T!6K]'RALQN^2]"K"293T_@W?
PMI$,DQ 7C<8 @9D^C*#J N:(6[&;=@PH"7;A0QUE_%VT_^50_X <54YE!NC0(X+G
P@XLP%JP/?A=>;S"SO&$>(O09OC.S"1#SAS'[OW?2291 RU"$1(KXS'V RE6VVN,?
PS]R(6CSRGTXBH5B33%UG41"B9?]8NS@GTY['MMP8M!71DDZE4]SS OX$X]=YTAK!
P#$K8X\J8FUY'D_>%N%T>AD(FWZG/H8V<;FYX(:% L+F>N#GZ2\-CWT@P-OZ0G>_U
P.*D5PIK<^T%&+"*:=1;@GQ<BBHQ;NQ#TCG7:]V$?ZF2-B]C18J"U1.?+IT//BHXI
P0MT7;^0:@G:\OLJ^?;C$-??UL-5-(>#5TU,W-;#4#$\O ?<$IK5!V2VL-GNX_>FB
PQW!$^BO+[TH3K09M'KM5Z1^K0S62[YIA$%=TK\IY+C EE>GX @]3T+Z[1WX0;"\?
PCR]NI(S#;7#*R!MS;3%D^I.^G4EC5??.5HR'H0? RQ>>-\09;&[FUAE:3&4$Q\L%
P8_?O56LB5?<DJB?'S;^B!.:R&A\O1FIB.F+U<UQ<,$/N[8.HEVG3'S;T@;F$NVX4
PUX%HE[!EQ?O2Q\DQ(%0Y-X9]Z+OB1E=B'I:;H]M=444US\4^P=4Q(YR>SH <I_=S
PM_=-YR7[2+GTQ.AT1<0>E8..= R9N:V&3<HTW-,OM@,+[$A(K5\NO+H:^(A+7B,N
P_XYM<C&,M;,$T6K<T.9&UV/>VY^NUT)9^.'[O9!GS>K!>*+QZL6!=(7QT/:+7B7=
P"OUZ5&/E/.TJ)GVE0 Q NHV0&"HP8+$2SV3=15B8A,>$J2'YIJO0]!#6ZAXU7+W[
P4L0:U^%\+\15VVX:S_<A0UL\*<#%PKL4.R&?),:GR88I[-0-] ,EYK&P^^J2 CVJ
PF;J\SO5*0D(VF>XH7KSLU5(*13]:=&GRMQ4"<62RP=*!7=.@#;DIAW6-46JQ\.+-
P3C5O:*U6C R;XV%H2PS"?N1W&K$YR%>"S3)R;SL![FB"+Z'+,8C]F:^CE)IP,958
P=Z59*D2Y/_.0G4=O"!3\D[@UAA]JGU>N040T-@U$?>F%V!;:T2.&YD<^;S-%B,?(
PGUP.L&7 '.Y?@H.$!L,E*J438K XD N2_'^.N;"Z5IB#-R;1U4>KDLV[<".ZYU-/
PA=KS^0#!^T1GX$2-8H9$.(J%G"G]5IV8!"3! <MQOM[MWSZ.VF^AC[OY"PN=9'77
PLW+E)6/HPU_&8K58(;\^@I]Q5:H<EC+R,5[[_![I>VA:EG25YB1%U1+R-\VP.2K 
P7'^U#H"M.&3[R_9\D=KW?*;E;G-ZA/*U!INY,-\^%,[^C5@15E^6NUV%HNA9B9CW
P;M]]/,COR7PZ4<96:#\EKR*H?M;=W/MO3VQ5(!M8)5(XV0F$NG/UNAXWEB1V6.<[
PLSDI*0S.3M[QRV-3F"\GI"&C&3)7SSP;1*QXOS=7GK8JD*(J3$5CE.15$:,CY"<?
PO#CZHOT_3"B<N9MB?&0KU;F%D3*X6<JOUC8R9SF.1#$T)]$1'C%R1_07"2BUP:"_
P1-_24BY"P==B7:Z(Q,IF_&SD5O KJPWZ4T^XHTB:$'>W^=O;[E*W&B]B!SA!^R]Z
P&P2RB^T<?'2)ZZ2JXFIM'2:ZE%[N'#:C1;S(PIE'ZPE)619?]&;)ISLV-?QS9XW0
PB*'M[ ?B0<A(6Q%PGDD4S\W!4*KN "(Z*.<B_T$F&)&V>0&DX6RA6?EMS&+KB<>;
PN)Z\_>_P JZ&0MY\*X =<\D>ZHYS&3!4YW/LMB9J'9+3> E!W?SW0&H(Q/GU. 7G
P!Y9==C5YH:+M$-QH1";5XY:AS1>*3 B&A?V?:4%CBB=ZF\-Z*B"R[&W9LK/PBEY2
PYKJ+L:I\?\ !KR1?BD1FZ@LW&2 -=XJ/XMLQS@CQD&?-F\'LYDP1>]$$:.XU]__>
P%.:C[T6F52GKA,3DUI$\:R5AB+:#@2=+RC+8KQR>[>=FM:4=Y>MW46YT5D <N9N$
PCKF$X0=P4]CJVCIMN8K[OKF0C?J'D1QU\PNX3ILCT2.MB SQ:F ]#J'YIKG5O+$F
PK6((L91W0([]#-!W RU7Y*"3P(V^&7FI"A=J)@K/ <0.8NKSR0O"W:8*..K%/QP@
PCRER6? /P?\ OSPZ2474BYU%=B\HB&=U0'_6I6(U&T$;)"FJ9FW+XF-CN61I/=K]
P-9DS/M6L#!;IU(O[6JY-I?*Q<:8IC1AE+>SC%R//C?9KV"73&%1>08VSEI&<2]<L
P;5S>B6R&Y7KY0?42QD*OL@7,$<LHAI,$$!@L(@(BL*?P;7@4<S2 "=K80_-F=*A^
P>VYI%C7:+".94'\[VJE+Z^CRR$)5L]NV'X+<58=NO]5G;$?R6;D\+@-Q:^*HKE+>
P5,IC9#[%V5JD*VTK[X'YT*CI6@^ >GPZCC\*J9.J(S;NJ>(M09&I36=M#:O2LY'P
PW62( >!3;=X+ZT[P^XIG>?FPDTMQV08.K?-;_6L(F3,#"ZY"WW.=^85_<?ZMN,^Q
P,^9XY8'7CPR14_"OG<DV67I*F>U%TPI&$;V*:>C8:B$,>VVE5B=H]SDYA_<J)349
PL]]UP.V7[TU^R@ -]L;8]*-;HA>0ZS9C("!G>'6FA;XCD])Y'X^OPU1Y0T9HR3YD
P[/CNJ)SEN8\)JRE=W@62B7%_9L23')3@20'3X,9)UY70UA8E>]815[<79GU/B\[L
P?SO-?,D&MF0^E@ Z0I0650]"0'8-M"$R92"V&%/;"FE_70@0;&.6&="SH.PR<F%O
PV,I]JZ'_PG.A36D**'Y'GJ=?-Y:@F*=QFM!?,^AV&F\8,D,=N.75\R$&ONIJ1&(0
PW1Y^/I @XZ$3<HV4TV'?RLN5T^%V$"JBT!5"M*YLV#9&L"\]=AGH!:!\%,_GMZS=
PH_%Z6JJXWQ,'FK=B-/5UMIQFY]EEM3B5)-3UGE):@LL/<5;H.N+V[B*Z2NA,'^GH
PK!-KPR/4;K/S?'<E#QGBFLX%MX]:!CY6YXS,9$RR;=EK,O &81;LV6!\3=HPK=8*
PO[H$<JJ0];%I7P8K">-GN_YRU$J)3#5T3-$:WN\41>_WI&TBW!)DDDJFC:C-FY1E
PXWWR3C BVE.5O>U/Q>1I&AYN0Z"?T_<[5K4(?MH$%M-/1NTM VQ#>0HB<CZ);XEX
PC>R-?[3F(U#NFGT.:G/R7FV>H1;%Y>DK$P#-E(39DQ4JJ=TD< WG9B XZ@&_T86E
P6KCV4$T5*\V9;MUF[KM;A<7N^9H..IS%=ZHSB,YJ$EY4. 4N=2Z#5YBK0[ \B,M^
P>Z&Y67Q"B4V\HBT-##L8(U) (A#MG95 +BZ7#.],"3,$K\^"\92:X!.0@S0\O2.4
PPG9VW]+CM6Z&J*GZF4SY1Z_4$<J;&1I, G?EU>D (S.E]YK%D)QEA#Z#8@^I=3PK
PS;7=53#"V,0,XKKH#')P>339WWV62G.ISFIF]OR3/]<(!!-2<'VKX!)W-]T;U@05
P*D OW74BM0G&/G,E&-7,6#;!>;DG7;7+ ?O&21_FFHEA;T*YJ'IW4V5"3(:ZK EE
P+@? (?[ B PEP!PQPQ\&(2@4#>"@;R\@ +832%<&1&;OD_SO;UY8BR#Q'?0\_:VB
P?XV &U[MB^*7->F5J\8 *(VW%JF Q9:YAE1?$#^L2O37@&NT]?A>]<JP%HZ5Y?;-
P=J:L@P_YU9P(8*'N&3)#(($/7=2 H:ZB I[OSD8!DMH?_)ESN-:. 'F3,DF#N5PE
P#A6Y9A&0JL]Q=>=G: 8D5N/1'. 6K-?E-M6=O(7MM(JD37-1^(WJ$KQJ9FHQ$MC+
PXI"L$\$X7$7;^V>R/<4"A2CU"[0J'T\^+_5VR535:;,?'B!_/988Q?%,XS*IQERJ
P5 ]ZZ\[<2A>+?U:&"S;O(M$@ZRKL7S>$IAH0_S5_;+Z0=:T9*%^Y%XQO,.+?S8F1
P1\9C<MHF>/P1^MAL,#^S9A_B'R:Y. &LE?FH(D=8P-&2P ,D%IP)Z%5F):R*/G9K
PU2DP3XS^RLC>S"6#[BJ_[8%%2@$MZ^96%Y*H% *!8"TTTOXI0VP^9S.%/H9TRMJ>
PE*$6G'3F=QX!.BX#>#OO)1B9$JA"6F5=H$=R.PLW\VE31]S"B:966DG5P7X\#[FS
PAY=%+='1.@5.C%&_C0\_OG?M;:#"V<WM!21Z+6%@CGCVO2,"!WX5!N=EU)^:$&))
P^YPL0D66KMTE0+@3AB"E\B_7.Q>V--I\DUZPZ+.5>P= CQBL\7\E'%T?D3)'<?>5
P%-$SX+M_+]1-1N:8)"([DVQJMM(/CBJ#.$A\#3?]4A:57GU\[5[T@QX!.=_I7^ P
PS44^@0\>#)2NN.(_!%,):]B)O@"H!'-WZF!W!I$-^C*EHD4=:9WD^F>)#3.EK$O=
PQ-O<W+S[3OX2Y]RB751K!XTGDCJD1PC_/UVWVI?3"A_BKWGCSY5>[C:'39J:J'J)
PO>D^^ZSQ@]3WDCQI;RBYN"/A*,DESHRUGNL%LK*\JKSU972[QU[*Q4+]O$9-#\!^
P^8)LH^J2E'+8][B*ZE/!0?>TNBN4IK_D)O0'IR8@RIV28LXA[U0A;FBF^TQW!1HR
P:#R8PI-/217Z?+DPD\JK#Z'?^6#?:$-*_'Z1Q=!$Q\F.0M*3::?:2VT?S:O_;%23
PU-&UB[AXO@X?7?IJ%D& H#=^T]T?QLRZ'"_XZ2@-?=@:.>:C-Q_]1H&S:>O$=2<"
P4YJ5)UQ;'M#YQ7C$,0/<,/3ON#_!#:2]+$L/$:K(#\3[JZ<MJZL&I9XR!Y&>JEC7
P7WS1W_Z+Y,.;F(-9D^F>LA!3)TBW0^@=VWG7M9B.WZBKA)8R%)2ZZ-G@,4268Q'Z
P9=(H3),(B\2P/QM-V32BXE"A(PP"LPDR=0.N+!T_HHQ*NLE"3@5/7R&$7/G!%D:&
P'D,0QUP)%B8YXQSO]BTQ6:4^B>-C%+$4Z[ U%8VG/*V/G53<BM]0.5(&"GL4"/_Y
PL@&VUE=8,7@R%JJ*)S),HH30DDJQ3!4)]O*:GZF:HZ?E1_W&#+ALMLS(TL1 8,9L
P[0@MF1QTGBLQ3R&XM$1=LAMOJ@!+ENB6\.BA!,ZPB$S^3(H-%EIF,XA3,:VWZDFI
PN2$A1&<UD$JR1^'U*]@P4/C!%GR-$X(R'?H\F>H#)D5T<C(WDI:H$(68]^&JJ8SQ
P_J\2FN)&\[\JD2G+_OQA.Y)G,Q \D>+Z'YH8]G3&9?VCLN/ :F]SY(O:$YV?O!=^
P6=^:;1H[3G<JWEX/.6N?M".Z,#FVO-F1',,GZ%.8>4O5%"G<>NM%T-S:7N092<B[
PX=D?<5[* T\'X656&:,-B?2+5(L;+K-E6NE^U]S7G6D;\,("]E6&CI6/ 1G88SX-
PF.Y'GSJROG5I&'6)4_#-MH"*(DXF&@+WZJ#TTTRNR_:JJ+=T?)H= <-85B-8RQ;>
PV.(N"UC"PFEU\K<[-[6"N[G6M!U9S>L(P#12@D& >SJ$[#\B(+UT<A/BDD8$M:1Y
PF_8WZIG'ZS$Y,*QPHD.2+==CWK_^T/O="J"A_2"69]67$%BQG7&'!6'WX5)SI/<=
P!2\)[A+NVA3NP\)LY.PN";.U^(4 M$4E+-#^[2! &EYV M+(EANJVPAO8*OH;@-P
P[4M-?V8U<0=RZQXX_3_T0+J!\H:?*\F_./'(\L%%Q* X?X@YZK;'@$IM;+^$W=,D
P$NJJ>IV%@[&!EY\AOHQ.%LD<<W*($ KMZUD%&V'>J^X;2I+3A\R&T 5-@\0?@K,'
P]H37XW?HZSG3&S_>@6#*N3 ??C5UR>0"EU/3<*LV_W7Z ) S$_=Y%ZB3*OLIKU!9
PX]][.(J<+Q84($Y']:G!1>*$U]Q1*(-%>D:#YO9E6@^X01SM TRAR96C?V]%W'&D
P@HC5MB;QJ')<U'1ZYAZ;.I3HLNE:;762-1T6CGZ;D.-,-%>RKMI"W)Y/[W:N*C5*
P4V>=:V5DY1TD_?>Y/U /:C-!8F!;DX/,@P>%/&HNZ(DQGKKZ";R:SXND(&;"#+</
P@4@%QLJDA91;'=""H/8[YQK@\KJLE>/U;L@ZN#[A>E+T_(+" &5NA7$Q[^\%(BG(
PO(A/NW*DE:ZUX:Q"O YR5>KYN/!],,XW9X#8_$O_H*7<&UUN 10,+$I,F27 Q;S3
P;_K"9K^X+VH5BN:Y8D.HEAQDOH1;/=F@'F,W_[N-!%^Y7W'>%>=.C#$,YKCL]X-:
P]S(/?PR(]#P'8W2B^]TC;)*NIR=G6:/VR**:+FF@0\+V3@@8^UMKX@]G7B&;_]9@
P+;20O&MV'(_R:T;B\8HK(=F7[3N5AB,_69(?O[);,+JT+A+8Y-'@&_5T#L#'3_L*
P-DN<(K+WYZJ(+R$D3'U+QCV- S@0GS.CY68*J8+GU4,_[5PFI'6*6T9,]>C/(Y5_
P>G,!36"BV1D6:)N@UB!S$E*8ZTM\' $YYR<+!]X5Y*:7=1_^0OCN_PZZ A5U<;3H
P;K+\#0@+?3;P[I^(VO7(O,&G'U$/)B(4>.SD>[F4/GP\%V-T^1<BRR@?H#BE]=!*
PNMF/Z<@NPZ[YK3N:LI<$VE^"]QE^>7QT2<^OX]*''7TPCE/"P]]BO4J_3BO0_#=B
PR%RO]RG-QLGXN(S[W%,-1GYN; X'3I=5UP&<AF!-]E9CPU/&3F>X<X>7[;'H8Q16
P:YE%Z,0CA+_F6VYBB&#)4]QYT=FA/4P;,<M0+9V=2_4KWS'5ZX^U?<<^#8GC(W.P
P4D F..8?ZJRQ)MU(O>B:,8+W6F")$;RW0(Z'6F#&M&+,":44RMW!SQ#/RTA 1?>+
P>6W7["V1#.2T9P?6R)'W!U'1R^6-[>$G=T C""H/F]D^.T20*T\X]A-9"('5JL#-
P*5^WX.5 !A:)6OS<P78B<FG7HHBX=VMI69ENL\479-U!AI]_ZJZXV6J6(=R$N;JC
PI:^=V>B:)0CODK0P_[9(@FS@/;\R$:RYCA:,YCH-Z2K];;"ZGQBTCP8<4T-.AY!=
PWUALW)@U>-51OQU'^FMA*3DZ)WIZ'\* ?'?LN\Y>3@$%+WN*P:AXQ$\$5?X@/'I%
PQJY A9R8J^:!P5X9^BK=\9^GO)25AF-DX>>MQIH82>O34)A6 !%7M!-[^S!\A^F/
PAZV:&D<85<;Z=B%%7@F_GE#(3H42JEW.;(=+MBR;H [;.31<R/Q[&S^BOH[5T,GX
PY,EEZ5+=0G:&_Y9!W3]'?.Y!3LWX1_,$?>$3CCMDO&I'8F;OWCKIQA=B8>I 8P \
PQ:<A4;Y?HD:TF>^39,)_V#OV$3TQ[O[[@0MU"\?K>IJ3K0MO*G6<[_R_-?S>V,3N
P.XZY@3 )<U'ATM9?-I.X("@ZPTC.SJ :]'%>'@.^^+)]LX&45Z$W/*EZ7=+/]%?K
PFW'0=K4M9,;:")5!$?T<=I< ;1+0+0?7_3E1,":=-$Y$5WL>K%SZP,2,@NV*]($F
PI5/U?1B\G)@+36T>9'V1KW_P ;[,['RV^.THS9A;^O5^WSBBJQ%8D=Q)X<+2!90Y
P]A?\!]8/2&6G314Y\/[71"V9W@Y6)%E%^C82R@(^/J^"AK93 HVZW/;5_PZW:B'>
P8(O""WRT+A#CPZJ>0+]<C=>9:-IDSX@[:YF*]I-BR,I1.-RF64.\RG7-?:_J!]/)
P1^OPZJG(%P1)?,H80VH44)LT>Q6G>G1%GM1U1RYN!)4U[21]*ES1ED=HEM/@2C9F
P-:& \Q9<KGT8%I X%NPZOEDP!M?:1NJ_SJ2JC'#!>@HIUR]IY0%*SG4Q#(\<N17/
PR?'_(.QY8CA8CP;U:1#)(_U=M%>8%A^"J8@\S%$X/2N>0*8/0_=W?AC\8K%S^VT<
P^-'JS=G+^DZY"%.'K*5*H&(&UY[<; \.: 9THJI;BRPMD) ;B*KW\D$M'NHH:G?S
P'6Q(2ZHI,@.5:1V.1Q"\EL\RI/-B(>_"RLV8IY8O'YKC\0F_U'SY1+$>!QL(#'_U
P\$3?: @]+,IN9YX?Q.1YJ7U_VL%?[U*(6$@17IU-'EJ7F;-0:&G'H)8NCG$^Z57A
P63W "',FQU$(!FTL%*Y+<UAU7A]NA>\\0$EO_I.:>7VN[NV?O&J)!D8SH@%[#\\@
PY?>>I7*MFJ'W&0_XUL<0(2R?$Q-N\UD+$W'/7RG07]#SQT*?<=2NNE:C[#?VKO>P
P9@"7BQ/F;U.Y-T>:?E8GD=60Q'_Z81\V1X4@9S]5(65TY7B&YE"[G7*WG'7:,M*X
PCD1M-+<@TI,T[39I_'PT<-+CX6?'V6:;HQC='PA\=&!?!#GK5<J%(N61>-)%+K%$
P>9GKD[7M-X?>.ISY+4]SMC& &SHC^Q]1RC+?=6MW-;PO59F25(ZHM]]M]#I R(>Q
P3?QBNNM?8/Q-F%'QZR,@-\@^D)NM!+N.3[A5BHH2H_PYJ,>]%Q=+_XX96T.M=#NL
P15<5&P]7Z&CL.K=9\NVO5"Q'::].T,+NO49!QS5I]I//K?7D-Z1DQU7XC(IKZ_H5
P>% -"OZR.*^=*!7-\"^ ONS*1\$2KEU [NC#0/4BDQ^7P<K<4OZD>59@3N'8\/#1
P>V.,<E,&P\:"&PDAOBN'(:%:W8*<!>9;FY(ZTXST,1V3H3,@.VWQ09,MVHKX,2RL
PF5AM[_V"6"\XXPN?6Z?G[GZ--DT(Q1[+WFEF51]86N<>PSG/]I3Q!:7337GY%?]7
P"*V*'#1DXT@N\9//295H4DW_HGD^T.V4A.;QWF\B/PFS;"ISXOLX5CP*MRZ(Z2KW
P@_]Q2H4<W[->DOW>U(<'VE5^-![GV"H.HLF.I7:&S)HBPNCQJ:?++1V]E#9>= <8
PSU.5*NLSC7N&"( .3"U25@@( )<BY*75>4AHR(V8DX:;*I*%GLP^" V!$D;9T8OX
PMYI&JX)BF\7-MBZXEJ2XLZBN ._N\O) W.)=\>8.GX4[?(#S>G\M^4J#A\\>!T.Z
P@H#67?2V:4PVY@H25\!<">;V=G,Y9[=7T\U3C3\;VZ!R6O<_=J4:7;1C'*#_9*%(
PA,.6]170.J)_/O^\!3OF5W1Q;;S\EMC8?V4+B*@TF1MWXB+5VV&*"65$RAVTR5SM
PE?D"3WK31^13U2> KE5QOBV?:MJ:HI_B#V2*C@N"6H;=0C[C'"ABQ^DU:R_+XO?%
P([90W.&J31+FG\3R/1,3NGIE1/]^B9!AS7"(6B4W">%#)F]*A\ _30;^#0[@(78*
P52X2RR$V>/&+O VJDCCR_+I]W$8IL95!.="HSH$BR3@+;U9Q5]3A=%"EIL]0, !B
POGU6=\76E;VOV2X\%J?/JO3+2.#CIHE]D]EQ3NX,R1OEU'EL2_=L<]/PCP&V+TCR
PL0WN!A%F\>ZW>&:7P5TBS.@568B1'"$;8-#RF3-;T+S!5@*C!!CB!B)@@[#CZZ:8
P.G*Q4TOV%P;P'J_J9KT$]-LR0,&[7(JI*+!VPN=/U D><W=!\N_1@-?K]+9R>7ST
PL\<\\"%UHK0XX/-S,4:(S)$.NV*B\";(72;;,<>>*]#\O$6H>I9"7QW2TB^""<[D
PTM+D#'[?Q6ZBCZ&/:']1I/;T&OB&FHL+8 I'P]R15E X@>Q4VS9V&MOR^R#R>ND 
P)]FLS< &_TT*B<"P\FA.6>%&MA\D+J@I/ZIO(8ON,<1X6OK.*+L8=M/.F"O,VI\"
P-\SE!0Q_NK).3AO E.]J Y. X4SCESIT@9Y>6<8!55V<6R;;Q,$'*M,EDI9]6[4R
P\D2,I[>.Q?X=W;M!ZZ:L_@N.-&:2ZDF5AV%*/7TAF7:W",GE:LIP/3X"/HJ$*_O%
PYC_VEG,)=LN]F?S]W+_\=\QR5_$&.3^$8^H#1SBT(97Z&%:1APEZ%>)$DKGF&3A2
P<JN[W(KT^BU0/0%WQ?GR!#7J)9:("!GN@++=.\X=JUSM2U83O2(15+@1#31[\#=;
P=\XK63+!9%6'#B7"[H5W>-6[;GV=+3+*=:G,>Q-5H\_ 65BB&*O&K/<+_>AB>5RM
P-?(#+2[A>9+>'4%--I-2M16>/"VDD_2!SUTP3'7KM$UJ*8,K/%V:+N)JGJ_T"]AF
PV0*#ACE&"6TEED-/TYY,H(?1$UJ\U^GKY-G3,B[D$70%4K@B]8X84<B,4C+BW/^=
PRCE? 6"J&R+;F2*'&?P$X%:=E>"5$L27]9]B]G.E^LO;W$A@U(N96(SO=:GQ# <Z
PQ9-2@EE[>;R6  WI+> =""3RAW<*UB.C?IU#24PHD89$%QK7;L=)S4$#M3O7AR4=
PJ'7_V*J1L6EWTQ2=;SEE90^U+#A'.D4?^%$2BWLJ<770D4VYX"V[L=;9H'W;V%V[
PIP^C3,[C\/M9UQ'JD!YN%'M#M>6:IT4S;T$9P&PIJ%ZY X>Q(Q\4KD@_\F],'6]U
PCAP@QNF(V(F4,1K2)RJ:#(1004[;A6&]AQWT#:J<?BPON ?%,)C8U2O#R$W<CZ;>
P%K#IQF2?_3T_7O<&?OQXU\05!G]WE>(0I"33!B8[:D*)5'N2DA1@)>(518D8.'&T
P2MV-O 006PBP$'(*#<WS>*44/]HQ!$F<R^(+>N_;@/NY0$'QT0/$LTR:\4%[K0#8
PRD4;>LUZWS0V-[Y ;PD=)?MWD%ID7Q=@>+E?I=77$)B\VZL0 UQC5PGM_OQ> )T<
P[)\B2&"BB\E!T7](3,(A :"V%8';J$=:WZHUZO\.6K=#<U ?M_(VRGG+A?\."PZ@
P=].HBT53*&)TWI9,CN[_SP[Y-_5(X7F4Y$;7KLB1T<FDX<0V2M-;^K</?+W??;Z+
P!-(DZ\&W^A@RH?8@<WK)7-\Y['R.VP?F^/S '!G)"3"JR2$C,^D@,D.?P@W/XNC*
P)8ZV6=-X$Q1(N,?A/"UIS^3;F5Z(W[&\G\&K5*<Z]D#W=?'!&3_/%" YK$D"MT0<
PD0-7$LSSZVT<4BK^T3_BVA2*/S+-3Z4P[C\4NJU\+=^%'-7<U8I5%=1]JK;;[,!Z
P5N.6QV' [+8&WI,\%U8*UJZV$0QP-- UW&E3A"6 %#>Q8SU'QR*2\WD208$?OXTM
PE:8DX,Y@4._1B)5>$]!9)NSVU;[620QB4 WBX^2[OW"HP[E-D&]W:(UQ4 ^KF67A
P!]4%CCZV>(ZSJ84/5]9*B[+Q_E\"MN'O'(>QV\[G,0O5DES@!1AFD?#;4M'+#+O4
PZV:[!(EX)X$K6HXKZ)UD>N<.G)+^1O"UZ^OO_."0JDTZ*$EULO#&>6#MX#N58X)M
P)AAR/S5)I(/D6T)9I>N Q%)I,7K*T?H$?L7DYXG%$[V?_DL>;C[):0,7Y%;BUO,#
P)(KQR. +>)PMT.U.A0JC_-!\;K[!?_XJ%#'KKW8O61?G.=$4BVS1>^8)PE;$(QWP
P'SI9#])"TJ!3O*+&:R%51KYY[TL5./ 7.&L:]]QQT8/9^#ED'W@"[+]H9N8LA=4N
P)C?,FE! ;ZGBJ@(/">X'I9EE[L8;HD&TI!4OP>>>#XNY.871IL$VRH^SM3XL8<E(
P4CO<F@,U!F(R]8.$NW9AO!\Q?34'+M.PSUSD7(*3;"/-(3\A&_/?G)%EY4XSV]A.
P'F2-9.78A=-R=GT)%PFR,=74<&UYB(E%3%-]R2_P*A:FV7Z:W"@X56.\"3L/T/7R
PMF?H>[9\Q>MX<?I1BO?;9/CQ,"]>#-_B0C^6SD-<U^@:+BR6:Y8Y$CXM:\21M$;(
P#') MH(&?O?Z(;J]* _[%X!#LI9!B4Q3PE&V8T2M(&V3.W*ZK>T:3R0) S6O/%P.
P&=1/D8/T][Z)2L5-9/2W6;.B_Y1A,C]&'KGQE50@N$GI@NYEDY A"YZV_:AL('5>
PP5)%46N2*UC.=[:.1]^WD_GD<U:N=$17 /RB-:&0LQ/+:AA\^5SY";QYR7XY=[W.
PQ!FH/<,$.HT59-W>0:-=6G6=.U:2@P=MU9AU_IU8N]&W&T213.F5]*&TJ9APH#QO
PL(PN)IB[\+!(S:FJZD(]C_4E@!TCS%;!=S;?L!_3X%?$&&L[&H_?(CZ0 MI+,L;R
PIUBD/ *2-Q5"[N"_*]:>=H;(D]H /FN2LI>(G'>>_6-K';/6(S#79WR5JFG\ +\;
PHHZ#59/$:QKPQ;@<X>$#;9D:]<FKC";+DV?J:/8U?_V%9,7?O\?3PEG'12IP"!D7
P0N)\9B^EQ]^\0DBE<FWM7BU1K\Z(8%G",W@\!IY5* 6MFD8X?Y=1;XEYUJ/1121&
P5\P,OJ4" ):KD&N3X**C>]J0C3VJVDE/^"^I;BA2Y_P_1%A*]K@(,PJ]@8-VPQ%<
P'V%8VC!G)O0G#<;$[)D$";9?A(<FQ-$=:*94^M190]"L,"@*P3!8>/,M+Y\'8QHO
P1:=_ 'X5*7;PE$2IH./".XDN)JI,RA"ASL\'(N]VEC=@FYF$SB]S]@,4E5=<R\).
P8XG0S\*-..C'B50+M2"VN/4,-3'"V206\AV5818*^=G)HK5;A,_I>U6C:(]&W,EF
P&(LXP%K/*.S:SZ?O^=S>ZR-J"+0O^CUA)H:/YJFL$=-PX><&E]V$6X\CI?)0'ZH(
P8]YVHXU O9WGA* >%MW"KQD\:'=:9%>OT9/[?[:)?I-T@-US!"3(.*Z"*ZRV/JC:
P</ AF:,&O1KU<^8$W)8$,AG4^(,66CDRHX3XIET3)J:5P-G.C)$TV2NR!5)3TAE.
PMG IQ*8\K5*B0'7NBVV))>>K(46DT;VG0<3/=+Q0&K8 2L.;P3R>1L0GT_I]0:R 
PG;OUEH!'J5=<$!H7(=.PH;L(WV'YBMAGWW$&*RI$F.^<,@)3Q5-O[H!Y7#4$-1;6
P;H-8V1)XL"SZ'K_!Y%RXV]<0[>F3S5"]?.*3:AWN7D5W4/<3#N 5LG+A; 3A)^$(
PT+8?(8+_(?99D8\Z%R)D]BFV^=VG= N#CH[?KIT;\U\L&\9H,C18OY9!_>.Y^SCZ
PT[-[Y(@N@Q$JP6)%JH(90)U$!8BWPIS0"RH!C)/H<M;^C/OZ,&&,KYO'@YL-I]S:
P/S,<:V4P3'(P?C&;BR)^VUQ@N2=L3DO>)&%S;BS&+C2B^Y<F]:V=L%GHC*-4>T_&
P2)#E8GF2K%Q=WV1E@<FPG7QZBKG\*_=7),X?^1YR'&%6UK9@6^Y\^D6,2C6?UQ-X
P\1N,C\5RG!6EHW ,0,I4/*+8?0G*SB,G$*^.XY*AN8PVUT2X6*KKL/ "9C]VA-9(
P$Y"46>)8/,Z%O^J&S'O@AT] V]]8X+.P)+Z-$V"N#!&/$Z%@X2=U&SQ0LTMZX/UL
P1/IO+*B)8"N0%4WFVG]NU9AFLIQ_)_9C?]Y_N@O][?/XY4E;;ST4/Q9FV/S L;=0
PO& ';\QMACX268Y5=%B;.]:6#C9_09T^]+E8>3+==&E:.W'*7$4@*MC_>LWV;DYQ
P.[S/[('21=/LMQ.V9:M<U"R ""O!=^O-'_L\0P1W,<W89SJ( "WYA46$U>[?-F 4
PV8:HZM@+2"IK2U^)D-H02T,@H/G>\;PND)B\E!(8!_K-PY8ZI@UT*BCLN2$?;+1F
P*)G^"W#MD+PGR%UGI?9'5GS_\4Q"C*\-LME%,V;%%*JPND+:QP1>DJ:0YF?.^)1_
PZP^<SGI#D:M9$K>W',F9,>;WZJD)S?F[-*27G]$/N[Q(-6']X[2D!&U,F<]F+;X_
P5$"<KSOC[U3F0=>!ANHM3,O-FR@9L"%ZB_I)^=YX'QA\!U/S%8!)_BJR(,.M5;=R
P!%#/VZZ ? JOTAW4YZ/A6K,H!:HNN@&ENUT."$W/GZ'*D,ZR!*E-!I??P![))Y #
P0Q(^.LJFB&%3 [Z2"[Y^23N@RI=O,Y2$EC.AOX8BC!"/2%D"BCY3/Y'W-L@[HEAC
P85H+[CSGN4L]+KZ8ET41B$ T)572>'E3;BL9.+"1[_-A5\189N!Z=W\0@@A- ^S.
PT'J6K6@)HDC/SL)L95^&DRW;T.<06_HOH&-13\1?4C4&&#STHP2'_+9DK7SP!0$K
P8^5_+1;9E<!A%#JK%@_C4S(]B?N<@,[@!]7G//"W4:'E#O1D;SFX&7%HWM]+:6I;
P>U6PQIJQDVY@T2(#LDW/W*(':"(N7T@U92V+OEUM($K@JHZ$4:)7TU#DUC8G;LJ&
P*4JAI]:X8;%/3R%@PA>_E+[OOWQ,SY+!85])NC_ <]_H/UD^!JEBF(23_KQ#'[J"
PR"CJZ&KSFJP5T.&X[1VH#@$<_;?CMF\6OQ?S.IZMJ<.6ZN.-W&&]ZE-8H)DC/%T1
P\YQNL%\NG&9MD\<S.N!;PN%+ N8U=:(8*?JQ!9&OW+[U): .J=D6>Q!X8<K]TV,>
P3R-*YLP^WX(%]8]VY6[_@1!5DIJ8D#@@?GY3S>AL%C?Y4Q71!#.3Q57=)L>,E&!Q
P?_Q1%H'*!,/]*F$IF!P^PZEM;%F+@?WPM_8C@:#U ^9^GZBR?(.28V):JQ//P:8Q
P[:^#UJ+TT:'A<'AYXJ+KY^]!1RY%VG3[F^H>.BGZ2@2"I%V"G&03>V%O!=/GIQZH
P%.2:Q_<2N*HWG!WM^!?F*Q[J^9S9F,3RI(O[%-R2^P!;]#NM*C@ES&B '"=4H/QM
P2.""^,;2=8#/3,L*.CMF][)66[IP90P]XS:4'S3I&,?CE2W4:R7(MU-GU>5M>K &
PJXWX')S0"/063&1.@&XI'%X M1B3>^P@YBZ.!&%Z3:$\F95W@%YFZJ[J@$-_Z,16
PQ E2@DK3C7A+&!O\5)I9<5'G&KVK'>U'%I\V>M,![\IP<'P)A*.3EMI%AO.\+8>)
PZ1KN+T\14>6AZ<PZT&,W6@W6*GK+:UTA.5M6;3[]LW\33@K3WJF>DY]CH$M/UJ6X
P[!U)E9.L4*9(\<[T_G@<R+7IJ+NY$FN [-;$LDT%FF!0GW9>-65D^Y.( ?RO6:/=
PF]XA='>HVI?J,\%YK>]C\:7S\-U+M44DK*TLMBH>,.A<.4BKG)#TTT' TN2\O Z5
P 5(4U^WH2K"7]I 'D6YI4S('Y*,2E))TY@7F2I9-ZN^6R+O)>X9=,EZ,_SU_+ '^
P=(8IX<F$.I2.TJR);Q+L,@>6?H[OZ*.0Q)]:HX"1RBJ!,EH19 X!K_0ZB2+9N(Y"
P\6V'8_)9J]<]< +$5!E9$PTONFY.E:Z]6(&5@>:FH$&>RZ0!0JB+#9J+^&[F[)-G
P8548:' 8Y_]ML0]M/>D3E=/_[)@@(0_[7T<H5?/IB/20?=D$C-N]X?9G"F[&="_7
PL#WKY5"7!*9^N,]SC,O"JO)CWV8JT-ME6\#.T%@EJ$?[-H&$S=;8"5=FR)/QA0:&
PY(;?.)@V:DX%B">QO3RY$>H*]6"F6O+Z4??:<(E$%C(R=8(**&MVC]@M\*E]3?%J
PN559'_+L1@0G=RL*2*M% ;6I-X,VLI\Z?-X GKFY0=FS@0:8)+K*X$[D0N)]-D-T
PT[]#J6[V^3=-BF8=0YL/[8SE2UZ>:=MCZ>JTP'=FOC"M!E]6\]S==6-VG(O>?BU8
P+)6*$'D33T["3"/JJPN.</ HB+U7<EZ:$E'SC JT4"FE^%?%G=^B,B;022@\H%,'
PS'%C\(-!WX6,*F[4%>%%)@LW'[HI&;OF^AW]4W["]Z6A=%/&M\"$I-!BP14F=O_%
PX!7V?94OFE:59&6I+&^@A3;1)'K6 #V7:/&[;@G"88XAOA8+Q*5L;A^C9ZXT36IK
P4:\2K"*)3FB^M\NS6591CF61<(,2D8;964<@8H.=T*M%1L^%+( (&ER52M<,OJKQ
P)[R!^.CL<H<\M66/B=7R!;N[)5XZ/SU9/%C=%$ZA?N#7.EW=!1*EI"67HIY.A^QW
P[3.'IAN&"[#'2#'AK,MEWKS>-@2%!-O!ZPW_J37;-GWN__\>3@CO:%;Q<YHI^:4!
PAZ3>$=;]V>-BI!4?Q\*ERNWPJ,:FK9TBJ6:#(&6,#RK1/T$I#K<]V%+ !0T!-FHG
P:OJJNL+BKW5_#6!H0QG<\5S,BX5N3I:+-0/K%7D3L5FR7UNO,_[0%V/BP DMV+RS
PUEQ J=76<@ NZ$IP0L*G$,"K',W=G*/2-WB*6O%CI$X "$.0TT%']):QC-9-75GH
PVC2<!\JL,:N7E/C/+,PF,&>JLH_\]UFBMJZWBA2[M:66HL16.M2#&V]9,_0XY@]3
PW2K'!I'$.2FI(&#,@V\N;L:F$ &<OG:N43IO3]9"M'+I.XUI7C'-LDZG^J3Y'8!#
PL?F%Y7OU99J9W,A<CJ^"K!C\% -VO>[$9R_BD+8?MM8^BWB;##2K=TI2'#;"*OWR
P!P8:>.L/#QX:I 0.$XE:N,I$7?^*W@[=!P^38Y>JK-W)FH,]*SBMT*B3 MD#4@E*
P](5L;<^F==L_1$<1W#.25DY1["MOPCHIU!2A#A?NG\M\.*'_(6^#U(DH08K.M2'>
P6 \C:L?]L[6&$KK\U-[.B^GTU8JF]4% OC155GAT2LK]DQJ<!_9 \H+.(VK0(KVT
P"<B-\8K:5W6@Z^AW&4;O96+F9*7U&&E!JZH2?A?NA03I2-9D,3JODC,=[1(;I*N;
P$-VD,!?3=IF C]^T"O-Z4:XL,JY.VFO[#H9$Y?%;M;OZ0#"^NSGJ8V&O<92+KL$T
P GD[((&*M:GO@-H_%!G#H7LE';3D+,I!7T)"JU=E"1U0R<HZ:X)7.-<W0!.ACU+M
P]5!!> D5N.O1ZE^F&#PH =&NFR!=MA=K6T'Y>"OW?(LUOGT3/ESJQ56];5 :[W'^
PD7L) S6N65YZD3<<RCES(ZDN21!CIJ8@E6>Y+%[%\]T>J#QQ7,Y0H>4#Z4\NC[PI
P:%G$7%=@UN6"_*Y2X_?I8KC8W]&#"@_.Z?S$J$MKO5.6AGLEL@\5M<5P.3NHJ'"W
PB_/S:Z029A0?1-\T[R!D>_!"7JGC%=_20<]R\'4I6POF*%G5VN:3NN J-'D;S?>9
PU-(MT^"30"-)&L"1-G(=M"*OH"=^1NWOOB_Z8T74BL1[PT?$]E?UC5@/]5<7MG+<
PDA&<T@[^6_]]GE88VAD4!%SP*OQH@%2_/W4_;[/)LS9UW+L($9!/Z/VX:Z(#=AY/
PRX'30V(P78QCAMH> ]&!2D"I8^2(I)/VV+<TS)7",M[DOAG%P:;WN#QLTD?!]-<^
P"6.P! $@S\>Z.(6_\HC\JP4AHQG<;XJ=RXE->Z^H\&_+\P\"HN5/WI-U]([Y).&'
PW"(X1INPWKX*K7",^D62XEM?_(<T'T<,%>[8ON5CJG)M4=>+&S2)<:VH*":K4X@_
P_-<'KA8I,,, QNN"X=MGTK\3!(BB1W FWV9Z3/&_7'*=E[0Y)XXL2(;G O()!%_2
P=%>=LDS($/2&BV1XI\2VHJAF&FE]M*)DB@6.B'@6I(W5;S2J1^E8T]?U7R L![VR
P792GT=MY<G#0M"X,AH+@.7,7JZ.X">!8[69@P+1,XE7XH9DN6*U7_IZUS6N)B15\
P JPO=:O0W-,=.&;&QHUH5BHWNB&D6AQ9[LG4C7]F:X>VT_#, 8162LI$8JZ_J/9#
P7ZIJ@:?2#BV;>G_GQG=XSLW1IE'"8 SC[R'F)0HY1P8T6DO3H(R6P!7<.']_#,\%
P6=SH9TXLD]I.LEL[NWY7WD46U]W)-MI08;1NDLX(6)U+OV%@P;DC1V*.\;M$;[7N
P1I)J @[J*)[D";[<.D:G"=G&<-UXL2=UX0.\O8JQ0"2^7L$45+?G/'6P93^;_#,H
P^IC32OUIWI")G%56?&YA1$JF+(@I0:>W(FO1QCHVF-L3Y<W2\^B]IY)/,_]I02XF
P5SG!%TWL-@%>)#MJ0):B4F#KGM)/?/A&*3F\F;/P#CKGF.(?,%V]M FC,&9<RC>9
P3ESB"<9)+%0\81QB9QI]Z"LC<$<A]QJ*&)=G5@AX1Y\W2+]D6ON?4# ]B.E.J^2)
P0Y6MP17%-S?X* GPXB?I%#0JX.:TB=7O<E*FTC5@-UH9FSTOW]"&]O/JEEGS,O8;
P!B\9LQ5X,N4>^RO>?+6PT?A>,Q]<6PLB\'QJ</>T?F0C!O6M;#S,5X6@2=<OK^$F
P=>W:7"^B1VH!T6-Z1"&6%]W*?("""DZSS['#M'MST9$E;0'URQ<!<B_4,K-7(PJI
PPVRS8T. SYK7M\&[H%\APETLR[!WXS!B7M3KHQ'M5B=!63X9)"^ER^I #;#C)Q2=
PG/T5IQ9O<,PPTRXR,3&,R7(ZD+,,7U-P"/8X_;LZGAO+6HI-/J,,_\:\\$ '%FUI
PW\98JZOVE:['ANY0'1;9ECIU! !@OV'4A7G:;2I6CP]0!@!DO!*U@#/L3Y""$1H4
P)%3:3;2#%B=X;],[C""#JT;?@*$BDC1EK(7DGS?Y1C,]+%D?(PEKK*TU_5A ;#RW
PV </O*9/8]F-(V:!OCT@.W.S@S!WB9(>A';]]O*6@WZK'>U@B?Y+GP[8!WI<'OZR
P"*V9(#B5$8N5[P/D!QL+REND/3L\S3:GPJ*$#Y^Q$5)2:.'J8<@:QP 8ME4E1.O*
P]#'X^N+P,\GDE4!-;:^(F'NP3D85=/#@X*KG6G1S-:#!^Y/T&:DB)5U]OC<6YYI$
P2PU,40V73Q ;"*D16QQ,A^#(!3*_7PW6*G<4RRK4"8\JV$C'NRC'C)\PT; CT7#/
P9O\*;@F ?=H::R?WW1OMXBR6HW (V?B7WQD=I$08C5*W))PDGL,KH_5S:QH] \L'
PUR %^@[1=&-E]$U$=UW9>MIA.E9+')8B3,:YOVD7"GQ7E!OYP(\:RV.+(TTYBM/#
P/6)L(G!39T8)/<T&(M<0T0.(1LZZ?24/$3[XX)Y.OA/L/]':^&J7]8P_@45<5LGL
PQ;;]/UO99,*Y&;*?/R#<%'1>6>=7/L [Q@*7<C6N<HP[IGJ6>" /61S)/J(Z!Z!I
P@#A)XT*#K-7P10K8DBYQD3W+2H2*G$76,H1TRK.9 [I \%0*&'LXHXXS]1R8=[J-
PI<_U&:4: W3UK2L$/JJ2=BIB)'R8D$'I>/Q@J0^IP6"%]3[9E\HRH$FR5+__6U)*
P^[KD'OC/1G,$0%F3?SIRU,L$:4-!XDI[_V%L3453<^'A>"T152!-X1_L"M@>!+;T
PXE:B@E;CK_HG?#KU3)]J+\L@''?->X''#^,N[V-Z1"<HZ(#\O3:=UI-P>I*L^"1]
P*R%=A2B'I'[VEK^$ M4+PZQRF@GFY$#+7NVX.0K]?E/9T!H-EIJ (Y-W2L[7@O*S
PWEZ?P@/Y*:M<TT!A+X%=IS3%AX"ONFAOMLWB(@!CYR)Y_ P+O0S=Q)_LS'4U?C;?
P[24W@NUM!/_U^AD<(Y'7EJ,)93VJK_JN)-C,8O$R7"G@V6CT67P/KKE58]HH?X]9
P^ED*E8=YF,5D/Y% ]?OU=\>7F.!*)9NU.R_V=>P\ L)>:0H%TX8]#']-KD-)9&.I
PSZ=SS-0F;(7+9KVQ[<5:*7_M:T Y#V3:#,$J1B*$>*U6MIC!**6YDI$Q\">'Y=7'
PCOO!,  /;!H#L;J[]9,T1W>;N"$SGWEN@N,2@)Y4@E>&OSD]PD&3(/!4,6W5*3MO
P3*F;_>J-ZB\&B??.>;S*+D;K61P=2/4^302SGLU^G\;<2W.]:+ U&]F<$_0,Q!.D
PA5;4)!)Z7F@VW* :PW"=\72,@LVG8Z0RP=XO+)(2D#*_\THBJN8U@K5.9DQZ3>"\
P;-7\&2PPP(%\X$"+XFL*B(<#F1^\U#RF:M$TPKAT,AM('5TZ-GA]==2_N+<*B'UH
P<Y.<)AX-H6H>VZ[I-)8QWJ3*+!N2A<R2-"H(^'W4YIA9.M$R%V_XNQ.@8$2F.].I
P- 2MAU^IPA BE2AYWK'\%?V/YAOSU6/"E_&XS-#WH^0:[= A+;Z?L?>-FZF"0B#[
P27ID&\5,-2HY'WJB+00YP8K;.A1.@3$6G8E_6^)V,II[)V,% =%X@6]B4H[17-PS
P&7-X:/N#?,533(IE>ARIW.W.OC;.4)[2X"3\\(:N9"2BF[(P1'FLV=(/8, U%I/N
PC<H9\D<S%CGG"?;'PK#%;OBK!U7[7M!+%D%D1 /BB%8JB;+!,,>>N?JVMY'/TAP3
P6U2&3=)@WU'0"J4" Z\GYF:5<<N[/ Q^03.XCP]N0[+&=_X17'(,@9+LR:CE7MJ]
P*)F3DA0VBKB\$E3B6(@@@NI-:U@3O&7E!.9":5V903?!KA47'3XW3^M"^-N'"V]T
PY<,)<-M#!_JMU]A0!!M *ULM-]\'V;N:=N&>K1X&T]F.K.^C@K1U;M#>X"PEE,BP
PSH%>\<#'88Y$X_-'Q,94[8PI"3]JO#:TO^JQ<<<F5T5). <@:I&,!<%G!.97?:DY
P&.)ZQS%E:Q6LK0;N#EV$,&=P >7$YX2O.=STKAI(JCJ3[VBM3!:_X5*%,K,A(9QH
P%<GF'H0L%]TKZM.'W(W>UGXO!GV.,+=RQ"V+;BJ04F=*9 @#3C)FF>7^!WC6>'P\
P]'&8^"6+G] WP?R.@ E<$UFMJXI*(4N9.%-,8C< .?,X4XKN=.OMRQW2K:1I-(.V
PV[?^9F=;ZVTHH=PT$K(?)5)+[RZGGF;O_45T!WI)3WU#R&B5<OR)9P;:69D9;F3G
P35I";<[Y#GAZ-)?RI/;L,)DO%27;FO(B[?;3H F*/K.  2/>Y3.RLI1.14&HH5-Y
P%A +VPY)5<0@PH:P^J94N=&%5"%[A8%+V#81)E/'@]>1K&X[V@[VQGLH%<;H:6.'
PQN:0/7'<1^ET"A)99"@?2Y?S)?UGPD$+N5H^ZNMQRM71IZ]:>;3T8"C'@C(:LN]%
P>A(Q@FEW#C.3:U_EX9=P&R6SB.\M 4Z,YJ7:]/O%NDZW*-Y,E+R-Z;H+[;PC(X9M
P\$ [8X\!M, GH.[<+D^3ZC6%]4:[GQQ 9/:Q-H72?Z*)-I":J#?3 ?*]&K\'=C%6
PU:CHGK"@<(^J!Q[U;;/F(N!N^QH?[@Z@E%TA0YPCNK2Z"8:/M'M$;*Y\R_+7PU !
P J,0E-T0P"G+*.47/Q/C@N:$$=B",>-$E_'!T7$".,&Y@QO;]]7(M<-CH)8MCAW 
P7]*\LWO5LQ7,!4VA2]U>@-)LH1C\B&0-Z,Q+L[<6 <-:<NPR"'P^N,ZC%$HH-!9$
P8O*VW*J7:$EGJ\%!]*L C 0"ZTGO:K-G4'W(*&6D13I2G=X;[WZRP\ )(T@H[6;Z
P!F_=EYGSN=_G4F.2>F6VX%FO%WXK %%HJ9+CH0M!4JHHGW5BA8#OOL ?"YEZN3M%
PSGKLQDQ?BS$PZ#O8O#*T(^54<;'M*/-U!ZV?B#8JIC2+Q5%!M19I/1K942 T\7%H
P5*DC2H1HXC%F3M!<.C],F\J>RXQ0<].Y4TM)-#J$,W_>J_D7NE'?"9ZN8!L<YDRY
P/TFR:'QIT@OQ[B^D'<&2Z%7P:%\1CDUJ,V*R)@X/+.NA++WPG=C'3Z;R8?]HPIBP
PN/XG_K-B%_29'<JPY%QUV,F<*HT#9O0A#Q7WQQO#9K_Z91@*,]^UA9L-DVMHICZ<
PSA 0P3W[1ZYQ29#,EXYU=EW/+F.)1]ZF]"0U/+:217X2L*-8_'/3MRQ[:X)UX+R>
P<P+4H,9O)CB[WGK]T?+:74<'XX\R.D5\D#?@SR>>7'Y'T3,L(,7L%(5LAP:$T]S)
PL)PH"YRE/>HCEM[NA'+4";?F_8/!&W\*"4Q*H?]2T[SHG!9]!V(@%L G9PEB+S?A
P,P4^BG?RU7Y4A)ZC,DC#TXX2^A2(%0,L0?2O&V(-%7_]N(]9F&.6NT6ZT92VE@4$
P9!HQ)K#6DCNQ2#,I"G)8$E;;D#W OPWH1X=RS8*]^>0G$Y6?.LF!3O^[[1.A;D@&
PLAG$DEO-TYY8,XL5R((4-[IYI-H0GUY099+"#)4P(7_U=UC^+L8K%*9>0QK3J'TD
PV6#A;"D%P#I 4"6PBX$%0;4T!;_4_%K>$*PBHUN/E!T/X33R_$EL6.1^/8T)*"=$
P7V-WTYS<87)ULW99?2'%2]D1^^4ATY_")[H,Q"*F,U0AQ6#<\/L[05/-;4#-:CN:
PJCL%*%DA%G2-A\;/0LW3H_;3-9S069O4IDY!",(@0WC.& +S?CN?"8I=:1+"RYWC
P^V/)N.P:Q9C?)"<3,&6)/7.]XKR//J9_><)$ N@[U__F/(1J:0GZ40J,:?R6J=E'
PWD\]1T543ET03I2.,Z4N+\C% <G,&?#R;BL04L4]]&9P@8X-T\+>%">4S"N^ID*8
P=UPA=#P>0J"ID+Q#(..SUHA+8O9>$-4>Q$H1:B&$C]=='%(PZ^^&5\;[;HD=(MT9
P+19B"$5:3@"3SP.S:MYZKD^@'@B*@9: C:V.J,Z#T@#R9T;:PM03C58V/-WM@HM9
P15,:"./[9')Y*T!%S<(UACHBMX!^[]A'5E#Y('=@7R(>QGL9O"6W879C/WS6MO&G
PJ;=ZX1W 8]FD( O*(];D-!09@3A06&SIT6DP)*:@[!GRY:B0A[M;OH0]?9-87V;#
P<J]L:SU_Z_(%@701\;$/7@RX/RHH]6H74++(C%#-:$T<Y*O]P=D9W;M^=#')@*=C
P0!@D @ 4O !R,X(TG4^Z6_9=-GC-"@]]] 2K6Q*]+!%5GZE_GU*)==NCQ4A%^D_6
P'HBIADGO^]D'^^/_C$LU:=O&4'T_- 0ELO 5PT:P. F_"VW3R=KN=1\T)6')S1".
P*[U>\L."<#RLCJXZ7E/17[)[3NJ^V5%AP.VV91O=$S)>8&7RMK'KW^T?=>6Z2JW6
PV7[Z<1UDDJYQS9Z\UUN)KV25^;(R3[^X<DPMEJ3<U6&8_@$B@$CF 8%%@W-S.EUJ
P0Q)[+,8;05DQ@IE;OABL)R4S?])Q:/I>9J.RI8*&IA>UY=7AE,W_#X#X"<T[?O5Y
P63[14Y6@I=O1:V[6R 0Z6V(/& 0M=X;<1\']VL5PX1 @V3Q"MV!Z3A/'JSB,0310
PSX> #;-(X%:GEG]VJ[]L 3OXU%J^#4K[VDEIF,Y=C>)7[K\YMYD'"WMB<A78R\W6
PV1K+VWY6,3%_9BBC95[74E$K4J)1NNZ:^6<%+[T=S2CAY&9LT^-Z-OL>KAZ+U.&*
P*C_O2BE^^!G@%8/$3K3+C00$YKL%<'<PP41G:[Y$J]>[V*V^KN 'E+&W#"AR^4"V
PE7^4T@0#J&(2GU3=%CTQH@+9?T&3/?=Y__E-C\0=I71BY><*/>"KN4]VA50^J<*M
P[R6(K].Q58?,8XI^,1TJ,@WP5LDNCUW9-S70R R2T>IZA-^1-BW?S[S@F&<"C?VC
P(&!IMKO/!Q,$F2"%:Z0)$HO3/44-H,$,,CR>^R6J/]R%PK>!'<::'3A&&EH37>N(
PFK=;\8T$?G3#LTF\9T5*MFIVZFE@":9$\L >0H=&#1N(K0-OGS6GRC0-FJ8Z[FY3
P;U^$[)W9-0 ['U/GB+B+N+AMJ>=AA4\A&P(#("/*K#7W4*\D(NVT <UQ3UL5/I50
P:MBKTX,SS"5"[)&L*);I;Z%3\-04&+4TQYJ'_H=.\)*ZPA%VN';8*N3>T)E%X9(*
P3Y'7&KMI7O6RN*#WB50[<2_>LE6U\P/R$6!@^NW^7TZ9OY*&"7?<4'Y["8$%*=.8
PHU/M(83'<]Q5[DWG.B<,,'6[[1Q&<EO^!:!7L5L4L"PAP7ZHK]H3#!'AJ-N$SC6T
P7,A]_T,\(*<\R5Y5W]&ZM"Y4>MW"7RM(@_VXF78*CY;9#0+.22<[8^CL(;Z_(>QZ
P":&Y[U2]<-JMC65KLR#OD#8S0+R0\ID;NQ?Y>>H*H2#IC'O_%= :X5[#*::_$4?5
P.K_K;\SN4V-Z\;[3B+89!I&Z2,X[OS1#=GX#7SS7RPQX:AE.G"$&-RZEE/:&,(RI
P[@J'DP_ E:0Z-V54@G'-UQ&;(7*^$1J5?PG/:_[T<T"<>AE?*C]LM=S>G#C2:*UU
P#)P6>G4RP;W?Z.TR'0?/Z1T89-;Q,[,1HI7PY2+.;AOTV_8QUCH](=.A9.-FR_X$
P6$\;<W4A<8,S=YEZ=R5M-@\ 4MD+1.W1OO@N5V@)Z)7Y)AUY_G/'9!C%SF;=I4Z 
PSV-M>S>V,X&]>/!_=^+_?O: #/%+2GZ!*;7F 8.:(4&[GGE.)8!^K=<_H*(1%%"R
P+QY>X^SE@I%2;;E/?MYT$5WU;J5:$I4IZJ2'Y@XS&C&$I&GP.B31*5Y?7*-<_)V+
P;"*N#3%,ZNC>'#2980K+'<FS@H^B'A=&LZ68(Y2\C1BF3;?:\1!I624E_C,Q!:P"
P/VE;U5>W)[#*@3I$=;V?>XT+"8(U24#\E;#LN^G%>4J65@U4KBK2"<+L*O)'?#,/
P11J(&H:03V ;FF14,9*!> 2JPDOF,.@[[ 4Q_?(W>M";3]&0GQ7_S\X8X<?& WN7
PY!:+$R (:!H+_$>/H OI:]:28!IJ'=]F+C &4/2+:6O;< :Z'-BBW'F<($MMBBZ5
PJ%;$W9W0.)D8WUN,)YG"M\#ZU'[3M=M70@YJKXK>Z$;0:KW5AV;\0^DM$!8Q&A?2
P8"#E'!HB <&,J8$+^]Z-)=$WXAC^A_A2 &@D4]9;EZ1\NXNVPF.#XZ!_N.K@6(C%
P3FDRP*XUO?6@F"&N=3(A$/_A"\$Y1#L00V@RFQ//-P926?U_MH<LLBG3#X<GE2D5
PD=)ON&>R2T* DZ8C[67^G\19828.5>4%&O:BQ:C86_] &DM=?<6GZ-LX:8S?OJ"I
PQ/2"]6+W@#C4]. #NGFK4P'/D7$MX&+PDB@;W^T7V';_;B;('2.#@.(-' MA^N68
P  2T3ET_WB#W&R$N[6,9H>$WS-X\M%;R'ALH8\ <^R]P ;(#IT/=9*OC9)S 6FG;
P]M %G,#LYG_O$[-67-X&,JG[F+_4,"J)?YKVF)$/\Q\*QRQ*;4X!8R']!;V>UO/H
P-R&D%]=8VTI:VBS\:X;>#R!GGOQW$C1&/0)=;Z[FF"[A #%H"=]I)6D5KLZPIR@T
P O;.G0-=K70N4@^4[\,%"@MH!]X%U70,B+TM+=6D!UCK,RATS$'=&87+DU[UEW:;
PDC:VH2G=N&7U+4<L!<N00^*D:+Y;1C/$9S+5: V5%Q2]I,)\A+()VM^SYLLQNW03
P'< FN<<X1/&P=+0W7@005"K L@5W1#IM(EDNE.7E !(3Q#\DQ!%%K]9!91J_+\\#
PP163Y3G)9\#Z^?/S'1V1TMO'?K&?T#P6\+MQ*BPX6DV"V!Z]/ZBTF'3X*"ZNC-U[
PP[#I(+_6 AN2PMU0L*^)5R)^\$X=R3JII-"199:T3G;(AM8L)'G[1$ZI2%+*:D4V
P835\6[K/C6;#=QB,GJ"IU4T<[C&)_M9E#2G(+>TCH [W.X9!OI-)L_GFJ3&47<7Q
P!<L5NZG@=Z&Y^5D*PIXJ1$<W6J+_S@#MJR4:GGKMVL0@GAP,RP =@6TLY=]$$6_&
P!1T;*C[<_D/%:;*3QHT.\JD/L>GJS %]_N0P^&F_"[[W8T=7W7ITM>U%8\MR?YDQ
PAC#D(5%O^ HI1FD[H,DC!V]S.L8O-5'K,'+TNCW<7:F/QQN1S8OXH^O)=Q:X[\)$
P@[*DL?DXRE]VL44:XC?I9T):N^A,>5RFE[]\+<XGO8*T?F[9;[V^-)^X9,]:>'<L
PT'2NW]U<?$B7T56([&QLPJHTR@T#(WQF'X$X'G^"CACF(%AF0$S6!SWNG7JNOL0+
P;&W(].'(50$N:P.X&;WUPFD.]<FOE7['$J5Y2&-N6G;BOFXO+T@"LQ6:Z+%[QS_%
P',BPUD19)$>]%<7M;67(;K@KP2AD,B?R4!C#=:;1KFBH.G]+O!?ROH$V,ZDA,-W!
PN=G5,L1#]G+YW N2A)&B)D^8T8-;(JF>[.!//DI;$$%RI<"C4F@^%86V(Z?U1$$K
P6%=V*%'3O^;R$".N,^<'2(>GY'J8R "T=IDW0Y#ZR\@BK@UDQ_!87U[9WFQY06?'
PE4XXV; _):L+R@"(H9@:)L*$E$M33M)&,CS3R*2P \7]V62TN<G7C V?QX"+Y$@K
P8HCS&_P2</ A2Z#<J B87Y,*V;YP-G<EF!"Q(VHK,&T58;H0;>VJVO/G[^?VQS$_
P1PM[B*GTBQC@@.$ZUX6&S DR 8<S26M,%]+QGZ.45IV)MG%V:2R*N@?4L8W+M!QS
P)")AJ.IHNIA+;LS.TRPBT(+__J85J$OZ-73"O=G75C^/^]"-!;SHLHDMF\.'O#-=
P.TIX=G^E4JYDQE"'/="==3>",(W7M]04JIRX@#=9:Q1I[BGKO1M)1N/K7![ L$MR
PMENC_,_3!S6*8R7LG$ 7T-LZ-'8#>\!,^H'U(,+K[[\#[\&"\(VG=(>Q>]N/2O4O
PH<8^>"!K99;7=+C')7:88D(<(-7E<W="X'L1JD=ZPG:YIJ]&B'UN:-:+@N"CN48R
P^LY_OUY?:PSL:E+-?>=?1_>4=#;@N.RXE)B+C%5)DU(E>6783'CJBR"]1^]O;(,Z
P:[!JR8J/[\S):;;3=WL5)5J?-%@6RE=S,V/GW;%^"&+?VO-UV3(TSFA!XQJ,T+<\
PF2&9EJPW\AF1%Y &QR7;,LO/ZT"PIC@F6U65EU.*AW?M&#>O#JF\+Z,L(K7-H',;
PN--'^P9HR:SV5@DS"SD6&#[@#>%ZPH6P8_NIB8_E23+_:$V@KK$/!YK:@48:>[DR
PWF*S+'5<B@(:?W#QKW4U('/C?K:Q=&T-T+HS)E#Q4:Q7\40"U-11JE55^_Y0 8W=
PM=O%1B>[ZUHWYT<Z41 ':6;SV"8J]?$N?K$Y/!F-O:EI<1"TD+J(:^K]'&0 8L*V
P:L29"?WG&5H&)/R&XN79/ ]U&_^(K+;7)3=9 H<*>GR(0#"*83'P[;I8>?WU?,B3
P:W4E])J'INVE>199Q3#\SY/ZR]LXV^@9;+SNQ.3M8HPNH2LB"*&OSTTMK "-/XQ<
PJ+P'M_88O<D7_R=K4D%V(WW4 PY)D'Q?6:E\11 +@&OIUEO-0*^J0WM1#(9H4\R^
P<!SY.45I;"X*^,$8<TL_'E%7HG12&I:^V\ V*NWG#:M+<V/(\C++%W0>:KHFA-6N
P  :<FA7>M$UR:HW9N%TR<\WHQ03K5C+)P.I232CYYR[>UR(V2OJWRH91,$0/'%;>
PXHCDJ;T4?.Z7?+W8@0U'*J.&]@;(<]EYD43@,]2$?39*-HF"Z*XNH2!O.Q@E54WX
PS]<? $&'RF@Z$-<!2C<]=\X+GO2D$8KI"8C%^[Q)!OUID1QMZO*^O5$OA-R&7AY9
P,[M44ZCV>**"44I"SMSE3FP:]<H6>TQ4QKDA&A-1(<CX2.LV@<0XX1& 7YR[IZ4W
P'_!]*LE:B38?WU$R:BV=)<HG9+]:U<$!<RK.Y)2M+?1H4UFCE!9M@I9H9HP2]"Z2
P9$3DYN':FS?QR,%Y%*#<HW#K!AYM\30\:R<\TE6D')A4E.O!UY57+A.+5E&+O++F
P0[N I/PE57=$P6%$ ;*QLIB<BFU+A(/3\%UKF/, !J7!C[P\V_EN]81ZIW,93,DS
P?A*O@5>W49#BB--872<C,L7H^DK@KA%(+]LDZG_<_>T1:WUP!\=D?SMB02/W\:ZM
P-(%OE<SGQAP)P7>3QL RE!#.O6V842JW)<2U0%%]>[N?(S/?H%D"#H0%Y2K5,R-^
P5KSD!+^VXCA-0I5]Y)  ],7(C8J@/^Z5E/0N5V,M-4U:]QG\).P$3IL('-R^'"-=
P_B<IKRP8/V?D]!1A2^ M2OXXZX$*5%VGKG<OE(HA^G QF;IG8QSZ20^<56=*A1\0
P\T#"[WIP3U<:BV-ZTR4;$"SE@K+9BSZR4QCF_*-UW8GRI8[-TG B#<!0HKXTC:T(
P'-2=DE]V5^TL1V!<- W]YQ,FU)'>R[#R <?]$!"+ME01*C%->Q\-;^MA LY.0P W
P9HRUN(_:]4E9_22E%V&WNYFHJPA6+7T7C&?=K>TVEII*8BI)Y^M>O0H@?)+3]Z#'
P,P6=74,=Z$M[X6H@++/WK3D_ $#N3>0[\NS;U<'"BO:H!:_<2=LM )#('WTY ]*C
P)I(,(K:N2G\HHK#6(O JR$N2*GI<Q+\V+N"[2BAVZT=)I89O:"NP3.X08N%N8YY%
P%[9!A_I3SNA#*DDTF_DNB7U:D91BT%^0D9.99A[%B ]1"N.3]Y/!&C,WDS)AZDPD
PB88_P7'16"LQ>^H*G:";3-!G9\U4,:Q^>&_C@(FVKNI(BTB$P($@L^*27O5;V!LH
P+[C,>M'%3_0OWM+WFF?>L4S)%3) 5'JI$XS5^HAKRM))5<TFWAM./KX2-,0$?DB)
P#S]X2K->YB52J)$G:8>OHREK( J^:.LBD?PMEL2_]0';^".0G%S'*4S5_[=V2CDN
PW(_M 7C?!PR7&3/;5Q\GP9#?HUX[?X4_2\(>\H4TY#C9N2;$-4ND?O/'(N4/<UFN
P[GCT,ZZ+?"[2L+5:_5>7M!5"([%)NR,.YQK-?@DSQL<AM^3>I$E:#Q22X0=09NG@
P2^O(@WC4@%\>0'IZZXA\2^.W0X+=J*?+YV7PS=@H^S$CH48"&QV25@1A[5653O0;
PTBY,LV;$\TI",M'92%F)+&UQ@Z=Z]#T=K-V)RS^*^/.9.(%AAU9L[U-J($O?"POU
P-JI4GOXKWQR.EL9YG]%N\#U8.8P$T>4M[<LGW4?<4OL).1]@&[LD/'!(J8YUM'HX
PZ%?2U%"2(*U6(.J'61,7R^B+5-"8^9E1:3/-HE$[GO1]")CU/74LOC6G6V_UXT-#
PTU16BF06"&[1%H0XO&7 PJ<MT@]ZOLK\O(^L MW^5$@$,#Q[&^.66^M6HOD_E1:!
PQD9):B^)U^:J"%K-P?T^-@C.!;G2=PEFFO/>Z>*ZI_SU(R\@&V) H #4 0G<.O3R
PF;B;)-TY'<^[1P7I]MPT5C-G+HXOTG& 9(:[6QH_MS_Y*U\9KRH8;'6NFQ<F_2@K
P2OVY74'N;^%@^F$FN5:FV2<2P-AQSXO^UY<5O(%<"$ >6/?/H_])>Y;S. >-&A!0
P#I9T][(@WT.7G3TG!EX_Q>93&-"$]6"J>%_3,(E$C^YS<N.9B]LVVT$^[K<^Q?='
PCU.\"'MF?WJ>*0[)\,]34:)BVN#%CU'J!N3]]+,-=%.3%J<00YS([""3("578 ',
P2!\_J<'F:/_$=_QP;O9J"SRU=.A"4*":UCQ5*XX*20< <EGY^QVW/L+0SH.5.WUW
PC:,#!J>\/;(.B\+5C<EV8.(I5LT*!!_EFB4R(1^'(MV(?4?&[^&11\?D: F&8CWS
P><?2I7VMUU[\^ 754]R5FK _S8(L4B(K+)([N0NE(<IK53NHST1U^6G+U'!BC!>.
PRCKF6_3=RH\V[ ?VEK3:Z&6=,V[ONL@;"EG.(7L-P- BV_N(17GX6L*%>7LKYC\Z
P,+FDW09'A;A6%*E$P_TC!-1UC5\'[.G-B=:PU61Q?TJ=V/3_7YO*WK)H';2J; '5
P-#DN+^(5_1UTFIU\IF*LDD7^%WA=MQ*-&DJ;_85Z@7-1^,J7'<Z$2<<N6^V,OA>A
P]\9_]>C#,5E?<-4#Q6GULN[,C7BGM[>XPGZZR"[&7*H4NV+WD=_M/M%SRMDNI.#W
PWC!G;?)<PJS.86X2H28W.6 N4$5H<K4W[7M-KO@R0R;"_F3=/J<?I,;07L7< IA<
P'*-P0D$I4B;>QN@N#$HP!2T7]R;U\\6)G^GU:!\GQ?2L\HU]=GYN(8?8VQ8U==[W
PR*"[\:F F?OMIQ4(3F-36 ZPA^F_P_*VQ_XXL^OQJ$%Y^+$WNCNTK,>&C$X^LN4(
P+#<:AV_P]K(ZG/@OK"T;FN6/30M$T79Z4;2;Q"M5,R;N[+09_[L*?72G7'.*A3MP
P"E.N:'!S[K]6J%\:R-4S]H2>BK]D:Z13 ']M!>=B7YPYG R1_\3N,N)R1"'590BA
PS_9")GQ=0F&@U"4-((3 VW3R"D,Z!9 [\-"@M?.ROS6 9C*^<O_>-G-%A5QIVFTC
PS1#UD.6/G+8M-I54P:*BN )<?/*3*GDT?<]_M *NGLF.>-LNENCWV?\<DGVR32:Q
PG71KN)*OWZ0!%3[=X@W LK5%=A!QT]?_L5M;JG=>Z%<D-\V."ARU]/@BR]-0[!]-
P(ZW"<E9W?=&:Z;04?IR'%T=S/>72^%84)^Q#UPA<OIM$UALO?=9K&5V$_2!W;P^)
P1UEKMC[)>9%SB$+++S23?16V]+1(\ZDYI&/*LR#8FQBE]BL"NS1Z:O;LV+VC,&PE
P2B?R]CQ5BQY1(D3'IM[U(6$R9=M'HUW:.5\Y!IH@YJ),&TWR'7'VN1PE_\B0'C&L
P\DC-AFR1RE?DV0N6N0)NQHO$ED '-CTC(P<EN_ZO$R_@1,YYPS!55$.FC2]>O2D5
PP6YSA^&"_BJ_":9%N'Z!&'43WYLM:"&U0-8I-T^?/X=81DKF8BK;XYZ\OA7VH&%3
PS9061JFG$+3G_BNR%=AH2ZN"8!5GQ:I?2/PM0 .R I@@+3J0K.5DZ+@V_8F,$DIJ
P[ZI4?:.K.?>Y1QKNQ?&R\;R=E 0/O@9E#>OHU;:I]+6 <NH^4*&WF1^H!@E K.?W
P'\\6R(@/0ZFX%>;4UDLTF-R1?,-HVHX9OX='L$AG?'I.<41L?_/1R(FQ3@^TOE3 
P:D@+&@/.<UV8WZ(;N; NG>*Q<YQ_':(M'C297XZ3*))=GE=< 3I[+.N$F61>;^:\
PASZ[% GY);[@U7>J12+^IF-_O+1]MLA[8^MD^-]KW3+JPBZ<IW'QX\*K2:>+)Y=(
PA9R*75V(W.*H&!+J2C/'8"NM*S[6W%2[@8/.5O5[;D?[S2LE77*Q';#*.T[@UJP;
P+E[6B&;<Y+#B^/*P05DZ/O5ES6S3J"'V!D-P+Q8ML\+#]JV[1BLX:]BK>'+7,X8-
P:9(7Z!@%_]V@(:] 11)_X6D "M#]:QZ'I5MZDPW8],^E!$\S;IO'SU2V1,SA5]S(
PN:*KX:4H92YQQ#H\'N+)^!@ 0,-J3R#8YZ<N_)K<+_UPM;A #ASW+1@W@6Z^PF:P
PKS5OBT\C'/>[(P]Y@X2]]90-V1=6)1U))P?#VD/]/*:0@FQ%);$**-)M1KA#-MH[
PT1TGE2"Q^A_(0A7WH,$157#1<*]8;,+1(VY-)*>E%EAC9@HV_'^.U@S\5?#H068B
PL*UT*0$CCS08))/,3Z^+1IE\&J=.-'ZAHR='H6##ZLLFK[^>#EFMOTN4H.KUC[X2
P_PA@4-ED24_3W ]=O>A&F;[$2/@^,=-84[SRLTU.,U/RMJ*Z/CAD<X:MH*/7<?2M
PNBP*O):-;B?]U[D ;O-BL4E)!C5>S6_AL,F'C\$L(_?&4X0\0%@#4+TDSX,+H5;"
P[G&WUI8NF6 44;1K8/#FS674^4<O\M4YI*D]35Q-9;[IP&HQ@P?T_?QKCI*5@U05
POZUAJ08WQ2*BH2:\42R967D369:1QC8)"68$=[B2ML+X\XPQ03<]++,&,15#OK6(
PUSI%3?@-1HMX*D<:WSR)%:FT$X7MX@\KJ/-9)%H]J*B;&"K(Q0W6!J5<"64&&/+%
P]4__AD)VO<;:)-@O:0V!;_2BY;-+G'VPY(]ESAFE5*X^ UZIGP^N8;V_U-'GMK,B
PW^SY81WY OD8U5LTZ0=1C['!])2I-F[X]Q$S1(A1ZF4W@^->4@BVR YO%,,%8;DC
PD1#NY_.(GEC&Z0"A^P2Y)T5V/H^<ZXC:##NJZ9^)%"Q]3%K52K/9K9_#&\= 3JA:
P+[74J&FUOZ1U8JY_*1+^]![TQ>JR;Z2 R')K%6F3T<P9?4Q5#PD$XP3S)>;T$]\&
PT%;83&JUXQGA%XF-[U^$!,;L+3P TUM:'@W9AR4W'J]\?6A!1H*+KFW@7IAZ(E>%
P:!_GWMRV?&H&-'^X:V5"&&[0^<^MM('LM5S).W>N%$ .7)%!HP:*R9S\Q?R7YC6,
PCB?*9%80A[$(T+$SZIH?*\6-7MQY:B79FC]A;6?5NQ1P%WY!.Z.^-(4I*%I-)CDA
P<S9AX)[P.P@SKR8I8A5?.Y=>\C!FUXA+NS8!ZB?%I>W >WYMYRVC7M=XJJS<ICIU
PLFP0S&&-M$^J$&8JO)CC\V&DIM5W:&[52&(=Q& R53LRTT+@B^:N3G^)NPJNAXT'
PHI1@O=:1G$1B$DYN5NK;^$1S\<-3#O[Q$Z[=*XV^)V@,#9"Q);)Q&CA!Z_TMVEN,
PYG&F>;/'X1)D![(LX;6DJ2K4,^ >>*/\T/4NAQS=TUZ3''EZO>KO> U3Q HKI+%E
PC"EVL.1'*&B:;\VP6'&8 O"ZPZ-Y&%&68W8<KJN65#\M\JG<$D#_%&$.;:=# .>I
P4@0$_]:+52@-[N#_,)>3<#@:?;E@KMRICS2AC#J@_DFA!"^"[>:'MSDV"'WJ/"]=
P"I-#F!7Z9Y+?J&MLXNB)'B-,:=MPQ5J1BU 10ACYP0:VED.6EW"9.17V^?H%D0LO
PG[8:A&DXT<"K(L59ZY6X5I)5EYLC."[B,*7YJ:(DK[=/H6V"<Z'8\47;=9_<VMCL
POX\1@T_PT\S 6>Q3E6U)JZKL/Z< 0J!H-[8TKX8O&TX(J:2*DCW;FK1"J:!<:/&O
P?SGJ,]H5-7/W&/@^K)F*- JAYG2&J/=\Y[?>TZBT:GY(."K7:_B&K[XK+)A,@@V7
P>[6H.H (\.ZTT.XA3'OI->K/1DB4"\-.I7!G0Y-DNM.F$W8&7D7 M6.L,X2_Y>-.
P.4\E@"P@9CP_,\94,4SI RJT+:H?IO-^::=MPQ,^@G.LL1Z)M>M93;_J3W=!89SI
PX^3(9M(;*>HW?_F),FT4F.F?M9AV\;?Q@&B^LW=]G U;:?'M%MG4TE<G#-:+8?B<
PPX@S50\5ZT1L=#1) %_MNVPCGYV2Q.G.9?,FYI^9D,5+T-)ZB"A?&7AC"O#"X#5M
P#\<H5([.Z<XL/!LBT0RM1%8E;2!'+BV74]LJ=9')N"+HN.+)XB-HGKT"%H:E*N>E
P2W @@K-M*^-1)W$5X 1TEA7ZP32$Z';,7!6%T1H8";@H.7D)88#P]X7(Q\VC\?)2
P1*KZN7W>SSKV-PQPA8#%<;5,?^)?Z25#,42 7P/6.<Y4-@V][*'JY2=,>7R0<JU)
P':"B\W^M%L7GBD6;4D5^3'R'R)#UTK:3WCQW]#;[>+8D6!RH3HA?YDU_W&^020[@
PO!#YP86R(O<P]K!"$P$4?YK9')=].JX4DSEAM'M "Q$[NG.@]!*7#@!G77/S>I5;
PM2V-9];JO5"7& U 9%:S?+F I/\2R71$W/Q OU)=C%DPZ?'[:'5#PA#!"ID^GV=$
PG=^:\(N+?%,MU&4'U/_,?)<%JJM.JAZRZ1\K\EM:I2%5UF<P<J1^:R9F>\VXYJBB
P:?[9,'LDK3"=9E:3!9;%6WH6KWROS?T[2'38"0L&;O871I(8X$HEQ*_97<?&X>ZM
P7W$F*'"F]7[<BC@,7 8/ G;K[UV<)*^LS)L;*]4M@_,GH9 K?D=*HP6?J0M, 0JH
PU:$4XF_ LQ[U-39Y_8[*L<7DCX"8K6A5IG^I&5'/K.O?*PH//]$?'-G;2&6]+R7@
P%H5$?,9Q:_1L=8FO=H<J&C' XI?'\3,'SDV'B)H$C3SNKY<N$UMUJJ7_S$]%'LJL
PZHYHI>+__+H;%T$7Y0FQP2J"54*!IAZF?S^P$:<=VE'1"]6H'%7*(3]@&8.@223=
P!-ZR"P+>URL[(N.>F[K?\MAESJ]BLX)]EV:2QJ1,7B&LFZO6T?0;X&LC/E72?=%V
P0(4_8++A2]YA(@[[$0T"X5)0G1P[H"1\,("L&P,Y(8\B6.)E.-ZB_3N]3!PGAVOM
P>+[&_I$C_*O?@EVMB\YU=C)RKB0,<7P;R=P-D*C('"Z5@[N$79:"H0\ZCON@B5L\
P>W<@]5LO$%4!#6]=T+$'])':S>YX;&"^KZ,]P8@J:SR*[D/>Y '5=#;W-]&:EJD4
PUAM;ZL?8/=#+:NP#Y+(5"-4#]>1._A'--B0[&F^#U/>W/1_C:],E$E*PKOO8.X?&
P[@]N('7@_= /1;1=DF.1K8_"[K;! OV!C%UO&IUJ,UJW40"Z- M]&)V0 >D^BA$5
P$;4G!)5\*I<0@,OSYC_R*Y!CSC4W0LO1T8DS,KWIEH%D9B)SJ9J5 /M94OB_$BL=
PY);+VIF_.["VSHRS%\G#N<$ZBL-SAVA;/6IP!HB(U/\ &+BJV;E 89C8*CA-*"K+
PX4HR+A./RNG#R[+[Q\;?VD]8S4+[;3PD22HNNF3(YG F6(SLT[D?XOYI0(J<=>$+
PC-F<,1NYZGIN, .DZG0,0/2,]N6?S.%W'4V#8HOG0_4?FA<DCV,&A:!4>=&>[;G-
PM<?[">!_=YB^\>6!F+%H>[,UE%R%432"8;D#7!T2D NT6%<*_($0O-%B=0"0J<WK
PSU9)'Q.!I@-6H!%29^#S/ZIV?IGB_%!$3Q.9P#H?)=1D. '0?H0J!X/4(36D4N+>
P%S<](.['R7T;NSKZ\-U_%4JAMNC1*(^/Z_Z( ) BV*=BRKSC$T?6BS1BKD/%T]C;
P+EXSIQ_7"_K7.BX=O&F8J?+'^TTYA%S\/@@/4%)>7QWE9E"9WQ#K2G:!.Z%Y\QB.
P4 8QN#:XPA#$XY%BJ@,8+KC"-)/)*4 JAJZR$LG#&04R_* Z6J[KEOGLDQ<\B"F/
PWWQ9@>CU 24EN'&6&UR)=VXG)\&7L3HO\E9J[J4T8 MYL75%[A!>K@C[05.#6^#@
P/5LJ=)X\851NX;OHQ4S$4BA_  G+BN)JV4/(<G6R.]$[? /'6$J@19H@3^/U:.;#
P<1JXY0:'=CB+!X&^MH<@7G/-7Y$#H\#U*:X4DAZ#3NRC'P_-B,NG5ZBPP*D@#2@Z
PA0,3ATH+!0=._[S6RM$\,G?3Z;?[6/K8G+N=#K)[>+T]-AWNOG>_"K<C>XM"YOA>
P:\>:I'+)ME..QI-VN*$.E,RHCTS'H\J&RD"-GS9JZK7(_8& A*K _;B8*H/-7T-7
P2=@Y^J>U/C;XY<3:OUL8KY<^Y#M.VB&(@BZ"P>CG@(\(9JLQ+48S'TJP ! ?U;+8
PB@@\\D9WZK-YF1.8BP57HB"2^9=A)M5B]2&W2W8N[=N62QY<)P$-$;'^3QY%>GS=
P8-!MGC[TG,X%I#ZXW=CM%F3Q]D00>;%P?ZG.95O&Z?*>"P!Z%1W@%Y^@-GYSH4X=
PN7ZG TFMW4')(Q '))OT^$&OSV8$K4JKZO+:ZY0CZP+7G+U$Y<]":B&? 0D.B-Y.
P"5QF'=A<RDTS_P*XJ.6@'C<GA*VH5: F7K#C&DKFB50I&5SA35HI6],,=1WR?<2R
P0I8P*1<773,:;CIZQ^E%(M529(I$ZLP4KQ63$DY5 _8&RQ&CH7:]F[H*$,H*"FM$
P $+WUR39<#E$B@/_<6B"^4IJ%3B:-7[;^O5'?1U.-;T B$8%FF!1+ZK!0PD$Z;@=
P=$PR- _8Y0-]E<IE_NN*)<)4O9**\]C30Y*3KO>FUW.)%+A%W)G  3UXK?DT'41=
P;J!\UU\&JH!QO4/B[1(@50<0/F.1) E\T,H,.9_/\7OZ6+P8X=JH\/!%/E>SV*^:
PTI35+L0S>#%;[)5WH-8*-/%I6ON%OUKJ_ ]#PRE[7;V#^)[TE?3F31024GDJ#$HY
P\SY][G7)3>N#X=^2,>Q01@9V30G-*9/E2IZ5+5H\=LHG:XIC]F3^8:JC, L%K>[F
P,4A1&X&YU5BY-3LO-5_ZF5G*^0;\,+BJOZ+'9LGH;=O:Q/V@2>QJ\,1QT'?TYNN(
P"V6BW,?=_)<GPO0D/K]R+4UYWC1X<NHJZ<S7S#B!^F*GO-^Y&H)QTA2Z;=0F?]^W
PX/[4!#M@_''OJR6P1E.FYP9 <EK:=\5L#U(]I1N88J<U'ZN(O5>L[E2,X9)HCL.*
PWT6]RMCCMV6NO88A%U+>?)X7ZA OSP%"/W:0K>W<!W09]7\0S_1\,:&!'[$/JMIL
PS';"J=)#(5+OB^=7^MKP=P[&9AG]RYL61Q*&"Q87I0)$O(+KN?\O_M+&QO:Y[11<
PX^.XL <6FX/C8+3!%@P7PZ.U SE&N?J5Z=05L5RXGS(KTCYE0(+YDT5Q+MG/+<#-
POZ)@<%DX'J4<3W0?!TKTJPB<B(YN$+-Z(R8<U=3C%4$'3J(7ABPUY M$05U3K:!5
P<7G%%QQ1PGXV!9Y9 @!H8OXC<J7#FJREG<G<?1R;;O/FL6YXD^!; ,E$4#8\::-O
P&+ :UNR2TN87$T2K0O>0G!#6=W68;Z5UD>:*Z]#9Z_X-*-JQ#BFX%&0N,Y0.-." 
P*9$GLED!5WPE')K11>$1^$28MWY8Y!?*D[?5:V)15:[S,:*'<OY+;V>>C<K*UQ#T
P('G##27&T7\.'4V_BP'RE>1/??!Y XTL^\QQ=_Y=,T;H-Y]Q-C&!06H?JKI^P:\A
P&<I+62,_'4L_&3GZ3>R71\.XC--7QI,:$!S+>^.Z!NF,6+5Q%H+[,,TNH&/3AC$M
P'-XS,-J[&%R5*MB=A^:_!LKW[R/07VJ:Z\N1?4 #F':2Z;:.;Q7>'9S6?/!,(]5Z
P"R;<DJN\(.R1,N9W3$D0U+*0IB7\_M<^]@37KJD<3-B7#@*4WU7"]?V@O\T:7G&6
P;A* JWT#B%<61Z*UO CKF;A@'7-<C.NK.SG+&OBCJ)9;R9A'0U*NK/._L_!59-;9
P-38;?$H=O9MV%I!/#+FIOVED99DV@*W&R*@W4O4'5\ZM*RI6%-2Q8;#<T=KDIE7G
PB+Y>*-#/5JK\,L!D [1P87%K>-^UPHB<VI?:+M?I9P\!6R9'35!QV)HE3:5*%TBO
PDW\RC7\X8_]0P1S"?)5FUF18N9!S"-[PXSIB FD?/TUC@R IT\:-!@[HJSIN6)F[
PC8<V6:JH_:<CGK+&^NLS9O[E@YU/BR50(5E['=.\VC**;$5QGN8#%\0ENZ)^H+VK
P:"<OG:D]%I[4)C'@, F#OW&N"\-Q8M+NB(M3+RLR#$#L:+>-B_&0U"F.%"$A@K25
P@NS%@9(?%SL-<.-TH4MGG\Y-F$(_GUY/V"#I":'+=OZY'F,+Q(WI@M-WI4R  1\O
PQQ/SRSAIY.86^;^UZV;-\*][\H&1IC'6=H9R2\#QSR]>(7<>P($C#KTZ-XE>6*ER
PA89\-T0C ,-64V0R&6I6BR6!8FL7"1[ZZZDND^.O(1 K B(DR((+KMR(8"0>%?IZ
P]W<2A#?E+%<G]@,[&WF*"EH>Q)A6[ECZ0" XP(:95Q'9?"P.R&[O,8+YQU(!-^+N
P]9F?E<OO*^^-M9K>L--I=PX0!"W%_3.#).KU4OXB$ Q%;21[)"Y/WZ!5ZY#$I++7
PBZKA^CY>&Z[W-UJ2U7SR'U&QR .+MS)FUFDZ.]8T1<>PY[B?'E[DLW&]L@/+VD([
P[IPA"+;V)1-I #[3+:)NR$)5FX.N@W[V6_KQVZC_B>@&:/*LV\8BWGD@$Z4ATZTR
PQ2K$8+C1IR5VY4);P)C?K 5] ]1O8VK<'M\RN9/CUU8[X=7H7861S9"FS2I)(0)@
P'8DI2)?C+2QOGY53]9+20]K 5C1D)P!E9*#C7O28$ @J\#MB[\>$75OHATCL*P#!
PD50\%YHSAA %-OUOAX&2/\ZEBUO7@ ;4*#TOD^S2 $C0_;D FG^P!3:$V"NK7DUO
P.^Q4(.$:$86W?!"U69Z3%W;7)*[44XX4R\6D QZWC:5[)Q'=SWP=G./V.OX)RG0]
PM\ &*Y@M@Q@'2F&G.T<L/#"Q0#]TB*8+WW+ISO2$_V57/?XZ0]BY-Z)L;I0'$U94
PB6.G\H,>;.&[Q\J*&QJ?Y(QC/ -360WG_Q.?XV]-XGWEO%_6Q(11?+CMR?;6O[@W
P,!P>T"4L99R.VL+Y2I&:#9CU6@ZW3ZQA <& 4V+1A<U&;H9?,"#NV(/SQG<^_4A'
P!E#U!V4;I[6G/-<^U _2,.L!?#]R?2H4(\3#NR4N4-(?J90]&;.FW;I.T1?95<,I
P5OS_@-_=<'##9ZA/-:M/,1(@O06B391J/O'_F)3([V)!8=/D0MK'+D"^9AYS[L-L
P;=>LMLW*39'F.EI,*M)5:?JR1T?;B>4<*4VMM-#TF6Q>1M&\Z5SOV,Y_\:/R\5UK
PA^1$^($H3"W>>X+)-;HCEM\K?+LB$/3-= (0Y'-G9=C&!I*^... >7$I)LK4'VV=
PJ#Z6P^\:<X0R$<4SRRY:_=28S,:E\<IKVAGJV&%&4087D*YF( 9R\^(E\&@)*Q6T
PZE%#!Y!YX0[V8Q*"7V#T1^9^'-.@Z^V4?N1@T*=!HF!YKN '9-PQQ_QXYHH[X&XK
PF:),@@5-G?L:*[[Y)E?_PK0+X51YCWJM7#52BJ25[$]<J6?6J-&8NLD&*I'8&7 3
P#CR[N#C(7!XS-FY,%I-U%L:<'J%]2#)6'59$)B3,QIG*\:2:>+LL7,#D.1M*5D6/
PJJ,'E!TL_@^5$!S5A<JL*\U.FE@.XOM<1%[*[XR]F++CA^]'31X;^F&H?W6QDGEX
P47Q>]B";S67CB!Q;2=Q?8#ZG,5^?N@6U!0#ZY-5GBM6*##BT*))J;;?^".UBM"C/
PK'>8/^GX)I I-#)E<NVUT.1?U!@7HX>HU?9[/M5VY82RXCY;I29/H6H(/_[\ .^9
P](8;<%(NW!-UAHIR8U1X/<J-=W>U(WY(B"-<RX,>ZCZMS6X)^@#X@?GNFCX"B0'#
P,?Y=0>2.18#(W1 =;>T4!?8!G$ 6-]9D-Q_*EWKZCK#4^4I+<WJ2';ID]<I>*D3U
PKN:SY64?3H([W7'J.Q\"%)HW6-/COX+AS/7&++RVB:'XB??MY?A^:"G/"9 ^&21O
P'NH[V0"MUDU\GO>@CC/I-_08H+L@/V&/ZHK7U=EA6@L2]H[U#P%3/CF+H'@@BU*2
PFG,+TI8-K0G"?:Z@#AXA2"D8_$L9&<8D@]$B?6A,UXT&_LLD^,_(/.[(5Y^N\]F 
PKY2+'AD^DD\::5B<H,E\#Q$ZW\7/($^Y>.[G'4G# S('*VOC?-][IDJ.AZ+XP!) 
PH1L<XC<=:7; *S[>ERRG!_A.G'2O<"\4/8#&^-8)_CS05+50\^K ]NP:#3T$"#_I
P6!(#WM#6BWM_\9P,.M_ZF J7GQE@>1;<]I5MIX^:F^W?W.92B*5]2C)<>B'Y= :"
P5EN8A&I_FEA?,@M.#] W@%'N$C3#EC::1FCK*VGGKO#KQ,&SIL!0+Z2#_!YU_Y6[
P COCYD_OYH57L893+.Y9WJ:\*)VWY#4LUX'Y,*O*"-458:&R Y97;L>MVS756E#7
P&?QD?TLZJ0U=43%#C1JXJV$/O +O(5TB.0=\(*VAW*I@3#-*#ZT;2X"%0GEU<6P%
PR1 D/^Y]L-SP4L=1#1M<$_VCY2-?J:[]WW]C?JO%N'D-&W/,<^92W.HA<>6"E//P
P-Z6*N)0!G-^I<X7YB_[;9>576;W/OJZ6<&\N):J-72-45?!04V\N97JQSC'[(+*A
P<2IL8LQ79Q"YDZJ%%V%"ZEB^A,3MC\2H8BI8NKTL[R=KBBNW9[MW5*WUG77DRC/9
P/)P6@1P_JG_-,#*#@_/7/EZ.'F-G:X0;/3M-U;O$;\<(Z/BC1PYH]Z72TAJ;UD5C
P-BY[[DP%L5FR1+VA[[1##G$Y*^X>,(Y(9&E7AYH1W&TC='/A^FV6JB;ZON0Z5,O)
P(Y4:,1"X_V'R9_VP!9+DGPAW>Z4-%LT_^JYP36"XU2#4W,C:@X!,%#MDDWG?_$CX
P22UM'$CQ"_P>54S'OC.[QC^.%H&LIB-35R:B?7?HCS4?;'DMNHS$=A;%4@6-Q_@[
PM%"]^Q\28NH$+W+]F*Z1H-0%# UAM_!Z2;?1WQ[DG14;(,(OC"'AGIO68TFT]Q%2
P9F,;0)97-$;1Q4M^^@[5F\M<2<S4$(1\'M#3W -DI2>E";?:7T<H]#,@Y\NT1C'@
P"LGUPL<;!M=%0I*4'?3%@O,2S3%U0"$-NV_:Z::BR##I[3'N&P,">6&;_L.\$P- 
P%1?%6$;9QX)S?T*>^(&;[;SO=2I:_1HZ3PS04&K/[PU*3K$+QRFFHU>A+EU&;CXY
PF9Y$,MMLB$@,Y7B39-V)U0U9%;YR_)N"-%\BK^0]7-J_M^[2QCN\<Z._:N@W3Y\B
PK1^3N5D%7!O];_;U2![I&6X/UE@?&54?LY@X&6VCPBT\.E]Z_M0KY5^IK2R^CXE:
P]06X3:/N)5P6P57.(43-,@5C7VFE'7&8!W"CU:NETFCM2^9C0?X2DP]_K3>'QF?K
P6]N>[DF A#[L50./YL&NFBB9;.S8K=)XZ@K2E _]V6X*4%@W?(?$#%_B0FFOB?A.
P$<V,T70&:B6Q5.=?&A]T4F0 *!AU!NEDI+Z'+P[91T?@AM?5_&;=SO##B\B:J<4B
PX=MA:I&>5,Q^G?^UA1(WD5D?K-/4V<8I'O#P*MJZ*;<+ FRAZILC@(VL1[)7>NU,
P$?E0L_^F3GI)$V,+\;H)!7(G:XCQOQ.I,-7"(_=M&(A.+OIY<74YA)6N.G!#W4:8
PQ52D%D^GL3< ]\EK?5H\[UC*^,L%$QUFNV(?T&9(TF=!'1%KI+Q%&9Z"15()XG>'
PFMTFQO2O;Q%!;'?[+7U++4ENZB8@'</**Q48S**X6V*4L7D(G7WGADK>-*O"38J+
P(R,FC<OZ!^ACUSJ/[H&W9JVF'Z/UWK4 !5^$X@R;OHP?0GR+D@RBKI &,(=H%#!A
P8:9S;!]M9_7SL1CXM@K#8YB0B<$[N!:!1+EHTWV,VB4W&YXNL):1#ANPV!!0ZN\]
P/8BUTC(;9HJ*G2E_:?W;J1C<'[??\\39 <6ZN1RD4 VB7G@ZH/C"J^O7?O(2/S;N
P3 &]!=.92WN>2&"/[?\YY?X_]H4G9W 3ST9,!;ORBJE S+DK<IA3B2'M:Y[4RW0S
PQQ'X5&R#W;YD[V&BW;BM+5Z/M]\=.XRG.1554R_OF#:-[U9P@(#'=+QC<\?T!<)O
PH8T\8-\(-,0]W1(5MI[8(B^9:G/??@BCK<_WHUCM<6?+G%7KL.=7;92>]_8L4.3=
PC@+Z>0.D?N/G8XO]_+BP-Y)J,+8L-(X:!_=S4F'M:4NY]B._X-+J0T8-RTH9ZL9_
PG3W6<S*NTH0-RJ^\=ME$'5K>'(Z.2;T,&,/B6$&5TC(Y:6L.6JVE8#R2Z%/%2L*.
P1*8C\VQ!D[B\P1PG4ZCF@H=6LSE[IML@#I=RV9G9;@(RNY%>6LA*^8R[>LL\2^$4
POJIX4'71KP8N_+A+(G[0#/;FV8.1JH<(WWJ( >0:>;'%8P=TYIM^*/P^Y2;-.R9F
PP*;-",R4KRW]0!1:=?VS.Q2CMVR!B2W%W."%(L;K7(!OZ7 Y.&!HN 98K=7-ZG\<
PA\C8*9U!D B<D4=8)0ZNZ0Y/CRF)/@<RNGI_5[X A+$DER&*WA1[Z/?L7EC! -&Q
P7+U_"/JA\:K/V+;.CC1MW#!?^*D0DA4'>*?HS:)ZPA1IH?BIWUTL,#3(U2Y(PQLQ
P#'\+0PN1GK-!:ZT%?C,:/ZUJ8RY7FZ72+2F2EC_6,+<;E_25M-G>.U1.335)A803
P6-N+E-^D([*V9S59(Y56[I4<O'<W>Y,<U[6C T=^2@8 RA'M[*&&6IA/B0-]V/X7
P^ \'TZ%&PN&#CLB/2OV&5YJ<3T4L5JU5ANT\4$(EPX@&C7/1*F>;?@M#UR\&$*$<
P:I4O!:;/W>X :!H,*+SE-CO%A!K80O)C&]3AD7>UTH G@PR8!#*81I?-]=R>\LM@
PG=S1>/DNR90,MT->E,FY9@DR9,QK4NP$*IWE0_^G;PE.*</ ]6?/< ZSBM?S915&
P2IPXIYK+"U5G2\5H.L*:5V VV]]XG@Y'O^Z?/(U%N5?D%)T\;-NKD";:+BC/NT  
P->L$_[JZ%'>[6VM%2P:F.IWW,8GON $^&@2',-9G6/L=Z0 FS):P[&JG '6.5'I;
P%1@+C[FXVGW+:8,G:FO\$@OW;0N=#6[&]B<8FN4/;C]34*L]37^0&O?)^A@BF[>+
P+ZJHDZ0/'^VM=HYG@PS=2I0MM728O@>6EC%J\7^M2U1AQB#+)O2'?G$3+S%-@.P_
P$!:%:]%<HU6*KL.8D2V[96(G9]L<Y3B]7"R/3)'.-5Q!6F.J@\'VJ77*V_FDBSNS
PSBA C@FM9[-KXA_#^R5U^&.1 P7A@;O#V_+(31G[00KW7VP#T:S4-&"$RX:K/8C5
PI5BUD3%[ZTN/3$12]N?_/=0_3A<H3D=;-OUGVKN'%FG_?#*OP $3H<TKF21]"-$8
PV+R\NE_]:'=<=/A41.DNC>^40D8$9]G)M7QC5VHW[?M"8JD)^U  ]>BDH>=F!Q*+
P#DQC;]R=,%63\<L(LUOO[^8D_HN^T1EN%/%2"T=\322#ZWY!-F7'Q0$HG \K3.Q1
P#6!E'I63+W@SR8QAA,(K5&/GSX+!R FEH4N&Q"(MB,\/Y4E?7!(@Q@$O9*RB#Z]\
P[6BG)=!(M\$B'>!3@:P#1'1T!SO-7]3FMYF.;-OXS:OV,R@ZF[4M*.UY; .#\SI#
P"7L"YCW(I=!@([-@C2E?VQ%O"%E!B_0J.;Y0WP<PYM'T8^/"&P^5K"5W*!.O>K:C
P0.(.!LI_2Z?S@MT&*2&/%\=B:]",[\K1JY"^_"XFHYD&YK>(@K?8"&8E< ^K/;@9
PL!I#6JF3]3&M#T[&)\,<?=H=!T[#.U):I%EUB>$PU3D\?JQW4,V5)SB,DD])&,B+
P?MW1&(J-3 U?BFI%G>._P@(YH+G.'=2ZW[-A4HY<2C?XB93*7A2*KK>?F&N:60IM
P%;!F4_(ZBN!E\KB#RD$(H)]H\E^17]:ZV1[XEX!(S/LX0#.3\^3P=3.<Q"$_7+$S
P]6J()A\A7V.;*JG6" 4PI+5-M=X36[D T.VZ;7ZS?"C'SS,'O>XN==8@U+LN!.3A
PSKP"TG_0G3[?'+/#)8N.H\US-NE"VQJR$!56GD-I/AX=<"VK4-/^$]7>-4M5W(TX
P"SZD_2(&.,79,M5G2=G*8^=%OT*T+ATJ-LT7&>XRZUN?J5*P%IL=BHNC(-&SG\\N
PZIVOL!, 7TC9(QB_4P\+><9GB$O_@M<9C5;DD<$F:]Y7:R,^ />3 ;)?]WF$UBNE
PB5H\G9Z6D:8,P2:0(CWG:3@H!=67RC2?7.XCM^Y<4+Y_+8H<9,3 % PTN^7"^M$K
P@SDN/PM&-0\/;(6+J2C;'/VS$>G )?RO]L%H#4)Y0C\$D +1$D23[?U=<;C%THQ 
PQ,9WR= @%5950>::[&;M/4^I65/4<WRZS(_?_UJL%ZK"I5G43L^)[LIM&=[%'ADT
PM4-)4N;/6Y^N=K)9+Q"DL(\ S(P5_&QL'1QE-HLOZO5!_T0##.!3B!=BDM4'AQ.U
P6___/UB<:,F;=9'CJ9 CM1+E$\9J35)7!X8UK)>Z#?S'=^3GAW5A$R &>0>Y96Y,
PX"\6N_ZF4@!6&_H9C<,<>L1XNJG+>X8@<8D*#^?*0$M'*(XFC65EO7_T5WA:7FO)
P@N>FL_X6^4SU)"0O/*-\S[G+GQ53]#,C=*@)GRJ#13_]L)38BW2&]_9J+KT=8<S\
P_BW](=$JGLW[Z:6.[8CL>'CAX^@UT:!6;;P6I>5& _(F'8#LC:WY2T,+ #TD+V!*
PQK8B*$>$@"$,LP_T:W"]0 %<XKQPHW!?:*7[71X*1WJ3E^<K"#%\XLEYWM!@->3 
P(Z%TQ *R9*X+#NB["9,()(SQC/#,V>73@/$+!HG=Z"Q'.!D^NASZ4FP\_+U)#<BR
PX[^)$MY)D6KO$L0V<9C*Y%.H,XZ?$WO$*EK\_O@$#<A@K3\RH7CB)TCEAJ&4AL2A
P"0"712ADYA>4Y@+\' MWGE2+!\-V^H][?48/\MC ;WA1M72\V=& Q3(/7WM!7BN7
PSR(9#;)["%B3ZZV^:-_RFL5(CH6.[HM6ZU/'&![N=K!A<A  "A6CB#T71#[-#O=[
PG#D7?>TZ+S,?F3FW6^0C_NB2^!.@>&07)ZJ!XF9KI F06?CW'3(%&%7>S1H\6E-]
P](62[K!/=]86",U*'VC<LPQRV)!\FL^C90-F4L)FM6I5O%RZ1#GQ]=ONE&>62Z4+
PRK,, 7"4U)X,0K*5UKWZWA%/TR2,@"HG@\C8!M5H[P68,Q10,6,[D:.JIN<.^0KZ
P%2D1R/V;@L6D]'OJ-P'3U[O1CI8LG&CM? P5!_ X4.?QY@=_(T@/S(::_R:[.47C
P?)HRZ34&N*^(E.=&74@12HQP5@T1B2/;OP-"*4'C2AX"7/#A;I\N,&"I1*TL\#>F
PHR?"J]0HM?QJJ:@U1XP$YSJC#);P$:S>W U$/G5#9*&<G?*A3^U6-T@"I5\7O?NA
P]A<*@Y =R\/">"'@3U=TGWNZA]O >)3F48IR#HK,J"J-]BPUL>#C@V:(:-:VW(-3
PWX0 CS%U<TYG6-O)R]#"'<3WT6!X2;O4=[<:Q4:Q*7-GA6& +^,>\;)TZIL1#0YI
P<NEF_[_ZAPE+XG[MTW;X'J'[#5 :/4.HV;Y]9LS0:+N%6&H0\=UY0>)Z(F!+!$UM
PN74P$ ORY"W4T600\+R.GQ>NZ5LR"N0((-N.EEE>M!?@6R&K'=JY[('E?HPLFFR\
PES K6\L,<B8/@@F&]E++_*=./D#L)%7M .5$3<-[]5*K%;R-[(<Q#;=/KF&3Z'?J
P9=BD99LP+?>3!,7TN3A-"<^^.<!=/#5]EMO:$S?0=@9CS/NW\:R6+'Y6)\N:5P_'
P4TWU\2T_[>^GM$6\=;+]^^SYJ"P*#-=IX\4HWHUVU:+EHP43N=6)\F>/KN#I+'F4
P#N!@'0D/LX1IW<OQ7KP,T,!J;:]27JH<_<!T'U@K$<9UE.G?^JPDI>DM!]"FYQ8)
P/F)T?2G@@L.2,G9^I>5]F[C5RFE69AR<AJ<8[1 DG_1"L<N[<&$1Y&Q1>1-[VT_M
PE(]:N@GN=YYP].A^(F09E'H5X$?>3TCH;02@$*#V)B+#V9\6SXH>*7SJ+$:5T %?
P^#[!CXA%ZI]R/:?WSCS,?P9YFF!*/TDW5V:/U%4,'6D,$#@UKXQ3XRB4]>%]&<U'
PUY'(P]<E=-D9Y@.2DI6I1-GY*Z :%D9)K,)D04& J8]*')JC)LL 5>K <NIU1 8-
P2=U[> 'RM.X."S48?H*&PV:]$G(5'0I>'D5B\'8.Z?=PL\05NIO=4C1@%"I$)!+#
P2?I[BS9%SR G@3?VL<FA?+22#J$-NS@M^6$S>'L;!#TI_Q5+X2NIAF8M3+#9B_<(
PZD+63+M</ %RV=)37;T?2('Q3?(.M/0P3NYT:Q7ET<OMR$Z/VO&VI!O'\'R7Z_*9
P0L,&,5-4:U-9D^KY;Q:W'V#5"],]Y ,84>7IK(O-.%JF R*+$I6M%><;L_@%.1+S
PUVSY7U'$^.&KW;:V^.;CBL6[,F-W-QLVA*LN_8#C%076);]K897!;125R84*4T^C
P5X!"_[ '[D6JW>$UKQR[]IY#&GL&NS?+)EW/E;/#05I36?KFW*PJ)U7PQ93> 53F
PX&CR@!EH;KRKR&9[ _4-MI6Z7RA2@>Y86%N;M*)'1]TBS22(>A<((E?6LVUJSY!(
P8]?D-Q.+OI>D7/$SYNWGT?SF]/$6E'P(O9GY-8DM;3"I[9U/\HD<2VT0*1J6H)>)
P\>GTNMK%UB@!->-6I?J@<'M2I5.YU9ZAV/@C+WSX8O'_V\4,(D\=FE<^L_XBF6H4
P(=2#_*5CX9\5XK0U-"TW)DI^L1!<?:Q,"4-#NQ,<CJRQJ=?MV-1D/"$F. XQ,/,X
P-&.(IA1=[Z48&J:(J1Q,;;:%^E,0K@Q[L$'[E=G#*<?M+ 43H5J4=;-0.5@[_P; 
PMZ/>>J2(,&%4(#""8.8U3&@%A9Q8LF\E!6]!%R8*P% <!$J:B+C0K;JLQ$.#F@OO
PYTBCU\[N(+$2\(EPB: B4J=V@^YD3]%[<F0FXF+UK5G_^,%P,ZS 8M*JN!1_DMZ?
P[!HT5]) &><#VF!PM@U_MJ9$TSLV[:8MUK1 J;/).]("YG*C5ZO'Z=':IXP4#$!-
P"..^#T;HWX&V"[Y0JW:(8I(5U!S87X9(EL/#--G0,F/AU^JG)>AS8H!K*9*/@*@ 
P$<*O<IB-DITQX>+U@\VF= PGT)5KL'5LYN _*72C:6C+8#I6SR0BZVN0L[-;A3I,
PX#>]/WX4F.01;EQ.;Q-:7_6G<=.I.3'F0[DDOWVNM[:LCRB>E3T\0R)^(=>I2M-D
P96_CA-E09R5?[6';#JS0[=QQ6;"[G;*@'.3/5GHQQ(7=GL[V85AN, \=GZY?? A9
PR[8,QO$-$DG39KR/J(:4WNZN TY"H6NM\SH&<^R!8K '(J%(L: 4KB3<!_C#3)1:
PBW]88ZTX0(5TDO-K%+[O3A(Y4!Y9;3?9LM'"$=^MR@8,$W0L":H^,>7>[R%>Q.^Z
P["BEG14E.]NM1)HI$#3+IB6#'-&H$+%>UH";%$CZ)U : _7E* /N"IR=_6J@$I93
PE.Z]F)1JPQN-TCN7LG&9'@VQ620EZJ-YY0GN+.\/E0F&HBQ.5$Q(*-^UHXD\E&>H
P:QA^IO02\$JO@8BZHH[YZ$DEL#<&-3=L$[UTVI.0C,;-D[B5VS@K=P.LS[U6!!%I
P<4&I!U:,;!<4?\Z93[2"&;)--S7PI!&%_A23YVE*M?..LXVTPY[.3PDGM]K^9W\M
P.9L?WO3,U(,!ED?S497U+27[P1Y]6B*DP@$K2P4YS_PAR7C(">5PHN;-%-O;_^CX
P.5#$A<+]LSV6HT?^MH&?A'+CZ<DJLL/^(&PR,4&$$AK]M[WMX1FW:,/E=67S"?F_
PI638P.HLL15!Y1XQXJX>@=DL&7.R]V]F?],5N@]P-#AL+X0L?FV7>+-0"80P/[_V
P0S6MI!]Y[BEGHD8XVH51#PFR=39(V1)0KEG Y+RZY<2D9JCO&GN56<=B]<;YN8>'
P]NLB[, BD2;GH[+:SZ:O1(S!!@!?\CJ3^X1GI]:[Q()0#O5L!C)V.6<KN.OXN+V2
P.VC]:D+%LYOY),H('$[*NLVX%"K$;]W")U'(P_^MG9)@&OW-<KYUL5"#%':*'!5L
P^6!1GFQ]VKT.TE-=,%3,4Q7SC CPK:1M27?RP"5'62E?CM[Z-:,CQF,7@_67O;)L
P(T=$)BV,Q7YTRJG]]/U'-)U*07ZYO>%RW.LB&CO,A:H-0@QUAO#4WGC+2OE4N-XH
PG&+[$MHZ/!P0;I>A;/Z3U4 [6WK#0!;S+8A=GFG5!%,@W)8ET@]_+.'I!R6Z6*[,
P>=3O3HMO?DE?84E/9.:-,U0@,6VGQ&X"4*UM.P$0#0_9SS2V[-_V1,$ &=WCJ99^
PLOP2S;\I)*I,64F>4QUY\>JV0S6)R,[+V0)"((R)&%Y(SE<UX_N-@6D6_94FH5WO
P !;>H3S$5YHU)O9!/-/;OS6QY_2=$U"W8R6-G>\]S=Q9=#>X?<'5_=T6=I+CUDCR
PD@O8RNDBO<G8SQ.07WG^F*V1?3@2S>0ZDB:-[D?\5GI/HE BOU5P@^WH>FUN2U(:
P6NEA/TQH=/+/MSB_*#G_;UJJ*FT)KL@C5D#4J?,LRUH)<0K/3$[R[$=+60E2_Z*A
PEZ'/!P<==G(X\>-L*<8X+-'+CL7I/M_J8?5!G0'3D9OWS]?^@ARK4L>6Q\.?-P\Q
PNSSUY9%%A:'=D(S?&M>.)W8_QVCB%F[%D\-(*-$>V;ZVMN,\U\BBOSR27X9)KX2'
P0>R1F(67B=]Y,[^-^D(+"\*I'J>TXG5RJ<'$4=T[JR_P0^9V<OID0R-.P'3L;2^^
P_(#4B?)@7P#SIIYB>SIT;$ZE_@[IL0U2S6S9I,?VH!5-@=\(4[V"NOU1R7 *F4:C
P6\S(T?J!)845+KT-MC%T3N-J B<!(ADQ<LM3YB!_%&=,\;?K,NRAQD? Y?" ; 8E
P@-[(^5R!DZ@(5^U \K9XV 5\H!;G,*HK*J=!E^64ZI+HG(E2O^4Y"E.J&62M(=).
P>!EQ*^4"+^QYY:49SA&,%8!E++\R-O[6.4/&M)**;#U*0H[V?PXDI[-*_EGJV+7.
P[6*_HSSNQ")P_Q$:8^(/'("-JWYA_#%/E958%HN]"$F'/UY(R"GDI45V%^+'+NO1
P"?&FDI2MY;#E:FI;RZ(4]C>)\[[6JDWL0OBT.VM_&64N-H[=3M,K=^.#CQJ*!-KW
P[)BE(F(+[;-'^I.=]0?-SF2 @#-)EC)K\@^W45^"VWF[A\-Z[1OJVO'.E:M-V0=4
PW&9MO\FG5SCBE>@4=W5LT30RC2-61]C1E.^%/+#'63*>,G:^PC'2.<S@+<$G_C(Q
P;9U__Y"J5^Q3%'=MC_O+;17-@&GG<VI+3OBT8=^<BQ#HHF@9%N?Y7"C?=<*TS-&X
P +ZY^#&NU"CFIDZ.S'6XXO<<_^@C*YL+N#ZF*><%<+LM=EA;!3A&3(3RHKDYQ=%[
PG<O$!$!B2H+(VND36"I#VJAE'76% F@]I:-]7,<SQF]_"'2 *(_O98#!2$JC&\ /
P?)'7<_GJK]P0?4H^U-O?K:-)#UI[P0 07+'IFFS@@0?]VD"*ZAOXHV2D %8A "G:
P&I:C,'"<1P'V7.\\7<V!*A7;%J/I[53B"RW8N=)[M$V',WOH5%D4#\)RHVBP;L1B
P,L?OMGFVN6AY*N/]A"D6*-RR%&I/G?6N/5")([>L/040F*0Z\CCK;17QZ^>!I;'6
PY1Q>$%V.6TW0*H^)B%PU9<8H-1M'MS5J/@.7)".GP-%?966<SQ2YSH,/X-K**:"T
PX[?=WW&Q[AQWGCRF271PP;Y4%K/#.X;;\>]@ F7INZH3L27DX9R3PF481F.M[])0
PT)[LN=',;!CD^:V,G1=A4Q0N4DNKNJ*R6N*]&A3"(]&+[^YVPO]7QC.4)0EE7$$[
P ?;Z=6:1(HQ,#>X5FX(9FZKH;_]R54O#6L1J9@RNIDWQPM?B&AT$.'SXNS>E ,CM
PL/F(GO;PN5,3 BZ^@\TWUH.7MR?=2O,Y"5V:TW3&[%6,!P^4!AF.U0]SDS4!QGM3
P VKEG3YPI=CSC*V?.:LC4C7\[)CI'D>GT?SD=HO_,4&^*0!J;-CD84U=HRD;1/79
P"\V2'PDP;=V=3ONE00? 6]C_I+KT-5JI'N+NGO5:!/-9T$?]6ZPU429DM^;A*W-]
PVXYJ/^2]TZ$D8ZS0VN_++H8[#U\8-GB@#]ZY2*7F[]]P&H,>Z4"7"TM[8V*!K=SI
PD)OJ",46&-AL[U+FD@#F/X@M=*5A#P*^ XIL"!4<CQ")XPS!@I"Q$B<D26(C">V<
PD7#K)Y>E,,=(&QI&JAH'?YM?4AY9\)K +_2 BO1\#)J WX/P+A/+"XI9)W4^\[>^
PVDA">4Y><5=BNFJY'K'B<)G6(T [/ L!$0'.R2A)'K 8WY 3J[NS"0&$L:XXRU0N
PUSNOUS=B13M),I-AW;J2CV?#J-7K]CZT_;B*(>9PN1W8D#5H;MLP4YV)G3*MF+TQ
PJL&GN#Q'0T$W-(1[_,2<TF3&N0XV6'.#G"%1>+D[;N(QV[<D$H]/Y'\U.Z&'B4Y7
PN%U,_5Z]VHVI5WHE&_/1A99%K\0?8')439H=A51=C<!W:EIH5-YLFA43-?5W@(>%
P1S<B>=D9_#N:F!%G?>0:V+*WR&3%D''?4"LBK,H,&3'=CS*/O?GOB95J+]IJM:.W
PB:'ND2]^U715@(QV2LL*KUR/69M>Y&])8FQ]>N?0^A)W5?JX&9)]GQ_HOF&JK-31
P8V7<PYBR\&$KB%A6D59OU/6'H&5+W+/I^<AOH0R.8XBI&!7.0C0F;)GFX[OROGML
P_QZ<TA1PIJ:MB!EC.;AFA]U#NVT!PVG:A'L\?,G>E"V>$$\:T>ZA9T_C^FDSFT=P
P_(=0KK]5 L!0XG;;>+ZJQQ_K$TU97AE<50W_",IOG7%;<X?NB+&D,N2W;V',M!D-
P39+JH9UEV!P1R\REG'LB;4,>-Q6^_K*[Q1BLBQY_57N_6EUZR2MU.RQ9II8A'\\3
PJN8%78YGK.S*/AE4^6<D:I*1;T7_(0+&WP$#U;K"Z+-L/3W4=)_\H8.I7U!6H$';
P3V"#]%Z94+&QZH9QF-ZQ.*%UCIC?RX6!.?F^.JW9 -TFCHM[)RL8'ISYM("5-.K,
PE#+[C/R"F/HR3P@LAVE?ZKL80,IBE%, S(^I0?V?37(RGW$;:B,Y#K=UMR;G\=--
P=H,-^53.:RCVXXL<BP)FEDX$8>^TM*DON'#)XD%X6[]U?O'[V%)TO&@;^@;A[*S.
PN/.ZS&*9PSR(/WT;;F/+MNA6%IUFZA![[,?HFT,Q-B)4638[ITJ,>"'T'9D)3Y!]
P(69=&@IX7Y;Z'O,'4&43=':YZCX6-[MA.7/4?/:+H45-1T."=^(U'^A]ET_D8-X/
P!F@X&L042T/N739[3(0AO#Q05#>C67TYU4@T]0=Z!E;?I+N[*W];R39 :O X>9?J
P2MV*%%_EB6"?M1/$2F.@ME4!8VXZRO=D^J6AY_&B:7ZWJUJ]=@LW5)ZZ^X/:O?Q 
PKU+^QXEL&IM!^.HM .G'3KEQ)V=,T70%'G/^%B$;BJK$<G#P91OE2R/RE?)A[C$Q
PGC1+&6R2'B)VC/!DD:R^JC'N%=\Z@>1QT+E/HFCTCO^$&8%;=C68>D65W)U6[7"H
P+_+3;EW?_M.L#Z=D75;URKGZN+^&W2,#Z[F'EJ\IBOY8/^@%EU0];C3@W:LY+[*D
PFU#S1DDK-MD,Z0AV:*\['OR:E#88> #M&=P1)%G_K\G&%2]JJ#1.=%O0P,>G()V/
P%69+623"EBN&AXEE9TO@F+O]N:13RN^#7E'FCH]-Z!/,(4W*F[=)V)Q:?WRO4X."
P5_M7S@X$H[RE6VSDHW''?J\$"S0.72CBN#QH )-RP[5?W_'JZ&<M..FP%G@DO1,F
PQ_3L:V9#0!Y-X$LG_<4W5.@@X*W\3[;PU)];I[DQ#5G2_4^[3Z>/PF ,4[/0'XH'
PX,671+@^MA(RSN&LIZ/L/ >6E6^FVAP%]Z]WJ6,[@N&4E2@3O@UX\]:_CT&'R-$]
P).\P<W,(T1COLYR!M:=<4=^N(:BXF,N8[<J4:!8;FW7F&_"9UAH@Z*+U?B52#SFH
P[3]"]>9A85%'7O@ZI.'7##'?)N'8L+@VLB?$/H5<IR:[E!<2FY1!UVSJK,CU7OF7
P:];3^RQ1KI/.U(ICSV*H>_#CD>_@6(MVFS?WFJW>VP$Z_W_74/4\QNE1FFDH]Z"-
P)%4RT'/BV [3R4!?E@!,X<'S;M]M OG3SUKO)<IFM;)KG L6BSB!^*-X6EY&XH:3
P;_;NMR>QJJVZ[)B>]B'=V,V,N+E7LJK5@O:3]%9/")#=\61<(&_T)Z/N3<H1H2R]
P5")\:@N]FLL(8.0%UT,FMY"[U2:E1A@X H]9R)6F&SP",7I>2&^MZ@\<?%/<J1[]
P4:PP+:[#*CP_N:D"DR+5W8^*$:B.K>VO8\XXLPSQ_LXA0#/_-5_<!@%:"2)0VAHI
PFOB/L*NI[2T'5F8$A19>L,MP5\W/>/W>==7S]9_GATN?&0U-/5_IV08T-$KUR;(=
P**\:/$U]YS?ZEO038Q;112KG&46Y',"B1VGA0_MB^Y:TSK3[=L13GSC14].9O^+K
P"0D;$'/][.G7*(')UOAZA?VQI,N4EBV&#/8U$86@L[ '-#2%=T >F#+="#9MQ2Q:
PU,GMIHJ*V(=X_.P1[M:"T_ZBN?U.RE.M\3:+V.ON5S7@3:0XJ('H:"SS9M::SO1D
P;8:7)6Q&%>OE?;/#MICGR/;<RY._W1Q?(I.M+ =/QK<: 4UCXM<:CPLTG)Z_>U2M
P_W-F (1R6;W?[;I?7LEQ;JU(JV.1(+/:T[D[E!T@$VDLI($)]IB<6]VP:LN)O%X=
P=M.!J&YS*"Z++FZP!/'ZBB8=1T</U[>H>*5KW+0X^K%(Z@_?TMXE7T@/VR6Q><RK
PB%?6ZMFH::&"%4<LG'U0/6/2B@#F3_]TV^ &P!I(B=_!!/U<_!ER2'7H%DYZXT1F
PGVDF:('ZJ8,2=19"-OW0?^)!\LX>P(+OW$>%:)"(Q!=P0K%V+H=/U)%?/ 9U4@_Q
PTU/EO_%$GM<(JG+2.+]-$IV&]D[T04D7M^6B/6+I/*#/&(E9H!@3>#S=?QAA?1@$
P%4[N.'!9(46&3CQ"7(GKBLO/&VSPCJ;5M@'"86Y])'"@.CJHJ;O:TY6C0)CU=_1^
P&^/?:+_X7YO'WK\Z-0UNMDAX$:,HL-:=@UA=9V%G?]^&SEUD#:% 3W"(@N+"X,NK
PT=HR84DBTRY(W*8.KX02"O$'1%@6+8B+\#4S FX@4@S0MI'^F0N!AE__MQ@4VFEO
P^JV<W(*>1*C=H/T.Q7IP:!QO@XN$8(C:X[&B66P(.%2UZQ/S!VF\#DB8BP3R0*44
PM'>X@8*+XO;@>:$YD]X'P>C]TJ<*N0X=X^ZDOSPJ9,$&4U!>5_455J?#UP6KY[[F
PH:V^X(:@08+G&G;,G71[\VTC1$$/B3J^'4B1:5Z_T#!\EA0-[^TRVK[1OX4(B@G6
P=UO'N)=\EWN3<65 VP>26,@%$CALK*^1G*^\26B/X\XIS$:9.I_9]7)29WV5W UF
PUSY"J'<*/B0"0.9;4T"+-+2/^^=(YCH&A<)W6:.<FRS?W#QJ:@R",CT_XK>[9##&
P-=&/*!<)^(92/J([453_6,/\B+M]W"3B]3+)@,TDR7:1QT0(;JN0MN0 &U&^:C_$
P6F,.K2!R[U_%T8W)[@VLDS62I@R)XBG2)L\YO%$#5"=(%'J.%_J:?!%TO\(2W5D+
P0[_Q79Y!89]DUKYEJ]*I%/>:8/Q5;@S (Z+A161!8-[D)+CK-5ED6US[V@S Q]I5
P<W9U@C@K1&TJK6@K<R,T+7%<V$L?)%IT-<PBWXXW?O>Q=-Q?.W1"F+[@=FP,BF1D
P^>SDHIF5._-Q::]'[=2Y@NTI-91Z>0:TLJA7OG+86^@WI_/%LD?RTE^]I]TG950L
P#:\D&JZ31VQM#3!=U^?/TE<Y)3U>',Q;5%*O%7C*3:)3!="80]7)VZY/XEVJS<?B
P_"@ 7/$3.D?N!8@>0):0&OX&$I)#"44T!JV],QJY*<4"%RDK]PS#!Z.$I0Q T]5W
P+LC-3!<X8!%R2OXF> HW7 ,C2V8$[)X2V/UT\"0#'5DL3NW]G Z!IG=_I#J&_+$J
PC6T\"ZV>4+&PH9_LX7-''\4?HT&Z3"GP<&6G"73%MJ]':9B_H>T*?+:*;5T#K\79
PGE(W_5,N-K*N@)1!3D@MIFEX^IW2RZZ3K)J6E,8&# GZ5-",QG?O4[KZ@H@IIZU.
PS")'._:]C"LHL-0]]X@Q/G!_\)-'1)TP^/6SKR+AO84Q,\O;?M9.Y0I#U8DZ8731
P4VDJR2J;'7>\!I0;TJPE14DH+5IV;Z?^8'2U [T8@%>1<%2==-;14-M,-;RS*NZ)
P:M,AH@UZ5LN=^Y@RJ(/7-5YK=D2BOCZWXJ1CUJJ?')MI/(DMYPEY_OX5JA,) 3GA
PU/G7*J/,?QOSC"DA^Z/JD!RHP%\]S[0.;O<ZU]ME9UBV[+(YEOK&6\KX!F'X+0')
PP=$RW'\)<2Q=.UBBRCH/ 6C?]I28[P/M!(GL?NC[C=")TL48"0Q\GUPJ-<Y(';(3
P>18PD'9O5G.+SI$?_%Y]A-(?'WMJ/EN<@U/F)WXX8Z]H_WAP*6):;5JL(-V[LL !
P""0P+-NSE<)[4E,#-8J4C]!I_,AE/\*0*!#RPKFD4YTZ$.2$,*\6V%VX'QA"[F_1
P41[/]*K1LJ"?V/^W^$JLM=@1I=W(61&=.TEL+,>:VEJ_$J9XKJF*4ZE]E0-CD0'_
PJ7,'H,VU F>;<=.U3&+B.>5P<RMCOM%LM#81/;.4SPF9,+^7H:,\U47#\0-;'E36
PI\%/+HJ)J$\*9%XR3A/!X8:R[V=L2D.]IC.RUW%>=KX<J9[PHI,)W5>5.7VR!L<L
P\?\R15XK;R'TVZFYM)"GW/[*-K+;2QJ$FP^4DVA7#-8Y[H;JV**7G]@IAF68R[?+
PX*5]@)D_@OV7L;M14W=&FP:I&H['AY5?2#)/I/\_D'_-YJ5Q/J_!8._BW_Y&Q.IM
PU3NBIQ!I:M*,5VG^B22MK ?*;EV?T&IT\G/>NO7:;W8+GYM^Y+0S=G 4W(+UK4!T
P8,'&"J$^A!DR725H2E:"62TWT[W12NY[,=-U?3^J!LI97?]^!K/^D3/-+NFF.;>]
P#"P__SCUCB3RT+KMCZ'AF1+5;(NS%5@5MXI]54Q]"S76RS&P*F#5-C-$KZEUS;E-
PF$&=>V0B*/+P\&RVT]1,E,Z!0#$;[/XI[-A"X!4H<T<!A+.@UW%"$3!6?1%0?4IL
PR9R091XTLQ-EI-;"J4L/@01Z&8[O#0.KD7EW@]XTP<R52*GH*_N@;7D?EXSE28^?
P>B>"ML>\L>ZN";"LQ9(H)_RW:G\^7G7%FZ(3[9B\F:T]]Q9UI47HO9V8BJU];??W
PL]+,-<(#TV885D$65BI]9F2J$I7?W%'.0">?A>KP"-SU\<Y)\5CWWX=;;(/TG%TE
P$?V>$YH4?ZP%$]ERT%Z0F4K^\$E797N=3VPM-+6UQUEO_7EA+*K 3UNVG#N6Q702
P4U#"N#6Q)"*EXL55'RZGL["J&.-4XV91:9R<XTW:ZJDA O#6F.20'!<FBC&!W/\P
PO%:+1/&&F$[-2=P^-9'T#/'_L&4'G'Q]=N% (/4WZ?^$#< 9V_U1;=_3Z[^[8?\:
PL)!J&]E(^G^"53])FL@Z/+2U=8J'5W/[7M64;BWDH"4,*8FO)BN,#2&XLG%-=QXN
P11;Q?X&6N%*%]'I,LF;RCYI=$#@1C-+]PQAWD-UG@2B.M1]M&!7@BS"O7.:B-6=,
PNI(X.-A\ 0%J!X-%5;F+P@8Y$CA([54BVG@F@B4'AP'#P"'S1;<)03\%6.ZFM-T*
PC?,$P9@4=BDOVTT1OTJ?X"[DP*#U__82-/X 0YQKH+^6N'!8->E1>6-66=-Q5A38
P7^BZ<DZE:++4;2@Y=U S^OSQT&BD4_\V70?V!=0":SZQN&MG35V=M\6!B8XAL@O"
PG"?\\,9_YNEA>J9[*DQ"QS)A'C-<O#E7=-1E<)J_[*X$EV:HB%6=#'M4F'>>D<V9
PN9%0I'>I<^?&AS%ML0XCL^X+Z2[6'162D5K2SH*:C7?U'J2G'J'79UTRP,ZON3,+
PP&+][;: DIPV8=:\&(/HP^\+K0T0ZE^0J=D)-DB:$A8!X%N"DQ2]VL4"Q:_D^F_(
PHG3S+S>83>+/HP=G3/J"1W,1F^>V[5Q6D'-"LNQ;8#55=IT:[X$I>N_B_?#.)C)+
P^5P4@U0@.G][3A^"93[O*BQKWH:G& Q)E^Z'A5WZJY]TYAR;R=*9;'38G(1;T\<T
PO"=69)SZ=4'46Z'<K[=5(;J1TJ%-YL3KG[-K;TPXPP1,"ZWG@/>B1#N,USQJ!!OE
P0[>!^%H#+>*DZ>9'7D@ST>E/+3$ZLEL*JA/ WC9JW84I; =<4(ZC_*)WXV3,]'*?
P6#+-9;T6V[(U,PNR_G.P2((-G1^2'IGHG%I1-==?I[^:9M*B@OYFS[72.46N:+N+
P!D.>6,:@+)8F+WE9,QO"1A:.T2X_HC=50G)$6L5,>*S8"(Q\8":LZ+"\P6N:!A=^
P:YPK:[K&&-F8APCN>V#0'[-GU4 L!TR8O<[+W5=?ZOFJ7U"3/1G_0<%M8'"C[P25
PV4F^N?.](:<QI.2C)(?S>RDNUPCE"S %NAHH#TW:ZTYU1-X,E Z"1_EU59L?6*TF
PS[RD#PD206-@4RF&[P%\PPK".--9E:*C?&H*N)X;OKP+N HJJW_ZE(\<CB&+T7E<
P)J0HVHAC<(E+41>?0UT9%@=%"B?;TLD@Y):5[8:I=M'6)2AUM_SL@2X&R[ FI$FN
P:P#$[6(#E<6\+DN6"C6E3\ Y/Z(F."CHU/0$IH=.E[\+8)KJ@W1F^[_>?F&Q&U2)
PR2;*&ZUL-5!S.V&M:L81VWBIEO6C--7 +ZO>KV!2 VD9:([T\HHKL(I_:O5JY70:
P1-.R/XX=]':RV@(>,O/!\AK#C+MV"-*W-] "J1WOW-*7:B\,C#@=(<:C43=1HQ^Y
PUNV9*0TQZ'*];-CY1A>S'!XM&H#:>]Q:/JXL&!8;[Z>O/*IYLV'A#?WC $U&?%U[
P]-N%F_OY28/SV>(:(C%PR/I\(?020>NQ+O0VE,B_ "]D::DD4=PTM[B.2'RFHK79
P&GH"Q"-*XY?BF:,0$P<*#)YU-&@\DS8@6@@N.Q-C=QHW.I(WEGXNZ]A!S&4MD8*'
PIW4>;/*!YALHQUQ5T^MMB:X<9:)BJ:64X.&[E$R1)/A9B :4Z3U8IJ/)>?SOH\3"
PY5XX\NAX&( HO3\>J']V.F[+74;,:3N5^P[-?D  WO 5]?(8.SM)O7"+%L[-WTD:
PU:L:V[]@\^2^!0KH&8P=L.=_?]M2?>] I=OT1  6C%R$ 31VWS0Z.:M/X.Y$;)-(
P5%T.!'9JTZ5C(7IF "8FXJ,0U03^) 88O4DC#*]!Y:-TR3Z[=/9%M+7UOY@P$BU<
PQ12C!7"KO:Y6W>TDCY.C"RKYM]O43ZH!_ELEBB?S]="K'$3Z))%+& 1%SL4RDKO^
PO-W"FMIO#&@P@_7JFR]_QKWB+E:<FWXJR ')<9<K6PJIX27)9KQ _Z/P0/HT])S*
PR=$6M_W.YC<N(RU24>7)1PH5O7!CQU#^APPM4CD$NH.G,R<+G$@')5<R<\,PC7S(
P)7F1#'^D]]P*70WX'\ZB/JO,#N2<*J+Y-Y P4S=9[O51Y'PYOD_?PH&%]268V6PK
PF]!!W[&>R#?)NM9\F;&1[3<@X#6/!)";LF671Z1'/8BW6[#!:\P6#091.Z96NRD'
P+71>B?+K1NTE"1QF'8HFMTT4(0>;;<Q68.NU45L@*=Q=MWVH0-]M07^64S0W=^:'
P0:'<DUSEI*F[&*8=87>-K%AN!F&P]X[,3740-/X6^3KE4R W2-\QRV,"&FX<"G>M
PW[\&G0Y/CK<QUR\#2IF!5=,>;#8W@WZ_$[Z3,*()S48$<[W797.EZ(YCF1KQBU#$
PII#B*$=-09?+@\#ZQ%#+'Q(Q:%$KQFZ86M6D\R[E/0!JSZFGJT1\8@N:$8G]E*9,
PP+[D/"-(.:GD?.#]6:*,8:2OG3.%YK:\=AW7).58I3T'8DK^UQ.D4R58<)0UY'T(
P06_"4QAZ+.K:^.5Z[T$J+'XSJS(HMV_,O05K']?4[@T$K8+$.H:0W<#)MP_@3^CE
PCR?N/&GR"E+1LQFF7<:J(H$N:J)T11,/JY7QP)2A,-5W$Z@/' D?'.0LFDXUVE;4
PF6K!]IR-#0"J'<W[[>H&"S80J4]6T3Q,Z$!<43X]>)U/I+I''8 PM1PYP,S4T'.4
P>MG<*WAEWHK,JGRN!2DI!B;J%U7Q7R@K@(/"A+>C3GC,]GS&887CN55^3*>LW6J!
PGT7TVX57]0N<^061"-:;7%V)=5-;390J+'.&??"6>.]'U$?^J>V0'>3.2_@KHAO<
P\W@Y!0+[P#8[,A;MZ'\&:C1BI1(GJD@:8)I3XR$R]T:-$$R6UJD1)/AI1O1I$9*:
P,RGY$>Y<SF8X.]CK?@L\@7?8DA9!@F"?=4O &E 7WH%:*O<DVYZ'M"AA<TKNS:7)
P+(P [73L37%P%/IUI7?]L!:XB.J.^$MGB3(.6#KI'K0,3[@X5 O?N2,RUO(6@3V8
P7H]J5]?YD'NBXE4;%QZ+9OWWL5A$?%W7!WK^6,>4U\U$C?";T9%K)J3=[TS%KO[=
PL7?_=^<YO$6P#=_9[$:_#-1SMS_X0WHZ*$GZ?<[A^BLPN 'AR6<LX$KY$7Z@EX#R
PZ?2U.*$*M.I^%*:!)]S9]9G"HLQ*3FY9+%P,D1%SL%(V7=(6J@Q]S-++C$%!E96W
P)'2?%]2=RT+ABP5\'%=A\7K@UYI0(  6F.D-( TM_.S946]BH0L[1%?O'3-BI17T
PY5-3HRCB@GVK+U=<6UMCDXG53B;!+Q[S+& ZJ*LID#P6AY&;;/]C\5CSEY(V?ZMT
PYM$RT=6')I-F,/7;!\AO"_9O"#O.P@G&CTZY#V=J!@A0/:1/.-$6*/I?R[%5ZD0>
P7\N)QD*PK&P*\GIEF4OAT'#*,(GUZL'#]28^RS)SB2R>"1^50-N7 4=.:AO$&[F0
P9F_$>J5R\A$Q!F.-EJF5* =?W[;=#+(=&?Q#]F0@DA=3K3V4G2%CR0HAN(/UVK0X
P>0^294(D?5OH5T+X(\A2GQ6R"5>?S*EL ;"H3#6F_KVHFCD9%1*TU753GUY95C:*
P4 E.62--^NWU/YHF2=?J#H<<VOX8%&5;W6:05;KAIXB& \C5C9TQ !:M.<C"CK@N
PU&(=&:O49!%I^K\;<@3)IB7NQ,Y<UX^:]D0(MR FX='4:[$/#*#Y-AD-F/ T0P(C
P)KR(!P]E;;HO>KZYX&P)OMVUVU,E"R1H$I);/EJN[[T,JGY>B9!+ L%$Z"RV@#W1
PNF^560FR6.LCB%,,7@X9&W,BRQ*PKC>84>8V"4K8(!GBC19IKK:5$S\WTC9K0!$H
PYN//1G4]=N58.HG;#HW_?.3AP1U=CFI;QQ;7YH1(RHX0!J+M$/'8"<-IF62S8?P6
P![] 7$3]>'^@\+M2BS%60\RLYG 1HQ$R87)J\>@?:6D7S85'[<'>O\W1$^U."DFN
P=YC(/EYZ73U8M&/%ZQ^T,7D*ILQ)1.@M=G@H2WW319L:8V@RI65N1BSFI:#!J+0+
PAAD_P&I[ A*CMSK"6%U*##9ZA17'1B7+P3<@V,XE4D=-W2=EB4A6ZT-59U@R)Q',
P7J[B<H7WP\8F%7Y':0 5RZ$/N9RY@-S=S:ZX-<J5[+7%=TLFJW-ID8LV'N!)/8!N
P79$L;SVIN&F28VE@ZK]V[B;#*:(.Y]G]4CF2-X.()GT(?>EF?-]XL,S<$)+]*3C1
P2)[7/CEF!C1MW#V(&9%K6P'\THH4>8F5$)E?)<Q^%;7F&#0I,A?EB:#< ,)1Y?[E
PPB$RKT3]^I"$=0\R6SPTH#!<7#EAPNI%+!GT+?1D5"TUT8[/\QD-71MS+J#D*E@F
P8A,YALH?G?W[[=KC!BK2?(Y08$J3PUJNY'3*(ZR6G.23.J=ST'<(QEGC)&#<:YE3
P0,5VED'IKO./*Y6B$@)I;FEG(93IOM8D0MBWTL#ZD;&.>N_'=NIDIX>UPN2I5AP+
PQW<O4?/&D/IK'+GR[[F6;[GO 83TWMG>UVM=G!1_16'\\.]8$FD>V/" -S!V#'AX
PQRWGL4<'5"YL$ [VZ7*$[&7<&KS9,X)_1R^X#P@#JL,OAM5;RX1-20G=)G3P"[4U
P08"QL#0*;'(?:Y#N8O%^O!;UH/G$^=F(L> 3B3.W,3XR[3T-).I96!M<K^)U3(BT
P1T48&Z")F+ L_LO%=8+U>S+4V.'#KGL0GA_,E+0U5Z"KDM#A? J&CDEO<OS.)T]4
PRN.>DF*U/I>K\CPG =*SHXVM>MS5D8_-TQ4'(_UT'FF+2;R?_UT*2MJVU+A!:70[
PP_Y6)<;;WO,VSV2*KK1\_$$>P*9.,KTQDUQI(.+PSW&]+';O)#ZO$>S'+$"J19S!
P7GL7?ECB41&6ZQ!!D-O31XMND(3)MO;LQHP#YZ@<9&/$!#14D!"-@#$%>0DUF VF
P%%;7-QN*:%Q\NNC!1T7Q>J6N-R"X1L44D[89_S9C"@Q]<V=C]TPER"1VEA7EN4;+
P,N@8D%,<'_"Q@C[!KQN^<6;A/3,5UQYG9'-X(O2$V5_F&C.KN AC!%M4O#5=8HY:
P"%'HBMFB:QGQSB&0>^:Y8]30*4+-(19N%AK 5T_"G =<_%G4H27&V'S\G_'3Q:FN
P]:NI+\^X8D\->^U!\!;C?#T*%Z( 3K&@N>1E&GO"5B,GUI@B6M>3,\XU/7:[+OOL
P%(6&R0P1WS?B"$F=%G"8C.?$*<11)[?/QH!522IE4!H#4'V1?.=@,(QII)-(T-%.
P!5R!%3U2_$Q2?H"PIMNV72,;X0R\ZH.VRXUPHS4H&ZA;QE3G\W<*X9R:DDGY?^WC
PS7APIRLTA8=(BE9;4I)L%EP?.JAFR-W-KND41@K)>G&(&7]"!AYPV&F8NN/\I&]4
P&GLYX=7Y*>@%V#Z1T##Z<=+RM%_=4PLT"I;L.S/QZ ;6[ZTUX7%"M^X@;FEE:'1:
PUSBI]K%K\-;#'VX3E?N0#-00"R?8MMF!Z, A#F2BJT0;*R?6; BGE1)M"(W14P?!
P66-R?*;5 9 P_T,RDL)TH/&Q'89A4DGELIY[HI%HX^0FG':(&#-(#TA@]8(R/OCN
P%)7"L%4Q!J;W\;K6&.([4%8BCR',?X'."AR"(5V;I$2# !+7E>@-+]=L)M9E;WC/
P>C^N 4%3"CYIP?&AHGZ],U8-)B[#9%FA3PL\8,(TO:;*R=Z"H/P[8*V:@\[*Q\,1
P_K3^.;60*SS\8';NLS>']"?[((+QA"ODB9,!TBAXC$<Y/;F3"7KA)FJ?]R<P!J1=
PHO"QG';4< :&0>8(S1=SYBGKES:W$RI'%FJ:Y)*XLRN2\(1]Y/XE0)M:>__V]ZS@
PC)8L'B%'*K-D5SI;=*W9W"V;J+F6^ )Q^NH-@+I47*N6I:9]DH,CD[;E<.S4#L).
PC_[-=^ZB4?P.GZ'%]K.1<)9L>G1WPB+.&G3B0]GCF2)77"0I.GN_8C)Z,,L&5<<[
P89L_#OTD 7)#KK4O"G:L+FGFRA#42_,C/YI^H\*R9 R-K??V/(2IM9V/_J2G5F1 
PXZ!R.$,SD<\S+[K#&3!&SK9': 8'^K Y*TZ*.MZ->$O=5D?U8B@6V@&Y&V&?LO?\
P-V<R%E>UA#0;@2R_FZAYZ!!">4C%]/?G&/BH19+W35W:OF786PZ[AEZ\1* \2A'[
PX/][ JJ=?[M^6?6DKE,I86-M:R16%9:^J/?99A6!I5R<0:43RC2D/W[HPWL.+".4
PP@E[3@\F6<\+2F(EH-HPE)4&A2.N:R,1+5.\4#2-@*4:+X2,:$!&J9Q>*2\&9%>)
P&#]^O,(D1B;M#<2P#\K5_=;6U5J5*+>H5Q,>Y]F:BJ[%OK"\:L^TO 1NW6*HF':I
P+_H<&8?QQ<'%D_2Q#"88!)4=V-TEW0?HE_*"<#.^@"5/AZEO3E\/]@^O:4%5%0;I
P_#J7EN>V%*FK'$6?NAL#72/5-SH'G"B2C\*6#Q!57J9FHRS5L[B;6W,,.O>Q]TN5
P+IZGEKK?EPJ]24#H;6!7L%FYO<_*"NH^,L[$*N1B/&9;%@HH/+5&)%;3?[=]6O3M
P'_N!OT2"?_969ELI9+VGRS91'C TY=B3]8>,F+L&6(K1107N<CO@;6@#UWYWZ.V@
PCS[-/):]YN,Q:[T_:@>65^D]TY.K&I?\;.%UBV2)#;KOUG,@++W*A#5H1#/@QHNO
P$/GIS1$[H!N> F3-8!O5>H#HG?^L"#J_C</$[^LOK\9IIN8B8"I9K-M9W.L7HCO&
P O4A3Z1_5*N1PA4*(1=E;BP.!J/]S$.^T>8QLPR]_.XT8OI"+QFDP- )#7*$A\C1
P,S7R[0!?C1A5;!5]XRC-@;3[W;OKK[?5V4#V '-=KI-.96OS# G[@.Q/J;2WVMS6
P#V^!A7G]7?)+*',1&O?D+$86R>=Y[)AX ,7$N$[9E6<Q_JM3LUTT/RKAO7GB1_:5
PB>]XMDTWN!TY#<;0#6"^6!2WXKY"H8E"-[/PQ,X+G?[\P'N1K[^/L2@?HF*&5C>V
PUE%"45FTM'+*73"L2=:)0W[ET3* \G@%4WJ6]'&AH.=+.J21D-][*=III93;!5\9
PUQTRU.4V[L3&-/V[.^"E*"_\GPVI5!HEC_FBGJK/JL<U8U3PP_KN3'< S+V !S,0
PQ*<M17)A3FRQ11H:O"G[1UTA$1*CX@60-/$0Z0)1PW<W 7AE;E^F.7F=[5M>3)3A
P\DSH!(>\>C=J$I,OHZVX2[[,%_](%GR2_^KKN;'HU@2XE?J+"@N"L,D305$#-^:?
P$_(U[J3"VY+/7_/O !&JURQ\LRN$M)D4\S@YSL%Q"75[K__-2^2E76NL&+#A^:#P
PPH#>E0R.=V\L*1Q'O%R!D0.']\E^F5T*,^//<RR0"&;T(K9T>^/9U1R/<HAY"5.'
PC&,[P"S'K%)6G\=(.@WCOT=.Z/ZS.*/8Y,^:B#Q&4G_[FZ!-/Z,9 0DU"C I(1"/
P^'>:)ZG5Q>RW+@'Z126*8W=EI]!R@1J0+R^'W_!;X!<@7;*"YDT3\(ZA$+'B4>@K
PYC%"[T]\ E];SH?;'("T9QY=CW[(5':]1$T?@'^7PU2SO^3!_>+ @EME>21A!2(%
P*\"GFYJUH;$^B4S>@X^']3]K1:N@?9XGNVPB#XBB6/EI.5M5K(?5?O3]*O9" L.H
PAAO_I0P6\2C?A,3-@]*[W%>8+&]>)>H]4J>!T8*XECL%'16CF"HY6!":KDXJ(.3G
PJ%^.F%W<WT.D4WI7P4I/%OHZF<7"UOOB5HF<CB)]%X(XYJ_1PD!, YZ6%<Q"<":!
P)7R"1@[]IJS1%S@9+%S>)ASK/SZ=*]G)U"AU\<SUXQR8;K['!3ZE)MM\EEPRGI^F
PR\URVOS/W7)A,.\G>TD-MH*,8G'=G>8S(D2*VM7 3U4(8DY6LI#S]4@XSP7($]2#
P<@8!]'"Y]63K&6+1Y2:+]-3%]MC@<W Y;'JJ*OVFR<I(_XRYCA&"?NOMC:#CLM-J
P^\ HQIAG!'D0;-^DH=0XFR8J)CPO,<7;6N*]&[\^+"SE3/DECQ*8PG.RN\LV8];!
P#3*A3ASU:7R):V=<)5$FL+5Z J<3*FK7Y_Y.;$]DUM("\26QN7_5M2%)L&^5TEMM
P#0%MIR"WX_8OL3J3UN2F_DD)-$,$SNKZN@3+PY['&U\WCYDAE<&Y%R$)]U%=7Y#C
P6X]9_!#!L' #N<SY$U)CT][;Y4QW*O!U@S8'>K%^$Q$,^9#0/ZU<\KD89'].KJ-S
PX/.\*=@Z]K;!WDZ@^T&BT6$2<8=,*2EPV:3_.')$@]13MBQ0NOMK.C##O!]A0K).
P:1IE=8A',V>QOLS#!4Q&S2I&(79VMR&2EYLMY$1[C&<XM>X6#VCJO'E".+RM7FTP
P$V\8_/YA^6G&V*>!Q]4=$JUZ$[KXE/[R %P"GF<P@EH(_]"R-'8ZK2K2OJ()0"J<
P:3Q%>-!.;>[1IQF MO]6>S8V9DG\JXZED5P'=47=4L"Z_C3F]_1@%+<R 0',J8[D
P1AH<N:[Q'F,+/1@!UM+]FQ08NE+Z9&';=,:*.+.OPR&@2',1JD5U<5F5<CF[6^TM
P>^BO3P0:3OU9WL22Z'%YP.=-@H*79FK$.L1$"'1JZ&&Z[^0Q6?VDVI[H#56/>.IL
P2+!BPJ^MX"[E#+N<^?O=HK0<)+D4 ^);'A2>+P&A<4RQZ9Z7L<F8L=+@70FF,3DI
P]SMPV 16$ K"XI>-2#-$^IY]N5$<I[SH6Q6B%]@3:P@_,M;J9PZGEI^5O1E@A==#
P**Q3Q*BSINO=]^2G^]-T>A0AC^04'BMX)'E4V!R5OP#)ZJN0F["VPXO8H'@(S92H
P5D ]8\$;3'0Y@B&:#)9A,B9_X-MHI2#OCMSG"2K9(SV'KYFIYAB'=0N5A2^$MU#R
PU]##*K72?/>1_R.;"J$#H8.C2I9I709)0K[+FO'?M*LW7-!/*MGG@:(P"<NU:F=(
P6TWB>3]9KFO*#_C2<KV\IKIZ_MQ;U442X6F#AI$^]4,S$J"2$A%,PL"3!_ *-\.5
PI[)P&?(>EZ&@;%25#JP6B0;#E[X%W9K+8I(J)T]I=^:S>GYOT8DLK69BL@II@&#4
PK_W.]8W&8!0R(C7#:G8U.K*@DSKQI>QD971S-A#_\Z\94?O[86=M._<A38*TE#V;
P./53!.@ET=.>6!#NHQ<(2>!@\Z#C??-F3$P[>.O&F3VIZW+6$]"F165HGJ<Z(]^C
PV*S&<@/W3F]H>+)]/6!5:;A)^B^56]IZ3 BDGWO_.O[X)_YKX &LH8;%[QL5LSK 
P!'V;ZOC<534SZ(!(+3?\USC8[6QFAOT^Z"W:=#5B,#OU([?&)E%V?/S?J*Y;OZA"
PKP>B_<ME6@193?(,PJE_K9(L>B"MY+6Y--Z*??EAI2?J=VYXJNTOZG$=UU+]@3\W
PM_K=XF2H@/V#)8=T/7OIH5>>8(=0:TH&U'T$<(C:NM\MWJ$ 9>7W,U/XI+RBYK"<
P:Z:89;:?KNXFT&9(Y%UA\J#6IB(_.NUC491A$UR)C*ALDD6NTP#A4!C"+QZI:F>F
P8W*X,:ST'Z%MLN$F\M$8#7.#/T531DR_FZIUS%[ "5[C5"YU.)[IO)P)9(":[O$3
PX6OW]@6=[I1<# !Q!]4A<K!FL&V/_^4&-VE?:IAHM9QN#V]G7RV0]U4;?J 5.>(!
P,[?PGN\=(;&ZVB?ITH[\5_8)J4ACIO)9867P NRUV(L&LH@ Y1?Z>$M,%V"\O&I]
P%%[5_I7B'<1;S$SDFC_AX=(.\D<,4?'>7=$:.\KJS)[#GB*.ZRVE7(M7WA7#+SO*
PH$UA%VBWJ*#DS->3.Y YD?T16_T]X-4?6#^J185*!5'(+]DVSJCW7H*SWT ?,'!>
P7B//%D$2.H^DR-Q4X#8'T4NZ+:&,%&>[(9?NR5[7(XP&&"?2<?,2AG"^#IC?#GLR
P8N,FI@X/?@LS$9U.V_S^GB Q)UK!;;_.VY6&+1TS+%?"QLL"'XM4[2'<@*A@F(\9
P51#3F]Z)FK]!G,G*Q%A:[ W'4\F'AVI)1!2#+ :$FE=4I3RZ&0[PIJD+3+#8JF,^
PP9&+Z6%P*:SV.!P%S]!2N,'!*43%HTD"\?U@:^>NR$2 ;JCDPR55@7N1Y6)QU@Z=
POM'+IJ>T:!)M6UVR2P>O[&F=$5+;\BB0)JH5IX*'.9P[0SQX4?MTC5AQ80L=P"@-
P*F)V50>43+ LIR]= R%  J[,7*:3-Y^&=7\$'0"EP$^7?/H#IW%0!Q#3G>AA?TED
P.$N 0N]&OGP]HVGLS!_+,.5.%CN(NE$,4_1#9;_<L$ TFD93(UBDZR'UC(OS6J3Y
PK ,7D5KX@N]. )(J58QC G?6]0VXU]+.<;REVGZ.7MI[,B_RAL3". HP_B"M%6"-
PA1X^V7"^FRA]UXSN]$7"&KNXH0RK #)9-VZ:'C9(/EHS<(4#$HIYQXO9';,]PJ\X
PGTM/8<%K@QEW*!&+QE-Q 8#N*?ZQO#'B#G>Q-'A,<6)1]56KI4.^=^++SOUTO=>5
P;SADZD]I^OU[:B.K'1Q?5BPG_8'NAA5\ME!?_*2DE7;[_'_=&O(P0(C@\GBEF;(*
PFTRQ[.OO?^"/_YW'KBP=@-_'O#G_.GUDIMW\^.101;]HESFU_W%G  =GXXK ;B%V
P]< :XCA?#)TL3@Y72BFY=!G.G2$+U5K@1#;!!\7F477I]T\=QDG)H;0S6$ OL;5T
PVP<S#QS<P6@/(ZF#N",7$F_VE].?;"?>-XUV 8OENDH18W_9M"'G528W+OR"IH]*
P/9[[MY*<SY$%08\W5U.TGHE:.;K+!"Y8CU'*HKLJ)TDIK1[(GA/:@KBH,\UPW\:S
P(D!AY47=SW[=G-](.3BH^S8IY#VX1PX!?PP3Y%.UKF:]DN3X7@)ZO%+[PHMNU-B5
P <4/T1W64]*7-/)QA03$M\^>X!V?Y4C6#D^C;C/)NB[X0GTM386\V4E"@-=63@@S
P4:U)B?5^,4^@;N$0_6&V&'4\1#:YGNF)C(8G?W)$FB^$WMO;[DIJ9N+(X6*13T2#
P.$KBFV LQY49?D'H,'<TR\721D=X"/3 V(XW+9%9><@:+= \O3=<<N@WF6DZ7\H^
P:$!^ PZ)!B^KT9#<P?3<9%QMX3T=;E(ZROU)ZB7"N4$0$?J[ [LR6TW@-=:AMP]V
P(0JD+8PHS\;5:]9*(SY8 YKDD)=K&B]BP<>>4S0ODYI_=X-WH:+;>% 7*8UGTGN@
P/!9LD)&A;'CW]0,M K'R7/EWUE<P:._]Z2J,M)SIRRI!K5.5D"J43BIXSIT3KEC%
PX22M*T?;8Z^[7M;B(<>3%3A'4KFE3/0HP '*7!ER'?]:TZ<#?]SO'V#YC\?LM8BT
P@YL<7? KW42"E.E53<JT6*B*;(E[RVH"P!*_M\(J_)(<>?&LYJ0'0_R)L#\"G;7D
PP#Y\Y+? J<$B[21)5X^.S/-.?6B*:++QGESE-W>%<88N%)*1U ,9B<K%)8P/Y$&?
P5)[W_1]8@/S<.27U:)GVG]MSKU).*>SF$^[TT:V]K%4R;DQ-]=X$I@KM]5VK];50
PAU[*_1 (!(6>M7C.0,!OQ.L1#.J01%,M,(^BIR6C.$>[/*3BGOUUSJ)_W0<B]1L8
P]6*<34Z(:1KDT1ZF,NNJAV4Y8A_(KHG75-!;!H5=U_BOB$S_FFX5L=>X3%_, YR#
P%%&TRF/.%[UR Z:CHN[7WYWBXYTI"7N& @[%Q,$%"2>R[D0,ZX/S3R?%_%</S[5"
P<,CTOFS]I2R+9P_#0'MQ6XI8)72$ZY)H("0FMZG(E6E.#=QMI.AHM+\"C1OXB^?L
P"F_N2H'QI*%93'U7'WH[(KS>EZ"6P .( W@V+L Y>#&,C(S<8%(P8S?H@2T[#[R^
PS&!0JSP2ZF3Q![1!8?Z(G[3CT!^0WN@GY.G,/[<*0S!@7J])// \-%#R'NC:NZVX
P +7!VE_Y/-A,@&CU".0"Y6NB\@AGI%OWK0L6&6N65&XD.WB'<]76Z\06UHA6-$YF
P_T+7]/<-%ABEYD]?II,K4JZ4O(8KDDA=] \64!L(&WBP>_GGB/[Y2Y!D,;";66^+
P3NVM)EE2NE </C4IP%*8L[J@6PA7H)*QDC94RE&'>T":;\W/F[^NCK*C]D9H ;@W
P*[L19M1NW6I="C7K%!L?X$#]J396^\+0N&Z4>2._)O_DL8JSXK=BMK"VGK*Q^6SV
P/NJ& %+P >C'37,GD]%Z!%OP0,[O98> D!47+$QD'KN@S&Q"XN;.]V/KC\0OS1Z#
P?S[*5[XGDNJSTN,T:#"T "E*V0T#PF\5@YB(R4L_SS4B13-:W1=S]BK$HH1OC$--
P+XN>FMX$DW[26=&AK&% 15DY#[#T0D))I-TA(V>$/A57R!1V7'WSRW\3<,M\++@V
P&D(4/Q7_6Y3)P*-GP#X@!5#D B%:[->@K/[PQA[?9E<,7T$3K6S6*Y Z?BO:MN\(
P=>@PDL)G?J8Z%T\S?&I*8O-Y/_.HE<7'\DZ\0WKUC3D]ZV@+T/98="Z+A^85+';:
PR,V4MK9H0)8WZ=N5=?:L]"YB'*H"3?J6Y^)VM*$M'6\[YS6 O9D;5GN@A9\@_Q^K
P+3'>F[']J<!//<T'M01YS)O<XK;]\I-():Z,I%PK=KL9>L:)'C[HZ37"L>7^*'2H
P8_4?_YD1(0DQR*F=Y6WUM\75(,]T^J&"]&\<O<Z4?-XSN]5J;2UK-D,N3_Q"WR \
PMGDU@V\C?U* X VITMAS?IL+8QC5^HR5'\.\.])9OO7Q'5O,N'1:7BD'(XH"2<)C
P0 L.X]8:$89LHKI=2-K6V?N@IDU(6LQABO;H36T)P^T*69'YF4QXO1G5M7(!W@B+
PCP9Z4^B!"4_@.X#GGN/9WE[-RK.W$OP"*')B.?1ET^YSTW!\GBO-C4HK.AA&$FS8
P?X0L+J6[Z!]X^A6)[Y"5-O GB78H=Y^CHG !GUOCQ!F@!\C74MZWCC#O$#QF_0#1
P^U'53.Z%,7SMW8GK:9]HPU>/RDM+!BYU9/)_1XQ%$I4'C6):9DSQ\'_=_. #C2X+
PN5L'R']5S/89LYV$0UWR#9_FN/F'!*YJSDB-DLWM; =RB([^(@4!G7'.5?'P,R>9
P.&@+C5SRQ$"E#@(\VN2(_D<HC:,F-ZNC1^:U-W\&3(E<6;<',AY_DE'=:B2*/*NG
P0(\<J[I/.KEOS9RX<>N2L="-MOM)%>CW=V/]C WY]BQGKE!N[#Z*<_O[P>S&-*55
P#XR2#THFEQ,;<_DC?9?+0:30Q:@1T$WJ-K?N>G(RAC+(_S(A[IIQY&6U)/.Y;^U3
P,UBJ5VL KBJC6EKSJ]/ !MAD1-8R <)0];6M.DK>%UB+DL!Q%Y=K7!HWGC?@O\1D
P#82*']C+CJMONLM9=/R_-W1#B7QD,<%R/5Z1??QI8#PB)/^4*:XX55C\"UOMK47?
P/X[8)"CZ_$=%&^!UE0R_G#/92*T,P*_Z-;%PS&'N>*O_X<J!R&#ZI</FWS%S_7&3
PA(/W@M34Z%<&O1WKX:*73U84_QS EQ.;7G68BKN\=N)CBI0<&_V%!NR$M.M^,<Y^
P1+01?'$$FI-5,0OL5A^WBKNK;_D_<T4:T*:Z/57J?F"'VD8-F&$,1,S+V.O*M@/,
P!+KRFC#/7P/'%Q_=)S%7=9Q \$)]L#UTYGJ9N JA*RD&GV-YSQ%;TJ6K$:+M!_/T
P W-QC&6=M,HFK5!'P3&JW)F94Y-;,0L2-T"N@?8[2,?3[&YOBF>=''?0JDR6O!QI
P@B3WPH=I>PUYM%6*%R>4,(I=9Z&SOZE.I/3H0'+SO@J+*6Q@X&[ R]&5?'L"2I+W
PW'@J1"D2B;@7&KWW&:\2_6$L:%B47)'PS)JG" 8!$H9G&W/FR-793\T1UL^D$Q]^
PLWI%:9LN9=<AX3,[OS\S==\N&UYN3RS.(:5Q>&(4WB7&1 3>+MJ(&#QI\3S[_Q]%
PL@'.@F8VJ"D)WKGGGA<<AM#)N7H'IB*2/_VEZI6&\:?UQ !]J7KZMFP''&[LNGBW
PJO?EX:;6$=9MBDFRAEP9&[:G1NXER7T!C8 2DO540\;-!P)BT.J/1W;SW=,#9R%>
PYG;:<83FR<'$FQ:27\>7CC==72G0DZT+'QY!1B])>T14QI2.0ARE0=ML RJR6G']
P]7S_%>$Q<*,Q M&EH+"CM="F,"U/;.'(L<//E?N(?(^_0H\Y^PN $"+%=0"YVFN9
PT*Z/QU77ZJ?P=<EL 9KV0P'0_C4NI^E!9XY'>N1F8UY%5P)I-5_(YX+:9E8J283:
P*7ZO0 [%B;/B>@T#9D]43/=-EEM<E(MWW6:,%6I,\!$BZ'56"_;GYKKG<XIZ9*!A
PU?EF;XI:&"2X+_"K(;:A&L^D.E:V?WX$Q%0:X*>B]KKYH9?/3D^5W2>/NGB@29ZC
PT_'0"^G.CT("L'-E7+KON2,ZE@E"$#;D@(>JSR-/#W+,)%JW<#EV1'M5Q>FVK2(?
P9Z0SCJF+^S"'&PS&8:^/H7.RB"K%YI9O]HB9G&.!VX%+!=]2*G[Z:SRXF;#S<E:@
P288M3[?&Q$1OJS 8V6N71Y2S+YXRP3+-[1O7)H*=HD%=&7.[?.;S\\XQ7R5<Q3Y]
P'#4U1;2T[C[RPG0) LU.,"[J9SHE#Z][WG.6A%W&.9"PM>?&I[AH6*YEUH-@]Q9'
PZ?#F[@95#_\'<1Q>35G;9T<)HWIL.$:6N,PQN3^,5IL5467R/KA7_S8-.V B,EC5
PQ>X001>%%8EZ5S(>;/>1?GT^/#Z9#GVOT^T0GSKM+0VQW'#:;?(#T-_ C^4'#^HP
PVXLC#FO>)[VO/CH^B09G,J#QY^2<(2GA3>DT3WF=_FZUQ0+$YU_*[%O'UQ=M SB<
P0L2\( *T=^7[/DMP3L62['Q8*Z*\:0SM/TC%@OK+I>U*FE4$)'L7-V5>D-!95#.X
PKNDN(=,8.2G>JG@&LY# _'CI^6S>;L2&X\S][4IMVJ$/ X%VPY"2LKL?,/=+9K',
P;;6G!V2J2!-C1:+-(OIMG(IO8!,7U\J>M9GB)6<WE,<4&U84?9FT6W?.2P#M:\;N
P]!JT*WG!/ZOQU&]AW@U9IK>*A=G!9]C*C/!HW; &>"D<(W-S6^0#@'KO8%*4 ]+$
P8OEC3'*_IN#&)< HV9Y!!WYBRX]=_"F:3Z=:#9O,*IA,:5YP8%0Z))[;"_'Z.34.
P1ES=?,E\R^X*H7'Y*,_"=1)G(G$<UJMK6%2&!F3"FE!V/9SR(?KXLE3!J*8#"+AP
PR+8X-&<,'&+ 0@[0HPN9L@\0O6).2&>%\CF986=F'GM UC=/'T88.'N<=$15")*7
P%QAO6 @O$V[++ P0#?CB B/A]3#Y F7,N5R70^B^Y2&J]\_ ?ORS>$1[T";Q#@T<
P"-;&QYSSFIX[7V<V/@)9Y@4GER[75Q%%)& >R@FPQJJG;$^O))4="C8W&!29\&M*
PRAP4^DY6@6R!7$O4;30LB'/W9@U"=5I@$0,THB @Z?60N<:.W-3&)"R!E>]UD+X]
PHP\DVRNH!RXV_9<:*J'SHH3 >DT64ITMIMRU\.4R;'T&:_'.I$:Z2M?P2?_*)(O;
P#_">'BQRP2U5?6&_20@N"?U5BC>/B:$HW;$RMFL$J:34C$#@7PS.Y+%K.<PA@LG$
P1C"=(>4#PJ@QJX@"QD7C]=/RG.P%S6G#^[M\/_"Q7MP*T!K<<-,=?:G]=;!MC!G/
PGXH2@._8'N^9^\52]A7-I(4X5CAHFGZ8DG.4 8U7$%UAI!2VV M0E"A&X:>*Y6)T
P9>W+(5DAMOW!RI&5U>1NCPF(X#A7&3L!!GPD/9#2ZF)4AA$&)G/TQT/G/=.R5L_J
PWE=R>7O!+1S6A%94K'JK'U;K5M*5[-&XFS[K7N&IGZ:*<QT+-TG"ER(,6:7-4@8$
P\<LM\39D77Z8.5L_H:^KS=\BGK?517_!A07 & _"C$"<%U_$IP3QM8>?Z'B'W+4P
P\'CU3\#+>"8DA,3_)(766&\]]"TXVL"O:GQ0-RO$:CTQ!UD":TGUI]-]]9IVXU2M
P!-24PCH0%VST1ACIF6/S(EA$BJXF^@35*HL.F6V;)LQ23>NO9L2#%]O#'=CBXLI9
P3_3X_?",5]:Q3.5B&DEY!:?D5=0%8B\/@'AK!=@&<^L*:WTD>292?MJ<E/ZMM#@D
P,WXIZT"JVFF** H[OWN*T@90TSP;-S6U,7Q(]UA9+5<LJ@)YI5K_5.C5*Q5R>/?]
PO(%L_KSN<&,761\<CFU28PU 7&?NUX,B.E\,BOW;A6O4<HGVX*#/7^VWL[P4H?BO
PD:!IG]S<3'/8:]]OZ5A\R4#>,@4<J A;7)-N2Z-]^5U7;8V2&]Z115ZSYT[4"*LW
POP<>AAA-'K,A==Y)!GW"P _EP:2L)8L3:@.QFQ^GYC$A]H/AK1H0#7?.^%\*LT;)
P)0P8DH/FNW^A,5UF#'*OTX](H?YA./JNM=Z:9T3Q@@2*1?)ADJ<>L1+AO=U!E/$\
P*7@],VH-@V1I)%Z/"N9XAWRRSG8$-.BQ16SX\C31YH33 J263"D5MUQ"^#64)]()
PK4&5STDK5?0PIDFDJ5*\B,\;OW&JF_H"V542ZLJ[9O!MDV/K^R@QUE@-0\A8XB"$
P"4BQ\4LG%KD8JD-WE!/5U$>'%>M1^VDU +IH0,JQW"D (M@>FFU';Q!7]SV&/L>8
PT$)0R?_R22;^=+^9A=ZGR!!3Y$M8U-*66S@4BR5^BO]HR3(R+'QAW8;?D0X/U(LG
PR]12+Z!&J+R_G%K6C)?WR=IQ'%7S0MRT^7:N8.K<4U6W/VZKA V46%9?6<U,73D%
PLM>L):]4I)!3/OR<,4C,X0 OWW2EXC.@]N[]9ZZ5IZY%H,"2=4;'T@OFUW9VV%O4
P)&U;Y=/*DGN#_3=ASO0)5:Z3DL)"WM#M' R"G8;WC'/$5F"91J-0V&F!YP4C68Z+
P/W$ZG:@3Z@UX#%F?>K+CAP"D4TE-7[&CC/C*LZLPA-CSI$:9U>$_7<!J^6G[D>RA
P?XOTN8W,)!9+CWZS<$==M%I<L.+L[++M!ST=88=LH514]?Y>TKHO.(]O9/XDHCOO
P[(3]V4*TJD_D]7H>0?L3^LE^$M[H#PH60OI"R,QA\'_V'!GO:",9Y'-R]1KZ'CY&
P!1!LL-0 U)D&M" +;8_F9_)UF]D_8!;-';$,$AVNX3P'%^NYNWU6/UH.\R/SUN9,
PZ4FT!Y(@V$=:Z)%:5]L[4_/ F>>YI:8O-NSA?0BRT3R$[5'Y1T=%%.TF6EHYC6IB
PH$,"3>V5WJ2GW]-38_!Q1S)O4-N6!580DNG/:>[_S$"/DX](!L2J@03"KXZL4$%R
P=Y/)RHY@CXB,O.$(5M3M/5EJO^<<<6838/F<R>%U3T"% %B5P7UVM< 5"2E"2B_U
P\VS@\^(8H?-4/?FKC9'P^NL.##.E^2:*+5'+7BR9PW7)S"R/T)1P05:-;6IJ!7''
P"2@X&;G^[B].JQ (@K="E,C]0]JO?M,J''L\@16C8#*;TB!P5>"A"QU'1&NRC1)3
PM,K0_V9BJ(I;"8\V14VT*61V\I'M:C)(#E36UH,%0?'L/41VK3CY)O53:]YD$M6H
PL/-(YJGX&&5G,$3DYK[90&28Z+9^L!^9_L!=?M >)!C_:B+Y)XAJHSR25&!SY)4H
P5:6.OQ^.K=X%PAJRYA;YA;.HK48/?EE8>>1G\ L_@$6LSVD]R+3B,@G%)8T;=Y+&
P<*7ZC+\ 23VB,50M$E1Q UN%F&-LNJ'ELI_\G)76),@?]+5J5.,*#\N( @(HXRWQ
PIT][BINKC0M<X%&F;XK.,ULA^5,5C!5>\Y1 H@259/)'54!'.WE)+#E0\OM5A#_(
P6_ D+'Q%!M<G5/M:"%Y+=A(B[E(&>X@9PD3\(\H_3>VE&ST746$P-])@F913C],4
P4%?$F%(Z#\3"N6D3R'K*R 7;X+0-K?<+':W),".-^]BG;T1FS/RG-LJM(I?]&_I0
PV*OZW#!]'$9DUW;Q9%F80BN#VHTL>+/D\A\3%T5T 7WHRW^R*&80?$6V]R?]75*4
PX?QF%L5PEX$MZY;P^V05"QE98EIQR"13U?@+)=;=DL5G\.O=%/MO>SFNM^C#.78C
P2E"!5_.:_HK!G7LU&<D1$#APS*^#U+2T>%0;)-)EOQEZ+Q)E.@)C;#THGFTS)\\\
PWL4H X5?X]'HC+T5M11,R+5L<>Z'WQA0@FL:+L$. "9C/_[_81W+<KM<'[F%3'&[
P&[KM(<9_&2O?H5]A:RY^1;U93>+DKJO)9_(0X+^_2#%C7$$Y <[$'. O&$YL[@?)
P'11V?$ABY X26M2F$^4 +N7\#'E* T",#<KA!7?_%+\]4U>#&97%H&*J D^P\8R 
P!1V[1!W43S93(/ID<-D_AHHX*XH]0A'D0MFD&'WGI@QJ6UG+6L45;IRV.U7UZ9JM
P_>F>Q&@ O[IUEK-^_/%"O"P:=7Q:(8I"NX*?!.7A_<(K\GQ!('[;Z8@YH(5VMQMZ
P]K^<[^;//U00( LW^D'?12'82$2TL#L++22;G"LE1@: *@\]%OT N!]=T&84@[,K
PJ'.U;Q4 06J*'_R4"AV=]AQ:SOT&BOKW-A*?X/XX]J9EQUQ$,TS[0L'$$##"R1A=
P$5* :;&^$)[7,L@;]OGL7^I^Z(4 7(%B 25(0:*RB>!>T[N]M%(\77N?KUBLOW'&
PQ/6OZ*5B=,_'*E&@D=M2$)TW ^-K:7U;86L"0L@*3TK>%:?_=%IHF'? :"^.WA9I
PU2M6JC=,RU*1& +#FWR[OK+<?6M55#?Y-(:LW:1V8KAD^7XU)I#= 7$#/=*?JX/9
PO]Z1Z0B7/W^F>DF78N;(@_?)8CV!32#+().&I]X=>>2I*>094.O\%FC;(2*S0QZ,
P3M!;W$*4"Z)0V&JR\3ZZ*DX2@^;[C/BU;'%T!_QD )CG#>-H^[GX^D3^>F @?B&X
P0F3W@NCO#_S4FTK= _1J+3!5T)+ Z[!U"DLD7M:>#@[VC*%S_6&F4.CJ&#=OEX&'
P"RN.:L KLCD9MNPSS,#+8G!DUE#(Z093D-^QZ@(T3330%<T8-B'3G5=C^?M6Y/^'
PUQ$4B1ZO9SVTX#>3*\N;'I($WK$CHP,Y.;EW==[*^RZ]*2YG$&4L>NR&&"]T">6*
PS\MP@PH<;))HB,]RD!Y7>E_4*F=NV#)JM\LJ\[>;J_1#&8%A5%Z8^I'U, 7%V8/9
P4'-68"+*E7L83:27&>R1:!BRT150,<'1W]15Z9 9SFF-&<(K' 401=Z]4J#"K#C1
PA@?E3=&^#:7?;VRK./+HK91V 9VM3S1>_FC?G+1416J;GRV(+.0C#WA6@J>/I*N:
P8]AMJ:.W*L)3J9VH(=Z2LAL#^>=K#.,BT,,E;IP:]XT[ZA1O!'I!$4^*W6*ZLB\&
P;H+?)JTW95*\0J>>JVPIV^I7'C^(XU%+CP8'-V:8LI"M?O@:-C+K3AA3OKIR9E&S
PZ[&&!]H01!*8B_-_'MAP#,K$O<%H*G'SDT7>UZ4)(:@O=UVZ\Q+L% -R1>8BI@8$
POK\8U"G'%H[6$D&C+,HPS^I7C7X,D/(6**)AR%LDFN%IU(!#)TC!'TSN#1.&#T60
P'2979Z#W.^=)ST////*4^S Q@]X,3EQ"( E0UJ=95DB6][2/%B?Y]-8RX)=!_O7&
P#>KW7M+K#T]4V!\]X):&%Z\\,"\A ?<I)@-%Z,C(<LFK81XC;@Y?NOZ;*P3(]LTX
PN=7WFE'Q97B3L[NC'7\57250P#:DVN,"UUUYO\$:]%=E6@-WMM[D:9W2J 6U:_T+
P*W"AQ'-E=(SCVSL,4)<0&8HIT\99](P$>><%=+B'A.1RAK@1J*9A/*/L(R__&CM"
PT5^0IA(,<%EUT$M:D=PLMY#88JP;$GZJBIVWZ' AQW(8TSY!F_)U3MAZ?LG_P>E(
PQ0?5GJU"BQ]GH]/:BB.%9VQ]LDC1]'E4$W,U]]>3W%X>:/H01;&&O!)W'5Y&VR;9
PQ+9:2WH/I=9\>!,MF$<0'8J1$V0TYD5\"FTNG$^0ZR! ^A:4J)FG-FE0(E [<9W0
P0N07CQ[0&1##+I!OU67;M^, D*#_@4)G6AO)[NE' 3Q3W59>Z<6A^*V.DNNO1R!4
PPVB/-<RO,O42%QP>NO)7:M)Q^F*Z1@/-PBDQ<3PEI8&L*ZE<CD49J8H!S^Z] J,^
P'K1J30 "@/:_,XQHQ%PDS'G,A(HL:OM'AO6#3P<=:H:J16VYLC29SP5X6%@FC_E.
P$I(LRA>6O-<)Q*\;>3+3D)>X&<;U&DZ98+@Q*<YO\G &)D926401;</RRPB0CYRM
P]ODGE[X;]AHQX9-#V8!(WIP*Y_>VOWJ /STW[AH).&UVQD0PK!K)D-<*+;LI0\[E
P<[!0WY/3$U1JM[D(@*UQ&B>RC579Z=K5B07&-Q1R::*QD2V\L%NDU)*^@L@8L1S0
P)>1ZU]%J\,-)X:"MG\5X3!7'76:I/ZON=[.NKE!OX#>&W/QQJ/ZWKT?#2ITRNA9S
PACM8F+[R[7SK,)@UWVU,Y>H ITQ "0N<=@,,JS:%"Z!0>I)4V$1^K#[0@EY"(BH\
PLU4L>_IVBF[P#WXN@87XN@#OM:^^3?5ST[4NS%J/[=G"UQK7+2-;J."M'[] (VYX
P"P(8RQ@AI]<<0.+=!NRW5?.A-L^@7LN$VZ?9@+N@ZVB'$*S%:#%9DSJU C,$<1/_
PN-FK=U^I;S,/-OU"^^F/Y-1P3-VV_\"<()LO(.8&07(-TR?-&*9QKV(-K\L$(/#W
P=V*RRV??M/_>W!VDVO@A#;9X"R1*!#_ LK\/ET/WU./!3ITZ.8_%>9CQ@>*%GI I
PX/;D<&NV?$3>GLL>^+")>M$[N;B)F@OB_;M.*WF^+;LC8&1^60*NNZ:QMAY@^$$V
P.W>YK%L4@,UGP8R]_(#U=-[WZOKHN< 9>]H2DD+4GJ%WYFEX$<_>\";N.8K3]E =
PW)1GYX1*$Z57(II=K$"6<U(;T@NYC0H_4@0.[!EONA$KQ.8RB& JO#C_0:<$P^90
P*"9KR7J_V47D)K\_.Q[/AX ")%+&<89&&KW"5RHSI_KT=_E**#[M/NSD?/6JB>U1
P1>/JH/7ROLXFU+=31! ,@O>M>3R;P?"HSRYL6%$P8ZU/I+&BO$W_^#[0PY@9W)H#
P15+S<9/O/FC%8XQX>I"#[U&J7Q7.D5HB4XW!06>BN:Q;B/=<R#W4[!UL[\2//2GL
P8)EEJO^?EEOH _;TN$H864?1YE*@/,'FX*NS[]V!=&X)%>GV;HYPB^Z$0*T_"2";
PF[@MHQAVL^C?WWEC%[L/L29M2J;UW79('XR2M*C 'H30UTSC_R9IQ/:*!Y[KQ]Z*
PP>@W.N#RP;B.SU]QL+Z/OS!V?;%N;:DT7S!#'.CF>\_Z#JBHE<RAH#.P0IPF/2O^
PW" J3\CV?D;2&*OD63$_G+6^:J?&D)2DGH=I-9R<2AZO6PT 5.]0=N6 ^::L49CS
PK*ORVW-^9S\1&@RBR+?'0<UR8*Z9*F(=[5^*;/X$_H-%W[#BZ 2"JY<27UZSEI%B
P%[SR[CFKH.%G83Q#"NK8/F)I#S_N0**>E)F.0W(M!J?HG<?D"V-?=U"A1\*E!3WF
PJF H&NFOJN06I:T73S4'R7%+#-.OM,%R6"#@B<!,Y&YV#2##%X+IG;C:E\L]3?#3
P2+Q$\I)5"RY53XN@/H2]!NT%==(+/4P1?X4$P_+U4UA\XH:0]+HC*NJB_JTVX';8
P_KH=<'#)#]SI"/,DE'3;]Z.RBZ:RU.>AT4&5SL88.A834X\#EZ<J (\\C92=_5;C
PRSV:6IP,K2M>:?!M1TX^=H2@.6%1JEW6"NM/.%!UK>=XL. WGGFP@!?*O8!T$.U,
P O2HC+8E6BCHT(G/%&0E0"'6UM^:%BR:BE#"4/Q47QL;]AWRE66>CSPXKH02+01N
P;EG.CV<UP&2YEI7.-7@>L<A)(HU&I)<^2TQ>1^-1AV$(=?K%SJ7UL(77!<7A1CX$
P?:T.48U0^J*4J0GIF(JZ3B$E(;25V8\=<K'V?:Y1)H Z5:6^E35.&ML<'H'%E*H4
P/\M@P,9->,KI-EV=L+MFL3A?LQ_QBISIL>[L>H61+LZ!L4+EA0],WM.=\&*.Z3DK
P#YA2YX2,N_>4^WCBMP503N(S%L #=]8CP3Z)T3&FJA+I=9T+CORO-<A??GQ[%YW_
P/K+-'IYM.U]XK8[1,+N/:'$<@9&V,6AHV4^8,YYL&J,;*JP^@L(<7_MNVF4KK!FJ
PF#*&2!)V.0:^&:P+2(Q 1CVHH=5EE/5>85\OR$YJR>FS.:>^ &=.^Q4^:0\OND%.
P ^+PT;;?)4YM/(W^8T8<LNB^K.D$Z+0(BS;6^%E?,OT2.%TBNH?-Z6EAJ5$B-L+D
PKP%F:$M<L_90HZI4I'8UE^5;B2TBV#AKR_>BZA(&>SEX2R@R B1@:UJEF)C!Q9!_
P?A_:\83<S*&7Z=_K:J<JZN6JH\6-S?^R\'BS2UKV+1W2U&USOK]^M9?Y>)7$YUY%
P[]Z%])*#BDR.P?HFMM!K#2P'C&ZYL7@^B"Q^I!S+$ZF%'&"<@UF2% Y"L(@7P-<T
P.7RQ%>TZ4P'82-Z@C(Q' %(A @PH!("2XE.GZ Q'\-;UC9$1=S"J''>[BOB-4+SJ
P07>(6O1U _ DAWK^3T1X8XT2C9HNG<(IODZ"1':OI]@*:T6D9(6SSES/<+/8F]=\
PC+6XQVX4&+K#!+PL()4+R5H&RN<N8-N7>#7ZT^WGLR7USD5A6\#<YZN0,&'*9T)S
PO'FCD&N8E,DL,Q!0495+MJ#HF(CCJN32JN14<.LXXT?7V9< ODGT1/U8V@D'<&L:
P$A6/-D&?,FN0O?V;,VF"8]^=296]X]H#\D*FJM=:1/"XP1&"MCC0WNEF089D0K;$
P43MND7)LWV'\R-; "^^-;YKEKHH24?]W;:8"EZ?:+&FD$I ;GS"@SW=@(VI5R8"O
PX=!UHC=."IM1,FPR)4\R,4K'97M'LM%T1#2 T<W6@1Y8_!"C!K\G@OM#A2V]'C+^
P;.Y72/:+YO?W*I'V!!FW)?(#@*/.GDR-P3+\<-Y4J[(7_87$4DRO9RU@B>.>;?NN
PC"&%*$KB?EE6A$%;"W9$XEB__P(+<#')#+4%:Y^Y,S%NV06D$QRC(>IO.?TG4,M9
PF#4 7[Y@:>+5*-%!IU0BU'Z_$_F,AV]1:1O.DRQW0*F'>#^CG2 2@PO',Q'!7!\1
PR&T';5KZ@F/2QHJYX_=Q!0F]^/\7&-P1Z:?H1[QP1;? C267,\.]D=;&R6ETMY@_
P--^3O_"YQJQR<<8L;71<U=N ,9P=3Y[&R6@AH./0F8?2=E !RJOQ26V*=S[+ "*/
PQ5E6<UF45:=,R!Y'-SA]XTW7%"+>>$0B+HBW-0@=9YS9#BY2Z74>VGLR7)._GK?O
P;=?8^OV49[G$"2(Q_85KXZ5),!_D=FO*:RJQ(H3.6)MGYBN%-O<[CCI\^)L'(QFS
PWQ".+5B51S:ZJ(\5?0X_"JNMK1?ZF5V_0^#HACYF^,V9,8>_E.U?,^U*<DX)@FPP
PD>/[!"U\@IP_PB(T3C<^\%VSERJ#O*U8HK]R@UG;.5B#Y4!:_-CBY\DZ3@) (C_8
P3R6RWUBJP&:$]^#D/B4MB%I-/@P 'B>.Z=)X*(A&<M&%^\_$</)1[P]SJ"OYQQUV
P64L.GA*M.JI:A:F!HM[51+%LV[Z\$%)9[4&"IZ\SG0CTH0GA\5CQ?+*]G'3^WZ53
PY *WFAE1&$"]LG2 C(J*',-T/2]1.,3XNIZZD](L@7% @<5P^[S(>XAXCAW=K(49
PK33;7E#I!LF05WN/" ^:WMJ$=:L[577R$HSHH8QD)\@W#]IUKTCW[HF16@?/&P3L
P<%=+CPW)1+[S/>8"@&D<!VB9:95Z.6RF54',.1'[$5@A^:FQL)ZKX]V2Z40J(OLX
P(I58\M4AD:EUX":K+Q^\A+>^:=5<]7A[?Z2/G^VGI&1/FE"!B3"N)):"#,)S25KB
P8B?K]M*#_RK203AX@18NJNEY&$'5[7ZL9 9%S7/NOJP:T?LW:[W:Z.(#/<IR.Y+C
PB;;'>W X>:#ZX@SRNIXBR&H:9CF#=J+0\07O(G?K$K;(JC\?FQFTCUQ^C-8P>J%%
P!;T29,>\]*?)0PE39\.'/J._DVV7TP%KMIU$_UZ25,5)1LXZBIQHO<>E6L!V8M]&
PWTZF4JI_@%!]9#4!1'.JO$8_.O@OCWBT.SM#$9"LDJ8;$L],<$:QKQ*;S?[!,)HV
P1^[2F @DGK"*%LK/ *WQE$5:BY (H2JM':WO0J&6D+YK]8DW?F(;Y\\^%,*KW7M?
P#;S4-"!SYDL[RHO\+:QUR>MQH ;X2&_^D='3MSG"H$@J2*<!;6Q)X_W#<0\;BM(B
P:\GY1?_+@QZ0?.W1%Q!V<_]GE6YFQO^]@2-A^2;J?H$[O0\LMW:R7:WC$[P_D5]M
PNI1U;N$WR!V/@&LI]S23_X9N*NT!Z1_/E' Y,/Q(Y#M"0PUH_Y\281'\I;92]:IY
P"I.^EE"<3 R@57B?_="))4*?L=UE9C1"HC?IZ07[:L= Y:-[3$5N80H%U;R*:3-G
P4ASLB(#7>P"RQ#ZE+X&H#14SG@&"(S><Z,KSA+0WD5K,"H38Y*"D'/_8'2"H8%)K
P1%A=Y-#J[YIQIR$'6;RZFJ^7<L;[M]&)U;T(G(\S5D]BXLGF'W!9M:J)WB%C#4];
PFK__UI@AMK,'JLC\BI(Y'>E[7@[ 2>#:$1  &$VR(3?Z44PI>YM%J&2PI3W<6BN!
PUGJBW7T8J4GZ-1LD;:^QF_RN)Z-I+$Y.KVHL[B\AF!.Y1FYW<WY)\IDA_C6HXB>+
P,L1E:5JLD\?I4O1*!);]1PKCLY8XW<GW0Y+16NGCY[ )8_Y^JF<0.953*^1LF:&E
P)@ZC4DNT!"V"_#YS#XI#8==8H:^&$?*2G>L:G@GBW4AR[>& J)7(%SPR"[EHQ2NW
P1:K=< @LAP2VCT%U#M4=8XKQ<%] >$_%9VQ4QL@9/<U<3N3(]$!Q$36Z[B:\')9Y
P;EAFC?,:;^? .KQ'W) 7=N&3X[==_UCL<4IZRC,7W]AM(,BF,UM22_H[8Z_M0"B!
PQL8TSOGYJWH!:?8L'3_#P60=?% \TYNRG99ZN!^ $J:W\!\MAP@R;5^M(*+;F$I0
P5R:AY@+LX=2<&(_DF'E3[!\RY7#'*KFDRH+;E*)\!5+,R(I\NWU*"5M;ZC3> \DW
P\/'NZ-!GW[LPD/PP)N/81($6&J/R'/086H_'6;X]52C1DMPM9K *2ABO&PAH8!\N
P>I6!,XV,-58882\$OE !/ &^?*,J7O+F&7E)9(+?\@TWHTOV*5UIJ7S[1CRKPG(*
PL-'&]&=URM&,6)9N6UL0#\,[.$;#[KZKA2?A-?\ L2RGHF^ELVM@'T(W^,7;< Z'
PTXTJV>8<EZ9C'INZ0E=/A]1@LSCA]9KJGVJV-]J VTWE+S8('Q8$LOR-WG8VTA)0
P3/!E,V)(5ICVV<K=>8B'-++@ZGTH94._DTU3)T]^:]O>%0R9/NPR!/KS;O;>+,S$
PA96C1=!0Q#6L^E-%YFAFM'KSAEXD3R>YP"N+(X3)B$8*$=?SE]#\D!AE)2. 9=Y2
P^^<+7E-*(N!$#HK8M7HB4[^0H"Q&P[$;P5YJ6G:_!55LQBC,<V'?_\9H;T+W*_@E
P2_2^!)L4<W@?T1O.B&FARD F:3/T9N_STDGQM.I;+ >0<+(?G?@IZ/-&;1R+%0'E
P'M&OIK.KA]/O6:8V3+WH 0^W1.,@5\U(@Y'K<7K<N)=VKQFY>IY0/2V#-DE4HK78
PF!3Z_<)S.A&>E22%62;NTAZ;E:8M%X(K;+OZ,]#9+]&: 75,<HI6/!' QBO4X:GU
PMRCQ"<D&A=DO*?H8BO0<PZI$YF00+N[>"G$XY?!Y^8'\5=TM"8$,FA6&;P$MN ?]
P6)(A9)*AO#]\PXK9JC)N02 K7<H>0TBX5^@GH7YBT]ABY-^_K<//F%@Z&E31Q>XD
P$C%,+=D^RJ41+Y%*U@00]?VKE::O/ATUC7*BRA\QKY+7V/EGB7>ZJ.8ZPGU,6 .R
P#0,^KMX([-\8/ T/5DGRM5\H[,TX:?=K<9$(B#255 VR'+3\]_;P)/@#EY/_Z76@
PZ$=%(!3@+EIT[4Q,W(?U?:H>;JIOETEGP-KKS(.@?;&]9$$/8E*:FGZ4%N4V/([O
P?X;_0N@]#^2\PH:ZD1U'GLCA _;<6&.U6,42N="<<"+.Y"9EBKJ->W(MF$,-,GI^
PXZYQ=47_6%;<YM>*+<]I! BWY_.7CN@N8K= %8NR#QA."%^YO,V_W]#7O$RR6(+A
P]/$2?UR=#=M<3&\W2HW:EV+_][/"1%5#"H>^M1*E8J9R:80$->;1'&Y]3>1H]2'%
PV,&"4VQDUSKS[#[UF]AU_5&NGL?EWA<P:YN0$ QV<U#PR6>XJ:P5?HVE=C_I1Z!T
P,='9FP]E-1*"[*D+OZW*3MO[TZ.:!L2*T$:,.&!KL,_VVF"V$PQ4<\W:H"6:#A@5
PL//9";>MA*VX9DN/I@H7@A0 E4V)CD4 #;Q)P:^CCPM!HSKS*U;Y.Q=@9Q:W:X_A
P/&L>,M_+0"KSK2DGCS2+[XSH*1QNPD79._)[]LZ5!J;NELR72DP>FK\,XG 8J?8A
PI >(*D(L2D*U.B0B%5.[P=!^QI<0.AZ ]T!P(+''#'/QV3_'1?F3$O 2%_89DI<$
PFUTFTM5A!->J,=BU37<@:+N[%IICSC 1LC>8&^.L"H^K!HB,+C<DBCD6_282XK<Y
P QCXO[Q)+]V701+M7)#J[W]W]9$&CW.YK(7X5F;=\-WM5U^\;9DJ8 >$O;';Y5'[
PXQO$R9DZZ_D8J_E4WKI$6&B-1;"6'O6_.]"N"]XO^_=]1D2F2\J<=TYOT89.L#G*
P@7'^\_&FM'C<AF9=$#2*;J5;ZL5EQZ9\'XQX'.-MY04_4"967E>XV3*'L5/$E+J[
P2?O A,.G'X;.1U$^7$E^A[9,II_PPHMQ&CTY"N@PM2C36?A/Y/:2S^-F 1\P9%U5
P[RE3Q!HO,R!=4ULHJ3U:?/#A'('E8=LB/4/9=C;UMWVAM8B"8/7V+O+>:7,-MJ:E
P*[!#RGW1%0&,*7:@?$EO]Y7PY)0P&!@MHV*9PIK<,!LAM'7>P3QW=$5ORR2+YB&T
P;]D1+]YAXQ))8O9O97 ]WCRF;W_18S^XG3%-R&,8.KRN[;P^V$I:;A5UJV?9%J=+
P,D>TWC;6%*8N2P26Y!/.K@(R-+AR1>VZ,0U9X+""<F*K F3#N6-QCE*61H'9X-^<
PPN!Q?%(M:X?Z48.<M&IZ;(4[;VW^EKN WJ(M^F7:#  A7>=)[C<X3DCUV&A^+?8N
P&9>(>3L<]W%]5=XYGUK]^+[&MWN-K2  7^2_H(#1.K;M[+]FS%4%)#20!D*AWT@J
P'&@>-:$KT-\+ AF65D\=C0:ZJ-O:R'IDUW;^,C"OE=+L$XAV3I:AX$KO:#2^=96F
PI" !(S,;^^5FI(0K+LPY;CY^&/9@HXQA)^@'C;]QOKRU9*(2CI'J[0FR7)C)ME9'
PF8>I J?-MO:55OK_R1[45RDGG'!(0_NEW<K*C;\2<!:*'?(3.ZFC(IRIC8YZP[H$
P(3@CI^+%Z&#PX1G%L@- MBF6;I&+&&Q[$X*_^<!DF44US8_OJ4WNGO<_Q'"?#0KL
P< <[R]VY0ZA*+BX*39#X-I4"OA##CYGFT>O[],PJ/GJRT&!A<*6J6N6FJT2T246U
PZRP=0DJQOQQ"\+(;.W1>!0;*F'<+)J3?%'@Y[\N6MI8KVFM;U>7 T%3PR56A;_<@
PCJ$7P$.06I=/(97+*OB)-^X/:H#'50_"*(^OY!3B:H+$H=5W/K83B<)3U24!/U -
P][A)#W#-2MT5:A7 CU=^</_O.8NQL]TASJ'0R#P!#4O=X]Y#?S2&>VXIAKK SFZ(
PSU1(/5A*!6=?W!HIMKZJ;\0(/6*(4-<%*39\=J+GJ>$[A^W 43/>G9#U9XZ @ZJV
P"KQ^IVF@P$0D$.Q0+@OT?!HC2A\<] ?H>@+!&<UK*$S=7M[&IG>$2:%$B5;H0 ]-
PS/TGS_PG[?R?TZ>OX.<?3&[XAJF[]^>B3ZN^HP%!IN\4W8<)F.5@UZ96'\>XH>5E
P%B;77BWGR%0IH2D7_$"T%_78U55C%QO@='OZDK&QZ6O5(OI%1NZPB3MPFRB .XU6
P/-RA1"MGAI.[,%PD^#SS-^;7N@DI673_BCGGJ*@XWZ=%L'B92VXQ3  G(QV&0V6"
PB<_X_=[O.C@0J$;>;&I!M!28KV$3B1L(U8#G9D4?EC+^+D=K._AGE^SE@)>9 @N(
P[U4E(G7$;Q;:/"[_&)6O6!Z8^#"9/F<:Y[>QC\<ZTU3I=S7ZD8)#8_<*).2(0=!D
PWT0/I%BIA8*32F37CAM.%?)PT%KN$A0H]J%=O_IV1H+0#BPP<XW%PIN<N<4-2=$K
PED#\M61QQ+U@%ZH!U->20TA@,B/IJN&7O;4@\J;$R,1;(/I#6@>H?(BAZAFXX-EI
P'Q.R6!V"_Z,01Y=MJ]BSG!<C )>&^XL=;VAT< @UKZ[L59EAL0X7(QHKF5L8F3 1
P[2NBM3W^4$Q@\8\@!?WK?8\QO-JN>1$(>JLWI9_[S1V,<RGSV3Q!(+=^C9KI :JN
PK%)8UPT&AX[2, < <K'S%J_IX@_Q9RN%).ET4C.3&;*^9$.!69GJ- (>W$Y]7&0T
P!^++R\I* 05F.8P1QYO$+"GI%MB(O*5-2"6C321BXW2%ZARSQ9D[GSY.OZ+E&&OI
PL5L0&5IVHMBL*/ED'%)=6&-%=96&ANVC*6NWSA#W^2<_\FG]7KS8QVXVB ?G"K@$
P&%YG$SK;>5@T?))9*D'\6?O5..B: #4CEJLO5O*1J4C3AJ((,WKLIW/A4E:B[3H"
P>^,Q@DE![A2;L'LK$^<QQ$GD/'<^H,%A15X3@H[TN:>:U^J6A"./AO86 EH$')H-
PR])&"0NLX!,8DN'V'"A?YA271XJ[;QZRMP>>?YD771^1+T<T.N] CC-_S<[[-8CY
P@- &SO!$':*5;=:53?E-%J C#G$/BSB'$?^2>K*%T0^83Y?71[T.T4@V".XK-SDV
PEJ_GD: K%5K=_'A%]]*X;]$A(&M^#[)Z)(Q>D\=AH$<V-1<0NC502\3 A4.4 *(X
PFII\_$+[7^'G4=8!>BZ:CPK^$4^= ZK+-$'.]DR:H"]+U,VP\*U4)Q\,[8 ;\;O*
PCE+]:_:B6GIZ*>VVT%*NW[P0C%#6M*O?3'RDE4.VDR%NUO;'UZEPEU#<K]OK7^H5
P)2F]_T8Z!_!A=:U$0@SZ5T;RY[7YVBN9@Y&Y@&&NXM+V&21O:I\&7#LKO=(^ '&G
PY.88=;8.8RW?_2X/IZ-8SSRBU?LJ&>02*JD%F'83D];C0%RLCJ/K/ZN$FHI;$ ,=
P2T1A9B2Q.(YR2$"?PQ=.L2^C%Z#%T+-BJD8E'%J<]U;%9%S@3E''!B>I.TAE6'$.
P1GJ(2AO,[CYJ]#P (NR"P#^9J<X?^C'$/9I E!C:J;/F6FJ_B@00@JS4Q@R6(1:L
P>(O[^2-92HAE"M"0#\. B)*=C3P2 D^+W))WH,V J6N,[OPU(')#)51MZR6CON!O
P*;?O8XYN.O@1%;)FX1GLFUAA]8%%QT-:/C4LT1R;+UK\">!6":$N$^'TU89Q/**1
P'%;TF;F!KOC^<R\IRF7,&SYJ6]OXT5#SP@$V=3!XC66^>!G[F!O#BAUBY'@/#VT>
P">D]*G#W5;C#J,S64%%P%Y#0$B$;(!S=:0X$WMC(SDPV>HO?N?]HG;6K<X/\M92!
PAP?XDPO A!VGD:I1750$]@I?Y012&Y_RP=I9IGF[R0-M :O'[5L@I79 E*EE*!TY
PBA>#9N]QC(=]H># JO<]$)0ML:G0:YF3YTRD5A)S(-;FN)2KS#]@Z$W2F[C!$(>D
P3RKY$40]"Q"$V9QRH_.V\L"[I/'8G%^W#2,JNE%UKVV--.-9GUI)F8$>H8>&1#"G
PI_"<+>Y,/S#%W33JC47^%<J\D?2VH3?_#* OXO8*3QS5]*.I[8O/F[=0A ;083QS
P%AOT;&^89<L,CK9FY.2\J(K+):D1X@ %2HFL,0'@0A_U :_T]'S?,-N1P-&M2U?L
P&'PLZ?X^E7'=Z%H_#YVL71*79+*G35@7QF2)]KEPL]?@5@W8><8)?9?J=U&NU:HW
P7BFIM2H7#I\C15]C'AHT>*Q<5*<YU[B!M3'/+4/QDHW8O?QQ"PL(J"4@U8=LH)Z'
PTVU:EVEOO=)ZDDB "=/ E7QG(U4PQ _>P=U:NLZY%[F5Z#Z,684B-=0UAV-=\K=J
PIA"<JKK*8CL?\BE(L! 77%;MC$@M#)0 4$WH6:6??4,')Q%U9I,G&I;F6M"E@B("
P8/!?7V](GW->QA;*);VR?J$@QAKZIO#7_#- FF#V,YR*1:O2>?WIT^M=GX V@ [<
P[GRWVIS=!,[PC0=U4CX'4+"Z0C/^QV;1_&I@XNXZ0)V59MR*^GF2>%!K3O5C@UF,
P[@ODGBZR,8LS8GN-@%M>(BDH1>FWHE#@P^8X/XU;)$+?MQOT-_$!SHB>R3=_,Y>T
PLY(5U!LDC"M]49@K'A9A94B'[W9 (P$O-WWV*]A#_HT'7ZD>8,=S<.3NL:</!S/1
PVFKP%[+WCN7)3"""1H;*$,;^L:=T[46&N)J7UDUTI.AP*=@,G3L.B>[B*%(0&+\,
P)>H-N*^8+E;^X9V/3-UC-[Y5)J\75^TDDX(ZIS8TC':<T8.XN+GQUJAB;0Q7$OM"
P3* UZ=UXL 22):V@&]\Z^T"6TC+[!M&U+@?\YX^K$%(S<#/7/$#?%DQK.ITX,[:Q
P)(3SJ1H+\(^ZY#5F&+2LJ?>V3T2.GI(O&.;1/SGI?]J4R+#;S6/N_-R/N*54I>7"
P_SQK]NE&>+?6FQ^ 2M[/'!BQV<=UTZ4!2BK3$<>]Q(D$S6,_^IK5F>1M9IN08F-P
PUM1L:Q+64DF=;P]$_YZ!:;BRW?3=JVPST"306!7S6QRD"5_529I9QU9NT.+"V(?;
PXTM. >M )R>3H3?O,YNF3NNNW#$>, _.^^[:!!A*;5;Y!H>=W>R#>@=YE+5"ST-_
P]7=66KGP'TA++6K4BJFB%:M0,*W2,$<!NK]U24^U OQ(P"_W/!@)F7?:,$29#4)U
P];,<^( 84ZYDR1$0*)@P4X'Q$*O>-W1E]I1$!X\4-(AF[X ;1Q&"]?ZU_>L#2LJ@
P[%Q1V7&3,_G]E,UUW!D@&Y3^,1)H"%+?%V:.!"V+X+_(FZXY7^/O/^4[C2C;[K_R
PGK+74G^II&X'?E4$A2=ZPNMIT:A3PP?2PGN.&FTG)[@M7710HJD[E-ES80($7#K;
P4]:?@/:=Y @'*_TZ'3Q]T+(W?=0W=5LK4-7I$TV*"?4J\7&3E?I=_NMGN/>MX>3)
P$I\C QO%;K=:E@;[NA=:0N*8B]0G<''P#F+"-;'QJ<&0C@GT=H#M&LVXFZG1!D3=
PX/.\D?']X#V !<H+U[;81^9R)BL*;O#25!]DFBT).QMO01:"S1]DK9FW964B3(J9
P;<0TH&Z='DEW!.C%(+^\:O7P*)5PZY$FJW?@KQ*7[)6]=@S)S*K$#.RG;5<)^\5>
PL^ D.WU2Z^WP]RB0[L^$5="+REPH&2EI7Z?RC=5F^\@)J-A=OG%SFUU*=+@J)#5*
PI;E44VT^5/ 6$R-881],LWBC>"$?V;@-WM%+D:'-J9?=LJV36A0:)>@?#+6=S[ )
P/9'L#F2GY=T3QZ4JM-' 5PHDT)B&9J'48R$Y2<O_(.%5#2A925+!9Y0N@1T>ZZ+I
PA5SVO+VX"8.78O 9J DH5&D9"!CG]G@#JN,PF7[  4C7<LIZ!R&J 9#YMB>AM.JI
PH(/82W8DET*2\&:T^^ &OD<G,;"[JF[:WU19.@'# F\8+&+3:P[OT6%<(I^#D3"/
P27^SBWDEP3=NY&U.?+T-[)97"]<1SC/LGQX7".NYC/H[_593[2;(!J(6$6DCE+-C
PPW2 U&4<DAIQP* R:>;=FR+'XA5:W]<UDV'I( SEB=^']=GC/5P,&&8Y#L&@L@%?
PT(1DOR58/:PD,7C.)4Z@H+\'"39KWRO6_NH[^L\_O.4/ #H1?_>EYL$W*.DDQ)$C
PCAG7ZJ.R7M%Y N:1 QNW&[X]1>+3S92T.C_Z.X:5)8RXWDI:<2IKN!K>>7F7!'CD
P^4R;CS*_1O<WU8D^O,R($*>=H)/MO0-,5H>[%QT@HK4BB.>'[(-EJM'BC'N_G<;5
PNJ-MB+5(!V(V6D^!3,,&, XQY$50>[!)M-^1M:WJ.)D 9D]_]Y<A@O_"")GAATV>
PUM%F#0[5RI6J.B&E\6#WW-A&P2>RJJCUG16>&99P4!#N Z^KX:2IF3*#OD8L#YU2
P44;R_8/?('0B,T_SP&BVLOP2^.OM09^**$W&&3K^?T6:IFE>$3RR3",$L/;9VK=U
P+.L\0P,:DS(B=NCL(MD,133!W+3O4>8HYGMQ5O'-_@,UI]TH6GP"49?"@V #LB&8
PS\P6+C)#Y#/9G_#^_<Y0 NRDDM(%U+SUK-#H$1&8,$<$U AX)]?#(\5UHM:E.UB#
P>?%,RW%:'\'QK<:VU.=>3!,%7JV,JGT\\LGTX'&=T7I?NU0<"@9(+X1_T::Y@O##
PHV["*H2MYO[WY@LMATR0M(]OI$=;S3246FQ98LC! /^7B@: G!3'& YF[Z^;F<W9
P9ML30O*>7^3E/R:Z240ZNWY(!P ;B:'!$$4\FK=1L71QL(1/($4FTS*WLB39.[IW
P@VSC'!ZD+WL92M\$^[_+CUH3%[(8G_JK8U*E9! I M58(.9H](]!4?2SJ.ZN;^N3
P.AXL,4[5O:GD_^PUN(^VO>'*JV[K3: #'RH_HZCHR+K +>G9>P8_T=^Y3N1V:"'N
P_ O]^8I7U992:&Q5IR.*EM[^_*AOEG>-PL*W 8"/BZ(Z8(\%A2T2Y* #>+*=!PM?
P&N= \X)= EL/96%/N'H@\<ZR31%R*3OO)'Y()?T,/V/WEO\K2'IE-[J!7:!FW.!)
PQ[M[R_;3#"_/,9?$P%S)5AC:75WC$[<]?8 C7LSKO2WH@U;*TZD0,032 BT$I DJ
P=:?6AY!HY !)Y]VR:W-&Z!&&I],9U\;<<;SWZQ_2B,\I(PZK"0%W#\K %!0]8Q(D
PH+4=^B#M*#E8*)-469)3;UEZ2'G (X&#_N3F=IB$8X"RSY=:CO]O5QB13"MQ'.7"
P=7W/IZHU@B XYS-/07)5CBK?UG*NY$:DG50@T\+^B9:WYYD1?CW7ZD74 6H6(]O.
P;7Y!,76*3VK:B>8]5ZX]+9/)BGHUCE)*E*I%(R;JK5ZQRKBD\TN?02OI"9K:M)4$
P2@2<]PO915M6NUP^S &/Y'J1\+V,">/G8]+YRXH !H]).!#7!<A75$@X4%QPZEE#
PSOXCT^BV]FKT&D.VB<S]+[U#R+$)*@Y7)[9'R=TO+TIQ95&@(0K!F L<,*V)G /4
PL:C'&\A> "A(\65V(2/XHLS."!PF0D5:3&LSGC#WH+*+:WXJYGL.XI00A6Y.<Y=-
PDW"=X\:IQ,$_9%9F=ZQF@^=WSP/^_403R&>2M.I D?Z?PQHI)G=W 7R&N*6:8CT3
PRU3%^-Y,EHG7OU3^K/L/'DNT(*@*$*L8M#_<N\R6NLZQY*;7LV^;X/ %3ZU^H5$D
PZ<Z_8B/$%:[FH%YY+7=1^VH[@5H?KL@;;7NH#NE;<TD 4G&/W3=#P(42*:;LT$6(
PD^+)&R>864TZN0YCP<F>S&T^U"/<UO_B[H%J%5#*?/=TB]\S @/2\I(0)2]3K]DW
PJ[R-()0ZB1:MXZ2CA0P4?(2@^/#ALF0306AY[!4,OZ'W V]JKGVRERQ1%5G#W.+-
P@*]BC9:XG,D><K\YJ @_X7GEO)SUCOOMK0(:^Y+X5174L/K/&BE]/%/+84.VXVID
P1$N%0)*A) S&3_4O^*T&U7L$XZX+QUW?4U 9-SY_=HE'7!K5558$VU=>?>F=1>?3
P9DUXH78S4]T)0^^G3\X/&^2 8U7,0[U]L'&_[DP'O2\&>CGV_8?E22F<157P.KA,
P0/VQQE^95QFI2R#L093STVD#G4)?VM\XD-N0SRJMY\N3LT&M"CX. AF,'_40X<"@
PHH>"D4U>0.5>*^=T+K[##&18!P<Z[N93D"%H(T,CFD7=?L3+01?B<NSL3&?#H-8-
P[V4A@L[4M0:M3*=<=0G8O*Q[C,$D<KI!*)5R<KBXR'^0IJ'Q6EC2=S^5@%Q;J\T\
P=.'P?":%>FR4O=?U1!\6B0OO,^N$?;-J5L(!V2$  (%82EIDOO)%Q'Y(3W=4FI)!
PN.4ZT\NW$'L?PN4AG]Q>H%J_\L96$P.DCMSK4&7S-0MC039J:^.=E=L"=7=*YG9"
P(:.?Z=P$[)*K<XI@8NR@MAZG+,PEJIB"#ICA#=SQWOC4(TEE'L2_S1C#L_,XZ0,\
PFM7^^TF*H;]_<5U/3_ SJR6JL'=R6AZSU:S:1(&^O%601[&\91W(X@%.\#WF//[<
P6_^)&A\.S\2&H41DE(#=:,K8Z*(O$W%!MN'".C8I,A[::ISX*Y90KB$K_80RC6)@
PWVP/U,B5.]W9^?+(,5F%%YK%<0\==0F KI%6.!:UE)-.%/*R[-^0NG&--K59KPV;
P-P^ETBVPD3*H]\>H> Y\>="*6,Y?D)RH[ON$$65EW*!!542BP;L>]G%CS*Z]3,G2
P3Q2=H7!%8KQULGGVSX[B47.<@!6:J=&FYK]W9HG>&L=C2%(D/.'D]KU\":7DDM^-
PWAW9EN4VJ&J' "8Y$=T<C9@6E-%.2N4H\A1P*P1ZN7:"?'M]%!'.LD' ./A&FB$<
P86J$UM=A=S.KT< 0]2&,DC9Z[Z@1A:E%=PB_=]PYE)0^Z*%Z]$?"6H,Z%4<P>.W_
P\\P#G=N";P0NCDL_2EZX#?V92;_Q6:#U8M,.C%WAQB64R<TP+,ALV:1*%\D-WAOO
P.&#M:,2-X0VH?"- C=C=@$40/H.L#('Y2DP+VQ)&;L"^YX\(R$?5;-_]F\4,FL&[
P/%K?@5-5&V@\[IJ$XWD&+#&( IB2F$\H_3PO8!-\OTJBD+^OZJ$A3<NBH+8VI]W3
PZ8[&%,^6!X($19)(LXR-^T)5O6E*V7X(;3\%EW^=O,IO764#RUM_)&*R=JX M05>
P(WP.2/ZZ%GKZ@82IHA=@LV61,AKS;S$$4N#VDHQ0YJ[+NSLZL%[[5M[1N?<'9IBV
PA?J0MXU##U6SN.>N#,9TLBJW@>O;EOWPFT=G]VH(3N9\U@,D6 A1DP+\O'UV)@SW
P X_"_->-1R(!T$V@E@"):**0\,*F7,Y8,O$X9KH=E6->%SV@W# F8>DM\-[H)J]"
P5$V/22P/B"#N/K08S\:=KVZO&;3VGL!59_YQ3$!X"" ,V8>5XO:V1_*[G9_9N/ZB
P:R0J?)P"V?G? <%<*J2QFS[ G=HQAAH3LXEQ\T2Q5Q0;AWK:[CYI8@&5V\WH\OQP
P7I9([ 2.T0Y2, S6?_P(?5E 6N$FF4?MW[S_.("8&P:X44H60A#WK]7SGU:OL2E#
PPZ!!I&HP?L3$B'Y:2F124!E$)]D4$@D]//6M%K$CQ=1^%-LWX)_NR-3SUU&#D7:U
PT<:+#?9&2+ELB='/N8,4!E:K)XQ>0)8?-*SH)V<</_7]#IRR\,_;KMW;K4H0Y:QS
P)[C-0P"01RR!B@R19W'2>Q5%TG"A!.Y^M00G'B/?RLG7$T%=,)A?TH7KF5(<KUK<
P=-$CF_AB46(3DGG"2F+\@5R,+/+C"(4I(S.^_QE]BIE:T@VN^)V<%/A 3)Y0-12T
PB9^,'4 'S((*+SVJGVED6I&\/A6D)?[#Q[$L_A$W<[VZ-65<6#NQ__[.P<](1I,'
P4\/,2KG;W9<^;>&W:,Y=BFP5$VB=UB5F%NGFOO_5$WU'IP[94.S[@B?/^)+S26 .
P,Q_H':1U,UE0 4C)]C3@>6:H21/2.54P[@-E8G:"LQEXM#;]C<N5R=0&,(B3K3:;
P8*-RBR\C7 Y>M@_J_('D([_=/_)$8Z"C T:R_<." 3R8(;<?>R#CU/06.*RZ@$/?
P'P\2X+]KST;*^>C])!AU(TUV)<A+?HM"<6%\O'J75P1$8D@<;S,B(JBIXB4,T7YJ
P$IB?E.)C4;?%FTGA%&ZQ@B/%(3DPDV4\C\J9UA_5+!I?\+$:PX32P=U4,8% 0H1?
PA3/P6,KV1 ^^S;,=%>T QM@]L( =DHLK[$3L);$[567"PBW*/(N0F'")%KJ>=SL#
PUR-/) 9[JW-X1 4>0V(P;CME'+9#\>L@QC37H^VVZ3R'0=B[3IH2*E]5ZH$Z2B17
P O@ECBA1L2?!E"*DG6@_N)CFM\C.I:K42QY!=JVZV:?@7N6)!WVH3\VZ+EZW:B)*
P4;U(CE#FH"U[X1EA&-"1Y?2?U61C?X*? <+Q&3^_D?&70,Q@!6B\<) S;!3R-0KI
P4TU5)O_VY(G63'6',-(RSMB#5V2._<'>.'A,6][89Y03J)L3\-L& [16 [J\.41!
PD4@3,H)5T<=6U!.6*.T5>#I\99<C623.QKK<G**)A164U %B5B&<<..#MV;_W%**
PO8G3%5FT4E.W?W<WEU/*<&3=\Y/S<8/<CA>(I<BIHG2;%M?,"X@4QB30,S$,T[AG
P#QQ,I:^4,'_L2S@F$F\."(E O"MQXXZ+V,D\;M(!@<I?N\U1L]P<N-D>PA[A01WI
P %8)%)YF-3]R8JK!F"W7P4U62<8_%YGO?@2K"<TT_U>A@\HQMVV;6B+;X!ZU2^O.
P4 2K)[>[4;,3IWAW!Z_LOI;BI[4 W_>5SX^^3V_G?9?E^#^E#S"8RR;)- 1Y[GQP
P$&I/ZFIFT3_C,&7O8_R=*B'!B$5,H/O"5VGZ53F<N*#GDO6/M*3*YC<V!=7>HJR1
PB@=&KWYL\A' 7D_#XG"NO._6MX!-PHBQ-T%E*!;^_&3RI'IB4%_(&V$.':D\P77:
P/L'TPN*W?(/.5:E*[;'=BS@58NX^U[+'[)7; W6 D''(?7$U-"T'IP'9D$_<5%*E
P2W&V2Z&[=?DKV% .O[>&KJXS=5#B1!?M9BS!B];C52%S\1H*[H8Y6:*$K8IL(>.5
P>T@ %O+,=8C9+:A%*03![>73 C1\QR%EZ>IS_BG7^)TL?Q@,AQN.C%(&GSJ,]2W+
P@7L]L 83]=W1'W^0FBJD,KW3^_IDGHO>BI0$9*_Z>4;9JVK'$ELZ\9L[L!W7D&^V
PKL@Z^XV01TAK?/,&I!7^ F\O]O$>'4RB"(.S8_!,?8EAO@,U%%2 )-B,OA7 977I
P"_G#PQT]W'8A \S_H4V<K_J8@2#>$?63'#2IMTJW%%%PJ:5"XQ<LK:($S,CA]G#L
P$4)5X,^AJF,9/=8($?J#HEQP"/0 SU=:(!(!FUS:NY>_"R40& KJ4IY0+>44.$Y%
PIX2L0XQB5VA)Z,\I>::8;:*Q\./P'S<X+[(>\7T6[<P"ZU&$=-%,YK5\KL&1XH?S
PRHQ"J5V"0L9%_.T?S(;SGMND+M<;?\5E/)D]2;_WOZ0KA'1Z@NQBZ3XXFT_VZI05
P5O40#L 2Q"\&XUMWGY(&'#PO(F._T/-1@__XDJB50QH<NS<&TO_Y:HNH$P_H['JL
P8H=.=^[U*5HX3Z+_1*?6U)I7K6Z-J;.Y0]RMVR(\V2N08HO1%!104!YJT#:9 S1#
PD]Q7)3H.^1P"#79EGDE%K8=A<(K.>'0"ZN6R\^$V95NENI5L&REVKD<>$#1[?&N=
P.J3S5 #TMI!)-"T[:J\4JVC4C%"(@U9C\HU]%D*C.!C:-J$9PZUHU\Q]K-OZ:39*
PS/PO?'8V0;^'.0#>"O7.6)/D';JCT?!I O-5%8%//U3* 6L2D5_HP 19@ 4G[OI1
P8_M3DLV[\O9:^EECT#53T%MG3Y>"!M.:T-P$KO&Z%+!0GP0.$HD3]LLQ=)?(G"[X
P>Q8PX?><")LU(/7-08N&$%R+++E#X^3\%1FBU*EP29U RXN8<!G&%3.Z\$K%:.2X
P2%/]W=R5>?G0N:IBHJ"SF8DIFU9-T.QY@(IP_;CRIC@J(*.\_K]-0%9K0UL);&T!
P]UHC(NLKD<\9"]DRMW$@(3>38*WBHXG$3@T\*@%K7@$*JW-+$GFH_?EZJG22M>RF
PQD&!*]8NN>?C_$0@)D8H2ORPA4QS7X=!!W6UT<:H)P6K D.[?-X@MN=Z[@H((S>3
P?9<.F%%.B<#8DRR +?>:W3[Q#1T+EUKB,'MLFN;IJD5K;KU)W4GS<<5'KI4QE8;M
PN0X+Z#_]]H0;'S;@P1?A\F'>4^I)"'C( YM@<-D?-0[XPESK7>G_?F <TWG>T-*>
P>;E)KAC^3!5*P_-6XPT5J']_U$I*RI?9&5GQ>3SGI\+-J4<ON7J)YOW331R_YM>I
P,8L1W]Z\#.5\/1&FR8&^*3!1$6\?4Y1F2\M0]_75W#TY(O_JZ KZ'OG3)K@4ZX7(
P(B:AA^0R Y0@@';IK!NZOUHAY3;5#P:[NN=*L:=(YR-\^ S'QU6?!V>#J(4+?M]5
PAN&W"-!UAW\;7"8V4;9".MGXR7>\'P_5_@>=VC0BSW,J8_T83SK/9O7';.F[UK$/
PJOL@GMMKP2YEX<DB%8_$IE*>AV<@\GV+X*WVQ3_EL29IQRHWR5Z8V.C$TX<JRCVU
P@Y ?D<GC\_/UCJP E:\&GQJC'F'&Y,?\DJ)6L:#3WC=DXLV$3\U1>22.CV7)WBG>
PK)1@>PQ%KGB'HT_8"<@)A]'FPJ(?!_@D'MJ ND_@+%])J'Q7I(U1VFH,Z3H"#I3P
PT),.F>7J$*M;(V<.'J-I!Y9R*.+."I)[5LN#9V0S"$LQ[=V"\=$IH&6:0(S9YWE(
P",P]<]OTPCI2XP!WDN#W-'$0@U:4#/H\KJ:D*RD ]DJCH;V__T.;@+>22R6(#FN>
PPN-[&C'?>N>;+-;(H?03C>A=W?'5$'(RJ4A-92"LJ:$QQZ[=ZDB\T[P"P9V(G>"J
PD]F2=%%[]6O#,FUTQHAA6V88*\"I( 5NG>5.%X&4,1-N&]T9,\9@O_L!OUB<"=Q%
PXZ"!@-B8U2@C6P7=Y:HK6/. 'QG0'#SH"B'LR8Q=F7.HZG,+K1HSR;<XZ?(*-X>W
P]-=K(N*KU01\+*23 KA)J"RQ14O7-P=F@*^M\L[9JUIQGJ< =9"EJN-IV36OT43*
PJD"HF-#QN!S:$]L33''>#-JIFHL[Q6!D\LDUKZ#@^JLNWO4L5#^;G>MW"VKP#$)S
P ?Q8':-C O(V47+XLA0->,;7\W_D;BQ+$]*\>%U4N&SU,1WV=>Y[4Y!F@>9L^]/"
PZ!I.CXG[%&'!0H;J1ZVOH2?&"+4FR:0_@A2%R@U>V3 *AA!H$OB+7)+I](/<L?VN
P8R)Z?/YM5AFW0))WT*W0RO6]K;6:?J$<9UZ()XWPW,,D]BG)#WW_+C6:.GMDAR+'
PGC %[!.,2*_&.)K@QYP"@)U5"S>2%$0_Q0SVM'$=**>,-09*M%3+*5\C[+L ==]0
P7\B)C6]$IOX:6/4J@(BBS.+>K/,,,YSA/ZLIS5!F\4O#_M)JH:G!RGP6'XLP!9_D
PV8KPB5#5/ #[_S$:5GC1 <CX?*;!,>Q:Y-4BFNHU15"B03"):^A*(4=A<)!TT? =
PLR"4M0A^E.B4 H-(A2EL)9[.G_#Z*>=GD82;DN&++;U6'+^NZ"&V-7RO4'1M1+,@
PJQ78&P#KMQ5(CX(<5#\14F?!7=$5E@\51UDV9!P)'&VS;0VOS"2&N!>"9"(VZO0O
P>2IG*33,EXF5D\$@G[40OU,TW*K%'5KN3=]S';[S[^L?SQ >>*]17&);U#V@Z/C"
PJ>.6 $&3P5*!(K7'8;6;:I:S!-U!?6&ZHIG(J%6"EF^W@)<SJ?3\;M\%S1+/U?V&
PF83S *[5;:/B\0@YE<9D#>"P$M,>%;7)3I+/)"S%+(,<(F%.7)OV>+]")CC(U<@#
P>UB%N4X+X;\:(^L./O500N; -[D<M(&@-JBANQ>V@8;M4EQJ$Y",/^<]. -CT$1*
P5ZY?3WM"=0,=\AA"*G*05$=?A"@AY!KP.Q]R>P-06A<KP7:-#TYYN7M'-L%6!Z]Y
PY?5>Y=.<A))E8"FC 8>NB@ZO;'.1&A(9G;V3?'39OO7Y(OY\OI%B-I6KS2'I"@!A
P0:9O"E[D<""?6XN1).>@V)&.PPX&<DI0 "1/9FE3)1:T?WD/+K Q\U#.QF[8^A'T
P>_.F*\\\5MJ[H*R[S#S@!XLNF!G+[<HQ)[9YNU%JWF/KF'&S'JZ<,E?[UYZ(5AF!
P)Z=!]AT6QJ-'$9E7TK#HLA..DKQ7C$4L=)54^!=$Q>X8MI9$T=RNY:C9>.S%'W=&
PL>]'P:UIV;B"MI+ZE9&YD)B\;4 MA7!0-Q5U/D7Z_Y$G)9B:6IQ8]2?@V@'UB8\3
P[V_X_%R*7$31\U]2%ZIMF:5FXSTX7ZNI=9B..#Z:A#Y1O4TS:Y=\%*.LM,J6HJ]G
P<!%OMB[P%>X]4S'NC3@/\TMQOQCM?'0B K%9C+*WKA(0X,31N?U,$9R"4^P8\A(9
P;X<T"B@0F1#?='?_--WAGW2N"RP6/(;S"0D!THYCHGS6HDB[[LN*3BE_%'/_E]NZ
P1QF9Q6 URA42!0- ^ OK$35"!PZ08F)#U=K;0)B_L7BT<0HM70F<(H+KN*.@3M11
P8FK?H-;2QM*JLK6P[/M-Y$)VW$IRO1I- 1,*$):]J')8:R)C\]3C=Z!GI3HG2^]0
P"$#E]T7;UQQ3-41RBK>> &#8[+;UQTEW@!CWQ<&1 _Y.N[>H]ZO'[3[MW1IR 8;-
PV)_/ISNWK<N$DVYMSO/'K^K BLR2_G7IFB9(DP5TOF'GGNO@<VRG[W7X6L<B< 6B
PCV60YU&QA.30EA$$,R]9KIY0H95G$&*10GS_A1(+JO%#';8?49L#5:BN#S%-R1R^
P9A-M)3N0[DDR;4V14M"=/^@ (C+'ZLS5H[D\\UWZR;/FO%1_-88W+/*4QK\,@Q2Z
PPB68*2HT<=@<^$O,<EA)+.DYI5+OSFHW7=;#*#!R<P+6_5NW6GB(&</B:">X-TA=
P= 5[C%2QU63<5[(=T=_7'=<E2<(N:O=G-;MBKM*X'&2@[/>B;L#15O,,RB<8X2,K
P1.>R,^D' [,U+'X&I0<-4MF1U3"( WJL(VM!.G_OOMUP?'>2M.2UW674'3_M)PBH
P>&PK#9NSN%Q1J=CN+4JKVXVK91FL?C/^6QI2JUI[+8,GL_HCET[IT[>KT=Z75",N
P:<R-]J;=>*IXD<=40>+@&U,K]I/1>QPP):] !G5E8_"9?"K29Z2,HUHU@U51"#3Q
PCNO3&]:<I58+^CU@X]'6&% M;TJN1.F*#RM()%\I_RK@N@I63(?E4(&_-LYR^T>^
PF47E+91+7'?^07OZ5W=^.LC=2OWG97[>QA(P7[FM<8<:<PQ-)S(:2<^NQE>G)1:<
P++=I;,9S&@@4KAS*BLAQK6^2JF-LX7;%X/+0OH]VI)+F.]^]<KBU]X7SN95'9&$:
P7GRNBEN0KUHRJZ"@M*H@CZ:&1/AHWTBL@XRDBIR:DE[EF),=M/_8V@)^%G".H81%
P18[S7=WY@EG1M)F3_CZ\R&6V%,M I[[,[U-JOT5S'ZA0(\HRYZ1+I:I4[S<I8F%;
P#[,;3E47,X'(Y<T:CC!,\5_%.HP_3P0V<%VXYRXPM;?)[*_'0JQRA:X= ;\)H=@@
PG+R.?7AV =R$ZRZ^>OTN=V,))L5GC;#9"XFXH('#8 W7O#@BWP':(L#%K1;G8WSZ
P;YGX1R>6UBJ:^;!9J<31UI7%'%VG'#^K98"N=A4=;:R8Y(@.HX&R,4%V#630N/V(
P7>V-.+K3!)'51$9F/7T/;!^-L,YQ1IWW9RG!T'JW1CN7G/^;.-EBOI-BE,]C=BG,
P(^":$M #^RAQ&\N7'\^R)1;S=REFD6'4&Q?[[?OG 7L;!<:43^W )[>RDOD0_M9_
PCO[(.;:H)^DHV($$NZZ7UH_W^)-,/96K)M80:MB!I<F65#?L$%C2E=IW;'-]#CE2
PT68)7Q+80Y,L3] YH_OMR6Y#$G]R?QNB$?:$UTJ95K?PRM^5S-.MFL0ZY:YPT-:Z
PO$*3] "'UCTIF3  F5Y#?.DD1$(ZSDQD"@+-#VX>\[;%=Q:*,:]($#7]3'QYKK [
P5%T(I##?G5O/4S18&@"/(NU*;I<=Z175-.Q+9TSKO%C=KSJ1GTES"A4_4@HG6?7+
PVH%*6PM)(8X=306EHM-" G?&YIGJF\15GU>"Y! OH0'+I62<'7T]>ZVJ(YYV4Z<S
PS6WN*;/>B^%8A>8V#+M@=]5!8?U=9F3<"M6U'T$\-K>3F;E8^%WVT&\8,^ \:RMP
PNN>)V1O9I$Y<W[+D/,=$N%TT!J7;@I' K.U_L4AKIF3Y%=@3VI&W7687Q!W@8&/H
P%?:_Z""@(+'+F*CF/^%_3@$$S5*Y$ZF 'XV\ Q)B:$$>U=7EC  50M_P.C?ILNA2
PL\!?]_Q#HEY$;$4A)8S1PJPH@.#V'8(J$5BAR4HB_\)D,@7@(DH!YW)/> '9M!7_
P0_K26[J[\G+)Y-?FU(T9I#?5KN(D63JT^4ZBKEXGUR%OM]S5;6>&!^X73G>I,D<]
P!#5\(1(%*R?YJ.K3R(GQ3/@/*[-3V:4G!3,/=] 1SY%3_Q-$[!Z&]P$0KS+CC#!;
P_9+ ^(%D;0UGJ#7X.T1LN7NPR'*'DG*;5F=LQ@^:F@ V.WF>'?*SLOX2)>L9*GYY
P\ZN$R/PS!, JR1I#:$J\)BI]-+=*,"/2NX $ '(N7)2_THX[YPO(PI3_<9%]U%)#
P/@*W;*!D QQMV$]+ 36<V 2P[A7+@^6L.U&V)SJU7]UI!)Y$W ?YL7#9@BXQ@ZDZ
P5/1X%&7/NLW?XV %"\#WOY>F_ &@Y6SE=[YU7L XPG>>]DN5LW,)H\59K\<FW0<G
P0+PW 7/TD+8ZK@;6< $/NZ 6-^?%K!H!<JPT*PG!MI!6[:!PPO<$')]N*8A^A,YM
P">1*&]_?ZGDY7M8+S9^ 4!^P$Z#'HUI=,XQB%GR%(%.UN:47MM>@#3/=F_&7M39^
P?LXMMNAS0NSZ$1\]?)1&K876SEM[?E5_:)L=@@VRI11-$_.E$H8=)OP*)*:*A_38
P7,"E1E70H/^-_3Q30*+,=&$9=Y"FXT$P,X;+]PVATE!Y![(SPMV)-3AT:.O&5D!=
P0$ZBT$-(C.A#T=VAG.VWHES\&S;$'+7=PM*J8YGACY1^0Z$GAWE-$K%XBQX)@DOX
P[T.UR280UI6RTM7;A>0=S4:F8B^:\>-A%Z3@N]1%*@P'@ZW:*1ZF6(=:  #^**;'
PJIGB\/ALM3Z5UXIAMB>PA&Z<Y/5ZTN/XT:>Z5:H\-PM@3,R0]&9<S7/[>]V!:&D+
PU%LO?=-]S,'GHD#J0D5$..+\ED"VJZALCE(7NMM2)I.@,:A'.A$U)AJS.U/8=G\*
PI/.(N2A:]JZ!BQWP5%F15/X?Y*/>-#YQ2^U3!N.M3CHF=$?G&^SU;9OF]0H'Y#2N
PN6T=4\"+[+B E>D/B"ADG]L8:36V=F!:%P\[*U92V/C+> ZN[/?<T^R)2--NPO^(
PX$OVE_ .ZT].@]7 DF/1WSL[1?0U@ICEM>4YX*/4V*=S 0TTOQ1D+HDI7+G+@9#:
PL-L6C\LF\$^=0D AK>J[C>PM<6XQAM#VIU'0AJ8-(*0M4E6IX8CY]O=)Y\UPV/$!
P].B04S99+Q[Y#M7IDIZ8TRM0PV,L^<>/D?84UPW6UNGN4Y%TH7%:"BBM%AZNF:GJ
PS9#_*O_#MTVP!,!IHWR'WC=(=XS HIIK4(9F[CB/=A7%>>H0RFN,=0XU$S.Z";@"
PFS*E?G%SX'_'*JQG(;%G.\EF#*#J5_RYZVSF3F%E,<QS N4;?8!@N)G0U/1]I*R]
PWI\"V%4^F9K"CC0:M$!Y4(XT\]#56#6EP&[W/H^&Z!16H)./$1VZ:ZF_V2(CNH03
P'W\^GJS!4!AL;E9(),VJ=/(NO8TR#%8,Q(TA"D2"J#GCG^S73T&MZ=(!_-0#1ZOA
P4-'/HF[+#6=ZJ68:?'BGB\OW*Z5Y9!*/PXA@G=6,$ZL >#$50 9T_IM@N;-IOJ0(
P%V.E-,!SWA[@$SKR,S1&LU WT(Z[QN14HQ)E;\_<UB,=/HA9XR$99I\DP-12;I&?
P- 3>H+NS#O2./2ZND#K-BJ7X/9IVEYZ1F#X"Q6F%3>\UI$C?65J+F,)IA WW8)V\
P@U>Y%[G#\ R*HOQ#X/D&C!+@?MM^P@$9<#K*-]UM1]NQ9H7*1L3'ET+Z+; V(M)Q
P\;W=+RB!D)R[C<[,+2,,%0K=^R*UC?3 Y<_UAT3 8A[BB1D)$F_:5QJ.^Y'K M9"
P>V$@ T[WF2BI:PL&7;FW.#(\U2)\&]K(:T_$*OC.)$4BA'[5W"[JVV]!NWL?W6T8
P:$JQN) /%Z6YHEHP>WW5(89UQ<UFMFRRN0?EZ6YS3/Y#TYZ<\YRU&2TU"ZMDD'>3
PTP6&4W[9-@EX:I7"TBQZA!UN4'EY35_^+?7S:)@-CPBFBT=?T@>]JM@*/JV+Z1OG
P<CYV@R+07K5\]%XDI++KD#0>@YH.+P%Q7BC%,!-%8F\-!)Y0GZ<C;YW.0Q4;*PB%
P#(Z&:Z.JA!HER.O%%ME%BF-E$13NJ_,; UY4-?@^$W!!6< =.\%[ VM!5?#@WZL;
P[V+,G:W])P?X3A[3B7$T79JZ<O*\'Z^[;6WDOPEJ5M-+LFY^U;4$9[(-Y#:H.Y @
P@N@&+XN?[6TR2ST+*I7/37F&T76Q-(1R@7N\YO[MW$E10PB 2$ZVVL)ROIK)GNZ$
PGZ4QS]!]8%OVXA"*2FR*_:TB^;,_YH7U4:Q@#;FUU,DR\_@J*+P+S548U3]FM=#:
P%FI[C'/,&*BN/BLVP09C_RRLEV\45Z!"Z%FTN5$[WGL?QNNSQ='1^KA5I);=@E5D
PKJX@=*:XB!^VSL N8[^@W-L&:X5>@?B$;-"F/ZU[BC$AR[MP:%9H3M;%DOE5%^<]
P3'^_]HP?487'!;?9-!?Z.F2_:6G(=N\H%"-F7B&&RWEU*)B4Y5P0)%*&.LI"^H_I
POL6X]A:HM'XP\ZA'Z9+R.5Y',4H@'8?;DN/K?R?Q:]4L0>CDA\D*JT<^V&]B1.%S
P41T1,3(Y_R4UGRX.=1:@O-+#?7CE" +;!<&+7-OA0D'++Q[]858?)>VN2V=H8E]K
P9I1NSGAP$$#VB!REC[#XO_%W O0*]YZV!F\(RAK"==M__*!F]UQRT0 A<$&$@S(*
PE_ND7])EQ5ZBQ_5YF-%(I54E?I[36P7.@"/<V8[O_# Z3-POB96M#-ST<PD@RD2C
P@&"GIEL%M>=BDC-@C1D"QF2]H.A6,+(I/@Y9MM'^I&B<)JO;CST8)CXXLVACY/_8
PK=V0*PZSV[<_^8^4A(8\?\ZJF 4+9:OO"[1 5MBFNRJF[.O[4*4*BTUOM&]A.4Y 
PM9UO":L0+6-BA0(_U%M^/"+(/ L-AV@F&-CIH0?V]9(=46""[3UCNP&34RAR!@#$
P]:0^#8,)DJ.QLCNUGHELFLC@?)N5N4<2 K%FQ, 9-ZV9_1DM.QM&"/"VH E<C]8Y
P$\*-([(ZN Y+Z(4!E._F]>&J8EYG0F*K1JI?'MV[EH%=S# .A56<5%[CRTM<A.4)
P$"1=1?L+R)(.J\?^?IE=_8TP'M;"<2ON005_# 5(:HV<]15R/ZRK%?2ASJ[+:^!=
PQ.&('.W0NO2TMT$GVZ1L)6=&0##A,(/-4LWMCXH#0OQ&P6?J\U:Z*?YE)4VG7/GQ
PP)ON-1+9L$VV/=PNI!G:$I$Y_#C&]KDLE?DR+A08I9&#+8V+:DHKC>ZBVM[8O8__
P>4S(2!$"MJ"%VP4K3B%B#1$I8?XQ<1.E$<F=-9=U7K# $&R4=QC*#79!RCN'8;8S
PKG[]0==_/HD^#N,APY\ G&PUK U=XWL)9[ZH#76QDG/&GC(I4]2R$Z+[/HH#E]V[
PG[,J8$^-#@11?I:LR*WB#>>VONS[9--AJE:$+ZGKV[:(UP+:'CL52^27=& '>V6&
P3-[=>US:!X.4K]N[%\E\4*0OU=RRU,]G1J"6L:QY;XNP:6XQ28&#Q6T(>'I^HWX#
P .UM^5*A:?;FRU6#\M<]ST  33M:76W<R9:_*Z0#'Q$7V!ZKKB&.61&\BD[QE<Z)
PV3CJP%.:#)"D$-T,<Y/!$%@B[Z2[N6J;=,X_-F($<):"\NYR32_S[TQ /G^UEPU#
P\VT:PFC2T!)/+9RG8^[BD8[!_WR7SVO&5 :%.54IS4F,EVL_QB,BJ"<5KGJT5N7)
P%X]/'K1*E;]2.*-$0X=XE'6;3V=HT1WJ?$)6>P/_E!$YXO#HR]X:&\A)401QL;L8
PV#TZQH:\BYT%3N>7";:L09C\X/G]0A0GXTMV7)/EOR'UY 1)7N0JE$]+1[3%=$=J
P-65147>G2ODZ;A:?B_O5OAD 9&(7P'$+^YF?@]CICME-Y#J7DJ()35V_:D\DNT$6
P+ITL+/(>BJ_>J)R-8_K@=!2QGYKK_$U\P*2X\UP\GED\31'S EN71P6C\, U)4^D
P=D<(GNV/;"9QQ]*]&XIR<1UNXE$O$'368B.A0OXF-%ELH.8A "\[S>.1:I+Y#[<S
P166JPU?]%TB()5)U5^$-2\(V63E-\%JU.'GVQ3+I>Q3I*&ZL/XG>=S\*U)WUGYL[
P28R\T35^F#(V#^#7N4>+(%S6XDY/@CEXT^B5G86X,<,82R_H&5*-"V/+F4'/!?OF
P;G+]R_FD"K(Z"[.Z$G?;3.;YB_&PPFSU0C'D7\[P%D?=X-B3DZ[N,;I=7D1Z/[4*
P5D*,3$\?UNVP))>?,3;PP<.U ?/6+,=D1=YWW,*#<U>OM<YHVVZ5^N,@= =9SKX\
PU'#G__.ZI'U5,L*EBYK]^0-R*'O<UXR@DG1L;4T;8*EAX8]"UPXP4N$F-7#L(7_5
P3ZL:=J3TX=I-".0_9_@C8>N49L=!N*>SDB6(_$%ELF,NJXO3@70XNJM5SJYX8K,8
PGQA[8M.K>U"GK<P%C/D$$#;[C<V&$H7 4]TJ@&>EDK"87,LJ]IB9P98SE\CMM]RS
P]'9XT^;]GB1Y))U-93TBZ9L[1T#4QI[2?135T@1::'(DKCO6T\T;<[T3>]?!:?AY
PE]1=*AIUV=DOM>A3]--KJU;/R)#.-%M?<X+J,LY^;R]@K=X#W*"YF_NDK_4#RA'V
P4-P*0DE0+/(61;B^DVMQUA&Y^>2!)V.Q7'6?6#MCVKU?74V3BNZDC/NAW0V4^L%T
P.L)LS;17,S:G/&5_*_PMP4;U822O^!61EP$S$="0Q)Z.E#%(RP! A2VD00U95@'M
PHBD(GJ)A\]-^F.7B+!,E).U!H]3WC]H&'>ICCMTZHJ,$VV11Q:\,MH8X1517M(J0
P!$M__ 3=+(IM:ISC-L4!)J>#MN8M8]_'/7JE7);*UVNCRR1A'+T&NG1:!@+VJA%?
P6VB5'>857<\O/"&6RH^CK_RA#GW.%4/?4 !V:W5;1A#I'DJEL*[?Y$N< "0!K<!&
PVW[O:Z.:&C(T[08^.(\P*B:3+V:\- 2^!,C35J^#@W;B%%'FKG5V:_#58+"@+UK-
P3W,)5V0SF$_5-"/J>-R%S%&V,& KGEYB5W>I9>%H@Q=39["VY(YE4P>Y$Q_P)I(A
P DSCRA@'-YTT_KQ N?+&(7T<''M8.K1<B)MJ_"F#KJ[OMI\ IP_UCEM$,,C-A@&[
PBE[&V8D/[K5Z'P@KX4: (1O<L"Q""TT=/I52?>VLQ<+K,&SY"1J ]O=9]5FD_+9;
PUV\YY4$P?Y:MCWG9]_V:RM8!SM')TPRQYOL7/&U5@IT1>-V=#-.0EB%@S(F5TKM8
P'"QDQ%L=RO1T*+]@3S/^+E5+*Q0JILU.HZU%1(?R7Q^FW[G:%R3F:$[7[/TNRS%_
P?03<"@EF^[,QLHD>+NB$%AH>7J?WY[7._,L$0J%1SV<*;F<X!5\GA1FL1<;RE=<5
PP(K*%1RU,NV:P34.&NMIIX%3!^4/(5C.?3N2\=!IU,>SC5F,<0I?KE^LL;+(.M"V
PHL'H*NT7)O>4J7A7XH*H#TE0QY=KG"+H:-8*Y:EL_UC.2#*BBX7A# T[XQ'4DQ9"
PV7L^#[XY> RR7)J0X1 J0V;';;#_'/N?JYVUY;&KOA/>T-^YBJ=4W0*;H\PAVJN6
PV@"6 I%]3T1&1-YX+9=RMYC8]FHZ,99#E%A7Y849&76]1YC5#NH.&"SPSY#EH%)@
PC<'4>P&]+K$TLN?OB]N+G2T' JDZ?$&'U*</$ 6)QK4VG\&76V-Q'U_.IU&12Q3B
PG2VA$"8-8:;-<2G0OA2G5#&R>B],9ZA<P>4T#70K<QU9H0#PZU5IHSF]1:]TR]<(
P.99F_1+1+!#B-9_Z@X*.2P$&/5LA;U^I<)UHDK,48.F(@1_GB ?2*!>Z=3O<^I9T
P*0!"V#++_+D=MR]$I=7]TT74INV#5'T;O_$R/8_);I"#G/!/BT!4@O2$7MRL8<T\
PHRF]V']%P#,Q,'OW;"6KDZY4#WK4CFX'26#.RYNR'TL/5V.T[_(5^/RB(GKEH-,:
P!P.]%?P M<AV[ZP0I^P[8I4%C>^SG2*9?.=D?KLLVIOHC==E(DN/8-T=69O74=3U
P7%[$YV]%6#=XI=:?:N)<L.R*\)MS$42<NB-[,:$,SLN8=7!Z OIDLJ3N*K?;0LC?
P:K51" G+ISV/Q4%[G:2C\TT_A9LK#Q!)%M)4MOL%R,A B1]$@4 D-# ^_L*Z_4K/
PL[T"D*@OT^-^CT&R(#*!/F<.$Z,(;<*4_>RB,7BT^)BI\N/&P+6+YG#/V%BHN")>
PUQCI"]N%Q(C%X5MN4VN .,69M1_]<,QQE)3B^,9?,7W3,3\]ZO],Z7/ND-_'8O2L
PQ!=HM.WN:Z)DY4%3E3%?'R"!GX>5,]@SOTH#W_K+4)?686W;S@F%-Y*^D#N<L9Q$
PT\X4R]'9I>YU+8+)=!)W4IN2JW:E3G"!6_W;/(\C[L>I&)RX$'8-S5Y0SHVE3!?8
PJ>$]XFH3,9?7%*LSC=PUJ/ %EOKLF&: ^7^J],I2PLW"@._SUHBB$6!.(K=?S;*N
PC9U;G7:\%M!=/) SHA^$WO/0L%">QOE"HW@3Y?/,VM%RPY%V'>X!2;UY\L(CE+H,
PJ<Q#MG<H*C;HI/Z\5U:EELM(N6V#K-E3PU'>HLE>SD$K2?>'W:#>X)#0*(Q(BV1H
P<0_6OV=0KED@KE*T-&RW#*;.ETAZ;2Y6]6T^\M7SOM2TEJTXC-Q@Z)E:JA[21M7"
PL^M(,1G;LIH.>?1JFVL-ZQ:BN65#S!/[')!W49N^[O@_\E[*6[EZ;+L#@D(&N_7>
P&8J[W/XRJ= ,E#9N[72X6M-S2\T$B4?N/<CQ7EWR;K:^+$1-:N;S2851S NEWYYK
P*AAY@M!;Z$N8V&*%\0P-Y- @]XIN(</ E_Y1+J2C^AWR% !@ZF,^KLN?@(0N\2M 
P5CI"B-FYL\N'P :BQ#LU8+YUY +QO)]5:Y&C*1_D._"4-5P7%?L*%QJ0C^F>? /-
P&0'[LW=+WBG]IO'S(UXJ8(*3KNFD<1'-<&72.3P/ZR=!A L5+]YVU+'PS3&E6&2U
PT=5NP*;$2"H8R2\U)G+]-%5\9H):6F'OI+,HQYD>[.YTT2&45Q5$0=&H), I!#2=
PV#VYRN#WGUG165,;6A'5^RYH5J]ARVU.GFPEP/G'<[>*,D*61WQ.;3J$\(>CM,%Q
P!XR9?U<._RI-^-):9>&S@QD1EM^&0=IG(E$JR?P963^VE=E)$9V_GM\[SC^C)W)@
PE+A/&9<.&'1\[[F>7;JN8\O2&GGS8!W2]?#-U^F=XUAR&:7V\C85K7RDGTDZ.FAQ
P!OW__UO7^K=*<J _]I8457*<2 >95QYV"2=\' ?BULDI"$U)Q^O&3PLBQ-0J8PD7
PAO&/U-P:W^+XKCX&GI?VKZ3\6WE\( B/34)O2LF,*:=DU%%655R##?8CSUBU[6H,
P,EH*@;"_R3Y0?OH3EK>M=9-)71@Q[AHN:MH--6Y9PAO[SE<%J (XA#QV5$6!R+A#
PHLN8=0-4]/%W==B:)"MHT6#8;<^*)?;6\+H46"*'.Q" )\#0:)@<?9\2(3V,M(!A
P9RY;W=*VI7LU_%4F<D8I1)6SN9_A1K_V*&\GMJ=]]1GE[7_X(VF'"$L)#.D#XA"T
PYC@09QO?IM@V5K;M#(3S^"9O5P'C!8^#\ 87"*W#R#\+HAMT![(. D;S;9KF$*NQ
P,-3A^W[/C0HA_U!'BCHTP:!_YG<O<=MJ+32K/?"JB'"JPB77[-".C%'+0LX6BFQ6
P9C^4$)D76JX?9IC0(-TLZW%*\<]59,2!+$OV)\&BU8D[1FKF)=@13*!0DM?'P5W.
P*290SXL*5_'SBP#85%J7SPE&9$7:#(-),E)&MD$9(G'?#K54@A -$Q2>8G!@&WX(
P_/S#.2,,Z]I<$.[1>-,;#V -.R:J@8 #HQ&@%2:;EQ*^#EQ$['-=;_A@'GP_ U*3
PWIYHY<>ETS(TV>$?94_SR,<+)6S]GG6V;T4#W@NP$Q8#0MS%#S%/QP-^1IZ6$5K@
PP80HRXSBUB*7^?[GWG(PL8(V*A#SAT@*_G3W&_*_\2+-;<I\V-8BWX<"P_1=0X5#
P>"D;R::VX^[@;^.$HHM=&^I"0W-?6# A%]=D,(>4B3/@>Z:.GMA)/C4%EL3GVRX\
P8@&COU\9W9-Q3,\<$RE;F*%O6.3H64QER'R<0C_'N35I6D32.<,(0%TM+[S1ABHP
PGLH3_$"^I]KH&_27G3\\_\L@/$G/S)5@RDPI>5G<SN+B1^>DTDB02H(*-IL9^J)#
P5B94C)G@0:@VMR$H*>-TN%F$!LZB[>3-"BMF>?[JXI+MN@A1;N9$O6M9+;3 J?=0
P5Y'8Y-'K#C7V\Y*-&>^@7UG-C)-U-WTF1%DN3Z<P5'J7;!2:M0KE8T'D7+@H-HE7
P()A15U\'ZO3^;-:[[#)Q$I5Q;+8Y'-<@F@JKBCEH6#H35V$SGR4#RU*F=B+$F/2Z
P_[AST<FXQ#X>V-O@TV"0I%%F/UJ^NOB[*C%._/#<ZK=J._4X','$A Z?:3K5W_62
P4IE'QZTB<OPZDE89".EOB+Z[]E<:%-CQ7V01VQ>6,(IWQ,_=&G1K@]JO++7T)$%.
P I.$PJ@EXY.W^R"8S5+/)LM'($E[/A(G[A4W4='P^-+?4K0\F>P,G,M_.*B 9EB5
PT?_*?-[#RR.&Z,R!:=/M7 /^0'@3 \A@*&C#((^.AS(E6$7TV(D"$//-W0U\]VR3
P /)AS_0R&-BX5$ _[+7Y[5XZ:VE&$CHK?,]EI3W\G2N?YQYMC)3G":$%.\K=NGYK
P,_2S7614L.8 ;<Y0\FD-_.3QSZD_[&2"J& $R0[:QT 7?"F%K_+JG;^TT:KFTLXK
POGKXU[M7@:+IHD4VC=J%ECAJ2!-/[%%5*B5CE<26.+W@'@%/L].%8P3!DMVLM(\%
P>Q)8W0$X1&83_5[SJQ)ZT-:.LS D<)81@2?23/?K^R?_]%LE7XJ*LC8_3#DJAKLQ
PZM<YD&WQX>_.E5#JPRTCER7%Z@$:R(N6FVWR\C<W8-G=[>%F%2+)YHN$!#$"C:Q\
PJ L4R<I5?^9<Z/I_!^1$/UI("3WK68%)&Z9N<T40F 8?[B.E9 I7^><9S8_,B+1M
PSCD+.N:K7Q]7I?T*EB;D /^S@<&Z.P.Z;/ELAFC%85.VRV& H :3R-WNL&5MN*8:
PP\BS"&%>&29[6F7"=*LV,/,6_TD&!%)O8&Y/8"&B]@NP^[NNL[4SJ9>2B\O,G(4B
P(E.7UY$.(7EC7;:0]*5@F:H5RP?+?\S$%:PX]FU-V3'ODB-.&E29AV24VMX_A1?3
PQ]L[/1S>#^E3BL?+%DFG89;YZ),,5"<\#SV<1QA9TY^/J7+?II_.9^*#G#O7Q>PV
PT;^&S;SRTYH4A?$'UBO9 ]]75YL,U!7!<)B9TL]NJ\Z"&U$Y=N@>@4E218-,/V8C
P%=<@"15"$[CFCDQZ 0MJ4\BU';""8?3\@:Q2R=EP*:KQC)<AJ<[R!$9&Z,Z\KS1@
P1NW ,RHPOSQ+O\+9IM:#0W_@&0HFM+9:$E4&Q_)C?];J).6.C7H-QK:,D_.FHG7E
P.Y_\JB 7,0N6RF([^N(,*]P%*BJ:7L^7]V%L"$4UEZZK2D'\+.?[Q1[M@=ZD/L2F
PG=8+N.HT:\_E8@%*P3@(-'G&/:!^UYOA?OLG2#?$DB=!)]T<(/+EWI4-M&P%G%P;
P,TA,+Z.JZ"8T_(V;?4E?"/?/,"/^DCKOH^ YN#Q@5O]+_=NG_B-Y(3A%3&!"QH%K
P:!*(%7T\4S@V;23:@6&SNIRZ@G)!ZAV(#;:K]I;605G! ;'XB4LZN@E(S1(<:[C3
P-412)12J2 RI>6C%'LE2WJ)VKJ;@[@DN^BUO*)]#'2X*D^]*SBUK)_*#" T9$&.?
P"H UOC6]C7P%HE0S>TDIZROSV%DQ@<D@!(L."03L?8D-<])B(]1U<6DT?&$DZ5J/
P=P[#AM%*PVA?0%JW7^3T@3WODOP:_G#.R@A/<P!CQL,&&W5'P>@APVCYAA:A<^3D
P3LZE?#RU8V?>R('YR2<?H<]Q!X.775IRB>VNH+OY<)3_-Q.3+;1!>JDM:DCWH)55
P%KC/N4[=_L%*GB#8W',&[?ZSPD1TVD"MLIP<7*7*VC8/0R)\2NC?*,Z8DN$=5C7[
P<%*@):!YE4K'^P6&/Y=VF(LC\1$O>"I(MA+;%$@ME\\=\RDFGPNZ,,:<=-'J_IM^
P(^QY*7\>IZ4HMA/1[- L;%TI<B$6" ?W551#5-8Y4(R/ 2N0(U4(\X*/-F,"KM::
PL!Z,J=\01/Y<*?'Z,V*B-P-AJ%I[W%/QKF5DM 2;U W>H"K:8;HS7?8ZP)?)P"^V
PVJ[M(F)"8I&IT$DC:4A(E:9-M0G[D+N>%V/(YEM+6;7_N8]@P;85(%2R:;1"$*]>
P<70C%.<< CSOAN\'GAX#O1L+TG"(/-6&V3DQ[XX,K\/+9<T)%/3KV%?JFS;!RBT[
P,<[MO$'[-@Z9%];2>'J?'+\Q$%8U+^5L8^E&'//>/TI1PU( F=A(:U=.I"%XXB?*
PPM>B0%DWF"+[^"$41M^51AO/LDH,'T(#$M=_W)9(T8QY.]_> XM,WP#YRVH/A==V
PQWVRM0X [BOX#QT:S/>%"W;O.YI'*V ]@CUT3K3#F1E>H?\&,$OH0);: >,QF^4,
PD=1<S:Q>$>TUV;Y(6P2WAT3$5.24''MB7,Y+/9^[%F? 9:R>LT]#17^]7Q%V!3#-
P!9']^IE_0%9G#".!22[Q!*=$HE(/ )QR4]G) =SX*X,T5'W79.07ACLO'>6>EI%I
P-*^SKL"X@R5Y(8J.&M6<U='NQ^WXR__4EXAC;X9Q22HQMMCPJU-@O3?$D&XILQY_
P3=R/G1#IKIW<H^V'L%,O'=P?\"'[7*M,'.\NVY>A77V"KW=6DJ)"=@AK?[Z5O%-$
PYNM_UP+1H;O: 09?H(8%)?,&/N.':2W(VCS48P.IMN)B/*D&^\),!--7WQ]D_D]!
P9%E2-;?"'2?[Q*@N$ (5B'PT"?,I'($ K]5#VQ*K%2")C1"K1\PEE]^\$D #Y30C
P4WK#@5$F;?'L!F;9%JN1RY!NQU#I2R7L2OK.7R/DTX8&(#0!#=D8_N>?*KF+(M]6
PU2<2%E>=SM<2P@S%PL)4@]MBI1=FC!J+$HG20NP;45N:[L[@PA?G<6P5T LE9'DZ
P6;72("!7G3F1UMQ'ED04[F=%U-Q*X)Z0WS"T@;Z9+'E>:,\BA8HUC&*L*(U)8*J9
P47Q8[3#SIW[D6]PW0 WQL?$ZSO;EEELB;0FD CCXW Z&3;[%PA:R&WX)9E QON*Z
PUQYNMH2X:EAK,8NO'9@I#*@<Q5 +@PQ,92NA9$J6/(^F/S$3-WTW2,!\\G&F'_!@
PL<5BL6PJ^8F_@HO']H!+L^P.%F43_?%P-N:,><1<E:O\>B;-+K0(D5PJ9FA+L,4Z
P?JV:P,/@9[I8YNVJ2BO*LCEJ\C3,S5&3QHBO:*H4AKIF_LT@,K0DU3J)S!. GWDK
PM5.&H<_ H ;;K5L=)<6]B&08DL=ZT/JN=]>AE$G'@P(52<S/M3<9*&+$<@]]0WN%
PYR9<[*,';^[_UV?UL*LRF$)Z.J];F$SZ[*4 AVIHD=.6=!7-4PK7Y+BT0;Q@N5?<
P/-,/N@#FFKA#,RL4OMP_VG+$\Y)B/N()$N2Z8X[7?<V_W'J>,J,W_.'Y$8/27@KZ
PESN.-KP\&3-@';SGHWUX8,D%H*M8I[IF2QI0$\Q,BEZTYZ'.4A?1TQ1Z)#X*FJ?8
PD/8=53?4>K[T3S2=^C+D^;:J+ZDAO(:"MZ0KV]+&(#M1SQAG( 6_G'P6O/B>B4(/
P$'+\5'KGF#^WV6<U=<MTMK-LF8(8(&P&?50QVEL2;W2=IZ6X^5G<UM27/>A7'NN+
P@@?@O/,6>5L_G<, ORX9\>Y3*VLQR6> C[(,],_4_;(I_M[9@)6;4G0#^4(CL82P
PZ6#6/]^H#9HK@\(0*&8M*IVU$27P!U^GN(B#O!I)4>V7CWL\9!51$#M;'TMP4I"C
P?Z?LWVXJ5I_U <@I0*CV[5?3H 87T454ML+A-R-/XU5E;EL(QO\$-K^^",5Z9FU"
PTDAJZQ4O+D0%$S)217R-Q?.D=8J?>F=&J4JCIP@V=-X1]]8@1(D74*J4<73V_,Y'
P#D9NKC-[9&MX7M=_7C (7K!1O32Z_W*?<]C&Z-_710GAY-4KF5)QN:2[  __L%Z9
P4-R=["XR0MH>9 \;"Q]8_&65:HNAX._YJD2]TLNR!1Q;Y8-,5WL#\05ZTK?6@_!W
P2[LCQRJ/K:&D-_X0<3YKLA=45;E$!_#<L$EG#7YISR2Q&0=B^4CU41F;S\#S0[/9
PA:9 NWN"=?\D]"%"P?K=Y6&V ]MYVJO$P=>N EEO4^'%N62ERDZX?1#(=.6OM*&@
PAMXWUAC/%RQX61/'7WW7;Y$>[J870=85*"/8!:)UV8:C[:8+\T=P2E(N/(@K"H@P
P)G-R=7*_1]1F3JJ+R&.63<'[\O^$7FU-V5ZV /$3'E[X 20,9-(Z<%)>!(<8$D+_
PK9)B0DP(0"[4D],/ B^#1R3@HR\$W29A!!=E\\R2A#4=-P744Y83<M%FKA%0RQ6"
PSV]]=_S"KZ3\=%!Y^#DL V=MN$QS*#C6. J;;<$+\EP4(."-:RT  %L06(5/#2C1
PTV;)+=)1'TN=/?.S4')D21Q+'Z AP4$LX],\<.Y.LHU(KW.BSH$*R_X#]E?.^]>R
P:U4Z*SIR>=7#(83OD^44Q=*Y!%7_T.LTQ=H7C3C,5QS.8\XA(#S/14G?_XEDBM#L
P"0%;CG5;XZ;$L\Z5[BY^QVMB'$,1V(IKK<#B8UOWGF(>6^5 )6V6S<3[!5R0(K1*
P"0 ,0-<*TXMZE[$A9Z^T1L#7'V4(DC3TXA452LC2_PQY<N.(1KNT[&P5W"4H$[IM
P&H8XA#> 2\5G#/">+( ]=DT88'V%@RY,O^N(B*X.R2_#8_43OX 6PYG"!NX>[&"/
PTBM:/]S-'O"8O\QK\4&SS)/J9FA"140?X?RDEPD1"ZD&@L! (;>HD$VO*\+WW3AA
PJ$E_[^\F:NC9BBN2N& X;WZ!^8LV'[6I%5F&F)6-U7\'ZTG]_;#WI(C>K0(N=2(S
P^MLM>QRP4*A&;-F]D8GNJP7;-YC7(5""!06[SDWA(FJYNV^4H(6J&>J#\H2MT@:U
P%D:N:@/#:POQ@O=,+)'ML/@P7RIJUXX5;AY<]\JHX-F,X3BN"A!.7:/B@+GMWT3!
P212;6HC#+SK=_]<%>G,61RI\@VKU)Z+<F@#-:G;,H?1T=1J\$3'$M=5!,*66TKVF
PGG&CCZE^3-4&&4=7*.,FT',HMG?'5"O_()YM><@=//$-' Y9L>8E*R.#PW8_WW<F
P50QMM<$BC-W<A2WW.-VGQ(67Q1OOH_!H$3.YU7H^!+3U4W]7&(/.6;GZ2&N,;T<%
P:C(*18?N]\V<Z*OWO+Z$Y><O7FHO4OVTJ@_S23R.Q6J?OUG.R?8%IOU )+WPG ()
P57+V,GX&X,#-]M!#KGI/2$_\ZIW@__H 5R3'[0,\?V8=Z#Z& W ZH(G\:<B1T:*T
P-D@^\TLEWK7MK#X=UI&G5/-53*$1>TC] V6J,%SU>6AHW+5N+#1L$BGGZS7?KGH#
P3PF\5CZZ%?&49F(:N+G]26=W)-E5HHCG)II:B<3/SCC,J4.76 2*Z"!,_+;"NJ#%
PZ64S5(7=)H8%^[T@OHM>G[%41S3FE+18KFKKHT<G1H*S(00T<(Y=5GYW. +JC(N0
P(-5;*=RLETW:PJXFK87$FDG5R6060RH V[.>_11 +''9YN3V3$GKRX1U-JFBMPZB
PRGF)AFWG8:RR"+B[3X>D&_YJ.W<+G; YB!HU;**:2%+)YI73A6&%HBZ%<O"R%HO8
P\ZW@ @_04CH-A (+YD*"U3]15S4N#^E2-&I2RF2)-F2>@(3IKY;;G(6WU:K'E0+\
P<IHN==]%3&!-*AU8LJ%JS.&14:!R0 7:BLPK%OK]&,NHS.LB8=D2 &DUF:1>#)H%
P:HDSE>,S*/'6\"++L,Z_^;D]H#0BB<Q9+HLAB<?]V$9T S"! AYF8#&0C9T)GX%7
PB2-/Y[U)QE9 [\Q0G+'L'\FSQT9XUKH 1R <@'I6?<1#GAT9&@@-!B^-Z, (\TO6
PB)7S'GY,)966)W_>KQ@2NMVVVJ-RY&+'T4)K/L!%MS/'2:>B,OQRH2 IV2VH5WQ@
P'+F*SF;,+F<)UYN296\RQ?9[<^Q_[[W>'BL$1<#WYE@SIGW?%_96<!$*[?8_E_/H
P] 4QX>=R_V)Z>T&R9R H1QK2-$%A2+5[I+"4A.CS)8 $\^K\X&VZ2<OP@HISLE#Z
P>>F&PWO&FG'/C+?8<0FRW_.\"B'2M]B2\]V7YZ9>#>.6V6R+3UKP\[2DCK_5M*O;
PGX<;7G5;6_-&@84G/MKU=]#WU%'RX=/: ^LG]R#;K#;%E9''&>$0^$IP,HAK<^TY
P;YX[^8"_!B$;#\!(GVE/&MK]M->YV;/>B]A1?$L6#+'.5]$[;I&@1D=^_J5_ T/1
P:J:%#0$72/CI.U%_W45U3$(UJ/!_6&8)!>D%\1OZR[>N E@N=/&M9^8T]EX5R5V*
PMU7=PJA5NR:TFB4((.)[6Y!6I!(.)M!WO^WNT<7QD=1F^ZBL<LMESH8";.;+V48K
PJ>;K6F6@?9TYIK35N(.Y8+(,NR6<"H5*@K9B,N,[TV'6-VCV2E%CY!<R /DB9&IJ
P8W*$K_-*M%^H@WH!*]6K!;BU[KW1"FW,J@RC!%8NS',;_C2QYGGS@K) 2W&Q"[V'
PLKNJB#Q+YKZU2]?^&,+KE;"DB"'_I7+,?6$UP2VC_>/P6'/:=R* $5>1G@2?L$\V
P=O&!#/51#4<CZI0CLZ=#<RKL"++J2X#FU_( .5=B3JVY"+D%>]?#5%OM?AWU/RC!
P^N23*RT5IUEFNVZGU\Z+X>:%U@2_L"^/%@+M)T1.;.D6<)I_+PWX)]#A2>_2Z'P!
P[*9Q'PR7.5"*QD!<EO*IS-&-RIMC:MID-,E_TC#R>/ VYCV7"[^5T#0J5]]YZZ"T
P&HJ-AQQ&TL8P)"%'U=.92-H(@;H'/$A3(/%A#%++.BK0:J84_Q8@75)^*!1DJTQG
PR(\BQRD+)7YZ>BNM:QI(]-\P5XJU0O8]>*L)#Q_GZGIXRUI^)J&[XXE\E:Z<5PF=
P_&!_2J+U&=JR*MME9AX*GXH"_H8<<4=A<+#;4DY^H?#!]"6U?FCO^G4;T@ S:-V5
P!/4 K=.Z=SQR?M*X1P;E!]K7Z5U,F9LHHH9;T:M$P=65Q3(0PO5^4JPT8ADL6 B%
PC7MG0?C>T!@-XCD5U!X ^")D;EM'0G8V5;:BH&4JC9;/Y([,A?3"H;7^$/@7N1YB
PRB,U:?23^3S4L%)'+82[PUXIR3T?.ETCV18S_BO 9UQ$*P]:'_"^YI8VV'USN5.U
P3^-Q6)@KW;M>U%:W2LMD<_J>S=UZ2:EQDQ7_M;94UK'"/B^+&X>C\9R/:L^OQZP.
P%G<$]7_>MD&HRTH2<]PLJ+NS[*5U] T#[#]/_*%XF30E'E,#O_-9FPH%A@8;=$GG
P.G,.C\HGRT5E8V+.;"ZXP<>7&#\4_$.E#:'PTU+GMH1.K+^MA*]D@4."(VIN^]28
P=5+W&++E7P042)!H4GY;$V<\0DR"'UH$Q6P)WP4*)>[Z.(\N1C)-X*73F>[U6>O4
P.%..4-O_TX=S:M*4&WK15)T#VPY1-<N3!ZK\K.@[+>*O5%KN:E)UC)AS!YP@[+0+
PU7KLS?0(8JYS?&,J%B[3(CUZZ1*4S\**1K7P[<HR<B 4@4X/ICBL<)LQ%(V!3+H[
PG1:G\C0 J:2M0SL%B61^9K; ]"^S3?+4MS/F3^P7UDC%QYT<C+V0%@E-<K_ >H)J
P @$NJ";1@Y%1*,MT2!=J1^D]#;]B7G-BFN==?]AI*"28FIN!^UP+VHF #%T988G?
PT%EA8VAF!EH"GWM6-('"L*)&8+PR/JFAUD;WP.\J'+Z3_OSNZ!.>$I^* X$<WP;;
PN .RZ_J6>PCI/&_AF&SLXZ?*MI&U^H,MX?->@GAO&L6U.]_3&VWN_<R^KS3E5MBK
P(> ]NI.?BT(L!]RI)A#8L&U^#RI MNKKLFLO%I #=Q[.]4<<!S0L=O9A!:+!]=KE
PU>"*VNN!-LEZY&R27>NV\P$%&JP9)(2V (S#WK2'));QZU"T0%]/>:*BHZ5Q"ST(
P;KO69QRUBN3ZDQK1BBEK07XT2RJJBI(LT1A^>XHJY,K[@W%_K^Y.'E?UY?)S*> J
PT0P9LH:8GOM=_4&JG@%P>9,<Y378U(=I0!LZ)"X?'DK?[?LU!']U1'<8T+> *>&B
PDX-* :H01GE[IKDDC3JJ+?@=W%*U/_GZ"'+A5+XCZ[_[\:E<G5Z_XJ<110\K@I@$
PMMT1UEH/>X ^O%NYYDF$ <3*$MH7^N5FMO-1/*P-_R.<LXEBG&/CZE*4*QF:NVD0
P_Y_?L'-2R%+.NM OS7XK="]B:]//\/I,%'%@.[ -)82$J7]N\0AHSIP<[@<VI$'/
P[:E*+"!N(PDPYZ#6/_.UZ:N"^FZ&985   B4HN@J;$ZA'=1>2IY"O'PC*:&<R%QR
PZ2_=I@A[,"A\P>K"F4#3[QS'2U6+YU<QG<E:.^]R\$,U&E)HB0]3MI>)X6%(&D-'
PM[T%/@<W=MJ"3U6<O*1EB2KZNP$T*=TDU80;FI:FI=M"9*ZA:>ZV]]%HP5,RLD_(
PUQ?E%H;]T/7Z8F@+:;X'WW.G)-S_?(AT=6E<)O%\C.SLI1!(H"$RKZ10KN)F6WU.
PXV4QHT=[,KDJY*8: 5$>XQ[R@[UE70,5"7IU8W(V/'N)A0.UQRP,Y3(JD!2[.>@Q
PM<:(JE.EP4P6>G\NGW+.TB>OEV-%'?' L?]=U!F@MQU^D."*[5=6)-4$1"69RJD/
P,PW@IN-O90NTLV780T^#9V0<= [ZA;=7W*:F&P%$)]ZJ2]E,J[["GWQGH7'/EH3R
P5Y*(Q<5'XEJE"R?#18>H@K,9PBUS]Z#U&'&\\K9Q+W<><85=(ML4AITZ2S9L6BV2
P"JJH[J629]3NJU2\$%PU_CM]_ES=W.!@V8X@Q-VT^+EQ!TS+BVK>J]O[<IOFNL7D
PE.5GT<D&GA?"%U&O<!.+VU82 _#W=Z=\@G[!Z9\#0PM-X=O ]O:3Y^?YNX\E /2@
P[&%+K$[M"$BN-;ZA/Y+!U0]5CF#V</^;XZT4\!3[[2-#CQM;__=.LO@-HLL_=-O<
P1!^/!H:[,D?"Q<RZT*A=QW=Q9.RPE:2Y0& E<_DDRX(4_TA/+UR\U7=ZQHXLV$2[
P=D;]QR5"\@]\B?0H91I;IZ/Q;?R-H=<DPR)6\7XT_X6 [FLQ^TMW6N5,/02F5"".
P-92:#FOJBZ/GX7B3L8^H5X=3F0=HAMBX;6#F$LYYF>F5@ZTS.G@]#-94F9&H\Q%"
PD0H54PNC;5WEH1A^^"X^IVXCO&KQ?$0,?E0-43JX=Z\P/ID*@..7A'W@.+1"&6"Y
P"3C 6^D 'R%8;D2:S33=WO?6\J;N+6A2+(,L/2$)O-@D:Q00JA A!J&%):Z'_&!6
PKMMJ,FH@3/SZ84-M"TR8Z'+H:%MKU_HQ*74 4B)F@4A5E;!SE "G+GD7 :(II911
PP8SAU6W8+ML5[O47!9NKU&C%1P0Y>!%$3!M:Z!YO/DC9Y0U%(+LKZ6V74/ 0R7Y&
P,)LP4.A1GD@29II&O;_OA6'$]2CZ?:5]Q1*FM:;Y##X%O]E]XLH]<OPS_L';_S3B
PG\AH=\?M,)5.OO>"MHH"AK@!@XY\]!9WA.T:$&67BSOX U%GN.I(JM7OA!+>;\F+
P"M(\I"W9[#[J-&I@(YL'1O.Z 8,TOM[Y%CI0IZNZ-CW<JR14P^#1L?(B%+(U>GA\
PP8:=>(?68+# <Y7FIV!<4V8<>X,M#O2J1(I1*/Y%-79ZD1ZC&9JI?ISX8(<.KY[.
PRA<[[]/<#[^!9GKW365;D8B%TO#8:'#P1:)1RGE HV-'4VYV@.-J'B9N%6^=%Z<L
P2RE*0\I#Z? )E8L_U5?E'U="]V]DWP_'8$MU> TFZ4YN+/"SNN/.J:Y34MAZ&7<\
P(W$U1C2 OA?J!*5RNN7@:*JU@+!<=04_N4P)R1W$K)BI/W0NH;>9Y3<PBIZB)^'2
PVS)R44WB2D>0N,WPVROX@%3_UUN+:D3T%15$I-,Y1S+ATK-'F2REQNN>/W+-@?P3
PV#\UC8#$)52]3N *"8G1+B_BU<^4X4O=_=,18Q:@5]Q)\/=SRDLUWU89%Z5&3=GZ
PJ9/!7@:".+];X1:%RU?5VNXXZ0Z@X,8(1.M9@L3_*!$I$WZ4>V0]EV';*O)3G%0S
P5)% 2/S8(#-F3V!AB<0SV*C&IR<VHS5Z8*>O,*SF6)(N#%"<=^U?6K5,_8T.@]6Q
PR89#Q/B3V^SI3L97&DLM9CDA;%-[0'X05(Q.*$%<3IJM(^2BAS7,H.A2DE\C\,;>
P.Y;17''W*8SRA=1B:UM0'C("O[]4AE\S@L]0@N!JY!A;?D+^3?*N>=FM]>L.K_1!
PE"#K B^F_PR'WX?TMU\=@K0UM'FL%C-00/EPG334YL6IYAF)K"D:?MBD^S2V)HJV
P28OD[:<TL_%76K-ZCW7BJ;64T+EB &>O\&ZRI6  :-!_?JC%FV8]R.B'#!9:M-[4
PXQH9[I!S-I27W6+C%Z*U9YXL-%H@NJ?T!.W)WP75G!,,/1+ UKWU8!\: LP=3YU 
PE??2<:A=>6LWG@QUOS-/X?:MQ+(F:FQ&;>5AA[W >YU_['IE(3SJKUL\YSQ4: _S
P06MGF4PW9DJ9'WD##%(A>?B&<4C&?>Y3_*2U9LWW( L<^M:>CT@#H^GL=4Z=!!QM
P3I_ZC?'!$U:R ;QK)N7QA2_?%:3FL$K^<+F+K[?H4WD4,76H$W))?(@=5?AC$?)E
P)];D<*I?F+*P:M6'W;B]>8NKP?:PU%XB[2+47.^66N]7*"=84C7//S#"G?#+5 L8
PS)NH)*>$Y:T/K5]2-6VJ^WHCA#N,3+.=Q-(EW%;&DK.@6 T71MK5\RM\F!Q?*8I(
P8?)L(N#0'. >A,VPGRA,QZNQ:"L:L'C"G "U=753WN6L^W5M+\]:O3E0??]2&:D 
P%)37P)?9_W"'P[M:Z77]0 G7LIN5U0PAX20#@6QC2^644YU8V-S(A+H^&'V$J/&Z
P+#LQ0C?L4>$? 0\YO\R/"N-Y!S6@["_ ?RS4Q-6DZJ[M $I^;,V^I!97/"W< RMN
P7T[+_A/5ODB+)Z(:@ZSWK/FW 7)J&E$BQE]B_38E7#I5(HNRUV^_''O I(9+U8(N
P?9Q7TC#YGXUIA7NIH%7;-YSM;,->94(PD-Z< .RXBR)!0DU<"_HQ^@RA8H*<5URA
P?A?_$/G7JY//%KCA) +[VTB'=91ML)/JO8((SA84OBE.]06#[<) T9J69C'7%T%N
PJ@MQA)<4T1*W6075S^RGYCC)#Q\ O5O-R!@Z85$1N-+N\4!D;)\ <&LPI0Z<QI4Q
P8:0,KL<^19N>Y]P>19]"S'4R4>=>QR):II0%"7)V(,WK7318//&F/-:P(@V8GAU'
P]B@B=X5Q+,X1$A5Z@C\,D8N<47'C>!&CVWL3"E">MI64]6A\>)W+QF&:MXH)A+NQ
PM'=(+#^0%'DO1-H6NRR=T&)F_ZL0;Y87-]C'E],L^VMY%<8 ,D1E/B3IG-;+Y/%R
PJ7;]1FC6J#I2?L=.Q(#I"FOZZ-Q,*TOZ8-W,$(MYM<LIZZR/XLEWM9T>1)4E@[04
P"SVFZF2\U.DB_J<>@-\'^O/0*0MR4_6Y5G C'3G(1^L=='Y=<66HUE#@C,3R%64*
P^J,PX"SJ7F"2R]\T*X8Q7A9FBPA0$#H$*-@SNB(J*W6,LK6)%<"EDE1"PB@G,.4C
PRUCD-R0+>&9]=FED5"G*-B*X//'QCOU4$Y(Z6XBW#M=':@EAA4YE0T(M=UKT,:WC
P<!H6BX]?XOVYXJ19D"4 E1WZV59K1VZK1;5HO=#=1G"X2WR,35&.B\M"COT$TG"Z
PN3X$B5A_@-K!]SSBTC[4%R3(RN"#)-HH&I5_K6TU(F'.TF5',=\Q(!)(B&+%<B2A
P[\A"%0)B^EW-0]JK9%\[U>CI=2PF&\W\,5WV'MCS98D1@Q#,%8MX5WH40T8CRV[F
PAXCBVO@9(-5T<O^$,M%^3FP"7.C]7[+S6'\/LTC^ 79M U;]J8$:4=2+%,5KXH^I
P'IBMCH:#* %C1NU;6QI[?N'>7!^Q48IB_S&MJ>(EOBH0EE@WG\GC67$D/+_6_D-N
P5CS<J2E+9"B!)>QQRD.P(6&YR_ /GZK"SE7YQIH>=\UI97"]GY;N]QKGG#KH2!(@
P:!$U;6TI&M<4F@\,?]J\06:8BI2KGW&</%:$5[P:X*N6?CE :TXV;_SG")1#MF]6
P'RU5FUJ%9#[Z'<,W7T+7X TL-#J.Z"<U.0UW\T:H]$>$TX;O?"PR5W9',+5FZ5/A
P?*@,>IE"-'_.E6V5G8>B^9-UD+=QM<X%:_6&]H)"RN_><@<)O/%MF+9ZW^@N)8K=
PQ(I-E/Z@$0NAM<],O]S1&+WMXK?W=:=:ZR76W'$+"Q@=V&H^U.BMUDCY]4CMC9D\
P^0HC:&:SW14S1)%I;S^GC#3G'_,4<PY.MA *@?X";J(__\1D(&GQ-)H_6P?Z;;0^
PY7N#M#I8!VSR^RMZI\_'T)E.(O[4"2]Q?I_VQ4&]#L5$"=G?2M2I?*'[1S>FIXNM
PED3#H_\FT5&$\5<N02JB.;EXG!H"JHYAXX*!KYLGR#RK=^E<DT@%-A9+"J <_OFY
P.JZH((-.U:7<2S :>4.&G.*R$1*OO)U T%"]]T%?Z1&Z$X?[72,/$H1<W0T.U(8Y
P"$,M,+B]!-+D['T@80[=SQ^U<CJREW_LJ')*[$B27VE_?[*8[G1T65>(GTH92D.X
PX__R@"5RJ;.<F-Y+!GUYX?]/^_XMLZZ<*&I* (:M3:;J7?DT8GLSZZW@VUS%8Q8I
PLS2$3[-^RH%XIW>D$LX@"4__GY,K7J\!K*"T,#6J*126@B&0QN0X;(%C578JU[H^
P(M6+>\]3PM\B-[BPDA+ #RE:_[#3QM$#&@/L7Y3"7#T((]KU!N5^2YZ"<]KVY_\3
PD%Y1+Y"^8=+*<7:NI6T:P14BC1_0CYRB:C]@,,6*>BBH;$E&%3\A(<2K>G.9G=!T
P96W5WWDXT!A;O@XD\4P->T&@4_?#@)WSXSG%\TBKW2/-ER2(;:@>Q?T>R%8PQ%U9
P2+=(S#BSZ< V/4<?B!I0+H5LR-0MNR4JIF-CF'LS]5Q2:\7O\G8EJ%;X^OE)7?Z0
P\R#!.X AE$->T0T ?73(C7=.*Y*3(0U!OQM+FQ,>MW%)>,$1H#PIH3&[%-&Y>U!+
PTCE<J7]29Z%:).(L?[X0%8M/GRQ85*W:/%4H-$]0]V*!$<\A7X6ZI CK$L#JY&(0
P'?Q >[[_->WUF=Q"WS_NYK=-]]>#RKI,MPZ30;7D8F620+/HX;T=Y*@8QQ=_S+P>
P_A4VTO>Z+]9&K]!8)K'I%O$?3:3$@[!B09#\QS.G(L#ZA]O5"S*4^<E0L%7?A*VU
P\^SY(5-54+@JMS# E_VHHAF8J)><4)(Z!0XI>5Y\B_R0-QIYR5KRJ&B#%^KHS5(]
PS6X31VCCF8,R(YP^S9C_!'.7!]_F>G?AV>URT1[IKOA9I0%0-AID>[?QISD0645E
P3[15P3P(B$OM%A Z[)L+9D@"(X(R\,S&W_7YSRF.L-&S^6:*KZOW7,).DH-+/6]2
P^IYR'98ZUV$T'N3P.UDD%LWPLL\\)$7G?9^\@'S:LJEI1?D*(A3Y1^&@3VK=N$6=
PQB,O?YR>FQQK_^D9X5] Q?&P+5X23=ZR7K)/&W9^-GU/LG:47GT*0+/(T0L%90PI
P727-Y^,:?#*%K;N"?TIAKE#?66B$D]09+60!KIU^MR,5/D;S\1Y/#$P"NTN;$TM^
P9TQ*8@^"X.(8I>A5S4=LB)[NX7ZU4B.6>P0\ N^3[2@.(8)"]0T?#X$-!6*MCA:\
P0H>^A,/_F^ "]B*/ K\DVMSW<.SZE%\L-XKRB^:/#D$_@M64H^453+(PJ$T'T023
P[)8:1^9FQQ_Z2IK(F:$$5A-;Z8F_7NF,U6>V< >V,RJI'?PPLD_=_VIBV"%_HA?B
P9BJ1=)'*[CK73S@)Z4\(?G_PZ/T-P$MK[D\JOM!](X#^2[J=BE8"KHEG5QPS4$!2
P.[%_?P3"%6TN8V39[O+ -+P"3?X)8UY&6OGMV':X+4+?:!IB=9X$'"W1[21,?TJ%
P+?9)FT[;O9FX4\AD'09J3OG]5G$&RVD$S IW*Z*<:/=1XN 5&6H24Z0M51GHZ#9;
PQ6TP I.I+VKG/&FK\,X[1CS?A$I1]18*XRF%#RP#'$7Y90>Z*1/W5?A!-B^=6X;"
PL(C2[H#-Q&;;'*5=,S'!R_&O6]ANC/DMT,JD.]D'!7\^+!6]"<2GDT:X,_X>8$+2
P\& U(_.3RP)4DS7-@-*G!AM7SQM*$J*8V%T-#=CQ<Q<'FE9)_USHW'F6$MQ?VUOR
PB^JEO\O)6,%3G-@0(2?<M))2<@ZK1</F.A7)L*R$>7^80A720>]3]083$&PH!_MP
PM4DI5L[G4=\2S16T/UBB+$11)N]8YL&XA;WBY>$HN]!]<6JN%W,"3SD_N&-I %<-
P?"O[+ O<>DZ>B-[H-,LK4$(;= K(M4=-"! L G3:H=C@Y2H?$ Q5@=P1[BTQ7KXM
PSIDT%3YZLP\;W24@.RJ$IW9ZCV!ILA<.\: !%Y*J=^6!'%&Z;E^()8\H*A>)M[YE
PW2=V:%3&T]#"NR6:(.;&3:GYI\OM(.O08"@!UVD+6FK58*.UX)8TS[%RS(V4FJ#B
PX;U#6H@33W4FCSD#4O3-NX!JH<1FS<3<;8*!1&<\'1)?@IH88E4DI$$8#!- !4+C
P[4R2DK)Y>*[0![3ZSNV^X6VR[''BF@*I\@6F*9UE'<+1UF++B>8#L1QDO8B]SJ1[
P3"CT$N^Y\)]^!G]AC8SN7_2*6)DL_!)!NY>+M6X)<AKW?2#-=F)I^V[O\P'"5R K
P^0A =5H\\BZN'C7JN2<DN#9347S"YAF#K#ZD6^4\ -8VK7PK'_ZA7[O5L"LT2M_!
PDM]#[1Q9[0L6+W[21%WP4H_-C620<]7H$&9WN^-R:6O=-0YQ3.[#)1*13@USFS_:
P"Y\=)LX>=1A<;DH;ZG,@8VX"3"_A^U"J18,/-H=DXVF!W&P^[>RZCKCV-Y<U(;J1
P,'/;>[(QAH1M"KP'-@H@0*.&>J#ZIMP')X^/%!ONAALGLUP:,"O_$C./T D@DW9=
P%5T9P#EA@;Z NGFTL[.?+V$5B,>T^'?/5L'7=.+0VS:->\EM,: HW)B$68)M>=\C
P#VK54Q$/&FC-8K/P4D^M>]U\S-:MCEZ^_3$4-I(>,% ^-'&O7:S1X]-SU6J.&-.Z
PYH.LG]U=)Z%9<:8-Z[13+T=,DBJ-AAO&L6 [O-FNY_B49H=B[,8)(&Q'>.PR@60I
PV("SB91#>M-2SA3.;Q;]^8D\X-8KW+2J=<9L4W[/5R=WAFT_^+8MSCT)!UKWX0TC
P?Z69+'5Q:=R:O(V[Y!S\%IU#V.!JB$"G_#&%.(4S,J,0*.B+B_%IF=&[O39NNLF^
P T?2/]H_.ZE6T]B,'#.XA)^+UG[CV&<?;+HKA?KZ'I!+L[<&N6?M-)T;,:@/ /G]
P=ILX;EXY)T.<)T^+]S#?)DV(S"VB:,2TKRLLANK:899C$G])9.,M!+23J(\2D, &
P1@BCB'AYLEB4)B4+.]$#X4$H:73RJP:MJ42T#U0>@0'F!! .Y8W+06[N/%A6QPQF
P.X> E.?;%R+4Q:P(L-]&&99UNPI3A6,8_(]QK:#H3Z7CRU_S^8Z@B>;B36*'P3QU
P/^!5IU<&/DU(86W)W539PY]YH=U>4RL;?6ST36HK0XNW:SVQ;B4=&-:=KFET6L8,
PJ=>'LE(V1_C3N:&/P82!J@6(;PCS\"[Q:%&7KG43%FKR\Y\,*#O/@3[V2E6]C$EJ
P+*3ZO=*(O)M7C(CF=Z)7L8(3K.@XL9^4"?/C-"ZW7.28)!Q/UL=#R#E[^520S&"-
P>,;(P%4K8/DD6/19X+1HNR"[2A[[J$PR6HFQU@JGZ;:;P&7.'/+JK6*<HS8 =?VV
PL$@ZX3,E$KPIW33AOO*GQHS'YHN0JRVH[L#\8$55KSS)8^'\6FA* 9,&PX@=?0!'
PZ]7VU%\W-\X)LBM( Z_F\]10=B]DLL:PJAYLL!(3,-T"7\?^+ 9#<LDR_(=!L>'4
P.Q<68SQ0&BV=M . ]CA;#>9"!]2:Z8_D#KK:T=N7FYHM [WQUE [D,<*W9^!\@&*
P)]=!3/<FTQ^.E0^UBRP-)6:T"]#TC*2UO+)!9G8$V8JS0V@;O)=S^%!E.D!N3[H3
P++O"./>JR#F?WU 0%09=QL1P8OQ+Q8,%K 02;! [(,/!+](/-&.(N$N4OT-K+.G%
PHB/ I9^,_OF!6<\*5'--:J8++]<;.F8H6J,[53\(@1:4"I E6\.KA(:']P6+C"\<
PUW.5+O/]))HJ>&+@\R.J6(#C WWGJ06)2!?%FMEV1DSOJC 8O1+IOLC,O-OT _ 6
PS>[-#7O\4-HAJ6W#0'@;1["?J8HL,--27F13^'&7(IK<?T"KL*NV'0A3J%2!\7_'
P=T6VT^Y]OQ)Z@.YX6D:G<VAD3V4@@5N!,NQQ3!3JO),TU>=89;PWQ2$2S95=BTSH
PL>D%$7((8B^@'>*8WZ'M=_13.)I:A5]I:*54<;W4R57"1B4%_7M "#-,J#0M,X+Q
P'OQ8049W0,,@;^I-EZ2O3VT24!+^X:.$<H=+?M)&ODUD1P_X.SW3H%0SMFIJ,G:%
P*@<0LM&?+G QO?YVWC']4>E)1MAE+_]J<^ JC^I ,I&3/#>W7W+V2D@&SI@$R7Q&
P._PZS4I/]IL-,4]8>7=##Y?<8RFEA!M'X)_0-=K9Z7=+ZGE@@<0]B]9$;74/1MTK
P:?%5:8)V@0'DN[6)NJ:S[F$Z7#9N-OLFP%PE(C?&M/$\9%L9C19]2V7@J(3!\J.5
P*1^&YHM6/;H#Z]_%95BZB;@S:T$RHXHSDG_J*-,=GNA%R".\NZW([R.?4)"#W2+R
P4>'5;9V$H=:1V\175D 0Q-_/QPE!)J,##>%O-'0?.1S84>LJ#!OX-[D?FTDX?Z:0
POJ[]%O<R#[ID=CV03"CSV);25Z@8A[25!KUCQC7!,B&$H#5[;QE? DZ>$"1-P *U
P&IY;Q>@5X_^OHCI728N;;2%A8(U[7E3."?570;1\7&\$6)6R+[T*[T#A?F F=2Q$
PDE"51M=THU..Q@_5_,!)[LWJ>$;PI)(F< L7.*?"*S$HVG%,'(C\^(UA&D(JC<N6
PH2\NE1V^X@?WQ,G^I[\27-G*=A(9?1Y(( 2[327TP*ZM93HP8J?>2GZGSV:'5D\O
PN=:D(XO].%:-/BC>D$FJL4JO_5SDR[VMK=I5..NGCN"T2$:3A=L3*V841Y\"=H<<
PW%%:P*CEI>^+7I=O=>@3:ARB5[HAZW4$>QVOB2R]M_A*/;\GD:T%ZG%A6H" R[FS
PT^*$$ADH_<2DNF!DX)=6/-4ESQH;PI.$;>B<>O_^P\]@:K%(LQ6LN9",D.N\TH?B
P],B2E<O*^<+OFZ4MMI6MC^_'IYZG\1C1> 5OXLV)O?)%%X:.XO *1ER<)S<5I2 7
P>"J]^9J]A80J.C99YDP0899*BKR#'(@WF?1(UPC[SUX%:-2\+8^H]\ V\G[]V)?+
P$>%<F7@TIYJ@&8NHU[YBFR,0-7@9QL9A\HT+Q <82<0?&H*W+ %SSP#3@[ZNNI:-
P'"N28=YU*6(Y@ZG=.$;;[PB5^Q1NB@+) ZG]<$SY:$@D_93..0\WJ52RSK:TC*7R
P^,>)]/.$4 R7W4:RT64^>OTR@QJ')=YDW$G&6PK6#ALF-F.9!M _K$PKWQ25N<!J
PPHS*2*;83X];/*JL7*33U$%'OWP3X@\<A/]8V!V9J.X?:4#VJ(MVA^I=XBX[IO[<
P;OD[I:P66_OR**R1^D^H/7ST'HG?SQ,<4/O;X8,AXAC+^YEU:]-9FE75VG:A\;($
P9#ORV+[60GA:U*^GJM!B1TD&C\"_5+ ,#7S6.G_WI.X(AF&%ZQ[V)ME5HI!U)=4K
P])M'FX"0VR=?C.;J3EY0.9;2:9#2]#)[?W(2*L07 ")=HM<#S^+71@5-Q !(..VV
P8%] K%]LD?O^^"AS KUWLJI#U,KF1QS'4"B[F;[&&+SB>:PI:TC5>;&_DEKU&(7$
P[&&9-2D"^2IM/-B"W/3 G3\.P/!Z)PB'ZW(#(E?BN@RAA^-1CXYAY"=4/'0-.JC$
P[FL.57"=6%,67Q;'&_@U6"4* _NO5T<M!F,OB>&><[GYDYN7I;LBTS,MY$(/B#5P
P45O8%$TFEE0PZ\C, O\IY.C'(I:,!WYY:EQ-UKOJT>UY^@Q%?,M6(J+77/+!!3FV
P@Z3V>LU=%G-QH:UH8\'@M??QQ(:[/=4'$C>#>W9"Z7^W7#_9O)DM^K(-N\=P^O-9
PR0#&?&(K?JVQJ'O6&'_,B'>HY)/'001.RWA)G%:FDA73 U(WY*!#Z!5ND@D<!'<)
PW6J/<OU_7:D#'@S(F)(- @*9T*YC.Y]L]$[419KJ],AMEP0]VE3QA.F(0>N-(-!*
P=W$T?ML$S('TVNZNE+1_NUSG?3(&1O..<NK!2(=[WV8IWWJT(^SP&P3,EQ&A-@)[
PF>"EB0!9$8$,2Z8&+<5M"HS:5ZGV5"2RY=-_G34U=ZBULE^BHT*UOMS<'BZ[5M>&
P7-V6X6ANX7[N^QHKG3+@/!T@V:X\<$9O'O$X1ME^DI?E:IK3@9E+0M0; #KI"54M
P+-&\#UZ[BE+_>9I'-SJ6WWWU;TP$3\NXIYRH0VRF I 2A.M-M/'6!H_D'SL?4"G=
P"_Z@3$L59>4"4*:6OB_HA3GZ.&Z9(/WY/$)A5'TJM7\8"5_@G8:\H""P/RLB14 3
P,]=:\Y4'99#%33ROI',C($; J&<M"<=_V'UK?GE6N * 5SQ!XFFS0$NLA(-] E!>
P:F49/[%6P!QBM,OL<(BQ_$J_!)4>0OB7JYN09=2M4Y&N0G%L%!AB'-GS;WU?95G,
P$N>3K*0RC(5T+:Q;<^U62'W^.HGT%"!42.]*M$C.ZYN&MG4+A-C7?,'2R(1X+<-1
P%K*FB?6)26RFQ <%(%.[]&.Z*?2?JRO02/]:D]M3_N!ZA,6468X[,9HYN[J<F/ZG
P_X0QL'$&O&U .'V#:;)+5LG[2-$.<FUUSL(F-OQ1T;-;\4F=R=)AIJ9!SD^+'RS,
PMIYE+@>X<XYENT^GKFE<.EV;[@IKL-[ 2?O9X#^<=;>JHD-F%(=@K#7RZ)7K\-[I
PO]9O3#DK/;. "!0?7-_M4DP0=U/GT:#MIWKCA)9)E]OD_*N)XT[A@V&2#.4M_\L^
PS_#F5W1U/M>L*6V1-+C52&9I6(]N/(""H1^F=I3,O756MEW=N-;)?F@7/G:-.MJ:
P&C";B,T1F3[F(TR<2Q_5HW*?%A-E]>P.>0U\6K<3BE#P; ./''= G2 +H#N\]\PM
PM3H +6:Q;&)OX^4)'2E,#YO1)%[X!S"C1#]HA</(6;>5;T&,?IA?YW0F;Z]-GV1U
PC]Y\,!8('>4<"(8#M^FI1YP^:L:=+(ZTZ6\9QD ]S)?^KB]/4+ Y]65=99@YH/Q:
P;PN6+K?Y.GB)8EC=@0MTT@FZ..A W+IQ"LZR9.9,+/.M&^@2R*O#$/;IR""/,I53
PV./M+!%!H@8EH9)'Q:!C!I83)==GNU':/PZ_:_MF#8UDM\5B'<=I7]6@B-L#5+8T
P.3B]SCGGNA<OO3Q!>Y$_14 :]Z2ENOSB85WQA=C_=_,#<EMM%BP?#FSGQ31-&*1]
P+3_$$-$L.9@&98]%6*!^A ;BR2@ZO1?[6!)[\ /[08'(Z+:0Z'\VESREZ[#0*2]8
P)'/3Y(WP)XU-KG<>I\.L/A6D<2BK!B\<D-B5&)\2\)F/W[HD!%/(=K ]WT6@ZXXD
P8:\G:;^SH-GP8!.>F8B@@4'I8R@&E00$ZD'P6M%+G7C/S0&OIFVNZN;"J[>%.#!@
P+^GD(F6GS(4?;N:%S%C2ARY^953"^XB ?609=^?+QIK6+*VYB&*S&4V&PGRN,4AQ
P\;_&W+/YHV37]]#5E2!.\^[$<2,,B+BF<BM=$#9\FWQ:7# WI+R?^*YR^B:MBWB>
PU.?^T4<QZIW@C@=%T%R=*HM(ML8?0V'FA/3@6J&N:V.[[\Q'@ME:4<SFB^9*1P =
PQ+GZ/"7!=+IJA87$Q/I$)&2U*-?<[6=Y0SBOS>\*93I,%GD"=E\I*(PR9H5L7=A=
P&HX.WVQ;)??8VB\^^5)N Z:WW:EZT"V]TV9")Z=C.+4*!L_?'A"6Y8X4\;+PGMW 
P<.AKA:RA$#,WVQTR,"!<,+=W[NI,?^IUB)^M^..CE3-\S_8[L6:[LA"9-U;@K;*7
P\G8UTO5]=()%C+MP]RRE;@]EV]W\!5C"6X%<X5QZ* ZY_6=$>J+)&J85.^-)DHGM
PU3"F ?@."#;K5M2I==$;FLC9P(.71X#0YCB6?$OH9[WT-2*</PFP0+'_8)49$9$2
P_]@^=V9B7?H:B]4[ESB,[C"NN]$(CI(:<X/65$?"PWA7Z_&G1PQY*L.6>JQBWB.-
PL-G(^*OYUDULR5WZKLQ861< S'&^5JO2SG8M:Z@^5HPU+M(8S1?A.<R>9,"%\LIZ
P=D*9\!$*?6$@^9>)T#^E/#SM$?9?B_/XVVTP+G_=%40<Z'H8PCX/&[P_!S!SU1P,
PDD@XU?D"#K6'1H= "H,,JH:6!XXI#:+"07X#N[7F;55E2#,T=P>\\L44C9_9], D
P8,7.LM#R<C*6#^0'W)&%X']4YL*D%[_5<X%LZ=+"28YWM>MAK,X^K;."I(!<_7CT
PN$*>C(58O^ '&<HQQ(A0.'*X<5V,[$G&L[T2EJY^F8'2IM,#V&R+UOAAU.B%I A%
P8Z_@Q*J[TF-S%!)L;Z24G=&N<58T;$?S[4='#;^,(;2P*%FCOV^DLP[FI#(S^^#,
P,U5"3:Y:Q3/GQEL/)PT 96R_>HM<\G:P"4TAO]E,0@:]#:;_0MYEE6@WQ2=YFU!,
P#3A"B)"'#G]$!?TTJ,]_6/*O\CH['*1S"Y8=Q"6BZ_Q2=&:FV$I%GS%G2>QU6HNS
P;OJNO AX%LIH(&X949Z]><M,%C";.$0OXMS2R%<><D T >9&/U^"$[4#R&=?U^?>
P>]MN0!XAE6 )&8=<64!1;7>?)$;@O>IS#4J1(7(G3.;P,#&(D!Y'9).XV3$G79US
PM\(_98D=L=&:=&)I]E+N4#DQ"!49A4LUR8583K!,GN [LQ3WJ)Y5$J+FX(/GO.?5
P!ZN=Q[FN+Y&094J*C\JBP+_?<(B?M&WY[#8$>][,5:>Z)*LD_XX#T%5!= :Z>AS*
P6?6*VZ'FLV^9+W;)E1#_"5/)50JYO5SIMON.P;8T^X^PYA.O PE#E"=*%8<4L)1:
PB@KY._5+.;T-L;XKS;?Y(=V$&A_T@&E D@UH[0:EQZ2(I"0J1LM7=G1J]>3PHP6[
P%XL2DX6W/^ZY\4P0>;5QU<C%<:EP'1]QAX%+U#:8A/9QM)B\$#]-CFAWH=PG..OT
PLTAA$5WW^9DR)['F?DXZMC]=0\- 5+EVH4XMH@PY^R\K"<P/E=/$JAM4X7O;=A!2
P)@^(>!&8Y1CQQ/H9P+1@=I]( \*:)7M6K):+K/<?BOT%443_5@0EU6KU='Y<+ZIQ
PF?&_E?2*M,S3H)<\R,]I-&6Y+^ARZ=R>T:'3KHM_*:#%:LA3;Y4;45D3<RE+/+P_
PR*K&Q?SB23%ELX^:>5O O91./9XE9+*FEZOD49MWR-;C?@SNZ/3)$S3O/X/MB]!$
P_H6LP1W&D//UPE[;LN=0[J]PET[SVUD6Z67-FR6V:$$>[@3G ),;$\R.4+I\$[+]
PH9%886?< =H)MF'T K:B*1U@A_Y-O"HNX8U],[@Y8LRYV8U/<6;7*TX:1*WW]4IN
P69C-[K2RJ:?13C">U@ZYP6 0F[*\]MM530A,VSZ<WSWR<]O;&9_Y#WNR5N^<K$Q#
P=..Y/;;H$5U4T?RO<<03)<^"7*3K[E@[XM$PYS!IJ2801Z#W0_$17*,( [U9(0,*
PSP):72W:OC16<QXX[G*GRJM/+"Z1,PM(J:DW-P-'+:Q.Q.,N<%4+/V7Q I1S@2X=
P&5%V$%;4DW$]WYV5K!,*@>05WY:5GD+RG[5+QV.\\.M*;/K^^)M8"="[_7R@.Z$#
P"WDS "6Q89O97<R7G&+9TTUI0!#$'@@426'9B/M[5<L6N5]N1&(.-LDPFQTU$$&4
P(Y=_?+-I#QFP(S!E?]1HXI5ZR2%R *-N>K0 K<IE:%%LO+W@17AV4:?S ZBONC1,
P48;P)NQ1/C!$HW 5?^XETBA3Z1U#X5+&@;=#*.9CJR<P0R_2JQ*48G_EJ%R0OIJ+
P&DW^?V7MZI95I6\W-USBM$; I=L?&+71D9V?9*AK!.'/O0=/=CLUL!:NC\B*L3J<
P=E@9]MQ9/'9"4&G++#4+,*K26%4R<Q(A=;<EY"A9VY+2KI6EVHONS/>E-QW>PRX-
PN-*P8QY,]U#+]7D6>KP]B_FP8R1L3*C2DX#O99^<?[/\L1O,*W>1T-' Y@,-^EI1
P"@$@?7/:Q0<V 8[M.Q6>[ZW._7#^ND+?X/E_-<]9/!M5']I@0I&%=OB]V'CC<5M%
PX%+]+RR=[CT0^J#WDO3KT8F.3&G ^O#E)RB#;&>%2,=O4J6/U6+L>D[R; +$*]5C
P!6UR!%,LEXEL?7'_M---\C/1=!X?"C")M^60C*&RZ]JF:[>NX"\ZN6A]/&J(>&54
P/S]:8RI,.["GC86%'DRG]S8WSA@[70RF24$$P*;M-:'](*]ZS@+.ZJ40- ID;(.-
P I'?)G'Z%VRO*PA(JJG)491VQ;@4.X-X(JQ.,C35C%XH+;.O=06_._=5&'H[,>>"
P+F.4LD^=T[V[I0=PFIN,U3:%<F'"5/0Y.-^R@>DOZVZ7JH<4R&IYTJBK[X%R'$.I
P#W,XG3HRLB5L 4WA)KOF2FLW!H,!O)M[/<QN?X[[E+=42A:[8JFC\@J'D@1)R+'Q
P$V&%N.)6>'J.0AD^R]'?;F(Z914RM!ET7L;5,?7FFQP<ZST59? 3 83?]PD%DYMQ
P!9T#D(L]RAV7]TY5) W\!")8WY0B67CKN415Q[P]T4V"DJ=:&?C#^:E8ZK[TU-_Y
PNM&P9O^CPWXF;<:9;0V@) O? UEQ1QY8W\W 7@0B"BQ."LH*-U"^N(QY%<=QD1!>
PM#P F1(.$!Q=[V0[72=.<6D5:OSA_3,96E'M;YO+#IK?VG(,Y/W?<63DJ[86@4F^
P4$=W\74D;F3""8WX#525CJ@W4/C$<H9L=Q$8XJ\M!GE\PIEH4.!A.;F9WX_7L66B
P,2,F) 69XSON)?LA>0@(_8V(X(S*89>%UGB93[T_!"$=3^(N K#H$_&_D<B:K\)I
P*5?&!:UXZO[YG3.9Z)LYA31 6EB5-"C+*(E1X<5]KTP.,2\B*!Q!1YF76@,Y@M,2
P<=3""(Q;[QWM/Q:"'9#8G.RTPI3CI0OS#4[.ZC.3DP.XJVPYKQFM(FX)HAAWO ,H
P#8BRT':;F=1=3_/KEM;!$!+ :[MHAP_!E'0@+CC3@<X%.WK<NMSEQ9 H]O\HPAX]
PLCJV>">5+>-KG5Y3AC@G9(;$,,LL8'GZ3_% ')-C[DZ):0J,C\7RA!W2+C-PYX52
P*I4B#:(K'F-X^@5U[7T'D3(TWO]_D6QYE7F@,@EY2$9JO69TN,.U5>0UH>&48NF.
PBO4^2E2#S!I5IM"SIY%R%09?,"Q8;SRCNZ\4?^#AI:J@B'"37KF>HQH64Y*?#+UJ
PR]G6489"L)\6AFIZ;X=EULLK,3>')2CMIIE9 (#X0Y:M%7J35T ,I?OX8T/!?&S8
P_9T.TY(<F\C2M5F+574V]6"#RK899H>!D$X5^?) [!>4E$A=X'\VA_;Y&#T_<?G(
PU!Z=X(<Y4068'=@\SVC_'+=\XQ@D? 6T"T:> _,YK)]\ ?@=LV$W"FXG(#4(_N_M
P/W_1L8O=_M$HBH(Q5SA923)!9Z?9S[RRE:0<\!847M4V." +H'A026;!10O%XLN#
PX5=28I1S G3<[ES@QKYUZW[/35=7:]:<Y9O3P-!M4HP'F=(0D9O"2R A8[2CO,UY
P4')G4V2X0[*5AV@4!A;USA7F(G).7K:S<O'^&5^C:R(<=GQE>I4NMUY\+Q0E/#X"
P5(O\ZQZQ#6?CO' _S&-=>H%K6DU/2>O."$Z]LFH>"O ,3UQ6AQ&26/X0GCH\_!=H
PO:3"9&',V,%/9+-",ZJGN0;\9:CU!!Z$>42L)IW!YOOR<6L221AU@'='VR>X45T'
P1&OLK;\$ZG.'_#3T"HO-V7M,T>G/JK(M5)M*<79H/ IDD2<*2/"2/JY8@<TAA,.A
P@T+!..>KI$O<J6I9.1L*$QL/[L>N!:8_D@%022_1V&RV!ZUM%;*]\B+E@ R-E>$Y
P5K9I3O2%[_\&FC*M;N>3\O\A\DYFT*@;[54 DBGH!;7AI'R%@'\-A#J/=]&+-YC%
P#N<"Q]EK+"LJ'N=RRRV# 5@? ZX[324LX/^O\ZYX" ]/DF=:7A)12@IW*6<H/BA<
PN6D?=48SZ5#+1JUC0L&32]OQU1H#B2ZRTX@&_)Y @GN#)L1R39V3+STLZ'4;8Q2W
P\% 9LM(VG$?"4V.BIJ*2RC:RJ:J9^TZS\HL44!T!STCE+C$SB5[=J8*59>4-KP H
PE.(\)VMR@%WGK,OCQEH&3GZ3V%Z@U(\K6EJRO#Z2/W<0!C;FRFL"9!+5Z"_X@]6$
P$M[Y)V#QD$8B +6>RD2S7I"9#0:A)$$5L<'4^JO>OHO-PNDF5<I#GCD_"SB=C9\5
PD3]CHHD"UOE26BS6R8,,JRK(RVFOB;+&)F:R.W#:0B>8Y\3M.*/UT2>#4SF"I24L
P*_C[72<\M:"#\MAW.6TPX7@DE?*-]T@D240%F);$ 1V)_>=UM("LCGSV)?:D&'(H
PT1<*&Z:^G]?3CX:\2-[.?!:6 7!52(:N7A.';FYAZH(I @SRM&/#=P@[^?UXCC _
PLKTR,J+]>4Y]YQ#)OQ$-L1F1!#>WPN#F)G6< ^VS<>3O,P\#^:R1=9(M2U7%]K(Z
PT\&GZ%2]S>["G!?6Q1DL7">,\ADW%3Y)'M\T>*$CI9I_E/G-@FRS%(H5Z435.#GF
P=I#^FNOWXW2:B]M2B=YY=C>E,2V]&.F_/XLONP>5YTZIQN<XA:V*E_P!$"\UQAU;
P:V?4/8!].GK+#8Z@"BH@7)T#62FAF*,#.JNR]XU_C3, 8>\4 ]FLS$#=!E>%7K'%
PY;R+K4X8-YMN0+3=C/7\/0N-8CGQSI:D/G^UE]D=D._)%S,-K7I3%D3$\'/?JGN%
PR^UNTAB.#UN*SN61*PKOMNP4S1B$E7"- X^*-$:(HV@B,: PG <SW4E08I,1D3 B
PD>*>Y%(&-$V(EZ)J-P4QS8GD/XO^Y, J.L:*3:7*2*MF(48B?-4X,@&9G!X7U8- 
P?"A0:BKP(_W>_8HG<K>]Q*#[BL"NX_F <SW>].+,U&+$"I(URDH/HME>5GTPT>7-
P-YS\/F2F)+W8JX=7_BN&F-DH484*6\\^F3=)!$[.RI-S2%86[;<(BM<.LVU!7SUA
P9M*C2-,'CM/OQWO<?%1,0&^-Q,]H!0-#,N@/IC=/(WR7!8ZE2-I<),_"CT)S7E8[
P-WT4E5P-.PN.JWK9A5JC0JZQ>TK=-BJ*NV$N&Q[NO]XMHZD0&12_W;UX6KKFJL@A
PP<$Q1_J,O0(E]M[KZX"[VHD<AH- S)4NK%_=]9(+W)/E+!@A>#O2?FW)5+$][<6B
PC5E7*8V- X1=5O9;3;2.@5P*(X'MZ7??)=0LCKA5-51K4D),=8279J%JJ+$24WM)
PQU- @GLE3N ;[L+$D*7T0HGRV&'.HB-!X7QYF<TV?,17UX2: X@1LVKN0'3=04.9
PXF<ELM_]W\<)/ZLB^%#;3&C/3-_$J7X=T_N']'&&&>01]@[N00.=*S\#*3%@<W^Z
P^GN&5I]R ^NMK"JD%/!_R'Z]X,@T%"WZ?36D@UC'68"TI9>F@-_8>[?B:"<0#$&A
P=#I,GD9L]^G)WQ0+PZF$?J%DU'[ODOMR$97#W(D$83J$ 6LW9_!N0!4FXV;K+(7F
PO::V#D7)9;"D?[)=EGXYW231M/U(7O<B7]<,_^=*9^^0%SI!/X0MM;.F[D1P5<[?
PU0W3JQ%G.,"*.KJ4F+23]")EV;_>X^C+B3%V#C1@WI18<I'.&SQ]Y<(;+#5WQ3JX
P\;\_.Z]3-BXDZ1O 7^83A$06*7C?5"?5@ KC"'.HQ_]RW"^F(N!\X4=:G"'A/,,5
P%(WRV\UG>)5S]-4-Z6/TK-5H*R,6[,JGX]PX/YL6B:.6*C")N*4\VR)(XSZ\T(CY
P(@Y0%SGK+97*]Q+OF&&Y2B#D^!](&L^/#PRY#D,/U&3 _\58L5 ;99.QO=X-,G@0
PZP.?G1!)YA>KZ!9;20'7S+9J0%9L3N:TGM,@T:LN<0<:7KG@XT=>B=KZ_BJXYIT.
P^N_2,*_>8>ZZ'@XP>:PND3@%9KB*/"_,8*H7C_-X'\&UV:'_I'14THJ*<@N1348T
PI3'%U8@ IZ8,1%7-$E6VA5SN#"9(V&. GS50X4&O4_[/)9?)!W(IK$UNX$?DV>Q2
P=I&97T?=WC?X%F!)&"&_B 770U+C&<8_#VUY4>FJM&S*"6-@-@OFI9/N&(-YQR!(
P\[&??S 6F5AFLHE'EC+@W @J9%/!L(X6"PB4C\OY>E[SZ\Q141-IXD?61!G,1)V'
P<'I(X]6MX7RDX!9%").BNYDI (H_5M56P=ZMXL:2[O'>7EQK$:=( 5S";LC=X!DF
P;T"PT?C3G7L[R/KN+QT#MO>DC10R4TWX T?VKEZ>MN^SY3:(G%@1YT-,49;/R@Q&
P<_M,^9.\K9Y-;G3 XCV3LR']H[L3M'EU&"P9W(_)K_C]28XB4J7"TG#8L6:@,'U'
PWWBYRNG];UD:ZVTE?FFO<]ZR$4!&*&J_F]EIXN&[H=E=>TJ$O,KB#&[G'XH^K%Z1
PR.G9^#/CW'0K:@@WL11ZXXYY60VLP[XPU^ 'SR@3(G;-%B9XFR_P3,(9%#NQ^ITF
PX>(O^'FFKQ>G<@C0 >(A6,K9L.EN!SEAR+<.2%!;? X1%*<$?1'._(3@AG@AUX\>
P!]-B?_8NI5]>UDW@L6>MOUH@J-KW]P?.H+H+:G+CHJ_"'!=$^H)@7-.(GKY>#<%-
P<[:2UEWKP>JB[65K 0RP )%<! FN2QP# MT=P:ZI(N*K"2^K+^W4P%A!6Q7+B)U 
PH:F@6,-IE=:IH+N2I-LI7I/&U$3X.H,<K^8[E*AG>.^ #WY4LY-UG4N5?47R J/0
P\81883#<'Y)ND(J1.M7U(SL5)<(Y5N//'Z/@1_JO$A-N.*=6/;A_Y-F'5M>+SO?P
P+H>Z>*>H%1YE.3\"2'7O'(QLLW8%%UCH<ZD ))O=,L.61,7BC;@330 Y;)4=Y'3%
P:L')R/[NSDM:GB"\2F&A]T[[H+:5L !=;W09O%$Z['<&O\T-IUH\I^N*,HU%H%2C
PM1."<J3_HO@L!R^R"98HI]+994Z.XMP/MLX<>D"A;+/%29\7^#2]NQ\OEW,4B(#Z
P@[:=7=V3R:R# 1K3[1N@=)?M"M6V-3DQLX;* 7^?(QC0"%A[")9I;-/B:HJBIEXI
P$A%47+5"KDW]X' >MF9\Q=L; %9G4-179ZM]/X;O_6='9C96N9^*V' 1&?6?I+Q_
P=F7WS4J6R >:0<MXU8-B,NS%#"Y1RP]0D_HIRV75<DN90A%#(?>^/0$5Z\X#U^49
P:9[V;LO3?SOE]V*B" 35I:6VRT;+2;").^A?K893ZPLC>/+\G7@68'3'=K-H%[6<
PAIS7U8$J2'"+R$DP-7R$S,"'+3^0C\*]PF\([SQ WHE0.H>N9PRK'*E]BR9]!"]D
P5@6WVZ3?:<&4RT7_PVT([,\$X_I#O8L$+[<U%=M:#<]1T.&MG;."M_<X9[_-OR5?
P$!W-31/_M?1:*!D2K>7B<C'G><JM$N.EJ[G$NI93UV+/F@DB0MSJ+U+)C=>:G&!R
P [Q-3:T(!5'6F-G-TU=>/HH0 ](V=1>J.4+R./7%V]A[VEYZK$EC #E%W'V"'0E7
P2V9MSEOG947TJ$8A!HB!F-9AK_K%JX(Z%,^$MJ*GU^@$W(;5M?B]8HSDS[#MSPR8
PZ'J(QPCU7JMS%5I^(N%0/(3$'OK+(6U3:[4G3K^&!1..I<O2-L0V2/0HJE.[KVQL
P\I%D1[%T;YK&UZ^S70T]-JD 19@".K@(7[5DU <G0&RPVSE>HD6OEQ$5$B[WA4?:
PM*8SV:>?O3K30$'I[@T@P=0= UH%RBU<H,,WZ8Z"3)=N' C?T]&C$-+7_-*.."0?
P819I.C.6:)E#.26]/DZO>CN8 "X4$7Z_P'3<=5;"?329!IDD><MZX9\!I2PT7\#:
PBX*Y&H@AVL-)\21=F0 ]QZA=J>6#S#]WHZP4^[ZP$=XH]^\PII5$Q6.&V]XM*?+J
PX"(T<LI:S.^/8[6;^"Z%L8P.(-A[CDRWR>Y!]A;TOP4\K)L\M!6BXE>-M,;$=6V9
PD>HQP_-";;GW1&OBR3;(X@(J^$$=:HFZ2M5\)'#I5'7?U.2K'5+KQ $EY==(YIQ<
PSTH?U9$X2J)BW8"(<])FE'4T102\D!-G!C9ZOAG(1!8.+8N?PS)'=(8V#&;Y >SR
PB#+F,=3K3QVX<,9&CXH.=)-^/]43E@=YLO"JAA,I_CKVG/\3<*WOFZH;C%3)#D,^
P@RZY?JM/V]2V1/!ZUGMY01\%4N4MO!'IN')?KNZX&4:7>-VX%4_#_"BL?/9!4[=B
P7J@GBU$TXCEE(D$]$K=/@K>.8KZ"#+KV4UG^WL<'Z3*C(2@MTVP\9$F4<*K-3VOV
PE,CNU$:FLI,F_^=5/CGE]_O<9)SCVHYA+B?=9BX#">^#HI>"5#[=J\"%*RIFL2&C
PJBK\<^)YQ>*Q_T+8UOEG:<7\91?<5,FB5QR!>W9=._"5Q$6$QQG MT7ZL@IV.;IQ
P<OC""X$ [K%+BEB,/83;2?=<+!YKLQ_W;:+P\I1#*BYI4%U_!$/U)(N9CO@\P24+
P?*WLWV?**/4D%B#ZU>A#Q7F*7K5HN\T44_F]Z$;)N3(,\[H/EG!QV*B+*L<U[LMP
PIC)J-I.+=44ZT[Z8AQH96$!Z?L[4Y/3JZR3%XB'3C? ^HH'-QI3JD'@OWF"H"_'I
P;C)<J/&([0)#>>[&<5TMJ L7^I(5O06Y5EX[_9<Q.'U%EZN9WU_X"U?C0,H@^5!@
PV<H5PU_.DSD0!%6:YNUJ)[J*U&;:#62LQS-I3=.Y=RX_*H+%Y'\X.Y ><UE\TY+.
PK3)<C61;NO"H.V9*="W+ \B9 Z3QB%<-J'NI0"QHD,!W^EF:%RG3/9@'78HR+L?6
P,P^H#Q#&ZT,& \K2BBP[XP+A/H[I1]D\V'!)N,)A>9[5"#N+\R=USP!)O0XT7(?7
P-9(5#!^;Q@+$J^X?G&MBRUVG)-1?X6<+*JL8$HX,''G@!XDV622BNU%H-[[-EYL^
P'WNHVLB(P)2*2LVA&Y[D/4.A67LFJ/P$^C(;?ZP)PX1,N F"&:<%3 :J1AFI:HFO
PT-\?\T5_,I K9.>(4OQ\^R MQJQG$!:_F*D,6:K/0K6L7=OU5*VVL%2#]LLL5M>I
P^FNB[8"9-$F;R_#=]IYY##>_GGE5619B]\HJP'48(6KQ!H"^!,K2I+KU0T))#<4R
P&[/>A]@I_<&DJAGKV!P-LV?2@!/!JX'^5R,KKH+;V"G>@S'WJK?$?)F8D[E;#]@D
P8Z+XL(<L? I"5T:?BNE,*I $@[X$ZS[OS19()/?D@#[LFTK2J88IJ@JI5,4(IKM:
P(_G9<H;E^W#J:*<(/@8'.,MP$;K[;[ *)XZ,V&A(_*5UKHMRU9*?YF,/1ZH:<D,$
P6?+[(N_LRKS0#5;05XU,$<SMDLR@#8\-0D9=\QP]'0>?'<\3(#7_(QH7YZC\NE+$
PT& AU@"R!>-\7X%;-CXCXZ'6.+9P\*7X_^*#P_\IZ99A#%OX769R;;*7_U#9>7.H
PW\6VD?\ O1$-2LQ_0HK$@F]M4X%P:>8Z4JV"-2M$.1":.7@O1?<F$+HP^K[(N#Y<
PG2D;P_-GOVY?26O:^PA6G)L-J_)"DJ'/GMN6POFJ>['>MY6(+UN19"<-HXD>C$ED
P_XL$+E4&KD,"R';X!"B6GA_)/XC%?1O7YHCW\]K5#D?-T\V9AW_[]2;$NS1HI30$
PZ(',X14."8ZS\-9)BF[.X,_@+ ?TCX/B$XKW30!+3*>1*-]L9K851F/ES[T*0FO]
P&5>+7= "!T3B.CP>!C @'@BXP2R-H:N;4.7)^Z94T6IMV<$3X:MQ_0CYT'LBS;KI
P2[MX7"M]M<1LKD6<Q MRWZ4?N.&S[8L0./03>HM0.*5^P AC[]V6EC;-%V#D;^Y"
P)9P-O&R=R9A"N0=Z8C#7]CK4MPD+_.Z//491WJD.$LH%!EA#)+^49#(#M&?.=L]C
PV=SFT3YYGUQ2LBU:OJ@"LD?@452661U8.U)' )RTQX:-!6"23=YDC>NQ4S@$!SV1
P 175='#6QKR< A!3C,%,22[\CD$ZY<!<A;;Z2X_=T#4VD+WETH)W@>Y_!4KI?ZH8
PD[\5^\],[.[&0[V;4"9_1Z1+XH5.[T^=1PE$]:%#K]H_0T:)_[\Z+=A)"2Z-:5C@
P[0:#/?)>3\HJTQ?6CBTI[9;L;C_QXP*^^QA-2P>1=V2IWL-%D>XL&@+%>G![BW&+
PM9#:U.Y/R6T,T#F+,!>-.@N(B1"A=N *#J<3):J.\"D]]<<;4@IOM*_58,KBOVVQ
P=.ACB>H+&H=GHT#Z&) $'+5XVS2%N8UM,QB*_CV(1,E]I(3H%FG]K1;#J7G8F755
P,9:'5F[X[;]$FA<KJ-4;0(&+<@))/AL.IY+;,NO&N$R>%=Q&QMJ(3Q&_(1-%Z+ 9
PLVZ5L:*&U'.8CR0;#+U6K9@ %+<C_ D I:?XV-)S[6<*%4TOS WOST6SV5X!(R0E
P%8;?J+08-))PZ+"X,0$S3XB7R5R ,DQG _RF=WK+#O@(J]K0L*)BWEG;F2^6A.NK
P("RK&_/<B7%5)3,(KO6V;O#PO,4R<M'Y]3>_^6JF-M6<S!T"\?:JQ#[T%8] 1NT[
PJ/_0D:6J,3MCQ&6UP0XP0T0KS-797M[V\?8^S2L@ VG1&6_$9_*:"@1W]S"RY_&Q
PI/(.WF*Y$Q7PBW1J*QA:OIK5@_"9OZTN*/)>'44 ]JC4P7124[XF7*C<KW=M@VSX
P<TM:<1,1;.]AAT_!.'(G.*!*%2PI "RK0--?M;E_=.,Q9?\7N\?H.>I5B^(7KB&V
P)%2I )/],]$M#3&:D14*JH'!S/$XI@C_\OXES=]84EW];PILK=69OD$!ZO)=7D=S
P\K=[[7N,0>@TVU'JG=/8#SU%"?#D"PGCK5,'#I@6IQQ[4&I,*4ATJ0%E>W;.3GRP
P_\Y^U*?+5&@YY(+XB0V:P^!L#Y+H$^ J2(BDA"G^%<&$37#RV%!*"&"I0?YEFS(G
P^"4^5^EW_1Z?Z(6^_G$A Q4U*4A_EX<MVK<U.:@_20>Z-^!"FWJVU)T>><7(YSS%
P(9E+?GY?!=&!^6;L9P8BA-_W12$(FDQF.Z+K5%]AL0=73+W>K75E;2HD'Q3?<(U_
P^$<K5N"6\ FX8R.%HWJWLR@ .B2/E[?;"FD=Q8MZ3<()MU(89YS7)JC.7VO!@?;7
P6#*TX6C<#['3AH%?!'\F_YK3_'[8V*7@;VU0N!PH)#!Z ,,7.HTU"N>.>YS62(+H
P+P:>>X)QP1K#\JO@WI#W?9PP[<0G"Q=+,LKB*F,HI56S9JIT]@:],_)FQQ@(X832
P_U^@X[ =)NZ(Z;/2(%\6:&9\;N@T:HWJ*42J-!FYFP5-^B#&WF1D-/>T2J!<TAYM
PLWZ"_]NC*HS&$%SSP)/K?=3UE<H/OE7H\7JBQ;Z'Z]>+IV8CCM2,=W1Q. _2EC=&
P6V)A1.<)U@5B.HK6?58E(-<:8/L+>.R)GR7TG%3T,<2/ 5<9)PW]GPSU.P1],AKN
P&5<H_H[P],QO6IU*1<FR,1454@=X8_0GU")()FP2B):UVE"LBAZDOST6X)P<=%D7
P;-HA%.U*AS(?&O"1]$B&F[5LY\$.;+L(DX,8$<$9LT1#0=-6+N(=_K$ULW;-0@^@
P#X[NYK+KTAP"<IL4](6X@:%01FMT@P@HE!%[RJO#TKX7A/C19D'$Y7QN "EZ<0DU
P 6 \>O1F\BRW_;P'+TP[#5=N4!JPOKV30(EP]*IYBU9BL/"'APJM:JL7S(64!6,9
PFD?=$'EF&-O4G]8X3%L2@+M3D:3O,Y[&>HH(HXLC$6VNC2I*@J*+L/NX'RS_I N/
PXJB; I*^$7Q!RPIP%CV+0<Y*;HI&0#U2HYO1NC%V*NI4+=LKE/_NZ>^D5;+RZ(U&
PI@0DTO^5-HN#H$.SL/.MN.!I1 OYY/1'GN1_]SCI4T$,DCAF>1%9[IH/8G%P<9Q%
PBR$C_UW.@L073EU^:-B&D7LTC!!VH^UC!SK2]1XO_-8=9$D_);0-X,534S8]4Q=]
P?/:!UF,[0!+"GKOQD@##_B48ST^\FC&2/,0T!QUHT#!?W,=5D2"GLY>?'+Z!JFD-
P;]1LKK&MY(WGN3?50JH+SK$'#M P*LO8984?,VC@<:3$6:ALHQXL!F?SXU9PJQ2$
P[X$[%U_'",XNLS#,V_K>INQ9D.")V_5S'="2A6=&F, YB0_[")]4;KC);D+&/[0%
PE=OI2\JB(T]ZBU$C*<P@.O$I6& *0G!EL\RVX0 Y]>+-K);$J>T5Z%"KAO1%*L&R
PO]_-N(WF^]"E+DHF#KIQ567!#9;+KV741$::EB%( P7,#FDJ-+ O\HXAYQAH&DS;
P;W(?/',)K?EJYEJP[JTK]:3O(6>?;)]],;)K/-D'_C+.FC>U";; >_PX^RPC&2F%
P[<**Z/F>"Y(X)^,#@ *B L;MKO"\L%4ODJ/,'QP$5U$<M#IW/\MM+JJRQ],XQFP>
P!E7@DWX!<E2R?0[EN2G:!)( BXJE6USJ.I(&P!QF0E@D2Y\>:?0&& VD>SF:8--B
P;1<?#&YP1:/'68B'6?,Q1"4=-"[\MEF1\"!'_0,\XMSTXWN C%JN$6,(J1![=0_#
P">$:M0ZO-C?6][L0 );9WHLQ_M-! S32BY^W_TK)7" P\?65VZJW@."W<A-VE3K8
P3'-4V7Y*X 1PY/B*539ACK</8I<.<YP3P=FJ-I?P,8<:=>&:HP&34G]CXQ"_K+VZ
PUC;=T7T<_V2^*70R0[!R1AMD0DN?IR(CKM5I72GP72*+1)6,V0NJ!C'GYY14?XM@
PC%G#Y$U_PN596&/P'"H>8G-$_6_B;P0MEYY%%C YUVEWNFI13XIZ]*PB%,DT/G).
P@F&(UZN.IU4E+7 ES&[<#HXL.,8NDNC2GE6+W3ONQ\8?*%$(<"']3K.'-Q.'H['*
P64>>_)'K.O85V;I@;V"Z2X\ A*X:+=R#)AC4:I6D*41&-^1T:F_142> KR)#XP/6
P9."\ ;&H7"L" X0.Y@TSD@)V%U4?0W6P^*1Y8Q6>V\?437T*.^P!)]02!WA4L)/X
PD%O$_^N%=\])(^EMQ* QC%Y5CYX)#R^'<2!#W^Q[#%LP[).U#(?^[R;\0^OH#8KT
P1[569TV 7H\L<%VL*FI0^8T<G3]EJB89"72W=#'+67ID2ZV@_LI'RKS&SC2^-#1#
PPUVZ !H@RB/SQFP^\B)'^(8&0O@FF5IJ OF?LR%EE'L.H&ESA?K(;_@!EVXNV%).
PS";<('Z1E2<8O974.-,Z/CS)\V3+;-[: #!*X=-@ ]O"^T1/(.@Z_@KO=%^:7N*D
P3"+2\TF=DZKUZ5V50GNQONA/@NE?M/Y(['.;_9W/PD\O4I9J!ZU5"2V<.WP@[F*.
PC-DP09K,0XIT=71^2"X,!5YM0TO<"+@TI9B#^ACM>T\Z$>^3:W[A7U6PHD-]KS-+
P-0_) ?ZXMTGT?G.K049'P9'_#V0(C,])BLXA(S^6GI%?AB$<E75]MW9P4N1,97.J
P6D<.:%+$G<DZ8AQ[L>,A5,.)UDHN4%S/SX]QP;_7W"&L:P)I\.-_7 EXAW2I)N]C
P.GMZR^$59R[_C=!6H@"^4ZA@2P4J&"'QG^F,>!MP?7Y.Y!>A2P%*'F<86PR"Y4\=
P@7'4JK0"-@ P5!54V,]D( E0VIXR^\T<":D%U#VQT,,L;E2_M01DS2Z1INIBK5L0
PF";F96:D'_=-=&1CTYJI?R^;(/ZK%IT#V-39K%#?X@)B0OIS-@AC;"N,M9()\=5N
P,,O(+' K-@[L'_\']0E5_.,!?%0=!6#@\/R862ZW[*E$YJK6N3Q(VT%[TY)2(0@Y
PB@#JXQULKVDICWJ;F=IS[RBTK6T%&"V]596T_BZZB6.JQB*=(F*X9*U:/:(\P?6%
P,.-7!>G1_LDHU"1+ZE<0#V\77)A18BLXATC&A845S&A A>9J JVQ2+4B"%<ZU&OP
P, ^N9#5%2%';PXJ%@E@;23R^*._V%N:7K+;>;Z?,QT6Q"OPUKVHA[IE"WC19EPF-
PKW:E2+O8[T 1YUA&G*PE*SD@!G#57GLI1=U/&>!''%RM-3M06=\9HI_O ],P$:U=
P4X$3)W&]J"1,KVIL('7;_YV;9&5QBS6C/:!Z<_4(C/(GNTL*B;2@#OJN2YM"?U@=
P5;?MK:7Q'5<U9QR/':B_7]0<_.8:C["+V^Y,HW[3WV%T[+#*FE/Z8#TSR_6+;5AV
P>4?4,2Z.D!7B !6W*8-17RK\#9A\2&D.9P2FH*9$CC!%8.=O17%Q*(E(_C,MA=M(
P2CEVTF+7FE,OZP0C 57L:T?,<Q?AJPN5W:$3S)QHK'#B ?7ZE 8@E!M.N_!KAR7K
P-GE[M'&/:;Y:%Q)RL8I@$>*6'A7V]!SO04%]<37# X2PMP]05G6)Z+L 5$VKS;IO
P[S:3W ^/#63D\/QF JI20:-AY:?YC5CQF!<*V@U920M?>W3X?(D4[. &'#BI]Y44
P*JA[SN[BDBX?70>F_U#7#L8(?V[K;(M2(*OT? ?ZC2M3^?E@J85*,HFWF*64@"46
P)P<N*"?A/A<6.&QA>T(HW<Z7Q/8.:KCU,K<T8*A_<K]PB'4X>*G5P#,2;S5__1>Z
PVVF*4QX(->'':K$T4:?PL10'GV4<-"7=CW+1P%2RE%+07+JOBP=.B 7L$-0"5N)W
P[0J*;& /OY83[,XN.+^M1G($F5 @_96#=\'9,+F!XPMXT$Q^R'DF C)-8K>-7ET%
PE>2U_HS_0OE%YH=LE^-WT-#0VV=Q_QG7C/1?0"? DA8:_X=+F;BX?2DTTHOCLZAA
P/BW#>KTIB"-4SX"T'YQ&7,.78S*X=]-A)V_@DB8Q4G.Z+OJ5(I)#<O">2QZD43V(
P#>#5XJE/:4LL;"I ?E@_R2-O04V-V4I?8%.^94K:S5'8GGRIT*=_5$J35O7NAI$L
P.LTG+ FKS5$-=R!GZ_BCP"L;H UNE."3C1NI-C,5RD$@N9@,PJS"E[F/;8Q .^Q^
PY5?=>6C2OD;;!""3E^2@APG\V<U-B'U$E'5&)=Y)MJ3OHJ!@G<OT7[KRL&L _2O@
PX_E<C8^=UDQ4^%_"2LCE4,,L95T(YD_/+K0!RF+;I]Q(=\_KF_7"VWMKG@.QXHZ*
P\M8H[M5\^FWMT!LA&N.KB>G@=#[+6C4A=+LBM9<Y<[\M?KV?(0!L.O<:=925K$ *
P"%#%4K&WGS@-V>6.7,'E#?96^. "]RRS<AE :GGR=^;'['?.=I;NW%8@_NN>E<(R
P3\YR4R'B*$803]"DSC/=CQ[% )J-D!%_VE.(A5"G,IZI?E<18'FNOZ:.R\5"AD*1
PE^X!E?K?+8X[0[U4;! R+A^Q%&I6AJGXP$&/%U.%@KU:0NV<3E-5J3/)M64N4KU^
PTH*$1-3?BK4T]%2"%30('1"%2K*HVP ))%1Q':/%J-&#W)%,?H^AH82OB'9PWU70
P[9YIG@X'_>.4S:[%USW5:\@.#%[IF3$<DT<0-D(F)9V+/*W"-/&R(= V-%<6QZ8S
P7;L]ONODPU6U?&H$;<<3;7=H)X?==WAW_4W$[W2JJR%]Y+=)G0;+DBY\!#0J<(V9
PB1F2<4*@VPWI6ZIJ5%P=_"NN-.?-OFET;+@Y;&I:_X)Y?FM'+3*/J=>UY-GS6[4;
PHKE7=L(J3MQY4Q5JX.G),>^0N0ICB*0CM[?1D_U=,ZEO]T*NY/8-X%O *BCQ=-.+
PJ?GLV$L3>=TQS4I:6_!RB/&DL9;8<QQN@LA.V4?BVZI=TD/9%PW.^52""]S^&*G_
P,2I9>>((?#&Y#[PT)J7" (.M>2R5LFH@<"<3R-87A5$,U<[$,IT4;\H-'M+%LM'"
P4 W5OZW2R*'M9.G"#;#"W#.!NC<E-0MF""]A9W+K/' CH5  $#\8[+^N17!920:E
P=F$DVM(-.:3XA%2=1FAZ?:\M3>EQSV'?OPW[F4ZT8B).[HV,!9#][)N/S4[$,>WJ
PVL@<R4# M_3:$ QEM3WZNFNV!:;,_[SB^4E+:J!I9&YAH_S6;C,7 9NNE4]CR&*Z
PB2YN((="VURQ5STKW7V%9XD 1  MC![]I;"GS>=Z$[#'U_K]YJM4,!EWK+'+6&W<
P* 9,LW,B>'5;#4HW/:)F_MKNE'P4DD9M>^#N79+)JD_;ZR>F#LE%?CQ4!$H9$=98
P "Y\8.O=K7*\KF>!P(X=O!1J&W,Z5JV^%J9PKF&.&_-_.&X1"/AC9%> ]MAW"^/C
PZZ ]^U9L(AC&N\*-!>TH&(;Q+V50-:X)U?_K K!>8T,0 R5E*\'CJCC)4QI!4";A
P/!GM;S#S8LRHN\F)NW&K1T=)93N7%W+Q$XZ?-J%"VO3HO<95!@QR>%8FLH9G!$>K
P%89#IKD5\)IR/L"9$.+?<_ 0(K[?%V5^F!>8BI:[<Q)<X7AF=,OUNYDJVT#*CN/;
PXNN**_C9%A<U>2!'&I]9V(MGC?"+B^A:UX(KY-(%TB/,VCD%.PTL_.G%XZ""S[_:
P5/EG8'"-\LK N4CS;+G#RK;+PXR.3_%^@+CQ3+3.%FEIGI]ZGOQV_MWWE9X:]OF$
P<<9 IQ^ L%VC<5(#L:C(2CYCY"@M<7?;@7?"PVZF2,PF.2>SXKO]?9GJEG[\#MI%
PRWQG9,]IQS'7HQ5]00$_U6Q@B:I$H7L*3GK./%+ .[ Z:!@2([.L!_@^2:W9XM5L
P-MI5@ 0#]"?#8'=+G(KR!LEU2)"I0IAM=;G\N(<<7!R0&!A.OJI''FID>0$_F>AN
PNDS3)2/1K=:NR4B]NF<\=*'Q1P :'VAO*HE?>?:I76).\4*?QIWR#7*?FBT\FBC8
P&US3MG3/9JV@<J!B3A'TGVHMO>"X9_R.4G#SG*>G!A[N"PR@B:#^!X'.1W)CO]I)
PX _'>VPP81."ZXE48UIJC@.]']\QX#$_WC0PW[6JC5_4#.T$;UB(YPV+EYH&!-R'
PZN_\ &5##7SW(\XW01WNE4 &T5"<6MMRL7\6_;QW-H)O9UQA&<R=ZT#3:8'XJ6CV
P*2I.9""CTKQCO20QI".\JG&6F"GM?YL@BE*&[M:P]G ;3!6[ O+?K)<G3+X7U:6:
PV>4:W=3:+-$9@372R(YU/FHX;/J&>KVZ<?X)B*]!Q=3QBE12X) 4U6C=U)C./651
PK>.(WO0"FIF!3G9UF+9TQJJ41?,>P-MQTVZ0.CDE*+=-1A3QL8G(W0$D*+;3_KI<
P\P?Y+KEP6C9YO;H0 )B&*#+PZU-2ZH\>F8'X56/]2\BE$V+,Y;?^DI8=CE=%B$24
PAV5$8U-3W5>=5S1<=EQ?7P)N;5[VM\Y(*5G5EEVE@TB$_-P-)8+%@R@$OXND7Y#G
P;ELF_A><C!*T:"[!G.7I:)<&_\X!,YJ@9C&*79 HZ]?-5+K_B1&K59S]UQQ5 2\>
PM7CZA[3,W]AQV8(8W?C?KTF3FLRN7@Z6M(%!E+=J_IE2NDO2XR.M)-55\0U:3?T)
PDMGGH8NO*MK %\L 76"JAY ^+$GFSH-GBNRR!>Q*LU[X6]X43"Y-!.K&IV,97K0E
P/&\K2?ON]>8J1>>WH842R/$LGC=X5'<KY^.H*^;CQ53/:D)PEX2?O3XG/UE9HMYG
P+$7JQZ(V;$K^6_KGU.+*I'VZY/O:X.Z  1WS:8]DI;9JK<&=P?C(04,9MB5#_WE(
PB;Q]&VFE;[HU22X>JFJRM68?;C"Y823,<"\S6.'GK,YD0V&[C^5GVT/*?C&0TWW^
P9W!5?;ND.LN=V<\A8+_[#M'/SU'6P&Y.2.B[>7+RX00>V!A/C\O]Q_[\B9$V7%C4
P9EO@PD-'-08<J4N)MDARA.:9?WL4(/\PT(VU>-9?$L.>4/4X]U[9[!J.73F#2$^P
P[=O-9AUG=:,RU!F#31HH2!:2''^ -!FFB%/_FR:3J_84]^5;*C4XSHRM<:3Z92>=
PK>DM\_6TF"S_L%)!$)47W[W=<1[-BN-A (L]&YKA)+[!RH'L8VW;84^W%,^I YJ[
P>J\02&SH)/86D#\(LVF-:ES-2?D<03W2E9G1N*$[5% &"[P"7,C:T]2I$'JLU8?I
PZ@0$0@%G?2=[*X?Q0<EY_QMI9;XC9SHDKG7XJ9@LR3RUC]="4,\^LZ?40XXIJ='@
P_IZ[&:W9IMYX%E<*J(VA0V(#)6AQJTAB?0#>B0_]V4E[O<7QQ6,S/^OR,BN-T) P
P+YQI+1Q-^24]]69M%5Q'.XR'!+"!&TKF^A93\4\%CI $.WT_V'*?1=35*I+"@:H#
P[?F('0U;;&3!>9P*AB:,"8+#\>&GI[^M.RLQ&NT;39MVB'DEYA#?^(*W3RR0=VV4
P%$,JK"/MKMQK*25#*>\$30.;[YE Q;*%>&V/X-4=(,'[A*1NR6Y!!W;)QQP,PYB^
P$Q@7_MCYC\)+8V\:U54*C;-0L(/U\P5X90 "7',0<-T&717DSXQ5E*,.0B#"RT=F
P1>KE,"@X WX9$W=) PQW; -Y8;4@#KX'N#<=0P <?70KA]5X@K4@;-XP)Z -%06R
PT>Q&!8%WEOT#(^BP\P18!0WU2;A O/H 5],RJF7J5;-2V2V%N\),GR!)IDL6A7P2
P]D^2W$,3KC9\*%BV'MX0V?,JOS#13MO9J5X\X5,:_[?#Y-VPX:%_4Y8;7,O8ETKP
P*AQ&UF9O^7)PQ3.VBS[GY2$;*N^E8,(/0X1?DF=QB3.DIF ,3 BM#UMF"$,^!0<V
PT5"4'(.FZ9(!+YV Q:D)T7VM4D52;3#M&$![;YKS?#W, UAY[A5'BPE<1.I8-%C>
P(:Y-U?=Y&FPA1".6GU>##@,UK!8+EBF^(6IX7BM%7C('D%O]<3HI/F>: I[*[WP!
P?@>($1+H4/TO2JX@O82.Y4 KC K+Z[?^?-F/&*R<8Q]M?]SZ?,8ZA$YOZG85TK:'
P!4R-F5\SP(N*#.\6YT>F1*9&WM>Y1E94Q7I^9Z K.3T<%#NI-62W:]3$]&T8Z)6W
P5%4E[1K,8*16ZZ:+%H%\29"8+$"(FI7+Z](57JUU"CQ"%06]5X-!.'L"?\1VAR;.
PDI(R%J;[/PS'ONP/[<(=8#$#B^-0BU >L+Y?X:CNAD4S!<.,;2S-,7?V6WD_PXH!
P]I5P9S:DT!8/9S8_REWTL+FO($O R..=!2(5.C[?!W[XGE)S_B5N:@O2KSBXVZH#
P'14=.^]ON[,HU: LFA61_*=?VKA1%V9]+JP+YC!\,AT,:.@BM"3!*^2.)S6)*JLX
PK(#![#?TX,9C(/'YV?%W?.2X />EG)H136[0&"..7G-?QTKP+^9'L)&[A!Y5M=*4
PIM?#TY"8W:X<X[?# D</"<4_!U!<*M@GL%%IO ED(>>O:,L.M1>.PC,<C%Z1(T07
PIB#XKRWU]:AW&^#_Y_ZN.0?!7RITT! B\V!KF,F@Y\=N6W7!W#X:_GEZ2K[;389?
P)3Z:U,<LC/)AQ*N^X$$@J$&3OS*UO(_XHK[I&O(<,!S\GP+%#EH%<SP-OG,WU&,7
P%68]KBC=V$D]DVYMX%M6AVS;]GCM/-@4A<P+;+?AK/\?VS>'3ZH^42JA*=(N(SA9
P:->QGY&W)P?U2&8S(++=I8&ZQU\Y4!43:E2]%0WD:_>3.F29_#64]0K]AV!(VY[7
P4GM4:V3/J:R2LQ: /,>6["B[MY^@,[#9XBNTI+7VE*N#=O$4\M4+DPAAIHL\K ZP
PW6X0!TP5[L0?)U6!J:2LD3(K09J<;ZI0/L:M3#I?ML/^^)MC&IR.,N.\ 419" /S
P5D$26O:J 0WGX!8CT52SDH73ZR&QQ<8[A\?1<,S7VF+'1YBH!E13&))O)US5]@/E
P86C5EP Z]"7(P:SH;F%[-TXOK9HZP2LPMU/JGB"X"C$OG;V'Y2[;\0R@5\RI^4"@
PA<(SGAB9SB4?8""LB;WN QPI[G4O>,-6F&U2M0>%'FEER\\;?4,H(S)H3^6U\F@:
PHF&:O!;80XO+O(YZW;VEO',U UDC^:":YP3L)1Q9R:%!4=->!ZI$$;C][@FL2B:H
PGCXB[A#1C; ?0M=G#,;&M/P'9Q5X(,CKP-\70\0C_U,8\B08..KFRGW.TD?K@$HW
P-ZHJ!'=YJ_7%%TY]*:S Y^UN.F]9B+HFI3=AS!TIF6MOX8A94\P3[3,[Z2:G!+=Z
PW<QC@@^WAQ9*D9U PQ AMDL^-3N/0T6 U* [$.1?4W@.R-4_/ =UP-FQ.EO' $7A
P=2QI?$G0#JX'$RBV:/D9UU_E2<?+:@.H8Y84O\E T;Z@0+#]9_GSQS+&8HOS([U0
P6+9WXU<JXBH3"Y+,^$MVZ?)61R-L4\ _#7;[GUB+6S [^.LD 4D-L&@QY1^.YU29
P=[+8PA-"U*F$&-\._!@6=64*4IKF!(@]LZL5O#PS$PKRV2R3P0_Z6'T%)IKQVWX*
PC@/EH1#\CIS-/2@O/)7H>JNW@"4'2,S%%)U>J%.V0&M0Y0L[X_M<AJDOE^9@&#U!
P&7<2BX]"TWEQ V,##4UJHM3T*"*VDSK<Q,HWC(/G=YE4KGZ4/'-H1[*G MU);_ ?
P?O^R-\<1K!>BBD>DF'P^";AAB(3I?.)J6Z4C=GY$; _);B<DXUB4P0?>(>R6?840
P1=#MDG ,<NO='S-UQW8IY^'ZQ$!EG:7+?_PXOP[Q3O4&(=H?YS:Q*C5*^NK@P"9J
P_0:%3Y[><;C]\3RGS!X'EE;<^;/)G<-P^\HBUE?314H&&E0DZBM4LL3 9 D[J4*Z
PQK/XV\2];T[9_#61T'9TZ"SE*ABS.9#.ID1*YG:()?='_ZQR1>FO;^*3HDBGE-4\
PZSN[>&-'D=7.^\Q?S\;RR<_8D!,06CSQUK[_L,K]LV\J6_*HXQB;$S'$!U>J<W"X
P.[V\ET[Z%.G)',!>OAA.!\7B:%LM./;8HXNV 3KKMLH*JABH8 9H88TN"L2<8Q6[
P7G/82PF'.-OTYN2\@7P8[?[(JTCO\U>F8<";6+$62*>N-.*66FR#.W>9T+^:I?UP
PA+_S4H3V5C$\@HSRX.45M*:B^4EEXTYGM%[8]'*EIO><FFKW<CC"+I(!.E/Q]NZM
P)85< MOGM, Y!K]/^D68-6#I8'?7H/<,UD0+WIAZ%*L,B0]PBVE ;V.WMXD.CZCY
P_[1;(]_YQ&>E>#P;/XX2:)0;VXABULOX+)DH!1M2J[<E:IL.EPQ%W6=T<./_F#-0
PSX0M3:(TYNTVKH_86V)P4QAM0O<CUD_E'#$-M09Q11NGE_P_G$\>8U.H+,S@(A;'
P6?VQ-#_GY+WR;*]\6FBWO4]?"5-@ADJGR*E'5Q7SAA4)?7S?GP"UE4,#&N&Y)4Z)
P.<9BR@@I[P 'G,OM1_,E%G=3*.J(:E8="<I&(_=:RJ,2FCY<^G$";D.5_ HEQZ8^
P:WW)^:P)\P0FNEC[0WZ-:*&JS;>XXR]*C!1O3NU?O%F]VN<-A!D20F@:3%%'N%FT
P:@XDIC\QQ^P+KX;>69])^,.6#@+M,/P@\SDTZX+;@D+XQ?"I4HS*\1P_Z65R:$U\
P9]:HF2H]%,V-DW+UY&HDVTU2S/!C\UT(-0=$6/@I,2%KT[C"-OT!]@C60SV.8@C%
PE+A]B_&'26WJ#%Q^2]_"8M/0;F''9>BV_3X"1+!G5@7)ME)#_R/-5\]"@PZ()I(*
P6AH"0-.&>*HKEI:VG@#J)LPU,O=F4V+8R'_:T)9_RNO\4Z&32 SR_N-30^=_N M(
P$L>JW"EF40)47U@ZW7+#@EY_C43+D0L^&=6!HI[<I_G0\*@&9&_G%(.Q>+#9POUH
P?D,OVOBS@G9$.C 0L%!')GA%3NA%1K&V3*N9I+M&LIOJ!P,!\S ]LFBI''\PR-B^
PY:"H&?A!NZV:YI#\CG!<A+;!8:)9SZE=C*O.6A9WXU($D(L0QE?3"?^P T7X;+GR
P.27LZ34C*5:([Q?25'F2W<B^H.KMU*?EY'Q(MVYNJ]<%A.>'0V><_9UD!/)0^'ZS
PQ40X&*B2O@+Y5UT+H:'+9WS["G$\(L!4-G/(EG_VOG\L0?HKFVB[(,LX &JEJ84S
P86L,+G:53&F+0OWI/^C63'+<3]HWT <&@]B,6#E@ C:[B7N4NZ&JAMR&#5E5'4P7
P:K7$)<S*H43SN\LC8:KHC]?)Y%N\@1@("CY=GKCRY_VJ6P^Q +M[9?,*(D-H$9!7
PV]Q2U-AEGQU]#<+?_LA_;0A1[AWE$34=:?Y4+&JYZP@3R;2>].7K0SQV_SW+49S6
P&K:V#(2_-.\"T0+PA8]^"(Q6'\^06M:^\MZR<70*KM6NJHE4Z%"A[WI!D%>K"A\S
PRNL#O<H18LQ_C]3B4:HC24J;Q<4]-66Q?QB=_O;K@=DE%-^>=$9PT]ZZXO_[4(4]
PL.W&>K"N=+F0H^QQ#<GDM7-*MN5H.'H=&63?QPQT5:J3Z4@Z'X_KKCD1)P\KT/OS
P#J?*R#8NP#R"XK3V--VQM/FA](H6*[8I17-T;O$N\(/=,G;K9A]O,$6BZ]I\QD8#
P9FZP,9,AR.>,'+2)NQ\[#NH$>.V9W)1'XU(-2!@Q.+IA2$V0 Q1"^T ZD '  21%
P2#J_J]'Y@FQJ7'F%,<S'F(0L0P560)+N?K<RN-&]YSOP6W?Y-7"L8?@N*$C<,@DH
PXGPU>AS(ED@3_T %1>8B352]ZX.K>0L'3%3;)DZK%.^$)N)R$VB-))^4"=WY7:K@
P$+)I(-.>SBL6.1&3$[B"*GE?T=^=FK@ME6.DEE&L9#AO>U "5*XCTG=/]LF4HV1A
PUZ2I@0\?!S;33&,^CVP$E%\B0*OW1^4:%RWX%$^-T=_?B*U2T?@(L28K,DLW+XIK
PE%Z G2:XL6Z$E$>PQ"3&IC$V&(#YL+JMI2!^]^_>$V53&/?@S2$T^5X%(,ZOZ_^L
PG\8$.RX42XQD[;.4"-"=Z_P79@YFL>[A\W7;_.CU\DOGKX4:?T09R70W0\EDA,)3
PX1=^55[QRGGYG/>'.T7+5-'NL.//-]'50QQR$/5_*ZMO+6G'5W $,W6MQ[*S$':^
P?$S#M($^7(0ITGTEWLN@F4]AR_9M9\HP]5)Z[:A@@I):+WKREU7+.Y^E8XDO+><>
P+W7!V.J<IS8'Z0D5YM-_M*1[\1F@8^V[.BO:GLS.(Y8C-843N\$/YSEL#'F2LWN4
P2<@$4:5P<);R[W3?N'02^5\8!FZ52^@X::*Q[R<T?'MLG=; %\K@Q8L#FL*^,TK;
PZ7!Y'8(8>/:KMMCJ- MS(/N,S#8)EF@9RK7JRVK*\,UN_;KADP4=&X#M'3E&\$C_
PB+#/F1# LIWCDJ?910C=Z86(PC>)^;&+;U@@'$G #X_0%#?0KT%;Y6,1_X!S4.QP
PCZB]HE=QNI95]UXQ&G)!<B]YX4E5AU?_C?^3UAJ5HXX2[+!V K'I@T^3_QEV>S@=
P/099ZZ^' 22 2YRG3D@OECJS:W1<+PE<5LJ <.%5SZ;)8M'X+?2"?AZ;;4+V?8XF
P@0Z;B9RJ*QU<Q=G\55!1K8*7?E'2'6)QH9+EYEJ.I= D[Q3//,SS"UZ<_S@ TP!0
P5<;'2-&S_0=^4$]7A:V=&:\B-DI2/%,]F2K=P#P5DXQ=FUE&#DR3/X8DO]B,X/"@
P@5G9/'S;OOADU;CW\#034TYO1ANJ8:F,D-ER@3PTP;':UU0TAQ3[) 9?NX!Z-W"E
P@%[>)-X,_MAKX?SN?[@%]]VL)G"3>"H\@604U4H7VXQ/S-D8EG^+@8++-[H ^G1Z
P,S\X?8_#:WX& P^?+Z,_/,O,[4Z(#,U\L\!;6C(%I"BF7*D$TO2Z+26K9%"E-S9:
P"-5"SE7TQT7CSO96PM][YMH-V7\4M)#KG;$DQ7W^5G#4##D*5_\66FZ*U]HI'QSF
PW7N@%\99_(7HN(VC,9Y%.$\D$1Z:Z-;A$X\6(R[UT*,1'[H< 6)L\ND /IDV:?>U
PM*PDO+;%HL,L 9U!0=$FFD)MF<,I&4 WW\,8@BW*JU)OYA=$0BAW[OV5J<4!"ON1
P7QNK2*7@LEO(LWYC+AZ011=(R0OI9LL&=6Y?]O=/@=DKK]0]%+]I NT 4#4SS->:
P3?RA!7;8[@0Y*SH=<'(K1CU2I49KQ3 SZ3>)-.'QC@,BL2'=\:5*\HDM-NCA3O<A
P;^08C6OYFM_YG$M*6A]MP@:HC$>X%==;,DQ:'V. D&;HIB_6N)>.MBF19KGH:XEA
P*ARIH71Z+81O-28""ZQ/6TI';:X.UC>MF6!7XY3 '"<5!SVP[)MX8 "S@#0IKT;]
PUM<#%Y%'G[SD@2""&I/05'#?, !97U2A  IU=0=Y04EBH("XJ0>=>4;C;YP3*'S"
P#;)\V/X.-^E"['YIQT/>K(9('[8S^)UB._J@Y?>=,&O<8%#A5]@PJ%1@=GIB)R^%
P(#[1 F^V&O(UF/>2PD (1O=$7+-JHE?CKW;#:&\0";:Y=Z,F*45N%+4&#ZYD)'6R
P+8!9H]$I583JK'4^/]ITQ=$;5>!E-"[$F>765KTC[:<QN3(^CQLL^I;C+^]-!4F"
PM=8=KR(SA^3)97]@'>!-\>F:2#&R![>EC$@!5F'GHL/YS+$DF3"1&5">=.>FV3RZ
PTA<C_,=Q9$1%QZ6G/RH/.P3E%6<P2+D:7GQKWX$3 :V(1@Z5OYTF/@8:<A$SAE!>
P+7H@-NW WKZ)Q@#54;E0V\"*SR9$ZM+;4Y&?&6)%7B'H[&9S]FXOJ5,=K9B*RDW\
P?J) @"SOE$U9Y_[A_)\C&@Y*D5,!ID<V<S'=J/SRZ'KQVY8>X^0)U[6R,L;]PV4C
P)ZD7E-@-IQIVO9A?R[;-92@_XDKR3'IY>=*W\>DWY/&\N.&3@W$H5' %)5NX)S==
PWD!QK+5"D!K*$44C=0_?@$-TM-(.Z;HSI.EW,865C;J("*0*5=RHP]7))S;C*4*=
PC;>\)MEMDL)E(]PB>Y:.,^$H]V]WT0E!DO7GDF6G,?*:QON..,T3"'6Z]%TMBYZ4
PS-ZFP'O?[6Z57*#"3'U];WI+'14]WW2G.Z_[JU:FVW?PGSJB4FM;T4!H.D#D/([<
P$C>;\5=$?1/J>KJ<"7C334A/<;M==U:I6Y)SH\0A04G3J\ZF7(J:'VF0&S(_I)'V
PVF) EYP1)M(C""UU/2Y+,1I0,X0/*XWL%Y4@U83;%5K<,U-8->BM8U3PBLEM"Z;S
P!EZOG^"\,DSYF4]2+^;-U,=T-7<!"U-0EBZ0SU;CG'*M!QKSMP>U0:;!-/X'Q#\,
PXRB)@#V1Q=/%AU0;">#<=#L#54DO/*'8&I:>DM$EO4E8&K<>,$H8:CX9N]7^-.Y)
PW5FC(Z?']$7:J'4<KSU7C.]'0ECF'YFZ#OQSFE[A@QB%[^C#C-G:L_OZ :1L@Z^F
P']@I/[(.H]1;8A&21G6P@?'?*]HDH8@B=:>.8>^]5.:5M_:N21 _O(::\9N8%J-&
P'2YWR@3P[I0-9[>+V7CI!J\C(KXP'Y8 I44L8?_+7SGP]#!/G1,&OCKKM$R._<Y5
P5K)/JB.XZ3B.E#CR'*E8N>+3%4P.UO9Y0A>D]0Y^GHB91O0JK,F\]MENG3F]" 0 
PF'*JYE/L4G K[7\S:+)?7JJF+GJ]"@NG(6W0>48^V_QS60X$SY4-9Q1*E$)YF6_6
P!+>A.E$]I!IG4#[<$-]8[?:&+CM-'4(9?OXO;8@JUL* 9US:.1"NP)@CK&5BDJ%B
P5M+1-4UER_,/5JDDC7(?[WE(!0I4_"R] R<X6#00.I&HLMU:P?-1%00/1(;%NL2!
PT'[@0\I$33^O$A0,4;14/?DL55KW??\S5S(.*E1&@1IRY(C\'/  0TXGV%S?/S$O
P)ZUOYSTZ!E:"?. %38MRRP$[\HJAAF!:?WT5A=X*^"8<HW\+KT7M:2\.0;@8SS#*
P#%<%,>2 G6<\O"4]M'/\$<(2TMJ,/C^O-Z]J0O*$5JI !AF<ZP61GPH,FMT1]P%#
PHG:.@==[C)\3]CCI!]B*1 ].A/\?'B]*+?$"Q/DN6#MLZ="A P)\R7)QNI@=.0W.
PQ;B%O5Q=61K5T*!)F,O=M(@Q.T9O:Y/"C,<'UH0OZ-?\[^3"['WQ\B3 1HC)5W_H
P/+^1_^=BYH;IFPP(8=94$VTJ6^R&'.&48P*UD)*0&!->OGG.7/]QJZ^@*)Z=H!>^
PC@\$@\7K<J1^[56[9OTVX9;'F7?-2P>(ZEX4\:K&KX">+'@.9L/6HJIBL+U+(.=D
P7G$.K2C6"(?7%0FO./Y.= 8S\]!=]A@N]7@4:B@;1YS[UPG!>6R\,O$PZ.>&G@9,
P-]" 7KU_PH2@]78/H)BO7TK@A*U*O55!I/.L95(LL'59#J_4_&;*3'G+)122W"!M
P"CUJCR_2_58C<5S ?1Q'%9'VM9'Y8E9A^U"8JY'@G'<!<$.(-CXD*A>CW%91KZ["
P7*6;%G7..S^C*<6<!)P2I@V$@8.)!2 B7@REYJ0Q2!LXNU=YL#FZ<C'!EB^B&?'=
P%XB:+6<KLE4+[BLNV8*07T"2P=U_BEW]3]"'H\]10FO(=56W[&:HF7!)>6?B_!(E
PE\E7$L(O[-8VQ/ZAK1(PMP1/8P(5SA/-*AKMRJQ%A-BD^,$+OAVCHN-$"])9<$)P
PA>^O1_(:X8!9S8*$&^FAW[M)S4))-^\O%QP5)"/>J!^%C:!W9IYDVON$>)(P!Q8@
P_HJMO$.J?NY,/Y7>.MO&,_1&F!$F1E02)][67#,DH8AITZQJN19.Q(O %E1?JF@>
P8A;_%H;CO+8O5BA07L[LZ[C<#UB@MOHJ]UI,FZM]:2B!QSUJAVI[5:91,Z3#)XA.
PS_NK?(MZ/.%6=Q./GB5%M%F!D)*5,"5+(^8YF=2LO+?1' 0;>51URR'+)RF@*C6Z
P7VU9!5K8L%>RH7+6W,5F+561*7J^-56G?Q$8 &,JM8>:CWIE_U3(/D*]R$]R1'LG
PR&WE=7/$2S3X^<M%!8YI"*R_<#T,%O5UV1^_>74VZH<)7]-J]KNQ[9A^V(;MY^N&
P5+BJ1A3#.A*S4-N+33W(,TLZ\[&)JJ]F)PPQ>KALA)Y#*S#F+TQ0;7=T.G:1HRI4
P) Z(N?ED  I2BVPE,WQAJ4$ZH=9,H>6_6+S/7^M/7,PO7Q^DK=C[T;<MI,'0;L[N
P=97W350O$'!N!@?!8.ML 8*03VT/\=MZ<F >O@12S_TN%%J9 ZOR-VCU],-'.Q[>
P[C_X$ 5@EJOG;9RVBZ=!O9)2\?^#)GJ8,V40*"X>PRLSR:4N)_F%[%;!*H>85-XN
P&':MATBS16]J0LP?\-V8=-^=3+Y3#28A*O&PPJ.W;M"/M-;!A:ZB3O/?VH%21OA\
PLUF^6KW!]E;@S@IHREHO8F<#S=:@6>1@ SAI\ML, I_2?)DIWD?DE*]'*XV%[$Z1
P-V'V;)A.A=D<=!-:4>ID;YHP++ZB?-Z@>A9DU@SE\[>L('_C91BI8$Q/]\6&'6PP
P+83D(1-YA<E?#!Y!;</DCV]>\LLC7BLA0X.HX#U5^^DD,1-Z9:D.7V[:.E;;X\[;
PEC2HOJL>N(>;W $5UHQONY.ZUY[0^G ?V)2WY,U7Y#S12L=&D _(\_E=9?*@9TV^
P/DBRM"'&$\YKZG^24:Q$X>)?0S,K(^O[GQ^>4BI[8KM<+B1J]9;2"OGKLWEI"B!#
P=0IU#D!VIY6HR6O]B52ADNYJ\,W05+>\Z-],GP#3BI1FW.?D(*)]-ZT2B4Q66Y4%
P'Q8*"OYUX0%<T^^&F(AO75>B^<G>D@.) &L/4P)T0GZG_;62)TS-,/Y#>OAYM65(
PG'LG ]^EC6Y%\'FU5+MR9!)$IG9R4(;4Q\(^MT J;8L<:=J$6>GN(C"KL^KV]M3^
PO,7IFK3L^'LRWT4*MVJYR:ZPN\[\;]E4.WY.9ZX"0_B<Y#<KI%?C28!PC4C<3Z$2
P93,2!Q>!(XWIQ4A8?[*>>:S?<1[L"-LOE;JKE;*N++6AS$4VT7A [*=XV[2:K+VY
P&@H-2QPO"4*V2ET0\_E/4VT*ZJ_98HW%IV"P!T(@.[H>203:M>$DC0<[ 72']%+X
P10X#6A3HV?OU82KG\9R @:K(+\VE6M+VA>4@" E>_0=,\L:JV@X\6O"P*X098]6M
PJ*% 8EI2$<]ZR"2S19WGHOCLO:*/8U:'Z,UK_4(O;;K2'J6+.!%]'0_VY\!?B@\!
PH/_54W$L2AIO3.D!( _VCUWZE[%\G"ZZ Y3/\"0P=V)Z=+/9.B":D.XV$"<E.G5!
PE &Z "560922]])2+ B-R_#"S%.IT!+IM/"4M./]VZ1H80PYXBT'KF9#'BG+T%2P
PV\,*VJJ9/5B4CPH\J0*]JL$4EHR3#&A\ VCZ$T]T@XEPF(+Y(VY;!/XJRM-.=G/9
PGI-J?9W8R0#*I8CM/%34-?))Y%C?!YWEQ0O6*^E5I>(4V5CQL71III_L9+=/J^GF
P;V/G2NF?S:&IO$1@!&IM6_S%H^736G$>0&*%1IB?5R]BK8 "8/@M?$7DL\HY2#4*
PDIU-2>V!B06:/3T<N^9,N!R!<-XCH<1C&$^7%5(*VHG_.)7QDH2<D=8,A7;*=1'=
PJT]?XZ1RQ_=4/?=@A"Z&T6$\!.XHFVUNL3:R5GZ=%J I;?:E\@17UZD<(&<*%@S1
PO925S&AL7*%8R@A;0(JC1#186>\*&C$@-[P$*)=((F0BG<==6*!T 7OG?(FHF1MN
P$#-X 5@GJ/+9GP^ZI:[%Y&S9L2&XPV)7-FF)0MYOF>-SKF!.P446%0IW83'*FO\K
PO%A!()Q!JI]5])F X6.Y/>^/^Z+^S+X>-"C.#Y[9:P61KSK\\X&=Z'*U?AA =>G^
P_7\+R@#^_9EDK(:RK?!.$OB5-,>.T]ANZG[^W*E2NSWTGFGU1WEN&G(7>HTQ 7++
PB^!@(/[9Y28F\M>DTH*T[H^06H*$!^T)9E4AS!&5'\C>DQ9J;)$D+Q<3OLKFW3E7
PD"X"]=;#^%Y>C8IZB':'?.;][3CJFR_7&2Q4JXHQ\T["F07#K,]?78!8Z?OBOI'@
PXW(=0_E;67%.M#T:XG"5_2!R7S>"D"E/Z%UD8/FJD**SH:8N7O[2WX &#E#MC@[$
P><1@UFU$"%L+ ,+\6?T:VC(>.2O_1XF!W-&;9B4</B]N0_H^5EGO86$Z6\F$&IR$
P1%V@%TES$FQP#EGWM8O%+=9N#\*Y=E1@8Q?HK\I!6OGY1;,OENBJ+]IW2O8\-TG*
P_K<V:[N(#7S$AJV_]Z3(8Z E,7+'Q,<L2K3H'\KXWW^\B3!HT^9.*1PP*!\E2=H,
P<[,PS4ZJD"=17O]XGRA"A2L>=]=Z#^+AQ_<TQ_'G"P_-A[J_]P)S3'-U/S)/G,<F
P2VA<7KB8MC!/_]!Z@ ,&IA=K5V;2VQ\MKV4C(255R&2YL;^E,!^QXMJDH].6&<?7
P.YGO =]9Q_$<VGB22W+PVG+=#<8^3ETG-GZHD*EN(P#>ZG2"!>XG0QCZD%7GM(+.
P8[TC'5!)C_K6N\FOC2\4*#03750U7#-P#7XO;(/$8=9N1&W.+T$X.8Z/+9QZ1>"N
P7M0&GL*>D1Z8(%3OK228#6W<\UXDJ1Q$48T>1%2VJ_ =*'7UC0MW .AR/\)!I&;L
P,QB.O2!3.2#M!XZT"!3+E(#.UTY%C+89K#[4JQP/ 8 3US,?/N!B+)BY!H@A/78H
PZK;DY/A7^#)E\9[)@A?E_K EH1#5WZ$XKEW1!D>4\ECY2<Q"0W#_H%KB >3'+-TI
P JA.KIU^%%\Q72W"_?D(B=K.=<1B<A.ZY'UWG(3G$^R[^./Y[)@TBP+W6MLXAR7.
PH@)56,]IN@!.&&6)CJ "A>+V#UDP:3"M^SC3\:)4,&."'OL)(*:T1)!91']%<@:%
PE6< D"WVS>-P_NH]9FWFMYBJA$T',7%CC)J)( ?G:L5S8QB&B&,<T.>$LE]_)LAO
P1"?E2]RZSP(?W>(_%6L#JRS\KYABMO.>\NV_0:N:;OBG63 MZ2VK&G2Q\+K<U7/H
PS%%>ZPT4+QGLAX M6. O&\BJA!2<NJ4?T).-=L#FO!>3F 2BX=1/=JMHUQ8T5C&)
P)Q&J$B,(VCW[I.Q28R2P64/\O+G*+0L4V)8O]1S[>F,G=0\P3TS0:.<%1:Y]DN-*
P4939N.5+?/*$YXK0"@P#1,8,O"^JA,B,YZ]40;QOWK316Y4QYT,E@V;XS-S\Z0*S
P4<AT@<N"I+L"D% (9_/!I2&E FZ+7@JO0+&\;NN;8D66$H$ZTCO= HQ92%ME )<6
P^-C(Y6C/+G'CF!_=$*L0\]CF@&791#*QJ4S(P>DZZ]^CVIGY<$6:8W4F-H)%KY93
PRC70#ZWNC.U)Q:XOKH;\W#Q4>;:BD'5UQ[!X]''&$WF.![AM.V>BJ.!4)'=)^=C?
P4M2:AA6:'Z"DIPME$<D9+A:B@S\[5(*4"8[RDH&1Q_F4%WULN&'7B4+TUK'L1#-Z
P3*2(H.L40(8.QYG"JV+CP.N5594G?1:^::ZP&*RQX)P<?9IEA5N*4&'S?,RVRU,;
P6[SNZ>Q)0@=UY0 #6P-[0"2_'*=HA%D:"PIWI?=,N3LM8-\8(5V9L$71?Z3^G4C,
PM71@K&HOY[<AJXU;[T+H7:%A>(G"CA<'Q L_+7=@4'BCOL4N46BO B)96BIU/^)9
P03'2)"GHC3Q$MQH6H5/$5][FY.,=<TRD="&@IXO>:BB4[52\GZ;'.GJ'%K(]4^"Q
PF+4%'K]9-GBR0Y!VPIW)=8.FB%XLH9+HK<Q +J<'XW!Y?;W,3)>%O].>+H/_CDA,
PEF?@!#HZ5GX3'#Y(?)I3:VA61*2>;X. 5]4-9BKXIP,(Q@UA"[J3*'L:' BQ((PF
P];#?JC)N*4D/WPVV+NFDC&U8G.? JQN6+EUU" GC?KD$HAGP;%T1\'$3Y"0)7NE,
P@"@=3S^WGZ6PDS9%:Z\0G#H<OS1E];D'L%%$B8YP;:YN))2\?PQYMK('-(6 BY<%
P>GZM,$)-XZM<#:WT \'H(P70MC\NEY.^-2['/COHWH89A?X!6[E2S,QI*F:';W#9
PAK HIY(W\/-+6-,*8059Y#WAYO0=5M8HZ\L1"+YX,?QHN\>5"&%<9K4)%G$_?$T@
P^FNZW04U.>K(:>P+J[9?H=&IJV"S&,?=IFK="?0&\OKZ8501C T\6<B\QIBMER&0
PWR&=)ZH;\: A@C):>&9@[]9%V8-M?>1]FA;@_V[EBF,$8Z-,NHT7/=M:([8X<W&)
P!V"@J7R%D[7))D?JTHWLW]X9YW!5:;Q\F<F[&&A,]$AT5>2\8*V)@^EES%63I6U9
P$B"?.:I*7L%[:EY;FMQJ9M.KE\&# 9"@3>%'%%5W/V@RHJ1L3-2L-?/<OI&*LG49
P@4[CAM-F4!KCQJ'MG524:!O8:*2+7TG6MR@0,: 1B! ?>+*\<L\ I(/54@U==\CO
P'X\B=3Y5;"6/TUOR)HKPN>7E'!JCO@/E^W0.9D[[/Z]ND5JVS-%=927X\.;C3!;!
PM\GP0[=X,0<^W9E,#)UGN8>7MK9CM3<N]A"=I)'<:H'7\V?2AZR.KQ,W:BA[3+:.
P3(M.(PXS!,B9E]H80^W?!7VZ0;6):O/A/1=,G9.:ES>*Q#[]4C6/[W *$J5I/7]0
P V5Y^A4"BCU3<)%J_KX\,=H[D)R HML7_KFYNM[D=E6:H#&INI/M^]CJP?ODE.X9
PQC[H7WWZ8&=V&Q)-XRP*_#RDK#CGW/R*.K2 *Z2TCW3V792, QSC3QD]GDT5&UD3
PO-U.?;U^Q<*<)RE/R\JBOAH*Z6"H2BF_<9MI M=MNY-9FOC:0N :-/85>Z"KMJ*Q
P;!*"\AS9!%F]QV!]":24MGYM;QO3+J-JCV4W^((,2KFN*3S$4!RFK0")S_/=+A#K
P 99J3,)+9NFJ'G'DJ+RYY^FN>, Q;)_]^BZ60)(K(,]EA#X=)NF6"+@M< H=699%
P((PQB$$(;X>MM;.\23B@7N96-P&K2>MB[V\Z\WKTGKL(]"GE?3KKNBN<?>QJ\J-J
P@TM2.,P#3]J7 ENE,_FJ& -LWHR]0+*LQT)23 I/J+78 *)97^;*O9ZS6V$!^<D?
P 5CW3RB6L$33-73=FU[;NCU9I'[*3"Q$7Z-'DGH["#]O]J%; QM#.7]T3'8W(AI,
P%=$^?)/_L[[)$KF:QX5$!"1$;%$754^W# \KE-8)Z&F"@J#2.KT>ZBI%?(N;MFM$
P"D\M_\A;GX:</G33Q]'/[/+^[-3!I,(8ZX>H8 Q0Y[K;WLI12;KBR"*E?%()V$;G
P&W(*/X,SL_C4)2I-EOHUO/I.M%BZ0W73P-J4MSY%D"RS;IT$NB>VD[\TQ'0+WTVZ
P& SB3WI#.**@'ZTU'K(;2K&VF^&J(H^U3&K3F2]UX!UUNE@_D!-"VX;P ^3TTRA!
P%/(3_,.B0T%22%\CHEBV1Y0*_[]]7:;%A\@W:PC6*#'M-=6/9@8.2;M3S&PMPHQ\
PT9O1AIG<5E"?_D#T,.F"A"8,/*,^+2]%!>74+3-6(NC_\UKLQLJ\@4,!B::M,!@D
PBF_88Q# 68B2V?<\QHC\:(L>(FC+IHPUJ(G;V11I"N2 KX^:N+5[;VK3$RT/3EMT
PJUI3Y/NT"4<JI]S>;^#;WE:@J;>()D/P94 E?'7&]S!>U-#']F/92\ZG!4&&A'SR
PH,I2:2D)W.0;$Y&2/@,[/XDHV0OKN!*[HRK5DM#:B9V7SC"*G+L+QZ'W)J2RDP[N
P[R5TB4M]>4*WVCA^]="@EF&;Q*%Y^Q/^5H050UV/"=M;J&161@-2R<(DUX:J,2]'
P,4WEO=_@\"]4%&N?>XE!7;KVX0: O%OIZ=AB$K$*+WM8[2#H!=SC1135T[1=)(6L
P4T7\R*L;+E,BHDN 4[7.B.K<>QNEM-KDB4U!"+G^);B&RN#9WXC$131E[9TN(SZ>
P!E>=#?4=I?+HZ&-.ITQV]ADGKS!@QYQ'AQ8\,:ET0N,L8O(-57PV^ SVK\.G.?CY
P-7IPU%^V&;5>1R9_Y=(+HH,0_]6&@V=4*X05A;"+:)44JY'Y(T$&&"Y[BT(U;T>T
PQ:S@PZQQ_1Q8G>BJL66Z/X05^DPM/$,'/0 59<H!+YH+)8SS6RPFZH9_-Y/MSN9!
PW'\C4D6U8OS60:!IN;T2(8<[X][;6+ _3!MWL)^WU237'I/YJ)B.<CE;4!?_N?I3
P[6 $6J[.C^+G!;>?>[, [4!+?J(87N?>"O4J"L)BQ]2$#H<XBD<5*Q*Z/*-!%K9/
PX(A<!1;CPU3!.*4 B(0\E&HJCKM@*SJP&%RH2)1J24H@]A&5G\J::J_ET:HF[92W
P\X4WBWF@%#Z B!+$.OOY)2<N96GNB%(7Y2;2L8=30L@)(AZYJ0-(<W]K=ZK.>-@7
PHCZJOUMHI<[?"KA2::R2LR!EQ9Y2QZJLIA1:QLZ'D+ &M3<T7_=KP18:P2:]#C"1
P]:M>>L8E/W4!Y-@BS*RYRGQ!NAF(40'@-?I34$$M"NIB]2A:/#0/JXC^.,7NP[OA
PV[T7QN(X2]EP7&SNA151EE+_PRP626A^.L98E+(%)V8R/2+R\M[ ,BU$CF9@U8%N
PP]MF<;%$L:=OUY'1%4D& Q BW]>'X$#R/Q2&/?IVKVNF>L2?'68[ %7?8BIM'(*>
PDY_&?T$_K*KOWZ91SQTV*M1895K'I?Y3/%$\+0C(6 KC A"7YZ'+ACRGQ5?#DS#0
P:,$=?&1S%&Z;2.ANYL$\UOAN"NXU_Z/I(%B,8_XR18JZ1[,5$%5 HUKA);4P1[4D
P>=.?<UD9>W(D5MNT'\)SU2TL6FT]09 2P^7^=ZXA35*J'_3_F;C$PNPD\CL%.0N@
P\R"[2H>EI'QZNLJ^\WRDN9FCNQ-W<.H$MYQ*Z+E?-2S[($+%WJ5!.8PY_6T2636M
P;!HMC9^:[S%1@E%_9 0X;<\IQS9(Z6/Y7Y)$+[5#2<%VU$0R"ELUGSQK%[7QMBK2
P/C.J %H5K(N2^IPP#I0JF]8<4T*KY>XG]L<_1BT0_><XSKW2G_9 H-W]4_B:%/N&
PPSL@O0A4^4MCG'BTC#B>%9F!Y'U?]L>"4GI-J\SY\B\#Y6QHWE&<7V(*;TC7^99F
P9F^H&Q[C1ZP?GY\LE+^"&(\OPPBD+,#$.XKP:F'/XJ8#</$P'%<6XI>@.41/63M.
P;4S*]R>Z>YRL\/[AM2U1_@^-%3(RX\7MSO/;"F-+99XVU/#%V#-YZ-H;394@\P3]
P>N!&?>;R"?OKP)82M,5\.[M*^;(.YD9X.=<Y)6  JK9FMQM[4+(2#;/>4HV0BP9A
PEE10VAJ+@$LIE"S4J7)>C<"Z:MG=DL'ITCW6L*,!Q8S8= 0^RJK1\8H!B(X0#1U-
PT8>\YUAQB!%F1)\[7!M..F6CX/K1<;;-.PK1 JR\)!JI XI'4TJK%&)'8T=N[VF,
PJE69*(#>WI4.I/WWN^%89-U.8;Y9+U 7L&5--9#]I@.;2%.$L [&;6FAK_9272*H
PKX&WL-B8EMJ^ ]C&CW?W=1-(67S\"5KKI4;>&301%L'7O<ZO\2*OF5UZ27XBJ(%B
P!T%+:TEO\0SKZHNWB4RD(B5!0X3<3;ARU$6S^6<B^!N?[%V8(9ZCE"G47$J"."I&
P6(5=?B9FN,81@2DWU&X-+H/T0#3/4,HP_$2311UJ&?HQ>95\$QC;@8)M*T:/$=MS
PQ$>UV ?-)SS-L]+NESH5A>)P;V/G  /"BFZ<K].A>R5:G\VI7RGMH/T; ]6Z#&#M
P#0S"SLV&5@0=&%43P>VL$9T=-B#WS"<GO"%/X'>\<^VJ(_;79Y :5_/&L)HC*CHC
PP,$Q$*XZ_9&I,75M /&F%++CWXFLF^E:A<Z+)@%3<!'$\_BCNYJY/*E;2^;6#%"$
PO.<'R+@X4/ZQNY_UIAJUZZPX?@7%E(-8UI58IS][XP@+\:]EERY'?#"$6$J/YH$4
P%C)QEQ_("#J[>9VMHYN".J$7>YVJHB<D3B\SZ6WPSN/\_A[<\ .2'J?D2W;'O@,Z
P$(1E59'WZ;(Q.#+^Q-G%XT\FXP(%2AE[I9:RM_GQB"W"/N&D!K=7HW@W+G;(F)97
PD!3I$ '/<-]K/XAVJ'#^XDQFG3E03YTATHME8FF#1FL<\9Y712O>R%T&7C9M(0.+
P^>/,1*X,-@!]LE<<U?I6X@H8)E&VD(N+3"3XY@)S-TO17X0QXSVY$#;3<JC:W[2&
P\>YG;W8+^J7# Y7ZXU HP%@%-3P@H<[R_YS":OZA;*)=MQ5I$0&TR/-HU:L4?:U2
PP(M<,H0CS81@1!IEESYX]5F!J&TC6"G-9% &V:R215)1IW.>:4PA6R+'8WNCZD (
PJ=0(BO/DOD<.2!6,;/YFX'H^KF /K2Y09GTO)22 35HRIT3K._##>*C)XYXPJO/!
P?F 6:FA#-ZZTY0(I[J17&T9-S,B(,==Q=T%HHG4%WG0T+PQ_<YHVP9(GEN_@0:BV
P&HQ?'*I&J6^?.;VT2P86*!VW;B&7+'&CJW3]+YA'6YH[!3<RY)TG/FV15Q9@/GN]
P0&>EV>3N6! 3SLRMLF\D"!Z,#T'.ZO8DXFF"IK-T)AF?[XON>/54+[!!I66K)C*?
P^=)C^Y]WQ%=D.]NQ_9D5!B3$E9'';>Q/Y0Z5TV>8UGM;%%^^W=5XH@Y;4%_437=-
PTS38W-.;A@M#KM@JXE;M?QVO[DX97-G+YX^W9LXM]#:44NZ$T<S21?FL+ K7N*($
P8=[#3.[>)>63SAQV^FX\]=+CBGL2C^?LO<T18FT<U6'_Q^PZ+'12I@0Q.PK4@TXM
PJ:9JV;H'H7+)/Q/T,[CB @YJ4(X4 <]'N'SM5O;2<0313T3R?[E'&)/@C7MAE])3
PD D1]719J1AD;2"[>G1!1S*9E;^6/T2().-J!/!;5[IC@T4MHC6I]@1ELVP,(&A$
PX5[G^)7E8<?E3[IJY_7#6)TOFTGSN[OK1$!7-/H/@26VJ=4!^E? B SMWR<!IT1W
PZ;L30.#;MS<V&[UE2PRVGE<\M%4W*O=NXZ\XVAWF3M@'2D26)^Q3JTAE<W[QT<C(
P%ZT7&$) +:UIQNI@ LB>]E2S^<V)H]2HM^D#:N:*71+0%_<LCS9GA[$$\2RHH"R;
P)R@J!\=[TTFKD0U?E7Q:- J5[]]+4&:I'/X_-UD26,P68F_,AYI0E$V(M&8+3'=.
PJ"&(";-F-:2MR#;=YSI*D5LTDP5W%1^SH@(;I=/X[,&;5IU-T@L*56R> T*(;-X0
P]W\\XJPZPAO4.>KFDL+ATW:9!U;Y_V"I2)WWA@0 ]U(] ]4(>^=KXDC -/TD2?L:
P[A75=6&7M5Y!:?D:ZDDZ (23?'Y(G?%#:%EK+-RDQ,X<TGUBG<#W2?TL^,S,,V?O
P )G #M56*[2YR][@[<FR72!W);C[<"LR?/YUD^;#+( 4.=MB6.@*K;7]NC[<*S^S
PLB!KT<25-BGO#2+7@B7;+NN!3R&D8RAZ#[6FM&.)R TW%ZF.)=6)+TW8IN33:5\M
PSY_K;[:#II^2"O\QQR$QFMM599L\):;"JKA><+O7+!=TII)A\:@<-GR=Y6.NKNTB
P."4^7]*GLEAF!/#(#)"*Z/S@;Q'&1+U@=YW[_@2]1UQ4I,!0!\/8W'>2.5$D^X2O
P+)1Q-#P>#?T)P-D^!P6^OB%EQ=7/2UE?,UTSCXMD#=;TA.]AWU>7CA4+9:TYV._*
P[J"DL]-,X.V=Q+O[TV8)U(H)C[E>P5]P%*V/7YJ]1S5O"]NN"E>SWL$"P *P'W!-
PQ:#,I0_Z!DR1G(%;"P;TQ7U*^'$\>K URYNP>Y*LF(%,_ M[B'UV<MH"ZV%%!8G%
P?Y[Z?*T]:J4XO,1I0HWBW#( A0Y7=*W[5(ZR>(=F5Q+;5QSI60HU5!WE>ML F?E2
P:G;>?#*GD)+T5CB9&L7&&_8.+.3U-WKBTR8K_?V0Z##0TFQL]%T>7&/T[7>.#6OI
PIC-S&39"/,5:IY /'?*Y[B9<;?]H@03-&7Y0WH]9?1)$N,@YF8;9*ZTG:,4L@<L>
P"=XG8V$ 5IKU;ZD(XXN[ .7&[MCKYQS_1'Y<5?&V!0%4A])TD%.X.JI.?.R-.$V%
P =Y9.FW8S[D<T4BAA)_J1US.LH.-((4\'+TUKD$9,!GK>.XS=1U,^3^:%ZC7E\1X
P[\+HV1Z+M3IKL V$S0/\4,RZ"(32*21HB4[SGY-K0S*V5ZIS?XLHA#*-_WP_0;"+
P2(33GXCV[#1J'1*NC^<'&.( 1"0/3,R\@]=6O/I0%DQ@B*%N8UG'O%,'R4%3,H01
P,P2 CF>(78L$)$=_#S&]+98 4&]54XTL;2_>&^+PG]0<M>#7GB(_#"]B:U]N3 _<
PNB9: X$&',\1BL8X&;.NWNK"L'Z6Q, >"DC,'+P-;:2;F-R[YC:7'2SW?Y3M%<K]
P-#RSX.4_[4D;K3\PC<BAVN1"8';,Z#<0 1!6=TECXM4RO(KA.FV9F)L8?:ABV].Z
P+2AJCZL.0KB^4<%Z%344[+MKRT.\N/88ZWF@Q-L!MS@*2-W:;YR^^(.UZ#5;ID>\
PTDC3+<>.G_B)8_.9-N4TQO/(DLO<"5#CT$JB-34J:DY( *!UM5BWHSVFEA4Z?78X
P>_]K294W1\]U&G-#@P+A[G+)$O'\^G1?2\*ITBJ]"F-Y#[J>9O-!>7CX %3-J8J>
P^SSAJ2=,$VIW6P_P?#Z_058'I/D#W-M@-#=<1(!B8HZ$WX]1A0$$]:CKIBLT5>6P
P_,:/SYZ/KW6!SS)7"127#A27.Z&M,]XJEFW]DQI^YW5+L$I2+L2=V6 N;3#?S0*D
PW%_2WN*7ZHARM.>V%.J2GM2LD5!1<TX8@]9V)5[8)2B;@NL]!S(2=(<SGI;4XEJE
P=DK#.[*K;8B8%3;C^.!3XC1^RQ'Q'A)C5O'\"JWQ=)P^5)>VZ&:_"<KMYU_\J%>"
P9->C<.4%J'<PIZ*!;5\YM'ELIQF/_\U^Z2@6Y3F&C8X:"SX%ZK^8)O[6,A?N_SPC
P15"G )]NRJ9%U,.O1)X:MPE;=<<2U2]H6[WZ^<F.%M+]J3RQH+F*MMPIRTC#E,EV
PED)1_*G@P18]=\73EZNV5TJ[T$ V9LLAIDTE0%S7D@2LY95/PJJWVX.I8BDXBMS^
PT^#35T/\M4,EFR7*;Y+GNO<JUI8)H$6GO$K1;3,P6-J4.:FX:R 4;/>PE>AI@0VJ
P7)2[Q-VF7:^NW4/L8L:XG,YG68CN@;2,@*Y&0 XTW=I)[UP85_.+1 PC/G>/RT9P
P>4,'I.HD<J$(L\M$6>_J4C"YOBE4G-=5D$9AA_\?<]M:?TS1-2OS< 1 ;>%^SN3/
P!Q8X(@3)[0%N-40;XB1@3P"T0#$6&[/?92K!>3;&$F/JOG8H:!:??.-PQ@LN(IP&
P4\=1&;-=@QCI:#W6SC5B*!I>[7(]CQ'-EQMT,^%!(!;MO67;&BD*1.OV/%;7Q[IM
PZO.AMUYDC0@3FT^KE']%?4J4;%UUEN)_K)=*I+N3JKS];'CC/L]0BX4PTC\5,<HY
P8)3#]?O(X\I2V2<]\>QOFQ]M!BB74LU%$TLIW?P4IU;3W(!N)3*;$>.-?7//:LXN
P\O[ PI+UQF7$)R,WQI_82Z@@\TTJW#7OHG3V4 JF]JH-=]HW61=F?OJ2YW_O/.B+
P_3G!;[R[^Q%-RP3U#^5E+LS9>,#!B>:1F@'7^_%3[RLW .XG;FLW#DC4%%#<JYR@
P3Y?3>^C8PB&ZV>YX+Q0QFJ6U]6Y/)KA$"';41DT$9@>D)6<(NZ@'7#W(;%GAJE?*
PB< !=#?MSH@W[5MA"F.3$:JT5X2OPK:7NHB>%GNM209<"$C$E;RE2/K!*O[9T%YP
P)'-<*VQ,SLG=O%J<$JF_.^4=-&<B/E4P&\S,*TM+ ]!D(!2]>NO;L>0Z4KG>)94G
PPK.]ES<UB8._T>"*C7A#0,0_V$_IZK]"0, *#ZI!I8E\EO1P'MCCS$?6 F$&F@O,
PG GPCM<&R,=9>SJ@[T*)D0>#U(05AV>EV)\ A !X2.\Z-Q,Q7KR3%:.'&]@(I<I*
PF-1*.1WJIAB%R:%;,J,41%-)L"'?J739,:DEJZ>=AFEAS5SOO+ $(^88?.@:#%],
PJAS"@;(B%GQ6_1/YVL,?I=WZ=$:Q:Q==,:%M58-.:]OB1J9]Y>HB5\;!?<KLGTI[
P*1KGZO1NONL9"'&[;B9<XVDFC\7[.><R/7^Q>;JV3LW010H(@MK6HZB7$B5L%E+T
P:\RI7?@628U9Z;>[!PJOI3HV<4-#/6$27#4KM9MNM;77O7;W*5>@$7<O.[/: [C'
PC]:P=,7 5NY^GG/$:VP$'.S$;*[U,67+9\>\NP6<<Z/1!#/ Y\#F<B6! <7)BSL!
P$9@R)D8SY"T;((8',BP^"><Y7E[O+UI<CA0QM"K5<1$Q2.OWSJ9["77W6+;7BOC@
P ,5Y@S6F7ZG=^E!LB2&A%YZ%8WC4(CZ..B?ME=NJA[T(_N^<]J07JD4Z'7-@M6TM
PN!*^1"RS?3'' 5"\N,4%.HHM6BK*J&'6Y#V)U#K^$3](4/N#[,,=%E9*6V!XD1_[
PNSD3 ;'@+LF/B#/'HG8KD2G.*>[#/OOPMNX2A$\"%-WI;/7W*@[@,VQVO4B%CPE=
P9>"Z.U<0K7!_0?MWO>B>6$OB*XO*Q<VAMD\B!? &2/HC6H6PH+L6]4&\<75K1VW6
P:WV I3-#*4=8,7',]G<NRNAQ+#*&LZNLOF6H2N$*^+E6L=X'^0BP U]Z"F=/@#N:
P*)D2S."X@!=E #HO)VSJIFT_+4G*S?(U[DKJ= U831&CL@C:X#8S"N4^]:^2<*1I
PY-/=<$9EXXQ6>++<,@_B$N["("AT:A+_R9ZI>6%Q^*&O?9K$N*I*21%AZ(R.A4SF
P)-EME(U);!.+X]H;/'PEB=9D 59OW[=[7=6,CL 5AQ'-.O"72_DDE6:OP5 N85LB
P!N!]DJ"WH:X!984=!#C@BCDB9Z:J1/^281=A*_)^88@:JHW3-5?RG7N;491%\I["
PJ"!TCLQ2!B+2>E '.LH5RK,$NOHC%++[2T-7KQ.W%@2],6+3103X-<W.,0<?@C)[
P[_\ZOKN$VABY7ZSGT9-\@,1W^A]FZ0,YQ.F8F"T6EOR-E,S0.A>M=B1FKOJU+D\^
PWCX[6S3HNSHV4*W$1\9VI6.&$ZB%2'L 42(SV8<T#"<O[1"!.(PW=HC_PQ:&=DD8
PZV CE+J^E)V?+J/4V1&F=9FW$FUOZLYTVY6YX/KV.PZ! H'\ZZV)>0S3^@78=@D7
PZDX !.3LHTAQ,LB0=:10])C#_?P9/T14V6@R#HL$V0^ $OFL3* *YH<K_.RM<3A8
PM12I_00DH^Y?"NO+9?L9KGM\)0^^WR,5_-0/<">&ZBJ$.3?60H^44S>%2@)RN*E^
P_9=658]>-AHG$:YRUZY48+Y4<D:J16C%C?L1L]42?C= _WBPRJ/L"1%.^AC*,!-X
P]'GII2LPU'PY%X?*5+XOC7B?)^;O,T (;*"<VFW,VOW- FH/#V0L2;1\\W6X_H,!
P["%8Z@Z?%^7L(9]ZY1MADGOHO%:YHL"RVFEQ<Y&\3<2EX%75/<DWO9+%/V*2L)QR
PI0D>3?1,:J<AUG/KFYO<R-U-K!'#XA2"@[CDOMNYG+HQ%=;:CN.F $,HU'N* 5[<
PYYR%#;'S?X8Q"#\VC__B1#0;'VZ?U-34EX&?"/B4W7"G*V/?[ND,R%:4NW$DOP]P
P>Q!E(+:\!#.SV;AT'<Y51$.JLAY$U@03)W*84'V=?:"(V\WKV)_$RW>D(Y<T/::?
PI.< /FFI9JJ_DF-=E<]*E9]F64Y-/L\<%PVSML(:= %OP>W!*@5?^HUS.>U-*.FY
P),@G_>=A2Z;9!\1+;N,$6JIU_W;,GPY(_V:*N/$N2WA:?RAZL DD5+%.!7D JGT<
PS@,&@YBR>(RI1UWY!#R.:DL]YID]4A=!J)&]QZ&S%#@(K.KG9[B"[! .-S7/"%[1
P:=^"AQ+<,Q"T"V;^G+^%%"Z*M0%]']!O;[+ .V<[B!<%N640D$_,'&C_QJ7M&<_M
PP: %XZ =;KO:%(N;HM"0>!E#DWQD63Z3GZ41!^,2[+LO5%C.&Q!#]Q!K=[G,U;[6
PW<A](1OH?>8LW8Y)'JP6%CAZ$MW$#T<18DN+Y!(Z1SRLA% @5@@Z"/R"HK686(6!
P[A2CWK^>BU<K9@Q,5*(.:)NP=7]CO9H!T+G9!#0'@$CHH,PG)]6B-4VUSS"V5WF3
P;'8(,<(26EDI,8P(GQ2\VN_?:5O \#?88I\G>C9U=\_B09>X[WJ2L>4MD]-?)C2Y
P1;+2:!XK!PO@](R8-^0K\,2BF-^":YWW4A88!I)]%(2P<LL/_CI10<^#XAM_264:
PBU+SI86H"35O&<6W/ K5M[6^[OTFA%A7H)78-"WOTE_H'X(2U%1]L@X@<#\0.4"V
P2[M5'P_NCE7VT=?@<6[*WM6V$=^47Y:*TX_(]9>US;Y.'*E(8>9?."S\D$?1'++,
P5:Z%#[O05OJU.,+MNCER[O(;/%"(WW0?E<!XDSH%@W82!UW>A!C'?*^+SQZ"T45Y
P]U\0]B,O9[)&/V3RU5\7%0"#/X)#>MT]'3._*T0]HWBQFQGS#$0V._CU_)(;%6[Q
P=E!]9-Q0$=5(3[_,X.M -IAI,K) 49 #-N">MUJ)%X$-?RF^&L>(4HRW 0S2\RV4
P*$[ON[D0)L=S9:9YV>WF,<@5U(.^>M,)Z24".P3)D[=?$=DCS.$<FZYAW)R[NY7*
P+ CMW"EK]Q$J45[C:H &<WT66,VYAVPY&/ -)\1TI-LLIIL2-]N"?%ZO>=@W[W-X
PL[IZ)HYQK*WT^L@;<U?:WOU(_;D83&1:+VBO>V66+1:[8E*JC!YYC<K*,PAY*2#2
P3W>S7EOR^!SJD)>0TB])?%=;?CJB4)? ]_.744LXS_]ABEY?RV-=\N2K7G2R^^<V
PY)P/N+MCP4@*I0*+SNUI1?^!8&4 -<%+;XNICYJ V:@#I4*TQA!L*B)BH;U*@&L&
P6*KLR>L/D_ O,C,H?[BJK^45 $68B539\I.2!%OZ,LEH7; <,0*XM'WMJ1M:=]!G
PBCMNJ+%QI0&S.@L^V]S5W^I\%\W9 N.G%2?S]UGT221L F;PG2'$++6F5D0&J(R'
P\8A+6**43-XP!FSTF@X9\,[>W\VJ21FY>$160J2VH_@'A7)%0:#O(F@XST8ZWED/
PS^?I#&<O5W@-I$)Y.V1%0@^VX28$SW;4+2"-B@_2Q,$Z*3@0$(!F19P9?G/-I$)G
PVZ]1']_*4[QW!7I0,L04#QM\VG1J9[)<5%[#I7ZZ@P*//+-)\@8>5>?P@VZ8 GY^
P&[[@7D&-RF^5"UQN8L'DPCMH1%;]8)L!F7<D-=3F=E,T 3/V5Y^6[-#;ISOTP1^;
P;W:;R=[7Q&Z2=LTWF"A'M$G>S^WY%!XZ_W*L61&. %Y!UJ-QRJ#D1[OYK^/"D3I^
P%+HVI0%.C,220%I(RK@W57>B&',KY8I,"-W\Z:%.]T#K(80Q812C%\+_ME0*LQX!
P&?"A<>-$74M7B@=&_6K'';[>E<G:,*SR9P]AE%_S+"@HHS!"_,%D+C>#3&V,$<G"
P32"ZL8585GSS<'P-"FL"-WCU*MQ$0K'>8F\^[&$K3J]<J8<A['IDY$]O#1I_7X'K
P,P:@^&W66]>E!-E..B3;F+QC, OT\.]-N$4,!$Z@>LC<-]2,WH$O\UO\<"X[ K$Y
PG[U\1O?1>/YO?6J:46HU>3NW</MEE4R7-+7J^*ZLM/+LYC9*V-I'_!#2=*_(/59A
PZ9>D]92@X8 Z'G*^BQ$39?T>6\;9*"] $W>EZU\HLG3G<*(4.?ZZ!)32N+:JUIT9
P[[GI:8PPN_SAQ'-%LHSN&27X_-=@C^LNZH'>C%EJM#E%W3Y!MZ_SO$A1+:J"L(;G
PU$#WK)J=KL#.B=H*D<$@AD"6+L.%(67:Y5/7K8)&N0$)PM^<'W'3W!/55OCZFKUQ
PG>%(SD%_?237@D"!ZS(!.!]Q.SG.S\)8JZ7&S;1MP@DLM-<#NAU_J?NZ[).+TV#7
PXQ$RTG7YFH':,EN=+:,P%99-;)LH#<=VVK0=8WIS--J.[)0O251</2_G//6^^29S
P[ZK[/.S" QW9_ GN8X/Y9:'(A<&=?XP+EG"WEQ!^>I3*:NE8Q%J55U4;_Y*<K>[/
P>?YT0Q#^(Q>U0IN'//BZTI'XI6J:!"$EEEP]>G?<5<+ N=\9E,$?<X,Q0EI6A>CX
P%4!9DQM3:=5]LU[6K,Z<1(:/1'HPTZS_!%\S,30BJQ!VG' -:+DNO:"SI>WA)#SX
P"CRC@KZXE;D2F.]CPH.NSMP5WS;&,'<C)]J2N%,.F+ZO4PL7F^?!*/ED'"[^K\3R
P/"8K9AQ237%149TO-'=\?^PY0*.?NWWV ;CE#; OKT<L ^L&>LF)M_L$1.J#2$4M
PT7@,9J>YHJ#(NHS,=K!>4>WX;B3?+]*SWB8R.1T@KE-F]Y\:/Y8[9>Q)L[($4"?5
P9=;(H&QA?_?9BJ#&/,7\7=("TBU<S=#,DE.&Z!B!I25H-%I0 SCA%R]>LJ+E1YWO
PB!?_)_:6-SF$+0 HLFD>L"O=\:)H$\V+I.C2Q.O%8(A@[Y6 K;79Q_FM7>6]KP#L
P.C;<O;[K4$3TO(DX^8-3WODHFX>V0-:H 2@]9Q_RO.-E^Y%3NSEGYD!KH1Q^SBWH
PW0]I3[L86LS;R_S"W:JZU"KS119?\CP6IW?,]NWC^SY#)8!92K.QD5]SRB27^S,7
P:1*F>W!\\<T(H2I/RZTOT;R4@07;&O;0^S_?ZAX=*L/,<U7YN1,]KJWD5VTV1B+\
P:?Q$K@63/M[.UD$#UQ[7)\ C*B"M)RU=Q'!^H62AR"YW,3V4DI ^!>TE!M[!0B&2
P?0.P>'+E#NLR@?S%KP^M C@L(DO=TIF&3 LI3"O,W@KXDM](=W"-,=;AXL^K"O%"
P\0]&,NR^WG+0C9<>02*9G>51+G=]75O9C /7)UXG0".EV4A>XW6UBMD6#9'?J@R0
PR"?:HD"AZ(%MT7AR0O7X_[@JTVI_:GM ^BA[-3<S/2NGON(XFH$DZ=KD&3*.D OY
P-(RQ^3MA%X%92%USLVRM-I:2YD*IK; B(;T[)V@;<O0@X4Y!YU?8"D6_YYKN3*9J
PWTYFJ=%[F8C[\% <X4*"K&MHZ-T-A5Q^FWQX3['#]W&C<H4=F"+ CB.B;!W>$A]I
PR5W..AR1LL-P3_S;%!N$>]FXN.,/X!"W7)\GS\XT\%'?\$H6=+)O!XA;[!GNO.X]
PHBP(-[Q.A@YJA.^9^!MM=3H$V1K$%+EMT.V"S!_,:)U!Y!*%@W8O AA8!?LX9*)G
PXB]L9=-S%UA9OZ=EB?=8MI,<H;U.Y4^710I\IFGFJOK5YI6ZPBK\6,R_[CY-"O-S
P^X(S/E4@EW[I2&RG_<1@SHLN #*GM-T3&1T(WE(\A0EEM\07\(2[J+W(RUUAR#+<
P-VS?%E'NJ6HIZ?G#:MQCV=0TU5FL^/]E'+8K87%?DE+1,CH*6IC#[2!JBRY/^[#$
PT4*_4P6!BT< #]]*ST:?/Y9$\*A3-6>8-2P3B$C&W2[);!UG!W41RT]T90B.4F-0
PH%XTM/OCYOPG>HTU7;I*7/T\SB7,...>]@T07W6)TPQ2871YOI$BC$,YK6<J4N^4
P1HL@%Q7O&Z*D!8O<',+@:"GVQAKE=VJZ8T>!VQW,@P^)5_78SJU+0^V7.52'5 U+
PAD#UR/Z3;H3VL_?8JE8)J;I!WPX+ED(';##NR"6W.#\P,+O3#<#0HS)%X7CJCFN<
PBF3J/E_))5^DWNJ><< .I2C1L" @F_%=7U-'!CKM^<"2='$TV&<([435RF[" ;[O
P&H-*S?HP)N:77SD3%A6YLQ."5KX*VRXKR$A[$?M 0B+$TL03#+0P7-DA=14C./OR
PSN%$W$R)S=JW^G)8J I]+L+JBZ0C+@8[,8,,&KXCVN8#R).UGTP55Q"/R=<QGQDS
P\+OE"2MH316@9Z2YQ1/#:$HR_$4_J4\*U2'5WC=SVI<3=Q57=4;UEYNA8B6PDML0
PVQ-3>WBA']XX^K\3NH=PR6V/W#H<EXL$3?9?MXDH0I5V8YB"JB*%[,7N'DHA47Y[
PU46_2RG61^=#T(]%K105%H_[MJ<P'!"$D/93#ER"RQVV\62RNB[\/\:YN\,K3H"2
PY)<!H,9<.B 1G/-&2MA[5FG'<NL,(0B ,3B@E HQ9$6-<V?$<,#(2[ZWB=JO:>+(
P'_9,\Y04\GW[]9B3[?%OM4:8.@XMS#V+M!P.;'LE"KG(BP3Z&Q#D9/ V@7H5>+>_
P3V,W('1K\TE:M*BAFOT@EJ*(#=[F4M)C K&90_@61:ZW2.XNT8O) 85S-OUB$F\7
PR"%9D]_T<0_Y<8P@D?A'W"87?>TS-YC@&1A0!(0?L:^#:9L=O3=W6LS=3':4VD6_
P96YML9F\UOQFI-SMP&1O/Q=>Y^!""PH'3C>.*LPQ$#L0:G\QF6 $EL#M).%,Y>?T
P[+'3T\+@DI"8YO2P:T==]9"L.244-TYHLJEX-CX+#IV+N4["$_HU30P].VZ.HTM5
PPY(]>8>7V7C_?L]_-+<S>Z+Y/O-(PE[G8XII%3?($<;3.9'[F^\^LW=Q"2PD7G$J
PG%:9MV?0+8;@-K^JQ/_EAU7I'9'ZYU\]NMR8\W0F8UK#L1V8QK2=J/4->LM=DK:%
P4?7($"X'G3'R8/#]#)#":JWCLGB1&UODX+RBGJ&/W\Q@93)#?#O43KR\V)T.<Z/Y
P/5Z>Z=1 '-?^P2G2T^Z-1]&A("6XD';WLTYOPEB[9]_#;/$Y\<KJ_\34?U=22C!*
PQ7U%B,]P,.W/^QC)*PO1?C]/18LW!,J)<VE@ _<L+I\Q*++>&<]+@2\J?J2ANKW(
P+C2]16;FM/?6HS*AATPJBC9%E5^V5;)++QQ+[E*</("&:-)F:DCS<$YF,TH[QYZT
P=_5*BF%S, =%D^Z2F_*L1(*Q.,T@\EN7;<' OD=^_FF1@MS_7/;E>IOIMOK9*F\P
P0M;/G+. PMXQ#"%U(?2T-:* !YW\:9HQ$F^R2"I0L?:RE8LCOP$UX>9;U335(+V4
PD</I$U4 Z*Z[78?><]&L3X&57B'.B2TFJ,L9K<-OO$5L,Q-J*&K0.'0R<?F@A[<T
P]TCXW>F><W :'MR5!43U6>"90A[0Q+KA80+5?&E83K1P!!V6HE6 M*ZHGAY>N6M\
P%()E/D< L[L-36)^>^//OCC+1"U5%QQ"G;'*8I/8SL>N8'(>4%9C5)D#^!*ZA-:$
P,W-1Y6TRYEXD5<M)=:'CY&6,A4(RXE\I74$5]XS5M$"0#(AA%CLQW,YLZ]\N-U'S
P)I6R)W1"[H Y:FG,5@P)%^)$CIA$^_ 0(GT@ME,Y@ -K"+& [A9W8UR] H;ZA/_V
PA".Y(V\/<I^B7MQ@F7X:I3F'"Z-RZHYAI[!M-#(JC=W%C$9BYVF_S@(#8!\Q9NC-
P&[L;_XW/7HV2C.[E1\!#4P1H N'H<DS=L)O&A>+6=F";L3XZ0L8=MW)%"[\8G+OQ
P;'],^RJTR,TEPEW'*L]F4F'1\V28CK8V07Q&6LGOYZ[%U@=QT@]A&+MB(QIN]CG>
P0LPV(G@MSN9:/E"FF'" (.<$^6^*&8466'8'T.Y@X[D>[76'G_<)+]+[B%9,:8D>
PKW%?^E(&_L27E_E9;<M6WF/AV+YZWAY\:"<W:2MX,7,\3>EEHZDR7"G O$6#COE\
PP16GK7M ?!VEX,^/:^DR+@K;9S]_XIHRB/-UB\$50S7Y!$WWSXM6_,0*/B;-49T.
P<>C[3&PZ4EQ=!E2XK?.0K7U(7&0 (**[/;BUHLMO0UGST<8U>//:DP 6.&VZ 8MX
PMJ.)I-J4V-GB"7C3PG-)8W *&=-:0SN_?-OII6:%50DC+1L$IT49/= <CS>TA(JZ
PH^#^5<7Z9L JD82;M5^-I6A"<HX5;P)N.HS^D".Y6DZ*S#E,,!%P&ET$9'C)N:( 
P"\^X!M*K,K&!>:J(M'!07V*770.MN?1&F/)BMPH28@^E9:M5BN[# <?M$!8#\$H5
PH1BUVS/^P1/[>6?87_?8V _N>Y.#N.1==B"*- .5I73>8ALV8V4@IYD@AV(]OYPY
P[VE DQZG+PX:>#K['GMS@N+=Z:ZO>'>75U-.4/#Z+K'UQ5LP-G"%84AJRB_+*ST&
P."N=NTJVHJ"?Y43E&+$$HI.SL3F";M64[Z*%!@ND@Z8!NP&=KAS75V/U"Q2?DL )
P<,PBKQLAJ7+T'SG3'L>_ ^@%FII[VMIQT[H(3(*ESB(@OQPLC:HC]C221%*NMIBZ
PJ("]#7AYU5G85(-U.JA[Y<9,:;H?N??LQ<2S!JQO/]+6@+2;,<KN7/>&23OQ6B#D
P R0LAUE)SUUD,  -E1JAJ<JNH[PZ#QR=J>:D+Y7MK+?P^>&'8YDDXGM-3M\9X6T(
P\%8[2B>037P7Y/@_K>HI2#PG5V/J 5^E%G#Y_<PVQ^JE[R!1YR&,G6N809V $Y8E
P&?G@2$AA9XB-89>+>))!"(I$\).*;HDFBQQ; "^YPII[^:6?;"O@7)Y[@5U*4QIJ
PWO%02"9?*J0]M.\=Q(+19M558KV+YE+*6@@4I8'!6YTT31 78; #0.P>MS<]QF R
P : @2'=UOPH;[70F''GZI:SL X1,]5"LHP_R^LP)P(,SEWP42?X'^7B6CO/PO#<0
P?[R@#;EETE@8=- \,*5QQKU52F>*1B+X!^@B,0&V*%[W1_5;Z1MQ08O$)--HWR;'
P#CD;LGGRUYM%\WW6"JPLSS,?J*6NNI;ZAM[=2>.K2R&[.>)\I9]B[FI_HR9+_!?A
PS?2_N]RZ1G BA<D=V7NUI4UMH7MET(&ARWIOI;BS(+6WQ&?*$8,%.[;3W(0[R2EG
P>2ZR;U ^AZZL3B/Z4\TT&6',UZ:*A>M?[^N[^)EN</%.*64"S,108GN9,?F!!46H
P<:J99O<?D.)1CE;V^"H,PZ_"X0@#[B)+]L*62-YI-1NPK8^:.4XS_N3AZ^2(^ 5 
P%W,_0A2PR_6:12IW'*NN.K:\Z(Q/8 )N$JA/=%3<4_&W"Y"KERQF?,F([?+Q-)T\
P>$#A#@GG+D_KWWZ?N#N=8%,*[7Z-1-92]@1#P6Q<Y&*>S((F<$O,URX'Y^_A%AN(
P! %Q<,A,3?P./2(:DK3"(;%&,XX%=&]JN/@WS-K3 .6O8L+\:(=_2,*$Y&;%=U%J
P:4WGT>L#J4%HYN:3N#=*9<V2%N8-QA\<!-5,']3=;O7)6+ S9-IULHXB;0BJ2CY'
PZJDZ$]/G_BXJ[*P60SBC 9SD_\9R(+UXT@=#26=Y/K3#4PJZ("NB87PGDX-UURW+
P!_/'NQA3 T3;\/:$>JU2K/@HUI:&NQHZE@H,W\E11IY5F@1,L@V/:T3Q\(&!%Q9[
PNL7?<[-VM52=L #Q?1'Y5;W_R/( Z";IEZ[UB<VSLS+A[]$^?FM10HNLQE#45TN1
P,B3&D(,8G:[ N9N0ITMVHC 5\(M+KDWR-'N[5X2]/)UJCYD26KQ '7;JZFT3T>T)
P$7I('JMI69D!!/()%B-$6\)YW8!PO,0G\(_$'+/H-ZW[&P:7$/YOV\MUZ\3'L.8F
PG8-V8UP3-9*_'D9/T[F]"?G6&K^+5$KK+/#ZWV^.&*%0!^_HX+TZ@KWN^H#'K#9#
P]?+F3ENI;_;D6E&.%4!@M3GUF/"=&ESVTG#D=7 ECK,2[=$-)>Q4[OZ"N+&0*29Z
P1A[KSY_L^J,8O-$8<"A7/LB<&:6*W'*3#:=A5KM*?G.ASFH=0*%V/FWXYR_PF. 8
PT%'PR+BPV!]F9.&H;H&R8%"VX@.\>VZF5Q P=)4Q@*4"/,D^Z&(WU<"0B [Z<C#3
PQP>>;G_(8>@2JO.CV9:$(VR5#)ULBR*/KDXB)"NSXXGWV7JUECLHB&]]?Q14_>V5
PF8^$FKD1-1,O(0WE*M9OS?NS0%<"9^?1$W6&.:OMJ@F[,==W-9AP8EJ4<2BCJ!.!
PF%GX%TU[BQDRP5YKW4#Z7?)9*C)R I/U$@%_<4?:OBB)_4XIGM+AM[7Y![/RZK$C
P >EBHU7_F>ZNQ$>;_^ZD]UM1O>GMYBQRB_26Y9T\[VD+-*HJQW+?;9WZ0-!2B_UZ
P'&FY5G!V/QJ1S:BMZT!05-@"_';QYE:XL;[:2>^*QVO]F+4VM5[=!TA,V3;1[*0"
P!T+6_/YG$HL'Q]3#]&DW,!DF.!"J$=)'CSH6DJX"O>1G9+>(Q/5<EP7QSSQ".)\#
POA)TOA+-T[1#0_:#F0_HJ8B*>M4WS$PC(U9 BWDXG( 9^IXVT19MK=TASJ,)=#@U
P0L#JD6E;H7.] _<<R4]1BDZ1!L-(.S-E1$7:5C= G&PPLC7?YYB+15^!W^.9C%,4
PS9P8$6:#&\NX?0,5Z!-[V :P@1\>0F#'YO.S4H57N$*<&+VC-RV2_^W;>\:'?1PO
P>KS+B8;F_N$,_R^M<'YT8[\FUOAR?$/,@.$O^6=6"'')Y;[#MW3:G^[1+MF1JJN\
PXNZ[:PKQP+Q,PI4VE3&E_".XNA]F9 TM03H)0;&KG<5,'**:!)*Z.G+ HO],?O^$
PY:F"L>@4*O-O<I<8? J7#Y,-37&G'/;9DX6CO)5.LMW!D/:JH9EMN(^HLA\4?9I%
PH^&WP:=6-R7UD\$4$'*E*#L'ZOW^*?+H_0N?/0Y.;<K'\ =&+QU[L(D'R&R<?%+A
PONPU76V1D6F.'RPRR]W@ ;NA.K,_<;82-H^C\_\ 71\) 5>-&0L[>P>]3 ?O6L#(
PW"Z[KIE'VI]7P:]^?M%D-S8TMF@?'T(&1MBP('/3N]'NHKF(BT]7@Z:!H"BS7STR
P>-O^GQPM"YU8C']C?';?@VG(F98.UFT'[$WHM>MN\3O<)=!>V?C&4PSG1;"PS7"?
PUHEAV!+TCEV]ORY_4]VW$YR*<\+W?QWRV%N\/9](R]]W7U+8-D'2;,H!&&Q)8)I]
P5:F<SJ76@.TT-,4" PM.8Q&#.LF* ^U=CT!8C$/8U:G*^KYI@V06;=Y6A@H? #W>
P*X(25B *P.%[='4(2$;K,EHHGKA?7//8PUP,D^MF.,\D#::JVG"BZ[$Q]I5(M?7L
P02!T(T BVO RC2P7^*Y9:;)",_Z3)-(*"WJ#/K][*(9NO[T^)=I]_4.MS5PPL&%G
PL.,\]\WJ)TR"=-U2 EP?GW<KVQ;FB9'@MV$;?*T/YL5NL(ZS&'R>P(:-<]/;?OPS
P&!(30HC+;Y1+(6//&LW(4UDS"JKI\[#<6O>Q9V=BZZUXFLW)EZ7="-:XY?5TW,\V
PEK7PLP5G9Q\VY&KYK\P<'QX8OZ 77#^2  9$&]7+4!D!/2XU8T?= 4=G/&2N).0L
P7;W$-U^1NGLDCFL.@[KT?P58\'"8FU" )8 )M=K_3(M?NY"3G+QP9R67F1+@U<LT
P@"1ICWU!%O7F)'"RY9Q&@T139>%PFV+([K?G?]C1=#TZSVJ#_^-[/.)>/@!&^ %6
PF\KKKM"Q,(H+Y\KG50)SLQ[G074J89Y^XX*QW7J.8*+I"5<F\PW=%OM1_U%FV*O#
PF2IEYFR&CENF@O6@[R)O:T-\IO4B8$E"%.7BZ4'9 ,"="4R5K4LZ\1>E$R;B*M"_
PXJJ[!MA-BV+"/-W;FSY/G(R"R/6,)9SF=7N(5Z3"X<![?KXJP1]9#&9JGQP_Y\RK
P5?86H=,N";!L*=GA1W7Z='_&=M'G$"8TIK3>T#2OJO,DG7GO7<;RB9Z-?G%(P?DG
P>2Y9/89N0(3_DD9QK#5!\.T6]2ZV)] YQI8;DE40OE8B(J<79VKU*ED6[H)#3"[Q
PU/![VI5;'+/P%)L,I(I>4GW I1S*RK5@!B;GX53[-Z_G8'!@3G_-]_ZS^CJ;-4G;
P57<@:)Z?!<@/L9T7++2\(>2R1&,J^S M /\ELFU7M&_:G,:O&3!3<ZM161G,/A%<
P? (N[+,*BU36W]IN01846E:#@DM>QUUL YX@?%F@@)6J-U>C^?:DY]YS,HVROO,)
P <$9K[="O_^S(3$')4VXUBRLS#E\:CYC@_;_^/%+;NI%,<OZ;;I)1PO@H2^_*(-J
P,)7WW6*_QJ\8#ZIV A2&6C;+:*HC=;^)W//"R?%8K.81D7X_^GMU0-/]N_.G7B3:
PC'[!BH_'D./?BXH,#!+_B;(Y*:RF< CK5^_W@XI.UR;XQ# /1#P6+L*!+=/(+^&[
P:AGE C, ]8&!5L&9B0A3N*:J_"X?IW?0\1E2NQ_"\UM'DF^\'V%X#[[6 #V?PA%Q
POM659LUF?%*U/(*3;.AMB:GJA;.-JT"W/QC$7/"9G6FG$-4^Z$K)+=.\.F+71"B3
P\9+N0L8Y(D,BMNQ?2>5NIR@"!7EH&H=ZT..T.18N)Q%O8Y69/%CWZE-+@&:J9;3)
P;DIWSM39'$8"^O9_X .Z2KV@@TPH%@OUKGH$K'XUBJ/R_G)8<'S-[J%"]I"[ED&B
PB%Q27ZSB6"IQ^#H"Z1-!1;>9Z?4;)XE)NNS#9&'(1F6+:F !-*)4_ [?%=QV;W18
PNNI4"(>Q_E$IQV]#-2> 4=NVR72&\4 ,CF6-2*:7,>2Q/,C*@A'"U9PT+;=.M@S^
P$;.YV/*R8::<0"H'?.U4?WK7&# 0A)#1M'K*GU\"LKMUED:.&?HT&:&*^K_+*[GM
PQ'@PQN0.4(<V*%3/@55;2;BP"3K: L<&H1%VR<L#5I&ND@4@^*>Y>3J,AFF1C_,2
PQDJ(XLOONO<L%8HD#%P+?GBFOO-ZQ+,] 2T-]1P!?'79-OLC?GKR& \\I*=#I!%B
P-1%(@YNAYR$8A.7V+092'31#$RZVXG_I[->5B,+>+6//)'O9Z#&5!>I P/B\$R'\
PEP9QI\P$,]5&H)>-5)B\@]4] 3OZ"-"V^/1-&TCIW_[*O/#NP$Q@+R0M-NX>\:AX
PS-?XL-3QQWV=J>KJ!8$!/ 9(4*_9<WSZQM9+Z[AV15O6'K47NQPOS%/05EF:BSWW
P++9DM7DZU!*6. C(L8THA[0O^/Q8*DHH1;.@$:6,SC4P=2[,#,!DM)8WHS1#N6R3
P^Q!VX-,#.H"K"+Q;^M!UXF*\L@/RA/&@0K 755.=%JKHT@"_JR?!>-ME?K=#A:+%
P&]V>90: N=C;Q;$N%KJ#ZJSO=Z0CB3WAU?M2P$M6]#1-8I)D"9:S3(F/4:F=G#A!
PZR+\U[G!F% =F1'E,\Q<A2,7+/2L4+ZIC3X$-JM"I!YXW.6'2+LMJ,! #G"((2%-
P'ZH^4WMC2G9YMTSD(54ZW^C3YI1B3F;I!S@7O28!!T%#PZ;HR_M=A24R]N@#RI8]
PH)2"MP9&__H"W'YZT2*!I)=E6#64\[^K<EE"LY#J$=2ALJM-O7)@@GGBH=Y?PX^$
PJ<X43#JZ$:E_AMR2!GV/#'GN +=<#%O4TZNK#=2IJ]7)L DYZB/W3#1N$WZE<27L
PX4AKSQ!O;R*S^RB,$,V!I093]VZK%3G 62KON+]48(["+6Z%+L>L?)&4I*'F"Z.G
P:(MELQW$C,W_$_T*HV@VN"T@O))?7)5(.?(HDHY*"P3Z3.%?DGM9SWT6@=6 W;WE
P;HPN6EB?BMZ]#OMUJ<$-471,_&0_J+9KF1=5[VLX^71Q]'Q25$KPK]TR?%K<R[S+
P\LE6CD5)7!S &-02B6+08;GH.K:\^RJ ]$%IGP^V>R_[456%C%Z^+4D[N,YPFOV6
PBWOL7,/U6<KQ*L,;2R8CH/4O5'.'0AC4(0+46R!B5NH>_)V':>WP->"H!-S*Q&)W
PRZ8GFCXBK1QP5C[<*&PXX<6>RJ[W$IJX^)'BD<O"*=K+PHT*,3)AA2FN (3*!!"#
PC8B-WBSMM621N?LA2O0\FSN/ML!1/OF<X*-:\4K[,+T8T8&U"YP#!52XK?1JI(MH
P(0W!H3$TC4HB.*H;&H4[4NH_ ,P'W=(2#G\&C>?(3NH]>WOH '8&S4O-;1MFWA!<
P[ =Q?V["R[8("XJBE/8U0=ZX'NF,P5U$+E;:P:@+$16R26L%=$/"::3]7SP>&PBH
P!(4-"SW;:T#6+Z*<H.,4JL4=/)^!3_I<T;L5I2%$6[&L-V.9]9>AR[QS$SX/U%\G
PHCGYG^E.#X$4.N71[SDN)_]"CG$ YFWQ*[$7^"9T0$JM>SE/*X3:RO<UIE/8WR:C
PVI1QTL(/#0NSM'[W LNMW(6CPV"A=+Q*;CGO.J'&1?DFF=44V2HY"NP8%NP57B+Y
P/@_B(R-(2P><C4ID5:C>=$!4LU[2!E2\EB]/<B)50MN4@*\33[MH#<6:[#!W0IN*
P_G=366G<;PO'?FBEL3QRZ:BQY$ [AFX0OBK'GCYNSKO7D-/HI+^)Z=;VIP.I&)LP
PK00IRY<N!B9>+KQ#8+)@^LE8UO *RU&/.00KRL_6> XX%KZZU)!1)MY[6,"K6@7 
P+O-OP//&C7B+!4L>R;NFI1' =D_,]Q^4H&B?5#<Y>%\C_4&I3RLS_T1B'B;=PG;%
PZ8*.FLO]!RK_K8&K?[Q$NHUJZNT]&@20LG1QT/GAIXH<0_.9ZX$/B+*D.&\D5V51
P48:9-TTUJI6Y?,,(,Q5'DM+,$&-J XMP^M 7O* ; ^X2M@9?V^,&0_H5$PFMO/>5
PC.Y4D3$TYB336Y$A7SEW^5:8*V)@2Y6O_- I:T/\(P^[P[C;0TZ,'-=4<V?0C./.
PI?63TE'!]7I7I-WF/+C<@G#$2@/ ZZX\@J4K*11%+8VS\L#0L&]XS'")\(T!(5(]
P6X!]U LC+ ]6OP\VZLR]:RX?"\L,>JQ<?@=C7X8Y'=WZK+JV8=>JC4ER#A;;2;QD
P,Y+Y3'GG6_KSO@YD\_.$*GE0I61N><.'J[T-'J0_5Z3<M^_[[BG8+;BO%5T5,BTO
PQ!.*O86@[N0Q]>*W#6+TYL5 L4RY[$\HZ><(5_HP*#=* -6R$@M<J#22/HU/+I]S
P,?TV4#[LHIV1HVQ9AB\'\*YJ=H_?Q_NR*E+06C,N17G[=J$I.21;N2T%YT#!8@6;
PUFK#MK3$YL+VMT*AM;UC5GI[\X$B6G1&$WIPT* %>="!>W,R1MKF\\H%4Q\0A6:Y
P+WN-8P1PO\SDE\6F')L\*U\VU/ZQ;5SLJ(#A"\'(#E($;0>5@/GB(Z>5:045_E3J
P_)<]8SQD/$<Q@KQ<7%_;'%5$TS5DJG(J7O#(4'_>1EL=EN;AX.8[?*/)>]>*3J:?
P+X6@Z#+-6N:H9PK!T$_PK,/[>0BYZ*H]V_,Y_:C[:#WDV"O<T[;(PI7Z;K;O'\T?
P1M0!L"&HOON>4XEVY\!T[GO+H09;N*G@J]H;;^UH)'H88,CN-T7J$.AH9^5+EM7?
PJ1:-@A5N]J $9:=!,F:4 +"B*D!;< >&&H=(IT:4*0^ZI44?4^(']\+AX9*IEQ;R
PC>.%*+2$[%LFP7Z01H)!8]G<'@;*Q[.@C9U'4JV()'%SQ_V1))'D>:"9=(J\]$XJ
P(RH+H,=_\LZF(T$G:6KBL0W:B5Y+/+6_7&5ZR^H9TB]4:])?;3 @QTQ$D!2'[KKO
PR6"<O5X2_XU2%$BELU49BBZ0SQ=Z'4P @0":E(+'>.C>*\=5'U_/XHI6V(UHN!I:
PAZD_Z@6K8F@@!*%S :0N>L=]]&0#A[9U8B$ A,-JQGZXBCNZS2@O(54YOVG%R;+.
P/)5+L'I&I4%(T6UV++C;9L@E^\$B=C\7[@XZ[1W$G(T B4?J!ZJ4Z24E%8#HB6$!
P_(W6YS*=&S8X0"GJ-&.UE,=KX[7>@/7?I,XW+X@ FM0W.EF+"N93&W,I3'RGF387
P/BRL5VK<'4&=?+GEHS$I]UKYNC6@9C\_W"/PIK=% HP.@ NXA"&2_W/76;5UBMT;
PVW%1?EEO83N=<@RVK=;E<WRT2' P0^NW.;B8WZM@8Z))@&C>5,98K.FG/TBREM+9
P&3$"&J, 1HRBAV9 ;;JW: (9K;:L-;D]*>[9?^BD3S0TUE?_ #"-WN>O8\<A7;#"
P9>] <&^M4&7JG K)KOZTA+P,9B5CO<S=<2=!JB!NR/19\SDGC)3#IM?6__($,/,I
PG(V<V:BX: C?47!3J(";/7C I1$90O<3'4RD/\ZHXQ*ED4UR2:TZ=H)-$WI(*-,F
P][XW]@%-ZAH(2LDEDJ'6EL&!4Y8# M=(RRX#1GR[PA-L,@]'W7M@#VJ]AM_/J0@R
P^:CTSJ0)SX/U*N3T>8K J6L?YH/?JDTK(AY@-E4 P)SO5:B8_56CW$XK+AC)DWTB
PRFY(T#^* >>)6,FX0*]?]R.["YJC<=D2Q(8E2J ':<<,A=*M7@7GQ8>>FW\[.\['
P[R5+UH76K%906"GZ,S@GF&U3ZU>G=)R'?#->/?HA&@ K#O9KP?A)>8#2_L<!I$V\
PW6#@Q!2<NID<J>I7=A]G5(8"CCWF>(6R<WE_]PF&]@M4-;=8AJ-P 68\]XHD+)E2
P//(.JK3''@0U9D@2;1,PFQE>HJDG=5[J<B"2SK.)(;2V!&_-^HKTVI9B:;OHNP .
P))%M*F?R@=4JV(0N%"*17(Q*\6A@Y/$.ASBWXT?=G]!W;8B&7RMN"D+7BO^\*\++
P--F"1X\@K*<3Z5)LQTMUG^ GF])3F"$Q_*_I4$KBYZ0>%V9MI=<LKMQUA>8A^G-%
PI_, FQZ(+'].8"\0N8!/"?(*0!H1G>\@/P7ZUA&QVK:26=XZ S@3&2*)&/EF7/^ 
P<]* LU3Y*X7T&&F6M"<WM_E<Y@+<U[-A4/GX24/*DF5BHST>A/0LX5(*H4L-D$P+
P);N(A"<4.15\O=H RRZ^C@YRY>>*:##Y 0>C<O%*<Y.'UE=OJ8S42IUWQM&<!S\R
PNY=IZ)Z4B$=R:*8"6-/FWC6=SEZ6RA_<4P0-I^'W&SV_*2QODF<^OVNJW*ZM 8$.
P=-]!(D5+ ^'91=)X^<^___%A5WQT<50)/*X%@[P)H":<@8Z6IB?(=@9ILP*DGT^2
P2I8GI,OH 65>E(@2HN\31E#=S*<6I+QTJ."8R"=D%X]O^!6 ,5I-(FLD3DW@F+6G
P961;2 B&U +Z:!7CY%<^)3\<&;?KTSU]G9-O5O6!I!+4W0;^8R0I!GYT[G9T'P2!
PD(-2R>@?5RQ=0MY0V4Q?0AUA:N12B8!^4(:2'3M0PF.4UN\XNJG4[C)H(E /882^
P-5H?/2(7#%RO;> T'[[52>$%=NWK+'O5)G1=M1XU1=G&;EQ3:U@FKNH?:%X3;T0$
P'^W2#"1LR/6A6UY,;7C?D[=H5AD*)KJ43AH T8=,C,KF[](,-4#^N:XZD'T%\R_1
P+6*"-2?I8X">+LPGU"B:XQ3Y9H]C^;?W2>8HJ[)1$PP^^72%PFU:P4/FYA&Q2Y-)
P(/A; U:9(QI_:DF5-3*^NP1_@7R'U_(O$M?R)X=$L!0!'2\PHL[S<G.JN6JBY>F[
P9Y/6$TG+DSU_X><3 Q.B2:QZ[!OVDS\6T['-3B.>FKGL)N&/\(K&/<,H/&6:=<ZC
P5J*;FTG<F#]*!92OAQ@R.%MZJDDMJ@DUT2H6))MG(/B*L?U](>3G&9T]HMH0?4X\
PP* @*L5EI5]:0G@&89\Z  D.P#F^+"MT(=#%H2UV0(GV)*>O>%4&3F)__NEDZ4,'
PL[[*=(,;<EP-PM.GCJNN[GO&;U5()/_!>*]W#$]O?+XE:%=F'IS+AK+U%8K1(2$+
PC?+-^%.4,GIF.HWDA12\V'U8WH&$]J^8=$_&9&0^0NS/M L9=]U(#>S4<<9.E?.3
P=.G]\"YYY$,4JR (;=ZF5>5DQJ,+ ZK?F@9O"MG-90X57_5>$&X";*&-HKZ1^%,!
P(NQ?\7AOB36J;WI@8*OBBT3F1P'GM#'TGB=#[R^;V2O)9.[;)32JOA^>NNZ<=WY[
PS]?&I)K"15Z_T#(Z &:.R.F,'$/6M[L2)%S(O(<TLE !Q%(ITDLRT5>\XBO#!V@O
P,/XQU88;7B;Q V=.T2%B@WRW.,5DNLYY<,.U /:P.U6Y>X-S[@?F^/D8X74"F0WD
PK#4637FU?L$K+().82GI3T6X;<]8F)FOUIJ"HU[3L6#BM-<N@A*?.CY:6W],$V@?
PS!B4[(]G]K[,>7MB(C>$I5>QO:Z#QI0$,O!&I*\D<UWLL>"X19FE92ELLL@$FI=?
P-WQ\U$]P>)ON)BS]".]XL6NB4O)['<%9UK.&D:DP6<>UX]M_8699#7RZ$\0A:!KM
P>6:*]:0W\31X"G<S 2S?Q].73.*3:,IRQ)LCAJRI62$):;G7W4D)&)2H9)=SXR+0
PM+(3=Z-.#6%)ZOAS[RGWP?/Z*LCQZ%BV*AIHU-*6<0;9B<\__11=N]0UTROE3<FQ
P4SMSTS3GI"X"5-ZC?J^:J.EX97YP3VIVG0]%PEIY.&H;OB<7R_+'=SV55Z:+EB*O
PSA5%P!DE2L GV][ A'N)R]<CE;#'6[=1>DQ%DK./V(J&C27(B8>7SGM"!+51&3Z2
P]TS <NAYU6=YB+=7*7N7B$- G$F>@45GCHJE,9L4*MB58-VVBM]LX[&W'C\"3W8'
P8"X7Y#'SIK%@MM \'>,&\Z<.;J[7J*-6Z(_%K+V1*<\ ."Y\UP-%*4 $74C<*"4O
PGZ?9?Z0O3<M&Y0^]?VCTH[;\^%C8QDF(FI81%T6>$0EQ<4-QXP"O#BBM65Q9;?$<
PWY7006*HUZ^ILZ T7K*=,//2:MK&A+:AOS?1+3ZO- $;\=%DIYFC_L]OO=P1L0[K
PO(,UM:KT>ZU@+[CPJ6.U=CVV*2Z'N$1K2X<QR22.4O81^LSVLGU/PIAK'=NXO^[F
P$V**"OP-GN(OQ2>,@/BYS;/5G/0M!P_8A#S74+C-HR.\6&:-VS-92IHKR,;PC/Z$
PM9"7[3EI&J7Q:!24"\1A&V_<G-Q')P*N!-6^:H"*RNFJ,V/$_XQ791IJG1SPW#VC
PZ?295PL+]N4N,G8%L(#-$MJ'L9P6E/5 CH=BS4*IJ5I,+(EI,G'HZE!9RCVCT%*T
PAV>*B.0Q.HH3U[3Q5-02*LMM4/YHUT! .O>QZT22G[N8[E;1?4F/\\7;\77BO&) 
PJ3(9MJK]RSB<),3\:(P+. :&#GOA,R'8_,N6"5L&Y]NS')O.K9)_CV\MI:;Z^J;-
PF^\YF=[)>_]TT%-V0!(CJ*RW%9R*@"%A$M?^J3",-&0.R.[RPM61* [_E;:*17'\
P@HR26U#2%3H^4@!D)L#A9]3;129+-J'L8_?527_YA_6%2YH7VJ31"V4E2][:18-6
P%5Z<\?>/X-^.+BP$ (#V<.NA>$0P.P=U]*TSZ)Y3*$7LB[SAKLS1A6_0'0?LJ_-<
P79/+OQ4,4+;/Y-8C(UDI!EJ!F$U#Y.2Q5]]SO,KI_&)V^ELW&*ML[:@_NR1[^"O[
P.4&A.CR\2-Z+."CT/U#>9MSYWOWHJHL4MF8D[%5!F!O=_/$V"UN54\,2$Z[<T?1X
PE&E;Y+V;7?>/ [I)T6(T;&+/Y7],?*'+JL>!2V@U64-*ZHS66OES%LGU$(>Y%R<Q
P^ #87':.^E"<K+QP.M56'W[P>9.5 U+4]2_55-A=8>P5CH1B06,'M$M@%PRY5C=*
PUI1(I@7C,@ \J"?NU8H04WR[-0R%NH8+XT_DD-USRG7\CTKXL]IV:I-T]-5PSOY5
P;Z0/@KO%A.2:\($0OI'V]A5F=):-C &)>IBMWAC^CBWRPJ1E,4Q00Q+A 1/Z;]N<
P2@U:?H$R0MI)>]\J<V;%QN-V>OC"74 ? H=B8(:XY-:6EI@;02)35AZ$GS5V$.=G
P)C%1"'510PB_)T3T?M$Q#8NTB/]"E$.6RA9=RTTA+O#*&^!MG'?>\XQ+7274T[K>
PNYN$SKCF>#V=^;.N2=7D1P=,+[U*%T$"D"-]$ZA3X!\\0[HKDE<KR:T4'VI 19MA
P[H;:AN SA]*IUXAH5S)#/>S"X-7XZLT3B@8=9%Z^P9/8EQ$&!4)6R7$/J=?<&_"9
PM9W4*P0\O8 RIEWQZB"=-?5H H^BWFM(];5\WL,3CFH-3@I&F74/[,^M9:F!XFL^
P>:OP+^9892@35CJQ0)*Z) 4KTZP$VBGBAP&=85+W5T_^+(VNVYR824!@0C@@9*SS
PL2C(4&R4/KNN;A&"6[*0:< JE8GX^%[+O^3Q\#"G1&?_P$(W[>[1C;W#WTQ(Y2P;
P)9$J5D7JMM**7?6W[WZHG^YM;+]J775[M%DMD(-,(R,QW:];<RS_YKT?_8&/O4A0
P+> AU;KW?Y6N^,'6U*C0B@$B*>\S,?A+!0*:B..)LV\?P6LWXGA[W6>K4$N,WLUP
P_RXRZ/,"FKI[!%7 <SXX\C,_1)W2XZ:37+(T.%$&VI5(4S]QL:EVSN=9CPO5A+C>
PF<LX1,7?>)OQ)$,)%W6Z.D32_:Y.=UOCN\BE@F%?.]"6>HOB9_TV@^Z94G31K2BC
P94"_%36P55X5GSL/@P1&4Q9*5=["5<U,5X ",X_W!X.M2SI@7R9LH: .HM[K;]J)
PD5GV($L:-"?@Z<R%[C_+^9'[Q4F+"<5%E;K3U2ICW3_/"#&Z(7*._T5BXWNEYS?F
PB*B;E*D8@V@7J!P)E;I_B&_,4STC6@:C,-U=W[8,Z+20R6-^]]A,=<?RZ3D..$3A
P'6UR'1_J5V  PG[RSMETF8KO*QPBB22I!%R'.>0!2X.?1PV(VV#O1E$4,\ "55EC
PZ?TA\$"F]G]&="#%+,"$B]P@D3;1)EQ=?*" O'Q3G# #*C;@CWC=NZ!H>@44=G#;
PIL&<&%NFN7M!Q1%)L<124%FT?^2T< VHG'-W?)O/9^N=EN_PSDGF+=(B//%27B/<
P52UV<[ 6K30[.Q?T9]Y)J6Z\B99OA=&D^7B(YN:-^93+ II!_89&CZJ9[1OC4D>S
P=U%$O>WMU(D2B!]$#RV>R&8H=.PEC ,O5M^9),99C6]AQ]^&=J8J.5@A1#&/9IW$
P)O;M<UW\DE16<7*;NB%_!(L*Q&IF;:=_.+\44AF*0GR7HK ;<T1_LYL+X@ #AE_#
PIAI8:WO'Y!$,2YM5T&J%-6DCE P]Q2^[UPG]T: -W/@&W_,]\M<HNEK:YNV(0 D]
P+*6;L. Q*L"/Y*F[%'WOYEM3U;HB2]V1MNNK\UE.*7MWGK,H'$?E)@26'5&BII.9
PCYR0F5YGKDK\A:CF5?_6AAKN68@Q\EECUM9,<1I[=[2.A(-!,8RR?K2*@^XBV]<O
P?FXU::^?ECM-=>GD7D:S/=9WH84XOQ*5AX)L#,0O_.E*YS3&A."ZK<E=CH56)QD9
PDK+M2,_3P'#1:LM\E-I>_?N5"'6G(X[(,$WJ!.G"O'+;6)(&'$%G\6^IM+"[]R,$
P^[N-!%QQV#<,;'<G:OU;#/ >G@#-I\J+YK;_&<P6RXD,I(%QO/KG2W#O$'#P\2FZ
P^E!$^XO[EGAM^/=K+.0M8U<A-5%&DK;T%W(#MI^UB"C#>?)03E_)EF.?SY\:E'8+
P($QD,WJ.[F/XYY"$==N&8,.1I83*Q_D@_ZY(O#(-++L+F/R0JIM)%A MGLGTA1'!
P*2,S<_0\K8GT*(8QAM,EPJA0=:4$K?_R:+2^F2J09TU),_F-R8'P(3\9\BV@HJ8(
P[8TEU^GRF:PK*DPS&%^R_B%$?9Z?.A[I9F*2$8MRL%'O[S;\=<'X.W^],OD?=37Y
PTE=%B]>/^=K9DB34(J"S7>&N&?%Y4 !WA*YO$,M/@E+^$0DE34*H/ )57TO2JKS*
PS>6T((7R=44,U=#@_1OKO'93['04)8>19!09]P#(/'ARK=UV^5N<FQ)_M_X)N8;4
PIO\6EEORN_M[/]4P0W%="*.%S].BXS+4T;2^ JU8MXMHD/^3'Q1Y.U$%^8&*+-W#
P@X8;#L7.X]/1=T4=_DUN<S:I%>!E7?">#&9\G[S1XHY!ZCY@'_6DB>&E^#12E_G*
PHT]3.GG1("?N,G:MH15*U@E@T]-[U&L%N& /VKCZLQOS=.K&EL;DD?-(S?PQ"JQ%
PN32/D\W$TPL"%IBL=](YD9%!3A:M] 7-5ES\H$*#+:'_-9<=7NHNK=>2P] ZW/8P
P5H_:>\QWA]?0R%GU/HAIF$,7EBW#P\Y!N,"V6\*BZBY::[@,(9Y99&DLL0J+B^Q?
P^C-BAXW"3Y-)5#,4;X]5>W?(/WT6N(=79+#_[@==/E5"_<A0X %4D3DL TI@F(7^
PNP 3[1L)];TF%;+YZ>KIK'YT\!?]AA[CD^U&:"O:L21IIG P!L+6N',0MBC1?P#!
P7,=.UJRR4/U8(L<),'<!A>!I$P\<*K&I5118:;.%BZW#[R(8^(V./%-;_(1!7O8"
PU59UZ9<%Z[QR[/G/9R%K6V^P[8_%/,6PVHQ8-[O_[S3C%!<)8BS;N+ROJ?7^K8D@
P;)&%%JQ6;G(G"12#*)D3,2J%8)9PG([[-"?R?O2+9S ^A20 '-[D_$UH3=Z='#\-
PG%P[+Q5>[4"8WE=_'$#\ 9Q1Q;QK.0._9(V@GI4MP,IM"6#4-)>BQC$S18=KSKWF
PM??"J<_L,/[QI'ZTKP-FF>V>JZI^0$&M1HE5&:TVO5O[_P8,+ \65SIH@8@23KXP
P^)5-R9M2F]TRWU03S3@OHNYO4B'PDNB[[X:9-ZJ #8ZI+)=M*+ZP4!*2[Q"ACN>'
P]:\-[BT@EVL^<]OXX4M/\.Y(+H"9B*R!"II2\488=/_7.<E3;8>!B/EA+H)PPWVS
P;@P$/)),7D<MS6N-9Y];P"N%_"'U"FV0H/Y2I$ \T6\B(S :QZA<.%$JP[TO;)K.
P+I+0@U\)8*%C%C>4Y$M_#>IB<@%Z^)V?UDK<:N\1ZHNEB_MX9;1NZ<=CW-^5^43E
P9/B8H(%C9;OFZ7FWE[+BWIM4+\. 9F')G0&6Y]!^\+3LGS)&6,V\QAH[AX0XQO!&
P7:T(Z_*-?./-TI]2\7>M+-F8 D"R0ADY8R^W)4KO*'C'HH/ PPN*_$0UCT=5 *CQ
P*KPMUK'O XBO+,,WW>CBH^P7R'O]3UZJ+X6?9VF@J>A!<I4XB$H)!_*>2K(Z3#K+
PO\&450#8BYM0*'#G!5O[I0H\;A.+ 5#"VU?GE$\5A;-=U>= BKCGIJ]P'"&3NS%U
PG86[O'&PF;Z^ =1XD57,-7IJ<#+3$2WP@PW.VXMZG%/XP"8+/22!;:9)+7*Z--V)
PW*K9N>"GGMJ4C3$2_1I=51N:M6XJT1/=6!%[LX_6N+-TNPC9K!0'9Y6Q:IJ73O8M
P](((J.\#XCO1TOJ:\T$VNG1_H!G_.Z8F?7=#DJ1,0, 4TM\)D99;E:)8N\<=><H7
P=Y:KERU;G"GL:'_Y"F*LAU+<C$G ->3>1OT*S3GMW3Z[?+H[<HD1"8*R_TCV_",X
P[8,>2?';)\'W[IK!;*P1%?]-%@ _DBTC)*I3AB.<S;VMMI3?TKX?TOBVI:M6O(]H
P %&,Q']6?VG:Z]:OKH@X,M'4'<;7 <@CUHB';(,HIE&$G/[ABF#YGZ,\D+KO)A[;
P-\BAV!C2;^@H]O]&"=O I6LX?L$,L(G1@)A=>*]P^!07K/>3:7S^$J&NF6MWX.F;
P#;(25R6?8RA8ZQWJ>S^VXGN==)YLNE?S/64-C$65N[I(]"#S;&B8X F'=[X7XO_7
PI*G;!,4?YX:(9D;P"66P_>LBN6CWXO%DNC.@.VE=E%GP5B(B.6AZFM$YG8B&]:74
PSHY?[ 4B=G_$9=%Q@ZW'\_K>2O\*B3L!.K39R.-I12$W:$17@5XH*BPL58F5IO+F
P[KD1(^#_$5*'Z\80ZZ>+Z6<*DN]L.O"G%'&"?0%\)%<O^ +)?3Z 8B>*$E!>TGZ'
P%:SQO U+SGA00[:+\F()V>"223.(Z\9C,R>=U]>-O[T<H8/>P56-_#*OT62F_UYS
P/?\@06(VGGH3T=8JH-EL+A K4!*:;!4,J=K7%'&:D#7<%?C+>'GXEENQH+?[GY)"
POMH]@;?T0R)>< KVB>)RS2OR[&^&AJJ%'\N+P"K7=70ZZ4(W_[P700'K)?197L&4
P#R3XF'V>&^.$MNY8*Z'[P^35^$5?MXHY5/;LL774-Q,/"(*W>OD]JGY2\/XN.,F:
P_"<KJP1/[W0L%(9&GNW&Z8LD %'(1IY^JD'![H-J$,QR5JMH,8QM_D$P;@W@6OUQ
P"[;$3P96$FDRN(2';O(X*U^/<?O!QTI6[6HE;4[SYRI<-RQ9I4"4>K5,9 ;-!;>=
PLQF*8"-JF*UY&WR 1 5KA2;+\B$,<4^\XZ]_3>$+X_N+9>XC;5R7!8"ZL?N0TXY8
PB_SKY-"SF3KT/;Q@IABL&(=.EW.>L6)1]YT;6GX)TLJ7^6>S;>6E,\W4Q0[.RKV;
P/Y\ GOTH3K;+BCHO7%3=M0 4LQ4A3]R;62[8BOB*#70?I*@WA 8%1,2T R4VE:/#
P'\P^<+MQO$J5Q)5M!.DW8HO\\VN;=VX>%_ HH G0IDP2D."8*2N+LY<5T_00($5B
PB?H3/4*I+A$Q=DT@(PQLLNA1ZS7@'R 2CW/H&"!GG4G?CAB4*4)6?T7W'@=YH8%.
P=\L$+(#\^XWVE_"ZDBHE/AZ <G'5:A#0%*]=6(=$ZZ2P34K)L/&"UWQ@FFT.4<T0
PVG'#'?K#_]@!*%=S5#2;-F(YB2+M=4GQ5JJ <[/G6Y9DU@<R*-Y@4QZ75TIY]+#K
P(6BE_&,>^\['KU]6FWA@?V<0N-X]<VFCC+TJ*H+%_\=T*7]._=,L:.*6!-176'2I
P])W3FBCY,-CP?W(2P*-%+7J;!*J>VO2Y\"_I0*_"&23G3D1!:2!$-R>TM,*CB2]9
PJ,ZK0==1Y.:EZ1-\PI=2$$+&OUWD@F(7.\$ #ROCS3N!)FKYY1IQ',K^^0%MN.#\
PRDT_/":4FHW;A="IMQ6>2*K2WAWL@[:T&8BB,Q)EZ9]KM S_[UGK2*57L*#>(JQB
P<XW[3:'OW++(K&:_J75#/\,B(I"[V?K_P<#G(\6 5 W%?#MV@4 MD1[G'R?#PGYI
P+ZYH$V'(PG>V8?QC]XK"\+N4"&B:")-M![H0H5/Y:]8E,M"4E#,< 2(I/DA>/1A1
P:?)N\4FQ.MM;T%Z%? "L3)>DKGX!9M7U+8=YV,;GCQD&HJBR1>8Z2SD3S^LR;ABR
P*<]<BD+_*L\\*,\&VCPP]4RO5'UDJP+XF-;G;M$E<0A8'YW'$4<J#V4#P47A"#S_
PXH7GF66%^I C%&"ML=47^%':'H\R_IY0D ?\#*)YT^DX&3P% 7DB+[:7GQM?MT31
P;8N"1$/T225-WTFL N8UI'5#Z&6S7W1(=N4(([K$@!2KLXI\E$ZD;=L #>S12K9=
P;?S) ]8X,*TI*:U*5+:*\OD%2_Y/CJE.6J!A3Q2R G[/\*CL&3,#P*ZNH+K+SG5!
PS]:>CD0&I4J1M9MQ3?VE=C03V$"BT&3.8#[/V^H<F-=<[V^LO%+P>10R]!I#; Z5
P H\Y%L^)%R"JY-BUEO68?_QMQ'\RE1,Q1Q@97R\XVCQ,$(\SH+&(SZT@A(.YZH6A
P/_Y:<9 X-K;X62Z>,R50+_C\<*&VJ&D;3A3*LA0AF2YS^D0,W=H'>&;/33D5TS>K
PB3I9,_92[WU%B?;T+'#T3%J;C]0<S=COT7";J9^$:SSW<) B5:5?DU&KZ05_-KD7
PZ;&?U0:3"I9&0W-CCW8P>[D"$1_ _">R>Y"YC%:WB7&0L( 0UO$I6[4Q@TIOKT^5
PC>J3#T?XR6#9J?Q_+?3;U1EB-55:]D^.*V4706EX?6CIS]'7D8\[:<ZP#4=]E1CZ
POX&^2XR#]MLLRCE]@)$1OYMQ^R(0R7?'1-:\NZ14[$DT+ZB=0&!P=WJ=F<>+NBL;
PT;DME,>DR2!$YTL>UJ(^H;RF&F!,Z3$(C$?IO_X/>:;RB@7S0(=@&>QQ@Y5^\^1*
P8'AI]FQOWWSC_)7O@2&K7WL^$J>,N3D/</A/.&%OG/,\JIY4E94:RWL86WG3.?P@
PFD#I=3TD+&,@+2LZE0>VPN7!*M-90KX<]TI2X3B_C]-6/56S!M/'9@I2K5WI.U*"
PX_)3!0W1,P4PQ3#41LXL/K&RNH]KR$Z[A4P[G'9, V$*+"%\"63HD;XX^,)Q%!(?
PXD'%<@+CP@$"V%ESWWZNA^ 52\O@I!=DX+KY!B:6M7ZCPIKQPDKF?P[=C/6+-8CE
PU;F^2J+R5:ZX]0CC>-4#2+WP$ZEG3];?&'AG*134=5-CUUV4@IVQFP,F4@#[=AUW
PP^897MM!S2^&(W,X?=7$?';>.!ZZ2JBPF6Q, X75Y!@NX"-]^,25 UOP>&VF$,5T
P><(^OS@<YA')-DK]2-'@<4QYJM-]+<)#^_T!2)912X_H+V3)@?V).DXT @2;\.WZ
P@+=&8X6CY-*JNU'\:-G6Y&*K7GJD_UW V_G@<(*=D^?S_*H-(LZ=28GC2H945$LC
PDQ!@#8\"S3?&PDF@1[BPK0:VCH2/A&KY=8J1,P/Y;:KWJ!\3'W$MNS*8],]=+!61
P3FR[_6$'$(%,)SP6W?42_#SVWAW&C&)W/_K$<+'K>PIAJ!1"*P;JZA<V"Y6-RO>3
P*-+?A%U;\B,GM7,L(L.BV22'VDB/GX&U,6%77;=L2-H\?F_A7 ,N.:]EB*W2#WI'
P(6_UX4??/3\YO9DS@_:CP6DO>,1EBK=I1513HB!V>':]D0$&5?<2<_-4^T1X(.[T
PHTG22X)Z<:B4+HEV;4^M:1X5H9BI1$R_Z8+18^]Z9Y@(LV5=:%.FE!&ECG,8I)2_
P_X?:YQ! 0[SK*C<0;TB=H,IW1XS@ .:UDD<+[:X!1&]./X'<U2:,;0X=!#3/,KF@
P \H3A/7@MF^*V$A!=,STL^(GKK6\!$N==<MP1"H3_R,K^R0==E?:9RZYJ"]X<XY&
P"0]E0GY]7LP3Y,X);U013;'/+E<>14FNFB_5&R(*F3Q4+#,+Q9,)24^H6$*"9Z$<
PQ"F\,E81>-;9H"81QMHF(.T4Y0YGH.UI:Q9 1 @3'+=9"Z90&CF8G9K9Z&2^]*#$
PE7ZLMI^W)($ORT/9$PIK]QHZU"S;,,O%'G5(.<129BJ;6_$Y<ZWGY2<]6\U[KE0J
P.;H/;:8KFK<]L]X1?FHZ_!E2_[LD$&;Y.O-Z:1?V+M ,%/$;<AI6NS0Z]44Y+5(L
P>;:N@I+G6,3=U:,O36O#POX/%#MX"(?54258-'FR^[+_U"?+Q 6_8QFL(I%9<9=P
P(&V]?@2@*2U.[!C/!S4ZMARTA/0;?ZH7\ D2%OJX2Q)[3X30.FX%CFCC?9/@Z&,8
P5=&5#1(&Q]SQB&\<C]X@S]Q#;]K3AZEZVG2Z N?S8XJLD^KECL#QWA.0AW7CRHL@
P..*,.!*GF\#7@SA_; 64'30 G.! A+A9>LJ?C\"=7W<VF#P92XTPOD?^.YH0$2AO
P"@PE);'%$D&?(P_:I6G=UGN;W)=QA:$Y5O!>Y,74M:''4R[UNY[79/5!F7"BWWE[
PAMY3453*IK0)?ACUNZ:IX!6KG.'?MJ8KF+D=B>H^LN:QBH%_&$3'!QM>(V8+87[B
P+/:@H"W0&C05[&R:_/N&5-/;DWW8;O@S/F:\U#'QG'3%::&X PS?UOU$R[%.V#38
PRU>KB%E;D:KD3!Y_0A,J] @XUV>Y*-?C?\CP@X-M\?\X8!9VU\\H:+Z,LD]8\ OP
PCY?DZS0T5UU;\J\P=&.YO\ZLJ.?AY3\;VC*/]3F[OZ&NJ83!Q>;]RJ6<L!O22MB,
P90I)?XA0?Z[L'_DNN;HOXN-ODZKFCK?IQN:!ER6KX1)ZCON?R7D;.?;/A$+-X,V<
PCGL'JT4M:]"7E==[-8)ZIO'4\O@ WDY._4]IZ=UO4=,9;2T+-*%>$U 47&)]@:/\
P$#I("&:?BNQ>C,?3:U>LL@B;F>)_2V4*&-^><_'S9[?+90*-_-539,F0:3""R"ED
P!5K+5 <@6EMEJ(CPI3#2OG_%X$D 5^<,F6\;9J:.=I^Y^P&4#*KEBB6A>91#BP9/
P&T5U%AUB]F@^U]>%Z\1)4)-M_S<%^L 2=G^W;Z,EO$G\-@;SQ2UM>O$M.D@A"TN'
PU5R^FA/OMZ?I)X>G@WQB0$($:CIR WL[D1ZH"-H)W'!8,H4_P+-L(BDN?.E(_<-Z
P-#.US(K!.R'L!O -'EV+_4*2@)E8G[.4L=#F'<'/DZZLDDB=T G"#A?CD2J+;>C5
P=:AH6ZM6$O[_6!=[@/B/N4-6(CBYZ#_!%-IUH7[M4\=U55ZNVVW9H?'4DR?)_!++
PF(,S5\J_9<?B[T*#-[Y4>3<<,C _?+14(C%\/Z*36TOO"Q>8[)+H#PNRGRT"8A5W
P333D0]ZA.GU3^[8%NQ,I2@GR_/S]X)L*1/O^[?!;J<CRYI]>4X";4F[4-.QPUZ__
PHM%Y/V;&RDC4TN GO?>^BQ3$OI=/UNQ]&T%+M(AJK$J1W7"%">P2T]@>$?P"VW4M
P&H(L*S\)NK!EN@'2HJY>VE/E+B$[P:?$N95.-5M,(3@I$N6688WW/,]CL .1]D$U
PE29R,4W?A/)89ZY,/3@^!YQ+M5^USX^GPO8*6]:L=HL;9A2LP@8A[EK"5&XD@O#>
P$,>53L^F12I;CY=EJ+H5:E.MB*O+":^[/-"9JX%3;]J2[R9XX'1BGW.N[)%#9@<5
PCZ(*S'IABK:O_;N:2*G'\)K"&NHD8JB/F)N9?WA,')EX6.4JT^<T7D;F_?V.183M
P>(;=OSVHR9KS&2[&HR19-(4D);PC_<OZ)\@(,]W*&FKCM738@?"WS?=&:QF^ IYT
P;_E,XXMZ#?45_"G80X>*>ZGGP'51*PL5-424B;2M22SG<]Y;U;C<O3&;,[@OG'(&
PN_.D'[.9^6:]Y*3B G@(*.OQTP.PK8X/0-?1,-#Q2QOM5-/5'MY:8GZ9X*=F=)):
PK@F22*.,[9\'5&K3J3S >[_5UW:P,MB,\P:U7/9O\[JK6V65<5K^9K5$DRR=2UTY
P>.<_BHO .QC9LX&RGVI,C-!%7P(,V^:$TNP[_^0*P ,H *H4 +X,9^T:MSAB.&!9
PU&52N@152\/_9)_U^_);@::0EER?U!<+4A/#&<[?!+#)N%T@PAQ^T-AIX,4U5Z$3
PV##N'.'X^;6W9!2X4&& X,3MVP50^Q7/-9)ZM7$&0A9?/\0/(E,(':P)1"LOT[LD
P,8;0T@3=L:+;.="C'AZ:JOC1RXH-EAU 8]*MZ\TH]<MQ5IN\I!E)Y#,DLSK(,OJR
PU(0CNGTB12O7-D)1S6GO4'!JQ%U>YOR3X1K*P_EZAD"[][1WW4 70?_GV#>,-7K3
P)HXI[96O H9SQ F:T3#]6>FE,!MH/792G:C"" ;]N_QP?_)+R,Z!&_ T5#6^\Q4M
P^U"61\G60Q195WY33AH']AUQ(&(1DL05K]4@E6(+,E[R34Z;0-T?TVBZ:=/_KS7,
PD"6T/BU9LT!7T"1KU16 $PX6=#J;0:S=*?;>];A);9BG,#GORG.>,'8\^+!R61ON
P"=_/PI/^B;A?;7-N^*%4KBN&L/WQ%3,K  C_"&047Z5=H-A52(1DD[W1 M1JC%D$
PN!MN(#O22W21U0.I!L+Y-G'FF9J56G8XS<:Y_ SCBD$B#2\&^VHO089;C;JT#FPY
PX:-V<%$=[YGG;:L8!+#F"S<*W(.C\R+4DY#4;M6D;0L@P& M#K@7LJ9]9%^-6N*S
P@QSA3: L,N26V[_M"T_%$6[D#SK?]"]4P[D^9I&PCU48!@$ $&/GYT[-/Q??YLPV
PA+A M%.;:GUY(!BBC$DE9<Y(F*_UXZ$$<CKB^###FL0BBSI[A4-,5"CA%6/9I_@"
PTXTG]V7&<1DG"1"LG#X2B3R)IU'IFB;R18Q#VI@;?"FX71I&Z+W,)=L^OF]Z0P^;
PUJ2*J7.@TN7BU)\8)N3#.<3A.2&)]YSXT9@<CA2!S-<"&-PG=R'HGI@9,F<PZB!3
PT7_@=$\C<<%>939NWU Z*ZUUQ"*-CL3*:O6YCR4L%WO5LP538J)>EGZZZCXI+E+Z
P6\"3@8_XG_ML_+CE8CS>S77!KR&W8$3W6"P_&*O:TF6=(C ;COC%?290X#M4D/:G
P9G*$C"2ULQZEA-2@BKMYY;CHG]/L'_>%ZHYZ$B2N#$A79VC!_%4N3*QP]W'[_67U
PC\:.)'GRB<=*AVMDK9O2==,>]2> G7"YZ DR\U5JDXHS@4@MXN8S1U=@ 3EY[B\B
P$G#D3<YU?]_[#>,;A>7;/4HU1#WN)=?9,8!63>SN+%E?"_^X/)Y-$(H8)!$C->X,
P0*OVW#>*7DGYQ:)O/JC-RZRT5SM[B&T; E+.V'_RS]S[5-+3LNTK87A[Q2^/+GOE
PJ&Z:[ &,KT'[/N!-E01O,F5CMF'.IU4G(3E"E9'AN<O2:KH/;J.W%T<\249J>.5B
PC,@J.,?2($O&(.<$[H_?R24;"^WMJJN\#V?KC0"NVAT@CCUE:/U%?E#DU1/^?I-7
PHU*7B(1Z'X;-I#.V@\MI#3DJB'+_M67C>N](FC%[9NL*E68#8.=*YQXV[8SG_)\^
P2CE]@+)T_$4Z:,MSP^Y\<IL=YP$$@)3Y@.QIS(4+<S6J34'7D.B+DJM2L]0KI>RK
P%A/O\:" BFJ Z0%FG*W%VGS'6;2LU_>$0HCQ793MZ3R&BI-K9(($$;98$\EGE/-[
PXX3*6KBOH2(\L.G%Y/Y+4!82]"&[4IY0AD5I04GZCUT/9M^UJ5@4^HU_'2=:!4\_
P?<MWA=@*=@RU)R<[XSIO!/A__2+GE) G\ I8<*R1'L+.?0=KW1\)0R &TG_Y#!'$
PY<Z6GNX+_XU'1P6\TP"4@\HDH?>P]UHU.%9/D_-D4M@>S\!K=9&,7682M 3I+D0<
PW%=MNI^+8$BE..1DW,?^B[AT#/ 1=[JP?. #M=0ZCK,57=7"[-D/J4P,#1KK^$?0
P/G$1OX,</+PBT5Y.:?I/)]5M5@.</_DT>QPM5J: IO(^'T6XUG%@OX8-!@3Z;E3=
PN)QNZWQFYH+FI'@D[>KM2#GR:3]V0^"#58=4%4K?WL/Z0\M1;6P#?11_F&PG(5[G
P$:W-C8K-W%>$R1:B&JXFP%XXH*6&2!7L)=P":L\5B_H9S'L@20$9G&G8Z]+]D:N#
PY'I5KP2(+)L@ZYT\H0*W7K8G@O.ZPL),S<-IR(_O"W%/,0V*%:HN=2K;:; G0"?D
P.'U&JBA>]2#/,>YL#EKLE.&#ULDR!E2]DWKM+W_>M/@M+^^",X/#AVAG"T53)[P6
P<$6$=<'#1?I+KD]*[B!">YM4(XR/O?2D_*\ @.MBZ<C>G*>W2_):R*]3?*$\9:I)
P+!B/BHKJ=AI.-(^3-EW.BA#2]!4!6][UI=RX( J<L,!@NX5%?T\<_<O7K0!/=M3N
PL/;&G&$G#G]1?+P2FVG*GZ//W6.I(BVF-2Y\L[.(U'_ &^9BWV\%'T.@]V/ &(SA
PW!.['-"XVC:_<I&7+7,6I5'Q=3Y??09#@ 6CZ:Z(=WF<3TSB*S"OHEIXH5GV;T)T
P;EL129)P:U[YYF)39E=J=W"W7C"V?45C%^5JK;@_Q1L9,05F*U1'@-*]J-MUL&*7
P#RQ ^8M.J%7OQB*^.+1 %GEAF;?45X"<0.> 15Q/AD3@!JB'(ZD<$O,]?X0;3@SC
P+D%!E*(0/P<P+R4\V@T5X^FXA!*:P@PNNBWB>-C-&U%."^9F 0$]*:">A5"VSUR2
P.H5<Q]<Q:F'!W.(-_2F8UF/BEO;8-@ B>-FL#D K-I_DBR1Y;#;;(L045\8?(#!W
P!V&_"\R:$0:<:-!%&ST4=2C3/_,;WX(-%Y0DO:OQ:K_2LC>8#>;6K\<E[B>QR/R@
PY^,,4M;?YH7H?[K>NFV5_'Y4.Q$L30VM$DNI8/6_6&3=D&/FQ'SZ?'#[O)ZL%[>'
PFGVH!M<9IOU\\C^SE^&#.=-Z\Y@\B%UAAI:)#F[4:B!>V4:U;#X[AFIS@R>#X@$;
P)H5@7"\#%G4.'JWY.&;!/HY*O-?1LJ2WAX#O>?:?>>)>MFG*\$5I(W%LU_NLRXB4
P1[<+AE2X>@/4)/5^'9$NLZ$77H/-Z#S_R(/-%V34\NA)9V@+L"?=^US<\A$O2A"?
PP6@_>]\>NC,&I@M]2?Q4'EUF(XWM?UJ%>60:D%W_[A'*6]$5#6V8MV]Q*_WF!AMJ
PHB 2C.@9F7+Y4CF10=-]O/8DXY(T-(H"CXQQC6/E;P\CNI(=7_K\A>->0Q5OBR)3
P5A4WUVDB)'\G-Q&BGB8JT<_Z9"E^Z7!BQJOI=DNI_:MWJ<#Q(+BJ2X3BD@;N3)K5
PVJO%&ZCLZ")$\9N9*N($674CRPY'2^\38MUK^QX>CUU6,QR@-6DDR6H;<UE&;\X2
P'"!/+A!T#'>0O)T %2T+O1"A<W9C?!, %G>,EMWH'02^>*32LL5),,V#Z_S$E)!T
P!>X2E8SM 9E\ 72VJUM/[&"UW:H6^EIR&<"N3@N\][A9WE+2ZD3W*])7@5LR>1_$
P+XF&)],Q=<P9BM9MDRG^CX%LO*N7.T27C03@S6^7^"._-ROY?B@:(58!9XI]O",=
P/'D6Z57A']"^X]X,@!SB+A#OX%:;$V3A5Q/SBW,>RB06](MD!1T_*DEG&._O)1W0
PI@4.H]#PF-D^D;26C+/D!@@7LQ \+\E(Z)KQB5H_(0/82:SD.YZ9H_DV'@^)9\4!
PFZ:G$Y4=Y!NFE6-I"W93[LX\RRQZ&T<G"1HJ2:TD:BGKN/4_4CJ'<_^_V5FMH)\P
P:;O]-!>K@9[VHLI\M43"W^Q3@&!60*%K#QWE=K,AF'5C$GL[A26:<BNT)D="AB7'
PU?II26.*.BF25&4"INCG.SDDA'WBOH'.8,(N:XY*Z.0E3R0M3[_..U&_>'A -R^G
P+EK9,=#4HC^.7K8,52GR6?9N6D=!N"8B,/ 9",7]]Y?/D?]*$$X0DF3GIHBB6"-'
PRV>3J<GCWBEC:JX"AK4KM#] !GJF:3._1VITEU*$SY>=(19DW'3)J4!P$3;UB\N(
P%]XIFKZCT]Q1R;\N0M[R.GC[20G\7\/I2'%$?8K'R>5%CJ%W/[R8\0%R\3=;GC[M
P;!6,#[33:%QF6C#8?@WA7)9F*R-*<8!HX8/Y-\O'4BS>^WK4K>8^%4"(L@IL%<54
P?@Q)PX>6]B,PK7+&="]#DB-[^ +5CXXP1>->U&U_JVTWYR?#GJRJ!L3:? &9Y,:S
P?:JFFWI.Y6\5FV8CK13ZX]'$73\IU,Y6GBRW0-[:) 7P64,FZI!@YH- T ;V@'L!
PF&=?#:H6TC/N<%EH5 ZP\QG3%T!DMVJ<'R@+R)]GD6/<]V(1J3+?L'&U8%@S2[9>
P-Y 4OF=B?E/$EW- XZ$S,2*[_?%,6"2N5--:R2-F+4\T%D1CZH9QV#<"S_^3,2W=
PPHYOK<)XY]D 1CLZ-L!-;*40];3-!P4.(0*J6N63[4[:$%5O=UP"NOB''_V'7D85
P^A3:4Q?2+?=F<]$IULL:'Q7/2&_'0*<N-W/O/Y[NBE@[24&[A#X#A@_V*X,5.(,A
P07GU\.7H9]NO Z^O^LXY>_C'JG474[9Z<'A+$7?%QUP0C39/=OK"KA=<1UZE-,P8
PPJGF*=>!R KN8K$1'@"Z'O'OIG#7M->)K.GCQ4\_4)>1_-?4 #&$-J21N+^$6V[ 
P5W+%:#G3^C'\ZQ^LD_.W]$USGL>*LRB3IJ/UWYY31;(V1L3 K3&%3Y.Y;3"CU?SP
PN[_N'JP(50=TD!-N6)T (BLT@:YYM7/K.<9@=I<N03!?6H3.QDK_I)WFF;<U#,4P
P7=0]6933).P+PR"V<GHQ3>HPQD[K^_K0=ROQ915"Z&'Z"JCH15KWO,SP_78CE'!*
P-I/8^\24?.3JO?$1EJ3:21GIF.IS#2)K+1$J2&[)"#V=&#A[:6MJ2W@6',-\^!V"
PP/3FTAT<WF[=<NQZE#PFR'&KXQB4.J+G[!YV-\I+PKM<SQA9 EIH3<93.*@QFXC*
PKHT2X($_$!0*5(+<]#K,4:\F18JR\[@WJ[]DQS*J ?Q=@6JT,8F#;6MW^AY)<=B"
PHZIS<%?/PU43P[7>3$"%,-<@A@> R+]"'UJ.YY,KJ$(W>\[JK71I%6C7%ZOM5/GA
PC'#CGS<'T:2=],W,.+]-L#/.(K;S )V_0G0>QTK>168I?ZB37>8I]1$&D"<#Z<G1
P:979_J:+>3593E9T4#?I!DJQGX\G<W?65AM;3QG\\4@JEY(WK?FJ0:A6#/]VJ7H@
P>Y>Q=S-X2LGI@[W@#!E'=](:D7)&VN0)AJ(BH=?,^#T;5(6,@\!SK5P_Z$SQ+ES0
P>Y-#,$UG[!ZNE.D[CDM-F8$+B+'J/1OABJ9M$K5\X[>P*Z:DGA'@.R4.%#\:A![Q
PCC7(@4=IL]QE4TGJW\S?XVV4:G)H<NP^H)]'UWG/0I'TDBJ4P85<CJ.#5SH,]P+J
P.1#'"AAU<9?739/1&)0?FBR(,+DN_N3CGD<*RH7KAP4W_9HWJ@]QD+$*'2+U@^H9
PY/VDP_Q8A7#UR?HOO)=CBD&HVGON=&V4H8+$/ HY,N[B27?MRE7VEEW-DJO)*2K4
P&P0]%.K@:9-__+;+U<&Z4"V93-4:H)F#Q!$S(W\N"QLZ#+3*E#4Y:UG4>6(>5H\+
P'=5AP]IO5\N2!JMV;8YD;)[;.]ET&D3 G(?C-MUT!N=E7RC'?Y5&DW[IY32W^9VU
P02 SV40G/%\Y$9U1?FT N6(_MWF73I3KP?Y"1OUH6T-.88*=%SO08VL;&M;H:H0D
P G:WY7<$T:N%D2\[%(-@KS?B+>3,_&%I7"91V1/55=MXM=,KBM\#Y(M#LVT"X*A 
P9T:^%HV.A=]H%X;EN\3%24"+9K_,YL(E<^G:]3Y=VJJM2<#WN'U2+?Y'(!U2C!3Y
PFWC%STP!R(YFW><!R1]*P+2B",(LQJPME6VW]VM8:AN#,PB.=C]#YC/G41Y6MM$^
PG6,PZ<.ECDUH *NMZS4WWP/.Z267I ST5R'_-R1IHABUWB3H-O,(^I]JN1Y(J5LO
P@JSS:13_.[BRA*"F60D74@@'T\570R)A 7$,<HN<. MK%TZT*L^\<V$7<BPB('F&
PH@.=*2)^C-4L7-;Q)S56IP*'.Y@-+B60U\(@/0^E5F<FZ\O&'63ZUW"?^U^]-'GD
P_[)*1NVO.H_-R&**JY5J&D[]9]#[20:<U>BM*XQ>:*NYD$;P2-*FC&6S603@K5$T
PDQK4=4+SF!H(@&E'9JW&]F 6"V6W1I5A[Q#K)R@(RIY&5<.."/Y5K8Y/!,K0L2V=
P-.:5MV5YA/32OO%_>B#B2;<&"&UQMC_#TE15=T]CD'3=BLRVK28\S"T)Y&MJ8$)-
PQ(5EW1N+ '5_)*N/AMLI(%])WRL@6QC@C,.O,<'QMG!1TNBKWF.&Q1ZS^R4ETW+:
P@:]Z<"E</0EU>@>; :S$"VX.PR;UXW0<2H:L"@5>,8O_=%,$$3@/X/"4(,&P#M!S
PE:^=,TS:9VN4^QN="U#0W 0SJ]NSR"TQO+,.CSNS?V\2(7T[6*$;3#=U ;1$Z\F!
P6D=*4&0:UY-06OA9PJVJG=JMO>R -'ZRS0*43C#VJDCTIE>G*X6(PV^+KDXN3VHC
PQ(@^;31I0&$-T294PG,PD-_/R)M(7E]>]4+<MV'R16,=O9U:<2S/!\6P>V]';G@>
P6WA&7E.O1:T-1; ROBN+J;T)GXW6J,;4=>N8-BM[!PCRPBN,"J,[WQ\3L)&46]*&
P\H3E18;9IBOM4"XZ#V1(>C3MG5M[N&U*' .#)HLE1PU+&N+DEB-%_'*/=>6T]R*S
P] ]I%>@%6#7=.>E(:O_3MDL2+EFN>H,V3ZS_$KU"S<?-<OC,G?%]I,G-G'T-W;X:
P37WD4+N7](Z?GXG8UC*QM.Q!BMFZ08\AS.UMTR)]@=.8']0U*E<C-5.@?*6,( WJ
P>LSB(.WT!R$LHWT=.!S#=,$7GUYZ7$6+H:P*S"8DJ4_EE^=@>)[+>_P1O=80R\B-
PW/M)1V0:69 0OIKP5]R#3.#6)[1&*-TV_AJEK%'G,I'?)C&[_FDF-6.0?X)45JJ-
P0^VQ&OIYHB)A(PH4T"XE>H2!@$>!9Y"[IH+3B;D6D4I.[]&NBP!(6\.TG?]I=AI/
P9R.[<5HMFVE(0D=K5S7P^'9%+2#[Q7+6W& -=1]Z.O8FGR,(&&6$L=:3C$NN@NC;
PZRZ^*=1WM/G+95TAOUS0([;%ANSLC[D&5@R#=#]<9^^^WKV^=N$Y(^Q>2:WJ=@ G
P@YET6)2D9&_Y#],[FRX8)53%;5W9&V7=ZH;NFV-//K #/>$UDQ1^>NW6@>*0=8](
PMO?4+$U.A@X+OWG<2J2,Z1;E:8V0IF&/%U-<.Y\T7G*_4'L=%: V^_7]HABF3:_#
P>))IAO&$7BT_D40+SK1EV@#.VXWV709PSOV_O"U82FL][;Y4EB\Q[=+N;B-AM1"Q
P NB1>?8$=@8NQG+=MUECBA'5-VYZ_$KL@44HR;7F.%(V>6&7%=[;1HEEX=\J/+-U
P7OZ+)*8( 625TK5!&4F>*:F[]!0YPFOMH=GBC4UJ@']$)KI/I-4,M8)&GO//=D90
P2-<+&&=I&Y/A)D"@P>H9 [,N])[MVV8!PM#'XE *)O#]R0[4;R"1G>RZ\R:;WYM3
P3)S[X(<.D;M6E5S'^E$L_BCA2-\I13R_J@.8+^@Q7&^&T&DLAQ)98D0Y<$,BD!M_
P!4-5RG3+)IT;B*L7TR7,9U$_\00O#;N5/EHF13OF:L1MX;K2=^B86D+FG-_<6F3\
P@RQO_2ZU!F$Q<(BY=KQ-Z(!4,&+[,JE]22'#=X#LBEX!ERD*;"^!"5KWU=B[I3,J
PM."+ O!B3*:_U4L)^T+$TUCO8"W?:IJM(NTR?#/D[WT+(*H"&9=:T?$&"P]1'!V3
PDE";V'%'5" G^@T$DF!'6LW78QB-/U#-(YEXZE2J6$57FG(M=(2AD(V\$M=3S7B$
PT@>,$(RL>(E'S1"*==K2R-=[@</41T#3[;PJX7#TJA@ K(L6%D8]C0IPC$4P(S89
P)$H^#""\V,!KB+RY:T*A$J*2FAMPT%I?BIZ%9PBL#(S\",1XQ %B3@ D0YQ"WN<N
PB@K/(D4/?57-H]2Z"6UJ,*87.GZ">Z^7'!=G713EL].^^-^KLZX0ZGBCILCL*= (
PXJ$_EE$!89$0ZPCKQ\5BQP@7?JS#2>G"I(Y%#A>/OFAEGK PSIK94SV,9QR+')XD
P1@VB0$1NH@/4_P$ZQ7D.U3!;,("O&FFXSQCP-IM- 'B\B$OL*(UHDEOYIFNUW.. 
PQ'D#GXM)JJ2/"G82<Y\3 )=7)6GU*;_0;QQ0QN@11XW.M,Z"#<:WQ,0DN_[YH[2I
PA>:,1S=-Z$J$9CX<H64ID@RB!2)>M,%4^VHAKM-]U;D)W25@B)_2E!>2/G#TY"5"
PAT5FG]L#3X:$E/)]M[%WAQ_R*G'!EB!C]6BLS<5C4U?/''$,!8-H2D+:V-*=>-!2
P%F47 (R+07QZS'VHU*C&!BQ@K-'$!;M5:/6? /]@J^#9VI6;3+*3MVBLF8KF1(6[
P/(YH6Y=QOS1*F+_%>?M[4*GYGM:Z"V?4EQ TK<'&S]6=#NIXF3J.@1Z6%0/I!*5)
PC>K^^NL;027V(Q>OW? SBNQT@-/8[4_,K6(,$_&VH]VXHPT-89Q[VMBQPCM+?@E)
P$L6VETA&"N2OX:I9!+=.4'3>-!V"R H05_<&Z',R-U<Z$81)J&GZ/1!JL;K^:]MQ
PE1M)I9^\P<0TROA9->,-9;M2#>=R</)I(#>@?@@->5I)QD0#Y)[NV%/4J" UGOKG
P6:WV9HFVS0@8R^#:O(6\U)'$)4"FJO1KI>UKX5GM2^3] E1L@04:.'#/6@7W0?5W
PZ)ICJI/[!/"ELAI$% +5HQG!2=J+1Q)_CU\_K67<HR8EFXT%'@%E0E:I@#])]-!7
P&L%]["RHM<OW"0@H(E1ZWW)!B6P,,RQ.E$=&HMKL[T0#:H+<6&^EG(H4HCYMB(1/
P(;]C?2F&>&K.':?WO0] H__2,#1Q_='"QTX" Q,ZL!G0/ ">^3U1%'K8<5KILF("
P3&BF6=D]<"YN:HJTN!=O*:MRU*#8./+K3'5?)J@F3,^201;>D)B2\Q3>JDB+:_Q6
P(?G2-!OP#*:QW]K=2X#?7WT\J> IC;B'HT9?7,1IS&/?/LR!1ZEPOJ;7LA6?1T*N
P70!5\]NOU&R+\=/E[%@?>#*OKW U<XM:DZESV%;V9U&101*9("+/1#5,RI1YH]5]
P_VTO-8]D@)L]4_>MD@ 4JNC0_*%&P,6>CAV1%ZXV@[2C[42A#-&V(EKO:M?#RU!@
P\-/MNBE&2.KLB^9F#3^D_!92!8/;#Q^4EG%ZN09!9[PS-6H..GV D+?[7]>3J#5F
PS/LQ0,0B!H:<2? +%(UU,&@G&6\FP3;J)C$V[1W/44D=*\(V<8NSL:64O"U?D0=(
P?122+.CK^A73N]U@1MB=Z/QH/5O0G.V(K"9^H00D0(+C@\>.P0!B^XA9J8 *^D(B
P;<D*-<\ZS!]Z3JO31&4N$//AWKE$ZA&*_3-NOK%9:FIUWFQV4I&A%D#W=_!,)QX]
P#<@Q?6_&%8M&>9S/+_\OHLY;G]<HHK_$4#E5TP8C(+CB0TMC=16!,IT53^/A^+&O
PG' ]W%I$JF=I<"S7G>%P5Q?5JH%SCO3O[8B)';R,L F#QW^]ZUVT@OU= Y3U5W&\
P,D@\( ^_\Z6 W_8@0GVO?F+3L;.,[!TH5+W9U:RM5-'5G-))F-]PJPSH72(<=?:D
PJ)Y@9;1O?3O%SZJCG89AV&'VX=E^'$A^+:TII<_>6N?M$WB;?CX91%DIEY@7/$'Q
PI/?B^@U41390!#&MCRNJ902$"GD>0S)XBLD&,A,K[/:C4G[>*,8]A@LE#,Y_[=]@
P^9T!L\#8)_[&/7.QQL>I!_<-J2\JI:D(J#DY\NPSSW/#$N H10FI#\[4D$]8;3L!
P(R/JWQ.!Q4&IWQUGT(&-G,S,4.'S+$ "E[D^M6)%9LIOL ,3IGLZR/5:!](W%-HW
P9PR&WYL8PG*?YW^,;@.GS L>Y6/[=1W[^3:5_O2?"Z/7SRTA+3TFU4-U!@%/NF#E
PWD=9DEG(*=#NB^< 9U+:H?,+WS,LV<UR:B1X4L>6[XRFQLI@@F#Y^_D&."M8HE0_
P'%--7YA D;>:V"SG8L18W NE)R_2/TEJIF:]% TW$_1 7-]#(%;U+K^:,[7"@6PM
P>O"$[^OKFNV((^7HSB"!KKD0U24Y'X@%63!3VRDOVC3.UOPMU\#T#BO_-\!X[7I@
P5UFWUS0RK2.P,0/8*W#\A_GV(9F<'MYQ T$Y@EOHQ$BWPQ/PF8H0(*[;U,,95?DR
P?@UA0H-+$+<)#2VH&4!4,1-?)/I:";1=\X?GGSNM"GNJ(,56(?23@13()ZEN&&%T
PW5RV$#=V$]3G<35#W%*@$KYW[>N]HGL=[)##I39- 47.:3>92P/)IIU0=U2I))&7
PL!1X]G\6%=#0*K :5X4 D FP;.96(%+/V9P( NY\##XDH2Y=+AX$&[H=*N?@EPJ'
PN\B_]VX]X>?(C7@Y.3(B?[6W=T;B>^5] PEWU.6W\A\R9$T@)N+[.,Q17I"AO#D@
PC\V#_+6%?EX<1TR]!7'.19N-/_[E'V5A-[J:HXL5S\0ZBJO /FF,A9?WK'2[G<+3
PS2N@F^A2=*[V*E)Q0"U<8=)'/FZ-\?WL,)N\!B>KT/C..YUS1"4S>/M]W+$OS9GR
PI"0^T(_8>K;!N@MC#BL@T$8YA4=Q 8'0I'03@!*D9N\6C$CHV5T=XC<D*14>QJPF
P%WU;)S'03#]H=2 \DN#C6)LF+;:JRM329!ZB8_+PF,=UVL<;@4W^V?^DLQ_?OZ-;
PY6EV/'$:9(2>/DIHU2(%V2>IS@[H9-.K-@B E,2H7OX/ .&QX4"^W''=,N_^P"S5
PEM!=36;Z*ZNS5#9+USV[KR(P[Q2D%Y%X0:7O#C43^LG'V)O"<)'WG88:KZAB45N5
P@8'"UEEUOYTZ3:<3<)E2@44+<]82F?"/R'ED7Y6%I>\(NXH'\5BR-/[9R>EV8GC,
PGHC=7?[6,WAWJ- 4)5U 2JS,Z)"S6HRO ,]2()HD  _FZ)F7&7'9%)GAF(-B#E;O
PR7;D<2L*Y,XF;\G95K,U9QCA+69W'NGXF1%MQ,5/^'TX'^]"H7A-Z-GE&(>WDA5D
PVT/1@Q0);851\)9 @+SLPC'WIVS)["(X! ?A-7FA@FFU@LRK#F!G<[K#\.KT8>O)
P=NC(:>I?$9)/20I:T0U \AECLR&:4UECR]WO56I@)@NG2Y')B)9V+#P=&4PRAM[&
P0P_DKQ%)C4/*^-2"'_)G1PZ#_EA_VI]ZOG'$".E&_C)6+7R72<P1TGK71\8O(VZ$
P(8_MW\DY@%F/*/[5;N9*9Q%:XM77[V3&9FV!J*2I?(;_K- > @[JC_@D"1",1K/I
P&>N]2Y+V]V^Q%<A?MK/5P&PG3*3VET\\>S%: ,P_Q0?:G5[8!@#--^R9:Q939\6^
PUVPK)/4S;Q4 (I*\LPA/;^%19<U9B[?7T9C^X8+R9R.7Z4$G,]7@1PS^V;V3W!6/
PFXWHU946M=@OJ!MP+;V;L_'MMY+KPS&EH1\RCT.$R11VGHM;?/1M;72Z?-^:R0E%
P=@"?SS%IY7FH]3>>M=EV*!F3N%F%LWJ,"7!;BBVAO1MX/&?KKF@H\-0^G+-9<EA2
PG7))'W8U<1]7)$A^6@])I&/ A%9H:CIZATV&(LN6T+^)I,L\CIV$1@V?$.9=FR9<
P(*'[FTA/)L\6'LG?!\VE>VW\3W7'1>ERP1U!]GL1]*X+$>P3+!U*T,,1-E,S'OZZ
P588SYM6Y]?&#D[GX13((=YD 97WS/K3OFJN< 0CCCG8HF$P-5>7_:$*CT(31!X!Z
P=*CI%"YQY&UH^-U)<>U^O+ >_2)==V.F.H'Z^D,S_CS[30E8T(\VE4J*&6'J!^_/
PU.\SY^8??8_1+Z$&]:D]@YE3P,I,R\62< U"CJ1O#:$6<=Q-$B>KT@?+OO5A^,\5
P<OG=-))?R\-RF4E6FXD8_Y>:0_45#%7YC%:S3R --#PQK\C4^(?MH[19F!"ZTY^M
P53>0Y! ?R!ZD3=VU#;2ROIK+H;R.;6_$L=7:3N!=XH)5Y:7RN@I?6-(]#.#\*!EJ
P-'_S7%G[4RWV8HC$HY_KAR 9LNOO:D(Y?\&KK)V==-O E_.>33K.3:981P7R[V4M
PZ=@WZ\L9-&L%041-U"TV?\M'R,#G,,O'>APA6Y*[,*?1%B21W7\&$)DB,UOI#Q4^
P<! /U0QMUN^N T12 MR2DC9S<"JAU#EF1S4E]N>XW9=40P]R<GC%U=&[=>QT%8'W
P6"SG4S#^':!V1DL4FZC(N'Z$JIG24/$\E.6M](LY J@65(G&H-@S3E/N!L\!_YHV
P=KN0-XMNY=),6[;Y$!X+T"ULG1)BY2-GIK_Q[W):632L+BO[U*4NE$C?0)"166D:
PV:MWV(X6NCJ+D!5*/<!<C-\:ZS?4$ML/L;I>(R 0,?L&/13,@FSC_2Z)_0PB2J9)
PL[=/\8QE0Y% _,T4L;02 59C3];E(&8]7:'Q[H\_)ZFW#]*@ELJ=GL$N>*;K0W["
PN(">Y:\.Y\S9X1T,AL, &*0*=6I\$K3X-76"*S4H_\W*+/INDM%(9[2V2?*IETO+
P).YAL#Y0]W;J FLY?=]8B6ZX;D+M-YW(+S2D?#9W',OS!2*2U@ :2>2FOI^$ROW6
P5M\P?&WG$2V_BZ38RNP;4\ZY$.?#/"MGZ(U]DC-=3S1M+KN\^6G1,>6(;QW#PCBI
P\GLWY__S]!;:3LJV&J^K2.J<%;YS_/XD*;(\^PTGWTA#!2PE 3!0%0,/)QEKHUW[
POR20N']<,_T)?8'T;K-?*-'?ZYC/'VA=1C*)O'6%T GQU9RR<UA?D_ZS@R<),QI+
P/F)H;CM/6<0$(R9;6NU4+-BXU-$7Y9V/&'4?J-P&;5Y^H:V<V73F?$X**5;1MVB7
PLQ1LV?]P%#;VW*F*<A 2)XB9=8N9!>=I@+SV#OJ<[CWMAJ=8\?>E\72[-H9?ZVQD
PPYX<0X"_46V]42H+-JG2>E<6]:PH'4B>9_)EF9:!^(JVA2.S0?V^=,'PT'I!3K]N
P(K9^!)HS0"EFI0O/]/:791O9K")]DS_7/)DMHS0<S&-%5&B;I6#GM_0FM4\?LX[3
P04"3FEQ^N/^0;)$Q<#Q65&L\J557"N]5_QTO4$( 0+Y>-J*L\^^ FQV4OW]7KB[E
P@[T)82R56Y)TKP4K1_I8/G.-%WU!T2ZV,:XVNPRZF;(/^4KLHFB?>#1!N4J(U=&U
PRH0MDKZV;: ZT4^>_QRR9G7C 72$W4Z_&\:KIX1&1ZV]FL^B+$R1N6CVTS8VO:U&
P3WG2K_MOI[I80=9.%.EH, ;TEO<!?D+7"!Z@UF%9:22-LF2L@!(*V,[4RW[Y,=;]
P7&J\ !F3D*P PN!LGB']H9,.OV5*;[46^@3;.I#P)0ED,@NW36?=),D+?N+P6#Y1
P:0W6=0:UFZ8)2HZ)-D@:_)].W]N_,\5]>EN^0=D]3Q@7FL49!7A"9E^=F8\83<XZ
P!C3FT0UB."HO+;YW?'!HFB-Q?04ZU*!Z^D!_]HE7!"[[VT;&[7+'5O2^@U^>JN0'
P'SOL32%)/9/S=)(*ZC;AS'U/"/+^!#++I6/LL3WGT= 7X#R.>/$):I[+8"3BUL_\
P];@00+BVG!^@'Z?)QWXQ$]Q'_JGOKPIQE+J@> 5Q$CMWEZ4)K8Y]*F><\&7CDOQV
PLV#M8$^#0L%M*VCG\)Q<,R7KX54V/S+(Y';^\Q81CS9*PA,&\G]^[WH>P[(;IH@X
P$TDN6_:XA5ME.S]V"I$VU_:03O/?9@-G0<9[1N? <Q*NQZL+N66KD?3FS[$V);D[
P(=E1$9'_< AGGW>#G&)'#*1><TUU\#M7 K;$(.>U=HE10$]C7;UU3-@W:F+#NM6X
P/ 3(SN$2JW)H"8<RE*V"$BG<=$3E9!G$8=C=XW:8/[D"B3:2ZHYY&MCSND6IN>?&
P,VR$MZ@S2+,&8=J?7Q==#.7LS/@T]/*F;Q0([)>KA\RV$;(/%^OG7*_S":_H!_VX
PN2"%QY#_;^#D6=8F3#OBC$8A&D70+5UYDF/!:-W_'>#,T[C<[!"."P\?(18==X89
PO<%Y++,\-X]R4I7_>/?&4 C%<3)GIO\]=1G?$77F"2&!71R[S?82NXE7)BNH]C,]
PNGO5/6 IH?K8//[6;6-(-Y\<2-URZ<'EPZ&//&=B#$&/&,7S;,DXGQY78.YJV*&_
P01:![/4&_\_5JJ[U5P$?>N/$$F);%^^.ZO= FG M*+@#'F% "C &DZ#';+Z*T;I:
P^B,2H-HH,(#_9;+*O6'&.S:3Y<(<4:@LL.>2-&'^R0<IM^;JT1MJ["(I_$JV%[Z*
P&LD[)\74W?4(\_@S%:AF<0&XVWD_7@2+BNR6;>32+#'5Q,M%W.TSIY2I=;FW"FT=
P^A0X/Q0N3CX@C8Y)1!&&O9X6@N?VJ09DY>A(F4>JNLD"BY)H<0 DJT3\@&)[^U71
PQ#](M7'@,_R IA(Z)M0 5UPQ1:3R;Z>$QS_RN)ZFU(G(9+5DSB%DA^Z?<(O V1U2
PV6QQ*,.X,V2K!ZCRG2TDL[2JC\21K[W.:D26[$HWT3T>Y%@W00 O#*CEZ#9R;;3C
P:L&93(-"Z=TJ!E08>63U:->ARH)<_=;+ [RB/K)""/.G@UVWUYRKQ2<D!-FPXCRM
PRPRCV8%. C/EM)]EV,K=:>J<N31DO'F>8*:O^& R_G5%3)L^GBZ^/[T^L<Q4=IZG
PP1QB_Y\F;<N@VP=?;87]'WY#;ET#80\\(-F6Q!K3\@);-X-R$;&_>F[_9Z,3X;Z%
P0XZ"^I(JGRNB&\:RL $?)6-"&K[SDZ:J0P<J U.L%W;_X3L^V^&X-Y;:R_!@X!CC
PPCQ,IBJEKU)+@I[_GA*Y[);?Q^-/V\ !Q:UA<LA5/\/+O/K4HS]J2X(0_ #N[S$ 
P;7:BUW+IHQ0$NI7-[/O&*ATXA'=&KN"C*Z8H4N<_U$G<U71R04_+#SK7)("\P.40
PZ6Y2<>,(+1-$^"*J&WW_"0G@>@.H1WO3Z(,(MF:\+E[QFFGZ2>FFDGULUJ7BUA3[
PS^?@\;/>V7^9+8!$SE/&NT][<UD!U8?O']0L\(Y08?+: )*$62C,<"7H@A&U2N(L
P15X9J3'\$,2X,"[]PLC>/\ELH>S4=CML\!R$\#T.ZE3+^X)KUU(-&%T %;U"%[OT
PMT.7/?HHCL6)ZL(<G.@H5]0!H/(S$%=)?";INL[.F2:7]V;@P7H-BX'.<AA5!] 5
PRV6*&*XPF:32^MENIND"XI>?N81TE5&8^=QKP!5QTR-I\V.US/(8@Q4&Q^EL,D@4
PJ3.^E.F&149Y*./X7#H>QEYHQH#P'KTBL4L^EK)!]:96'&S:'/-K1RFF4F$9UBM0
PMP5SM0K(/R9VW'@%&W/^6M_HJ_\)096V5KG2[G1-4F=;-!9*UKUR16"4 NRS;<EJ
P@6AN$YL3=6K8%&6T7/^WH'+=B]MM_6IQ#-' 9^+SSR\>TIP3XGGOMAM4F85AQ^9<
P F:[[F.&R&<XMNXU9,2G@+51>M:AT,E3PVS/>L*?SU]E8G-,1!UK.SU)0DE#:)9$
PP%=&-TC"]RQ(LG^$/UPPT!RT%MLATTM2A64:; PN2>J!>YT223>R_+;+F<.8IAD%
P+92R"15.,P!5PR-8[4=5PEM:T9T)0@7*5]U/0;<E-(8.XE"Q2KJ"?<G PPD;B-$J
PCT;C>.NA&,2)^6L2\Q&"I[NXZ7Z[VXP2I%O?"S#RJ+/E@)[EK:@%6*Z#D4QS!<!H
P([^#:.860B??Y+T/K<C26)QM(,VCUI)N;(6TQUO8OM<&*<1F!A+?M_>'JR6)ZX"6
PFU.?HD7)RR).1@L@ 00'YM.X-8A"-'P??$4V- &U+?.MHY.]6DQ(60[P?BZM;TP_
PUYN9DW\)5 P1E)-Z;F86AZ*LTRA)VB'JK#'O/+OYCU8\!W%S^VG<[8X_#>;?[3:X
PBF=DA-)C%S%,9\+%R 3@0]U+>'W)BG;M8R#0KRAH#QQFHZ6IUHB8IG?"8$DMD_0@
PNYF+]6LG\)@=]=UN^Z;#$^:;ZSU !+QHH*8+L$;@:QENCQ@]OG52.TFV+" _NP9^
P(":.?-\\XQ 73C=ADG&ZON0\+PC"5E:,6VH>@]^%K"&4)BV5>M(1SM1*H=2G;OAT
PR/X/\RG"9"8RS]&97-\X/: ^B')&S$ [2FGV29';?%T0^P]1FHD'P3 E7$:N082G
PTW,D'8&(G*HDW\KYXGIBQL5\^,TC2@S:QPZUN+P I*PV,0A%DPTO)IV.:;YZ+T1H
P=06DQ:<6R>4P;A6MUX;\(#\887Q@C&I%6XI74+4!MT_RO=8OI]0 2+:)&J<D>?TO
POQ^^/, .PN]#0,UF#4O7'2*+5*_[90V?/7"%T(JP_@D/]+66N'JR]4M\CNQS;_0O
PY5Q,F3&@V+K[/*A3@LS">^5^^JF Y&L!4T<LC*&O7>L3W[#H$D*20+63A\PJ$>"F
P0=X_,28X B))7GFA$F9.[DU&;P='(N&T(H 2HU?#&L)P>/O-/15 H]Y5=HD]>%+8
P'!X)TYSYB$Y?"(O\L4Z41@E4)$K9,$^KQL5\E)KPQ]EE93^S:_2(2,PS=>$\$QE>
P3,N/BG=01#4K6H*XX<(ARJ(DC=F^@;\G.ZJ/U?K9= /()1<"O8V20WSL1P@#BY E
P%@,S#W/&2;0N<9GXYC_S#MPO?A7AO-FVF4!7>GBV"<VQ?ZM"'%73Z:2Y\L:70OO^
PS\%QA7@>WL6_HAX;[W\U7S)[ZB\G;'M;\YFBW^A'O/>F #Z2R:4@U\]M_-E;&,:X
P.LZ,>-.YJ8BBFHBOKCZFI:O7,%^442"8F#[Q?)JP\R$-R:D$%?7A\]JP9:U?QQB4
P"L,PJH%0:P Q;S?*WONP/U<.L-2RTCT)$O:U"\>T@=Q\\J2,/N6E\:R-L$N%711\
PHVV*,Y$G%[7,1BS:RTS\N^7"[>1JU)ZV6 5+6*%G9J:>0GWZ#T%XZ#KACZ1SRE9?
P!V<73VC"+._CK=G*KMNG"!C,VYL^5@J*U;@^;2%L)@C<6.^Q',77HMJF7B+OS@MF
P8H3]%\7/DL,J$""M0F4T2/</M8>3K1&[AJK'E>;=CZ3#$40YJ/_76!D NMK/A* .
P1L-#L-%>/OLU74O'@ D(>N^Q7\E;&"U@R/641;ME0>UPF-!DO/VM9L@X\ 6F -]$
P:[F=HC4='\]M._.:C.B^V5-;F6TJ+!]3@\PE*/#7Q5Q5M@JR,1/"Q L;03T#JBJS
PC4 G:X>-1;QJ5\Y[T!5CVP+E6P@CS4Y8V5>"6Z@[@68NXA!16R6H14,A#<@.PKND
P30T_X=X\!H&$_/P$_M<-!<X0B:5?FAM:Z!<X"24J68HD)>0GQ(U]X#M/H.D2_? C
PKT=Q &PE-O"4PK>J*0JIF^3$L)Z;,@P]9>5?Q?*W% Z[Q,N_YZK'+6A--/B8_^SK
P>C<'L=F\YCI!4S26_EBO(SR[ P6SMDU[?DY*]P4'5@7HL3&_0"]U/WL-WKA2'3PU
P.K&;J<3>BBFDV 2US_]%V<N9'D9>R"G7V#B)-.D\K:7W[G\U9/]66:W'%W.J-7(?
P,\FZA8_0V3,O!@V76\ZW6B0E<!1/;0ERD3[SL(P<F R?6/H6:N^#PQO]B9?I;<NU
P(]X743[@I9"?TC:GMB(S8?_:L?Q#I>G T=6R&1TC]HA)@;<Y:A0,W/]@=]0,4]@I
P:6Z(X^MRZC]A.?AYK @%]V4&TY7 J=&Q??DR0^H"9Z?#?4#OY9$SY>W(?;37D>@J
PSD3-@7ND[(\41Q$/YA9^%,!LWU>-J>(##>,U6=5?0V1\3JW2S8.+-U=$@UP'&1CM
PL%ZO_X=TB97H5%P.XH*IPATIS(%_QIB"\@-U0#FO>5X.R!U! 3#KW*7]I]_^Z/SX
P7"3[MWML!W?TM''"KI@\Q 7@8A"&4&=(U,[F'V_:FZ&R9_W%*<C+7#W^O?O5I*BF
P&ZDF7!1PXI,BL-J 9O[EXF@SR#(6M)H"R><6;OUZ)6BAN?>\W-K<L^&I@(XO]H]+
PYCKL:9!-(!U5L,_SKS],2UWAF+,,J0B450\O:K8"Q6=<L(AR8R)^#.08)81_S,C/
P1HBCR;0]M &H^*L>&.AYI,  7)3+<U?.NCNEA@KBS.=*)?CFO%%7GTK<6#P;PBK)
PF79*/0]C!!5F&WE122?"-)="VCT\KDW0M+KY#V#< %N<>4'?<U9"_D IY?8$";;V
PM3SEXA9<R(/G0'WW59.%9(152RKW9R+XQH822WW<7O Q@ON'V #!6K?CV :2R#BG
PQ4B?4JYJ+,&Y^L.6\4\.3'\2*B%XEQ?$HX#N;+LN!]*L>895,N,;*5*$&ZOG.NF:
P;:O4EU%P9ZFSQ),C>E\-L=E9$@#6C;]9BC8[N$V2Q &TNE <=$PK$1"=L-K7F-]V
P6X@GMP1&'.ZR3(_,8@)X.MXA^&2]J?'^JW=R< T8FT<N7$MV-#]06Q/EPPP)W/(G
P!I=E ;K0SB%%I+P^R"&;';1;=/GIA9<_:D/@[RFS-"JJ_=_:1<CT%-!7EQT=P %3
P1Q=1%@GY)PN;2%REM2V?'>2 >-8J987(1)03AHGA&-57F?D/5,ZZVK=#^41HPRJV
P$;.86FS-,_!FO8]_>[@V3 HIR46R,-7(8S@4[WLW["_)YF>3@^Z#BBM!Y1<MUOYO
PX(JO70<]$V3[%OD#3H&%J*^YKV]_)3[:>8T6M/7M:B2HFFCN("C!>,&>JP;@(5>"
PUR7I\A48Y.44:@493AY;*X+23@UIGN'%Z]H6"M:R3ZJ@%-;1);=E]V/< M-(-J)7
P;MK<L>W0,IR#'EMG;,7LQ%=<-2?W@3H13!_%5"2#0WVO5WYF8..YBN(_C9=IBTR(
P-( 2AV/26RM:N?#9>A8T#2WQ%HZ<CY:FZ;+R[%)KQ"E/R(32U?#YF+%)GG9%B$/'
PO]9_ W^"E[M]4;+I,XKF-#W!&'KVRHDAB!M=/-1A<>E-5GQHQQ($/[(,7P[0"V33
P.N#^D=!ZL70CC7J?0KKY'*/B9GP")G1J%/.. B19#$4H@ZKJCQ&9X<M4I)ZR8Z<V
P5)T_!@QED^5]B(K $0JVB2?/6$=+#%Q.7#GL5)FFKN3R_!<,S>HI&Q=SJ',WXX-)
P>4D9'\_B('?8F,1S@Y21GA.\O#SY'$4Q)ZV2PI-/[1I]ZDM%!M&?-N)-'L=I1X;/
P=5N\0S"TLX^\DW+_>AHXM*-9AE>(",8,^O-]:T^($J)?PM.^JHG=R?+=@N<0A >'
P_&F%P"F0/V9MG]T?Q.S.2^)A 9\E*NQ.J"N5N]V!B(MUO4%GFC_#XM;B:I5N/!IA
P]@59?LLA3Z-#^)N!6VGE:G>TY@A.#$.&P Y.HUK 56?776U&A'LH[8!**1N[58#Y
PHZ/$HB>=(*DF[[.9[1H<JX1&YGS\/EZ3A@+<"O<!"VH0>H5."@NRP;.)A[1:R)X"
P<D>;'5M-C6 XP.K<O)76",@#*!\+&7YZXDZ-!N5\T/69_FW<23<I4,DVK11.!T7+
P6!O&(O,G\*.[$Q=UEXR2$7-0E_]'.C EF#*9Z4IIRG?+S]:WOS%B^\X8&&6&/'W"
P,GLR-'Q13YETO^_N%*K^U!2#?]H%T(EOLT<C:64@*P"H5NR0RIT';OG,Y'"V'%DX
PH^ZX2*\A+<YKWI).Q/;6CL$ KKG7SF>*!5XNNZ/QCK?KU#/9/OM$[ I6.Y:/-L=E
P";O'BW':O\,]U@TR2K%BF]UG5TT5D)+9? "\+&KGZSNVK$L9'V36MR[6Y)SEV;=Q
P[U)*2_Q$B31M>!UXP@2]\KVL/UPAS%=;V)-IQQ<MZ!W=:#2BXH&U5X1@HXI=1BOI
PX3,A4T1&4'\8(X,-@>1^"GDNM5(/8QG,!9M=Z(0V(SA:?Q;/O["^OGCNUHB?1$&T
P&(IDFF131A^^1OQ7.(\73MHK</;GQ$8&'_:754N<+%N 4^TFA>F/^I()8&?6 ;8(
P"$>+7]TR=!^'?><85R2^.3*=Q1;Q7X?YDEN#5/JV$'GA5;OLT_)U%V;.!-Q<-BS0
P&-S1*FC<V!',O9W=W<-W<-EFK^(LZAK@A@H^UV?VGH"7Z*)T0\SY@=V_(F-1C])*
P"KZ),S8<<P$3N^SWLV^S=$MNEUT=%L?V\X$%AV&(JW8I.W[5#+:99"25'GC_4N]#
P":S$<%*V[@SE'$BP!(1RH/6V\#-JA(A#1:U.]F,X;:B.GK4KK]/B<>,UK$CJA_*I
P%9N_8PF([YJZ SD,:Y91T180>/ K==RQ%H8S,GSI@1L(PTB/I%(.$'%R$-3_K?/L
P*$1T#[(;QSU/E;YAZPU3R#O!7G]*#Q+PEIK(ED-)PF$,!&V4C_!,,<<I6^".]-_A
PM1=:BU*&]B+QQZ)OUO1W\T>]"*$/IAQE.D\4SYCP^[$[I#7Y/JCD\F*'/)K'I$:Y
P\F)<S$M4*<XW5D168YJ.WFB69G><N \BBCM07,-0/1U7D+60@^9Y?4R_&%:[W S_
P_Z)R?>6MP2#LG5C+<63X&"4@@WGY+VM0+!?FI$B:($3C=W4\PU@=<UC0W>UX(HXK
P<,)Y<58WN*M^[:0*M ##V;!XF"E0E)N.5>.U'*\])R9.Y(BO:@5O0\_SX\@M>'[B
P>*8%]#'^*]^%/O#:%P&Z$$";SMZ4_G!QPF/*EREX0X-4:X+NGB"Z(D[HM_GNZ)$>
P:MO:GP-Q8/:V-;[?%3)&@"TN=:"L@!,S02V#D,#ZFW!^9-C2JX]>@1R3<3> %W"U
P3]$(/RK7OHRQ1$I8D3N:PV(<"N,+3.05[B213MSQ$EQ(#S?Z$(%E_!1G'CMM;N(M
P[E@W^9X'CEO\"I78-+KG1MKNF9L6F%@&N9F:]*=QDXZ+T&C7E7@TB;8$U%U_E&&&
PV(:,,GG*+T)DEH0A;#LQKRT&D$WJ0U?$O[O"A%+*/XV:>XJ&5_Q5"^96EDZY;L2/
P9G5 _@;38B 25^B-[&*,6&2UPU#O?4]=$3HO!\U-G4ZU#S[_MF6N0;,8]BNL9KA9
P[5+I@DPDUJ=>[=O*HBJ+Z<L=!)*HRS6$]&E1P@BV([]13[#3@[;S5-6&/G.$[4H%
P27G<VH[T8U8]S*(K4ACM0H:+GL!FV4N2&JY4^Q4\86!A8"Z:[5)3^..#MKG7QUP+
P% ]$AIR:QE&SD?!AG N&K_J.!E\;5-<F.G93AT 8R!98I2M>WF&L:."Q:*:A(O3J
PA#U?ZBS.1?DJ'H=+_2LE93>2;"Q\[%Z@.6@\=6']<]<J)%!2:,<CMG+<#!0)/U?!
P-B-CV-;G?\0[>,;E9RQF'JMA)TJ^[1?%Q;W'Z,PPQCH1"^>6WH%,[NJ&I!?2JFJ+
PY+F:EU+^YPHD=%;:GVCBJU1W)&@+BR57#"&PW[#+HLN=,\DZ0T  /WF(MPW0^I?U
P'20&:8"BJEW%Q?%J.U?Y03DA/WX<?@GZ@TR'@?Q*Z1A@2.QH6I7@L#P/)X3UHT2V
PO1CN$PMP,Y>UE#;33!9%?2_;:R+Y+FO1N^LD^\XQS@?C2%K(&#Q;1V>^3]]<O+P<
P9B3#9Z41JU%_521]5(%SE2[MRPWIFP[NC,(7S2S;<HY_B^N51X]/M^KJG60\H[*6
PYL]>2<DE"3QW[&0[9R2#G@_8_^5<GS?U,I2"#V4*^D__4@8-0M@>272S4^P0U]_>
PS(JY:U].LXY5,U=8Z8.7+]4\NB&*LG>Z_MW9/R9@ZY28& ^ 07H".,QF<AJDM"0H
P=$(SL\\*P6^H@MOD[KGJN0*J=(Q%U"_?1WX*&%[=>R=,-E]T4H^H?FRW;[<D,I/M
P?^_6Y^:]\B]0O:%\/I@,F6!T>*@O=7JU?3Z=Z.1/J3T1+T<F&D_ :O6Z[<7JUI.G
PJK/8Z4GP.8P--^:3,M##,3G^__QL(D2D+&V76'&\R5\Q3)*Z&S\LI0^>#"9..=8 
P=5;(DC-%'=.6O(2W 5K9:^\5]7]1H5?G]//L4D-*'4??.<,,04+3=N[32OO.IDIF
P,-@6EHR#C%)>>WLS8I<6XB6TC/K>1T4"8;.;4)P1*:6,:4#-1O%H Y+/HZ.MJX$2
P>4,!UH8\]W3M6KZW=BM?12?76$>\%Y=-0 'F?PS>]78E5G:N><A: 394[Z$I:"F#
P4\8<Q7(ZZ61>_ /KP#2Z;K5WG.[-"WB.)#T> H)=NZXA[LSFD9U_O@K:9-^:S+&N
P]Z7RA*51SF"<^S4#JK5&HNG\F]V?J0_E<W/!1:-T+US==U_0V*_/76$@<XQU<  R
PL)!O.3!%S*JY6S\E6.SO<D:]BXS&UF$SL._ 2'.NVUO &DG*I8\]HSA-)*/A%3&E
P66*?'N^=FYNGX6$?T-Z1<KF#Q#&7Q-$41&F=U;_W1G [D3=!KL*>K8U+O-FA:ZIT
PU8R\@9^72@W&?D,WGU(^VU3(AA#S@)#"F+&T"%6$J'S41U=>0O6%9['1*E,SE10M
PHW(1^T6M#<D/E$,9,BK@5R4*24J1/A+2PE9'X=;71DB$?-@&U(>V2'%," 4-(-JL
P-;9MII]]=]:$)D4A[ZIEUF6S2:T+BB>"G-UZ'Q2E&?L211:D07ATF_[Y2HW8/9A7
P-)S<REEAFDK[-9+&[":D%L5+R1FYU&#UOA&@32Z@<F<SG@W!L3"]Y2YC]MU'Z(HP
P"@,R3RJW9_-:=+SFFXU[S=_;AQVI*+<Q_!3:'@$ O?1&(*BW5#9&1WK]95M1& AI
P<^(3P-\:,^US?&H"1M&WW/_^[#7C[CC$/D:_5I"+!]*(>@=CV@3Y.NKH*)GCM2+F
PJ*.5/D"QUJJ8&U?ML?93KN6)L;JB<K\TAHCE#0%98DG-"G @,\!.QNSD=ML3&;XP
P#C':%SE> :-KD?I[ SR42?^7PY(A>1  "?+UUC,U4_4.SRA"@GPSS6@(TSQ84R'P
P\F3*&F"? 9\$+C*&\>I+,F,S\A-J,_'FC-X+3+7LD.7$E%-0>-&3$:[2IYA/@]PL
P_F7G5="9:B#U"6<"T>>L/G+>>^8<"EI"43K9' Y*#/8MX9*6QW8A7T$;U$0]BJ_[
PS].#Q:AZ588.?"JN<1*NL$#0VP#)Q _-!Q)H4HP+RY5M)>YS<GMB/Q1N;UY'?,$N
P*,4%QY"'_N^+D?@N=QL$SU)8CHE8Z5LOEK=<(AX=V>HA<.UAR0IZ->[!^N3-LOEK
PIY8?^#JC<<SCRBQP@B?B?1%VX:@7/)-@]Z:#7KYJSS=2!!2.M*OA]@7(QH'E'J[)
P<N/O7RZ.J<N[PF19-R5TU;YS^N0I6MP0CK-WW-TPJK16>\N@\5X]P<A5T,;>%%W"
PZMNP2 V;_D\7K.LCAC#]0^=BP2]Q)6SX$1T(Q&10[$Y-,[\2TT&^[#UN5UP85ZF_
P>G(^)( N3UM1?%8I<F"/Z$>$9F9NA;XU_^+ P.GRK<WZNQS!VBA%O@NE?V%MF:7M
P1FN'F()UUJ.303M&YJ")OO:/V7>Q!%F+\I^C6;_G0-A"5R^P'PG2^N2@ G=Y^#Z7
P:!VB;?T>4P=G&B>*WF8 S1)!_]/'FZ_ R;,XQ>7W$!Y3LK9+O<_0,,UWQ>X8[KCO
P!"+0R;1! 4^=*>O$6\0K>FXPKU+;>-S<D$B2"+A&$X!M T@D@3(N9<%Q,KG#.&GG
P'I"".:%P*>J^&XC*=L11MJM74A?_,"@"Z1!C5[I/_9&@( O@*I:B&WS/00.J%Q Q
P@I U0Z=4%7PWYII01=(,C+<<DEK8!,WJ_Q;RU&[$1)KE[ZM!O3EF80%;WV,&![.C
P >DBAE@J)_LGK>S7*ZWEQ71&M+.V*U\AYED7/E'\L7 *GT!_X=5:F/YC8V!_"_!-
P_ZZ)H,8U0@OUJ_MRB::-!B?Z<2/,O8,S>N5.I+NB9]AM09^]A%Y$YC7_@CO ;\(6
P"K<S*H&*E8[I+7:&WO++43]5"(=][OD46-4*6A\%F23,$>/YVT1YG,+:EP?0"W=N
PD$LU+,BL0T+4$D6_P5E2'8<"?FU*>MHSV[L]0NE'PE'NE>GFA66 V 448H(<?FIF
P!/X&EE[R*<(\Z:S:CZDN\[6;;,TKQ2A\>)M@N(0,9)HI(?'@9S_-7IZ<%%?=)>N!
P'Q)P,OI.7HQT;<CW)I]T2V3[P%HU[#V?^U]_?-XF_)BRE2A!X1(>EO%QX->580?@
PLMXFC4/M$.#EUJVJ\<5V/JR6LAOYM.%V,[&P0^578XV!S$E.$S)P=$KDH#C:D=?3
P'WKLYI3V-E@:Z;/7AI:J< NKHP5\+X,QJA#(C.49M7GDH-_:"V0-2(UY9LJ?F#9>
PSS-E/IZ3#[Q"14GC+B;,4QIE(.D(?H=FU%$B<JS8JAF2Y)B)&N&\>X@)]KT;*478
PEKA(I0<L\BG@=<$,Q 76,HX M[-\ V!YT?[0P7@B7MVR!)A*.6*^!P/!R0-%I>(\
P@$X U&%:J%OC 7Z5L=A:2-T@3:@].S9+\38^<.H@OC@U5T'P-=7F7WJ6*^XPD69Q
PVE&XH:"A+S,VR@P#)W%E.BYVGR_J?DELC51BFQ0%9$T+?%2%QDJ]PDY32ZRI!634
PY=1K.TK46Y^&ICD(JQ]^9N?@B#)?1XNX,KAT%:+H'&K?\V%^ J0UWU6G\E2U9'>6
PQ7'Q?^UKN,/79[)5>*COD>[,(]1EK5NM6M2CQ5[>,%A\L0=[>O$D'QN!R6W,ZQ]-
P(%RNAEQLI_>,JN+K)C?E0M32J-5,'L_W7==>J3CD7)U"TD_\9XK \TZM9UEWJT9T
PH#=N5J;M;$X*IME?5PZ15P>]2N!HD\L32@R&>3H:!JL3A[U$ X6&MQC>AND'H)N2
P"9#>8\C0V+0G-L<;[T X)L :V# 3"7Y^T^!(X "(4KAKR(SN(BM>H\?-F;Z.^[7#
PD1X.[O,$UN!^G ]LO.O*YJ$=BKX$;=VF[VT8C*=(4T3U;CVE)[R(?03_$>JEXK7V
P/P%8L@AXV,E92>$@5B)1F;:@(N]*0 J5(X6.I($AGU2I\U+=U;LW7..4PJ-2\K34
PY11LNKHP %NI"'0U=X'NUB1##:ET;"3HER_020.V2ME!($JINM/J;W>XLLODO$W;
P->8+@+YB(5S@"NDW+'K^LRIHTT$/-JG?&.4<M<YOA=!!W)A:LD;?EJ%,@AS]8<&9
PHOM]I0+T#%V'>=,/?Y1ES?D5\7U^@QA)?8V3 \+,G4 ?DC[,6I DQ\/+).#.1Y/)
P[M"L;@GI2AT&7N]X>9X&VI^=C)^RL?IOU?W5]?& BKH!X]MMD"B;#!983Y:5?8>=
P,RF!27'V!3YV&]#?+Q(^K;%RK+(/=*39E3C6/^_SIPDV.9?=;;@$YW*7 QB$,PG<
P''RP1TX31!VH$F)_94(,;O-SQO7)J<Y;*;,2" !AO\]K%38C74>1KC^<L5_R)%8,
PI,=KY5'XB[CQ L<?%,Y-\]9:0ZG#+%V 5.T<N)((<W<H LZ;DC3@&,!11CWV47PK
PT#YR .!4&K49PDF]H#6K )W9E(",!'DZ R;7:42?;]78UE>$'W-20PBXYKG1'_@5
P9$#"&:*E/?65QF</#@(HJ-K22R249K^DE 5)9>JXVW8\K-9XV<U#"8,SUK!:C,C]
P91/P3LQ" '"OJ%<.OA71W6$JT*'O7-EL TS$]3[4"EZ/=3&?IP>EH\Q_X_NU P9Z
PZW0VUQ-:VM<<FK?5?=]:WRQ#K$AS"\.88U_382_AU<)]^$!<>IS" ^MNB7!%TW^*
PTX8XDN59PYTZ^994GA\\3]UA1J(V[G?$)L K>NAXI[-C8?YOL4'QBR90TO\<WF#%
PBJLF$Q:Q3?$Q+9:Z'!6< 6E;89#]0]KK]SH? Q:-D24IRB(CN$C@7-A#Z^2B*H2L
PW7&\_R:?LD?C4:7G@9:02K*1#.:?51\CKO>'5(2B<PIAF[F>[*W]7GL5/.>FOT;6
P9>CNU*.:K95@[(+M< PP@N1J"F.#\>CL8L<-PFM,;7QH9@H,@LR4!#X>NQ@+L:7.
PFG6$F?WB345D+3>TEU4$I@\81Z)M5>0U $F(WYF]^ROWA=3BE;;##/),AN.V)IM"
P2R]D ,&,TJD?W9/\YN D3RG L&!8@>.]:P'4;OU5*<B@+R9;S+0C'>Y0>C@O2A&/
PM.-ET5R1IN6T36;0&HOMU=N(?Y8 M-Z\7L[$%D!GE^L8R:&=M'#W35^.RT! ,E#F
P<P'FQ 7WQ7'[Z<H/JS+&8]L4R.N@J&O8A01 +C/]DH+2Z$)),M&6CV"5&ODC1-[4
PIOU=N\VVC$.!4*![7T]N07M\$;YX[D'H1GBI%CZ2D*Q'PGQ@MN>NE84G8.; R!.,
PN?02K,H?3@O-1L:N+2L"3OVZ'899_@PKR]'#5JT!FBE!LV UCV<_(=O%@ M^\H8%
PU9(W/-S<8D9CMP]"J3"H1N=:KY;_\2*EO(F=3,.#HDUU31WQM4(0I^C<?W0T"J:9
PH*\:W@\;(GN88JYV%&-D5.+%_]-/7^Y-XA.TW0*,%YJ7HZD1<#:J.3)T-<%36-.O
P>2:_;JR$R.1@GFC!=O@=_UB_<:"HN$B*YH4F:UV.EWD[DAZ!O% OG/@JO*=UM9M#
P 7F$KP"EN.?*E@/&8*@2:$FW>OJ3F%Y"L$YC@KSH]KUY:O[^PLWZK[^C +J,-*OM
P\5(ZV$P ;14RA SX.YP9(NK.5?8P<M=?IF'25/W62@FUI+#FW_5;+9A9ON -)Q&3
P'8AB::E? ("[SI0:[5B*&2>5>3Q=D>@EY%I[ !*6HT1I$<1#7HQBN*QM&,1?P*K?
P5YGFE9H?R6P]R4!"^V[K[XCT3 I '"<2H_7N?- Q& "R@#.%D, KQG+8Y"7^L#QU
P1>A;]W$ ^[Q6F2(TX',%(S(=,GK7G7_># RCUYQ43<\00H=S_G\);$U"ZE>1/?^>
PA($6QN?K8&A^N4QQ\O*!3J[_1YXQYUBTML[)G&;+\C7H UC6,B7D78/IG1##+0N<
P-[5+D7%U-T>@4I^D6UB2Y-4^-E5@M\ER=3@2F ]MG0($X.L]L,1.Y')FZ?E!QT55
P;NR"K393/PS,6/!$75&9DX]#O#:MCT*])N=E< WB-0L[02LXIG=+!\R2"'P8Z+F)
P1,"*^[[A '[4W(3F0F(A?T(!#LF18*VG#_H*M]8K[BOHD$JC%P.?W/4"]+5\[_KG
P%6M;^A= 8]SWZ8G3N7N6V@Z*2[0!'!>7*R%:)]BNC<A24W#),26&J!XUEVXC<F(V
PR'+/B>Z(AGWI04W1H7W;+#=,'ZU).?0,W $CNTMM";W!B[("O,8,0WH4?M&MC[.[
P/3>HR[-/?_WF6=1TQ:)65T)5%IZ,%KC0W/O^G3FX#;3@D&L/# 6?4B>M_H(6F0NR
P1*LWV3%]G3?B^BL1+K;7A/.:^=MZ.GV-=A^,'2>-"Q:V58]D7_^Q@ O5F*'V.VCW
P##2Y7ND>KB.W#]H7MBQAQFMJ@F+N=+4,WPL11T2AVMC)/96S,'9-I%V1LO);=DA%
P37A.$XI(^?+/O7'X[;GA,99EL5D\XC\O5W249MG(%F/7!78*KO4QSOUFUFFZ1#;S
PC-X8'C]@K2UV %G_WG%/_\>:3!%I7U^; AD5[:4G>Q,V.% :=IS(0ZWM:/ 8EV+D
P%G[\#7[%!@%D=TR73T#S\M_^F"N3$/BC12)](CB!:=M<,(Y2Z<C:HO!'TK.#P_*"
PZ)5AC2Z.6.KM=LZJZ;/PPPJUZ]?0B(@(4P7P&U +?BCA79.6B2>W,V@$WKY_2##1
PA:NJ>=KLXP9IT]#M7UM0_>.;H+ \#)Q_,_RFZE]9++QO&#/L,%U 8K,\:1M<Z#XG
PZL@OK!7':4P_BB<]9L4P5*/ "S#[;5E[W'7-]^G3B.2[B?EGFRF?IGK@D =>L,ED
P%WF@4_N ";9]38=52X4&803+SAN$QPQ\7P0!C_>(-"V^X8^%18$\JY^K2;\,VZNM
PJJ@)MB4.BV2A#+;.ER$ )>BL^R1/MEVLT75ZV)FXQ:>['=_+?R)C>*A[)0F1WR"D
PC'#,*\F#=0Y$*Z_[$G-H%K48QI OU1HWL17($Q$V59W:RI+SI=1ZI*KN>KL *;(S
P!N.C)[]_<L4]CD'ZE6(9=Z:Q.V#V^VAAQ>L3$LS+K3'EC*:CM:. *I*>Q,1P2J^)
PXUQ=%_7K.]EF;"(4W+\NV9W-6U$_'YM#;$]H6MD_@3R_:Q1H7]D&O<?=V7;@[FPX
PO)F'PPLUD8SK";ZTKI.-L, NP>O]\U6IGE)JR4@DUCB"F>%9U#*@9/M4EVM&[R$P
PH\;ZTL4MEO3&:$/VT!C@LU]]-?0\\Q$?^'^:E]Q>N/&S858%04Y;(6<M_G2X\91L
PU(&+\3*!]RZ!O%(XCLJU%N\A"U2GAC8*:#7\F>/6XB!,5C/R %M 5Y*"=M[6P-+&
PF=;"L8MX;#<A-O%$J:Y[QQIL\Q'[\_N7[@%A?4)V4>J!QEH?+$\U-C9!L;*@*GSY
P1B2.@OGUU-^'@@!-P\>=F<GJ]5'H7*&&_ G8GI-BS1GJ>V@/\X+#RB5V>]7*N'W1
PES0(-RF)!-08@(N Z[13Y6H84KG >2$1W_(4AJMO$WQ^'VIY NH0:\ 7V1^.&Z^/
PH@\#X8]H(<2)GH>(M.RWI\'H+;GBMU2!!OB;*J]N31OI7ST'UT]*!,%0H:'GDY>V
P^!HMZ/=SI$QWP&#RSH?6N^%NJC O,$V!A>;TP"[=-5)HGL89=5;I1M,_ZWOSZE 1
PTQ (#PS; D=*5JZ('ZL:\T:.KC+?]E[.057(RZW1$ 9R7"509 5,G4U2SI*7_EQ$
PG67.!B8@0LN5Y!2F-5_9HJTD%R:4JDR;E[8\Q6%#2]%+UDQ9U<K]1AS\$FE@/,,J
PI)-,O2/8DN],@=;!.@]Z1OD ^"RB"_ %D!.E8QK#_A5I.>!(3"*EJ_</@=MGFTKQ
PL1%,7O5WHHBIRQV)K-^7DV< 'W A.43QR5,FAZ-C$>8 _M0*G?#,T,T?V-GB7-])
P*>J'@/L49IG6XRBQ1ZDN$JA7"'0"NM>>4A5QRV789VS[EJ9=$1#/:2H]W<I+DVX-
PK-VE7OBDP2P:H^8 NG2N_K[(L7X^?E?_&_N71VK0M/_>XKZKDRK;["=FDT2SAYZP
PDG2C$R(U(JU,T+ HS@O;C%A--_WRSWT]SU#?^W>1K%O[^B"],+=%L(> [$Z=%I!9
PT5AM$/EV<W:NTXC&*8 'G<-!E9%3.7&"XD?(1A!5O>DG;()-%^FP>$U%[)IC^]]V
PG6X!P)R ^A$N5K[6#FT;C6@ZE5I;:P.33H.9 J0??S>^6@[3BJ"6Y_".=[>MU ;)
PUOR%A @F$.L-D%%.KM" I]7"8?J.MGG%!V:6<"+H-'WYVUV2)V'HP@CC5)*&9CLV
P- ?<+0*(T.J5Y^IO$<N8YB5]:L:NGJ;8\+*@MU"/NR=:G3 NFIN]U3HXW1PBJ]U,
P<YDT6=H/DI?O%*4\CW]7QGN4Q,/(TBO\E/#?I_EDY5^N-"Y'E(H+#Y0HOQ/F0SK@
P ('U3#ZD+D#OFKGK(,HD7DCF")^X\K3I=FUHM)C]T(CJ$U"KU2?CJ=X"+<Z#?.%3
PQCX]2B)6@36$#>!VVT6LW%_UH%R34RC 9E\/L/49NCZ$E=57(MS2V/ZM=MM =HPV
PH6_JE==?4CGNH"M'_5&9[,,3&=+VN^EMB:\(&#Q'VA#^ECZS%QA;,%7E\3W"(&_1
PF6(#OU._?.95L+KGG\GQ!WDO:^G WK+*B4R:%X!E>V+%BSW==\P!#1!VVP@KP=2&
P3N] 1/\<!)_L@YU^('3S<&H3C]H&*U"Z];38<J<C"7ZN?F[.\M/[-WK]EX9/ GG/
P0@H_F[)0'19'M.A3=,>D/HS83EUDM=T=^0KRCE?T4\YHU+_I*V8H<>3<9QD"1<Z:
P8!G;]8RQA5*3@6EZ_"B%:6T.L-3)J"(:]D@,33/([?99TO>!$R1@MCH2,1HQ)\!G
PS,?06]/$.<Z+QQ%/$?:_UZ8) T=CTCN4"JV^=/HAXY5SSXW^4O:P0=+K+ZR+@+!K
P!*=[\;H5R2YU)#7LTC/'/8M0]@MEL@^,\!"SJY10_SL17_3"+Y/:E2;U#6"0]11'
PHOTOA.+&'BLAH,X_H32&6477#EU*F'QEL'<\)BUXS6L!68-Q\A_%JQ$U].$J2@II
P[,QNZ,>6(UU,'=8C3L0.TAF\]!::2L&=G8_R/>7JF*Z$:K%Y(Q]L43*@KTI W@M.
P+21X+:9G6,@RP* QDF/BM6SZ^</=4+I:?"]'RAIX0MZ7GYZMOK,.B5D]7.K@/5VH
PBE(18(Q?G.&LY+OS>Y1#',;!,+T>#0\=2H'>ZM;9/J^H6/04^[*,DNB#VS<4AQB_
PS64Y*6<CI9]TJ B_RS2FFUC!)[SZC"YF/2H\G)+7-]2L '?C R64_)MMCB'5:J(B
P=:5+X3G%*$PH7@@KB6:M1V;/=)QNX%([P52GU7>7<B6 &:A9!VT-U_2Y#'_T* (^
P.DM7HD/43=$J2@V9Z1"B?2.AKG\XOPBNR=LR[$"XN&I//++D+;LNF0AT:GIX?I4C
PX1?B"@,@M$W<#8SQ*,].%BYY1,(K;G\PQ;BVA[TQ^/J?P'OVUL6B*W#ODI].;U"2
P[$ >KTH[)O#U!(R^Y:*TDJ<]41T)!I/[P0M^2*H9;6"DU1$UIP^OCY^JSF2&I<G?
P-&2-<F9B0O=ZXX1<5TZ9I3V>WY4ROTG9E5\OF?P5O]5XCKT*D^]JT):$.<GI4._+
P RI;V?^6H>'Q[%7E9[,SBS/7HS(ZS'AF)7[E0X?N\('2I9-W%Q5."J5[54@U[1)P
P*-!/*Q[+G1)\)"&#ZTZ'^FD868JR *8@=DZ:J@Z 0FKN*V1+M0:32<SY>><<8D=B
P#$LA"D;UFTL<<6#%)0\]A!H[LWM)JG[Y!BJ5OV)6\N>/=PKO0MV,M>H;"X&VENPU
P,%+^F;^*T.O7*@JO&V)T-G%G.&_<31S:%]WT M2:@=0T_TS^R6/-?2/NND05>"(9
P*:2+ EH>_CKU2@LHR54CB0.@7,.Q#>Z@/!2TRRX![(P38M)Z+WEI_ U4,AGI@/)X
P04/QT@#D#*P)8?I)70JS,6NL43N?Q2;I:5BUM=QDC6U,E!>7?&SL].>BYJV YLBB
P3KU&?#9HXQJ6NFA%^$<6Q"<%GEB]1=U[&=V&W%6Z.K:*WP\^8PKV&],:<W[)^PBN
PR>OJ_^($P,^4_M^GA'N_I@#W/HF*04>@(^^"<-2@T^2"D!J$OC#V[MH ;AIF:?$C
PM766(T8S$136,H;>"SIUKW;ZI9<BVV4ES;AM#QD9" ="S\3"[:U#-7>0]%679(^A
PLM? J06=_0)3J1R6+@/<%.^$P X4 WD0C/EW6@XH6NUK<!#DHYZD36TJK3VNHKVF
P3<O$]>/B94@^,%-3_ K\A7_4/7*&1(JH[7IP0='C]-#RJLP_G@(;E<GOI^UXGP7H
P<G8VT6-5$VV%&4/A%X0'W$<,[VEA@@UQZP5LS>^AS+7K#U_(7X1\9Y?W7O]*4@BU
PYUO!=PO2.GJWDB@3-QR,?;[GY).>-+D,@8%*:!R]5 O8]+0>593GV$H?EEO01F1+
P)QO#T*>KSE])ZIO-:;1=?JK'Z?5;(68P$K/)P+.GQ> :41<F*A>)DE"[&#?*2,R\
PA2D75>#F,*Z&HAWF5&@)#MD\70KHCUI?]\H(\L\*5(HR'AX+XHQ4*L!QFDR@:[ZN
P=JA(OHG?;[)/J'.RH92Q\G/DF%O'M)-[_%=T/X;/:5F6=T=L/S8%J->0_TC)Q!($
P[8Q:ZAEP*),FY4^G=9BRUBE*REFX@@S]X5,=<3VXZVR'XM4E($PO<TPLQK=ZA+2G
P-Y<!655!0/,,4%#3-<?5( &OB&ZS8^TJ9YXPO\,80>8ZW91<_T95)C*KYE [5Y"(
PUDT& ;HFQ,1^,9\BJUJD[#FV>R[6RL&/MO3RRN 5FZ@+,'M(9,C7MJ S&N$1#%&^
PX1<7C@OX8*P^;C(J3B^'6BF%>=[I5?D/: 4_%_]C_':?-&UH17$PE@.".AL41<?<
P&\A6,@-:PV+),-1X@7J@BVV >[24?).(C),+559++_!G2UP7.( TY67MT76W>++A
PT7<'W2B$RAKU&HEQ1KVS)@8<B'$D80QJRRBDG>/J%Y&#/J,3(;'1P M06[PYD6T8
P"V1Y9LW5HD%O'_&S;E:V)007/6J<R4R/ >U.?KQVR4_":JH@O)1XR7S+EK:F-T.I
P[1"0ZM3RF1S$393C2-.'=^7,O[*'BEK4B>Z>6FV'8\HRH'%;3(&U=MNFS^)TL(9F
PKT X4HKP>50ADA,S^>*37]*!0::_5==DE,-/[;D(O*A)@^Q_%O'.2Q3L-\!W92P)
P'EI9;:E\&^7>OID]*_XHM0 ,=?UBR!.^'%6F_'^KS=#MRSSB/WS+NW>K&KV:KJ'L
P$%:AW(NEA,^V4,CO8%.].>^6-Y6Y(S+QK2N)4OHK6(=RQ*-Z/,UX:+CH1[TQ8*V=
PZ*_SKFX5!.B?+DVH/0"_+&:5)C0ULA5X;S/P7 S6KWYP8N52;?3]^9/'D/8S).V_
P@5/@KW+AH(F2!PR//OQ@$8>8LC;U?$2(<)844S:%MM(8WE!$J)/4^MDV#CPE!\]0
P!C ;6<GS1&JMQ;CT.]]VGC_W(PH)G#TH"4XU@%V7D"$O,8G-H^=)>&7A'$?.VW%)
PDN@6E?TB&/T>)AJ0.>* AYW= 31QY,$;2$K)7<;"2JH>4886XG@R: NT"A&8^V$C
P0=OC_OO=W"G!U6M::N8/YOB;?46>L,*LW(0G\^>%+@W^)"Y'_O>K8_V_F%\*O:TL
PSVZJ7-,5^-MGM^(Q%QY#SC4KM'UX1:=_S>:XO<<U5Y3&EAP*2Q E1E4!XARO#+B3
PXK$T,9O'/(EF!M!I*GU1-)[(YAT8X"# X%K@669W@$E2-'<B>8=E8@F346.E.UH=
P8N;<>%/T.J<F>SW&&,JH+QU)^G/E92!C4)3;[\<E;_Z*[0A6)/>Q6KMYZF@[.L<6
PX+7.VD.&#/!E&G6G;=H\>^'>54KM+8:G%.U[GL4L8P8V5,46LU_CAH^P]VOR@:HR
PJ74\V/L@8^,*/"R#EA\_K6 4 /-%RO-709;0NEX27'=-;V]8JQT83\,7?>U1G'+(
P12G>-U(_O4;=@ =) T3H.^%\*,@OI";-UFW(UD W7"IEPH!C1%B<U3D>!#JA9L<3
P<L00CG!P[8(CMOON4/97GR8B+*.!RSZ=R[QE<,P!ECAL!ZVFO$Q<65JVSCU97YF%
P//:-6)7.M WS#D3,LA.'.W3'"*<0)0%/$G@6)V%);Z>A;F"28\^*'8FFYRRQ>UN]
PPM_LKKEHQ0HA?9[\IF8?*F*TB >!M7B#W3+F\;EUV9!,FZD!3'>D*],XM>G:K2>'
PQ-D<Y3736/L8/,$#<#4$) 5]R)M7UM;H3P!TNH O\=:YU=7!:$8$:JPPJ<F@RL' 
PW+2=]"9R67[8C3J;_+I1_K;=SH.;>I=@X6$M$EAP 0QK)0GFG,E50H=/56:J;^#\
P<'!"\Z$?A086:E=-' HZ&]X60Q)FO#='F9$XTND 8+-K:,L;328.(*!XL=1ZYV\-
PV;0UNQE)6NF-)F@K9 D5ZPPI'= **H?L':KC>@+6D$,K*2-%"?V2\Q2G5YZDE4<3
PK:7^M#)3((,+&[![]'!V^D2NN*:8O):61F3O>*<\H;XR2$#$=@!F\VOFU3'EI B4
P/J;-'ZD!&F MM8:BLVS*?A"4ABPT\>JH!2'FW[R=34_!8P'6C8("HIB7*,_3)S=O
PEHPZ+'=RO.M>Q3S_7[E%+T-!\4N5FM]T_6,@*GK?/AFUC-+/0+>+OUV&>8L0:?S6
P^RS><K22.[L#>W/Z6;,:(FT3PF/J;[F 3V8B1WG"'*^FWZQN#I?5"6 <NIR%P<0:
PR>&%F$\[K^Q+]7Q6+OV;(QE',CKOP$#-Q.I 4ZZ#M'FB??(I=(4JE@=^A[J=UGO'
P)[_A^%E*TE-D6*TQDD<'CSUE4V&5Y,^ATL[R&W=T@#@S0QB".I_GXN\@K(D8JN12
POL3:/\ %]2M%0E=Q>Y+-J>@7MO[HS*9S3;2S/.F0'+A(*EZS<KO%<EI?/;@9NHQN
PQO3T\TH<1T@<'57K-$4 EV>9%D#'TV2?:Z.C@T88G9:W*PCAO7NQ<+ER52MH&__<
PU]+#Z?HDY1@ %AMBZBG1T3WF0%YAIJND11W;UG4( Z6AE*V ]9@EK_ZP*[D/ DJP
P0MKK'EB/=X!8G) T;),!-LA8@F@>)-B51;G]A_Y.>?+OW$GUYFV)C&;(:;<'"K9+
PR^G5+*BER\JVW*]L"XNRC=_:$$);[J&CN3A,74E3M\W8,0<"N*_%$WM4E"ML7Q64
P>4&ENYV9]#ENNH[_&I9*A@XC,P#<XK3UD'RL[RZ=X'60#779<-<S8IMHT<4NFM;Z
P\-[+'L"6#/AWFA^FR(=?I^FYP>C7\OQ_]A2&[I9>OON..V!^IP TM!:RW \X=X.I
P(G"$<"#+SG*H>OK<C"=-IP6H$X#-G(] H9K7@HKPX60  _(E"N=4<FZU>+F\NM4O
P2FVKS.:"KZ,L]MSF=EX!ZJ;JE.IVBQ_U2\*$+]>#$*-.DE5O#4H#ZVV.B]'7N6D*
P;5I>_P&QI<N^Z+?F 1WMMH=;/OR'4%^.N?XDL,^EYSL4JA.K0_DU1E0.2(BU_.,8
PYO4B[+RM/]-)-+!M=%[XE39*3R4]</3C75RVP/:-0LH5AL" BN!S4%/'(*5Y!YYB
P:CL^_ZV!8UC";.> #JZTZ(6I/X65:W4OVDP'L^]$UT<]=E?DP("TZB^R^KT+Z@\3
P/' 07A/LPPQ$ D7 +1>**?W%RKXV<D8D>ABV/3N6%3=K$BA,-PQFIJ2A<ED*A $J
PMH&6&G&G:9*IQ?=:TN(;Y+G$SASV]:$G<=]$;PEYY[\NPI:1>WB&3PD[VQ8SV'VB
PWIT,OU]-0SNN:LUGMG7(G.3MGN$(2J!;8LL'WF1&*T[-S4X<@K#[='"_%J66;\AA
P],$5UF8$V,,8E%(K@CNYKC%I;\6J<BWD:>;214+F/5';$D_(J#0$?K0L\C29OXE0
PQO6!W=Q%L.DR8%E^:<YA?"5:C&GW[SS]C0^5\""#T] E]IX I363W$5]CS^&P=TP
PZW'[\S-(178U\L6!%;=5=#)G[""![Y+,*/DQ_:<:1=)%$!(L4P*EL4)A1ZXL%,*[
P/1B?[E/!NN]2RKUHON7$.!ZUXV+&5?>]Z)6D(=E YHTS_SI=Z>-^_*O21%>*V- P
PY[*T1+*P*9PY\<8*B=<5AVUW;I_47Y#=;;GS/R_1.K9_X/B'ZBN>3RE,66R)TFLS
PTX&!?2SZB(L$S*!GIBD^OD-?+H3\>E>5N91E"M\0R4JNW,?KV#,/(:Y^,R-_G\CX
P2!-=2P@O'% 9DP]OK#?OW&B"4GQ*'<;M3QQ 6TJJ].<['$2A%<8Q<L?W+@"J/)-C
P:GQDA3K)ALG^54>/HI2)A!A6,MORG(LLL0! #+[;VZG.$G6!V[\4V[Y'59P35$_0
P\V'?8I;YB L2!+1ZF\X"))7U%IY@Y\X59OHAQ1'U7A[+&,WMJQS%&/Y1%<&<;SN)
P;Z6,@/')N3>K)G F,X$'7^.#)-(G^$AVZY0JH[B<?#PD*N7,1?X,N6LR>L8;Q@X8
PZLG14#[&<Z_*7DP(-GWC;/*-,1J 6I1KQBL^@W,F*?W)<#)%V(R4BX&BFZ..K6#7
PNW/DA>+J:RQU7#5V)ZK#/.0Z#]H 9,-K]ZRU&#X-.D%4EZO,R3P5J"M^#]7#SJ[I
P\>-*9T]]T;EA>N=K95)OE,7T#%M'_5'6*Q(HR]%MVB,72,5\&JL6Y+]=1%.",(;H
PRO:/77=D5)LCUC>R(4?P#'RT&UD*6.7TXT=+DND 1'$^(W<8G&9,39KV:SEA 3?#
P55)SN,7[L91^E9('E8HHNXF@L5W"/-8$Z6,<'2HCT#O*@A78K&"54Q/[L[MQXXV9
PU#E<L!=.29!#IWP!W#TPNMT6G1)6O>.TXPKR,+%P<LI(]JY&8AE6RU:IMP4,ZL/&
P4Y1LN'/3QHFR&6?'Z;H6%;1[HD\/\D1[BEH419&50A>XT $<E<BMH^I["[76_N7]
PL.*H8YYGM"E@.FDH1:@)89_KWED%"J%*]2RX+7Z?S-JH1A^HQ0YKJ'ES/-OCE^+>
PQE"FZF;4ID5(Q;+@:53-3E\">JN]CQ@M@K2_XR$M=3E7M#C>E;E#M8\29JB,*3*U
PS6&Q!BQ]IF6-@H&,[#$;)..@E66)I18.0#6.(EYNG]/KGET=.?WC5 C([(8H;YXQ
PGTLK_^1T+J!5M 5!/( U\%8F]&9*:LI,Y.$E(2 ?/E;'2!?4DXCX"V(?J;VP#AI3
PJ_VF"KRK2(AV[W<6\Q] /68JS9L:-,%<# L)RI5)9J 9'F#[PD8GNI(K/46TW:&U
P;+K]RAGSGTODA\UDMY^>=N'4S3ALU!4RCNV5/2($7QOY[[/Z+D"&E<JKMY>T]#M/
PY1TML&BYH=7OB/$#[ &Z459;T("7"<D(PZK:9@Q$>S5--:\0GP4BPVL:7#MDTHS&
P>#*LO5QE#QNN0Q\8@U*+IOMXV4E%]3 HZDP=0*\0;41"!^+J0@T$!Y@)KH0G2#< 
P$<C[2GC477W_:@D!/,4'^%!LIWF&G7#1AI*)Z<&>=Q*.5#J_BE!,N6F7S+ZJT_"\
P=;KA9ME"/Y&<U8Q3X]8UM?((JU%WHY';;7+U:A8CO^7]Z);:B]2+>#V@=^7W/R<^
P?LQ>]BZ]=I&?=&RA_[(_V%[^BL'?/>C]@3'*/D)R:A*J^0] HX722]]_UAM,,J9K
P="2EMU;#C62DM=!)E[L:7!+I]I\!'7J G&CJ@^_;"ZPJ ;VJ>RG&K,G/9*=#[H#/
PGM;VT2Z$<&F10(BLP-2UQ(=3U_9@9[<D: 4(Y40.'E(X\Y6)_7OW?_I$K[)JZW(\
PJPAIFPKR$K29%4*\5":/HO*K&]?QW^5Z54Y%/@HX=8+H^*,(\Z?,"\-$6"U_VTZV
P>#>E9^C?*KC@B5\A3%8YG8B>U6#;OP:!T\6XFO?1 !1-OI&2@K(3N&+S5>,K9Y.-
PWG?H]@R4U"757+ U0#ZMI'-+'IYZ2[L'E!7/:,?UP[+KI'P5G&X4VC5?BD<Z$-"!
PG6/NN$/!DPV.<5E+.BVWL^L1FI8I7UGUQ4LNA<&&G8$:"NZ$R&I:KUQ6-"D,0UIT
P>M I ]B9#T43R^,GU?]1)V;?M?UG7-,(X.Q9VJ>/G^@;-2-]F ;&10-$MW'9%J.D
PN%J>:A]?M3&'(SAE)D(.;S"BR!=R6EQ0/4D<_A4XB?R&,*H_9V;EH(^9%&>WVEE8
P:%O)#A%#SCF9&HH9Y+-M<,D^>EF@CW)WZ;>&I@5,KL,WRTG7 +0^.'P?(/I9Z+2&
PJHDO=GKN]#AEHK@ 0%"IP&H[#6BVW)#.CC*W<9/X/!92:L&^TY![T6HCE<LDAO4!
PT_1*&;:W^7PN81P8/4SNZFHK:&@VEE!U\&#,,8)$TA%<F;+(_3>VRGO!)9;R>A%5
P#GJO%=,'4I,UUG*7VJ<BJ6E(&KB]2@A&H=3.I2[CZS0RQ%&#U_5W\PSW)LWV/85K
P1?>NS%G,);J#/,*BUCDU^WOQ"IC#+_YNO=!!7NOV-:9:]S"P!M"::P#-L#P+T#SX
P>!TV O/&65]<!<J9"9P+W?T83;^PJ3J5C,7\\['% 2&$;%X)V*M./L\^=Z+YV%VA
PZ+[N)^=7+Q,#6+@HF,!R&<-45W*WN$76/^5@8V=>_2"'P2+$!N?SI\X/7^@Z0IKX
PXQ9W_*Y=2F(BJ'-7=("M/ KH_FG>3_XB%K^F_W?.,B\A1$,FG>]H#)<G1&>UED9?
P>?XQ5VR5Y@C4WSJL4]DA]^2G;DF:2&X@<0F'R5#(_:IIRK=_CTE3N7S&[4PN:]D>
P>I&#J[[7! 1R:8E%9>TZ(X,22+1:=W[F44YS4Y:-Z?SO!GV2V*>K:Q29=FDRIB=9
P6\53[Y:L .LTC$CZQM>R7C>(:6S> '%L0"JQYRF?1\3D*H:][B/PN.AG(W6US/;,
P<%7&538U @SJ/*IC<?154H@>47.>BU?]J])IP,DT!)4K*Y<F70W6VML2GU$Q:7?"
PNA#26!@K_Y ^')D5B'2@^1V XSPS8V>0YTEZE7E]5KUZ;;;_8'*!#92J_"P6T^(R
P?*.S C[%*$RQFSR[)^F)^H2Y0.]O@,P"\I*)14:1]0Y'DQIK9*F726@E2&JQ8A8N
PJJP696V0W'=HBT3DN3HP8G(%=(X.O>3QFM8SV; ))3JX"PW@X4A#ZUP ;.019FV?
P/O>J78G*3Y\9V$Q'+3Y41J,!Q^7W"EPJG(XGO$@_(VWW/!RP"@27WIW96?^'K>(7
PAZL!9OR9'N3.1V-4WX[RQNSD/WBF[4>OCKJG)GWLNVDSF:-ONU9#LJE:_!__(C7>
PS789P8W#FD%F)CYO/E2=>UHD!^Y2>*;5T$R=Z18K]D]]TN;Y8&]/)(\6DV&L2@]T
P&,X;L?1H*S!BF:H-9*QWU-]_K5K//(JQ^3"3<9\(IFF"1.S5G*@)B-51YL&Z$(!8
P/G#-,('!*]IN37DZ!YB8LG)=]W]%/6A.&O^8I4&X<F:>?1@GVQA*IZQ"YO#-K*2B
PM/#,G+XR]YSE-7+C-?I,'O>Z2PJM%"F$B?,ZL\;;KXH0JR ;MT-:@5Y0BIMUMYP%
PD_.#L>GE],9W=?92+X+BQDU.ZR;Z*5 .^V%:.E@.8VJ["9W^I6_] !3YXEC<F^S@
P1"D$(G#HE31N7_-M.XL,94=;(E-R*I\^>6\+3S)H3(GM18AP.[+4SX1!N7I;SF2X
PB3.\<EHSRSMVO^GI+1?:/AY$@BW55(G&>0LYU2\OW1N@18U6EIFJKSF/K>S_\_+G
PG)2DQ6VU1M]S\M.NU@Z_51#B>_I.B7W6<^08*1GH/)AGC[TN[U[&!WC ,0=8YM%U
PM4=0'L6T8Q!4S3:*%_0EH:>=IQ.1,$*,%6A 5-6%KY@ .QOZ>BT>L;1EYS.<W&N[
P8S<#-6DL#"^<W#PP=%(M(--VBE][AF9\@3S&C+HIS,X.O%K%&7_$,5-D4Z]:I0CC
P667BI40A''5H'=17)%^;MTJJ(%>'S"@YY(N;F&+@&%/L43=:NI59/_YM0W"F C_\
P,G*.)[,W8YR?2A*9QPE) Y,@)"131>%QS'X=N6M,1 7ZA![*9Z+[).?4O;#Y]T0J
P24%_Z=A@W/MUR\15_!!LXW./M#IS6D,P;1R.)*D498DE:T6N1*'J+](S[64O;RF5
P@@/1JB)=GQ%Q+(S1K6) 1?H_;K?S\UX<(?G_,BPN*G2S#QU?2J[-&Y+)>%V'5N%L
P>PAO>EI<R)HO]@%9Y.<Q/XS?-](UH(M6\,J@_R"CE)2)L>"82>U9M2=IO'U8[LQT
PTI8'O?T:Y\/IU31"$NDL$4;R[P3#VB'U14;D/#7^YSN\SQH0B^R8,'I_#ZM%@]MM
PJD8$(.Q<#KQXMG"3[&A9VM$U"%%[A0PW)1><1!PPJC)Q"]8/*EO*=(6A!6!7ABQE
P[!=[ASG:.9>Y'OO$S8_'"'YH0\-^-K<6R. KJ@Z';]8XL(MJ5=JU_W,(!:QYCUC>
PCB=AB1/<DJ^9/XM4]7;%P;TEM. /Z36"@FN"34L[Z]\3*"^  O!;:F(!O9S Y#6$
P#VX#V3+5])\'T80J';/2+0NAV4_XJ6TM:"HQVT;FTL"<-92I7DI,L^KDQCY]QU!&
PPPT##W'8M)'@<J8:)Z9CI;VM'#,ALJ)F]Y??%X./TKBTARBQ]+43R9"<$@Z I1/U
P).'3,]!>P2M/X':E/9U"H,1X.F7=FCWMUEF3\(^692R9HDET@35Z6K&'&\H9-9(>
PAZ(NBPUTX$&JXB20Y$^H;)K=W"S(4@9.C6MM_D $KHK,0O<(2><,XI[@V!#H@#HU
P@D^2.VTK%2V7C*@R8DKJ0LM/43+Y455HFO=EGDCLL3N!.!@0YK\H6J-;4>F".7=_
PR,M;WVN7;V#?<7QV+,'ZPR\)BGG_JZ*UBZCQC)-D)"'!P<O45+4(CVZ/E4.!A-V-
PIZH_LV935T*QP!#9@^.6=+KHH'D3-4)<HN4,$X137YR-L5!V?8X-2QFCE@O]*#EU
PNX_^B^4V)H J3KK$#+F#503002VQN4S#%%OX9HY04;"^;]S RN.*%[W"1HFNZ$\)
P@(5[H7VB$W([F4W?*'V5,28PXR!.YRC)6FSL=T(*!)DJ3Y)->T%'!._DMMM(XT31
P@^N";9]I4"U?2,# Q+O6:@JD0+.4^ZGO]*L,HZ,BHV#MIU-(^E$PI]5;Y*]1&T#;
P2]U7(_Q)#-V96)N.4)OWD/RHZ[QPW%F"$9_Z^9>[X/_AS)F[TB.(NOBA?N1G7K$ 
PO^RFJ_O,>K2;_OGCB72D0[+><ANI)I,U4AQD(QLF57:(D%KKSS4SO*-VZBQV2<\_
P1UI,/O?MM9FLRZ.*'C9%X<=E+!F4/?UP=").5\_K)^9MAY,OH E(, M%^J\-]3YP
PRX>;FPXR]F2>CL6I/-*^48=,K 1#NA%+U()(G(9'0?9'0C;)-20]'N%EIH9HSWD&
PV 6%[F.3&H1,$KJM$C$Q+EO;\"LU3#9S4>)O= URZXP_&N.%$QT8&\[PLE<#?V^%
P+]5%XZ!-YZ#&@*1>>A[9G;C1ET6 ?XG/RNH%+2?)N@XAT]^$&Y=7;Z#)4[&52DLK
P%-CCXNJXGD?D?,=^Z#G>A3XH6:NT6)-JA#1LO7,L,&$'OR?+VV%+C=55ME^[G&TD
PA=0L[9 TK_OQV'JG;V5=);N!92GXE:I >)199EU.JJBLXA["[?UNZJ*'?COQ_4R;
P_BPB"OX"GR:A%^:\%R#M=/BUKRS\$DB27;=%<VC4:GI:PN?0]Y^@R=\06_Z%,&KD
P954LM2T5V;9%5%N/T08P+TZ60%\0T,E^'_37D^ROM:!-?U17</FU8WS_+GY2R29#
PQ0YSZ;ZKV%I@DG;@O:9Z< )DN9LL^P7F?(&.P+G<.<4<(CH6S ?*? 4L*_E7BBHP
P%N(-M!315X%76#D4#"=YE=#_CX$$E4\4LG?G0IQ#NV[DJ/:\UJ?344<F4YXN^\B1
P@;,*4&C$IOS[A+7BU9](=?"L40?8DMM]]EXQ'O^?/S,-I06"I]FUX@AI:S?\&B@0
P6"'+CLC!G@I%W5NI'&@P?\-0>)C?;$=?#J/W8QD ([S>$*-!HM? [@N7NYF#_6!,
P,:DX0W0L"H4?1<%5!%5OGKR0Q:Z;2:/.6O\G^FM0F6-D;@^C3ZN-^8<\/:17](.!
P8>M'8OQQ@+O!+"\5$3PL<O#FV<O#B19S"/*P+@X[A:TK];=0(OZ%CVI3EU5T)!EP
P7U9HU2-]_P/;J.RQ&FHD<S8"N:D=+3"<C<X[B=VGIS!]QYQ@:PA<9_!'MZ#XR_XM
P21B[T_7M7S:65D ''-<>K6@G3CNS*VY]4YOF9R7+8AAS:!<&F?:W%-.1S8QN7,.)
P/^;1+K/UTU[\#V6<W\C)@ X\%A:4^X\1F 'AN%Z7*^\U]"@:IQ?I&7E]Q;K:FH0^
P4XB(X\;3>R/LE>[(ZH&8W[3I?2[\?S70/PWD;:KJ89;.>PW*=S&6Z.GUI&P'H1!D
P@FO=FD!2Z#\RH74@79!#6^]!EY5ND)EOG,;+&5J36PE1M]Y!'*E&0X@8L1,;&:)<
P>,:SX$;58C$V\_PA&P"H ZCE(=*9;P*0+#.@.Y4])F[C*&8&'SC0L:38-I91 /$=
P*U%Y6O5:PES<OBJR%M/YEC>^R/W=^V8_C(C@,X%TNBW'A68792>7I\7/8..-Y W*
P$S_1D"+V]F6?FP+SKC8=<-]S#FIK:O1:-/,067#W-.1YK<']1CQ/3$CC]0%E.\+U
P(IA4S3/+!62@1TA<ML*Q(T)2!@K=6>4TVX""(\K;N;HUL.U'^XX#H=\KIC6 Y7C1
PA$7@<*Z5OAU/J4=%KS/@CZA+:9!5]VDA&.)F8#"2Q\DLFYH[/U]^$;9&DL?25?"C
PZCH/]XI.L45..?8S>9OPC2W6TD#+-M\ A:$@G0@6&FL=K#1L7L=#M4;@=B+9//6P
P_6'!/F)KV*%\/LQ:'!9J?]SX@CHUCEZJ@"BDU#_NMI9:!!4D0[.443S..NW'H(_X
P0 5E*%/Y8JC:(V<@?=8'*$1RS-[JG_?\SI_F\@:_FFT$SAQX!-W0@W(TA\:%]4VX
P:=I *L7?C:F YK+'K/B9>[,;Y;Y="<?\/P#UO+,KSILB?V;@6Q/QE_Z<<-52?D_>
P?8,A-1S]U<1I&61E[S?+?FXS9[&D!>BM5;ME3)RDEY!"_"TDJ;-Y=A\L.UB9;#;Q
P<I91EI'OK)Z(<LPZJ\V?9)VG@ ST!$.E&M)1N"QP<L^J6VTH\R=;]83RDO;_$P"C
PVXFS+G-E*-7"QRT9-VQEIZ*"F+X?K/+U54I=&K+C28E/*0Y:G,RE&%0FB9FL6(0@
PKJ,W^#_MW$P=I?XTP)AR4^,)@A+SSI9HK<WP<447QT57VGP]BNB0ZOH DUI1JTY*
P9KS;X*BYVD4*+P[1 M.V_D](ULU:8PZDDH30Y_7C^ 9T5PV@-%E'!_E\C6 % UP#
POJG]'[TZSJA"(EH#MN96&;W2C![#Q:_)'W?D*#3UU$>Q%%R0\>CVCM63L8:THV_D
P7E44]S(IBK*9]3ZOE+B(*UZ$8(E'02_L_<"9JXM->B?'3"3 @P&&L]#]6<[Z7+7D
P<%?GYEJ"0'#N1N&=%LPW.?*K:"AC)-\S+%NDW2%87N;B\'V0Y0'6N +Q4X;AZ+.5
P]8PL"$UX%V7XJ,"-H^77< !_!%==CN8<E],=#JN48C?$BV'V?%7D,UK1!.-[F.E<
PNJ )E7^VUXW&'9:19 !0B0\B6>U;,8/Y.WO8STRK,RM5W%(+4>NRO8=R-B!CM# 9
PZB)&?["OIM[])<D3.(^<^%(:6\6%"&)'"0+W'3<DC56/>R_CBXPL9%]IAEM 2:PS
PJ  D* 92[I"-K:.?A[A2B6N)A#R.'JIR9I_N I'('&;ZP[0],=JK#F5SO/N0Y(V(
P_=I[*R6H=P$-B_6V"HZ&=.Q,V+&8J ?7Q-9>X8+L&R1^:4D<;=_,W>BA5_A8HA1H
P:NOAZB!UFZ$-UXNBEX5*M]I^;?"\RW@2PP#?L_"-=U9:=A6DI :2U:I"NON=O/JR
PZ804U>;VM=KXXY3+)ISN(<D5SCFXN]^+0O_LDOP7["[3IR>>8QSD\+PA$=*,2+BT
PQ+$RVPH+ )F@,.7>).OI<DX$FDR2H-H8&MPQ>:DO Z^<)GO\+ .4+%TVJ$0>T_FH
P7;&HP[V[TSI-0GK$8 C@15#09/+!#6*D]MJ-2S@I ,6^]1N&N/P-!>I!T2:O_\AL
P""CCXH+T?,6T:=VY$/)/2O%9=NJ L4+HL =/3O+_"<M!#@?$$8C(?2 B=+&' -"9
P^+YV<;DV4;_16I'0),RQ>91H2B^VT$TAH/1<6R!D=*T2%_]1+6P5"C(O<FOYV;-K
PCVX=T7_;\?0C\0?C7_^O*D.39Q<I'O*L[DS!'N"8/YE.CJ?$A\(&^T(5Y)435'<N
P5W2  T<N2?BL7:O7Y?"4/O"]_/\6+IXVF4#8"9 W<R?RNJZ3$;F\:1^.2=XXLV:\
P 9<(B.?Z$1*=6M[@-5PB*GWH'< 4>7[UL!AH<GD.E*B 0F$)?=^<\Y6((0U1Z:29
P8?]EFKH5I9^VA^8UH]]&%G9LPR>G2(LF\E?XU\3",2P70S9,0R<BD^&QJ,[:2H;'
P* =S))4K?GTX.2A*M:9G-Y-U=4?-,UMUYC-;N Z!]U11\K!K-T<,EU(.5R.)F#VK
P:GJ_"BOC*:#H8O7F_4+3,9LP:[EN7,U6/%WH8U8'@V))7]!G&SF=3SC_9BP8R2SN
PC.ZK*BC$O.US,[:,YF&TB<@!P49[[8^O(4*T>+\HB1%?OGFN WG^[QJ@&HN,\;EC
P"_E531CL"$C[14']CQ$!C 6V*C?%X=#ZF0_>4U9&KGBDMZ_E!KH7?-V=U94/ /N#
PN4E6 R*IOUGX<+:V="E'01<J+B0=\<F*$0RC>[-A4+HVBX\V%>VW;,U69<)4\:LM
PGB1NQRV<<4 X/(<PBX^]0,UP*65&L+_&Q3C?Z=YI/)%4\'-T'_A08J:S)):Y%YWQ
PHB(LPCIW!_70MBK ^_W>16@LI[<CBN,]\$<#_)A2A[ 'K7;F/1L>!_BWNA319-4:
P=9]NK):OJUH:,(STP!63,U3Z#26ON+<>$2H4V_ R;OU<@^:2![T_]G">"2?M*G.8
POF$Y4?H)8?'R %*2%^"799M%2,G!OSXXVLJ\56>+XI*VQ/4+) IS[90'V-.?Z@4O
P^D;P=2:R"YY-.I 0N\DWK^)/#@=AW+^UK1(OTJEI&V7C%7(C $!>+L;YFRD(HSR"
P-D5>HAV9Z:E!H06G^ABQO^&^M&-J9FSI#2L%2')48VA5)WK U#O^B4_%@PMC_1DU
P;L_V3WX%C5K_C/$]$<)@"10?.J)!2;V?A8A,-"]8E>FIRE(&/M,LT$]U8D:5C'%O
PO9"9M^)!K5<BC(+/@17*(\Y'OT3@D0_ZB,*43+%P,!;*)"-\:[TI.57S%^*<NQ.H
P"$5HY[=C$ =B8\4AQ1GNV3WJ<FZQ_VNOG#['%E]Q\UDT@,,=4<1N_RY7GH<L.NKP
P8SIX"RP?U'9^80LW?,VQ:TK!R.;#G1_I32V_NFZ"-Z1F^Q4'P$?$:YI+4)Z@R)&[
P_BP'<7SC*W@, *K5H& :ETEG]CH*4M9#^\"(Q<5T@1'VRI8N6O/0T%!1F&>][:'J
PLFEN5NY *&V '$-L%$; [W*O44]QW^ 3UC2;P.]UINV%II:*&8KL=F>J[A$XH%2B
P$!+#0C.B3*+;!(>E%8C8HO>H$P3?>'YC<<"<F[O9HF]C+N#;^K',^QDV.#'<SU1I
PCK9KX7^X@+RN$2=[4U_J%AA1'>'-M_!BG+J]'"B4+&Y@D$6.$P.ZR<A&KQ=156=E
P6;<$]N./!K>(;IL[LBD9(W;+\I.NXNS3#O3S7?'>&8ETG_D3!P)I:;[9.,IK,80Z
P:@ C:@K45<<Y$8D?$8/%0OZY4N)/K3 *.:.*MXTY8<*<"4T_6-#Z2Q#1XNGTN\]2
P4U2*<OY^":_XZ64T.&6+=1AA_M<:-TW:N13:G[>7M8O$XWTM#H"]:8E* B%G==)X
P "A]A&H;RPBS.@0*=4,+XFQRC8++]L8U6B/TH!D:*Q7O33%TL!R4.)/$IA((*J-0
PNMBVV+_L*I9X85PKX(AGS9L3=[TJJNCD9UA 'U$;FM"MU1N*ZDUW- /1^(W9Z4!C
PKD,?V5>$@2J.2Y-%N)*UM@+":9?I2J_U'F!S&=H\A>=46-4)^>"@0/ZHEMMU@?!X
PMQCC,2@0[\->XQIAR7L?M%-5CZ3[;@+"4IDUC!A<-YB6":_3])/_>F$&98'O=\[(
P\SFOYW4GLP"58,'3@.PQ'@8TQ/X_$6C6OV'#KI)@HUX%NW98G%EIS W&OEEL1]+@
P@7LCF2[(Z(9PH48= ZO"@N.502><!G]&KA/%*E!M)T88X-,"I0N'MDJ-B2UAYC:+
P&LMT;3023)2M>48C)Z/)B4P[ ^DF20-@$)MK[Q3(\+7@$D&OMQ^#K5&K:&WUB4_F
PZ[Y5[?'12V=5 L7T)C<*0M6CM[><(*C]%KK57Q[[8\=^^T"!THCS4QS<!L<US)[;
P55L6;!J^6FJC5V73QU&XU"W^2+,9.*BGR%.3-3]8Z\P$_,07KW?JJ)AF9>HR0'K[
PZ=T4 JBVCR8>RO9"-9)F:ME4$_ X4/ACQVMY_1[1K.8$C6M.Q?)=C/=^H['"W?E5
P4!,[49PT/_3" \(?LNX$]IYF#N"/*'K[#4ELR47+]QF<>K=]#>,B)W+0%Q@NW"=:
PL9>M"6$3$[9]$&]O?\7HEBD3:%CJ/.A,2TZF/TW,![EL2EV[L)/WOM^^ FGREQZI
P?&K/0%\N,Y2=3%?/1-MQ4N7,P5AG+D#MMTZVXVTX 3LT<(QH;J?;<6W[<0C#D\Q[
P[PE0Q]!3@UMU#MBV,D)- Q_R#QO*X1//4P)6NNPEDHQG"KT+M<@@P5?R;[C3M5%2
P0)!0>PSB-O>LXLB8TI_W$HJBJDL8CVN.2O?V%-T1GBNQ_LDG+* [0_S,B:,BH8;[
P?HA,D)P6M(FGJ5YN%0J5,^T",#>$F@G#YLZW/R$S5*SCTBO087+ Z'<1E4E]90=I
P-CK+(T]?FB9C4S,F2])F0Y=8%CK9#-EJ>BNPY 8T\]97DHQI\1/B3CZ,O2/#NC#Z
P4 2*[0_/]*,OQ"A.'57@4U?\A<CH9_$3 NAJW(V&T!>RLZ"2('VB3&YEI ,["TYK
PX?.Z!':$[*32$6.0KG[*+#2D_5HD]Q.S'+8@.VD<I4_X1D6I3=S$)0>E)0&V;BD1
P@BZ_$)F!5[KD+H&U[@,7L:Y<W%>$PG9>R#F#B]C40]E7_P+8C,5Z00XII)B7"BE^
PB&6 #\H\5T1(&HR^VAOTZ:78^H<G.JQ6*TY'.A]KO$!(%7OG8DY/KX/%3JRN8^"#
P OAXH/M#T JS $)P'.H/!=;/^67"3,I2&[BJINGIN8EFL0F6'1JM!:A+,I\JF3*<
P\8_KWS90ZAD1.!^.PA1&H0&P'QVE%/;ZKY++"1K<'#H(I%?^DJYT8SZ:C$*Z=/A-
PUYTJ7'=]+28"+]'K\IBT K<ZIJ>*N=YORS!?Y^8AJ"8A7.UDF.F^"# 3:/)?GUA?
P0(@P0K ,Y9>/L#X,?;!*^_1 [-S)N1+)9&OK;II&.)N"+>0S^,$)G[F?@\?I5F2:
P<^+*1;?H1UI<C);J:I4J+9W\Y"QOU*O/,$L]H,J50>,\@[R8(%K"M"2NJW$+%R2Z
P7#'-MZ3Y3=D1N:DGMH%KZ*T7#3D9@PG_.JYZ"Z:@K(,6D*#]Q (S(5K'GH%23EWC
P-H?K"@]X">;LUN0SET-4AYNNRAQZ$$#NI'\+UT/GN\YO.]J+P[[7*7%ZUMY2>KSI
P/6L9@?/_0Z;WP( S__@S7Z/B#"&SX=B3#!FI<X&J\+W8_ERBDQ3(J30M$[N5PH.B
P7;ARF(W.5Q"H%7[PF+$<^^E^(N!8AY>[((O6+-,-D[,W+LW77KI9>.D7I3=LH.-2
P^/[,T^I46"+OO@!DM>Z4AHI KME$TC^" T-//'AW]C%GFW4E/F>S::@(M^R4;J/5
P"QEV9=,%RDS,X.W;MG6R555/7-&SN->=\2;>.4G1NJOY0;UKIO<];G\D9'BHX6Y*
P1'_F+T085Z3>>Z^<I8)F,RF(=/#$$#AZ&.F[WRB9-KZ1&0!4:B"Y>X%5M^T(#G6H
P]0=1:WEU-E5ZY9Z)0EAX6L[=:RS?M>1QR9"8NK#6F&PF;2'Q'!E'5A[@6O^CXO_K
P8K>JE+2/3W>UH,9\O6!_?C$QHO8FC">Z&#>6]G?>VN. :"JLOP2JN)]X //G.>2=
PHH)^RB#$K'J/F4T;K^L:&_IFP(@)]DE:[+:*4 XZ(Q'G!6ER01J5FNTRI14M#4H(
P[7.BD)\.,]ZUT](B4_Z +-7LQ6#BO.\)D[7XW41P73(5'W&EI>XX*DO^7(9LO]"@
P-HO-I"]6(&+#ML>+.YN=QCD:9J,H_=<<^B+&>R[ABCJX#6),@&_#RFN[S\LZ>G7R
P)[+9<8D:' =#F,GBHQIM8XBNV6LZ(%\64U*C*&K1R*HFQ+OHUUU*S-8QX9_;[6Q%
P9:K?1^_/+=YIKW%QG#\_*7BUWQNBLPHX0[?G'&I*J,)4@0YG_? >>J=CV5.=L]?_
P>O2P]X\"E.TAU^/NO;C&2L0:;P_L5\H**ODRM"<KSMUJ\*T.G)W\Z7>-;I<;$G4/
PQ#JN]'3  J7-S-O#URG-DU0M5ONFL*&<DU?1%4[EX:K^$VKN_ BAN9 FWV*9KE;X
PK@ %L_8T"LK[W(.%?U-\I_#UY07WN#8ZGO96&V^X$]2 5:!CFQ6KI=!>A,T0J]P6
P<OJ3'@'[M2)*#+E28I?,=U6LK Y%Q[P4_0?_;U@"M!&MN=2==.L?0P+VV07_7YHM
P_LN-L$PN/@FIDJ6VG(T'!)P>@$*:MG3UWJ[.SL439.PA>D_NQ9QTG#CKKO_<]-G@
P\I?CIVP6K,HZGDR.33\? T1(6[_M-@JB_.D7-C/Q:)7[MMP-5<D0C^U:2$=0%C@N
PK;TO["K-+"=X,8841W$ERV:4,B25=-G28\AC&CRGIK0F]!78":QIR,F [$LG$:*<
PQ,">O[ /(D^X8-5/B(8*',1@?<ZG+EQJCM>E\6_Z-7N1='A0Y3?HDJANMO%$2\B?
PI.$M'PCE@KV"RRB[_77%&9)?%QBB(([*3/Y8.AMWO\7#F) .]GQ\?=Y<6/>[=DO!
PV32NP!/&Q9S!'*&G$B8E; I(X:AN>(;<P2!!!#H;>Y>?>5EVC@O[#Y&<AL1R]KR:
PT+W7?-,T DGLLQBC6019KL(OA]'P1M+?VW2?MYUE\(I8K=EM/.@/[ZPJ\.,9W]:5
PQ$!(KK(9DG?+4#7I9B+<(V#---S\OU=!1#4V5C#TF6DY)7GX(+ 9;1CRZ9A/>AZE
P/P7_8>_W^M5*>[I1IZ>.%ZD._SJ&&FI3L*?6*/%\T3H7&U:\&ST,JTMGQ!>*UTUY
PIDDEPX),MI61&Y.T#'O,MM#;^(.[,8/D>@FN>:N)U?IM>\'05*W<\U;E+B[>%MZI
P*^M(EY^6UU]#RL">SB@8SO'NI/]>N=,J["'ZEKL.L9QTF(*RF'P0>7T)0G_5J?)Z
P^&J4V84E("R6^Y<#FU)9#<$OVAG]X&/J4X.1)YGB5$H 8T6>AF<[0#N"/,"NS]YS
P=IV08CN _CD$X&PZRV#D;&Q,$)R@%^^IVPM7M-A?C2UAGGQ_W0&*9W^?:L'M3+U4
P/-;KTB*UF0@4^VAO4_DP/T$R2Q+HE]B]1\X<95 Y6.O*8N,Z8?E[X#1<:L7@R;@Y
PMT>RG2-@5S8'J[UJW,'4%#P!R^E%9#?M46S^F= #TBBIJ89@?UY.*R/#,SK '(.6
PG+DU579N8O[#B.E"APIJ$8%^C87V-S3X/7,BCHDXLJOGS%-A^1'DAMLG-_@O%OVX
P,FJ/':,C!+Z]CF[8&T+T<J>O]/^M?PNDH5'F.J>(-@D\YV$F(4>EZR7W#I$KO,*6
PF<^QT<@:;+M6?5O8;Y@0V(=/7&H<(\S3DL6QS U^Y54)#/"%T2>H\X&I4)"V6QZ0
P!38KHE=SR5I*C2FR;M''5GH2'8V)%-\ <+3TTM,5.'X0-H;Q]0XSU/CH_2C&%WZG
PU@E*TJAGC<!=9$S+YEI+8W:MW^'I.AK7P):I96D")'L&I=4SRG+HGEH;&IT\S,.T
POE.LS#G_XE5!]I,6P\0<2F#--'@>QA>L \=& MHL:AF4BD#?:WS]B4)JB/O\N@NP
P2E7  [D'Y$1-Z?4W#JVPQ8]'E:FKY3V@+V*#^(V$6W2/@EBTAP#5@_9;:!M,9_!*
P$2@3*0%&^6'JAD52,J+2 IQ%+C&-PR1PZ+]ZV@@N,YXL!'38CF8!C*LAT ZZDC?V
P!--;' %R$JGKV$S"O!_U5Z53I2T Z+'5\AZ7=Y7I*0ML<[W]>"7VTA*CR4VL&Y"O
P<)H51BHWREAS#T%'LPM^:UUT8C7I\J*M1+;:Y"8[W]FO%0].?DI&5->IZP9#OC<.
PBI53$9WSY-D $2J4MUA=$$9DDCJQ]DADH7Z&#A8,";084C>ZF8.)&&G3T[Z<).OE
P/+:*#8IT5QZ*9 ("BCCBT>+M&Y5_4=B3J5&2-ZKCU1G=J$77':U+\MH@Y[E,=5,=
P;40/DXA\BG-.N\?;T5K.4)0I]_TTNQ.3W@0SWL/4BR6>3Z;8J2'>&8!AUBH[JU_H
P/KE.N,Q5*_M4A0FIB&'$V[FUQMVYMG,Q/"]4PLH0*/.=ERZ P,C0^2FF'#(Q.07L
PK1,1K/!?VR74"C"-%OV_W70$*W 5,@$<S75\:Q_FC[S%T-:5R/"[1O^D:"YW/D"-
P^'>ZL#CQ-8H"E<?&G\< 0+T_(59G^C3P7D,]+.^C[PV(S-8^[TX+R"K6F@(]^_"G
P-<1<^%RE"7N8%/8JO,:!6_V)X:U[%:#OR_9=SKF P\R-DA>"?6BHI(S3&OF-!V^K
P&Z_*';E@VRW"$(\A= Z[>?K"=XGCJ,W]*P5J34\20OH^$')T]QAE^!>:G/U%ID))
P?NU*V$_[9VIA7EK\U_)&E/W6/,-B*?"M"T1EJ$W6:X4OBAB.L'G=4=$/[J Z&*&1
PWO82DGK,L+[-*/SL:%UH)HFU;:Q] _NJSY./:4//0O_MSSP:ROI" H-]Y'1LR2!W
P[[1]TL_"#4J_:"S=C4)5?LRUGX7$ZV5S[N^'("*.8']2";P.;Y;54-XRO7=>RS>W
P HWRJ8-J.M>797U;*!2-Q%&:4M]FZ;>-ITY5:R[H4GO% @_.^@VZY+O/#^0]O;(A
PB_.J$+=S0$OL<KM1.$WE(D D4/YL,:O^VPAJO#)ETI(WPS&7*;[Y@E]W.AK6&KED
PQTIIHS(V?:!1V- ! " [GR7 5E17O6!\.?,$IJ1);-R=U.'_77N N]KYED,-#]W&
PW2"^2&%=N#.!DZ.Y05-=4A0>%TW;SPNJL&Q^ YT9_ MSIM910&F& (]'1!#Y]PAU
P4[ X&S9R_!$&'??APJJ*88@2HNK<\*VJO0P/Q])%P ;&(!GZ3\%O5,3(QRATUT3J
P:\*47],0W]<P0@G8C[;35<&9+,727NJG[Y):T@_6 8!,]O<@P9LTP^SV,@$J"$<!
PY>^ E-BQ04HSPEG2B4V==ZZY$-3>8CT6FJ,[^FPB#(KIG'#X3>^@X*MWMMN%1-,;
P^AS?3/T!E,V)*F]CJW[,Y2V).E5!>^/%>QNX0:L.0;7P* 5P7J&4 J[XRO4XNR</
P(2VJ[V4Q&"\($U,6)(_-2_=5Y!*EP.R%PPY=D?U3WZDBB/7YAJB[1 J Q?#'=>(.
P+J^:-.'MYE!(D SDSG[EX&KY%-!Z9;9]!B@(9!(&@%O-'EBS='\CRJ39U/LDUY\?
P&AXU6GXCH,+3%.E<LF" >V(I=^2H\QOG5-BR79U'YQP6-'*TCQ[B:2O)#[BL9$D!
PH80Z.)YS!PEQDV8C/HIH^V]6G945YQ4ZR)I2()-91#W/A%:D"I=E1?&&X#[Y>!FH
P(N";;<?LSR;R>8P!S/82P;I>.SI_=#W.M>JK!*Y1[P-)^)"I1$8AUK]%^9'V@=A?
PHV[X4M0:EWOW#3(R;?5RF8?+]U$<*LI_27@2#,EX>Q_G!U!<_0TQ,C2;=E<$HNX'
P#FL"$#(Z ;FDBV&[1W^#+0Y&3\T4K=R=";IGA9IT[SX5W0"5Z%1 '!>',*J\U>UN
P[CC0:7^:>94$4#UO3[+>/^T>7FR5_V)_#UW-B\XJE5(4G-QN^F>*//9C54R#+G8)
PT/90M"/(!Z0KI:+>]AR_Y!X2ORIC4I7W<,9#O8>N0WY4%^:TXN)=_J[@N9G^\G>'
PZJ#Y$[Y']USN+ZCQ]:XV*8CGD)HUN-VFX%LF-;.N,/CE )1*=@PM1/L!07G<N(S8
PP?FC!YGVDZNBE]="HV@>8VM[YPFVV"JP3>RF2Q_%E)_9NP'4(2K?/+M+S6V+8QP(
PNM&%6T'HE5[A0;J011O"92O==:B-M8EG&LHOY[="%5UJ/G.<!S<OIXO)OCUD"L]?
P,GZDW#Q8*_+JDAT#A$H43*8QYR?;PN9!WDN)[^9UQ6,WU#GTCM,V;UZF4<:9E(W\
P*6&K.EIJ] *+*/QM\O&F\'*_!MRFM3@L 8_Y!B3D)?*=KTQ;>1WET 5K>*/ST]%G
PUWE6W!CLI:TK>A5%J6=V@H=8V95N.:WY-X 3E,P/I2(+#!_A;*ZG1><>BM]>J73_
PP=M=W8JR"9HXE*J6Q:DU'J'4\ZCB=G&U#AG!SR^2C0CF4YUG&]8AB14'%Q.+,)EL
P?A%RIX!4 N8NL2)FIT..6)^X=(="1 $&@;+&D]E<:0%>4W(!<3/_>@)8G@YRYY1V
P=0A@QM.$'(4ZA67A,@0'O<N% ;WK,!#\L _P -@N^92\X^&0X**#-^9,78#6B>J=
P#RJ#XI$'EWV+!ZP8>&]13%1KG*0QA3<S$>+8TYF7V:*,89 ."\/YXYCUV)8PAV:V
P,(")D<+F)X-EYARQ&I6<F#7J RW^J+W@,?99'FL$]3(D(SVP('3A7WE_<-'^$T'-
P!OX]YUDW/Z$@ME5^4CGOXX$Y+JCB62O2R(5I#.1=&4J>7#=JL,J"?!9+SJH_6_W#
P4IZ]W?U-#B  '*(^#9R7P(X1&"\K><N<PYG$H!778Y=IGN$IE?C7INOY":?8G8W<
P007T+NWH[<Q*5X$J^X?D4B#5A:&]\^95:QHD9D4H]93$""+&OR3&DXG51ATEASA_
P;FE3RFTN>%A:!OG'!DBPCO[]'F-C^''!V>CJZ"";C+_EBQF=U_U)"'0V)*: :&?*
P"@<;!-\S'!_'MTYM\G4B&HAW<:12_H[Z8[E%(4%]POGY8XQGN1:<(0%$L+TBH%4'
P?7EFWT#W=M3D"(<=.F[^BPZN''S.*5C>I-32BL:1A165-?KT]SRR,U:Y!M5,=/BG
P='FFUR7V 5>X(=!,&9K&04K"T0$0]]U;L/*"II)X!%X>*(W)_TZ9//2Q&6EX3345
P)K'4ET8LH$OI?<\DU!#EU?ZR-@<0X"-WP;WT.G')NFU,G85)$G % 0"W-KX49UEV
PB%?9E74$Y($&O>F LKS^X,S2?+LOI@EG/#Z91Q2_G+W6L_%Q/,.^0[W\8VY-1>@#
P_AXD.J2[):XS\J2SI>8,P(*<>ZQU/'OYI#F'SY8X&UXDK+;LJ.&MWO8))"6, *48
PQW-T?;.+'V!MV/7?RZ2: \7+*#':U(<BY:0!C$B[MFZ>K7YSLI,0V24[FW=DYD$R
P'['-^1"@(0=VN@:;O,V!79^/I#27@ZFQFN6@I"8JTGQ,9U+1N+8V<HJR2'QI=$G7
P]].RF9.:9CXB)IUAJEWP, [? 'ZF;33SL*+*"QM/D$!<9DD;(AFZ50H/Y#ZA,%?H
PM)"V]!;](UIJCGG/+T]M,$3[YYPJ5F,<^O^)C+#+:_PI! V=C&79#>4:.TW:$.L@
P RP D6OTR6VMSAT_=:Y',ZB*8P4!9@IA%VB0*"K;F<_YDE.AL")Q"C$@;&&\\A"=
PAZVNKWZG'=+U70P#S"3X0D!6EYC":26CU&G[8 \J*;S50!R:==9O#!^L:HG^-SJ%
P=ZS\5?:!;US/BMS %?%W4(XCDD0^$57-&2%CB)W/5O-M@W?U>L-C-4/M?=/MG\UC
PM(*%A3]]/1&_'<#5 M[$ NK)%H7+;3ACF':<\+ SQ:BPV\QVJWX.[W[($[/=H.[_
P'X J"3S3TXVPLG=HD>V)2'^'-RDI3[4BU'O(VH2@<!\19HIZ<7&$(CXZ!RDRJ8+4
PX@>M4V(LU#0W 1_H\,A[)(8\^I6Y(SW*CEEH] TI:U(==8+YKOFVQ585ZLY]FF4K
PWJ%0>Z!QIQ*]@@=O$JQ3#FVHNNEFLZTWYW+I^:-40S(;*O<MW*N1]2;"*T)65/:-
P8N#<& -2TE/8BIY0==]6?TI X[YNUHKH24V[BVE73&(V\UN$_,R#'/>"_#1\+&JG
P7E\=Y&(E;;:?U&\M@@$<WGH)I]W9FYP\HU'4,=1*UJ@=AU:@!Z5&A@\LT*8)^JEE
PD#MO<L9OS)"%B_DRV*\?^) _'>+,W6RWOG_J \5ART]R#! <DC9S<=+=B_4C[O0V
P;'Q$5G^\.K+8*[Q3-\*T1)(N2ESPAT*J8R=0DSMW,3/F=S)1#L#=CZ9('AJJHBQ5
P0F5D!2-3#'AHKU6+&U=W3+&/I[BC_\P#9#[K?U-RH7A.S1@=J3A)<COM5LYI&H.Z
PR&7EP3QNM._UCDD:Y-L6ZMD>35@MVS(ZW;/@<* _>97E[C1,UAE6:?)']^'Q04.8
P^&W3K#&>[C\8P>&FX7 _QI<:IKW-IIDV)J2V?;<#:\GNE8;/T-/%92DK@<1'S#VV
PYWM-CLG +KZUYZ'3Y7T&;7" YEX5U$M5CG4"PPT246TLF7;)/A\/+K^_>-1@0Q**
P3HRU2)!*OW L!X?Y1+25?/O""8@ MGZ%UNMZAAS@S\#.0FJ0_WD2V3&,.R-Z\7&7
PRRQT=:^DO34F/99#C0[IG8)1L*48$K%?SY\')?XAJI)49.9Y[9_'N >OP+5A,Q5@
P@&!W1*,LT;0 ("_;%\=2N_@7+\M>[^%SF!@>L"7)#+CORZ):;*WEZ<7L(Z?YHKZ&
PD+\WALZ-+'+NHR9K/J)^#XF'N;\ZV-KU:H,T O-@IUW Z*Z;F0]3RTL_].I7N#D'
PJ+C+S)[=]Y_;#+R>)\@4V"6U;W!J!UNEPNJ6/\I((I854RL5C1W"#+JF+TEZ:DKU
PV9_;_E(>ZNO?347E+37M5A-^9YZ<I#-K="'PAZW"N;%EUVD5(_%#3+)H_H!7CT&P
P#^16L:0ULX?VC>3ZJK5)VLEULQ&CX4QX^7_@E;B%CS>DG:N<V>B"]'08!9_J5N1E
P:7*RJ,G6MOC]^%3A0\"8N;",$B7S5]8-\&">R>.R_!.S !#"69-QX5*K,5I4X!#?
P\=OUB!G:__3=H5PJ7ZP>;A)RX;>HM^#?UUXJ'JZ4)5?U+PA1XP0:&PDN<7_@DK@X
PA2;,(0[IUA9Z,YBZ?T&\@Z06L>/DD4H.>G$L?_@-T2V7'HK!T3,;@TUTJ6YLJBF4
P>.I&A (F?I^!*7+-7=L]KQC#)_D%<VJ7-&H[Y)75^LZ5^<J!TGU5<VN<*$WE01=/
P &9+/81X# R ]*B)(FEL.&QVF5M#YQ8U)I+/UX_M[[Z$Z /;ZH>W4"T+]?15FGDE
PMNJ:B"#4%Y8KG]WBF7%#9\Y&Y'\:5'F=!\&X91R/,$S8Z8@H>7KY]GN#7)(MA\)4
P$$M9%^00KB-\-2;]G>144,V=US4(X#^J/SBT8I2TY#NL[QL22$0N"B+-2J(!FSDX
PT*>IH'Z_N7GV10KWB)JP[J"LG"8GO L;"5^2HD8DAK?(G(]H)0=:"98OU1?[CM,C
PHE[?[S<FF(%A28;0NI.W*;"8V(\KQ#02P\<."!.X*/?9=!5<3$D#NF.1+1#LK/BX
PVP*Q]\HTP* PODT6X.E4U78G(W]"RRZ>1MZ3@1,CW.,B,MWMD47VQO4)R=!4R?7:
P4B6]93OF<0L8W3&EM#(G8T]>$P*69ZHQFZNB*J1P@Z@A RC5@G.YM=C",B%U-Z75
PMXY'Q8%WSJ0;(G"=7<V4MY%47I%'(L+;N$\/$\W=S6(0/=>I0*:;26-KJ +<\-Q>
P<6L;[Q1V#G0M731%P'SP$/9-P.G1>XU?S+N0;/U9IK35S:-";[DAW8F\,X#"9]$A
P@; NT9G49>-\+;@U;MS6>G2A=HCQC@;:I#*0@A"'4<'O2F!WI.$V^EA<BK51S405
PV,8)H7$V8$:4-#HOW=? <RSKGZ)J4G>(C9_ '2OCD2 /UH.$ ^3$)^YA9C4I36WU
P?G& "[Z$KN/G%V>-*I7W/%(T^6-,: 'I%2&^-]HHTL76B^Y_T%/UM2;MY0F/WWY^
PA>W'9XC>[N?D@71QE/^RH!/-S>6DIHBJI_^Z,# ^7A]WF5R)(//M2&$_,:=M@BZ7
P]G>/4QCSKH-6^C,Y9G-'U(O/VRJ=6$ TY)?#+FXTH@7>AO1\MS;W(O5)* >V_'4#
P+@_1^%\,_$2T0J62-Q-C"\M_VKM>8!@*K]YO&^1,>[5D$EVC9-SI=%-RY^H)R/J!
PV\V41FIB=8/E?R%G=:%I=+ZFBF D/,<ZQ#5L$+6_HZJBV)/_%CL"<"V+YY(.]V^S
PM#H%%FWVT$$"S"M[3? E% 9E"3T45!X6'5JTV5EZ$3DOYN@Q9WP1[%)J7 NW=O/J
PR="?6-)BK!T&M;&-MSYJ3#0KY<?)V4MBM8ZM/S%<KV.(PM/:=R1>E[1IJT@5"ZZ)
P^Q5[!/YRLO>R><#TV%D"'D^]7;P#)7]L;"6QF,6XQ,9&M7'A^R^A]N<1F/L\9VS5
P @/HJ382BK_;R3:I=%R_$'8.,'Z3Y!K*-HH01:7/D3XECE"41U >;6JA$):/9.W?
P?SK>)79;RAB656$,<!^$=D2I%[6)LG:6T@KQD ,J)9RBM= #D,J.!Q1GS]+6?V4>
PQ"<>3S$I3:'TFFD)?D&?AG0U8]?JUK3[5;D)E2EGW(/;4VHL/#'0K>PXH*]F#@I"
P]1<NB,[E>OZRH[(O]3N7]9CP>=,HV3!Z9GY@M-X= B\0'K'1BMV&">RO$_'@YJV*
P8"+M,'R@SLP@W4H \YE"6A YS/Z)93_7*+X<ITKL@R+I,RS11WN=HP+M,W^/Z(SL
P.?FS:TXVG_:!U)@[CD&+2'ZHT$ <FKK(C= =;83(,3AW <Z.S>XD'[?D =Z 9):;
P ?'-]I?;319^O0XVU&!6ZR\YV9"]97X:30:LDQ#%>L^G):%A,EQ-TL3Z:#OK>;#W
P<>)-=$A<+/$IT5U,Z\7J'/H5GJ-NBQ:#18&X/U% ?"V,P6ICKVJS+X5K%&SZ[;8\
P94[VJSBC!1PB&VNZ^E:[L&LVI5LDG.+TAD?90.*0LIC8>(-..S>2$QO3=14".--C
PO%;\/5I0.A^%.#C5?XS;][IC)\_UTN=Q11!H%P=?:+CD.]M(+=@U;M[R_Q:U[L'B
P:,7:EGC[H0A_)7QEHMZ0:&AR9H=T@YC([= KBN^Q0ABVAOQ->(P.[NRQL[ !J[\E
PD:0&YY1M#PX85<7++/T7[]XXL*C&22!%3G#:T!!6Z<;L!^C=AL//(U.1H#GV_D#,
PH8@]1AUG"@37C:" 0'<IW9:E0'#@3X%S,8&%\D\G0Q?9E+)M7O#O_Z&O3JI''YLL
P31R^MZ$_[E,^NU@T+EY44?F?=^RL'B!2%#L\M03A94;UA@YMM_/XI,3MQ+I"- ?K
PC.89,98J!S&ZI 2?PSZ)21P#[2G8MK6>HF6AO2"8A&"F]O;<7FZ[BR?M[)U7A04/
PLO,F$PO^A68[M=^BX7_M<D9(=CR=>+)A($ ($* @2IC $T(,$*AK[//YF=4AOVMS
PJAR%%[B*8U>Y+L?[Y:"^YYD=68[S87@VS P"L[#>RQMH97"D74N\.9Y!A%:BJ*)!
PW< '-7P.!T%[FGN'CHWI.0BUB*=2.+-[/ =J[8E0]7AK0'T")M+X;+;@5N<;/A/$
PKA4%V*C')A.0P;#'30B7T<;Z ,?DZHP]#B00.)(EKAQQ()G8O(+[X#3UH'@\CHEU
P6:10.6*HE3B@,IZ4UHQ_%:-SJ^).@Y_D_R3G$ZQ,1HITI>R9#<=)O7)HF*0':]L2
P_*!93WJ" H(FF0S?&_M?XG+8?"?0GENHZ585&DZJVT/7$;$U4"CD K8.2ZV:SP^*
P5R FG7^4LQ*=3\DP"J_5Y1VR(JU$WF#LDA([0$6Y\64 >:[_1_G;CX!ILD1C/AI^
P;M#HL1,%C<4%L7M"W!=!.;3,NDB/;F/-@7Z/%(8-3"')C!UK$PQN- V<3D* J!QJ
PC/ZF/WJ8\HUQ*3+(5>2&I^#6"'3IZ1%LY9)_G K0 _5T/YV]J,GVLG?F;G4U6T-N
PS&MRNDW.P- <:VY27S'W!5^Z"]S]/HEXQE\*<J!A4OMW=*@Z.L#"!;8,C@=>Y90&
PQA>PV;I_'W:[IOK:?)ITP64S>S-Q.<YPA,#"_[*-K$B ,\_#4^BR]I8@LP^U_0]8
PN27%_8R8?"<JR0X%O+U?[<C9^"P:>P/_ ZZJTPUSF;D[K3-(P2SC@O9_WL0>D!2/
P+^];M*?K+562R=(X.2U)G],(Q_7&>I)(,DKE+%R8BR9)'SE:V-"#Y&PRC,')>F<]
PGJ=\;7:06_2M8F>,L"+Q7%+"[R@0KN=/&8WM(CV/.IPAIT5.\GQUQ57L9K!6X2'%
P-U\Q4'=9C<JZ$%M:4S+,+".P>.1>-J47JP1YTC%2%M]TTL6S:YE/Y\XP2R37!,><
P #H>: ^=I:7M1J[RA^-W0W>S:\#XX9=G;^L"A7'EFJM2!Y$87!5B-!52.(4*R/N]
P)T7]\C#"UN-4L]_&DEH#).ME+5[ U8W,B3T=_%MH;8#*=^4MF7J+/9^4(!A)T])$
PYA:B,I N'$IT@^\ZBXD21^MCJ@KGEGE^0@5[)BG=HEAS7:?_N^!A0:A]H@]];AL)
P)A,P5-@5Y5DI5EY/Z1%;C=E_-F36M>;RM+=AC=<E:=>.9F_Y<_Y<)]VKC^;IF\M$
P97\;BAE'<#?Q'_<'0*OU>O(W<<F&,=^^)RF\>0J\7[ZX A'V.@_:1RZT*X[A=MEW
PNJUK9W]XW-B/&/[T#NE'C\,;&$'D)1),N'?&[=<85U?XC "-:\HO;YCHR1AC5N0#
P8[>.(%Q55#W&T;B=1S('78S*AIPKZEA[MRW_#IR5N:FUO@=,=?F'[G?W. '4(5/@
P]YPOF!8G$/8;&&UT\[P=F3*7EXE39G5TN<TA6*[5$5G6$@0]+$6_AY'$7/9/"]%G
P4H&B/?8;I?G])GQ_6YL>["[9P:?F<M4]RZJHVZI:[V8G1Y3=-/4%6VQ"#0?5AL/M
P6RZINBP>1!H&+$F&M#3<-#1NMZ^&/4VJ_.G7 2S7;IU_B3R-:0N4DM$75DD'.-'<
PYMM4NB9@M-!\&?S13[ P@&= +.8KS#>NG"6N'( U=&=EZ$"-DP1CSU9$"FW1;W5)
P=-8(G.Z!YV>U (GZOV3MOKK-A'FB:ICP'Y:GK^=[!5ZU-<-#<FPTDO.G:^W##S7P
PTT:_U7X4ID@0(.@1G8 :X7#W!("-0=JG1($2&$FS3U2\8 .:(6GEIZ[ZE9D[<FK9
PM$?>+\K9ZS$^8;C07 @RD,.LP)OJ_EUO_=OBWYX3R\,BS+5XR8J')MDD-'B-Z/F^
PB[K^MFL C!YK-EM5-@4WA%-\C0OXZB;025= ]7E)0W:)*+(MV0,WB71)4E''@,=*
P8J/:4P4M$4F-H3V.W+1(F^6S[Q-ZBB?&TTBD[EBTPJ3=[MM;=W &?2X#E!,H,4*_
P=%+RI8%5OZ"H^ ,F0W"EQ\[!*!KSE>:2^75_V4JYF#&+4QD>\JLBX^1\O3AP.DV[
P;Q0IJ:;QC9[N 6\VWDAS!3ES$>8XG1QSD3J]>R_2$" A&6E42W1T8BER6)K>[NH$
P88JCT49O1"OQSG7EYVQG]I <^H((2L0Z0/\A3*_P>_V=*:(LL<6%.Y3[NL(,N/S2
PB7#E8Z["_#LER504)"YO;8LR!HBF(M#]W@%LD9I(?U%:RAA%J2JEZQ-;9GUC4^J&
P$KFFN]/<L0YR"3XA.G(P,)N@J!O:,:2H-@.D+^WWGN>D'+SG]J6\]1#?3>_W8L2;
PGU>P+_&8?*?=60Y9C&J/J WHZI)&2=#-I#VF+_M&GM*"9;( 1)21H[6"S+G.YU37
PPHNS:EN7 Q>YI5\-!LL=,C6GSRS:N*L'K:6"YM-X(+\3'$S+,+S#517LJ:_F1[I2
PO-:VN\^-46KVC91DY^GKZ]ZPTH&]5O\VRKC] #7/O_K]2]\L\K$'98E E^3,R_$(
PWY/TT=T1:&>X/.UM0@=OJNPX^AI!E>UR=W%"28P5Y.W&@X+SV.09L9\Y^:RV\*8R
PG:]OH!X9K3U]!I4K"13F@,#C=3 /+3XL"1NNTA[78-+*S>\I&C8O"E6?MXLU:I.V
PM%I%Z9K6F=+)%CN'\6'B)#)Z!&L][T@7CV_7J/8Z^>S$O[N5>D:)C=\>]=I"OZ/7
PTB$L8.9:?I;+0JP%5,+SVSF8L1WZ+!QPV'\SZF-W(!MLO\Z39-HG14YGMZO8*,R<
PO#?7: TTO<^'(MWU?Z]W).8ANF%C'@N R<)!IPD-"C^WI?=+9'=[Q;L6B (!%\BZ
P-I1R\K!$LQIF*3PGIERZ^ PHAD''*!F1O/Y59($M"[X:@/9D;F87X??W9T4E!. =
P 'T"/))M()=_,_"-?QUGFD.^.?;# #;(R)./V>;_,&\F,NL?(OASD;E]AG#(]DP%
P_$:"LCI>2N$,\IC(FU+>VBT_[X^(RHVEC'P99"L:RBB\QT7V4BQ8KO'M(]L W9FJ
PDH6;3LV93]ELU=QY)Y;/,A<D4\M9,UM-4*ER>$&7T$%D_U?K 3;8$"@=<G<R8I-'
PYV3=<-4^5;0-HN%09VG@OJH>HK!4E[H.OO=PV!)NQO]IG74,-VN;"4HNO*UEE1):
P*:4-GY#!OX\5Z,"MA&*<B(#G54KE#E285//WH SY0&9+VDDKW"8"^YZX5"P5O]\H
P9@<E8PBT1+Z*6>]A78+*1?ZTSA13/PXP0X(\ICK-$%?/3[U"IQ].X):]IZ[B55^7
P#V:HP""/$972"D1&W?ZZ6&Q1.?ZQ89:U#+V(\;V3CG7EU8",:ED:STUL[D8#7)/T
P;S/UFK%&HN@<9^D%?719A;ZW' 8<.]E08\.[=01=AI!PP#/,](LA+,\/S)&KN3&J
PX9T\X3M6E\.=.AZ9 ,HBO,SB+:C@)E6FOIM']S3U(+WC.R=P2/B=*C/PRY^Z>4["
P:8A:U!:6?F4O8V#JN_S$[K7BO1+L(QH/PVSZRNL4@[U&X>E^4(K[*=%,PK0GQ/_3
PP*/Z][*IU)9,[_S5-T"PD-5[_*7;*"1(U%#N/:W4I65!@&.2&0S= %U2X\[*]R\2
P^HX*'6HX.*9V"]SNCDA"NV.G$W$&U%C+;I *9KT%>>P[ZI:WA[@*E?65_(OW;[PD
PB_^,W%A1''2E5!M&M6/PS(;9:B--@=0I#BG 5_7ZUE,S&O<.OAG43TAXQ134K)'(
P2H7I 1%*>#=W:F4XHR4(S@T,>'J=]#IX3'/?88']NM:(][:L.,&L! ZYT5J,+Q1$
P)!6UDE6RO]NJS]_(PJO&#KW^@I@.>MKD[;-R%2U&PT?#>\S[/M]W--M%N62U0<QP
PP[6;H%DI$W:?B'WZU>)S2)3? ;Y]=GYV%YC!8.OUD<(6Z@+M'D22J #%:M=ZI@(%
PN9VM38>"KV-7/#(RT61BLNZY.J?J4Y<O(-&_C]'ICI8 HN,M*^ 6&T <7.31&;+T
P"!&A1GJJ+)^E5U6#IST6C.>9Q30V2DKDNE>;_< 0TCENW6[(I?0TCA13+%=2\BJK
PS/(*M.3;*]J]&TJ$!F"+:3VT*:W)'95NHE(Q/"YS(MJS^Y^#2@&[(;4,V+/#R"./
P>@/LE9DNTFC3O<JT3(OPB,I>I@#W7O->^3?,56][>G0@6=-1.%;.0?7 E(8QN8NA
P3:W57IUY/FL/TZ030>"%V[C]YAW;13OV\%DKT^-FHPK)G&S_-Z9:;&=\G*N!<[OU
PP )+Y4QL+I$>2B@^[CI+5+)SEMD*@2R2&OYHH3UX?%2VZ5G^<=/"E#%#@K4L8(85
P:+V<COSMD!<D,Y_(OB&55L8N"-H3RLF7%EE7Z+YCQ95W48WI XO2DK?(LVWRQ_0Q
P76H?T,@#X/%;B8;T8+@XM^0\Y1S^896,ZP7:??(6V%1/-*,P88'AY6[%F7OP-W :
PYCO\7!)3IR0 UXH7HU.]\IK4!)APM",4X_\[+WW2$WF^]E;,-!G]A G\)A(BK]$%
PSIS[AO\1FSJ033,ZC[0T3PYEYA VE9D"D&E57[]WU,EM*R1D)P&L$P=V XR\F>?S
PE<S2(5']D6K#1"QF.)T48*,RF!M.<KZ'<P5OL\+I@5R&@IZ4WI#-%]P,D2?@/O/[
P.RR 8R#UY.C406 2W*M*9$$Z!.]Y4TF(>VS2QBV(=VGI/%!M""-TB239%1EB"-MK
PC%>R],=79SHH:N+NW>1-@V7"HVZKM+IJ7LJ/9+M[KW,.M/\X(=>)W:3(![6I#)GI
P+J88+.6.<VI8NAT[Q*-6%3GY1&,D;6]VY+2BXE-VK6N_5E[B6W\[7_2C[&D&ZXZ&
PX"LID*/M=I[ZS]&L>1<,,\Q&VL48Y D<QB1-M(!L30"J)&-%'A(O4;_$9ZT&+_7W
P#'TI]5A-^WH"ALI-^Z67P>8Q7%6:JDSG6/$NR@7RPK2Y7Y;AY\HBDDGPVJ33%!<N
PYLD>2.H @.M8W(4M5LN[Y6":,:+DQ")?X<XXJL<[>[I4BEF1M?@WU1)T9V]CJ1(-
PYAZUBF?U#;930--4J#"6/8IC"[_U$)+4$_"83;*#U TF&-;2ZA*6+V@RE\:D&192
P?8'+/A"[1^N4?H^OZ%*D0QHXHGN<!YC(D-I+C2GI?@,>@6]>9PUHVE1T"L%<J+GE
P>M,\<<H#W5!\+Y18Z-@N9*78,H]-5]09[@C4**@'PP8&>M3Q>L 4$>D0<C<OI**1
P/=+<^OAU\)U.Q6$^[*72[UTBJ1^E)PI)$*:$\:#UZ[:7G&JLY!LEJNF3#<D_91YS
P<&LK\QATMJ/[])$_]F,/&)L;0^(5_VS5E>YYQCV03V!P9P6>ZU6;!F$<14[& 6H_
P,P]\ 1Y]%A8D$<Z-:\ VYT6E!]^@>0:6;?.Q+_S!88:DP[S;@+?.V_7)$,Y /8C)
P53C4!\RW^<F9@0A[TS-%\#4)%VTF=F<?9/6TO44E]NV:0YZ_^<6C:1_ZTE=.8%)^
P1Y#5:M%>X]Y.,IK!;"5+A1U NJ2=YPN\BHFC:AIE3_ EXV."]WH^2\V[O+'97]ZB
P9J'Y AJPL\LD]#Z7JA)T9+>_M<%>*@.(7&J=NU&!K'MFUWG$<K8)O!\J,F!H2BH9
P4@.NG@Y.$Z25,GL)_6_<-D(N3LK#RZ74ZK9X0JL]1G"BY"42MB>=TLA6>8=LCPX6
P]#*,,Y^7G-E+2*%*/1*,LJG?O571 G/KD>XL4)ONLICD?9R1P/G&A%^]7>%2JR<Q
P*PLZ<@P0%B*APJRZ/SY##ZFV!]$(\F+]4L@B/%(CB5!1)37] "43?K3#)4P\2*UW
P,L6>@Q;8S./,DN*0XLZ ;(ZFAA#?\\=?[5@=HV5/2_2HOM'\$R=,SN3S=%A,= C/
PSW&M"YB@U98,#C2BCX)W^Q&HP"3F>BL<XF)C'L"Q YX>#^]C3M8BF8%B$=]%XY.*
P'C'V0FAC1&>Q@IOC-T9)BM%O/X+B] 039==$<C;<78Q3AV)Q7[<38B@R]A:?TF&"
PY3S-<'*_M3+L.T)A^A;T7HC1<B@@*[VJ"0+H+\Y7(WC0=Y4<O7M^2L;XTE!<X*$W
P/LIS_1#22C?";%\0<:A-.(18/?I>II@W0"PK4Z=RF8L)-FFQ?C9X!&UX?A"H'J>5
P5",/7.@W@W^X:.V ',8;DI)O;X2F*8JAGE!'CO)S$$&=H5IC)T&K&1?L+ILS2PBP
P6Q&\0I<M5C.?X<]K4X??=E,:&6FX0S/3<*@(P=G84- OLZ@9&HQ0*(2'NM40H 5(
PF3;:.@Z=\TE?+V=.U/A.]W=QC6O2'W&?T@6LJZ"""\$JP=UP[H>DI_.:A 5 '[PY
P>%1&(%M&#*Q@<&4T^:)0]7L2?HNP@#U'%81WV]-]Z*7@(6+:A\\T;#H45&5H&(_>
P6]B;>"R/9\LA#DW)H!Y[!(&IZPT)FUK,ZJ&QSRJP:F;'J67G -P6%4@$ U??]$&1
P64X;K8HM#I9;$=LW/WV-0(%<2Q)_9\7J*'41JL$6-M4P5^J\=3$_DZ"N74G%A6O]
P[BHOJG7R"E=O7A7+-ZY2O2EP*T[\7TR!'!K2 #)>X[C9+W]R[D5OQI*TV$]W:EQ/
PW$$K*1E?LT!*2<&VH#,9)=&A<3>UM$7HW_\#R9Q 2DR,']R\_^N@,]?9-Z$CPZ\ 
P7<;&V9IM<$'R!=?P+"0OD9=S-.Q"YKF!/\Z"BPEQ9/G[6&>N21UGT];B'EGX:O(7
PYFI-02SB X)9(7;^&M;9-(_>L%.*"BM&2K=N;$C&,8X#6 18T?E.5]2N$,2N3>OQ
PB8#H=?#\/=P,?B8:Z2_M$E-S3]\&+VZL6O$ ^("O")"M7%&""E.7"D]+$>]AJK-0
PW9[0)WB$KBZQ(1+<0"TI^V^16GR]6;FTZ[]\+2)C$[[_YLF7Q&"RP+6/EW4,/C!B
PQA.**ABMZ\@7J<0\Y# 70J>*%V;S.3RQMW,HM9YPQ:7)2W,[*-VB8A$X55\:..+7
P.0#HSH#+5CR6U!T;>%VQS>.>T>UNRTA!F#HZ![;_J$ODC)^1BEKK(A3<[7M W6%?
P=2]2=V^4&^7^Z"EV\H)@7B4&"S#KRQ\ ED4FM9)^;, T;-Q&DT;.JK"/$HLYDSLU
P.4A4TP(:P.')[SU=F2.*#!AB\+?,-3\3J\41G(DV6..&%,7V^ZM'2KHW<R.R>4@'
P^<+*L-A +J7K,G>B&MP,_7O?%UBAC?N7[P6R;.4*]/_;_VM!"39P6JC&]VG#GOMY
PL9(C'#U546Q]]@]5NREQYX%1Z80-'*MJ-^-%Y-B5VP"@2X#'_?M]W/SK#E8E$#34
P1!EEMT ]?W1T];B0.)!/8@=67AXNQ"[%?SEO5U\10B0:6$"=HZ4LBOK"K#N2H?0$
P?O,!B-QN<ZQ\,UFYNZ!2&I<H  )_]6+84(><F-'YK3?0D"W&=_*SS>=&$+@S^VJ2
P\(TOO''=V^D"8:&'^2?B6H8&E:(3>EDF)<P<8?XDEYE!L9\F .^0L>32*^WV_;,:
P?:YS&*;]A@$G;VM0EK9$T%("B^=Z.Z/'!-K(8M'/CN\W1ZP.4I,A6#FVNAY'=;'#
P(C)/2[!;>/Z>?I][7*Q<6=N/_@74P"1,6JOST4^$KR;AP1G<[NJ+6H(P%,<*R1OU
P4BVEA$>,>I?0Q2$\?LH%JQ(I-BL;^>XE.%,!T3N4-Z1)CK:40K XX-CQ/0?I:/DC
P2%&--+'(1>)14#SL?E>U/$@^5<#W)3OB@QPMK9M6V1G9'*/!$8>:#HI)HZLE^KOS
P-I 0 5=Z;W?S$$;_Z #UKCRC1;LDBW&N+&,2_Y6/,?H$HBRU!X2C<M HR6,WBAB^
P'GTE^YE6?#T"M0.0+.ED4.4H:/L^X*UM/%IF9(/NB)+Q6S ;ALR=W4_UY0BXI.6B
P!RK T/]67J38,P$CEL/T)P[$2[02EXJ)3A\0/,,S\'7!K/VJIEV;@_QL08=>&!5 
PX/75.;S*S?S3B)'*>IT',"Z(Y%J07X*/P+O_$F7:M%8BI_O=NGZ5"IT_U,X'W!4G
PF\DZMY-S>2G$<EECX&D#ZCLI&?-)<RYF[087!Y4GK<FV;N\,U+),:$1%-E<W>@PU
P MC$YV83>Q$I$G\.'M%>52Q@A*[I:!LUAO1A?]_;+G2M$0:*4_A4=VHA ]JI'6XC
P%YA84-BV//HOE%4:DXV>ILE=F<9,*8N.[GX$;U$L@N:;W/W\<36B:@NTIQ_^C26M
PR#:6+E!9:XB_QM:I 9OBT4@"?QC-&]YNR<5>7.?Z-+5W\/]I%G/KTF.!%N<Y^R?D
P/)@\QS(.T7V84ESJ<2FK*Q+,PHI;:SG$(YPXMLG-XL#5]74V2JT/^2-3T,O(J?1F
PV8C-.)N3Q)1.F3SZ<%L[?^LC*\I9PR=[N:RC?>ZD062NFE1U/;3E1".Z1':O#]-&
PTCH_'A?V?M/H!>ODR6$SV !ES/G7>7' M KC"F(Q9=AH:'LAV5[SH7G 4+!'L7M&
P!<),+I(!37BIX#N"^JECG;>PNH\+D,FZ,>O_68L7;I9$Y@I VZ/6;.".:*IKK  ,
P]DS*QG'Q2CL)5 >@A]@_$;-]:Z^%453,CR_ZY"Y%VW??I[3@>W=.)6GIKK8H^!))
P\--E_(6.<T!'IR2"/6C[4+Z1N=FPD2!-1RB-MIWN=:JD:6QG;WEWUBW^^14:KI5A
PC\)HM0H.WL!DQ,)7P&I_#Q?FPS"'Q87#-VK+AC0QAL!HN7(MR=-6^K&H$CF$L09$
P/@+,)W-4;Y@WHL8-7!79HG*>\!=(XLK0!+NQ9# _&#S5&@\CS%$.?AZIG#CY"@U5
P.Q3GA"((J=B ELW6^=S&<*^J\0&UX4OE_#SB-_HC'[OI77GIO_IS3-Q3\ (.0M%)
P.>X\(N[^2=G,9F,%&B=LX FV"G__T?EL\_BN:@U&9KT&AR$WGF(%C06%=*<H]H6U
P6BN>>S;N"S0$@6U_@T5ARY7?((HP8<IYT,_EO^"W YFFQ4.V]SHL4</699A %@P^
PNC-VCS,)6_]'#1>*3!)^S/R5-%K$;6&1M0XL]R.A\))3X?UCA*\LK^<%'I>A@M%6
P[V_V&'TY: XQ.-?],:522HN8BNP660<SLJ,:+&K&.D25/'HSL(LUT-+;+=NZNRW_
PRAA7K()_JSX)6\OC&(,^#>0*>&MD1/?BU*5[JFQB'Y9VR,D68)W:X_MJ%_]#!C)$
PU4HZ7SZJ4<3KL(F'G0*NK9U3>G:LX@YI-B!93FUHOAO+R7"%)\+'\L]?Y2Q#5'J]
P=)4U"1OI):=7%0 -ZUZD65."&TP'45* H/J+?/)4M?EQI4'$:\*37IDRTRU!(S7)
PPZ=;TU0@SM/.D6UWS@A2O61<^H^%"2<%VK0BCTLX%].!ZS(2E5Z#SOWQ(%H*5%[]
PVN/'YY[ =1!W\7X[\05VK'K?@M5R:&&K4J?H*^:V'D]_FA+:6D6CUB'6<^.L1GFR
PQ&^RM>_'1&"Z8"GPDX+U7S4&Z7+/HNP#YBX0/,'=.UD/$$O3YOFD=AR9#O66BGPZ
PZJ>K'8.ALPQ]^(."B%LC3WPP,WF;CY7GP98*:BB5,'627 [U^(-H%/A$Q";QETK%
P+ -><?;150E+P9PC^E9<)E87XH3I7=7;&XY#PO06Q(8:,U@OZ2UXH%TIQ R/*>+^
PV7 \AU'863'?EQQVQ<ZS+K##$B$LYA Z/06Y6/KA+CH<I]WL#*CW9N8Y^*YX@E0+
P8.U+*Y3^RC7X#XUJ0)F)TXJ18U>]CLKC:0(4*EJX.#=N6KQ$B#Z2!"0"/#?)IO=D
PKS0S;=,IPX:(:M&C?1UZXLI#FIA,,@JB#9A];7_.-+N(,-=I1!T#<Z*)U/%K?<K)
P:?_I_#AT9:C9]W A(5KN/8<Q;;(HUB%*[#R]1BA:5=VPA8X*34*U?2>>:'#,$.36
PQ(D<> .&UG(@F#EMZ'BWL%^H0JN]>I[Z&H$CA*X/<NU\3&B'(_U.<.,N>ME^]S8>
PIQ[8F1&DM/U,$^6_$RZN\,M0.I%JNS'M>R%S(6I' 2.,!D8%B983SS+F.R*/X_Y[
PHEOQ&M)EWE?$<EG'HD0WL?LTW;,.]H#.2G3)!@ 1/ \7J  ^9U9"59E5-306UGP3
P0ZKOE0F&B#05P&WDY8G>((>]*9Z&>8S-/I0D670'$KEX<O<-.:5V:)]B+(>KLWVZ
PY_K_[GRNC!.^*FFEG$LU]"[= :.WS X!#[%F,4.T#KF/(6D<(*PF;H1#X\2IN"+H
P-L45]"/'ZHIIW)13MG)_7!*DL8Y:4,O[I'674-OM\OGXCQU*"KC0<C92_T/ #\AW
P'?>FJB>X\!=JQ<8^9+00*AXIJO1CD3MZ-;JOZ&M@;XNZ^D_&=_JPC8P097C*QN./
P));TKGFR%7K=5M4EC"37I#KK1S-.M=A+'E&BTPNK*S1P'F[ ZG32G7K_]0%[DN]<
PEIV#U:+]5PAAOP6;7?IF4C1UN!^!L54Q*YVM7 Z*L@A6X!!7RFYG&,)FFLFGQ-E7
PEB/RFPJ+$]\K$JGHTVL4Y>E!84<I]UV/A'87OO48,,-X9(AL"T^L.%*"4.%B&KK[
PO=]^-QQYQ2N,S+/9:1E0O6;J?2H903M*D5+/$\-1$-J4"I1E_Q0#\IM0I<0X>58F
PT>EK!8>7^5KCU2>VAW2L^H:6:],/M='L+-@D7:O# 6VM(* _Q^ZFMT6^;5SZ_KQU
PE0R\,BDG\7+S)6T9J(P?QY_M3 WV""=A,(+=5!1_V+O5:5("XX/:6=8TH0BPXV7T
P[?.Y:^GCN:==^U29OU[B16C"C])2"P ["+#,J*5L==DLD;W>DPY[U7T2H.@Y]A,S
PA':]#QBMMK$Q5"@>+_28Q+*W!)6\@CU=3(]W<BCU9&)H;-3')7<O?RJ]=$G7269K
P$1X,"K98"8T=';34X\'&_9TVP?2KOYZO;VV%]NA4$[X.^(3GEDP(0[P*BI7D&[T?
P<,! TE3"IJ _)@W,@$K[,E](V7A]-O[(ODFFC0H(PXGE74[UNQQ&-H3RB.DX$T-]
P49=XD$UV,72<\" )[?=NVX4\YR"4$H?HU2#$"2&-&";4=EZ]+&,NCG-1U.8XOW]<
P(Y>TWD;<BCF(+*"1' "?C[ OXVH5R<=[4;Z!O-9T4#'_^&*1"K/(R4),& 0I.0O(
PI8V2UK/.A4V]@^H]?W;LH^)UXT6:4F9&F+W/O>X&ZP\0FFQ OZ-S1P7H7@$1+H!B
P>&47L[5+"%%X,R!)QAG802-AO0P64P7EQM16:$2*&P+ARU=GLZ_8/U<.A.[%,#=3
PX*XH^A@7BIV LID0L\MU>YA:]I(Q5/^;9)35@+?D=09EGB-)'\"Y,GSX/U5_!%$)
P992ZGRKL)3\'8[:$.>16%8@!J>DH(N)HFV]GY=CEX5>JQM%EC'T>T0ATBHAXR-[3
PUXSSCOF[B^V3ETWWH<"BVJ3+%:@V[F>2(%DC@SQ?O%E@+PE,1>\WJH5)2+J2]<GP
PSEO)#!M852C?.%R'[;NW<-B3XE[T[CX4T8"67RLP!*<;!:>$"I$9#6E^J'Z]+!&$
P_EG X@=L* 7SPOIV^\EXO,/6JK=F?%YAK6ODSPBI\0',E7@-Z$?)?O4&:&* VXV&
P%VVVVN_0)SHK3X^,LUIH$UY6/9E>A.&5L6/L"]E:>[>15HV5Z_*E\ZLTG%;'R)]/
P:E-Z&M/ ZK:_$7N4'5G;NM$HZ$AS"NQ%6,8$%]"/JXJI0#:)6DG")B'XL@0?5%>&
P^-]^K-U7[_WMJ"Y\!:>Y %,%UJ"EY&=]C+S:)EHT ^Q.7<_3B6UN\S.<'Y.2RA3[
PT:RYCT.FQ=#'?W!JGW^3K\7BZ+!,[D3;;9I&6:S]&MT#9 A 8;N!>-$]F \%U9A!
P2&?TH!YK1&0.4-B"'MP%(Z50U[(^FXXV4"4VU,4'B(%'O*0.; .=ZBV2"^9?-G0!
P?PHX"#3GKYV:Z2^9)"3FU7GT.!L2G8P$>M?53'BGEN][?&(LA/ 1?K24:YG6!L0F
PR'$,YG?3'J=TS_I?S>OP1CCOC5DQ0S^(ZD)*=4=S  B;NSJDZ1Y(]FO08S<W?5BF
P2TKE@5$!J@!'U5@XV]_V^W#CJF497'?O9+O[RZN)F(#<:T!CFL6FSNE+=AC%'R#N
PKQAUG!M)HIG&JW 8S?PFZVTT/+,A5XOZ:=JR+K&*,% QJRF&BD5C+_!1EY)V]0!U
PB,]I'=I].@?G<?@A<-3Z8OP4F?Z@V:OHD4<N#Z_46\P)%16<;;HH3]@HI[KRW2AJ
PMT!\0&G% !I@*%>^B2^=Y:]1H"F (8T12_=4*,KVM."H">=4CV-:W/YE+';FQZ:.
PBV6T%ATZNGI/P38@+F2/3UD70PGYR&$#-/CYWX)J8O%7N34JUH&K"U<&<'W1\G2_
P4-8$PE,RTN \=?AK^?<D+-M+[D>8>R\$2'\$>^C-BL2M4P-MQ*_<7X%G&N(<-?<S
PZTPA@N"\,.Y6;?>P@.EC4?K6?/:<A!1H*.NO8E0SF_US +5'A]PJT-LS*4"%C-[#
PEQAR7KL_@7YQGG5CRZ?7=2%79NHIO<\;];&S%(<VIJ*FIP080()A *^0Y&:T:<> 
P/JW+#0>P3>[-G?V7DX'+,O05!62]<'6\N7X!O=?\+7)-.-S)//M\]X^%=1 1'6&T
P*.B(P?$ ORW98D,*%7H8%MLBH^;9?%0&E6IET.I7W@P#<784].Z+42UNSR^R&XOR
PP&EUTG 0B)8)4)^]C*_.__NL+: $P(T0&_I82S_1O:RE#N[]-Z\G%G[^IV-<<5)M
P@3V8FE1<8'4:%@^AM*P=Q\5LF3'3TBEC%8%8R6;.[2._$@=B7HFDES?9MHSG"YL%
PBY?VM38SI2(>^2[\H\;MTNDF$NN$+_$IA_,W(?Y^(V:88/JY31)Y5F$)4@%"9E@=
PI2G+"F"M\%>QL>*69(YW-4(MZ'BNC0"*L0ZL].4!S'>S)@5/R+L>JMCP(DI^5S]?
PYG,?M33DGE:_DT\S/\Y3FXDRY\0JN-NIM^CX,5?("TAM3U^K9+;)/'J\VX0;NT%M
P3K^+VEZ4_L4UJYRTF5+"D[8E*G4Y>+0H[0C:;KO3LY%X5WA$Q0;RT!4 #E*/,\UM
PWQDD87$W5?7M?[*V&TNFN#82[2S /*#U;0*JGE,R#SJV G<9DF?1F]HV%O%LE#,Q
P#CD9[DP36< C)W3X.V[\.XR_>23>9=>(C1"6;6R0^AUV;= 8P,'R%H^(C"#KU-RL
PMGSN)A,>\)*Q+XQ89XICR*,YBS;5#;^,Z<;86M#!CJ=B"*++5,"^K??!U7WWB@:\
PUDX?^M7KCR;H9%=>3 [6^;C/[-= G[X, %'R:0A33&ZWF@N,I).]-EGB"I8*8[EU
P$0Y,UOH2RT+-M#&=8/'Y:'3YVLQW$(>G_+B($<#P01(EP5UK!4CBM.2.H.#R:?7)
PI5 #O,A[+>QY/3 GR;SSPW[^0IQLQ8$B4W$&$^N",:N=V8\Z";6B]$=H>F.4G4U4
PX*K^_CF1@VBZ#<D$47V;P7!?2VJ$)F>]0ZAHEO<V/<%S*I7D:$YEJ9VUXZ (=P2$
P7%O5"G'>C&LKZ<%[>OM4'_3DT-;")1VW/"Q]T3B(KL@P^=H'ZT8VA6R+]CKC73;(
P0FO4;MFJ<908\%T=,WV^&JAC$5-.G1L*. M9O#Y_:R(?")K/[&X LMR"@/?+^303
PX.-FTXN[>)-+2/]LTFY3DX]^,(GKJY<<&>ZEX$I#70PMQ]3V+\/+,O88%ET@IQAK
PYNZA>]E&?5Q/EE[8$4,_M#1IOV?O^3C, WGRWDF(<,7LYWM?GN34Q<Y<F<1P'JJ\
PL#/[BW6O[ /QT4M3.[4CV9I<43CE4"D+C8+5A+K8)B!*??XWQ$^T=/T@@+@N<C#W
PT_@$,1P[J (S 31Q% M3F[GXP7-/@WNHAQQ+L3#_0L/0#,/D@P8N-852Q6#"4GA]
P+>L'DW4"O&,I2W:M['5A:O.DGF >5A_XRFVTS7L?W(B6G.182!C(EC";%^X+G1V*
P:0[M6P-01R[7H7+H[^ JWE7 7^*=DW(7SZE$"L$J?D9,\Y8 -13!F)/9Y1@L)2T\
P7EUDT2*[I%(USR&TQW^_#V$V_#ZW@/ZDU-7;[C)[+]BFI^$*SS[F\U_S):FZ;VJZ
P)5K!D=Y*@.[KRNPGI9"4)I=PL%6S=/A="X,@K?0FH58\;:='+CUW++B1)2]$/?&<
PQ[H"5@/ZB(EPPJ0J2^U.8Z\-MH^\U830QYTAYKPNF[/3$Z=%X>LX>-'WC*T'*I*U
PTSVF".QQK!) F9#@<"65%,@N3G)@MZ*- $$11;+VW[A-CB2+^"<UEI-O7:K'T?!D
PESV.1T<DC'>4_PQE@?<*H+F2QD8ZL0@=D27!':&$K*)//1'_G%YKDTB[*3?_+;E?
PYJ?06U0?9]/([H7(X9A&F,!-;.D.9Y+03 _DWQ=YL'1Z*'9A'ZRKJ%\Y"S(!,85V
PS>&25C--Z/8#XR)O#J;#8P2IU6@?+2L%[K-6:,>;KE&9J#XL+B<!&Y <=M4,%L:W
PX4418[L#O^I 5_A0#">X(5:.*S[$D4U!PY FT5 8.V$MC?_->"W)PHO=QHX%Q GV
P_/D1$T& ,4<X'0'_*Y[1LH-O)UX?!A^-]Z?5*TJGYUA@R4X>,H1^IUI%DS?3BVI6
PNQYN- $&<<Q%P5R>I8OL9V#&2HQS-J9!_?,QHI(AC=;PR7^ CQG;GH*1QF9[L%:%
P)1-Y)<C%NFLFIH$ ,#DF O/0@^Q$8&3LY4&Z9#-FL0*2#W*<]3B5CEBF1L0+4[][
PNY?\HESQ7M00%AG(4.7S]:/F9Y_KQ1C:@2QO,C!+QVQ59"P%GM!/;76]36]O6S/'
P)F]8F#[ED%EW^43#H$W"J_5-B:V3[!ZA/PEX6J-+Q"+9"TL$JE)W,"[T\2W^4%MJ
P'%U>2FMD-HGHI]BN%[+2SE^ZPJ#%IN&T/37'UM;8 E^E TEU'CY79</]M%]H[CN0
P'KXZ@U#YF2IM:8Y6<+T87F 1&<;OV@.PC8":ZN#U$"*@*67$NNVQ@@1>S,EF@%-F
P4IMBJ[DZ2YAH7;BH(%J/&]+,9O(R5Y#O(Z+[)M\TUDKQA*7THCU#ZE],6C/9$"C]
P3DH4*F3VE9C-0Q_A77WFM0#\=_96B&%>LE^2HQBXYN^)T=B^U.+>$-HJ_'7VNT>9
PB%X@8"ALQXD5I8#2!H]Y?1$FNRMKO39CY6A1B)<%G43FQU.'+O[SY%2M&*UD0W._
P3JVA"_%JSUS$1>4^][DR"6,O7-MMA*0"X5,O1QW Q?W<:O:*M![ZSB0@""W 0:;U
PNB7X(=L-:"B]5;IIPY1R0L?C3;?1'-LLY8K*ZS3_<NO6&<_;[&OD#KA$ W&ZQ.<3
P= %7K.Z&KGF'3%@NK.W.S1R) <)=J\;(01.<LC3LRE[B5_%@%W+F?*E[L*R02\P3
POP6,>D-CT?:<Z3L$H4A% TUL^G/,.#A1;.@J;@W*&SSP2E-Z)(]1?.9X;Y<=3!/)
P=;L#%-$._QV\##_IE/._[W(-9+G#+*B=,06C-]I8>'>-,$6I 73V3D 84_BO+8<A
PP4LJ>L'9V+%'("+!8G""I9S[#9__(,Z+V9$IVL&)!-\5H'X!_YDW@4/F\V^%U0]5
PY+QZ<&*FEU$G:)WV>]F]BF<4<L1RR-0Y TC3T5 TRZNV;LD,FK5)BUX-#Y&5**##
P[9UF2X)(&,X$X'_RYKJ1LXW.J\<D<$+Y<N<^QVX.R;:"H(T4:.7PT<**%$<8&3''
P=33'_8K [)48J8.[?CCP*!7$DX*?S_X4)0O+DP\)TO"9!_DPSHC%H>5ZS$HM@!P$
PAJY'B9O])8(?H YHF6UZ#;/VY(+\X'J>U'V!53L;@<+K\YK8O*])V!"0EUD1;,H,
PKD\=.]'"TI)RXQN#^S.U->F7 Z%(:2Y.)J%%H3P6AOQ1>'+RJR"$F]O"JZ\I]N.#
P&&!>2.RWJ9&TI\]&0*P* J1U/YU=!&8?'R-@_I2?#FIOM[:6MY67"<[[^':_@$;\
P6T3C<<K!_[:A*8TBX-*R]:!R8Z$3&=IY?I+5!$B&K5"4F #3J HM]=C&QQUZB(/ 
P>-I?98,'RLDW_7\%Q8-FEF>E);EGC1G]"NDA,0<! /+S$3R[D6^3R+L,X#(;(/?+
PH6_F%> B+5Y@$^2[@Z+E7P1H42R8>+N6[LJXXQD@:A"EPB[A?%09T49V6"02O7#+
PBB]D *D!W*-(9;PE8?F)]N4Q(1"G"U'^_PQQS.ZG/_ZEM:Y1)D%J16WE2UQBO K9
P: ++,6RNHZ[]G9<(1!^YG?2=72K0>>U6["C2 X]KM7=:@ ?P_WW.XWOI)?)C?\[;
PXG2O5[($Z1C]Z(R+H#15%/<WN6NUST8?T9^+5=@ H;$TKL[L@T%O9E=I3+\=D2V!
PH8R@W%_1OYHD;)9Q;82YDP&:A"8@U<P4^IJN1NM>N,'H@U:>6P?\1^#-UZH*D,B^
PY.@AEUGN+FY1@1/JYW]>N7!'%R=#>U8NY72=27VCUP@BO)0NB2$%8R<]+]UD+]^[
PP1FY<A^ 8A+"4('UM3WH OY=61B+>*Q>7))4 NNPE)-%Z2^+VPC8 K"$C+\Q/CR;
P:VNVS11(<=D3X>SD-+4=M-I2,@16YF+;F@\"09VH]$6P<D=URJX_*Y*!YQ?M_EMU
PBXG\]3YR, MZN.C<J<IRG!_8O-OV<O7]<6UI41M\+><P+30F*K@VS&%HK!$FA;AN
P4[GN?U,[<N@_&3=3#+-@1UO=\Z7>A \[:&T :4;7VXA)?#5__RJ$'7KJG^_K6"]E
PX=#N\Y[(+4,ZS;BD$(T0^$ATF6/C?8^5XFHUVPOT:"8.FJ+.P<THM. +EE568-@-
P#)HP2BC9]"%Y-?_!,1IE<A_%&+P.5HZHI3T[K"#1L;^YLO(B;S=!H3%-57;INEY8
PVG$$$C^JGZ<1NLEYCOII"W=^8&K_#T5"9T9GF#X/[A/D/Z)@3#]K'H*9QD(RC3(C
P.TD?7A<Q+8_;''V([WL_1CSV*P0Z0D 2M>MN#NLYWH(:>-:&?:=QF$+TJTZU4(O;
P(RH^+KY&4BF:U-0 #VS8N^PV!_%&V><:IAZETX<.$&;R'G+/1K")"41"G]4%/BR^
PY2:QC#>/2LOC>;;N['N'5IHR+Y7C7"X7M4ITFCUS?<M[Y3Z,3=%Z +3OLTU'J\F#
P*O&E+N&,;Y=LD\7K;((AK:2)/WN%"?U\<9N:>7XJ(B9S\ZVQ1= ,U(?3]/23_\80
PF9L=*^--/4;4F]*XAAZJK=/Z1B5Q+W3&>7+^*1;YJPZFD;ZT-[<C"MV77@'E"0<F
P$$:W/FH?%HSD.?L2!2P!,BB;.MBA&MW3[I*,UW<7DN2YDB%\C@G]^2<"!&BRVTCP
P!7P#[\II\A..(06IS.308I#SB8)0J"G4H%^GVXQV34R_P(D)SI-&?CQD8^DI]WT^
P$W0+_=$Q&N!AP>JMZ!H0B]USFOM*3=9;70\A_J8J^.ZZY9C%'NH4%JFV#BGZGNT<
PF653;HQK8_M6V)^@/&:G%>S[0M*K.U&J\1JP?L[MB%W!^FOO0T(F@ @H'-(V(QWI
P@CYKG=E8Z;EN[;.B8DJR5'65S]G8A^QWC<ZW1,B#)"$FG;<@BF=M26[*C-<1>28Y
P2G7KMO,")SE;'G0YX>-:U3%>WS.#.(6 UU[_C?Z@-[YGL5<L)$+U@H?)D#  >UTE
P:!?33P:3 ?=1;U* ON+;%S9',8M37*G6/J,^07HNR?AG8!>6SYLYWQ'T.1J!'OT/
P"4=/,Z:"OO%QW>%9),LE3I@V<NG%N2_+[A&9-)#/@_AV-!3YQ;P "JHHT>XV->S5
P\&B&'[C"P^6T3F>@&@H7LV#:F.FVYU#%Q,L8D3IJ7![B@\86-11]3WP$@)*YK"9X
P/DN;'( 6A5$)+$#6/''-: KXK!0^E;J,^$^1?)1HN4+:1LPI:J_'?TH[.N>3B;E,
P_>*?*"*L_'C[V'^K3;[34Z(3W/3?D[6VR]/<"M#6]-4P>R#"<(270JFK ;Q>!.)I
P@NR'&>3CPQ^/V.%69&?>6VTZ_4;]<%,93T]!+O^I\Q1PMG GWU7>P/7H<@>VZ(;Z
P3KH$8%3/C%5O:P\%W):M^B^I[ISLS&A#;E!5WI-1'?ZT.ZJ>(J,CA1]>."UU,=:[
PN>XTUR$1 ]F-]NI5HE :@<$/=UVXJ-(/07E&\?M/]'WJ-C]57ER*^-G8>(<%A..O
P3/$ [4 ?EWK@_&INDUL0\^>O<M9O7:+?U-2GUT-V8I^DHL6/.Z9M,BC) 1L V1_)
P)P\],.H"NW":KV4*0VFJ2*T:S3K>KS&+6X&:O<F3H:G$#]N)5^S"FQ./@*K, H+(
P'^V*#8J'+K'%ZU<'2K<T,B$\FPK7:5!BK!@;)L2*H/PZ,&P+2G:4BH"3:TJJD?7(
P98Z]W$.BOA;'K#">__+[?ZM]&CZ )U.E85!- '-_\4:8JRTEJXP:9H+J-UK,9T[ 
POG;+M7GM@Y&;:/K!GOOEM#9=3 LS$33GRZOC8QQ89D0^\L;@D> K]A"=NDOV\"*X
PFQ<"]1K"*PB8O _P?K@*<QQIHBKI]Y E@D;#D;;F]I,[T JV*MO(<"E6%.'O(L4M
P*[L$27#\0B#>[=E2D0MJ^Y>?+MR&B<UA&U/< 62:9'K8#7J^LC_O+26;Z6CQ>\]P
P&Z?+A?.?\:DQ;'G GH=LNA-OXG%R\<% 3C@$FT%L%P6.C55>8!',F)Z?F+R9%-),
PXY]46LAE#@%%)/D+/-.E[8U]1"1P! @T]2F;#3U3]1-6[NGSWT"[7K],:(B@%T"L
PF $^(%E?O#MGV\IH>"]=K_6[:KE27>ZF,B4AR5L[$V"9+DH&'.TOX4PM*YVMD=ME
P]R0Q+&+$R^FAV+*D=GR^0!REF/=>JI-G8@8&PB[ 92@M_#4TA5:AOAYSD[-RFM^#
P5OMLH0?5T81(B4:Q)BJP^"7V[T&8OB&XF']SBG8E/K11^ZK$F176CPQR1_:3F4%M
PL<:TR!BG7\GED-5=L@DD]F3<*A+H_30\5AK*(IW>29@[V;>^)"N%+K\XIQ&0AH]"
PA,\"4!)*FN>A+4#XJN9)-ZYF0%N%2P\_(6L\,_85J[7NSBO\UOSH_<W(#&;+P]_'
P&%VR9  G%R&JF1LL1M,O%2 ^1OV@JU_83XJBV=:0IMVP<R&K!<IJV!TU>_TERB00
P" E.Q'41Y2APO0G"!=8T2INLQ)F)B03!/2!QF</R"I3^-P(&!)4D$K)S."F:44VM
P"S9*2*/\>2'62J!B=ZV&AH?GMN7=45!2Z*0+@Q\^1?7Q*RI1?,$)GN5E\C%U:KD?
P[)[];=,9#]K@=5WI]_@NX)<W9[0":1+(4H1<T3JE]H,%!6Z3@%/KQ^@%.H.AF =<
PHWP^VW'#OAGXC05&RQXMWC6QL9JU*C*.L;7WZ$.!)-]:Z.V+@I_%94N]<>K)X=]P
P(?91NI@'B4*E)\B&L<0MKQ']+)D%QI/?SY@ HR6-LO#+ZX.R$P:UT/I3EP<IEW.M
P(F"S0=PBS?AV\O*9ZTR"&\)'ZL!H$!Z7 3K++(P7Z%12E42?21[Z6>AI'U7[JGOV
P7&?<"U+(]=&,5)B^T9#XL[8[M@N6E)<NQ;B92+2!A>75=OU>/^]T[@-P=R?"%8P=
PXDC N+/<*C"GY"II^R!TIE";/MW@=<.Q5=.' 3X?!0=\:O% 5274>FNB56-=NN[P
PP30$]ZGJ@O HL?H/6NNTVWB<KN'/RR51\JP$]4GPZ:*18I$ZUW/&%]00LBYJ%B52
P1\P,4H&!4;<G'%)"YZ,QF(#VGF%CF\';;O]FD; $:6<;XD,N.2&7+HMK](9AGG.L
PL],B# I;P&_@ZB]!BU;B$KSB3_D>(AZT6M5&LUJZAT^NFRBO P)G-1!-GLG-^.YP
P>QZ*ZO9-Q;']#,CG#;V.YJLJ@+'[ D.F++/0]"=M$#72)!TI&)F4LO($E[<;D(7A
PNM53BEG(9^\[2G3V%%.SW\[9O*&694:0:LI-E, ?0Q8O2/9@5^H=4DUX&9IGY"1.
P Y-U!;% ;^N",;T<2CRZ8)A-ES\J45T*G@25%.IS_93E:19&.A9\),ER9Y3"2B+J
PIV-.WXCHS=<.=:-Q)W6V/52YS'*J7]P4M1 9Z<&-83D<@NY*J07:HJ\<PNKJLZX&
P&=*NZ5K/S:_3E]%$!7V$EY"2DD]13=SG>.J"O:)VF\W"8HI2EA_O%VH?^L47.U3K
P,]9&*G5W3M:;)^["-_CC>;PQ.R:OT\ ;YG)<'^P$A!#LRK'#4@3 V,I^3/R%M2)D
PTLE5I694JX;7/7PP2=LDV04N^X-_?"WC^:=T+*5L:P50LI1*)8*\R1K(5]K4U_E6
P>(E:5WS&: UFN<!7UV U0$VH34<X$1*]3N?'F->+?#3=@5)(G!C[G':]M<)^E?4J
PN<VR#7I@>J)PB;4]L(F>"[BUC@ZX8_"Y.98'-J)F]-4MGG.:KXK)2'Y#156,Q=TZ
P>"X^Q8!:Z&6"JLNG+/%Y0UNL;*W]H%,VDU*S++L[]QW__9TC&!A_$_!)(>2K(&9=
PWQPU6.A%S^:@U,'7/-<-\TIR:[,VO3/XA44+C*G_4O>5E!FIP3<%=8EIRKO:A@^;
P;)O_V&M7..O1A.+3-MJ";R/<% <''A#8U*+^:FFMI()WA6V@#<('AO2$X@N-TQ?9
P"VDZM6'K9 *;', :)V=-[GU;2KW*^2M,&.G[R0CDUP7D@0U@S(].-<WX:I98VR@,
PLQK;P;!F.252R\CYJ2J">;$BKR<UJ%BSRYU1F/+R!S#J[SW#!HN^SH'"$G?OX91T
PML%LVKM>S2977OC&9&+<PAN]Z8]D/5C)N#&U?V1TW5RYT%1P1V%=^FS5-A^QGM5.
PXQ29P*JL!N!_4Q:E$$,8*>&NW[4Q7EP0@1M''(XN='S&'<_"+DRW^.OYPFJZ4DPE
P1Q%YGW2P'?X\ORUVL+' (K=UQL==C7ZXCD,'=1$#[]]_M-^1OGWKCC-Y'[ .RW=6
PK@RG;SUGXDXW'>JW_@+6NQ9]+I_-O:(F]MD.C:O=MGKLD."Z4.8[<V+/CM(7@:&Q
PI^.$/C+=M1:SV&/XZK4D2UAX2>$5VVT;/?6@'0^FCH64&XY\J&6\ZHTR=WQO006\
P@]K?#(%CEGSHP,4NCA;#PJVOGK/_32(#F=_=$7=G(P-E^NT",5#&;D%A5-"B_J8Y
P:$YOTMK^0^M%\$ *IHAT0,484MMPL/+I)+1M%9C+Q/ICG^7*/&"#Q67NZ_?-/)*Z
P,/,'=GLV[ ^I-+2E)_L#Y<18N=_$OL30G!VM(;\6VV<0>'!*"%0:F\UGO]RZ 4J!
PY$G?+?5@H??PLP=-%\IQ?J^(7VN5_6([2!_V/J2YVV41QEI4!WJ,%<"(^I4#0   
P!"!WNSC_"+[VAF "J2FDDF'RM^@#V\" X5C&N6\+C36N<(LB7MU69C]Y<T"T4Z#@
P4$7HJ+5E :*9P-^(<$YJ_BZY@2FLFD(-\=\GR07F'8^;>+*P)9YVJ(V9*9FY-8 A
P>R72SY9+0?\C!L*Q?D"88EVP-IIY: @PB7?Q*W(8C$SU7ANZ&(8M58T/)VKZ#^%3
P\]92>(WK1H)T:1!L/1&'("01]"S'?YEXQ#$D^:T'4<U!$13U[?YA[O1Y[!7R 2W2
PH9&Y)S+0Y <EG5-W+)NEYUP%:ZO/#N\!JW@=B9P]#_M'S6WHQ46!^&=V]"G='/H$
P(KE<]\7!K=<6@BP3'K"W?Z3GC0LL'1C&H2]T00=7X./6L]S%!M6*X3,5DB_C3[6+
P+C@R/86)-P9DMBU?(8NW?"  :Z.LPY])Q=5EOQ62MCD@M63-WT2MG^'K^6U?I\85
P_P<>D]3<09!+4Z.D3OTXL%3H8/3YV+5&I YOO[=$]0O0:((<+S\V[M: <JGR],P[
PFY2%134C7BNL=LCW@E,Y_#>9%I7U"]@+0:6[V1]X8/$H+]9H/_OP'8J(@!R/7D+F
PH$*-O@^$U.M1K(!O5"<36?XVA5C>_6T[9MS!^XCJA.;.?_?UB88V4K.-.%:9F=8;
PC=Z+ [%?#PZTB(,Y1+F68##L4LC<XASE292^T%"MQ3.,7WEU)G\494@:6G,!$O/_
P8%:9'CD^Q42R$6'C3C1R4)9LFTBG8\,<>F L\ D0:(J<NM8$&WXOQ,_<!T&"<1VL
P:W*5TLF$?0?K0Q.<0S\:JO3&$2)#42866!;G*R"TL/.K^KM&48O;E"^4+R-0;CXA
P0G,H$(A:$6CW<N7YM)7]RWM6HC/%&>]4>=!7/!2A!:^&1R<I'6:=GD^7((.N=36E
P>.7^J:>U?1$%I5<8%C@#*4%N=*X@MP=7"[2<NJ6)2#],J%I*T))_[X)V4+",U??9
P?EQOQ] !_[E:"4SD=R7M?2D+S_9R?^<H W@9XB7ZM_]PQ$2+3$6=Z0J!&_+E =Q@
P+V3/6_X=XP?5^T\TZG\^7Y)HH3=$C[ZH37]7<9NU* M:N[>;!<A/E6K+UT?#=PW6
PB<U(%$)#ELJD:RJ*LL%D#@ 69 '&:\;<Q!3DJ ';=9@Q[-P;-74QX_I<M;#1U),C
PC_2\B4X&@3C,7_NSC,6VI=IE(6+P<>$TWO7@D>\Z&GLWD8-9>H42?M?]PYJ8!<CN
PRQ+>*53VPO OLI-L*+8I5@7JYL)^4@SQ,Q8"MP-H3TDNGX1!/,Q<*I4U0H*F@ W9
P/GCV*I4.D4!@IFSI4:[@@G;Z(Y[''^&.#%3$D&^]0A>G[@.OT7F@B8F[?\O)9#WS
PC652@NF1U-X:0I"?,7[QW7A%ZCBK/QORD>8TB)==P4(1)IA.!I=:L#6^GRJ0"."L
P8YDQF@J>@+/!P1T5K4-7J9(+8W] +KTV#H5""4HO%OZNVK%RN:%2'C&.ZS'[2#'&
PWK(A9"UU"\<SJ23IQ[NTL.X#YYZ]T!3^>7V0)OGPVI-^QL<4M:5>0MDGC678_^+$
P^^_/3+C,TKE+]*DG\SE3.0S:!X7E_2Y[%N>7RO0D],A@/[M<%9]A6C /=.''Z8UM
P@EFDH:+M.T: 4&]UY:I_\0ND4:[]IHB9;(JP(NXJ//6/Y#(MF&DC+9ENTB]DS@#Z
P".8F)>PU9?(0:QV6M?OQ($@;;NY68\2-<(Y?],Q,LUP@R$AQ!UVG9:\#O@/W63]T
P>NFL%X/KIPY@X;B-;O([?@\0<^5':4OT2(%>.DJ/T0L=+$R^X%'DQ [64!TT&L2V
PW'W3J6$/6#)RUAB;V/=$N+<M]]G\I(2$;['60*0>RFNXF+,*=@&*HWOFL?.@&;SJ
P)JV-7>*+\, K?'V]EW8KY<%/EO]=%BQYQ'O'/Y.=X9/V7+89PQE=K$)8#[[K'Y*Y
P] )-*PEGAE\TE&Z2:N<+QX'R\N/\&R3HL_290@SK\Q1=,M%1K2ZUA0F@>+T^H=JE
P_@SZ& DWX4<5"UHZX]?!A\$/U6&S8Q"7ADZC.>N]\USS;NW.))\'XO91>R[UKE&O
PD.&_F(IWM#-WLAR0<.&@N5 \,SM.DPO"D*[6!KO*GQ!$:C9EEELT9GV. OIWR !A
P0[02^,:.;QTMZ/<C(>1_+#( ,J J5&H>/TA4NO+5VCO-*CK\/AS^[EIV3GF4-FIN
PC?0J*'$#W;T%G1RNS?+AR8XDL&E$ZB@:!&0#H*]4L("D*>;F+JV\M13A-8Q[HRI6
P-6M/F,5''PUWMD8Y=B"PB63<TE4$.<'?TT4(]B[-1#6U[5*1A;$2![D>;.*&EQ>R
P3"K^&)-:E]Y>GM]MKPE()(98WX.<&X>G1O!8 :0H5/+U[.C&<?/2QM#SH_+$=';^
P3%NE#.,;\?]UJH,>X5F21%M;($W[)@I2 Q0%"@7D(CEZIGQ!1&2[8[6% <KTX3&8
PJ)5>TG0^.*[\7LIW_P!]CX< &[[N8BAB)2R_UV[<6T1$M _C5[,LIH/&+X)UMG"Y
P4WJRLOM%4K))[#C\9"1JR/;P55C1^YT4Q1(YYOHQ54\G A]408M19KF<;H^?2GC>
PYQ'^JVV4KVY[N*3?U,X&-LUD%G?/_N(+^[+!\^5H--(<.+KGAMM?\+/<@ZANSEA%
P^IK/"6.TZ?$*E F]3:%+ZE"G,,HQ KWT)+$1&7\FL7$MSUQ2U:C?@XW,=$&FH**/
PI7%OIT\"CB1B)ND6 .IROMJLI3#TM2U+1?]S+P:E_56T93]5ZSYGK,N<>@B<QU.%
PUU]5-!EAL["9&2QB76:KR92A)/Z7O!N$HH;(9):Q)[JF;W^WY+ F?G#T'CC8<['Q
PN  U>)1._$:;F$8G)9.+$>INK>ACN8;Q'_<B9E?'DA!9>V_:B\!4RT_1!]BWX>L\
P\"*#OJI,'U92R)\VU/:<4; ?]D6HY"QUI%72N-U$#\\A&IG/)4I& 9)C-+ZX[+?U
PRIYB;SO0)Y  0)ZI_SZ8'2H?L_K&9B^<[RTN'@O117?I<ZEI='XX9TEI5Q[!]U[P
P9+5U"]7/U'Q.,/[/W,*8WJO7O'>5VDA<+,X)!>.1B=BN!1T;2ZU28^]'/0&K;S"Q
PV1R=6F,)U<AH#8110(V^O68:WKW]"+-8]OOK3KP0Q:=J9D9<*,>P.XY?W(V7XU5G
P8C,N,@;PK9V4QSWW39\AN$=@9;/;,_R#4-Y37=G:8+VN%C129*="[$\N)/N55-]B
PQ/D55 Z5M=#0?JBGF3BU^,UL/V<!I4B02852^A"7G96;?A.6#!5+#P3+H?A752L,
P9!D%N\,:K<>(7F!ZN:%-+;KD@F%1"BY</0GJV2*%$P6WZM=2F]EH9\./?J$QH7J3
P1%6P^I[?P>4:SI@995V@2Z/[<*!B1'-WCJ"8":WG=W??J@WKTSUKSC@$<X_%RK,]
PY>LU?J_?%=(T:QK$PZ/5@,F0WT%,\U<T^YF$"; A%^%)*)XV\]WTB3;L3>I]M?96
PTLO41H@Q+^&8>KX-TZS*:UZ=!QL9/<;U)0'2Z=5,YI5]SYNI+U3TU(_)^AAL#:OD
P,Z*C*;?N;=^6V2BV93HY/,S.?"=$[&^R5=4'VZ)!1AB0;D9RU@G.XK!%Q;%,3>L4
P7O'4\IV(&4->\?OS>XC9J 8[<,V/V[@]0ADOX">:-Z8X/GJ9>1RL>*7-+Q(7_$WU
P&@5GJL>O6Q<3'IR4Y&PWSEH.?L1=7O?*(V85=U<@>^;.I]]DAH$FBI)3W$>.4V[V
P$^_:#K1=L7IRMN/-=I1,(N%M(O!3P!RV=<FKU])UV=C9MYLT%>"LD)K2.&9+^2:"
P0$&X3)<W4M7:5HG$U$?B5ZJ%K9EQOVWF:X:;\,5]"DU8V#G+R:#[H7-&IU&N=D,@
P_1V7PGIKW0(<-?Y]S[AX4KX91X8MZ5RGLGF$=R :HT\14K 7S/#[JOJRTL1?9)TB
P&"%*F8$0Q<]OGHYAKBNE*OMGBJVE>(.M*>0N =)@I)M'1" ;H]J5MOZAU]_6&"NX
PV_VH&+BO>Y@CA])V+!C5IL4$)C/)'#@AS9*]_NRF]5HW?,AD^%-\Q,*]RJ#JBQL@
PQJ#:&51E[/0WOF7$4BK"O&[4O*I P72P0%=G\@I^>G,PVIO0:NOU:Z>I%;CN+P2\
P0U6_W&OR_K5-FN/=VPE%<K5?$Q>O,8V5S'^)7]R?I\7KFIM,1%[N^1ZYMC^K[<T9
P6>/.V4*#:)BFJ]6"7L1L7:]-M1,RMW6B1Y1H:6.O_FK%IU83=UD2>D;@,L?E=S4C
PN""UT:RP1&@_5H \7N]_HP"2]D *&NAB_<^!XLO 92I\D;<O_C*05E3FH7R@%?HO
P R;A06U/VAYF%^"?F1CDHWGL$&O-,A:&[]0SJ'Z* Z/?%D4[)T'3/!*[DK'_7;KE
P]K4Y=HAM!GS=5$;M0MY:Z UHTK8/7?>\N='+B=%,D"*36V''@N6B7H7@(U_H*5) 
PD&[[TY:]LBA&P\I')D2V?JM/!=_+.,0TZ?4A0>6OPA&I)AIL84@R^JDX6.QJ-I:6
PHT.W218-P[M5F:<'!D_KU,/;*51L^,+[MAB7'T9T$2P5,5"!B)BSFZ * BJ3U:Q2
P%[0 <Y:,B-N+=STF?H4W([262+R>*8$AV038WSY//]0W=W!2R#=O+34TH<?U+U]_
PF9OJ_NZV;>/6PYXEM*9S.=?,+P(:<J&.3%J#8N'F+W@]\%YNFKG+QCF@L[H<U!A,
P/OQSFN-'#9NW2*0%$8F=K]$NFC474S=Z(UZR1=6VT7RX.9Z*^1)',>5(-6_6]/#$
PA:D'-ID S$P*C?\4Z6[!F:;\/^=,DI!_>#^L:+'F0BTW118=$ ,\#U)9X*%[[9[7
P8SSL#Y?L+"W#7FS._[%C-$&Q$#-,Z2O$8(1BE$'X<L^Q8]<0 '@-E==UL"R2<T32
P&2"4C80?]4 PN$POB?-[,OW4@$'W[ MH,]C^]K6',/(_#-+O#/!2.=XIUER8V83:
P1)%_T.9TZ& H/F_JS.=B/\@A.?&&AF5E[3Z4CNB7B7(,)V-8*"SG\^5;$LNQO)C7
P&/@Y:_J#/T?QYSZT6,I64Y;/K^1!@%_Z3.! ,@=G>UL@B(^E<@M?Y32Z'98U-5K1
P%"_SN-70_L:_S38=P>FV(,7/,48HLTJ7%^:RZ3(((!S;N@+&_"<GD@LOOWD%E:VL
P#2WD/I\O_"I&V6,;&"2M,CI(*,JFK!OJP*LJE;:<#M;6[Y@3:OMOQ+V%QQ:/8.5.
PX,@Y'^W5HF?+_(U[Q30\WZ+*H?Y]8UN'/>S:@ME&Z;=&L[EN[30&8J2XDKTT&$.)
PMQYX9BJ9OJ/HPR,*,GYWU&GG!G9/8&3C"'YR BED6ZXL4-5^:>;E$X90>X[Z#H.S
P=N C!\T0=[AQD,YWX0^Z!)^&F/O<9T46=0AY5&7.\EHY3G3K5Q:,R/'Q_?I$ 4C%
PC0#;:<PLEU] 7-JM9BH7*P-^9VPVWR%)YB"(ONB%"Q.Z".N\5CU;&+HGUE[=79[U
P-/W-)JJUN")_?*'G&64/CW[DNZHA:I]3;ND488")9A<5JREVLCSZDU])93^[BU$:
P\DXU_\#IL>R.Y6V_EK3\E'P..0(O<?+G-98W;9JUI(NT-QH*'BGGG)ZH/8&9:=N:
P%+"@C<4'Q49YH] QQ0S;UI5>1Q9\0OCMT.]O1(1ST:($Q]@Z<O 6  H8K&WL%3Y7
PY=8G(J/Q?$BLG(#Z 6549<LTUG]H2?S3&8[&.Z(Y][5;OAM"NW"<6$]@I6QOO!(9
PJT?@PPE[\YE%29!;I^!A]6H$)J-44VCA#Q776SG0"%W@'&:.2MG&Y5%!,XI;=X)2
P8PRR=JY<K>%V/96=0#\#Z:;P4MZN]JD>=,E?A*G_7))+ IQ)6/ZIH"5!.]D,0"^9
PJ2"J1NM<VNP]6P(/M@_G^;OL&GCQ:5>C=4 &T>"B#/1\FUK/7/,&4=9C8L%/44-5
P1:&=D7-]M)U0RU^F&T/'ZISIGE0A.MF*= BV"<"=/29<+MAHT2B!Z!73%0JJH 2R
P$_O]%S8HZ(*C@<TYT<"?/ZSU5-EBZ,U/0K/:(E_D:.VCYGC\J"#R^M1_8GZMAZ#R
PZ+R3:^)A";[M00<%D3^LV6<4Z!,V1O>MN;P0__ WRJ<^K*.#"/H*%P(:@Y=K&M>B
P;5 )3!1IXO\3"HG_G3^=__"(&7J=AJP)',N+9(?)^H%F+]+M,SAMC@_A.:2:A7/.
P965/93W*48Y*U[HHQ!7U3TB-_1,C:%2/-48P]#B(^(&A;,8?!XM&&V?NY#][&@?+
PBAS>Q'S4,SU^G,8:O]R+Q5YO>64Y/_#M?7$V<#PPNP024=[PR_^#><L9I?*/R#@>
PVS#/\9".A>T2%")+%E#S48\/EU 2_RZA/=RHMU59R]/- 'ZD,IN2#A&\(U_I+.K4
P?R-!:Y[&JZI/PJ#CGML@FMY?&LC(4.@VIK43NJ6]6%N_3C^[*3!=9^I9RIJ":J'Z
P8%(W+ JJ0BF+%87>)7(K0RI=]N69FGS;E'75/(LG^;N&K!FM6-W_S8^4)2+4C==J
P[[ES0@D1B\\.Y5 A4\K(W51@A&N78?3*($=:.O\-+LV%IC4>D]$>?]HG17Y_U4V;
PW-YQP)[K[2@Q90VJB7!T^I_IJ.'KN%=(X$("WZJ0\&%C+PBL'I50*=\+C %K=Q!I
P!MUQTLL<].SK6N4N*)V69_^^1>N8\DS:N$%, R3"&G:H-I,-JD2FO4IQ(USLXEMB
P/IIQ%[6<,BU>E0P0S,EG.EC2 3+?42*P52%/ZXNH"7%CK6F-0/@;S8EU"F!VY=2Q
P;I:ZZ-.7/7^!I*\';N27X7,Y$$(C>9'LQA!X'/>"P3XGV'Y6R?1LWXV7N1EN^>WT
PK#F^O%6CL,-<#8@>$I8,*H4?900Q]ZG_MJ 85H(33"H@Q5@)3_'3,K6"TI\H5CZG
PG9;N*)'E4@)<W/,U/=Z*6*\=$TU^9[L*+N8"UFM+VX;5K,=?4V<%?7C"4?<WMW0H
P&8YBC_?AEQV#C4K=E)9@Z\F9C6NBC^)+%7;_!,6=#2PO5:HS)I!@JH>>>^9),EIQ
P#PZP#'IGID)=?)^;C'&E22+@P5F5=H48EJ;Z6H[P4=SO;\Q^LBF-.&.2"^S)A^DZ
PX;3/%"0D7X]@IP2&!?[:,$<U($%LGUP =*>,&%IZ;2GN91Q;O# V:D]*.S&W?#!-
PGLRO6B;-.26#U7>D/!>"4B/A^UOE;A!"4*%3X$A;U@";V)9#<4-OW"U#QVK[F @ 
P4-B>GS[GVN4V1I&[7,P]8D$(('%+[OEJCGU%$VF=:T(?,HA,@#'.EG#K]^U(4<"P
P6VHB-?E$TV#]2[A)Z  [#,D?/F):8@-?[L;6-84NZ]U_U.BG3J9.N%2NN1*TX4>T
P36S"/H- ??9K[0^ Y__4!DRMR$)@DH5M,<&2# 6\XY#,OSCVC@>69.%SD$R/C_G!
PI39A@3OC=:F61^Z7%;I)Y+LR"+K 4%$]<V-=+V#+V2>G\W=KB8BQ)V_-T0]M/2?,
PA,D]3MK0( O*K:]25Z #5-6P0\@7:#>1&EY@$A-U1>Q!IBV=]GD[LPCN-$S=T.2X
P46%/*75?AE4%=)RY(#+,CHB%V3J7H!N@K!K?5J^+8=\&_QT2-=[KG1 ZQC !TEK 
P3JB9)1]J\H$[JBX1_,8&"\?AEP(KK_R@11GA#&<YE*#EBE-;NED=0;L>Z_1\ GWS
P:V^)]Q@'^NA>J@.OJ0,9QQK8]L@=9;?QJ4K8A=EJLH;:5_PCFFTI^^04DC.R)6?#
PO](=%);/A7'& -7<UZN:8SR/_@O(R<D\%! SZ2P\8+\4&.#D#[:5UEPM^;O#QP4;
PJCJOD=!D-6@> =/_Y6,:1QT:)?6S%8[4N:8R:8U50O_%IXOJ!IX"NLU"OC<_T"81
P"3F-;#I<)6.$,5KPZ597TK=&\H>6$A1@L]QS:GSW5K^@=SW%(L6>>NR3T.RH/#@S
P#W3*8$76=V7<J8C <?A!@C*J8L<DZAL9.DWG 3:^+]RP[M,:0O2GZ5"<&,1FEJD*
PY.O#QZ\ L'F"#RD0\4K%%ZR7$F9C!^^?'M?C1(7;/^+![VNNNL\U=DN;T"NJ_#%Q
PZ+MW=#LX@?]XM-?JR.E#,I-51H8MBS_F_^K93.E4RZU+&??2N^4P!*NAO7IR3=8M
P6\PB*\2_;-]+G\*ZCCBB9ND^OX:D."(<@1865146GMD[=$I5HC-X CH2/0#!7,@&
POM/<>1,!&$#?0U.$Z MV'HB)HRE((%GBL^3HX_#D(34]Z^UY*)7ADJ6-$J4))B>.
P(O$,ZJ"E(MB*I82Z9$F>R?UW5L)&97,&8=[TP5C'?NRW=W2E?XFPE!!I&!P(3@2&
P8EX2N+"EPH:/L]R_Y0PJA)_/]ED OZ<J6B_RQ.30<S9'E1*$RY_@Q'X^WX3RBY1^
PS!$,U N$ >6CGC0S/V=P*GT32;";^N)+$QTKH+;@2 0_H@C);\E*C@.7.LQXN*"^
PE=R1-RM=F'/*\8Y]83D>M:%05*\_IMDFYF64CK.[*9*KF^^P<F HZHWO:%@_M&*>
PLB1)B:<'V.%XS,;F,&A"[V48-/[1,5"^GT(,XB3/N'4#NYKR7<G)==A_,<]V/#"*
P2?PXBV<CME_.1PN[^(#P@M%1/IZ**8R5^@&B] 3CNDY.0%[(HTEC0>&<?1+[RF:J
P #W"@<9=9)W'=-'USW_*7N5!TF\\?"^1EW4;5U9ZP=1-IH^Q2-X"R/&Y+%!53CWS
P$&3EUE0P@.7J&#C,M#.V%0MO[HED"-#F+P@WMG#-QY=^6F7W_'YIOG ;L+8%"\8L
PM\CHC3B%8Z5+]4'U+9O"%6BP04/_O[%F6 1GY DHM^SD%?J,,SKDI2R9:AN7._;A
P_W/5NGN"2J,G^X9.==+&..QJ/Y6V/S@%%3^\7>PW>O5J<WS*#@JU0?N@SLDFKX?,
PJ EEF4N$][U0 &U4$\[ST"^L[DT3)8XU2YO@9IN?2LHX6AQV?T!2-EUYZL!0,I<O
P7+*URJQ!AB<;0S9SY*S9==%:# W%I _5S\RL10.J-I+*!?L;OP" [ W+ +CI:2Y>
P?$Q*>*K>F9A/;U*=FEOEB7]HC3A9B774KO/T-25IGG$CZU(R>UXFW4%C*$XQA^02
P0#R4N1:C=*N+PG[/0?)&&)F>&<Z;_Z+*[*R&9X>H4#R D5JK T SF<D<?W<U'[OY
P06SQ+LBFPI#=9_,INY7"DWL!P<I.B_JM(@N2]0WJ!H"],E('&:2"+SAZ6451J0/V
P6HHM[!D@1>B8-LZFCM(5SX]TUB<E".MT7]Q@Q9,#Z@N$.(!S)QOF9B^F=+9J7=_2
PU'W:6M-A5R$/+[,/AR]D<98N'M"W_LFNZ)G/=[SC&2R<QIEQ0H1#HO5)(]Z0J&$?
P2Y%,+T7J[1@E%\*Q6-@C1.7;.Z%4&5>]%3)$TG3]V/)311 [!?;.VY+"4AW.\TP 
P2:UMOJ#BN*-[E4MYFD ,RSZF+H29XJB6F:%67K>K\E#'A1HNFT5Q:5-@@.A_3H2'
P6<'[PM^X#/X<*7\3'[#\G5E",IC $^-.:0HZDOV16]Z H60[SXZ2MIWIVO;:RH=D
P1&Q[-@J#RYQ,8$9',6+?5Z5_U)1:A \2*14/U9S9]IO/,7-1U<#%?Y<P"(H]+P7\
P%ZL^.6?+/6^90>B>5"6+:@E%4&CY'FT_8@B0%&\E*XE.>!L+:%64G>PE.R=?$^1>
P)DF<:U"I T (+H_6T8OIK_FYY^@5U'3GM=K1)O6JO10_ A(;QU8!YPGPX;,NY/R4
PUKZJ>TT,I":B%=?LED:_\=IT17CQ@VW6S319:O9/>8=0?"):?1I^-C95*W[=W9(E
P" >GJ[%X[O9L[RV@>8-;%U4!.V^\2^N=K=-$7KA GZ2$_\@;V;_&),-UJ9I]XBSF
P*^RA7F^::^.#147EY-IZ:<2>:;F+<\KY[%SUJ(TY;=,+)C?:T-(7.?)ZY-;.(O'L
PYK'DQ?4R#-[7<V(77J0+45E+/^U#JA0\@F5^RD#<?4L8H*C!! ]EP%#:,2 <DK?O
PW* 3W<0S]HYSQT;6^;6=\ 8HH $2!0W6K69U<4OU/5[O>AM-ZK?*YY+QV>$ERWPF
PRJO*Z_/1!3M!F48#MLGC3MC4*#4V\PJ@G2M!37NP&L]?"DW\R#1E>L$Q7=^4G=".
P[X7"_!$["N0PQ[D\?;#O>IIMFMUC,D]M_CY*3?.*@/*I6EH49LRREHRO,:C8"'(M
P!/O%Z$W?N[80\ZQ,)MIBVP._I>9*U6N"#V M#->%["ECX_M7@PIU(^F!^6KD?/KD
P#Y@E-A%P@CVS=89D7.90^6Y;5]<D!X.,>2-'K0+ZS5]9 1>E'!PY('*T]1()ZZ>-
PW>"M1MXZ_I2;CI5F?MD8.NOH7XQ9JPX!_N5ZT.JCT-?_CI*,8QPUP/9VS/Z(=@!9
P$:(CJ.0%I!WB$@-U!@__<%_PT34].*P8ECEL08M$CGPY[2A-:#.2<OQZ@S=$7-4"
P^/QO.?PMH\_KT/JQW^9#Y!1>B+(;.&*-I\;=$C=;@IV_@ZO22U>/4\)1^V^(!:#$
P'Q[;*?K:YTO^].JRA1CC:,(<O&CJSHZ6OXR#+H2$XV\0)#F]"KN@>@@K&'9P4\[$
P/J^-9G%4P#4R=6,@>,VA;'08I .Y"-SK;67YLRPR4UXJ5X9"HI1G7K=:A$27WZM8
P$Y@NFAA/N>J(TU>67H'N'0QZ$6R\X\'9FB?,U,2K0)-,#VI>Y2'US\+(>ZP582L:
PA](87KP-W.L&L"D#^VM] (1@ Z_JA:]=+=1PICCV2F6BI.YA[3FA1[\)]*B$L?F(
PK?NAV=*;M#]7VRROLS27L%Y?*6 10(RR:3;Z ;N$&K7Q 3HSY .]&5^O_K!L6$+=
P1=1Y*%PNNJ&\6)B=ZN[ZCH-5YCZ+7DH<3G*=\$!%+MN9"/[ONK"6WP,DKV*!>[:Q
PQ9(H+O+AI*Q&#)W-:1$#046@,!3D="C]Y152CX6;E<<>S"X(;I_OUS[GH>;%+H<(
PHWP>3RYN9MJJ2M)()J?NHVL^@[?O#?_M<1(/K'ZU@Y+T$@Y-"3>_G$BE&MO@;-9\
P]O#1=A#_*?V)&* 64BIF:'3F>_Q%?@*"V/T?W*^I4ZQUN8*/<&-3<S#&#KOT/0J-
P^"ZX)3N+&+J>-(J,&1*(XMKH;5)5@GXL9*,(T]-AQ&=49;) L)(RT@L:YD5 4$F2
P8UB+4E0VJVEC7]I#":?._WLI67T&OT,L*D(93Q(8")T!+XQ;K(M2XGT>ON/%7*G.
PWA,#H?8BS'+1JFRAKU^X-<V"@(V&@'Q^_75Q#:B[-:$W^Y6!V8%R@9]%1*=-&#-9
P_+Y<G&;JI0;4AMG2J6ZK+GI&[*8> &,>@/?;7QB +IJR<SDI=-\Q/;B1PP^O12&@
PN]M,-:&GV LN=*)F"#I"/H]/-N]T?8!?\H.:D&08<<5,C1 O!08%5=WF!ZCSVN%&
PI;;:?-0'&%,90F\87T%A;-=OKG:F<S'Y7<''#B+'0D6HZX/8@6!OP=C7$PYLGRX7
P^S'R\U5S$5JN?N,(!T;[21P$R%0[362%Y/L6-RC+&TU;5<Y]\7TG0Y%IX;5_6V*!
P(*@A^]LSUN-L(ND!OOH;+D$M\^N\>6O2X#<(CZ,U]U4VR+ZXPG064MAHY/@,<,,=
PJ(4^:8;"\A88R[5;#1P$&]%A]/!0(+QG,U\F_T#O6^7:@OOI]5O>YDH*] B\AP;X
PY;6U[LHHO=7(>[0+6&7S<H;[844'*[4D)2/) V]A:ON;S&KJ;@\>?4)0!C<%A[<,
P7Y(ULS?_!?D/.W/'WO>T-%4E!2\71JP$NXUN02HD4"KS& :!S6%UH(21A_X(^ ,<
P=C,)XR[3$]ZWYYU38;E0_YQF$V/K.-)>R3?Y\6AJ_+^>D?2[E1*/W&C.J6CO]$7$
P^ISK US-6$&B??X%'969\<,3?&>SJ*A>N+\,J9L/_QRI_+5Z<[&1VRR) S'J;ZLY
PJ"T+T#<V!<_')JZE<)R/T-!9[+@#A8]_XQ(WB.D?SY(C_1C@62LM>/[@J!E@TI:6
P3 57))N E>!GJ%DU>8,1B+1YY%F0(0Z<X(>W:&5S^F(''AT .%O3W3DI"KT:I!:L
P=UD:WG 3%6QY]Y$>/=4.9//?-R\L,?SG"SA>;>X7+^1$N!BP\/'DY#L%>K[J1;T:
P49]0R3?._U^-@)RJ-[*<<B\>YZ)+0]!R7"\:1W:F_W(SL&/SM<S]D@R V+=\*.+P
P.4IO=WZ#3'\V),SD^6!?,^/7X0V&U(3\X$X)4JE-SD!@0)V!028@KY796O"O9G3%
PIU+D=)<MEXUW6"+'&9WV*@?HO=%&'@WWB\H'KU^5^/_I.,PUKTX;APG^90.]?X%D
PR9$=\TY78FT6R(I@1<L$=!U@[**MA?42@5Y9) KBX"4(A^X&KV!8'R^4P1S$C#O 
P&GM6QUX^/P''9-Z0T/%GLP-)@O8L**_D9XFV2IT('NF.44?6ZEISTQ@%(KR[=1[2
PM)X_\I%[>UAW&>/\%A:+9A<:-+E9ZU6P03T2KM<BD2FFJ,NHPVG6_.B8#V@+\Z,N
PI>I.3OST5\W"4JR?/9)LP#73AB1IZ*6;R1@;RY'7S"Q;X^GV07X7O$(!:$Y:1,(,
P*?3@O6:V='6"]N>D6<[* [OEE'WDP)4"^*-=+?7 =6H+4/F81\<]'<,(D7QK$8A#
P+&DOW8V,EL;\.C8@(O OY0RZ W(GO-Q"_I^^IPF(UE-A#@)8%HNR!2S'^N<HPQ;A
PLZSX4NK#$G)46#HG_W&%L\7813G+[)3=:O^'@4@OEUW?4N[ ZO%&?0I"E;58.@^E
P\&:ULHO$[(%;)S; 2/_+_IINAT:YSYN$<KO ?M9F]^\O38 .WU6D: 2MU^7TB)%D
PF[33@[DSIQ+7*]R+Z=VR2MEWQ/LZ*6)&S"-"P6A8$TAKX0#0!L(I="Z:H%=B$B[)
PTCL2G4JY?4?WI'/4-ZFK-EX)WM0HX?T9>S*6=*URGVT4@[_1J&)?5"@M\K"C6S-Z
PI" P-\"<%1X#1-F'M0Q.8D*?6@WU1=AQC $]3@J6Q1M6 4#*Y/3BC[:@ZO0_.A#*
P* P'"":!@7<LUZKULPSY[-2#MK),158F\0ES<4G46V;O]VL-N1=A*2D3'B$2\+UP
P\Y[YAA@MO1O-0!C,6BNSK5/N7K14_RHQ3(7CTGHOS,*@;H*+.[(!V(D:#9^Q3Q 3
PC=4=(8/^W0J!#:0OIA1IZJV87'KDA J5'KB (-60U+A*A X782GL50*@VDGT7S"P
PJZ4!4,!2(VD4+_R]L5>1XC@CFPJF^*ZC:R2_HS+.?TMB_USYX4N@][T/V2>7W;0-
P%/X3Y$Q#<P<)%0DW^'EF_\L,.0)+!A\KOC]%0)ZM8YXBD<S?,Z >OD*C>A1'4RSD
PK+AV3NOKG/]$:C.(O%0'JIN^@RZ^BB#'2MD!<A7C"RX #S%4/+7HA@#C*=2F:SWP
PVJ3='A+OX !?6K\;<WG*<"GO8;K:VV3Y'=UUU;>L7R^F1I8^T">/AYX_XWWHQ986
P!J9'K<^9,@[;A^# =C47O:&C % Z#=>S>W*OU'5_2C$U9,(-/L"_-ETH+Z^@0+5T
P$;?/TC@B!$K)4&X33_6W8PG<C.YF_++INN8AK#_;\_Z>G]_R#*\1.\SY=U,K\D3^
PM*Q=.GQH>#"6.O?+BG/#P+$Z]][08S14@5RX><ZL?5($0+7[)#/$=:]]YCYC.2TP
P+54E#W@M<@6M020@E!L@Y69\6S-#Z[UNTCS1G$JQ*"\O+,HMGXR^O ,7^(#C#63(
PWB[_ %N0!YZD^.@.;4RDA-C&;0)=HDJ8],W@Q5T5,7F_C>[5CNS77AWN4#^6[I2:
PS0;Z-*C$KBT8=,53_)H*0I!Y=>*9IX-"U(K.YG/Z-_AUZ<>FDG%LLY;S-?I="I=3
P*@0>0,!BK)H>(IP# .+HFV7=P58PJ:Q31"TSMK/5&]AQS*@Q:O>U=-70WGI"993,
P]'\@4^R)?!(Y-#="J8(/1$O\8(4;('EV@6 'O?_*ICFMZMJ57/P0AIA@$AEO+''M
P4UP6?H^&V/.A<(<M88G&$<('JAIVO>X7M*![Q!^4LO$WI$=B&Y8VHI,Z.C3KSL5/
PN,0!EU[LA\'7^&_7YV*9XQ">IZBE.=,L["OH;_8:5&2'VN9>+\Y(8G6,_30%0><B
PA-VD8-YH_F=!I:S=^<T G&D].:,_\MCPW0?$\BFL^"OZZ5?/.TOHMRM' _R\K[]Q
P1![\T94H,DYA-H9,M>)N]PK?G%O?)$'7=;X&Y)23W+X@H_Z;*%T',4,7P(2W/L 3
P)'\[)B?.?]#O$,S+.=6M7$>-R "-+TJEBDF6UJ),936'L&T'FTWV\SP$W?R6$W!$
P.&N:6LZK17H>NV6]T62@.F=U.Z#83+05$?VGT\^7.!BG"&"'HJ0GS\R[P*S.8:PG
P:M[N3F??( 0^]L/N.!R5U,!'<Z(X$J=*X7(OY'AH7=$;W8JJ*:MAJJZ)V&P]"$X5
P&W' KKHZ 7X5?0!  *VF(#;1]//#JAV\;FOJ\VDM>O!MX@Y+"V^QY%:ZZ)YBBH:'
PX[.5BD6HOC<G)#N9HZ<OVFA'$CQ>WNVP4(%N^+Y:^Z?P.U#H3J92*UFJS56W'$+\
PL-W8<2]_Q4NT ,/>=-XE0*PCCS@KFWJ=PK,1R=A)O\B$AGI!@Z*OAH"=[!\R ://
PL0.$ HF[57, T#Q2<Y[6*U54U*M$H.]"74.Z\HYO=@.9(-WB<Z1NE!>)3#@GW;VX
P'$)P9,E(?.P@5]DP5SZ,#3+I02Q*/X89KU[[I/6OQ-V%P)H5 JSW2<1,4@OTE:7<
P#NZDA/!ORD6P2&!_RH X8Y*UMH2)FXF\4=JU>"@W90 =;A*FL^L 3-(KG]&BI+3R
PG",!?P#7?G6JQD:%L+9=D"T?WZH9G/R_OC="-FCUN+MD?9#!)!HH74DE 5XUO9G-
PX@RUEC,K;O5GA#2%G!M.)HCYY*2Q!ES@U!&_@(B*IT$-DR\$ *]A^[-^O?1JR<I;
P5(\<A-'63?KN:B^PB>Z+&R^J_1)%T='D2AUFSX2<?3?70*;UTBG>V$(8FW*[9\:+
PK55^B.I7RAZ92X_$GB'7PMJ>DN5)]FV9 H*7+Y3FS#>$U&IH+KBL&_:+B8+#T]XZ
P-N6HD:G_VMKJ9-L<3?Z:[RJXHB\Q=J0;EFNSE'$"5"J:2 I%KCX$AL"MX(>\8F*X
P ,3'"^*'H3A$:R8'C5V*4?2H,/O!?XW((L/6YJ2AREJ,(=QI9[ZFOS'X.[MN+SRN
P?T!O*9$Q) 6T,$CS6@]Y+,9I\QY$5]A/7Z71>(*@<.T66"U8D-:]FG-0EH2A/.I!
P7F1H">&3-5RX\DYYL:^U9'?C*>ZN_08GB(SSV]$2:((\<'.30ANNS"PV"D_OKK;T
P0"](27>ECU[7-S4U^%M+U>+NT(Y#C7/9=!X63YD%&Z*H.LU>@*AB5 ;)QX""LSV8
P-.,GQ1*7KS^U\'1#GS4H+!7US/62;7_\H<9GDT;)0 %U;,N?#C;]+V-5Q+MN.X*-
PH#A G^F(1<&[ P6SG]_1&U>&(>Q^DW"N^T?4/<4O8*]Q^;)!8X4(E+F_G,\>KU@M
P'"4$M:LT"F*V8V4ZT^1-("QB.#W1=6#GC X@//:QF&7"F0/(Y1CT>:2;B'/,W)WY
PAJ'@(K'^!:W0"2*""+ZWV89K>.WX*S<X0[$%DS^"_B9DQ0Q,*7+V%Z/D-C!H3^''
P4]]V1O=X:S,,P6BT'.&BMFD9BUBU/K:S-]/?X.MM:Z@^^)HD?.""Z%@QF_5'3J&_
P)[5NAJ7<S@%2-;SX+W&,$7[N])H:R2/DUC(YWY7V\I@@(=5[7U.0KU^7R4ZL&7B!
P&-#>.H-\LHA3*Y_L&"#9KHJ=GS(IT'?44H=_= K OI_P@NU!;D7DBX%IF-LS>PBR
PN\EO7'T#AE ]CR "VPE,LW]&;F"3%)%'588D@0_V'DNID3"^O12A&(1N-[^E646X
PU^A+9XWW#I(/9JB7UU/'S#6%/6TS$LI >,S*P'QS^$7=P3,\V2%@(N/3_^!?VO4+
P^8?O.PCTY_!>X/0356$GZS-&PNI1IEC@@T_(W6IW/8.GX/ S4\\]?*:SK4J\OH?W
PO?0\>]*\&=2M$W7ZF]A=LJ7,:JL3[4-4Z#Y:(!^0X%I1F)EA#Q:HP1,+J*" G]SB
PD@:"V$8U@3N):!N&W6H#(354CS#(+24WU^W!!W#C)>[QF$ LI,^?@VZ#W)PE3P#A
P#]35&^S>H9IF7ZR0.J 4+Z8I(Y6PK\'>LBK&^O/!+S>L+>2QO+3 W3DOB2JV5/Q,
P/)$9WN6; 3FFGA"C.;I>#<9H/P/$!G,/"]C9P@'6U2W>$W=9E3:\?"8],]1%X0LH
P,] N'K-C(>MMEA9VQ:BR.GM61KFJ&D1 KSQ#,O";%>7<EH(NAG'*\KI\/Y9W'@K?
P)R&4[+ =!=!PF(+T#8K!A(87<P((G?:?B^*X7*^I'UX4?L,:X8GZWRS*^)!;/XJ 
PM*F!5TS^0!CX[K@=?S,]Y8S^?O'@]6+&NPEQKI"9H];.T0&WUR;J.L@_*X+'QE1Z
P89L&+7O4ZK=!Q?R?>[ 74*6S\#35QDJTFW[ZQNF &1LT*#W&-HU95;K)8NZ]7>Q0
PY&+8K6MP/%GCP<H=GM*AX.;7)&$>;&GD492AW+&C_NX:#F5EQ/Z9^MT6BYDD(GHC
P^&%O,^YS#O/Z8G\3 IX/!Z7?4-4)5"#W ?H])2:#2_L+X-C.\.)1(>$3D\N:,SRD
PG1ZZ^L=2TGR"9U0.,3,$\P R*(X*_08LB3YJ;H<$Y0MZLT(C$EP-S!/,4O6M!E]@
P40[HR?$4=MU?8'_'8_?XH$ .84 P-O@U$=!"M493[H!3EE)' F\[0Z\NR+Y&GR,8
P-"4Z\#C6NG^SQ!6_0L37HY3*"F.+[YSZ)SM^*TBO;9X)*%BU<,=QZ>>+:<E%+?[Y
PK<5A[E-1(L0[H[K%6+):'XNWO(;X<@E@!_?7L2WX8-"T@\FSN$-63R/L54.CI^H,
P>+I" &[SXXSDRGI0R2KALNJT>2.S9P8?==^8+'7I=99"6S$OO$ VSL?W$;1_E5F4
PR1)7UO^EB'F5HKR>&+ 8Q*,AJN&I6'D$YDCG[Y]H]&T)I*4_XT+BG!ZB4[5+Y=HA
PYP6ZT_)R66$YG&$$%F))"=8&.Z=V!;FA&>\AMNPN64N6O^K!\N(X?^>FC_$Y3CQ4
PUVVFV>ALBKKD"DM[OP('"\^I(^ZPC5*6&.^FB&JLO M+@/SP?R^SRW*H73F5_5H(
P4W1N%;_0ABS:P=R]\^*U2U=UUT?3HZM]3]$+U/.^7@LOE&6YVEI_"1+,;R]3F!>G
PTC<=U>(V+UU7Z2%7S4(N*)^H8')3 $7$>_OWT&N 3 5J57R.?=UG>03;,>AJ-X5=
P^IJOQ>Y"0(>!^H..U-0J//UV^K/Y2KU$HBT/5N!\6><J6NGO[/$M5\?DP20#_#%6
P [LFYX!_1KEUOQ]=P/&*LER[]^%[[?Q"'Q?J)6P3CQ?8)RBR&C[Y =1*TD*\:RIJ
P8' (PQ*?87CC=:1OM$;P"MVDI*.;9S(<Y+]J9>E0D6)J(<N&G$*IM:,?:UY7OP;_
P?%'6VQ!%/< 0)NB/WJN #\K9PJ-\<K7BM-9#X8\;$_$P?(DBOTUWR2*>TT4]SGG-
P:H&Q(F&XFEAO3+%LG9&SO,8%;P$<7WI"V[.WES<Q"XF(IQ.C8<T(SJ'["-Y5BRX'
PU1#9 B,,1CP$58'L7=68MH"9-&20\8F_O E,@6+GN@*V9J(+:G$[@@)LN,UAD!<(
PW.]TF?:@Y50_T-JF,#.9J\<<:.34)!!71R R29\PJRJNYDA8Z#Z^^JU!TL\='0X6
P9SS:!K]\-X29/+09#=@FAHQZARG-Q*G7R>YBC[*1Y[+)Q+(\\!,Q(3'7?(](O+_(
P_ZQ0.VHQ#\#$A'2HD 4=7JECE9)@TH1YM@43C!]8$E\#":*-]1)#&])A.M>AK',H
PW:_C%GY/G-/<(U6>'DO?1"C0'7Z\1*W)J?:&E6G#3[ND)D=.K0%";"MO+0 U-^$T
P18XILX6Q7Z@N94^0(_3TL34#3+*E1M4"_412A]6=Q'BEL_S8&/W.$2>+@@E'QBP7
P_&_X&#",UB^LNWDU<MR'[SL?G]0:TO#1,Y_)%;7J-RJ/\-<.W_.GX]DA!*B94]\?
P0*_?^KE@@@^W&P_]]3YO8)4ZEM02@=3[+HE\5; L(^2KU2D5 E&^5$.%"L^UK$\P
PB39P-/MACIM=BXDJZ>* *?VN'A+J1H;[\H.XB*EWUA@EWA'Q35W-JHJ]P<E6'67<
P*6GV,'()&W[5(%I*950T#^.R-?4_EZB\,JW[T7@XU$Z'UFW'9AN<\SL!?4V\T_NP
PG:T:?F@6/(PT\Q,Q9$Q)?019->ND7RCJ:",EW.5@]7UE,M@T@1TF#!0OA"FS\3V'
P> +[LL((?I NZ+EZ BFR+PA^XQSZ"%^/S;CWL=G1&24W/D5FY-2FUP0=YV[S_;(0
PL7ZHQ$_^7%UP5TP4DBI9_RA#S9#]<^(WS07FO?0\C(YQ\#*W*Z@;'7$_! #8FS2I
PR;>C%4NJ1Z:NA;B[C5R!L"\C9/AR2(M^9AVA0NPP[1DKW:U$V1HG47-.8LJ608P3
P#%M*_*PIZVH.)ZE8_PHFN-M4$>A6AUZK#\AZT;E0!9*M!)X\)OF=SNPP@TISP(%@
P4M]3E"W:Q8)D1"L:UU; V-)5_3A#TS?<.'NW\IC'?^H@OT7ICYCGK-)1*3 F_,K+
P+:9+BL%(!  5MELS[OB9"Q%Q:U$<W^+-=H9AT&$_(CBLI&\<]K \D*NPAD '?S4#
P7/YI'MU.0@C&(;.Q5%UK&LC>[V1XYY(\F'16?4603721SO(1GP+[5%#;[:TQ527^
P-!I*XFLFH+\@,TN1'8=2-EZP:ELZM5RL]<*F^/PZW(X];+XQI6D" C">%/PA5S,8
P(O]K2A%E4)G>,MY<,15)9BJ*+Z%. K ^.;N+!Q 2-+B'">!0H ;=WPVET\*,2[8E
P^:,*1 %9NO$T39S^AO"M3I"@/W(-$?!4*-F93K,B_'*]^DG<BN'RGN.4>!U^[;@H
PM;)Z]?S(Y(*LR;&$US*A5MJEO [R>Z$I&6 *YVFJ:\8H279_NEE!4:!D3TK$!'>B
P9,%6^R7&2"[WP@S6#6L.1"\9^)2U%@<_"WU?S)A<B#,3MJC1X2(L'C5XAV3K#6S_
P2$U!OH5\63N/<\MP$5T&T\ --,KON2AC'Z ;F[_EM;S1$T"<B T8<)C  BME/>'E
P%9QDA9P/<UZ+6!,67/2KD,!MC<8C4X"N4(6J5,<S58H*5:VY[.]&%L77W$.@_]!,
P([4E)X!*/,I^^W\"W@#93?E*>ZBE6\9+]KN')I/6%MQ(0R3-2FG=IFD/1"7>JX6N
P^8;N8UH+&HT%-XQ=<B4B=QHD60TL?\4$?31^IR$+5"XU[P?"F#+4WLB2%I(O+<>@
PDV;\G2>;/4/:L;S PX04=4\4QTK$X="$N,P2]YIIMZXS'""8A$U-V-^WZ1!P[@J2
P79.@=Z.-+"/1<]\R.HQ"0#>[NKN5@SC^$JUZG]R++D09A-QF;U?,B"MXY83"+'#W
P)X8Q**R;L->QOCP(L03G,\#BO2ZW9NE$+?OR:X#E<L=L,9K= >B3]=450(B(S\./
PXP);/E#A)(X?G)2%7'JAEEYOCF*@*N9AJ=."-5'1BI?IK.BJ:I8^:+0DA?;N_Y3Z
PM^3[[0EWE5%4JM)"%(<V>^BLTN[?Z1VK.2J1ZH<*+65PU9:TA*K$LA)J>0V;':UL
P#67GYMB:'\#?#06N%SYB[.]SE20?PYZ#C&:=QWU<-\=9U 1/CJ-?"GOU'BR2),9+
P7CH*-"33O6(:HWA6Z89Z@X2]![+=^(CFY!&]^^D<?)EC?,&"#V;A7"GY%T-*& =S
P@NS\^+[J1BS:D+[65&7>ZBH3@V(W<IK*2_:.83C8KPH.?R1'0AH[(,Z3H*?+[U",
P[39'FE,)[JCU5@@ MFY3LY*OA;'I=,2'X,D4-Z.C@\V]2:\312^50*!?6/UB 2+O
P<%K(1)9<9 V*VU_-D]C-LW=S/Y-N$0WFI<JZ?^FSJT2CC.(VXJX;)@67=$O,JE;"
P)O/V"D]'1+%SG5!0MC=/DLX#7Y-->!P",G(G_I0^%9\X(: /(*D'?7D!Z& ^+C%W
P(8+F8*'=7K6[+?GP/<]OAJ(Z[,7RWI)^A3&[!AI@#9M,<9'X*!>NQ,U\!P(I-\.7
PZ2FHAOB.TWCJ:;S;<!Q\DCPG%0=?VY.8X?NG3X&%TP.-P *;K>1H]!Y,$J,8E-"7
PS:*?LA$< #'048X#+Y$!^SQ_I<E+R(\[9?S%F)*U\]I<>>G!$J[2YH-TPN7JWD@;
P8J[MT\^4WP.-3/2::Y+*)1-4'#0,-+LJA8\V^S#F+*YW_?UAF$OG594:*](@MX^6
PE:K^ NBQT%6JD1414,)Z/OI1A:.T4/EER?E8?';, V%0:![)8\J6F,!(CA8A^4W=
PIU52]Q+R%%*R!0IRR?3FB(^&/,*)4W9G+5KAA1?R4^:&325SS98XS(:Y)&!<-GI-
P*$4QMK"?-7T*I"CQZ7&T!&A69<&#G3Z&HFZ*]=T#,&"0GNJEB=W08#RY?PFYC6"-
PJ.:6VS:_7)4+IL $)$)&\PFAP_2/V/?_1T[ \JV#0!!?5A^MB>QOZ1Q'=J!VL=NN
P:V#9G-&7<V6;=@.XYD5!HA#E6E9[/I%PK8W?F8?6P\AK+LT1=K)'N)=F2R2.T68R
P2VIG?MFU_".1_RZYIAMKYV;@1GSH]YL;54KMJPB#K[VL ^GK (C8M!"02':5.T?@
P)\? WVTN,^DME<' 87Q.YAVP;[1@ANJT)T]:34WX JGB6LRT'2$'.'8T2G53:E6G
PX4K+VC]F%6_7T5=?O\-?Q8YY5ZKHY<+]!L:N4]FJ>>Q'^^9!M=]DE(V#1"!Z2^B0
PM.0TY4XH#7+ H@;T?"0/.N*VQ7[H&;"/:V#3#T^@U?]HYO)>< ^_E;(6/QF@HX*S
PL_WZ'0RVO&O-;.2@3Q!.*?I3(8F2&>J=&C_8_*2_UD\\YPQ:E-DS?)'9XHY78MM)
PQ+K/6A/0.5"Q3>P^%!<CY'U\W5+;J7)&E'D 8H+=+F2;8\"7A!7\M>82M>=ZGC[S
PY<.>4DG[SB]1Q "=>W:/G0?6%U.^N?D $C7^[)-E0.ZR48E* ('%?H+@Q!FXE?P8
PL,'?1)P[;?_!!8^R,0['T/V )YH,F"(/D)RD;,@45.$5^*M&!8%^IVIK#R.M9HM^
P(*$X&J\6^U!I*.I2'C29P^7(0BUD"EC2!GYEUHH.D>2E\UM>OV4X/"JI.YF[_$CP
P<MM<)MJTXN_EN=E=5_0$*K#L8%/HE%4U(YK*%Y*;PZLN8HI5?Z>FXY$*&RG@N)(/
PP._4(J+.\9N#/.V*:ZVR79CAP9&5O%4('S/:#@*+M4$NGN)&E;MDPF",H+ZG#:CS
PB(V*9SWL!>3LG$2*(,-P*=&W1WH\I'=\1,Y2\.@*1#TC]BU[_HZ=]U>B9.6&9;2@
PHH,[F>]8&#"1V( /;,/A"H<W^QA(+'DKZ*QOE#,#I?"L"J&(MIR]S%L*;8+#;(H"
P6Q&"*#='-UL6'+C%;2!)X'7>?B0VDJHFH!_D@K@0VC@ _873C5UF'D$\^]\O0%2G
P-CJRC\EQ;MQB-CQI8BSXZ0T <&O4W=C(WF1<I713+G:Q*WP9.W_&R-K*9'OXV_O*
P1Q<P*45W>?1;)SLZV8E<KWTE)@W#.J+B$)-FO\XN._=Z65I9P#V1,NLA7>@"\9R\
P(Q =:$T.S!\V[BB$]3"ZGH*JUH815-\_2ET8+/6N6G+9SLP@1HC[DHNQ*#FDTI0'
PE :,G(]1G32]^NC1PTEYQ+*97CA@J+1_D\2 XF+"PVN-&<-,G#@FNQ>@GT')F1TV
P,VBBN.JDUE(%DX5])X/\3&=Z8!J<S;+13$NB%<Q#TSU\9EXU/,DM7$0X08)YDXJ!
P@,[U^PU O/#BEV-%K=4-,6ODU=#-W%#@L\ERYG1BN@F@7?_['^]T"L&F?F^"^6N,
PG^E 0W1!UJ'1VD\1P%R2-V'GV\FYPB[Z-CZE==B<(1=(T^_7E3$4F=@<K"XAJ6 H
PA:33 WF$"%"K7BT+:N!R$GMJ?!KJ_U>:-LKK3=9^0_ZF?-V;AO7'/6%Z87H!'[1$
P YRW\J"'X<<B9V*%:-<FN=Y\J'047P#NP3B:GO0-^CD# &;H[R]5H']882Y&S>QC
P/*=AZ_$+F5(%.H8DV.!-Z:DY+8)S8@XZ;/+&9=F9YY[:SV#UPVY&6JD7_@SD>LF$
PGDRBM->B!%E0UVVG.N.0EF;TJ-UEK2Z?LLN?MVPLHZ,&I\KWQ#E713M)4:>;00)A
PSMI1M8U=.(,E5A)7D*'\JZHAJ9+5,0)$:A4)@0^$@!C.'6GZNZ]_^MYM#\WDKIY8
PZ_(5RGJ("?D<XVE&8"[QASFP\9-W%L^F-Z?#F*'T_B#V!:DK(_)XE8E[J$%59''A
P=.QO.1!P+8RYC#@( +DU>M W),*OB3S_"5N3KS>^BK-LLTTEEO]G\B%]LTI@BA:Q
P*7+O\;!\-IXDX?HU;QDQP\U8?=ZHTR*'?0:)VI6(%#RDR6X#HO9UTY*1FDKQ==0K
P++.WM-4RAZ%'DF1R D3"HJU :\T**JO\!HG!:[L%'CESER6;-A:^ BM34R(UQ/+"
PMC&7Y/;SN +?^CP 3CH2!-8NRI.H0WP3I<SPZH,G)'I9>RRQ;H8;5^(HW;.-=<K2
P )VU9C2UYS:G\C5,.S<G-M,[O;\ _NVQ_G5ZL/>#4GJE2A('!+ B[T=2U,?FEDTZ
PQB%;.8:"8UWO 4P<QN0K1ZK]@R8SG2E#M7[MG4J^4JT:\5\P+H[CQOYV4IE.!A<-
P<,H8V>TH(X>#BDHI?YCP+3]&(-P-(<:6_#OFL9\T=9X#/8&IV$W7K"YA!LE"*USK
PE4=9C2>HY[!?3-C<_>:-3H[G#7;"N+YOUVW]Q2CHBCDU/RFVH+CT&5P#C2DIYS;"
P4X/.-LZ:5]\Z_N(7.-XP+)[E\0!@?!_9?,EV=#)L([1U8VU)S8=^V?F*]BH;Q;AN
P3&SIJDNK>R,U4)57RO3M8D?]<F>*_;%^I+I-&NH!=HLC< "%M'=N*76XYO$W@RO:
P_<1>*M5X777$_/X5*OSKM0%?F)DTF,Y5WN#*IM*1C,_:^OX;PV!?&)@IUTTQS-3:
P(HPH&.+QK)KX_5\H3;\VHL&O*4CE/.E$VMFK)IIK?Q[(#5<VARM"G%_-19+3 ;6H
PQNN/($8655G]HP3)_:<;Z,L@X_).\/F>X836#10HYKT+QHSMNG,Z)ZB JNS+:78A
P?WIVK1S,9,&)AK5OD@/301;[VC0.QK5C5=\@RJ'6X:*YU9=-65V97U&"]K.:.+8^
P?5O4Q-IGNQ&V-+KTK,Z<>LW#&_SS &0SI:GN65[$B5(X)'OR&!3T$LO,CZEX2^Q&
PD+CV<@U [Q6CQG2GFTG':MYD..B+3Y<B"2<>GI#S@N:?4P<BLF#".\#)&:0A3,*?
PPJH8!TQ2H/HSU_]\L,;..,%<K_#;#L8Y8Z5$L^> JK#)/MN*Y="_["SF(!LPQ(QI
PHJ0 1/FZI ?X@EZ0 *K_T<M_K-G<DG95O9J,DC)2%VZZ0OT6*(<7:K3N:N^E?P <
P)J<U(D%6S_'CUOWRBA[R'S%=<H&$+T$E!^MK[(.U<&]Q1I=W,] ?]M^J#DEVT"*8
P'+-"MM93NFS]%6_M@]J D)81F-@X/_X_>1R_&@BHVV(G]*+P<XNZAZE@\FH>LM?>
PBC.JD)^,TL4"AQLDD^< W7\])Z,136.8 3$TUI[XYY:1Y)KG&*UU//-QH-<MEU0Z
PB& ;W/QCUXO",W96=B9W%X<,_VT!+GSB[YV:49*+>I+PR!'^&@Z_<^44$GGM^/N+
P_QO/E]ZMN]UJRVTYFZ9OM!D??.87M*>Y'T*"\-A),K0*I!ZQ'#-,?'7_PRYE*D15
P13JYR"H\J:] ]O8N)H8.10 \.)K74/AP)5SH''C.>))/C>)\,^H^=6C1.!;!@\.'
P66KL*;!&(LW_"JGFY2J^.JS-RJDDXBD<?=_6;UEK.B $O3KI*5":4/<;#X!['P/S
P3U,V.#H$Q*D&2I1)<)JF!:2UJ.E]\>/3[I1EG:1&04M.V ]K+:F#OX">X>NP3@Z4
P[ #RVZ1:4>Q_YY_1.K+\\W_$M?%6!\WX,JVVNQ/L4 7G+_G @GF08+?>^1D7%(NI
P*63IYY6!BE.L6=-MYA24&<9]7$H7_$.#3JR3OXT,VK94M*LT>E @*4SDV&*GM/ D
P6&D]-6/5Z+Y:/I#2R+[PE*W""?3(0HL3*F-X%KQ$XS+^>\Z_]\LWZ1,F0MK1J?#J
P?D8\-/I+2?AIO%^7\>+R+SF[N<5N1N$40;W\L1J;DB+D>>O&]@'!/UZ9)/4?GP?W
PRK)#[5"24FD'BI&'3 H5V7PM]YL$])+!*;D1?<>]OD>:S>>Q@[B"Y5. ;+(VXZ.\
PSP.@7M@3JNOBY.BI)N=1$5#Q79@LD"6PW\73+/FH Z> 2=,URVA50)#BWP4F4M97
PAL2^,$]Q?9)^$2CO*/==\[#09G-^$/9O-(C^)9L'XNMN1GJ%6Y_\9-DY*/BSER]2
PRXN6&K$HL%%AZ0 S@Z)R(KD)FYI*S?WC.&B@428JL/( C*UG8 ?#_91/4&FOQ:[X
PF^Y>&P%+53[+WO@/75D+6*8_+6J!?#<LF8]39E8[7HQH5_L5 S._>X-%+S'OE >7
PIYIP2!Q*\>-M2&@$"3$?KE;@UG*PO7;19&3I%W^M)7]<-72"(1BPPE:4:^3U<,K&
PZ)FYO"8Y>@-Z(C\!Q1*Z,N6O$"?"UJ[..AH.&47]_IOB[&[2C,WA-RC'Q7:1!@/?
PD96477] G=1 85[ 9_BCJL#F)1;VDZ/I3>^_?V;XAG>S4)>6]8;G24'"LL+266V*
P#4@7MF)(T(8V!TU23>>J^*AFCA[9QJS]"9!BJPX'_!HB,!BR[)FFFU4,7XPP-HND
P#,M@#>R@T!:+E,6?DT%!6^SKC+#;"H6P1_VH?.]J!_F9M]$\GA-- K[)#[P/9%,0
PU\;>)0$B)P3BY(W;2_SC'=]8>B*+/:H]D4MM+AQ90NCV!,-!V!$=8KQ\2N5$UMZ!
P5IW8'M-Q'F^]]"1<2 VI) F=\V7Y'K5%X^\34H+L:D4YJ,(@@3+[FQ DK!&J'L4N
P<787Y[EQ/H/(YM\N4";D5[[C]=N5:5BW(;18E:N,4LH%DE'E#LZD(O;P03<K:8'L
P(63YYNLQ(98&M\;#MXA+ZB$T;2'%Q&_-<1RV,.@2$8JBYYB;=J&C9Q"] <FC1>R&
P6/RT;!TJ7?RUF.E9D]..#X.KIM$+WCHIT@7PO$8-^WH>3SP=(FBV\<5&ZT/Y9?M^
PQ?7?LW\Z $J4P8*#2LZFZ)I-Y(3+#["34-6IK]H$DA60I;%*RFX?)9RP%3RU@^O0
P!.D5//+&T'?DEX$:/2.<(NZ%;71^4ZT0O:% 3;>)2?3RB_2H/0.,XPVSFXQ!2#GU
P8F4GC):\3;T2-[^2V.\U_7<Q;?GNYL0\$CXI!1XF=6(A(Q"W;:^:K!]\9%X+%0ZA
P#,7VC8E]GE7W-$@X'#3EM9=D]7,70_36 9"JB\Q^36SS:KO%@C(@)C;X5BW"7#+N
P 64#[&K^#NDW7&5ENLXF5H=&!.8:98)Y5WEOR(\P5H(I]17<>[&5AJ(P5:5UG>O=
P.:'BP'6Y5[U.%HO=L1$XV1N@R@4!>=OR#1DQJ"RYQ1&F)2=6C$C?KKC+F#ER9KN/
PRM'K8:@>43F@JZQ)H!W.O9JL$\Q1"G9&AD,!Z7#7L\[*=YY D04HU(3/XHP9E?(L
P -BS[_P32&Q(;4-H-X^YQN79RA\$,@\^"85<#XF_G;:_YD'CCF(D8C(VTD4HU!^?
P=%F913S!HT4"-&F@$,>GB=_[2-0$71]2C?>AO'_WD#.4C,UFZ0.0)S^!6<$9C;3D
P)(C6DHP-\L6/3T*NQHX(_%>@1)"KSJWC/MHGODUN*L^W]2AUFOSO!0>[9M#FA/$5
P3-*@!')[FH2V'H*'9YR8X</NT^G^A]?S"W8RBWH2<K8[(4F8PPIR8YSPE)%<9X0+
P&_W3%S;C/>'  8RUTNHR*>Z$G., @<8_9VH.(E0#%$*^EW/C"\J?[/ O=T%0"#=C
PN1]#6I<*M:TB:WN(0,]EOEHKT[;7S.!-FJO,4L.&-?8%V(1A?6VCQWO=W%P+6KC$
P-S8]Q]!& :O<0NRCX1W4?,>0M1]#B4Y 1V3IMX7:![5U-@4#".\C,LCAR\H/9PG 
P<5,.5#A83W$R,< O*/Q&"W4?8=%>O@]K>8;( $]1M;8CS]),8M:OF?9[1P,;B_7@
P6W1!H5D9SY2JBGEYV@E6--4U9[42(X2D,*]G#3'&-<VM^*\E)L _]!\?MXK%#T\=
P3RE*&CVJ,^D@*V03U=9>+R30M/)V/ROJU<9#FI<+,)A0<_ =NC,+JT[WCF_Y[Y'<
P-' 0?!S28Z?JRUGQBC*AEYX60U0^B9 QI_N+K.I?M8&]F@4N.J&U-AXY+[EO]@  
P/<0+10H$'BZ&>[[ &G DGK)CWJB>_WY?TW"$I1SO;(V RW%G[$_W)YP -C(%;*M=
P5UCPQ__6HAL;A6UWV]]S8"]4V5EN'YKI0C]MUI'PCA)4)*3A F 1.6A EJQ$;[OZ
P86@DZR0,^(X+JWC>B9BOAZK!HHNJF!C$*U2(CQ$',ZBFY'&S#H&%"'5'7C;>._9*
PK",9PFY3!'R_'@/LS_78N+A<*1-\FX[M=%QFUW=>(LT]U>; NQ"Y/F>KL1\R&U@]
P0]5:DQEY];EXF#*@6JWN0 JI,)'CFF^ QK%X6F63G1/$8[%M)$@+5.)09K#<(/J\
PE_)+O#I3.<@E_1 X3.U+;9RSU-H7S]+R%SHI5F)H]/7I5+!^005%_P'./C5\1Z'/
P,SRNPVE[]GXY4?WTT/<-\DR#"_@EZ$]=UPX?D:EP"+ 7V?'F5LI!I\L&@]%1'2E?
P2K*JND$EST)H6UOL?Q^ 9,GJ\S=I7J[YX@K/=PN)+24V&<,G:L?3MO0L4?X:+T)/
P" Z*TJYUS%N<+9':$IK/&FH3IGI4S9Q^Z>HAVSSVL:9X?"9_M+HX;3//GY ;'7^!
P.)>K!U73DIG@2"#,V5->+\%SNT93>C4"+.ANT3]:W]8B("?6\'D=W?4OKHZ=PX?F
PA.)F <^'S,I2<N1YFL>H1.D-?9FI2=6^AO;@6."NHB'_%<A\@O1V&(?W8@0^1K@(
P*#8_N^H@#=@7HLRF^_(TS?_K<8#3;#!T/TN0(ZVHL666Z:6]K9VD44#+@9,@P7\>
P0R5N66<YSN'21_O("[QTK-,'GK,:0VV)7CWZ3OZN57]@G<:"]-6N8.M/8WG5=SDG
P0\3,9ON]BFPS)<TLE]"S3%BD\PY<242WQ#S#1:GO /=1?)TV;9M;RL%90BK(U(TA
PICL/3"BBE521AG. QK<I'B4 >]:[R @Q_:(!@AX'PU8.NW&\;[0:,D,4VQ?]$<"<
P;G?+DL.%O!L6'27^:FED+YV(->(4 4W#-Z)J<H]\='@8$>=O=[?+&_!ID]4V_K;T
P#BB(4- K2]O.,HPX2R*HT5]D-A,P=XO4"2)TMT)!MIYU D#U&\;_Y^4\=PAA-FB*
P>>A3LZ#)-V]*A2D8$'LU^\->:R8T9_"[R*24TGOM["&K?SIMX2E@=J#9GCQM\7XM
PA,5.)3=[7FN.?'HKJ:B_CMNH%[*]W6*7?_QJ]+U3&=P(XEH_IM:[O9@N\[I_YU9W
P$$_"*C^14=RY)TGS%=>6IQY#[UZLJ2?+/W/E_"86+M N]UU=P4?@'B[-Z8TX8ZH 
P4(2TX?:L,PW95>"^:8 U*7,5-0^$+#7C<EN@XD.EP0[NN$X2TJ-%_G;\FS)V$UM8
PE5-KM9([;)HPL-=1?UWK:AIM9)'?:.%)JO;%MPE@+F\'J4K05 ZKAMV$;KUG&9A3
PRMU$N\>_1JZ)4*A_2*(PG/;CJ#+GFIC@EW^TRW=)XZ%3UGCT,J?#VKDI[9,*G24D
PR&N[LU],RHN?;&)CV,J,EJK5UN'!-D*HOZ"NT4:Z(1?*P[)#.H#W$"[-GX Z6^F^
P+KC;.<<-,E@'?0H3(4E>4<X50;.O0R5XI GC(9W]RY73U ZI"U'+;3; ZF_%/A9.
PGR08O^HZ+4\HI@!3&_4:H\)YK,DO5;-W^[W!5O6/AVB%+?H[#CB*&DI!GA;@'D!J
P5@+AVFA*^2&_W<Z*:LY[>Z[K1U8':ONJUB< \ Q3/ TNKX*LFIVKLZ> 'G_K([;E
P'(D18C]?FHNC?E/LQW(>*G#3X!X%'>M:ZVT9]>(YV ?"^68'3:.?.W:??0CD=3K;
P>RQ($V=T;5:V/?RZ91P0_/-"FX@D:*TQ2RVBH3=>S*;\MS L 7.N<K8[OR7@8B4Z
P<CN)HXV< D$X!.]X,RB#1IN:'L_V(H7AL28^;B2P.E G4=XJPXM8'(P2U_:)$6=;
PA;5\B?EU)"TG&6(U\N;LX$U$.8D4[FO5PZ*:IB/0*4%#C(U^K/[CTZ#H?((WL+ Y
P]?..!E\5TOZD#QTFEM'6KJM\.4=(_]D<!"KKBCY-[^_#4',)<35US%0H7?L%"EKM
P\1VRLY-H+=KV&%&FK,T0:PP^S<05DJPXR7?>2'K988>_T16TF<A@:< .7YTFQ3,Q
P8%I,%('GJ%9YC4Y<Q0T2"GTOZ5'/DO%U$7,:8D\F[#%ZP<79Z:+LBC!6>Y-F:(F"
P]V\#L",O09.OXF,NOJR/BW\KMSW?F;G7>S-WK8HNA641G#R^MU8Q A0*DSW?<176
P-:_NVR.&O-QINYEAL(0T((J#BA\P51;^+=<;"QU<*+<WCKK#7S4O&/#VP1E."W8&
PQS$)E^-;;05L)_*OI%4!.@IRD+[QJ!(*Y(00C*"$C4;:,=_MMO"]WV;@U>1'EZ]X
PBL; )$WK9?O?%%QV4LHF67SL3W)AAL[WR9+>1M_HVY0^%1(-0HBIJE(MIES'W5=L
P.*MB:?PX9:)7I65,"I$3^K-]BFZED_ R2/$JYO8(N32<MV#]:\)![]PP,:5&3)C4
P9N ^=I:G/ H0M-;&^1 "O1"IDH&?H>3U>: PDR4%_]Z^J(+D &ZYA,]0]G.99@FN
P)+PU6BJ,$4K8S8-HO0-"$GT!AT1>8+WVQKDO19PED6$)PK,?4:+*4!="OD+]NAF2
PFZG.$*,T\4:W7#]B1@M%37S[S:+7Z=-LWK&^K1\:MOXVF ?JK W\)>YX5' ;YT3F
PV.*:@D/Z4=^T'I!,8*+/'X0H660"O82\1BKX+^#8.]"WSZ/$,=)HW,NL\-N)Z_Q8
PV"53'OU0O!R'$8NJ]\[M^Q3J$J.9*6:D;R/CJUGD7YX+\JK>#QCU"8[I]/40N;(Z
PI+<#$Y5<UFE_RU9YCZUF@B99Q$X&%8*>X7AVR8)GWE(#UN]OH!@[6"RN9)RR+_Z,
P,9++:5B4#+:.@I3JN)>=]%)G>'?/SO6O&6LUO%Q\"*'W$M^G=>)HV67$X@SI$NL@
P@.KT"-U0#/U8@=L=TT"D(JW%OU45*,9,DUR;U;D-EOO\%["QQ! H/.K&O5O]#7%G
P\H,^+<"$GT]I'P7:GFC#4C6.F82:&@)T&C2Y^J>&Y_\!/7WZ7;8WN K6><XX6-FP
P!.5/4N*S.5:*X(5]S4Q7&X8%](/9A(.;B*]P=A@P<1U"L#7;87-B/=6Q%]@\@UG7
P"*21!X_%TZ9D[E#(^0RG8I.EE/,/BH &--7*AF:#ORI4,U=8[!T]*P8WM[PC0#]6
P',FW&#;(VO7>*H;B.!Y+$(J!9'DLV!(V+D :@"P)8<0?=$LRA//0Q\Z,RPD,)_@*
P_>&(AG>89%[E)3.CYNH$.Y!*:)H^9GD%P_XT%Z PF[=F'+Y8'\V.V5WPB&=@;_6K
P@'GV%PN#*+&.,J#!'47I9HC_0*"UE#7%:F,I0>F4[8B%I0Z]@8XF4G34_A5<Q/@0
P7,.APBFY@:=^+FNV%%DUE1H";W"*HP]!7DVC9(H+W4IU\-/ELX2'+DU>\Z2MQ2U=
PMXD_.5&++F#'PY_%I)NALB8OX;BSR/WR%$8="C; "!"7B-088O;LL8#5D\GMHFR 
PG>/CM0;C7?OWC\J>V"H4>2_HY./66M:!&O!&%WQEE!\_GOJSJ;B:_@7MZB,]#UJ^
PB4>A-"50)L=UD]2BO3,&'NI4B*SC@U+!>=CTR.Q\-<A]>7.SG%*-N+* ?SZM(2N\
PDLM_5!EYVP3*PJ#2"YB+")=Q1S"#7K(Q^+=Y0P->S%.\&9?_5&?M#.R&'NS7?<%+
P[TAAE[HX;@64R]0P\W"6,.?3?[<0KY7\"@0"$2$,N7?"R]X%AB+ N]K_R]]\N$!T
P9>+L7L_?6!I_(#.$I""V6G<\^,M0IXKBC!0*.]<LR.4W-_KT)^>L.AEZXYV?TF61
PY=G)V&H8("C'N>O?*AZD7@S?T=D0BO*9U'>: F8XIS7U3-7_?='R*!2<M^^]HO20
PAA,[7S4S/O</#/W+=JOTTBZOO&"2NOX24YTE NK1DQ8.!NDSZ%9VPX-5*T9@1HS,
P<\QYL4'D,!RE8SLHI-[I\RDK#-0T87/.7#2V/>ZJB_ PF8C=1[3;=89<'GA89BHJ
P]:DMS-D;]7Y&H/%%B'4HK*FG=0!J\IIG0K,2?SR!SL>0<K 5 B:7+!K_0*Q )=K@
PG 5M,UX+)V<:9<XXU;& G<16_S?'OI$G2MSJ]F&I_Z.;KB:2/;XH9S*DD?+W<SIF
P111IGS<XX=<]HLD=+O_'^ZV5=5 _USM;*8JSG+$ZLIYRN1ECZJ+.L%\/N/A?,1:*
P=5/*][S4:)Y=_,/?[+<C([XTUV]ZN!_E]031$3+("/-V5D#3@5,<&]_17[" +, ,
P9W*N(!>]FE(;,,MUC$,PB+8LCT:]M[3'1V_K^_NE%'4Q:T8?#%![,H.T&GVEB5HF
PS' J7M#UR$+%.^($;#J_"I6?<]XDCC&<\A#L-Y_:>7^0MITR$U$I+\>K#;N8(H)9
PZP:,>;XL7L,41J6;6KW@#XN.#@C0@AMJHP=9](M^YMG$=Z1Z6/G0!]\=TW@&/'VI
PI2M/@*4->E!XTW-#A(UOGI<)DYC,FN*>91$."QS+E(M6)CLT35/U/*&!D]2%^M] 
PIF4\C#22)081A2G/%6OE#^P,REZEVX=/I])ZRK+85XW*G23Y3;0AIWW*U+9YZ$@W
P9(OR1!F&8'DRO9Y#@S)_"AL=0M^#G'3!NR:].+C>OKB&Z[=7JMS00(,)$<;?*FNE
P8KLYX+*][VR_/:H=J) 8+VWO; %[B'VHQ1=(/$(#Y-!829'2&NWK9H9J0V%8VKO!
PAJLS?RBEC+U.N'([AT(]A=:JZ/_AF'J!7^5=PE\FJF9/0QGFR';B<[8X0+=0])"V
PU55NH^)AH.WUO7?=@KY!FW:"(*NQ7F5)ZI[8A^VUSIM4@#D+E/JNRW7PB]ZS21%Q
PBH'_>Y3&IUD0DW]OK6&L:=Z4NC770<WVV%70<)>RF$=J%;&^/>:]_+0MJS,8?VN@
P^@E3XBKQ[L>Y2N Q%@ZC5?HDUMFXZ#;@Q?(:180%Z:Z47$&PR;C9,+YXZ/NRD(P=
P.64Z%7(X<3!*<(-B1&4SYB\E:(/3$Y)./F;'WZ] DIYH2WZBMC[=OY+%3GQ::4J9
PNUEG_PUZXM%RU A\B+-QR:39C $\,0UJ,4),SK=?=YPU0[YO294DD'Z -QDR0Y4:
P;51,XE VE)N4/?2N1-1:FWI6-2Y!K*_+!G&#^]/7S:=!U,HSR_S9SMNK[=?"<C$C
PI&/F0Q]1NE;=(P/XU+L>[FGJ S_IY[@QI1%.V;L[/7>1/WI"2N%A<6<IFQ237>@?
PV?RHF*BQ)([,.]77]*R)*?0NKI%;1QW,78OU>_VE/@-*YW$VOC>>E,<7?$F\P%GY
PF()C 07KPV1QEK9:@.<$4]E_#Z;IEGL0_56";W!LKC@P2$)%[3I<3HV=#L5CLA<C
P*;UAR2#!6PBY=%B7=>S1_^YQ8^(.^&\2J$_5>R5FJ_]P4FIIY40S>P32[368DD2R
P$.Z7A\3HKG(G\I4.D;OD-LPM/WMZYQ]IAB=:>9"&9+?Z_*JMH$N$\5:!'Z,,@S8_
PZ0_DKL9O%NC4VIG'@\%UC3T^$1=LF3\#[7V\P<[M/S=:CDZ\Z.(83R&75%?-AOK5
PV*)#%:.E=*/*<,8>T*PO/Q@\'ZGAYS!Z<+DFE'1KG;S7 O$"]\9SK_AYA4'F]4"U
P/( ",D=.R(W%WPQZBE4Q'([+31 ,U_T<S^C&R.-)!D7B0-LVIJK*IB"F/S(Q5S**
P*^8C$&.1F38@T]R\5*G=62' [9SN)>;LH6PJ30N0Z57>/K?8T+E0&,[^:JK9R2:;
P[@N\QZNAIZVFT?\0*'.8C)[7V0[ST^%KD#ZU;E.-(X-!C-?;V&WPC-8WG[$$6DF7
P[)7<0M:(;) ;3DMFE5E6P)[H)QT>)JA(1A@V8QJ38;/\GF YS2!KMBRKEV1# X!>
PHE:9PQR.?6$?(HQ1JI=L[OIX0*7YY^^!YP.C.*Z9=^&]D5Y0V VMHR=,LY]>9D41
P/+\J3&AY7Q/;XO^4CNUASW\$YG8P,P!"0 JT=GRKS5DC;&NTS2])1U)_CC<$&5Y=
PRS*PI?2#(J8OSG2_EL>S7&3KM\_Z^LB.0#KC.+0\9-,338+6X,3D9<H4 9MMG)DT
P2,6MXU3?2H^>HJ0P6$*!B'*.$6OTU0SKVS?)QL=)RX% @G;@]/\U,UPF>K^*5"%W
P&=;FMR@!.'%BAZ]'=!TTA9PU:-L_<;DDM@A(.U/A=7*]J9[+DXN[ET05DH:[F4@O
P"VNT=^_3:YG">) ;*A1OL^2_&C)<XW:"(9.A=[!,SOP)MYU/C (NBU<,C*X9NDP?
P9M?/:N_I#<QGV=DZ&RBZ>VP/^$<PKC9 KY4W&FE;K)"@B7GY1X0YP,5Y^+ ?7+()
P30X\H  /"U0XF@#ICF:[C4Q#-V_]W=G0N]-BE'.S(-V%4L[+-ET-9\L*1[CC4E(N
PV].4WI.<>1:6(7AONV>"PN<KUI>;5)1U\"PBT!V:X6=*,&1@\<*+0#RK0=U'>&.J
P.7"36_D0,:]((:D(5\0.2>42=+5?,"9/OMV&@",<JRL#D26=D=[3MS^2C9*WBVI/
P2!&V)*FN.->X2LP$_;D=V8XGO)9F*E*PX:C 5@%9GI5_PNH@K<HW^-I4ML03AV6S
P1UN3>.0I5J:C(3+6KJ!,L=Z-VTEJF'#E4V\_@&$F1ESPEM<B<^%+)!8YN\_YFP'L
P*G8DW"L"WB6:-_;LA,R&PDZ.0@F[_+I !"Q['P[F)QB3\W:I81-L$CBZJ7QKU-:E
PI\K>%$NWH-=TV,PR6(.EPN;,5?MK, B-U1LXTA%/N^E@@!G=_1C@%?'S\:_=[[]S
PZ ?6Y)&#8A89R5G]9Y3HO#!A1.\U'Y97]%U%;>+Z(M9^'XWB'/<\@'93WN27>;;N
PG_5>D'OAP4ATZ-NO!$ *$J@)]Q^K.0!/"9&OG^V'?C 8W(<5_#S5OE,-33]1:;>]
P#=8ZEX7C\1="],#QG3E)=SQJH7XZ?CLA)[(EJ#D2^K(ZZOX!$$H4ITP\;/1(IQV:
PTS/[0_=VT$:VS@*UR,18?DN=NLQ8=_U@M\F@@*X1?&IIU?<@:_V=_#/14$P^Z?U-
PJ(DM+]RH:FOIH\4#)*,V"P@MU99M*VVN]L%/U<VWP*6D)P,#?(7UOLD2??;ZAJ64
PAE)GN&["08@ : *?J=T[0:=^\S^XW:M9M]QS2GC,8,/WHKI,XGCI\]0R1=N-CF?-
P0PMGA_'$P9[D,^C;J"E 8<XB"A#DWXSN9K:A^OA"GK.Y%%5LB"85X5*:(QM_*DM*
P[Q444\1')4'C@5Z)1X0O-MZ</? 1)0_(T<5"<U>-+C]SM\,\VQV"Z.]N>T8WXLG5
P8F#(IA+4.M[K2N= 3DCHCH!RQ?&'2VX7VB6 2:>6=IV4@JMM':57]M?!8ZCR*K'J
P)LK;2F%$^VO;2GFNIT7\= R#+AIU6$=7'^F9BB31SQ%S*'B1[\;[?*Y8RBW5(38-
PIYHE>M;]&K,1W*]U\?M=,.U2IMV@T9'O#FCHHC-\TUH^Y)MLM&XI"VN=V5)G[T)]
P*+.UJ-JF_YI8^35>3GY]8HU90?\8<AVZX<N_1,/98BIC,M<JC6<]V52T8<(5A18X
PLE4;RCSW8U^3FF$/3T"JW:6 6R\VR(Y(5F"U<HI]/E,/,68KG45H7S9/;ENUDEW:
PLB@DH,H4*-S<*O%U_B^>@(:0-D!F";M)?P"Y?QUGCI,/0(.>^A;G)6D#Z]_O.3R)
P[4GED90(%0B3?>F9KK7]Y4/SEJ/16)VWZQ(YO.B?K6BO6-##<"+D<K:8OU>J,"PN
P4AT86:+S%8R<P)($E\31QY7P(?C_!/@&*16J&CR'"!_N>:T;&1H(C/0<KBL]/C&3
PWK[Y+EQ%OW7>/$,0W-C[U0,CIE_?#@*Y*3'H6X\,H1B@2.0,4K&'3,W6WL7-S 9<
PHAL(*6"P(A:2P LN@CE,3BDZP6KS@JW#5UR/^LD-]^Z(Z_MYYA7@IW%FL/(Z]DWX
P7"@3%P' 502MI4=P;5]@QB$CW,6OA9 ]9V'"(3>H=<E 0P)^35#;F1M+6BG>!9'X
PFIY;_$$_%<LJ,QO8#LOJ=@M \.P7M$5WX^@NQ\KQ/P2]25<G/?O,\U+DQ@C,\FOH
PWQL/:G"GVRU6!A]IY.(>@I@U@RE7Y(S_:9_AJ@'&.JTI*Y83J\>?<\_GB R?XA,Q
P0/*1'9=S3]XZVPLBLAA_#4X<]%\3]69.2BZ%Q\\;Y!+49U<O0[JJ,9(6O\:MK>&C
P1DF%9%6H";#BD."<ZHQ,3S:.1*+[PX71">=**.$1,%+:QQ:-SKW:_WZAG X>H8S_
P).+0IQL^ U?VAG#A,M&-@J?G3"9*D<\F\[MP4S(_Z*-L VS[RO;<J=1F0/E?#<G"
P8B;D[*]19/WUVM6ENZI_F8XCA\?AA*X=+MB"K?+P@*:4&-#/\B(0GBJ^4-8V7NR<
P&#H$-0)Y<.C7B%-(J?.I,Z=;)A=,W2M.QDO)N AA("JH)&J3MD9T=U3GGL,;X.0(
PTW5C8X23RT(X9(\YF\0J\9SR'I6=PLC*<YE-^Y/5GL&#TI3R%6- I"BF(/J*N*CI
P[R4:XBG^QM&H#2)(P"A7T,7H]<=\%T5FZJ1B_ V>:P/F\KPYMB*-MGY'(WP0]=7(
P/E1O]8J1:\.PC[O5G,2$B*M RS$C&TG?<M85Z0"1D^E<8:F<4OM<MNYYN[ O.[7 
PQJK;R<E?Z'Q\\J8X]IMSZ?-7>X"EN/ VU' ]US1Y$NEC.L^87I^^<@E\!CT!U,,\
PUEH6W01JD0W"[YQLB[G'Q')Z4ZR#L2=^XDHS!6;-XJI)K#Q/P(4_B]'W.Y+)LC6?
P6^$;9OW)^=GF876&$%$9>^_=##PAD)[6_DXV;"D2+_I29?12Q7TRSCHZSR:>[;8W
PN97B>V7[P4PR&4W09C71L>-\U:8Y=R>KK"BZ+EM>PJQSDY! F8U="[ V XVT])0*
PHZ^&IW3<ZVP=- &L\T1KNY,4Y[3LRC!)S10QA.L?Y/;X9$)RFMWT:.D3+$+PF:HR
PH-\G+Y2/7'THX6%NO?1WJSF'^WA_5SG7KPUR&.A"\>UF_;].BT*$D<0,$^7WT1RR
P=^$^W@%0@H?!TW] OPL_*'DA0)2^16/8<D.@]/^FN:F$,_%_&NWCR_6$WN:@SQ 6
PN?[OIVMSWFZ*8+T8H%V"AGPS/LK'(?>M,]K=)8Z2\M-JJWI&B9$_FX/(U\*N6N@_
P7?TQ0I?+H(C5';4/(4'*BDCG\3>.?%V9S4G"Y8*1M_1;A'M*W[3T2.-Q5=/+E$X]
P$VLFI=G*5C66BXC/Y6&=+ .Q*?8UQA72!%+A%)XZX/HTF)Z_FV]N\]?@#]+(:75K
PQG,D8)"-YH-0XDJN#:4JK\&<#>=L$*D6[H@4%^E4:"-ZO $9F*Z+#OBA4#,#BXH\
P@K+=GIT3>,?7<$.<]G4C\Q;7$FEF-*5/0  9,NUBX!: E<SX04<7RO@A8WBA@X.1
POQH=SI3W=] B7(*1<>C/,"WU"WU!1;CTLY[_OBLZXS>/YJ?A]64-H+._AHZ&PW'N
P3>$9&^=%5T]]RG$Z?.M3O;?!78QN3.?=-;@3=(N\::NL<";Z*GL"MP 2R$O@%WN0
P! 2D]3SJ=@,5J.?N]QYE$6"E[3WTA/4;JY"72;O>-J7 +QK#3AV\M %A$8UDXV6H
P <"!,[^C>Q!D.U$"3M"$^&/EE\02AV/-C7B-$XNY<UJ KF4+FZ-<_KN!SBZG9NT7
P,IEYZ),X[F-"4EV2;:I9/%[II>,C;8_!<J2L*&ZS53L3E36_:/#N11'N&7I0BZI7
P@M'^B.Q1P,KGCO1S9Z72>.)MT$C@KE.-=T3*"<-F4!0T_N41N#ZZ;]8'5"3T_DTQ
PQ:JBC(+8-0_$#E<1G;!XX)9 *NFBQ5/:>9TBI]\J\X='/*L-L=EG5'_+I-VD[;C6
PS=EC_7R&'8&&SV%^$,:75"_*8;1557S'/=! E][*I2"?U7?Y8$?>"*D!.=0KG&.6
P5+[=$2C-P%-E?D&2JFG0[P4Y8=6X('APOG[!)*ZM0?LP)<,-R+^3K3INN->L]M)6
P.B#NPWB:PLE'RS$Z#'EVVR+_4/IX- :VH)P6&4? @7WRTDYSD:W)6O)5;#S! &X.
P/E_A6>@$EN*V2VS%?U=(08;EW8:?#SN<VY4<2TX# /:4:N1/-Q" H?,MNJO]_/P\
PRAGTS1M,#Y8S;6P/O!.=</(ELL#O4@IB7'A@$I"#\W\JV'T!:;+U(,6KO[=O)Q5I
P24AQP:W:(S_ZS-6<Q2N :1=?,;H:8@D7/_CZH_(H/-HEDA-"78<K0C2>\!BP)-&#
PO%>:V.-Q<SQ83N8HVT\=CRUODF?%G<MI-ZBK C6:I$-/@EZH')'(T9@4J0G_E#HA
P)=I3)J-(/9(D)- #6,(]ZX%O&G'6!9?_'SE,>%3X8M_3Z+PXGL-HTL;#)P)-:KW"
P*;$,<&J+73YVE"J'CA)S!/[WKG@)VB$1,T4\%?-3+8I3!9/)O8-']X\EYA7B;FMP
P 'RE4GK49;KZE\'B/YG0T8U9$(4@G5DW^K2+%JD(D#/1W.@X%$-]TCA7UHOFYZ5I
P5X=TG4*/GCO(F2W-B[1W3G]- T3G/;OU@2*J8PC?AYK(S%0V[8N6[;[JVHG/U+"D
PFC5;:@K:)A"Q\O842S_4.YMQ8A7S: !J1UDVR_AO/;_0A0,^Q(LXUBUXVF[LBK'?
PSF=\_ L6_X YZOSG]LE8YN37H64ZTXP1OZGQ8^6+K61;WCC!WP#88U6+?W_F$WVS
PSS.(UVV'RE)[I+^AD4+<MRL@%3&%$*?^-*3$T404J,DDRXW1,*GN\5?,7SM/9,!G
P9(O[>XB3%.[AGUM4) ELQ; SNTI 1LVGXDD%U\8(AJ%2_?_^\]?8[3H.^ZKIF?NU
P)LV3K^(X;=.+UE_3T]^EZUA78@DQ:P$K48G-- 'RYA+4):$#J.OHI:NH5R5QE6*I
P#RA+,QJUE<XN5R!:5!;WC%FAXW6#_J,%'2U?>_ Z([E>!E*2A0&+M(C-3YLU']=8
P0V4LEFA7.9&_8[_N=-:_PI*%%R>R' J?;=N1[HKR.Y(WG\=86^;?.FQK.FD?J]OV
PIA$2?M==6D\?AN+5GU4W&QN'+_%:E@463H;%J@*]-2*_N'#JX"#6//)!'%RX?E9(
PAPMW-.(;H:-Y#5D>S#F1&,$XQPCI-9F8.6DIK3WA(]Z> LYYTY%!B5>*54%RD(\H
PP1ER=.[+1@VJ82>1 )R<,[\SQNJ#SOUO@GWPF!WFW&<!RMMQ)%)5O;YHDFO$R-G;
P2PP]4\3K$*TL;="9JS'RA,,6EX[D9U2*&)9 #'),]]76)V]<%@5YQDC4QF@S.K1$
PYKKI$Z;(9/0[:$03:@Z_H!.=&F'9.Y$=-^0[T?Q[$"/I#6-?2S(])?MPY"VV7I4^
P)>8,'.GF%B<.9#M0R"/TV7B+'HQW,Q*7_ZZR )_M**@CM7;MVR5=T<F3UD^$HLU5
P=RROFI3BG6>16LA7FM$O'<'S#52"^0Y7O'42(R+$_ZV8W&?.=.$6X#A,@YR$PF7!
P2:&^)H48(2AS9N6TM)315!)E^P( 8!=?=UJ&S?FI 8?0-K2X%(]O RSY' 48T9WZ
P[SB0-PQ]& MYZU!-R3864D-=6?59\XO3QN%$;UXV;!5P*F-T?]OKQ24&V:+I(+PB
P?QZY4KT8GL 0^)IXQ?[7BI87XS#8F"7.T?&\<%I&9CY0O<"8D1YG9V_U.J673^;]
P'D(4H#NXA52)22KRUX8FSI.:KM?BEB<^]HS86EO#58NH5;!7^W"SF'US'LZI # !
P5I!\2U4ADR*)Q7Y?*JW0=&/! &9RL444T%Q#M9JC3WV/1H"_<Y"%:C(SW67P5L$!
P*?(%RL)-W _(LZ104<4276W/QC^=0:_'5S$;CX2->K GZZ6N/,+O;ER,+B,(#\%9
P2?#^TC>[#,[IDAX;0Y+-HDX4.AG"RQ;G9GX<DAI9G8K/AO^D%H(3P+_<&GQ/?[2F
PH"3S274L4"U$+MAFG&_39HY&(#/_$Q-0@>11":ZQ^L3A[PNB\KB@(GH.Q5@8/QOL
P,^0@GLL?$NC47G!)"I-C"T(O(SB% (;F^V0F.JAVL,IT5JO]#E>@$B8<^=>2D:'L
PI&*L9F#Z4;6&Z6)#U-KO+E![3='((CCC;\O8=GYOUR=Q1 EZGP[3-)/>OY]-$KT;
P"D# ?[\>.IHF7;TOU^J<3M Y^>_DB<ZF3MLN=$ZX'<=.% ?O95-A6#J^?;>$?O^(
P]Z2_/M0\9:&6ND@>D!!V*_-.L^USJPZ=CE ?5QENA%GA7$A90.(! =4U_&&'"(O_
PC#G1K2/3*2B\=DV+2"L K)^9>XXOT:E%N4'I**N]; ML=2V7^F)Q_K+3.,&3$42>
PJ.BMTC]9@5(K/O%.)9Q_DCI!U#28TF=CE#/Y@3U)!<W<G]FZP_JJRM7-$M<@:?WC
PG_7Y]_N9IO_"Y1.D[[^SW24VQJBCR?X.CSY[*X7=!="NJ566V[=^<&$ISE/&U_SN
P'QDJ!^7O06S6P]RR_I(A5%V[%,CQ\W=6[U2(F[\5P'^34&=S,&NJ(]/BN3IL ^;F
P%>$G4HA]+D>E#W8&0?,9/7Y7:.9#V1 ?UQ,5GVG^M51 .G S'0#Q1MZP W:L>13O
PYYF@4I'6G6!M45PKWV.L7=1IW/I\B7=:BW]?/[\1'TH[*/H0EW$U?7P, F%1:^BS
P:=!GTC1F5FYBM7XXWI]98I-7P)3\2[0JD/O="YRK3[-Y57SAF$@/@<8%BCTIDTV1
PG+Y_X(6$$D6 \Q5-@MZ%J-9+L]\5)33,IVY$:,.F%-FN!]&4ZHKBS=WV077>S? X
P6&%N@!]3IDC#U\5FA55\<9>"\\T*;(%//C#\:>ABK$9YS403KVM;A7>3_)1=LHTZ
PBM<NF4X@O=+P_$^0.*1@V&XF.\4^*,%NU]V6FC72+6?(SCF '"KQP:-ZRK6GKK&#
P/3.,/WYV24H[^?7!*;&Q#XYGG]FF)[4 +5P@#0/PJO_$>(<WG'G(HUJJ+<ZQ*XP"
P2_M^9-LT,H\252"<!W.(7MCG%7-/_) B2_O76H=AS,8Y<TPV1S0']]!GA.'Y!\6\
P/9 $*YS/>[,=$RP@3.?;E#Z0;M:+\5V7D,%4C:JJ"?NC?DVTY)Q[, 2E'+;\88?/
P8MU(H0AXH^_&=I;Q;F*4YH:ZO+T%3E;[3# VNV8HG+?X\V.&B02;# ;5#2DNK?+I
P3*)A:VQ*()R,AZP:,X67_OXH"0C4'VRF2),_+>MH1^$4._!E92!87]W-4[-46@?)
P43!]?2Q'S9]U.U@V0F0NWFWD*6& 8UA=(7RH26S_I8U-VX#Z)HB4T>:99 [4^%=_
PQ0 6P[>G#9H*J=FV>**FIL5<%J_K@1@U#!3_T,2(IZXX11+,3/",?80IT40"H,V0
PDX?2D<I05.SM'M5QWXN2].>#7F"B-Y38#P'D;RU0 O5 H:. @)P<@^!&+,5U3<EW
PMMED=V!NT()+:BQ/R1TP\B+DY2 G5"7QS )WHWY%[%7&'.)CT_\?*O]Y8B%UV7P"
P\2/#UM:T@ZDZAGT$H07@&29;B-N[*E3:#7L1.@=#5Q;2P[\4D8B6WAX5DS!T2X4N
P7R"">M>9DD=F2)P@2S/+!/^NFKVQ6<,&@)F)\F=EGF&#^P4MX'HW[0C*FXJF,F4#
P=U7W#/,$I4(H!: +S8(= U??.\?K% 7O?#V\PKQE'#TQH%Z?V0E5:6\DF\5\_H]P
P@IF#'OC8 +X/OHVH;K<5 CY">:^R7P$O8(E2I/WC^ZJ4&6-Y%5WN2KFQUWTFLLYA
P-C)5<M1/P":7H]HA.F(1</7A V$**[906D(9$-!9FT2J(\8\ L8PN1[>89=#"U;I
PU64Y1$@(JY:EFP1'5/2B($QW00*TM-?URB<-VV_?I_RX-+9^T0BJ2-V/7'^ =6%D
PV=&^1<,@'B7=)-#V'*-XHM+!TOGS23_XA#WTGK/BI.5NH-_NO.18WS;;+WJ2-ZKA
PF>*3;K/YR8/C3&8C2(S]5?(/H#^V3;%RIT>G1C^?<$?CIU=+&Z_49<&/M^IK4/O2
P+&$KE:63NZQBHI6X,(WW4UO"G (S 18SK2O#9$?S"-#*:X03%MF@_=ZC01!=#;@A
P7GS<&#/)Z6-.-$=F_Q"-?"UPOX/<V>8HJ,:-$SS_P>GM&Q8S:2W V L?.G@CW4!Y
PII,F/[9%!*Q1=;NMUCA<4$*]H]>0:74);[?XNNSG@'Q2.)X.H:Z%:'N+0J79DW,C
PI1&Q)B%3F<FCU.)+2Z9 LDRC]GH_ ?)@-1%!P>@?3&/W:F5Z\(G1?&6'DZS;E9X5
P6QXY.UV_10%+-L(L3K!NX^0?80ZM=4A!T1&EW)#G?6/+;]+4-ZENN.H[1M)=P4)W
P&=8^P4P[>F(T8MEXRB[.S4QZ-@/C^]\QZQ@]&MZ*@/,IG,(GKR7]V%XP!$RO/8 :
PBSDHZ$Q";=MC!E]C@DB!E5&."JZ3;:F\J=*(":T]86: F(']E&&!G[I=5<OIL=V 
PK0?Q^C88#B1>MH&)ONOBJ6XO#F5$N<?-GB*6X53BQA]#RNU9 . IVN[!7[(2"8D3
PN$G?YYSW[W// MF>BRAY/^_VCI\L<[%JU@\YM#S0_4KT-Y5(@@*>TEN$%H(L[H8I
P- ![&G/D,=*D=UI/OF<#,R&2RO_R]1B7E3CK*8"*Y#D;K, -,+);LW%]+ZHR-+FK
PENR?O.AFQ$BP'77QNQ=U_NJM[!V[OMQPFO7^<#K;]J\/S"=-0)'I.[D8E92B6;31
P-\ RQ+P.U $+(!7CQNASKG+07/\03PF=4F+Y1!4A.LK7 QI]0%3C (?1;0=[LTD#
PP'1T#R+< "U9BXB-??S]RS&6/?_$ -*!PKSB=85J?Y\ PVL7M#?R4UUV-RU>Y4YO
P:_\=+]Q\.1=9HQ>^;\QI%<Z^#<Q17*C%Q6H5D$47@+J:/?_F234*67HR-LU(XSQ3
PK+#+ABSRY:H_ H9YQUNL>LR^\P9Z/=L=XN1U:[?M7:C5.003#HE0N3HJ6SJ)UPX>
PY'^ _#+9WI[_TZ7RA+\&*K>KF&V\N@W[AV59@$Z. ><)@KJ GA5;;QGBCJ *?Z%9
PN/55_M_Y% T[&I!520BB6:T2;R.%(9G<CQT79((-Z/5%-2I.L((F,B-LJ80BOV-9
P$)R8D2=2!M(V%MDD-X6GYHABPT7'WI2A[7RBQ9K+T&!3\!]G,"ES"A9R]T1)TI3<
P60/A<-1-AF!T/]S\F#8QA"PM4C5S/'P)5%AERO%30+2(8-Y3ML5<C7<UW-0XGTF]
P2\81U6!E233?R(N^S?*;! SIX_;FJ8U1'-KGUJ)AB3822GYO,+0LD?X?0CIH'7+1
P.*PN@-#1S$".8955CXHE0*DQ^HC<*)F:VH]G3URN+T8EN-'( CM?LA4AAU,%&#WY
P38A%JYJQP_@!(B=;25TZK2<X"=V%%)< YY *57I,#@YA:]L'VE$G!W/(V" :E4ZA
PG98[D+-VG%DAITFXB8FOYWO]N<@>T $47@T145NXEQ2.$G*P%)4[N1 I_F4,>H]M
PI7D"^PS'(^M#,(.&./+&LZA%'B\@.:*>S7975QN.I3(^GZQP;8=7J8I$G6]&=3I1
PT4AB3BKX9-<;6K]0/%V[5\022=$+G/A919B:1G#OQVKPYX +9U#D)XR;_-8$-^$Y
PUJ'^?[W:$UT1'APZ=1&E@1V/ O#K:W\AX [< 3@W8C$-8/^1F?%R ,X75"Y8M:A/
P\7+#SU)=\*>4\YF 9),:^P XG3?75[E(M!V]GK(%KD! "](/W3@[3XE6HP>DXI-6
PF&Q_P_^ KO4-4%<N>F#0\FP0ZKMSU-E-\Z#E817C+0!7J/S!1?=IPL#K$[0,4G.+
PX'QH "!X="^AZ+!X%4CZS:%-8DLS?O]6*1;FF?C4U'A1A(JXABV8#\5X6+9\K(N^
PY426W 3<#WHVV4R5D,5ONIDO 6D+^&,R I&UXS9CPO?:2G9$?DK[P][TG81)9SQX
P=0PI,Y,WU6.UXI&0 <@NP53592&<Q95*FA53[E'**4QV96S\9;],JO+.T^XW28[5
PLZ_[_R+JY"+\]2,@7^*"&)TS9NW,I!:)TW!U:IGG^/)S\'SD-L<^QYRDI+,-JNQ0
P;M^;"2DI4FQ@T1!'K/;+M^?J]CM+?>L70'2=#IAB5E/N>;M(1^V(D"/QS(QR5)ZZ
P%^0(*OQ\K6$BFIE:'[3MX4AA[(1W$!K-5,+NT/.KHF6?+[_08),E/M(Z5HXLB1B:
P&^MJ)(8#)EBZ>28YT";!?GO^2)729!CU)T&'"RVQ$I9(@ @Q.C0-47B9H<9W([=,
PMEA"U@F:1" --S$,71ETR!=G19YQFXI6*%F_$3W^*D.GY&>HS<CIRK2=HD,<?Z2G
P\WVF8>Z^\-5,G/DKXFKQ%_C1E&'T,7]J:8%G2-3V=>T%[& BLC;H7K H[<F/+Z7.
P]MLF6:)%)1M84Z]!:%M4?[Y C& #6OAX8QT4D5FU([KE]PIMD@C!Y<)"UMEPYEY]
P=UQV-,E6G=0,B)@-]0A(\D<4 2[9SC8G(\6[6,W^?H_U?O#(^8)^X'NQY+@A;Z,E
P^!8_28X72Z7%Z:+'_"LS7#D3>/=&GEKN[ESLQ_:64)YM,7!W-GUT06T/ _S3\&VI
PIOS03B[;FOMI25S7!M=T@R:GBD=<S2"O&M\($J7%8-SZK@K9,<B &487QO 5 !Q2
PA%J,SCV5UNNRTV)9%DW#-1!KB:<]RU>28YH<5HS;[I_KPYZ3VHIFZ/MTRM!X=0:-
PBOV#XJD^&MU9!1F.)Z8PAUC#$$0(C'D6\EA\T@3A5?'Q>5)?^$@9,6VHJ\]\#%ZX
P4^".HHRNC.<VK<U#K8%^X 2T$/3''"H834<\]B=92+SMY=1X>W$&FZ8G^NL+B, Z
PIJA)7*_9 )4X;"Z#IQB4)QJ2/+""FW?@P-6>3;*_0C8I?Z:N'),+,!+M8A#X_0_Y
P1&$_4BL[0]+V5'UYA*GA>\:(3UTIR*I;.#(IFII84(7J]2_>T=EOF"SV+:=P0_,R
P84:P:)XR0?$?;%Y<I7U85F5KID%&J$OC?(.,(- CH^D:HA*@W*ATBT'? T.:V$#!
PD!_RA*J78Y>1'S>%'?,\6R/"E;IIOP9=SJL_/@OIO5\L+?>Z#MU.! _L:RMP5^L#
P<Z@?*S,RO^_CQ)9IH0 5K^,7?IRX6MB C5A U2B)>+C*G=I=B9A80EE#5:ED)"6G
PC"K8W[_+\W$?G,H%*Y,JAWU>AN@<=WN$/B:1SZN4S/OS4%.J\I.S -5=9TJ:..] 
P874)U@YVVQM3 =7O1/GV27T6WWVP*[7,[YU+!QVH('BIG N3)RSL3!X7U8F4[Y)^
P[T?U<=X7NIY;FPAOJZ$#)4[,S(8([YH!T"=MWXB1%S\_I=+V1^Q;2.H@-4F->W?\
PE?3-*/URCL>7V(-_@ZM3WS\!-*SB,=%@)DF<X"XAWX5GBR(SM+XSXHD,%VAH+8V>
P8Q<M(]BS*^LNYB@5!8LJW#/3Z-"%EKVXF_!K%) &[/$4><QH;Q1R-DV4WARFTL(1
P<-@QJ-[(_"_(,;[Y/*%=< 0/K,:<UPV8NIK382\J4PPER@6_ZN$E.0=>^5Y_]8L&
P[G_CW9I4=*,>@QC$_]OR1P!22&<PN9PLK!;B2KL*(N'$@5XF=^55.5VHQ656@8^O
PZZ!@BOB3[WW->RNH=JGBH3#LJ)=KEV4&NLQX&\M^:[J:48'=?;FORJ^[49*[S&R;
P)PW/(WH!F#VJJ<UG^%@7H\!_WULO*IIXCP?(D*R[L<@OO TAZNW3[$6(E>"8H,B-
P+9V<\\$?.4]_1F'6(RQ(302Y;3W2[E(;FD793&/4LXP"(24#P;. JI@5=(G5/OJ(
PA9C1P":9,# @ETR2$V'1TW10<C4\SE2(X'C1ID.!<Q>Z#8TJ@R3]L'WP,M!'-M@-
PN\Z9)@X<"_[M@)G1SV;(8+-+U9[6#"S";M(@[%QQ=!*=4I0G]R_L!SJ@YNW.EG9$
P+@&>U5YHO;S+2%M\.*U*^RE-EF1)"Q-TM5[,UDZ.(5>9R#!:;UH\,552+;6_6-2$
P-(D[$S2$(V8MG;V7^]PV:U1661G_DE;9!!LH*9&.S=U;PDDW4,F/LH!*0"DMYVD#
PSO?A!$G(:V*KNFN^04"G.&<3LO@C_DC-]E8#-'^3&B6I![?DX="5@JT!!H9%VE<:
P7R(XA(7 .G7="PNVGLM76F8D\H)G\]@-_P)I0:Z;MXP\F ; 8:8S5,5=NY&W-A\W
P$.=N6W/C3 N@%<'X:^PS^(H05H61-$A3F!Q#MU0Y'+X>$-?\M$($_L@:$C*7G!P6
PQF^SX3?ZYTFQAA!@B<^,#&CNMP4)QEH^(%V)7;S'5:?6!<KBHN#-/0K';?^&+#,T
PQS,S(W'ZBTN,2U0T@O%C<A)3$.#PJ+:YNVU@F-Y!=YW:CW_@A\MBF8C)*+7KVZK1
PFF'4M0@T4%3.PN.Q;;W1E<6B)GX6?]5UTMB )T-"O4K[5VT6%#!"-"-H%;EB"5?)
P5_40,KC_4B-E/)>LG)^1OF_Z(-;/@3* Y<:ST!H*T]NM'>]O/('+ Q:]8CYQMI/$
P*?H_:)]+5\='CS"[[@V^]$^?A2I/&VJM.+J13!C0?8:-*O<RNV"YV'>14G"&(EAV
P4<Z4?D.*BL$YYU?FA-'9$O2+FBFA! Z#YJY99.N39=0^O(+UB3G4L^/^2'N_DF- 
P".C:F#LT[JX(T-11D1PR?XQMOWOW5TDYAR9-+]F_O KOR?K8/K?JVE*+PI/K;WI:
P%C54<R(0):Z:)4%*?^;8N6_]LBT?64/,X=/2*NC^?>G@W"! @9=($*Y+5%^0'.IL
PJ,-R#1K9V=Y'#%T>+NHL%-@]:LSI]/CDZ&3Z\DZ#_D()&79^&"PY%R]1/A=VK09,
PU5UL!D'/3!#L_BE3<!7(Q@;F5;7^T"3SI4>^%6Y;3AA>)_79 S38W#8ZA8 6:6]+
P9+D@"8;OWL(F%3P@_<U'HY<1DQADUO'7P*.FK[DS^S52C!1K1"K?E26H:]$"M8Y!
PFNX>B:D2@00(5)>CR^4S$3;ZPMFQ-PR3<\1,,^DXH1IZ#ENN*M#QT+FF24@/EN9=
PUP"U9T;-#81I64:57@W9__*:_Q=@O;S;8-H"GGD!\/;C/Y5*U$;80 FQFF2_?ASG
P9*,/YF'PG#];OS[P)R)96"!\E-LK-LS3O8\\0(&/ *J['B")&:U\/2*T)TNW&0@[
P *G,Q2.\'$JS_QRNO..SL#\6^F6W$5!Q&Q->S.DO.,$'J)"FSW_<;"D3,)]%POZT
PS\->-YC#@8Y>3/ZA8DD\K-,,X&KM-J)C(<DO>/M9.]%JV@A)?!$E++K%W//.^B[V
PG-OHJ+(BB!HXE[N%^/,TG U63M&+(ZK^..JHV3$9C[.DW>N%\M=0Z2:'"WV3HR'_
PWV0!0C_XH&#6[O=S0CE1O4V9]\%85=A$C$#=02(9/A]N'ZV/V1C:PU-DE$?(=DA!
PY'W,YBC3T6J1E <YT<R9I>;?LM0_PQ84"=L6JBL0'>*<JD]^-2R&/7EK>\G*'E:3
P$!MN!HAT?U#HSTU!;"*?%%:L4#O>#H>4;5$%(;EJ)ML5J?_'RHXH".\HW&0;TTDR
P,8)+K#(P^ZV=!C1OU6ZS<YUDGI**(7>$#QZZ*^S&&(6)RTNQYN&TI[0$:Z3/*'<X
PH+5H@&AV$CN0R8+P.T"NH_@DKP4J8:P3@^.P'^VYW\\ANK@V[@3!Q_UG]T]>.CPT
PW!*IR2^J,"Z6P&91&?K%#IJ2:XS\N8(-ZSFDE.6$I!NJ,*!,5RO4O3*JF]A4HF5=
P^MZM.0V/%/VO$KM$S-N14S-1RA49L /5M2/$3N-S>MDA G5)T70+E\EAR'/8<711
P;XK(7Z5M_M?H@=!6N5+U)<H8X\ )Q*<_">7CFB:P?P1)5?1"_):):]*!659_IGP3
PPCFNPEE .9CMVQB*,FCF5K'IN;._L.@)9EBHOLO_GC-;C#R23'=-\M&^0$^W2?=_
P#59 A;)F0'F=QV >*W8O34%F?'CE)X%?A;3F[I#Z<G_B8LLG+ZUXOR]=2YQ-%&KE
PG'#LKH0&"?DHNOPY28>RR)Q(*]K"T\QU.88>3%4@YJ5@2WMR@G" !(/+)3$=EVN=
P7K0^E\LGO<TFCDK@JWH='Q2V7GNA>G;5CD"#D/!U-4?"T@-WQPUDY]"Y@)AH<;CY
P^6(,ZJ\=J%!(6L.F'2+2W#8"[$EAT)GTO*A[*3NDQMB] H9>-X@R5;)'4U'9C<F=
PHO_N0)E#\70+6_^66N$L7O&*,MJ0 52%3_";I:949/3>P*[$<>Z?[?:OX)R2)$M5
P;BFG7+TK.^M:VAOWXF,^@/C4RA$Y/5A!(H8!PL9ESM@_ XFM^Z,)AW74?*1E&ZT>
P#Y=JE^W-YER/%,FRB>21,C?#R DGDG\IX$/*S:?"SY9HH(:JB/6,US%=JO2K@$;A
P.O0/F78D3X+[ADF9)</1I5@T=W<A<KU\:N\CLTHBZ(F_B(L]5_@UM?1U8J!=EW_L
P%F-KQBE7<=HBPA^H2?9Z_;M3(3SG-9NUG"-ZJ*E,#S!:5_CT#(#%3Z6^7_%]?H #
PPX7>"&%V98N="M8&Q8IF<E8=&W<@72I 2!_:G#X7;W//M+\ZYCBD^3G#C\>*>HZS
PTO%*J&(^J1$X7[0"F0.G-2Q+^_Z@Y+04X=M72"+P41^&[L703PD:'RZUJ&W6F[*)
P^K>C!11:-_TOD9UL-YY]2L=.B^K"?^Y2=O*/^M/S!G";F R=?:CXTWP>?C' /4Z[
P%U\ZRMU=STD]1)(3L!6[(G$:"KKWGK506XB(U)Z 7:W?^69&L,;9$5(/2H68D&74
P-?6ZUD5YV!R\D;/]_6H  >^3)1OV$K)%Q _J.YK<$5!(QC]"IK@LC)%*1-7&LZ:]
PLD:P;UF45A<PU]'2AG.!;7$8-U\*%%GU BYTK5+AWSO";IYD_HLO;E8_[UV?L@$1
P?V&[G@09 *]&GM#L@0-WY28Y])'( O<(S.MGSS]G;;P_7,-N6-.A9:5#4N[_?%G>
P;7R7CTY.9K9IQDC0<@+/IY,6G>D,G$!]T#LV?S?B?#'>/U_7(N;Y(:(L>DG@Y*RA
P!2UEV*S'@X<7KU\(Q5T1.(6J^X*@5=NQ! WAW?!H-Y;+V<[E(6IZ+'(4\- >@ +?
POT*:S)Z:.&U><'$Q9YY2]+;3&-ST&A'9<#95S5OUKIUY?ADQJK!U?X54?00KGC\%
P"/F-K&1]A-]F(4^(%RXS]16C:;5D%S2#0LHB+-!S(4M@&6!J1"FJ/Q8B&HC.5_D 
PTAZ"KIN-GYP\9WVU4H_$ ;B/('!U0TAT4Z:LQ878\<=F5R&G29$?ST"7MQ2\?5:C
P EMG6H+ G$F'U^*!-QZ-"O%M$^UKP=K,0:XZ@X&-$[+A9KV^[70$K[6"XL!J<V:V
PR,C\;F-G;O)A7.=#D0PEI/=4J)$QO\801,F;N 5^\L]^IXB_R5/4M+6X:1)>P0/K
PC,#(GG'Q! CZG(C\W\M!1@U"GLJB#R\D2]P6[PU/_!B /@7-)'V[S9*L01P(W:K<
PP.C3/[Q+FNFX0UU'R:ZKCX@(^C0\3VXU_)D1*AMN=P?+5NRLS7T62*XF5;.G6GW?
PZZ,/*DEO6)YRBS*Z S\5GMRI'*H/36C 5&?,@N6,7,DGVPB"42BMD8M7>\5Z*<*M
PZO-:I,^=3 6^6=;G[[="9/A%R*F:&9J1=649R3HT8SW'"/JQU_E9R%G2>;B^=ZVL
P!A_S732K BV^MR4T%#H;M/P'9=VDH:.76D"=TM_JA;X GM(%TV#$XGH1O/;V\//U
P#J =&]6)GNV+J1Y/"O&;["\2?1O,9VUUJ5?!NJPK-UG6#5Z:DGUR6S#HL\V+/.LS
P[^\?.QP))%L>@U*3._$V*?TJ_() -"'S?K<P EZL:/'=2V;5(&P!?^ZV-J/VP^?*
P,P_'$0U^C)Y^[XA0R<^!HM3TH,[S"Y-^?+M80%*B$\1!_(QM-^9[]?H8$%3O*^47
PQ_01 T(AHA$^PL:6289]D@,1!/&5P?"P/@95%,.J[6JR0T--SC8_,X,0_,RHLL&I
P!X-[K+")H(LB=**0<760B44DIRF$+;GUHX!)@'=&M6G/>7UX;AM'IV= W)UU^W2;
P(<^@9K;PY?DDT @ FGZ9%^;(YEF$Q[#AREB+GY%*F/G5PQ%$RWH1=,?#@$+>Y1X=
P5F2Y=2?*$:BY99B$*.!['T$HR)7[@P +4R5KA^$(>,/^L*YJT RNU"$LE@%"*T:@
P I4(V&L2H^S1N OM<SA7:, WSR/X?65Y.Q?3N%8DB60OM$<"C6[VE)R7W&]V%5^7
P@EKW#G"*U_Q7="6(V9Q'AM=F.83AC:WB8;2/T::]4FO"I-$&42RL#QQOU[^)G6O$
P)QFEX<+YT\R>(SU;U,K<=O[C$:+U8UR<7%$:GQB93;:MM<<_UI_X]O\G?^%O?M6"
P^(__W"%'UYYTXQRC2.[F2T QO_#!/!+M 9MV I&T7D\:D,:&7T1%JZ6-( \Q8'NG
P=D@]D?\F?QX(&S1G*^.S/O2]YEO[6SY;:$Z34TC<QKWO%==4\.Z(B?"PLCX\:%T"
P&G0'E5M71"S8Y*(_LS UMHX5%4W"+.S /#=Z?S).SM\$NL8.FV*JZAK6_;Q&\_T!
PH..>H7 LS\.[;[^@XK!0]PI/,OE$7L:&[K#W8-@3-[KGLAD/GR)^J"DK,[1!QV:;
P,5(K8'SW&HNNM[%+VU.EED]#Y(.5;D)+C)X%=K#$/&:N3:XW4DQ3?/M+REA;=;%3
P@'LY@.EP:S&4)G.Q0*U7B42^_7 $.,L9HL9( =SWP' T(_]<3-LK'@"&5[Q<(Q86
P'R.3^ZM%841"VN$1B(59*?%Q]7-J?]&3 _,/C%[1,KX,K86>_G0'NPB,&:9'6?<\
P&^2W)84<!OF>3R6*>F%H;9]63J9$C")Y43=\=XI*78]YR49J]^C?RD]2YI9E"T(S
PRJ4HW\PPC*>0$-A\G%MKI>'0V#6N$TH@\5O(P#KUW-]"U42QLK2SL9-+^M^0\0M%
P&6J(G?AOO N)71]*D+CE,R^(I!B<5ZL]A N'6V13*4<NQT$7')@/_QRQD0O'T] V
P6<\*/](1X>K+JQR)NM ,KB4VM4"'PNCT10R<(<:1"<*6R>&B7+7OA8:I"GEAK*J.
PBP;=UPE$-"<'$JS=:PJZ1RY$60I"_TE&3A,:9&9?"GWZPVQ&J'."0Q32-R-J#A5H
P^AC8)-@_!6;VT9'D[99WL@JO+VB"D/*X.+RC1W=+W^.UR@;,,\$V/!3N>[-$8J.(
PX8\;G]Y[[D1U.LLDUJ7WHLB-DFO !>GV5Q/R[71[EE]:]L2&-1_ *0NW^CQ]_V/3
P'U^BX_=ST/_M+]^Z4A"BOJ=L Z?EVU<0DMJ]O+Y\=_ MJZ>DL^GH MHW.;!F@8=<
P_Z7KBH\&(=MRDJE#@VW1%68J%S*((+=E=SF)X=E4D?Q/%%%F R+;H'-Y"9R3+B8W
PQM7:51W6S]>/9300^0LHA;1/ C2^E8S<Z8I0ZC< 3;V'%@K+NZ^*N_D57;7]UA;W
PIENXALS.:TEV;#.U(_A=6<N^/4A#E$Y3VUV5+3'&W1-6G4;2JEM%>H%R P?,+\_F
PA.>$+*^*'VUH/P_O \$*+N/XM!E'3,'L5 *)K7Y%9N@$9$?(IB'Z#%15MD<B]$CO
PJ;96_C<T6L\S66V-S,:"HS";_WN8^X0#[9.GXE OE]7R-2[4A$?L[;%H.0O5A+= 
P)7GS_LJ6!"(+WCAZA8)@#GT1O<RWL,0VS:UZL0-?^SWTC^,6P99W[3;LP4F;6EB=
PG=L-%R ?Q887%A;\"&/TFW\\2GIQP]WNAEW"326N3%.#G<Y;U[$%6QMZB!H%Y5!1
P1Y*-UVH/J_A6\ISJPRB]U!XJ1CW405\XJA[KSNWKN\)=G=+I,=M%3O8WA^&:*"UT
P> NM^]XC1I%\+.T'W(,&CCS?U/HR("#+2M9G'01SK>\&RFWM51)7$)F5,JO3K)GM
P#Z+1J<),#I)4L#Z31#51+&&DU>-T,%OVRA0!C:.E5G195"L%OBQ_H6JUUGY8H^4B
P6\D08X#EA(*691Y5LXW(FPWXS'?IU5%,Q=[N+8^V7!&HJ;8NJ>B\_*@%9!:$P+'=
P1:[X'+ IZ94[X+(@J(<NIRP)%(EL38./@^E28QWB:,DK\GU4W$<$/!B17< %OCT]
P$VMPI4%/8>2:.&' )PLL,WD6>"9U"]?OE=UFY\7,=$H]S<D\E!#3-49<-@5 ]$BJ
P/$165?8S98+ I#!2($LR/,-A4G_!@'8TWOK!UUGVU'+;*E.(C&XXZ"R/1BABZQC>
P*#,6BHM;&9Q9N_R<,'/F@-[;4I.6V0:[,;-['WU'7)RL 1E@L0=TJL-A@5VC%P5-
P.DTLRF@@Q=)GKBZX:Q*#=_4Y@CPO-N+J:BO<Y^(:P'N],8 ID@&$];A+*Y)!EDFN
P)SZ!D?0&8/)LY?V[%KP3H-89'%!1#1!-SG%W.?,FSC3O5K+,NS<CXPF'1\C-L:@=
P"L5*=,+'PG&FHS82>2M_G:,\PD&7YP0-"78I/3PB#A@H1.1;\N?%2+I>^^WP(3H%
P@94/Y&RZGHE8/E!+D4F!.^I'2'E$Y6<.LR%;4YN"QEVJ?YB6*ONKE)I%@Q:1M*1T
P0%P18@,$<=*1C-NM)'[T'!?2MH=HK+OU*'U#\$'8+;OL7 U'%MM(VJ'B^2*JL9Q;
PX;&C(.%+MX=$U>G5##"KT-I?4L,C-"QBSL<X%R>&QN)T-T/)T_F1?HA&JF0&IMI4
PK5?(D[4GKF68P?D->T.D0RG=?-F<B/!%L< J,VG-JO$G#YRHJ(0Q9=-@V>C$YU$4
P5,E%=>"JY^9D^'D<7XIQD3@]8"PA,#/?*%:E[@0;SH6[*M9T/1K,483M_^."9_'M
PZ/[1VLIA+[K1P;POK0]_9V]WJP,I-OZI4D8ZB,4](V3^SK?,@ UH+(/%HTD+HH!-
P5UL7N!_ID.GJ$<8@TJ&:1V5?47<\E7ZA[28GH4+R5,:.@.DVA7@B45.YN^@FR7&E
P:"T0N*+3 1&D?P1)>F((C2LF.'VKR_SAF#$\TK[[1$*5ND]PGIC^H<#$*VY%M<-3
PCIBC*J -.WEBR.Q]V_"$_RRAAH2BPF<8<3ZB1SHW?-X;?ZI0TH'+;MBPT>:9/<&^
PU]H#G3F7_$:>!O-9\!FX-=W@0O5/+'.ORH/RN:5DEKRI=N, Z&T*7B! ]GQUQ$FU
PT-Z9GC$ VR\&RB90UO#R$/6PH+RU.2I:]ER_!4[J*@47C6.X("]T$HZ*5H#'SG-'
P7 !&<6JA')G6A,*4::UJ[Q>C'>!*T(RG9.+C0,"?Y.*65_;K&H$7)G/W .NX#>W*
P'IJL6?T_%9+[:W?(XQ3]LUS;3C;TL;OO85MV;6C02$4O[ *)]+PU3K'$L*8H'.#Y
PC,^=F?>T:;FKK6!I;HJIV0Q<AT%S(DM$GY=X:/2;S6FUM1(C15Q1K/!J[DXHB)43
PGFS+RWX+J!Y%R69+LR'T539+]_\:>E(]&01-@N#1YIR9.91D]FGX:'1')%]U6<1W
P>VQTW8S#F@]<$""%Y=3O&?[NSYI/L;>UEBS6W(Z1@6V#?",'HD;V!,\_21U&;C!H
P1/3!9NC PTUM1K@,8_(J)U $M8]"C\ZN1L/=$,UPA#GAN*)-F)@<7NE8VDPE,L$P
P#V/#ZM, \0PROIM-*-$\QN<_2"XD*._!AEDJMBF/6/K)HFCL[1^QZ*0'61*NR1F&
PQ&D<OC-LWU9\LH \]%90F/<9>^O#R.B.1<)]:#ALF5LA0%*V#]75/JZ&[9/5,6A&
P7@7^5:Z^%@& I['H>NL25S6W!T >@D&'SDFCZ$PJ9#%80O-\-BY-5MKE*PBWZM#4
PK=BQIOS72O@/<E]CC)H.!;+!\#Q*7PCUN_6.&F^P"YR#QT5"H:**=Y*K)V;G4<22
PM5O2'X1"<87_V?#RZK[-00#=, Z'*$]1Z."GO'_PT>PP\O,UFA7'[('FT&!9Y?4-
P:N9 D[IE(6+@$42N7X*.#0I]K<H8)E^(?:4RG 59&P4ZZ:)E!-_/@H&3!JKAA77Q
P/=T34UI&8F -V:880NF1@H7Q?/C .Y9N6 F&ZF=53=';;Z$SF7\A7C%P@4;IJ+M9
P+;?G #M[?#=!W+./RJ//V#147<[O<B ;F. 99J OP3)LI>B]Q<5 S\&#5G+[H,U?
P^9( Q4Y9 H%WM ;%PBE<&D:2;I0Z_2;_'']8?K=Y%2VU[TA^)M*B&A'URX^G9M.:
P_T2;6#<K2.\S=5_M8E'7F>W+%C78E+0= JU3LM9'?/];KJ[-W*#OAS0GN)!=CCE7
P-HF82(%Z_XE=2=@FN4%DU4P$4$F\'=1?="=@#?$)SX2"%3GTK<(:44&)@D5+/M\O
POJ[XV_[^0-)1 *7@,.]Z#&K]N*0GWP.*J,F,N+9J8]$@XA[(C!O0>:^NJF+'G)9U
P1L)$L/I3@4>8%S.<")I,6:S8 /%WYW$,,%"W:>J7'>\T?9Z#*R<)VG87W R ,A" 
P?2*% $SLI"/[^":5GY+CLV_EG,&IP>;?MJZH62,8CW5ZZ9W+2.8=![;0(0WLO:1)
PE2O+YPFV('KV+37OJ(0A0W"F>CGN^AGMF(GR# ?[1,;N$_#X:!L:;]U?%!+]>W H
PNT=7CEP2!> C ";=%(1PG45E/Z;,5O,$6QP1LE-%Z2\3T/T@I \YVM"41%8AQ/WC
PR.HWBN%7O\\.:AQ1L"041;@& P/#04QW>$_A)+&#=&X]EA.W(Q^W+837">SWA+4A
PT"U7:Q'6%(HF_U<IVIOX FIS_=W!WUP*I//-#E9,RCNS\'BP%X7'BD3Q0290\/ /
PI>^:02U?P%\^3=5>O3.  \Z#1(!GZ3P:S0,3DIV/48<#R(0/X__1+7WULPP_+758
PD%)F&FP+-!+$^&Y )[N/\O2%'0+OGL@M>)!Y>6]VD\H <%/2%G/G&6OXF/Q)P$F<
P/*<=88<5-:1RTSS&I:[Q7PI<CE44@,.,.(R8[QLW=JLR\N\Q2Y\6H1F0U0&R44;0
PR=5@=/;]9\I.Y:)M#C;W $<+FHE0SI"J25D!7T_<M7H/8.9'@\;I5 *HO;BY!#>U
P,3.P^N5&^9!U3-=^'K7E&'LV"*OUXSM].N>MTR'ER@^O$#3AQA#?<LS46WZ^J]25
P?G4K<++;;P\HCER>'O.:_G4$&_<RZ7?)%*#O%;/:%95,HU1S^,N\F2K;A_#^)G%5
PS%8R^IR.QB64)XG6M-Y>5!&>B[V C%SD?*M(]Q[.X\WN/-3OY>$M*J;8#W/ME1$N
P3EVM6Q)B*09>%8O8K:-8.^HHC'D_R28E%]J?C?2M3QGFC-,"0D^$/R&HD-$9LO[$
P"_16OVS4U:[-'+5V)U)&AQ?I_+<'\!*ZCJ(B,A"W7YPF3W-C08P/,3DK\<OD1&36
PGU*+9 <6>6WTM??W!2LT3A:%R%&H@GJX[_GL-*R)V4',!I2JM,26:#81,,O&-=('
P,"4,M+O77#C#E.;[>ZRO*$YIK8F^!%MK6!T[&?]OIRS'C.S9AD,#=*E[?,/=]33E
P;/9$1&RN7+):^ULQ<$3Q?C1L'.RTM:C%7#5L [C7DNW,<5R-W385HYO,[#TM"I%:
P0#,FM=]:P&"G&H[HV'W2\Y3]-/$*<U(-^RL2K2*.ILQHFM)#8.A(@14C2<[(YD8T
PTA!P#.WQM90N>\R24EVRG16?X B1:)[*!P(NM94;WNJ=53!OYI)IG*'\'/.Y26+U
P>ZMI:C.CG"/YH*F<&;^I:BNV/)_!$6Q;KD$G;S;./=0&_^0\XVZ>5;"CPO7$F-%<
P![T]V(<'.Z[^)X2MO[.3#%A-/)AA:""<N#8Q%5NFD&I3@>5T.O U5H\TLBI"14D@
PA,!<& G7W*0W"]JZ:(.12%J!F+),NJS 41!5TR,5OPA#2$2,2YU.I9YCR2L_]7$'
P?TN+.0.USY;7B-' /AD\G\]UB9.<6+!OH[/>+1^]JPP\LUY"PCD/ -$/?9CD4#6@
PYG3!F;-,?<5=GAM3J'#R,9*:_#O)AH 'M+1NH9L&.5.%;S&RDL'=JSZ>AX#U*4(*
P&HPS+>CKX1=!)_;I&EXPB)2GM%-*OW%M4*DESETN[6!JRM[ I#_*8@L723"TF?'(
PXG(.29';ES@NSCWU/40.L?TDI>\1#C>;[85FW'%;\F$NO$*5.A.A93G2/&,'*VEC
P?6D.PTNX9K2T_VWLH!M'JW4283K +'\%M,/TS02U-\B/<90TR;2+"8>FE!T1#6>;
P$7H./ZZ[.42@.GDJ4> TPV;Z0YR?#??9(#&VF_3,G1U/^A-]N0'X^U-+HG\22W-N
P@^%*-;-E?&$G-0LM:G.@1NBU8@^BX2LG0-0)"24IC=:5EJKH^5B'"Q714!' TLE1
PD P%#@P"D-I^0Z]6K%$B^)^M3G9*[6*C15,X>6=E,2K#U1?N07^$"2T-UJ'P"]"P
P@ID&:>7]+//K2!+HH>DA\,L9Q=L8&!5<P-M-TOR4W(,M?6J4\+="5EZ"1BZGYRK>
P]K <B<]Q)]1-V]@E@G5$3-1NC=N?"I:7[ANSQNF]3\N!+3%2HI1_-SBNG*<_WW?C
PZ:7;S'G<0S%7-P37+;[BVR%J^^I$8BV8[5FRA =@6* 35@QDGT487@YF-/PDVR_,
PPL"%N<*P+KF=5W)QF.>KE(PO>#-4S16)?.ABW@.2">,A4\>^DY*X>MI^*Q,"=?\9
PYC9NEDXKL0\!Y6<;K?&ISPSOC< [^-PWT@YF?=ZA6#V%(D:6E#('$0G#F?85^+[F
P9M]!5GW0>%6@RCBW>QE98D-"!#Z$9FEA#S+^4XA(N$M(7-#+_&&TYO[SPB("\!^,
PE_!_TY(K]U5:H8F7UNFL_F[KRW$F:GE$N^JRO4H/+UM<E*WFA?BQR&?6X%ROEZ&/
P0!J;V&5K;-<!4DG\;[QRN%3*@PCYGHC2+"7'0NN/ASP^,Q+?5T\^8H>*Q8#YE/B^
P$]\1*H#Y"3A8MS.G4XKI\W$ #[S3/ CL:Q?*('G(/PD)_< [M&A=Y(>7,UEET7)T
P[H;VOEO#[4P_&#]8QB&X@)$PGMC)5&JMW:$4?MX]!60T(],)^SW@E(#$B7CSVZJ0
P1QBY@:IBA=(0YUBNC:UH"<-W-T'"ZYNAE($(IZX^5&?&[S*L)R-;@5'6 J'&:L(A
P%%60[1$+L/U LX4@/L7#_> /LL_P9UBC'-\9R1Q#3-X^Q%>>@2:J?>(C)<'=+&\D
POU(2H?6J'*7U0+%<Z'-B+*)ZCKQULO#RETCYN.3<M(CTOT-NGF@9&^F&O.)D&K0?
P9@^DE:* ?]$:>70^-I70<H (QI\@3TLH0G[#3 T7[@),7G2 V*E96%,OM"JE90.G
PJ#NR^V3^I*%V33CBDW?*D *.A[?J.AJV=@9;2YP0IZ\E"-QU]9H4 &]/CL_VDF=7
PWML%LZ,K[H9U3-8S 1SAW>C@G<[?=:VFX&4.Z)[C->*![_=/KEP<6>:WEO!N>_PJ
P0)<]-D/0T_4VV8*)ML9!E<:U#WRNI+Q6YDTI[\I6>4?.,V.$K=7+I(0>W,0]F_A)
PN5763J[4LG#=PEEV3;3@OD]'?*V_Y(2(<_-#["[4PL?-D^<F"<']6#S@3R%=_IJV
PZ[4!W3DU.Y)'WNQNZ\C>";$WD)F'/<9O[-$;Z^4+(\0^A,3H0_R&J#FCO%:"% Q>
PI>Y#Y2?5QHDFRB,BF'6$DP)82J.[Z]6S@7K<#<X[WI-TT2K_+_ XUKNCS5O;DFJ!
PWH*ZP,'JK=D[G>LPU@\/'\*0-JE,;<_5F)J3*Q5+NC7\;GB2%>I#/#T<V4<X[" *
P]' J7%<C@YE<4_AS!-#9(=\$[I!0,WX-5DK:*,N2]IW1&8B2(@]JX:ZYHS[-!RXL
P^V1/E/X/B5]=3A_>6 -+MF%4=AZ+ 3XM)>FLRNJF7"$O^#SY6TJ']FF,DFN>]L!T
P$)JI:YNC=[S-M8C573+,%UF?\M2/!,'OZ]+&^AGC*^:?4M+"YLT&'I+]W"B3C6$X
P0,;%_VB[V8N$L@VL73X>J:?FU-WW9Z'GF&[ =<>][@*]UJ)CIPNR>L%!K\/^PRXR
PIWJB5PV11ZWK\WO*:>5EZZP-J:T?+-;89AJ)GN!].[)H9=6] C)>#M&A'RKO2\6U
P>(L:M<OM"X/Z8DCS( M_!BW! VJ&16>?J><>K]RKU3 ^ XC#[F7U[Y5G[W5+<HCN
PXT1#4V0^C;";HQOI T7_\N/R#)J9:^^B'"J>8AN 1ZW4;4-#3!P2^7=%P9RO@)$)
PECOK&R:R9=_IQ<JU<13/HOI8V#0S=O)^^6^YAW$=I/T;R&Q3B:[M]NIMKVHGZ?A@
PV7SG3-UEEYINN:OV ?C)6#D8JYX8&G%J6( 46C@=#J(XS.(4 IWV,6IXS<S5<@48
P,0 U0# QIGA=4HV.RP0D[ -6?5:2)# "J:9#>W;9N%W*@#>G0+!P=R/'X>B!>GLW
PN<*5NU=%I6[3NY>T1'P*XO#@L=)<4 ^$'HYNS$E44^F#_4MPE0?:>FFW/93G_6&E
PU6L5=E=;TF;-4:,ZXZ#UD<"O<K&:62A>;Q75^&T60*%P(Q:8M%#+=S5O<,N2QOJA
P*R^D>*;2L;51W "U<36RWO7NFK;39#ZJ6;JS_VS1:*5F%;6 PV?5_W@J"5>L,9UQ
P;WI65;R-Y/GO#V@Y)LC8,H<$HL_W+88+1D/K3M?Q.$&I2-YHDNHVBNO+V87^6 94
PS*>O+^+(A"(6K/1 HU'1>)8EX;&[%FBL;8&9U,SEJ 97<>]#F\!8=^*M2IL]7$UG
PIELQ?@?U8SP1CR3C WAH&<%.[W>\-:L7L4G)JL$YR2FGA[3IZ[=,V%R]V9Z Y>6+
P*L#.?'YY&K,\IFR^NM;&07TGC;<,[7G[.D _>_K@-I<P91R';_H',^#55]+0G):Y
PC!!('JQV_">>EE*'-D%GWGUUYEB83V^G=#<Z'7W?Z7#=:@!3).TU-C-FT"YDS"?#
PO8CQ[(1!VGD286K8GF1Y0[7=/45L0&5&J*CL8JYXOW!9P*YBM!#K-KR20(R9<_)H
P.D !,<YOPNY]N&1VL%/_(KPN5ME M\\C'?=6[/6;M@ ["BT_&/TE8VO.?^L4Z.#W
PE*'GR>H#PYJUMK( .VBG_4]G6#>@1D;ID)I0/4C?*'Q/R9%--@=+8/)V-5%DWTHR
P30^V4</GTDA,CO6M;_@=!SW&1>M2>&\2(NU5&]_-"J_M3"5Z#K/7N5'+KNU,S$@@
P*\24!LAYLL,R8Q88#(R/MA;-9<R5Q@O8<)3*MS7?]K]:B?5+)!?<K.,QR9U:9(>@
P)[Z)U8MVA'AE? GEE._MTT=(OFA[G"1-^EW^KYPGX+&0#+?T(/?$?&_P;["):,XV
P=Z?]3!\FKQINQDR EP)#&H"YRHU\]K% W[CUYH!U(<R/6<H/V4F90G +%5';70?G
P*'GT-S.M56!:PIB!JFF"![UQK D%7;+8ZTP^C6A%W(71K60/C$ZOR2(8PUI\R.<I
PU.3KWWR%!!5>,]5O#/,+R14T>=C?&7EX.96M7ZT.V["D1[\$H:1 :2AT_?)_$7-:
PH"3(B^\/I3^7&BS:ZP\9"39);*XS$A=V'S#K3M]ASZEZO')SXP0_<JOB<-UN8I%,
PC4W[3+.!"\51P$?+<#!,BB<[?K(KZ9.:^:K?<4?$/:FPIBI /8V^KUX7B,\U**[D
PN&<6E;%'-I\>E[&/&2L+A\&Q&Z//3%0ZQYJPBD<.\L.1F?HKV89 <F9U6E%R"1T$
PO5(P%O<T8%%-Z1>J<;<IQ=*84+OX_R 7$-(4; W@T-%#;$4+&F)XE><J'G&Z\#BF
P'Q]F&)BN?,QA##$O,)(T?+M.&#P EPHQIM9ZX7U#D]/NK"GI V/J#=1V(6%H@HH1
P-&=9XN9E%:)= 3FCO"_[1>R&.T"#VP+C"8M;_E[BL-M[^;VS:O8O8GQ3_Z:7:PS+
PE#F57Z(R@]HU.FU' #(JZWR2(>:MV7=)OJ(F'##P?_@//ML0<;RI^BPZ/"%[.*L*
P7 ,P;.#PXE(9VQ'EX"[XTXW<]UOY[2M^JCV52VF//,Z%[BQ:K%-RNMI:&=SE ?LD
PVA_M?(EZY]/JL3.%7)C(9>HZ&N';E!@.5"4;11&GM] !(1:0WQH-*?JBB#.Q"]9'
PC58JX..P$T3[ 0OW$1G)^Y$F5($<O8/B<SP,UBX_L'5R>;)PO2[?[B  _FLX =IQ
P4*,34O)6""UX5#_F4:I/UX^GP%HQ1*8@'6G^1[-G@$J)7'IQ0-@9KPUCWXUI<R-Y
P^8/P5(0HGA,&4OI5%8VA:1$^,[LJ-D0$(\,U9P0ALX-CF\?8(Y.'^(UIH3ECQ^O:
P3QJZ[\90Q%#&&OK37Z)K(-8L3PF#:\VOPPQ5U\29MA:"[MZ4]$1R]YE)I7-JZ ]*
PB*FM GNHMJ KM"TZ/K-;WKS@<DA8^J?<<&[ZC;O@9YR+$OY\+M]=(8.J*9XZ&IV?
PGOG;["_?8H*,IMTG0R^UAW#3ZYHQULOEE/MG>1XJ(17 T$! .[YDH9>.!4+8U.3C
PD"N8-%("8'?>3;@6&-I"TLO3E'BQ-##!44S:W(5O0@S7!SAT*3\C+DA.I=1U& 0C
P@2^!T@FB5UV51CIV3.W'8HH"82A> O<P#%7IA ?'!QK_SA1\6#)[#59;K_)?5ZZW
P5V"W\.74W%]S%!(V322$%]I@Q!'J0R!PJF+_SW7(F[%]]0V]JE;?0J3AH)D*GXAT
PGVXAU#5%RK-8NC?AA\Y5YF3,])YT_ 3=N%/ QQULG@V]!7'#%/_Q2N\6?J$/KXM&
PCNNHN#E [X6X@(^T,Z%TUV0:O8'1 ]K[B!)8P0,"H0291XCTF\<55C/^ G^=%2EW
P+I;?7(4"X:_U27JA I3Q]3Z]ZU@@Q/7Y !J;L,@FUE- 0$BX&E2-4XVOS\\&S.U[
P,!QN0A_@1N(5+_0-@S<B<*UFI.\(N?]#3 [SG )/.'WW64/8_/'K]\R>V,G7B'"H
PWN9Q$]%CJ@*5:3K?*WQW%L:OL_Z,/;QN"]C90%9PH,NJ%Y61A%NI![NQ'!F%ERAI
PUN[HM=J/Y:+?V*Q)>S?EB9.=))C(&F#^4\TNV$+V3DG1_JL3J2GF28G@778-WD5_
P\%>[2X75ULMAB3F]84 AXKJW_J,P<C!&O>PT6<(1X<,-D5'0>;%FJ#!C?FFG/=@#
PZ74>%Y[K"PNFHZ^M;MM_.@=*K56CG2!5/QCTZF[$6F>)HD8PY5(EF^Q'>8;6\IN8
PUAZR+Q'L:" \$GU+AUMS-A&G58@B1]ZD^.LXZ@/\Z &:8Z.T.*:NSP4FOII#W\I-
PB5)IOMR%JI7T7,WT9XB(@? C/@$P-.KW7.,]8MT69/(88VD(;0:+73UO*TJE(FYA
PJ=F$Q'R3%PNMS%8^P=N)V_+Z,'X*,SK%R6=/+ )Q+/ 9F?H(>]TP0SJT%[WL@$E=
P;8;L$:WIV2Y\[*LV?1W'^V9F0U&EWRF K;YPO+J];1D4XO4J=*/ZDGU=!D^9=R4+
P@U4!$\\"BO7$MD#\]]M1F.1>!@P-:X@GMPT<3"0%'+)]IW](&=O%*7J[B;5*/6RF
P'6DH),QI+XJ4A3S3$/V=;KKQ#&_.^8<M$/4./>-[W2;B!_-<5J(5XQ?\20TQPDX7
P(DOTU&6.J*R<T1CR#J_B*5*'+1&H!V*>%IA\BQS?@D@I3%#&/OW,"M5V.Q!KYU!9
P*YRG3>WMM0,#!FO@)9SI;<%551B]?/&6:D-96$ZEPV5B&LA!=*XP[9>Y"V<&^=NM
P"!K8WP6,G8PE'.,[<IZX\T@ @HF$F!M=H#IZN)67($7_]M)GQG>&H'#CYII@4E2Z
P'5DT3"/1ZE/U)=!?<4G<I[C9NO>"<%,U*7\.-RQW0YA8>CY5J;V_VQ!&<9:?Z3M;
P7$+8>*[ $_1BD8ZPGI"2]Y155]^:9I]Z#KB(R UUN"L(LG$:#^,!IQ.4<:FSI3_F
P%AZF;PQ^HV_AO>_*+DAY*09-2 H0:[ER]L^5+.C35EX%KIX[?F&^NVU0F]BJ/@A/
P$$T3,T17R;'_ ?DS<*$!C)S1Q%D8WUI0<G"Y \_AH:_B(322F3TX@X+6TO&"PB*?
PVK*;].G'<BAPVZYU,WT6'N?;;%,8Q0$V]@B"&GYAY#_G=S,9CF^7$F2KTFR2=/H8
PY6[VI8P6;OJM2-8\XXAQ4>$"0M%V NK>UV@C3&_0)[#=+EWY,=63$EHY!\XZM8(+
P2UFKF9_P!%!\KB$7=4#8W&JHM"+KRS*EO&Z57"< JYXNQD@.?=5>K_9_(!#[98Q*
P)0.RB]!IMNF$6@IPX>ECVNN/V?'*6K5%"XS32%$,*O G/..;&S&%Z+XIDKI:&J5,
PV-&[^ZQ.K1UT<#[PRS";$)]:G"!!%*;&J=YO*<2>*T>[ZO+)?38;O/V?'_J="WCT
PE/W8I^VNO%8MZ:6_*^RQ'R@(83CI10N&#^SH]0":D/\NLBN;Z@;/):C-]*)ZG2^G
POQ*B=M14K&1H62\-)EP0R#.=&L)O9QL[JSV10X83!D6R$HY<U_4=?R1.)^Q+4$9\
P$UQ(Y5MJ79[[H!HKV2Q?5.O1GOW'CXR2;SLD9F^$"JK;*+KH/S9[<O0[DD\6"P\G
PF6230\S>WYYTPX*'@V%,;G+1I\,JI_ZHC*>ED$<X)AH%5O"#O^'?6ZAUN0\PW"2Y
PAJ1D"9]'ZK#!'W*BY"BM(P9\R$T$*[TICQ4?S(7_M%F!09X[LGTWS*QE1<7NFM^R
P&BB52 _%VA+XFF*]/M1?XZ>@WXBB5B6*:]G)2[E+VFFLN]UD$\3F7JE=L(1@O%&^
P%X9U[PRH3T0(]O>[2<\#H9N/9G(3,CUNAG\E$&H'KQ&JR"HA5RW7WD0#$ON))[H,
P$(UF:RVMJYD@R:IR\N8C:,A\+.!J9M$E\N/EHTO?KS!529[3^]Q)P<X]W':_9D4Y
P%)^0T-#<3<,;"4,X$3VHXEN 6WEU/F4"EI&\=W^41"2MJ&T3);5]<I&;C:#86'*+
P^;HWIP=?^]<,6,)-YSY _E!!1H^*Y@]HCKXR:3O1[,D"T&DJ69X)YF'G4B^OEXCL
P59IXA&\$$=2C5.S;>L,3Z:!#+1,?.1:%I-;M:J<N"C;J%YR1=W*;%?G45NP@H<6)
PY]9)V3WT0R8*$?U5&0$!RI4 S5A3V!9^75M!0<9B25B33;BOJ(=_!P';H"5(:*,%
PJ?V$0@,%3B_406Y;4S@8M(1<B<R=BF_F(V!I,\HUW%@X]NR)\U2PENF+LEU49O5N
PG;X=,]]UA&<G0PAJ!*&FX4)F92OEVPT"E]#C/L1+'\6YDL^T"GR4!49K_JC:[>X"
PYXOA$6^;"CW,,R+)G5/#+.!D*O,P6Q/#F_276V&#0F%/5?H*B[RP%[$IO$;$HDWI
P1F=)PO1.H*H52*&S$_;ENC:%&[@:%M,?5[+Z!?!.N,(-;!&+>Y80WDDO"N@JF=82
PDDI'LP?.!Z#9D#?2"VU[%D*Z9SC^P!7Z8VK^>CE/QV%J[=Q?,-*2 H$-<\Q#\A?8
P\\IA6B+'MG])MBL8)%\S^-#P2"-GTY//9OW*.\;Z5VCPH,\?V]5,HJST5RFTY!4*
P/@(1+8M!&J!)=L>"$D 5+JC8#BX]/J8H/K*!TI?+<XY:A5CHVMT AO_M,UA?CSY5
P3(Z<:6H_ BTF70U<T3_Z$"S[+,B CS_V=L\SK-JHQ'.91DV'[C>;_N;.\.,_)XSV
PP"/5%-,Q+@=E4TRT5L/7EEC7TR \"[4HF^_@47U5F2P.^A/]0ZF;)C*41H]I4C4V
P[663.D5B-Y0C^.QJ.PS+H#Z55R<_PM:;#Y<@.J]#-FZH4*V!4.#*I*9I% ^%0"15
PP8XCQNOG;][NCSO.T+2(M_\-A(7L,BV01KLO+G6K6=E.) ]^@;MZHH'(_-R]DV%G
P#U?D@#Z'EH@9+G1(TER?AN#W8X6;L'\.1BOBS$57@28=6IU5#]#L-(J'T4(C<[P*
P023WL3\O8&E[>?+^BM1]3"/-D";+@@&,MGY+TM+V9J$Y,B1_D!@/8FRK@8X;V!65
P*]N6P&]_.&HHEE=GJ5 !TQ'!]0.VV,"DA38S/970KC4:VJ64(K;H)"U:W(3*6NV'
P=%C4LI+Z96UV.>3O#PHVI$ITP)(DW>*=/MGK)K.K0"AO$OB' EO/U\ZM+@_RK1$L
PG+XV=#LC;3_Z+A+8:L#'HIDJ2BU&LVQY)C=TD&PS+Q(4,=H9GZ;KQV+@<LC*9FL?
P.QKC=9FQ"5MZVB;JU3W]/"I/*_YWY,"('#K8 @POZLM*$*7Z[XGZ1\!<J-8(?DZ2
P>Y *_A['U\'Q]0\Y1D=5MHZR&Y%V.>>Z+.FFKYWF< Q#?RMS;]4C?<E]YW>[%Q%I
P@C]@U?MW)C&BI94U;>'SRHJV(EN(FFCT-#O5N5G$MP:3+($)^JNM(:7Z5H2SPROA
PK)LLB(-]Q[9?;7 T,?Q!K,H.(A7 -W-1&)A5/P)FM>UR&2W^2YV0YOJ*(W1-N3"3
P8M(!J<X*,_/BH3'+&..++GM-V^(P*(D@C3#VU9%/>^PHSTK0IHYE7/K*?IXN)@18
P JSC[?%%'4LA R=8MYRA35/0 D[,+*66YQ-<3>F<DY#DQP5_C GOF98AY%X\SSC4
PG@^/+M!##*^UT3J5YK75 E\[%EO()^EC3==%-GAS*S^EL:ZSAW]4*2B*_P>4F^=X
P19CPRM"Q!6(6D(59%0VIS!'W<_PE Y]YWULA,!LE31A?^\IT/[R63&7IPFM;5*$K
PQ>W@TBOSO,;8BI<OGKEA_$A@=Q%NI8O'FB)Z6G]^2(5/4TM50AH2UD"P6$+X'A8\
P3PS<-TAPX BFQ/L2#.\H>!A711J:"I0AF:KJP4%:I:2MP3YV>Y UV(-RS,Y!OX5Y
P8S-<O!B>Z?FFHDX%\"?9P/RA[?$\8@]/+!N D,&BUIPR0$(&-=L84K:7P-;874\I
P(^^>;ULE6Z!]_[SO3/_M"0+!W+0AXR! <3%5L8I*_>>R[DZP6B1B(>$P6])9.X!_
P?/"GBNU<IB,ZHG-B/5W";GYDO*O@)TOB>1ZO]@04NTOI:Z<EN/L,<*0,IY8QY3_"
P:H6,DA':^33+,B%B#2>:TX>X"SW9SQJ8"$O91.&U-8][D;=U5A*RWNNAJ[ZL51;2
PN"*Z+?S(-W;K"-RF]@K5.@[RT4<.]VVEU\@#Z5>?XY_^$!\^T7.7R3D;[= 6 C3@
PXAK" 7NLB._^8(#MFJ:G3BXJFPSTMA9F]&FY;[JKO]MCI888($<+H%:V,J6D9> 2
PS\R,,7;)$:]:G2%;UU,YBYY078JX]BRF*\(F5U(?MC%[_-A3I:[XH$\E,AK2VV^ 
PKILLH>27D%BQG;TE?.98R!(9:WHC1<+V*P.A*)*'=\"JF/XJKOHHQ3.PCV@91>$%
P"7JXWYU5@OD&BENY0W&:ND/'V/C=Z;_WCY"^"U&!X(B>-\HQ;#0R8P,W'[G868/;
P_;#_(U)P1=$?&3!*LV_#BQ*75K73>'HC:P$)L(:'?" R%'-:H'4Y=_/!?[B5>@J_
PC1Z_)"*J")!Z&"@BJE$]1M)^U'GI*6>81OSRL9\ U2Y?3LQ#B+OU]5RA=570+1VG
P6T#T-LD\VCM5R=[BZ8## TV[R69V106<@U,K4 !#_D]EQOOG/+%1%R[;]W03CL7'
PSX1KW%$F,L@[*O_//PCL^0U-[U)QO! ,#S,EZ"!LTME-$\S3PW!@W<: 38J^%.%2
P.-"#@W9_N."!$Q34@CR]=D=TD9%87=Z9W'1',<K*8\=V7>[E#;Y=55M:Q?@&?5K$
PF0G&589!HYIK17M,E'8(]AG\RX W:Q^V?U-:N1(Q.2=^MSR4?B>_W2GB@1KIL4K6
P#7LDL(*!>_1@S03 7 6.37=LU0FM^!LM;"H7*^PAJ9FW1NO"^\KK>;B *3<EI#Y?
PCD::G5,*$^'G/>!%COPZ8#@'G%O7-!([@WZ*K;]Y3_A+XZ++266%=LBT$/"2/DJP
PTM'J9?@^QLUJ<>0SV,9'&BV/>(FH'-]HDZ<?P*14&20E001'6;SJXS@,M7$/'!W[
PD($0DO<,G?BN+1/H!-,Q9NN?B_.J^50YK1IK*V]DN#,Q*+V)?D%BR)7GEV9[/(M>
PC;VH+3F]VXR"3NZF$79X<LSHEC"CY^J8W5%9P?,>?XJ%*,F(!1,EGW$1]FUWT+D5
PUW,.L-6Y'/7816*$Z7O//'=6M='<\X92Q:R4(EI:WMZ<5MKTITRHUK:!B$4X*-1_
PU8#<BMN;Q9CLPJ%GA1^8+-67QEH4SY#<7^>ONK!69I$Z5&7I9(?3%YB#Z'"8WL&Z
P;HSP)9!\RSV=*?KP9*K2)$Z%H,Z$<#]GNX50&09HR_R0%H$Z%S.Y:5PH 0W\KVR;
P]\9QA4-K9D;4*=%CYM/&%P@79*IP;,7'E@$2$D4% ,&G)-'71=B4F6G[>\="6B7$
PM^#<WP!L,)SMJ27,N"XE&%"2()0T"G/P#3;+%.I0^'&/AY^@TR(K*.0I C?LXM.\
P/*@3J=]].G4>[LDC@[LU4<8]/);:*I83O>G-$FZLT.7_=8205,MVM$A>K"VY\S%E
PT_-15[C_-27&[ZQ;[OLYXN>^)^YP_+I:LA$;])],E2ZK-0"!:@G<79>%PJRW-9NN
P[)TB5ZOJNO47HUKLFON5LZV1I/( /0>_P,QJI3F:U2.,4^J'\U>9<8/E,V&<_ZNG
P*6DG*B&]TH3;BCQNB?"> $\28>&5.%B&#[(OD-R<>05(LM:2=C7]UZT$>MR;MC;X
P1@JJV!N,4D07A M(G^I07?J1[QV8N,I;),,U-MD$#$)7P^B*PL8G0A*AW5FH"2YY
PW%DE<-<%$MO/^<"7^MTH'>T)<*S@VG :'VU>E9-6 *YS?'Q%:G043M%WL&^8W#TE
P,@3[ 1-Y5*V^@$1L'+B!\3[M@-;!GXGRMA=57]KALW,25QC,NK+<N*8I/Z^3(_-V
P134SSUHL8 1X\,/8D7'9;'K[3:5!;^>=H =,YI83<"7+QZ,QN\^:V6-A/R;U]UW7
P M,!2MJEWXB!=W.C7:'M\*J*M]D&W8P)C4UBK =& 4:DKA36IE#^>VXZMK=.,3+Q
P-L9A?#B3[(91I<4[W1U.652.PQN=5LOYL5Q* !MJN49I'!N ")R<MI]+6BUN/?$X
P4N+UH&K>X5(?TTV?DS%N78XP8%G;+[IET-9*09%6OE*X%A/6^]QR3WE8^ 2XVVZF
P?:QJ &6%@V$O-*W&KI;.X5_L%Z2M>6]%ZD5BA]LC[L_;TC&2>UG1BU)_B5R"T8QN
PVCE'%7H_4N"H60BNO&/I+_+TN#4._'DRD7)RXNW.NIK)1+.) L[V3I<K+H$OB95!
P>J^EHA5^P->JC>;%J3>3YG?YD2J$&#5#_VLP*YE>&3[<[4VW/ (H;O(3<?.ME?[;
P5GCY??QLZWO_!-GP5]L&^/9"&@0%_-?$8'GJ+GZ\P.+"Z#AD496.+SCR*@9[GOBP
PW[T!ZP%:GSHHZ"P!><B/-M86F%Y=-#VSKTY]Q$^&E>$9 H2/V3<F:B+ZEOYBHTL;
PI%(W &@6 )7V$CRV>JO%@#ARR_:V>J4_4*%QK5E69]\QUX2\Z#2!9(L"(OMBJF[P
PJ"7*3_\WU&D9R',! \HI]D2T"];4TC,@UJ:D5&GGM>RGX^>WOCUEZV(4_8VR_-,>
PC3B/?QATYL>\CL*V<WF'D(X4,!4#&G+^R, 4*)F][:3?M^!!A))GI0'P.O$#=T.\
PSW?87 DH:6+Q0K:([ BT3!Z;"J5_',< T0DBP7/B&D=E8U'T3#_3(\=MYBDP;X_E
P6FRI9,A)1&07Y=SS7S*8*NT&O4'R>>S%0FB2KJN98D=U;OF3')_3M3[JJO?IAY-U
P)"_J*NG#/% /QG8(MX;7$!'_10#VQ-,U$H.TO^T1.LIXX%-^E)MF^PD]2\A%<[^S
PA7<;V[PZIP/<^7F+@'UKCE*]&F=0ON*J1G!^!L](CGWZ"O.S@!5:SG:-SRAN7ZJS
PPFZ"NTM[5)Q_V5?[3_TVJ-934:7_<Q8#2*E@"G685J<BNX9R"U:AX8-"32KP.4?Y
PSPASX\1/H(&&*UNM"(PF[:G8>7EC$2X(I->-"W)E!5-.@.NX+3>Z*B\Y8V\-[9I\
PX9!;K,\I>U^P-A6#K<D\&06G^M K5>0EX/Z_5[:T/1"'(E[^YDJ05VD4#W-:^*KV
P %U084K7RW[+6A<AM7WZ!:>HT$JKW-B+GW?,[W1]@;%O@B\;K+N!C]E\E7=\3J,&
PL]IC4C6[Y78T''_'.$0@Q?3)1:4@E%VOHK=S+IOAKK&/-52UQCR<LR;@^W,>5(#*
PS@2TL]HWC_Q3N0B 5O,0W9245^L8Z 4X0FQY8[ 0&A(FU'Q!RE#JSX4[3#J >M;'
P7LAG31S4CGWUFL^$T0(#.3P5VL=[7)Q.C<"I?^V>[LA?K4Z\LM]XC5<UD0BZ1_IJ
P\HUXN9TEL5:$W>_^0=N#OB8:B]*[]QB!ZA#RP*1P%E&*'!\U<NEZ\<OS1CG'_]*P
P\'?]]3C+3U<@[HA1!&<ZXCL ',$9-&D(L,+^=87^_!'K1=G17'D>)*?ZV/1ELS%(
PU/WX$6L [Y4UGW!%5=T38NA-#(;:?&WL(0=0T?[5+_\-.7;3P]O0 ROYBTK'P=)$
P9($5JWRQ_Y2&6@3GAF"DC0NQEVTBTJL>/]^A7#*>W+BN!=>4%7"[=,IJT"(7IS/-
P:;[H>-@.0OPOO,.BQGXZ',2O 7;/P7')G,#]@BKU=ZM,O,E?NZ0)(WLAZJ0L/>F.
P02,EI\TRN;3O'QTTM,M.UAF7LR:1.:!AIN'E*X^H&Z_5%&KT'BL Y&M(P=,H#M[;
P;>CY=!'3%%[G.PBAL%C.2J1_716<@C2'WI5NNH0Z[Z!O<(PL$)QC.";C]?S^_T\B
PXO/H"MY;&.B 25&BGV7!J(XH_^H2[329E"F]$#X=57D3ARMJWY?SDTHU6HPGX6YB
PU9Q<O86MY9% -"^NPP#QBRD]=)/N\CUBK1K;O-5*%#2+W\R)_+/+E@YU=*I]V-FG
P7MN;_GTLP!:.1WK?[\AXGC1UK?CNWJJ.086;3[HN9#=W)G.X*<_?>[,%$5?R&L5Q
PD=+SO+%U\:%0LJR'0]5Q>0XSKEF9%D(*_98PD>M&1$OV8P,2HIGE)_ 1L+XGG%7:
PV(4:]K[/*LLN7F$T>8O:Q/GE"CSFBN%<^?!3@'9)H!1MJK5*+#M6D2230 <Z^N@D
PE4#U4<I%)C6=3U%!;38"IFB(?OT"8O-059%F^Z4ZU,Q1FRFS(/=/LP8B7]0]'Y^.
PVS UCP%>6W%C\8&U, \[#AL$(/@IU@GNTUZH&[#8VJZ%(;15&E897P],>.U-V#!*
P#]E$=FJ(VW/5[])V[=UL9+08Y2:)>J$+L0C1:; PJXV%H?4YB@1Z,D,V7EB8SFYV
P5O(Q?'>@['5P*,Y)=[$DP/^DZ"H'\=*$8]&?0^@4=GF\'=*7*X"DW8:$:[?_TO"I
PE^4%GM;:<2A8>H^DY"01$/7@:]WQ =>6\+;3Y3V *J@X,C0@E2#VH(VT^"/L:_E,
P%]2MH*EV%J9F,Y'B&4^S;&9)%1#%,DD%&0,,KM>SQ2ZS]D2$-'E6@%M(_/)-_W0#
PCT/+2IA@]/8F4#<!8RJTJTXK'FE@<$^N_I$L*4J\5DIRD;MH@=:BV3B'7,[8II? 
P1B?_?U#>Q#U64ML @8?70XAKW\ VQ7 $4'TFO3S]IUXD9-AA> ) G#E1TI>,1'I+
P,A25:+DZK"4',Y?B&<.#3AYM<[F^C/*+F[@S9Y!C1,H X( FS6>VU!+^[]5?A4_#
PJP3O<#6COC\Y#.TRC?57/LS7G1U_V:/$81K&XKRZI:?':@X8@QHF)5F<S8K*51TL
P-XQFP9U3^37ZAO[C[DH!]BL<"Q3$X]M:AYF[TI7T&&DTVOJC)3@9IP-8U50_&A*(
PIF&%2T%0D,G-*A.#YV&I?9SW;B0NCU"(7A9CL<YU&K0(^DAC/9@BN6_ 9R(I,![ 
PWPF:S%1R66?@5IARB41]@H6%XI>,749F7P4][M)R4J@CL7+I.%97J,'<GG(_Q;+2
P&^,9#)?C7.7J*6M)H(\\U&+6J[*&:MXV' -J/T>7FL6(PXG:9<C2EI XM6SAC(<O
PW<2.]<L+E#U5+:W'1=]YZ4)][X+X7%/HGE$S5UW0VBNH/ 7>Y@YC[VB)3PMEA'H)
P#F3$W6S0&%C-@EH]P0"U6*0LZR1H,3*GQT1[*3X5PV#XY_GFH:M88 DR+7!36#C3
P$G)T]]_K#\R(*_HI0&PJ>$,U*"?%^*ER1% 8P%I)L)5N+D_5H4J\+19A:&3U5$I<
PZO0N^'.K583@L'J0Z G:Y]39#\6G%[.#6[DO=00-PC YK.M;#+6<XGLJ^^COT=;B
P+D2 "-6I:+^[1_W6CY1,*5OA4=<L\7B7^_UA26E&56<]=0#JR)<J15Z@W>HNI]FJ
PN;ST_5KY4[IAP#>,G(V<"RBQXZ^2]T;O9CM235<@==5>GZ,]X1R%=55X6WY)'(8'
PWVY3(VJO98Q@G(]<@-F573:4O&!!E!_4JKI*/P630,ZZKHJ-@9V8T'\D(\]XEDT/
PK[N#U\6:@9>/?^ZW=:?PM-<S3RXUSTSC%J=D3PM"L2? RXKD. MQAU8*M<U0D9JC
P-*RL9;K:9^YKKUO DK2@R'W_$XH&FGK!^9,8%UA[[M=G*?6'ZB,7LXSE%=53\N^3
P*> !5%.G-A!]!5*9?AI\M-=?'K\SWI&YC)K5F>C_>$T57M]XH!&A.PZ)C-J$&1QE
P.R@&$PVQ"$3-/68P6$]I1BY!^WV2-8 /,B6Y9.FKV+G!B\'< +825&:N]W-YYK)Q
PY#'5;1JZKFFS#5MG^>$1X6$GCO>0N\V';Z%H=LO$2TK(!QJQCD,F#Y#TW#\SKBT#
P2Z7AR%_&D_$B&"$66,&?CEYZ,SV%&:4=.]X0LZN340HHK )@$AE@N+-Z0JIO1[.V
PA>WWED#99;K=8H",#?&$7,$2D<SZ[DR5O4&GN,"+'4F8Z]Y+MCOL#C<1UVG2^,PW
P]])^%ND_[/;U"FAWR1L=K2W/,(..S&8IGSN^=[3[ O0H=\K>)X6O4TNA3O42'IH_
P#%1?FESE564WEWLR49OC#[IP4BH*%\U]HI,_>Q7(-')\?'(7U*5A,TCD3HBPLWO>
PY;R;9],:-Q-32P^;X%?F@\'N](L]\W##M1+L)".,M@R-T1 ?WM&"!8S-C$QR(CV,
P$,]%VP'90DC2NHB4.] $^JQXONW!"P!R_R=O;B=\&PP&LZE>J4?RT**K'B\&-QJ+
PH*.KPL: >H6".)VS-R\/H]()0X<:T6]=)?#!'HS1L"9.T@30E\XP[ZDWO\EBAT F
P1X-%).^:.IM1Q=]N%(=R]O+HSTQG2\0Z%A1B]S=U]HW5_C=8^3P[X$!&W5"5T1#9
P'R%XU>U++ \\N-7EQGC)@H$[<VK46%S,*/YA&[Y[4^D3UATG#07+W0GV"65Q!Y4C
P3R@#PG81P8P-]CY_L$O('[(,42)M?NPKPU^V(;H++<O&:R)Q*#EC!N>CJ^S.E_U<
P21<+"$549C^7B++G#>7 H,[%0"Q&,?CNM"U'JL_\$=Y'F(0;P!"<%[74E;:('LSR
P=,A]+)S D7?I.EYU#^NL//;U,D6@&/H#OUSJ9'!L=X-;&'N45&IB\7Z@N C?8#Z/
PF,=2G7V9(81FIC<_?T?T9O4%V$O+=F?H6D^DXR.&P6#O\7"##VQ<G9A"&T (_)_?
P\GCZKRNB_$K,F(>NN\ $[JG4:6,[.3O2+J++0OJ^?(4+#M6J>I45'[1L(B>EJWHW
PARYIL6"*MVWN,:DY/S>ZB=A3DG?C_XJ,3":H'GDG#J'$0/8?7^_G\5(S&^H$(,$=
P6,:M\<'<+)!=]A+AO<W00SH:I^R# E+#=\IHEUX]2 L].FTRF&45&4#N4()/+9N%
P-P'V@72Q*53'JQ9C!D//]*U]9I=J+$\XD'3Z25<.+Y?#TX-):J$'V;_/J*/*!=UR
PDX$3V?DY&,T+ MEC_(L[D% -.5WZQKG/O+1BP+N^=*LBL_BJJ4Y^84^3<*XPA+TM
P29]HW\8#]2%$ ]N&]M6SN 6".MF_;VQ2!Q#K^<Z[_S(@$X;7@&]>GHD(*\4S]2+0
P*.4^O09RVQ4]^_^0 4]:)3X;E *=!T$O9<;*^54#Y<0T&YLC[TR,9(DR57;5YK-<
PVHJ;I2/50]<0PY!)[YNS2"R@*X+4.>6ZW".!U<YGF9'MP,72%,<@<L=0W&I";QU)
P[]=!$2ZI:D<O$AL^/I6'.HEU/!9"JS<")/% =<;946/<^1VK]?AG>6E+F15\[AE,
P)5UZ0IX)\X8MIS0WEMQ9"SG&O^>2>EE@,G#">_9D95US(MTC#&#:4YD%6>FCZ"*0
PU5QS.%_'S.T*W^!4L./AJ95"5)*#;S>"I>A?;:0O3B[WBC8_M9%N]4IYE9WO[,JA
P)]K..%[YVK,3X8]%)KZ8H-%ELO]B::^&,LU[*1P*,U+ I\]WSH(':)_#]\[LK6VE
P949OH,9J34/B7XBB]+QM_ZWXLA;Z9@**?)6G#"U[P*1?XG[< BJMWA.Q9FDC/?3 
PVT/M;@ON.>$9B$?=PZ>KI3FFCD2WJKT"!>7<EA<_S%Y$U#EX5UC%D9:U+^>:B$EE
PS5MA0//8Z0ILFK\B%%=\86S]Q%AC(!:XN0+M1=L_6).V_RUH_U7TR&O#".%C)BQB
P9KUD98$5U9H%PDD3BDU*LVL!<E2QXZ?$I"=Y-.%(<GU\XQP8OM;#DOYJ.]$*L7:+
P;O J6\D3C*BFH=F2HO19,K)^??W1/EDO4=+SZR+,O(A/R+#ERJ.5#"X5/7ERG'][
PE;-^&#QV.W^R'15%5\!8:_JQRF#OKQJ0#[5'UE$<H+/)1([WU?D;-*(-TH.FH>H*
PS[;^"KJ(WM<+9=B"W3F5_?^5]>P^:,Q#Y(E-T=(*.W)C.8Q]18UF4?Y)&C.);9H9
P6 LHVM]I>.*ZFU70Y5"_+HMS2$[BT6: M4V=?0IP##AD5L3UX"( TRAY8QV@=WKO
P<B^@FZ5Z89D'=$0O1/3!2NO?8V2!;.SPW<PTC!X)]US95$"\@=5^REV=;_+P:/R>
P1._>61D=)ON18BB"JDYE<ND/R'R$/<P+K)M=+Z9X99Z;4DL7?U+UFE6=D%0@0Z5S
P(UJ-:\BB3!?^$AN>37FW86L?U#.9 !HFJL9X^<G:/ [OG14^ZNUI5Q"/\N5#VOFK
P:%M]@#VH+$\2CN85:XMF+PH3^T?=6,NNK5:,V,J?^J1'$>FC_$[$4L#7* T9?XXJ
PX>SR%>BD1G-T).._$: $16\60>70-4D2YQB?#4E_YB=:=&E%@.<YH2-7QZ3Y?P'V
P_,(MTDL''5EZ[E4M(Y]T(O2#6K,J0&;"9Q)+"&&M/O??-IT#\;\N[^;<SXK#\Y,9
P-:D]W:(MK>7LSE[9\\1$?/>)I?C&>YB*K'V$1O\;#_MS-B>MY4W Y2R3G%T4LH1/
PSF7,,YJ$G82)8!4GVPV@;T/N/I5VAYI-))$(,Y:Y:+OUK('_C*^#]?@H*Q)TKFA,
PTQ+G,#*W]KN@']_]6&.@.'9Z%S9HWNE!EQ;>93T,D=>FE@WVZIW);*GY+)!3S??N
PLC!283)W)1)9#DH,DO!!^A'>2IK=S3O_L4!HE4;$Q#9E1J(Z"1^QT/&R5]:'_E5!
PURH-Z!\$PSY!"XLR0MB:LG7_E"'3+S(.(V:5'I,0YV^?M#;, 5IA>7_/",,661#N
P7LHPIGO<9.R;.EVS7=<<ZA>W$ZCY+I&4A_PM+B>J3#+OZ[??O-'WNM"BV:";ENH=
PD,/.M.8(XIWN<^<&;R4A=;=W'S-JI&8^YH""N2R\]*96)WT7!KGT4?%OGAM:K)_*
PL.?.OP()U,BZ&!<'XY9@2&F7,M]_B;WV)E.?UZ-@;_ASJBB5]F*46X&+2';1_7Q6
PR0:'\9NG# S+TQZ3D_][ NNEDQ,X]05SBH.Z7PP]8:BL;M2W(27*-4O^\7DQ#@00
P),W\.-:B'/_O;KYZ=$@59Y-6)T+X&L4HAHGC9UUL0],5N;)3#24X*[5L_0.,'CO]
PG4) X$::;9CG4;"[9"4?LKKYM2B6K/27OXV[!>0DL/79:$)DB5P<>*BO_H:Z H$C
P\/MR0W5IDR:;-I...D4B!&CMFMNFQ9"FXQ"3#-Z",#(( (GG_F=?3/G>"FP?H 6W
PAO/L,*+)4T&7)!P:5G\U4:HWFNIO3ZWS?UAN($ZF ?1. "*P36 YSFPMDKL7%[L&
P8A*=Z\6 876[R\]RC0XPZS&<W&N=-U2MJ9@:>\G%3/'Y"?3OJT/:\KU?2$5M%4C<
PPSL6U1/6,6CULV9K1OG=- 3AUM7$_.YS3 9*F7LYQ=*%=>J@I.\W.IV;0-Y@\5RA
PGG)/9K +6PJZ8%7%8S]=Y+9]W"M/'6*SZ)B)(2<942"47NIB=?OHMT,;&X89U*V8
P!FKJ+];$^<P)JAT9XD9*5V$M /3F<2,)3$]T9^PH"'M5Z""^5?PP*@D]<^*7RBN3
P'Q61;^*@1&31*^IXTG<9VN[2FOM@7VLO3VBNH[^5MG]"4M^08CB0.?,NZ@ '#$7B
PUS07]L:C=>KB)_)4M2T5J%7O>FZ4S,6&@ J <-@5329I90-FOH>"Y(W VPZ'P@[J
PMNZQ:#T-G1Z[3&GS3D1*O.=XW;9DFIB!9[!WBL- O\99 #_EZODRXI"<,ZBN)$^.
P(C!Z5/Z* V8&W=M4Y/&P,VU755"-E+B)F?S)D/R\:BIG/*NTM^$V\;RX/'+!A*(7
P#U#7.&BBS4X?L,']0/0J6N9X''D:)P3^E&P[*9*Y( ,3BH)BY/Y/)(WRNS]5XN<!
P>;@G?4$B^*0^=Y0-O:S#K8.;#?/E+@7%>HPO[/1N_<*;SE,X\M=K^CX!P>X(FHXZ
P1U-HRO4DQC;_!&2:8R??1]4_K)R)KZ,[V;AW? [V$Z(VGHT_ "@&:1;+Q5*(=3 I
P*)&UFQHC>3:29D> BW9%(IZ9@L PVFEC <Q5(D),.DX:.8'UA,N2ESZU!YJ_7O#*
P%R35XO.9;+X.L8YCR5D3^U_CS]'.6^)[D;<S\W+&CHAKJ6&5+\K#!YRNLYY4L?2'
P"@.F^%G0M^M$]IL?)>\_N"?VW?-G%<MM7K_S-"G"?/,TKR[MJ*Q=_K"8;1TVCKFU
PM0!X#[0"<)XBR!MQT,'VA/O9EH-(..L\)=1T<9[:#&W!U[-Z(V&B;*G/2!J'C2% 
P-!WY7=H 05F-^#ACR" ZPQV&JVR$!4;O?IK?9$XC[(</X&DE@K'!>A=IQ#N(Y#)N
PRPBM7?M?T%0RPJ<;]AU18(.^>96X!3%S1NI9@K+'3E,Y*K!8^F_1>5ECBRF<8F3$
PWT-/>*"L9L-V2&$\V<G(N_#^#5'D!7-T[-#".DKZ1,$9M<(<:SYO(]5X8%?%;2G%
P2\'KJ?OP@R: >]JAAJ6S:!J,<8\T9X]5%T6KQ15'3YZ^L_4X"<);%K5Y^' V8Z]*
P- '7.XD*KIV$X6?VR:,-LZ^)&D.@X.S8A;BFT5<0M;9$/9[:O'&;TF[;*.%=L83D
PBD"!VP#;?@:X:T0NF9PA*L:><;<A6&?MB&'(39['FWQATE) -4A'$(9YHETB0//9
PHH7S&L(W4\Y(^5O^-X-_I_K(@_+=^[:AUW]-DVJ0;#@H1-V1=;K;Q(H$)N3?X++J
P""+YA=S"790(;Z7"6FA9;XQ7G9JJDU0UU^O^N.LZ#D6K/)W<JF#]S.+>QY7VMP*U
PW,BB,C-7? T?*]N?^,'#"0=%C- :%L0OA94K+5GBF8F&HI<+LR@UR0>P3_(GZ!*J
P/8V'K>?AB-+&)N&OG&4&2>U1L;R"4,WP,\/5C1:XR]9[J-"9@Y[__2*/UH^: *_6
PSMY^2DP0"E2+Z0+@(S.V,HR,LS"6Y#O*%> O3+2/3"UZ&SHK&#4!6F6#-M1I-J2D
PZ/[AN)5:)0=0C"0(KO9AV.N< ?5F\DF!FB?G^?<INV(].#SE14=TBO[L(LU[MQ]F
P)8!*:HM^.[M0.4YXBK8;&>[A@[CR*DKT>B[P55=68SA(=N]AP9P$^;EPOLZ_8_IE
P/BN&P.Z^3P&FV)N*/X$>$XL7Y6]&DM70R#3H^.902&+7&GB8*H-9?B(B.NAF^JR]
P[P7\.A7=B&2ILZ[*FU/-[(M5PN0U$BIE6'ZB<%IFS@'@BDA<8Y6T%INO[./@32\7
P[OG[%=H59)M;J*'$0\1."](W(2ET _5]N:=_C1N-,[GIOLX[]:1Y(G$5=ZB^W44%
P\ !=*(8:9?XY+?@8'9"4=D\//H'OQB!L0<D7$5[+,4SQ0:F6I4T>/O\U) -=0C0*
P^%(O_QXF6')ES1JSWES&/D3?7\%O! Q%=(7O&C/SKE^9BJRU#9S,A7.19'YTD>A*
PDOJ;8HU9"8VM05]*8@(E<&)9_JC(:_/,)A$HFM!>.F1XBD,HBB$X596MO-V5'J^#
PJ1LXU9WCO/H@+O]K=)V/7$Q-;T1,6%[?1A79?/FC@@&A8SL++,ZOIQ70S=V\Q.4T
PE5* ]LS'Q^%Q*F-,W9&))!6>@[_GB7P5$)>YJT45Q\J5H'(;H#CTV'.3@,G(3ETP
P: \%A#?2WD/%NFKWQ;,R0/S7!%P%_*;B[D]/&'6&JY9W0N>0)37+W_%X&X"*3J*=
P.)!K-G9N2_9 *$@5552WQFM,Z""<'5&LW8^;F%'D&M/O/$UU:^,\C:S)*Q-A5H[,
P83QQHXY\$2:N;L$^A6P>_/WH2F$X1>)\EOTN(^RW$JF>&/]VW(Z7>'WC%AP9)8;W
P+1<2?"EK-6?8RT>^2D&THTV!J!NG]JPLE!Z3B'PR;5E5V8KP5S_U,LZ=9YO]GXK:
PT^1WQ8<?4/72!/NEB.J[:J!))1]%ZD7#ZQV^)#'RU7:%42DGC8Z*$5!+0JUQ6'G8
P2@*6QC9=4,*K+/%O\IY,4^;,+4C@S]8P(P+L4SR-HID8;H21"=*<(0/;%-B[M<#2
PV!)'4G71-:XBR<E.^B^6>B+-; >%T%'G ]2X&7^&]N7N%-SS-O6"] BVZF+$)OG:
P9!DSQ"N5Z%T*]WN2I1=+H1FZT=NM3;#(?"Y 9=6=1PW3"_"W>PC/^$N3QHPM^7P,
P7SO%D""@CV"RX_TY%*2R32>'=T788,:6C?G@^IA@T?M$]LJ?/>X0VQ[9PZ^!?!-2
P9TEDK5DB+V#)5X:,98_QQ]/*.6*C_LA;<8V ?BF"E;9;&-W^7DS94A,\?U$.WONH
P*+1(%63E5C6K1"\,7G12%U+2BX-Z&P#0YLSB$IA\>CPKF3.0+P:F4XBL@&EED)C"
P8PA&]OIG.]N\V.%NOU2UQS'ALH$7[823@3$J0@6@'!WEO\2H-HS4X0D*+IC$I^YH
P;9O%CH-F.H0:2((4G@2= =$.UZ[2_MS5+$9Q^![PG+LU(*N;6(83 A&3M=OD+$66
P^*7S31XYIO=: =X"_3*MF!M'!8#H A8D8>WA9=^^0(#+N'RE? T#P[B[ON,DU+0W
P)XW30AD4O@VI^(YG?=!8_:X+\8GG"T8I.:">4EJL268W_8]78 FPLC6[)/.;QO/7
PW<W_)ZD(NQ"C:P\0$]P1J/-:,DT9HDMW3W(2HL>1%-.L[2T<UX' ^07R3[<.$VT-
P"^,CGR 5).%ZY*S*G$!'BIU!OV^%2MM'%(1_&"L'>ADSH9NM4IN:Q::\I7G^DJ,W
P5114C#[W1+Z)@701RH$X1M;,&F5AKBR^R]G5%BPAPB O9^.%6XD3=N]8>J#X+-/F
P9YSUSI*=;#3H8.N$$4@_B?VN*Q35<8USH#I["@;D@A?A7?%R5Z@&NX-A')PP.PZ\
PEJB43058W0:A1HH.-5A5S)NG*9KWA">!#AFIQM&#F>+8F],H.?V!KB;L/28F;C).
PH+V*7DKR0 #/G 0F4*%?W)^2S==6_)AT]'381CS_._+J,+\U@VQR$WISW#HS5FI;
PNJ_:U!-QZ!;30@5F;EDJ1].P=9C'%8I$P:-NV[?M/-7?HJFN;QK+50F*=Q$]6SQ,
P)%FHD22<V(#6[.C9G\^6/C<O?2R*LZ$IQTL'J22;@"\;<<".@J "/ X B./SYX# 
P5VA70\U5=1GD1BRV%I>?C+B<6O<.L?[[PB5'*JB*O#U;B><&!0L2#7W+C?/OX=7=
P:X'YY$N W7"=G;1?,2ZM3<9+(XHR\1"57S%>.O3'&N_>@$TU.N*Z'P<T @[/%OKU
PL JL(UJDA$*'@%Z"#:,NJ0POY^6BQ'YL'L-MU@$L^M!^2L\'6A#G9,QR;Q7K/!8%
PBK=T[:S&JJ/$L">Y=4I'>]-DYM;?-[;I?-#2LN(W%)C./XB2GLL>^ ^K_YS7%^&)
PQ_=;FWYB%8H]GQ$4_;7>@] /_0E2N!:B[(K0447%7 /G#*;VD<)U?;^1Z@>S>"DL
P$!S1U@.=-QC53T*:?Z#NP$#?@[WR>.)X5.W[684;_UPRS2I-4PHI'-GS-=.<AY,!
P&54-]CF]17!B:7PA"V])= HP_>-\^<5#VPDF5A2H%)VE*PV-W';PJ<FA@$JZ/%N)
P'S/&CN+FX,9I-]ZZ2IV^E&=[V<U6]-;"K@_5L&_<]H#Q4_Q0J&9V<IIC,8;GZ]FQ
P,IPAJWNX(3*$!UWOJP.[B3EG<9Q:8^7X"+AXGVZ3L22G3BOOK2J^1Q*"(>M/K3:2
P%-C&^QM\P\P\-?" $AX;IM;75J:JHB9$9T&")$+!>%(7_>8R;'9?+(C!)+62&^2;
P,K[Y )W+L. =Y_11^CN<'7*4H7'LZE4ZZU))*7AWD'.8!T1>"079URG'X^_F#?RF
P  7$26)Q+C\U^;#G#,2,PT+:U(WV%NXR=<>F>?8X[Y-Q.3<<N-VFW3C NHX*;I7D
P7G"""J83 ,H>'))>YO(T4V22#SJM*ZP?:U<N#SDDVBZZ1L?/3WI4VGOIK>N)OQ@O
P81%)/&WJTH7_@F#SF$CV,](T_QV]&"4*CF8MF0J."WHQWKE(+T^_]/'([/;2?^/_
P1- %":4IN/QZF :O(5,>]72F"DG%;&AC7P<>(-$A)@&=QHD2%MP)9[7[*M/<ZH..
PA3G7SII3$+I@^A$JSG3:="S;]H2<\D32#R6^-]YYJ;R$33BJA:6I=[4R?S"Z!B/:
P@_YZ@MW?N=J7 B$L&40"E"H]#G]\ZPX56,[MY!/$36K0OCG@-O8+Q4H=%Z!268(W
P>J\C>&LHX>^1';! Z37H2/SA(XG_WR]&FK:D/TZ!N0-M3_J)TSYI6J9%MP-6K1O#
PG=%D85">G_</G#KV8M%FGK8;]_K@7Z?=SN<F!'0(#0.[EY7E&"+2<%#^]YM>0+C"
P<A<C&T?CA'K$UHK;&VT 1ELQ#8'^*?Y+2RL?19[>BGNF+\2766I/$&_HX8:F0U!+
PG3O3ZWETS=S ;"S'_4I>-6T"5@.#3U@ SLW9B-3];_/QDTR=VAI(-G4 XJCYF#7M
P ?G+N,?*HB(A"U#L:_6'C6K$,13LG'50RY0.>!U!=]V 5?_QJ<ZG)?W,GM$C-\*(
P6H!3H%PU5KS^:"@$OLXW$8E*RZ[9:!>%&UQCZ71I"<)4V)!]"3E:Q 0>T:0@*QO/
P 3GN]4?"7!_Z07G$PT7WS#KNWYA*T(O0 /+4[V-U8.+P$-\,VC@B!,$\?UNII0P^
PTW/#XQXYH@K_@7\5V;]B-M]+FZ5T49F/R=G+/]6:P>@HR_E3Q(D\SM7&YDMF($NE
P)GTKFR(%9N7.]NQWWO4*C# %0(-5!LAP4"]69/>0HBE[ZMB-[PER<.Z&"";"36N,
PNS3J.1HL^5A+%P'2GB\7C#CK613L,%\E[&#:WVU?9KO.XY0M(.C4#W*4/F;I2M58
P\Y";VV^H*J<F@4YIXG[6OC#>OGEN;PE7#"E5R=KE7)WW\7".I#R^L[&8QJG!/1#D
PS]85DVZ<,>PT!5X%G^K"I=L-HKEU(C#O)_F21I(=,6W4(YCAI?&>^9M:;QM-O%Q/
PYD[YB)K+*&M:ET@.SL 8(H*F^F?3I=?2O/0:'5YEGHOHDB%81I+[D)B_1ZH8=W'E
P8C6N+36R*3K-GJI/;F =MV>\9^Q4JR<U=V0KO5#OL/,:A(5Y%P7[[WCA%90NB\M"
PV(;M7X_T,S0B^=&,*-AVM\[H)(BHI'*^_SN;3WT :^Y)BV/?13@9 HS54E6$6RS$
P(WTL' ;T_U)5ED)<:R@X>?>ZKJ%/V'VA%.8GJ2FP>#Q^*%=^ &2?"X3UA>W2D)E]
P8Z_3$@B/<4_"C+>A8?6TKTD9BXFF02 PH?X9T3(Y/&Y(FKF?Z>6N8:-*MGBX46Y$
PWU.#5 9I PQ<JAP[T"")[0^%SKH=:3%VV[7T!-0$SSP;P"F6&(':)FIPX6$1@P_-
P)2^K6QAR^,FE,_NUN#[5"DQD>FXHY\<''6!-59Q@^OT-AK[Q*R?164+>RA5JPD'9
PIEXA$,J8!+(46A=6$"C\[[TJ1P26QQQVSVW.%_E2>2:$.!>0^@AVW=#%V>0Z3P;Q
P19?.>G6>NN$")7^ 5E/_GW=_!R?,+-DQI_%$1%%-+:N_@(%-9NJ=W&1MPW ANE4P
PC9\B.8'_<UM7]_VOVN"X112E@7TL0O.YI,%R.J%=V^&G7\GY3=E,J].\ND_TQFHQ
PO%%-EJPG!;#<.@UPL_M+&6D:)TBI0XP%QAW(A</A2)VH"C_QU$."-K0+4OKW,G$M
P.)FHU0+HB4A^@ZD]V)QDA @D>\TO343&).K"VJ+T.^?S[)RN!X-CR<N).YF8$Q7:
P2Y91>^=W7EXV96EKVEB=%'J22(W/T#GI*O]VM:BL$R6SIZ!UC8OT_/EFY &5?_?R
P%/$<_+!'"5/0T$GBG LZEBH!F<P^#KJZNW>N4U/#B S@]J?LGYHM"\J)A>O  D]C
PMR]8/\5L:_T S#UM,6%Y*YW^$M=BW58 )NNH+ER!<RAP?P4C)X/,.@ 916ZOUJ?Q
P:<?HPH6V((GHU6"?\_UO"\A3_1ED:CZT<76QT0^C+)W2WSSQP=WCIJYTP?4<45DJ
PV3OPL]9][OWMQMV=9_DRY0F5<MUQ()WF5#IXR&K_BELVOC')MWIF> +:?0:]/,*$
PBE-ZJ%TA@H/I'3RS@W&BKL4G=BX/AZW8LQAOP(&Z$T?<>U&2>/Z79/>N?CGHP8Y+
PQQKFG7]**9R3@LNU**JH\3'54BN05_KB5"C62C?9$7XC:A-+4]<WP,702 +H$P[>
P[U;B04!-> R,418:R]3L;]1ND$D^79PG*I>,BV ,*;ZAE$D9KL($/;H7[TIU>P,L
PD$H+. 00%<5TA%4<ZM@T:BE["Q2>L5QU_['C,_JV,+\TE 10OY?X"KV0C+F6GT@#
PM^]4\BL+.GG$A(RV]6;$M..9\DS=E]W&JR"%>=:SKC/^E_JJ":8:KU]';![U9^D)
P0:K59W[8V2XNJ]5R;RD)U^#AXW=#E:G;0/G4"NEOZZ#<R8)N0N>APK"R;;GJ#OVX
P:*D!#MEIH\H-3%%HJ&C$!4T_'PO+K#L?1^M;,$#(E1!D -0G"*C!)T75TM/9@V"\
PU;5LWOEJ,!XWGM'YM69(>36!::!^PX'&G%5F-*4IB+X\>$<=/(=U'$V\E$TUV4X+
PVV64*'E3J^A#L;7<<19VP&K*Y)\09%CUGP]ZFX[;M02NGT?H$:T<<BE05?Z%O/KY
P)$7K$F7SF&%?!B*;_%]*YXPAI>FEC2B>+"%@OYRDP[YM;B\R/7)"Y+K(3G47ZP%_
PFG*:^+'AZ*0I&N@TS^J0IKJ,4C)4#<)?H,3O3CF."AC3U7%:E>5X*^<K;8F: $YQ
P'&4(!Y3#YF3W] 9D&0EJ_?&(YEO]+_ [2TCK*!_L&=*/K'3@CYNO%PK"D&G]A#S9
PZ)H>LG\V"UM1&DH[?^*K4H%<\%\:"#$/P>(W]0 @>V#)M3T!_"GU,RQ(UJAUL,O<
PI'^V[\9[+ QYF_B2WU@:< \1+\(1]W>KH#Y$78FFC6/QX-H<-#.^$-,4WHLE]"<O
PB9\N/>S+<DD6D=-]]R '.,BM!_&)HTM5<,W=*+[A\.XALSA0RAC54;@G*V,)Z*8+
P7YV44G1>HEB*"F!1_RH*!E[W+"B6]G7:LC#%4J3C=:!/#>;R"J/@I&TLP<=WAGB 
PYZ;?PZ]L*3@3C\'WWI9BI3N9*1)@$C/[7-,4W0?]1\>,.PRD3N,(EUWNDZ221Q<K
P>0@35U^*J/J/+E5_6M-)FS^L,;9K>X113,FQAYGNUZ=C;G9R5\<47NN,RTY1D)+U
PJ>9L&+;L9=17[ R7GZ\HKC;\KA=4QGH@9!E#Q 8I'.#K\%;4)!"AX)/L\!<O)BK3
PV;&FI1%YG?,*8QVM^F6V,E?3+_X93XRT!91;4Y&J#XUE80FL=%DB+:#191H F$!*
PB><@WU\^/Q?&O_V#?+'P47#,),Z='CG?XAX_&F= )\7ZO>;&%_1L'1NQ>&JE=;[L
P/L>K]X%R\OCCQ3[ V8>PO4"%@*M]S .G?7-O)]YKIJE<SN7\2FP!<.3Q@0NB7T?V
P=]BSG51D9X]QYG_+A4:<>0"5,:-F.46'\A:15G9W)/_KQ=;11'(#4$Q+E*'S_KRM
PR'2'KID[CK!Y+N&]CS>Y(5 ,(P"2(2 %P%'9^C" E*EFV'$(N/AL>#AA^@8U6&IZ
PAY4O: .*XMK+WE9<E+)B8.\Q>::A]0&D]M]R_Y5[=VM$L;.^J:80'KH5\73X":Z#
PP0K9V4D#2]2WX(/^#^. .7!2 >F?EZBG@/]!]!#.WDO7'VSV"R@$,=(O2^$;%D$#
PT(V#4XY7:WV(1_Q1$ID[';LUG$8?$\]_89S$W"-IUAK[%&KU\4H#N ,0/4-@FN= 
PA#ZO9FW'0YZ<11,E6'0-M<P6QU"?]=3^KK5U(](K+R_7C&-AFAD4'T1,EC7P1-VR
P0"G(Z,D":^Q]5CZ2YQ0:JXVAGJ>6OV[!S_:_&$F]!FJ=47]D)#CAU=*8<-67JOT1
P^4\2BE([5[DP@[\(XB>E$AL #14".++W.\Y?1G^)M%<_B7^P9YZ=YCW(P>)Y&#,%
P>C9C(*J>;;Y:TL2=4XF.V&;/M"Q\PQE1D<.#CO;8[9,0H%75H>E?$N7G.P-?UAA#
PKKTFQ^Z8;=DNK?/F6V&Q2%';3,#P\G2#LP)>N-B:[!7O.KRMF27S@</PV[_*O]EC
PS#N.059K$4FI="[GD;->84,8C4RAGVXBU'-H?D!48VS_P^1-_T[U[O9>)&0>XJ:J
P2TY_?=*78L$24Q&%YI*2L=/C!.A8YU9&[4>NO6?R/@80X#4 >&_8?IRU(^<2N:68
P:E,Z'KR>A$M>RP&Q'*)W9,_K@HO,:/!;E$XD#N7IMEIS/7.-?YP[)_M_@=%N?-PE
PU#S^3H9S@5'5L<GM\;5Q) C;F![=FG=C?^)*Z"&XA259K)>QT@8FJ+5\$\@XA0/[
PHNI\< 3.>4Q%7F4AEG>7BD-%3VWX5<NNTV15/Q3)S'XF_R[F[O8>>$6OZKUK6H<>
PW"?Z26--0PR1%_7P<LNQVO>Y8]Z4D=)'TKJJ"_*R*7N"E=8W:="]TV)\G%HQ1U<T
PQ3B@V, D&M'QLP.X3:%" &^_)' CS;+=P'%'I6UHLY7XL'2FS22+KJ^&./Q- T<O
P"V:0X'N"=!'?);C25J":L;-MRX*B-C]+6A59*3+L)#5[(@P]QFF(G<3JEK.]RK B
PSH06N$;@RF+O<<B/W@UNS9?[ .MVA;X-$1(FV))L6A==BX&EPTAT[1E.!/8\Z*1?
P6<=+>J644?&:SL='[%%FY5/CYA?1HI?)V7-Q0LK"3IKG!]8P3@8^QYFSQW[/>!S6
PDT5GQK&&Q(AIL[*L-!M.[TW1"^W9NT%S90\9"[7,C:Q*XP&3M-:]O;X T(DOG5.0
P(,PU,G0:AS?[[:^;L-0_P2QS"]R#].7G1#&6#?ID%10#?2Z,Y9(-.\\.PV;#"_ 1
P&,#WZUUG,-</7IJ)$ HKU1LT[#7HF33WG=$97)ZNY??'@ID <77,_GV=J=]ZYP(K
PH*:,?:B?B;#:5O2];>43=+!5KM8AW#"4N#6DB.X&LN%[=2 $M\ $\<;7P N;^A1$
P#'_"'[U3.W5?TISNN,V>SZ3I%P"7N7"\C.S^EK?I4_N^+M% !83"K]B3CFJE<R!9
P+'8GAMG8DOC5:IUB188<-G:YY2TS5G=1$7< 2RV>+ER"LLG<1OYHIHZ53UAE P$Z
PK[ @!D!&TYP^[S'.'UA!+[-QH!LI$'CIZ!KN$-3JN802[<T]9"0)/XM'<E1(YJ]/
P+-:,YCF"\UY#\/W S[&]+A, $-MYTJ]"Z<&R*C&2HJ1;43T81X";U<$ (;SZ^W07
P]?M*K:$NEW"-(_3^0J4"BL3J"T@'(.L.>HOIC9;FJ7S(W.L&2@@Q2+8$[DG!]CH,
P*>')TN9R;4*! F8'/B]7H>NYWM6,X+FBQREJY5KY;TJL>]Z5Q2S@NNQ:0CQ%NF5G
P1S@J+:T0E\WF;0(-[VK\K^ I4)&G PN*:-YO&>O)B9IO8C.F_>@LC+Q+=%TH]CIS
P$B,WZZDB/KR:03;TI6-F_V?N)"(A/F#3=C0.X53>UW+8ZNY5SYNW+V5Z49$=C 6V
P3DG!<QR$*E4?VF?CNT  5QG/UTX:UPUZ\' (@2;5'K]@-\L"AA"USQ7R:@7B13JU
P@#?ASKWQC\1L8FF/KVFTG&EC?SEJ)G0%/<)Y:O8.^P9H2HIZ>N2@/-*):)3B1VN!
P8XX!7G9AA/K0^M<__0YRJ4P8Y884[[* ./N#,36QQ,*%A0:V.$B;++V]#ZV<QM0)
PPZ )WY0PK[1PYZ4H]9_,;&7 DST>#3\@SAV8YA)'9/C0CB$=WU%,7Q@YK!BWF#M5
PR 4/L;1VBB70V2X-F7>3I2@J1IMD#",J^=7,1D^(K5## Z!#" 7:S^+O<G.0N,A*
P4C4,=3\VT&W"6=*:? R3TX/84.71S8@^4*Z;.&D KZ=)L11B8K,5%;"<N*F6:[J<
PUQI ,1-$TY=;SA '#Q2Y(?S9R_N=L<B2N.@'";7#HT0]5WRQR>"KS?^AB/R.B\FL
P>RAO.:^_,^>#&UHW ;8<_F\TS(.]:PL,;)FV#J:&N3][.2J+2Y22GZ"G7^H:%.[U
P ;OKG+5%Z+IC)DM,7P%9^.[2:YBS'4ZCZXZ8F\XOR1.(&%+>WM83G2)AJ<3A+CNO
P?%]^S+\>UH=N?6X2I<[,R(EX#M!R84BI')^K3F).=J[)K*EU -IVV6_&V"]X*9ID
PPSP]4'<_W4&&@[)XR2=-&*6^@9ET6UGO,&Z[A@J)KXL3LQ&SC_BN2NI9]R:+46=*
P<*TW.2VQ4;_,_N+J//<H*33,O7;M?(LLM:[]TUQA=E\Z>COB <QP,@IJQ&5_;[?6
PM]*=@@<QKO6W$!8>!<NN=IM"GWA&W9T6E&W?Z:MR&+2-:Q.UN_U#(4RISD.<__M'
P[K2AW(C7W"$3QJ/L?JO!D+@3C39#YN(#F9;$Z2EP[^*,S'#]L/L;C^%4(THFQW2T
PDL'!(3KX2S_KF%R1YM1BIA98&FD9RE@V-_T;);%8 9P[MW,Y4_#MC1W;V:A738$M
P_1WQO@!UKP/0I1KH^7#C*]FC#9X&:;J_,X=E\8+-41T[$+(][@B[P0U4*#8:L=_\
PN/90;_X7R'B0O(X6S<1(9?&>,/QLD);;+!PFVB,@=J]H*F;Q3#OG1\#YT1+K,Q+:
PW$,!/U_HT<$T&,C2$!'%U3K"3XVGS_>YR/:IO EP_Y6X]<?#.AF'EX/-G)@P"$!X
P+<<2 [#230QGO=>9AK0NX>PW(Y2S3= (\)!OQW9]3R,MA4<;?+CO*A$;=7*7@E:@
P9X9/)@SC=F.I!:ZCD69I,BZ3D;-L>#Z\L#Q_+6F(]? S=2T14 5!L/H0KD0U,.[0
PT"_]8-0>*Z)IKJ?@WV>Z*'-\H2'+'QM10S!#XCRI'WL0%54&)0L>3S"^!K%FH<?"
P%2B.QK),D=2@R%R<" ENG-212C4$/L\'LV0EP[O)!'--39AP6FLB79VXY _%L(06
PN/5K9X5SH5<#_W)6Y .R_QN!X9,#V<HF^:S",]CJ%YL0,Q$QQXCMSG)4E'(W@&LU
P8^FBS4M!-P9O[JIO8L\+=]?/1T%4-,MZL$Q/J+RU)LSIQ'SIL.*/J5!$HP2H4= A
PI1M[N;U6:]70V:3H6_C6)V;B!Z57G(0OHQS&5^E+=($"JG7\.:+^/QH5%)?M< 9 
PI_C%6=RLSHK8VG27N7*7I (.!"36Y&>G2K-9-):^-MXGO4*7H>,0*@G52Y01E@^R
P_VV4YTT]T^-DT*/>^#CO&"&[!BFRGX$]YXFN2 6B/8R<M!8!')I;)M/]/%%?9>$,
PFE9+]>W\;#I^1?K3\E5&7L$)+$V_WX5D ^27X!2R YH9MH*FB<+_A^R/178],;31
PV%==JC:C':8V;YJ?*:H=(:9@(J<.I@MZ3L%7()ZXW3J X7^<4*1HK;[ C-?IW14^
PPK\IL,P/JT'&=@^)NJY7OBTIW508U+Q*43IMA=DBV.].Q>\OR&QTUI/PFNV':->F
PW)[V,)ZX#)UNZ?U47%A<>X64<OCLV?H2NEA @HF9!7;4T >;&+>NV/J(.6/O5.II
PQ$70QC#@ "8;C-.L5+R%1,2>\H[ 5.SV%(*(TBD0%+3P:O4N-2>=_>:H%HDNG?4>
P77Y!6D&[ 79L$/@GR)2=]9LPOBE+4$;<Q^6B1K:C!OS0#0E3+HG$RSZ_IB4@, =5
P8O$$:,1RAU228BNE&V, CUNH[(HY]!6&[QI$7%ZW0=87%HW9>ULBO4"5]A>>1+C+
PCCJ"Z[]$7PI([_)\EY.YC&R $^TL%%40PS9/A(Z7F[.XMJ?*&F/-PHW+J5P/??%0
PL,;9V,]"3!["?1I+4?N'T0X@%G)HD!R.RHR=BYFH$<+ *)^&[_SXCO%^MPEZ;.+'
P+"7*>DA[OB8%:%6BD%QO1*(-VJ']O[ZI@=X*,#BQUE'T/.>TTX!Z !I,=M_XA:81
PJXVY!*1%-R.H_0G0T*XX86%FJ:Z"]1$S9G(F] UZHY%<G-5?1HX;"N!$AJ@8C.;3
P2\DJ!:/'O;QK5PE:&CS.@@3U91LRH1P$_C+[8.&P^!>NP!=2U8(G7TX(.M&5WC8N
P%)3]O*HCZNHR.-)Z(O'2D-.1[A?9'0HN7Y";C./HJTS(]^YXBZ2*X%IGVD<)F@\T
P"%?5(O='=T6OV6Q9-KY-*J9%8^-Y%R;C\]>QNU\MK^K^JL3\(2HGA%49N:+"MB^"
P;<$2,B8%+Y?<;O5OJMS+K+AF=#*) G!OX[]ASDLKI=W-/[.;M:E9KI,$NA60+5T^
PLNH0Y]HGL9-#/+XS0S"O2\7<LA;U^D:YAZEG"A^4"9CV )HC^BERQ5K,2E!Y!7/O
PO'NHO@VH5"WXR L%6%.B"5->)R(DA0)-IA14\>JW&O<+4SGZZK2Y^;")&N3IU(4/
PB?F'\"?WE\>H3PV61$-S;7.]-/OJ(/B$Z"VH%=VO&#< /+*VPGP-[KY,&!GNW32&
P8^L3E\)26@[>W&PDR,TTD?<2*[)$*149MM2@PM+U==?K:JZ%0)<\WYB!;3;A+)(+
P*8<N&=7P@8>?C-]VT_).ZRT+IOU%^F. 7^B"!+U!-R4*D$I:6>QQ4]&E8@KD$B=I
P-.KPV?$ <.OW4F39:L(ZG"P1*:)%X]Y=55KQ44)G8TV%[&I>W?W$!'8+UUUGK.QC
PN]>:J3P(@(LB.HX96G2)UD#+BBY%Z)N'K]?'&54RI-V"KQP_H]_F?L941>BCS=:7
PXTNILQ!QML\0,(F@A0 Y=8PEQ)J%@=\23*3DNTD:!?MTP]\3G39;.$>^WNYZRHH8
PI6%/(<BRT,:[3T"%L!9]$R"/G^CO5T22"BKUK"6?ZBYP '*I>K+";VT3'.ZV//O#
PM-CJ:EO_ZF5Y+\^Q,:$%XC %)JF4I<2>_83%>)O%,L"=R-.YN)]+5V>:WPQ 3M93
PP .J/_,Z@^A@9Y^6?0$R\+44?V#HVBE?SK54KSYO(_$/\0/Q*$OZ%A1-^Y=P-8RF
P >=;SB.4PD.OV"<I._X,MOD?FMX?I_;DT[&(Y+B,\1+%J)YG.N59O/(<5,2S6<3X
PAE^72BQ#7UM3N''>$'U<>@8P>)8P'"7]L:_JM(.CSE_=2A>B?PP,R0([7YLL=9U0
P8[V,QK4:7__)V6I3,]F-[P18']@MIZ[:@5B3_8M&M$V*"'8.P$8:SZ?ZU'?ZF@W5
P_]]!_8=UZ(_MS;NHWD)\Y/.!>N;*D.D&D6=WPGX"XG?GF8+6DIUE U#=@MPZQE!%
P=LK\EK2OV[G6)9HX4_'[0;FYNA_3N*C<NCV@W3X%8="@?M*%+=>3H&_L%'F\>,B]
P+XDAQ?2+U<3"!T?+[8D[3>7P-;#<!)])>26X[U3;9YE8DH/G<=WA>/K+]TL;-L3&
P;LD??#68%4<F+DJ'TE#@0>US&3D&:4-=7)_C1EG45KED1>VE*H0*F,,<JLXLUUN3
P>I7 0D5WT% (ZASSD,$54NY0]O#7[5!NB"'F.P?(XV,M;W#8W(#:P<?%G+YQJW#?
PN.60'U6:I)"BE%)& %I8^^LYY,A:J_[,^[)\5'*H+.Q"Z'[<JG0MI#*-,/]LV=IE
PHC8.-6\R0TBU^;GKLQ-YM'%QE+M*MT3 =YCE/ M:2DHR217T4I#LB04'AY\YB,Z\
PM8-4]5::1MDP9JN4)@?]E:T_47S(HZ(LDYX@5+FWJ&^'LCJPJW.](V@S>=O*BAK&
P-XGZ)'4'\VES/,#V.77^+89D!C*RD/<%"+].J'WGE&+=Y23:C(#U_4U<S83KQV8R
P@]^YY)>QC#4=04_G;TD\"=2+M;I!0?46<];\#L?SH:-GKV)9L><#ZLLVQO@[4'WW
PBQYGJ\&'X[$\_<2U!W^,;6&I>#U4_;)I&R#B(S6/PD7GIJ_8Q9=\4>H+W"#@:_# 
PY6+P2?3A3EHHAMGI_V%<H8*X:A2QCSF':$EADN7557[BF6+C$7QUTB8]:E<&ZZ:K
P!'1?!F+Z4)K]2M&*H-H?YUY"]EL=[R%8+$4XJ".Q\"E!Z,QDKHC+2?9M9Z6SJ#7D
P#Z7T^M63P1V-^!;26B#ZI=5E;)'+=?D@EPM?FN@OGVA+.#[8NQD88#I^B*4KA0NO
PZIKZ]Q=DRG;QM+V*(:$)GN0_'RLEW@P_/?BB@$(RO719>I4Q+$BT&[+;X ':>,2.
PX]J(8*<ED(\P5(Y@=H9XZ9D_=36U^Y-DFS"0 #2\'=&5KKZUWA8@;]!.,"S%=H<7
PQ6-KOWFM<R\<,=ZUEF=F4HSO:U0X3X+DQADNQ]?]1)XS-/97B<H38SF/'YT=3[WB
P[)=@)%L;<AQ;"9FT7IK"4+^V2,E3<5(C\]C.:1@*([7B-1R;/SI/2)]LVM[T;LXJ
P K1U#.\VD*2$.B"A'91>08D%J[&.+WT$EK33=>$E4&[;RK])_0L5)[+8[,\Q !T=
P]EY0SY5#9BFNJS]I]GIU]N6Y[-%$5 ZMZ'O%/]*=P>6 C3/M9!.B@\VH+B0K#FJB
P+?Z?"SVS>S?+=5_" AST[_3@P3(_R6UHC_"FC03RE;34*<YH"#4P^V%%[<U G(VU
P8N<_EHN\/USRR\A4M ,H".\*X*#F%?>I[!1%#KCI55=0U=P'F?GG[T,);:34"(5Q
P)$>D#^AB*B4!\B,];'3!;^A[O2ZGJ"*(Z"#10$5FZ'X9Z]#D'PJ/EGP\H5^LMRUH
PB!!%W!NX0DY@X-9D4!9D5]$L_"H'$S"EN!<5%QVZ8ZX3L)T]UCD0X0,"<9)GC%6C
P*X)7>L#2K;Z%H."#<I'.=071INELJ[YRGUTDYB?">@0AYF,!]G)T.:1O0662XL(-
P['7^ :E=++GV%]7.:<:B(:3T%+R$^+H%K@<"R9'2>Y1V O0_?RDG<_H>[&8##?!6
P.YS_$)H.8>Q8!\6H U%TL$#_B+&Y,YEB8LQV^XVN;J:2<K=&SXX>QQ]HU1&50;+E
P"]P/'T;;963U&I-K%:O"KEP^)AM*?&_F51!L$!B:9BY0CO+S.K5S_(5-3Z'1[A\I
PA) >BEM-0^K[@VOQ/CU0W7X6 "$VJ.[W!]W1AH4* CLQE?5[%G[\<16CLYR"XF*Y
PTJZ# V[PRZ^4SSUFG-=:K#QQ6KUDH=\\?4SJG/(!RU$9^/'VQLO.M=4SC&0\.7LL
P[F>1@)9*WFN/8^U_^@*4G"=C0(1+D&PJ^J3]8-$O4LMJ2*3_[M*+2:$R=%NX=[E6
PSA&WKHTX\8BH[WHMM8?ZY@(,4GG]M ':FI41C:09\M!^ A1$3#9!9>([,:\13M3W
P+H6?-E;65,!0%F<]EEVRPDL\6?SPP(N:FB.^MZ41^#?=Q]8ETC22DEW$.U-K%I^&
PD'<S>+PM'+?X)]F8-N;VF<401NK#+53U&+MH!\@(=0$E?>+D*)0@QQ!4! +;UA@V
P<Z_3<4DI0W%VU(]0"A0-^QQW#-GYNF,VKU3YNN]^PY+Z6-4/_LP!9@JR8% S(<2:
PM91U[&N1^A\H[-[-SZL@?_J I^C-SU[P2U7<XW6E<V[T"5[L?[^P/DX:R)C9J?.U
P=UT8PD_/I3!\E7U/*,JK_^"M+"Y5"2% $^0*9<][?UWN_?Y[6_B%_GN'9RZ:>BKZ
P4H$CSY-%^]>I<3ZS_K L4$#M6YAGZ_OMKXQ_S[< R-8)A>7K>_,2I0;)4[)CR:MI
PBQ\Z?(]5N@MVQ)Q^U+U62)QIW&3QQQM%YS;Q0[%/AZAD)"/TV6W]\Y88(0[.<SBV
P.L(<M,W7!,.QZAD6?0G^CP\"T-V57^NN#W?+HDO#2Q':;OX2:2MV>2X_^8E'VX1Y
P'Y;3# .;'5@:D![I?LR0I#EZH/9-!54T<YN82SC2U:^_#A[C%3AUMU3CIH8L"X1J
P$[B*,S@< $4*N;BC$JOZ\A">QL??V/5"7,SGVYB,^AK\[!+I#'9GW^IZ]9#E='T"
P3 /I4JIRPUAAF-L0U>C5\W^1OF*D*PJ:>#-PPS ZZ=G8)\QT43Z!%QF8Z!BUEL ]
P7<'(6.=?&'5<[WAV],$?Z(J*69HTIT%U6EX5L<5;AELMHO109TE6-&H"#%6+.)KW
P<9\%T<W<6) \\GE5J_3;0V(R+"XBRYG,, >-^-DB#1HR9]^C6/'-M:O +_)(,V-Z
PDL\8*SO?2GF?6L71+Q<9D/PKYF#*>4Y2J4+QF=#)1.?\TN2R6.7)8CE-SN+7*.94
P(:6X0H2H4Y*IO=FKL_5P<0C_:%% #(3Q 37B [D$VI.:9U40<6+I05-M+#LU"!)O
P<H@F+7,T!V(7"J*'56UY@1:$HU!]#HZHJJ# 5N9S(0&\AVK=9:_,SR_ ' S1OA-<
P6-9:13>PW-JTC\*QPQHF7RZHQBAMO"]"OT7))IQ6[,5'N6PBX1<RE.T]S(4<P0_9
PHF1S?A,) FQ!',G<H[??.08)V8O50LQW$7TA8:FWG&NN#@M;)Z)D<(7Z@5T>("9K
P,CZ^VN#3, UW%'\7 IVG@&PSS#*N,3V>WYH/1%%.\!B!X!C4Q*)*:+O+.2;AQA\?
PO+__P9]0MEW\RGRZ.>E!L[VGGEV)Z=P50(*"$!(2)M0E UF+9L3C$'^0F[&AK0-\
P>T8UGT]:KOR5(SD;A?V,,1+KFI@+9VL/AV/(JJD9WM"C.YZ- ^>((0&E$INT-+!S
PPY6M#:B/!IX,F_W/8TY["'Y+ZW^T:ME!?T-&^NTYQ1;HD+S?*7\Y L]W&,/JM;G?
PN)@;G?\LC\R"Z&>,ZG[U[K33A[^KX/O4)/J-^IMR>S:([EIKF=-EZBB[)#B!JX9'
PY@4G@Z6E.Z;"P^XCM$.PX^+0:G(PC]T40MMU#/GL77$9FZ2):K2DO9HFY[2+8@(A
P+$)O#RP^MM?V2PG>D,U137/W?$N;$<DJ+P5=F_"XMN'N5#59!7(0H\:M+9*3@S;E
P)'^S]A^D$F@S9;+/KF'#.: SYG!.5=J_\U4PSP.Y$.<\<&K^CN[$%GRO\\T[5(XY
P?/\-&.S$/U:L) SQF&G?7_4"1$-O.Q6IGYWJVPE4S;;@TR%-RA,0^A_'3#[/#5'*
POQ*%+9PPYOT:]+FI(A#?T* #),LO-_6UXHF2B>8]-UN"9/46G?QH"0[0//Y)!/?Z
P2 <#R1&M6^_Y_TD6S3_ I0,\>.(Q;OI7B+R&,Z8;/DKQ(F'%>YW]>SA?(@DH*::(
P<S.<C$AA\T*C61E;1=M'HVAJ+)\RC!2435!>3B*D>U892M7G4"HF!S9PMSNA>)(D
PD24I@FVZR39<6YPNI8I]]I<7@N0!D'6>]B7_.> GD,66:*&]NZ@MO@=EHE9HK*)4
PJY^#80E/41QVYE0</\4[M2>Y'&Q&&W=FN$Q5".GXQ+'0R]RV(TD-4$-CVZR,.IP)
PE$G8[V+67.HU+90!/M4P14NI^3([?DR% HEX119.# 994A="1?[D!V!2#,\[*>XG
P3Z<8Q7#V#/MM>WD^4#W<+JFDH;PVK1F)J71ZHD7T[)1-SLCD":GJ<U?(;&E+^<\_
P;<K^RY>^7#*E2CUC$0@ECX>R?=2DSP>CE\&L2 +?,^]\4QVK%Y/TBF+SL5^'8?VD
P!07H25DL;^<$'S)7>7*02S!$E/W+JQ0^!KW/W6?%%_AX:\0U60?D&O+OHS#R[. \
PG$O&?.A-W"G:>-M8:"=6Z<QZS*ORY8N>I8>2=BR 1#,J'+C:EY)2@KJ;8#HD?>1(
PRZTL.N3KF)H/8<H,>HC&T912,_+YJ-3/_K<F,&>;W5].8G3M35Z>6CLGXBL<([5"
P]%JAX?_&8E9X[#FF.W"T1A;!V+)@-3_[\EP5O0@S0^F@,F7-TT"7[V6E)M:SO:R!
P;K'$A]'DS6X>@OMJ: W+#T!/T0HF<TFAN*#X(K7R>;I)\+65Q>^R0LK[6D9JI;5X
P1F/C,Q*/58'*^*XW_N &\0W/.X8L=F,4U-^TIKO7XY+(:=MV"5G#E;5=8>4=$%-G
P*6(T4U4 ,W?Y91S((DDS=8-J=/>@@//5"C0,,(*0$U82Z@S3M7DSS[:"MEXHS=B@
P@#:?LW_YHGVJ[#7DZ?+8!N@&?GZG#?V%G$0G4/73Z7U.PTQC4S^N4 3$MQ'BWAJA
P'"L^_%"1X.*7>4R$7G\1ER@ 9XQ).9".E^1&LCR#1B 3R&9NX5!HU^5,QVNM%5N(
PR-F1LGJBFR3#]O$"O;E4G=L$SKLG24!N]8%E_.D6/[I-H_79-#5&)F ?R<(_6YRI
P#D>'CB=L=C1P!I:Z?O=/WLU0DY/7WW7\&$+&VUWEH4&64/LG/HA?WU!OV$,!,[""
P9+V&1G3F#7<[I2;$'^UX8M#V8J8VN!^374=7H)J.MO9T(I[4$-, 5AR&&,&N,##*
P@A3)]U*05&=>X/QQZ&[$Z?*C1]Q,61CR9A-@S_%$A- D;S%-=[(5!CA:K4:%%8,D
PPE;Y=BOZ)H*M0Q^H][F*@UH,K+A((7WK3N 6A>9?Q5 X+%+O%';;#83JO$&\,JL+
PK@72E6>6WDOLATT"=U#:-G2[.86E\*-]B?I0-ON8;)![S;N%/J(NYQ,OT-P09;^Q
PBUF#O+F>B@5*X:E :4SG5O--:ADH!!AT\=)I=5COR!O@H,Y,^4J8[<4.GCL$:A<+
PVU1ZI,JTH385.I%2?Y'8CN+T7!JUL<=6COEB\;N2+R"=64R1G!#BSEV*VL?W,:K?
P>TU4!Y4,HO&@UH4<BM.BB["3&6GHOTUVX?\M/1B+\X@]YL:3[1X9ETR7.PX7QL@=
PPU O@/7XK8A,3NR0'("QZ$^"="==C:G:@Y>^VPJ$ -J^T7HE 3-Y%'GNH7Y@QO5N
P7\44\ G,=<+ZHFWVB$ALQ6P 1'2Q)5^RC9XOVIM$M +YI.S/5I'+&U[)R'_</RJS
P.2:R-1N/?D6AR\&AK(I3_YHK?$!R"2.^;A:18YT?0[.H[+YT)FA,6VG=>)GO:I*8
PPJ%>F"70KGEUUMJ>^ZYL_=?E46ISP_RLG;^JQ@]":6UIBGJ[U;/,+)X1?T92LO0O
P:R<>3@XH=Z-2@SF"QG<,@QE:WH!L*W>!X_M?4D1N\T&&)5KD:J<6JM.$U8LG6UOG
P?MX#$<1SXAKI9BCL:3_LIJ9?L_N:I&Z@Z?T,K=<;736V:(=D;8USO/]8)57O4=_V
P1JJ7 #Z<?SP1:XN>L_Q7THG^,2-?J*;T+RIM&++W/P3G22F[VHHFZX[R6SRL/&NW
P5=%QYN87*NC.T/%G.JA5IVL]."I8KG"A.G#4HX;5JS]-7RQ>B*ZDVR3,U!/<?BI=
P3*D"20B0PD,'Z#,/6T7TOAAY L;9#2!"2[$7T!+)EH%?Y^D?FF"8[P?V&AI(FMY;
PX7<&TVN\7#M#MVI<$Y0@#MT1-6O23'.\K@F.-[).HNX3ZJCT_RD=2A_7L]_[Y-C%
PK79)3_FJI8W>"Q1B0M>R32<JT2\$"[E[I6#&O4P#R'0E\_AC]QL0:"(,Z+B>@BVS
P76(/G(Y8^SAQ8A>%- [X,!VMP4+HR_]W "TYHA7%TU2[Z[5[=.K2X[PEI$XGR4^3
PU-OL5L^1AL$X#9F;94&S XK0R;^<0,TQ;HS?@@,3BY"_TQ=B !N1?LXV<T ;1IJW
P5N*9\ND8CU8330!F9(EWG#M)]A.R81TRV T=7]\%1 JT8$PC$5@4A^*MW8+@.RB?
PXH\Q] S."".@?5W;;VDB&XD[X2U=;0JZG;CE*Q"WY>D25B!NA2,0LB,1RZI=L&J,
P_9)&GU,;#<U4B %/6VX)-@_$<3(Y2[1>D]Q6BP-7F$*XG5%V49B2:XBI,E)8109$
P?B <QPPNPUI-^7')GGX@ESJ>GZD)?:.$6K=O)VUQBT@5L\6E\<W@VA<VM8X?R?#=
P25I2JKLD%LS"=%JW!N^$EGT1!U1_@EEJQR*=S<K9C 1) L"+K A^C2GM[)214NS9
P ZSV."NQG20YO-%H)D7@]"#'.UG4<[@&4CL#.;PEV%U$-[Z(9^KBV'[=%BO0A"X^
PH:Z/V/_-TJLCONGEZX[4>5/465R6QME#C#OF\S?B:DAN\74UY5":SICQ_Y6XV56'
P$B?'A7+J:\R3#D/EW9>#SIXX=1<X>>M1(=N]+U(H-@3]D&.Y]ZK'<<1C+07< !R\
P'=A)(/,7B\C'A3)TF)_,?]S7&XDP[3%I=_T'*@X^-BH_7Q>:<'&ZK:"34/R.8ZK4
PVQ8CSZ1;Y[I4(11'ZW&N/(A&_]1&/-*O0;5I_/F(+T(Q$?/2F6.DQY#*&39V39?%
PI!I4]5^\0.Y9MV4'E7T!ADN(.,N>Z&.]V:Y@:<W*/PG\I^VL12)WB9KSR]RM9"<*
P2%Y')]=X%,\'A:-E]Q'[S2=O6P/LN:L6.4@RP(&*$0^K%A>6*&QOU93IPW"$T5</
P)0(9KT9QYF$_&>4<[;G69CW7Q#20):B>C?)MC%W6"(_.DK=->I,Q*N^7AA570DA%
P"HP%Q>2QPWI)(]NO#U]E! E="R\J3Q7#!?Q*C>")6&]83/5.,5G[Q1T18(<= ^ES
P^F!8E><IRT"(L;%THX/V2V[V!K8#7D]- D+%!#0%]?QT.W3G4/H1L0RN',N!.O#3
PPQHKL34!(>KVV0H0/4XE=B')0(@LQYUEV""3"R.B$<27)=!2P6#E+@8^2\?J#5P9
P[QP*I+7?+*)8V.OGDO;NA/3_^@+H_F3R9W3=LL01G+\;"BJ@M"E157CQDU!X88+,
P(T& =AE$]S FD=<OT]62_I48OF2W(<P%=^)TZ2E5/TFAWHN;DJ,X1D+YG>R][ G4
P3Y1<(<Q6XBVT86!=(2,3:(YSH\P_;LV.OOQYBR""; BT+/3?H'5V3J@(4S??UG@K
PZLB]NG=$8 #'FY".U!8XO#R4J#9?\8)B:0I1P=6)/]9GH(+-::F_=EM =M-(A(N1
PI**M<^596A]Y_PG1VZ(#I4;"!+@^AL*"HZS"2LQ4:$WXBW176ZMEQB;[D8#+U5EB
P6Y22W(7A*C2B&4MM6AE4$:SKMJ*W">O*%D4KQD%,'O/#STW6D,4ZQ/<AJLXQU\##
P:%R0#C$U)U",GQ;%%W9+?2KR;$C]VY"Q,(-3J_=K>66#P5F&!KTTA7=/_=6%/A+K
PE%UG14E0HZ;<<68F]Y+62RRA]T* LS=:>7ZD#&'&I'U8%\R]3H'S9A8O9*H:"],Z
PSS0PDA/+' 7WD[3PP=4[G"I7_8>V7P/Y)-=IAM>P+FK\QB)94M.F3EX7@^Z05LA@
P." #0*\Y0JER^\B$,I&&(7)!\;59+VM%X1O"_%JE!L3YWJQ><\'BU*C^$X76@[@S
P]*;*21HI@U88M6NEQ08:-N"QOBX>I8)?+_<[,Y]0>SZC\#E..@C2C#!1A4>#VLZ(
P44K#LP.H2:YFZSW*$?M61[4N]GV"5+)GI:8[F9I$82N&XT7@"MZ'[5XJY$*8J_FK
P'?I"?(#'[.HW*43^?"4&(9OT,OMSFNR&U!8V(ZAP!B;LI[=*/ 4PFL@K<(,SX6,5
P1)DV^1+*%[M[+-2JCU<4O;W?-WX_Z(9O#PS_L(G;$:>R=LV;0 ]//=:/P]_8?U@&
PI_I"7M 3+(.(;OR9\8L1H )2+.N.SWI3SND]$(:Q^BVT-:+Z];6(WIV(K.+1Z9#*
P-P0$+L";5<T&FR^!*>S7VN78T=K%AXIB;1:D<@QD';.G**PPEHQ+?9'TJ VM<YF@
PO5_QQ4U'Q-03A3Y1 ."9:%*/QV,U/"=.$M!D\<(@<'<Y'( AT&C<.K926 YJ "H/
P3;.[?L#>B*YF?GDU.J2.CZC,(;='&FYF_U[E!)NL+Q'L(2B HI+6X]'U?/LWU$9O
P)6OOCU8^;04GYJ'91E#"AVJZG1ADEP@=".'&SF#AVY+/!$<?%<GQ_IZ)X ^,VYF^
P0DL=S4+ZK'W+8AH&&*<<"0)WKX$#\T2KF4'/7>N9'1<6=XL [ #7%"*K:#[^6T\6
P2!WYD*#!9@^BZ/%%1F, N,Y6,%#$W>;0\]K@_NV1*@ 4FTS-F'=*>6_QXM"O#B2$
P\D^F-Y'CDK7C?VB=%$:R0*DTRHZ=3MD9+/Z@5B\>'<"80ZJM3X*=8XH_;&O8P22D
P(MA\SAAG9KG'17W6:LT<;9B@T2[IM]?8.6)=8+[5@!RQ.@#;%5AO(;W6J6]@#CU$
P@NUULQK%H'.S)'.@/([&=-;241<4%R#.BX+4)T 2),EC\?EL:;U,&T;HYTG\C!Z8
P[:VB<EY]$VK.9I@DO:1<[8U'20NR"FPZ.ZNJ@_ZK[3X S/="NF]V<1KWIWX!V\RW
P(FRC=%NP$'JFKZDMGPD?HSC9ORXWNWDE HJ.7GG#C-7,N,2.5%=M;0I'6C]7?@5&
PV8 3,.K\)ILUT08TO%R,J>KSH?'8_>?@&T*TA-C)B$!I.-K1>2T*S7>.=+Z!^_1:
P3WC)$&Z/AL&"^3K[HL\31L'&^/;H*PB.!D2.[-.'460X'-7K.I4'@[QI3G;NO_&,
PZ?2!A"N6MF-N6=<>-0;C2CL!/U65;N4\$U_/LWKZ!4"N##1I7LK[5N)0MY'+GVC[
P, \Y5D3?@V8 24S&_7W$3-9!M??Q:(,\U]!)'=VVV@[H0Z70I##80:YT@78?KW$?
PY_--FI8=V^EI@__LT;W U-&Q#=2M!/'()P LTQ/W[V2,6;Z.EQ,*5A5C5"*=I"P/
P6!KMUCQQV)0.ZLO!U/L<B1>CRPZ%&Y="2)!&*@<B ^Y]\[(B]PQ!]!_#!PB"TN@^
P]F!]>B];0L)H*Y@PV6B,F[+-<Q !G_I&U!V;S %^O[5Z#>#=D6Q!;&DDZS5Y)7N1
P9]_LQ <?1VZU5-?A)5%W(ZY6Q)O$S?).>(\4Z$C<ZH3S'>T6;?,Q$YB8<QK#BD^5
PVP.Z>J.@1R2=<V ID!Q%JE?]R8JBU%NDG4P S"V2/#YWW#4PB6T<5*M*BX=JUA8D
PC+:?VE*BTO#IJIR<T3F,RZ'9_I*Z&\K[."<VA6+5IILBV N IRZ%Y&YK[2JN4](C
PKU O@=L\]1X7&5!#*X@DTFZZ?)KZ!&Q*Q<E%%<T/6J>5>\JS9"_L]M\>.:X<BU/8
P%F4F<;# A?]LI5_(YGXDV2I.>L9%(@7TWM$SC4J%Q([:R\MJVY[15W$_TV)^:A8=
PMJK#;P8$T,?$IUV2)3V2T#,P/!E1(A,0!F5_O]">,XMGJM 97W?D8E;\Z0EHRH#6
P'=/#_' ]HKF>1)J>2AQA"C0"(<(%C-FF4WUZ%1O6WX9*^*OV=;B4[^!W(,FCB=M*
PHB70%0H@-'=,_SD)A"S_G--FBWP\'0<^?#4E;;=AF,C^Q!IV;X31R85FUM(V5]^W
P#J BVZ'9K'42FP76618E1+Z+^N=3PL-4CW6=@)N?I$4V8J-6BT< #W+ + "4FL>0
PPVU, /\C]P%BQ,P0NE9^;?M+0\BF&S7?&;'[9_;@16QHB:.1\:H._1&3M%&9FAIX
P35L!NA'[D84DF<Q]K!76>\Y%V<R0Z;*?E7T-PT)@NAG @"JON:R\S0&N$'(^\FTC
P2'*\<24AX834%/7$ \B6E:ZQU7:[AKV5(K#.<G^G)]_*K!+54WYG:$AGA&:/17.B
P LMOM0$W6;*+R7,V+R;)^.?+DI]SE(0PFI.=_>#>3U. F7?XVM[1>-439&**<8RW
P^SNF"V2D\VB\8GN1.0F[9'<,$^V?3K\%Q+P.9KTE!HCBW.CWO>6'S+.//=N^PAE@
P><3UFH%-4_ZQU2U,-I=IH-6U[WO_-9U/+#UM9IDI+SSJBW60LY EBBGJ$318Y@J/
PW24E,ICYE: #@X_ D<Z[(ZN]#'(W1B<L<O,2R%CP_(:>!M7@ <,I9W[X&((FDGX1
P+O^ZK'?"V=[G3^Z^<1C5<;L?#)<GT[@C8$L.R/,U*M_P:R?#S[??N7,,,2JQ$]AL
P5%;"^3J%)\G;:Z'&X@"1_4 $-Y*UY5,"T4GQ;UI<#NH2E\>V'8E&0[A'>>7P/"DZ
P-7N3\;I*D)=RP1:-6TA"ZC=-/UH(D1)*5'3=Q^O/^/(M..4?P)F,9($!SSADU"VB
P3M3F(5*=&'5LZ1;_XPS_?1]9Z)W!6HH5+L8XJ8=IG6IG%ZB")VGG3D435I-!7XA>
P<R<MT1\;>PJ,J?OEZ/3!PS1<T?_HBB]MFL6-W-5:)K'J;<(:U"#JQ(N+,1WDC8$K
P87TT>C9+'&W PJ8RY$]27JTXCJA<RS9J0;%P8Z>(=SXZOH0;00S,T>]'0%H&.5['
P90L-LAAEVQ;2/9M"VY)#&SJ@1>#O$J& 0P.@7Y-X4Q(DU#1R 5:/:\G9'%="2\AI
P8-!2RZ)+F9%M7[?&U84GE'RIOVZ6^Y?1M!A##")$RUZ=B!.@BA=\Q$1]!M.Y^5%?
PI(+E,Y<&;?!FCNM#A_.W ,M6>ZY8N-\RX]4OG/9G9PA$!@ZC"WEV!@G0BA? O6.0
P)'%]?;;K<F!E(E4&$:"^F^2:3A+%W6Y M)A;$L1']:+[UYN*AV6$I1"8KDX=BA)2
PL#16?[*FF(_R932K!GM%IBT$!2(*'A1NRY\VZGLU1;IA^+LU;DO+]26KHQC6H^-D
PW3!&^+%2F)56Q=Q@C_ =3T;+'14"LM@^[?XX3[CK</*4Z!T1$JC+*G$:&E@J9?J!
P%LS:!5/C\*.$#0FY5G1V_%P1!26VW@'#"K"AW%D[W,TSZD91U?*B6.A6/N+-E!-S
P[K@ Q1GOB;KU1I%>_BD[KC_4VTH=B^5:M6A'0D\Z/G,&G=T-(@HN-].[W1D^4JY\
P/%>OBL%(P&_%+'.-6:ZV4!#;YL!1N7B)U']Z\:B,S6ZGEP]*<6X]HMZ#?)*CI_QR
P)ID5^_N.R^^JD\0A[JP? _R@3.@ZH)I$NWL#_J)MUV-&0KE,"O7^^V#]\Y=2FU-5
P_;+1O+ >=R/8N7@]9NB[BM QEKEB-Z9'P<'#;272L'-7+@O%^W.8]032124&#IDM
PF KVOT8K_0+I;YI+=6Z"(BA]*^:<9R,6N@AO#J@Q6PWQT1V!HZ?+,< U&=\[ #&!
P^2IE,; 12\\E!:F!8I+)H0R<HTN3S9)3+\PTIJSN1?]H#Y OKI1PK5:/$!.[,)QI
PK_/52*YOIC.#P;9-OC+,B3J>Y)HDDH)@[_8L;16WH\6R,D0XPRV01CT)[O/5(H=/
PY4H_(XU)Q<Y%5B+VN<]8S%C9RF'[%>W=KSN%RSLA*3KJ$%KNYJG5Z(",B%3K75'J
PA:;M"NFS<E?+^0E7WS@^TG7I'B^/NJZ-D#N1LI&_TY'K2PO@^MLK[9!%0L-F1W<:
P]](6 ,CA$HR)+O*[5U4IZ<D !1N6Z:%\8_T+3<3S&!*L7CT2RSWJH)-'+Y3(Z0)<
PF:[@8^'<YFMZA"^8+7:C[='.CZX!*QKF(NS[L;?DB&"M:M&OV3X&1N46]<WE19+U
P]],)N!2390AJLOK%I)[FOL:&!5Y"'*W+<]?G?<7DG.[=</=$<$$4*2F?^2-Q+HI-
P:0^A5GH-5G1);7!JP81EDE)L%MCN9F/KOB[RHY_4GRS-:WF'AWFRRLT":D[O=0G_
P!4"(.#DEB-+[[\E;_.V 9$WDE01?M@X#*1F0F<4 :)(EZ^F:%W?6Z[^.['?SB!^&
PX@"CM\_8^P_3-&8;UEM:*93.#VR#2NR_PA O/\8*K.5MF' 5A(MMEMJ*SW0."6(*
P?U+:V#?/K!;[(]5^-SCV*C]5L=])4UY^CI!%FPY>.F?\?>*78D?Q+CRO3L8HW$AW
POV]R0B,8+HF0@(/RF^,'RQ.*D=N)C2.(_2HY$1<J6+A[BH=A\Z<]NZUSIS-7S"(]
P[R7P[;9TEI'?3,Q<?CLC4 N]$ *4,D7[ATA\]A0B5*OR]V(J!_HU-N?,. #U (:T
P(-]1IF,>R*#3VFR(_LS+7NH@AA.+KO/J[00=( ]VM*O =O'[PV?&8CB<35S[F8 9
P'8$(^%D75L52UF 5*HSN<?4X0=,N^-(?4\L?^)(D0;6S><?8MN$(S"!DO@$4&6D[
P9Y"&P$6-=$RD4\,>:KITY0$L8+=DYS2@6C/E"6CX-G<[]""@P?)Z(7>5HD0:AFQN
P'(K,[Z;B9\_587TUYOC;=E_XD(&H:W\-53,=(B6;JK: +-CDW6P]*F@_!EQ3282A
P8V#C#O]G%DU)4;R2.%N8FRUHGO9UQXUY&=D-&CAN*'K8OAG[+F4E0<M9\"$B\,J>
P'\(ANK)UEX-7/&&?(5%[OW0.U!O#T@7U:\9-.?=1&>&FQP>PF><--_B98=^C#C[O
P^A6,EI0A#V"!VT8=<F'/4AL<753_QNFM]=@HE%I1'3O9:O?:*Q^RRN[9*(L_$XN;
PZJ$J[^\%H0)$AQZWKE&]1N=792N;[N2W+?956D2N)LU_74FI_U8Z)(J\HGP1G0H^
P"3#@#&",R/]$"#]I!SUQP5CNPS9-T=+S#[#1G*/BIFZ4=P=K?AT=KR#R%[-&]%)M
P]<3R>5V!EKGB3?R9>?_!@%-HDI3T-EZ#,FG&6BE.1*SHSBAN2_SEEXJM_P^H7T8\
P8*(MG3(3#60<K)-\8C($@+4A -?$('LOUG';U.)JD/5=Y//YK2^"O4Q\\A0PK[@$
P.C<6);.HKYX 866$DS#7/L7,$RS2 ,ABAE=YLM/PI0_=[1<,!P CSH"K976,@]3E
P#[&$TH\TK+88ECP7&T#](-.()\;6MLG!'5;EP@(G@4P=$H%!]_I,3QL.]E\0P+#@
P"AG:B[%E/OR&Q0!P8-&2STO)5?5QGV]LW0/!D^+09%Z'+KC^S0RL4C_[XX>#E %)
PE04[H>;#=9)L[SE959#=CSD1#&P7W8)]1#4) $<#[>!=F^&I?=E:N%X7Y,\9+Y.U
P8TZU5&AU5#NBUU#+3+U9'[Y?%R?:E:)$B51^^.5-D@]F'^WE'\C^%^"@PF7O TI6
P9W4=Z51['8KML>5)Q;>63+>+%OSH9)._3$>>DR18->=]J<!6IU0K,3-B=!W:S=;-
P3AB!<@:.#,[M;B9]&)BGMXTH-UTSF32!M!*#2@.T;&;^A^=2JRD?3'.G9 C(RO@>
P3@(6)_((.>WPQY#2?!KIBLX:\&:T+U9V??KQ+$,*.(6[BG/BH!(P2.S(69'@Z'D(
P8.99N?Q3+%V-Y&UOD3R@WH.L6 1@LP[MBK:MPS;YFV^7T[SB4_L<N2"%!KOB%& [
P;V-D'I\Z03*A,O+X441IF(V]=E4&32_18M]>&:/@/")3-Z"0HE%5@N,&LJE_3&WK
PP*W+DMY^/;^S=R0._KU433;W['<A)/Y,R+03VK0[$P/8QF%%S!G_=>N^3.AG:P6L
P*C2#EZ803\Y3SC4#6F*!2*MV?\Y]M>9,I<78FN!V38T"O,>0A%OA;:0%_9BNK2,C
PX>)7.8_MZV(&V@1-AXIRGX2Z_"KMIJX^:2T/%2QEO%_"[DC/.[Y'B-1._'V"#WF1
PF[ =1XN/H. 6CU$+.^;MJ81G.")<$14(CQI"FHUU%!*]M'BQN>:HM1D761YY>6ZI
P%T=I4XI =8V.'(H^V]'_DPT'<<15-\,ER'7:VJN3.0^7X5P-9&Q,H%=RKN>?'YOX
PYSRD+\=_C8^SD_W^^\@P\O*#:V8#/\-S#66RD\!;\/&2RI<K5>  H;9>LY*&CEB9
P-B5WG' P4B++N[-^B4/W$$HXC2$ 8->A3?<,D;_\G YXDC#*#JJV7< ]26W.M?MP
P-\("\',=YMT(=2Y$'_7;58_<XT:8EI?#R>[5LO>=2.]%K>"2U6,H8<>Y374V'1L$
PK4%P/AA.$RO^V>Q7<.JUOE,H21T40IC)5[:[+'7O6+]7:]J\O-TS 8#4_31Y1-1"
PR++SRG=4-!&K-=219UV9BBW3?6<+A^I[8:8Q>T_6P2LRC*,@%<IS$Y7;?=PO:0L.
P8D3 S8L'C[N+ HK:N5M;![]1K^-'$W6>,NQC6X_GC?&Z/D5G($I%R.*M\F!_)U([
P3X=^M6<Z\G5%,-[8=ZD%N01WY9HRVV>;("[3@OQGI"R\9V? <I!QYY;L/#8UW!E6
P"[Q>+$"<U8S+[(P_J:.<Z)(5)93=)_I[NH3I<^AZU9FE(:8C2!/_?!#O^#92HQS2
P+GM>=!+K2DV><<0IBSB."AA,@A6Z@<\<3?,'<*3=.@@I14<^GI4,DB<T/ *CGH02
P0>/@GG!K"(&R9;T@']%!T[6+WO_H<<D*,$MRVC(@3?3#,=P/+8=SX638PM,\!M2&
P (BF2*.EP?%K5;8KI82N3_$@4?A4^5B^F['4_JHO5XG4"K[$0[%BEG5'=XEAOUAL
PX_W&U$1E@%,HM^=V?RHDL$=(51,^&__>M>R^;0ES7:3=RUV-C;0S"RF$=U.\_C>8
P>GZE#DDZ#SOF93V\-_P^[P";[Z,9ME?,F.$9R5-\?3#/'P7Q=7)J,Z<+KV%87S$)
P0)PI=6"R!FT*B^>FMDN'MBZXJ![V7"2O$&6UNC,8.L6(E_(6UI*<".>ASO=1OISC
P68'<0B6HP1+J+!.S= IM/:T&%T!X5R,=RO+B4(C?:C"G !*%BUA[]CMB=#R=S]U?
PYL8SFJEB(+]=$,B\\#(,/W;YG]U\8I<AF"M:A;D$V+GBMDXN_4_:A1,%E>\VZ;ZY
P[/1]Z,E]1C#YCV'N_VI923^QZ%!+"^?:T=7\W0WS;VWI;%(XY4"0?^DM4PU)UIR%
PLF:G7[@+L:W5L@+!DD?4D=0)50S<@ W;,MA.#!N/,\]EAK=0]G(E>>P_P2S =<!B
P47JKW;M0/8]?<!MAVVD)_ZGU#;[/-E62I(!9GG5CJ1WM#)!AL1PZJCPTOL;@$@Z0
PY.2S9J$S0^"<QV7Y3_G&W6LKIF;V@)R>3<A#8/4@4'>5VS:D?5LV49(/COE[8JX#
PT_1A1-X]=>ITK<A?+R['JK_++G\1N72=18GH*%MAI-DY]H+0R>5'#(WDXQ%=%<IX
PD,/,').D5E+8H)*WS:O^VT!CS])SJ38TT;9>'+8B!EN1.&6O2G))5(/C .;K)X9Q
P][D3TP789 T_D!5!I+Z;*]40*><=BT*5M2FP:^W;;>(-6A?!K,3/,R&;TL8,I G8
P:#CX:LJ6S'-R8\N<^EW,)L<+3GN$Y<0?%"YRD1I0-DF'0:*(H',L_&1S9:)M?.8Z
P(FO9;''X])'@XC48"5?%BW>#1;5>>1B<^J8Z2R#K>_N!]K'A\.2;:,)0&N*\<U R
P98C<+J#&26&T:K#AY$G&W,FLESKR6M!T/UXHP^BF%I;W+8860_]!D.]8T?@^#9RA
P(]Q^;6<#HU/.$*O-";XX$I]AHI'Q;LH%<4-5M"656J%YW!T@IT]+=@&L"AG126%R
P:/JSKFW / <I9 ZLU-"=)$>-QH"99OY9Q> 6$<F7)$[N?:W\4SX5=7C=R*)ZM7JS
P%8"Q963(XF; N2O(6U^-4UB*\[0_!49@4YM92HS2QE"-K,>LV)EP:AGU!'GK1G-^
PY0Q]RV]L: [94:R_^%0\<1#:%O)T6&"8X$<C ,4V:B<$&83$M7R(H58ON[WY]U>L
P'B"FS-7$(]F2(0@\(F$E5M<%#)=[HJ"MM3&5&;QL/)->65[4A(8N>^;J\L8[#Z-1
P;,C<8C:#P3VJ$?X7;^5CY"^&W23P^V]CCG$0 =<I.<>>*2R1;HBEHA&8.M^3!C.Y
P54H+"/0+"@9XSQ.+&#4RPAM*"JUQ0%$0(,=^1R*V)D(GJ%=-]6)IM6CF?V:799;S
P)-)I'1:84H+Q;AZK(P8A8J]$)ZF7'(\%N46D[6+%R ?Q-+K9# L==!/5=QQ#8T9A
P.OR9W@G#U+\M^7?0M=&B OMWZ%R_!Z8YL+X"V$9]B@6N?2N3W&IX94-),L'T>=)T
P\T,&9V@F!>R9"<$N(A3#GL>$>"LE-F[[.V&ZH\0D.AYZ<F%VW<A:]!!Q^MMQ(;V0
PT5ZI+MS\6>4]U5)7^D1F%6)#F2E&\F[*9'WTM.35$Z7P76D;C_5WZ]EK8'%Q[)$E
PC_]_<ZH$2*!#9991SMS36^[;[>_6TVBN/55#B_16+9$)((VY+"'@>.P_O)YS"@3G
P9[]YT&V](.-9 <B@I&IXS-I^+/=][,K))-CG;=C]*S+:'C'6PR.$AZ<D<ZS*\7](
P4UX1LGB:0K;O)GR#^LL;X+-H!39+@YV3H,IDV3K%V?T;9.VWC/<H"WQHW\F1G"TE
P#T:^^$>+KI>"B%7E9;H'RDD.IBG:W!9(@F;7R!4'^>7@WKC<@JXX6K,C;[>"C4UU
P+\V#6(M!KV81N*5(-YXF>SH:>(FU#BF^H"KZ4YNC)9I@F$F2K:EMA)5LGJXVBCCH
PD7FR_(6?Q0W3L0T?LU=S4&]MBI*OA-))XX.*<DU"$R]E#5-?98QY )3$ *9]C9+&
P5Q87C?1LT<%WFC$[4;FIXZS<Y9[:5,PI&^<,<ZN()"21+;]^]['BJ>7H% !-'1!J
P6("7S<2G%=HJ;$"6"J\2J,P]-X(2<I^EQM5'!A7,*PU76\-8POM "2.RU%-G)^UF
P#53%B7R:OGVXEVYD# .[_TV[\F SV\(XX)LJ"_;YMYB/5+/DAGJDI*'K [U:1>+#
PS..0W'JVEG&8'PS0[(-EQ/\G&'UO"K;O=]>^IF.C,A04&.>^+BKW:W0_?M&J%U6]
P.SP ZP;K=J_I4E&#,[[J[ODI:DYY17$3FI(A0-,(P870%HV:L),GKL=]!?7Z%^1Z
P:9;_S;*D$ZL>:VM_#=C,P260=T2D<2",WR@("C;]L434,'\/7G@I\RHK:V"]@PSR
PVP@DI8L)Q+U:S(U#0Y'(:TV-7?+PLR@ =;LOQ7T'@%F?6XD<>I[;,6#X_ 3";5Z<
P3P'6@-9E^/:E=SKN@"X_%JQ8Z J@ %G@&8)XOO?_3818L7/["FC)@;T>Y>!/!V2F
P_4W@?5U3UWHH.R$+>;UZU/Y;E)(K#RL'I]P7T$.'^E!T:W8A0"UO5J:_.N@B,'?^
PD"_2N9DWE#PY4[3L^ '6=J?J2B+BW?;A5J/WC*"3W9XY,I=H. KOP@[15/M-?S1#
PR$;B=+]AE9S?CY SR@@Z*[UN+W[--]\*'DAXC[J#M0._&[ELAL ;M]LS,LEATK=V
P40]!)B)<;I& #)S.^G;AN#FQBYDYT3#SMPLJ#89&A2Q 9SM4KZ9(S.F,;5RR_$=;
PO2MW?&1Y;=/#-<[[VCWVSV'48'B_%I6<T$2WJJ%T"909];HW,9*5I6'WV.PC5Q7%
P[L6\[#6\$R6.PK*F3N0)WA*TMU;K ,:8YYX5?3*^2&G\!J4#+VH9JEWK9X9EQ-^?
PMNJ(1HYW*5$3!?J%ZC$L5I>P(//.]3:/($""JZ:!D5RE&(MGC6;YK =C;VRO;' J
P*>83SN&::75RE'O7=HM87<M[GU:N_9ID$<X3*_C18%MJ3E\1,F5A8=R-/"CP_&T1
P \3KB=E(T(A]BP,R-CP@&[;DN52%Y+@1(R)?]/[=!SW?_*?-$HHF:>33MU7^OTOV
P)W [2Y7K/_I3.53G?-  HM(1+S^:DBXELIL2I.NU[.=$>^^)C]/?6,A \T;?]R&C
P2 ';6/SZ;#>+_&=3X_]<!.'D1CVB8:D*X:][YSOLQ4OD!S._N#UGPB3S=@/=9140
P[ZWR2/ZK'T1Z8W?!6P%E1K]CR0!X\3G;Z6A]G;98\H@\7KQ@XMN=C&Z/\[\>U:WV
P1S\X_9!=GBZY6%/Q>M%>88/H^/HX_&N(QPZ=/(0,K3%>0G4\4PI#:]8K%SU'SMUO
P->AMDY4D/P8U>-4:]Q9FR?,JO?AOL:,]*J7DV&>V_5GXL:LM4-:T([081?!P/@!L
P@ I,K0,2G#O?EX7O6*<7L\]_V%KJLA!+1V")<9(\,_-W 6+P+@47QTR[!4)P#FV@
P7Y(&M?0O];/Y'$M,Z6\!&//Y5&++V3)'B\AJ[-[_)5VA*DU%#XL@5VR_IS^!DK(R
PA?#B[4:.G?CL9(8"HOFY38N-!(#;O0?V%\LWCUWL@7_1'NTB#_2@0)<UE])Q 1[H
P15^M2'6*$_];VAKL+D ?P&09D"6AN)-[?M'7$M/FD'8/3ZHQ4FH>L-<YDN0JS[MY
P"Q#"DU=C8X_(>"M 3C';OJ?+9_Z?>)(2E+'50X<G(#ZLYHK,05^41'=#I$&8G7PG
PVR+EZH/2V:)U>K<<W5-RJ<8S#4R9"T']W38>6M_Z-]3DXSGZG71CHLVV'-V'[4#.
P)EIV$8"ZV_H?E4.3*_K_4CJ%VQM&+O>^R)8XZILN%$8J;6X13 TZD3+BR0=)2P5I
P1"%W"(\^4=RZ_?EHMA:@H4%SN-@C)JAE'U$;A*R\R,]V;'^6EQBC[6O*MBJ2?C<O
P+#FQOHHRANF;F8F7F?09+0BA%@7O$$,LT7M!D)#,J?Y?$KU(7Q 0BJ=HGNAPU&[/
P>'*R(*9@=U/=!4_^=0F7&_CF%U\Z;[;"Y;(Z'N\]\76=/L(IT:6C*Z=<\:4.MB'V
P<9VBL5()J7T5#B4#_XAT9:H/ TO\XU;[DUS#R%,Y[H^O5V4SX].RT_3BIOC^!I)R
P.?X?XLZ'CL#+F?#,41KV]I.$EW@J$$0EHJD*MJNOD0=<6M+0(=@RT%T@5",!.F57
PO=/LA 3+MB!?_S8(C5#(>YI0)W)9I64KCEY!\N1\U9=SSQ;;K15QDSAE!19@4K1/
P)_AW@A^[!Q0G82L#Z!^FP7"P^9I>=5-/4X1<#,?;>:F49%0FUG&*VD"74$<#'8JQ
P65['#W&I(^%2+T> \$<,DEI(HTAGX/6"C"V^<36A7)*?,XQW:O'L_W%B,RDIUOM'
PJ*MU?.N/>YC)<F6&077R-77"Y_"MXDUZA./E\[H8!%Y0DGMR6W9GW.>SW<+4O!21
P["O\#=F3+.E<4K_"^%LLL)C4=WMP.*;Z_&@;U?XURIQ ,IEKCH\]V"MW:Z]A<:[!
P*O3)2'GT2H2NG[,W=3EO54_/PBBSE1FH4P*9,WD^7=%\.U(#46M7#&)KH,;"ZYJ^
P0V3C>(-Y:W1*J-LRHQJ8_?G):ZG\9)HTZ/ 0C](F7>]R[@Z;9/362/&]*T0R3IM_
PFZ\(.%S1[Z0E&=6Q_+O7=?9J]0>>.5*CSFRE-_<)#@M[!GAD5Z.^BW8EA>E.QFB*
PBSH+-NOZ*U"E@-SDKZ*:]:EZ-)2GSG8B_I7"HFB"BC+:&X:5)EOM*.2!DDP,>=4'
P(/;R2%5HL[<#[A)=ZC7Z^-(*8//,XU4G%;YU5' L-5E"6.+@]:]I/G5HNPZQ05M*
P<?S)X.NZ\8,^X,(U,)@:W6W3@E,16!"M%3=>\&E;OY5.A^W&N"?/5I]4]B>D0%+7
PY6]="I<7+OFS)^B^X,]H^;8LB$676FFW\U&.P,J>19)RU?F)Y%+ 9J*<AV98Z5?J
P9V^ \Y.QPJ$(Q-F'1+ZM:=.LC71\/3/$(?(/JX^TTSXQA4)&S?D4E#12?]K"<SE[
P3#FH[0,F8$O,7H2U##LL^L&:=]4).A:M9ZNC;AB6ZX77_SM.VV42 ^N?>$HX),07
P!T:[2N9@B4]6'_"(O"124&QD*F Q90+RX 25X,+;-3,,S;9,W L0_T5Y]LO>=NP#
P_#S>42WV'3!Q$S=(3',G0MYS/RG((COR=>!N5XU;#,Z4L>^!9T+'W0#H=.[R)84S
P6K8;TN9<"Y\U1J=?::7KWI1U).O&\Q(7U2EV6&_LR:Z<=0;AS=L7B0LYR_!T0\$.
PF<1.]C'S(]I3=YIF"RV#0?H>0:SXPA^5P9N(D16,8(?85()9@J?=@82#Q>3&]W?N
PPD,2/\PU5Z0M1 5R,IH>*8$D:E@;@FP!+]-P,4YAWXL66?IHV%-=:]-6S#0W!"1Y
P"GQK\,A^-FN1HF) S5.T*9!0%3;('+H6*Z!F)04HV8F *R"S$5!P[.]3%'GE#IE?
P#;7E"'<4/U\3VL,Q<:(L0))T[F< Z''> )A-4K,O0S)6;$Y9%H R.23W-TQJ$7<#
P+9\G&+TTZ;AZ'$5*DU/KUI>IL]ESNY=)T&!\)E ;]_A0+TQ/SMWF5IGT@E<SK@]T
P%S(6M7XF1RF)1])N1V,B$:+:'P1CGGZ).P5'<OY[3K) O+X!^)W!@$./GJMA4_%-
PZ(O7]*G1@'D+MBHT@N:5AWX69KOS1E:BUB8,-],OS (*A?PZP2?ROVGT0"F,61#*
PT,4G&*>7K[Y.A=G;NI]O<!F2LF*F?%\#O&>;F$MN\BYSR3ILKYQH>HMH+WNR-PX@
P$]U?W"B.\<U+QQ)VJQ8XCSOC*W3G-/Y9R>GL8#W-O%SJ\O+43R%*.&D%6K<P.;(O
PO1,#84RI@SCHW,O^J_(YEE?OHS>-:=S%K 0WP2X8G)Q-BF^_]4F$Z.L_0+T2]1:7
PT"_#T<*F6K$V"J!^F@5$TE&H_6,YA?]<J>W%'Z;-<G'O;($"N2:_N?B@GPTO0?+@
PYJNW:M[JENC6SHE9^>H(KR&5"4CPR"A+7>ZIDZ2UUJ(T(.JA0O'!I':%5;+K%VW;
PX*7[.EC=TK.XOBQO1(E3IW-H7-< HT3V&FH3GR((\(F7:;>&<(9NR>92@U&4\;P3
P_3NU2<C80((55'E&,UI 'S!P0>Q:=M7L/ <1U@\]N!',(7X-T(<>O<>[A>Q+QX\ 
P\@5 Q+AF%8[%3,L%-RS&;67=:E[@<7 <:F@.UC-;GHW5JS"_6= P4"C!DT0"1*UX
P7 CFAC$Z'*8D9;5]A;%\@0EU>_@E[;8QT729GK6L'K(> =TLI<0#BL[CJ?J?0U['
P:PY3 G<Z=<'<]*'^*5$NP6,JE^[\RTK&NRXYZ[>\SYSF'K5=Q#&J*"(82V,YV^*4
P1=JXXU"TX?.CR@$T\N]TPS?*I[YO? K,07F>8NM8_LES:I.1\@>._%B->0&;6D[-
PI/AI-Z"3>3*<H;-X@?*Z39P>I0URZ@DBE%9Z&'S4.$GFJ_[.'85E(XH4?2^V?FT5
P*=- /TW0#YPR]L!U(.D7RL8K0HNROB(;NN'P!6;;*-W1^8:?)&94*-@GO?Y[PAN-
P.Z!=_L0QW=.\S!GDL2?Z,M&"0SC #56JEA#M+5=#R2!M,VH6F[92N[RY 4J_X[Z]
P?VG8R(X?SMGX?T8;'NJ.>W-]R/(#%&6:%\_8*)!R:5O,/[+/SD%R7LHK:52+ Z\?
P]U%X["E?TL61*/'W[F*()=\82;KMV4D:6H?6 -+"&27OD)"7B<K]=_B7$ )B3Q1-
P%U81^,#Q[%UU^QX*8-S#?RC*6O8*"'A&<4*H53V0U'GLEP\=K'O]CM/P?T#\R(?%
PV+%_\GEC"J1,X2;9U]?=0MP=S#V%E7O;FAS,A23&,,XNSM.LX@=DDN4!"%;O&1M0
P[Y,A,$7'=PD%AQ1 ,3L[]Y1A#<YS+C?P,GIG2[MG%@O6BOB)W>GO)<1<W&PX)P=1
PZ[=J7 4X<Y[>0MH3/IC-!#$.J_4P),7A'0!]@%(P(Y5/TBN*:U;RUM6./ RJF'].
P!A*!MI1R+W3SH^QD"K+#9DLX$, ?(ZE\"XE[ -!<VJ5)A'K$:K>*ZT,S?_,L>[^I
PYUBB ,R$LZV7Q6>T:SP2M>0$#R_*_<A6EG'8:'][370HRER8@S)Q>-[U4NJ$VLGK
P+(Q1G478=8<$=(<3W9,R=.TX$8B[B18AY:5;J\>3N"'<83I\Y2;"WC(*9)BD J+<
P[?TGCLN!JBIP9F&0DIOLQ>5&XD8_:*7OH[5;(Q_:^Y"EGU[(B.YG<O$^K, 294ZO
P43PE57-R3]V(,ZG)V3?F$/FH[L;/<#OR:/)*UQ=7IY!4P_.YK;N5C'MT\BOJ!3*J
P_IE6*;]D!:)Z)Z;PPU,+4$VYX94T3?:#U&"QBKQ[\_M^@>J_ZE&A$T\WA:,3+^I+
P(J]73\\B:O M%PN"/J= =="]9'FOWQ66);W$J'T#%"[+5U@;Y')<G7(2!NXT=&56
PD][FB&'(!#008"6FJDM@+&Y26,NHUBP3UD,?3W6WKX<D<DJ2D;B14RJG(?%&XB>7
P7ZH8M =7X^X RC#BK)C7M+WW;^0S+2N8<-LM%U0=IJ.<]GZ!"/ Q]6QX*_O.YMV5
P_#A086Q":70 =^+2V?%]"-X;)\'6^X8-&$(7&1"%FDI5YH(ISEG4+^(R_YUN?2\,
PR,K'S>/@7'WE.AB]B],9MHG,D8*)?Q:(NXC9WN-FRZ<*>>U:,TV[@J?@T-)CTPVK
P9G8*:L2:5=\J.#NTZ9_0;(9POV2SQ[13:\?B *S3?5?@&U^^6FGEC5$?U4*AFV]+
P<)9HLE&6,TZ__1=U:!FNF^+B2LNI8_^@=(W"BEG;B2--$A?K8N">@*PD@YFF\=0[
P92?(VDFOO41S#<<BD'VDF(S)W_I/.'KD4)I^VJ9(,-5BQKB<<!&TVBN7T#D/)%<V
P7Z#N'?I<U1XC*]/9_&<^.L%@V ]A Q#[_$)(VJR/JG:T:.RE2$P'T=5-Z>_[8W6 
P_,R74R#4(YGN>O<]F":IVA\G>K-]DCE^A^VL^B025VLUK'%QE5WRC["=<5SUOXWF
PC08OP0)?@B^%QR?ZZ&+MW7R61J'_%._[+-*+P0MJE<E-92 9D#=JHA"-3,H2<BG=
PXJ8"LE/+?$,&@NC-M3@Q%%Y3708L/BH;1=-;;.:%_,^K#B82&SYB_L>_\NS/H&9/
P;%1 F0?:MQT:J1CU![.7]FX8^VY&'16SBC>FC V&/J_[L^T@/;0_NLSWO0=%\;I 
P"@@]Q3\>*NK_!-84;Y;_?K@=_ T$ ]]QCL\9.]3LW&P0P!.'&6AB=_>_!K8K)BI-
P"N!Z%;!0G[_"+1:>BW4D_ZAS$<A-MKJ:2=L_AF4_;/VKYNATG)3 W8#I9JQ5POIX
P%=>@0%^LMRW'KD.]F.*VRGY$R0E"LOZ]MCUU@7;#RMVG\V30VM!J:B^P&,5Z H[D
P"1C6-LQAVRT?&\@':]U8V'#Z _#?@B+'>86A]PL)Y7C)AS_POGE2YFQ(LEWQ  S#
P?GFYTM/A?!\HA#/C\=>?3I+E5ECR#9-< -<O3E/,R1Q%#O",B.M@$>I#V[U*@(45
P6XR$F$Q2V\E65KSHX%_8@*TT/_Y\;C\>D&I(!SU[U^TH#M\((7N\_&ML^-E>2F \
P <;7.%@@84<R@!/>SJ$B4G+7?2/"+U%#D(\IU^<8[2(;7Z[^V#;R&)$J3)3I!=?_
PQ:Y0)K?9IH,=2"=23=3EUL/K"']:YN/=!=?&WY8+BT5ICN$ZV,L["&5-Y'U%QM(+
P[OI%_;=S'G)D%;TV5KU%!B282%.[1%C\#C@810?HI"HN=UA3<P0F#HP!_)NM\+H&
PD2*:I,$LSDW6>N%E1EL:)/2EW?MH3HAHI'A_T"@BKNS61M($BXA:RF>+Y#1F\'XC
PO0.,TZ :\04+Y@,3'1FQ-TM.9TO=XE524E.H9U _3*K;\3*+V&^+4J%OR5;V8C01
P"$^64T2P]S'S_^K*S2U'GD9/G;1H ;5^J* W%YP"(:JD>%9C57@ A"BP+)TH9N'8
P9FR9Y&+PTB:%Q(QF(6Z=')BQ&W35S3QC?$;M);SD>E'_P'_Z*<Z=6IS\YD"3*!W;
P:+M^QC.4PYFE&1AM33*I>[_(:24MCWLW*9XX459"N&4;GC].[(J.#&L1MP*&4S!+
PK3<9-SQOS: HX/L5E 0"7?XV6 >70W/?O%:XU,MVAY3_&>T$+>^$3.T=7#V>T)+H
P*V-)AH=]2(MD@<3GKL&G!FZ)(Z<<)Z>V<WQFZM5994BW\#KX$"! MU/*76WT?')8
PX04*5^9K59#$-DZKH5E5SFX. L-C0E:W>KB]3=VI-'!I<_XY&V"?[_=-.U0*M<'>
P@ =?2J&&/<(T43($S60J?/JZ8X\;UA::"C=1F_%M[!T[_B+*EG6A,$JF'R?I[K_G
P_-^** YX9MXZ=$FUC<*+(4GDB7:>S.WIR^2!8#&$E&P;Y5@:9RG1UXM:_+_U:(B\
P)*EFRMEQD3M90=$U:TH_G3.3@.6Z3%,D*E)R++A@C,[DR4U[JJG)2JM+ZRO'KYJR
P$S"]8(UEEFJ%K-M2IEYU^6D*8@Q^U$]:*E?Y5'QZE%P\ZY5FJ.BXEGT=,,V=&X*%
P<=>,4Z_(_56%5PJ6PXA*X[)%4*<2JU,0V5NZTX?9>E(9 ^XO@>F_8:7@\%W522LY
PY"Z8[VO^;@JQKHX \?^00=+?(_3!JODY+30^FH10.VFFMV7 L, ?^"4,Z_G7JB"+
P6+]@A-((KTOHIAOY(&_DLTN3_I-6@QC,1WJA3V6>"*0\S*@R*F)#JV?"GC RN4X\
PKF _R%KVWCD5NFQ$:!^I:2S-H2@FL^6!%^T/%OIQ!VK#*!03UC;/D OPQO1KPUBO
P^X5^S'T1M?'[7GF];GP?GA4=F:"A/*<1_/WS2UX^9P$>D1ZXU7-' AGO'&%C;DF@
PE\:.M<#M,Q/A^Y>9Y.R=SEX"DM'1T#I]&GK!5@U/] 0G0X<59OAU8OE2.Z02A6VU
P&K@>[-R5ZD12,98.W+C9"L6N3WSCD'*D\.>(5#RZPHX1/5XD@Z$UJ<IV.L]66_F<
P'W&9%:?@I,ZD $X.B@W0#>((:0NL,^59^H9^;+ZY!64D_TBE\_02J!R=N>X*V :!
P ),5]M]Q\];Q27U3%+Q4T=[  0?%D?7H?TPX'\%T;[IRG<D'<$)('84F)EO<;*SG
PD_3K!J61A8DDHM]FY-(?D>&(2BW8%]8!^2_&'P33Q6-'XY@8!V0 )[J#O$[9=ZPB
P?3(N@DJJ-5;%!SI?,ZTHC\?($99D=]OL.MM3_-J$'C%]R!X_-R@6Y\?0"9ED,.S'
PWJ8 7/U]B)SM2FD.*K#%N.JOGF%T*PM (L6Y#6%%D;J$#G:I!\",C&&#3)D6N@)T
PZ0&!+S?O&S;-:X<]4W*Z%YQ74K';OA3150S:G8E*M#5M(;]CF=V \+O.WQ#V1K"9
PY<#PI%2I*Y18Q]^2CH_4I(3LRF0$+ B;=/2-8RNLX2,WW'C[NM[=9-I5'\KA6"5Z
PP56!&8[MI-I3O@M.(I$PRW8BA?LN]\DW.D_^0G\/I[C(!_] _FY8TT 'T Q1,2S_
P1YV3$X]N?<>[_VDH/FP*>O5U6%KHRV .IU7/_NCACJD/WT+3%UJ&<-REU[TUT.?E
PSA'4-8NK7T/X87/ V+M7,941E$VV"3413^6T]X8 J'N-#)3^R57[UXWD2?RL>G$(
P1<,/+,(WC%XK5+:^(QF2,-26:GLM%?,D$,7"<6W=M6P%/25 SNT6;*\CSX2&"K7\
PY52_#8WDV^EC=(B>=JH&%70D4+Y!<*$+F;ZG1[_[@-U<1FE,DYPN8>#1.\_TR.%$
P!B\M&*;65[ND]M5'I%!#%-[6=[E_",+)/?3</TR[L^3QO(/L0(-7/7+VZ='A!4)1
P:AM95YV1KXH_LJ[7GO.;QHX</8#YC0F'7:18RIG9FNT00H"\E[("IV374GS*=H0]
P4'>"$6>^@IFR\?(C5:R S=MEFMHN2 3  H+"$Q-^J.$MZK^[?F%#S>Q[X[-,%X>"
PE4ER/A$L[$+G9>(KSW&7(,M#XHR %$1W3N(R!_D51 &2XH3L0\+%LF,R&U_02.":
P1(<$U@+A$HM68YVD>:'6'&>S70A=%28;GE@3E"94I.:V2)GEJ1F*3JUCU=QTNSJP
P!+F8/%#LD]"6G+-=KYQ/?WY&"HMMM\/O::9!Q;1 ,D'4E06>QX]_07CV9)_+[S(T
PRJ4_2@/*N($!A$:E\H-$X&M83Z79P&BI/TQJT4<(VU^M$O[W%QCGK8/ZRH9 O=S?
P/ZJG%_I 2L1K+R\*HO.)3#74X^[(+65(MB&.(40V9 _>LF#<@J.DT&VU$*WO,8Y]
P]8">I(^MB2R^@4 '!NXGGX)V6L3\&=$:]W;&Z6\O@LP=$<Q?VN? @O)5>?RF[2[X
P/_-&WA>>QF#"L+D-&-O+W%=/\+@"WX6.M3BRG]9.4(_F;HE_$).>J(4I)+AU)O&H
P@)#%^!OT*GSLX=$([/.T+8FI92(IR/E)A2X2:OED&A)3[N@*!I<;7;GND'=Z!4ED
PY#MH%&%<"3[?CKP>Z'=7^Y=[LE+<::;QS8;I.OU9QA\#3>.P25DHA) O7X##B'/(
PL7>V8GE'?L?#*1AJ<R\G"X4)?FO.Q#3TQ6<,-"W([0\Z17F?OMZ-&U\6]'S_=GFD
PB_*'N5T?U9X]/X07Z0TC@"362?J2JIH7[W&&%LM9AC1*\%^8O)6B=DO;Z;Z((4Y)
P?K,*!Y"3[:3GHRMIX :'1F"><=%F1](&[_V27SVV.YO8&VK-F'$3[] ;WK3[.JLQ
P+JW$4EJ5GZ=KM)']DIG?-\^FQES62@'28.A/["?AARH0.AS)P7AWFQ7_C6L<*]D6
PD*+TU;E3,,H3[9S=PR,[SD)=%Y489J&322P_C+=W"I/U52Y%([_\1:'ZS/ J,1GU
PB\+P0=*?JR";&_.IDJ/AEPNHJ5KMUFE<?$DICBE?. E5[FH5-3[7AO9%?S,?IRFP
P\7>Q[H)*XZ:75V\]=Z]2%FN'[TOF0RJN']U$4KDRPI]5T"3*M&O.B4[6K] 0[L</
PV&Q%<HP]F9''T= QI+#+P,Q&Z7N&U$W&"6*0]T:B)>$6E_L909?([A$MB)<<,$;6
P-)(2JD559?&PV8@S=>]$)<, 1H1 BZ3*5FO8?R3N]5CJE(6> J3XP(ZJO5Y??E,Y
P"J7%.D)!:72$>U2#68_-\ ,]>$V+[<Z35*^,N+ +;3'V_>QM]IU8_0Y74 "H6R.A
PWO)8LORG22@F8I^D_2X!PQU&G$LV[_N^6#9$W-INLF"*JE!K-EX#CAOKHV,\M!F,
P-_9_9$<<FU+RPYSR(1D[9*'QR$'F0[MY]#E(H'6BEG>XPJANY>"R7LV@Y'<&G -4
PJO5Y#9#N@1*CW8RF<#ZX,/Y/M/5VKW;MFNE0H=5@A" J,BV]&'!8U6GZ.EO3.I/H
PL(XJJ24P^C.5QO!:F3[6KSA\\(BEHJ">?1C%5,IGA0_+)VS@Y_X_5URZ192L_NQ!
PYHF4-9-ZK%6P)=+,-M3_'^ [W/3I5>+VC!<M<LVHK243G%O\,.I2U7)X[,P.3L/A
P:#$4+;892A\ D;KNFFV.54][AB9UA-$M&=[DFL#=1SO&9#MN_CFZ^0C4N9(7 I[$
PN;/I?W2X-[X!1QW>_0+OED+$8U%A*/(>>LPVC-<(78,P[++CH!U[WI6K2ZDU?'<&
PH;:"[^5\Y")U,&/Q$)+]NFX&A"%F JXZ[YG0*KD$=,CKEWK2IUIR2=E_S<9H-2<9
PJ26[T_RQ$B4@-GO 1VQ%P6&OWX.#*,WW;W8\_@7<OMY<!KVO^)%;]>YA*990SVII
P6#)')!;"FK<W%0<IX#QHO]'W++^Z(R$>&H#X511<%DB'@85;*S;8C%00#'=E%F"K
P*>O/Q[Q8X'G!LI3UG0VU-ZZC#>;)\;B3%\CFW?-L4NW9.M%X70'AU"9/X'&&P/<?
P/'TR;H +L*%"$H'-YTPR&X_M%>N= S^$17S7KN1-R#=1'4I+)R?R([A2!#<.@O/^
PSQE; 9\%;PTP-AIAN9#Q0RJ*YMP'%<:)M!JRCV/19J95%C2-"I\@;J:CJVAJVR$5
P$OQ$0\%#4A"YB!(VU/EB-8ZE?07J=5ESK"WAC$W_(V#Q"_\_)#%--;L9%,X4X _R
PN+T;P!-8\+]JT_Z]/:='!<*O1SH$J;QA0JI>CS+%@PW_#>]12%ZW <#].S+ZYQ-L
P$9D_^.&\W"3%$&VMW1(/LH^C$Y)L$%>Q/T(.W#/35I4HQF&SR2UE[^,DMTECL6GU
PTUBB0@^;>P88JZ7FQ!N7;G>"!+;GTA#3,GMS&#E>F&B4E80'MY)^6[G2%ZD+W$3U
PTU;L3?[*D/K"6EIG9/RU25%+*;TY4+51 77/F.?LLKR%J@QG"P"__C0#/X@"'L-D
P5[M32Y3<ZH2GO!PK$,%7*['Z*CC(#-8 XJO18TM/*0Z$-1%&BB'FOS?$XE^&B_HB
PIR070*>4)BN"_(LK9K[P7>!93;@\;'\_C>^COM<Q$=0-ZVO/^^B?WP9B0OAW( R9
P#W'->A;M+/%^44";;KH=LDHSV$WQ-\VT-YD8JK4EEJ>*DO2DC*/PS.T:I>[2ES%$
P:DIRHC2TY,T]YJ*(W;Z!'"TQ/XPC&5<\</6[#SA,'4 ^8VO 1:=Q^0]=$6&RDW&I
P=%MI,_G[24X' D<TII,Y+NIR;.QN\5QCV@$W=&\!LDT!J@[FX\4\JB#F^QFR)SYW
P1FSK>1@KC..?&;R>K,YY-CJG#]B%O&Y -PJ24+.W0&[YCL'7B7H:^&^P)^B&WMBE
P26J[Q*%=X.)GZ;2]GX;%:2T)X<1@G<K]36A((O UE9*(UA?H@)'>H:LT/.&WBF+4
PB#UIP"T8E53(HH.(0M_CSCX""$;JLD4YGN[6I,:/E$NL?F8;&$W^9G,&'V\5$!L_
P:VQ#&1)INNE(KL/:3G=@%;) :#Y?'D/<[J-2G*\;L7^YR+4$JWFB7S5O6TW%CQ  
PV1_]"*O\JTZ''N.) QF1I1?H1E!+$530Q6?Y4OIUG1B\VZNK5O:0LT1(B$H>W"(7
P3S]WS<2Q6,EC*+TB=RA+-,TGUJ.M>\LC%%M"<(6[T9J2OS=;"6R :"EI5IX +^NI
P2 E[#_OC5?"J>ZC%'=CO1.?]@S22C2,TJ=K1M/Y$F4<L'YNS??KH^3Y)]<2J&#07
P^/F,R=VPAB<()>&55?SN\@W"L>=LP[NP<'0**(E/"#YHMK-+/P0<*FC0D;&%281[
PC:RTNHMU-8_\\T+-QRE&AFTGM5)%,S.UJ;YNIYS(:&L/@6>_KY[[GKYQC:>RA?T(
PGC;6P@B?W3Y?+$Z1=\=$.;=-S272]N:Q4+F6*7#,R^IS)P_:C2?4Z94L^C)7A K^
PV1&%9G**!4=L"W"S6X 8/A9[DC[AL]W"1".L,1%?W[X'2YHR*T:>6U^2_MR')DYB
P57ZHNN>;!D2]J*SR^D=XIV>@/6(6WZFWX;F&2+)_U@$7(L0\ 3EKF.E#<7^U&R*H
P_QP]0J8$.X/]55(._EH[F8J/]'7K*9<IZK5A5RSW^_7G-NTZ6:2G1]J,I..OZY'N
PULW@6R?-(@V6B;@T&T]1?W.?"N#(<*/1C#$=?J^/AE =9U!G.L?5T7Q17!Q(#'F5
P$R\T]+%?<$/JXE:ZGN%SBR]&U.G@^!+W[DLA;A@*Z($0R9'279,0%^-?]W??IOCW
P/(=GQ)%IW"%]8'PZ,>;A$>L"TKT_ '/KBE0YIA>V)>/O('Y_Y7>A_U2K.HXNI^M2
P1E8#X&)/]^WZ;S#7)Y\SP7N_>;G#TM=,"84<%<F8*S6U2*_ACJ^[I;A8A@ 7G>)+
PP&/4(^9.3AH^*N/22GMUZC76>>/RSQT6 F/5>)06X(F;WM U^H5@=4<<&C\Q6'DS
P- G?:A"J!Y51ZT)F$3!^/%Z(J/1K/Y7X^J?"X\OO9!4873;KQF&IK%7L\Z.=0X(4
P?^A(;\R%?!\9;%_C.0O9"6,ZF"W"R6WS]#F-+5XP5&%3#G&2/YS?,N CP[T0 !_(
P>^B!ENX8F/SO"PJ(MIE@25(<U$1R 9ET)P DC(SLL)(Z+QS:D:WJ[#_A3%A!M)K]
PWXZCP:)/KZ#4E!O^[6J3ZC JQ;.]_5*"RQ"[^G<CQN7E.0*XZJ)[/>D^>83YC<A(
PF;(P )P/KV/;GP]]NE8Y!'&.\O@^$#3FN4W2DZJ+2F;QW;@[!:"E J>L-^0!O/]N
P.-\.&_/:6[)WA=J79CRUQ3K;(,WM8N'5$BGI['0Z)B<A %$L7P(+P27X*Y04F;WR
P"!4.Q^37U%]JEHXWWK9$Q6<>)5+A5M8N4;?[=7O0&<"/LC:"_R$K:6Y_:OW3L,-S
P*S]OAQM7,PY53NARKH-O:T=G%T82R%2_X->I4FM[V.0TA=N'QF[??-4'F[)IQC29
P*ZVH:(Z06?B;(X[MQV?T,E](A"K!.6!"LAD44<\DH!N?DX'2\P>2=JDSD%J145[#
P.7=R2J!S)V24[J#",@MI'L_A:@]2C..S _BW1$2BX#X\EO-[47*W2+Q/87]7Y[;%
P;0PV]NS%9:-PG:'Z_L3MS6-CBLH;[H#:/6YSG0R*X"OIV5 #" >BD-;% OQ)BP&T
P?Z"GP5:S>@1Y G)W*R6@YL"3 >OD:.ENYBD*?)=/2/8E,U)P!Q&D9@%@H%J]]%T[
P:FH]29I%94DQK;G)B]!@W".YF ^*WONU1'XU2%//C]BG7K#)\Y!#HA6K?:F>KW8-
P$!E6Y26F/<38[(D3(^15]886N?_37V%^>T,4);IFL\B7BEY9!1_6^XL;YVZWCJX^
POZ7:S/;V%SK5FG>I7C^LFOEA'%;IHW6VW.4IG P_6\Q04PJ@$,*$]_M+Q#5T.1PM
P@[;I=.889<B4G2P)Q>51B3X_5?(O>'BNE.]/\'@]V!T4!FJ/8TJW/]MNI7?,XRCZ
P87V9FYM/G7)6AM$@HO>N"=GZ:%46-M)XV(JQE,NI:Q74J&E7.+Q;5,H6=LVV[@(8
P08@''5OL$=AO*!B!=UIZ, .]$R]^O&-+AA#]QBENRF[?$Q<M=;(9PH"0T:7F2H+!
P4$@8MVH4#X+9-HA>?'7AR7&=AZ/B<&E&0FWM9S6[DZY;V?=F@F<)F"Z##3V .0\3
P!AJ8?M)7";[$X89S"?PXSB[?M:/(P($-U.LSH=SZNB-?0SV.$?'Y<*#L'GT1N=W2
PLYJSW8A(MKA!L7-H;>YW+NXP=;H R>JO!^BU3C514F2DVGG.]"SSCX&P^=A'Z!3B
P)Y70S\'>PC+[@%-\OOKGH22V'ECA6V^^*F!IE@T3 4)L,.83EI?<B)<,2[:YTTN=
PHDFIY(]&&8:9+YM<2O1HWD?=2=JJV&:TE\DVV%Y??KM9S+[>Z!T *8Y66-PV>\95
P-FVIE#BZ]!V]IGL)*TI#07*=2)GMZ*;*S^X%%9 PW]V7!7U:M4>>_+TYP,>594$7
PVI0682A-)XS+GKQIC(M"[8>>!4KJV3\;IFL507&IYEJ!-1F#P:GZ:_T>]^RS>XRX
P))MU8=Y&D"+[4P-_1"/#G!^^$-&PQ*]MBBWRSX -+QL;>^3K+$D JWW6>C-3[@TP
P\8%GATA;]^ )M!+:I_*<'MQ:R!OVYPAUD<O"ZFLHWSMSRORQ\JAOC7IQ(["NP9=Z
PYH0L5;-&7KU+%$9M:I3MQ.[9I5DM-&^^F)@%^6[=M5MDT"!\G*<D'1&!7EZ7R4=*
P=8**N;BALQNSQBP9+2) #CO!'%FGWQ^IYS*SJ#ZU) 9J@".MO)603<?V<BN5= N8
P9MES..[<4'[^I,>\+N"Y#)]/Q4C:['Q@^*4)FM9@3$TZ4D:;7\% B^-$!1: TO#1
PPB9X_]&1,PRF^XR^FM($4!R4[+_.8F?0DSIG>1<YV<6T+@Z&/Z)1",JT9BFH98BW
PX:/NMU<<;Y 6(LBX2KI]9S[^MYSN3/R;%RB]]?W^V]'O8<5DJV\1VIHC>Q,)[#B:
P%W-".HXQ;CS$_K&.SFP>7.-?YL4]_22ZOU2WUZK#^CI7J-4K IZABXWEHW."!>BX
PZ:^P!+SEP3)?U&$YG^?H]<(#1B?7++O$V&+%D'Q2#S5K56DKIW [2%YC_)T%\7FB
PU8,PI;JA2A[*J*,"HWZJ<2@T, !@U);6J7MD.%0+-A1I$E.Y3RN1H'M175HK MJ3
PF?K801&], P\':61+$FE$9U9Z#B$:1KW-A,OUP,S?D*X5791>OGF)T:*%9"2+_D)
P"MPC L78E[6!]$&_EVI92;,&:0<5E%;8P2DHLNEX8X;<E 7$HC9\+) ATWK>"NC>
P4]ZTA+16?K2YL/W<67GFN+TGZPWX]3YG.0<]  QN+:5!@\'/X9-,EGA;KLH?;_^%
P>J1!B! DC/EKA>6WT_NI6;ZOGZ[0-ZL3)O >V0!*UN,8XX$FQ3^UAB:]N$24\G6A
PT)>WVAFSZ\#M'M,V%*5OB[%&(=UT8P=I5K,J,OD^D->E5S GA;&UM0V?@$^-X;P]
P'\S8XS[^:)1,.70= Q#]'L32S<IK)<XZ^5C?^O%T/-&FME=X&'T7U278K !ZJ2A+
P)B"%8ZOS Z0G.=VK,5I1H3<T*<;>6>HS"+C=;]Y@2S7I XP^!G5.OI0 8Y0EI2T=
P*.H Z)PU/MU8"!X@%A+RL*5L>BXBG(H#F-_; 3C!96"\JY\4(IV2D(J:_!-0#A$"
P[EY!8(3WO61X_AII@%>?_UY$'XX!B)?<]^.6!K.KL%#NZ,U&XZ#<"1)]) \/XUI=
P#7A#RKU&20V+"'XQ>5Z'@&"QVD1<*VWS^(G>,<+2\#_?/0*P,TDD<'4W6DXYI//*
PJ5K7IT5"R0)H"(,VI7#&U1VV>>DOB/-B *2?^/0T2MHBV+66=8H0]9_IZ3@D61KZ
P2\X<UB)8P"'A5T]C&-LU<([4E*I>"?9 Q64#30KTN/3KQ'4VP#6HV>29@"E@E4P)
P6GNS/PY^50H'NPQ^]0&,=.ZN/HB&U6LL%9PNBKE(@>!*T;O4X[=I6SEL1&K+"%?O
P"* UM)D0L"[80:,S?C%QD04/&0,!:SR?D2*N*/D$@A(SR>$S  K& $83F&C8B=Z^
PY]D5(2DB^*G>9.;R4(I!J(JFJX,K)ND(A+GSUT/'>Z5%<3PHY"\XZ/LPG)$O4,2/
PZ?Y(?EL1O-PCJ?\,0J]54I%!*6:@1 H]B#&?RKNP/:&4UP2QHV4X,)N.<K*K4%E?
P:5W/'J,=96\9>RX7;=NDZ]PU#*&ZG)OL?0Z:)M$H,I-2$P=MF<)T1.U_#T>&AKJ8
P1SDIH+*8$8%Q!>8;:^Y#1]2FZVK6V3=6*'!)5AXGS-:C8,/TDGOS 1$<C-ZU=!Y>
P@+9?,0UJ:%\3,(V[[@Z3ZK&%BN';$ ^Y2#Q$9GFU0;9)8M1_R0LT3O$I*J%%[PS[
P>YQ\O=;PXC$I^*XK,)2L#=,[WV)GCT^?TK/M93[IU6BA "C;/K3V1RD\?YQ9$/C_
P!G/,Q#$9E;X"F[$AXI5_S&W?"C?2-C:2:NUXC0@QGP#-GJR0^9'J0 Y]U#,MNPJ;
P\SJO^Q'/\JQ.O3_CLO+].SK7]NQCL$W$V"-52.A.NGD;:J!ZAUH&I<#O!RI6CAJB
P@HE9,421V4^/GY5#S;>U3HC:^>>)X!12)BM@W$HY-Y1TV\( 8,P;6O"7>>&>?'Z-
P\][/%S-VRF!S;G'H>+EV4Y: NIE--"+("<:ATMT@!!LFB53U4HRDB&+"!8NAP%A]
P]"_)K- 'X,Y3;PZ'3W'KG-,KW\ZLUD4\EP8J5T,#4?:-D]LJ%0)]N:3HYS!(F-;$
P!/5'Y 7'8>R8P8#@&%"?>.3[2\_4*C']/LQ3"W?W/<4>W-,N[(>^X[RXQ.  \8VD
PH;83RH-4>99VK&L+0X]@18HT[=C/*WEL:F[4@JNF<)1@ I-MDJ%G";Q"= SK.O$3
PPAII+"[.1T&.&-4$26,4G##N32'$3_'PII=[S*;IW3,4FS4^*=#.WW+JQD G_J:Y
P+SZRV#UBFH-R;%L%]545@^>)(A3E-+/K;]J@S_M"X! F+<XR??N=I'0694.S_8#Q
P\E,/J 4CEL: ?%\4X^F@)[R13@3Z24Z24F(2EY-,3-%+!E>5I<%8H#F#*^$(@[_L
PB,Q%6U.PYEA$6:,!;_;8VO:OOWP2"4H#":=Y5K8YT\=8R KU*"$=_7^BU\,6NK7>
PBT>(*B;H?5(L=#Q)I_/H;[[@,TNKQV!6,91=S<9CX)]!WWGD49FR4G $?8M LE)]
PHW](I2<5K:D+)6I7*"PS?#^'L79@<#&:6:SXU!LYM2#FN48VT*$^KJ1@VPMHLG/9
P:-\R0[!8@%LP-R=V\: [_")1GWC[:A\*=H]'VG#M0*I3FQ7^;&GV&K9?[4RZ)MJ0
P9E"Q.INK%$O%84(M0[52970NE00H**2"%J!6.[1.JGEJG^>%TB[HN),84D8^W==0
PGMUE?X_D18]P/%$PL7.\A7!F-\V0-YN:T%E6'K2GN=<.(<<D;;)X 06^KN0\C8H-
PKL^EC:-)42W1/R;-+K5EN[FV66J453^U@=0C#.D?&D4@E_MVT[RW F\X#-5>5?5=
PSD?&J""FZ);9R0OEA+=$TR8^J<N^VO:/N2CJZVF+UJ#HB7$40O*'X]2Z^XV]GVCZ
P4[8F+$3N3!^F38[%2\$!/GSG:D)LS7C(IV^'=?.G&OK<(R[Y:FYQ]H1[JC!%G$ *
PLFF:7VF ;;- )XM*QCW)^X0.6YHW2\=0)'1J9A;'FK5OU"R\@7C0?]<;R%=M+5)W
P-OAH!4]OF87Z$F3@O)]HOA*L#5(-CZ+P^@\,=.^2:TWIO_M=<93]O^#[TTAIA]HD
P9!#XA%*6#0:4W+@Y MQ=E^5/"BA]>BERWQ@[:'-Q4G^O%$@+60^3VZ^&K\"KO]]I
P&-9[>TYJQW0,M#0%Z^PQL[% OU9;8^@#B8>A\OE\?[-D-R^Q;X97 9F;Q7"_:W**
P=AN-2_N^O"PG'3X_AEGG(;B*&RL>ZG:7J5O@W2**)/Y0[9SK36>#/]+7I<E#)8/J
P-I@)ATZ":[K\&O3D"^'#?U;Z=KON8*OI&^L9;4L@G_!Y 0[J(09B*1Y$ZINXN165
PMT>7&,_JB.W'A)*&RU/\&"R;EU'X4#+D/*ANOT"HS^H3OU9$0Q083L=.]"0:H#H)
PWZ[VYIVX&BH"KU[TQRTQK[>N.Z#IQYG8MC[0SK[C(LP29G*?JO+^X:)S^V[@BH?J
P=A1]ZZW9[XAIOZK6HN)V#P)^A3$O<-BI=('^J$S5G),7(Y9HJ30FE&YM45T4V^("
PKTCU\*_)D.$'2?"L"#1YW$ YV.=XX\!*[GPMJ):W;7YY='SMF7N9U-\3]6KE?UVD
P=*<SYVJW.D(31-ER[H6OG0#?; BNR,C_+96[Z;F%V](8TUFEOSDN<"5+O?$$$/2;
P,A;"[,ASE9[M<@90K[UW9[OT=35D4K*+"ZC-6_X05Z_NR']8@$JPXUCL"NT%JM&,
P2,<FLB#</!ISBI1U2,@:Z+3(/KN\[ !50\=&_"+5LXCL.-_T#O11C11U&1.99UX&
P8C\HVWG68-IT*%6VX:<$N_G32WDKY5D*_&3ISGD6(N^037#-;I&FP^V4A%A.29!+
PXH-5W"2Y4 +K$TM'12<CED\Z:C42Q;PD3I.K: 3$F?\">A">(Z5L9!0 S![EJM\.
P76QIE!D,+Z"Y=J9WLF@K>OE1V!0BEGQ!6PI0*Q>)GT\"LR/'<<ZIIY_HE5IY/W"4
P7J3B=J(YR5CU+8E) I::SLS['(RR)8@,>B/;-1%>.4K70IXP:@!J3H]I_Y6C\<X$
PEU]T*E']C+YKT?W3]KC;ONF[3'5Z+B5],7#29SP=-L+G"AP+E8(/WV731AC_!!TX
P;\Z.ST#?9<]S%52Y2GYX(PGHT]**-#Q(>,R$W;] **44?391EL=EQQ-N^V9!,R^8
P%V ^O5\FLX7SW3PMO>5=[V6F6UONQWCP&H;?U6/=FX5(??K82]\<UXOQ.(07)+H:
P+4;GX/1X!- PT^5(#M5K'&-C+SG[>-6 ?$L_;RU!\[_S&V>J2B0^?.2\\+>2BQNH
P.L-VH(V-0J)K;EK+27__5#BA\ 8D:%3N@'E"VT[*55%?7,SY/B1(B-_H,!5DHZ&?
PK;#QLX<$[\*[%+4<Y)4;F#9"!HP?1(,.5NU5PY5V.JO,(F! GTDJX8Z"\(O\\*9'
PWB[8&/HXK"5KWX#.\3PI[O70$EGT52,!:OA +M>'L3MH\XEUJ;J\#7X0&S'"9']'
P/ECY^@=&O^&Y( 70R[,H:;A$]K*AB6=:X(K)-Z.;+_0T",11H ?4B_*1;SX32+OC
P0>?=]<,]-+24)W++94,&55KD&K:NX[D\"X!40HHH)F*J,5A7#)E1PD&K7/Q%4FB[
PQ[4$,Z]VU]]:M\2L>%,[VK>H*Y:"<U)'D^%\+"="&<9]U'RBLV*I"/*]=;3TCL$S
PC5QWF*-:CK.L,$%^'Y2<_GSNNP*D"BGHC6%G;AY;N4,:-V\WM)<$XK918.<@HPUF
P863\8XB/OAGI.M1F@W6K-(H90U*F+!%:T*[!FN (XXKSQ3L$OBPP8*MTO>5M9E6Y
P>DT(G!#5VJC<QB1_AX0VS5I6FA+$8?AU(,8-UNDXX]&- .GQ*ML3'_O68*L_<3O 
P$K*,*C'Y.=TZF\]NPX#=L@;$22W^P4NZT57ODFE2^>EOBER2D_'TSHH0&>MZ(=5Q
PF# "S??S'RY$TQCJ8NW0-)%T4$&E)]BA4.='[CNV$C U8#:Q3]3=6+B%%V8I^@7U
PT W=?(HF3;^'3B\,;L-G3>,0N3<^DZTQ^ESN;83D%)&Z'+K@4Q?BQ3BP=Y14!4$H
P9+'[76"Z@'DP5]K7DXLY"D0[3Q\BL#/JR0@GC=-U!QZ5RX'8YGXF1<Q,R4T@L S,
P>0$@@?\-7YY8&@&%Q:X8PK^Q=](&AE"+"M< (9;-!H*&;L?#G;MT^5!TC1>#G0*W
P^TYFSFB$ S,(*?-E/7SE<@\Y.C=HD7F,R"5AD4. $4#"R]V9V<0G:V)HU];KS.Z?
P[.Z$K>8']_2]T>#Q%OGE,PA!\^O:>Q?0_B1"G?(5<KQ^W;1H> ^<\/:\SRBF1)W&
P8OL4^Q=V4-H051#/7CCX_YQ"[#>5LY!V 9E0R"[]XZEGZO2( X#4W\M@YJ=AN*2M
PIZ49F!(-H$=_%)QQE0WR(063P<JGND!3:6PN68C]S?FN$8O %R_^5E<$&L[0.^H%
P1>B"<HRTP<!UVJ^]@!XA<HES U#X%LLE("L*7DM[=33QB;!B]HX%C$&5Y!D1!>[W
P2["'73-[M31,M.G"<H*!/OQICUFO[&RES"@N?,9=Z?>$Z-O=*P98'Z]$&!G@(!^Q
P8M*K'EFZ>A1\&:7R>) G)VM2<%]9>$;>]D1_UY?XDY;OPR3.G6I $!]A:/"^T ">
POFM%/'FA7-3Q'[F#$^2 ;9X%:1JN$+(X&FWW)NVBH+1(T17J[+9ISRS0'(I*O+1 
P=N]B*6%%"D<HW(R=K-LAFGMO.%>4I:9+N^WE[R84@[I3:\(@,.UBS+0VR+ITU):&
P@2^8->Q=;:NIHF>4?='6-J5_:B7*O7,)AQ0J6&NX6J<'S4">%D].]E5#-<Z\J$>-
PKH+M"3*Z1*,;L_J.' T["X[9U[VP)0"L3O+#S%D0$VUH&;O&(?&FVRDKARJY%?1\
P,(H%IWZ^%]&]9D%JPN_MTAHOJPD]Y[J+]0XCGX (H:FT/W+D=7A<>LSN2D!^&E!"
P44U__N^5*;IX"*YO4&R)M*N4S+9-XE;ZJZ2#B 'J$[U DK!!)^Y""9OL'*\6$VNP
PJ9_+@K58-8IDQ?4L>=U;26@P*9U3UB;.L+5'\W\A.HF$6;&)^9],8S;O"?OB((:*
P:MM3^4'*GK9O)VJQB",!(;($.U ;+L.3:=88(#2)%H<$\.H%[3)9"IS*#%?B2?U+
PSJ[0&LOBCM\.@"SG**Q!T9UKD[%U/L>\)30QNE?I3"K.T=^6Y9RK>:ON5$AKF@&0
P_QW>5  8[%!(K4/YXQ]#6K><OI&4H5U(.AJ.E?58:YY6!+^UO/ "KZ#9>(*I[3[,
PJ/P68=S*NTK/F$YA> %]U:+<!?9]#6S*;@2E!CSTR?1L_J[E1/G(<\)>Q,L6 \KM
P%/H*4._(QYEPP"98*$@[5> B*#VS%W3L<<MDBR8@1/B1&#YW72)P]U:.$#J6(J#5
P9Z2J4@_7G<M%V Z<\7:+0.?%$-]ZCEM'4CU?=3572;ON(?U.@'O\H'C.F-+72RUH
PU4G%_:6LD%Q\^L:*)??3NB7\243B#<"8VTB+@V.P(_%Q()B>LWOC<\_Y##("*S,;
PKTS2:OB:7;>PK_H;N1!@/FF7ES(';E5M@(@#26(\?N1-;FS.+DT?\)NF&J0#'\\Y
PI$(4Q;#%1C$+WK69#T7W-S/:]1CIU&3ZZ!>;YWR5)I5@0U8+=U-8-G$E$O<7)V;7
P:+>S=[.B72ZKJQ7*?6/B@*C$.;Y=D6&RB*K0U! >H<0,;CZM.:"= 2_NG-1Q^JS'
PU"HRV::V\8[FZ$-R#;@Q^PV^98D:1'2#X&Y?VK["'\^U"H1I6 MI4&'JNH"C.+!W
PA7W-[=/&Q" <S("QQ;#SJ_@(W;5L1ARO?;<-\FH"G]PF'!E^IWC,LA&;\&&QD5-%
PEQ /FFPFP%J_RUA3*!]@MD=$;=BJ6NWIA@JX_>MTIO"1@$3\#=HH9]>D-3A3N8L8
P>B2E6@#BL"3PR(I2G2O?6>6D,&F%3>"J0Y;\ZN=O_EV/<_JY9@9N()1U?YT-V])T
PL+(S^8\N"K,>(@O?]XT"2F&R5Y2Y>)@ /S-STF!V&_;?@;VE_VY2#N<#OX_ HR1G
P#(M>*EDA_LY ]#NP^HD\ICXDN&/[O0P?/'5*ETYOQN"HY<"HD?*^M2;+-G;=.&IR
P/X1C8FOQ3JIUD-H#/?]#F1UH3Q6WIQA-6&183]F83+YMPJ<*Y(=H#F_N6>3)_4^U
P.OYVABN$'X\(O>LXI_=_QL&* V?;L"Z>M:=[YUW8:\Z/2A9S22),4Z;NDS4T,C+[
PTJ6I<?'F&'#T(JXJG-/AI/N?B:CYU:]G# "(\>7 M((PZ2D@W6CC@-5U Y^(P'(P
PD-1#I[_2^6>P5Q>7C!O*H+YXRT'K@2;6YF')9(N%_];LQXQEP+O6W+1B6IUVTGV@
PH%7;N8?^+]XU\<NS7THUZQTQ9CRK'['SH$5?C^3Q[RU!A\+]Y&$J#^HNT]Q+,WPX
P9-U+D:0W!PX:6/1X>]6I<&8NA*A:7) @F:SV,574RJ+D:ZR63*D"T-:T0]O"^OJ2
P,XKFE0#/2MB!Y!32IRO%@WG?=^@K1 A;LYZUFS8S2OJ6WZPEK?:O@\H*:)EBS:-,
PGA!<=@AH+O!*9+)XM)B)\/^XV6H7VL]5PO=PX2I0AXEMX*BAVYACV5@@OY60H'#*
P2LA5)LF^.P85+ Q2-CD08 %JR(&4P'YBYZQV*7XYWXKG38CWS>$C)OEE->QM;S[!
PA^)JLZ([U#O/]2WZNY3J\1+H) E/\.(@4IQ8<AZ50']R!F+=+C&KY63=OVTSQ&M?
P/?K(^1I%MC@>-QFHML:+S9T[H#VGQN%@!!4A+0Y3G.?=MLP(Q8_Y*ICR"E.>JX_Q
PS6H?_[L;16.A%.OLYX3?>O!-U*-_^/+W\R0_X?1D.RA[G/L] R>I40^">EOK[:;;
P8&$=]LL_BY.OCSC^3-IL?B^@GK U>+Z28\+W_Q9<CML -4 W,2)--LGVDC/,VQ"W
P\*][R!L9_#WW!<M)Z$W_$6'$K/U\AW:+ DXNM?/<&=??KRK,DNAXTM"M^$27ZNZA
PJVT\1,XDJ:G4666;>O@]]M](N=2)+[JF<I.0Z%2>M@4,42Q4$T_\[,JTLI7J,Q@%
PWI0Z6I) 3P4 $"4()W1\[;TH/ C:[A'%G[<*M\_87_-\\BT1O:^-CB[!F"\FBH-D
PR2107LH[HP',R64:_]@'X]62WH;+S,)=77\;LH-1)[A&W?G7RYOIC\\OMY@CS= 3
PZ:6_[&/7[KC[^<W"S15 @%<Q5DS&8][%I;2!L3QGY@GG$5-%+FFN3J[U#88&GX:O
P'^MRG(MRTC4"_E\.DRY4\#@)Q4>JJ@H'2LX6D!VP]H;UQ\#7:R+T523U*G90%9RE
P\,$L?\VV]=^UV^9S?ZAUY7TON @+<]H9QBA=DKXC !SK&?T*6^\L_2,"-@IBZT@3
P\=]G8H:M8AAZ=;229SCJU.^C])\8&)9URT145(/-6+N?2VDQXTS9X0]T  9@I,'H
P.L]Z#,0<3U<?\OLV-CY(0QX7CH[A)A-0&#! (0RI9U\*X2>2NNJD[TR\X.W-*DZ.
P2**6Z)R)>'=12EN?UY*/R:#(&1-.C40AG90C.X)/GRNA]QF[81/X/2U$+)H&3Z^P
P"+V4'EAPC: ;-[Y*2O6T 4JU0S@:T.$:Z@LU)5Z5C5K8=W.;% P<(Q7Q/.'=U9Z[
PCSSGKE:76XG6 ]ML/Y!&_:*0<1%E."2935<?O:VY=F9 !)TM!%O_",S>G4T@7D1#
PS9"#KRR^@[WG@9:X"@,PY=>.MJ<NFJ/U@?/#N.OXCK53:I7W]XT3@.;68-KI1B-3
P;:FV\$,'!OY>C$YF1*Y(_G1^;L> 5N 2TYH&UVHK'[O9^K)X*T[8J#(7F1WWXE*M
P !7X_!,'&-BUP+0#KAW'HHM]FEV451PP%E6GXKS!)F5B&)MC%+)W:^X/$<$]+4VA
PK2A0C&@]I&R62;D&BQZ)NQ[$4YC). 5R4GQ4S%GA[63+:6UE @L6D)KOT0&QA*=)
PJK&Q*+!YTL7V6U-W$KMS8F^I>Q!2X$QT%#YQPX,9Q0 %7QP;H )EN!K1S+ZB_JG[
P22:%^?!+C4.5]QHK( A64-2DK*J$/WHJ718[Z38B/&4_P;%85HX^R/ZO-RRL"SPL
P$J5(Y\U2'-Y;IGFY8?VB'IO:Q&.@ R]U'"=!F^CL+QV3HK!:KJ]R_NO\D;B^#EC%
P2R6?N%N^Z[3&G-6:0T*?1<] !2VFK=01*YJ#%,US:=TB(@77'U<2R@B!I8$N$5"\
P8@X9B1)"BQXH"K[Y)=5.K? W/80<[K4M8IM#)7FL#@U.9<AB,F!'GXN""9P59S>8
P=P?GL?>X&FG#H$$U[7D2U ;%P2!R2D%]VD(?'&0)CMFK);;+HK=O^/+WEDQ"DF$M
P\I,\G1%43U<!/KQ"4':U_[PD,^5+!%,R1>F*?+ UU:R<(<\2S&FUEC,VO9OH*'>7
PXI$.75 SYFC=RG#LR$XW?.H(&GN(-0XJ74QPNN$$<=H_)7GG=%(?5HI20@*4Q*)$
PUXCANL7*&MGKJ'D<.3ZQ@RE!4]TIRE=2U1BEKP=S9E3K7.VB-=FJ5M ^-:7*2NYW
P$N&3F%M!VA?FVA[444U(3?ANAV8/MHOB@3"O?,-O;E38>/5D"%KVR"F2>BA4A(.%
P5,E%_&6% R)(EG^-[S,M45$6:JZGBQ#DLORGB<MGKR?6?@!JCQ^2(56FK+O+$G%C
P&<.@-S*NI4R$F@1 XU_Q**0BQDLYOYRZ%8K35W_QH8Z VR]\>8@>CHS^UJU1D9 U
P8LOO#T'VAX*51VL1KCVS]1@R3@CXUD;$1>S.$9^>U?Q4@700GI<8SYT0PB/WS_BY
P#1T2@"A?Y ?_CWU&C/;,C(GW..$*A#^LYDU@2%9V CJR4/TR$7H)@V,SM4Q[YID^
P5LH(><KH<HD/?KE^_@]L':B+!AA;WVC#=P B1U@3?L^!*7>VU&GV )B8P/F]-MY^
P.-F1%0UEI2H E397.(:ZK_6^4+VO(R=U,]MF7D\"*5&W\Y2A(#),.L[H%&YX,.)*
P0T-&LF>K#1$/V*,HU%V(+S^B2HH@+EEHM"N^+)W#6UP0+D%9A,TC]MBCIJ2BDWV\
PC'1K(# G':167\2#K*L?B]N"!"\X*\U?*%7AD@LC([)BI$@[!^T!XC% DB(\M?#Q
P^Z0E/I8;#&9^ E6]X=.550"FU$F6 #]P0MI:S&VV]6"$7YQ O&WLHS[D[R+E/UKO
P3%>TWI?^;S!,+SF.@T?%V/SO9$QD0_W7<@YB+B/Y+ 3.,3Q2%#"M,=))+TR[P<Y+
P*"=B(]F(#&*ZU9'TRA>PGQKD:]H2./O)/O#*K8QN;0DH=MM7+C0J'YC>F!%0R(EF
PSG!&4T=[>C)1GW&UM>V[63VJ\23 #I4J^"ZM722_I4'_6/.<M\F=_)@E%#]6&I[$
P?F2]/?B'7'#2,7!40[9!60MR^3$86F%>PDI(;=AY^R<HO])1]AQ';W^<PN2SCC>6
PAYG!VNHC?CL5Z)[XP6'KY'WQGG@O[<W &T%N<[K8:_D I6'5:S=]*+<BXZE\#2_=
P_G _=/,9-GC(48L3:1.A@&G%6=)2=CY''*^EZI>8#4(9$H]V8<N>%=@_X'8NXL$K
P9J8ZQE$0IXG=@.TNDK%"/*]_U8A^T,TJ,0H.%)ZGC;R.;%DS'ANNAKY>CR#:#H/X
P!H28UPQ5^)X19N =W]D,Y+8A,!B?U"+&5&U>SRL*D'+<G\5B8>Y8K<L)3!Y<N?3K
PBFFC@WK:)CM@X/(,_U6%N[P*^8_($#]1\QN23.8TB4Q>V^%R(%/$XAJ^WZVE#J L
P!],;%.HA)S)/:1_$V]0%7R[QN-'((52OI-GFK<%[-A8KTJ*E B'<*U6C G%[ J\?
PD8T-0I4]4B;$29!M*2H?*W,I+UYP<<2;IO-+QW(50GTXO.0>H_8SDG(I=)&@HSI$
P1IT2EZO8&*"Z_7@R2!O.B0XTUA!_3&"E>O6>?<O>39X'9Z'0$?JS+XVG-Z*W=T1.
P8H[F45DMG- 5E9(ELX]JPYID&1L,.O^$"7"9#['T]MORTGXE[Q.O"UY?3#;'$@'+
PQ5]?-E#E&R?9RQVO2/M+EL'@H2J:3V4H9*'RK36Z?M5H.1%O<$.$?&2+8 >JV)MZ
P$^%Q<.TKNU:'I4JPQ;U<$*36P'XHH HF#R[-HU)F >NX*O9OR$INI>U%;F[")$AL
PENV4R'59+")*/'3J>O*SVQ%I NS3#><K0&R1C=5/XSEF[014[(^.Z@&I6(EY46CU
P@P-")ZYX$:+#-^"&Z6=/.7)9W/)97I)]L+T4(()F >3P-_KL5KT_QOL$YC#0D1[8
P@_KK--"$D,KI %V^:<0SI=G%T<43RY"+;67X>),-FOV^9XB6<\%W!]?_C$:6SZ2[
PPL\G&&9??Y"JR:>9RY3;4$QY]5I*8:_^9F2"*?CQV&U+#W1<1/;XQ9/1A.B)HI N
P?M^,PESV\N>UVOR72#97UI9N?C/;A7\*T-X"MZ@I=K:'RP=:+.7 )4(SKG!X5;8/
P8[X1@%S*(,ZE+(J1@H5^27_:\"P\-+E&Z?^Z[:Q Z,1T/$K2_<ZV]Y##JLVBGA/3
PSC"-;%$8+7:"+*&NP64]YG4PG?J4?V<MM9XMNZ1.I4-3-_ZT?%M)0_5R-##U8N/Y
P:;!CBX5Z!*,,\D+H3_VB&43 T!C$.$9)/KM)FPGTFA4YVU ('V*L60NV0Q2F#8JX
PZPS1G*+3J&%]XS(P_D>:C)\S4LA'EA7NS NV.-?(S]2S;]RF;YUHL&P!=6@I%28A
P1"+_+5"]'6OG"0!L,5+^>]@=DS;_ ^@9-,BE!J-\FC7L 7$]C.@>)L=;*'DQ&_DU
PQ/=?VP!:'-)W76OVKB3FA0.79,U7^.6!@ 0ACYH&_!G;@3[>(W.VP'):9?>IV@Q7
P1[*I:AQ*45]%ZL)_\Q;4ZKTL#W&LODK/.\GVNK-+TLGX07B[PAM<C7<%+>+_[&)W
PTYC1U;1716+&1KY++#YN%%]C7O"E7NDAY,<]G2 283C@4&_LQ&/5(),,+N4>:; _
PDT4.(9OJME@)%MCQ0%O_WTITB>-Y1$8/-[A'3Z-3<^J[OY0R_E15\!%+EU$#L7A$
P)G:Z# ;?^O8!0>TT%Z(ZK/T[5!0329-GY(2+P67!;BYR&!C=A;%"L!DI5G1!F"&&
P4.B8^^B;KQ5/AUR/BCJ2UB_6VD <M.$H?<'P]"\HC;>?T-GY*6&2BIO(15? 5JR:
PYN !KT, 0IL\B(=W%/6+>22_,4$?>#.W/!LL.*Y0NPL.K-B.^,9ZEB.R",'LKR7J
PFKZT$241/DEF_?F__.+0QZ9ZL:K6Y*:'\GBZ@>]6"YNNA<#!KF0B?E+F1N5E9?!:
PRRXUK.(8GT7]Q-=F/[EY:#7-!*_F^;/YC'86ZQM<E=E:!;=-K$\'J)W_:>X@97M3
P7I^1/M73-$,X/ZP_2S:JOA_ TH'RYRXW5MCH'KZJ>VI2&SN!3TMB(]#1U.#>: /\
P+5@"N881.=8C>"C1D7BL[!+J224"MM^2M<:4#;!Z8W<J-;]$]MZX!?VNRYUA *&&
P^2B/T_,+VC24\.E!7R[>'[TA#?2$UVTW8!;JD'9XX7G;4/UE/A39+-TI+226.;^@
P,8BE<7Q]3\\&M8@\D8VO/\7%_B!GQ&3%Z17JC/])^!>&BGU <- D:"]A:699PLRW
PC&K/$MS$:<]Z -XZ;TJ$8,60O"%PS^]*/%I.6(SWQB$/F/H6V3)#9S#A$1RKC/TL
P)W_X16GAI,-A[]V'".P,ZLRD8.#JD\S*;WMC+N<JR*4N7B00H,?J>P$.S9>>0*:*
PNB%%W/Z)@ SN%>:<^/@I:\I'=X;%,B'BQEK7;5W[JC-RG@!T^0V/U(HO'6R9V;^P
P.&6Y&RD*943;,0^!E"O\+!@.]) ;6T5X#AW@1<_X)?C),_ZUIH1EGQML)4@6"_2X
P6OG5'T33O6Z.YA3- ^SYZ&9%2@YA>\]^K*JI2:?*(_O_91_+KX+DUNVCS95)_*+7
PRU+)\=W:8_,LZ["H,E!DW+AK^K0H#<!'R X)"4OG$)\^''5MW7TLG$0?%Y\1HF^6
PLK/T'_MXV!@M]I':QMJ'T_VNI\:K9EH4WA7ZO$(Y6- M'3 3]IT*75:3%SYEA'+!
P[976G%;_.Y*C>EVL1=,4=MK)PL."EB*2M?(HMW&@E0]S8V:U&L<G7@&B0@$\5JU:
P=O?M,#JE]:2)89K$^:"'Z*\+*P7@WCTB%7I_]C"5.W,'WE'SV!+C%MM$??@N#8@?
P MG$BCU1C9-:O?TZ<^7O4^!NKY/<L'!*489L*PI:@IAJ4,N\LH!<!#4-ANM?/99)
PHX2P3ZC0,:?XVFL@ '*.7&_(%K9DH;R^)PH03RO$ H!2,1L##8O0-]USG>M ?+2T
PRSF7W_'PHPS;$?'"X&BPG>M,Q=G/'I:\0 6CELT8-1U4YJ/I\\5O"\(9;%U+A/FJ
P<!@(M)HGUJ9[E] _+]_(0K5&WGNIW%G>W:=CLC'3[P"BP+.1@L%&.8]GV3'_U$LR
PI:;T]3WK?=30'T#*.=E049CPV/IVQ?C6T300VVI@\@F>%\,3Q8ZU:T:*I)SR629Y
PO5;^(BGI]Z2[=144Y?:A%!&%T1K4Q@(B1V?:J)GRI_6;-AKT.M+WIZ==61QESUF]
P$LV.$%>M(+"NGN2P/J;F.R32PQW6BC(CXJN2C'2+5;+R48P4%G*V_ A51L__H374
P.6H/^ZB>^B/I9-]<6UY3PIVJ 7,^8"1TEX^SF[D3QAZ>\6VT44-K\=K?)D@P',)6
PC /P.8:/ XW:5N!+:NS)+9G\P90T?V3%!3%X8.(W/.D(Z7 CN8(M&/J3%"GR/;L"
PA!W!SFH@9=8\WJ-;-I,;C9J"D G*^\O<4T.N/[Y F)170CH&H2U_ F  .68B8K3?
P@ERVG"<$MF]L-R/V/>/B:#&CF#78 P!]ZE#X,-7MO_%1RRD/>J?@E1>9@@QX JYS
P*FF.3ZCZH)9U&.O7PXY\1YJB=6.+@38U1KD+?\V/Y+:(E B>>/M'6CU!4S&C&AWR
P3(C$.@G\[TNLXUSE\J;9Q]08F;$*]C/4R'7U;C2-4(/ *4+"62H;RP.'^CG_0R62
PT 6IE(511MTB9=49\B&76[?Y$,@Q++^N'+RC1=(QL,P51=;\BFV_F%X/9<%Z92\A
P*U/S91I_!15Z1._%J@8">Y>:P-)Z DR:+Q[789Y0P5/J,VUU< H.\.RX9 ? ZOV8
PM:=[.61];9\K!Q!N'*_0WKFMC:%QN&O^2!2:Z.OCLWW"LLOTF@I!3UQW\"7>*D#'
P:W4M!!DKMH$L5PKVA\M$UAIHAVP:1>Z%O# 4H4^-;<]O9F;&6Y8+^$6::S!>A!+W
P)A4V:9^#+6%'XJE##D@GK:-]7/H 3HC5>RPQ;%CCQ9Z5L'&)SO"C%ER_\+L%DGVC
P&1?*VOT6[_^E9<0 2SV/<:SDSNF7>7'*!C-'N_7! 7N<T8S)NA9BV=<N3$_<9PI$
P*/XD,^B2%8\G9REHTF]&14B#ML5\8OR\,V&$/5'J-?R^(0#NY3'3Y_U/3J'RH.I7
PSUJDP)0XE!P\B[V*X%1S:\NZ%ZX -V,Z$[\12>6"_.1RT+*US$%&51G 6#!R"W^@
P4TJ+*"]/3 B*;1ZE,<+6Y<DIT&8"BBGENXXP=__+L8E-41%ZA R.-]5_J@?8",5A
P+\OBP3ATM'7R!S_O3%FEFE9[7&7Q3 W3^)T[4/ B\@8YDTR_\G#-%Q^&:!3,JW&>
P$@%?VE]<J0Z:E]&)H;BQ8T5^DMZ\N<^Z$*MC&6"A[XTG=X$\<9V7V++.:_2';*L5
PXC\S="8)B2,U05UMP"=\QS7._.O(N 6<_1^V(>$?(=3:8][Z'N,N3<N%SP(VW[]I
P]=M[&YW!^C!S95Y9<WV]':&V+2LHO$]E=*9,;L8X":ISH&^?A3XB?Q*U)C6+N.5H
P*8(>/[;C*0R+=#/C3!CR#C^*S",KO1!T39R8^K)RHRF+19I__N>@$+]OMX?/21'*
PK450^:L&)@89>)O.?TV[O1.:09J&!@O84X,*V8QD<A@J7)ML*-+/][,L_W%'YRUR
P4:H[4LGC/ I:G=80Y!#NK['7W_C,PAM,R!\*\=Q_;''_Y_L%HZ"U?O&75BOH+R1J
PBR"6'?_.F0;#SY[6<K0+'=/8EFYZ5&>Y?#,Z:)-6L84N% BH-K>5)NKTQ-#R@F.T
PF!*'KK?'5;]H>Q#G8AHTM@(7N_:+&KBE]T.C2C!A(@X30,_\]@(G\K+A1-6GD9(W
P;2;B4_L3"8=$.+F, 1*;:*5N[Q5@J1"Y!V/F0+90(GY,QYQ3,3\H]QD8FCB?S>'<
PN$:DEY1'M7WG&'DW]Y?]']W:5C0SKWW<:.;UDQX01WHHC@37D5]:Q;ODP?P&A,X0
P<4%5SM&.Z('J^7",)'8>9,YQJW_*#BJ=TGBJA^/:QV)B].M^3GB.?T#P!XW.9"*M
P-;/CY"'0\@U&#B0K^EI@+U'.2[1:EV/ B_^VL4'XAYN_31TS8B/W1B(4G-#D]'9"
PEQH;K?ZK7-[EE_(=] 7_E#/>O+O@G^V3VHH/5<NTU>P]XY>M- "S7YJ;!;TAXI64
P//BTX&>?JM,R1%4>(>"\V/SZ[/:B7Y\''RT\"4&%/A"'&O>=GAJ%0:R3>);T\<$$
P-LG6TC&+;XE2C4+.'G-3G$\L_2/V*J1+Y[=?96=Z.M[-J(+HTPJ8RU_F80^C2%OP
P1UGWJYN-O[# 0:Z"[NR<YH&!&X#S03V-A[Q&+?*R.BU_E4;>K1_)RA50$5NZO*MV
P ]CEU[NP#.1I;32=4WM8NFK#P3H#I5L4&EJ7_*;2]_>MKW32=-T6987Y><:OM<9V
PL&..L,Q%J:",C=\/1>TU).C> 6]")'904?]H:KQNK?0\*^Z,IHL'OFH@5K'4!_./
P&T&W8I1";9]GB8'CU'0<4-/+70DG9N@;A6^J-B%(M/DS)?!EKGK++CN8:, >/<K3
PS$,ES"A*<M!JJ)E4WZZ#"6! U;.RU8I&\+(A- *\)G[0[G)OR\V1]YI[#!F5(A_9
P1;1$$M0 U57R\D0:R%/XDBK1RN]XO0<<Q4@K#0P:LDC] ![?2';J*JFQ^S:PEW #
P0Z9E&S$PN<BHND^>LG,J"#G(RIVE,\VZ>GFZB_N4ZV4^94!FVAQS/;.HL]CFUY59
P!"+4TG;!S^U^>Q83A(<!<#+W_/;4#T,E4 =GFDTF%!@3?T5"[V,7+[#NZ9@_XN13
PS_F^\T927?*2@2U@(@(:SBL3 _K>%N2UAOB1IU04846WA$//G 3._?& V0X%H#ZF
PR$5>C/:NJ+Z"DN$T9)WASHT,!E6D4OV*-; )-H3DL73DALS6 >J.8F%HC&:"7[^;
P9V6Y,664P!9STQKN;J!@6KJI6W6$H%:DA>28]*NK(S-KC9]YTME/0TB[URJ:>457
P59J%0H;?(8[BN\3PR9N%!=RMR]Y>6H#QF",+XQLR7Q04'L,&7\1P0HPX80WKJL:W
PQIZKUL&Q-,P##,8ES.X;W+$YUB-2]\--@2,7\=%<4>>1H0PYEXV$0@!30ELJ+H3.
PNR\@5]SN53:6.T?Y0*C*EUK-]F#YA,$G!2+Q"9P].0X#"/']%[)>XIF^+/W\;!-"
P2'"7DUD1S0\/*L5C^EJ2%'^HD;).:=@,$C^\9JM-]P5]<XTU<11TX-3.!(J4M*1>
P&I;FURKY_25XT(:GY%Q55W=:34S40.,0GPQ=Q0K!"?$MXWD2(V)U(G9'Z-;661S#
P8"* ^E"=NM:^@RX:U!@FG"2N(M=/ V9]D&ZM0S&AG$@=]FQQX+/%*G%/U;<^J&G-
P]M;\Q_OB?W])5@S*JY@@MT[VR8E?[LCV D+E\QNZ5,AO?CD/RH#&@^2*:,4]+FE<
P(5VA3B;V.<",CS12T#2Y^/$'*6P#OH7$_[B/(+[5RW14@\_[%R-9O2)91;EJU'+-
P%W-:%.9,Q'<SZ0P3]L!BLWYG13%;GA<#/R+PC9](13TTZP"%%/X[QYH!!%S>OR^!
P0AO0EEE2HM'[-B ?=Y*W1UZL[@M/[C!+$E<,3B75F-=/PF?<B@*%3H<X@X,&N(PI
PVZD)P.VYC8;DUF)V*$?&*"-E_A)Z8@]=V\X1#B\B=W('>,A_!<:2]ZP! 3>A(? .
PQ+^A9,>I0)%XM*FXF4S GM5%6SJE)<S'V)WC>;B7DJ&O+ 2Q/ $@7[ 6F$E:K'"8
PZ/<]<JKKE$C,XJ@3L_DB$_=UUT#U=>8-$*"V7*:(IA%XSI/WHMW:#?1Y87+2:7D1
PBL2PKGIQ*1AH"5^W9FM69 ="PO8R,F7[==D\F*9 -Q]'/^]'1PRQJ+6A$UZ$8^\G
PXPD#P9[)RF"1CHBT^R</@"7>9D/U.C$&9@FZ,L8$I'QD/U:W<UE]/,>LB*#!9*M-
P_)!7%\;D@^$=>DR[RD=*E"!( +NF,_N',^(G70RDL@D_PK"HKV>M-_EF5IGJ/>/B
P4NPM@@(0X7USB?\J<;D172<3VPXPW %#QP[WRW!MQA^=>.&B.CSOXB1:OJ[4/W/%
PRLVDKK!6R<(VZTCAF[8U;\H*<M('9,S^-\J);"6@23P HJVM%<\')DQAOX7<S(=L
PD\\O^?NA@ETT.!;7GAIFPV?F1$9&R9,H"5>HV7<%AOPWC5B;GBLGDPDU0&92.H)&
P QUGSQ?&F2\(ZG7E=M,A$JW-NYYAD3_7O?ZI@>WO"E$@D/"S+/GO$M9.4W:#J\A7
P]N?[M$/XXVM+_.KIT>%"ZBLA#D5,+/F=L[,<KO]2PQ@"+E(US_"(I3$1<SJ'.9^C
P)P\ZD*X"_"=4_OPU_AS@#^P@^'( "Q/2/3>GWW8T]PR^.-[@K/Z:;Y] P1 T #FL
PTZ*LN%;QBMY/SK&M6:C//(JHN&JC>S\),$%J<$M\)Q/>D+-L!EHVN3!G,E2^<+#Y
PECN!-&$:!_@@K=W]H*3F_U*-&T0FK.T((QGJVZ7_[3PU=IVPLPO.^H6$TA?D\?U$
P"YN25GYM$J'W(_9@WC8S.^G;S)C@%92C]YS1_Z"_6YQ"I-,6M9JPB*&ZN@K;$P8=
PYY?K\D-T]V\/[^5J*QUY$DOFB+;8CIY!ZH?UH1 &&8WL1UL!S@['3I.6',AJ#TCN
P 5.P[\49\%9U%=ZN'ZK?X]K1/ &G^L_S9#8*\>J[(RQ7Z+V^)DVMMZU"6U>N=?,J
P<?MT)J;9AHR'O1@(#%A)R%26^""D_OUJ%&5851G/G$MSH%J.6)P=]BK^'GJ?8$M/
P)ID(^[;02CSR :G%\Y._&6Y;Q)_M=!GWBM7ZQF2^9<FO=AGS6W,][U82@ZHT]]9%
PRD(Q.;)>24-_3]F*$*#K+V>>(%&]\RV^-4YB4FT@J 8Q@E,D_W("?M(^]:2!W'2"
PR:&-()U;IL;KBF4E<*\L4F?4M><NL""<;-<W4&=(/X-G"=C?A2^VV.::-2=C2#-W
P3B_4>_LJAL/4Y0[?P+ST\9(?Z&_2%>13<VK-Z00&=MR'R&-X?6/;YK:[EBC>TQ"=
PC6%'(]E2HB,Y0<@'KKJ&WGK,_8PINJ&=?!P4'B3/:HON0*P*'Y[0-J/A,^ /D I%
P?6HEKP*;]SS0] G-7?$2<N8$!L@W#T9J,H*YA54GUDP3])$LESG3W\-#L]O>.2#C
PL=-S4ECVCNA_I)^X8XQ?OO\!I+.Z@=J T<I *@-B1*N2B-*^E0'T24:^-[XLDHW'
PUI2[X*_>PG&1&>1/G 92#70@4 1XF5\!V#E1Q.);!C.ANFF!:E]Y6[0>RV-($1Q^
P[;D1F;(@LJZ<0ZJ/=&1/:;Z3V !>FTM2QV6X__RHF%FK"D1[F8),H2CZKG'XVN"R
PK4-,<N:\(QFIH2536N/2KU/;ZO@P<PP%[$2DNF5-G/<J4# NC<:=28L 39'82V)5
PD+B@"X>+UD-X\<"_G%*@6)9M-WZ_T'A&(]SRDONB)*M<T82N;_SX1JD"2.I9N6W(
P!-(Y= "%<8VIRJ-(0Q3H[-DAU[3-57O;/*\#(^1C_B 3"14LP#)='W=>9JE\]!+,
P@@'=QJXR+27>U5F%D6:W\I,A(F7Q.A_3P<N":3OHU(2Y1]I=E%%I9N[^BM[^&[!V
PEG GYNB;B27*\1T=CR[[-%K6Z2IMB$9PFE< XRJ=A;W6X7.66DZ(4:Z^Y-T*HB=6
PLE[=VP64#&O)TR_FDG96RZ(40?Q..M:U*KZ1I\C,V:&52D(B/$/+%JT_2\E'2C[O
PQXTI.U27.1SB1MA>$Z-Z4_KVEYW^!).UN>71OR7W+13PV!_I:*/&["6FI$[$YR^E
PKL <(;8N@J?:/-3R,!NK&*85X^H9,J#1,K%\TAI@^[@_T4Y)K;2 3 L3]+F= P96
P1H!BU]BO@*!/H7%5HB&.REA5C^60C;Z6Z.]G\,K;YVL0^CXR!H\^X-M JQXVN7&J
P(C!5W1V6>ZD@;A_2?M0I;3GY:-D*RF2D])H%G&AFB8?0#N#.,D>H]<"W=UD!SXW?
PN9ZFF>4;?;V#,Q:"V]E($*:.,])^TVAAW9_>NW_A4FIDJJUY_ 0,C$=99"HWA*TI
P>B0@<0*6R@_WVS_)AK$QPR@O"MZ[UL'PX%Y0>4'V^VM^:E:BD5Y;&0L9H"^FCC>C
PQIX&LZ!_QY:3R&@[.?2-?;_EGU'^<QBGHOBUG8M'["(FWD^N('!OQM81,/(6T.*+
P._SD[;%[#<K#$]MMDOG^=B<5C*G2V^/X -I1I^4_T^W.AJBUZ5+E@WSM]S,1H9@:
PI61Y\.77'RTAE;''([H ]8/^"JFKR%2><:F/4!M'+?QO:*VYJY55N'<=]UFO@7P[
P-0(*#MXF=J2_C>6$#.T$5"UB1GR/A1IN,>7"1$\*6D6]AQ@VD*S'GI'NR!#_YU53
P5LC8[+[Y@F>++_1*N,[02T&)$SF%E@\GU1OF=5'[#A2KP:OBP3Q-OBDRR ?([?@O
P8 #18;W\W?49/%W2@V9-HJX.A:?+[S)V*?-8QRDP@#*%\KD_!Z.G=$&=I7&'H_0W
PT@SJU.FU'DJ;\7K<4S0$ )5LC)(L&1?Y[V6Z'%] _XPKP&X>L[G@8$M9W]FY@LRK
P#(D7&J[[W+9HNV+(*[*YJW_I_#>BF5MH#M=F<)7%^_C?N5ZM7I]TQ?(]\^Z/.7FM
P2E//M[$6NHJ9JB4B+B*P\]>C%EAASZ>P^WKT_>#J- >F<TXEXT#!#4ASP2FTW3I#
P:TIK32P?LQ%[@N (^V:8]E4TM!"0@*TJ8U/I4YV940V):[:WF8N$)8,,;^RF]]:R
P<ED96W5$- /A]55O>4DD/,_N=8-]WB+%AG]P1&GH(Q+#Z5,ENLB+J.7K.RZG'1DQ
P0(NK4ADG-E9-@1_3\V7_'CC;1.TK!XX@$=K03.*UK:L6E%LM@D-2ESH>0YD;M-,M
P<3#2AG_\S= ZA9RN<%RNE3>^.(!>2(*&RW<:4H]J!#(4I+]"]_&*;R#3>B,O$)2@
P06$.I,X/DTF!>$[79/6:/==(\2,G $768Z1PN=U'6I>(X3V$RRX:!A\26=8_N!RM
PK/[<\T9QE">KX2::PB4,GKI.4%V]C/?(J+"=!26A;S]9(6&NG6^+-%@>*:FR*.^G
P7U;9AV=''D[8&H?_HDH>&MW$86TL?]$#,!DO,Z 3&S<^)(!NJ[LE%-;PCI: U"9&
PMJ\H0T(]2TT<@^LJJ4ZGI/9D9\XN'$602-]T"!,UV-_6:I%!. PH_P$(]Y, 9VH8
P"/LJ@21X+A.&Y/LXDE,_Q/:O<=TSG!)<]5+*.MV/*+D1_XG/*@UT+LUX)K!0PM?$
PT7>=81-7)TG5!IT%KYGS.2"FMQ++1](_]K?WIRZI=EB7V]3&.(/T3P.G[+W/LF#T
P,Q4MHU@A5W9XJ/<H+5PJL[9+>Q5'K$($B.,KJG?7&P"K3Q'0M6K,')YYM^O.9G.^
P-W$#CJC-,'S_'N8$_\YUJ+8!**XT!LEILWJ4[1:@=[3ILLBG\ ;2UNY9T(S4G!C9
PV9?0Y?'/56*EN$MHLR!7@^OC4=H![?_'-:#'Q5KY]X?C^@1>E(I54=(SI>',,UP 
PF@^T)K0)A])HE%,_4\-%<"A#03D;48RVMCE2;1"$!LK.,.$#09.765M +0PVK]8X
PKJNEWQ'7[K[$-X*7:!@3#*.R9R?K,86]I@Y'8693XLC]VV95 *]'WKA:XL#(RI/_
PC>XAJD4'YJD3H$$QK68X3@C^66:R?%!'9!AH+%)(_3XS.0^%OQG&S0Y1]7?=XLJ>
PA9E8D0TS>(LB\.&>T]G,>FT'+S$X]M0ETEPS%2-^?++7YC#9A]!M/@8O*YHT?H&O
PC-($*&94CNSGA)/)LH?N@D/]!DG\9%?@"8X&WW8+0M9MS4OL#KKG*+TVWE?Q6:0\
P(P=9J+V+?$@DK>(KO<!-SHTPJNF?OD,58+35SGCM&/O6^T0/=5AB6MD(Q<Z::%56
PUZ!#,B)KZ$*#RH^H=NE"@\0*D[/=5^MFEY^KD&1]68B?7^FUL3+Z1J<P#9X,\7WH
PQ91:_M!%V#DB]*_2"=O^_90W]&#Y62H5C[[OO2(7>.5$U40!K9,?X^1Y=;'>67<^
P- EA?OJXOG1GP]C']':I:4,GI"Q7WB^(-814!H7H)LW0/N;.@+04!FK/A]'A<S/H
P9:MC?EOXS[5.B_+(.6;KJ&F:&<P.9>#,[VX-C&'AYYPKEW5Q]5XMGK5>&9R9SE2I
P1X+BQ9T;6J&V;#@>XO$! %;H4.V[PSFNO1.'J=;B*%6S0#(AE1?9@@3#N?HD=?!\
PDE_4(FF)OTVB*J=W_S.W,SO2*Q9$Q<7NI_"Q),(1053:%AT\:HKSZ./-JU4:9?08
PAPM5>N!V- ;'@AIR@RC8@#I9VGK$0Z-Z47[VJXPQ2&U :2X94YI]#L;AWOLBA.+@
PB'X9X/[;7&Y0TK_H6\4+P!B-MMHC'172]"CO:+YG@R#'IEW6T)526KR+Z]Z2$P^9
PC1;)7W2C]NI.5!G[/!!SS*3X/CB4R"2=4VY[B!5D1-"W?0,0VEW\*Q,7]F6PDE?)
P(RX>F0@0H9A^>?!:#4A3%W^ #)"X^UG5=\\@+',Q;>RM?PUWYU]**99E<0GK7*OX
P)E9)T"H*DO]T(9>QML<37.D'!YCNB->6]V20/!65"@OWQ\*=:2=HFFNN\5Q8T@[:
P$BUR+G25D89-;O/HLF5\['M'2X7XCHK-#<*P0E!*6--&[L],-O&MI37!RXBS.@"-
P(2U#[TSDR1<F'_^:MCMR"K5>?$VN7J+8OP9[YH&C@NYCDT7^5]Q*+^>!D$P[*@GC
P'S^5_\):43F\"CLRGM_/9B(U:5/^7J.8H(J!2O:]*'QB:14+Z\,-,,D+0IXY6S.K
P@:PA#/*QO'Q.ZF8 7Q6A"^-20%@+8));>31 ""M#YQYQ>JQA7*^J%,D:<PL!.;U[
P6X;I$5AXFHGGT*$^ F_IZ PT2GHKF[F)FZ2-4. YU$]^N&KLV5HRWXQ:@OK-N0.6
PYCHI]*Q>=8\?KVN:7-<5:CSR*#TWD&.8*SR'CZ^8SE?6=SZY7Z8\<!O[B]:];$WX
PWGLI*6O>;DS^*67CO%?CQAM2NAX;V>NO$LXR3O@$(SGQ;08Y31?**[P>.!&EDH[Z
P34U)03S+YKGYBVCH_J6)N'"UM5Q1A4>DT"IMI5\2@B'SYCF\8NB756_(TXH$:Q<!
P1$(&\F]J*?L@E Y=RS?2T[#;5DM+F$H\9X6?8*CKL *9DBSFC@M#_7XQ^<F]6]S9
P1.'W%X!;5Q@HJA<FY%M+_Z@:K(O?6MKI0.!.".Y5A@8(RS7:O0]+]\F,N.V,"1/\
PSM0W9)M;UV8DK2@F$OE4%]NATT9!6JT%-,J&U^L4@%BB#[N_N'B06^*VM7NQ":%$
P*$>"<XY&H8*TKZEH<@IQ8WA36Z(@-*E9Q=0MN%@==RT8O;:XNVY\K^^42?#:H&,>
PI7:W\7_^'W1+#D?$ 5OCS7K%7$N"T''#R>W/R69%G$8<I</SAI0CZ@77XTUD]M2B
PS=,!BP2#!C.HQ5N ]A1%%74O<>='4ZR>4Q/*3>GOE 2QS54>*[]!\2P1 ;3B-&RD
PF/[<I5U>F\?3K6*AM9BJ!R%X._8"L)VIPZD^P28T41>.DB1 2(W:RTN4+*76K%@@
P&9SSU9R<,>?,66B:FAR&A0V*"HXQ_%6.#7&;E8<P73\LVK6'K/#RH<<C0%S/64'$
P/T# $=11'+XGS(TTNHC7LF8I(M&"S+21QU+Y=QC#B\..%]\]*Y;L</'&1P;8+XU 
PH5XOEA@H Z"+S6I8R(H#,S7E$X+S3(F;'K1'ZS.9QYDZ\AX)K"$%-FW\IMTG N9!
P9O#&Q1J'A:] >SI:4TD0]54[, N)HBUP6Y$97[_%-]F2U1WU+TV[4Z@5U[CNI-:[
P2>?36'<&GK7!;W U=['F*D?O7RPL+B/^J2+RJV8#.^#(N;8[M!I+*FA-O[5] H<=
PO T5Y?9[\S\HJQD,KC<C1DTW,=W8E$\^0DFM@S>H) ?5> ,6Y9L>)9$EU=)-OC[0
P$Z%&!')<=_H/X%FM-QZN)C6]"+JT+5[@2(2=PZ<R(4=93,7)J>#'_?;#D=Q2)GSG
P%HJ,+>1D:$1[R-X6B^$8]^=JFR!6/P#_$QG"73.$RC9[BYY" U2*(@=_H2_E^2MK
PUIS.#(II8*FN%?&-P02&G AFN8%F3,R8Q+V4_7,C"N6@J<$JSI!/FJQ [F+;S*T]
P)_;$Y#2934#>=_L=5Q/ O6C7_=-]*:_/M0^+2U<).!^ZO$4\\OD[:"BE>%!_&-]>
PW@'<CP/BGH[1B,T5RD6_5?@YT)U1"O -1GG(BWVK-H6REKK:HR\QHI=$F.A+[P#G
PG8<]H3/$E!-E5O]NZ6_3M&R#L;;D>^T04;_0DN!OU/E$O>R/&CA?N3ZC'JI4Z%"^
P]\DESUHI3I0J: ;GNR6<'3Y'^)/K^<7JL>$#MF0/I6#3;[-CM7*IE>'Z>T$0)[.1
P=DK1]QU0;_Z=&]'-*E&!P:R1!6YG$$K_' D*/)67(5VUL""1ID^Y.+L_/OK]:=Y.
P&VHQ'V=ME PT(_=Z(;D#IV<G3LZ>\.@<("PE54"\/J;'"MD5H,'0*6"/T$F<RN;>
PHB(7?J>JBYCB\K2D>212IUXML;+J&X3IN&BB^(=/C32W0@'AG;YAZU$G: )(:Z?W
PA8^QZX6'.$S'R8XD4+R- <A6//2^@,7PA+.:OX?:>I1.D<;95H9MHQH+4D*;*33*
P6B?!<FR3Y=@=@Z3P=+-? -[@="+]4U (+N(W&6,\%U*\$)-63=K5L#6/NSRE:6YR
P'+^VSFXW'FOS7\80N"/L&J2<1YZY\\4*HGRD\/GY>'XY!+B]7:C"6E5:'R%N]F>;
PA&1*_[\]?_J.ZO+;;+D+@'[G2V&5FBRK5DJZM:SR0@J>J*3RK0L6=<=V%[7<42%%
P[RHJ&RDT#4GKJPU6V@;G9[NJ2F-QX\TK=Z-L]QXL/R((@9:N4NI3\!"H<BI%^H>P
P7D)(E8<)93RYV_/:^^G'+:MC+I2T.A_J9@J;'9HKC&BD6O#+!.+RTP=]T]^^F(XT
P]@[0NB'C,9WYOVT!WO8GY[[II::D_/M*9LV>C3+!'1L,29)H$75Z&26=&],LG^"7
P)K.5?L!4B*@,G/D%20*K_T)RRH73YPDT9R8<GD11J[UM&9P\C+3,%%%F])UKG6<8
PD.O\V@QF7_#2!6\Z4KZ3C2Q^%YSM/) 9;H'1$#NP/["S?>;ZL8+ -2/S"T\B,L1?
P/Z'HL98JYC_O0ZOS!^#@7Z$7;@EE]BP:M#[5O2+G)I5U(WSG&71NL0+3OR$A(^8C
P)D&@&\_[-)M85L):=2^_Z.F3UGLXTQS@&EBV8M@?BC4$RBR3=J0//?I4Q *^V6'A
P+;C7 S42KAS-A*F2.[PZ@L4#MFUT<%0#ME3@T--;2CV#(%2^:E!!>6'0N1Q.S351
PD"&WN3AVJGM!FE!X6)2P#B5IPR:U3D9O+X?(Z&_%*]IDQ<CDO>!1S)$9CC4SMAMT
P4-/V]/4&$YH;XLD$^LQ&G]./H7">K2\V"$"8?[W?8 E)1;8"LT$]50O%2LPL:9?W
P5;P1I)X=PLKKIJ+G1[&DAR"8H?4<1?4]@O8VCSD0\0*&XVT+NK&(%'G(J)[__;P9
PBM\?C\8>YW"PRAK1XDMQZGTD;EU'%:PN3.3<^0XOW=<.GVQAM=.Z4FP9-^93^MVW
P/8V2C;0W8Z13#E)52NX27^3W$$7;S8*D $;A?Y!W]Q<J+-<&4A<:/OVXRMV 28BZ
P"MI42FIWHOA8M$]P036UK(!BTU?V&3[QR!,S&RJPFX:8]C%ZB3X3?!:T[*^=6&3 
P]WA+K<=T2ML!5N#=W93+_*  $?;HR_<)\50LB1>[O'#%!'Y4XDS\7H'M?15"W),S
PP-1ZK.=%D ]FN+0VC//V.:H^L4Z#7]KGJQC::3X1A;8/._#60@H.&O>OS5F3T9:)
P=:?*C%\#F1@V7P]WXW.TQ6OJ--+#7,0V(V.-;!7X'+ZS4&\X1=:Y6F)J%ZVIZL"4
P@9T,<]GGT=&'-3AP=3BD;P $^0(%P :NCK?97K$'GY,7;O@ESG,[*IW&(_P(I!*E
PE&3H&N8P(>!M8) O]'K*(F!-5B]<'T[B:L %\\*P=$^]E[]C[T%7<MZX[HU7VHQF
P=_2JI=7Q)I<="UT>H9JNDTA81X'X_\]2L[^T16'U+<VE79&Z%RE/R84@>AKUQRN5
PWPU6I 7B-B\/ZXU0^XE<4>2NVW/"*' W(/I0-K;CG>-+&1R@R1SC!#DHC18+,0-S
P)=/1B]'?;]+L%L>W!OJ8I:R)T0&>P_$."JJ#=)-Z [Z]\W/=O%ALWM2A4H$J;56L
P3&0:&(.1O$Q#T\KAC)W.3WE73 A5_=U*E5HS<[:A73^K_ ).:XAHIV0._0_<$QOF
PL4G:0$CY&9J1RU03,Z'6:#X0=_^3%3*T]TN*PR6!BV)JFV#=4F<N;%*0--HZ!#I9
P,:%@7OXYE26Y\K57A+@6/20X"UW\9=.-/J,[_G_[;:[+&T2;(G1:=:S5(OS9H^-O
P-F"(W/F1(3?U0M0U_K(<YPH-$_7*EN\&B?;V(;<S_[/V7;RU&;NE-Q@F^$;P!7C1
PG(4CV>\7!C$A2]U/:"99_-J3Z$+4&D<?CY#4?#%=;O6U0&MV*$M;*UL>WF;LI,/@
P5@(0C-]PJZ8?,;66)^A'61^T5<%OB4"E>1(+N2@V>_T"OMM^I/$)LLFL!5F&$U-$
PXHS<<ZK6^1WO_&<<Y$IF8/_PK<=X\8A\(*QJTH#JX4_?8LI^AVVM$P8D<U$P3XS<
P5ZOIWZ=9&K<7!%LP/^JS([!^R/,#385DDW(Y&>FO;:CL;/8]PU]CX2MF#8UZI2)0
PG D&:]%Q7CC?]L"@SFY4["%""Z;E%D;E9_JK$XI%'\MJ09;6?_RM;/*AMYL.^>)&
PF)AEV@;UK._EU$+EV$38'5&I.6J0[./O?5<+[8:[_K8]IKW*;/+9V1+AKN8Y%98M
P#/-JH])+\4K@&=1MHQ_"J$(DO1_G5\O3;[7 $D.XFF9*7IN>+OW"55',N0:(7!]3
P=X:7W Z(3B\LV5>/=U5]/\_$*;16A[I!]_"3UJIF*GI9XY,SZP*P11@L2Q^GZF<,
PS?AJ,DTMP/5IK3Q2$#XO5]9UIQ1RZ=VW6V U!O+W1)C(4]D8U-$90$"NP9^PNI8H
P#IZG>T7-J4[&O=W\8L"*UK\7(4@ 'XO[[4MB_V;=CP-=8!Y <XGJYRH=-Q0)6<Y?
P1M4^N'H[$$TA[)_F)S^9T9WG<<P>WWLGTZ8VY41)H>EW::+_M%T<6TA)E0=UJNEZ
P^9JSLG8[KE-,:''R<^;M&+>#D[,.?KHF;'2['G+6<,UT(7#I0FTXU$,B8CEB*\DJ
P$T>!=\'/02*M(Y4$R3Q(#>6X!37Z'7XF^S&FPY81+KFB;EG;,MA08@!Y?O/UB:?D
PT >3_QEJ=>HR;[Q7 L2FAA.UIV,)FNL@^A_<@U4_R[^ GY-0K_WEL5"I@CE5<"[*
PR;M^_D/ ((RY9^]E8RE8F6@X];(ZF%S2X-GA-C"%V"[.,%:P?ALW&[]W'>U3W2/@
P$F"ZU;/+(JQ5-7T^G?X"1683>U2%FC"3'G!$I,L. MX622'M65C-R5&H.J*7.\'X
P )V(Y:QWN&.\T^9O_H>5)&*H)6E6[6*6GO#4<S&P*QU<,40O)("2(1_>(.D=)M])
PLM4WVOX3Z\T=!^;+3]\#NTG\+]K#+0__W/9[F,\\RT?]7+LTWG:2J''/H\S'YJ0V
P /-!/1G4QDTD:<HYK-N/@@ AGGK _I 3&C&C_[OUQ29)G%&P9X^LQDLB^.@TFQ J
P:U.*,I+B2K^WF[3[:0P&HT'.+8Z\(]L^,(#FFOA,L#X1"?/8H43R9;T[3.)<7$W_
POX$*[U99W0Y=+$E./6L-^S@#:Y3CK#I[O(GQ=V>T(_T.W[R_O&-U,+E)>;/7/!$7
P]9MC'0H# P3@J.H=?T5S04(_J X*-.A'E2+FTO*INJSADP5YI1,_**$I=2$)5-#T
P.O9YD]5'=V^&4W-4SC[XIH.6Y_\!&JO_D,JSF[H@!E4R<J%U>(>I'$0V7S]GG ZJ
P/;FMW-0U$$E^N7E*6.*R49A0I&HZ!ZHH2PT \2D^C:'M&+#]&]+=:*_HG ZCEEN$
P-U%$T"@Y&CN"+D<8G(/DJ-[C[OT?/V(4ZJ_D9>LW4G$^DAN.&;:C<XV_3G.2?>92
P>6@\R/R:YVOLRFH+E%3)3X5X'QW\@J:P5*O09DG-]6!;R)X_X_B]BCQ=EQEI:(FU
P2L:PDLAY;^D**0GQ$@(,,*]THM+K;RWHIHX5*J-U,P*@R\43CJ0S[>,E$:ELNPKR
P.0I8+?6M7V):]6'FMAX(3,UF=7QK507$J+$2FP+9)'CLB#W 5GPU&.X^!&&%SWM"
P\LWYJ;\T1F[6:ED8<__7\Z&R*-V6%$<?U4)330!:]GG3 QINCZ(=+J#"Y,O*IMHF
PR*CP1&C5%"M\DZHI2]_NC9\B+\K>C:UADQDEY_D[PUHEJVJFBF].+M3'?)E1@)^1
P$=BUE49=A.^QU'ZV#*3<H3!W#"Z08.JSQFUF<F#<N^/L@JWN)Y #:[>YY,FAH<MT
PY8G_7(QF=8ZR M%1$31%T%9ZS4SA+FM6.CH2=+54"2V[/OXF_[X=H\@&=A;&N#L-
P>L_Q-Z\JA9'Q"\NG.BEW25RK];I7'I-:_$::'^,/0S_B53U9/0UE?^IC6N)S1H+>
P46 6G)O=?U^A$Q?J]HQ5' D]?&DYWO]E;@7(@@0MC0;'YWMAG" '(R!\%^XX9\[D
P="!&$1V\-A9U%!D#T<\@4BE\B\S4<1NZXJB^1!9-@1C'=:6?#\X#!+605-,:/1G.
P05+ZY]IA^\1U@IR/.+[,AA6>HVK^@J43#1S1U&Z<OZ:2=KA/1K)WQT%W50F1)SS4
P3Q4'-=$M%=YT!*)GD/!YBJ61<97\D=E[@TDHU#:OB57IV<<:IRFD4&(]3.(1%GV>
PY@!^9!/=6%>4!<'=T+ S)C2'F23Q$4@.K QX/]:18@5[:*:."@,7&XZ!K1LSC\#$
P(PQGA1;A2N<O$A;/SFU%EKSKI,+_4,/ET 2/Z,.\U3O^WE0?6-A"+2$-,+.$YNE;
P+JKC_"Y=<[ASZ(*A*G@X,%].XSK6&"&$6RPX1;$,3%A1G2@GNK<!LZ^->H2P>U-E
PB:I^^;W(U*\HY1I_'>;-I!BRV;,TNLN$-IXFJNJ\1JBEW?G6,/ O(+:KU?T^2;A.
PVQ!F=?643QT7::+"T-<KY^SM=D 4F6U0B45_J$BWZVK;=0PU]5M2]K909ZLFJ:=9
P=\"1H$$_X..^C"Q!L\#E2:C2&+\PRR]7/$((Y:=MT>>HM6VT/F3_DC:%0+RA"%@U
P44"".0LX2/2):PL@LE,[69\EKQR53L YIXS!0H8X0PDE6*Y[_]737>E01*2-$"XD
P*"YQWU6KA-K8YSK9O%\=H#:.DMKD@T)()8,E:'&5'U#C8I@5:;.PFMA))<N%K?L"
P6=5= =@ 8TZU,UGX_^2E#LF&AN"T=$&5]76GXDS),24)6W[W9WFWS+ZOF6?'0AX<
P*B2^U*<(/;7(4K_#3,&@:@OJU!DA+?$ID%P1:6P9'%GE6VW8#,:8.F6;J;8W3;1E
PC;D:.8:E'B$E/C6EQW)\4NP+B/R6;TJI=(@2VK&OT;0TVI1EKR B!>W@+ WZ?4M!
PJ##+6>Y(NT*"+\['U\,M+ F.:.Y+XI$R1Z- K11PSNK'Z6=M\MTUW&?4CCIY=9".
PG?;SP,_[\9JZ?#R>[PBDN;@H%NT%TS^1]90,T@8U\NP6@VH!]&"2KVFX-&IN9VV6
P!Y\JSWW72::12-(:8H\+)%'V,D\PP:!;E&,$TF[/'7#]+H3QPUI8M%HCLX!])Q'4
P2@<UG\:=/9ZJ4@<XN0W8HM[:C>D)$#*,EB1[ /\<RE3H&#I'G5@91F$?0J@<UFEB
PHO(Z>U$&<,[/^^OY#S;]RK8 "D%C":UN\2IPL=U$]45EZXN9>PXZK&%19[:HJ!5*
P8VR#!H3,S"#>#&GVCQEN,O5X.>\W(UQO __7/)&U)UY/V:17 SO>3./<EQ%S&0:J
PFW'664FX,]>USV[\;20OJWU(H&BZ&NX-?/\X6U@A-8C>4 FR^OM'</UK(%EAIIK0
P8/;#H5?01*@WO>8-6BM[K668XP_!&?&*M?A',;H:\6_X@M]@E;3WI6SJRO8\&38H
POX%G)4ZI2MR)*>V'!T38,Z&]L-9X+36C4?8T!5F,;/",$QK 2NS$C7W#LNV_Y2,)
P(B.I"V36^1^JY2-7-LKZ#P"" C30ELVX2516^1&!4'GR[I"6&HO=+F-+5'D ?-&$
PY/ IW"5A.[25*%\O'$WB YP[[0/9].!_VD5,0YZ?H*GJ^[F,]AP=X QE1NB$X/W=
PY,NM.BS).=G"41A3*X4Z6"3QW#Z>TGS@(4&N05\!=0Y$@I$SW"4,N<[$Y5IK-$R*
P_H%=4+A1+V$[W'L?P<A^H7/;TIW?C@K/)TD5J6ZOR^VEC5)J1 ,+Y QU&$-ES0-B
P  >V->-N_RZ,9LS"?^6!EDFAN"ORL=Z5'":OBWC'&^B/[1E)QH_RAE*I.!1(*]&\
PQ-(4!E08^E^YJ[82NZDL2'+LWAJMF;A 6W!#Y>X1[GQ'$# 0YM#F0GKE!C6-8Q@J
P)4-8,>8-IE>&'EYQ(]W-GJV4I:LXJ[E:K3?4&3:D<X3*M>UB35[2[L+\E4R1LV*C
P;+XT2^^%!SLYDDC7[E'.'J:I%D P#FB@%L7^\#'-_FL3,SDK831>^R2],B7*7XFZ
PZ?CPLMYQ:+NW>;4P>RNG'RK@)$J"8YZWOJ2S)S%T7(O_[SA#0-\V[E\5(M%<?D^.
P@V9*K*^7>K3AT^<VML4 />GSA>,1@];0R:T+$)56F^K@WW9RN$8-?Y'3(T^;FT8$
PZA(@8&=O>D$Q9Z8++X^@A'L)4[@3MSIR7.6TBY1:\AG:_=\+V2/)V^\V@#-C\ =8
P-O3I7K0T&*GU+_#R/: &GV 2P6E5R8-4Z[I\)2U)\&&#W&;L3QL40_<1K=_&2KIZ
PO8*R:TR>'2M!YVGV.J(Z15WKB(7FI"U/B.Y!_^.3H=E%Y'B)A,I.B9&@A3 +1+="
PSR 8[L5AGI8])^9"TTC@D6]15*JA+.JJ%43=R- XVA6S*5HM_N;0KR</@%%)O6:(
P^*-3V!4*2&=KV,:['!"%0TKP.M#;I?KE/H(&B*B-_ 2R1SSY=I(.RZ->!#(X^*_5
PW'S+.,PY'UQT$)X+]1X+C0O6,5;\V"B>D-OD$XY@L+*SKYBCB-:0ZIL9&,#ZOJ7)
PB;L[[7/*ZL</N(HJ(4F"F0@DVD$>?N^;L+'X<T!+CWA2@:?I-KX]QM9DB@QAGO\N
P28KJN?5J^4L+O,1HA6<1RX-2\5^X#&I.8>'.J)AJ=WQ/*:3_2X[O$^"K]\TZ.4B.
PN\0&:1V&DZT=Q+\!.VA"QL+&Q:45$%+2<^TE7D=N$F]!B^DT2(;][<'RZ=I]4'C?
P?T <OR<!NY36]] SVM@\?M".JB*]%[M\RQ3EB%M1O+N:FF2._((PET_^*"V1-TQM
PWQ:HYWH_,4[J)?3PC[JO> GZWN&,)D'D???+X&K,H4A ^#OGQQ.V_>7<C @=I5G]
PXP8(@4FXZ1DH^*=%^+I]9[-?&7Q9.U*KNZ.5. &KHT=*9)EN_\3%IB+#OYDW!Y+6
PQ*IN6=MF3Z^0LZSD!2G07#V3K2UW'!@NAD_H\:*8 4UC-P&771,=/J-'(H,4N*<$
P96LJ*JV]N7 5[@C]\E2BC0>G<9?1MX2?@-H'-X4?EBIA@T/<7#N'Q%HJ&Y%PU,\G
PN!'(_/H0WI;Q;-,+"6QSYT0[#S@/S/H$B 1O+-1MPF".LZ;C(%\7BX-TN4U)*GKG
P*.+--\MP$_H9[Y#[%;?Y/;UT9E/1\OHNY:CJL5]IGTH98KT):=+S!ODS"SSK:=//
P\2<8NC;M-OJPGG-C.G@$>D;82[U6:'GLA4FGQK"Y35$SB7!+L*(4$5I4<P6/DM'$
PGN@J.-WX1QK9R;R".P?SE:?%OY9*&/PN.98_*G]Y6)(IU'560VF]M<*X6^ 2E88+
PE9[]2:9;IQB .;ZS<,;*/BPV&P"=3EXR+YFC[:+1UJ>R_Y70M].M_?JA#GH<;KN>
P!)UP!26]DP!_X_F+<*<3]13C.QRB@J=3R#$'NVJ]:XIS 3(1<]X==5%.$J-X1!C8
P^V&504LP?(9(5(6I:U! $N1/CN<_OYE#XETUR.8$<);%S*@SU>R+CBY]C7ID%L">
P7T:]2^[(3.0M*@]/?)+;'F("E FA=UC I2:-D?;N9!4.=<JSO1;GQ)W.>%6BRQWO
P 7]?;F"'R"EJL^.K85Q0Y5E%G<(B?*.]/?'Y6D,>8DYM-[L&COUW-ZNMCS_;,1QH
P<YB3YK980H'P).7,SR?#!PU41QP<<Q+=]859/V1OW3[KSUS#^XICKI#R].(S+ROI
P,OD6@T19&28N#&=5 F@M+R37?C"J@I.:V'_DL^.Z\B]46EKXD[6QAZ:NKOI\$0KL
P'*/Y=M_R^<$.RV5F-@+H4#GO"^CU?JZ9]$5NY;EP@@V=BQ"1[P^VTT[K'@>B[60T
PY0[9^-3T/KZ)0<D/.&JYS4\$WOI&\%4".X2;+$!BI$8/75H4H>_&I=-<I1#S**_4
P UB6L\N^M0Q7N"7!JOUY02O5:%B/F,Z^_?@JQ+G1'FR;3<]R@!%,U>J'M4VH FHE
P^%KEAZL*@/>.*4$&W]SBETB,2N^S]];Q\4G$95*@/&N$'RIIP8><'*H9NG*)V1.^
PG"'IB-G@O7Q-0?K7$/]RM&%]OYC=BX]>:)#Q4$L#E.!P7:IY+)07();:*8=6[X+[
P5S*EW:%-XB6IYZHN4L*"C*0<IS[5*:->DI)FC+88"&.($(*!08HU0SK*]N.L>Z*U
P#_X3:S 1MUR*HUN(,=RQS?N5FJ?:/8Y:+9^3"X,L!N#"I'SRQE$NR9=Z/Q,!GNN!
PF(*; H_'-#GV##[5GZ[8BYD6O-09^.8][\IU2L\I=0F=3;LS:IN2RS%D.7I;Y1OW
P^Y'<]N]9BSFG.^<S82*$]OH1;SDN40]W6[(E'0I@?.LX&++*,7*E3^K0=T+SYI2R
P7"Z.MV.$C^SO-)X$-A:D7*(UCG=%,T;<D1FYUAA;R4C]MV@=)&9LL%CEG^SZ/'([
P'SGH#E"3 HJ3#(7Y:V3KZ4_!3;_N!YX80>Z\@U)L5#=(55J(%&B172XI2:1!G 5 
P[\3+*ZT<KJUF5&I<,2!0;K@42@FGDVB-!U=2D&D*.!!#%%Z'RS:N&P1"]X^:$Q2^
P$^K""3_CHEZ8#LK](++T>I;IL(-HMZ^$<]',U>?^]$73("<0L9_"J^OT@*]S72;_
PY(=HJIFB+GB>B(UEBMT/9(?0K;7G'@3_S$24T*X86ZC)@#D]'5&M+/YGAG%_*4N'
P.<%CDG;-K+E ^'')E0Y3A$I26XR./YPBI%T:(#P<=P'MADE6O_$_);FXF?)=E6 Y
P%=V:W#WOVA([;Q<,D-R/BHON@N)6"E1@N',J=D''3.T6#\C+V'L>K3&3DB^2Z]_I
P $''&9CSNU]1L13NKL!T0C3E $MW_+AFX&/$X-!*@*;E,-^T!FR>%O@/RMU,9E?_
P"(;)Y!:I+['I@3Q+*:=F?'R 0T@/;JSE'B,I)*I*^$;CC [2\RZ\+)6L[FM(2T$*
P;H\HD#F\S2A!!MZ/.(KGSK0CAQP1F+4$\.!%^7H.1!PK-A:2TL8$G-5+)-"Y;TX=
P/7^N,'%6Z)Q:H U&(.PP:"[)5X%M " #!AG^]9=KU1PWA-9E8K H":]4:9+"I8=F
P"&8X7$(!Q-4V85R'A6BOAP<'YL'%\<+T,RTV>(JI*+0'MFS7+R3\;W45(H S:C >
P?Q(6OR[1H:L0:IT_PQ6':(M?6_=F:\!76C/!]%8B9,KUS[E;D&Z8J,N8H7#W]?1(
P)Q&_>L9B[>,L+4? V HX/8MMWO('O4.AO.DLER-LORN@\\*AF7PA F55?U' 0J2!
PSEULH]QJ0IZL8UTW2"Y>'*>WM<S?^]\_R!C/!BLQ+'SJM !$T]*BJCGW9!FYQI$/
PT=VRT_/*T1!!EI\A38,IT3="!Q^D$28_,%=[>>OIQ]QH_QXY$6U,/=1 Q^:SYU\+
PM?PIYFJFT#IXRUGIL%@\HM5JKR@K3<6B/,:=.>Y,V82!U_"&6.OP+.>&$,&>;_^L
PL3C%D(J>QQ3NSE,FH;I:F?$=*^5B.MJ)8/D&\4/E < %1CTW3A#"(#.5<7"D91.Z
P0*8_B(Y1U9XFX%GU3%/H+ ?UJH*2*&(RI5HJHMLR-Y<*OMXVU?C/5%%[INO.5<*2
P7<<RKS4Z 2K>+.1<O].?VKR_B8%/:N$]=7*'$4'#''NW=RXT#^2C5 1UJ[U]N-(B
P=QV4F:"C=L%4I6:M/'OE\-$[C)OFDA6F!Z4%4+*NY+4+Q\M!U][TZD5.L87GUO&>
PA^/2H4?$75NA0^+39Y2:NW)FME.?))FV;9]F<S'WP;1R5K:AJ'L_<OI&02-&$F"J
P(CAPDT:A[N][!/6YO*521#BR\^Y8]#1+QPM#P%D>2=FK4TW9M$4#E-5EQ@]N1^?T
P%;"V7XV-I?'H_\C%ZD"7WQ_/:R'G=H8E;S%AU0&F_X*$%/&::,-5;+XKLU)4579F
P(WD0&SB:CSE[6KW9U0<T<N$#+F.>B=&:DP[$)1F7NM"ZFI@3U^@.W^E.!FHZTWA(
P)9'TEFKL!Y*L8$=D0^%;5A>.19/TV _D5(KIX'\MO1%_',86_#?-TX7GABEKB)E>
PC3Z3$$F-5W!9J08K%X,V5O7O01+\&I]6=C;QC'(1I87@;P&O(=.OZ-!GRKCAO1#Q
P-P5G@;5ST_D''@T+X:*RE;33VMKR\,-<O7 H"42#N1S:IA/]9]I*3F<ZW$4("J8@
P^/$$%/[4DA*\S*=@B@'M))_KT<%<<@<1BL>JP5NB%R1'FDUPMUF3E0B;)S,$'N*L
PYA%5K"/6 ?,<)[&[&0U719/2N>";O7<D:P]]//+DI=(3V-!);$<$R=XB2BB=9YHL
P'+IP]D2ROI,B-/F#-#W('UY#1;;=#3(=P\P$ +#E^YS^!S-T>P@6&W/9RYR[SE"F
P&4?CU <:&H\4%@W#NYV)\6E:;[,I#^"'@ZE#.=":I#/4]S#CQH>@(_EZV,^)<^J(
PZ$+S3[FY/<8MF"7/J*5RBUFX=^]Y0\D1,RCO[TK"?+:.L, JUIB@B$IQ[V#T0EWC
P 0HJ_TOZRY2W_7J K/V.<[[*PU[>T%4MGS#3MYU=<IEMQ0/W$F.8I)F>8#",KG$@
PCE^TRJUS<,LK^ IPD%,SLLUJ^@<-3K5=(S/_DW?YZR/"]5W>E/8RA<KB(G1,[I@$
P[3_111:)G'4T+Q9SL.2H7(:  CQ<Y0Z,)(YT!D!*.YWB/#8RETU6H_2NA,8?3ZO'
P)%,8DP;D>CY4I#,:&_YJ$)N1WK05!ED" ,DFQFR>C0$,R>-*GDP#L@:XI=\YQE4N
PN517J$-4J8S+#?9,WJ (;]F9XIUC^PT7U1Z*3K9=R,H?K%UC7KK( GD)38-4#1M$
PSGSCXC66)0B*MPV&K-6@^LVCR2L"Y/99J6I&G@G/9#M_>M+NPR2;LDNMA.#+Q9;!
P!0T2\ ;]J:JLH7[WC#?)I2J /GD\:&>[*]R.8#S'4]Q<DHBD7#@FVH ]@/@T #PX
P:IL+$.:21VP9I']F]XD;*H59V:ZR0]LOP6=D@<WMSB3,]* 7 T(ZL)X<LM]BU)I9
P*GR))$^&R@_(V//<YZ'Q5"NZ8)CG)#&HOQ8'"$6EG?C6>OHV0B=V&<FZW1"[K7KO
P [111<1]?\H_QWN8VO..\.JBH U.^I$SELJ[3-N%>=SL/8!K-<!D]S_/I3*]K%_Y
P//5R"#-,U.DL'*C7]IR"URKA?N-@Q_CH&'\W2I^M(O#;2R,_=T KHGJQB1- NJ1R
P5-O?93PQO=]'DR.#:A0+W_&QZPTUWHCELANY=512<8/*LO$IIQVQOJAH6RBN#3RP
P?9P:5JR:-8A4VY2W,B,7#;;DVO /T!(S>%8,.K,?@<==]Q6W#RBY!>W%[P(P@I *
PCU4OEX-14G8EWFX+,SNT6-2G+$-.]H=.H:4"@E/QC#9CMC(<@9!VYSC[;C]&ZTM=
P'7?PZF"KSILJ#+(1%;BU.Q:6#F]B^7Q5KD4#I<\KT0P_%Z?!3_-^) V27LQPD6RK
P(]7U9WPM"UM440@ZH:F.]YJ.I?S79J4<%CO<AKC[<J9[Z6YSZREZ<EHZ8B@IOZSX
P<V6!80SW!Y:0,/TX'S:N"$'U/L-P!@Y))/8BY?<AEMXC6Q5"[ 7O$6DD8XIK-I[G
P4;*%2"EZK)HAN??CX)E< =^$_\J>V%\06N_=[_C5BL.(Q0E!^KIXKYT,(2F'-WJ>
PE_8Y Y^WRSKS7K@%2U=]"Q2I,=3 $6JN]TNA;MCZ_5_0@8B_[1"8H5X$[=4R%-L1
PJU0Y0("<2A=+/BKM;1-SZ#&B#Q7C<(>$PV!"G@DQI>:7=-^=[I[-?M>LK@VF$D7,
PM[*> WVH4NM]\B_(;[$(V%G'4_?B=U#PK([H P^)<CWP?W:%%6&QG=LV&644I?+H
P V7&'NP:8PS20*[-(>KPK^,N65V<?56]V2?XU&)7/H%PIWA$K6^@Q>Y0JJ"R'*^(
PD^'H(!#]+ \;M!S?GZ:VKQ78]<6;>!>:[,)QVDRGKY(Y&?O9TKW,@H0P ADE:L4I
PM/$Z/+<J-#_IV9>E:&1XVH!+<]!LY34T)#/P .50_*>KJ;HK$!,CWD-;G?/GK^9B
P21XBE:_SO2,R8*01,%$M2-4.021V@XF#GQ32%)#XVMPBUUM!A9U'L]NV2\A;_2,Q
P^RO1#^"G1]@>EN "=OGO8NS,Y>.R#3;0EMG2,G=&J"E>W4A<7[L%$K5ZG1RK@Z"G
PBPT)5PWDBR"DGX>+D<T$-"O;KG9P)SX( UT"!JX<SOB'*6(>RTRJ#VSW,UV\QBA\
P</!!'O;?A(SS;9980V\\L$Z^=>0[16C@VC&'I=,'@ISVMA&P;R_J3]CE>QP.(#BP
PHMH^8+;]>[A[CX7)7,>+*;[@GLV!4GLR=[@4.YZ07 TFF)@9."Q"U,CCBT]X9Z11
P^W>0AB=[0#I.GR]I]NDM&FC WEX!IH.Q,;M3=854]UII)(=&( 2W;@.0\#WH[NA;
PPW:&E;MTV,3$5$]9_$(>3DZCSG9N)SLD9V&F \0FI+"%X5L+CFB1X\_T(E<6YK\L
P;>$9%4=L][,(G3IQ7=\^51R]F?1MW5G:(.4S%:<WA[)F5'('\XZ*'[7?2T+SO(%"
P#\CC])MRUAS B$$:\Q$>]]X<\#=P\BRZTC%#)AHD/^:?HT-_4;:/E,I1THY*[+]2
P*H0>82R_%>K_=R26_+F-1QEH?IQK&N%4T8 H2JAV+DE8:F(61=9E:X0>YVY,14GY
P,+VD0>$X%+GE]#3%2055S$UP)*0V2Q=9K/(/J0:E@M[LE9,"(D[MU0XQT,(:85QT
PYP77UUDW9=EA%,0]9PCX03<ML#$2,," J;//H5S+N21(TTA=2UA1SH!$I)< R;(^
P6"[;R'KGN;.+'7 %L(H$+-T2:4*<:5WC6)HY,LR[EL 2Z*+I55YUO=F^%#:7^-P[
PD:404#AKXE--BO-."A7F4'GU0Q# D^Q'.'$B*V.*&U(T__RO?6<9SO;OD)S_@KE2
P%2I<,9EJ)*5WZ%:1\LTB$GZ-?!;>%]4LH#P!Y66H;TL%_8T:%N0;F9C[>',OJLM;
PRD[M65)K<\!,)J+@7B2/>NR@E*8M JH;"H_.6@)8UOF+GLQ>@CQ+MXTZ"^=QT-6 
P32<?$3J8LZ.W+)-F"_6W37G2* )\,4\?T$PV89B_01<++R5)(5O2"""/9$S0$R1/
P@VKPZY+GX(;1 L)<DJV9Y>/V :\ '')76LH8OBC[%)O;'!:PS 5NJO*1F-\P>#&'
P#XBS/? 3.8+%9*(</KV(Z"M:)A>4=+4N(1C)UO7L\U(#'=6U^3/5>8W="[**;GEN
P7EQ^)Z>,\B:-0<=_-G'?I M1%6Y#LB:W?0O895]/XTW=1DUQOKW7?%*AV6Q2IJF,
P%CW4,3_4:%)-5_21N<D$^3XE0<%5T+SJK_'^;0(Y>X#[69QP3)HJ1Q'DPJ0V.D22
P[4+74HI('9@GP.;*)U+^(O_0 @PQR418"8C1]66OA@*CLV;4L[SOWI]Y_2(Q\G/>
PQAMK2>@A=^)77V>=ORA6J4X!8[G1K102!?Q.BDCEU$/#\54\@WE?L=2/9C _G6OW
P*9-!%,]9 G=D,MYAQ/KEG0L84H&U01B@?(-ROG:F?*C!'^0O<[F QB@!/?RICO<8
P+S ;.WA-K/*I18$1RYXG9YCD%G5_K71EAZ&1'9SEPM! U"%(!(R %?[LEX#O]/CO
PV30DCF8HC<(<[=#_H"R>NW6%=VAI!=J,H0@;;.V]P8(MC7!W<W6VUWI:3$9GF?7$
PS++S/15A>FX*3B$XH(A0]5$J\GT?]#"K.IY$209VGKT[]>-W79GNN;A=#I)<579;
PX.WPP_[?+GTD9OTU>J=B<4P9\IZ=)KT$?0?KT4.!73H,H%W#++LME,U^:P3NGKW&
P4;K^+3F!XE'*,VGMIF))5U23U<Z,HD4G(RXAQ<]/J\N1/ZI[@X@.V4_AJ1ISOD>+
PP(BB)N[EH$9\T-0YH%N0]%*^%>.@H;^*N+1JZ$&Q^^1SM] **X,>-)P=;Z]=3D<C
PLTM5WHW;DTG7U_#+RY<<^HK]]Q3D?UDWSKD'+OOU+:&CYMAN6$JQ).1\IX6W'+/+
P\ZG#+:\DOS(NUFX862&^\P&U)4B\?/\:PVM?IEF/)G/:WDZL21,9&*J7NQ_O")RH
PIJ>1L/QX_I<%^=N+.@SIR,$I^IW"J=*#UG9VE 1.[^90G432UV>*-AGK@V<^(^]&
P#L9JDPV6T/1SL=OC56BEC)"D^Q2V?W+)QO(U[G ^2 YM,8H6GYBD(5XZHFLP:@PS
PR+,/Y,>/YS2X14I!_1Q D^[[QFWSU1'5$K*O[F$5/J<"R*3^R$'N)Y+@$SLWV]'"
P[#V!%#F=*(SXYN$SA$W1YG7[)S#50.I>G>#5%:AW52NZP1\+B(-#D=S7,KV,Y9HL
PX39>'E1PMR3+.V21]'')Q0H*:DS:Z[%*OA]%+D=T'3C%RCV0:TQF_%M#4<[W] 27
P^_4 L!54;:5/<O:] 2A3;A8]$G9*Z$X&9G9^0"R*LB1%;/D7P9(GO">24(B?U/Q3
PS2IESR"+3,A ,C ZCZ\932[UQ 'Q'T)KS QW<-];XG WTQK?<QA.L%T9/+,Z5CQ+
P[\P=E/DNHJ$ >6_'4!/BLH,+?28&BVVWP5%%W:<G8"'@3SVO2]#>"Y3/MT'M)>CE
PLI-11+*21N)"PK^+=NQI%UTWG+>\4>12]4\$S  C,CI20L9%W2PGD+!^CP/+1_04
PS=5S'J4_*CC+/YT.Q,C]9R<M'/\QQC]\9SRDYX?V^==!O"TSPX&M-QN8XCF_= G_
P>M>CY#'G4WU&+1LK]CBFQ_P,S7HFEA>((<8\6$=G-Q_=@@[][YC5/C"=:HBUVAVU
P TF;G1PC5KS.%![9Z>"@%X;G'J:2Y J?J4Z9G[_'2B:F'#J=Y<X(#&=+D%FTDORY
PX5%\2#6'YO%A_:RE0Q#A[+VJX6<HAPP&<?+D#Z7X"<=_>#TZ=F,M'#-<&0N3 Y"D
PD\H>D4*_+8RQ"W+V&]0D(98DN$3ZHH!5O5N8 X.(VN+*7G%Y4B[5M "/8HU('(5?
P$<N;+^(B6<_E1+UY*?STM"))O"$M,"LJ57)ASFMU%C!0'#K_#[!6^J@DMD<="/RP
PH&J820,%<?XGL8B\[E_59Z8( (@N+:)MMR4-G"F%11V*$*O1J ^1'R5JR-ETQPT?
PJ-26U09PP%[+_?T.9XI<D1BJZNZ+Z>G $B5I?,VH#XW5G.S#F=2647K3;U.8!CY 
P#/PLH@H\)_+!/S@LL1B.[\")0JC8M!X>GGB)N6TK2U>28X56N>MDP2,?2\GX5O7N
PJ6:IX23^WK@"\ZZ("@AXB63IY\H5-N6MG/D5-26N)J3N853,[?)FUMJDP+A-K/FG
PNFHKA3?=?@AH/:QG:\>U)2#%*4]D)LTQ<X',9@6DG6-+O)_?%9[T878-U;0!_4[U
PVI^BF&-OFA5Z[,/+3W+3O6"#6U =.#H;SR4I"I&1/E>:=WS<Y=^1TD0=DP'@I 7*
PQO.C?]9%B+IMGH:_<N4E],4YERL-1%U__T;CW71^^4$[-KC48-OS#)Z4^='_ONVH
P=."?S:'L!,$3WXBA2">=+B<3L?Z9Q0A4#/-]:@S:R<\U=;?Q?1+%RI3 J?=31-X#
PD 23(R"0PK#8D+=?,2" H6VPG1K7QM_BJ!A),X%>ZK]P_8I8Z>,<.;WU LK[T3U^
P8P>7GV%.\9NQQ,,>1&,;XH(JX"9:NI70SI7Z:]5BGHE705.^BCP:+SH>11)TBO1X
PZU5%>U=@8$ND3T7T2T*N2Z_+/$H26=J?NA)V2O4E]MV3>X9IK=C(33-:U55G]KV(
PF,[Q!9]/%']*96NN5D[#6#T OO67";B^RO=(,(8.3DHT2IDGGL9L\7]K?_Z"^"_1
PQL:+&< K? @S2L+J#=LHZ!S*:3J*I?0YWCI2'FL^4?4[9A@:^3,XY!(7"N,%;<35
PWL<5)(.;'_@H<)#)Z.L\!\=KOHO9O5LC<JEZ+W43(6]#L<)-V$:J@ 9,HWX#I.65
PY[;A0TH!_X"\;ZU@0O+X<_ PR=N^UR";:8>I!.NBJDRSX-(&NVNR*^>Q1Q^;8&M=
P&_7?@7L79(7+"LTV\I;[.B:UJU4FC%N GTGY(?N0)OWUG_U @]XP\TX2*5Z\3C(+
P-DW@E%N,/OLWM:!6@@3YL8G[B)\]9Q,US65:X^R%R!?$1[[:<]M#FMJ4FE]7@N9\
P$8YS-@0\ G&3V YY.UZ,^JEF9CI,T;*12_T<Q*L@0R$3$/X'RG'"A"E89)M+8KOD
P)GJ+2;=_V0K"A,!MQ,<L*P.GC'('['5E/Y7MX934\8(^Z!<CR8$YF(.'J,CB[/XI
PU?FBAHA$^;W;&3=&A5XH+A; W0;#*1WGGTR0LF9D,'8N3CGG5@**<\=Q,-]LE6<T
P8I[.TZ=%6/JRHO+4=MCQ%GC?11(4*W=[)%W.%JTB;<^UQ\4(^<,$=88Y0DV8$9,Y
P1E8OZ!%* CE@*I54E6WA4O\MT%FY)!>J!&6JL)YC6_Q@U[$%O*X#P&9DF1'*4+U3
P^.@)/&C_: <*[3M/_!_?<@LJ<BJI(]@":1(VO:V06%U<?G*N]O-(JPR%VHIEW'Y.
P+QLB:1=> :8)3>=G+TM?!/&94$T X)/%:QANIC^!).'EHI0W:MCWWL>:2$X\J5DL
P423),;,M(+=88F1[O*"A![W;/@W=%-&.)%+(X"0-M;VX572]SWYJ=O)Z#WY>QICW
P,#:B?$TK#$&)UP5!*L>]N[I1).%9 2!Z[B.X(^"C:+N15NOXBR3'9=,Y:&Z0>>/3
PHS <#WH9(4@)1[Y"I>"@" )2%W-,?@D ]H3)D:C4"=*^Q--#$,3@,,*3\WPO/L#^
P_Z-[<Y&&9"HPZ BH4/44NQ/CYZ"C^CZG.Z-H@/I@/\F#ZHC/NRIA"'D ,2A8^ B?
P[<XT<:>"&_Y[]!U(*T6RJ@C;5)[$@,IAME@ \<L/$RHG\:$'?EA424N>AAVF,AM&
P3E./0DT^5C* GLKN+M5RXW6?Q%>#J44(:> -JJ_0:#+1D)8T_IRD51'S9,P#V2\5
P*MSID)=+AL)\MT/8=6G="</>I!0U1.9R2!8X*[O)<)B0D$[ ]C_Z3"SC@79&(WQ$
PI;K+I,/'H0T!<RY',46]&_B.;&%1"MY.+&7@PUF1209=:6I6$A@$6% 'EF\$*:P9
PKK*)R2#;=R_!_. #Q^PC*FW(E3.7 I(H-.AQ#J30__/)O!M+,C$+?)E2W44VI0_4
PJUF%/+Q]MTW\>6$4;26[J[$";G"?W #M_NOI>/=)!70N-.Q^^5K!?.$DPF.HE(C%
P0*0W,!R$)KZ9WA!*5#@(6\+ P;<])4X2F(2!-DU01>*K_;'YNK)2U$W>P"]D?+DG
P0_FBH"]>OWP^T6*@FH$(H$JS$YS>_%2,\-_[8OE43MC\DT!.]2]3:+N]"%# 5?\3
PQ]9]X'H XE+UG 60A,Y*X89&<3\9KZPCO=3.#6H1H'Q*Y9#HH14OU#6>I^IRER,;
P2@,C?)[BHG[C4LG)6+H)NT6KR-3/"7@,M$*;S)::?<8#+>>?04!E^A(#LY<0<@4O
P^&!C>Q-10R:^F]XN?%[TN+JOJ<]*TVG7!J<33RP:*Z'18K7>]>C.0RX0,N%ALH,+
P6<P0YA4PQ&NM+'9 :JPH0228^3.:UCB:(E0;[5O9CGG77+D@IWU]YH+6Q0VZD48U
P[V!/>T,:F+9/?:"2N]?S@RNO%19!W1",;G[C_.#%:<'*(^UX9GB@SO>7VNZ/:N9$
P??DI%D-50NE *:>:Y"BY7XI2T!>^RNZ*?E32-G[!D1X?&H7F+?/[T*+1\-0?*@LF
P<:R-[=<H#0WT<B'9?, YXI>GGP$9R6(,?4D";9*^]R$[D'3I.>OP#>:K%&:-/00D
P:^X,S.FXAA<.$>49'+:%41P4$C=VN=L.;C KP?%WW /B]L5-T7TW1E=1R;S>:T(D
PV0.R:<.8J:@#:O,!U\K?*R7Z8^I+"0<(.JABFIWM9:4<W$/+&QT<@Z/9MIJ"GAT9
P7^_57T4L*[OW>-ZPGUUX_JI<[F7#MIC!5@V'DV31'+/Z16E=V^II,C?$Z?AK%BFC
P4JKIN$].T!H3*R;1G^,Q'YM'I_D@OYK#8FDK00JM5Z7GPLS74VUO"5?:F>8?.</R
PS?]W<.FPJP-L Q"9U=GNB.R$["?C]$69CAD!*V/9B!ZG8:V5*3Z3IZCB@;_H_P"/
P% F A,3-4#NJB2_PUHA(%@3Z9N7=PY"D@L6;>/T25<NQW%FS<@X1HX9]\6L)3RX=
P"E!2*NN0-Q5"D?#MPC@4(8JN*S61*M1YBPH,J570<:)Y[V\,7;P6P;EZ\<2+>#B8
P<*?01X:KL?!FL74@RVR<!8_Y%3*L]1N66GRN^+K'I/1E3;CU^E3=3\HS-7@KR9VI
PE=E!7D=:W/RJP%4(O(_:?#Q8E21"JAQ,;BAOPZ!H26C6Y6Z-WS"PGRH)="O=![ZG
P-J&_="0[VG+?-^2KY0'QV1[B/G)\J6_32F(3S-+(2U>P[@X;J?LRLQW:6=-0&((#
PA,O.3-B<I%F1\GZ$>PKTQD+/G/=QE-%61UJ3%V6!H6/D]2O@U,UTLE<O63V! "J1
P2E1#X:V&1/1?5'\IL?);/S^5O@FEQ6MM\QNI?Y_IE!6;-F90B&V3( *DM'$^@P&$
P":-AHIRV11C2:[//,6^/##3$<&PD/H85(<(Y+%K2V^;2I [( L6DK!2T]Y0ST:0*
PSL_[21'!#<&*:M(VHA:VD:! _!.Z(G%,RC))%F,BPB]$9P++MR3]:N_QF;6!05P$
PZH>,8:WP>4&G"X<VP2\FC*CFQ<7EED4U2\ZX<4_)4\C@8&*_1X/Q5J+_S"Y8P"3O
P%Z%/)@7M4,=''ZN0CS?51)./@>NTCRV=FI\A80+1&&M?>C)9!+?Z*./$S2%\#U\L
PC%U%U5>LZ)L7_/,?GV8./26BYL(K"'NKY3PJ:*.9AT[D0T?LI.IQ)DAT,/D*5>^]
PK*K/E@E10BK\+#=A[!'AQ.QRG)&^*R4!V]^X01QB_;KOV1>\52=]C^ 2_A_/'72;
PK'P5&M_=$?@Y'Y;Z(8LO](UIZ$SVHDN/,SR*F1\HTV)F*,:UD@F)#SD$3T=.$<C#
P,T'$2%05HP((NM(&6>K_U->'[.#])FD:93.^$X")ZN3(J.9U6ATK,#1]%G[M+RIY
P!";^N\[HB6R,[F-.$?$;:M748N:TXLY++[2\*K5Y3]GV_^BK0+>1:O F#$]O\2?I
PV&XAY*?EEZ5:1BQHT+12XXQ=NZ0"*4HEH&N61!)SJ"^6K#P;FT<*?T%X,!![DNO&
PG6Y#GW9'W_K-SG[C7+=!5Q 'L AP3#L?Y,'VC\,)[:#D2TZZWT6!FBH]X2=W(3@(
PUI0!)A9772!"QWL<#I9]Z_">;?T^%BO4H;*2Q-\Z.1F0]D1?XRR&2W^MYR2&S,"C
PBYI)[X_2GF)_ (FL8<<B#C!_2?"7<*S%[!35N*@QJ=LDKHA82<'%RX>\+?0XD6Z.
P?O\AU>K[DA4'T-%B_)^YU?U-VBMCZ[R1L:;P#0@H"=8 E]H389CYS#*<!>X8,1#%
PYMBX#+^:.[?B4 8/Y;F_,[D$@8KHHK,OA2Y *GI'P?[P<IF B")3^<?"BEP*N_#@
P+4Z(]T4+3TG-D_'&'_H4E(P5NW$90,Y_CXY%PRIIQ]"81ZHVV+ :%D<R_\>AM$04
P%2?5^A%C+7YFL4*:=J-_B(0A-II$^BL@N?U=,:R]$@F"&'4-G#%27K*T)CJU^D%4
P?;>K,K7 W'!>OUWTY.;F,_FNL""L?"[LD0LG?\AT6R8XTQ"495.J!M:^ %M4X8\'
P%H33/;:<:S>NHYC9M(3X#HYC3%W9UE#'*:XF.4-*&@LC/;*&;@Z@8T8O-[/K7XO+
P\:95ZS?3BFGWZ!G )UL>EN*\#AM_.-^F!-%@1?S4N2U^(.0,'A4R@-#3N_Y(UZ+!
P,<W:: :+K"'N"G)5/1\/7K<MZTSZ,FL7LH&K@295K2W?VSVX<'W)()GAJH&A$4 5
PBV,5.F2RJ&F0E%W.<5P"P7AF [(>)RH3!$T&=#\0KWSX,V+P>^?YU#).F2V[VGN.
PXF-)G",1(F##"Q95&.?YYZF)NX ?\&"6[_3K [ZG*<3C+]250XZ92TPNLQ4-+H"X
PNZ4QBU0P=GL+3U'AZ0Z-O2FZB\P*B Z(/$&H0;?MQ+)4D=?-L.@</KC)+)0UZT<D
P(+";X7S%61O_L S'Z+S-G%;W3D$#X/?]M)?PQ&0O;(9C'T>]\?.7R5KQ MVO@OW>
PH'G5'0RDO%<EDGY65T07#R#9FM]$-^+YL +"%SGNP*"?@.!?,LYY_)1"E=T[4LK]
P8A:=(!R(/*.$_Q]O>\$6"5VOWVC-B3821MO6H0 DP _@()QVBM)N5(4FCH$D+S=[
PS>\EHD!-[LC/S7UK(N5UQ=LP#!Y1,'[QG4F')F 0P"0G=WI2=0#$A6,0E ] Y?!(
PSQ2.G%M@2EI+8]E-6\>T+5VSEVU-Y+M/>,NRGK**\,UH5U#'TIQ(>)D#$,O.^UL2
P;<1,49A(];UF=2:N:0>5YQ\3 32:**'[" HW]*\1\1_1*GG$6VCPQJAS/_2@4#4!
P"#N-<8F /C* U'JN_%MPQ@ZU0!HF2J-PA$/8(C3J775 9^3+*R%V)C<[F5L\2DIS
P.-E >.3^2&ZH&3MSQ?>3!GPSS>JU?%Y7R9*2T 8Q>D//*=-;O@$B& W1/T"/DDG[
P$=)KK\P?VY3OVJ7=@&K,,S7'C8=HZ;I*SU[U^WL/[GX]8$R>]BVLD!CNX1%*^0$*
PO=Z1Q^^WL^(JF1#<+=;)UN^Q%YUAAGQ)3XP932B:F#-H?C\>$K"U;K1&FT<[XZT+
P 1/,LALN*"2<14B[LG"^]?H!LH[,!-(X4ROT7UFS,%2_^VUE8+@_AKIAV-X*?UIH
P60&BMVSEM8-3=]*(/>$QA*VAJM)=G ;1</RNA;8)CWL3'YP8M8$4<;#,*_J,R 7^
P+Y!V_+"  _S>A#32[FP2 CK)BW'A)79E"25HXII1"(L5F&6K4-Z912=9!@%5W+H:
P/OB>^?XO9JC9/*_=8D/^72X"MP5IDUV6&S_'!=5OX(SUP5\E@ &N]\6OS'^7<-^P
PMD43R-5'5$]UPLIM1):U-8:RR9! A'" 'E!^QKK4];U]%G+UG4/*\<N>%W@H K0@
PK"5[BI0O1/7H?&1,S[OZ2;+:)))_R^TXHX4XMS..1%D*K1-7DEJ'>20?F"U:N4&B
P?XI\KQ#H$J@A$T[\KLO@EI<SV)BLX9R96+D\AAJT;L-$Y6GZ@ZZX>-<&X"-SAB%%
P?,7"#/\P!FSG"96+<61SY@/44M7!0:IB 01@7>@"'O7&$N<3Y^@X69*AV4!R^V?I
P(W<*@1A$>4J[P 2J1<D];#/EY!KF;Q?_8]0ZTI]Z$@CP4X[[%>]L&0MJ8P6XH,63
PX3<-P6^#WO4M/KETZ7IJ4V6:"?OUF;R,[@]AKU\SC)M7F<3*'AW-]S3+; MX2NW.
P.S<L"8CJ[?(!'904]K]+&V&FXCQ"3%TMG0A31.^FB="]C40/-99-E8[=Y+[WZ71S
P $GW  \+M&>TC+T_7S).$#-,<6M2A5P /D8:N(WH_6$]:C,O0A_ ^!=-U4LO@:C*
PPS 2G9V>&2%0CS[I&M9$K31>[7+7A9RK3B5%C+>AUP<MD%2;Z4B)2F*W9*"3_%WE
PH;,N)(F,;0Y[C<!>VMS-\!ZHKP>=DIP)7;_>;Y?/OR("[+__>K\[.* D- ;U*>5R
P@(_Z86K3/7AU%1N!GV^7J+EAS=]-!\8LRJ!?I/9A'\5WU.UO<Q4 502Q$U-DZ![1
PA=VP6@:DHN-77,W*O>%R'N5-Y'P5((V_O]9(;=R/-+GT.N0_2TAI1?!3^L>ZOAP(
PXCW]-U1%8H4,I$1MYK+A"-W4QR(:; N1K(;9@,.5_6'2"O''V)'^FQ!MT_GZFMW0
P13^X:[CIB<RK)]?_0N0-CMSHA2&MD%EW_ 7#O&'3.XD6LP1[DH>^2'3=9+=6G=LG
P2J\V.[S7DHD*H=XB_O!-Z<XA=6T]4E7.(_@.[_IL0(K?/< 8^"IS;$K<N,(&F9HV
P$7:S@4#@TJ+B)EE<MBL,+&F[#)KR5 MZKY1'"L-?X:,N;-V-(-%LW8D'3, I;/,4
P6('%]"J59LDVPY%/ETQR25>P4R865?\1LA@T*/RT-49Z#XK"FUA*P:I30/_!:O6B
P?657Q^V72HK).\1W%1.2HQ9_PD$N:'+7<6R6<6@S'=2F71& 9A#(Z(F1:]@X0JA)
P=+ZG!,ZBK&!Z%\4TU(CL4 YH0&NY!>12C"-#'&]KJ-]M)N2C[>SL'6<8ECNO?P1^
PNX%TAH5KD7C2%B4-5X2]F( %?OQ2S0.N+LB4Q6DCT-WX ;4@Y7U)/$?4^\ 758#[
PF+B6R]%.4SG<487C&&HC.JS53LH+O0#^S9'F< "(5G0AVH>!@?XL%E=CBB0RFA"-
PRR5[2B*"QZGNK;O*:;JGD8(@*B*K&@?@5OU0G;O5S>5OR!'J-4Y6'(DEN+MG^XKE
P%(*:CL+*@-*5[&EF[+X[2KKQ7RZG;@2JN6504PK1B69USU45FT *]AY?++NEQ#^[
PFZU\['90<*T(_ .URZOM$1]YP8@4Y0R0FP <=3!,%OO0I;X.>-6-*R5\7H\8UU$-
PV3-$J5T#$3JO)UCK2?'I8^[Z?ON)6 L\#AP9"9;!<!-Q62"E[.12=8)^)+_A7_.6
P#-R3OLU;76/#?"P_LGJ]1YDTW19!B,]IIV7>D4%9-,YW0M1)PMTHR,OAD+$'2!93
P>>@\S@\^8$G2*JS_=,7>6?F<T*EW=$FN:+-#[D'?[5/[:=;92OC?]1!-_Z]HIEUO
P?NZ1$;9G03"L/D1:;7(;:23>C'>P;*="U[%.PJ-UDDY1=EDJJK'[^4LG.BD/*'F&
P[C3.PO/ACQ%(YV)1K%2ENPJA( D4%'X^ '-))X;R._*^6@AA?F8E/S/S:"("W=Z5
PS#%1@M?X(A4?"G ]C:OH N@\IS!P]"[= ^_C)("P)QTD#)L(!R&CXD]D541E1D%$
PB(U3,#W^C)[K]S);#S<[*S&4:UY]%M&,>[H?CD6=B'NQ$9A3[_@>Y=_9KQ8CE*8H
P.(M[VG(9:Y^X:'#IP^_)1_=7Q\>S):5!*Z4G+4H3&(UQNQA:1F]DDSUCS+HLH5=R
P_1 +;1IZZ6T3[L0%[CNY'&MD>/-R#N:OC2;M"9"(<I!RS$:H:C,&/P$MIN3,N Z2
PD.G?NA.XL0B+Q'\B+Y3>>!8FL2%O^1L4_[5S0'I=51FHF4*&?Q(.+>?XP7@H>%S6
P)B!,"=7I)YW]?%4P40]K65N.'5 BU,N\#+;)M8%;WQ#8@8OKW9;3;1D; ,&=\#,R
P7D9VYM2#+ZDT[3\\X/,+]Z0@DW.=@JJ.[9,=;N<.XM-NY1/G#^PE =T'8#QOHQ,1
PNE0TEMCOFM@(GL2?#:RH(_.01(:\A2MO-#"+[4Y31BSK249V807:#JK4I"O9S"9\
P+@HT_!H&W,IPLF/*PH<D>+7JF.7-^WQY2[*;P?'8XUH7WGE[Y'UCQ>]LK+_.%SZU
P^2=]2PC4IEA6GZ%8D07#KNCBSOKZ_V%;6<]<)Z+Q4B0.!\=M;8FM#'^.&UDB)5[:
P*H_3AJ:H-FJ91O".I[E5_CX*IJ9$%X10I)VET1O]@$Y$L)0"355>5'AK3=%RF&#S
P3V4JDPN@=71F3>8ULCZL)OAX 5(R'G^^&G2R*0#D:.\#>?:#(R\>19BH"O)O45FC
P,OZMM\ #E\*;))4IPLGRBL>"<]/*]XLLK>=$\I)#?4L=IWI]P7>!_"NWULP3.;9\
PXF1S(%@Q@'P#3X9(\O\SVXT!9Y"^>R!A]:+>:OR%+&L"GP A%0W'G*)7]#3GF,)_
P\QL?2E-_R-^FV])H,4"X'PRV=:^U"/= ,] RPF5\:$@_R*/PSZ*Z9[I*=QZ6'N:T
PZ=(-84H58'_]Y0L?CE>*&?+PN;+FN7RK1[+-S(%.+LC.*BMWJG#KQ+BA\!,B5"MD
P[W_R,$K,)=N2Y1W!H!@'$#&3X/KH&UD OBE59TXK8UF'ZM5I)&*;L)N)0]-D\%-Z
P3'*=@-- R3S5]$=8@QYOVJP"O#U\>1?;[Y0I[.4)5!YF4VH:BT01[@CO6K'8<,OF
P@SEI&++<_?EN+(,]$@WL$M2U5Z#;["6:I%#4,,;Y0:@6VQ40^6&FYAZ8X9N5?CE+
PC7PX9RH*L=QQ];\Y2&IBW[&5/XB+S"N;\K?LN?@P,0BQQ16]MD_AR.0[")_AMH7+
P#XS7_5R'RU\DP)FZEO6<\?HL;?Z?2=\UAG@Q[@@2BT\F=,>];-AJB3\BV[U @%]?
P.(,($#FD07%.D#E=TIY+8$U[E+79F7PC'60WUTR,'8>:^->8U'!9^^R*W$9Q1D52
P->\%2;N4>4>G_UUAA>4;X_/ZC!4BL9^U<*FK7@0!1CJ<7[7XUFKOM(J+ [ X'V#[
PBJ,5J]:PJY0COW3I-25.4/R5%TZ;VX7^*+@KAN\NBCWE\)"R.4:D/F#8/OHDR"V5
P&B=J#8(;-8K+'!AY&O*[R[&&]6FPNC2&$WA];DP->MXN7H:=.\DMJ= '8)">&TKM
P=)P2XS,CD6=#HT MRPC+U_EX@V0@%'XT;8%WLB^R_VAD)FU['U4?F5U!9(#Z*B %
P^TH$15?!U'4$V>1!)./BQ8(.Z]@ENGD3 G+?HHIIMD_Y9Q _"HV%C@,;HBF2'-Q1
PMQEAJTJS)>)*AAQCXPF.@\Z9AT1?D@K/==6RR3!G,."* SL3<O^VT__^0S$CCE#@
P;GQREC=./&,WQFLQ_@&*];[4^Y:\T5GZ1A^OL#9N]CZ=+40.W/'!:A"S!W@P\( ^
PZ05.&B$B@:<ZK:H6='RP=;3SPYJ D#+?WKT\\0GF7,)>1K3&H]CVVV7G2SV\GQ/*
P67ZW? %K=M=,K/T8WE0SH/(^ZAG6M/\9Z&&3GZ]^"Q<8'%O'LRO0K&)A/-+]N $8
PQX9"*TV)P+!CY@1@3??Y>],..M:HSR=,Q[7\UJRW!X.C$S-)B.>OUV&90CV!JYU]
PA/M\G.)5FK/Y+G'N18*FZ8"2$5$BK1>HZ 92._MFA'WF_PF<$W+3>R+):M.>W"PB
P6@T8TIJFKA\WT!J0N^8&56X=M%&JPP,U#Z!O%KO]81B6EB6!"/6;T\GN83=TPCS_
PS!P/P"NF,Q)T2&6K"&W=-"JC,J2WZHT^OO?ER^6K9J=S(L>N9PQ%,/B$Q0R(48\L
P\-6_A7@"]BH7ZMH2PUN">2QYAUT:DSD^;G0518)MM+8#'1\8K9^NM?G>3*SK0L<+
P+H7W06O4%+D\D8G(O8L_#Z[*P+2"^E\+TO+IP]!8Z<P*0>W"2+:D =8#O?'S-M\8
PJ[)1P46+06+3*!(P(7]-/EN=3N8A3O*.:_;2,?2=YXFZYE1F]M945O^!.O0<=_PV
P0GNHK.\L#Q1ES8OV&.^8M2C_*CH#!/LN#*X&3H9W8KQ\L7F=#<;1<2QRJT&Q9J @
P$UG] 7,B[6?"OR3=E[\:"_JXLW0)14]NRWM"ZK80:@K/%<>B3?:N4A38T$#X*@R1
P<YMJ47Q,WYB)];I\0HN;]:N/Z74T/!RIS2[GJOJ3E9W-X0AS*,/QU7R"QP6AJX(D
P!8<DC:!X=/AUZW]UQ((\6;.0EU:WO, RT%-)<5LX'(*HD8]O?NVG^Q,#B(? 0 4.
PH.@'U/FL7_MTJIB_2?[L![BM6IKF,9F*3!*DG5,&<SU)$>K_8-V^.%@<R5;/\ (A
P6;,$'N*%Y9DCRC>@V\*;."^_E Q]?<%,V^#</D3S&0K0A.[\Y6$C>YC3D9 #)?/,
P^_(*HN]T>BSM(8-W8SD%(1KNAFSV'W"1;96NV*36P/GT"*(Y"/0W6:F-<TT=,4EZ
PZ?&K9@S%)# 6[1/T ?X082!J2 I$+(CZ=GJK64MG]^^($JPFN3[4P=K*W"CA9, @
P^?"R#O*;JH\X''^ZF]EEDSE]6PUKM'-&E(+*Q(/PD$LYL<P<#S!IJHO% L5$-(8I
P\Q6VNMY9I),_;K,2V3!U&3F0:EB&@<E663YG_<O 9HF*G<ZAW]\%3?+Q];&ERUHE
P"2(2^$_R.(^E++?S4BGX>N,A&%DD[5ZEWC86)SW?ZE\\NF@](GBO54)[Q]8(( #!
P 4 P@^N#@CZ0X<P'@[[V2YDYY*E)72$9B&&:UU&-TA?*;$CU.E0UMK8<MZZ]O7*%
PGVO#NY@"8S%,<%E[> 1U'M>W[./D?M0I9+-%;LQ>V,L[,]:VQ7#N[?K):=,<=C\!
P("R_)I<-#87&-JYY+!IA,))X<8D;WAX^2V'%>  !W14ZFTO+.:U!HD]?X&1>!NF1
P_I4JV8(&0!(^A'.KQR=I!<V%=GY[WX_8"A][B<B6E4NM:UHV%P5::RCH%YM8J.JG
PDRL*7[L4-?_@<T9YO+R*Z*36S;IE8I,VT$(L5YIV##G;\41K3-UDR%1GC3H5:?;(
P\?ZA[1)OS%BQK'/H$U8\!B3DEK'EU)"]D\EG>*0.PJL:]0\'.@!'0X,[TDS-U)$,
P,./;HBJ,NUB4H<=M=@+OF:4+\>!* F8H_5U8N=])8;)C=(>Y5"[86:I:C:9;>9WO
P-GO-BR:A.7&"JC*&L),T,&Z))QAA9&FTLE\R/5)10DT)"URLO^!+KD7M!O,,%G'9
P@+"'S)X&Y,WJ%6R"Z@!MS4+YM!MMN"$=U#\!5P262Y2J+L$1"'/IQ:LM!)?@/X]P
PW.M2 *S?_RY@"DNC9L]:;:=0G0 D2( 9V*^>$7?GD0=*A-&':SW^0147?:LS:-'1
PLV8($B[U$6CW,Z!T?X6$N*VZ54XG"(>.?UP:VKD-6<Y+43C+Z7,IVU8%<ND>]/VM
P.[HV- @+'.^YU<#_2)0/26F 9O? <TD\@3T^/P'IDELJ@<=C]$"XI^#7R< L8[?)
P60NHX\A<IL)73BU3)J]BT./H.;?V]'A_B).&7),V8LR//;H)-_*0SM<41W@H99NK
PA^5/+BVS4?SI[L;;GH#;I)3![.@.""PY8%WJ#Y#=;FSX3/]YGNII6W:>W8@P@IO?
PNV?C_1<*P'Q4>DBND>H3,FXRX&7J@PI(U+W@YSN*,;RUL=!X:\DKO3_Q^^+]@C?9
P\BE!:V.J!]4K.+E,=WL:[NXX7&-2)?E].>7^J[<,2A_M%MK/OOE06$:?,Y)S[5H)
PFZ _IR?^O"9MXK2@)[!N:0QMPD=&N,Z^>M%R>G+DVG"R6 TW?/E.W'_<;N.;RZI:
P^9SH16JA7_8JIO<YK,__;\X=7=\6FA'G"0R1-YG"DD6 8C[%UK1916KIS1*Y>0B.
P@+KZM6ZPS)'W^"PKV.IBVM4H%NTH$A/@TP[ ]=@?O"4K#8KM[Y^KBK/=\&]-+W-+
PL?D8>W6!Z,GM3JM6MHQWYI9>BN7]'U=IC\=TGBV/NNPYZ:L*WK]Q/9I[=56RK_) 
P5O^E?.+%8)M>W7/A_T,6%[*W3U9;T)PX@7J^MHH2TM FVRIM^8E(%&RAVGZ:UW05
PD\,=HMGS?J(@-@?@:1O9S6EU(-Z5S0N9VVI$$TLFN#<_YCT;]54 ?'7@[,)W<4QO
P%Y*YO'OSN>&^]MB)[EX_U2O"1V"/8;ICVUQ@F[V97_#=1[BF[%^GI 22M"]Q/CCA
P?(L-XDBXL]+J,-<DLR;.L<;N]1SQMY.U2YH3A$JOM%D4BR&$XM<C'NJLFSC\%[M$
PPF?N[_!;7Y)X83V]@KJ]/#; "/(1DJJE)FT(Z4'?JAD=G>M%W#<QPY3:T-!K-:IT
P&E9@&BP8"V&)'AD.\!/P\;U9Z0O/#JA"37HZ7)!:Y<W$SIK;$_A]U-485WI@&%"/
P@!+X7^TY(G2;,BUY[: &^F"C5< Q_PU@?OEY"B:"7")9/=$BU[_I<Y7?FH'SC@4S
PYTE^8/%(IJOUC9YQ\*#&GNBL.KF04Z:M9 >A?>6C+!1HU2OFJ.&\$RU\J[X3U?/_
PR[3K[<(KV VL32;QE-N&VIY]YY.@1Y_[4X_N$W<AF+^PO$PFYJ[JKHS_BV1\,HNV
P19,-I[K=,>"<M&'OD\L;KA(!A]*N8V](NG'93SL?SE<0>-)":R[0I>#\SE:,O63S
P==@NU6J<7;(3]F3-2J8>5L;%Z$=.!/Q;Q?PFL(+I1/G9/F158JJNM(J\/][OE$7U
P#K?XO#A6G5YYNU33[2&A>=2ZP^Y,.T6ST4L=?GOQN?L)BIU<#!#+"L'&MLATK>2)
P\U.CQ4Q_,R<5>)L@C>"V(NVY^]Z&:)HS8M2NL/F:"JN\=G!E>3=@T;KSAR1Y#LVJ
P4Z[!XU>=$RJGN7QN=\#/#5A=_[["KX_O/2CX$%>;6]'?"AJ"("L? J^S2A_+-JLJ
PF/J-"'\4CU)L85:I<-!*F9P5B\P1+&8EQG3+S7O8H-NKA36#./*_&+.'PP,3_%L<
P.'RTKZ4M^:W!_]T:ZL*KH%<,OHD.WTV<TP=N'F%+F'9[:^7K(A&$,-V*LJ:\<S C
PZL1J:Z%WSPI<06Z V',9=OV]7TG-F[)I@73Y)'1",&J2GN7..DYKW0,AY.UHJX^/
PPKJ&RF)YL/5K__(;)D>O:Q<116_I9*2.3R.(QY^MUW+O2#P*.[N(J_?:<-O(L(02
P+:M!+'O&<H6PQ^KR/J9J8S0QL]IYJGV-.*8^I;.#&#ZY:FV P_Y""DS 3MD2,/L=
PZ(?C>(3T7HD#Q%[?MGB( H",H=":)@-!G:%75P[I_VFFA/W.LSPC$-3_(K!YVZT=
PLM[R+S03XX-&)XL"3@2;MJC0N\LP2#\=R"Z.V?8EE6F!5BOT"R^MF^49E 2MSWCQ
P>\LTOW/U*J>:&70?_!;#:--'9$V+?TN*!-S"_<[!:QH#F3)ACI,7Q'#$"/\P]*JY
P/](=N2Z=AZ=^]!.@>$DB>)7']87H$_L^= .P);U) I7?I.DSLJS3756C7[#!FVK#
P;V8PKR.6I>,@DF5P#PNX20MNFGSP%CT\2DY"R=+%<5-C=(N#V#K4P5A"+1C$X--"
P\W,YWV0%ZXER@FBUTL:7Y&B7&.*+PL0K>R[_-Q51Z, 2*WR8U!@I3^+NT.[4^@Z7
P;LZE H9X$/-; K%F2<[F,8"2VXO>&C\9AVL'V*Y_Y3Z<2AB^?F([*(*='A2Y@6<G
P&&0:XRZ4U*LS#>MA+]JZT$V!I08#[GFL?/]N#&PSTS=M2+IW]-:BKO@H7 'A"R>Y
P:M<D[#&\@QL"UL!:CZQG@GD)^UK%GR$I^)"KGX#6_5=(/OT2,?S#R+80*3Z;D==1
PT%J31K68+VEJ-1CHX!?IY'@&BL!R)C\HM'V1?D?M 3/;R,PU&)]E'O%ON.R"X5BU
PI;%<1L.0I^A@'QH#7]1KX3R;/2,BT@9U/&-W:SF@!(?B@OVN:%5OV]PP^^V<V#UQ
P&1P2GTM"#$!F%AO9M/$3YS4B23?>042^)-L(AEI/X J-LA)SF>39E]HF[#.^YGFB
PJ)-P00M=Q.=N*9J,Q,'0LO3[],2!XQ58,U;Z8V2&6@U1)>1V\U'=B+P&TWR#@5QF
P",S@9\3[H\"4%;$]F^";AUN)(Z/Z=>_D&4,BG$L<,D4/>/]I;@K9) WE>-C;F%3+
PND3M&^^%V)GNP%%GO3I*-)=?5:4.*X&Y^*2=+ #S*'*Q<0;&?,0_XLR8 42KANH:
PM9#)3]$87[ZI84^J.G43F,UV-MA9%H8=N!!L/,/ON.S]KC!F5#(ZU,?#.)^,60^P
P4;"9<1N5?H;*2$BA38P_BQ7I3R/)U5P"A.F[WZ4<GYG=NZ)Q-FSCHBU^\4$K=RP%
P<_F>1#KC3&A57YR=E>>I3=D5/W&%]??-;>>"OZ..#R"*((IJ+FM>CFS=7"9ETWA$
PV\?AK[RB'X9?)-C=:BDWH,=VK8!YZ$]@)]"4;6+=*  4-QEO72^FYAW+4;R[8# Z
P7,H]A2'R4N)$^5T @0>?X.,8F=5'D#6WY"5WAO?[\(2()$ Q@Q#!(T?/9G:HO<;4
P<.(6\=1OY*/DMEO<K*%_J\/*L4V:M<)X1<I MI/C\$[P2(\G,(9Y8BV*4K8HDH4H
P<HZY9_A[]&_TH8RO;TMKXNH6G[+M8S&PR83NI\EL*H:*" <;W4FW5E>U(VBH'#H8
P!Q*3/KX7:#_(ZPN_9[6.[3Y0(#^P,^N\T$IK1I>E+IS=-.J<*X*09!//?AQ?V>ZI
PP:7YP9MXN*?[3M1PK-AP6G8W]3UP1J,=H8&3;Q*65OG$,N<X"X##3Q9I4VOGNY4%
P@[%.);!72Z/VVWQB6/@.9J0CO/3#OLW 7).6-_E/B\.FJ*B0"00P^CTF#D+L:VZW
PV'2*Z--46S!\0!:N9S0+U$*6+G<T14[T5H-$)+YN04H1E?H,UZ</S)[Q+TX0#* L
P'Q107R5IA$0RF4G<A<]JRMW<$O=)N0^M=?B3Z.@JOR/"[<)>7,Y^#I/RYC5!$K-5
P3@JJ'K)[M;V0W_EVB, [&%"N.&*V"0Y?C?[_^8=,,)Z'V0=?_UB5-2>G]GA@;U!9
P'8$PWQ.<TF&O\#P%^F9*225 W:W?NP_.$:JZB717CIW/BWH07VSK"+"D]?GM,P8J
PJ)(KY7MFB31N996J"&X)R5Y T_B+61$B#%:C^CC[G,"B/[TP!O:8*;CP:P7*O$<*
PA2^.?,5Y=.DDXRIO1Z;8+:&;,XA+V8T#&U^](*-[Z5-YX06<=Z4LQ*F/VCNLV*&6
P3FO92OJK$94:!-MDI#7=';VGX0;3?/<+\EB$,JXHE6.3Z8/L T2].GDC7!>Y&[GO
PW4!QTL.4&YW\-#)Z3GUFK,P-?9S-1NW8$TZ/_$W?5K,Z1NW^&:_+XEGAWJ)D>_ND
P@Z;[#U2G5*7H#S/ITW_3_=V.VC(#"ZI)I5I06/IO?JMM3PQ-U/YH]J!6FG-:P?K$
PG,X<>7)L>H1B3$78S<8SO9[_YR(^DN#B=M:%N'HIVF^OZ-;K *T<"4V4^5ZS G[H
PVZ57'Y_(M,@+ ;L;%VZ/N @K3M)%_8(<8 ME]Z@Q"8(#'D<)Z9R:8N,\%]+#Z8$8
P?JZB)RMD![TF+/E^1F"\1[2B,%WCKNYGB$LS3PZ>P]A-_;+&>X9??<?A_BZW>"JN
PMU48:/DIO-F_42$!!\#?7057'><D)3:64S^&?D.W".S#</],*VF4$14B!$6Y/SX#
P38DDH3B4A\0WILX'\'=9ZZ?UD^'> ,LZ-DR7=X+H##ACZEBZ#\)TH70C[0Y.I-G;
PN17WU>&Z/#'?^/)*@4C@\5+?(;GYAB^GM@+=6J&LR)&P3P2UUX[S6P.E.5J:S50[
P\*53=-\]K 3H2#70&B+<,\LNZ#N)\+KZ@@]7"8<.1G9?>?0ZRDP!3YEP@R]Z?U4F
PSQ+OI!W (.B_(/"=Q$'WO28A_J'-GP!P;\\_7?+O8;C2J"C6^'6CC1M2QF.4?=& 
PP_-?G<AJL@GAR.P\\YV> D3!?C#J;X@3"S'QK?9KZ]T8? (ZNT-LVB(GP3XC:]A6
P80BWTZJ0\,P'^]+QXZ0@LI1S*\!\PCY_L,^D)IYF//.,B#E\]\$A:6>0.6Y6<N]1
P\8,;RXK[55^FV?8\I"^ (/K\0A@<;!7H..P%/"Z9?S&9]<?Y/D\^28"0BWJ\5('F
P7>6PH"E "3.VFU"3N(!0($EL[N]_P"R@]"P*S(PX\8U%)]+&S$) D:W_G[^E(K-)
PLV"Z_"1D8 &(_Y.K1:I*C4&-H;J2MK=J8U^#K)@V,0=QAM3(J1<MX^DY6CN#0$OR
P!Y4GOB97I,+.*$_29_'LYS-5"7Z$2Y;CEN7U+@_Q\7*< *5Q3\"3DE+V<!B*VDZ_
PW!59\K2C+G_*[132>FK<()XR#YG/FDU6;;A.BC#F"-Y)6[53$%S]Q)T7-TH[\M/.
P3QVGB3M[7<A?:H_[F)BZ#Y'0%[B"]DM9)$JG08O1Q?F-[+G-+9ZB^IG^5 DNT08P
P!F*]VF@NTD[AA5"_AM#&Y3OP_(T7R1"!Y763T'(O'QFZXV>-IZVUH;JG3]N* S<A
P$3^TRW.C:%MH7F"^"('(">(KLS#.%14O&?Q/SJF.^Y?8<7Q<:\Z5NUJ*S4LU:C1/
PN$XB=5B5H?B%38D[*4SQ>%=0I%3@K[W[6!33ZXTKJMJLYD^+TUF?T!>-2Z 2LIZM
P.!=T6)<L2)O;8[Y^C]KR R-"TX3MEX+8C4#_;&1+./;LG+V/R9VULQ9M(3Z^%%T=
P.G]CM3UE**>SWS<CS94-<X=4\<>?+%K[!4G2HC5ZQ<3^@4D$0<#R(\(9JIB5%H:I
PDHS.YUCB@!\<0>%;(NU6/WDV%*?N?H$GUUL]DKX=%"<VMZ'BGPK&!8>5+BWHK(KR
P@;HMI(LJU3C2FSH8ILZ3(6YXY2LP1=MGI%'D9UU*""*OYBH2-+)^W:\U,4ZN,D4]
P"7'>K#3V-YS;N M20LWHHM665 FLRZ&%DACF2HD5&\BXL3QX&)F4028\\X( R$0W
P/WAK%?E!#2=KE3"XF&GZ6/.$,SOC5<[LA(P#B.N#@GV^6-3.SH-JL4C"^>!&391T
PB;O0FJW[$O+@/=WS7#B"JS9__CZD: M=S1Y7W?/V>1:4%H##M_C%JEGA^VR8N<>>
P"VO57.K^+#;'B@\]]25DXP487."HP_((MZD(]Z>KP@8QLA(Q\/ZN1L]#(W0AP%I9
P-S+0(9DBHQ[]UAPN*N=/9A[H/: ^8>>JFHUPG"P+;4)I@*TEC/J5.HNL"N]"=(!!
PEQ5%ZHG$G@\@P,,[D:RNN"7^W1S%=(,(J<CQXJ.S6FV]+595;*M?Q5&FGO5$V6@5
PW5,@ZY'\XTKS5,AI1@/5@19ZTU/_!=SA*E\4*@(5RK*$,XVWOY&"-HFO/^P$E\;C
P[<A)."/GQ-1$=]_>5C\=QHXWV/ ^.&];WJ&[K5@ZSX\:$Y\8.=6Z%5L8#4 7Q4A0
P]^[-F8I[%!++18[3%UWS7RXU6$$U W^)E3(PGW:M.JVOMHR)*%5'JIW02#TM,5.*
P][.#H<ME'*!V1?^/ZRUD\-BA07#%/;?Z^D</6W<P8Z]C\=(+9^"9]R&O$?+06NZ_
P[&&8ZMJ16Q33.), =0<3< .E=]IU4?!L1K23W^SYB9<AF]R[FR^MI44'LCLR=DTI
P+W7-+$H)!#4J/][*2?S<U2MY,2FIH8'D\4J')A$_C30*)V18;\6LG)\=L(G*S:H;
PMBL [G:F8:I:>STHLVS\<;PO/*_+*$#0*QU6DCZ*H#I<<MN+C9E^7$&PULD*324B
P>=Y(S@<47EQF$'K4XIB'3YMT,'5SR/ A TLQ@B6 AR3.;:9\9X,EACTKD1-+^SU+
PC(AA]Z@K\PE4PC?E76BOGH0+UK5>#0VKSLRH'-P(JYOB6)3>"AJ 8CTX!<Z(P6(W
PEO+8"E&#5C0B3#7=]JS-:5Y_(C1/U3/%V"(T5X?(3E.EUPLPQTB$&PE^JK0&>PZ0
P]#Q,S]WA:%)).CI=S<+I[+%=P@PE);ACW]9#@VPW+^V2@Y#NJ29L,W75I+ON5!-H
PH=]?,<_7UK1\"-?\5%?;^^TBP(WZ'$AAILXI0:$[.$!N%1Y> WIAC@\^GFV%C(IR
PRZS/L,/MIS=WR9352,\'-=K, 1KO0\I"DVGRW[:Z7>_0=M*?K?Z7".SQ".4%E5TM
PT"H3+^D\5[D6V M)I9FW+X<E%V=)!'K;Z95;*7Z3Z,4<VN*CT5&AI4-K@_"A!N(!
P*X=L5I&=]CU.M7<-*!H8.1IBU([(H\RM<,S$^2(>*P5-!L;JZN$*U*V[ZF59WI3<
P+[WE SIPW&SU(#::H9[QPGC!!S*NN*><<O0G9)0YU-G[-KZ[2<V'73()JV%__2,I
PP7GAR;P#K*'JN?[HVF[7PE$.FP\PC#AT:.PNSF:[6QP:E$0AGZH)/W=RR$M(7RE\
P@II9VH,CGVZCMOB .B4>24!5$/6\0Q7!J#E@,L=N682H;U6PGW6EK:TXPE[*0=$W
PSAJP<PW2!BW^95N(\GPB.(QA>Y'98@JRJ%Y$.B*<Q\S-J>\I\#4<I2K).UUY6%&D
P*M)["1"4H/$(&6'U^1Y-V?O%GIDIBX!V(=J"WG;<$G&3'#P5W3]6W= P%GU8UJ(+
PVV!G^6K(5,'(_@X8_'"#^R@"*ZM:7'FOKE">XD>["&?IGBX[?I<T""Y70G=BM%P"
P]J7ZNQ4?V49C5QM'\BC>U7&^0)H'/ );6^J7K/X8,50*@'3=]3#^^JW/EH!D.Y,\
P0(_@??P(#TW1UTSAK#B"'S)T>>8/N=MU(<_EAJJD%LE^\NI01EI7TLB_:V&Q@RK]
P8C-?(1\,PI%0-GIV#RI,#6/1CM(=-@)P9=VZ>M,<< '8UQM 2: 27&8., <IHWW:
PM3H*-0#,O$85+^@2U?$H]EGL-<G(XCJT+#&DE2O9].F[P>]9Q,OO6%KSB7%0H8PJ
P[=F1E2AK6_PWK%7P-&%PNZ,!3-BOEY2F\XSBH'^R_<X(80,D16H.RUJ\?E)/8_F?
P!4^/$W-Z3B5%V1333%&78Y4$VVU<*QOCC0'8#<@GU!3DUP\N;S5PN1?!1?VBVAY,
P"% Q$4[RN'HGL.4UO5V,XJC_"#-BL$B6PUMW/\\RSX:"*X\-#F//1]V-J\?@YU,-
PL1RU> VDPY;GQ+V_:&/N;>RG.,*CB!\?WD&64#5VC4X+]"&TB<.,_%T5@<\:9,9Y
PW,VXCMU1."+S"3D=.3](MG1M];/X?X<J3[PNS!#;+WX-4;--5NT[T>-46HR@.!!N
PNE0AT.7 YSZF2S(;_0ND+=@DZYM-^I<NS]?+75@W VKRH9%!SA"L^]57J'6LK_Z'
PO*YL.\VLW59UW)>(8PE.>RB;C=&B;$EVT!AB;$1>$)*Y1(D2WA"23 U;5U9-QZI3
P7TV A>W#T%21#U(#D04TE;C7&1N&<8+"'ZC9U5I.+*ZN?" H1J)/'XL:8,H:4RK 
PF,QL6WO#BI9!W.,M'+A<SZ//-C-.LVG\BS3H&@R5C65AL/(--EY/AQ'A(>CKHR0_
P$<B&MWS7SU [*>KN"VIV[G.R-7!Y+=A0I"66M+^3)DJ>(ITN_!?.^$Q+H$[+:T;(
P?%$T_ZW(@R*4D8]&PO4-<7Y)W][U5:S>I_BM[7//';X@%ZF=2,0$$31JN>MHWI73
P^"@ 3!(X2,*P,CF#&/U15PYEPJ H+75G ?B$ @PT"BM2"&E8(X2]B]$Z?80L^"8Z
P#(S>'X8(F#<.]OP9O4;7R:O]$T+-XF6"F#!0\_N%7MDPBG@.!JK$T:W'.?6[CN9'
PQ2< G31$@.2/:^7\'G>NA.0%PV:J%*I:G$#*"%AIN$XH?@+U,S_M"+M@E5#!+PU"
PQ0L:3(_! \:5,5W0C1.J).W_ZROK;<7)-.J#&<8Y5]CR6*@EZXM'G9,&23^')85G
PI/Y"31KS&W9_=SC6\J/ W8ZN)K"<'.0S-]$HJL=Q0GXH@D%<)Q'/3"RU1-9L(OP)
P\LZWT%\#O$H5$6[5[,@4CYFUS4'@4*7)2>!?^AK!DSUPX @1:C=0!.^TU4L>N'PV
P KDS4??H-$'EF:.;X<F'4YAC3N:<M]Q9!XF7H&C0^^I%'1#1 ;KF)$M"/!S^BOO(
PG(+_:I.KB_Z:[0('@@+WS<$)M;IQ\XG2_.Y[>&Y\"">6(3,8E@;>Q'F@_O9'F2[>
P D,3I=E9$)H@(R\(DAV37KPZN/FRE!533G3Z%A,+B:508U14C)^ $3SR>:N4S-M-
PO(G*GHHGE5&;L 1N511\#F1H*XLLZ(W1+0:=_Y5<JP6)FK]^C9D']N.+2R!]E>[,
P>FR=G;_V9(:"T$M3-50H,%N)XP5K.\\'I(?+#LMYA4MD(_JVF.:U_4^*I[T1 CQ1
P$IL/[S><>5\MREB7PRV'?=K9AFLUO;$1)M+O*1LSXMK]B&<N8 ^K%>]H]D,C"/BK
P*I(M(_T)VH_3!W*"72($<R4Q*9HUFL%=<%HJ%G#5I_[,0Z)'M%Y5Z>%J#?<_<MTW
P\UBA.5=BN1N*#KS9O8OZ)X\_&#NHTZIO&12EU)#&RO/=;PQ+Z%(66GC&^)XH8D)+
P@VPP.OI<\<0FI)5J.M'WS31V&J'TE >WM/%CX2I2;L_5,AP--8C2?W/%-T_=]UDD
P>%C+R&OD=\_ZVDE8KS*RI:N-[/#+5S=D>/8 B"M(<#']L'%?-3X1NNA!5P4WX\)L
P>VG4O<$'1-/#&KID:+,J%#,<%OU>7^_G-<K3:3?G D7\H1^SWUANB/=R X$[3]0H
P\[U$*$YX.*:=0MG/6(3P<7N%&%O*[[5_%JCL_CSC'L^5<%2R.T"EV.>Q]@1=W^YB
P F@6Z* 6S+EOVE*ZPAX*B][1CA%2?"C<JDV@]ESH@WR5%'%HUAA\9!0'MG30J$'8
PSDKYP?VPD@2E!6_&R#H5_"RUO7_?,#HW.X@!_3FXBA-BO!0L63G-3)H6@_,BVO6<
P!#P&-ECB])(?+[B[N&'D0#:P+9,^#H#T@@LQ@%)'"2/!FXTT^E(_)AZ&>UC2>3%Z
P08C8V[=!2*&K&SSFYX#2$J*3'EH.N*36CT8I> C#2?0YDO90>4RWI;$_)92L4Y.?
PRP&G[LSW2['^[MLI@EBU:%SY%9"I'K!+:N^MTME1<*?]IRV=:?0>R2!S0J7B7^LG
P _@-OI&Q0&3!@X8Z$ ;0]NW-B5$;I2$%B$7KD5%IR6SM.6X#\H4:ZW;V ,0%1:K.
P1Z",@@4SJR5:;E%E>IFS+*?Y?[MZ1MT$Q,JOP@F."_7IE5<;$ Y"-DJ7.OCF4E<$
PI_LP>RV6YT]4L38?PE)<T4"%;)O]J2Z3< BPVH55>^L[JNP,IOO1[-[%91D&YM;]
PIT?44AKHVB9)5-4&2DO31R\8(5VY^0$0TELS,[R?HZM,YB\/)DW[]Y[IOK[3&V 0
P:7N;M.,(1'>-S(M=)4%NEX*@X6Q_H'"4$[AA+B"@->QIZ[$06!-@/2NO-!T?7-.T
PRZ!JA#F:IL'J]"E9NP\5+_>MF-A>WM 1N475%3JD"4H[FU9E,:]\!D5HNU3V:(Z#
P/$Z[J*,W,^W5G9Z8S!/N_(RSWBK[RCC^ITF<^O6O%"+\J\Z,B+AF3NHJ( TF>D 3
P1?V"L/B4O-68H[OXXS>_ _&4,(MO1.1P+6($8.$V$<(6*ZWR03N(["9OO%G@'5[8
PI6*H)*X%_AEB3^!\OUXP8%7(Q)*"[.D%(=9T)MO7<*(76B'JH-,?!E/VF_-DX+7N
P.J>H"A8Y5^"?]'S_)29,J@R1;Z<U/!K(73$=4W3Y?E<;F@@Q?=2]E/3>5,7P]2LE
P=-[R70$:^\T(+'![X^MHK!\:[:]I9%=A!5R)50E"PLTNF-$ZC-0&"!9J^"^=@ETD
P#J?V.-=WQHC1L79( B.ZS?H5OD1*EBM9S^XJ6].1Y$],2L,M5HES-=/=0C'/*Y0K
P2D20/(X[:^LM<WRJAK!A^"O]L4&U#B710,\$I*LEJ[0-R4W>T_\J>8B'%\L6 56T
P=7=$A#8>'TN'.YD4B@&]& < @_GPKN60#2)6[ =,%/ C+31[O$!/1O>$;O)7^M6!
P3(61M@9BF=JU[*ZF;\5+!@W5I3H$1U'/P\-TEOPXF+:?]OU \D(LR>\Q%!3D2JV>
P(>\F4VLHX44TWF[[\:7O.,IBO>V>#@A )TB(#&Q';^60S9N68/Z2]#>7G\=_-$>"
PV"#2$W 5V/WF[F-W(PH8 I-+<02 U#5,DO$$?Q0<AWNW5FMNYD#/6<CS/.Z=8^)X
P:.]&AO/T,:1?AM EF;1$<C4<CKR5V*3X:=K=;M6^)+"+G<AT=R:9KTRS=PMP];U_
PC9TR.,(8[P9-&PN;M'!M?_YU/-N(NZAT+)4.27NR$OHH-PA0/M0@Z#33H=B G$4>
PT8$_Q7EVWAL]Q4HNIA!U#9U1^WPS X'^QGUT-%*,X22&=#MXO?H+(#6EO!7$Y:85
P?VDW52*YY4!N>.;[>$*'@\?>3B/#Y*)G4#58N%L[FRG,%GE- <9]C;_B^DYG8FG]
PNP>.4@:"*VCX*F,$YY.'ARJ_^;SP=&IRM_#ROFI/B5KDOJT,%/?R&Z\XJC)43<MH
P@-3IM?+N:03NU&X<!,I?[OD-X:.,0_FEYZFDOT'7O#=01'&$#4!U2J&#6=,:VEL*
P39PF"GKN[>Z*] LSBGB)>8?CFD'OTI0Z9A>UW"8Y<M!PN$)Y\;F 3( RQF8@^8T1
PQL0\P!:\BJS_;IH;@K77P?L-H=SD9]\Y@2-G&[A1R!;?+26&!O:Q(N"-P0 &ET^$
P1[$XL5WTA" &KSC;7"[2L=V0A:KD[[59_XK4X-5[^<D'G=/&WCQ71GG#?9A3&@P(
P3O_JPUMDT(.=4>?*H>A(AH"W::U)%:3D@J3+P<L$-2@DM?^'Y\%JD1_ 0 #G<)[6
P@3-H08 >9ZQ^D0)K^ =&?8U?Q:7<JK>H$KC@2_PE^"7-QLPS.2'CUUB[#T(!V U*
P54&E2L%V%4%R./7!:0"5<>18RJ0#='!13[3F=Y1>N7>9Q!-OFO'-GN=4GE[C#.+"
P=3Q>+C+AA<V-X)+K_DZ?<W=OLVRU::9-L?=!"[?ZTZ^KBMS'9;[334O:%[AJ25.8
PNK&GS7L0,=^:F<XQVOS3TM>EI@SC"]][V>QDK8AY)@&&?#R.4""'OS^2MT-<EUD.
P;@$E$P>\Z*G9-0JYYIUXSY67Z7UZ0"<A_3LY'>@:[%,CH@B6=RG.I ":SE <F+RB
P<6Y*LP@*SE!AGD_.8@5"WE?I7S=EU'^97N.=EWH;F)F1C;QYYWH$Z[SY$/U2\L0A
PL;%L\B4Y(GMI6-2@D@1"#X)5\KE9'"..K@'D]+1G'^0102);O2LR5Q*4_@):;]@>
P+"):5\VQHXX&X0L^6(\NV)<'%TPW 6Z*2$8H]>LURX')'LB[PYNT: ,FK+IGZB3/
PL+TN/)-FYQ;G@3'T7!4E=W),@VZLG?((BN?E] W\]+-M+X(NFGH#4LG0V[)E"D4<
PO2X3TJE.F%^:DM- %>QOIPY/6?>+D?+3!X SNF##49Z@>Y+DX.N6ED0N/1VA_#6V
P'3*J()T:2IE%NLWMW,K;M,VV:-=0"9,LO>]8_5BUR#@0Y6@&E2:%@%T1!,WX$0MA
P 64<VCE3\V0%1XJ/F(A0Y;!^SSMLK85A=$"W05KHBO#(#5'67OWL:6&Q&]&Y+Q/G
P*[PV!B&29EC*M3P&X6%6(M3VYDQ&']1%N'98;XJ^RN<'#9^_BO:10M$@*..Z@=JV
P[/6RWQG#1]PZQ&D#CQE,J=0V;[5#.Q#MFB+].<(OVO'A0'_XLN.]OE)J+@S8L-8!
P1,%KILX#QR(/HU/+V 4,!!CC4.%5.LSYA.C8:J#_7HSD1-';GGV/2A.R*0SI3EU+
PH"V!8FX8QE*7&WAOIJA2OXP+HFB:-K=5";]<O.)+#[:_Y6;E31]YS+!G,#*_Y846
PB=6@KAS?)R;VO7ZT;$-I!*PB_*^WL\,;_+4A0UCNK3V,X8+@3F4AJP:\*M:B"7VM
P4(P0!'>G_&;FNWIW0JS^$8D.303FIA<D:/F&HG$^YT'!\-&^A4P!\6LH!W"H+)']
PL",ZKUZG2JAFI^X!JO0WI&*S+1L@!G).(SKN;U595.0A'S"(FQQ"KC[_Q?>#E[_&
P]UT86: Q(Z=6&VRIN%YYT+<GN=/M;1\VQJLNKL+B5U:E^_K;0*O??<>AOI>@RJ,3
P,Y=?R^>7]XYPH]1C+G4*9GP;@9 ZKH4.A0ZH/NT+=<BE0,P<K?+_.'6Y5)0X'8A3
P4F@^'4\*#L@]6 0R$%S ]VQJ$!VD,&PAI043M^.8JU9=9E J=LYF,YE"B# 8S'14
P^6+YR![K;RV$?CTZX#+,'!/_C6?'GZ!6 OAA]RH"GZV!*+7Z9H5>L:+/2EM0RS4Q
P79J]8</LE?!#7_GJ*3TY(F-266:,Y>"<UB;#MQH!^H=7FN'?X#=D-O%K8N<64/X0
P6&?G\X+H$C$:"L+M.B\T E+G$$K61*\8VLFG;@EJPP' ((!CX+L\"0;#>V'SGWYF
P8,7JU"DR_A*G.;@)D_(Z54T5O ?^H$ >AI)G6#"*!P<8J;#;'%?K<9N(V&MCKQ)!
P&8#=.QXK" 32CPYQQ+!,\S)%&Y.(KP YG 7I54#WZNJGT<V+7NB;A*Y0![HLBT6L
P(XWQ9UPE:T@P:P&$:.Q;/&I I6]9H9U%O];$=YO,"HZ5/9SE2:\V]T9V1[.R59FF
P%_HTCTKLZM(DD1L5!P5TB\H!^$2&CZY)Z>%A!ZZU;@")UA%C.C\)6@U+D@+W$14:
P<H+N3N9#A:S:N#[K<*KDG%\FC^3;?__?>9$.E'_"?)EK]%"P2X( O226L.!M*-8P
PM&):KN<13M6#9)@)L=#=%$:'^NV')KOP0UWRF>!IAJ]#TN-LJ&]O,73:YS^%RH>[
PX^C2?UM&2?#6[ KNP]X @4<ACZ/RR7[R++@AK6BAL#^)?H,D5O;CZ?7>%OX].UY$
P?!AV54>]I&ZK,?0BP_!B<Q\ID8G>)R9D^/+O,K<H86L^QV?,,QQ5$-.T1YF#*2VK
PFXPM4;4JOSF*\V]_/"HD=_#1DMCQIJEV":/@HT/"FRLW[#NK?1/*!.&.0BPHK&:F
P<#FE'E_HPH4J:RBL0.^\]*&NG"LV)KR+(^CU2SSB;!8LU=;#6(-DS*GVS[^+BY,/
P#EZS,6'VTJB$/T%-%'8DUD+$"QF#GRKO:\)KNX3A7''_%XBQ0Y2IX=J%[F.-TF<$
P=Z<3CJ]?H&B=+*PP70I:\>6C"8/N/_+HT9M.#DCF/F50,:7G%=S?F#*96WE#,9]E
PLZREFZ:'UEPZ9I@ET'"59?.;V4^4A\E^33.,XQG9ZJ<YF<<1!YL.O@O4\F9;M]VS
P=/&]ZF)YY"L>5LR3<D*]R"S#N>C?XZ*0W K0NV6Q34/Q+$\&%^8O]+ 4[U]"F.R-
P7OIR=L X[5<_?\#+U"TY5],+4+<4$Z )_8H';0-<Z\MHXTEM679N-__6=S".(]F2
PS'0:^;ES\7GHPG-E+8VFZ%$3=0#SGLW;(_NAZ >MD<'NO6(O.!Y*,:EA%Q>WMR::
PY8LT?X=+MQR>9OT>BRSH\J 5VLQXV?)5W\"84AC5OH-#:K-O'%;X3R1DN,7KS8;"
P[\L"V$JJ)=D.!P:@"2;NUB)5I98?U  #=21)5I@I<KSF.E%3[Z>OZ!%Y4)X7V!K*
P%G6U^ =Z^*PN?F>YM8YR^A_0/68XEU73S Y2#E>K&=BW0S1"ZJ&9MKMO!&UXK*WT
P6OQ)A7]O[WP:@TIQ,Z5\RS'CKXBSEC_NZ&%X7?6UN5HO@P"O]UQD#'JYB()"QR4-
PP^3KUNUO@_<.;)N.!4VOWA)GZJ<:%__]ND";PUF&U7YLGB+)IRA2PMEUN[=KY"3[
P8;' 3+6_"EE*JJYAK8!KY=:V=EFO*'%9KC-DU'R([AC?7('^SU$DIMA 4>$DHX6N
PK-%@OO<!.R[>P\L-$SF##?]^#M_>Z02=F4JT*73 ]*% RA,)@JZF/FX,IDQS_T*N
P&'#O1884=%SU8$\Z2@Z/D&<WV=P\5PV]B]9Q82(-T3!677*A 8$OEM*_,))8I?A4
PZSQ*92CL7AQ<'8#66\Q-8ZT<])8X4U7199<O/OO3Q6%' @RPKZP4_ '$5Y"AV UJ
PEZK]N. &E%]")0@) >48BE39.KV4S?;@M+GW0J6/?H#& 8+;%+>R-Y1496;@1NAB
P0\"HV$:[M:ECG,^&=#4"-((OL+2=V1JB3Y_.]FIF;+4XMYOGH#K'L:L6WI4<@D.*
P88AO]RQ F4/FNX'4)"\WA0IG%GL:3O"QQCM*NEM #<2=GDM_<M )?7^]78$;5G/^
PI;Y\BM\^+4">^1?)MT[J^_(J?G<#\%-^^E"0(< [Z9?J"XQ]Q"#!GM2J=-W;$.0(
PB0560+S?4Q&W5LB7SG0UY/E=$ZO:63LP?6ZN54H'7H1C6B*$DV\?YHFW+03R82;,
PY=W;Z U[O:4I]I\_2VU$YV89W/[CE%(<MV,:$2CY7(AH)=#W&VT9;R$V<>W=G0>B
P\G[C?6 O87$MI$+X'>LHW]MT# Y^OV;P65A//6@(],;> 6,R8,> %9.A.9Y/F##9
P &SKW^4,N8"#TRNP%7>%-372\(3GH.YR:C%@D5#AY@R\F<IH?LY.JBL4+SDS8WB:
P+U#$NB.7:'@%B3P$=_/N>LTUR[04 ".[&E@3O\[TSZ>I"SO&W)EQTAT9"T.MKM:H
PD8W5MQ3S3XV8X\\0$B+8=OQ6W:1NN,*I-6K>%2=Y)'3(_I;UC:41E<8GIF4GA4/"
P)SRRQ85KF9RGW7JL^R)1F4Q6.>_"J9'+.@AK:POQ$DHSZF_TO8]/$1@O?G]G9U3X
PSL:+E76(\CVOHK"E8$9^49.BF'YW6QU6U-M_IA<Y2Z^-]<'HX?%%5LY!6[/'RBEP
P=4D6UD9V>[T^@J- ^3PB&%*]557H?Y5+Z5=:F0F@OR>UG7_TY*#,<3[A?GLU$AM=
P:V;VN@(X6570(X'OY%::Z,OP(A=$32==8$,%AKB.\$F<G-$A%6@S?%YF!TV;,AKN
PG.+A' H>)CU +2/6;G&ZM8N?QJZ,G"'/,(0-6AI!_H,?;0!3K(X  ?NB5H4D7Q@L
PC'4^3#XU/GAR '3AO@B$4^RN:JDSB33O7O&? 3:7$3*BT]AY6.L.H)S1?X!R9;YN
PE3Z)QR>Y(=5@@& ;\ $)U38I\D(28[@U0Y.&F3-)/:MN&IM$+MS$T1L@?4K9PSE.
PH-/R_$B1+GB=K.5\[($U/PTIZ(WM^X&"WZ&1&+%O'*AR1%_\ITC)GY&M)5<+3ISA
PRRDS;A)8"O\LUF4I-H4+\7@A<YGG=[U&\LSBUFM^UQX'_\K1[7%F]/#XYF!'(V4A
P^C<Q/Z21\(C8:I!6#U=]758]7PQ$Z,.<$\=!P"T!SP<"DBF?X5N^(PX1K?7R8+Q5
PUI8*CU[6TVA[&Z#86KP<)E>P87U-FX<!G".L48;7% /=?D#OZ--G65TQ,0#=%_KM
P<L'58?]0%5)2"1D*63;47ZNT6#([1!D:---<?;@:(%.+Y5&[?KMBJ<0?NOX:G$W(
PRT0\PE?Z;>009/19",9E^:1L.O[U8V8 [%J7KL2T+)CT*X>&'-=9,M\\TP?K^=\B
PD8-[?-54CU.IUIG$)%%2M+SBJ8-@R-6]0>E#J;HHHS[(L)'<KB,U,:0MU!)IRX&A
PU?CY#!WGME74:2E+5E;F,!6(WN]]B,G@=7T! 7O.,4OYBMHF.+X"OQT&]EQ\T4@L
PFV1+R,]FTWD!X1 ^2C7)9B>)73GNU5:.;0@HR=$S3=2D3X5EW(C%*.P5;^D S_5S
P%>QP<[UE^XKFD"03Y 68FW_9:;HR#'B;QZ;\GI;7-__MC3-'.V[R4JSYAVA9!\-$
P-*!6FZ#, 9_#(*M2%KX&4>/,/Y*[(H8>_.ZUXC\#+=C,8PZ\"RB_VZ C?F8A;:'M
P-ZD?GJ]*W&0?EI@Y:D]$I+?:*@Z^UAE.0D;^FQ<QY?,]R/2W'*- =_TW-DDEM.7A
PH20M%Q:M_46@S>!7-34 B2.8A,].S$'/12<V@-E3GZ/3X1&Y%TA%2M_63AW__/G1
P&SMX,?S,"94^]T]?V=0,BLIB[UWA98WY(+*%>K5#//2O1#-A=#2_S2JJVCJ$%VX"
PQ7OW%7Q7B\WI\(;!.L6) GIA@N @A2P;AR:O=/8,2@&FE]L^;/L]E41)T+PG^,?C
PE-;# \-4ZX'<E5G1F+BZ"C.06/)#-KH#=%K!F^2$]MV9K!]G#M[=^VA@2DZBN^-6
P5<V53TH/@K>1RFX.[2GTI&N]P>F&+KM<5F!5YU"K/.(;RK3#O*IGJ_IY6LZ.$S=,
PU*8H2%&Q]YSXWIU=-](JVL;#6B?)W7<V]AW8LX$>-C ,.FFND7@.RO@5QEK+>BE>
P+]#)P<<Z%_].6FXI3=I(Z_,OV$E,^7ASLW1.[K'FJLNPI,]Q]KN"D>8F_;K_XRXO
P^4*?W=BHM9<.=C50]PE;?^7/T5A6GF6M_X5(@TAGL=MDR@!AVT?Z6^UAE0EJ.WB^
P_KI6_J3S'#W7$0MVU3 Y(]G!NV QO6AO^EGI5U1&%-O:ANW!AJ8M-@Q9(6@,_X2X
PGE>A6YC]Z,'XF.K%$K1[4^[?^?X%W2!?L-V;PF_"-#\?6X>13(*/X>%$7[D1%7I_
P 1I8_<\$[T.LR"K!.23-(5.?2;[<[DP6?,-5D_=X"DYINW. !:?.D'Z_(^7J"IW;
P4M7D^_%_;4<-;ZH@2-2]\HB5GDM 4((.1$QAMUP$3>]]*OR=KOB&YKI^\KA:S+KL
P:Y)4"06HWQXU^Z?29P$Q!2!6L=V:?A#J74A2UL#T#1Q>[0;THED!D=#"X,:!O@N"
PT)A!G#X<^V]&G:F D\ 5KU,<NSJ,E?OW'NFJ(",&8^(]"L'_0<29(4>#(9'_G?]R
PQJU^2QK6Q"FWN /:U0%DQ$BAA9PC9L.5 >Q_\Y8/ST07;PB?@;CFCR],PX88EM7 
PW<IG*V1D]M*/C%(#%W]V[/;:J&*X[P@'P)G?W HA_PE[IH_6D/ACJLKJ&XO8GFA$
PH#83INQ_H#EE^NN]H&*I*^OMM^;[Y#(^'7U!.,641</+'FJ'+A7M@8JGV)72%BU>
PM=H%08CRH[3A0X.C:YCG_J[NW<@PZD[MMMN\?(X9!,)PV)13[P4FB9./*B"Y)UIE
P;EBCJ=&K#4V<>@AL#=B<^ [65A_%'+ ITM"?IZB@)S,EWBV09DE#<K  ]U0</V>U
P5&)?M_Z OQ D/:LV4T*JJ#1*&?ZI$E<MAQ574M(U\:NN'[%KV?KOF$@8G+=CZX2U
P"^D)XX=%%TEJL/TE:G5<&MAARN W_LR"--U&9CE#))$!F8M"!'<].Y7OR-RD/P^O
P=8L6(:L^FJW)]@-/V&-+^EOG10&%%H&/L873$A"!/;5[H_>K+)6<O_5L5]YSU^W>
P3V"\_V7'!\9E4[K\?K'!5WO3["2EE<;!ZC<;ND; :_VK87:\&W%9W2E*4_1W50IZ
PN)393+\+8EH]Z]ND\93)*.#0XH>85-']Y7Q@Q#1?G,SUM]X8NC%5<_NNMI[8UG6Y
P9D06#+M<=Z6HM01&X1?=MJZ,4]E3Q>=@7X(-LN/-KR?6+/<.G/0Z5HG(V"DS Y;[
P:S%M?@H4R(I$!G>&7W48?S'O!: /FY@UI8DJ'-R*MS>;X@>357<)D-))$,,#+"S-
P4R_@6"$OGZ0DTLP="^%=( D,]*%JJ5LIY0<AL=+. U<$"6/[;>\HYV2*ROH[]KOD
P;L LC[_N4CW+CPV_U13%8!R)OIY2F.'FFF"1KEZYO&N5E4,<-T?K*O9'MXM'5AI:
P%A+G)L[P(*$<4@,!^/KD"ZSG("ON,4[_ ^#A9!RMB(<=X4"VN(C?YUM1ZML! PND
P?_,TE_M+:2O>>K:@2J"1S$_5$IC]C[.U:%://_EY6[>ALE+JN.*7XZ!88.,#UZ5+
PAB#Q4-!)-&G%BKR42)#:7>K1H]&B!'2A5@).W^?&NF%Y1%;)H#<[#?B " S#YD&.
P]"RHJ1Y6[6(6HN$%S?BEW >"_YD>&ZDT7)+FU%B]K9D:RQN8;I7#5I[+[ZUA8]KA
PN/P<(80/_9CY&ER2% P=*\)UP KH@$>\+WIEI 7PTR:%%Q_*%\W0%1'6Z_G+]&PZ
P)>,)=0=CBM.Z))QKHH?/Q4H9-FH268-&Y>R_WQ0X ]I*0S;O+<E1R6(9I,T%*3E*
P!Z9Q?J(EBHX+^L?H5][=*!)1M9P<[<WM9!]TZ!_X%(J^%^/2O5<<KDF)73;X-X\"
P;\2E+MZ?/Z)AE4AL:ZD0@>4$RIF04;0J\5T5E]VS/"&X0\"LG,0KUH:39H0AG@MQ
P&U)7#K=M8HU]?Z[ "[8U]#J7%2,]\(N,7'3'=B@4-'B=6*.I'.'_"<UTIEX!*NXO
PA_<LF&8K6F34D=_7($V7^DS1@&< %9_$C!0ST)-@JL(WMC[@XQ"L+HJ]OK9TZO@/
PJ==]6=7E_30VD%&CH:"$FP=D)J+/;*.9H8V;C&BDC6)37RXP@-S>Z1A_KG#P1P#Y
PU(:ZPB:H9CCDBZ>7 8@= H!%LSV?WPED8*I%7\2?54J7 BB:_ 'J#M8 !!@']9YZ
P=U6BKYY8LG:1W9TK"AI #^^7&ME,!+%%BQ!BZO42??!B4%HPE@AN)]7@Y@^FM@02
PDA>>=[1^%'5OL<?S')?9RM[L<1(^5TDPAT/Z*:53V_'.(?2:?5$+NL7JEC.6O3TM
P:_?^^0*#0M!0C%[QZ2@I[2$5BS2J-*W:].Y.J12[>IF0*N(GXU8H9P(=46E,N-HN
P+B</^L_"-?3ZEKGI=34EJ1?+UM;%TBI.VXE% A]JC,C<T3M5:S=JDFUU2K?"U]BN
P0>/ 2&M'DC ![%27';[/!ZO51P>3SFW!3DY,B$U\/3\_Y-/V**$W5G]KID9DD5+2
PXJ/ *:DJ6OI1#!FSOB>_8MB3*EX3"O8UND]-W8B^MJ0^](H3XYL[[&LOQ7#6**#^
PAO5B[(@$AHY?X]S;7]('7I/AL^G#VP?.1)F'MN'5%7@1+O[@%JL#/1[%2>[DRH4(
PO%!(OEQ?BT?9&4 S.3'[_.D^]"S2J2Y ]Z['9(<@8A:5[XL/$"<)46K^]\X.SI8>
PVS1OCN<5]PL[;O!XFA4QC[)V+X\QJO]KH 1Y#2>>PB<EJ8VM@JYU J]B7ZI6U77"
PDO'JD./])VD8%1YZ;89.,MUEA-PPE6G):E(#O(3D&,JI.D?4^!T(USG!7/S-42S&
P-NH8 $"IH_;>FIBY &ALW-Z,F(VY(1N<,N\"7+R'!E<* >.56^%@-M,="6@O,1&$
P#9VHH]QY:!7QDWKYV&7TNB]Y(PP&0IU'6*C*N!L5QDT@F-HV^\(9)@THAVS5%VM.
P%,3S7_4VU=,H-HP%*9\ 69]_@(*I759>F#K 5HI/6_AG V-@EMT-6D@&)W ,.GJ"
PG *]Z#S#K!!MECI->OIPG/L8;/-Q=X*]"1BHR =*RWH3<MK\DU'FJ-9QK_+WMCB4
P2 TB01&(K1KCH).>Q)$MN$I74%T,!^D4#K[0(T7\@<$T^=I(AIL:_GUX#L0PPN3V
P*WW2JJWR9]ATRQN%4WE"W?U.Z'5H #[:+<<BUA,QRM'=D9-NC5[][]@,GP"WKT7R
PAQW]CS99_VN<KS<(@E_VR$,]HSYA)2<R*Q$!>NS(^7IBUN;SJ,L.OY[E4\IEE >5
PRW\GII$2+2''_6]5;!.3"E71)/D+[L=LN*J>*V!S_9L*,[DBW)_-%RF%<L)A2A>F
P0SHVO^WHAVE)ZB01#X+.S# B2^;S: %%WJ:/%!34(,&I'K^#&73Y>U.J8O_^]PS,
PG-FN+2@2*0]_1J._O-+\85]NI[SH5&8'=!$4#MH,_3CCY4+, DX]\,@Q U7Z:K&^
PI.!4>*"(/@JS::GJZC' _-B L2I(-^5),"Z:FS>XU@9W-8C@.J"\"MZRS,PID'L6
P/9&C^<G^2'ZE;'1\XCW'N6!+"Z U&[KY'RZMSVO ;7>0S@_&REA[,]?T9C!XFY^V
P7U3UROGKD-X-Q5==6KV':]IE&)#+ZT,$;>C*D][J0A-.'6D5_]'#]6)8\(6,-_&P
P\"DKN!;QPK?_K_/Y>?>EC1__]%72$[6:ND$T</N+WSGXHY#DK5B/P):1T6<_1AI1
PL: ?"\A3,:@=2V;(YH9&1.P[KA?Q;4-XI9'.1XK>VB<'.>%-\OYTG&K-C7:HD4]*
P]%*ZN#&>090 52JE)<RKL&M[&/\@,/)@JJ/MT3T)G](SKCYA)DP0%N#UO:B!#SI&
P;;K>GQ.@:5.!+N<D4RZYXB>/&UY1X:D'].2?X0#S_ >9LRIVD[7TGT_ZLL>,?5%,
P1$.M_,DN2O405:*L&5S1B^S;-]_WM:$C\;1/=N?46KSJ7H;IU6 2K&L:&2@%Z<$'
P&B2<F-Z<6^UTD)C8Z+HV@!)^V+7QB$E/8,5:K0X/"/-4<OB<1=>+I7\D^"_]O4;-
P G_K6XG@K ] '(-MD:?4P)*9Z<=V_!X#U2F2FV:31\^9N@:-?M9(R'8"YCC6^6SX
P50]^Z"G\ILX (QL4/=[3.=B9%>//4%<;>FNMPQ4U-W=+U-XMP:D&0N2X3L8,F$\X
PGD"]YI=FO";W?R _;&:Y!OE%7<)CZBO+,UI\,#DK08BB6&P>8W&$C?VE];1)U)\-
P;ZX'9"'B2%):V1ZZ*#RR%N!&QO/JHO7[MWG.-;6V580TN+Z_*-OZU.RYY9=+T!&S
P8WDGW!"7ZH<K]U8N*7>FM2XPY ^:"<166%W@&6W^I?.819;/@!+H(6 #%VFR6JBX
P'V\SY&,_0D3W$MU504%I"%FI&HD;953>NS+RR KO;H,?4T]XL2K&*0[$9')*YL=T
P+J.".I2KHFE*'73('A*$OZB$G>3+W+LULKKR\7+?7X0K"*BC_&_.-IE4=TAMO@/(
P;/=!_)?IR%!/;KX,H<1-;"S%RVQ_()]4X(?%G%(?&4C0N"N.$GRO%>[6]S*V; V6
P]@NU@CW:6*^OJQ ;\C@LPCY]MZ!_G7PU(>%\8T[K?697)Z)G"CC*CX!$$R-B8 0%
PCS<UG(+(C:Y$D_"8TO6L1MR$5CQIC]"0>T'K?O@Y0-);=E&W1+^&3K$0W&3TUQB)
P3R*-5[%[K[D=2((,&T+OD<G0)5$LI40L(0_87A-2Y$'F21?V(F,O'!4W?;0O,F2?
P6U3()L'6?[JKT>+IF4XCH-*;Y.5A15!.#WGET,48"L-V]PAE44&:S%OXD_GKN4NG
P?CV'T<X2J:SX$[R/:[^7</6:Q5',7HK"^ C"L/"FP78S3M->.9S380RG4_[)*"^G
P9,UU44_%Q(NLJP#:6S6>_L8QT.TBTYA  .%#CG+*#)VKX%[5T>/E?2T+I\P](.OQ
PK>/JMGY5B7LVLO95P07(%B;PCYIU,%2NX871]N$3_.4<_21C)DP]9Q,3#KU<(S-4
P8/WHLE>@'XU2 C62TDEMN?1!=&6%1[:C%\D[>Z.%TN*3>E0P]<AMD^<INH$EWW:7
P/](Y-!LS>9>T[1&0%X;;#G-C_D3X@BWB'-ATH<@2&-C)+52;8ZO>@TQU>>(;^_R*
PQC,M'T8HB:A6 0]U>\U81'V!P\.DU*=C#\/DCHH(;5O4)(<RL<I<0_03C+W=;J 4
P-B-1JN-Q:Z?()1Y.ZVM1\Z^^$EPH4ZX 0Q*CRD%;SV17>$\QFBQ:Z-V\"!_MX_W^
PV9+]1+U%%Q8( L&"XRA6KA.QB?=FKMR# PPOX>4 J]2&G(>-I8/!U/+'@GF>0B V
PDK\DSMXY"-=:5\9T5-<HN;I'M;NF^,)G0)#C1OL3*)5$#S42WM#Y^A87/G.]LUZ%
PPMCER\RW8FG>>3RLX8'P,P=P9P^(&<CLK:DQMK [H &+)Q5DUV0/ 0%P@!PD+AL[
P]K<HI$D,?86/C/V[C\B!^8_;&V3T(.CKOU!/!I._Q5G87O6+>\L&$R_9"V/KA.!S
PK8A-3DBF6^DS6(L/@834&:G=PS>2$_&K33 /LP0A",LU%@']>5FFD_+&S"P@T3>$
P5>E650#X]GJS#HX/FJ'O#%\I$<* EE_B,UOG]1]6T3#7>6&(48=,35_"',2W^:&R
P-]) TM%&.3J1\^;@[X(N=%^DD[8*V[%;J_G(H-E$GM.E\?E=!OP4?Z:'Z)O#*M12
P\_8R#F6 0S6V?+BA1M0"P#[-&Z_20^_DCAELYJH6<3>CZ4F ETM^=;\TI96SW8D!
P/(#[MQK*?FH(]H^Q3AX02>."*<U055+8%/<U5'..IY :S+)TMI;:$8"BP"<9[FH0
P4'AE#ORN;(SY8D=+ES!E;C:_\0\QO>,#WDK;EX^DM79B2',B-YKD6S\"=SP USRV
PW:%7>Q.?@;K"A\ES/+AHQR!@R3PXAH&_OK)=ZEQ2SW4'HGJ'I4H#-GMKXZXA4?E/
PU+!NF=1KB%'/F(.JDL.7,&T^0#6,C-^Q0Y-:7I^T(V@V":8FZR?,\V(:9L()0J:1
PZ0+E/YK:>=Q/U,J*@-5IQ;?K@,L-3,4M-=:,W<YCBI(\;1'Y1_L,0> ^F@7^%78 
P@9T2NT'X@&)^;^'FKX^P2G%Y7'>=,;!-@W86PQG/#[T*8/XH"QU7& ,J]@O%,R..
P706>R^,L&*YK0B"\2JA>[C:;1)K+YVQ3>#M/U9LN-QIZR0E/N K!K[6TTMX2;W&+
P3$!P8E;G_,RK!J/[,. ,@]O8F_"D2SY4@L]3W4&?FXJ-\[BH9X9S37/V6% Q2G+^
PMWZ9OCB6J<?Y_UHCKN38ZN_K@@KM<(4>B HSZ9]+IB!OGHH7?JF9$,([R3>ZC]LZ
PL_Z 2KYNCR6K[BBEM.HV/J9_+-2?9$(_E42SLVNGU?SE'Z I?VJQ$S<FJQ[YC,@W
PB6:PG9R@LN9[T[^.>7^LXLO\JFLW94#CL>SZ4TGM!"JSJ!![7%R$$P%0=PVFR'4E
P'&ZJ>+5^LH_Q5V-%$]>R.HXKD5?+_1HSP/]4:XR?]J YIQ@1.NKC:OI-5)NQ$#:1
P%0'&\GI.SMNA^Q%N3M% O&2<+IG)/7'4JC3AE&R96!O,6!A'Y8Q$N'2:D)J&_R$3
PQW;1$SFC%PM-X,#V&[C>[X]3*6"%=?V-I $3Y6/,I6!OF7$<^[>$R&E,[2\)?S"Z
PP6J3G89X:U/:/Q'M>!2S(SN58$[-W>@WMJ6R+4^6R1+G898!3Z8<!6[;K:.OY"JT
P]EO"&_,IYV2AVY5SP*CAAX0GA&^O"UZ4>@B1>F/!?Z]4L,XRF!KL?FLK74RZLK<8
P:(SE+X/+Z,GP#U5A^='Y?QF2ZC.Q1T'M/[@QEUR!C!%&?]1!*(B J*VN79<(*L+M
PV]-Q_"]@= )IAX'*1"IKL5O Z%IJ+L0!H3KRMA M9F@-0OHERLCYR/32_O[+)H*7
P8/(804XC':3*H7WOTV SW?L3"\[9&1Z-TT.R.=KC^#DVHU$,KV_D%0^9Z=0QW&7#
PPX \V%/K&6"<1RD9$_KS=JQGRQDO'\T'?^@ %C!O:"7Y\X4J=9(::=ZF6'QLM/7T
P>^-(SP6\V-2__E)G2!9Q]YG0[F8!CGO-5V3&I3^H?$WV,Z)$E+U2FAY/<AG+X4V1
P:[Z0 KT+W\$#$C1>&IW%@E8N+^I9)YGF\$W8;'E_0/Z6Z)A.U!%KA+LT!<>'F#;P
P NL-D!MAC?S@N,RE#5(*?3DQL7JTKAE^=I&Y&Z L$Y*-.^M9\T6.5HIN;\VB="XP
P2\ !@GTW/SAZC0'SF6%V/?Z8<X/'Z@5>?RF[=UFK5D&EXY//(DM9NR$&@_V+<W8R
PJH8&=K$6:@W?ZK]%@'-3C^J'M2U>S]O1$R*$/PP; Y,ZF#2:\@=2SBCC/FLL/Z;<
P,Y.F&ER5^C"/'!85N3(&8YS0@Z6H![-LQDY)IO E,N#X4Z'>:T$O(L5!Q%/VFLIO
P94D6_!Q?^*Y=6@3WM+A2)#AILK#B.^3<MR?,/')%/W]_[QV;WW:VH-[>.,1KW<:4
P=DB2&;JTU[UZ>V2O4%.+V(@0:9+/'N(>G@"BQCEK1[ZW+,8J='I8AIOF*^Y%+Q#/
P\D_J@*0FMF%QQ.;JWJAUE>$^6LL7WOK@OA35GPYDG*]?@Q!6?9GTZQS,CB]="0% 
P*C'F5?-[HTAZ]>\N%!>2JJ-6HQ:G3,A'YI[/^+!$V(@5SF3[S&IM@()HY%A#;&J^
P.'8(J<%CUZ7YE(?=-V*_)*U4^T@'8M'A G&M]@0AG]&, JZ?I]VAK0CRT0E_/V5(
PFLP4;I.S-.Z8Q$D6.X1I?^U<WV\"ZI27!FIF=<&_&8:_B!/C=X5(ZB=NQ$F( $G)
PS1<%(7197>7V (@4& E^=K#S1P!2\OE89O$*#_33/A;)Y52D91K;&XHP?VO-<9G@
P]$KM+&0F$O@9Z%N5_#P) 5RKMC!@T'&T.]XU!A?Z)Q1UC\!=^<F':TT;?-Q9-8RT
PB R,F('002Y*T3Z^A"48Q0Z%<RV[5J$G'?,9=T8#MX("]X:NW4C1(&+5&%[\9]G_
PU,(#(>*NR%H+UI109'<&RM:ZUS"55J7=1QY 0&L!"K9EUIQ-QLD_LD/IBZD+OY<<
P':WBZ,LQ&*$7?E:$MP1._-%'-;?WH]0]\G]V+U;R%_,<5^(;5#2KTAI RIB6&!7C
PJUEVLL4 "+,5M_!'+&(UN+2Q["+GS2T-^@9BA8*C2?GL-Z!3%&#LJ?!O'(L.00<5
P!B[$(J1Z#\<QZD&PYU>_&$J+ ^?:1WWF;54-^)UM59>FD!Z6Z:0 .QPG#&Q"+)]F
P+TE77JS]@1H3M'KOI6XL*BW58]6F;I8A*'^_SL!!7"UM*YGSX<!=R\2,[KV:PF2:
PJE5/YQ<L%7,E7O1#6]0E0&0G]"NBCP>5L!$$398=YU+)_T6"2>+LUCA#8+W3G.:-
P.6J=BH7 W0ORA>\A3F)Z7^]9Q"+5HUEX?10,1G:RT&A3'[48\JKRJ3 <N]DF2)=@
P"9Q?Z&-Q@__@C. I*[5\1Y]=Q6=[]X%=_V$_S\4<]A@*V;'U( 7FDDA1=3%) 37S
P-U>=J48E7(5PJ40&G1Q'CK!\4@?J!KOC)1LSXR;+RKC[2Y<-(1!"T,([#:?>IOIJ
P0/VF/'E/2EZU$^P/8PXLJ$_8ARQ438F:O#KTRS,3J<(Z";V0-#716C1  %26J!(;
P;9H2;8@=+E@]9H[S%+V4XU>7<7*DN2 _IBJ)<\>* OGD(*_>H,@A!^YH\6Q(?""=
PUY#AG*?.#^/D]TDYL4"518;F]*O?M>)XGIKG\ (TVC_>]4^4W(J>!1KYW6G&B)>1
P#"JJN73^5[A:I&F57ANHJU"%_H@LK"-,.3ZRAC+;Q1IW?4DYE*V9,-9O#?RG<\4S
P$AZ3$9XF]Q$#%7/ADJU?LZP1<1+Z?YG2W4_#/T:HW$GE$:Z8<?C!%>,#B#<J#,Y#
P   BM/U=C]EVOC\;X$S\Z6:0=S1_FM E@I@MQM-*W6GXGPHO_+%=MM1-+"E'%:.@
P+RV%TA*G$LL?#,X0\V"NZGYQ>  >F3+$W<Y.^1ZPVO^2+@[[03&/I2>&UK2A/G0W
PT'*4'4R\PSUF)XX%>6J_>$)P,ZY=]_BHHYO<3C,Z7>8%%DW<F0IMWT'VX@1Z:*+W
PU6B2'(97(,S"3'=R842G0OAV,F)8^29V^CM\C\BH;RXM@Q(XKX2GTU!_?[<#4\\_
P^R+#?C!JEPBV[5VK\:F%1C*2GN(JQAR.'R38'_BQ2H W1\<@^F&I6+LD.!QT#_)F
P+B<K<1?;7#GDX@3R8AX-+^ BN!")_C_1RLPOJ?Y^QO22>6#+)6Q?S" Y=+IQ>LQ>
P)0:6<+2F&PW6':]%=U7B>=X4@,E<S. M=;YXQ$(4PQAA(^YLCGR%RT_D*2[K>A A
PRYA>X09<IW+8W*0;M?JY$XDAZ26KR/&&#NK:0SDL8!9,NVY@M:SX9MR=DF'CFHG+
P5H"4(DAW.W?BV? _WWR&)U@Z:.\JO@#I64VH^\9X4USI&D??$G=X?I+<3D6!Q_L>
P&'^ 38M8:ADH2IOO\FWOE+Q]B1EH)!UT9<+*U^)G*7ZR%2TF)'MWAFCX[ A.7]!Z
PP0)>:9WR@U(L/?#V=<CC5(#(I1:DH=3.<?54^R;R8@(]8(1EC2&.;^"6$_8WGV33
PC--%0"-1Y2IJG)II<48ER#&!?G.8D77M?I 7 HZ7RBC:A6F"UZ12_A5.;E;SZ+P3
PHL-4:A].<A5PB-XDNX%M](9L%.&8A^+"-I3(2"E)$?=XI3'!BS?=NE>?GR*34/92
P$*O=%T -& <GC(P[U.M'YH%'ZO9D\W_5>H7A_#=AE58+XD*I^." U>F$?/WM%'G)
P/G!-!G;&)23X5*Y_<CT#2/?.O)R9HG 9^HP_A-##LWT?L&HS0^YGT]UNEP8KJMUB
PCJU[#4=5&>2(W*/*8'5$F8';NK4.)@*F7)[X@)G53@C36"RS5Y[CJN@:P!A3&MSO
PI@#4<_ZW#2:V5M%*K7<LH,_D2P5%XI3: J1=>6[ )!8CJ;&V@G>*-(!#92BYNQA*
P53A)-Y]IZ$<;GB36BD!K0_3FJCEF<:7V,L\ISQ'!Y)3DV];XB84!2;*]T/<L0X+H
P,7EA6UL!H>"-GPLE$=+APXE3TOT]DE>%?,@R5;*=)(S65\R-_6ECL PJ[X\02)# 
P7ZYQ+=VVBJPNI^0SA!<XI%?&L<QX]70#1@_X>E@V-8;D%JU?R<.??E"M/[<T7<K\
PPJ2--O8<-X<-WO-8GZGY<:M\-G'2WR@XT?&CUHW1"GK.]J H1QW!SS9'#]?ZZD :
PH?/9UV'0!='_JDKP*,05$!<6_-)A]:3BB<SR#_@0OJ#>C^2?A^>K$ZLLJO7COX!N
P'SEB,.'=<<?#+:SG):%Z$RLA_>KPA,VIO>_LL)/9HF-Z [:WAV5(+*.D+OUS=S6Y
P>!?-:04-H,W6=/"_3L1\ZHLV:&5(]D?WC\I!TM"'A&"U:YT[4Z,,?DA^#YR//I^V
P 1KJP*#7U,QSQTU%(*S.F@?NZR[<-U4Z8N$F&T@GHBBA#*NRG8P^6\Z,C>M9ZR.X
PN$_,9AM_H61>2<H6I+)2+2C2A3#LDB_\H<W*VSU\Z[#PG7>3^QM)MIU< A[; &X-
PCZ]7I35!Y6A="S@<3$%/9JI!D;XS8E>DK^,N71HMB>-P\TR6-F53SX([=U.O%AT5
PIBD/B@T_J='JI/I&WG:##IXJ*?=3@'[@H<PU6]^;8<MR%T=4+F1V]-A&U"*3@Z .
PCH>+O]B1YIF@KB(\H=-3!9;L7YR%ML%HR-]K9,A_$06^HF[%N&MD?(H>,P$!]UU4
P#6S)C4:"QS@D WV+^RY#O91S>+IHW%BPBT(HO4ACE +:43:7EC=*B,EZ]?0("'Z#
PZLD50  T:=^-$T3?Q3^6F-(.J:M.,A=E4_>Q%E&@@I-":TVPA+\F;=&&)8?=J6 X
P_J4F, /%I+D]/*A_637IQ:<&;)"%ATK^D$F)'B>OSWF9B<WF6$/0)B5Y#=B+Q#H/
PGS"=Q39O9K/FYD2':<^UK>]LOAZT;^%;/\4JVXQ/?_U'LA(_8L$:]D@J$S87[1\?
P,<HI^%@X<%BX%AZ$)8DN]'-+F%W&WGO4 ^6).>\VFDB1IO6\A)>O+L7U]2O9G'+N
PA&MM1P((,#\H_.06_NX$GF10/XSR_M&LS& Y45/FV[Q\N3Q455H$"V6'_'2<!1F,
P.R%'C;,=V%EWM.74G-KYE+__]A]$LQ0C_?=I+C]3-SEZ78H@8I&<GB?)AU GW\UB
P ?.OU1*N"S,:^8U( %SA?1CRFZA3*]X7.9TE9Q"-V'7!4U4)0;DIIBWZR.L*=@VM
P1\S[3EW5(F5_"4YZOJ!A!!=I;8+7JIMGRT)G@X;+6;S4N2VSQ/QLEM6DG=:O'"@/
PE^A&A#9P96;/A)*,S!+8(@%.6"W]5YL_776^RZ)(5WVX@S(*A0#,6(3 G??@[&$N
PB&)_1+1P&/(S$;*L8LE$19SY7 -]&\+K02<P)H.<(.VH<]\QOP@*SX(C81%IBF6]
P+:VJ=+_3,Y/K[$>2)#43CGP!+&M]6/XJ!D9(2![\\@[HSC?70X\^SUJJ'<GSV88 
PVCY%(;A$OM*.'D.)\&YFWZ@_5+@BIG>F]L\'>^-]UNF6F$(MR">HNK$T>IU?KP9M
P\$@H!_,DR6"$9$PSS#"75RDF,3*#=DYR''$5X3-DO,=5I0/(8R/S3<QWBNX_(="R
P"V=5['T![8;UH&(N9[8PSK%_;PNM1,Q)6PA: ;9N$,80"@D:G.T75]@(H![),2!C
P&5_%]C_1=IK'OLJ6]J2'#XJ\A:=F(, 9P.-J#%+C%[:M3I'K#ZF4G3?&HM-,U=)W
PU@ZU;"0R'P.84^0C!/IH==K:EF9.$[W.,CA'\6X,1,5HYA9F;^TF(X]3(ZCCW((D
P_+4+'OKMZG7X26H:05"4MA#I6\,4D&42RI&4:;LL\N_+95,<]Y^17[>FY0>C*46;
P!4+P$'9W?NWQU#/@2/BKA93:UN*2L0B#&_^.^#U]HO*ITQ^_I-5C/=-O:U&CI6Y:
P,?-2ZG<6U*2#$+,8?;9=<N1BHIY9T7B3<0UE[$.ZE([=]P.+)SEM_C'_"F)$J7>3
PK>CI\&==NP 0+H;8&0PW!)C6TT/]TV&8G*-TJ?!$][1CCM!'B8Q?5=*=H,B.NOR'
P/-7?4Y3X^"\Y2#T_Y2&H,4_-%\05-XMWWPZ1+Z!8=J&L'T.-K:+:4H9WBP?!\BS1
P;@H!:\B9>_ZN2D>BS1A>^K!08'6-W30LQ(&IG.L@ ._<9I)?YL?683?-B+%:3T@/
P#WBZ+.FP?:_\09MCDNB#SB^WDL'@\]TNZ8.RT<+ZB'X1?$)+&H($H_/TH?!]$(T8
P7<=0-H.0I6F3K7^#L9!>3VHG_XJQ\C=,5N%RW;U4ELZ,D]!@IZLO/'0H8*E(\+JE
PR(&M;G8/XE@FST9;O0DYB+3G6^#GXBL_PR61ZFB5R9.'YVJD8TL&J8AQ[N0['707
P#H\G[RHB&P%^-M [8L=Z3;_Z<6LRZ1.&"^O)4(^HNNKK^/PWI<YT9\OGR 1N)8K2
P:BUH<K)=6--RBX4:0L,:#P><<G5SNWS$,C^ ;F?\<N:*78]$)KC!HZB0&,HD?+@G
PG2-2 ;]./ U$5/+%WU98^HFU([*$B3H31S@4K8: \J.H_Z-)%,8FC6]<U-1&+S)1
P.A\R?66ERWSMES :87ZLKD@GK[+R8@,=;V$F$CI5^,V"8,2+V5<6 H QB!?UW@^B
PA&9@_7NDL!?10BGXZ!^;.3"-OAAPTIGF^L(LC?+1*6=D02-17.4OK<9#5L.-%S?'
P+!)E8RU\FV MBR 2%I.3$O-#Y9%K3>\"1?(KGB7";F9L(\0^RY2>)U=OFZY"8CRP
P;GWCGK,]#Z/)+4 ^T@?_4":WE XOM_Q>>\P]7(W7^>^14Z?DEA;8SL1"3S3FHNJP
P&[^;,'BBT9$C&B+<S17QPI""2>[#A;_VZ^U2+9XC!R$R'E[M/Y+0NU7.(V_/BQ>P
P'@C[3]4A#@E?],UH,H,';"(6L*Z:34J:V/6!?!.V]JI,DX7LVZP&XVN<E&?$.@XR
P^U%F$DEQ:B-)>A[4R=>T%C52O$#MCNRS.KF%/=CC^2&>-L+E(DOKA#S =<JU*@X9
P!8= ._+O"%0N!MH66&UK(F\SC/^:+78P?,I5\->UC2OKPP![7G,_QIV6(ZB!JKU&
P?[6%"^3I8N^F-@9X.<A'A_@4;LV "$A6@L33 *#LVO7ND4I!QD9('K U0X6%';ZN
PEK7E4?.>;\.:Z^M>/T$PF:G$TX ;YT)0X5.:&L8B/':+)8+C'W%T[$M,,JE"(R!0
P+$Q4"QHL12;(_9EI8&*O1U*@[M&CP^@$$A1@0(+*9<I[,9#35BT?Y/CE;%OKZ@J1
PJ0/HMVHL P+I5E@B6!-)_"N"HA,#.MJX&Q&\F_I3#GPJ+R*E-&!M5B%QU"YJ[V .
P;Y$%7R%,:!+(^V\I$"A;?=,8E-ZV@D,H']J>8\<$4[PW\@!O\[KW0388RS/52I.3
PZN"<62IN1H%LE"8S9V%D(F!SCG>C_:_^,#S6GYBP/,'HNU<&Z-0HT1( _YU@NT(P
P%?V<#X]Z0AVA:RJ;$5_POI<+-GZ)RZ_5##GOG\4JFY/96.W\P\W4H+IC'7)#^E^2
P[1;F;M5@0N25^0T??EJ]J,M[CR;=.ND@TF]*>7MURX4&7,==9%O@7*^^'16E3;R@
P#IPW AG75%8V1("PT08<Y#V=H"TRGG4]2YK%Q?G]HZ$SP+E1EE9P>D2S%PR<>F^J
PJQG.1(X@]U-9">$OQV6"+Z2Q:Q.B,^B'Y8X-ZFZ*9ZUOV/ AJN#_Y+J@/6\%F9;6
PFM"O0W+@;OH3O/L&O#)W;4>6FW=PYPHQ_X5(4K46049&Z2<G]V)^IWC6P5XYQSK!
P_^WW>E^U'@]^\+B;#H+SDAGI)33_E6RD= VC636)XXW/C48B]"+="_B'Y^;KJ>C5
PLU8CUF$K^Y>^=SQ(7!HECPZ64SL,8= U,ZQSZFL'TI.@Q5-&_K]'YIE)63 7DT>H
PMJ]_/LMJH=='R35[)PIT&]R?*8DT+Q1LVAB.*O 1(";@?<<TO.^1_"(I3D.HM& B
PRZ+VS8OTY6L&%<("DV&\?O+HEK?)IN$5NO)6B]4?%%2:M&\G9@]734FMD<:!=\9,
P]?\8Q3427"T,>(RG8M1<X;4-YT]^/+VS8_(CYA\?TW*!IU9/8.2=%Q-&MG^;[SM-
P0R&8O)[B)T'!G7E=^MZ/+OYMQ3^ ;3 7+$G$EJ6E$35"0JO6V5-T@RT5%,PN(+4B
P;$5Y; $IS<R\)*=#^2[ 3"^L:GJ.@6]O&"YMW5MT<0;6?.JELT7*LW\WM9QL/44I
P!&K%BMY[\\8MC$#6Y<39]$LM']%OBZF KE625-)+T.2/IH0*$G/0-=7:[T_3U68;
PG%#:Z\/*47^7Z10\8+8KU^M/7U7.T</'+RFYU*6\6XD%W*8DF%%@DD4H&\>?48S\
P4.X"/%IY5&IUSE2<DRWW",*C ER+EI8+=ZS3BMZ&,D/&UC14UJEYM^+MLIMECZR*
PD R=5PG.;1(\C=$U@[=XGZYE518E9"H51OPFG3(3CD'>E&&3&)UA%>)'+71"R/XY
PR5G"*&B<[3A&&_*V?=PKIZ0LR5SOP&Y$OEV?L^?INT$QNOB=)CO!2NR.3/V,>=1[
P?E,/6FV,H<!0Y_ G#=QD@PG]33[,U1I4BCHK+[N_!.>H6ES8<<*Q)H6DEJOOZ  V
PG0J]+Q/NN])D56"T8Z!(J1Q)I1I^CU0!JL8.Q/8XE=*0+A)$Y9#IH070M,+[\G;Z
P1+V.GBTP7#2-Z[/BEI(&5>!"MX'O6GVD.,N>Z]2-SE9J_@;<^2O\'8-$+RT\B#"-
PO>-TS'.DCCV_AW_5(:27$'1J[/:11;'(DOF:_V1Q@X85.@^HO(/6TG<LUL)H)C$F
PZGF+RE#\)_'-K'7$DEY6EDE5CN-$,4-[*7^Y.2):A7@F J#CRONUVJ8@SBJ;?; [
P!DA#Y*8D<+5[%^1-\]@20Y ^FCU[3-=9!QO5N7HPC?7P+!P9T1@J S[0 IC!$!=K
PE)@Y%$=Q*3FP4RS!BWJ"QCG_@&[N';R)>L8!M!Z>,$M9P*X C\V#K81&C3X(YR%Q
PW921C!U1%9@HXM;S:I.?)121$ RC&@T K5*0!LRAGE'.?JENH]=I%T03Y?]0!2<.
P-%:[6A-^D0=R2PR)IX>T?,+C/'-B[./KJ(!: .E,K:&R:..UR6,[N0P&O=12"==]
P8UO*J30V5D"@WH#A_RN8,E\([C:!#]= (HT: &._W98@=>6Q=-AV@[HZD$=%2FA#
P,!T@TFK+?S^%XUH^#B1GTU6$KRZ>GN0KA?#$P,T(MAX7:_$DC1"3F$]5_$41HE97
P4]$.GADE6_7?!DR2C]I*HE&E6P\8,AVEV?^84.M<VP"8D^B%-]S5TXZ#A+%.6GX6
P&<!\H<&I3QEZ3L=[]!:_--PK57[KV;9N6/#O"XNUVBZS0]6PI8<%#_%:O-D=,NGB
PZ46,PU(@V@0(1(&%'H_6MCR%R^)=N!8000R9B13K'DOQ<XUL*'WO%#,1&]"^^C#'
P4:\E2]<()\LY!(NQ!_-;I#<>XYMW!.-Y4XNRZ)7&5=70I3EW!5J<H&%*R&CZ!TZ"
P'?0/[VJ%'@N(;3:HM37KK:!2>'M[Z5)/(,NDNBF_!.-Q!P)B>EPWW5J4IK^SMJ\5
P_T7 FPSG _SBVNXYCJ5@V?':Y)-9!";2O;@^@#*HV4!A]J1$1%IITW ,R3VDQ;^W
P@5M?D[2E[G2LV6IC0S"'\5Z.=XHK+EWL\5\ASIM@G*[DU6VNKTSSS-%0MG_UO>VW
P1%WP3O#_=OSMTT%63Z.;(00XU^U"I2BZI5%7$L(O@L*HD5.G@<XE^=[M.\6HBKY:
PM'&F/Q1\-^.Q67-*18+J-9CS1KOO1[FV6"OW-^6\=^3R?)TW31H +R!$QH:):+!:
PQ(;:NSQUQ%"T >H8^[3#%/ZTG[4[>+X(<AS[;ML4MS!W5GN;$TD'&6X,!"_O_TTS
P.)D03GF=D0J<>,QX]F['IH/Q$L8ADM>X,M(6"07#UXY*CES,"9318\,\RUUQ/H_&
P40@EK([9WZ$&8#P4 PIET@F3#>2/@1@2E(3)72%7FU//5OUPD"=&%M;K 'MF].U"
P&I=<%>6>O_VJUX<?EHO!)#R:8R#/PWQEL84]^*FZ%EZ)C?0C67JO:H'B&!E)\%1G
PX=TB2$]D]01P]5CGD9\FP"G*/)"54!]#6U@0!Z>[6(U@5!B[0?!UE>R)Z8^< _J+
P>,II/.#!*MC0_EIL(7-O5F84AG_714[$]:"N8@5,T/F_>#(Y45_Z6#,P9JFNTCVW
P6IV!V6[50:$^S7.P;A'H=(33[3(T X!":9)U *J97X+H\$0BPPX9&#<2TVL5(@]V
PHMD6Z%5WJASFG]EIBY&AWR6O?!:[=?6[\?_UXS-^K;6$8KL"RU*=5].+H1?8&R!K
PH+/#_.1NL 2] OU%^<!6(4:J0HOE^_RX=@CLYU^)J"#,H2T)YL*22F/,+@4]Z#.9
P%U%"N%ALP[N4JY$$F7)/Z??U *U4VCB)GE=<F^2' T*T,M@L$&.XWG9 O]!POWU?
P@A/2>V$QR4@AUBEX07OMR<8(D,9>J.1.@<JFS8M/FAUJ^++B_TCS6C-RUL]_Y 7*
P)ZMMB-7Q&LHA6JB^C(#_2O"S89<1)F/O .-M;2'@$T1U< JU982K.!39$00106 '
PF@^0!9WQE!U8YK>1GPS\>0UE *#JK3RM.862-IAF%4Z9B\?\SG*7$GW9OTUFAA+3
P1I0UL' _J]LV)"?,K1@>?^G>J)O!V%7%_V Y(]?1G#I]MWPQ4Q1R_VY=>ER@DPY5
P_-5=E]YXDE0,#15K,X\TUB" %M.'TXZ_VS/$%MI'@-6Z_0T* ?UM^L$08X*>$C=3
P B9(V9:/I5VZ&I0$GA!?*M[ HL9]EJ)]$KMI(,E><2NY6AJ3C1I,=[1Z1?"]N35%
P6(N3Q!9N2$WAHW*;&F5NPNK0F\5QC8)%3BJJ%M[N40)?%>$C"DU<I]\"#93ZU&SS
PW69E^-52RMPEU\MY0:$X0W!%AF#&M%L)Z"OJUN.L81>(OWF2IO9;583Z0&=OF&YN
P,Q;92DFW)W';7J7?"I2=<>H_:>==H2F-=W/*-@>C:"".XR!U#_QG]%L@X()S"Y6M
PFE:G:-I,%6TS>5T B'D5CLQ6PY[J8'_6GW00=OK]372K:"'S?9_2"89O#-^$L.UA
PO1#X_^G%:X_V8OAX*Y4KXU6HD%0B:+?G%A/6S5<3M#1/"%H7P88#D?-M72P1V^G$
P*3$Q+6]C;3MS[ !^C8]6K1&1D:2D,4&B;+MW=J4C#DTA[4MOJ\6D%-F<N#M 4^;,
P^1G4:9L.NL^&PF7+Y3;'^CZ_WYY"9$Q!G>;R8"']D>7W4?M72N>GXG:]S'?:>ET'
PBYE>P7#S.&:QS-ID$U_JL"?.HHRL7C&X/=1<<Q+K:*76B1NN2>NS'A-$8[_IUM)'
PWG1DQ@[1P;/3.,*0JK=2^@WEP?*C5W#RWWI7&&"0_FF @]U))?0Z9-$DLD2/2F(U
P"LNZ.D6RE).(OI,(N?]H1ESXK+-W5A8L+7/:N@5+>1WKAH04#O;S@'%"MAX[3U>E
P[^*P^F5D<:%I4AC+IJRGHE_AXO*VQ_,U$3C^V"@87$FAF6IJ^M!C<Q\I(VE%P?1#
PBZRKUD8Z?5/*CO,5D$%-O22N'':"6737GYH==C$<%[JFWROB G"/&CQC/3/S$QQ5
PPZ=)CJ(V6PXZ90NXV\9Z"8@^LO:%*B@.'&#E"J^$T=T6LI#W/[8J^ J<*+H':G5.
PK.3*_Q*I?DD2>D;DPKU3BU*\0=-#(T'=>)8<W51O3C[-/Z 7VW"+EU"::U<R=LR7
PC"*IY QOBT-76%ONES+ N18U++;X\ *=0D59RH8U44!>$!?^)!NIMB?*K3LQ3O!O
P<SG)B^F"T&!PG=%C,61CN;5-U''+C #]+&GF;> 9-TOLR>0(Y6_W0G'E?KIWD+3$
PH4MS+)@%2OR-=$^F,NHK*VDO?0:A55-#3I>EZ985$9^%OEI7;RL=E[9SRT#\O;2Q
P8GT!GY7PQ]#5#"VUU(I.X"N_6_"URUU$W;50099.X7#;DY=B])TOJ]9O/5,>Y%IE
P4G5;.D3E28SERPMK932EORYR6<E%"9N@Y8R7G7/O")H'YD(.,4D=_Z"\L)\<;!,+
P,$\%X:TK]J;J@I2!QJVN1WKV /Y4*6B^VICPB9 UR)24%PU$0DVD['B/6AGCQ!%X
PTV6X0"8#SM$5 :='Y;:Q /\D#I1XHV5>E>Z_T1[MM='H_1AZUP6W,YM8X"N:S5XJ
PE*HK5([T?<<84&-C<&E1V)_7B>9N4$M6T;SHU]4QY@]_!%3-W_-J\''Z+>Y4+-^;
P7I;_!Y=B<712$1]*MA/?:PQ%+U$ZBL#CWS!7-17!X,(#TZ?>;:O8%C4??0#7R>S?
P$ZJ6XI$QL^.MF='!1M5:W%2J@?O@#6=?WHE ?C2\)\[#HW<909P"ZW8J<0[ON@8H
PP%6;TN7;GH)#U+()KM>AD7;R-T]*W[M_J?5GUR@RGH</*[83 4KBX2J>;S%RC#Q;
P-VX.:Z.G./;%N9F#7_5]:]/^L#(=@8=;#UA$_ D,^1CB$6V+!$_4.5@Q\E#-/[:!
PT[=48FA+. L^E0A I9E&:8NZ,<-[\_ABX@+"4AV>99]2'X4M<1Q49??[+O3NKVH[
PH#U;PNYXNKF!HC1=LJG:H-K=6^;C<6$=@X^*;-GU9CV2<!;QF/)WW=R[8THITQ#_
PXK>.& JS6=MKMAK;L*AZ^HWF]@*WY8KMM."[C'"?9+LC:%_?R_Z50<=_U4AP-RAQ
PZ(X-&+?MB9XKXC%GI6DA2ZQ8'.# J_$0HHGE6+#$.JM/M<[EKAS2W?_*LK<J)::D
P3>W_11K&')!C@%.@+NR.Q5QL!D[8;1F^:GMK$#PHXQ,Y+W%M3/ZB:60&FDV?O]_X
PWSC;8W-%' NF-69TFJ@OE1P=E"H=K%AFJ-K[@XO(J(W0@IAG^1LEI^-&>3<!V!'N
P4G2@*4Q?64I!@48"+67X!]M??QIZ[1%KNIBRF[@!B,8!(HA(_S2P="CA";^&'%TU
P=BXQ53#C>N4Q1)""[9M9YANSKO,E;UH([/\%_895!D4WEK0.V*K'K0-(ZGKNS^;<
P6N]Y^*N0)[E)E&;*2QZDIXO(B3-.OGZF<HE"(+T$TCH=3Z(65/&*TV":#B<A%E5,
P3C%5!93<@_?:I$@^2F@W;3!U>6OZO2>;+0&4<=KV$*"9)4P">KORX!NNK&YXI_<$
P2=W@72"ET=[<H&S^U0TZL7RG32_Q)U_0C?@&[-4$+9E2$W,&; PB_MNYB81WXOS5
P3.:?!,UG7$M31!EU]T P,AX0OK!G$.K7#( 9K7,N%?&TU>,VPHE-)CZ1V6L<I[=1
P>/S>.TXUFW-8WKHKO)XDOSK.C;&_AFE]ZI=(*;"S>/^.0]?E/D_@/]0-IGKJ(5AP
PQ0ON MZARWAML :*VEE+O*E[3$Z)4^A:5\3\B?*ND(K<G2"V@82O>(1$,_;E$=<6
P(%$S2H<9V)$A+HXCWTC%,2CK],4$VJF@S2I'XT(3C1[B\3V@_P-,05P?@_#36 '=
PGQ',RVM2^MH<90/X[0#[Y$R.V%P#L;6_ )1Z?W&2WA8E0]K41U"T7KO-MEMK]C2B
PXF9?(T+OJ!@H39[[[1,@DREY,9X![H66?+RSLY^Y440 JC],ZVDEKY "#^15P^@,
PAR6MH ;Q19JF&V.$PJG#4\L_2<H '2.Z687Q('#9MXOGULCV6!U/4R9M[I54K0![
PBP=&B[^K&<6>M/)]B\-5X"KV$OOMWN3_B6A<2\E"ZLR&!3SHU\^TNO%3D=6IW_8E
P^0E\K2S<,C89:[C>EN5OI_FW]C^XA?9-\T"!-@(-T"8P&2+(1B(>"BIG[&6P2V3'
PXQUFS5E]56P"61Y'[SFN<32Y "AN;+A9-+PFJKSE\@F6-C_0%'TMT!.C%8)V*)4A
PT5A\_/>+C4ON*65[HW^9'L*!R<7*OVGT8O#"[-P,556#]"LR:$GH^^F<SP6M3APW
P:V@5' WU0MOKRK0EY7'Y*00J*,_W1.4@_CP/@BJ\Q:FP?::)Y*&F#80XPTGA/))Y
PP?.T#R4,Z^)E;IN63Q8?".R3B]K.]J3VPJSAQ24&1598F.7CU[G);WV2'!/'^OUZ
PX=9")8C"TS7(BC 42L1M^T7G_3'R/.]@J]5-HI0[*-FG*5@^<I-B!HO+9'6#3=P#
PGLQ2?*ZRR#$0DA$#X_.1M%/TW3R/.YI"L.0K8-(OPB"OXU47,XDL^" RW=6'D)\1
P& <4L7 Y\?%TO@4EKC3<:1Z,N%Y<V:E@.YJX8X>5RE;I[@TLH^$8X *YA_/!?S)I
P0;""S'Y"(N2!M3X:3:N:09['RPH O'8SES L"C]1NX LPJGO_#J_9\I2&YG!Q4N7
P^D$LGNX(V2)/83H_]\Q/G>ED!GJU-$A:K-">EO&RBOC0B(MGR;PTA.3L*TZ8%C\[
P>YY12X+\36^8*GC[(:CG4@WQUI[J/CC2U_W#41Y0[@%%'3AP5E)FTI@K1&IL*.T 
P:4V:^]CFV?(>A-#*8K:;!YAD(2!**4C9PYB$Y^!HVG93#;@O,\Y5"\M/WTSP#+.X
P?_J,NX5@R+=',D+_*::BBOJ_VFX-BN<*8?+T0^^F,^>PP&%8%U\(V]T%\3JO%D51
P6G"+&CMG>V>6R"P(#-CAF=#AW^NR*Y7V29]8_.6.$2:%+LUD27Z(OA#07$J<X3+]
PS"#!3L7Z^V XEK^+,PQX^CUV9D)G0F"W6!+^SA-R7$XNQVM'Q"5$RFQ #-5K#^Y/
PZ?%$R,E_4:POG(- #,F[9CE6K>XW#!MDWW9C.X;K7$]A; ,,ZQ(C-3:@9$EF4V?3
PLA/UE@.#-4[YP@Q:RX-6LM^.IU=;=?7LU> ;E0PSJ&0\>M/#,>36'XFW&[J#KW'2
P6A*>^K=VD=9/.(W1[B/H_NC(I(JFY8^+TIE^4=M/L282H1!( Z#P6PY5KGQ%?#P>
P' FK4'SM??/#V!!JMDN_;.SL*9%W\ER[O'V@8*NQ5[4O>^#D%6"^6A#0F,E#QA3,
P=8 _G'YHX[^-78*W6F:14,G%'8YO0\/91)N$0"2-V5GM.H/E4'&KV:(8YIW=.,?U
PG<XNOMN#T@2R-3-_9A%<W_T@Z'+++PBU<WMYFUXNVS"YY3"MH P&5$=A%] [U">!
P\JPKE!4I\7<0N"U;@30X^3HQ(H<B$H012NY<RB%_,R<S ZF=G=E8SW\8=Y2$1'\Z
P_VS9W:Y6R_$16LY'-(<QUTL]_ZZOT\\3\;W_KV+A90QGBH4R!""O5_S(Y,">R\!X
P=I;U*1=H5!%=;P@(54>[&$SN2K+'R/MNN&5""E;5_*IE6GX>GP\(P??7/W5,)WXK
PR">F:4^7AI,CTQH.8.O"**913I=N$+!M$?'UC+;9WIH3&],TO-U1 7;'+-[*HD@P
P$V%EB26!B$63:!DX6E[H\Z0GB51?C= >A0=?K[QE'VL,0[ (2Q$6ZNX&+<E@]>[!
PS=0N7!:G88I2=D0O-4_7K=\VRU\#:F;$)NSZ7F>Q E 7V@YX:D^H -N?(=5[>X#8
P^39RA>KD8"E*6#\L234>XZ[ LSIL5Y_Q_XT$E2!H*,?C:)40;WBNJ OFJ&\X_JK=
PL!/7Y9FNL0JM,&3 F W8=U:;X'N.D-$P6%^![L=*$7BC""1)AMVY01*%%OZVA&4/
PXV9MV"VQ3QC"FU[:MEZY %L..ULN07!SDLJQ2EAFXAHGT[>#+!A/G&FR+B[L=<V:
PU5#K']"@!L\^438)K933LZZMI_9,P#^X,2AD 0FM.'Y80"(#W5.(6LT?+C\.9*5+
PG9>V0B2V/*3S#0,H/?*B(S>!_JYY(@=0A$UBB<XB<4! HF1#I$:_E 3,"5-!)'9>
P5#1\L,NP-'/RI>?/?BK4!YA7<4)8[S& ]]\)F+1 KT';]!,#1#(KL\@MN[VYO0>K
P-F\C'-\I39HZ*"V"2)0SKS]]<K1/AP>-=O=_O0"_<J??.+%1J*U5]LKHVU4^CU>>
PJD7<)YY)Q3TJM8<?E0&)<.22'!7O*VKP WAW4D0F8/E15IQ,AHOB8<=N/I8+?R 2
P))'*.' 50_L+GDKB2Z?B4NP9(@W8_B51#H!8F]1DDK_Y\=#011Y&7#8B83Q- @;V
P,(XE/D(C77>H-/[RG&>J"/>#H=LR".5Y".K*(JC\73H9#V'TNOA8)\<5/ S:<UW5
POB9:[V1^YAI,RR_#Q,FCO,6,>RZF%J5BY(0/L#IW>OD,C H8S/*'?@?4TX!2%^/<
P-Q%<G2D+X:C8O>F+PJQ#CK'$\=FM;T8T(\LMU>Z1&A3J@!I%3@"&*C47NGJG$!J#
P1"2AV$JN4_-;WO(6]QW O0=Z,E;@[-3$#%A#8@S+,03VO>A=56HG%Z 3&/-W4*AA
P=@+H&'Y='WD^3Q3GIBO+3B'06*'$2-(:TQ^S DU/'NO.J>D7/O#>9OQ!ADI0+U^7
P0'\L76V;H8= R21Z0:JG+0^I4 :Z_)Y#E[Y(B<S#]DBD$Q:\N/\,&<U?*R\6I5)I
P!?8ZBB[V&M]*Q#/404G0?XZHDO9&*L:NGV<":B?^.PUS"[&(IVEDWJ9M59"2C\=I
PZCD1EK _%][25?& 8<$VM*&Y^+_;)6%_$P$AYGNSLC#I3%GE]L9A-JHQU&[)L\GF
PE8XF>W9..<!9W8"[RF2\:M#KY61C"''[0SSYF>5*\4E9F$RR\SFD].>-,._\@>NG
PI:R]DZ?_WQ,U3@>Y!C E@@ M)>I1"GUCY-XL+O!C/.BV%)SW1$<T;C[6]O(VM0$#
P%4Y_U([L02]7G1&,%T62.&Q[9I7:TEVL?V+_3WH7T97ZJ]"C&]"<1*Y*AOA$B)+J
P;XBUF&D;("\X[$#CU!' C9U+D_H! ?,7IFJ@UOW'X:Q4.A#!E][]%.+4J06$?UW@
PCE[8H,]Z*%]0]]9\*+L;*TKHL/EN5E7-20#-$O<;'6\C>:!XY3<_8=D?BE[PH>5!
PB.5A8X>W*O4!VA"C^HL.E2\;TWPCT_-OAGX'0 -0FPVCX!FG.SU0+$O1:*CXZ7JS
POV'=0=GIU)UW4VD01RN$0*"3+@-PH67RR7P%G_)>13)8T@FFLLB8JV*D/:$6SG\]
P=1%X U?$1V@6X .89WIN*?3;B59,!E&O,3'T IEG$7D$/*689%,81:)8?8AGB+O"
P@^40B+I1ON'FLA(9@<C#]+.,B)>7 >-F2:4[TD=*GYF.861#S.+*WV:X68VU%1-@
PQJ&P@EMJPD& Q! <N9(=6YN&5?M_[ MR6(.KBIDJEN#^>_^B:^#_N?Q1)PQ*=JT^
POQ&8"S>0-E4\&#/=];CJ6=:Y#9"IZALF4:LH4%K.HR%=" HXFP(Q'9<U!8QIMU7^
P]O%*PZ5!]!4J6=Y;[ 'N5.A=;!+D"<VR,E#%NJR:&$TEC8/'+4:<#4*!LKWDM2!]
P?.(+\? ?H5KHV#E#+TXUU930:;#PLU 7L6M05JA?^^&0",JTRS(Z-J7O@FU,92HG
P^S]]BT/HG'9<7D!%_[N/W/WB@:930NR>8P6XOW="BME$ ^&*;1,J6VT=*79ZLSB#
P3!CD>T"9K"@5%?-$YT@UPD9EEMO723D.U%2 W4F.[V2SO_XFW^IL'F:D&&ZI8 KS
P$^>X[+;90-8<UM4TD%G9R"!,(NBV,>X96QSGA(5JJPT-0^&*L"1N7GDX7SV=U+_R
P_F_)C884EQ]UG\J@%^(G>_@&5'3:"]Q;L',)O=B-;>TRI_H+HA##'USELSX2J-8+
PIN/XW ^YV9P7 !REH+E33-X 2#OL?[T 6);N4:0/$,GB=/[:PF-0+JFA<GH!X_ZK
P:KE+I9L\[:O^NZ]>J,A$WYNXI+<SLCQA8BR/""&,\^FJ7@]1OZP@T6@LJ=JTGD <
PA"4*$^5=(!R,@#DF^(]BA,<D<0('(\OMV;4Y&K0^&@7U()-+.XP>[B3JGW+:3R<F
PD\'3H/,9!7T8?XN9 "8V3]@C'L?J%]+<=XMY(HZWZ43\4)7LQ<RG*CTX)I9Z#CB>
P23,W4Z=S2]WIC-.E*G?YR:"AL&SQZW@]6-N.2XR77!&GJ!'^4P?70L!?*C\%+9F)
PR4?)0LY1O83YU9*,1E:L$0;C>BP;(< +]NS8'X+*.YK$M/3RP71AWVR3\1*L(05&
PV=L(#?T"OTJ&F9LNR\PJ:=%R%,"JI!_FGPV).[@Y'MS0$%/=^?T$<RQ9+K NH,5F
P8K"^ P)T8A8XNOQM8N&.>R!M/_O_9U+8&[:DG_O9GNZO)X5 =;@C3JX$Q6#?GZFE
P +/A'_)>!:9/N1'0]"<\]R6+X"+OD&#$8%R5&F5UWTG,J>,A$F48<9C&7@I4)L=E
P3L]$$_FW<8/2GT([F;1J87[\U(OI\18[ICOSNF4F9S(;Z!]FCR.I4A7CI]A((-G:
P,V2TL!Z-;H;H6>Q2]>6R2,:FAWM>E)(/7/8#@MS(T)KZI:TP&P)>FRME/1J.(/Z&
P"P1:X5ZF:8'K/Y:5$S;$1T'_$@P0H#=RKX5)KBE"NCY]I9>G#[EP'R:0/Q5[5YP>
P=M/.B,\D]ZL?^U(U(+H>'34Q/XAK/-&-[B-#1,GWSV%^WDJ_'AV!6.$\%N]3FV"H
P#5:2B\_-CX9_>Q-'5A_$+=/HF!,EZ.MD!RR$H_<V5RN_?HJ%.'(V3P+&(J+[3B1"
P6.$S 23JQ;'7D9]Y/NQQ0/)KO-T['1N*&&"0\@<JG+*0CX>^/>(4N%=(WO:V$DPF
PT:S"8R [%[SYRN!CC))_AN;&'X$<QN(U[U<.]RU$D-^5V*IP\IG\+X3R2_3!RLBG
PU@.-W'<);31/NB7:Z5#T!E=Z;MN&<4NG9?*_E%?AME5Q$:%F"IT%K[5O:FBO3] 9
P"/:??J7\19?)0X7S,2D<IS<4\NN?@X&@\,%Y]JN<8F,4]Y-+=Y(^<"(@?5>ZF7.X
PB^6;XC:$=\\MT'"XW*+.LPY\.RLILL(Q>YLZ(-N,:*YJV8FN3F<>^%XO'10-;+KS
P>\BJJ91AQM'<SUR3ID&P5K^9^.AR+\XH]B^UU.:@!#CI=&RG#T[RBBH6/D!]V#I2
P]R9!7B<BXA.3:.:HJ0.FC/^CMD&I#BYLB_ !P.BO5NSVH[>> PB\90.=H.9(#HE&
PZ0>?6?(Y]+7@:N5JS+0: 3,#(^V905>FM!P\\;PO'=N!>',#HH<C!Q6]4F_0</&4
PC#X*Y(27@=W2,?M$R0+E,O?HE8F\.#U/"Q78\^-P;KVCKBLSO*=VY8U;@"0DQK]Z
PR(9F'#B8EORWV5G FPS;74E_2)KM\4TLCQ5/N9:0B62E_U)'M5UW]QO?LD9:GXBE
PF3O8GA%8BD*)%27(+NT_.XB[D=K[(UE\&WEM:Z'4N/S8$YC0VL =R3R($E4NVT16
P-RRQ2O&1BZ/B\ (9]T$)#NO_:7N=H\,YS;\1MYSNGI^Q#J_N9Z+D(%WSPPBYTB_"
P5!#.85S0;S$&\F4+QP\*NGY;S0S="_Y3N;PE'H*Q-HSOF[W5;G-B> KZBB?;02AJ
P=[$0 :/E/>Z/N_DFH7!\G26WLCG&8Y:]>8,@I]M*,APE6E>T&N-.CS?"]/GF%*CA
P^R2A!/Q<I7+$:96RYC3B2N-2TD]J5=A=X>IWZ!76^8YTJ-=G3(,@:&A0,D:F*@A:
P=C ^=YVRQAH-.'A4O519!&KW)M]>!JW-:'F?203%"A*#I"^>W_T5;+<'G0.SK?#/
P^YB0\PTB,*A+O1;.2.WME(6GMU;R0!@%L-V6L%/!4 /#>&4]B,0RY=)!6"W?C>X5
PW\+5F ZG# QQ,ID6B0Z,'I*36\<^@[[>D@R/.+!'XU27,D_@E@+P14\B@'K]1!BG
PE8+N-+,1& FHZ&\"XK5W0:+"\>=$M?J.#NSO:OL >E.V5RL6'8FG9.#F.T"\M:=M
P-YTV)F!.'"R\Q!2!W;=I?-(OO]LR%3,I;P!ZTP1*(6\Y"Y3A [0!3WQ)G>R8MS#O
P'Z;11>D[%@4*Q[\Q51H2U [!#LQ&!MU_^@4F/2M&=Z'$FO? HHH6%<(EA^5=[*22
PPA/+HYCDUJ_5ZJ]_U)E,$_= X5$'B-,R;\@^#-)&QM5,-.@+$ ^?KD"2A]^D*(R;
P)& &MX/I>,Y9/ERD:]K;+*@CNW1:Y89YFO6K>J;.N0?N_H6,@J$_06WWLEA0BG?,
PPM9F+<?QY7+<@6=4EFRMD/V5%?)]P*)TV;3:>L+NH\1NH<2N=3"_1W[]N-G2I?@H
P.9HL;Z5<*(>*15R+.A ?FW<XM6$7$/  @_I+R[P5*XZW?;5SZ3IZ^U N?UYWN345
PC$)<,Z#$+HMO5T+6PZ"D8GYX3+G=,K@A:2@SSVR=8M\^J7738JYE7FQ?F.%>\^[W
P40HJ(SV>0J#OE>G4)5-CX(<7"?OK;9C$!@K8E)YS,G=2$9VV4'3JM#$FMA"6B(J,
P7Q/6B7\ F<?)JBYOXP*/REUYQ!Z=,\>*@_DJ(245;L*YHL/4,73+[?0T\_T*1FBK
P4:%*)[/4D!R5UDSCN]#9QSR&"L!,4$BD4%X%:5_Y!Y!BYO3G&(N#:D&S95WDQZ,.
PR5\]+I:&C^M_R(N?Z@73YA_2.^>(9TX2/DRGHQL:+T3U 51/@2RG4[2(Y"15V08Q
P0JK^K_AT BD04J,9[S%\@Q<4==<H)#M9"F@D[5;,KM^B-K"8VW(KW8'#%*H1I@XC
P73]JE$YKRQBB'KTFP<M+HN.R:D5Z0*)^RR=CF]Q2)!7>G4\;L5TFT7,@_ '2AKM:
P?X,*.3%=&P!ML<];*\3[!,ZC614XK<2#:/-W95%8BFC_/]L.Y2O1'*+!!UUB35&G
PLDTQXZ\M!O)JKO63#I$2J8971],'N]WA.H70JZ]&&*2&&<OLTK?20&?U:L1\.,H'
PE/B-V\88U5\!ETB3^\/7KC-..WTK5&&E]JB,X+?:*[E@E;TA2Y&%'/J\$7[4[ZU2
PX%G 6>_M6.<H3W36'I282- 3XP#.P/P^Z0.F46J4LY\T25&N<@K18YCHQ\E3<N-P
P;S6PVS54+)<^]+[PUX/QNQ"V5,@SY%#-M W^T=8@@0MY?]-+'+\)3TT@,0 &7/()
P;U@9R>F#P/;)99W8"H0B9?"DO?>FY=UTSU'^0C(5EB48"[HSAOI.B8?_'VJ_EX7U
P;JGQWN3DRK^=!I=36]P\,)&M<U]EE$7-- 4!NL(NV<?F(;[C;?TFYCR/2[_X_.[6
PGX^G'HKG!)S?-X2CWF812+\H@DE?.ZC?U-E:?V]7"C"UL.TMOR8GCD&I7J(-YC=5
P$./A]^6H%Z7M'[ 7W(QL%NLV,X"G<,DCQVIA0[P258+(J$QT+PH2C4*2)HW$7"<Y
P$C]7A)EJEE3GAH9_NS=,=2/;$UPE0"_>FH.7CU6!DR2*BFO1Q)O-:B&35\>L%8_*
PT.P.??9NY53"A[3FU;^QH%YK8!Z(K'H!X^Y?[GHHPI-:4&@)E<^&#D3CD":"#-XI
PD?EV7(1979]R^_R?9ESG5&D+CJ,EIP4"&MUXV[3C)6G5( !<3#2+Z]3,=M4WO(G9
P+AQ.@XA7?P)=-7!7#4YLU:+N$K[,_>-&*A,S[U[$/F,7*"P:[4H(A179X3[/\5)7
PL%*=NSK\_B6CYM0)03A&U:?U8X0H@CQJM [W'\H2*9JVVBUQ$HT MZ?DFEH [UT_
P#/J.7^:J[I86D"?SRU\RU;LMM-@YL+K*^*'C'*0[SE";,,PBFX5[8\.N"MCV/N_,
PL+.\';/"#U:;,(">%'X\K>\T:9M%IR$NEZ1$<0#_PXAV*[ ^N![)M"3-/?EFRD;;
PR, 2PO"9[ I!A= <H@EM /H'P$*B947;PY9RK\<&<X\8EWS$D;)#VA3I>,I^I&K5
P&6'VQ!R,F8X O6_GOI#==K#H71'4ZN;U*J1ZL4.;G<%X72F!BAV6%)8KD')B/3T5
P+?LLF!-^IK2#I(]8L*#04.V#UY#J\UUX RBZ<X;?'( 7ZQ^  SQ+U)6I77LQ]3#@
P%HBR'I66Z*32 *;O;\?*)$B<Q7M:UO5N(I)&H<U6C@&1+%$<DH1S$6,('5'Y='($
PNN^_$' XD67NO?2DR8W%:XT&/1-%DI2HCM__!-N@@3/BZ*SNGLFY8-%/*#_* 1E^
P8I^=F6+[C6ZIW;YM:T?;"EXB<J'\J_INW?%W20+^BFL66O-Q'\%-,R-W^/!/ZD&B
P=F;.G8HQ8A3Q3]&(2+3]$G3IQVBD,1F U*/\HDD0'4 W>[##,IGXVO1S@.+!<2?Q
P5C#?H=XR;PSK*=T/#]HBYX9I)9GJ]HHT=6(">2TZ'+-)WAZL<FS3N_P_LTP>[LB 
P0V9GULH$7GTI45VHC4W#SO#E._S'Z4!>)!V&I,\)GD/J8E<='!QF!=,->9(&.2B-
PK1[990$[:OJ!,@C+']2"&QHMX!5?V/,,TWBUK@!6]@C$\$QS,?6MAVWTW>H]$Y<4
P('=O+'@*4.E@F5RSS&U/?X71EY5/T$MP"0@D11/@MF\++9 (YX6J:1:F03+.3HWR
P*W[3<4H2B)<4_%8F"1[24G_3^+(_OU,1%I^SQK9[A#3,;\0R#F=NZ5LGI!DB&#5E
P%J0PLDS[\V:K[^3 _,1,5X9E-VD,D=P4F G--_WR:,P>+W]:#EGE,BBOL<"^XWA,
PW8XH!]Q.MH=F*)]NPC7<&DD[;[TS!"+/8G*;5J!00#Q)8AX,]I\INPL+154BVB5W
P=>WL<0U?RDR+X!S;:@;#A<N8%'C<G9/9RWLUO9-Y8^Z_X(T0=)+"@,-6TLF];#'A
PQ)ZQ;I!.0/A)L_=C?IS9^=I?4_I#8"I8": !J+D_6VCE8%PZ2!;[N!5.R J,P-C+
PD]=O1K,6$@,DJ?G)QE3U]VKD.+B!(T6<TS%98@T0M3 1AMN;L@_7\3#+?3RB>F*'
P'G"[[.XCH'B@-@CHF\S(0#([PY8VK=M=(Z K-ADCT(=B2H;=D'%W1QBNI)& W^*X
P+ U*V5-Z('6DQ7)1&:(XO;#'F)6^:'>B0UT6>(6= S.TXTXO_[N3='=E9O4T")S/
PMQ-KB=O0M&@PKR@)F.A^<7.60.=_2>^O=SC13J$(? ;&T3.,6E<]M$&&K8$'>G#Z
P[),KL4AXP@8,8WZ;GEI9=S%O>TW_XFI#AWXZ2J"G[AK@@RMQ[6'*JLC!YS7$TGIN
PJ)&/I[Q>Q)B-)6/>K]9/KMQC6)-1?@.Y_PD>6G-G7B# =:WT+;BJ!!4/JIRA8)O8
P\:\G-G4"DF9O%Y FO#?MCJTL#75 P%.(EFPP! S7%MJ-K[!-,!6T.F#:9]]A:=[S
PMB&51#'XE$ZT_+T:9%NE6S<A)*>52!0A;P5CAT/08A7A+>9=CM"CV\ITJ8#X?<;Z
P&OQ9@0J,LX5?,(.1(ERX^N*+K71+WP[(PS&C#75+ DO5[-7+@;+"7:7XN:@V0<3P
P%8M\%( &P)M9(1%7.S"Z8UY9SS=Y.)DF]'K7,0.S4<R.&ZI"HZ22#%8$7\*T#&D*
P+>F;OE6SOOKF0[G8XV!P>K7!>VE2>8%RN2L/2A6LN5WC^HF2(AOE'"8FN4X"QVQT
PP_<B8?V+M3^UR#0;M7G;8E5HCAP+.JL<G?J^6/SJAPJ()#'CK'SR%]H-=P,CHBM&
P&;(O!PI2 <6Z!<0>%E8%F6U]X32':7_YC-67P:XCXFU%-1&;FU&Z2Q;GHS@OXJ?S
P1,L]X7KC9W',GP*E.;BYQ.&NOE0^":5?#>0JK@O/#,R:BS7"=IJR8)Y6V:L4PI(H
PNR9-W2WAF').F*S)X=P(T8Y>K)'PZPQ*46:V,3YN!]U9\RU-7,W7KHAQ]D-IMB/^
P6+;G26#HGTK(^T/_F2S21.1DFPT"?KMZI ,/_'BDM!N3]"-ET4*)!]$7XAD& K[\
P_*F&>&%JL>,G^"V2/OZ"_UW@%#YQ0)-/5;3IO <#NX':_P9_?$7:2SF%8S7TE,M2
PW4!!_&49XCNF7MB]PBF]]_(H5P<9SQ'\O9?GX+:WGT46S'X(RCJ$08)QUFA"+4F!
P6LS3 "[I3I;VY\V3G(MFY3.QZ1[J3M1(.I:M2T-<T."Q-NM>AA'LD?:KAMRL/4$#
P:7'U!:6+L$'T^EW*S>UVZPMNBLG$X]7<1PY61':!'9"NF^GE*)W?(1T24QML-WK'
P>;#SJ,UOU$DK^R*8]IOG7@Y^YJ6H+>KUB9R;F81<O]]')+4TV"'@34.>B8T-(>.;
P,IJ"AF@?,:6DI!6F9QA]KRX%=7?FNS;S@RW5OJ6T</4M>OF'M75H]5'\.]MCOFN7
P3/[79!?3[];ROWD=@9W3*9-[=N0^[O=>$(;[MNSK4;+_/AA 5YDX\M12&)=9&X$1
P*:]2G9="26RH("&!<83- ^W60(N5\-[]Z57+SS,.LT314(1U:HF+V#J!<>)/\;''
P= #DS)0->\JWKQVV-8N\FH9S>!HY.]K_L U<Z,/&[TKS;I@O,Z#[#J%:#RX,/\JP
PUBQC/0''>9X^7T@:@ 6TLF>S3S<)Y$<)8D0F4*?T"AT(>0):*NL,%MS5,GMPV#WU
P8(_Y-YV"3*;,1/$V(K:>@$,@Z; 47U$$CB5'N1]H==,+J4P"_9!?Q,F&#U*5<D%&
P!Z9H/0ADW$LIW=#&.;WK4+.#L&14*455G52$%JG_H@V2H#SO"$ $VR+KY6)GXIU.
PI2^2[6%!!!PHX!GB-P .MJNV=%48[^\-K];QE:0T%^0K7U'_IN/Z91J!5*RR>KLS
PB+_'MCTT?+$*U&$B('<14]B#JPCSD:1/'/[XA]:N2G]U4_,\]WRVU31YLT+D$M2)
P*;6:GFV B^%P M[4WE-#)KY5O[ K$*/6H)+\U>3AG?)P.M+NF*O\ 18)@?BJ->HU
PTP_I31[T=.>1Y?7]O#2+NI7Q#7ZHK0Y/?&O_8TNMY\#*Q-%!"W]B<AG6(P&4OJ8;
P0*_2S@B4BD$?9/I;7?B3ROK77]8^6=CZ1VJ-V/P0/'1*# W <T-,$V?2BPZF*+.H
P?E2@#R47(R;+VTI4.0GOXT4B J>Q*OO:V@Q%0>W,8J>(R$(6FRT 9X,#]Q(#X,ZE
PP_XH3QB59[:]K)[9I.UF#-/>1!D#VE&7SMQBO>/&0OP$9R*V/C]\FZ+4Q[8R4OC@
P4+'X9T"OPMHWZE/UWDPK4QD*0O[;2@B]C 3*FCW2&R*D.3QUM6Y8\WQN>&_F*D4;
P8B#.@Z"99GAV4D,0;5;E'97$^+Q@M9$H66^*ZACEK//Y@ZN>J%9V213]P(J7PV0_
P''X?\7ZA_DJZ)1PM"[:6/KJ^:;/9W>$US/K%'6Z/"/=,7+G!"0MH+7IV$(X?^J=F
PZ,E!E0VLC1\ _+=EI*BN<SPX6+"2+9&.[3Y1^.)E1J'\7;/;!*8?VUJ!F">8F^//
P_M3)[P[PF;.M$_%ZXFN]X>> O%R.J5??Q*C-L9TD]5'>SQ.3<J\;<,,&UZ:KBA>!
PP=Q[ZR" 3^B_9QV&8CJ[CQ<^B]-#O)O4!K[OXW;:C2+,$RUN7O$B%"LH3!4H0Z$K
PE_Q3K+V89%-W<G#''!G>+H0]Q>R\KF",6D)OIO8]HH+OJJX!"'O:\6TKP!&/M@11
PLZ=Z.2/$(8]ISC2L8&%"K"Q,[P+&R [.R\\F8 )[N/?LL[^<=P@U#Y=*]$_P*V?>
PP=N,M1WH#\G-S^.?T=*V<@3'_,B;*Y??JT;PG$%!]MC^)NLO0<KX(.;\8+C)[A=J
P@Q(:,7%IX-B#89@^05.W=N<&L^;YBD' J^=2%"4,VQ)WEQS&KC/:G_V3F%3(-W''
P9126CTJ#NF@'#&808_.%ZZ,9QL8DLVD!/447%GMFLDXV[=)-DF!IEW/&,6:E3.:V
P;E&"!DRL4O @2DJ\.)I?L2]CLT$BR/2?-F#@7ETR;N3,NF3=""B"Q$-YFP5G:3W/
PK]BID#7\M*S?M51Z/$H0NRM:NOQ?/:/I0/_^9_*_OH:;N^![?AUT$E#/:6FUH@;D
P35S*+:BUI#*U5^VCP92?4'"^IHNW#55FB1[>D(T1X"OJDI>-3&M#S%7/FMZ1<S%\
P,"ZIG@L&XZDNF$\?N84)TS14_DI?U6H85SPVVM0V&/!SM"0SBWS[!3>)XD&@4+KS
P@WX_";9UN7!/ %Y*C#M7$-%+#B&_^$ YRCF58^[7]IK_])>4N*D4Z+ED2VJ3E$(/
P#[[:ZZ274%.K'![7QA[!!66I57 DLM"YTJKY?H<EPW&+"%_K]_&M%=4I6&>J*JG7
P$XO/9^5,!!S0_-616K!TA(3;E/Z]]5-_=G2 $!) %\]^H3(IIPE.Q@*^F.C!G:(I
P4S1AWQ!QX)NT'T#902Q;MUIM?E"FX(@;7DP<:+AM)*?6[9\/1G^/C\J\CBS(&3J]
P&KRSV^X2FIN_,=@FE_OVQ;5W!TG5]MHS2+_-W8*?**NOH%W:@,_&!NR]]1OB PYI
PY0HE"*C>>?/.$7D(39W'^WP@0X/:G96Y&H'&Q# 4:B0$A&ZT+YX 'WU6.=$F9A*$
PSGC0KNT0Z%K$P,^T#V!_;0?^_Y+XL.")O(!%CXKQK^115))L9&Y6X?QH%DG/NR(W
P.O+R'";I2(#M%)5"=LK>7L%)AIA9LH?]T)Q5X,9/:/\S%!'D;I$X+Y.C)"NALD^!
PGCU4"D(![)58'><Z7>!RG8?SYZ'$Y_;UV7;$.#J+%&IK<79.5'&.R3802Z"1[+,7
P1WLX?JRBCO:-EMQJ/=C"@&"<+<262[0@>3:509.JI0:15*3<GJ@^51AP*(' TW-[
P<QWO0$62I2-MWY/!6T*I\'5')!+-@JGPI3M]*+"#]8H;VLWLY%PVDL97.1W,TC0F
P7T@O80QXF#!-2TL5?MJ?2[17!EAC2+JEO> A[KK#6/!E"OSUZZ8-,QB<3/RG!5.)
P]Q/FE=V8RS_@TBS2GJU>*:YSKY-!BF^(J]Z=#.$W<D66^HFSXWE0%&O")]]&_[CM
P'?NJJ8'M4QLMJS=7V$MYRJJK878T/H2;=:C'D1A:2QER'\/#:8 11JE-6F0^<TSF
PK0_[XA!V.A?H(+Z5J0@)3#F&6WK^JC9Q>,==Q ;.</OAO318(R#Y;6[&U+:II<RN
P"N&5%<#Y(_;A#^8'PE!5^6FW-8<0&Q$G .>59F-9C9'?0[&.MT:'&VA..:!NJ#>@
PAR(K^*91/&[@-M&?@@$.FR.B/MS!@?IXIMZR\!JFSJ5F>OPE H/*XB/I"&W[H)#)
P1\& .[<!< #4U7B%A*] K=@->BI1]7@.257*!.D"XZ#0,KKK+=YS3"+Z(EQA*J%_
PN?0KE_CJG53^ .7!^(?Q\F9ZWP'V7(H:IM:)BG_1=NW.$U@PP8]Z4*=E!0L:I+Q"
P48_%&"U#7=\6[IL8'!+BMSN$VG/<N[U<Q_ [,R=ZH#1#ZTS\).@=G[S/%X.1,<"@
PCT'[:=/'R3,N:<BRB,<HLL*3"\DL;CJ9-_4/+SK(Y<H_]-]">[U.U44SX4CX0J*G
P<8'_=T*X>>A^4[N8_"9X'@_J;+8"7-R1[%Q<M3A#:T5)K=V_B0IS8QF/L&_ /3D!
P>@IU!*IY%8EZ;ZXV:861/8:-H^M-D3;-U+P+C"<<B)T>C2>8<L!%78-\CQNU7WB-
PP1Y^>3G*>GJ\W4II&LS31JFIOJD-$F7H6R\^3F:%<DL8:EDO_D^T9I!LDZ/TASNK
PO7>\V%EE>='&(E.IGS\XT(+:^WI?A)4##4ZA7)W_AS$,27JV )HJM(*X^+>LT\D]
P,SD*242%E9N9^U":WJEYIQ).:L)6*'YW!;1,=5O$T'P_Z?XU4ZD)$8X2W!]9'.QC
PY%-<OL7]0WA4WRXN ^DH4FU?/!IS58KP+YW&2>1US_%D-$;<=K3TN(9^EU[N?8G1
PQ9PZWP\1K=@1CF^).@F21*H'2,TW2UQQ^C2>&8P,.PRG*\<VT]53#S06_.D.4;R?
PLG_'VA#@(5B[S9I42>T'L3YU6YK0%CS#]6WAEQWF%G-R/!G1DYU=)/IM-,C]430M
P&&AK/P5B(5-9X3QR\2.0=ZPY*N.':>Z^SH(FYJYO<!&3B>34%7MENW_PLT*6C7K\
PUVNA5W]R1?I[GRS3&PE-SNC/:$J%3:D^V1A5E>C$R'SAFP$LUBU/W$)E^G89#K?Q
PUY1Q$L%FG^]3A&[6T(USP,-^[TL%#L8-5=KU^<GCOA",59)<<)FU-/8X.1Y["D> 
PZ$DG4W4V?D#Q^+_F%7E)WALTRI$^C+B^LE/*G7,SBZ?Z%^R%D_F/^VB'1^#@E8I\
P#_E;CF'8*J*]H$VL"U@,3M+M5S=2!RGO  ATJ)X!-K$E4IF.?(O<A?[+0P75EX$T
P/Y7_I+7_3AFCTB;:&5XW^[C9\%RN*ZB)7D#1.DGK_]ZCIAZKE=XY)/KP!^.YM'60
PU2!:'BC[C%H+_[:GT+F7EMU#!*:J7N_T>MQ^G>A9.&M%DF^B2'H: .;2)<F8V*1%
P/TT%- *HMK&,7'.=@E Y$6;_HU'0(_9'J4M G@O&?<P=4&)XIZ(9DCR%PQ@5PHF-
P7((RTH.AL'&#PXT@3,AI_(9^_<T;6-9AG$U41W#AT AK7YJZZMB(5NLOO,HZ4LA_
P(K,C9, MIX/-TIO-P@-2,]52 =5L 3G\9ST33TGWD..]PS&&E*,U^9M=9--T'D;<
P'S+ZSRO1-*Q@S66P>I;2GQA20$XHS2_R*_5%^'LR3N2E$C([B/T_(1FLY)Z[A[2Y
P_]C^7256T;=2[M)>7V+=3-<69_)=&RV1KNVWLUK&?@*/V(SF=I;S>!S43B@.7.Q!
P&.4JLYRW#QN>JT1YY+93#\<UETY#:G $!6Y]GLV'\DYGD/EMT%H<:2Z@=3X07Y8!
PL\(4+EDA4<68;:_[;$*RH<9K DB0)G]["U "M:V0"C!!*2_[.<$%22W-8AT&S>#.
PC5+0_E88+U[T,XG29/C&4W[<HZ&$->Z4P"/J[@S7/9IRUDB",ZL/&"#$?,(W*TT'
PE-%IVYN# WG;Y NP'X! T[?5Y)Z#C=6![7!\'9-V:_DG$B@::Q3>GI+@>?08P(XP
P2$7.!$\XE:_@1VTL/T"0C_Z(^=C M^#-!/,H;NMA)RL+JAD?;DP%D<,6@'Q,%MJ]
P%A<+<P)RTJX2&$%9P7*RP(SV(*XUZ'+2>K/INR1!\<3PM=:C;LDS@)K%211!208-
P$;0=&AR6&:I'RH0#N@IHZ,<*-/\?>O?9,'RG1.>L<+T].]JI@6*GD^R\1:64\P8#
PQV6L>9)]EUZ"NKW=,:M7M@T? UN]<8>C=S@P,?V=OP$P21R;+S@2L0,V@N7Q#I"2
P,->-,BAQJ.DF$*54LW:261]'SH^[!H9<L"\DP=#^NY=-B)O)R>0"1,A<%WOI\;<M
P;T8Y11".?-97@@G1[W);DOA,2\3&,5>)W@5,%8N.[@";*/.+NPKPR3C8!@]5R$9-
P%UN^_\/ W//!#B0TW<&WKF3&F_N2(J'DOK9=8_-\=-//,>WXFIU5L=D1?*'4-;,K
PM[,A>$U:.U),#84=J#@'KX9*2ZQTC;=PF%X7-;LKPO=(B9 H#7".4^5,8.+>(O^*
PXS7!:'3 3RC-X,X]M0K@9-4=KEBD,#45#$MKE_WS8I4649DOMM]+"\WC/G8X"H&1
P"MC(WW!!3K.!RM#EL!I:^:+F L IHREEVT8?""\!@YE4'2111E,'(C;$KU:6.QHM
P+=XIU,:]X0T_*Z\0E@%ERYC/.Y&4JC?K]P^>I/:D%N9X8>;)G%8]_!]<N'49&ZHA
PY945BRP>Y,N5.! ':.9G?L&+JJ5!W%-^W;NF>XGP;=,\'%1AYFX+Q$_P+P@N6N.F
P^J8AV]YM]EV06PIM^5:Y3';:H209DF9^AB].P)=+UFK<T3%+,W#;<O2$Q2!S.RR(
P_DY:(GCLPBY[IH"J:KB)\7\76&*].1!;)B\4?:A^L#E ;S'W)7:2<>KVY+(JWI38
PCN!@+;GTHCW>+V;_0F'NEX@IUE6#$Y__42_,VPO.A=XJ\,ZK[4$M9DISKOE"')VI
P2;R9_KM/K[ 6$S,36@_#IZM/RD@&7<\[R2_Q:JA<1T K/ P$Y4(#!_9:3K7".S_ 
PW6[G<2SK_%7RS$"B50;[?3_$=3%I0+(T*J_,"F3-P%X-1H/7(H_BMI@/;2WLC85$
P_W5#VTY9X[FL(">#1!3,78X@3FS/Z:_D2S0D[;*[:$]X7?^?3OUC[? I*YV>Y9B#
PBX56O-,D=&9!:/>^H\K6::3*U8V#'7N[^,A?07A=J%P$SM*^T 1V> HWSW:LD$FR
P:VYI69KI"-KF',FYK%]@4JP*:DJ?B=/B,4Y";\]W_(F^>C(F$2#3V\?D2,0>_FK/
PI9/0&GYY%OF 6G?!(ISJ4)ENBK#>X>)23U7F(/?<NPB'._3  ]?M1W8*'V\M+EJ:
P#\SUT<$R^O5]O$[2KR0#+TF (IZ8:7L_>\D"6RKGO]'^F@<-G@3G:#=.MYF\UA5/
PG2P^ I0-UP4;'+%G_9K<X"T:JSJD<E2QZE'4XW>C8T2=P^?3EJYG.6RZ*&_BM<  
P/,I7FP&.B"DR?;2:Y7_M.@)Q;O4%?P]K8+;,9T@,<LSHW1#S@)W@^6.GDH_@(!\Y
P'\C:)Y1+T#EOFFV/PT4&WUT++@R95D89X=ND6:49.Z%47R+W2=T6"'(C8-MP^T81
P\\Q6P,[:K["7J^=7<@QY^*F)HQD DDXU-W8X\\0H*;09*=V?)X(\%H=/-A_U_/<O
PL?.'MU5NHY"AP+K(3N@+NQKBS!6W$DF:**=P@WD9^TFS0)]J?18V1]:8;N+W4I!2
PVL-?M =,;<[L@]XDE1<[':@E;'X;^F@-;)*&,.O(7%MZ& #/K#'9Q]3VWP2IXHMI
P<3M/)H]4DG3_>YO<%Q$J<5W-$1-M;-,-N38QB;0)MMKC\ A^(]N#MB[-9Z;RM<X+
P..$D<1&O_:&8T7L;DY1)HI,$4'^/H?6W=+0;,UX6#ZK!( 3X&UZ1W2RT3R& %?FZ
PLH N?<7]:32=0'K[+L:9?>!PT<UO]85XG<%$SRO,W/OG'J @#:H=!MH/ZAVM[*17
P7\%[!B-@5MFI&,1\X,X1,K8B>6'.R:<)<FUF_ :QE/9GYFL!"+=$8@MOAMCV=#%@
P232,D,':B#,+S71-S1W=ZIGBU+JNV2WOEXT@+LP5VK$LN8@7?X0J_X-/G76'Z^(R
PZ"0?AW54\!WSBS8^WYG!X/+>4Q379'/<Y1>/Q&/V<03-MW^FBRBK:D)N#GB)F^S"
PB>I-N5#P]8KI&-C_I)<6SH=W=D$*H]>VO0;BM7+DP&E(30HWZV ;P KV05!3E>5!
P@2\Y5?PW,;:B+O5U!G[[&3E(,YN./\WVH.C ]3"-7ZIC6(/(6)6"I1 _4IT"=T;U
PN-,=FKFZ;=29,26S+9Z"KI8X9<.]SU.3,2W/@@_>%#H&2)3$A2[Y;T7-XD/-G"!@
PD 38^*9[0W)L4A&$(&M!4)6[[=\U[[1>/*SRMIA@_--\9<P& +/<(DQ,/X#J@&IG
P_'"].RS3B?)86 4AK-F#"_%V3.SJ )EG0&5NP57GU>;W-D1CB[SDV_^]QW-Z'IRT
PW/8/RBDF#H#1N8 (#D$RM&7R%Q^D7!",KP7K-R<I#\GE42Z!4ZWI/:EW5GZT"W %
P5V?& %<*8*M"E+R"#H?8\ 9<9Z;SG%HBPE:#9?@YXA#B1E$V>2&VI6J]$GG]S;P!
PA$2XWY1<@X-I@+\5%@,,_YO$WD'N(CQ;IE<P(T0DB!\:"9JJ(>J6D(#%ZCL%:TB6
P:17N_9ZX]XY:T',Y_,KJ^46FG"<Z:^"W3&T>>9B&Y/2>Z[U^N.[F._O[S$*,'H/W
P'"?U6W*6EJ[=Y<#+]\ "J)XM09"5TM"8>))S8#B;7G7!^-F0"'C''=9!^KVUG2WW
P28!%1[X^.%X)CD$!0,E4SY$BR=F@T6^NPXB2DR:9O(JSDN>@:8&X8NZ(C92:!GS)
P+SK_Z@-O$Q<"%R))0GJ$'"JP+IK5$;GPHZLJ:P;[\]*OM]0IQ,9U!T,M,50IW$ZJ
PN,[U%.ME^OV6S/8'>5CGGZ5?MGOM)FT0RZ&DDMT6@7 I4';%G03(/COA*'/[9]]%
P[!PY."X'G^6H9F(T!,X5$@T19J+B";BP5+,8TE+J GDE4?B-ZB>MI+9Z_F3,(LQN
P\4ICKSR;<Z5>5XTXD\K(#UG/*'-B6OC!)8FC$RU-0+EFYZ[6NP.K[O6P:YG2D,N.
P@;L(5@9-F;!NN&!=U58*8(Z=(>)1O$3YX4TTIF1[#39',10DAR5:SB&X]SFNF6:%
PUEO88%A&7UY2MZC2E(_>^L7\[Q_C_>R"'T%*/3 NP/P1S:Q0#E)(9JKYSK_1FB5M
PLV\KK\N]%=JB _>UERXR _@G)78=X_U@.PI)%-J&T[:&K*P:\UC+Z+0<3L_-K6T3
PH*>;B3@KT]+*!0321_N@\,.'Q<' @;#VB1RDEF%'=4DPN /44<)#<7 72^<$IFPP
P1&H!P];H;1I%QL&;"S8_ 2GA-57A-RG-M80[5&X.;8FN'N3G*Y%<^X4(NK,3-/!)
P6B=[,>8OM*2[F^>ZQ80PL#*'DRE(;MO.<\5RMU :^J>N=*H@!?D]^Q%PF#K+[;D7
P5,$70Z=(CE0>%R&- *OW_E<JQZ9B\O#_(^D4U@\T=#52BLL0[+HT#H,:Y,!D?;<.
P[N;.BTXR*K>=68)02T/\IB:@9W&I"G[:SV<:;]]NH$^2MD>DRC3I0XKRJWB%<YET
PZ<O["I94P #=6C?@,$HG-=^1>QGN*2AFP"B0ZGP1E.#FG>Z3C%4YUJ/[N"ZB''N8
PESW,LWC\G6ITIB45*K[NR_.GTU,<27NS$R#5X7@JI$*%>+D$:RLD+)1W!6Y:J5 B
P$PM63B5^ZEI0KIPVE'EX%,3Q8T=^)50A'UKZ(FVI+N(O#V5H>H&8G6/OA1O<?BH4
P@%^K6'(BC>>J-0>@QN\/U+KL:.K:O52+^P:SZ9Z%9:HFI$^\!^2Z*(X'_0P'RXF[
PIM5$X,*OIAHS2!I2S$[DE>9OKE/CL+&3JFWLS+%-:&F8U_[WD6HP(/59T/])XKMD
PE^P[%[:\=TXB@7XE,\;0^DETUZ*@Y8A 5U)%P&?ZWLX=[HA>+H.H$;KKUR.8G]R5
PMV6AH:0%*CW9ZV<%_Q^%[CMHO>VRE/)B&D1K3U4>=>WM5AHE@NC(/:*GM@).F'=D
PEXSZ]+-O-'Z-EAAH8M]J71/:YCK=,4R[]I(@8/ATD;O;<\)B<[@.2^N#S%B=/^G(
P$[@3Z"S:D#C*%8:;S#07X1,47FF(V9ST.+C8WS^,#.-)L1^:2@'WD[4<!#+_8/**
P/C(U\ST_EFQ)1(0]IU%5:F>U$WX1PYZ#(Q:][0-97(!R$73[M@9&# CHA_7Z/+ "
P*1RAUXN2#["<V0484R=>/^U"$-%;+UH 8?Y"/ORU/ (GG%]6^>@7K$J$UD+G3)8<
P@:$:'0/ZNO<*G088*PT3]5Y>J[GDRL%0W7[]I!K(ZGN1\%J LWW9F #J%V='U'5(
P3VMOAVFRD.<P%42+#_1^VS]?Z^@G$;IP4EJDQ;VGNH+&$"YG3G\O==$> :XT[$/-
PT<(+$AC3+*PQ(4*]1UT7RV@1K-R21 ?'_(U^(OS7^L42I+H DW\W^[C\)Z]A*-[I
P;!XTG;O1 /LA'"M5.<Z2+ A&9]QYTRTH;02P!B?4@)1[6W7X"Z8W>H"4X#UP7_TN
PSC52X%'BY"3PM8C71/@RIC>T4 U%WZZ5+ :<]6I]O&LP:1>0=QLF[+7VKUK:1C\P
PXHETCEE(AI\IN=.7C%[:6AN=$M@B*,V.'Y$T=JX% '_7/ )Z4$E4H@1VM;N<N%\9
PVQG.K,$*XYA8+K<\SDZL\9VJ1SA2THO3&BH+R@,AO.O$/G*AZZ@'TJ7:$ >657A0
PX0\Z1<QI=Q]Q6FWX)FFF?/H_6C\F-L1V:,0NJER*9O60C?>TK%O(#*P#+3HQLH6?
P/CMF*0%VV*H:DNR[M'JD 8.N:.6A[Q.M93[0@_J#U.PG 32S=&*TO&F5^HJMD 9N
P>,PIA]U0*DP8_>^A5,[?]M7WN"VGF4/&3@CEM4V"M?'5H53HRM%"_5VDM0$H]4_G
PZZ$#949</-578NV%:&UTJ[L1>L<57K^0]G,#4%UQY&?I%D ^8@KP'ME5=Y<(]X##
PPB>-W'V*VEZ(4,3V>]L<9-38'@F8B[/K??'*= E*OK8&@>V%>9/DRQR$\B]I;$5^
P4>O[LS4==S@O*BR7&M&/B=A/6#)ZL_J&!&75%5^MH9H=>^7L '<&UI):**O:G_Y5
P(9[O#;X D0-%X@P;U5T2_<5O5DGIXFH>0W-'P,V0+ _\I[IRG=ZPKP9:7HX<;D80
PLFM(0(?NSFQ1%J.;!0G"^,3&31 0'-05 'A>C^T_XRH I=28Y([D@> #7N?3 6)-
PFK[9S/1OMX)AUVU<Y!]ON@:UKO+,+,E<E%:B<18;OS.76:T6"(('/D)$"+L&51F=
PEX[G>7>X?.6('K#D8U%9K0*3&=^UN[XN6[WW08U9HFZ,@\W1L?346DU*&[&'\JMM
PX1MSJO8M#M>1T[FPW[A\]K#+J?L@-4/+9#EZJ4\Y>^0WI0;8=FK)&Y]M T7JPEV^
P$D98*ZUZ_YQ*?O*'O+^5H&2;Q4GY_I8]R($CGK%-5"+0N@B]8?%%Z$&^">J]I('.
PD?>]2P\<HTGFA^JK!_H\CX0NX^[^?<X51F.7R3#(Y*PY3+FQ82MIU1SK'3^36U),
P$U@>,^%//] :>EZN\\) !HQ-$HEV\MN,#U6ZNB9,2ZHNUYOR44.?1A ?;#_#99T=
PINJ+/I U@<R-4)L'#[CL=]=&YZJO2OJ T\8DW8P\9W2ZHZ5F6ERX^A'FQ0UCHXAA
P$%%$S!9[6KO'0(M^UJPRR<VH) _T6XW4N?7:MV1!-T?7]V$;F1B/ZTY;^R37BW]I
PF#.81&Z[#1-HY= _\'3<5C*B8\Q3P!WC[U]0>+:W\?L+5("Z,L))*('DI:9:U+ZA
PFH2]-9B:4=/GE ,;#&X7AU!<Y*!&8#,!OL'G9YK80I6O8AWF&["L]R)+$2SN&[GQ
P!CGGZ1#,0XU2K-^HH1W. G;S<A$Q^W,@G*FX8']H9K5%1M \X0<6=A:DZWQ$:2,X
P*=>O$L'H11(!OMPA7W>+5>-<=+_1U1MKM1%'4"W**\TX//<K%UMT+9A)<%I,;+BN
P>"*PSQFKZO#U91G6 E0YJ]659C9?<7_/5W^K%=O*!K]=1@"I7V@WS?1KB.W>#^U2
PFFM V-0SA(64Q:*-:-3LO%[]M:([6I16D;3U@L7[I6\A8CBK"D)#OWB1;X$/Y;,X
P"W(S:+K*#G*@'>9@O6.2\CZVP4^L+$G/+G[[DVF%BQ+UAN5OK:*B/!Y+[8GO#+UT
PH)SW.-<6_K2'.%D!=,F(:K+57T%4"=MV3W8P0*IA??>8I^SZX#M;&MXR9CE1.*#D
P@JZ2Y^ =E4E0@6?9N;\^MR(2NX%5FI?D$MGRHNQ#]V=\0><X&T=[^G5P!P\>CI!D
P>4A=L](.<^EDFH/ZTI$3P2-!SFU.?7 Z8K9X),P/!)87;HH=F1:J4T9:G2HY-&;7
PW]W@*718M'>070:%<28,RU:>$^O+R,N)7J&;I]*H'@^FMF<HO0=@Z)\@JA(L(S%L
P60E0-<#KE1Y[PRF[2B'8KI*+,<2W-K!G%NY8KZUV^T12/D'HU*1*40.:Z/QF-JDX
P3!%8(QG;@[2HK/X7-GO4X2C]M])!9PIZV$RHW2*)I>M]C=5!8:4N48/?0OYRQN;G
P,@;.!!B(!)L%<!!#7Z!,^6%+VR]Q+O&D:&-K@!%EK=TC=V:;YI W"?,3CC53:MXO
P 0H$!YP1_,F%4[79Y'F<Z"A! -A97W6JNG$:B$W#(G<=P$LR+^F=M18%^*Q/ V+B
PZ[2HLH(]A(<G6J4,$)F%[$=9X*(S-Z:,\WM 8)?^"ZB R%XYIW2R<:N#YL?8LT5C
P" 2DU+'*G30L9!5[P,J^6..<&.H>GF^D/EK6I1FA&.1O8V371E#IYBQ&L <6AU(L
PGZ#K(3R":R E3C"6?&=O%I'E"52RL]E84FKVD+B]':]=R"-FY )6[$2ZE@GA]RPA
P/<N7MMV5L$2$P-8@>3=E"N9J]Z/]JS52?N[\0A>'WK,-A8Y[PNJ#BD",F"C*OUTF
P=[!9 0H7HU \?0+$TPE8_YZA+'Z<(5%EL[DCB3@%X]%,STJ^\;_L)G;0%=@3%[R_
P*,UA%;I/CHKI ;K*D.S<-$>;N\/ML@)/IK4+?:]("0@_!R0X'Z2_)^]?4][E_QVM
P).7KCE 2&84RPC.#16TQ5V>"V'[ 3WN.YC1F3UEH!63O@N^6S%:QMV(/2!:X3@O0
P)%RPGE]EJ>L.HE/6'(&J@K5L;X^:&/=C J?/6+ESFU:G;?;2<GA>$N$]F9EQ)[J*
P  NPP#TO_+*I"VV-FKX*3-:'[Y$.(1&>@>R*$6="7J 9+!:IS5H/2"L153+HB5@!
P7/;G-WFO^/DUSGG)\&BP3J]HM'TA1'-)V;INHI1:?<\,@=N3F!^#F%E*&%-6B_0V
P [\ 5CE1+W9ZIB<L0!1#XP@KF6SXJTS0OOU;\5[I(QVL-6[R_19'/O+.S],L(.R^
PDA.["_I)CA47SSN^V$/;C#\UU,34*C++E&7SCCZLD)-=Z[:G6X!47_,Y%5&[,AXR
PDH-6J/39P$% ITBQ96YSZ6.6B5V82-,;M(?EQ/31"J;BMO)R%>Y67@I$BFTY$ BN
P-WC'/[KOU&2"BRT[UV D856:1S2CLK U>V4+1P]"?^VZ2(7,P)(),?.,D;F:4O#>
P\E9X%U+4(!C;=N@9,-F!  TF]/0G@>V(;+CI/<6C+]K!C/PQ]6[Y^S!M\Z^=[WK=
P7K<A2MDTFF2?7M*7/[H_M;QIH+UQ4W=KUK$'5R_ATG0M3=98G7ZL^%A>P46OV0V;
P\AFF*W>NK37(2-=/UC)?Q.K.FRPI#^ML\Y:4UPWDU>;31CFA%1VTZ,JR!W]\K0EF
PBGB(<B6,4_K.6CW(WX$>/HH(.E&@UZKQ@YO8Y/19-P4W1L]T'[R]@Z,C=3!I&IV%
PX7D[IV&%7GRMO9-*+SVHEP9A@1BE-UG0A>RF8X E_/^$'<]C6$%#N%(#-:8 A,/0
PQ9989D-<5J,P%[_W<4Y-T.<,HPU"QNCN"WS=%FL>/'@H-17>=Z41>O'C1="C>EL"
P.O31)RPU!K.S]Q9K)TH!.:T+F.^Y_-7;I\/"4+LT*W,8 U]@5R?__;HT0I]_T@L^
P<22WD7.%MA>VJ9/DK3CZ^K.Y+')- UX%V0+NE=AEAMBA$$_*BB<':[':*"#81:BN
PUG]Q>Z.]"D2#"<T22(+=>["R*7F$O%2'/^[S7[&??,ZO$"ISZY*OG=5IKG.PEB<W
PCX!/@\-#L?](!-W/TYGLR?4R&!H@0&ZL6=\W>GXUO?X>IO#&.1ECLYV+9] _PTXX
PX.0&9)N\<)7*? 9[#-%QPUHY-+0\T34P+(H#0V,K:\FQA*.M3+&G*YXOW">&LS\0
PE-@W+$HJ4^?MV_,ZN]PJ4LE)OUGN&Q!@8Y;V/RF 7TU5L=D/K<+$MR!.K57$XR/Q
P?1*'#:7OG%QP!BD'PD#F_%(AL@Y_4,_]&S86[<K3W);=-U/]<D#PX3;'M<R,);1N
PE2A@X W' &QO'AJ_ANW-&JBB<[#"V$(I=[SXX@@N7V*FY]_YE(+%*8KNI3PFQ,84
PL'4B2'<9N5A%$W</*^ASG\@#4(0!2@S]B,R8)8$LP)M_R!_'T<OI>MN>J#6,A<->
PUBI-CGD_'E@R+":I2]4S^<7 19W$$HKQ-"MP_GX#RA, .#BLMF\R6Y 8 Q]N9E2+
P*T- ]M;F*X:OGY\KLGA*A#3Y-0PB11A?,.?>7+"?XC3*&16(K-N@+T.AXP@#!_*C
P*^U?=_G1 [TX5663;48^R\$,*D,=56F50Q15L8$1Z#BR?0Y:Q;S\=%)!W\ZK]12/
P-N#\]NM;63.'(9J4Z7 .?X-*33]"T*8BJ#_1!Q5K(U8?[1F/* :L:_&I!9QMCP2<
P-F=%3L\%DZ<M\/I=98+9X\I(*'5K?</^0XS.X5X :$FD2UQD[R&)'].L_Y'W?S7R
PO A9[EN,@*2]I@D>VEO?LZ C]FND';]]JQ7-7+J'@%KTLXA^P *!'"F!4M+<X=F0
PE6_X?H<J.$4\+.*7DGDUFUPE"X8""5-\FNGW9N\TSBIXAR^SZ*HK;_%0C!8B7BI9
P(KY-XLXJ[KE-K9 *O/*R<D:>"W+ />-\.G 1F<>*J)7Z2P@!']C.OF0HR7PF]&B\
PE1%"7GI#Q/_=R68A* I6RTV8^:<YPTS\5X40AKIX3]XI__]/R9021 E3 L7;O!: 
PM[G,X44);98.,XT,-CZ_=))*3,ML.;#AR^PJG;T5RU%$[H^W(4F!0:.#N%)Y!XRA
PE0&^P+L\A(9D5Y:C%I HMF0%1;]]N-Q^$+!Q<P@@&DIS61>^NEY&MK3!8GUH*S :
PA4OQ:G>N2.>%<)'T@ S-C>G(ZF9KK^>#LND=@)"/>@'8EO)9K);6J-C.E7IK>2L>
PELWBS.N']6P[\OA!>IO-C:7"#KZHK4,PH!PF[GE6,)X'&74TKOE!./!..C0R$!<6
P0A7A]6=26D0^,.^9[<R[TMN6_JBJ"V:,N-OA/C?EH: - -+G>9E/AL,TO%B90H%M
PM 5C5;:A%'3VOJ=!JQY&=7OH-M5%AR3['\Z7? FE8!VNM5_1T1<Q+-;%9!]@:O[+
PY^]:F0@:!27>,[!&R8?  M]P"JJ7-G?W@;7Y\X 2Z7\ O-=,%;*=T?0#1+)?9^>>
P8RZ.2(O%PC&?M?^D;/Y*<;.VIA#10HVZ@.%]G/#'52@YM!0?7/ATQG>#36):O$Q1
P0NY9NE#9#RQSQ-JSOUA@']4NI([8Y"Y\M1GD,'8-%,(TWG!P@WU\TTD'31(T]F%B
P#X3=N"<OX^1Q9Z$T<,GBTM=9KF35R\92\19IEW[RP>U4$#@K_W)]\@A7HJ[_H!JR
P5JL;>#=]((V^"3S=P],&%ACR%."[I,ZFCQQ*R61ZT3^%9IJ4 (OV-?5$S97X[K1&
PIGS98C[ ^=[Q6ROP:)W^KTI$:K['#*MV CZ(JZMKR;)BI*D-8/[3@%#O(&L,<;@"
P=DC*C>F*V;2P6F@T=66MXF4B^:H2_55UP6RS!4#STOR?*:="%7=Q%BQ0P?VUH"LV
PG+5,:GU>0AVK0/O^^*=3J_S??4-^J4"^*!34[(E()?\A=K[6V;J)^NP#QE?Y#Z9-
PJOX$T8"'<$\GZ!;[(8BQ'Z(P\KCNJ/=R-7=ESE@6*C%H$99$L='D<3[>N )<DI=?
P"!4>N&"KDRGPJ%<?E)82!5Q/+!"U6R[:+MY+"3?]SFLG]R"FD28LC 0@?#;ZZH6>
P4Q <9-\G "UH%)"(1XY_ "K H5$2)%VXV($G$^*.[W=N"D>L)?(LZ=N"GN\0SB3!
PQ< ]^G(8&]"0;CVN=^NA>7YAU0>!)J4\X3,XO3;/9YSM40A4VM"3=D"5:Z2OGV/L
P]DT/Z;4HKHKXN4+3+D/X(A5?Z9QR@&KIVV)>]NZ:J'_Q#2:/.Q+A,)I;8VN]Y#Y1
PJA9"QKA?\1'2,KZ)/>ML-Z?6+)[4,0&2W0YU'S4L,,TZ/SE]N+@Z]52U5)M,?G=4
P&Q\B&C=D.XW5[21@&MY1U_1+$\WV<5]&DW!<Y,587I)Q?1K(L]Q[3S# &Y4]8W(K
P.[D4HU-B>T"29@WL+Q<+UU0&BP44BDJM*SX)B#)E#R=M#7+P?MOB/,=V\.H.##UI
PGO>,,N*?-J_TEP_"JN.D(X_#!,>2DK2ACS-*A6C**'4T RR8*S@BKI]9YNT$'@Y%
P$'%,P2,TKQA\4[A&0T_2F*=^OS[C"UT]0=*%DLRMS;X@\SD%$!+;6<F0>I%6=ZQ-
P/=^KZ0D4DL!([%KK_W)$.CYE%5&N@#M7?SY]2!-OP_;'/[K_YW2DQ#D#M;TZR)D^
P&B,SP!I*)4R/#KVK..U?C8U]3 NY)ST,.S@):;7HT/^O47M6?U/%'+MZ.W.=]O;'
PF,A;73]*XG'*,>H/)G>TEJQ%E\8><9YDRF9,BBB6A61TH)#WXWYTPQ2QDJ'"W&KM
PH&RKVKTX>)B^84,IP_/_XOU8>-YBB='5,U_9!Y"=GH@KG<;.2"+]ZFE;2O61K#N)
P1[3^(H=9:/E!S?#0Q2UF^;I(G5E9YL.C8Q*SE/@GUGP[B %,?>'T<=U$Q)5!@M0^
PQN<%&<^4-9ON/K')O[?4[!84C*9 +,*,U8V=\&M6=T<%YAC!<F@] @=J^4?"/MXJ
PE4,-YR/(P\I6T7(UN^;Q,('TR1BIRK+S^F)Q+CX@5T+\^R&4A[FR/7E[@DX9"0[7
P.=<RT>V":L.5,G$XDE_J9JZY@N-1@%SKN19]5[AVP*Z=H:&_VD->OF9K5EH5YB:;
PPV2FCJKG^#LGDM>W]52_3#*B.$=:&G%C,"T[9SY.D[5HK18 ADB\SS D8N [+#=[
P;J86"'-IR+A<XU=:+,>X%CB!3I1X@RF:CE.O@<"B%%.H_$NDX<G(O0W#SY^)W-N-
PF(H?H8 9M2]A+W14-,_5/R*Z>50P$;=E113.(5(3[J&$L2"1\$_ N0:0M(ZV[>LS
PAW:), '.O-6Q&:\356%CA C2Z&'>!"[ "I.;$J)-S>O')"\:@$Z=J<G/X.'X,5/E
PB,NFI/5^U)>V&W\YKE+/V39_FKIROEL6O;4"5;B_!P'7FL68$H?]G!2UFXA^3M**
P,VOY,P!G2WDN(.TOHP"+M4^J!2] I@S'NEU0D-2W)0OX+',D#\_2@9/4R-?5=U-"
PQ C[@HE+M?'>7U.67IUU ;8+0F7 \X1Y5TG"P""7)^*[\AO'@RKT[W45)8K@?1EJ
P:?#N@V] %V1M+6 Q2?/EB.-CG&#F8I^F7[FPK^Z9K5(6!#KV2[\I,@L6:H>&/ S-
P5J\9C33<A(QTW@6OJ(_.)WB;ED9*30&*7\0>&CDYTGI&7&?QUSFC2(60JD0+T@YL
PYYA!@8>KG$VE,.)_EN)KB<2I#%,G1PR:G:<S'#TLJ+Y]CYA._X+(G]0#6&$+,^'%
PHID2K=S@M6K>;%Q-7WXT/LYMS>*F^^&RD!; 6ZT-ED$1/]5&7*\9&B])E^MZ3[J?
PV2 H_I+*I^+JU^&;M[S]UMPB<&*E$+W!*6G\2^YH+;W6.W<80!BT2MEPGY(#_&%L
P[G8.WQ\9G_G2G*N3?F>B,_[^.I0F]2IK.YJ'96@0FZU5#'E23SSH6ZB ,H7-]<?6
PPB]9;^5@LQG2?YL%GA,>,YPO%]KM-7P'[G27;Q"8?"W[94!7S.?^5:%P&M)'38&)
PR^=Q/*1Y9Q$86"QP-N'?^(YTK#\8AOA;Y0]WU5:80UTAX(4ILI7>D@6_ "PN_M-&
PCG,$?/C06M5,B=,M_=.K"Y(TC3^ ,KO7O!7[T,^:$QI;,6V99E&L-0*J<99AA&KM
PWC6?-G-O7DP(_+O_.OPR["O-U/<*!QX!A)>;6'WZ<Y19+FWX_TU00$O#F@952\NY
P).W(?!FQ8[J\F7SL!"'AS0CB?28$.U;UTJ>]:4!;'_*T$UWW_^E)H@RAB1,2++0Z
P\L0U2]>Y+?;XO->$_U)>\,S4VMN].%JTGM>E?&_;%?[75J#F]^:% <OT\&U1#"AD
P/; 1+@+D+-=HYWH)XSE/O(JX%S@%4%X(=#EQ7GPYWZOJZ8^[B/,Y@="ODT[?4!.E
P[3#U3;@=,#=-BP\,]_.)\=UH5@*_,L@(0 ,P(MP0NW!JQ!>)%#G*GZP\U3AB_3=&
P<&J5-CDV65;2#UB\;0G<]4Q@-7\ G!F;[:^I%WNI3E*#@BR CY-OHS _:<J%S#8]
PMUTR[_P!%QH^#>8M&P'/F3Z4UO!85L;U E0%RU+(D33>X^ *O 3Z6C'ZA4[WT=&D
P'*EHIVAO@LI?/R@!@*R?J-7QI+C=&1:KEW[3_4-+%Z8$BUF?@5E'8XK;3$\ [Q8L
P>7LKFLB+;'F&_?,:W8S0V8+*3024F09<]\I0GAF<!&4 KZIJ"\<BN$G''[1(PCZZ
P4E^:*.K(E5!_6U40^N%^VCX_ZFIH:_:Y,(#<)%H\")K;/NG12V*5Z-;$#&M;9T_F
P-YU?5C[)E[!0%J\+[7U9H#$[20=<'I]Z)=3UUI98B^2_O[HN6!M?A7B=;\<E1@3C
P@WXE<FM18SWI"*?3Y#KH >!>(@O=$!*ERVI&!8#B PX1;=Y07)(N0FLM%6)K:QV+
P)"&(I\I\7C#6./1G:-(![A<505?%E3(2L) 6@A_Y@3?IO%U"9%?H8UL1E^*4)_ -
P=:[K)G_=AMCE;6X(9P4946FB._\*<TN.B1!X<0$)6O6Z!<C58HFIA?KY@3V88L>K
P&P*8]+=+9[WH6*Z ;J($(JVN< F7)6SJ!REO/I,D,+PG.>SB;-Q^Q\ ;O<9VK-K\
P.U<"#.,,#UM90D$U&D-8YE-W86:[II4MB:.0+M-SOB:)=(?1@UKCW;65YQO8&*J/
PM?P>%#>X15ME#):P0?@-HI+VPI)TD[667E>6M=<?G#*ID^;(PU9""2_,8Y6X4K7T
P@2GZ.L5^).]@V@#2VN4B>7<",/</35\#5*Z*UY,]>6,0M0O \04%97GD")'NFQB)
PPE;@;I-.]0Q:V,6P3451 %M@8K^(!:$6E?ZQ /9[6&K$#U@OU'>^K4H6/2GA2W2;
P,^S,0"H05B+#%9.\^5(Z5(Z!;SJ$ Q:@)_8!;&<-UH7N2$408QRI"X#71SAF_1Q 
P$(.F;V&5TEL;H\;/7$*[H>Y(2,[&"&]GF+%%\5ONV>GQ#;VPIU-PM,3Z0N9VC@T>
P>TK;^--]=/K;[Q8_9[O>>O":'704M=3#7*B4[H10+?$HQO]E2\\9ZD9 !.5A:'F.
P"<* -NL(T*?BW;!.EP1CM.I<$O7XWJ;JA^>.AR=8H8#X)LH6)>?CM:&GAF]C1;4E
PXL>S<FM28Y\3[ '22USS//%K+,ZI'7V<JVDJ4** "U(WPQ0?^& ** &,#_J$BO -
PEG:,]ET75Z&-%3:\*2@VH\SAKF6EQY3 D4EXN"FG;W=MNEB8'=GX5C@4=F$@H=Q9
P5V6<061?0$%B$ILQ$)?>@-AG>L;PB.)2V(R#'\RW,2QX0_+?LE@T>.G7?-Y6K;2;
PE'R;R^(W%V6 _'?I#:VX/PE_=#LUS[;&%B4< @_AN'XA30F10P=KAROSDSC[]/(L
P"+F+:&!Y+XGE$,5_9CIRD'!_(7+?D$_'#9.?O8TL/.('&?1-5ZQ((^R>_:O>A@WP
P^1R4C$'%"@[SGHX)CKG<_.L5;@HKQ>285&HEN\E\1'_.I'5-Z-N\4"^")8+,=[._
P)^-H6"M^>^(Z$N5_2,-KY1.-ZCY)8%YNL(RM/V0!!I8-APW-D?ZFG88+S8,]VAC;
P,Q< LAJ$3X.I!N ;F.CLRP-J*@[R=@OMRG#+@CNUW<AP=]@E)4S$"8"9_$E=.K!F
PMQC'4='K@]JS"..%Q_=&D"Z)4&2*;@N/5X[<FFTTIN2'82J*!R0B4FOX:ILTJ=KI
P]F <2J#47-G@]),>!DX3\*.(S08/5 5@#6OCP?G:#(&I8'?6)"X8,FH8!/KM\[(3
P3'O/(B\\U'6F2VU6]9RC.W\M]ZT=+[,(5?GU6F =YM=K6S6AY+\!G4[=_7B":?_"
PSXFX%,C6B4&3R&(67NI"[KM%Q)G=?!V^&)L)<&+FBF1?V=6'*@(SGI5[5G _;R:*
P=4&:2*\#T[E7/((6B""=QQA1#P$05"J!:*[=OM_V0?_]- W?_9A_#!WH0RZ:YJVJ
PP3_-#R$!"MC\E_S3"! @Z<O5LA[&J9DJ+AM^YD7WL0UX=8H 6T3?<)S5F%X=M;]@
P%0D%RDZK4-K$I43-(P,X1_/!P^"Q>$F!5_*(+.^)%=M)Y3GL27ZX;2@1X#3P+!]]
PY,1;17H(/;77YLEJ4I.2+ZSSW/7]L*(P_Q!4#0>CJ8)K8&_ 7<W'E7.EQZ9UK;>,
P46C/W:*=$U>M1F+04TG-16HX3+VV:7HZWPOTFN\ >"*S8ZA'KEPTWK#CT4X_RJTF
P7\S?$MWJ"P*@=8)X@43<W&O44M)OY$824X)3IA-]#>,[!*-U*%:K4*;,''/9DU.I
P RN0.HB,>$N@%3VPRN0KPDAA#-6W((#3+K.]IC3A (8@%:$8T5\6I6!U1;@9#9C/
PZ"8N=.&!.CHB/\:SN3%[2:&KA/&<M3$2UVNN]N@#8IER5I)R@H@CG:1A!'NJCHD 
P@;:TS)!Z7E7,^,3(Q+ZW96F\6816%PH^!7!'H*- TCXA&NR6+SF*2F.<\3_O&_L_
P&MS[(Z)ON0=M0^1O5_WMHLT<Q>^18 IM$L+ZH=E*?5\EH?S*NTY_B&A*&1O!E%_;
P,"]FWU8FG8(SP+?%%A2153 I%"KS719J'P'^_">IO:ZL0L,VIK4\KNH):;O6P5%:
P]2:@!SV)Q"2U!I#)[93\ "$?>""M3\?>,->IT%G)=WO(?(QP$S(?^\M Y7.HPW71
PTYK6B/J0%29K-1XJ.FS)CSP)TM9"C#C\36+(-7YB_.S1=89'\H3I"Y)XSM&?S44.
PB?HF\X2QR?"D<41K?]E3ZK<]R)C7%ZVCZD+U#I>MB2\R:&-7T+[+QX)(Q3V'U;(_
P;)'A1X&M4[18(_.%_H.NW28Y/.28OAER";19,+D!<7O="[=@QEJJ1]TE4#] $Y6'
PL[?4;AIK'#NUL37='<,@3(!%'[MA\!;C(HWN'VG/]ABW=*0$@1K\K/XC!0'_^G-4
P5,_]-I@EQG 40Z$K?_BR\/O:]-FP0/$F'+A<K<!+4-LAGK-M<4(V>!=8ZWZ<<Z].
P(IU/_81FU.A5J"B[/ LIH-W'L+L0L&H/RD)AL(YAI':](391UK@#]_V(;*WRN5ES
P+QD7%%%8IN\"9;$C08[XB.=J%@_T1LH-6FX6!=%NO\/S# 4G &>Q9,U>\X@^@^"2
PBUI1M?-PR=I F8"PO9X<X-3 ^OA^@7)VGSN*D?PI;,@)GK47/CG\QE &8G*V2X,-
PM/U/>)6%[.I_@**@%[15Z ^M$,VK_F%B('U-K-[%=;J&$&9&4 U_E(#B)2B52S<(
P#-8>0.Y5MGUR9IE;MF"<7[W\F@78-PP5L&"-1;BQ.;ZB2'MO)Z'#QYM ?A-D31+$
P#51 (;L9L#^]@@21C5WMF[>WF<3D&&&!&!<FL-YHET.8\4P[%@;GP#D6RJNI!@IT
P!5+7\&EG@1KN@\5$D;&&9XK\'?1G+&&]QSMBS4.Q9H4$+H25 X>1#BX9PDMTG:F'
PL6*L;]_87J-G<KR609S*+% 0]NM-5XQA3U1[18&KCKF4=A.F WUNRK!IGW=YL\Z(
PY6[2&0FIS7P]DQ*H<D&9QC:BEN#'EG,N1 1KP/")X=^_JN='J05#]2H8C^<B3W&+
PI"F9%QN;#- *K.VXH[V6[DT/GA%0C)T#O5O^+#5<]:NM= *+^\*;!,GW/\>5%V[D
P8OX-U[T9Q)[EUP>*4(*_;*"9DPXIJ[)0D#_]H,4<36(:77.YQS @WOMOY1"@P>Z=
P3%FFM4A/W0OXEV]1].$\YBY*;[5 .U38_SQD<W]S68%.5W681)^><(_2N('$0JYM
PTN:UH,EO:D3$BM*<DPK>'ALJ@E1@C2CO+/B*0T='\250)GV$Y1ZV>G+EB=;7><X_
P65N<EX.;^AP:'3M0[^,5]TB5'OII/^'AO>2T#2.Q/D>9>]"B#E5+NHM(FU-XV')&
P;"T?8>OCBCRVU9:QJ@5>5S)E.+EW]42_Y)Q34 23>$F'1UUC7XA5FM)B_MS+N^AA
P$GB&[C;YZ7-M$-'^#'E0F(MLJ9!,")4XXIOU:8-AYTT6M+D5^1PUUVCT>UA"A7WL
P41Z6B#2<3[9\L+)6$;G/:W$$K&>,XN!*@R473\5KI\PR F\VZ[6)T-4>* O^]M1]
P.T&W*B(6:=+VAUYV>HNU%@NG_@FE)J*M?RG:U?4]08:V=AMLZ[*<O?3]P;M[;]C1
P(RZNS!]Y>PD.Y8@;ZQ(EMRE0(M#6:%<1XU?B.0*O.SOG7T?N]EWM?QL#G_'%B & 
P$:N9)9X*XBK=C;AH?Q<1>D.]IBK\W6#41EFPL,"W<9MHV)YOY93;B!>[E%D)(SQU
PX98KZ6P!<&(AS0GR'K_"&AX/I\T8[V<JKDB!>%ZLEZG.(G+Q. PS4.)**AH_,CTI
P2HA4!_8K;()!AQ>TA2V6Y1#,$XL!WDZ)3&;5B/RWH8>/V@)5L^47'IP@>)AM(P_G
PR%T8"*"L^2S]F@<<!B9W_6>6WD+Q#[94+<XPJA#36F!#KIP$DA8E;.9>"Z;[]8&.
P?V)YNP_CAL*I=,GL7:"TL,X\8="3B5=2& %;8?R4!NW$S=ZW-->"G'FWA04RBMG(
PP'F<(K ;A!PY,7S9]WXMS>ARFTOM3O[5O(WK%_![Z$/&+R;%_;1X'K:<I<X<&2UT
P,FT8TUZ@+%L%B][_GKV."[+_T( J(=# U3W)()Z L6+G=X55!>USX1M*U[(W62Q<
P&?8<6<#<^>A0Q3!B??9'RXQ/=A:J^V:7>F7C?/?BK7K"S&%=F'(+P"VM/9J$2]!]
P611,\3KR1SL7CG*TMX\F1N7J#\O]HAR>"U3E@8Y\6!=>^WW7(Z8?:2#92.).^ ?P
PW",0?2?A[CRF,I"XKIFP.-53_H.%<0P)DAF1GIA3Y:+@TV#KZMJY6"DHNP_J5L<&
P,[.HT#0]^& *0D7$.Y+)+3!M7AY4GPIO*^?O-C/@_-,P25&2T!F )U?XJASW(KMR
P\X!7@DSJ2RG_W82*'?0V4#<^6OQ3\LDZ&E.,(O$?FKZ*=[Q?2@N-+12$VYCD6PF=
P(\/SKG =OQH:LG'Q&XOH?5D&N2I\-@$[Z_]I#Y=&B6V:@$Q\:.-<TG&(ID:'[*7]
P.*ZATGP1*OVJ<EI8I(GUVZQVM>T,?@^!V/BN;U&;-5<%XG,W1-'I\L< 3'K5.&UQ
PK.%O_L0E4IA"MMC':/7MYGN<I@7*GC+B\I?K:AQ9P,G(/-\[QP\Z6.>_OI,G>0?:
P?5?0+QI(OU3ZSY TX%!N?7KT^%:S8&0!6P@748XS@CE4J4(_GCYE2G8A%X =*)VX
P)&?X,!]N/,YT8=B*6&$L "C73J(:JWO?.&SLP \B\LYIH_=J<'S.4)<ZBL(Q"C,<
P:F%)#9H >()TQV?2WX\%3/6D+6 9D76+6FP_PQUD1E*=3JIK)A(_$;A4&[1%FW3>
P-$Z4%5LG#F"K=&;U7:M<*ERT=.<L@""6#]WXBG=+WHN8/"RDG+)'1FD\E+5^V= -
P MH6=#N4CJJ2OYE5/U>,V3W_CB;*;%#+;@J]73BQA\(ZY 7MQM5FTFO1!<8R5V-#
P*[XEG1YQE1%%X*<EY.AL-H-OZW[ X& 32U=IDU\)0[DAR%9GB:[*;-RQT^9P#@_(
P"-_WS2"J9*47=GGLK<(RC!Y*HWK34F'ZK+JH>(&^4/L;"H-T8(!*N;_ G#E/U]\J
P_G@#1Z4Q7: <2P6]+=[:5[+H1CL$)2HV$G>N$JM5& 9CQO6V%)&*LN\"[*M,'E3)
P8S(GVDHCDUBL(/=;]S+57AL^EJEJC8G*R0KGX%83>(W$XVKJ[*?'$?3 /=4S:X5-
P\*_7*J_I;=.4]-#DE-UB5%4^S^:-79V, $X^F[3>'=V;XU+0$^$5]OD8E1_TRJIH
PXBP4>V-ZTX<(];DESTJFN#8J=!U=G4Q:W-05!E[>@;'EC0RZ7AU+[PDU\/.>4M!;
P;W"#JTHP\^4Q%L/S9M2GW1?UF>DUL=^O),4HO_1=#ZBT*:TY*I8"9XMFEI)'=3=E
PD:"*!V:=NH_G6HS3C\];14'+3#VXERK:SFMFG56V,QX"Q.;"M?1KH40X0IMM[MH%
PW6+"8<*_&-K&+':S^-CU);ZQ8&=7@B8:W M=M3++=L--LEO1!EK*#G>MA<KP*#"$
P52IA;29?Y:^T^Y^= +((@L$A8V"+PL^QGW55+.F^=K$/3M;T#[I@4!XQQ*E[1WBU
PN\YPS0HQI2J3[@55Q@.O?X-BWN%SG$1&@@D+]+]PBZ.ZJ$FR/<V+4<"/Y+A@B4R2
PXC\^$&Z\QMU_;>XI'[C#!\F>48I,*WJ M"^XAW&*&5I1R4BX?_G.ZS 7KQ%=*PY/
P6=^M892K=S_G.CL.[(S<:T8S[)9&AP'X[CF<^C[\U=,Y0VVC4'42-:S-LU22.J6(
P3@!58D>Q,,4F0J-Q6'&-YW?ZBJJ#9V#&I9!'V1RKX-A+9HNX2&0D>>>>:6J(E>3)
P9WVG^F% X0AQA%!I;V?&  _J4UM!*NJOIA1Q&CDP5E)L4TZ[OUO/3>9S>X5>^G H
P4R+?UMB5P3?1=P/6_)(D^73OMD]4M&1$B=!_)YG3U36&\\A Q*.3'-XL'I&\1C%?
P ITV1YV5/_,-U!RRBZ7V6;A5,X+5R)T,$N*IREILF:^6_9@/2[4?'GMCS!6!8PZ,
PCM9@S7*_Y-2MA8#F^82.O#>!'V]V@W-\^ZB'-W?8/_M^?!4,[CMLH<-F+5BG5;2*
P?&:@SJ,YCI]PEGS[&O$[GD$1R:AJUB:+MR@@]5VKF-%K9?G+55_->^*F"Q7X42G7
PX8<VY&,@VN,_#QE3UT([X:UY$<J!U#)KP5_[?WN*+O.?@#@#R&$^0YQ'\9*%)L>(
P2:^+Z/UI/];WI5#O-5M!SECY?[RU=B5N*/GG?)T H#*L_3T98["N'7(NPM.Z_K.R
PM_1S(TLAGV [E?EZ;@+"TMFH'=ENTZ93DH(C5>&(F0XD8RE^SE>Y*7[.CEDF*H%=
PK0\E?7 0>(*23]-\ :'B/Y$  *=I%*4V YK=T'7&DUS-:3PAB#YACTV9'3QD6%-Y
P9.O*<]GA[P!]!?O+?5K3*P))86*Q;;LK4.KVEA(S-(%6:( :I_Q/+)W*3GZ;_D .
P8K0XK]4+[IEQBZ2\?'0)NB9V.JR#P@A?!-^?=5GE?+.9IK1E<ML#4WXZ=A^0E"'$
P;09!GG@ ;[XAZ+PGK",Q82%P77J#0>5H7,Q<V3J(=P[)%U.UZ:>Y%T!-O8-W8(YN
PQ6(K G8%S+)2></!R$P4@NK^N=GL!8'N!I7"NKI._5:9<OL ;L*]"*A'-7['MB-)
P+U*U*G=^]\CT<8]/0I+@+!3^KDRC'?<@,<8(+BCY.KJZX^2[J#L@).K:T1*TO&2O
PJ(2]:NL>UQ!#5HT3^B)B+BW:X(UYV[@,/+BY4+V9W3:-!; ":<34L\1#YO<[557D
PHN )>G#3X4/_8%$QRB4'Q,ZU!FA(,O*\1:K>$<[I@2Q;5OU$4=6L,%CX@ /:HYIW
PD[9WA*.EP&J6P3/M4?O*)*L\)$1W%+V$CA#HHJL9K VPI.CZW),FPK*G/<EB"":2
PD/Z)GS-:%Z@?/DLW,V>U*Q#R3&I^>^@3GU$R#YZ=8S3FCP?,HN%/5?,;5HL252<V
P:?)2.&U8SQ*Y?#P*(]/(=BS\>$38EXS--[*T#C_UEG]&;U\]K$UGDGE14"0UUH[R
PM$8UD"#!$Q[ZY+F5L'AV#Z4$"^OGKN@Q>M9*,W:.3;LXMI>)X6\=K!^I_E6,0U#,
PEYAJ;PPQID:SE5W Q5'I2-GD *A9T?\_RSKM+OF8 5)6S4PP4F$2ZY7.B!0_3192
PS[3"A&T#V8/GY%!][V%Q%SL)2F/8VFUF"@>FG-X%/)2C6;4O&[H9']!!B]X6#WS@
PJ/3L]3ESYSA@/1WGY=RW;MYP<:]$3.?$0,7TY_R0V\ (/[KY!K'0N9>T#&1B[#+<
P!)(NYU.,/9@U'2%[A])^[[H\38GE;@Y1'8JEG:CL'[5ID9S!3 !2H@//(R'_Y-A?
P S&<4?^>W&^HT3@\Y$(V536WBYL ;G3DFW<R$VJQ($D64%_OC>QMG6/1:7_=M$M 
PP^^<2W=PI>#4B108A/,7@*C:,942D-)NH:TB#N?[N_JOAC2/;O31F@'H+V)'58;A
PDU^\=7%U\5+,!Q7 <S9.^Y\@H:=&,*M*CUS6G-@[UM)@LE'R/X7>^L5\:(O^W[Z<
P$8J'M:ZXOD[R0U5^ **Z6.GNDZ@'F$N+X$A-_3DNS_G4P;,C'!U\'QRQ?OI5 ">>
PAX"=#CG8,?L^/9-'OI1S_^YOLQ-ZBR[)M_I.5QYC5[E/OEY-2YS;,M!SRCFD&,+[
PKEAS!;1I ,L4,I6-3))[=3M?)O<LZ>U005+%$<0AM"J@+,.4=GG%S)9=50=\@:V:
P;T<HM^8G?G?$<BF-X MP7&AFS8&Q>,N*054*[YBZ?3!(<#K"\5N]SXZ=Q[G@U?>U
PU@O0U#'N$&O+[ZX(<$#P??N$4$O%F_>BY":^=!%TVC]U!8S^,*;4&K,9!=1@9:H$
P@WS[=^V>!>MWR9Z,?"99,.A$>%.Y_%ZFQ.YDI2PI$Q;7US2>7+@"9!LK*EG,6]&R
P=P I;VPPL8"DT&'U7E%2N5#O!7T#:-B'EYNI,WF67D%9O4><%REGJ1FK(]:PPF^S
P5EZOR)LAI_:W!8H";K.H=4!8"D% FI3]TS52?Y*=KW-.!)^_!V%I>AOR"YF8D_' 
P=]8!TPYOU#+]=O76S'JZR35QX1H3L@#/,\:WQ3TG*2_ L'NF/>377][! #:S+X-9
P8'5(-T?;$K'B^0NH[QQ!CQ4G@#MJ7THL//&)'XKKJ^R\%STIYO&"TE4^T3V%;U,!
P#_O! CUJU(.%_7+CYD'$#J[-)B;"+E;,@4S=^OK@O$/;K=$X12+;!LJ:(QS*>@*3
PNT"@5Y;,MM,CRR+F,_Y'G"$Z<V"%N_\FC[QM;<#,YO6,S7@X7RCEQA/V+2;"+M?0
PS?G"?*Y1TG1C:HK2P\R_V/SV/NC#QU5B[0 3 <D^ALTB.@;\O?ZJD$:C;!A!=]Q"
PC&%3SY#AIPV4+EE@NF0L_\&UMZMS\7M*Z%GZWNK\@N"[+^0<(!@;XS.<JQX[3JOD
P'I@!<1Q7.UUQ]&)@#'LEX+ A%'!Y>R(_.>\*V<RW/:1,03U;$%@HIEYX(I*8 W5^
P)T2N1Q&_2[0\PL8@24""O+DPVF@\YHKO0<<$[^>(:'((KQ'A48#/GOBR4%,4P<3C
PV.K;<#G26#^ :$-OK!%'CJ/E6/V8X.X)!!4@=FV \=)Z^!K0./X[0'7LL.V6,'P/
P A&(&BT[61EL.#:ALJO*.7G\A9B.;8UWDT8\HO51WT!Q98ZGB%W^+/\=7<++WD++
P6KPA2_9B_?!ENV, DO/T_[ &BE?0*MT-=55+G)MEC!P=,7BQ4%];,1;#-M,O5S 9
P-E8]9%:G#P33J@6)/4KF).*7UK=G&B<?4+QPX GG50CS/5L*"VUUKD#N4B_?"4 Q
P2'E8%,K,R.T5@<UZ7T60\X:\ 5$F=O!.9C![D;X<0%@I/*(35A8P*O?R_Q\<NYV4
P[F20/$3@(P<V(PF'B-[4U!$&+GAMO%R/0+R \5 XXKCE4-F<5"3$_T))0Q4R]34 
P4=?_Z;I3H&C#*H&K;SH?Z''C$*&[$1&=<T!0/Z=#K?);86 96[I@F5-/L7/V>/Q)
P7T6FDC SU$#T)4R9]JV'</3243#2YWW/-?34[$1M9&)L)2[( <A"%EG]^@'QJ91Y
PK*GHUDO*L$OM2K.$(=K8:Q=):8ZTWOHG.^HV;*,<?<U\;_8_'8&[,1A+?+H:.7YA
PF.40<1R)N 86)UV;&>1_=TW?BCB";_"ZK@CEV]^*@&=(Q*37$ *^MB<NPU3.TA&Q
P ZXBK(CM5'K>FXD]Z[]0_H4E'\VO!\9MKLC8Q^Z@8>XP3.)5:>?HAK23\KAY\:(0
P>U+<LDYI[DLK;T6A,YN]2R2QFY*2S1%^?+20V/(T3$D*X^Y.)I^:WNA8ON\SQ]FR
P9>XYO''"YE J=%1("\2N[Y3N>7!]U"\#8"COQ'[\TW8Z.!977\JLL?5H2MU,.&![
P<+0_[("Z'58.31N$6'".%&6ZGEOMB(O><5-KR+++ZS6G==+V.851:3O)=IB-YI/0
P:+:N&ED,-&@$QRKM)-)#@&N8]##P/J3WGOH_T+O^MONUM>.!+ML2CV9<.;T>IEEW
P/+6N17F2-9D/B6T"N =M%&]WE2NY=3>K05K;ZPS)!9DQJAL*2DH6\PM W=[DS8L1
P]ES=V?*6KWB.A/0CI8T3(3,*HBD>B&)I0?UDZP="(,9^ZX6*&J\&[AU[)!FN<!#J
P6=L*&)O#I#U"*!$V)7*C@>V=,PU8VV15+Y%(6[[IGC[O=KJV2$>;\%1>G;7X_7]#
P@5? 3^U<@6A)[=16?W9\/GK+*L+<!OAIP9LSTC:F6XL;?N@1/TAPH]Z-C6SF<_WK
PREB%VT#%]XJ%DP0@YQD?>2+^V\J6]##UL9Z"T-VCOU,!IG=L6;RTZA4Y$?CR5FF;
PE1-AGY2K22_UJ1#-&3BM:JEXIX9-8:R!Q*S)!N.D$0MSE[B$(;7&XRK96,L]B;4]
P][<D)\ILVSGJ:V/6*P:BQX@7L52U</,;3+UJ.DJG^._G$'/PU,X<'44OY_0-9@N:
PKLY0&F4;NO.,6Q:$101X:X?[;](= 9Q*,$]@B!Y.<G:$.TP!P;FW^O7:=KC/MFJP
P<.]F0,"Y'K5VJ79ZX\ONIY23TFRZ&L][ 1#H_/B5^MTU(&/7X4QX&#>J>-$@<%ND
P7<R78H6TK+&$7_:VE(!]S=*%]OP8&/C!([SYB9/C3+@E_=WRE&=X)(7*^4XH_H1C
P['2XJSL W)S%7HO!3E]<F3^=T*4+WBJ%  T +R/A,&A9'33"]V8-BH"V9(AVM0H_
PJ<; E&TY]+@!P*#)#(?=V0VS>-\7_1# D;=0L5P%*^4)8.!2+U0&47.\+CE.[M#<
PXV,Y^L?/;GKD<_^DX"$<W<2*+H(I4#^YYN?*;=?VAL.QMT:FY'/T\^_N&H&R+"TN
P/G?NH!!5XO!@^Y7G+W-5X"I02H()?7LR$LA<EJ&4).5>#H*>>U@ ^9ZX1S)LMNFN
PS#_ONM#]%%8M8Q;MNEN[$:U1&Y?'Q6H($XGF.@+<";-\"KX6SU!^0\&X;>)\KRTX
PP%7$?D^-&EYK</Q%_]E N0N'\1R7-UPKFX*Y8VAJ;&!&2$?CW!_[,CED'[3FM).A
P^0F[MP49NP.2'9&A6.PUN[Z4'D+(I$'QQ%@":9A>AIQI(+9Y\[*->/K_;F^M(V)Z
P=#.Y8HUS702;SW"-,VUR'Q90'!D,.:G8)\/3B1.^DAV;&?6AP+RICKT2!RC* H:G
P]V CL$-73P,HX>S1H?WWSGTEN.OG1X;VK!X 9>59VGXR[59XO$D'3DH;^@6V'&YR
P9__25A#$'&I(^!"R9H D-ASO0&8N8S0X>Z',CV+XM9+59DJFVT3XRMF[D[[=)<CK
P@2[ODSM$,MSD:9ZL6&V2*#A/K#VYK:]!#+LN5UC*9>;WIK08H!$;: )=E%DMON>W
PV8PB/F(N!K&0-K%ZK^7(J!CT> RWU5TDC<)4)V(8!+V;( X&I6=_&LU5&[@^#8L:
P>ZO+!YWKJ>E:6F::/M;V>V]BE:(B+BJX(/6#5GA<%IL_0EA=KLLPH&V.[E]87/UM
PF"L81_2F7C\VN1($J-0O95; 8@"E"N1!.]QH@N(\\^5U[,6:KW?XI. ?R+K=+GY=
PBA'AAP\*-1+,-0]!^P,A N<$(!.48K.+23)BD&/KA#D@'JNR?_^V\PC#SU$^"N"&
PWMSG:]&<CW4"&=U^)>F# H@;JI$E,=W^"=@!KEB)-=$GLIN.P%#)X-;#GZV@>1LJ
PD$BR0BU;$JP\UFL95G&&7$):QJS1%/5IC&8M1K#-IDWO-7SHQAO (8D[1OX4^#[I
P,4@DZH8(&$6[-![7:Z'3Q3'2TG2C4UR>4JR,["B=C1A5;5MY6N[=P&A5C&PL+>O:
P!K@4 ;+0G=M3)49+G?Q.89M;])" $$7!>8J3?1CG21)3"S7+[EM4;*)M(=N D#8,
P[ZG@]03N9<PLQ_RVV$JO3&F_6_>V-/$[_7&]F\2 M,7FH$N;'F36Q.!-B#F \*.B
P!-"GC Y\,3D6L9I[-[^69@17H$;XE-AN8]6<$FB#?G([:1P-^$%EP02C.DN3$I<$
P KR\.]==-5(','*K?&%S"M4\0!))9'[&).?Q:K4LCX)JW?$.6'1ATC-76Z*I0[RZ
P+X!%5EXY++P[PJ;BSV$W,QKN::F['&%JQ-<!V 01O<7/E \H;'PIX072U:-7?1:N
P7I,?)X!CT@CK="249R?$_&M_C+D3&>K&XJ-TL&4NQZ^ZTYZR!7RVA7U F]78G+(T
P7H&GS71%6ER?CEA]:PJH2'BP652J(',!V8ARTGM29^3.<_AE!%A$ [5)-X3BY3!6
PU<U'7S<N<?;7^B*EGI*"D83UJL<1U).R\V*"#E*<DN[^C";)9(8[E7V:%P6A\;.'
P1TE"J$*Z(6-(=60%@BNO65=[ 3O3ZY<7"VZZI94HHJT7LM%K-.33:0I:T_INY<X4
P(;OC";-7UDEG4F9:[Y)<Y75?"(8+WX"GD>5>G$B=0 '?C!9[HB!+^SH?S6]2F5:W
PD)QK0FYZ=B0FWQ4E@1].ZE^'L*RQ0$BCNYA->$4.4B= \KHW5O.-LF<Y/)B#XP7W
PBZ(#FR:L)]?Q)W17.DW[6)A@?<.KF!C%WG>QA*OT133ROC;?S6*VCQ!G(H?=C,KF
P: ^MQJ=0Y6FGMO32"PC.^"B^7=<F=$HE]4QM& U5CYCT1*_LGZ4$)[C79<I9L1D4
P-P'98<8S-N#KSYK]!:X1P2]VMRH(G  W,O\V47PT/8QCVU7\XU% B$$=\5LQ;8SV
P7HAUCI?O7Q@#JG@,03O;<3KR-J/'YG0)51&2BUF[-7']@75,%-')K&R9B*@F(H3/
PX:>O9B<#%>M96OO)P#P_HQP?94G28[LI4QNF3M)Y:$)=HL,6E\O/VZU17DHYWJT 
P:U<<V.=+;,JAS*'/JEJ,W!I]M3D$;^AUXT=!M79UY$<PH_FH[$TQ=C70+@+!A1-M
PE<B7.H_JM 8^*.,/!//8$U;I8[!!6]<0>LSN=TECK0$1R-3G>32@9$;W<%V-T@\#
P@9O\PTM6[$-2C)0NL=O*AM-G5Z:2M (4S3#JED6X-%K!@B=0':_+FG*D957'8E$7
P&!@HI2_K%C0V>]C60@RF5[UC78T0J*UV9T-ZO^YJOVR0J1*-+K1CUIMH,ES*:5W(
PL+]"L85#X3'O7[%IT+5=A8B$%I9D.VMMGI4,&NX27R-8@%.10(K_SUFU'N0ESHKT
PG"U?5I9*G!7A)X:\3^^*E\W,I#=$(U_&<KM8.D&%D@^/T5<NXGGZQK5E^Q;<6,=(
PG$12"PW/Y/73K@.YM :9!G-V XW,"K71>-K':E@@30@-3>*X0^Q&>B^&O)+(4^\/
PY\]AKRJ>&ZX=DJ3>N3K%?@7Q$!%.E4!>6,*M0(O6G ")Z<%CG]WB-V!H;+F8)ZQ4
PW0!_)?9%^7!0*]\,&@7]5F0N=_Z*=,(PQ1,\QDES&3C9HOQV+.>;&:."79H7$?JZ
PV1T4.(M/7\4#S>RO#76GQ7'N@.\DZ,>LYC6#_\'YXQ:VKH<6YH?&8A+K&^1<!^<1
P40D_]&3M'&;6'QQPKZ<.Q-Z#E34JG_@IU_J/2.#$]'-(6NCGU0"*/6AZ7RKU<B1V
P^4N0?&YI&A];>1V)Z @05IZ)&"SWUT>N]>B_$6.NTZ#VQ8E-'Z9"4RE#.%AU'*VC
PVC<*!9!D6-NA[?P_I^P%S&&FE5I3=K#5=;C*,_L42H6FV4!Q"/2PDRGTK#.U92R0
P!P4B[X$_QKTW;2PV,\&H-KO:P[7-RB16#SM1A,B <Z(A.[R_TBVJC,F$Q*:?:A<+
P:/9BE"J71TT)%B&NN1L0)H$L&W(0SM;.R4&A#5/7J:O05'G%3KY0=)%E$EO6XXX\
PJ^;(DBS LI>XF'*Q9#VN#G=T E_UB\:\Z. UV@@P@G.&F^]A:$A/'F,%)F!443GD
P<2T*H74ICD<&S,&T>1G(?)?-]!FTWY-Z7-U>K(]LRN16MOB2W0"3(WR;543/L%%!
PUP$EU5?'Q4G^Y J@SH-A6<D^G7_+RD!%$(+W4P.8O4>K#BK:JH&CWA30&)KZ[QV!
P'G#O(!UX._T-!*2R1Q5D8W(028? O?Z#>JQ?LY;-YWER#E%,A#%MEG[. 0P$@C(!
PK%L>4_0#9(.;:V>Y8?2=J35UOS1BA^*1O8T@UM<>AT.7EEKH:*9SF#+ZVQIB>B.6
P(,KB4F],?@QESHO2_%HE"G(7_/UF<2>6)]3J!IU^Y&(;)\.HNO7(L?H*=QI&5D*K
PJYT$@YI\4JG9,R3@S:K=:GOR'.B\(X7?X?"QEY!V2%A]*C.MPCB0/Y2)JJ-&WMFW
P?/2#^IIP_?.- .T\RR_PN6*5LDZP"_&,<;.7TNCP<%<W2<M6$ZG>$G6/=5^=E9%7
PY!TUK/'P*6CN&T+%64O/&8^.8YGF6 Q]:O7(\[!#FF%=+1HI%'<_%#4N*H34Z'WP
P:3,L9=^4M&=?/R"T5:?1V3=NMS;X,2R=D4 _LJ6L6&S1@HXH_(BDI18S=^5=0JY_
PB2K;9-A*6BV!&IQM,/2*G5;"WQDD#;6JH19)@I_H*K2JE8 WO7H04<]M9ZIW:%*6
P_E=]M8=K__%MWH9WY0VHZ$;L4UX_JRQ@*,%E3>R;!4G5G$@-93HV-%\!WIG.NHQ@
P\E/5'*7%AD1[,U@RT$'$JA  8.H)4RE/<K*/8&&C[RO-,DSKE JL.V@CK!O2<WH)
PX9XT.",%8%IN66@:J$<?#UT)WTM&TN=P[B/"C*ZK"^BV;#3PH6'TCYK=U;("7MY_
P'H]7B^!7$>2V,<Y[Q+OD=:)K.+!I8QJLE]=G!>3Q/PVMP;;[RYO5UN<7&4"_[&&O
P%+'0A+[TJIU<*C=O9;VGQ4\V: ;$UPB:&5+@GR1S;JC)3W!&W/"\%)XV#J_RI@,H
PZ>TE67$MLA6!4VF*SX^#=J]-4FUU]J$B62<K0Z89[2!&"MX-KP@AQ\ ?>XML4WA4
P,<KI$+5$EH+F6E.\*I-83?AW.BY^?,26<GDU#((M.M(LQ6_V%>F0 QS(3;7OCC/.
P$$1XH= UB:Q16@U4K%:>B6/)AX+J_+(@SU@R=5S?1/N%*;5>ORP+!-B5XN&K/]_2
PX[)^AOFMR"[C 9^V];5DW\TQS97W04]+6C%I1G5^<7/T0>VEE[39#C+ 1)!+5K#_
P^%5:VI#_WOEF@)R;YD<<W+&Y'RY8^]O+.A5R87NO@FYLX_)P<ON%F6 I&7>X*'E"
P5$K@7C#9@)+Y)JBKP^@(FP0JT5 $8;9^F'9)A0(LY=J+/<AX#'ZJE,XUF!4[$!YZ
PJ3FO8(9&MX>, %^0:V&9\+D\94_W<K>@EC[UD[Y:"P#.1>\BW#.@,J]FT(#_O;YZ
P=O\RZK[TX?E1/?86KHM=XL[V>=AW4VYJYSGW=VFY99,W! C 8HJA E)7?!+0J*21
PE-NR PW$6JV8;;I7YWI='IMP_29*<[0C"9O&,#1:C@DB+9/''^>X_7:Y*F3#\>Q%
P>,OL=]Q!;.R0M4MA]0AMO..%K\>3-E+R=?_Z:3.=N1M",M%3%(2;]J-_Z=,,'"D5
P%-AP<!2]31A9%47?C+*I<^OR=Y(=8NRZC35?9Y:HHBI.L'$-M GGOT 6,]?/!?<,
PNFAA/^Y@>W%_W:AA$1;:J*USR&<D=<"$A,/W DR(I\[XR>(N<&', ^,8'CXI-/,)
P9MC"235%Q&<DF1B:W_Q-#M%8\FO?0@WBFBU?3EHZ!B*#CE.0?>0"B)J1N50PMI25
PR$'-RD8//:NK[N<![2JOE$Z0L<7)+NA'IG8/@8+>EEKY,BDJI!/>DD:$JLA&[[#U
P%<^$ZY(TZEUG3O(\;6@XY=38UE^5Q-JB7FNS61Y$+*%<5IUX*#^3YX0[KR$P(,[G
POT]2Y7/'PS+QK&19?@6)[]^FK\S:^"(<X+E5B;*1U<\KA_NVOSVW<L^Y?C-/"-:E
PIK?7A?6&9A^U!>FTENP-7'8;2/?P T7\&>I XD* S"J4N3'XC1S%E6? ,2"M K5J
P3UC$"=')RP!\00EE?HJV(JI$(/8D0/+<::<I:\C'"#+2IX*,[7 XM[!",<*!A]JZ
P]Q_JN[W2"OMT(*SS5VR?\/D!]S-X9"2I-LN:\HJ_<&$+-AR(B<LRX&8FP<<9AW6Z
P,2X9])IGLYE$^K3(CVBPY"P> ;U# <4A)__AO\]$4T8!>PSBQ4XGQ"=7_"UK)*Y*
PW?6:TL*PZ$HJ4IWYYJEOFAF75+(I1?;QIO6?UMD;*%=SCJY6HS7&/$/+Z.L2"G2X
PI\\-).&P;WT9]OJ'T->I]G'INT\Z:.3UB]#RH%SA'S.+O5**XN=R;\=7J9:\.4I/
P1./( G HH5:.G;GISN]\X%KNN=X#\57@3=(3WH7]FKH3%3?(LD5LC&K/$!LK0,;J
P?L!Q6L@Q11.];;O$HG=$&A("'G#T.@&X'S$ (C<I.0ITUX(@YK9PMVAS_MJHHO65
P*1=5!W/V;*A*YH;/&76<[/)=7US$@@]R&7T ;[N(J/$W:$B::GV/#1INM-_\>A'1
PND#/UD-DT*2//8DH&3FVWZM$.!A]U1W^:UWJ>=%AZOM8.1.+FLA3'"Y7$"7-W$T*
PB7;>CF=K2$J0EIHFOU/.2HN*&82HTIXG3\D1G4A8'XT&;LWXF'JCMFXQY<\#4@ B
P.-O\1VN"MIFH"XUKI4"O"L;_@T+,=W+/<TS [WXKB,OYLR<LS0JD3^:, =MD81N#
P93NKV22JI[ ,0YNN<Y5NNE19,2 *<M+HDV%;M;4>2'GG$,<A^V::;TP]7I+=[?CN
P;K<V^)TV-2Y6O>.(QTL3OCF[]:F-RL*F1;51B'C']OHT*E)L"!]1@(1,II"I&&GD
PPN3C0)V!!277G^B_>^E:X4*,#/9&3XCO' KZDAGZ-V..(.>:8@:\M51)&<,['-+Z
PYIT$%*0^S&=I*"T"^/W;(^=S([7,,X(,C3N$:_%3()-8TKSZ;?E-P'O56Z$@<@SG
P9)5XN4I6O;ILW Y (A+?'"?S^:RPNQ=$GUNAR^A4NGW](V:01[13J:.W@<B1N?RL
P7IB(']]4?A$T3X(M7TO#85//_QIK&CS,&0GDE,JX6+CT\93K*%[6U,.LB.6PCZ;9
P[H*6'8EQOP+H/@0I95CIKT.L$_/78HE2[B:6MM:^Y48P(K;7A&/VL!*II0?RR/_*
PJ=PX=BG6-M$>I+Z"GU@F(&,O=OTN6FU_$1^X,]T632.A21"Q^1QX;C#0'_T0&#;6
PBXR[CL+'<78Z\4T<BZ-YN9#64:@(Z\<9Z^:_J2H.>C>-F.AF!%4PP2 1VSDR2HN(
P*<E\?=VT\SB]$V1'M^I@BN 9*PE/@*SH=]X'AEBH MWVZ=,$^=>8+69B>:MZDC<1
PLSP#JV:W_]I43K/)(^J6/SRSUT>8(T_?1&^( +!DI;5+>_B"J4F+<'<-CR\(H.$>
P),-\R7@3"TM2=:(*D_F1;TPWGVXWB6_@&9VDI*3 X]$P7(F GVR[[Z7XDP,(R;6J
PF..#,T2P(X51>*.B2-5S"QAJGGL/8GKT%# ?Y44<,*>4M[?PNM'_(IO*M&DHA[ .
P1^9G02 >S/08!>-)!E:8\U[4[K,;D]8!OF$$^%!G:;<.[W6 7T*M>U:QQ(-$%[L8
PO[8*9GYDJ4_S3S7?4:GR3/DT&;J DE_HCA)?#BH1(735&7[8?PUHU\S2>Y_CXG)0
P?F^&CFM9<KS.DJ4C-KWCVC1<@(2)WF!=/Z>Z)W__#I+C/!Q$$T[@4J:K+.M'B^%%
P<]-6P1(":;"-]*BMRZN9\H=Y'SCAHW?F;G+905 9/U>">FE&!1B80IOZ*2^I(8J2
P24)JMT?_7D9^W59<863,)]6;JKTW3D]9:A]IC,QTKYYO;BI^;#:!=Y%FCV_@0PE 
P@OL.;8DW?_D$4SW@(P<_'GF21B@ WZ/'-\0"/;X1! ^A1E4]>B:HC#)'*D:.&C\1
P$Z#"8A1?EM1_+O!)D&M$)_;=K7B+&!]M*]5^HX=,[?MMS: POQ",@0,P:)H=23/K
P=U7"KV@EJ6O>'!^N<?IIT/?8]&I P[@[/G<0]PLGAMRMFC18_1CK4N-,WWGB>96>
PK.$&/P3ZO+;I6A"\(Y/&C3+%*?<%ES\C,D,^)HY"W8A55:2[O!JKI,=F#X>FZGHO
P8_'R9.4('Z.:A,$<(-6GZ*@YE"2(FPJH4YV?8BS@;[^"K=JZAKFH;8:-=E*=MQSS
P5G:,R5*SW]3K"@O/"L9P% \?NYV5/P?4]]9:67KP<(U6L;.MZ"=D5+,,=SY33(O-
P!T,5]] R-7 ) >W2X)6S;6 ZI)E\N?;U-2@&*A&U'(5=P)U-EH(\"H=[!.'TK%NY
PJ-V^%<K6O+E0_+ZK-GZ&SU@S%]]ORU-_1>6)78CW+M;+V>A'3#DO T+:4)'R/E&#
P9UL1*4TPY5E'5XZ^1!33J#C^%4MQ6%&C:H@<GKT*)/$I^ &A:XQ9/2=3) 3"5[VA
P6LMP<(^*:W!Z=6R2I-2['?R1L4E7Z!X77? MZ'^OOZ_\,8RP5R'56^AN2H6S+5HL
PZ+3)[1YH_S?ZMH;JMXT"#P2;[F[$Y&UF2Z2/9*@OK50H2#W5Q.P \704YXP$8$V 
P?G-PMBSAIU)\9.7$#SZMR.K.KLX>83L^.$00_S#>EKL5@Q"F=*0J(-U$6W,EY0-C
P<C,FVN([;P,XG1RX6@_-.L)C2URMX #S83%V7O??DY^*8I<TQE8/"M]T?8M -.?)
PWL%D>4I4<Y%7I::K+><\%ZH@!I&R/TLJW6&<R2-^H4]B'5+@O6@Y*I _[W_^E<#-
PQ76:M=EJS2:]= ]E'H)%T$]TR//QZ4\AV6^K%-N*! 7*-JF%:HUPXWNR[!-MO>X>
P'S\* 70+1\,W#4.#'G\Y>B7P5@D"O.6RAQ#\PN$S75P4L,5K:8Z*=$<"<!3#L!B$
P:^KLHB"271I3Z!$D&G? RZN;$!N^@7ST!OG]7LEM/K:TYIM;RR3#1(!W'JP]@:&5
PG0K.&6PI9BW2;]Q"-[]),BW2?EW#E"]<;5W<Q"1D#V;[NT)VMV6Z4!?2G< '%@;(
P[WO0[L""\DW328<F76E#\Z.F9^6GZS+A<EG?I"<& EL!$'_NR&JM7&!XC&",A24I
P%I, \_SY VS8^T&9P135M)1DD:RM^JF-Z,1#"S.TB6+PGIQNFX:B7@XVS_DWH%S\
P>":R4-CHN61W ]#1-\#:,1Z-[02)\9$U&:E-)4;[@>%C[90Y]D*K&/R0.?J\%]@[
PJA$+&1M"H,',IR N] (#Q/UY^J*+W<'1&+,R4>Q2$PO5.T8D >VE\F+GT2OV[E3L
PKV!7R=H[8]M*NK+[M?/KYPD?'$.K_&S7.+&OP1T]M;Z-4 @G-9K=>N&XZQF@UZ3M
P0R(\K(N:*< +O1?)F'_6=;7%4/]8SQ%X0UP7LY_0S)!N?G!E";AQ?JWO"#]P.8?^
PH'^UAQ.:4ANW>.7;R\:*H+,""JH[:681T/@PAHJ7WZYEB>NV8EX[N'C0,%#9>0#5
PPK+0=!1@Q"\H>9L2PFMT,)CG,#62564*]&(+#G7(DTVLXV(4WIOA3U5&%6D\*J@/
P2.1WQ0#I3:>8@$+13J$:R0VP<Y!>%;QN5&Z+54L@V.&-2#TNS)<KW1I(Y^_0&9=,
P.?%TE"-*"V;I">^'T^8?_0V<*N\,-X1:*S.N:]PTL0UX"":23; &NY9,L$HF6(_M
PFFM?H="DKS9YAS+R5Q@0M+_M59GMH3I?3;.H.X/S$8Y2BN'!N!TB/_4"]I/<57A 
PW:WG"/40 ?-RB=;?Z<D^4U!)'%0V;CV4>"C+^V"3\*Y:\.L0WIL=SIR [2F7PO=1
P(\"Z=7_64U$Y]>,_@I]6K/5+_8\OJ>G5]AEL? B-]=D*.R5D3(CAS;J=75] P;?<
P_BUS9:H>*V;(:)U31>2!*O$>EM@-+NK%"D08>%$S-UCWVLG-)K]"*Y%6OE3"?@WU
P'1I]0%0 D2YAZM;0"B4BRY:VMRK-6X55-G+]OO\ J^FY=Q%:.2V"Z;@(C:+M']%O
P<6J.MM^2N\W1D<%7)\U);KT;1EC,#N=#+25:A#AVTS4 H Z?(9_M5;8M;IX$]%?+
PW\_(*34Q3#VY<]#@EI)('['_N7"3+AG %TXP3 +-W&BJ3C7W7GG\S1!81060Y198
P< B];X#W^'Z)="\56!^EK\-W/&IY;/I06"2ZK7*[G  [43$>*%<BC&MS]!(2>>RJ
P55RP3N&@ES]S04*I600D1]"YAF=\<%NZ%[GGU- $[EH ]*\G4P=1QD'1*EL,E?(P
P^5/'0MA)LE4#EH$.?"9^M>3@]<M JDL*30(F*RL'@@20+BJTG&\3P*M.K0*N.8BB
PRVYP';X<?V8)+#LR=%PYAW-\K[P/?(ES?%0]'L1'< [-J+,H%(HI@,5[C60 I] #
P\2:RI6">1[E2*W>;Z:ZT. H7V--W>'Z/HWO0Y&5@,HE]W(A%(1%>?4C [92^(:M<
P#&/M%,6*HVVOR#AM$#9XW19UR-&$F:@#JP702!*S5&RN26$U"4?QS%Z)IOX*5V=^
P%>3%W;*BI-#!A. U#S(["#T<A3)% '?FLH;)[DPBTCGU$JBO+WDO^%\A55L,%B?^
P.WH?@E=\RN$-W-4,NBN@4CD@]N2'8C6E@;$8O$;OQ&ET; __I[A!,1WY&V*LD?#G
P>W!Q;)IZ%]YJ6?9UE *_63-#E]$%NCFH#_KE'/9%ZE#+!\BVL^%'QVF [?I?0E<[
P&#!2,VILG(;HW34+,B!+*+9P0B:[O@Q/[UP:VD$I&X6%&/2U-42Z[8F#SVN(KMHS
P-D^4Y"#=[H&-)QW49*? 6L2DB''[LQD5*GB$4.<(4Y"@$29&!A8E"(V\,Z8=W8ZI
P]@,M::<I"*GAR?<VY GH,0[%2AHB-*7FL*L@LW:^@.O6- "B2.Y?Q.;5Q[*S$OCJ
PVGG6T;VN U9H-11O^@5QO@3!29QO."AS61>(@N5SQK@.>M73?S<VS/X2*T=<7,#5
PO$%6!C0=( \C7V&LL)\_&6B\)@T_H6/Y"UMOVD)5GH4)! &0G.MJ9@R7;3:9Z)"(
P+[L +WS[:6/F>#"6N^N%[:E8,QE2;>OA#_";-T6N?*MA=K_R(/%)$]!/P+0[(>:?
PQ H.MA>+&OAO:91\LJ.;ZBYS"4$\*[!*QB7M6/B8['P[32\4CGE3\['5)R$LB&9H
P%!DK6VHX11GG.3C_ HPTF>VN1[8<J0A-^^ *=SRZ2&R-^$H-91C53=AV$0?+;%W 
P6U*[]:G99*,2_:R:GCG7-+Q/"AY<T8$U8H81$@5&V"2=Q!RK1-_H8*6L/B2KH \U
PW<@/6@@F+3C.4Z5HH>.0O'XG8(%%)YTVF$X%E\7Y>1,#EX=&H[._^2*E3$_Q!US*
P7AV3W-^'KK?E*^U6U_LX<>#5.P%M\*53V@W7H8G,C%3+5TP&K;D'Q6]>$EZX6YN!
PM O_[R9!G&%?@L\N( ?H.?Y%7.Z%4#:4''-!RX7^(5QM>3&/WB) ;O' 8"H?G[9J
PR!A$3#O=W(>Q->SN31%%NRY)QXTU88MQYV#/*,,0K/T9$'(C]Z\8A:P\GUY$%)_R
PVU966A!'J%>CC"^.2B_3C[EW_3L*5\ATDA[W<N7E3-YI1IC7N9DV)#$,$T [C KY
PV[NDHJ&:];4"-O]AD>,E</5$QW8-6CX8UBW#8IE^[\7/8+3!=L1D+B]U2N!T.?6,
P*">P[X4^.3QU%W^;PE$BGTAT.UNOJ?(+!6WE*7+O[[R)*)%3MC,U4GHRPO">G^JQ
P=M^JFB_$B9:2G*S0+0@)_YLPKU6VB?QJ>2+4X^&4B>&C[ #0;MZ%<\T:"3T6HY6$
PB,(H(6U;-BZF6'Y=C-]NX@VS<CM_DH#)4$2PE?U5ZN!>%&^GL_."(OIZB2OJD)=E
P9NT2$83.=$4&9?>GTH!6&I._K&&XN7/OW\K\U42= MT9<%VM<%0(<M'-8RVFS/>:
P39^3% ["! 4E\F 0/!5B:U-6BI",-0Q@Z3>'UY+K'O[WLIC?$=8A0^^)8NR[3_.B
PWHE$/-=%PE$&>OSH6R&6RRP6/31JX\NEKPI7,03WMFPJUX&NJP_X,[>YY,[RE$\3
PEY2*-I<;EM^E.V/4S.051F2'#X]A*+W-=XV1JC8CLDZ8+=$WQ[<7]6ZMAR]FN2A'
P/8K).EH54H*X6I1^3!_QOTW ;'%LT]W7P#HO;<.V1UEM-8#R@-JF?6"SB,$1EO6S
P"82#=* 9#DUYCS0^9GWU$\\^EU(&%;5JX <-.PH9+!%BT$EBSZ5V7%,7KKX4,#)+
P[(J/.^(1Q^M./V__#)[R*V'\]/(M<=4YNM2%)B[JX<4&F$W@)5UK3OWTQ2E@\DDO
PP_#U!R#D%BFT&UA'PG3>10^1/Y[/":'>SU.-Y100S- 3?&J" V9);0!_K">=VE2.
PV7\3LF0./51JSZWS%6V^1) =ZR*MXBQ -Q!'PGVH2@;>]>VR[_25-_&_ ==E:X@R
PFN+_2(RZB*);;B!^C@:GUG5S)ID/4HL8OP2,CIAZ6NEX3R#=I056MB/1[8/M ,P_
P^#@0_:I((-P[B(6.Y4>^H0ZTZB'$8[=?>45+!@LZF"'YG12Q@-UPH/X)Y@QN>=GQ
PD1H.]J'13^.GI0OB03;?Z%;A&"[9D4;4/0KL.C(+A%&J/CZAF.&O=*)D-!O<)O:F
PO:^QB*RP2!1M8-1CPERTI<7;QIB)4WDA[#_6I>_N#JGL*!5\KP[5L.19G>!XXF#0
P9PHQ\@>&G*;W!Z\0!52(0$4L:S$JS1 6NQY+Z7KS2GE:;]CUF]Q-HZ8JN])E'WS7
PS,R*<3)2D)Q7;Z1X(O4_L4&8V2"VT*NX!&/MA> ?,6X^"[A Q$UO(T!(B*W5"2*.
P^PJY7T3DWQ_L)1FB):(<?7;3@PD()?(YMR-3@E8X-58?Q9[CV,D/7LG3. ,2MB1U
P+@<Y91D>E^$?N2]"S\LT5RF1'<H/.*'43@<GC^D?_?;L5&+\Y1<[M7&CPP)DV$.S
P8TE,$30HH[9%KH.\B0P%RZGQWW'29I"0G@*23@313$!V^*V6Z0Q=8_NX=SFWU[XP
P2VP\OC4:><?C#.NQ16CACHFQC1 $JIO3"EZ&VTD0#09T#P196C-22S]@%1#S.T4!
P"+-KI<:L,NPG4<)R$Z&5'1<=L%M#B8G$[O<;Z=OA#$7T-I_EC04P^7##O5;?R]V[
P^#/5S9P,1%@$G^S7&N$2O4)$6M'W;.C.H.2;3.! 0S&_3_V"U)31NXDN;$?R[U[W
PF0#^@A23SV-\ U*H@2S)/7&W>#@NZV?;/?7JM<NW:RT0QJ(%-;FN@=#USTY2/*YU
P.>V=H.A;T8W4NW FU*T%.:UTR<')#'1-U%.26"1>$+6A':Z!X^P4TD5.W7V_5Q*O
PL?X$.&Y&.EPR>CD"C3FHZ4.T0W9.; NDDZ6"9XI$K- 3KSH65J%PL8\DMO1)=$,7
P6V?,-S]/:>9O9KD"1O99O[+=S3S/!Z*M 2[THDA6EL0X#K)R[8I*S,3W8U=OR1NE
PG 7<R%4'5=A);,QP"%VRR)%-+38,Y;!LI]5U=<Q\XJ+<#GYMV60?8$XQKRZ=WP9(
P<%I2S-IML'!>;&X?T4=:1DLFQR)WU.;CA]6BB:B5F1>D;>84G 4ON=?G$N_\LV&_
PG@90@.57C=XPH$'"P:C;6W,J!7WBYC,,64[CE!H5&_I;E Q*?887+;_D=,GNP,RW
P*#RQ[.V/NM;,,QD\1P#H";^.S1<9I57X!:P.[R4DR!#<+BO;N<KQ/NVL8I^9ZJP,
P*N@2,-G3-VCV2RHQK.:EH91(E%3L/OHN"!U3F6'*-F?I/H89?:0SCHZ1MUUO#5OB
P?OD6$P-BAE>_B/0+ *[WV6V!ZA^UZYK4D""P"[WC?-Q-Z.,$BD<-U/)[#P[&^L:7
PS]E=YV#]3>+;]2IKTXLE')TQ(:DG$S.2JW*=5LTF4N(L%T(1NU(RQLKP[(A$U_;;
PC%VF^HB?Y,OXH$_A);K7QY>(P3B-4,!U!70[:WDC,U!#^5LB7-C2@XW<A>CJ:?CJ
PY @<<4M[V(.8N4^E/Y#5-/"PG.9OJ5T*QN7T"QP/#7R7R0R?MQS+)'EA$#I&1NZC
P:G1Y;HK-A:&,2K#(B;#=2Q<CH#2=/>>)J&;:-[H)D\0O>4-1^[F)'PXH,5ARQ>0'
PD.F 0A&+;WH^TSYK*J/.R62L.S/TAO)UM&Q[U-[X@,;R1=>B@[*3E2IK4)G4:!P,
PA&( 3!-1L^WJ/#P;/\"Y4F:*UZ-?EAPT63#[Z8+]D%UO>C28KD%>6>)Q,D7)KGQ\
PT7T> NBK$&Y5F96/_ ,?&C"]];T(ZV-FWD3RIX;V\LQ0TWHU+@'%7 :=G;;1&80(
P_I%LK!HT73U)HGPQS#I29 &%;-J\=\3O3*Q.^'&[K5J5TVVW$;'S&X&7@L)[4QX:
PB<RXHATD4ZB4N*@"23M5"9Y5<6['Y]G&!NM+,CE9]M@< !*%MKD7\GR+9Y4ZT.F?
P+>J[&YY<,,C,?=NK6Z\LU90X(TQ#-GZ=%K^">=;1N\F;\OTP#K;F1'#8=]G\7S_'
PIW1NJ3H.+61Z+U\%-E'JJ +V?=S"=Y$8R;9,^<DPU9="I%@+J3N8$%@+$U*<R+-/
PRKU':FE+@BE[3>Y=X<74$[LYQEYRLA8O)#1Y8>VY _2V@8+OV5)A>HT3HY)\$$_U
P>F*<RSX/P3YB+O5$N2NI5B_;X7#F#BEMM2"I9,6"\<B)FH9@4[/\^ Z]GP=H$G;S
P0N!XC*3?GMD^GO0I0$%&N\(+%0WD<FW<4:_BKV!&KN*H96EL[4I!=%=SH@-C/WI.
P< MY'1FR6YR!FK%E8F+B\9F9>SSG+. U*9W/. ;'@LSCA"]/7#\+0)3AITNG,@U<
P7[0%;F5/EWOF6F?>NPH8X&-/4ZWPTW0![58:M\((6+4Y6DA:4(S@AK@\QUZ</\%[
P_H<S7.R]=,@CL%^ RCSW:\*M2C@-#:JPV^1H'_T">Z!'&3$@!AJYJCGI8FA>?RQ,
P=#V5K<[5EJ^B7I:IY!'5W9:HGCM.E.-$46.=U/#6EDW#=VA)Q+8949:F09B$7>GW
P@2T935 <*[JB<&+']F$UL]_5%4@/Z-&_JI]&!H+0/.0R&'7Y"QXE"_^ /C*2[DJ<
P-91:W"<YU2=(064>CFT[LG$#.2P^* R+=]B&<D5W"[=:O<3J.T^%)[/Q,C,^(43<
P;7RO;+0C2Z_#87AA8^1Z,:/ =O09 *7.PL)<EO)VB,P+S&F\_XKBM(J4BC9>R$'F
P&=/YKC *:.T##05+<]4D @U.;>=OL>+?T(F(DM2;%)08<1*'E8(.8]>9V^)R:ZS"
PG?9E2Y@]GU:M\+V<#?V2"84=UF#^DJE_?A]1 T[$?LAF(KT-^^RR2>%:?V@@!,+ 
PWN),*OCC,KX]X+#24=6,8L@!%M&H&JJYHTS19JIPH9T"7@G=&I_=*,;OPOW95N^I
P:M 8TM1;1! HEMK7DT:$.$HXQW2G,TX5]EN9X5W'\L5#?DBDYJ1<;C7OXY#U:T$1
P>(VM^F=,AI 3Q_4?0.,40=O0T(> / /.*>"YKM1>-L^_WIF;WK+#-Q6XG[4YCV5#
P+4)OE7T^B8)#7-S^.Y\ _I9?MK7"AF LG.LR/:.*KJ_3S,H9&_=CW 7+ B0@D,9I
PMA.OS-^.:.^S-M!R<W/X-C"8EP+T@[X9(RS^_5SQY8H>DX*_?+X@=3!A>%O%>C&P
PY/N6A1\=_:K2E:Q'R;M";3AZ"#*MB09P!6N(S$A-\,AC"5T&N1E<&'_INI .H)6V
P$U&F"A <R$T[#AQF$P1V-10U^GX<3-@N!^[XU1N5>4"]S\OC <U'/R\U#@ZR)BIL
P9VJLUX5:OL)U=TN8+,)J%GW34L:OM_/UV@OL7IW9<K)H0 ]&XR=,0CL95\0.[!.O
PWQ+A@QPK]Y4&\'E& C@VTS0E5Q&X]SR#A2B;K&,BF,3^VACA)I4&UU7AT_/H]F1\
P<4WXI$? 7%B/0>3SWX!N$+E$EB^1XD$7^D)VZ0*B9%A"V]3,G<I25OT&NBL$K&#M
PKZ@R8PSP^9L(.4*6%70:8UT'.>&"@W@2F=]9=GMO?KAA0^<//-/7L=8,.<MJZA $
PW+Q261%A;H*)\5.0+340W=D/C7$.>_ )=;'.T48R>4D\WGHWMF 777+*2F!]]78]
PEM-5%R^5$;.1!FX!N.H0M48V:%$?@[1. N&*R*^#/#7Y-#_=$T^89! M5%[Y\B/O
P_[LI7?@:>\I^C%@6Y?Y8B0=&HT]9>7%.5J[Y*YC;*[IVMZR5F:6YO;R:%[/Q+/(A
PG'!ZR^V<.8*#B#\E,D$46YJ[)<?;B #)6$=\6'>B<#[S (&6 :1ZE<41?6$SE MV
PS//I0#L;B)H-1;:GKT;;0TW[*23N=;:WKF,$U2N=%QT3(A6(,3W#ND^IHMT8O$XK
PB-.8#3::C LN/$EGMQ_,DF";W2X +)OCN!;54_Z^RVM+YJ87")VK\ZJ<S-9G=0O*
PUE#D#P%!*TXA9QQ"RV5)+S-]A@$T]>Q9B@IGH'RR;%UW?+A27+?5T&[P0#&'ZQL)
PH-J+.!.)?L\ QLV@?CSOW<-T*/L)"JQM+^39[_;=&]J&SM>Y]2X;0 5%7D,&M]P'
P/>K191$;#YKUVF=^/QOV:6)K4D$ B\2>YRW=_-[HS"I+$=#[3KM.:=<C;/*.$7.=
PT-U_I(T,80:TT%^O+:3D$IR=0 'L2PR+]DNL'1&.6NQJ2'RZ3'4/24S0TAN$O3F2
PZJ-J7V(Y&OHN[ZO#4>N6N).O6)P^OW%I$E 5E$[Q;:=,6"HLD(FMN>\=':I@E62Y
PD8A7S.C%*Q2A.'H("#E\H65VQK;$STP+SX[\X9:91 V(>IDZ4Z59EM^-F7K7.0)^
PY3-;_"."V/5R!_]\[?)TUU)1#N++,'S15@Z)Y&]XE;UAQ E#=5H*>,U\Z'0_7S4N
P1*12@.[AZND#*,89EF\6?+GI<>!C+#IFU^:82.@GX$Y4B^%JJ17^+F6($?Y!RT@[
P66J*G: _1<:CC\'*6G"=XXEK$\9QL%1QO;1H\>.YD^LKY'W&[NU,NQB <"'&QMT;
PE@[3RGIOEL;N%OBI.:$2>.4G*BVE<3=*^'KTX565.\U"J>8<*P./P4R%H_YO/"2Q
PI#PSE;;Q;@0[BEI(O>J7]YB[9;@27HLZ;XG>EOG=D[;AW&NI.12J_R.GN7QAZS)G
PQ3B*FVR2JXN#GCG8@C4T W WZ7HJJ#7/=J)HGI0]])+J800RHUI(Z^<A"6YV@8SO
P-1.;2@.ZU/+\X-S<>8O]!?:2M]J_?6ZA-9DUZ52HQ"N>_5\*B;$0W['/%DOIRD"D
P2'A_ 57[$::[B!P@1YE)<XRR0,25.%\07B^+%T96:.]P2'0W49C\5S<DBN(X%"PZ
PH4G&#M\T?>7GL%S'WVUOWWABU2PS+=-ELFT$PGE]"6#5N;2#RT;B^6>BZA?/ZL9=
PPMZ2&>+W=\MVP"06BN)SPZA:E#KS-TZO4H%P40]R.-/DI+4QHC]#_R]B,!7.':M:
P_T?:V8WC#JRT27K_HX89 V#HK!6@>CH1TRHL69A3&T*'W5!8%5>*R>TF=U8:VU>Y
P0Q ]=DG';3.#W@OWDH5,HHZ[M.>[/9?Y'8'!UY^VYU.>NA9QWS$"%?HJ/ _EIZ(.
PH9F%',Y8D?A87%1+)MT3Q*+/[;_B*A-OJ+F[2YD&O)4=Z5ET"+)1PIZ_4N=*X5,G
PQ_F?I=(.['ZWNW?;8(8->D>4.K2"GA$'::Z1I1:TD!/J$"!<J?]UY^7^:*TR1KF9
P5UDBH[ ND<75DG)#_[UJ;'8P0[ZQ)9']RT3V@%W0/-E]BBP$+:+-OUI%F3>5#EBQ
PZ_*W):FUJ_(*TKAHW";XL$$R9-<Z>DSG08_[/<B7H;:W09=)[4!N5J!@Y7M5^ZC)
P 9=X7B.*4U9;%R/YK*;RDF.]..KAVQK]'-:S#B2U\.IP[*^>]Z@W;9 9C#I>P\LT
P^UW[$4O\D!=,HDDM2C913]D[S0J$.AB#;]"M!J6E<H2*XI8;/EXH"1"]EY_LN#4'
P-93Y,I%9$G-9E #]4V *4:?./CUA&T9CF8AR*03*\]9[P YE9\1V%*K1Q88(2O#!
P$=4\EXO8%:"W :9\+G_\U25D44751+RET4>4@K,R]ASA%>+FHXP<%'?4A["C#*S_
PN4@:(AO_4I'3V,U.-MM -41R,,+%I?R[%?C)1;YZISFM VB38E2F?JNI'4,)[6B<
P<[W LL*5?9D05Q)<1 ;HC_GFZV0YGO76CKAL[>1&&C7SY2KLQ0<L)VD,J\YC(HS"
PNX,MQ&$YB&B_9B<$5(;HAS^@?K:J(],CV:3L6PA9D')L3D920&ZCO.'""'3[N_6;
P)YXQ33(_O\2S.W[1U'EIP"ZO+& L?^[>SUKUQ?RUAB"(,*4^@8S(]DH+ZZ<BR+:G
P^/3K,!;GO PC?ZEI0O]Z;C@X1"VMF&N-:?R!ZMGS$4/*6E!4JOP?NR(; 8ZU(%;P
P9:CX5)%B2VVJE(>(3YP;>UPW1-YDU8\8E-2G%9.+C!OU\%7Z1P<2*E,4"=L='#(W
P753)01KM+ZTR1;/5U+PQINQ+C.I0\.XJUZ41M]R6]K'&,8,Y<H_'4M 7HUQQCW 4
P()0V.GD'D/:5%Q9(#I9ZU%W(KZ4PVE]BE>?IB@0I;6[J22WJ)+,_6J0T8\]3TF^,
P(DCK\X/:"$9&EFVI[$?&I8RY#Y%'FP=%RIWV\VQS D6-4@Y$V!4>16CO"TC.YYAG
P=>:<ZI! V^$;2[@+0?G%QRH >N#_G H?.KN7S@?#.T7K$A*%D(L'HIRI0,?S^&OQ
P;CAWJ[C&]76)_.08 BK6Q8#7I28&,.^T\I/DOR,.1^>($[F 4*3B;$X(G..BE9_7
P5B$9+P=BRK+8 QP5N?OT"_4=28@YZIN$(>D'/6:R%#5%&V^B VRQQ-^^14!^+!"K
PX],7E],GT/F<Z6R]_O)@ $3#=>&5VKBA!H'QP'?%T,_CX;L"43 \SQ C'+G]W+/-
P(,J PD6B3E-6] ':<[0O1<<E^/ LGUF(-KPD4)F?Z]*I269M[TS]01?M#,F)N];D
PCL:J"4P=AYG<4M)TV]XZGI=GO.*A9U^S",E+>28$'[+-R>&HETZW#B;B6:\!O:/H
P:_036IM!J]L5X/")#<B3^$0X&U=IB-?'Q>6E=?5H,C-<1_R]V(-4IIA?WJ5@4N$_
PK> "$R"-,F>Y%;+:.8@D"W:YM2BEFX,>=EA0?W4+.Y<XY_&(7+:45Q2O_-"+MQPK
P-0_=RQ*]BZS:4 ];AMJX+3>YF8W"F.^#:P'=0&_AFG)$XQZYV \7 MK>:;N2\ 4W
P6;369BZEHCDT,A-/V+N4XH I]\U:>$>ADF],O05.#3F^I]N!1TL:-;3I(C4FPQA3
PYHD/;%Z2XH?>,*,>Q2C.$^HCB^RH$UJ'HEZ8KVVZ)\MJDA &K:H$3IHBH*#D>[.2
P#8/ ^DZS_@]%J 2:)QY=;GN'5&Z<;SW6(-+?0)X;XI-?C1\B@G2S '80/CW +)QJ
PPVUY ;-;"+&*:%TG_,^A]2DW71?OAVL%"H?Z7 +K.EGZ"0E=]\['L#7A0]$[RKGO
PT[9T+,U '0 :XBZP/-B+KM$ &=X)1;/1I-1H(M]12II?]C.52PH D?2A%ZDY0<\7
P&W @I(!8YD=OZAF!K!O,9GGFT&FYC@F<$:85-'L)Z1*,@@[1KBG6$B>"T\L:$23V
PO:(SG7O1<RE5TSI,=B#2G;C?$,E-/U4'V1N K3UB3U"'Q-JM"3D @J/;9=T].XNE
P%3L^* \M7]"4>=OSH\F(4#AC?6L[T2*+]$[T9+ ]6TH[R-KAO!70>K^7@-<& U=>
P.I;AQ"EKN98-:?OQ@44F%&=JO+SDT#Q$^)>@:V#5]^A8M=>@XFM:KVK+Y#[S&.ZE
P8$>$5X2J).<WIS0L3F0J4R/*_\] =BOYAK^OT Z(U<3_"[4Q4Y,BZ-U=LCC_4GO^
PY$$#(FVSNT2L*V V80]-,&REM_2"<]K89FY<>[G:A VH"UF+^;R3^$O@V*AK&/@V
PHK9P+M<RO5_:^0@=*U._X%+E9.LMA:1Z$(\HFF$5H2503U /!/(1Y/H6\*45<[T*
PDJR4[KB3"/'QRYTDD@0E: F<ZCWG=[L8&*,7;&,*.(A DWF*]AZ+*8X0/\'8>!G 
PWC&HG,B,N.>$D;#5B@6L'9ODK4UGJ2=4%)QF\(5!XC Q?2)2OZVJ2_!DL']WK'X+
P-)C6]N?B.-CV:*5+$J)%.2D40HF[."![H[4?=.2'!!U8NRXG9UC^-A?[P2?B;+$U
P,Z$B3%QC]V:)-58ZY>3E+"BI*@ ,'\(D]H#&>'D)U!.97'UKZ !S68^IWSULKT/,
P]HD0.RFW!,BO&&.\ 4".^:SFOCY9MCV?D0')>)FP4,1_UZ=^T;7JW%&3TE[D1<$9
P8J7?&A<\7 #[3@>U!_?9W0WLJWT&3&TTDQCGVV+[^7$G*WUR"V$N"+O8#CV#S!;>
P;.A/ZC!C_<D?Q2@*EW9/'%2I1?UH8_YS,K?;DF8Y0Y%\P^P=5AP/*5?"B+B4[R^Q
P_IS;$R^S"-((^R)Y$/;T:7?^_^?F5'>N&$YCT4DOL:[6S[TK\5#-R],D$@LZ;MBG
P'@ZU"3P]DMZCG/1S;GH5[!8-J[A:C'P\3 4+5G>$H[(03/DPH_#.()\:!TI=*!7C
P10PY\/KTBI^>SGW="4S/,Q0(=4$VE^?[:WWS^A%W[EP&;?^KO]@U=OS0A)0/\<;:
P$,!,R[H3,^Z/[5\A/A98]U(S/+3DU>[VAE;:)C8HQ8F4W;Z4NA'/3M^"2M!W6(H9
PE^16?AV3D]+E _-48NND8:6@Y$LBR/K.=>#Y3/RTVO2LP:$PRYW@<>Y;BM@J!FO"
P)X/2I.<G)+"RX)VP)3(-?+2.]6W1C8[;/C[O? I<:K/ V(<:XGC5XBG8ZX,- ]RT
PWPV<0&MY#E[4':-J,9-J3YN6L3N?@^(T2O=B5:D:+]@KIDT?;S G$WXF]!V $PH4
PG2N,>=4!TIV%11@$7#/A0FD.Z&4HZJ<^#VDG]'T9S#:S*@Z&[/*[W0(44[G)@(MF
P$2ZX(ZR@7-%RP353:G-;/U8)UHL^48 [$\M,,=2,QIOBW6443I,6)GT3IDH1&@<H
P_J0^,5?O7WNKF)IE/(1"196^T1"UD)GK><;\(3UX8"CCN[SM<USBK6!MF;>Z#37C
P<!% H4-]-9E5R6A^IPY'K@;W''[N6O=0.[;[(>]1)>\XIH 3D/1A*\?T_6?%1OSH
PLLX?R3PY&TE)Y]&X].X&'(&>_;XMF.1<=)V_DS^A#$FESA1]]A/V5BEU1?Q?IC3K
PTN&UG-Z;]T6,":(]L.]7-W7(T31U8UT!B,<"78PY-QV?2MUOA!45-+BI5*O8X'?0
P_B#Y@<>#B25Q>N:8DVVEM")<U&B08/Z"(9KT]URFW#EG'I\^[>*.H7NKX8L+$%L:
PIJZ5HIBR[,XT4SF&XFU)/]@Z!<+984$@$F!6Z)Z\4G:37))M*WZNE,==4^Z:R%NW
P-X4OBR!61LYUK<!!6Z05B1]&+8D.(;S.(:?V46S[3O+QCBA.=84CE6I^_":E<-2=
P':$[EO"G>B$X1AWJ'H,02AZDS72!-1@A!!V8:^7?^W5>9PU2:@LYB'@,7L23E5M,
P9^W,KN;!O/^--Y0,H.89KLW,3$Z07V\7<I]I;6) EW)GMK5IP2YI\%NG)27W+B'_
PG:W'-S2 ")Z:/9V?^9*KFHV4SDE5 4T/AVEJC#IZXV<U([2 U>]2*H8;PL29#*\!
PB7*DH&-(.K;'K!-ZG1'O&-81]V!!%WE],*.*!]9=5^/MWRP&,)C>>.DZQ1I]6" 4
PVNEP9Z0D4FC@/;8J7@O<@MFEE>J,68N"^WH>J?0R7^31CN 6U]&_IRD9BAKDN/Y=
P%]'<"A]':S*0Z@-EBP[L#)@37#D:!OXE DF7N)&<<84-NU.QB$E&=RHN%A_('^$,
P\5TD6O[TJN':8]-\I+_+[)L6V ?AZ^ 2$8)F^%FWZZ(Y5TB'8R*6ATVI>/,M3K'I
P;N;<JG#E-S7JK>"F_U%8 -G$15-A^U%^S16"XB?5-I 9/4"-]<$C2Q]O<X&7= L%
P@F.ZJ.X.U'?[D9GLBFK"_@?\]TA6:'BW.)(:5KD_TKL]Y+;=/F8 BLZ#)#*J\YG$
P4GX1-$0""O=Y@, ?MP NOI95!*7&7'SR QC XSN9,OT3[)VT2G-(SJ!=/$TV_.O/
P KG!ARQJG(=M?K::$L?8T*G5.-4=6VDOKJI +ZQZI7W]FJRF[]#!J].TLJF;9GM-
P5O]!)%F:&;5&OP>..%ZFS:6P##%3Q3<6#<DQ.*Y]G_M^64_(TNC^4P3Q;_WV,6NR
PTO&V\G%5QVC _\;.3"W?SV,^2GFN9]8Y=AQ?2=@H2%H=' (C%[Z1I?T5\\F\Z)0Y
P"!Q^:.[TI7H54M7FF\%&I0^T.PIKPN71KU>4F(>EY>@6="U\%1^,R:QZXBL4X_7T
P4XT=&Q )L7@E.F12,12M?#^@6 H(59+ZK[DP]$=DU-3X5K< \/PLU$I)"1]/\=1M
PVWA?0%3VJ<72J]X;3:)@;F ZSAK6&-I;DRM^=B:>7]3VQHO\KX I3O,]8D5=M%DF
PICKWJAK"M)&AYAY]Y>-S@]47PGA\7-+NW#]H-=I5@GD2&8I*Q#S]&W3C+A7SJ($+
P0F, TV7TXWY=)\?VF3;*,@(EP#;)2ZQ5$5]G<!:R!K:UYX!KV>C*/:8)]:^?-TP-
P*(+1G;268*$S]"-]!>8;6H0GS9RL#0)1&6^1ZX'EJBLDUE]'JZH$$24:.G!6$09_
PI#]K4C.4XK)Y)A'I$9D*GO-A.X<@8C5(-'E%[XQE?&<45[[=I;2LYJ$<.4'LMB7V
PU4E]H*VZ3;Y?Q&>E$3V^$--LL<X]HXV8EL];*X(3<T)OOIF%"2>9QUP'DP5.!;V!
P*KI:&-GUP#2^"UZUH49X97F=LC^/J0^ALT<WI;Z8P#Q.T%*#MVJ.,USR-?\8V42"
P?F-@$E<_C^.!6KW0A R0"F1G(C+M3OO >S,U)=&'6@>#X$NIT&%=Y.O2D>-T)W 6
P/JQ%2%1_IYZ,NS??!(!Z<-;0)06BM5M1XOHU)"@.5*2.SE.XKMW$3T<%1&RF"#U,
P6:7LPI"=F!-;VF.74XT!+RI]'@+$=I@#SUS[9J64))?XH>W'H14;/:7#M@\K(]E,
P+H)V/GA7<E76Q)F2MI/"(+.>X:EF7HH(R?M(N4\\C2-%\^O^PEBB\D-U)>$((C]C
PMC,SV/(USA[WM#H!>^F$< [\ &&."Z2V[];[^#ATQ9'',:-N<H$O,OMU/>2M9OV:
PD4"UE7=9_2!N3M\,KO3#JA3D1LX#\V?VV1=^41!B(4QZ=L8T)8-,]P/A\"B\W@1M
PFW#,1?+I!4?5^2\1S*.[]B@WB'+\4__Q-XO<5:.7IG(EV$I@ E%SOQU,S_,S.VOQ
PHJL*!SN1^A2E<.94DKC8#J]#W*?:7/ZSOU ^R$.'-,8M0Q1B4?QIKO",A WEO8*^
P,E:C>1F5;1 7M? )^&-?N(;?410K!\H&W_%5VD%5ZM#Q4F7F"#'PAE[X6!UJ0:>(
P^ Z+8__J*C+SONF"[].W:E6-@+<WCY);;4H.BE+./,VS'.&QCS:DZ);*N-,T"4 0
P4;5+YDK#-;A -[>?F(";):?FMXBA%1FO3Y^U]EZ0>0ELC8^_<WI'ROCAAK_#RJK1
P"AL!:WS6U%V?\4[\8K=^.-21[;"T;F18QYO:D\EGN54J&F?1W)56W6D;>#12*II(
P_8.:5^!][&^TU=S)T+KQIJDN8*,=:=^DFQIF+%JSV"'J)@J._H)H9E)!AS$;A>[2
P-U&#+&_3_[$.U3T#]*C(O"-B% ]'?_,+;$"4N'D1(+,XT%)NZ,#:M=7U9*N:_WF+
P$IJ>.21JK6]_ B@,1(GG\7UA\!F5C\)V3=65.%_K7^/9D\#4+A9"F9@Q<CDP7T%,
P@6U"/,U:O'M^)(KDMWJWX=R:E""\NC!=S*,W6G^(MRRZSW;<#V&YIC(\L[+B"@=9
P[-!N(  7OK73[=1<8CFI0#Z$VX7PP2]5Y -XA$)2L[8Q8,KF\C$V?K@Q(#%4LWT:
P^FFP!@C8"PIE(5!Y?X+  /!:[)---190();N*6+CB !]9$2F^#Q*$DLGLDF0=V"L
P8[%0E=+>!AG;;Y'9@I!:GRPJI0L0610/.?AG^?\ >$.@LV:^P>5LUR'PBD<A2;/ 
P[60?WLEKS7V)D 76[P&D(]4IJ3CB!$S([>0<N+2R<^MAA[D\@$!!C">759 WT* '
PL3M0?U-F6M&_/XPZOU9@*[-N3@]VJT>X#MG-%LA#1AB53C5V)[XF8?NG?<KLGFD%
PT,GZP0'%I6O]0@A2I\G_UUWT<^D/TG]M>B )$<'W)\\Q"W_WIP+0_LKZ;_U+3O;)
PMR]V9#2PG7>S/^L,\,ZDQ!;_/Y[,LF/.!4P,D,7O>!XF1=0,(^9>V62YP.<6<FQU
P26P-=9']TL'4TD"Q,X"-I>XO']>);6!]+NY86T:19SM%N;#8EQW!N4'^;R:;P)_:
PV2[N5*LOW)&;-2WMD/ON;6GR"QTABY)%?X?Q:?EI4CESY%B1E<"QP&O\P^#K$[J%
P\!T0XNI7"?/G[#=-% 0%O,I>1\P*9&M8&<TVJ5TBD%E #OLI;C'2BID447]MN"]\
P>/6K/6'6/]P\K;"18"JEZ6<YF8NIV2WHM]SGULZ#.)BQ>=P.P:.>VC73-\KJ[E (
P%E5/S :94A%I.OLE1(^NI>*Y HDA"P>>*8>&NX*/\'*0;LA5;*GTU7U6V<$)3%<O
P1^YON,]:G7V;T4(B+?0C)=F:/ +1R!!ULP-KSAJ4@8V>>QO[QI7/F?2?'HO7WU5A
PX ]C^O='R+PI3];UEP#&+! G\JE[2X<3AU<;%3,!9F_--N_ EJC<QHY\6/S_EQN-
PDSQCC+QKH^DEZ@9 F:<C)U[)?LQ@SW72D ?+D] LN@O[#P!# <NM%USVA'12FG3"
P_,)M)Y-;!C(]NFL$N-,MC&%3B.'P@ ,-\+3!G,O)23/3A.T.S=B%@&I9=>%PL0B(
P5$3/(>3NX[XGS3'.Z*&$R.,T8(\IW!F16LJ@FCI-61>/8?2Y$"_(?@7L#E-%\4SM
P%'9MB)OSCY,,L0I=>5F-V(@8, =+6Q2,<W@*?UY.=-(:W#CW'+^/.ZEK%]>@%LWC
PMT?EQVC"V_/51WV"V'R+EU3>4!X27*2\>IAZV=(.C;D^YC.-'Q"VI9.OBBOW^$):
PPK/P^BCR%A4-[W<--M46 ?/3&&,-EXE:U!C]:N6<*CE-,8$$4%>.AT+ZTOS*H@UF
P"$#+-[3F?5'00\L/DFD+B5N@C;7BY=+K^E<JEP8U3!]Z@#"K<RWOUN&@I!"@01)5
P'*$*1F0$6I3XMJU>#+D)*1!Y.G,)IF)KPN(^=U?XYM5\2I:0*.LT58W:<;2KX%Z;
P;JDZN^$)P;U; ]I:3D(U@)Q//*#BXTL1'<R5&N--PG8NT@42?N*_PLR6%J@%!<F?
P!MX2W?3CU]%3]C2#Q8%T<F1 DSW\ )9$9,8K <>^VUAC3%W'=\&)B1X_Z=*W_L!<
PTM(0:45V887_[EFS'L,RC[[UC:_KL#[- 6'?59!:8R "L?=YX55W4+,X/ZLE#_-G
P,W/6<>WU]?^N>B5IB*DU]NNO80G^?!?O;/H:,$*LX6O7*$S%K/7["'>SKI0W^TQX
P)8ON"EARNPP,\M=!#BRGD<ZU<YZ!0Q*RGI9..0T"KK9>T;B=L;>Y&C9ND6W$#;5Z
P[++>@<;BHI'(3<-'4X:8%_<_0#3]?EVW6>\2^-ZS7L<;%!,=3L"PR/PWYBBGQ+#6
PJM0(C"!CP%3/7_=.*Z>ZU<%KUVGV(6B]P70@5%Q&9AR\5O!XW%.-0&[HKI5$H884
PT+9;J9S!N;6$-R$Y[<O!ENYN-69W^:CH6#S]DT1A4-5]Z(R!4'$$+@ZXP7RE>X4!
PK5J\\XB^E/"9@[:VQO\@PD[N HR7N*V*FS<9P/=?X8R!F1V*?/C4\,@/X8(/VYEC
P*3<]^^KKDJHM'@2H':04)_S9&]SFM1-&=I@VSX\+Z)$]0*(0OPW?&UM*B5F>C.(D
P/;3)AIG6@=DAE.CDZ^0,J3?ZY[V+LL]C9D351IU#H&,<@1@Z5J3-/C'@M7& 1@_=
P"64D=BT4N!:4^$6PUE/PDJ(2@NQDJQ64*X_*M_/4]R?-OD,_\Y=4J3IP6YQ1/%_(
P\_.#O.K:%-;[(!IF(KYJ)/V7!H6\D+'YJ>Z8LM^@(3#1DOV5JF"XDE['1_@.MFC1
PT[J(U% 1E^KP2LU4VK.!ZY.QMKZ".PQHD$18 ,WU6-PV*J#GYH&V*[<A69C0R%_Y
P?^<-+AHBWV]8O*M2;V)BQ+BX0=E)RW/)JK/0 J]5=]1PL26',&EQ(BF]7(.4D2RK
P\])FN0D YX&HV8V.Y_<#\BSR[@4)U4+.9 *,!%!90D<$-A+8 ODYSE(GVR?+S$OS
POMJSGY>2]&L&49>[Q8'KV.<(6/Q/JRG&DX)*Y96 ?6>70H;FHV-_? ,V]=VHV!V^
PY0+:4H@]U%QZBJUXH_[UUY7:/1$C?!AO=HV;08,A<+&SE.U'Q3&;;R=)N197:/5;
P0&<Q_0DT"(."KZS;^%,>PJWVGI<L/ O"3FA=VGZ#Q.#].)3"J*9WH^4I6YMID\)#
PI(UNJ&8:69G,U-=GWN070T0;2:;V*1'!+E2JRAYEF%R88E &[,R#>%=T."Y#Z?7V
P&]KT5/+<]DS8*,%XA.LEP[C# X*WAMW)*ZPB):6,T6P297/[>?02P2$NF<Q@9$R:
PYJ>SVST7W:<TJ_DQ_^T*R,A/)NV '0"!0^70&2^B%UB<GS8P&?'B7>:G7>W@6)KK
PV,'S=(JOM<\(^(3/+=RS=;(#8"/,"IV[XI_+:/[ZPRZMPX* O\;<Z'_(.=7*ZSR3
POG7K".W&ZMZOTG?YB];,%#UOP08"PC"[^*I%G%4NKH>'$U2P0$2K;TXG5>P60\8>
PJSTWBPXRGD>\?/].E%9TJTV$1!6Y>"M(P*>#2OFBJF-APF=.+7VW+16FQG.06,;M
PR[CU@SGJF*GA#GIS?>OFZ&UE-EZ1TB2OGRI6KT,.]UL/ZRLLY&L[G>WE4;C<X!I+
P>TYL<:;QX%E!#:2KM)CA@@LXN7_RI!?Q9KN7N)6)%(%VCY50\.:L6N<;*<,Y<"4?
PD,N.!$2=H7,!<XJ[3) X=BL.,QJ9C#>OL1R+8=_V.5B.Y^7"(Y9;[M< -"\5V&>#
P'5=V:@7PHP<3+4" :D-37I 12T.Y9RV-N>HX0.YZ\#E;\M7GGP81UEKB^0[;JGZ=
PQBQ19FKD9E47O&T):^KUB[5/!I;E%6#H"".SQ>4Y8MXKI;^F7-1(XXB+5$O3XGZ7
PX1["G\]Q7B-QQVR'XC[CN]62]R?%F /IC91IFK2D/1K73\6L=R>=Q">S\-3'YJ\[
PVR[@%@I5U^S[4B:.LJO03^WE:0HJD$'EYH@\%WGH6!\M]WRE@$E2L\LJZI5<\49<
PFJ'<5<7B6()\3DN3HC".<9O??.[+9^[P(>KCG]OK H?UD?0%QXY1GZ6X9VDC_%(S
P'71VP5:Q"=&Q$F%S-$\=MDEKCL6&A4:R[9UMN"OW</1C]@QW;:R+LD(]*/R8Y9EF
PWUKA&O9*3F4*#D*_/#T/*WJIG8)P0]5C)$.;P +U7'4Q;Y"/U>PO__U+ V1XSY8]
PXLX4&*5;>D' ';-(\\'#>[[MC98 &?)=<CFD<PC9T00*&V*#BLCD5?V^. !'O(0W
P WK3&K.[P<?A?1J8O7;^^]?I71^\=7^7/9I5"U,[W"H-L:!>9+0<U &NR%R]3:#%
PZ#(@9#9S\SX$7:\7MAH*1QT:2GK.4ZP&T-J*PY*W<+W<L;+!-^$1L>*'3VNO(>I0
PR!.C#AA !#.B,O*PAUHB- E*_6)QT_@CN.HF_3DP"6$(J_</.9D"L#+ []?A!":M
PM*#G>;ND!%K4Z-XCD@TONYGR<:<9^0V52_KO=HLA5&UAYM\8R@4>MS$@',:)6GF]
PL.F(,-P !>ET*&7Y!01+"@,X\T]*6>M5X!RZ+:G*,^/7V<%F39E716_J$)YW'/EK
PC:9P72HN@G]H*TO";66/KC:\DP+RR5AFX'PLM-?<&^NVMQ-<G]#0$I*ZX7,/*HEF
PI\Y!@?EOHL!6-;=_E#26@^[4\A4C]5VNG[YGCA=%@LJ3PC3YZ),Z(VHP/44A164H
P6GC%5)M/-6KR?VP(>7MF59MG' <^7<L!MRRD<"6[N%XG&=X'B0U*:D+27?,V'6S&
P9-(:U *L*GP%46H+;\:1L&7MG\V;EH8N_LO$>N0P8..H_:/!>@C,[KM@USK_V8[F
PN=7=:!.D>^G09N7.Q?>N7JL,_5-?E[#)>>WSK55(6$%DEL\5BX9&%0ZIUH9-+L:4
P;,K*3UI(0-'N#J_8;-0^HQA&SV;#617C,7*E<[2:9=IBEHQO6[K.<>@?)CCT;TTU
P=!(BO4LH1;NZ66+/YDL#3J5Q<6"+G%^Z<!>4TXW/(]R)PYQ6@;>+NHH&^=^.+@YE
P\V@IG4618Y$V+PXNCA!^UN;F6CE2>_M0%N.@)?$G@Y[!=AI?VD9PUX;I#?[9'VOW
POZ=%2!OA  S;(\O3M&C]+(O$GMF]WL-MAI_A]+YXQ'QR(*HDYM7'R0?N3M(CTAT,
PX+NOZ$!I3M2*GCOFSN-IN;0\Z#P$(@&\6[4B79]&64_XF*MAGRR#I+@-^TO0C:VH
P;\. ,#V9#KN/>NB[<V89F555QZL54WY-U])S,U/%_MP5H!)IS(N+=1+QMX(052!1
P7Y3Q)O%#YZ*2]V+B/0#:P$=PE% P'/@-DJ1LLS=<S%=;Y,<9$W11)V9>)04J+M6-
PLM)8]=MBNLK![C0:D#)X/]NV0;&SL)[,*+-^ O?6!DKB62=]Y04Q$7;I?L/GG*,(
P"2BBB-+@:K.!9(X*9=U8"VQY4B76I@EKW[YA/&BL0_>%%NEH?O].T6;C4N"*"TCD
PS):=WE]8)$4G\U^F:':7.'H9+/@>I]5DF(@OM.A4A@:@3"%F$5^_ 2&5X>XN@I:U
PIX3=6[066L3C&1]WMLSV@ZG0SRA9O!;ATUCX#^0L6GAS7G15JG55_NA'("M2I%EN
P$[NSLVRJ!?C_(WAD@DM@-%A"'*=$2N#=&5&FUA2[F0$1H.BC%!OSX1(L F%2GG\$
P)E6MM[8,<=9JA+0ZRJJ&YQ.7[5K=_W>)R@&-2<?M_UV, QIITRZJ3K@0%>/R=/V;
PB!.$]A6E(O.MA8\80IZ;,:*3]IE#E7]ZM3==O?!M5KY<%A'54"\2=I%"?X!)_$DR
PTAQL.\%XL%[@++U/U]I0.A'.%(H]@-2MAO#H@C4=3"S9?PYDEI-+KONM_$H1?'3>
P^P HZ.5\[%JYMSIY5=NICHI?Q-K$4/BX9?=-H)/)4D-#J*)'?"[U-DNQEP=W,VC"
P $R?\JI#W4^=<,'>1?OU%:F_W7,=I76XI(Z0_WQ[J;J;%P>K==BA6/9$DX>8'N19
PHN&?:JWK<Y-G+!T+@YON6HI\$V7D'4F'GIWD+P$FTR&UA(BEB]G99=Y2G',!@4MH
P#7M' H)/^_-VI.H^+_=01';CU[T;JIIDA^;U N:;TE)E5U6$TTI*/0.CSLX%V><P
P,*?:?1<\K'E@S^.[G7$1_!XOT:_+_2-?[:S*2V)RIPH!7__@%N+F'E[>'K Y O)/
P,05@GH<SD<EC2S7\&[,<\;/X^X^W#'"^&WUAD '[FG0?\J#*'O:D<%%VR!2PI<SS
PZT+(E?.V<O$^#*UF**5 5ISDT;3[C+"W%/AWLU65HWP<(TC-FR7%,:87-Y2+E,-D
P3KU2('O#I;/3V\ZW2Z(T%O[]XV'/"Q#@I^$X$I?:Y4<K_0:!IO#=XHCI@JGH<=>[
P=Y@^EKMK5OZV6\V)4BM%0")E-^PR-$!2%("?$E/OS/_2PN@&TF.ZV3US60N]LM%0
P+F:;'A!B_J8V50S=71-._A?V2_;:,- 8'P3D#'"(8F2VSQ2?"FD7['X2?\J,]0G&
P0-@CU_RMW=9$K$JE2V?:C)RC"7P:CR(.@]?+I@552$.X'XU!)2^/2WGYWFRASE=S
P] N#UI9#HHM1-L<_BX.V2-DO?H-\+PBND* &3 4!A"+PK7,Z>,T&B2%97&7)X=HQ
P:],356!"PE9M$+(BT,FASVG0[1[J-<.Z4&V^;,L>8N:3'4*ZKFP*W-5+?T?<K#T/
P+).Q:\O&3@,IQC\0N?9(K77^N[3>6Z%G.1"L\SH*._[Q6Y(G(BA;EUKX^*&[&!M:
P\.K)]C@YSB2T=J2U>Q8>_2U+BP($06&%YWA&?7(7L((:XFL=0KLAOIM+_HT\R9"@
P$<!9QG(<DP:$[X6SQ0RR=GVC6[5N!;U57;GN;K/*F[3<89L2;CG(:Z&F.UB(>8OU
P#(<P&7RSA;JD"+(/=2/!FT5_]L%II79+=JQL-;@3 GY>)9K$6Z'QO\@>.4<<!%72
PH>9IQI4K,.&-\()70HFR+Y37$OPY$QY;-22@.6<+/HVDGAVO4?0SI=)Z+5V\&&,3
P*CQ-3:.=\5EX,->MDL8[P\B^M_#36@S+7D=.CH?OF2[[V8/W>PRKV8YZJ-^48OX,
P$W@S+G484&-[6H[S4%'D^Q+2! ?-X*AEDDOC"VQ0)RI84?W%O&MA)]Q;0/RUC08 
P6%'Z]9NS61:7D?Q>RB& MDKWW*D_<"#+M(NWNZN1@X94J8;8N2- F/'PE.$HBD@@
P,+KD"J64Z#::##(?G"6?\]+OW^N^P'VY3-=FT=><6XK=_O$U?L4-'+M)4E;GFO+D
P?( F394:?EHT%J=K>-].N>P5\C^G'4,IKH^4H7!B[P<O$)T#ERN.HX93$/XT?X;2
PI/EO$78K8E^4[3"UXIM"VN5VD^KA\Y&$Y1WRMQ,"K[W#C51+U^/0QTQS(:V;1H%B
PJU6I)#N#Q+[[8:ND6=HZ[V>;'\(=-RRN&R4W^0"@;6U=B%.VORLC1MW&<?6PHY8W
P!?ZW>I6%N$%W4S-#R6UR'Z&4//",M_=L<@D< L]VFGLG)Q1;O,[SU^GI(MR!:43P
P&-RU(B:5H9XBVB=Y9R9?>1PWV:#A)0Q&]EPJ0@(='VT %UA\E+#0Z2'2DD5: P;]
P+:DI*$U+F3W=G#JFO"UHLZ8C<P>#X2"0JJ/ED)Q8.<09\G"5^I-<" FA;"\.RRXH
PN>H=NT5ND$EE0X9LG*"@-YA(MDZ9::82R_FUD<U\OSC!GY=XH8M0OM)M+(]O?^Y_
PX2$=NW\.C3#%+^FK:Y Z2G$)R0ZC@!?2 )@>&K@: N,PGAL$\!QV;6)_W"35CG:@
PB3O98YU&''8GQ.G]?V,W\29BZ9(^&-<GM2<A U>I$/HJ64>G4("+4%B'[:_?N;+C
P%Q%@]3MG!S I%P!/[*D@-1\C_SH*%@=%[&?B*HK)*A!!URA![&]25:[+<C>JX.'R
PRJ1_E2&.VQ7DQOEIHHF ;V51ON^U-B<I'B85*.HX*-0FQ/'5A)CK^9T L9_[<+V&
PH260[R&OMB1"QGE^X\)F:#;$+(D;3GF=^9HN++EFH4$M 3J8Y)(L[^7XT(\"Z50;
PD^_G(]&!LWP:!-L>"SFLY\#2.X7 GZ]NJK=!Q 3POS:UEZL0Q6<*CG#G;+\PS=#L
P]%LJI\ &5BL[K;T'F:O:)(_%$43(&*3L7#72$Y98]"Z8FJ:AOBGJ"Q$Q+GE<-U5(
P\L3.=5^/!*']B%T[3WR]1NVH9(@<Y%5[\0'/RKZQ^(TF4=VE<+X_?".)W'@"(9I$
P\##:-Z<";>M^G/?FB'/PU96"BP!7Q'QB10'D7T 55J!>LOGM#LT+N*OE.J/.A3V6
P%.OSJYRQ2&\SGX5Q=RPD)<*P2LZ57<#OP]',82O,"MS@//HPVD'H9EPY>VIJ^DCD
P>GAX[]A0%/X,7%.JILJ0EFNUKLV[%\O'U<8G0+'-/R&R"9FK$@ ()U"GRB;ECB89
P_GF#-FB$MU$&D.@AP^KMVH_*K%NF#CS?, IK(?1!)6WP7\FZA=IA>XBE<@J%,>J^
P-K\J.8,ZV?%</C[N9 )TKFE=XD':-?;B\YBH^'*E<&K?4Y]0W%K]^<Y$O4,-O,-0
P8G?1JM,/=1F2$+^D*C %YV[_Y<%NK;ZEMUX"?TS.)937?-)*7-+A\T.:R]V)RNX^
P%EX$X242R?(FXW@X>L/*8W]PA )#/FB 9@W'#D[8,R[2>YLT#3;'8_%'%O;U.-#U
P9ZCQV^1S?T3&XOATKHY5[4EW# [O_^HS3KNU9M4%%A/5,5NKL_V"\PZOD,E>9TP)
PK;^P!?Y@F15-(;RG\\']JE#NTAQQ98P/^=N>PA+:9C;F^;VWY$-*8XFS;;@%<T[+
P@B@<2YDE6-.1Y *DF["+&?ZFJS%?RS54SPAM/)^9'?6>/Y!NG/LTAT*R;JGXV2#=
PY4,%4ZCAEYKZPGH4X 9N_<NCRKWOM?$CU'C GO3YZ&D*>XTER"<8CGH>V.C[$4^"
PGDAK7*I!TYN8)P4@[Q5B0,*\1\F(@RB&.+*JI\6K8%<BS2E7?8T/N;(V4DS01)O.
P?/?FR&S6.[K?UE42_Q5*HL-SQJP7E.9D+_^2S=_4^UEXDF(?V^J /7(#/9FRBM3F
P&13:ZYRRDY*/\8#VZ339P[-A1FC12-TTJ"1FRN96(+>'_<TSG@$&9CT:0/GXPL]S
PDWFM=A4GCQB3GZ3Y;^^@999C*$2%&Y!/MKY;6EZ1A6KCF_%Z:XA1KU>3 C*P8GK^
P$3/L( ;O2ZL#,Z,K1$I8G LR2= <?X%)AD:3'NJ%F;K2ZNP[[%>;6]0FRS'2_#>D
P!7X(S=2>X B,F;A&1ZBDMN-\+%2%&[A1=[KRT&%(PS8T(#IXL70'(PZ3SLQ1]OG/
P%ZMV#,D,^ #&Z3>NK_L_6*1^6VCW1P1?9 1_6H9,08LS3!U6#UU5E+M *#/D08T5
P(!V9R<5TN.)5_WL3]*M[->';]%%4J9T/B9/S#4C*A, L]3NF<7HO<C )PXTGR^$C
P*5WZZB1[/E.S+2HB>$VD)91._LSD4*BQ/HPHK0'Z/&J"?;MUVDR$OZ"Y7H6=;</L
PSWE IDG$'^[YL.ZO?VPH+@9=>0#&[#+1?LW ZA)3 L]>@X&'X9\TV<S.6RR<R.2L
P6EFA ]5PGP6]W,^"BDU3K^MA9OD_[W)9GL>&2)(PL-?+*/JY"E;G3HV$)WJB'Z^^
PGSOG%5]SU_<=7?UZ1G9W_PKV8O86H&I ])5\Q]+GRAY7%GP*Q#_#=F8,VL&_"H5J
P,D9N+ER%Q?GFJM]MWI&D;U?]UEF*83!#LS.C-M;/<B7$1DY<^K/,F[.+6+H#C*XM
P%*VZ,8,;\!/G(0E V8PW-M'8AC0:M&\U38N)A0-[Z)]%F-A#&S_W>HO4I";9^/1]
P^46E W.:SSM1> &O.H4[!A2.J_H',2&?PB88,VC"E<Z0%'H["Z4D@>1'1&-5A^\]
P/,CH:LH1RE<W]W+CM< !YD3$/5..0+X(.N*!]K%B?6IDP .<P)*6(+O'+2"A2)^]
P= )*,42$J&U&]';HZ*N[JLJNQZU=UY$'!&K;4Y@&R,P.Y*@Z2QSJE2HNQE;%^!HJ
P0NXU9#/6.2%H9K75L;B, )K]/WREWIWE!+H[C[&ED T$X\!"897+.:##JB-Y -'B
PUR]AK/W+QC8T,TF$+\6Y>8T^X3*OT:CRC\C 0#[X%050]U/\*44-&K^U9$H?B;]=
P?=QCOV*!S0;DU@*'F^>ED#L.G4P#!*.?#V+[E'XX4QPI5"6PG"(H5JZ6I0RIQ5V/
PP)J-#T/XLF.(E2V;+5G5: VB_.*_\PU6=VZUR '!F0+APSK;LT8D//C:SCPDH;'#
P2T(/CE&3:S3@TGY6!0)4BB :?I WZ,-B7/;(\$NV#\!:V'5^\6FI5=8KL-]! [ID
PW0/R^FTF&6Q!Y !G5$[*^QW<OM'29V^W%B,>X7!9RV/P'(P^G8LM*P"M^0$ #$DA
P[S19>K(!.8";G@Z;WP#'+Q4*O,W"3)&U5EZ 6[^ 4@R6#EGS46+!!U2&HV#-S8Y(
P]$C$NC@6Q6XDISF^ZGL3I%&X.+[^3T\W%L@\Y!=\1!"[L'VK>)_X6Y'_=\>.9-U*
P,.M,$=IPHL-#!>*1P3\[5),$^6C+<=N+Y8%14+$PAF7\ZPJ%X-+%O0-<&D_KCQB>
P1^AU J;>3IL)X<V<[ 9TRF\V-4"9Q'7-4ER60,Q]VYQ9$7$PG,]=C;Y'HI8^PY[!
P34VL;R+#C>;31DM9[/8TS?R:[Q\KD(\4ABWS\^YPE)K]8-"F"0L $ MEY:PDLE>&
P#&3B/MU/ 7".PZ2P$O<'@^@$''V5[TR?AC,\AEV<M[7(K&'"HEN'N;/'![2=0RUH
PX8-J?IH5/YVIN M6D[[S;8P8#3HPKD2P;5(3K!53>$$Q8N?B#)Z>-WU.&9O:9NI%
PI+&[5-R^GH.N%9F283[%M!7R+:NVPXS3QXVQV7Q!NX-7?%T)%$J?D8(&+PV+2S&"
PVF<Q$"W](YCPQL9NSI5A\\MY#)M"$\</YI@RGNK.69I\IAW]ZS<DCRFG<:046.P^
PSW-BPI[L!\_MG]E4N5+HR 9C+ZD0GD5W'B<C8 \88CLBAX.^1A3)VX_TB\,A<^_4
P@#O$V>!&YS:KASVJ@Q&*0TC/1 Z7:+*E;^W,1DFU* 685I2=L62+ M16SJ]/Y:V+
P1%[ZSOD$E>?0K<N"H*VND)DF6W[%QDCC[Y[4!BF'J%[,0X+M4W,R?8OD"=.LOMA6
PN@E7K]I-0LBWJA96)]"!*U9"%%K99!R1CP;T9%YHGL^)804BYB?RKHZ2A2V+;>3'
P5;J3W&8T:+TRX2"9=OLFZ\G16T#'7J6D+NP300H"ZVO)JKPXP*0*',HXOGI9<AH,
P([*4RCW,+0<30B,M%$304(]/M,3IRZ%/S$6!(<*0T,O=W&,NZ"IM]3AVRL0@VYE&
PL<)7;$I?1&L"5\.O\XS)UL%E'D "PN7QJM\RG:90V@VJ &>N$(6Q9XOJ/@)L@0^O
P?H!MEUQ3UBNT+6K-R'.XD,'>VEP =?.8J\GD&&[V.X'S+4+-1BO[538XS&%"0(9U
PFGNC7H2,]"BJ,M=']ZZ[8II=UXG5\>XKGVC!Q_ /]<V1OYY5]R&#<K7-W]Z9[-]Z
P;6G*RR,K3HP&:]HEMOC7=[@5#)X 7"$DDH>&1K7I(D^]P05UI"!;IY_.3[7J50MA
PMLT8Y*ZY((JW>CNO4T'B1<E.4+%XDE0?4ACEK;TB3Z9AT4IA%=6AWW!Y^^KVS3NS
P3(12NAXDYT,X#W0UIJ( .<U&=-YLBJ4**/1MFX;_KML%,E(A.=5W'K3%Q9->;+.*
PK$/7>]=R62IYZ8(--.?1]U'\<;:Y[$>C#UF F%S=//!) ?HB0JXLX &S&'J-ATQ.
P \TFN%%X'1!.2]ZJ_GSU/H^,Y\EY1AK@\OB()^:*E921KJ\L;R]R@=2=SM[6>-OB
P+E:V2.GFU7-6EF_[?@&6FD:BWUP,GJ2EO-MF?TBHO4+4GOX5$6Z3^#>/J))D67!+
PL"G\-<.I.WFS^>TT^</#5,M;RNI[LA>@]<ZS_J+C 0NN0*9W8QJOI%3B3NE,*@.Y
PLF(&+4J1_^I?BHI\7C0-AAZ']Y$H122(P"2T.)NR\XJ!1$X3/W-T)B;8;T__G= 6
P>J22@CHXOE1ZTG;X>7P->VT9H"R56"=%.UIPB92_$.HGSB/12^8PAX6X5DU@]%FX
PI:&;Q2,.#N)8USHSX?F1"H";S<.GO9$:!XH37")9WC:CN4.R&'8VU6$G\HZU":+@
PFN*OM/T=+FAWLP1C="-OG%LY0GVN$TYU'HQG:4?480%@>Y/"1^V@<+T)1P@O$Q\M
P?TK #:' Z=ZNO0O_SFC)3YI6Z^%KF0W4IL;Z?OV9/SXL$'"]302:&R1K I]?+@UL
PAK>L4EH-)E9]IMA^PBYE8F >/)<L/X^'%UND766[U>;:*X7IO0[#FQ1WB;R%U3)A
P_2NAYW'9CG2M'>]4S1?[%BSSAHS2$,+S/PAJ[A.9#SQ _[.5%VCDOEQYSL?-1M;@
PS).]-6'KVC56OFEWG?)W49W[^_B4W?TF#TH/?&M(K)M>$4A!#P 53%3#+(J&5<FR
PXH:: V.J@UH>W^O]=Q8])25EJ%91I9EW[=>0OJ^#\Y.%40V#K2-J,FWE9?W.MQ%[
PE*=T;C_%!@:^2G:(5D&RA.)?:NQ7M7UDP7@=SA(A=1&$(8U8D@_7\98H"/<&P^7U
P:H 'Z/\:\IH"G\XTB;>NA0!$/G*C_ZOQ"0 \#<:UI2HIBC6[HIE#EI2X=O6$.< <
PI>SU:QE5MC[V#DQO9.PELZ+FM(\$0PC>;]NXWGH_KM! HTJU52=/<VTC_]#5)%W2
P<KABT8 F5-X02LI]Q4T33DK7>'^%;UJLES$S) \J$73DW2%]7 1K2#]2Z)+*D+V"
P,TG_TI>QRD]XA[[<ZSV)0V>Y[X3LS< ]-^@<)F&_LZQ9W? P>8MLJ6MZ!@5<RW^8
P ZJ6<\T,PQO!MG6YE+G%VKYG1M4R[GFT"_]N*C(W5X@*.4R'=YIYS-L=HMW.IZV@
POR)ECWO^"1,HD^W(2Y$8-*4W$H;A*"($#3D5UL5J)6O;J@C*Q.L?= ^^T*N.=5!+
PZ[:R.=#&3 (%H.6\Z>;DT-*GE['JSU(JNJIH<#MQC'/:>'K"?\E<1%C9"W1;93]&
P\T6=54C%B3Y@,/8Z#Z._4K?//M## #5B)B&]X<S3?$._*,%NJ%>-8])LT6$1C%H[
PA+;ZK)@MA@"XK<(C.9]JXFG6DG42<,=>!X ;6N_1'.&U>\7K-89]:V2A05)IM-+[
PTL[G2Z62!1_\L%$BQ5'"7WEJ2/XN1UM35U]<3P3M42L#EUR;V&0L9,[(X+Z0&P6$
PL6FY],4+/SH@Y>Q^(!2@KU@U55CFJ<!LX1K9H</ P1_\Q<R;>QNI\8_1=/HW- KS
PDK\VP";7G@R47CV<N$X3VD4_O\TO2,^NL8<55=K^ RU>2V:+!Y6A??<]E",7J(?7
PF/HX8[< M%]D2)RIAQ4%].8(D_L"R%0A1:BS\V_Q"9DQSS@!G>@,3:(]$'$)\^!V
P@AS@58<1=P6O!:\^),02+)D/":M@N_@AAS354U4YUWJ.3!^9W_DCP";A:T8>*M-[
P HD#&UHRQ"8=-&%B9J0W8$"*FF@@QTAQHYVEJP@)L]LH(=*R7]TH^)7 GM?"@S68
P=F[@V \5U$T\Z9CN4HG>$8L3PT3R"X2G<O(?&ZL_LI2=.#6I0/T;BMSC_7B;?!6/
P;D;VLJC8XSZ%88@84"^&FF6+7EW LZ_K(V'-R0T3BJ>5<<@'!?T*"0E5WA'L'*74
P,6]X^2=<V@L[JZ$9CBYMAU5(2[LT<1:S1DK4NU>M3?D.9"?213-\S3M$]IE95*?5
PF!H["?VC%[B]D*[7[-VE)-.L2WYM!HWHA+DA/>V$'U$RZZW.DY^?PE3Q4V+)E>@1
PIOMYLM,P[$R01665L@H>QZ7FE4-"Y_D4OC)2 &@*RY'8EVM2EX7V?Q9ZPIJD9@C2
PQ=M!*YZ*4-@J_S7KI*9/H$E)FCS3,B]C&Z?P5F1H 'O:%[N?L;;AAKGY>*EACF<.
PN)<]%19#YW2;B3_O6*22IN'12/VV,]L%*ZYL'*-YKN'%'YB2XNUE-?EXO1-["7@?
PUQ:3E?3IA1@[M8%C;,QFDUN?]#: (F7VZZJ8(FFR6Y.6.7.JY6-DZ'1GFEH='(R\
PBGJ=>@+3QYSO7./&Q.6(FD8;\7%SW)UIX'#JR"R^,RXJG?T)X-+A'WF#UI2;?4S6
POY.#GYTK)$6\<"5RQR(V.3HPB7('0F1M)@4K;9C5@[Y'DUV1)0(:.=6 K%OIT# (
P3&R'DR")J951IT&7;W+*8T3A7F&_[SXP9)V;2^.'AWINZ36QT:9%,18S0+[!BEM2
P*L^6$-_7TE5Y8FBS9#$CVL45*&!@ ..6LVT974H;2VBLZIZ-A8+7NRA#+:W',QK'
PYCS=*O*4Z\9/WDGRL%J2^$Z#"Z%2\@\0?WVA.GJE]%FTW<LM/H@4/='&9$.>< "W
PXZ.?DI#7>)17I7:)45^VWIK@!#Z!^D"NO/C#?8!:VS"18D"I1N?6OSAMS'N^IV-^
P9"\!,:A_#VLH_]@-/F#@L8_=E0?=CAZZ5$#E%PO.\_O1XK,=6@]BDMMW6];[8_&0
PIP$RI;]8Q6MLI-.*XIC0.YG=VM=F+=_+@6>912N:69LC1_R<!4.M!\###O,US@V.
PY96X&Q_&F./75I\MM*%]5KKN'=M-A@CLA*SM[1GB0]Q!'G7'*-G@1C0JS!1E70JH
P',EP?X_$/B<S @H(Q>ZUD*G3GYB>$H0ENL+WL&!^PMS!IJ1%K9OF4SC+V6!_"R6Z
P(YK$<O-=M#MX ;41,$D3&'IL8GSZ@09:J!R=2$IG-$7B5_N=$)3>"T".GE^1()-J
PU)-KHK,K /3(!L9*9062A2__GU-8H.;0L&9R*]BD=0\08[%RS$8O_N*FS,F^/>VH
P%[.+5%60,,,";-1X+':[4ZW?(PM0CA@S^*M7;YP]0Z4*=SR -^+8SR=W@#WK@KZD
P#V<^-2'KQ:%(H4H/HUX#=&>2TX^&=L'RN6,+?(2L8L I1U@>JF+G5/-%A](\4BY"
PFW+R[OB!;Q;7GL)L;\$J44;C'I+(/RF5K'!I(%1-1^ET>O#3DS"Q?1#50_P15PB6
P"EG8TC7DK;-XOPQ0@!L1762"#MV+VU]6:38S5SB5"-(<XS8CF$@A.W]X C8:S-$/
P'R@$72Z PFAA/,$9#(]*Y1']E5AU'$\'*6<;/W<3"?>@BU'8MPKK7[FL!\JG+&5,
P'1#]NV^YCE2NA(0%\(B*%<:^50'Z*:USNVJ&$2E[XP\E8)R<6B18S_D-7Z@'B"^[
P* '+'X=%^F,#8+W<P8J+-(RX]\<$LRWK^?X5B\=@8KG7QI=6,=;+P(0KAI$J0O2%
PI^V*0\B14OY#J%%\\6UN0TQYO6P/5ZXS9\Q"RYC)>P2LU*0VQ#X/Z-6)Y!H<53P8
P(_S>R^QN)/)M<KZTNW,)$T5>!'?P)G]PWJ8OQR5MF_JY)I$J2R1MDW^/RU^2"8-V
P-*W0CF>;<<CFK)Z%K3RQXTB##NL(L?H&#]J2\GI.69V%=+(B'%)6&Q\(FHX0WK%4
P2;9*"X*XER!6JOWI8"6>PASD<U!LTDM#+6,/44MM,.?]^SSRI$)2R\0>3,=7JC.)
P"P"V4)@GB. XRS5T&8[OK=/Z(.SDN_0AY,I'Q)(B4[&/M4.6H/5XZ$R";@(N34;7
PV2S"O" =)R@&08#3WC5;45]2"Z=='K_!=S<[K5+K%Z(K"',;G!)R<"5KW=*H;=SM
PQ:S>V(P)?ROCP_&I#J*0/.]I7&J+@4B85WW)%LMOI.M,UX$\4HF T@S)S;5 :+2N
P\6+GNTQ#ZQZN':559*9NM@X3^M-GQC HOSU5,XV%],K<)8>]CHAUO9A<>1/KYT1;
PF>N6#$K!'W 7I)."IAV$+J^Y\:4^,8RP(T?<8MJ<BT6(7N$_TK%1%/:<9T9;;TWE
PXY5Y (574$4/>]\$^S15ZL)<@_#L:B_29YQA%#68G"D#O7RN8S;=YYHJTFCQ>O$Z
P\-\DI:Q?"B^GQ5:&-VO^)B"X!P9..C0X8G,.Z83B&N4E(>S/RF0],=GZER(1.)S(
P[44G7]^4\YC[+%P6"1^^N8ANL5J1@TP&$("A']!.WK%^KF$_1^SW$R[7%5<0L">0
P#TC8@(_&ZXR965Q*"L7[ %>BK+PHOB]%'(S;<C?WSH'$JT18@226=D^\XQ=WT\=?
P3'6=$^,?);,.:E?WO6!-TR[GMK8WDX'BXIM,-DK&K$/G<WQN)5]- "%$<H%TJL;=
P?2CA/SF$^(KDX[T!K62#![N9;*9.&)ZN3:7-@632L7,<A-NI0Z:OO@-"=*6U5HF0
P805&UC6[UH,M,,]!GE/VH5*_4M+<YM'R96V^LRA3$9]C4G^*@QRPT#JK[D+I.KH)
PR!5WV@6I=^ Q;;R,(BT_Z)1Z\(+>=RZ3TR #&V>%F<)H=W0$2"^Z(\+SA<L4_#6E
PYF'>!+\\OT,LL: ](PBRVB/8<S^;D"7H;Y :PXQD[6DG0FO$YGF] YU/6!EFM9JX
P!;7X-[HG, +(5D CVU/ONJK3)YZ-)=?:-G6;CUKQ&#[U-T%78JX6O5,N?E9QI*?/
P*GQ1O91O>W,(U R4.,"0@>6'G<6YW^2R$1%;44V_N& JJAJ_+_0*?]=44&1;E1-(
P*".%_<_[V&-?&7&RGZ#'#-4.MJMF*D@'.-E5N_T$">V_@9H.X,Q'<3F-T^FNI%')
PO3_S40BHC2V2DXM0+S>YH?OG<S?5)F#)8-CX/L%W!:"_$<=!3L00 ..C6/,[8K3E
P\#]1UW9[>S4,=UJQYZLJ3!W!-X-)<'!\2CY7YV8J*QB9S+.C!&9"^D%"KT!".84P
PF(>.O8J*PW>ND6;VZ__^#.N="@DI/O_BVQ/!GJG,':H9)PN#)FKZ=[/)?-/'5V3!
P<D97COEJ@\6AC"#N/K0;R:S]&]9]!CH*$%@6TW^@25?2-NM9[K/]JY-J4ZIH[U8)
P*3>69H[#X]*'0;$66/GS%2(8 >0<Y(*H8N>M!JP\.=!P/G9.=A9:&2 2$--@M(;R
P[#G9TMO5*)]H$U(CEZR$^D0;EJC>9G2Y!$Z%C%#A&YTZ6^ K875I1_(@GU)I3KHO
P<PY42>^IH[H9A YJKXQ*U";M1.4[>I=PF!F('[5 VU9,GF8+;(HT3$0WC*4HX'>B
PY]L."*2.P?S^<D0JNAJ+,U^:D%;6']"P9["@E(L?(#R3RFH9VBC1?W?;I!?#Q!(J
P202=_L*A1<1D\+M!VNPHRC> 4:O#-L3GG%\=V7T"[4_%:LG)M#BU*PCW2$"&@AQU
PYF3 Y,:&UT8!.6-$AOL-)<_GGS=M.(NV#/S CY0HZ8Y/]R\_<(--RA=B-WU#$PFQ
PQT7B3]>=0GQC\;->Q+6@NU$O!)VNK )ZP?L]:A"E/S'$JOV\[+MK*VZ,-_TT-XEN
P%19\?W>)F^)GC:4AKM5,0L!IW* 8)Y1IR?EB&RDNQFJQ_Q$-(D)PH:SOV>-L. R-
PJY&=OM(VJ1Y';F^[%,[9NRNQZ#WTZ$&HJX ,IC>G\A9;O.ITFP;2TN@UR:2=&?X]
P)B!ZD7?0F<Z0.,\ 3V'MGQDM*YB]=<D'W#TK:Z-@O1JA)YM/,H<[T5X!W*\V =><
P871EY8M.1:'+@-R,Y]<2Q$007H$P=0-Q#&V'D;(/M?';H&8$QC$4LWA$, 8'>(^S
P*J/LGO7&QY70V76'$1JE]HU:*R7I1L(>#NY2!/A$EL,9,&73?-<"'8WPBASX,<?L
P?E#.W59F\0]6-#/24AJP8B-<6"[$OQ7?*U/.?6S\";-RY?(D[/BNU5Q8!!>'UW"H
PV<'HHT6ENL-SXQCU+WTZO"KM$)]#$%<1Y)&D >U>$P$X!A6!:-$X#U 2\"8;7RW!
P4V[+&[4(,4>-6_@GV280R691DNL)#&M5RV>4Z5PN#<;0S;:HJRGQ)PR+X09\OL04
P>/P&T.U(6[X1 H03!R@$?54H;T1DM6<E)<X%;T\6F0-HD-W.R]!E,F(,UT\D=.JR
P:B/+BX3@U(U.5-0<I'6/0W/[-#M9#4!#BTF]S3PKIT+IW9CYAG"*';\:/V&"_7H:
P7;!_?;%:!YBAX\_BN#]?7D3-C 959Z&%5WYK=8M=6+AD+>SE6B%9\*(-'NP3%QS0
P&4^<Q4L5"_+;T9ZOZ;Q[$UR!FR46=D-[-E?&F?-/MIC0696&LEX2\</6)G*H+SY,
P,;X*E D.1C@:ET;-D-2:\I-9''X%D:NX"(L8^2V>,7_@ A?F$\MU!RJ+=#HB&[IK
P! /)QR7IK2>PY[R><%P2+21R;J%#HS3F=?_R)T\OI53LM+"WTTVCL7LC1EG93=_G
P)955=)/(60D<T']UTEI!%Q:D$",VJG?&/;^-GY7XXS70[\2+S/O':2$G&\2?Y@"-
P:GM,JOU?3':>TW8D;J\]I"(S2]":]XFEW%:7?)F!LY (V06%E =#-UZ\,=@=0QD)
P^] X/^J7,+*U-X?1%9@0#A6^U]HH^R-M'@>9DP$:T)BO>GD^BF"C\*OTFEVE#E74
PW[\_Y7BI.V)H V67JD^ 68EG\&-![^?.+\01#[;0-U9',C\_511RKVG.W(A#T96@
P/HH UQI$G_B)N<<4'[ 1X#T=A"V+&?D4 <&P2YP&[GJF47C)=L$)\\F_F]V\R%+G
P&*Y_8FKJIO22K>,@]>9_%%75-/W9R/JPY\5_@P\L]0/3MT@9:72MS*-I]^"?:C,U
PQ3&B.7#G=0J!U$_@-(@BIV0J9CJ%.,T\.-#B@;1+D=NJK'^$RK%("+SW7TOR\=CQ
P+C/"1F\=OY5PSM9^8=NF *1CD'?Q5"930J[&H7;XGWS@@D1)Z<9]*XWS@HG-R$GR
PTO"P:)(CK^U"X!VI&)_%CM ]2)Y/(1WEH4S[_/$G3FDMUEN4:M??"Y*046A7&;GX
PX#ABR49>(U<Q>Z?V37EPCFRNBJ$79V(VFZ(]VG%_C-DK")'#AVRABDS=- 8?G!I\
PJBSU:^#6EN9Z4^W8M, V)<__\8I$+!YDH#G88KD\V9>@&=UD/,9RUVG\EP.IP4V.
P8CTMBRW(;-1AQ(8DHAIH]AZ7O(;)(4O[KNVSWD(S.W$AD*0I2=Z8LL#UI%SUX1G9
PUQ(Q<<'@2/8]XLY!>4O!6[V$_&)[I-'WWW:1_SF,+EN]I.9P8BSBZ9&+4=&X+L&W
PI2+1BFN*CPGNG!GFBH1! TR7N5D5$1!/1 \YZ==%J8$"NZ=;!W2K53W4?54J\/0#
P!Y.0#9>RYGC[3)-I>LMOF4T9."UWBZ$JHU5'ZX!^2Q!GZP0^6 ''R]Q">/VH"%GQ
P1O?/P"2S22ZQ.@\ YY\\/TK,L?21<NP?U3*#3<)P[2V&LA?@H!09QV-VT-3>Q>)+
PKZ!F7XAG56.G>26!9W=ER-!C/PU\MS\[  8[#!,#&4$G,23'A""XT!BV$?U'3WR)
PVK?P]$UM"G/VS^<Y&K*ZG>-'SJ>$GVOVO=JO$<2O" E8<N .Y)M;/%F4JR.-:R99
PX+:#W!,'#W'_N*/0?4.*W0_(+J<*R+MFT$2#!"H]25A)=YVMJ,RI!;&W>FF?9F#!
P__@3A=+ :0HT0]> 0-/=>Z2QNSV*6:W;*/&,:%00#;_IC83D9&KT_F5OQQ3-[>@U
PE<=1R-*C:S09@Y._<J)Y?Y?OVZV&.9X?X]E&0(OM'UR?/=9<K1SOTUB5#(65*4GY
PSH]*B.>JH=3 -&0N<I.G-H<\=0^YA4><3YKAZX$@U'$(&C5PJNTTOS([T_+(,M]\
P.5F"K-=4647Y1AB?X+:@ BEYT"7^R!!H'U+T7RR7')'L!F09N4:EN@-9!*'SZA!2
P#[]*V<A4(\^3^G9+!C:9RG(#70/B<V*?%5$GZ'Y46U0QE)4JI+S390&^*FDQ<2KO
PK<>1AET@UELU85R')%,,U_[J*^J*_#O.P@6XG =U3@\BC(/,?4@R=NU0>W?8=@I@
PP(K:_(5CK@A5]!642[XJ>6-;+H4\ (=Q4YF'A(^,BIA8KP +/J?2A<$Y/H.=>B<7
P(C.IV%;?"J62BA[8UC<S6,$]S4?0)*6,]8OA]C7.$M5Z+>AKW-P$G5OQ35.J6+QA
P!8V:9D88046OI[.)<N*8\#Z78(:S;@S(C\RS%$![R\E)46<8^JTG &'N$H% Y 'W
PU]RR@&71MTJD<@TZN3U\S/X.;" NY:CC4Z4R;?TI+$]!&^K@;7K^OQ= Y8UB>S/$
PHI(>8GL:;>T?VO,PN]9_XO,:1T>NZM^M%NU!A!=&@)/XSN.4VBE>+KE=7_7O4/>@
PQY[TDVEAF,CU9K1Y,"1<++^([()C) &HI1# 994(Y<4K[]M@!PPD3B36+X&T]PJ.
PR]9[F^E_>WCBC!CCR,(Z-9M'4>+A7Q:DU8 '0!N#\Y.W;4A[%>#-:J!VJ\[8@C&^
PV:]6:Y,M*I1TYM[K_D4Y^GKO[5[2UQVT) <!ZR4%OE!)(1 I!YI\>W(8.'B>A*T:
PV,TMC'<(^;30(*8-A1)D]IQ1A<3N?M;Q:IFK1!BNQSH>GF<O3-E$9S-AV^WW48P'
P_.=K6C/Z8BT-G@])XXX7UZ)NRU9AMX$V/E0[R/A_*L1IM=M0//&*/CV85'U2ILU\
P;U-5#CI1N7Z:9+.M#^5100FL,M9%,$F2 \*MB:A&7E%"I@LR(U&XDN98*<4<IB=5
PF@I2F#FGR?*84@OL*0/(!5&EJD@DGKX+TZH![^S(]^?P)ZAYMH&->.$7EI5J-[M=
P\TF9I)BGO+(>X\IPG"B<X4-?3Y1;^8#;+W"+4[/9+(30=!!K3^ID9G6=SOF.[].N
PNQEB-TYS/V_QNX**U:&4T^.XC%O>"@T=JBE&!*XCP'KX!I 0F"1%+[/.L+]W&(R*
P;$+EKUPT#5>DB@ U$^"H8%;<M10<Z_V'%@0KIRLH>]) #C)JF"78+,IACLO;:K3J
P8.9/:'3UK-YI#(N\-'*2&M=XMU^G^Q ]'-+HQ9?XH_62K 0YEJN4LCL4!<Q[F5K.
PR9$\CMEKR'N]JHIY47*K*#9B"<&FKMOM.M3"W_/%G-3J?ZCIQ8EQ9N8^_O(T-H4K
PV 4;_+_@4J7KDZUX2HOS$;NGHY@>?,I#^[VO#W>!+!73R2@^@QY/(P=9B%"7'\':
P> :1,3TEO* +Z2.J,ZQ':B LFXRC@1J!EGK%EAC ?GY\BR<;KH#JDDPT'G,:B)I^
PON_I'22NMR(ZO^T"T>"DX>O/0VX,M.RK(=FXV5 \ANT65PS7U9O8KT0-A<U0!K8Z
P!'],1VX7KF[G<S# U&JJQ"Z/PZ2#R$&@@> &8!/@_$\ WN7VZ^:D>[]9NS3##0<6
P.S0,1^NNT"W#Q%7G$U04<ONZ,F-?@+_O+Y@!F7K(TI_;:E19N+2MX//, P,>I7HC
P8*&@;]5L;F%C?&(8H__J52HJ(@LC?4CU! 4)J']^8W&55_)1V<ORN^!!=J<* A8H
P"N3]*5Y\I4[H-G"G \_>^UG)J-G&(2-&6AW,7Z9NA+$_X<TFZW"\ES=[XT<)L<"+
P[3QJ?,W3RE(5X6UF3MU_[!V"QPMNK>^9P@BU'490(MF9G,M"_^2=IK61]@\X2J6U
PJ>VG@RT]:1ZL)>4:,9]]Y47'TLJ2K;>USZY]9[<8F>V[I;!LCSWW[>IPYZ'14 I>
PDR45CFTOS91<4GJ%,7O&JTL%_Q :QKADY=YZMUO<]@YM:30?9]4$+,!"("67S+5!
PV P.Y5Z;3D$*3+OC*2'!]?J_B-D-"2#W]P0RGZYG(+.C95R]-0L4[(6ELKNL?U"O
PSJ0<M\4X9DL3Q\-)XE9A]NE=.(:ASV!-5F+YY];T<V5$4#D05KI^S4=$S%(&N*^+
P_3H:RQ8J!B$ $1[/2Y#%0Z(Q"<H&:_=CYKZSWU>MD[RH'3+SW/4ZU&B]S]&!*6@ 
P#'T4<7DR(CW<)6?V#\]CYTA4?3A@QU$_U!OB2]$G;Y@(?GK:7O#2!S&]TS(*W.3?
PG? V\*%O ?&7$*!*=9"C*IMR0C/H_O@0%20^,;('IB,($ ]P4G($MQ+HS=V6!17Q
P(-A U2O2F&G =3M-R:1&F%FVTZ%A'0['7@BR5H(^P!6PGRNW,)3 VA5=4DTLG9?/
PR#_8BV,+)IE$QPU'I"XL6\CLGQ:/0X/ H.F!'LY.TZ&_79/$BOP(Y8/PX1CYK^RD
P[\I0D.F:\SPS6 SFHB !)1B-^Q++60.?IIP)H U->)U/11 VC>#N<3<.PZ).N^ I
P$-"NX*^(ROI9S!A<1$W0-$8-Q%9/VPVS5>&G^C^")>]B["6, KX;ECNA=L1K?>LT
PV@^K>%E<H32(74]D\L50GX[]^XY>/)R'G /=&"C$ZFAVM6/GA-1&D"[N'T%M.&!.
PD'A 4!>'I%WY]-0AZ2  O.N6= P-$H$";/P*[\>66?)M3"+_C%YANVL _>"</\"B
PMYG,J1J_!*3<2MY2M8^]D=D*I!#$$J@2M,@'65L-F^:?V1U%0T"J2+EC<'I.N<H0
P1!(+DP_165X1)(*9,BXZ4'+]FH\^^E/!_L\X3*I>4<HT!025AQIU\2D?5M6ET5,^
P#*PCRR2I7,ILIVUQ3<T5HPD>B1@#AUWOJYV?XSXJ<:;H=P<>"V*VP2W#$4QA,54C
PU]^Y&&<[-5SN+8 X!QV!;\UH<KG3)TD%[B :\/+HK)(H)JM4"8LOM#,B\9AJEK/-
P8T+T/<<;N.$J>FTV;FY(-P65V=R-3X7C_H]1=/OMFJ'#021_;\&F_1TQ:H.0NIV'
PQNBVA#W49#Q0P ;:#MS69<PVGGIGQ4-EO'R#SB%4$0 ]?!SEM8*[P"TTOI9L7JY^
P^.XGG-6,+!ME KK\**L)\H8B[R]W6I=Z81(9A+%FH+Y-4I9@L*LA4Q##?F#3NO63
P*:IU,>304E]8S%564=*2D)A?V$-T)N85-#V Z;5/\$?7O\CZ&2V\D][3E9@/&I8S
PKV\[^QRZBA\0>S$I/2(K'L4SM$N105-@R84%Y72@UR<GICDF.262TD).9(@'Y,-8
P8">,PN/T]9NOBJ?Y!%MXVBTP9]6=M=>.F=1Y+VNB6SO40=NJ7!G;!M0\+.,0^0^=
P]&,D*3U#,%7:%85BB.KV__6(9^L#<GCD'@[E].]J=IC*R?R^L%F'A_FX(X+M#C'=
P2<)1G6I_BP+,H_)O ,\Z?\JKK*+?'-+/!)AC[B T*1IR-<4<-V6@S;'\CS#"HFE"
PJP6D'J#LOK_F4TK*-3C2/L"2P6:=$K&=PHFZU!3I4V5"T+X$S/D!-E 7?44?V;6"
PWBR*E3E^=8%?$ GM62!>P<?R%O 2#D5O30"'^JTU]>>S@-$B(Q ^X]ZC#77L8[4Y
P PDGHKXJWV#U@;%XA'Q**!2?\7LUZO! ]$_R02GOZ)=Y6* )CGFL PC24!/9@K2_
P>LXE-AENMW%6:AQ-%U\#E^":+QV#PIS3L1DA7N3>_JCZZL.<O$P8QY[L"FB'(HT<
PO%Y]\7\>S:-LQPDJ,Z5@'/TY5MH1*I#2.6I=D(8JWIBNW5:G4<W3]Q'T@O#^ZCP)
P=2\N"1.Q\$\+Y(5-(0]?)%@0<\;[(OXGK0_MG '$#9G3),\%"RC,R[H32PLV ?#*
P#[,YE%![#2AZ7:#9;)M)SPL#/OG4--Q+=R \8/S#< M[5)BS&"P3TITDZN=-W<C 
P<.7DL:DT_Y8EA&**L*0#F5VO)RZIP9;8N$)@4-F=YMKW?I^J8@Y-ZEG99J7\NP$'
PS[GA5K<%*EU&M=BE("E.?8J1!B,'B_USB(Z+[EP#@@2?A)>P[HD829ZHC*: M@Y!
P>(E ?B_#9JQD  $2<^*F\H@X1IW!FK-]:X@L_A0=21=C%*]-;G:J+'%__0$\#436
PAQH4IO/>BU4TOF7<TWCAV/MK3])J8)':<>+9Y#HD"N6A14[V=Z=%@Z$@:;1I^>X-
PLWZR[\*C++PJ>%[K.5=>>U^;.G?JM&-84$<MM4 <RG 2V5)[U %I.[9?W#MWY->,
P[)!Q\S?N0R-X9XNAEA%7#/Z+N2.8N4VFO\$V1LG@ONO8S*0?X@CB%^G(] //.B,Z
PH9M$1C"UQ,F_"O_U-[[8I3:L'#O=2'/8U"4M4&+7#/4>"K-&]G"!'GL-I5([6C(J
PQWT4W\,'B"S^5+'WQS#<9?-2)SY=Z*^D&>+6;>:UC)*4'EO>GCX(8PD)[R&%5]3.
PK"WP-W"]TAK07&+*?NS<M:H[4\;4C4]Z!.GG:5V^I!DN&4K.FU0LZ'Q(2E+0UZ<W
P5S?PWS'(+\F/1.C:-2XH7B3R&ME$>GS,-3 *9H91R_6&EK3]I$)JY>;<!>BQ)A=K
PJ(Y=;#\$4)=4$7XBTLHT8.C\):L-\X_I>P\A3K;I\\BR/#])@<?9^\:"')[K443P
P@UN%,,RF*,+MWRI*N68)&7MKZZ$<Q>.6]1GZ=0)@9(^P!I\.VHS+2"H&O=U5YQ!U
P%*1X7XAKHG>])*8&T92YB^;+Y[<FW*3*,I2,E"C_5KYZ=?">M;42'\?UZ4)FM#$X
P?:_A-%5O'=#<_>#7LJ:S@5WVE>/-C0ZW+FA4A[E.?\K![&-L'+%(Y(!=TB3[YTP>
P63@S4B4KUB>!4'F.,4=TW%LA]B=[R'R B=W7-D>#M9EAW#8%0'N"!22<3?J 2G2.
P^JM;4=JQ!< :-LJ#',%:V07!;2V[SC5ST\2B1-O\^PUB)MNM) PGNTSZ;BYRU@5V
P=94*!L$AQD6W&L_]I;LARG@4T*JN2[3%"4@?4] "@+@LR45W\(!&HW8)C1"#58$6
PWBU2XU^(C-'B'JF_N4@5;2.2D_<(5+O)H26#PY6"2\A:I,9!G8JC"$$+.>_5-:-2
P_)M\S4<,S*H#T<,ELHFG;><LM=1U])N]-BWCMB5[.1R@4"O5@]I_&>#,X"]O)LHH
PL2E1(DHGD(;$MA]EX+ST*N&'+K%OC'E8K0M4"F,BW8+&@?#@R#QQ\9HM_-(."9K"
P\ K VJ=Y 3!!P(VGPQF13J]NM-WB].57ABZ+=]T)_?5%98M_@X6ZSU*?%S]D39BN
PS[1+@IS50A5X=4X(U %9*8&]!'7,X;X#.!W;-N: :^F6+L\'.AF=FUW2?)IE$E-)
P&A$Q0Q]!4AAN?H/O/OW1OXG@\ZS\11A*YVVV'PUD^;_;_)H@Q4_6+<WCC6PLV$3M
P/E7GFSL$GV>ZJ9E8?7MK)QT?&L;^0<&Q33"^2#_K4N5!R*XG3SC.1ZP4=S6V!B%4
PUR#_]AZP^"0;[XED\>,TU(_+S&W"<Q+SYN(GF<6IC&17X:&G8$UX*N)\NG(>('RA
P=M\8HA.CO.WZM-SU\O^V]1AC>>^?NU4#BF'A/K0E$9:$%;F2Y4;(AVC*H( MY"\B
P"MT3'.=%W+J+6EX32^,I W"_,>Z($5ON#.2)G"=A*'I?LKUD+[1>=S2:B\#'@!N)
PX4P8-OU"'<N.,O=T/OYK;L@& #XZ,!XH5':?42H.G[8<_/.I3?Z&RH7 N-I2^G7Y
PA?(O#!_N^;45E2# :XFOHQ!K(*VE<VMQRQYG,Z-W6PW6_M79!#^\ND/#KO!G9+YK
P0CWU++#+5N?OV$@;W.=%=G3S+0'IQLTTB&Z &23Q>-D@>#,J1^U'S2-C=SH$(;0$
P]W#K.7ZO+2NAZ>%B*S<EUOH++;IR:N>]Z*;IOSZ)., &*0C%(HO!R;-,\3\A%D/8
PT0@1Y#K6 5.+YGH',U6MIM7@5L/H5"D0TN$#H7*GF +FO37:&;9S8AOLYOFRN'%=
PK7!MRH6QB8]IU@2T* @34FXSE+XV?*8PB-OK@EK:T/,9RN*0V&5VJ0QJDX9@* !.
P\1+.M(>Z:"DV.Q;*H @RHA&E26FQ8&,:I&RX[M^W4?28KNT*W^NZO7"MCD##7V?&
PMDV@WKE?ZH"NFN0MP/?;/U%-H]]_)R.NN&;R<G]/X^%MGB!ZH($*B6,I$F'-XZQ[
P6.2C6-"3HY()A,+AQ!"X"4I#@,,*MDR[TWJI,H3#'=W539G>\*CF2-BB.T;+ZXH1
P'<^/WL\4']B#HT)*=E='L34IVEQ%&:3W$8:;0_-W]FT<L7LC[:MMQAZC>E+V8%AW
P(#;44( ?8U)JZ/W#W]@&_1J*IH9%1BZ5Z*\ R7>#1G8>$M+6E-Y*7GK(OG6B):MX
P*3_]DP:FW@L5VX$_]%E3V:W_S$R'2F;7T_1P07</<P--!9[*S'VGJ3UB8HF8F8A2
PW/!^D)T5KK'3_/S2GB417#G+P984M@YJM9$#9:@H^E*=5]8+S1/T?R-YB)A^/8+?
PBJMQDB>3LD@\O,O6;Q)'0P32#]_'!;^@PRJ F7W:?8]@-7F8?.VRS>9EJ36RKB7F
PED6R#[NQ"Q#OQ_E0WT44HY%Q#D6;3TAO/I5D!<GI*,!GXC.O9C%\C^Z#4,^+^,2-
P3T,:A+9S.)X)!EIAWBA8F"KM;/OQL32V:XS*B#SJ'T-<'INT"YG@C6]**%IUQ?0!
PT_C@<VLI:OUI%I!G!T#?&-<KD*ON"U[\HST*$/#,-'.]T]A2 9+'>+@\HBD5>)G;
P& M$SU_&/$R^"#ZZAN&]55HVQ: PW)K\RI!2)5]?E)&ZE2I#HKGUI#BU$!+4GY9.
P1$6?(QUB*Q[_?-%N?O#L*E;"O#4HC:NC&1(Q)6U>45B7%'[*#QJ;A?(+U5*>W401
PQ\3;_*"1A13#%GU)G#W!]J0UMGMFA*W$92QLB@;UKX),<""R O)Q#)+4D$2;M!C)
PCW_#!_9E* 4#Z^^2@=&S@ O2Q^4.+G@C.TFD"&V*(V?QBS/,""F.6&=P1)>+J?&$
PN4F$ 5LC?V9L5UCG".U.M2VS3_)$_SRN'\@%.V(*[SR%$@URBY;C-1PCESJWUW9%
P;_0N)ZP9:31WG/ZL_ E'D_MDD<85_#)O&72=/:GRS'A3>J5C?O-%,B-\#3<R_@=O
PI9^GNDF&AC:8KZSP_<X%C0;L#HA?YWOJ QD*RS.2$7#<L.]..F4.>SG/<^//P^;*
P0#=DKP4DI9S(EA6,Q0WH>;%G]\O&LD$;[]KAB87"T)HY0V&6V=!?W>F5<6_W>==W
P:BSR#K6*88IW\0$]0,^J7@!/ OZU[H(>+H>NL>'>/,5!&'PD/AE"59,8T.L1$,-G
P+PH*O/+)S:WJZYP+V@%DRY9A :<F2P(Y:^\QFNZ"G_:SV9-WK()RW5WDPJ=)@7QQ
P;&DG6/_YBR(^\^':=J<*Z.&QYLN:D2:2Z!+KCDR0 \?E.N=T2<F74>0L.I1'\U0P
PH&I)#K3/Q2C_ SB_[_\< V!38?J<:\H?'>'X0'9P(UVD8>!PP^.U[BM BUCVQMVA
P5[?1I^DM6Y78E.U2*(EG?"C$"I("-,,6+*;,>+ V>"E;AL8CHK10JB=Y?JAP[77T
PN@Y_\[OG*(N##311UDI^MF)]!0#?9$%#[\F_+Y+,5H$<G<Z0O3(LS@OJ8NPO$J[C
PXKL.$\U(X3806^+6>4L\T,PQZZF$QWWV1C/=BQG230PEQ#<Z3&5G29LGCU=!YW6/
PW&F'R5GLJ-D_)9.A_5&<2^!MNZCO[3B*5;*WZ:A<V.P]<-+1<0?0Q'T0PM(OE/Y(
P6J%Z*B#X=S#Q7 3--J.;3O>^(462ZC_X.5-NLH,V]DO^BZONSG?$UZP_%!JW^Y3 
P8CWP'"6V+X?8J7J.SJ8<<PQ%$EG8!F%5JZNM,-"--QD60AK(QCVRV*0Y@:A5"?P!
P_-S('!2O_T6=M6%CCTX !7?0ZWW6((7%)/LN8]^75DLDK74<;&-K@0@H;+9*(!!_
PGL/K,#W?HOH1\VIF :'1I6L,G]\,G9"%RO5S%J#S_*_:5#7-0VW.+L4N].J<S,TC
PIVGIBL$Q?%XFS/!^UJ?60[M%]C) ZB> 2SA44W1"T]1R;$FY4XH+9,Q &P!'KM#E
P1_@?M3GV3F(<7FKG @T;G<>X-E.<6%0LEB"D;4:C\<P0J014!]@&8VXF:*CZR"&$
P$4&I!E7D@:$")2?@<D\4!N=DEHPNYYV3>1)*"/FDDG%GP4X$*U";+Y,+2R=V.Z'E
P>_W\+O#J(0UXG;7&)!#L\'HLJ*@MO&90<N1BB7_=-,&(G?K8\0$$*HR]6TWC-3$H
P!:W9Y&L^X#G@%@/6/[0R%,O>P#D8-!Z+S3<-OO9)3UZ2@_!:#3:.AP+W-ST+_AL?
P2&[R!?IL9+,F312S81N>J2X#(8_)J<R@.JQ='F65(RX$X>33N-PJ9D::C/V%,+#5
P$P9OH->2ZI+=W!1:O),,5@;U8Y=TF.Q&44Y[>RA$TI,7+.XG:-]8WL5_D^%3??M<
PN.L")5U-,H+Q4;F["Z 'I4M\ 0=33BEB0)F?F\\+3T#XJW7-+IGMC-,M#G+5=OU4
P3 ;D0J7*]<5OC%EOTK)]34@.MIZPIC2/UXZT0KZ(S5_=_23BQ]VCH+-T-E% 4R@8
PRHDX6_I3P[. 0R@SMC/Y*4]UMW<60Z%<EU0867LDGE'![=A>E(RJ%J)X&[4@]#.-
P G2>EQL;-[*M:RSX%;Q(1V_0:]<XF'XP,!=L$^1'L%V@F?W4OO++1HN>^FU2T549
P)6)"Q\4QU(4TTJX)_.MA,%)K/F U3,CQH!48%3 3@%E[%K+#8?LYC==2-+5WOX4V
P4?WYZ=I9+<)O[O] BP5OZ[4C%5-XHV6TM#5E_WJ#S:@^TP0/UW2(Q> CO^.(O1;_
PS8BQ45\_F=CIUO1LT@/AI5.:4>^=BP#K"0$4^K4*GAGT+2GASK8Y0 1=ZW3LX48I
P[UCV&QN^OEL/ :$O'>:-%QOV)B<K,JFACRK6/_K./??T%Y0YKEW*S.R!GV>$!D&F
P-]@Y4.&J1]-KE7PK*+6"4F4_\W<P^/V(:8^,\?EYT88%)'_L.!/+:CY5CFB3Z  (
PGU1?'*:T@3BGEX08Y%#HI. +C)K#C,3AJ5/2M-&DT$YTA96N7(;07((_@Y@C9 %O
P><MN2@CVCI]PA3D<VH!J!\[]\,?W">QUA*VT/XU%CMP_%KD6EALB/FV<\4<+?8U$
P6X6'E37IPFTM6U:"_=0^H"1\M#?_19RRIM3+0DT1-9ZN. ;D3AP_*G<>6=@"98E2
P1<^>C/=J37 *5,.J4T,"G>N.M8^[19KQO[$PQMIZ/.3QY,;,C<DZ:$("'GVRL@^E
PSC BAF$U/A@Z1Y"M6E?P_&'H,QES+4/FR$%^Y1SS<KC\90H]YD+5TAU;)25MI7SW
P)QEH,]FI-#3+"&D(G0Z<B!6NM)"L13F5!?VV2]_K&X,_$S)\]!V#71\3P)RT[U,#
P&!T5\][H^ZS/6\H4>LHQ_2<FXE=BNJJQ6#&:(#>@Y-XG.7,=-HG&X6(B6Z77W*==
P<$)%+'Z&(K>\():K:PBE$;,[/ "?*0U.NC >ZVU]!$J(B_62!ZPRW UWH%(Y68$2
PXU/WSD0FY)4")XC#L;9IP)9KS6H^!_=MTA,;"%GEZ78N4=>*E\-1QA/UL*]#"6_?
P2YR?.-+/);)G2>@%"T&Z?^_3@%]JF?1:ZK$>?.G5A1_B#JDPY3%GNS"NGV?%=EZW
P&KH_?(^T"P=CR!=4N 70N_\$B!:VB)XK!'47/L4V-&WO-NHZYY@WR2E0.*,K*2+Q
P^,,Z\S&+(2$%*:CUZSY,[)@1#XNS^WLHY^YPBH4PI)LDNEES(>3?&H&@8$1]%8/G
P>=6N]173:0E!T!: K23[O:_%%,0KE3BZ+;S<!+9W7-Q;T#*S_,E8ZN^EH:^V17!.
P0(6NF7V>.F$(=B#"5Z!R=$7IX?IQ<PV:%RNQ\<B\"4,S7DWB%7_*9:Q,>)L2 G#[
P/2JTSO[*Y38U20YTS>>85J:CZ.;PZWN&;7R<:R9&%J#6,W+HS;WJ,7<54^-'7<<!
PFP?^^G>\<[)&]PG)1$%NO%**F,=5R!$&,6:WU.R^[:4HS^QT_8%/V;%2NXX\C&W*
P-.%@39Q:M%1T^_YH0'VH6VAHW'+_ )NT%/*IR+Y*'<J". B=/2F],K)E984@?$S\
P)I'0"(R;$CC;?A28+\[Q[W!=D \;,A5X!L*1))<!1;IENUBFOUK>1D:21L//IU@M
P80:%@X4-*3-80-PZX36OD3C[8)YO.>%%(5 1Z.]'DEZF;F5IHEM3U4ZO>G_2CO1,
P0'YMM-/8@AQ[T3AK?"SJX*G16&7!.=O:?;OYS@/-\8>T+Z/<7M54S<H:+/21 [DT
P. )PN)U ],0GK_$Y(<J=HDR$ #P#Z*8>?P.#,_Q-0;VF R\>NME1-VNBYU);*_&,
P@009/KP15R! G=;K(XU09874[+O?/T5Z5!7(\O8$E50!?'^/: 70B5(J"AK<>,N4
P3 B;@%Z85D*T*:>5)2>QK02!((0B1#K/3Z:":2U1*(/6A8_6@-",[10>\;CE!WO3
PO3E<TZ?&L:6J,F=(MX*42PMN&T* F?2!:U$N7KU8-2TW,WAA9\)E&TL]6E+5AKRO
P*$?8'@JZTP.R9_HUV<G\+E)UL28CHWU^<$ *@:G'RZS-3-^FDC+KY42":<,S_+A@
P>U U=\TH N8*9.,:7N&M\^[Q&WM1=8/?9T(22E:?I-#F\"#;]_D:N9G(+&)T>..$
P<89G!9I>N$40V>;6)_@?LE.?=JW2]\][,[_TKB&)[^\TJOQA7OU8&ZV$E\Q=?BQB
PB(<Z4U=?(E5]^I;.%\ETYL^;\^37^=_U7Y3./7S\"$]QY7QXGZ\BD? IROQ?6F4W
P%C(\S6E7ARY@M=L[3^'N<<SD,04#2\"J5ARYF._O2BZ\*A)E&PV@!9L&PII6:@09
PUXKIC:=UFL<Q'^HXC>G4*%GI%]HIJTRRT(3EA 2M)4;9EKUVEJQ=6+DQO=Q[4[:Q
PCV=J\UW/@96U-S)5OX"/0\CNMD$W#@DQOR.LB>E%?-HV2H\LB6+MK23E],<$WWP!
PGWDA6$#ORL/E:RARMBN.C' ;X>E9VH#*T;5%,/,XAO7X@\Q'UPDU+L1AYA[A[(7M
P:-6V8,J6D9U("/N126XB8,OT$I;IT*"LLC.]./WSIVEHF@(\5G!/,EVSK<Q#I;/C
PH'AS=+@+88QJA(1VVT231XQ\,K-IR1?:L"]VFD[:)/CPQ)=;?(;\+@*%A+-QUZC/
PW$\Q8[0G"-Y13<,/:3*2(Q*$*D& MGU%A.[@ (//G80;#S=98B$BMJ-#P_93^B/I
P NEM&H!Q>5?JA7)/!?CLL;-19M$H_ZVDD4X^[S("B68C?\QK^)];?T$%(?$\ZK67
PP,X<ELE;IAHQ7**"?28^JUO0B<3?4$IG0:LEI]@<-+M -;>FH:^L[5/GFNA?-4VZ
P>],\$GXZP!5X0199DW>!=ZQ.ZF5DGX7)#CXY,)ZSR1T)&6F& 0PPS+^Z"^GOS3E&
P V>GT+:ENBNJO/UC03+,*Q :WN"<][AF,AU:4S10!OG:<0RRTCF=+Y40.U3%AO12
P*>78;6I' )#!X>":J/0Q8.E9_G#ZSX^#RX*AV#0;, _5WY?]]T-%8-4>L*A\J$5%
P5#S'VQ"CY>K)(";,B9E(T4BOAW$)U-%F>&QTKDR*7\1KQPJWF49:72/7)/69T$_K
PZI\*Y=&195S@AH:3\"I^K$I:"4L8%7<E^N"+E8#KDDH@N;O3E6S]!_AGVK);G<I\
P?]J ]6;893._(5 KQ/I8A>I3+CZ[4>NYF &G$L26U# AM<20.+\TFUOKBE>IZVL8
P#0K[",YVE=T1Y^&I@)#5"L-,I3[E)6V\L:W>H3\O1>P+PK@-0.I]25 @"@%\U>CP
P9%/ #2ROXK8Z#U!L@^\LZ.K>:U 4'\*\OG-+,P9^/ZZ9*'Q>\+9KP!07*@[MWD!*
P'T# &ZMP+FDFF9RJS,RW5NS(#@*;ZY*+SH^!K/RX[&EATUT[@0D-?.^B"MTEQ $U
P4$[BPSI]]XYCX;^XN,<Q=I_(TH3<K%UE,3QF+ZS,DF=M^6M^ A&#<HEY;5;L2E6-
PVGM*'NO _Y[/FV?R0=7(]NSJT'6@?=4P*Z+2[,Y$OFHLZRQ>I3EGPYFZ,B?H_S+4
P"CTIDPR $4/7BJU6YY%$2.TKW6&ZF^P/LC@_^JC^9@%S259G7=^FS% \URXFB'@U
P#A(R[S?':/;),M?@/LFW *ROR)@_;OIBG8[L]TW?DN)\"&=VM(1-VE<BAWTQ"<!J
PA@,'%(I7Q)^_"&$!A^=[CQD-D7^443QRL>'?+90^*;\27Y."![@H'IEX1AG@MY;N
P@$2E5+;K/G<+P'74O*P[?64N10DN8I[#KG&2C-_"O0?VREP%"E5-[&XG@?G0!OV1
PP/"^O1L2TH-'*!X>D1]7*ME&YB]^2#@M_?#FLN-*6X%^14[6\%QSM6Y^QR(I.6C.
PL]N<#E^&'!8&+?Z/@.,68T#8E,4C2GXE%:%><J!!N?W.Q1G;RU+8VPO<NNX&DTZL
P"/U2D1_//\;NUXVGL#-VJE.H@#DE3?.T-TX=0TNH$ML2@2^3Y]Y*GDD"LZ"\358I
PKP4B4^*@8,24'I1;1[9TD"R=5VF_OVS2B3R&0K=)%25T0(,@295IH+,&_./2(5F<
P@F6"QB*Q';;(\:ZZ)G7'!'<26?/@7C-]55($$'9JPSO"![ \VJ[^.\S4Q?+3B1VM
P6)&C1#?H!L()@4ZGG&]Y]LVS6N9.V?B3H)@^XI3E3-V@4RQ)<6Q1GG&'2+#O@Y8T
P40%U<V U)<%#:CI6#C_BP/X0CJ:^[$^=$,N#IBS=5*W6S%,SZ-7<O@7>?5\R4*Z-
P2* 7PTYIXT$98H)Q^,74?"K^@ER+WH+#;">1IR"8Y(X!#T?M)8-7ZD!-WB+W6X#E
PFJ7R# D"7J:?J[*4A$5.SBY*G=BQ#&P$CK@)-S)W>#E?:1/:7ZW@':,-^/ X0F<_
PH>^WO%AY"J[.U=S3AO;5&SQVV^SH+S2AJN-SU987J@<P#P^B"JAL5KRV9H!=Z=(S
PJAX$O1. *3H1T6&!!&=L[V7GM%!C)D?@($XN_/-M;&X;SLA6 M5*]WHC>-897E5N
P/3<[+<T#2R,*Y6M-RB("*DT796B-=?>I8N?[D\B+33N;1YWE=]^H"YY]8[IE_%&"
P9-2EG'J2 EH\14.Y1J0BVCN=AX/[K$2S^:5@)P+/)WZ$T1%'U4:#N]TIRKS/J QH
P>/^U&HQ+?QCF@X!Y5CT'#&\&N(00)VOT"M*JP.2UW.<)M6!(7!3#5.;="$AN_0?S
P2S_3?\E;> [-EY&2HL[?X;=D6^]A!&*A,^<SD-/+3VM"ZVP!0WA64.%MT&+I=8"3
P0"<M?+.S%>QG EF?G$;2FIYL\KWU.$0'AD<\PT=9(+@U]H#_=5^Z*?57?D[]BT<G
P!]5^,''C<QM(/?-7EH7Y__ECL2J]K^B<X48OFM<K**(X3TWE 23G\#3+8KFOQ&Y'
PQ**'6'R6#;MWHY(QL&3<H:CHDD->4GDTXL\%#HN/:!DYT!8OTGT?P)V6%7%Q5#-N
P<PH(_'\+-*9NU9O95!<BXT[A_-DV/^._W.=N4PVYYL*9['0J-OPJ;0=(R_M_02_?
P9#=S0!7;%^=TO,]YO6,N:M][ZDY"X!XPE-R>H*H9ZMM)(9"F[N!R]/@]=E=0 'HO
P_;7K#R>PU<Q+=EJH5\*0"32"W4J7L%L6.&E&/VY&K*'N*(MI+H_.,I6#F'=O+.IY
PX;YGFMS73+V'O>"VZ?*\3\\?ZPNT:/-8X62SMFZR':HMF&.V_K%[.V8LGQ;6)UUV
P:J'4_O/V'6MG%18?0,,0><'"=TN0Z[P?O!;XK S<#&_ -P<K#*Q=7@B-=3LRCNZ+
P-K_U4?F0;?(V%RX_G>_#J?;H*.R7$($(=N_FBUG"(R2KLTZ1?F0?$%PZ%G.H_OU%
P<*F]I @X+X1<M86<]T,^9M>1%+C:RI<T7@.;0K%,;2>T5FVJ&^N!:5O058\Y'<CA
P'EP6GF/BAQ%\LFRD2V7!S%/$LU&;E.)P4^:MS[,H#<)T"W;3%\8[,,\P*$$2N#['
PG.9/*P%#J=?U_Q@I7?P>>7-."?K"F7 [,>MG+CM?5&L%TY8,2(]@VH+G39+;L1T\
PN8CQ#S#PE!]MXC\#"9Q=DK%@8ZA*:L-S9+8P^[MP<(*H^O?75DS-SJ'+%VZ95TXO
P#,&8>($,0S1S2FZ6[ F>QXSG?G6%^H^\LN>X*V7'77%\/L9:.0?YH2WAM#;>J#J&
PL*(M Z\Q2L5W=@*7"O&<:-"QUH*T=I\%C8=AZ;4;FO7@C4R_H.OQR=2V9KCT0<52
P;2<*/>?)2#][JI]#&W6,=IAFC@2RB25MK$A:2?02<*H0X<N5A_:,GP].- RC@$ZG
P]*MPA0_D@K&V<JHNZZ%Y RN'3NG0HOW?RNYEL)RMBI"S=6I:6W[5:!O%W;.&JBS?
PFD5V,R<1@Y^_'X9LF=AJJ,Z2WG#229.W4J1/_C$9@^J"QG!E]N9/07.:)S%*9]-Y
P!8&9,G/IH7!-]#QJ6IJ$1'K]^$Y BH4'S( < #EP@:6%7+=%YQ_?1O)L-NCMW/+W
P,2>J4+8I9#L+Z$08IDC?-7;-4]Q9<Y<!,2.=W*YY^.N@;I5!Z5'CV"P,[B'"<IZ%
P%30/% 'O^?GMW".=@R97L4RSZ+GD+K\Q0":2*IJ'_@5\P&H03["&:G70)QAZJ7#/
PY=6G2?F=F]3QC<4!N\R)!,&)-G>+F-O8_9/BP@:%-C^\[@T!\AIHZ[$TLPQLV@?X
PYRG,\?217/^PS@(7-W9SN-H3Y%5/;80QH'4Z)U@3WR"HJ/'-8$(@3&\NKU9\\B(\
PF1S@W5-3FGU# (9&R5TL7U)5NAW/Z]""3"#NO:E#21?Q@5> @DS[ATCMMM0PVD7&
PV1CP=?BB_@>1\+XKI*R3\^8Z+L&X@5[3:D&3'_" 4A8!4?'$!V004'?9S>=L;R;L
PZ?RI">GG;6R>W$U7B6)".ZM:O+PD$ Y8*4/L=54#>LB/6$2V&:*]?CXH.$I*+I'_
PC18%J&]/$L7$#" O7"@U"P&0^FBEJ[Z0TT U_7Z7,K?27TB5]=PR35"Z2E<P4F.[
PF_H]IN-+S1!]YV MK&9"F"XY1RR1MI\] ERD$5CL),<L*@*U3NER?A^!L1V\3B+)
P9G(5ZQW%G*3! C!4VR4<8V_]WM@PJ\4T'>DJO[;;BCU 2[&1B<T*K D66K^^3T=%
PKN],!VL6_M_BL08JWW4\#/$H>2:B.T+PJ-&/P7&0E; ?N=:.;3P#!N"R?CW+<V##
P_L\&U%8"C)4_AW*=!U/MVOA&YA;J&J9CWMLPKTNA<=IKVW]2O<GWC"SF$4QQD:'/
PB$&"&BF'9V496Y:7QKP\?>&R6J@@/ME)M:HSFC>R\*>JWO5V*=T=U3&RO&-(=XK3
P,1\O.D21QT=%#4);?" "Y\-]['[IZ@E%&@5+AN40<:C6T_RAB^TML >6'?K_KA,D
P_-IFE8K=[P@1+KXX.6\D# @2;_7M?*]PY'Y! ,7=97G5]?P@@)H'JKC05>@CNA$T
PCB_"JCG^Z.T1&WG8/C-2S/Z$*J.U!?5(8!( DX@9ACL36#IKO/TM2>,T2+XP\7J5
P[S*)!)9H<";O ^@',ZLX6KNAPREZS]#^0<2IW=]+O/BJT3>QC:PWG*0GC!N5'(61
PG#A]1?)$:R4POD,F03%< #P:44!?X=X"!F]%VH(=OH+0VNQT,4#12?]14'&@.\B"
P',V,GZ<Q;"9EN-TWXZITU:>;"0H3-O$3L?)JWE*=21.][J=8)^:2NJL+V#K'!:24
PA6%I61;Q\H%YL#-TVI/Y_NW!KG:'N=P: @,O2QH0]O>=2.;BD22AP=>\LK;N=<J=
P.3: MP<#*0=RDK4PR_[!A"TY,YH8YB@WLSVM^^U:NP#G0'ZJW0M!TY:35RK\$1P4
P]"Z]#?3S)\=,//PH-7/ZPXS+:S9.?M):@=_3@+V$+%:L,\;9#R]JR8U/O_19W"*\
P%<C=$)Q0Q)PTD%H=0; >5-ICR"DB^,L?5!6YX /L->I:WS$1:4Y?5T^9>[14Y1_<
P^8+=79GQV7\*GX:9*')?U73^MP;;]EUU<NS".R)?>I*J F_N!P.D1C%_8V_U"_=;
P-57E]:C!JL1A>^G SF<:VQU/?!W0B.SNL')Z\+<,\&10V8$#[(I;6/):O]MXV%QO
P$*[:M?J#U?>5]/;N,-N#G\_)W/*9G,=#>#Q*TG0XYG>":ACY&!W!K2_R;7:G&@T>
P[7NRCV,$UZ:1&*@TWQRS1#NXC#]Z;WRP$Z[B1%JK--;3@-MYYIT7_/U3..HQ.$U-
P^_]4_>60ML+2QMX[H8)Q$= R]$.0*^LRSUNX;924U>KIDRT@V+5?F"ISS7/HDRN4
P%7QIZ"8D D] @XD([;8G=GR0&=<,PN"*D<1UDBSB4FRQH_^#'+B!A KQUYD(Q: )
P@9[L<;X;XG6I*1FWS\&JAR/V\^IUZ,Q%94BMQ3KXJ00/G_WSXUKZ*:T%#FG2QVFT
PZ:>1GR],J9Y,-0,6<=M!(E.._<&[+4'0]N1W=N^G91:O?.<W:O# #L!=7Z<%LX\^
PV5W0BJ &6%MZIO/J+PGJ*3H1&-L*,=T7T\A 6JB,(GE!<4O;VL>"NBWKB*\I[UXO
P42L)@X,6=%;2ZF@QGR?SKS^'-??Y3E'K_*8(IE?J:NVJR+.)S.+H8>>-@ZWJKQ"^
P0.&NV!I/3T]BE25B(<REAP5B,E@1OK9LKG8RC9 +IT!$?67PT%]\)S?F^I"K"JT[
PQE>NRE%,2-%[7>(;".*8UWW7#9C2(!2+3,_0&<Q6"U5PF1A+K2K#E=@,@?JN.(\.
P*/979#/+;-%DD3>A'C!6&I*#!.)[J?VPW;NT9IRBO<W_D4V/<CH]6"VY;<G*$[!:
PZ,+;OL;VX?60@SI*MZ?VR<M&,>O$V7EXI@CL4^4@C:'RYINQ:_:YH.BBN)['A5^>
PV[@9/.97>I]HZ#GU+VJ<1F6)[@!<LXQ%9N<G)))6F[9)\+E#JL/;P@.7\8)52AB#
P)DX0;)=.5(MH@"/'7G5WX&.QD7H#+9V VQD(=VEP+2&H#A]8"B3DKK^/7<(5&]I>
PI*70)Q1%[!X>"]2ND=>,"#)_/'NE&Z@\D\$,77Y2)W$F=[B&!2Q8K5&!?D]B"^$5
P+MH5J[B5Q:D#AH=7PTY-M< A1']9'+P"/Y:;968FW9LJ)E^76[^,VA8WT=/O3_@L
PD?[E]3JVYX[D<=@XB%* PPMFV*[(:TF[A-2UM&LG["-[=]-F@HVGK.7^5>^4]Z=I
PW=MS&"T<?HQ$FF*.BD_J=QV=?#Z0$@G(PMJ>]:0/!,\X,(6T@,A9UJ\^)HKJM#)W
PLS%8]N7^\<X]F_%JQ9XJU$I3O5?Z<K3AVQP48#6@2/:2-KPURW+2G.PP+HU3&U(@
P[TF14'[_I:PS:!5S@^U:[\6 )P';@:#]-,X_<0)E@*RK^Y&_D@#5DZ.\&YV$I**V
P,"MKJF\-_@.Z29MZ3N(93+GP:F;8UK1#-6H7H9@PCBRI(K%=YX^E@6_$5A6P^,7T
P^-@)NDB3P5'28>T8-+,@I-#DHE07#XU#PE])L\@-"R^B0^?@="'ZT-WG[#A!?(8F
P I6+\")[T$Y9"?F7:>_W2TZA_;K.U: "XPKRL,RJF]W3SB%(.0-\A/&8="M'H:@>
P$EJ_MHSR\.LT2U%D8('X8"KE19E?O='.38>(@DADW<;G<(-3HJ6$!H9Y']@8R,)'
P78BRK&%_%9(@&)I0XH*617MD?8>!7Q.*2^]-[MTG#S;=-*!)#?*D\35/\OI[2"X"
P&UC-Y9-^K=K7#J&.&(U']M/4AKCP9/NO-#L#:<J3]&VG^0[NT:H7\K?&CR6H+B'&
P-J4^P$P^>,42&WB>*X8XF=@S0-)HR/>F%-=BQQUJ*K5@&<TP=J-S:-('7H5IM#3(
P$HS+07EKSCLUS:T&K93+"O3/"HO0RJTG?<XN34:!#/D)$WIQ"WW')F?LYE'MFD(:
PE!4$%I$G'AU]"0:U+=C2E@@G@DP<SR@<O(1HS#9=.A?K^&<:+\;.%^S:%<GC%VQ\
P10G]S,VR,SDO_XB/M#'=#J?H@$JJ6P/FF$TQG,*9T9%CQ33D7N/VI_!^^![[LNRX
PI]]M('UGP4MRS'ERS_/<NK$9G$=3RON_6+YB'1_$+P)$'I8/ N4Z&P!2^4$5G6:S
PUK>W2P,[L>C(\$)PEA%W&J[B";><]##Y2W>_/6;?/ ]FH.XIP:#. - ?.Q4IBK8F
PT$6<5JE>94NERU;;93:,GC3XZSK*2Z%",.%,>.1_YE[)(YX*0) T\#<'8>%JWIOA
P*-#9RF>ENP&.HKW$GN:MS!T^K5F7K$NV]6%:N2>I$(QI,5QD8&"Z"",&OJ>ENB$%
PW(CLZ6&#(8!M$+E6/\7[EI;*G(17/IX@?V?_1M&'1?G&^8,<E2>(AM^_W5JL;K;+
P2U#L_ R24*]]V\]./:7K0_.W9,;.Z$N8OZ0_=YHJ'7,D_JYUP02$:Q\74\1KR<E>
P$U<>Q0VZQ;!6=1[LN^5H1<V':D=$66$SMXJ0VU310=&+69+LL?]4U<+9_8N#UK4.
P1H\F;6<LSR\M>I(>WD-\W3F"868XVVA @QZ=$HV!.K5A$):'>TH.W-R,2[J;&"P$
P0#?].:' -,V#V?V^78%R*PX;]);'+QF)#\<\MQ5/D.B37BA<GT);7IS+=8 QJ/%6
P&E=JI'=F*I:O#XWPU#Y0!$;M&,:2W=7&\Z/L(_@B(HE'263Q2>B5FXE_[VZ;PS%C
PA+ !Z6#+5ZNI\RT<MP'X)*WJ$F&WY#<'H'O)6SV4()+)Q>[+IO%VFKG\JKKCIMKD
PJN+^,1S]<"^#H\GVGSN&AA<M</D,.61<&% 4 (SN9JOS4X).@%#*)5A/3X;:CE69
PHT7R-A;]R[/>(B[$69_I BK:+XES3OZ3XYE[28VHE[1)2)-!J9N!^U@KH:^,G;.7
PO)H4\ADT%D5$\,.D@I<?$QX=X-9(>%]X,';,?O=M;?[[JZR2(-9^'FFK@-TT!/6=
PG.#8O!E*63C6&&!*_YOX\Q)GQ\P[4^[4 EX .O-O0QF1\0,<\GF1OAT3]G^K+EG5
P6@[I.BCGR);$UG1EJ@]%5^C"0(Z>F9CT- #P+(=ZN3Q1PFLGB4QJ]80%\&SMUUG5
P+8$28<ZC[+:%L1( ,F)@X74 &=0"VYO'VQX7G&+TR:A9^T21N'YSGM=@[C<3"?!O
P:FY18KD+.'XRG,%"-1_)9NVFR@U5 !*=?TH YU.CR29O1<FRH)L4T^F;HNPZOO&A
PY V,,1<Z%*+" A-M>V%D'TIZFDS9H'3 O_^ZWE:/C[MV7B2;N9Y9L0&]C@ /%)#!
PR9,='ZY5$:9/F883:E,6Q:-T1(4X#\/'2U%U+RTYK#H6@$=4S6OUX31<$[_$P?;I
P+\$@RC?_O/'5BDWNG^V<2"T,2E>3Z,GO@@.']YE*=;@H-B0L@=,/(3?DED!"?TAL
PRR_U4P-O[S\'BT4R9J4CT:$E@F*\+R2R373&?V\,G_ M8Z@H^3Y:#H<YN#[:%N(V
P0Y]27W)HU-&\*V>9,!2+:]#E?\$PU&B*Q9E).=*FN;)%SRP5Z^G"6YV52)GP@@D@
P/>I1=MVKE#2#W&6L-NY6KU8U=X(F$+CO4!5R&>VQJP 3+N&"AX**[>A%?&(Y//7D
PM>]_2OKVT1U6 3>R5ZB8AD8QC(688Z!._YT]5PJ02A)\E $L L9K9D255%Y$WA36
PW!#RU#8&98Q[:<M)3M2QKF)Q=K\ZF5@BK.'T10BS4].I@!/B_+MO\*C:B37^.>%]
PR--#'8F#3@SS1^<JS?)0=QQT44>R#M4P63&,AD@U>74NNU?B;QPFDN1>39*]O$1$
P(&*SBA;RL!-7GW%2/Z]%L@L(B=B],'VQ!>H[G0BK.KB8N]#/<11^VNX=5P#*P=+L
P3GQ>PK23ZG,1!.<42 ]N0G9#G'O%1?AJ6_)AZ&:)/MM'6(0IP\.R7?NQ^/ER$ 0)
P6)L1&J[;.@410N]/7GE-"S@0BF'/ 0T5I3@S!]I,I^@8[4X3+2^(KF0&6.B'B&;S
P8N?P2.* B,?;H#-)6+6.)P((%4.PIC)OJZ7!>Y1"3KZL-<N<K3;")O8D24W>RY58
P$ID^MFK^_8[LO),]UH=5M)5IW6< %X$JQ,";T[XX6J5CDMP!#>4;\+X\XH+B\V?8
P,8$<NRUJ:PXX$X@G? "HC\1<JKNZ:89+9TXAPJ;J4K&*7\-ZX_6(E\U,&Z^\\B=1
PH,"(G-!#WB5]P!4R+'.RA[Y8FU5_&I?G'>R>3@[)U'^:W4L:<9(R^I2Y^7VH3F0:
P8&LLUOVK1><FEX[M6!;RB<["J##"ZX'N1BT<+,GEULUE7CGM<FUJ!=7F"\,9,:P9
P:!%99^?Y[B: !%@T+ZH?W<;&'[WSA$&6&W"C%4X2\IBNY#RB6;7>,;NG?/&7!";0
PRU%,,)5XWUBT"_1"?U,6<IW8B<NK7U-T&[*^HB@\<!(JB(I"A>-!TA.FB!BM]9ZN
P38%MLA[[-_L*&I\G$_:,4AOYL+64J[*V*_W,ZQ%0MQ,U.N?+ HX)!,_SO"0Y?CBK
P8DRHWY5F2)+@\=K'[DQ'WDY!9DAM8\4DY]OB+N'"TZ-5QP40F1XU<,N*1L[CHFFA
PFO<<#YOGW?3G]U6];L9JN7,Z:^\O":UJL10"ME?)EX=Z>-(K!IRU>4Y64!STJ=C*
P+(Q>4,#BJW 8T-6?P=G1RS(P=SO[PLG\ F+E'A;2,$8&UZM$M^SH7_!7GQZZ9E/G
PT EDB&_55/1'>A-<]"\UIK5:6HQQCB2*(L#;)'0$M!*(X,,<! LFBRD+/6/@/4X]
P&9C-TL>;'#&\)LSWW1]0[E[2[D#EO6(#_K(,)#N[.D_AP="&NPT%!,PDOAL-]28Z
P$W%-JZZ@DW)I1AF@-+1VAD8/$$8ZMZQP94&VLWIEA2Q$!BP VB%*LFRQ 7FOMN]6
P7MRX.3LNBD'*9QX'"WV?HNQU'-9?$F+8_I_ +^MCC?FO:WN3%H^=XI'@OR3S"855
P#$]YPBM6N>2 ++H*\M*M>2>)O\Q5>R7H!?4(1+<=5,<#6.>_UN)-E:W?3HKA[J'E
PO-_M2)NE)LIV#0CFSI1P]G\ED9YS97,J10!-]@G50%4A(E_^ED(Z^DD"F\JNI[T@
PVN'7H,4U<WUD+;K%!HF0/=GXWYEBS-J$Y77!E0;+AP\]?$LWX$C.!!R,0'L8RD?%
PQO$A$^"!S)/EG0C'*,UL40,4IX3-W?]_48.5= R$ X+N"LQ56!:5[X(S3@ZFC6H'
P1%NX0^?]2 SX/E+!B\GT7+T8F<@+W)U#>[[^FDRMW\,)0LW^2O.0DIA^MRF9CB"[
P>F1^C/U+(JE&1595=-4A8NBV%[$3N-;:,Y;7E^"G6@B)ZZ\&W:;S5G?+IV&;W.<Y
P#W!Y&=LO3F NB*PV>&2@EM;M(@XE";4_(%W-JE9^96-2%E5U5*J\;F)X)U*ZOHJT
PZE%Z&U%]1;(XSFG>BHI;N9G?H]VA@TZK^U@1*$!L&P;CP %4/1\-\SW"FVV>T^M 
P#Z%]4[8'XKPL V\JL\%6TB,(WE6(NN?YUKH0<C2;O,\P327VPS2C\XA7I;X<U[Q$
P/"#[J=,>.B@<FJTSN<%,K:")O" ^"QZN'Z9O9H[NQKGC=TQQLUY#4/TNW7=NX%W>
PN^2@&5($;IX!&ZTT*?LILGH@J]5H[>R-"96?ZEP?672&I43'ZP+ A,#3@"4M1R>L
PTJ\>W#TTA3)FXMEU+Y:96;2?&>?.%I;J:N1*!92J%%0>4X%T^$H)YZ<7ID%[@02M
P7K9Y*=@1R'\*6,I+8WVY>Z&.W6CGU%F6<PND/PNUX%Q1ES[6Y$;$&#Q=6>[\(0IE
P]04,P1"9TW@YD[892+W9-THPJJ)8L2A9Y0$,?;AS2/%];;L[1$D.V=0BE#B_T,A[
P?8UD:%Y8JF;YZNWAI+9H?>CA-KP\!,UJ MX"&FO.\<8Q_O<9O^?-S3GT%MC$>C^D
P;^>MV%8YV\U/IL?A//;WTEOH!$4^Z-SG@B)_-TF+@0*.4$K.C8#'X:_9'OJYY@"F
P3-.]$>E3$O;S:A>(;92AYS4&KWON=#H8/"'OOPWMK8J V3>'\ H1>\W20A$A>:S5
P8&YO-54 CBX-<78"TWN$>Z/(6G1>L7_E\,Z7ZBYL[Q>Q[]7\'A!OI%T\O50N.H@3
PK#I%V3L)G3@J\\[^%@_X(^F/P!9AV)>)B4<7Z@@*N^'1Y/W]B( 3"PQ^[C:)R69N
PSES"P/"T:2*Y9(LK T?/G1(\DZPM"S8YJD:Q6&VY,W'I1;_WZ/+V%& Z@<("PZB,
P(*B ?)D)LE,^L5U !CJ0JMN2(K1HZ=0F9"RMF5W>WOPPA(1%/@*I.!MNM*F:8?#1
P$+D4AP,,CFZ,%&4:VQ=AE;L$PWNQE<=:S/L*I0XZ^E_2_KQE@?XX#K:^()7:O/89
PW<8@VS"'60P=#NY /ON'V3;T]QOV%.'8\'9 =OE*,4=- +W)5X_0]<W"E.$NCM0O
P1E-M^PM8EMVQ=G"*?TK*5C"S^)-'^Q[>3BN5>:/&H-&8@<+@L_EU+"O%X)4]T4R.
PZW-&Z)_\ZE=@OKL..H2%W_JB>!<K\IL;Z[=@;*=I/0]N5E91MZ.@9Q4BPKOD>HM"
P6C8Q$P\?3[$9JXH8D49>#@32"'RY3W_IF^8F:Y*5.=+N6-U=INI$UJ.2&9N5-K'#
PAP5TM*H\@@)HLGS:BDC/6NLJHTB\"TW^D#EOY<32FS@BN(V1;1A="[21/ *"VHT>
P,C1Q:GO?55SS0A5)4,SO\&=LD=4VA+!OB[[-?'!%:?0Y G6XKH@D9[OTW]?55;<4
P%42AU9_F\S4&HH;$6RRL%DK8ZOR^64;&1J/WX^R:#QQ2MZW3O5>O$T\$RV##SZ85
PX74*+S(P@U>_44^G:%MJ8(@Q^WD<8'N-]+5"Q2>'*1KP'YY 7T:ZX##YD&]JQ">[
P*X/"]\6V B_V1ND)^+KBSX&QC-Q!L1(5^EKX%'4@1.DIE/8^C^[Y4DZ;]9SE7.G]
P 4QHS&:N/)V#H+?@6@N#.V%F;$HZUTIY"&"6)E](NO9?I(9R:NG]IN@F@618AZ<W
P+E<=U4UGV:B-?& ,.9/CA#!#NMMIB1+U\_:<+1W@Q=-*D\D9I#0\!K6'3R5%X:W,
P2A@]E/_18.1D+MFNAPG&F5?'[FWQ-HDM1*;.Y#*@/4FG/\@"2D[!Y:4Y#G-5I]3,
PTZ4M@%/?@[,Y*'+#97;=/$IE4S"'6A88M60G_*!CQ7Z=WAFGN7NR/E7^A'7^/M>D
PZYL0EO8ADUQL_-C7>:T:7@1-0-%Y^8?9[LK7K^DX=31&U:I\"40<Q H36/NR*!)^
PY+1\=,4DG"F9/Q#\LE8QXS[8:-[/;>7;IV9B1$L3(, OV8SHV_#%N5::0[<T_MVZ
P6/3N ->BTTBLPR-C(MA2^6-:V6^R;'787O%M &^#]@(ZM=%?.S1Z?%JTO,["-6P3
P3!PRW0/E\XA4I ZH=T\SG9*"316:/FR%#/AB3!R$!51\IV;AS*.VBDHYK0Z*(I@;
P\ :;]._RPR MB_4 3\<-ZJ)!GE6Y:;N@0+=,EXIS8,+Y1%,AQIW"S'-4"8!R_A=D
PZYOAB.PEPF;6J"B^^ [)91'GK3JX#4JQ,-(48)(VV2L_L]:RQ1],M+3^,F?E6.3&
PPJG\O0[[[]S[[-PQ]D2K-&:7JY9+8BU5(_Q?V< -&EM0EF_V8%M=]4L!T7&9XK%T
P_X3",X^'L<(U^<EYN1%H,\186VX6\C@**&M=F/UFFB__^<%Q(!.J*F<FD6WZ>+8Y
PBD;)]+,!@[H5X7GSH6'DM5[2QH_ ,VM!Z;J[V_5AZO,*:15^35-/(XL7'8%%@3'R
P'/9!S(:.4*YR\6M:KLIQ=B;&KX%2938&X#!]BK-PS*I/G/@HPHS,]J!VJ$2Z^Q]/
P&#],6T&EKAEF;?D->R"K19>Q,/_6]O8O;YOJA&%I$I-+G\$J6GO*ZM&[]3+P<_J2
PYGMS=@C])KTBD\[[%OX8\U&DO<FN#31UY?,?1,AG4;S6"=Y14)V2&.W2RBP#L Z%
P=RX)7ZZ#XQWAG&?N+6)F\JBS2=J6[(H;:WDH[+Z&AP9D878/GY=9;RT&S3@9>X@K
PASWGX 44[7VV*K#E?I#(:J>_\5E9;^^4=6V.8MW)5@F9V(\!;F>(ARQ/\D9M%;T 
PIP95QBVD>$NB[<%,SO')%0.VD<=U*\[(@0 -($U;1*=J:3DW(8(LU X<[XBGN/SV
P.%$:0>5I.69PO/&KQG&V1D#S$=$/_60%]H5_8:8>.!9PQ("YOK@5 5UQ,6TW ZJI
PA3;SS-*BK6!?\I3\PX#EI(&^D]:$!W-M)$!^#G#M1>\26K"A][]3?U^#CBPS4S6I
P3[4"K7#E@#4HML>Z.W.4VV@.U_HH9GGQMI%0?_*A?DCY*<R^)REQ45 B'-8V-8G+
P-MV9WE9&]@-EN"R9U-DJ3$S2$'<^[[1- PY?6\^F^-12X7 _,_:9AD7U:KC9-Z 7
PB"!V!U6->M$2=/PJF]7^H8HCJX'F6S&J$FY!!J/8?GDG'JAPRC;<G!\:7=IF+8[1
P!F2OWM!3;:30-.K,4_W3K,& FZ*QXLHW%J+$$O/-R4/IA, &OL3)JGAOH6^[ (Z;
PAK6BA6NFY>#/-2XH*B^.-^L2NJW?R0$)2C""':FQ9H(,P]=P\'U6VZN5QQ9.?&HP
P:*Z[6D[V$,.*TRS;IP&A$22BL-QC;_?.2CSUP>V!)IM0D3G5M]>"C*.2.\O4_@;K
P\"&9#C_=[-U=:X^W: \SC\!LS?^J"?=,\T:+$7]"AEI)@,#29^WA9M5"\Y_GQ#[:
PR!Y32V7M4B_WC:M([I_/-0&$G5#G?NH6)@S(*8^L(;?U=JOX"Q_DDJ=873QW%?Z]
PF26-F"I6@(-9)\6=%XR)$D67HK.4U&6P.CO#4-27QH')U$\0D>$6Z*%KW^J^9<4L
P"/+9NY=RWIX\_^JH3:V2.61V'XXC<+$<U$M?8J;"@[> K2>#^75?>(HAZ364+L1\
P\++)+5A9!F 8PQ%\ 2N=0]IXN%UQ;K.33F[-<BH/MO:3 *;/PH;!$MPE(,8BQCK!
PNQA4B'<!_)D ;BEM95M=FJJU(Q.S[KC3[?S,6Q=$&W_HM[N2TZ9"_TDG,8V!.L[M
PPAV"UMPW/(*#QBR1*X,[T7O'AM&6?PK_TCM?@2Z8S2X&/"7E1!6;,CX,@QED4@O'
PUC)T'+-:BW5]8%DE^+>)\ZC%1;XC+A^C5QOB^6B.T)&11L$XD7<Z'H+49[+*5CR.
PW5X$C7GI[VM62S)5=*R1&4AO+W6#RS,]B"#RBB[ X&@S,3&, N9H/U@G.?DFZ<S,
PT&L9S!//4369_\W/O0VK4NZ;H[,+=6L3#&53;!J+"7M7/Z'D7=F'AC<N,E%W<Q2^
P:>U]+*[6MZ"UUTQP&8QY?=KXRU)PD3DOAJQ.AI<G$K&';^IG@XR^_ORCGU0//R;S
PF_1LLMHXIB5SMPN;@6.Y'?8C^(9-IUU/+5"IR=R0C9.><+@+B%L9>F'>)P$-<1D%
P:P)1@ZNF)(+T-=(KPTSJJT[/003JJQU7W'DQ4;<L[?O/"4;;>DG7>(]83GCV%DIC
P&&E3'E9C KLLD-:?'_:_RP8>C:R?8101WW0WY?&)E(T8WQCKA:S?(X:B18>HVZTP
P=O^6((3:S'Q\KBF8P_Z2(14M8XEVQ1<3;YJO_JT(B&EQF,: :MC"[4\F K8!D[%F
PDR=%UECM\/B/01(M;0=$TLR^_Y';Q,A/RA"!K=1#<1EW7H\5=.4*'K(1H8K^D6,Z
PZ\QBAVM=367?.*^_!".H@_+(@!B^3JE?<7E-MZW90OX:.MC'SW&*U.%:&QW*]"V,
P@L#BZ>DE2IF)MW@%[95/B+=M9P(V.L'N.+:>!:GX(V])1.26JJ!IT4W"8JG8<2[$
P"X%Z9;@0":9>R979S\LGXY/"WW7C]J&'VU@IK-W@,*4A/Z4&Z6C^]!7$N5G-2N_%
P#^^=B.Y;N#'&6W#RW,HZ#:01UH<4+MIW0)WOFIA/L=_.;E4EX(W2NB,>T4/^:Z -
P#^P+\OK<+17#N?L!0DF>)A<;"6]!;#^<\O8G!.=]YVO*H,#"IC/YL0]UF,A?]]BT
PVTSDTC4%!^JH:D!U*NX.AYT,+]*/8J-F=GGM?T4T#?YK7HC1"X=;1*A11GXT-[S"
P(5D-19_,DMI(QV<8A,F/+B7DQG/M:MCG._'E4</C$P2];DXXY#U*!Q^U$\0MD@5&
P /S11QXL$XL,6 'W;[: !2'7C7MU]5+@/;;EG<K8.2L%0MD7:_<81L]<?A?8"))>
PP5QL^;<N)Q7\G>1VE1Y)/9WU[OQ7*$]3<33E9=$"]1A6HF$%*C&,5<U4MF3^!!GO
PK_VY4^3$T%YF03CV'&>O3UHRK(D)U_QHU*/ ]/CU@<WM62]559Z7L*WWJ^HS$= 8
PXBVR*G^/SHP)UJM!=ON,[$JI:R2K!!L!4I.?>*8GI_!9&H()QIRF:RD/=UF1='YO
PZO,__D*<=<ZSLGW?LCA[NIRBO,"#7)*F,)*GD!GP>RJ2>8Q%D$ 7\C:!6>QK9%9V
P0NDQ*4,+L+2.4 %S^_ZLV76@)"9==#HR<S,Y?H^4MD-1\T_.3F=&@EZC_7+HD,D*
PVITOK2D1J5,]T-/>@/U$G,15P^'UJ*@&A3%D'"CXD'NI171A1GW:BVI>\K'$M[K"
PO9V><YG(\84L^!VH4>%[;%3;OU)*B,7PEBDN-N-3H^/Q:3\B4N?<$\X]?7J"R(%1
P?D>);4/IH;+08UC-Q43@"6>.B0YU*+K:9' +,Y"WE';%"WX69MWI%&_IRKFQESO_
P)NLTN/Y_FAIR_1Z%*:Y7Y.Q&J>E"5*21+;OLP/I3E[RU5R#0385<=C]'J"KB .8@
P(#X.4H< ' X';,>R"UKIOS8+LP#8$[8J?YB66FTRH5PRH\P8>95L,F0,Y[?)UQ:1
P=B9_]I;WZ2V.]W'XS.3T *!GAR_M&&D#K'S+4R#P."T,%;QXUP2@P- W[OTO;/*&
P3)+N_;XMS!=VX%\]7=3H)8"X661Z: 3GLL]IF498-V!U1Y@0:*>.#50*^XY3-XL;
P5!L;2FY0C/0"9=UDCY3O#5797O>9S=964] NG&//*&FT1_9KM#>ZT1D.CN(ZHTU=
PD,<2!W"^W4.X2H;I=32P(:D'>N :F<!?N:[]'@R4_ZX:%W9$VZ)C=',Q:OSE4^$#
P6$U@&(*+Q RG;!#[/5?9WEBT\O>[<R//)2,$J^L*3CV(^DQYN4#^D?0E86SL[:8*
P0.2(";P@'J#OJ2\:X8MML42Y"]1%"[QL_VVN!B5J^4+F@LO^/D1PBXM#*T,]WH.N
P^7.(/RJ(EY@E:,+,WBFN><INRY=4E)R_?#I@+9G&G&$QQ3*YA39M\8=3EE&12ZC4
P62C(N:G^;>QVHD2R?*AI*AJ@N F%RGRIG>N(3)=T@*]CJH5EE$F?);OD1.-RZ]>E
P8@!LS2KH<ODN0))O,4TM0H!H&]/Y5?;M-(!G.NNY(0DJ&[1\:^Q:]\1#[8P=G:'W
P+F04A0NMIQT6LY?JT-0L\'2E6)0Z#GD9O.!/FZ8/<,(D?<K A6?(CH1G=+-U'2-Z
PI8/(>9 ^ZW8%ZY9N5Y&O 1_TJ.&SP(+]H%&5.-72BD P;3S0B*-'UME2$"G_4(&<
PCRU%.>)%H\)80RP_M6#(UO%=F1MU1OQ'YQ,;KX=,>B(5B<\LKS%.'TC[Q_/_CQ;"
PF>TL"4,,](K^1WX7$65/3)&WZ(Z(5T=.9FD=N"#.H-!7V:R)%G3K[LR*XU==LAP 
PKX0]0*O_.X3AV3@9=PHI>M'$<98VA%!(D;..5A0=@Q" (WO(,$*5:):BZ((UA<T/
PM'0_ZWI&4SK=9UHBP=7XY4HDZ4RD0]&9&"3.[J&XR+C=-9@T>"I[LKAE"TK+HHN-
P-I4ZZ>'K;HJ]7#H2E6?NB;)/O/G^LB^@0GRB(3(0K>3?+J,J)7LMC6QQU.>?TP>Y
PV=0;F 8!> )CW'YVB7)E(2G] W9^VGL9OH/L!N@:G05:NK:N$)P#Y'7+JWHXITJ(
P$OE">H;;@K>CO?Y8<VR 2>Q2JUROF1<[D#AC^YH".>>+9$N#=,!G  _LTP6XI;63
PIZV&EX$'&_O8Q?"GY =9D18F<MC:HG2R;G^61?/28<K]J8VE#T S3+][9RQJ$P.]
PYEX)UE9VJ1)&N!0^JW\F*S.DX*952A?2I*NEPH4V21#1'!ROXV+K !_734[L&>13
P3IY>#9XNYB0][+-- HBWT$:\';?G();IUP=:#7VUMW_2A=4GXT+O2,P:^(R:NC_-
P!W(;3*;[7!#6UU?B+_FU,H+:/]%,]QQ'N;(KO^-%)\HNK:3$QG'U$ZXK63#G^:;)
PJ7X)12_(X-_!F^Q1V JT6S^M94JVO%0;\0VZ]-P-2/=KGL53MH9TD-Q6[C5RK(AT
PBRAFR1):9#3D_AV5.UR":# .3ALM07+.R(XKK%!W/ZYW<1:NFQZ. ,&?V6AT9.QK
P>>*)G[EMVJ/CD/2PDDJ\E;TE ]>P4:00\4GGP!STWPG41$<IF O-\"S(_\Q9.Z)6
PPKB,GE@>+?/EL.W6QXS8-'+K@*%<UK],()];!$Q\9J7*G994[/+@6S#4A9TRHT=>
P97X3'<^WIG3WQ0UEQ]#Y 1;LX';C&8CT.CNNYI]V7TN'?[Q/1'ZA 82A9F;E!;^D
P9#:A^@EG- '*&FYU7[2XUSN38WEX+ZM7=*.1))YY2^E"N,S[%J1RC\H=HF>#67-&
P_1]]##%]=FG9F:8/65*(VO'>XH<^5(L&)='=.1?HCP^&O3DPD>O&P8%W;IUX<@"I
PQ)_DT3@8X=_?B<5ARC,OG;D\XG1V'22VG1O;0N&.>:)!7=.D6:F3#J_R>&&;\N8K
PPV,(VMO+"0R2)8N0DA#LCCNJJLZEEEXGJON]%3&9P '0!X"RB?.E,>$=8X)5TK,3
P68FCR %6E>_"6%VO6?Q671HR1"35]@V:=6)UI-R8.+&QDW2'DS>;Y4>VNI,'I)Z 
P.YU@KT1%8_1<>^&X-%7 2]OYK5UZX\9$X$JO^MOF\YR"%NMP>MZIF:<V,(^[+KUR
P0TU&S=V\7;-%)^A!G>@$^FV%:_\V7$;7FL$8GTYA:5.M\S!?F_P4PG[%0 #;!M<&
PS(1?MK8A;F8A?O]H4;8M2SX)+)_)J]DPB&</V*0N4O$Z4-POL2QJ* T3)-N]#X6.
P]BN3QE>VX@H]+;)7G:YNGY-0/Q\F?VSXK_[KW7670.5"N$GS.J5 -XP38S3$4B?I
P3L!<CU])!4W,76YEQIG-6NA&JUOX"=G<A\T3:1:_,3DT'ZBBZ?G7\L?E38J_D=;5
PV2;D='HVIU40)GK,>NB !+?(&\K-\(2X*%__&?7S2B2'IPU3XMS@\2#'OVF54[)6
P%(81W'#P:Y0?Z_\:A\2B\%:BQ$G\0#Z(C+AT>PN_K ^:FN!F=-=SI0IU8U!9'IS,
P?>,W,_H&>*)R4H[[4Z^T5"Y6F )^?O&!JR-YB0?;;_TGEQD:60X:"4W"0UM&P8@<
PT>5'Q/@(W$5_T^AACU'Z2+/BF6:K5N7\K0+NY/!O<B=Z2GBZ>3\#@(G]%%Y0%NR=
P+"P&H?40[A=8]DE  I](!5 L H8=[H:J;G V8#"(E5Y$F+N)#GGEO;:U&UMFSO'N
P-=36=*6((PP7G/3#* @_0>.P6%)M.\R;*9WM(+ D:[_'.G=8<CH<6/B _&36V%X:
PY^B/16^%(A.B+]-O<JVTS2"4_=_]1*95.7VK@#]F-OU *9@'';4B7A6J&-J@A=4L
PWUO A?\OA[H);?V5'1) F+PGL,:4.233O%U##/"QJ(\^*1)\77HM?2T^UHJQ/P2P
PH)61DZ]S+C ,G,>I1T$86-F"(JSF)FPK%1%F.&-CLXRD#"T:FRV[U'U3+, JS I3
PRIL3B^M-<H%:T.IZ9V4>(/EP]V>:\;4KY8LKYM[3T UNP>#PIB3A'YJ/#ZYR7117
PH[B[467?'?QQP-><LPNTK+>,H7-B::U4=98C=75-*>QM9=7,0=LL@+0:3N<76H]M
P4.JY$3<EFEJ#?_ALH'RN;4 X#K0J*#&LN7O/V->PL!30=PS 2 A] KQ)_,R@3AOM
P2D6Z06JA3FR 9@J,HM_-TK[31KLT")6\[Q?4,WTDYYCQS7S?Y5=)[B@OE8W"J"!W
PUXIL(I,.V7[::N-W^,\$((Z3CNN%-.1E"'_55R@R7VLY^15P]P\ T10GXC ]@(Q>
PHUJQ-R/9A;>5Q"C=M+CH*):A Q@*P";\S=7\%_OX_=HESC>*VEK-TB>FU59'8FF6
P18,MR7WIMJT2 V4UYIZ0<?!R<\2ZW'XQYN+89_!TC**- JR_)M29J&HOHF-MLRM(
PARTYP.\F/[">"T8<Q$D8NWG ,&^I-"!)ZV%:WT)ZSHZ/"'];2".]?-[E.CX>97B6
P6<59O5E<*WDDP\[]MGR! ;MY#+L/-Q:]U\0A%.46- '<EX1_\91M,4A)\7O[K?2$
P47K^95#<!G?@XU1;+-?-,[:9-_M@N!%;*J\X6\(0(%-RT2\L*BPE%6E:A":RU\Z\
PT7T0KRVFP6GJ!\L6%.F#=58,#:&5)(RT3E$]DT,I,#196=@NW98=ZG>"U59QXCK^
PHS&JE#O1 Y033"ZGP:,E[<GJOMP*.)GKMMP[]Z'!B1Z'<^VZ4*5<1X(8W5DYYI+9
P5]G S.0P'8]23*J9;WI ,E/?>L" CEI>61Z*O-=1><5R0MHK]]UO2M0<G'^1H<EX
P-,KYC.?JWC=2P*I0]Y[V,A*O>'BT#W<=EW-.F=;QY_7CGQ92"L=#BU,F-$7IX^JS
PM4?!I_SO@TU(&\F0(_RORG4]?4.MCXNB01%(%_@_1?*3<>N%:$'E*A[8Y-CNH(U:
P/&F5F*2=R'@[WPL25'M,4L;%5B/OQB_]&08KK=>=:^WYOENO0)1X?2L/^SK:)Z:V
P04!!,1<C[R5SOA<FU[=JQCD-[N1N\2D>L+[/-G0X5KA@RI,&%['E[ UFPM_G*+B#
PX$Y8MNJ76U%P]MW#YM[7OW]#6_Q*F?+)F&$/"880BG!099D(QV'[-QB"%,N=3KHP
P*L9R>[T$K*FUE9D?A/UJ^?^L;L/?*Y3M'#_\(&!^Q0OM*_JD;"'(FK[$9]0.3EA-
PJ9$#?:Y!$U#1'_RRO-"_5_?K7V61$Q(91:S+OM^TGBK$ZH<&*!#%-S4NK;TY+H%%
P(D4]Z\-GPW_M^H2I%2*@Y811\U=[KA>QS64]4WH%#%'-#SY2=(8Z!T9-6DMVMY-Y
P59H$]:\]=6W[-HX3!A9^5,^IVR,,DDEY>2GX]-0*[H'^7Y:56MNC/*"D-'<NUWFM
PKU/XD5?A3B9\2E37%LRND6^2A-U10 F<46DJUX;+S)9/#_-!GAV!J4ME6R(?__:!
P7X_XJ=,D!=,916T3[B7N8<IH<?%+5TD,LY2$!\A&BYVJ"'\1>B''[4<HDQZOJ,Q7
P]%*.F'D]?>O[J OIG#:@Y+*]YTX_VA,>Y2A9P\/4^?<?_(*8W+9]Z\?.5F8I?_Q;
P#RXRZ;<ZUFBYG>KICS/:] K>=!XT5_:Y#'H^SVH3E)V13;2>5E 8@N>50#N\J G$
PF+E.^/(;-6"(]UE%<8DG-@3.V#]HY=/<7%OJ\R;JG47!4GM#_LZD!W=Z!I:&U6@G
P'N>D6-QH/@<%L>6P>Z\GYE[!_'Z@>6S_I&JV92+&RB*0-S*(<7#;]T_'LU^=DD"<
P4J2A(]9%LN6FI_>,S-H;D?NVOP8C1<CGH#2H%446$T#LV;?VFL8ZD_S691L#2"=6
P;T/743+2BK0.W>:SC@QPWGT+'N.!1U>;Z0Q@N6IP:XX<-I/. @XM^JT3X%+O]M@/
P]SJJIK5PC.^]%V_@^4'*CD CWVPM84G3L3AOM9%BT96E*V0=5LE6X.A,3YJ<)5 G
P8(4V@*[=>@7@F&C8VABT!1K9#+#G;3V$PG;98;D/N8<92,JO=Y0. V#O\*,IO@X-
P?'S_D6CV;A6*C1A8WG</WG;[H@F=Z>'U&J]'-P@SD]<+._U$^STFEN?VG^4%3:A#
PW<(7N2&,[\4 !W$*924HE+G]''H_H@#&<XBA6@0-?5YH6=7J3,Z9KVA_0&E9:@>J
PX36-7UG8.G)7O0"UJ%ZU;A#98,E4ZW""F=OZ-#6G)-D<';1M?\PP*T\H<UEE*&+T
P]FK Y=I;.*F'(9LEW>G*Q7X++-*9;>OYR:',RT4T',BQ#I]O(DJW^ _2.!YTZNU-
PT$'QWPF#Y\EOOVI,=8.M*]>\_+\=OAVV <M16Y%/#VU GZ,&57L&D'+!I^QM'6#I
P3WK- 3:<4'S6E4G>ES^-AE6"8$O*EV9A*6V\Q8/=U9VLGECIB<LO\7L<2(F,R-3V
P$L@6]4@'6D8_-W?BPCU]9=:TGC:5[/<F@&E/A8U:#B&"[P8#;K'SE<4HI1.<1>GM
PIE8+UB:K;&OVW.534@7Q?&_P_4/A)?,-W8BXIB2T"BD:$NPF$*JUUWL;5".:J+AK
P*3H<5[[=VB!:\O.O^K;?5$X(.%5&B$"0L)TM/>;VJ?K,R8(H>.]6P$02ORA942.]
P%>8QJ*MM=?O'M$ Y]4X\#0 9#WF:I-V]#"P!BL8^)OOJQZX]4; A9]$68I+<=4 4
PEI0FS 8FMG+QGN"ZDAD)S5QYU9#H#1>"%L# Q0G(SR<46;@^=UH5"I+:SW0"W0^9
P*.6$<XK]+TN]3]S?"S@2+MX@KR-UW%V@(2"FQ9ZS["$P^<Z5?CHHTXJ%+D*;';-F
PE.,>[D5?E6LMP;'_WK^PGXO([R,_Y"#,?<(.9XF<!<J,-^^VC M6M@K,0&:2-6 "
PVS:ZM[SX0=568IANSXJ6X2:NW#ZPXE&YFM'8^3<CS+# PZ5K7::_R8QIYZ(*+#\D
PI^-.KRFDLX]YYK +-)9^!+H(S!<]&I$B$K/--)G/D.E*(Z".%1A/."^DCE,"!!6H
PIR^"N=&<E7@5QR9N"7,;7M'R@[X%F1L*!T_;I_)S]:0\T\+C>^-"L](:FCN,?126
PW*"<<.K!T:Z?G#1=#YX#K>XX61H+G1MV59V8BJFOUA6*EBXE#MOY5K>W2G2.R4N\
P%Q"M\TTGZDU1'MCP9;:24M7>!:82%+\P#0_@3E]W=<$-SLT1H? 43QRV-L_GR0=3
PET<,E!<NOFTX257/MH.#!T(J',Z6K<_QA;B,$\E[MQ,:Y61<F-18VEVY204N]20O
P%'._ BDN<9/+&=RH8SJF/)CCFP ED&WW[4 _'ZI H+W_$7S=JI^BW+97SC:2Y [5
P/L6DQ$,-P.;VE_'Y%&H]//'OEL40$$'SD_V&DO; 0OFU2"'G L9ANTUQL*MKWW:N
P.6M)I+K+ :?JP ]1$;)'9$H>DO!\4P:?YIB;X] U5GZ=I-.)/7'IX <)@Z%7696U
PHM'DQ)NN<VY5O3:\VX>&MWZ'?Q<&F^,RX\SO3&:21_OF93QQ,X&#.XIZ+I5^@+NF
PPJN]B1RFFUF,T&BY4>P]82)\A?3O()!EG&T^9J,Y"]!E"> =I]GLU<WM%_R \B)D
P(A (GE6R;M'K7K2_/.GMK&O+D6?VW; N31N4(^]MW!'C;M!(Z#QBTPO<B[G2O^T%
P,B@%=I>.<KN-0PD!.G".RP,X'8T?_7V#-IIS.K::UM(L]8^Y/R3;(>)82K6;^((\
PV8>D$JF_=CF'IJE *O+2U^BNQ/0$K.O!%\Q=D%,FPMJ+.$C'*[1J=5YMWAN[C6:/
PX3F_%0!QDBA%8')+>NI^L63O<VO8*J[BN 5*OC)_IV:0K5W<PTQ^7Z.]KNAK+CN9
P$P"Z1#H0$8IE*JP= O/:W^>?GIR.GO^_1A,MD*I93_41-M CPUV/NX:KX_50E"9/
P^=Z'(D'WEJ&:2>LN.J];!75S@5:RR%W+*]?%^\4XK]$VQ8? _+/72P9V[<#;,P$I
P*57,G]D< &:'++^' +GTN_%#6QK'.FO^(W"W8&)>=Y<FKT?3:@TO=NA0K\A92NCL
PRYG&@] ;8CGOQ^+$%E:X1>M>RHGK<D#_69GBX3QDPU]K 6XTO5-.6B7M)X=&7 LX
P/0^B^6(VRE R,E_JEB\:8"$#,_9H(UU_*V6Y@\U_=/'>4ENH8;L %=#%GY (!"M[
P&68#6X'6UK7"@[>EJ')\!/=[_5 <<A EGB)V4W,!M]B$JTJ7-2,*%S4?(^'8E5ZP
P\LMO_4,5/Q((L4,[!]O,?(NT!.XK9':\+( YVR0RU/RK#A&5SC62TB<^84F-BFSY
P@Y-2-IDL-%]N35,"WC@D%EJMG/G+I[^OBQE4WK\U>S*X=(S;9T JL_)R<I1(T].K
P_Z]\N<7'7*HN 1<?S,TZZ1/*J8TI9U^$B?A^+ST<^:>!Z[(QIF&('>7Z253FS2HV
PQC&.R_S3E.&P.Q:)8W1HE9WW'J1UER=NDHC:<DXER^WD4^;/[BIN+1M8A]J#/5N5
P D,0&:QM"4];]_.SJ/:S8W&?4)'2[,E*4CQ&^X>O2ZWUD)ESI)TSMA2Y>^_[@(^L
PRDZ!YD)=.-SJ!7OKL)]F& /H;;X:,#8_)W;P108J^.\ S55AZ!2!'W$G/L%7QI\5
P-L!WY0(P<6XSD/2M;;BK[7D],++?M@MP9[>U=PMAD90&->XG)7>=6.-7B8B^+T^.
PWK]6EHI]H?+\DWYM?3+U\(9+9$!$,#5-4Q5M"5J0QY^963?<VCL"9J>0L&Z&LSDA
PX-/O<::9MI:@.83:&=B7SZMJ*:\<J@_(L4.P@I%J9%W\#]IW#VA%>9\ 3O.\G<:A
P_1R1"32>HBQ1_Q'B@(1E2OOO\G+UOB77.N"LGABF:K '6<RD=QB<N'%.46L>39@U
P%>Q>@ZT^!S!'O!PKEQ=?[D5L)HFAP\XJPF_3,S4=\^SG1$_Y&[B#O9E#0FQ'N#B7
PZWQU:?@=*.(CNP^P85N]V,DQI5K=%RLPUJ-T3 OL9!%CEP0IY&GI,7UXF9'91O#7
P,SOKY.RP,))V"7*IT35 EE(%2B#5TF%?QDFUX<I<ER)R%<,F%BXJ;ESLE'5NV/KQ
P(Z_D:.%2P+IELU=4G= 5,%<2($IJ3UBC8H\>U ?W%PFR\Q_HR1!HWM'(WG?(-#B)
PGPXX;_@8X.M]DJ%%U%&Y:Q,SFQ-(@U4T,<[,U4%.\=[E&?.Q%0:+O)D13.FT')"^
PM%%UR"PR#9RO?CXQ-F8U&5,*/00_E;RX'H;JA2U$<ZZZDD#RHV&&HG=^<<NP;B)K
P4:^#=GZTN&6#4#>%?0<W:@:IVKF'_167U U$#OD*8"W&O7"?%'.IX]X+B)1:1G!'
P:== W@SHE1FK#TXE!'9H\CT2$Y-^^5FJ./. (G,HIB^SQK8-I@)S*=)!/^C5LDXT
P<[]OX1Q/!2UF9W&3Q[X?^%GBCYU:2)SX;Y<ZU\$FG071CO<K+)A<]:I/*[S1"\H"
PYT]>&83+N4H+_%"$(*"#"))>S6.%5X5;P?EH(-H'1O@>6[UJ(&+<D5L71I2UZ/A4
PQW6L)([M@'(=#/^966IZH2+\Z>[)[\NV?V-?3UD.IF_8#Y71#Q&5-T_Y@*@ QXUV
P])QG"1-O\H._:#BP:C)M%)U4D&X&Q2.N.'% ]I(/%:6(8+H>TV.;!9ND7.0XL7_:
PON\=-L1QL)V&'A3T4H-_^02G;(Q;SH6C!/2B=1<43M[IP79H1XTY/F,C 2V1_Z88
PDGV$P!*TSP@6HSTXSRC2__5!@)<0U#B'K\(N'!X($7,-]^[L:+9]Q[5TI13DXN0.
P'K;TST0\Z0S,Q:J'5GPM"%$<R6WMCT2*#<;]+$HL'&LL90A%ORF9I(($)SJ_8 4Y
P7;#^O!<"KTX?$4(Y>#:/_53#3]7]]%,\009/$OQ^-=QZQ??X)].W7?ZE3NIT+[;N
PEVEG-^679YAR;+7]_9N^W.,N7932ZUM($RI(7#BY/J>LU"O[Z?5)EV8S*NC^Z%-W
P\0&!L7E92E32H;G\)[?;AFXL*J4>S5@FH0?EP .SQ3 [1OU3+ M:U.L=;O;+H)O)
P]]#[3G Y^*]&9.JMS)+F,EBH:6.JB35L^GW+2Z($\]%1C.EO(A8/G/FB9*6TO.J6
P\+G(COYR8_I)RF.26(YF/>I0B]3 MU>"4]:>IGT?!O];5*#=;>0LS\Y*4>*%9D);
PXIL77,&50--)).=)GZ[D=ON[>S_G.3A-S2="03.N.Y,H'/J%ZK(\^8'HW/2.8^0*
P6\6QE UU2YEY@\D_I%5@T&,>Y7,J",NI8=]FM7W<=D'9V[Y ZIO61$*A7EFXUGL3
PUE\;*/!>0;%>?+,C+JBH!7I (?P%T$1^@/C.VFY;<2-L$V[',"FUN<>'M(@IX!KE
P6;D +^*PXT1D6AG$)YD7GN=60@<:_GBW;DB1 DJVIH;Q0"LTF&QFBM'.B/EK('^.
P\JG5/!P971WH'5((8Q#2M)7)KB;'3M6U6 A_<3%J*K\L4Z=>:=,. &=!E_Z@LX%8
P_7Z[3ZAOW./ PVJ=]A!RM3G?^KK,- (3>1'L!SD ""0M/I,$6N!7_I!XQ*G\4TZ>
P+PUVFS$C8"$>YU"SNKLDMEPMYX9XOM@ZPE:@ 4F.E0!V12A9D-V3P%/@]S *L]_[
P 8#,R:BI"J,5+V3)V'K>='_%AN (ZGWPY#<9120.[??:9\:O]Z'^8#($*_I:?#N0
PLC "$U/.A=O#G<=%#8%H<W7HM)LD:>OD+TJB)R?4V,QFV0Y55Q\-NSA$V]*H1YSM
P.!PMA!JSL@.WF(61BL==5JW9PCU1.XRNCS#!2HWSUEL(VFWD1ST9'?*YBGVR 9XW
P7^*[ ?0K3J[X!:H]V?Z=?],;IEWY 4**AV;BME;E)3RK0VFKW0\?6:KFX 6AJ H/
P0Y#O&(AY".H_G^R=2X_2ZRQZV. XJ],:9X>:4O1+*Y%PL_"I)PXQ/J^G6M]6#;VC
P/"A1&(?##K];P5'J"7_K4:UB?*^#%X?.&+=N4W2W$(BW-% OB[+"&A.G\(1(3=]Z
P/'J+2E;4@<PLSTK>?$^@%2RPL_ZEK/M @7R9::5]:@3.JHK/K=CB67^TI0WW\[?U
PD[]D6ICW;6G:\_P;WLDV+8HO]H8]$#$@<<]NLR&J*1$%Z&?ZWD?]"CO]8E>-EQ,%
P((3G)10,]6:I?7O8C(&1CLU,3&EP<$RP,Z/,L;DS;&E-\>+ A0_.<^2I)N2* '(A
PO-:@XE[8 F1;,_?#IT4!@8!7V?U7XF>9JS'\@K+NA'RSQW3TI_7<?=4$$W9JSMLS
P&A[&V$:.[+]Q[8#]2$G6ZP:59Y*G1F1D&VJ=+]./]#Q(LLCT6L98%\:V:UI"6(WZ
PJ0/$J)=*%9/VB;3C2?LYE)=0YG0E'*9+/M&74%/&;KX1C$43ON0UU5**_S]>YYM,
P@M6"\UIA-I1V?-L\>_^S3A#WY1 GI8_%50%D2;%.D(7R^ B56CT1<4]FA^?9]M[4
P9GBCMOE-\K2]L7G)$,._;.8T=:<Q+V9QI?_=#L;VTHYANE1Z0"99]!L\71&K&>&;
P%G :@<5%K8"9!"T7 #:5@)#-$'2!+(*4%,$\3; IR#I_61=@==<":@F:TO?*T'\D
PC6NAW(U^B!)N\<T5L&WD[]$E7C ,EN=-5C':UK+-2ZN,P[_VV!ZQ&)UN\MB?O@(-
PA5+*_'-*KFA=%N<NT)S8E/Q/!0[B?&MQH>[CR(ODM\X6)?SOE9Q'BT8V2SJ0># 7
PZ0*MN&+]*372=)[ZF16LGV%1;WU.PD>S<H90$(@,J@WEYP=I3A4I@X9UL?ISOPE8
P"J/G1?;@0#(FE(?O7',8K)C4M\S-OO._I\/G76M4(.8,!"N" O1274>AO@%?(#%4
PLSLL&722CI*<Y<^-;N\!$H>J:#(*^[F'<7. OJ]OO_97R"J 1NBK)@IQ9'8Z&&3R
P%K^>5;U$* Z6!@*.)M(3NGD;FR$8XG@JZ^.UAY"$KO\AV+#&']?$/D>JO#N( =;#
P=G9[,D$'GGC%9VHDT// TKX@&G(@7,FL2-5$(3ND!&,13^/8WM<?M/= NIP;!K[N
P+'.<X67@EIYE\*/F/\@ R5&;99,2S  GK"*C#R^VH&RC.5JF,("RK"ST,-<(K#]U
PA"U3@SV2-J!YT*O%U2@%=VH*%2%=K?[-[$N5,@^[68:X2U4(EJ@Z/J 7+F^N>GP+
PN%W9JLIQ@Q5RB-W2*N*<+?PP65$S6.J^=R,\/\D3KHT/R*D-YK]Y4)+J6XLW+CS\
P7D 0D_?B702AN9*Z6>CQ??V'-$IZ29<5!?F@Z2%@]7NATROG4;S/8-14Y5\4XSXW
P?B5Q:IULW\PRI.R4G7!K?+&B/D*@%CI%;]#B3/BOJA3M 3X1=E P5GNF>$MHZ=[N
PCY><T37=="^0+%B-%WL+8KM1X-%0-J 5/O!6,EG*TB76G'4Y8%ZISHO)YM4Q/H"\
PR3EG](?P</?J)J?_C%/3R9<7RA:PR:UH0=)Z\#H-P,[Y268KM*T10Z?P+$?HEI!+
P>W4HQFG_7_STKP -NG;-(8/,)B9.9B#J1TB]2TV=:;T-8$[F+(-F.H=@IT!M(+F#
P=0CP!/%>#')(4"P'"*[NA'+&-[-I^O:=*%!1Z(3QTD$D-.0Z-#-,_Z'08:XH<C/+
P6'U5_&X Y?N]TYVX"GY,T!++;#$F3.V^ F7;=T.(F&[')OB$KPP;V9#*O2(D1&R=
P[XE+:;LK>?SN8KUG+5[30HA2?A%K[P!6X4:.AS[<LE9]4?C^P(4_?M56B<'8;WQ3
P[5[_ 509IZ[FCF X/CEM-;CZMAG:&:M!#GZMSP$'Q,*(KEU^L=M)#P$N9-]-\,!V
P15Y1RY>_].?+4:34YR@3&4HWLETFTD?$]X0.:T=ZKHLEK5/*K$WI/R39\XDKB*@=
P)TKA!Y-$A^.,V'>4A2:@E'?L"678(S5@DJ&7(XS 8/;.G&CJ=;^O&()VR@'].TL 
P W__&1XGET?JU=$]4X.FA[&U!_MM()!48SE:!BZD+!(:G)!\5%8"-=3.D0Z56D37
PQI&(K _P[\F5]U9DXS(C6\((3([2\%KZ[;6+M&$,8Q]LXQ+5[$U?](_E[YB&H@2W
P:#WS-]*3.5BT8WBT1V\O!^:@?>6C9@=.3JYOXE])O  "F=S.5YQ:#3!#=8DQU/42
P4XN%K8(SW?7X[TOC C,'FYK>/]=2I@;D?P\QH  ;D_L$ P!N]"MYC:*!*:M_K(95
PIM\>U\7YL\6[@7O3'3CZP"/N!9,:!K_2XRRA/9KMM)#1XA77W?<A8P%U!.W=EQ*@
PW4)I:(- DI,X-0WWEH+V5PDK+L!F_#,K7,?4 8S5^QFU?Z2 ?/TD2-/=!W<@T\VW
PN(ZNX%36M3H'E@<0+RK[P/YWX?T#O*:3!/4-:[[MC["P"&A2P"#XY^&EKP%-CWCQ
P/E&C)]0. NDDS5<'Z;2EO66EYV1E ;_-(2>]D6_-W=C[;^QH(P.2C^C\0UPF6_(:
P,#K'9 JBX3P/H;TS5XIZ4:!G?8\"R=_%$S/X4+)2!.65]Z8D=]K( 5?-\W%R-WXA
PS2N#1L$)@WO7'QSE:Y'4RT!*E)L)3"SE%4_4NB]31;9V0$ 3@T'$WP2W'RJBM3M9
PJSFR,LY;V']N>,YZVZD^]P&RPP>C[)#A1_MRYX9AP")VG#S[7RP BSKN)029W$XL
P)P0">HOP6"8B,!I];^@7-*FN FK,\^[]<3Z_-0O[T86X=%Y,,2NT$(&7]IZV9J?B
P*^_*Q^&R:UNSH/XPDFXOO*1-%0GX :>],[1$TX'O&R=BI<,U,^.\9K3 :A0,[N!^
P2P$C_+!MQL^-N=5KM2G9([AQCL@JY0>/,668*J&)>5JEC7&6,Z1B18&>LR0?XO+I
PR#L_?2XVB X#S,7\P>%D?""(=*;2U]=>.?G_,4UQ5?[C#M5M=&9K]*R\+)PQ8<D5
P.EH< FYG-ED57%V^<*FA(G&8:2W,&]:'=6+-:L'00GYNG]E88[[95K+-,+9JA_]J
P169>$DR"/+/8<1'S+V6Q>@BFLU!E6;',=E$?3G0D<&L"6VOAHH ;]TX9MW/S&?9"
P.8U>__: .Y)T8@+$+<Q$L *CV,&V#Q";%;^MA=@N4A;*1YW%)9N%]*I_\8''N@5R
P\K6(7[\F:[TPJ^!G7Z[&-YK!_[<&Q'5/U>Q=-$_8^&QM%;9"^[-+1SRTKC[ Z8,)
PEG6WQP^^4>O+%?LR&\3P4&X,OU]1N0-L@D8UAPH_I]H:11Z.02-\CC=>K%0%"CRL
PA[_7;%P?W01%>SD2R$#D/N[4**N0U)#?-N!67X 08#6TH[&\=+$A"[_EVA=^;3*^
P S\_7VEXX&E]FO_=C':4N_]6?"B03;41\CQT407TFE9B9F2' >DX_CAZ9;+JR"H1
P24\7YX='@(.VB_R>0."F"K5((8T?NDW77P>ZT274F%5XI0++LX0?^..<C6,* ]?%
P\V JMC9V<I+EJ[]_)C 89T'#X077T,EZ-IDN,!5VD\N(XVY+-]A)=,I[131%W RZ
P*3P3H)(QE*=6 O@S  _;RAN2(PIF[U:!3 @W3*@.O$3V#Y!W0N<LC&,1+JN9V+?I
P;8EE;HC#!J1WR4P@+F^)$JZHF9+-PXJ^G.I!TSX@MY>5B%7MAVDN;NED:$#BV'; 
PWZ!%\27*H]*N? VD5*WJS/XUX\]EZ3QCNLD&$/AE@\2N2U)UM2M7N5<-L5W_MU\=
P_U8*=X]S>/IB<.]F0*O_Z[[3&/?BY]NQATEAHV7$57 8J3(P&T*[X!.9FRJ),,\?
P/77J/DL\!;!*SY"P,?UG\!0,HD9S>KP4QCZN:<9.2!9'@4OZV#6HC<P _/>RHSL^
PTBGHQ/<4L XH)?TJ<+;$+PFUDVS2RD6I >5UQ0R$2PZ-9O!] TTQ##WZDX)YTQKN
P1(0#F(G?0)%^<AB/8B23%TV>ZO_N?DL[WG?N8G^7]"Z526]+VQ+(.YD^\- GD]UN
PN&)X=\8^*G8VL2<CKZT_#RXQL<@I>4CK/\5RG8O7QSMB,G/*4(5M'.CWY2P"M2*_
P<!%T?@%*=(<^^C,EEFQ7_X]:ERE^WYZ:/ZVS\#V/U.&NWX'2VN#?F?AY"J][J[#'
PV=GZ)3%IP#1;QFW+:V:Y-BVE:S@5?@">Z59.K':<D+87Q3AH0R_+ON=L_5'#Y+QM
PU7"SZZF-I+O_4/KC^2QO59,E34=+'+P276J=."DC'XR(?%XDMS+-7;6C,61^1_'#
P_\X+QJ+Z0S84IF-L%01D[SDM3CKF70Y9_$DH,IW5*)DF&JLPM?5!' <;=T[,@TN)
P.X"H^A!VBZK\,'O;@%";N< 2'&D[45\</T=MWD53<5:J@&@"OL.2-+!<.@TO\RQB
PU(UCQ-!TGD;9?/U_1<04(^E.P2)_SZ?!>V4LBX8'="12\<!P:L*4;Q2Z1U9 HIPD
P19)AMGE4"$NNH=;FX\:XB<$IM*Z/8C-WTRO0YSJ5GYF66J&A%CZ$2F4Z(!#2.?NQ
PW2#(TW>EIQ4BSR>V1'B1T98+\WU>NUI)RPK?6]:;)GOU\+X/8/UW[#[DK4*VT<&R
PH#/%R]GA4;4_V1),]"D)?ZX#59"CD166V$?[%J+7??SH5#BV'X4(&Q$9*"+AF9FJ
P>P CIJFV?<!#JKC]7]G7*8@O/[G9&X_9$^G>Y1: >C]RGP-$ BW%<@_90DZB6X#3
P?^2ZOA^U5Q6L]Z-"C@G0\YO3?R1)[S@L)C\PD9$D8B3*Z<;7;WM[_XA1<TUKZ<<\
P,E?*X^JM!S_BTK3[1(+E=D!H;XV]=8WJ%Y6.Y3$X%@AAG6"@J$!H'AG%2 YPP@D 
P2C:T N?F]03[XB'I=2&KBI'$\T9+F*54?.%,NA*4/LI6+VO(E-WN['OU8.9L>&9/
PT*V5MU</22&=E_F4U!<O@.!PRG??T2-VF;#8QS;A'--/>A'I#%6GAS9E<M0%ZJE6
PR+K:2%&;G#"+1]*J)*&%<)CTYVAX=>/DMI/!BA46=@MY@H84\]:\3E><[\"$6_VN
P+:DGRMZ]5W/E%>QNI^^9>[RE*%N6YH4X!<PB='K:WBS4NZ0HTL](#6VIQ8AU:0VA
PJT8-]('6$*K%JPY<Z!T1-H6Z ;[@ --=[BY8MJQJE=_ #!=B(PM^]I[\,5-GV19(
PE$X8X_P_&))M_,I8RH;ZJJ&7RKT@T[B>91(%T:!Q:HO/5Z3GLOBSP]\G^#&0!FZ3
P>8-G:PSUWFS>8* #08OM@E*H7.*R7"0D<,,(KZ;+FY^]8J8 :V&G//N8A0*4%,J>
PR7T<Q9*!C3">!*;&%L9[QH:,K9*HQEKDD'@R9$._* U4 X<*M6#R61PPW  85>!L
P@((J.J)F)'$?W)_Z8N?LF5,#:>L[-C8:F.\49X4.N.!OA)AWB59,/:5]*$('=M0%
PZD%=P(5NBC'-,*V+':\,A6K3UF>8/U7Y,U1IT=YN,<I-+0,+*^:.V15ED#,.P=3X
P""C;AL^GU@:!;' K._7AH=74,C$9/[)+\O F1DD>T 5]X!@=[>E/"1\4.:IIU0^5
P+4#!@CYWA2#%[8G^=+XK#$?(@]!F1,$8"N&?IK/HD$1Y^9[$5'<X1-(9F7=^Q<RF
P44NNO['$JJVRWT))Q'2N"PM+([P;Z.N\QL,OL#4T(OI*!@<\X1W=RTC@ %8TQ-AF
P:-(4F*I3>,8/G.[Q>"Q;UK=2\]-U5J:&HVCRX"G+(*WQ).S/]]G 6>["BYLFUQ.,
P'492;G+7F6+['6E(4QC9%A.G:9I=I'[5=G6$"\]-941I)SGL\\W-AL;:NEB9"6Q0
P4SH5]A7KT<703::_Y+SIO?9!'!]OYL0)>V'\0M+04ITTVS^(!4&>A<05?EYY(HPR
PZ0RA*H'C+JL8@?^WD^!TV&XI=06^#L[W0FAI+R"<JC^CC;!,T[$(!F5@VR%; $IW
P%E?A9;P"[_PB/N-)G%_6:=6CN$D'BBP!\%26.!QH*>6.!+F.T4'\1*FV.).335 I
P%C;X:TOQ+:,'-FH'N;@U$S2T']DY@3IK*#7)2FWMAC3NB)0:![P$38UJ7#6G4#!#
P*+FGHA-&Y9+5\J:#&$V:!PF"7JY,K\@I8>V2@4&(Y4 B=6E,L#=:JO*.1]38^NML
P'#U0,MI=QSV+N5T[R'\ !!1CIWRRX&PCH^_CISUO!N:R1/OA2W;&Z3DS%41:]G'2
P[_+?35<X.+"8UF+5IW9,M,AP29#O0:-0KF=_5;ER>UB^0S6&"FS8(ZD6;Q!V[$%&
P74]B3D8V+=]CSK+E.A$_JI(.2$;?O1*#%VSTC&^,X%U"V>W]SP],Z$ /?C,!7W)0
P#D%F#([4O1O;71-:+K/6<F", 0F0OFXLCV2U"1R#O9$F\:F(B=?'LH2]- !BH75:
P9/6SMKB](@QNWBZ;L0+9;>PV(O(Z(%PD(@'[Y46!+9L<Q3TBOIX/K(%7JGL231R"
PG0I!O68,(X=:-/3I,W[E#SN^:O+7,8G/198S/@=\%(5&U W K/\#)=*LM$S\>HOY
P.^!^3 *@7^%'("(FN 8(: .,G\?K05^V7M^SPOYX0D^!M2LFLU]+DG^M7-0ZJYQ>
PF)Y+Y0"?H%#@Q/%=$SZ5^9[SI-:I!6WRDWZ*(-UB6  G%R"/VCM=C5G)'O# 960A
PM#TN-H4 IJ^6C?_.[#'9_ E6(F@Y[-O'0&5+.GJ/T#69!!ANM!ABZ:<AD*%U[8(5
P4_*PP*&5CKUQI*7*;6Y,LF^#+S3<_GI*I:)LE&>=*ZJ%7"R9?]H*6$[-*.%'JOQ/
PTK]8.<;&-@-4W4J>4!X@U<)NI&!,!\-N,/W)#GHAPZSCQ2NMIL=XCGQ/.VJE^T&'
PG6.DZSF(?4 DDBC\=)I382_+M+).DEYB(X/_E04(Q)"6MK[T<X @G0?:YS7_<#MR
PZ?P_6*390Q><R RM^;^A*[KBR%]A)GT#VU(*!C]UD=H7>S!7S!*DBHKIS?0$]W F
P+Q0DUXO 8FI\]$=;1(B6@M9!/"7S/?-GAB3<EW1N[Q$5@9= D;91HY&>SY-1)A,$
P'<D=A0:(+"_.(W4:0 4W;ZU4G(#;AAKK 02]5"3#D@E+@W>KT5;UXT[2LR07[R#3
PFY3O=0TZAXE][#GI<-ARQ7TN=FE^PRJR#;])Y5)ZQNRH%G*7AS1HBI/NLL&,CJX6
PK(\@@^R!!L="\[7H_!;0.H$ X@IAA1;Q,>VVBWAHYELH##9S??,^\;9/+)1SR/+*
P-U<H7OF&"A+-Q_8GT6,/*( 1YLI>1]6LKS]VB6*Z:%Y59S>/>H"%2*PEDY8Q"3JS
PW*CF=!4D^/W#6B%5*M*5:_;9(J+F36J?S-+L_[38[&R8((@6\>_]L/V:P#*2WZE3
P<36'1G2*+J7_T3I9\+%:-WWJ8_2JR:,Z7_"J]D)5J()>9.B[[7)TI&6\0V''=O)F
PMA_27V@&U)?6<M[XAQV-5Q-:'TBTGU>O%(+'J2*]?O[5H=C!O\/2YWY"WCECQ\E%
PX-L3)-*(4I-=X<1CN=G.RP@%IM?F+%W_TS?WS]8WQ'/LHGO3Q-.>89'P[++D\*K^
PN-I0F+:HSP' Q[B*E1=[GP08C2K5+*)%Z,9PN@_J(_PE=Y7GL85W[Y]2")+RLP%-
P4;59PLTR@.D:Z3ER'"_[5+*++Z_?UPH?$-]WF;B#G!RC/>[Z$^PP[;3+FVKD ;)]
P,GC7I5$QGZB,<V"1"/Z>32,#S,E^[!8O[T8-ZZG+GZ)8"1*TN/VD%.#L)O6UMF'V
PQ=0*AY<2T:<LPQ\3T.Z'\B FUM#48Q-JDCV@'E(USQK['A DKX'^HD:3?M@<IC.V
PD"O:43GV_RB=.^I;JU$$ZV.N"X$>1_9RQ$&-TD\$/M*S<5:LY+[<AY&A-\2U)1@S
P(-[R-4_JB*8I:OCA;(!DP%,S)2W<T*%!+IO0IS/6@U;-_#[CM@HX!C%C;6ZNI!"'
PW5K@S[D]!.0JH^<0)8MJXZ!\1GK9]E=2?2%>J=]M=3(O7IQ\L2906)F.(2!R28PP
P@=8/%S:!18>GEFW=#$6L7^[;+B^]<K)T@A^P\IJ481HPP:>KTXX.)0(9MUB*5%&@
PIG\\R(?H$R5Y@2,W!%?A72>:L48WNLO?GH4?6&6^4QT:PB5ZAC<5'"\0HATG-ZV'
PXN]136L5#-$!P+BWQEFZV9@V>RF&69\'@^T7S<<"SBYGO!"=(:[X$!J,O<S59:;R
P_@NZ-[$A']O"_-LNEI&2CJ?&6QM7T(T^KP5J Y,+=?]2PD^4EKE<I/@&@@#I^?9W
PM;;^ ;PM:H7;<&\+\K1RKMQ'/TW"*,M&&-YL"VUQCE")AD)(^906N8C#G>;SZ(<R
PQ_YKCR0C@,YE6O/ NN0$*M^2GSZL$9]KE /[B=OXBGWQ/ZMC(QF\$S75AS46V1S@
PP/BQ3I<#9:BLL(6IW2( 5F.2,ZN)[H>\"+@(3]R0G^2D[I:-EC=#2N;J_(^QJ0:0
P7EM!-F>#^/ND3D2(X(=+F/'&?116&;F/9<;ED,+Y1P1XO;_R:W'/:?O E;4(?G$Q
P%L9[1*N0'\&S#^AGPR#>=.'S["N^D$VCK":R3ZC:KKO*I;57_.N<D_41"LIS8)HL
P8 "Q7=B0OAO_MTDYE(_#F*9$*R.Q4#;1U>&U.0WN+W,V%RF(B8#W;OB<G9 4&U6\
PZ-I9+X5 3:)?F_KL52[KH(>[:TE+'3VKP-/:Y+)60=L;T0:8\>&,EE7B<"R/$C]&
P4,RP$Y=C**%J; ,! A $P[PPI&03<-T%I@S!A&U0NJ@\6B6K^$K5JA(IA>D!;NM9
PI]+A()O<[H':V &A*]AL8#O;^$O]K*T,W+(4?'1Q@.^>NA/FHE*0^RA.,XGO"Z\(
P>@BXOP%+<#EM,2>!O@PJ'50T!UL+RMVS&4;>-G]U).P'7B-7T,5KUV&,,\@D*)ZO
PJX;ZYE77[?@#+R..03>"*1!!>U$-(RW>"N!AR%+=<P2/N<#KP9E+<,?ND.941#@A
PES!L4PJ^Q]8Z8G&?23L%_I#44U*X17?3FQ9T2B"K?*1:><O&2ZYNYH8?IE(HR &\
PY$:U!%=1!DYI%])HF-^E#P-/N<1E8,'<*CUDC]5%7:Y+)<4US*P9+^QW&37+;FA<
PA!6G=U9%8D!&<A)Y=-75A ]C=@+8T%&#@@+Z;"#9IXT)"_AV@QU61!=Q_/W2+6+'
P<">M#0E@5D%IZP*J>DO1Y*5/+1/:>H=<;(WI:4N9[2) Z%(;?\3,,]WN0IV@0 H2
PT+9BE.(.)M[^!$WS,L)W=FDOGDQWIQ+HU:A3=RYK4-%2I-[))V0,$'ZVVRPR1*4E
P RA7@"9@SPWZ-%[UO3ALH9B[UR6<R%\RD$("9&91\%<'\(XE3L-_0)"XU:W*%.2U
P(JP(Y,2PUA$N3+O7"L$DZ+5K.J!#-5RI$?S2OLW=PV$*PMX>$P;$?;N/X*W8@G"W
PQK0S4)]YS"/X/"IT_<);ATXJR6U,P:=\G<;T<N[!^=VMQM YQ#;HR$]OX:G'#.CW
P@I0+O4=(LP^SEM?%YXJKG+Y3"Y/X#LK F'IDLCNXR5T3;;7ZL 9(/& OQ0'(Q"$S
P[IO]6O#XJ I O7DXDL'P] 9U;679V.R@J=P:TFTR.,BK8+NTKHA9W>+D_XL6(H5,
P9IG-VKO%O@&N3W$N:K-[Y($D*NK+A$<%FOEJNK/M;)\.2,QP"AK#QO2G:B15[\QN
P P\*4.975[.D%]/8NY*M@%J_S@<?ZM=(&N$@^JA1LZCA=A501JB:H_#VX@S7UZ ^
P:<O>%IP NBA(! =S\'-)G]GRD!.LG_MX9K5DP1)-W+TT$L,&4&B5'7+4#1RCZVL+
P0A_35R&EF_+].]+Z88^@G6D%):7,5S;62./5S9N>D)'[(\$W/M"\KR7R\L'SI*37
PZ%S/X#LC#/F,GG37MX 4=8>^Z/]NTC\:K!HK_?,:.M)$QBY0)!##?CGNVCC*3Y#C
P0\@SG4<" E+@\C@_C;/ 4YI$V&)RX8?&OM>I=_CX*=(7>&%K74&31Z8R(\%ZI80"
PW:9#@$ @>' KW<7D:9 $=[43U\X1GC&%K55GA#$$CM\AOZMX=6D#MARPBOR.[_0A
PB,DQ[E_2B(4QHI?/=^DI@GC0F]PV"5)QV[0P)!GWGEZV+T%B@6&[+&]*XRE>\8TD
P)(*+&'WN>PU )B@0T,Z? 4S7O?&JW\);T?9,!SQG=CQZM;L:98?-T*FKSZ R:"")
PX"!H?5'EZ<Z8B\_I[#(J9GR^*,>O'Z_Z\1C\&BKPU L0'TTE>28O4[Q2J:Y][:-:
P9A/-"M!=5EVNAN"K<"Z>&DR.KA;"A=S:\MN0"#B-T+G$5W45XHBO.H/+M=Z4V%YF
P;U7J9I0F_N798H#V1Y"W<5@6WYB]7,?[!G$.,:UC8?"ZDM1GPK?Z("1/S0?KU;Q3
PE3BT,+Q>K:LRAO'2U !PV!X9G(,WV$%Y#[S,-TY!J*EEB3+9&9"% U/R:(L:!/?9
PX<Y8WT;)6-CN\[@%]!$ ?&ZC<_A'Z%;V6J[A8YBU8%T?_O/[*=^/("5X.7(FW_(W
P3#0;H/B$3J0S=[],[Z'L!/NT.1?S:YF2ZE0GY\CH1D;2,)QF%41P9 !K]!TOFR9 
P)P-QW,$^)*H4&$5]8>L9,R"]ZH_9>08_QG'&>%<.F%^FRVLLF$V^$A,'>(] PV8[
P'A-0>;XT=Q4$_EUU(<4BC_:,<GZ*UI=&(>"?N=7K8 U$@HC=^BX"N'V6LF,DW._C
P1Z62\I9^,8--4^!I%(%%%@,V!-]EML3ESW0R>^Z0/9-*DX4?7]D2W6K+D&'(:Q1V
P^2V&\\H6'NWWICTR!@V%K8AO_E1/ \JI@7=#+D& Y^H\'XC; #Q,)W5O3*#F^6S 
P"I%AW716(,J@ DNQGG-(4Y5D9*AL%F,9/*(1B'W]PF;@*L$P&N6FO?3@&\=(4YK;
P>UNJSDO;[65DE@0 ?C2,57+EROK>]IW?]B6P:6K$$'/42-&MEA";2/\1_ZKQ:?3*
P_^4>S$/H8?;;-$/OPR#_+8-+?QT.:8J>2HP_(_9EU%6!I'O%?9G6T]7#!\:$S8;"
P1<XWB'.T2TA$HSA[$Z%]++SQ4NL-^'K2D>W[?J EE./]6R7,^XPJD/VMZY-R8T_S
PBT+]61AD=]#V;HH*(V:8<7J0(J*\]WIBV4A#NW]/-O96@SJ/=)O)N4[(@GV(\C%(
P3;0"(('-9N)'V@38\1$$4A_D90U!8M 2MYL%%<X G8*J >H,$VCKR,,LFG[3Y7[E
PYM4>@X&=\KF@\/6UG"1X\V45'0=_27E.B<6M"QK,*U!HD59YRP"LB=6HIC.U!K,V
P8*>O9F;W6QSPB^WP6?["4^&A*;E)PCLXER.@%>2 N.$/9>6XJ5-?.:_WAHMYA$A+
P^)\X S\!-9.3)GZOI9^UD)OX5W[@%I9QI9"P#]Z6 >B*],"9Y%S\PE=]S49*-VS'
PNBC[Z/Q*):S:<ZK\'Y;9>+KA&Y96KA=]U1[]19MDR0G$'2#*35E>DN"'.1!@8AGP
P._D Z ^K_H%\<$IR^PEG&&+P7<$!(?Q:PIH<0NP@>,@Z<DM!S4"+185\$/U!!HPR
P_RX3,94HGCIZES"'L3!CDGQ,K&DDF4L)&X5P3_"B<,KMQSG&4L;S\P%L=U;_T/K!
PD:'#UP"165Y\2/NT?4FBHHE9O%/N(<W3N30]V<@\$8;1G"E$O=4+$<<"%PE&_"W,
P^H,$**9F:!H?42G9W- 3171!SBCJ6%2YQ) 5T^'ZU%OD]P$?5H4DL;LIVG$5AICY
PO39!:,;P-S4'K_ !_R3ZL_"]%>WM;_>@2':F:/C^3G\3@^#SC-@:O']T;(:L0QSH
PI)(VI2M'J/A#Y2\FDUQL.?$$$'A8X-+3A@0XD\J_F7KD4N;IM5EZAI@&3/991I&7
P0WE2*JX,$W9PT"YB90QZI@C".-W0-6U\N(@2T'^H=?FC[H]M19ICI@[I P Z%U#[
PA1G^IW"[T21AM?V7\6T/LT->\5GLW#%,?^ZZ/W_!?AW4CG,)._<!B&);$(R+5-OE
POR!W,CT*^3W >@T,-&UYH0]XN0UW XHU4]:UGB$1!F>']M4(\=@'E(&9IU?K0#L,
P$BHI?K2/3OJ2RV*TNGBHM,[S/0KAWW844IRDZ<H6D27#)S@)7H,ARQ_]<R5(J=]T
PBEL%>$;UY\@O$[AKQ B],DQ84DW#LHS3>RQ1'#M %TB'&Q"#/VNKO!YK3D4/CX"D
P U;Y\7C68!PJK6O9CI C7K4!PN78"8"E:%J2-%Z>?[!9MD,M:94AO$UWXS>;E5<2
P(J88D6):\H$ .SD7!?WGPS=HGGQD\MJ)SH*9EUO_Z6_04-8&V8;/[ L 8IZ,18]V
PB_\#SI#+T)KL^S]QJ::8G$&T'G 1TK4)OB0\ST.7FM,P>9V2/&^+J!84X'!E4KFV
PL/\/ Z[C49CHJB$[TUUJ3S^/\=5XM#]2EV65;V%'/3.A63ZG5JQ!':PNV <N(I5N
P$7X=K>0:ZSB2Q0)7=)YL/0'K7\]WUZ'%B!V("IPST)\RG>1S<=[F]PTJ"\EP=5E3
PTYIJ[1GO=0WK([-$ ["</P:Q$ !%IX $DPAO"Y#4%DE090I\K]YM%Y!Z*R.=HJHK
PO1/:EK_#_Y]!P(K3]F'$5,*";,:YB_%PG].5M/>I+8V3>O-!TW$-Q42I4S+@+_BO
P"F;F2-3L4,CS[3,QX]L]QIV+#YZQ6IK>XN@X-53MN/8@-GK@>E_>^(%-JHJ"+ZM5
PQL*0F+IC8E'N$^Y#I]:G]+ #!:'']R!TZ-&1:_LL6@GX?421%Z4; S5G#:G5O<BX
PYLQ(CL].B8(DHVQ=PS#[%M&I;H=!>3/ZU=)=QQO*!(YJ!?GX%P&ND##(=\>P[ L'
PRQ**X3/'F T%D$,SFS_4RLFIT@#VKU!;4@53'GPI),Y@W/Y#*+ZW]%5HV'=G<S5?
P=[&QF1Z>@3W =*@T8&3X-:D/Y>5]1PXUJEE8R6S>&?[4=7+I(K\('QUR+?Z#+$X3
P")AZPKB<VJ;PM*?+#.5C2@I\JZ&1/193E7*]3)A;)R3%+RK4$K&9R_UK:NN=BW;^
P@$X\G6PXOLJ'3Q,"(Y"2<T)Y>& O-C^8U]<EXY<5N >T0T^+S38H2%O?C_,7./ W
PU,NY&L_VKB 'H3X=#\LU@0/KK&@U_ALH ]'RV2!3<U .Q55.X:_K;%Y-4_683TZ%
PM=:)_N\31=!/+VN@$07?[:(IAEG@'*=X*U"[PB_+-OF=!:9"&:^Z]' /H*EELMZ,
PQK^X&(3K>$IEC>RA6'9^2X$$4N+)WG@@]XW2Q_QTR/:\M&^Y>F>U\UE&8[J=L=WW
P- UKUEM9T*5OFL_Y:&RE6!S'8.6F-=[4%*/]4FQN=KK>2MX+@V93,(EI8!;-TU5$
P[?-N,:EAT!Z,AV<?J*,)GT%8Q2Q63J(I;_AG9=26?D8966QEFCBO*_*N7J5-WM8L
PR^K.=Q@9J(_SYRJ.1,4AX)ZG>7R>E!*Q76A+MEIQ=Z09M>EEW3-B@)28*^FR)NHX
PA^'&?XP;M*50PK+0C\^FA:'!KEI7+UI&KDOHZLKS<^W"@17[C/#O5?U?7-3K E5^
P<]=;6VMW"@65,L*&P BY*NKW^)0)8V2XTFJOBDG1#D;YY=L&48'!LV/$%M8/HH+(
P._<**,D(3+")BB,8,I.B"3#A\T@/=?1$<LX]3(]:-IW"M_(3@ ^K[B2YV7W+"D!D
P62?X$A5!WK! @+K&2\(DKV9B+ \(MJ\/94I""Y>ZU-N/$B] XZ3%?&G:SA;(SGBM
PS[+:"I5!0OB^']5IMD5[*!IX9*ZA;VQ.0HRLDW2)A0=S64O_,!SKTA1'M(0FPLF:
P5BQL)%F(;M \7CD^T.9FNL69)YYX(_@3.2,]'$3B?TO;E"$_D_Y*R7IS%_[]0*?8
PJ::63U04Q?3FKB)U+Q*FN0=(L"%J5W%Z.9$'0:VLGP-AUB?E?3W$?]&<MH@'"S2R
PTOMAX1QX)FU'Q34J2<@7C+>6PNX]<66%I<@<24^0F>-UD\+U?^M=\6Z"U>>01I'[
P<F0X(I^7P" !:F:?TYP=0!8-7 _?WN",-1)&[*N<[-^)+I$IJ#-F2L1?^,A%-CK0
P[JSCG11H^YYW0*F--;L0Q;Z@]G$H:?.Y_@6XB'NK_(FAED?,8*SEX0]XC@++I?\E
P((K;KA-[B>*AQ5:<'@T3SK,QQNU;XYR/T3WP_<(]J!PC*AJPP3((R3HZ]!TWL$4"
PKO+.?&S%86K5APWXB0<AL=#MY/&\R2QWBDQO CC((<SF3#UJDP<OWXX]C/-IV71(
PD@]@E19?6.W,H$9WM:I/;E4<XW1G.?=:*=_E/],7_K!^<TWCA5+/T,"]U&_>P()0
PIS6L-']<EO ^PI5&BG81(C:Q&0SGL3J+B#I?LJAQDXR302BBKL"RWW>>DR$V9">@
P@H4AH&A6^>/VE#EGY^D6?!%IT_.#UCM7=-CY.E#O4I'FK.S!8I83^ Z410D;:)1F
P'C(BO98]TW)SS9Q!!M?5QP^"/66:6Y[VR/=#P%([*"D\<WU"Y0MC4?C5,J"BH4M>
PHH_J++!(D<':@ZNR7*HVGL9_O Q<"*\UJJB>@N#W=T?M$:OY2/MWI[H#\G^7M.(W
P+9:523BCV^/YK]7^NV_"VJ;TTU"38OZ,5'&"3X-Z=,4F+<4O?:W:N?91JT$2>!/V
P=()\M#^?_7.H9?LD8X%OOD1QA=5'NAQ3<E2/-U5* !WK(35(W^*(4Z37_,0B4Q1]
PL'_>SW;^M5(<>PL#M=)8&%W?OC<&=\E)_P04BBC_X1.*?LQSQ'S#=KB9@B^I?"Y,
P_G4=DN[P>3J*<4HA3ZQTG,N41YL6O!I47 ARG&DSW=##TM3_]'O1+?$HRX;Y5H3A
P2Q&C0V7XM+,K/B^#NR35OBUOXOPMF:$X*N'V#M1B_UGT5UKEY3.>O.B#^XHET.!-
PM.XF8^ER<DQ2_3''U-*7%K)>!G+;K5,=9GM)_A##.7H/)C4_;O->,HY"9Y7HEA<K
P$ 4^P+.LRVOU1?B*H(M#:*P,C0Q.N.-_)W* Y$(SYKM7\^TKS@'K[U\1ZW?**3&S
P$+4[^E2X#R;VTE':<9:.OA)A%!#P-"40^3-N@J0"#KGGG$,%LL;F"LBR^AGW6)UC
P)\*&I^P$?8H/N4NH=6[G-X=_X0)B8OVCS:U4?LHR()ISGK7CP4N#FY#3?^XSWX41
P_%9)_L\VF^,F -^ UQ2F9*0$H35^^M5K@4: +8/4\=#<01D6+K&%5BJ;5+?EK3 @
P<-%OCU#P^T',$ZJZ6U+1=-+N3-8?$6",&E?P*H,Z4XX39[,>B(%][-6K7,2M@76P
PE&YM!H/H);<27K @7I3MN0>2?@]^,CT^P#SH7V([IO8(2HHYY1GI[#"1-386J3*E
PGT^II'6$W.\$G2''%'P^2)6B>CXD90^-A'Q*QX>*QZ2R)\8^GVEY$#\^AUS#&M_W
PHV3/TK%AWNXXX;]X]6H1>R:X7FX16!RQV4V<(@]-8Y/0M&-W[5)[;%N]P)Y:%*K.
P+,"/L]. AJ.9V&TQV;?JAO(#UPCF'V4?E]15)%'%1LEM<;0:-9OBM;E]H\#K7&?6
PHA4P2YYP) 2SMG+/GD,*21S3OM<RB=Q#DRR)I[TEY/Q>,.UCH$G??CK=A[ ;8;=8
P,YJ\A4"V.=G&)^VS7$@D?R]<3FR6TZA%HBLM>^LFZP<'7?H<K47=^^!4/GDX;8F]
P#$!,+5S[=O1A#INVW^5J9M4RDK*%T<P7OAC/YZQRLF<HV8J2R*_S;X.TU4S.JW[3
PGPO NIR4D\=F1PHEYXAAV__T!#<WJ3%;'%^MHGT!>!17 G9".<R6\2$PLX[$  6=
P3YMK/ZLM-\"C7+?X.)<#'%K/G[+^$'=SUP.)8R,DNAWU&<H55=@+@O-M!)L))..1
P$)B\VIB@X80C#.KY-_Z,*XMG@K.\?,):,\Z$5N;)Z,QL04GY$+K1$),XG99,,+6?
P\<-@K?A&JVAFR<K7!S1WG5"+!OZ/Y#P/Q8? B:E6E@6>\ H!O_>)6I2]VEN!J>=C
P%^"[VWIMD#+(A5XM^X3)<0Y;L?A7Y#_H@*6H%J#P44A1U> 3>[M7 @6\'!7]4;SH
PT9'(GHZ0'V^C*F>A&/'.&BB["^Q(\^+=C^\_)+.8$AICV;F  Q3BI<"#.\?KF N8
PS*^[11Q#,!%+;Q5L8[743U;)%Q>;@N:T6M].;FD7PE5L8<*/[,VJ#'M._4<ES'X6
PG%0ALJGVE>4KP.1] /H5/$^P\TOC#$-G?#9*?EQ$XL3_T;X6-_\8")B("H&:_BT_
PI=R&!S)R;*3&V;25<D=JRFL/#$UMCR:T-(P)&Q I4UA&WNL1TW1_'61UTO6^QT%!
P=%CM)1.Y$3'<]E34M63T!NG5 7!8\DPG(MVHFYV1FU1S.NG*ATW2@T:E"#.WVTR3
PV?P"+6=474 N!%P9$"# 0B0()-;.LC !V/YE16HY+_\^GO/I&R)1[ON)^8J1+I74
PM(=[JZP_)IQ=K]9V%8+$6:4P+:)KTKD@Z)Z[8DS@7N:AWS__^S";9)Q03K;-4);9
P'KU:@4EB@S'GU;LG"E%-_NQ1P,0AV0.18/;R+;RNE#\!@$!M*&4'RB<E.?:5923N
PU[R_6.1BHJ.]X9=[L.9.=.SC??$S$4&$#AZS^IT>GWL?PSH.SJ>QP#FD&;5 Z_S/
PG'#Q?SQ^EJ29MUPW/\.D"G]$4A>7Y$3-\1>3*3HC@AMK]M0+=HO7#!+:Q8 HV2@:
PTKB3%.!R;O_7-RH.B Z,S(PT]-/W!]Q1N1-"+)U*V,W^MO:VWT7'P9F5B +5%-=D
PRPT\7LB_X*H'/6#ATK'3+F1-X_[ L;1YT"N3&WH_X"O.L'U;SD+$! =9$:9)J'Q*
P>>8$$9<.;,7POZW+]H@Z2/&U>.G2,-4<E9,7>PX2*YGQSQ8]F$;J8/@N*%/@Q(4.
P2\I$:'X6_O+W=>G %1$=%4T&!9'\RJA QX:]G Q69KQ) ;[H?=QL6AT,^Y/ ,TP\
P!+G?SW+4_9T##="0II>$MG:H!'(;A<I68%$<. 3/LV8?UU3!;^Q0/+_%;7A71&%1
P-[$GN:Z:$+7Y8_0\?:'-3PT+A]]#<1YJ/HG?GQ85N>8YKTG. SN*GZ1WL$P? K@A
PD]U# ^4KHEK](13:E49PQ\CN!$UEK)KEU%:]&0AK5 &"L,'KF5LD.O1FEM$#22U^
P-YL=QHDN86YH0UFT.O=7@*ARL.D5":^BE[6(4&(S.+RR&75=T"79M:0Z5?*_!XOD
PD=$Z8"(%6*+B7\-&-W[H:S E\!'OK.<#U3K$XOYQ.^Y.>C;6;9]JYBY%Q@T_+SS@
PGP&"H;QX47DABA*,1\28QU;?07!>TE6<6X-I= ?).80BU79Q=N@"BEW .D62%8-W
PK[9?\U?:92E&']M[7)RF#ML/7I5!G%BMN=V!/[O>KI:4O[9[3T;^7LY'\DGSP%8S
P'_220VK3G2TO8]]Q/4572G.Q4A++K)NK,"&\1I?I%U#YP4=ZG3]D^,C*28U"#COA
P$8QY#E6@G;Z57?%!;KNMI4GD"-:'7W8)[M]R,%=F(''!\/_@0KR?D9QLS25VWQ;F
P" ],IRB@?Q!#@BO*G*C$ZX3@5&S"_H7=Y4M'0M]]-U"YHKJ8(%'V14?,EI3V^NZM
P:^])J$<[P/V/2?X+4E[_%L$VU(9OTYRX\4-(K522:#""QR(24[@Q39U+0?=CFL)^
P^[.BZ%E31ME2^GQ/K&D>>L[4J&C]"QI4HW?G5' H7*VN_JV7.F_\;G@HPM5#F:U3
P&F:125E)8B:)^B*:(1F>AL&"M9\;DN#2P[^UMIUF:BKL-+U!<5M->[\RLS-1$%W0
PP0UV.,=C?LF6'-9J81,OHH=> /ME#'#_GKOLOH+:R.'D>/OY'XN":T#\['W'!%LA
P")R[R%&3N[(.Q2'WO<1:IDO'MHK88]E%2$57W&RQ9+X/= ?#(L05;&DQ@I:Y[!!N
P\:Y45E-4>_V5/C)<!3MJT]I9H+!DY3B.Z<?E:B"$Y0BTDHA,(V5=#1OHUZV"7/N^
PM^>6?);%X.4EC!(SOA8NWZLA3,::%BTY$D%@+7:RUP)M_!UG4K[-*I!VH..@X2.M
P]%B/C@W]EV/UUTQ <<O40(P$JYMO(BY@B:,>'Q&'<J)(6)\[HE0*T4Z#=WDA.N"_
P%,YA%;X?%VN4$K/V,!X?__COW@L5Z9==_4?>OL0PCTTH]J9$C)'V_REE+R4&Y+_K
PX2?Q4ZFDVR%3B!Y77X'%ZJZZ\:K>2DPGDB'DWBFWM918BW+GVN4G\G'?ATP6.E,Q
PF/U PLJ!YEJ*=0*%.[G7B^=)Q?:A(18MSW@VE'HNE$_6$I%.<;(=ZIZ=S0&H>FH<
P?@@%-7;G6>%$PYH9#'Y,8ICC?-CC@3Y'\WD4'8A6CT7KGV"#ZP)'M<6K$+)^U'[G
PIM-P'']:K3!U(S L.Y8&5=HX"GJUPGGSWL=2!#!258PV4;KK)!0* 32'G.L*8T6"
POD]:??R:>I K^=O"_"7WY]QVR3NT(58OAR'IQ<^OB_T%)GA:[E4S$1:NM@1]PZ6J
P%NL,>C73R?)1J=X@;1>XZR)1$52TNZE#TGZI:D6A[!C9J];8)^,,X$Q6!VF:AIG@
P+P^W0%',:ZN.J.U-ZVN(LV>4YDNS$,,XA* P!&1=-MJJL[=9FH^;@O/.(EG"*-6Z
PIB^2&HJBB/DIQ(1J_@AWH]C:O!K_,7? #.;3EV/M8/WD ^E![BT@,".Z)O"?FK.Y
PB%>/T9%'Z?Q*PB$[X"]4N9FF.E6LWB5N8]+,8#K?TBI=Z'ZT?IAC]_1Z.68U%,<7
PB42'1&41+W+DVN(/_S97L6X<!X][77%_Z3:&.?XR12]$L&+_UNZHY-?T5S][J[+Q
PH,+TM[89@)Q=69Z21G6W^%"5\UR8EV0RN"<0ISB!D->U'\P .O&6K]O\Q^'/J"/8
P\4^0B=WH4,?/LRL6!X)SU771JVOVY=FA%SMTSMQ,"OSH2<MOQ:DQ/P?%STE/JKY3
P5PS7&&L_QNQ#^%H#1M>^YGW<\47"4@X%=U^#N<WKNR8>0SETMJ.^X3DP:+\ZL[L/
PPZU:@\P8ZE:7_GW_[XW!P[\P;KSVIUN'*9"KO_].+R7'*T(5"F1^3S_%]Q26IC)W
P,4V<9;QNC);65[4:$JH0)<[B52#U]",.W",HQ#0G% H?1:3"PW**=)7\LS]%P7+-
P*/8%D"_#1,LET!L0?8<J%!64C3#/5)BM-Q.-.!*@IV%@5!&3QW//7M%HJ0$(3SF 
P$LBQ_%0EX+ ^^+D4+_R L/FBX*G2!!621QWA9.U"1DQR ZA&^ZO?*M6$1I0>H,G?
P5)IH_WTI$%$$0?[^:BX&T!6@+2<C,@+47^8EOLY043(9LPJS*X8I[R(56DNH:R6N
P=:0@]^I'20=6@Z<Y-^;1G%,?X6>LH'V*9XGF9XS*ZA?ATZ8 >FKL.@'AC=&-ZW4I
P0QI9RJ$+<6TS4IMRV[D?GYDBTM;K*>Y!&J5=(,K/# K%66LUT.7%K">J5<P6&AD7
P9=SJ_5C.&;BE+-V?1=(X?]*$4$KT9^B%RN)HK'UY)M!I[)S8JR;7(/)P1%(9 NBN
P(3>%P>ISJFB%-QT!]T/CB2['-AEC'O>&N,0[,[7@XP4RUB74@(]Q86B7.JNU@8=2
P#!&S<4J(K0'ZQ /D]5248&L:=2"<S.OACKQ^7IM#!V\\*2 =>59%G"VF 0L@B*#S
PI_?J^R& Z75;OI*Y ]"!?UB*/)R6H]S37CS^XSC*6/B)Q)9!!9,ESTB%#QT5EPK,
PO9^3'HGV'=T)@4+:NRH<.L& $_?F  U!3)\E4;G8^+ ?-0@M6GNBSU\^>*>2_4!+
P6%+P)@/&A["W.!@ID[(B7S:4Q6?]'/+J6F&9[FL+0MFNX4&(0\@CY&X6-.LIQ&DZ
PFR-5,+C['T2PT/:[UV:/L'6I:L;^ZD!=?;KB;$H3U9K84'G<4;$P5,N\!NV;7>QN
P',T<_C"CO2.B*IUN(HB&2 Y0$I\X9]NO$EPV>5@H+%U-PD9W8J07EKM1^#.POZ,9
P8ZP61=4.5<-#K=BVO%J;\3 XVF^*<CZ#.NX-;0XJ:WQ S;#79PT0JKAO<N>KK^.Z
P[@'05<4&@6+M&AC?%F4_W@.[S?B$SWUC;Y?8*N33/%E5GP? YRZ%S/W)>V-%9Q,@
P[3B3[V;"K5:"#[/!WRDG173:JLU]!9:"^8<*=L8;-I C1QV B>BRBHN)9*+BF30^
PA1BWXS2%RG&H4EI8\)FBX%IWCU/4/LDFAN(,N/1"2-E),:E[L'&8\&8#@3ZVL/>-
P''!='??\-;@)%!T.=J5-4-0PC@ IQ)9/>8HSE9@J"_%E-T&[4/%B-P[D&PR+?]ZL
P8J=&Z;NPG&R$]H)!BSOH&),AQ*H\7]!]< Q9_F!GY6 ,+PIK/93[%?@AH??;;Y<5
PN_ HM)[MU'I;(_HZKV+R?AF\7+&2DU;"U&F _F<QDKP@$C5HMY&YL82[JDL:-Z9_
P^73$_O2R_N+&^J+XJUV6T*>YF:KI7$I(ZFKJ#U6X\MB"!E%^%=/!L7?R4UT37MX6
PM+@\2_8M6(Q^;VX2U +C-^IQ:*?LID^9#^;Z0DEQ%UE>E%P"D0$5E0Q:?/>_8;EY
PKV_"_8="?1!JCW[HG*X5IHS,Y=<]]ZC)1B@Y!2-W742@0Y4Q[ZSS"'#P),\TJLK@
P.HN0QL,LY&F+?]8=T"3L7,[5).*]7KJVW4#/VHN?;ONL%:?HK B&>Q^9X]'MAV@D
PCJO<S],F:F0#TJ5M^%,.2=RDQ$Z'R^< U#@G3@=0)CGLV\-"$C\15.;/@;A-FGQW
PM%4:O5L!5Y/E&*H99#E?!4ASK9I>@)+G$=6FN!9*AFVE:%H^X:]_$^+>4B&1YVVO
P!7+H^GW%_F!M5Y?P=(,S-6'3\J;.C/FT!Z3ED!OV!XKJP?L[:X(V[-4HQX0)M4:C
P,Q!B[<797I8<]-TJ'2/R?5C"0DMS Q9+T8\W]!(@)^,/]U ([6CU'N0".4YX6$1S
PUCB^CI5A2;*$@(GZ7DZ%!_*X:WWR/C#T@?&A42VHB(?*N+',ETTS_'4;+PM_S)O)
P6;]K,0?U3RT>OG+XW2,-8AP\@J2'9HU^>J,8/H/')8\O%]Z SV"[@3#<@"9GF6 6
P$,%(I[;J[J*2 '>%=+8RRRDR?_11+^X#M+[L*$D$6GM);2\/$G+\84'V%DWAIJ%'
PFR9*\3;0[NN#^ZC(&DY)&16+?LQ%&[ANAX"=*TJ\P 5F=WCX@D7#6K;)C6$[(]4H
PL3 ^M_+RBHPCZ=1M,;_U1@B/Q#KI<J2TKO;CC6;$[M(>[[2#Q(<.5.(S_80!JW9&
P9^SI7V?K)[64LHX7O7M+*9&\$6.>H<I?KE76@=)>/9:-RD#&F?$I;]Q[;;"A]5JH
P:P,) J;%8<BZND3%0-VBT:Z&@5,IZH]%01HYW$8I'0I:QYYMN<^A<Q:Z)%D/;^I:
PE_A25#(5ZVJ]U4=9ZR+"*$?$N(-!V1OQ7-F\)EK1ZP 8!]\';J[CSTF#V0A>&:@G
P+=/:YC.D61G5%#W"FW^UR[%1Y[391AC_,3:@EQ!@X?V 84-KB1Z#))X7<V>(; CA
PB'KL>]YMEBY A\8H!G$=02U6.10?,M!73@' LW@P!,K<=2L5V$=@^?)FD3/<1C*/
P& J^WD1G,KG4!GMY CX<L+K/]?&/49N+GWA>5A76%FF*PWKV^K^RT1;8S(..,]M1
P<Y[L^]@<LBE B3)# BW&S3,;N:R2H+9E> >M!"3$T[<! 4X;(4]_5#KUN^D>:W[E
P7?BV2O[ "E8 +?[6_/CL_/:RNJ7\@@;Z\X66F#D62YCVWKMJSU>@&9.M' RV-;.(
P-X)ZOR'BC,^_"]LEI1J_MG^4??YT8<>*?96'J(>I,.P6UJ$\\!Q5=4*9"F3!Z3!W
P0%M@6G^"Y*\0;!QFU$$&_:"W> =L]5MLXL@O(IY4=32M5BWEP*KY_+=$BP0<RS)!
P -1W)LSM[<Q4+0[WF(5_TFFI]T9(P6@0V(S1Q*QW^&;H%^QSQ#5/]QPU .EKOH;A
P(^E?OL8@T?P6L^L!*<XASE_*^:\_/(M!Z?[G*!2L.(Q+#1AT+1[LTQBL2DL$B$>S
PZ!KM1)?1/KA4/ KE:+(T)8P[ 0\]K3VK='?<ZW.!L+P7;UC$ X:9!:8X* R@ZDS"
P>?ZG%E90$3I.R(7]HDESN!_FK\&J=A^H(QX-)IO@ 2X45 (5,;;EL3!0G-FWLA:M
PY[S/>#+TM1CNG!,8_Z>3(U+H _S@("4DX7ADB86H1ELW3CQ#$.Z>.5>FLIBX*1*/
P40H-*-Q-@Y+KJX6V?N/#A]LHW=[-[8@V!P$2*B2<3[<NI3<F4.06TR;^W%_7<!%\
P!)6?0R\01@.I[H6BMW>VL*_IB*Q6IN)_*&CO>IB/ KQ"L7LS+[-S7U+U'S@YAY4<
P/,N"HP10LZ> J] 36;_65LFT0118@E25GC4=5P@1-U'ZWJZL8Y=  W[4V7P)T-^%
P#I(.R:LQ^YV>/&A(F!K5EC%=<:7U*9ZIU8<[D+,[$>H49A9O50VUW.B:!JE]"3^=
PV:*PAWK0\<MG+J#/Q>9UN6%?V6X(D'F3M!FO.L7A%JA[[0E9[G+:KO'.F*^%GOC,
P5@=\JY3O@[;;QYET# \"0X5(FT,3F)B<W8JE *4HUN#!#'7 4@IXY#D13HN!J_&"
P0:X3.B.JF U-K6K/S[!AO[1/8[#.\P9:GA/%H#USUIM GRHI0DZ+V]3A*^PO=E;@
P,(4A%+%-ASLB*Z+]&X;0[- C]N#W7&PFF"H97@LN>:$TD*$>3_^CH4!$HH1/"&;H
P6[[HS%R+VYAH33<-;E/P_'"H8U!HHY[Z22$)?QC8V"P$T%V1XG[*X28<4@4<Q6,S
PAUD.-Q)XKQ(SV1-343R)#H[FMW)P^"OBMN.'2(MY2"9N##@4#W;M'>+QZX# B#[>
PAV7>M&B/N-J!%2J[A%<S7[=S%J]6+G&GI7!>S 0XL@G>NI[F1=FI"2D EG<1;DQQ
PNWV-8B6("JGB<T-1CM9K%!]?GM^IKCT >4:;KL-([!3H3JW4<0Z'"+[J]662V.A,
P+9_(3X3]C;18YIE,NG32,3GKH!4I;H0BEKL( I<_,[1\?97/-#-/<12=OK$U:P17
P*-/W/WE?"TF8Q6UIS:O9^0R%.C*ZJVQRG=2\0.<Y2T:3MS:HC'IYJME<EQ%I%)E[
P5+HK!*3(<?,^L)/G3"7\S!*:0"<#K'HTNI3NI(?:+E!_+[U@.1 89'[[C>2"[(%U
PN+SD.?BW@J'Y^T<T_6YM9;H:9\0[&5_MB*JB F7DW)+=3-:"TQG*EC$EO_J5K*9>
P8761C?9SUX1%YZ8L'AU"=M#)<"[]Z&2WQIZF1UJD$>(P())X3>@?D;5)_FT827$*
PXC%^H(D)^,J/^41/YBQV [/"1H\>:A.'0W4<FN09]#CUZ>.9=YF"]_$.U/X*FX"+
PCDZ(6O(9RP30G):*>ISHQC85-(ZD[XTR'^6K[;W-GPB4!UB+4]2<M@[T5)SMNE0W
P=5F;U?E4I<-N,,U 97%]&R1\OHVYF*D=][[C][A%BSZ,EL_T20KS;%_5:11J+=6\
P5(/-Q*0+@0"FO-".050,63H"/+\F444.=(^9E@O;AH;FN8HK0!,/PEUJ<N-#L$=_
P4? UW7W6GW?88.EC0X22FGP5EP/Y$T^'^/"4U@;><;X@)"^>XN>Y-B_]L'<<PISU
P, A)47@J@5*ZPG(VRCUQ]U ?J[_'A UB:M-+E-VJ[I8"0.:+8EYU.6[*4M"')E'L
PZMP/NS)?/J.,AJQQLIW#L'#^2?Q)!D]7_>*E+@?*/\T\.$J&<SB33A I_S)KBB_9
P#QDB!B0[]$1ZGF'LDIAQU*6B R4.-DR/\DLW(('N=VU[9DB,&FH\_@^'LAGKCMB9
PU7*]@ ]MAR3&?$#R6K$:C/(9+@GCG7>:A+P#CU:5+(M K"V?-?,NI.@5#*6Z2=B.
P_MC*+@M1D$.<0DA=F=2YC-MQM"5RPLJ"A-^15!) SAYB\_)^R!<J;>X'(Z_49H?2
P,"Z5,";VJ[>J[,1ZC=)\T$)M#_:3(SLI?<0287I8\)MKTQ4@)91  "NAJY@DJ8OC
P3PMD/_2A6- D?7? /AQIPJ??A97JM%HT.$S?1N7H] +*PUKT83)9P\3=E?63R,9'
P*H>;IUODXLI\N#6);](VC88I64KF&53<1K.+BX)'B&L" %39"/27?DL]??;FZ<."
P(-:'&_0&:7@@$UFE02RXJEY)7J_S-:O*_:Y<0W#UD4R8]09\ZW,1\%+\M.-:F$2G
PRF :&= V-;PNCT*QB;.]WP=N@S#N<E<I0<2_7T)((K2J,-MW32.9"+*M_?W$=?+ 
PB]GUG9QHSDC4!P,##1V7_?<*T9R[?B);;P.T")5'CY/3'19JHFTWD=CM".41X?;1
PD2N%B N$'U,W"FU.A[CW2M\*A-!D<'>H!^@JF[)_JE,(%W,Q!?&'41A>Q3BZ[TZ-
PD(+7KX+T;">T>0?BRBZ B^#M*"FPF3\;KTF-X32<8I:"@Y'[:N_R[+<7BC>(AH8F
P5J_S&1WJ:2C9(V_[$YP9HURT^2%R?A)TKE6U\>QV[\1%.Z-K&55EV]%9RW'[:S0I
PD>@I(=_ UNOM>FG[$>NH$!9T6V( 8-@_:_S[/S<+""]?OH\^%,]=G^S#L,FA!4^Q
PQDH1")+A3W)D=5UJ).ET*N?5,75'S71"2B>_Q@VR$C*$,02K*IVWEC*53W\F$\V#
PEP@/D%O<J;5*F&NZTKCK++Y8,UUVX;W,[WV>=MYZ6;[G;#$*GOR?S40E<BV43:<0
PJ(]$EYDE& ;-,:?OJZWT CS5HJ-NSGCT><8LPE6BVCRCS,OP3'Q6CQF^-4?\]$$C
P7?EKN](?&6D'AFZN,_<02)JH;VY0/S^V="V4S,RZH 0-MH7\SC]<X!5W6*1BJ-,$
PNI]E^&]3MKX2B YLUY('<^U]WMK=/K7."VHQOM3SN9F,N $)I1G\U&6)?]6-ZYS"
PB[6?R';L:Y#[)606$[?DCC+<O/O(DD;[^N"RA9Z:TY K6 PEXK4,:RZG2C@=)2N*
PF6IWC:Y#$5*9S"0=55#^$T4_="K,0?6_Q!_\=Z-/D'G1GVGY\,6UFOE.J1<7>]XC
P<^+6ENJ<0J3$O-GPW&%A$,+/V(*!%_(GJ5<A\^"27:Y9YXJOI-NJTPZ8(4U1QKUF
PVC8"4I<3@TM(T!SP=YS9+B<^ \_^+;<^]ZO?9795!6)F%1!T!,&^RW"'@"%]/R1@
PQHJ'.QZ3R&'RAW!W;HR%BR7:5N^Y*+W1:E:<B)=Z9Y/>X&,05UP5G8K4M2^UO:TY
PIX31!NB@?P"X<&28N!EERV+3ACD'"0G6$#4# MU-.CMO_[X_NBLEYM_'GE,%%3ZP
P0'J>R.I^<D<.&90W.E55\ESG9)X<^9$Q3JP;NDRM//E_6EBXB)OFS([W' ,^!*T)
PQ<7\KD^:"M9UA1Y(DP7%++YA=B;C:2V^=*@'1_JWS[XC4TH#MXPLQU"0*2P@2RL'
PNWXD?=QEPYME? '=2<ZX*'[D*#W;0*R>'PB*D\)KV6B[D7O]@1V\AE. EXE'GB^>
PBL,NR-:<('*,7CB9&5+D?'I[)TCUKD!N=LZ,?@YI!(G;YCX7D,NSH8KSDV* 94:9
P6&0K'TCSI?U1Z/,8W1G$UDQ64K)6L1.>@3//^G]X+FD!DSZT;@DTT< PK32H;]*G
P$IK3[H]885B/XZW+R)13YJAX^%"Q:W<LJ%^L M<Q>6$C""221-K2)>(P4!=,Z$B7
PJZEPDM'1G7BR09F#J+[;)^ZP"HEP4^@->RP3<R%G.>Y$SWTWE'&)FX-FE:P,79X"
PYUC!Z<T]8/&(-_"5-*FXA/-0-C="10E:*":K*ZXA]RZK""&_M:1!:DC^5W^D6!QE
P68!>02,_W!6"%'WN!FS7YU-B!;#<ENYV.Y>?LUU#H^'/-;G<@Q43BH[A[+Q.JJK_
P'=J!_4+E,1YG^ZX,,H$B*]U%[$;9470+3=$D$-*:&&6#7_]'DU(Q:&W][3OY/D>^
P_0L)=EGVHN$@N,: \C&3Y.9'/9N^<H!T$FZS^!& YXZ!?SNYYUQL@H/@ET FW4Y9
PACRSEJ+$Z3"P G*?B*.&GGH5;B,H_+#I#2KIP^IP8/$YETT!PM,'8<GF_R _&^,4
PYB;E9#.\,\2BW-#G"JMF84QFXMS,\EQ 0=0YSMU43V#W6Y#PR D!9L<T:[0Q^XEP
P!2=G@E!]8]\?K5X)SY4=PB!M-Q5FT^-[DMXB+?K\2=/B9D-RR35I[-";Y-YHO/_<
P+[#$/TY56Q+GM.^4ES[*S#(VGH:(H*2YM28!;M.6_'8L&2=GW63D_#5O3.ECM-['
PA.F[GN8@P\$R>1^EE21-W1U%[V3]9H@^H7%VC]4=)F[G)^2+6U]FK4>^L"?D$&/N
P,W9HQ" OA9U*-8-BWL#\4-!1"?&&<ZB-D0P-V5\SL%(Q:/'BU46^B?@/N8'%:E@<
P]C7<G^NXV=% YIX9:\AG^K]77S!/.$G0MK>Y924&O6I.!X$,(DZ8X<RF@69:U+Y%
P-/CDHB6&MW<YA0#].;:,J2%_A,GU\8I"?8-6U58DL<31:KQ#"U4QVQN?NP7(),4Q
PEA3!,,.-[,&1,@<ORY63#%T('2  A0UC%.#PLG.\IW9W<XS&0)V!=#H4<T!V_GC]
P]\ZXJXWZL8Y3LBH.<!O*]^-3=TX#_)L /R$Q&:Y"G>]V18DX*\,QB7=@5#_C\15J
PKB%XIQ*V6X7@Y(X;J]_H^=07N)B3Z5JKQQ \@V+/;9SOR'Y&0)Q:7\P"HNLT_!8>
PP]JFV-$FIW=!U.431/"AD1<'<-^<5R%.#.X&U/B5K:T*?KP2PQLLW[)CAE74["1H
P054S/R#IQ>#WH'KA,FDV@9^@+)L7P?2-=)G X3,5--#E(U)"3.P#R0,!?UP!'&WY
P]QH@D^ BN09$S<WC["?X<GNH744W;3M*^53QVX+DH^>+:6LP#?/?/11.[[F:=,SI
P"!1T)LA=+X0"?2<[USJG@M",W5E<=5T LFMR)NY!W3 FD,KX(]00%FML.)6/CCS&
PU&6$;*_,/S\]V2[ZHAAR+8M/ZDEF;&1]-$O;G*L_*TP91*CTN<)::$B-O+=JN0%T
P'"ML3 DN;SY7"QJ::NG9AX>1L__<X&NDRW0UN%%)Q1S_[QJT-+D?.A(1U115ZU>%
P+4#\W Q["3 D(NDC5@]L6C D:T:#/_LOL,Z;_2EX73TB?D[N[ZMZQC*(HJ_S3_O#
P(V+O9LM2=.T+J$74 99AW&90XBUK6GWM]+WYZ)2!#Z+5S#<Q/<B?3+)V],<*F/J&
P'R O^75M/S!]W>\NI!,O=) :[/?M*;2W:;JP^A[0&OV$U,Q2Z 0VWFLCH-KC W@V
P7+T(NMO6(DPO4U),Q7Q? G-3 *<%+,SZ3%D@4V&J4',+VV-.'AV]@Z)TO9ZPF'DZ
P3E@PW9%S@C,.]\78,:4+JUVS;&@=RC?<K6,'0L^*)Z^8)9)<R_'M\$EK0BS[D?5A
P->02S-+!&2WR(PPO,V>W\&-"'V:7 +"?S]U5:^'[>!L=Q!>8 [\B'Y),^@EAF6N(
PRWEU[VR@J:=X"[KL!&.),X3_($AQ19S<*[[.QRFO]L6\/M,B;250]L F/AXO68A<
P6N?^5T@61,<!+#;@3E&DP(35 ;IT<V.'8EUB75A2RWFV7;W06T%<)[E\I %!PU0L
P.AY7[17P,.;F9GBHFP+^W=B,$YT)$:+!]_X?6+BB&P1WO#B+KG 9_PK4/4#O5Q_'
P!ECBD;;1E EA3H,@(ID6!;1UFF_R.]Q6<:!=_D3M[4\/Q5NP& Q2HS_A*ER+LK]]
P,:%%C'G(!>JI&2D;QDD@>*PE+A!*[VDC^%^"IL"2ZR(L[ZK<I_@:^Y(]HE$W<Y.)
PT1G)*Q7A:NX>_MCQ"")R0 F""*]FDDX'<IQ#UD1I?#%=@Y*57$68WGAQDND'75 0
P ]ZD^SES\.T!QV=K/J577KB2+2VY%I"4Z92%N8M.*(B64= .)Z&\7#&,LTT=%L\&
P[T4FW$R/965:$"TD9AO^XS]%0G7ZQY:S;3DC_K Q/N;G.IG6F%OLE]?B(J5MG18)
P#MT9K(<RFAOUY#HUSQ'D)?:3X#'W+M>,=*M$#I$$DM&Q;P ]I.2N,4$+YQ\EGR"2
PC=N@KYJODI5@E=O^>2S8[J(L(DKGKW-A5H.%0)_D]',ZR0YO![]Y48LCCQ22G."O
PFN;*6-RKD$N MJ>.B>X9%X.*?J%\$U#&Z/8C2L*X7,L3UV-,M858+P_,IH@15$I.
PS=29/Q@;=+)Y0MB#'IZ$*[L5KIL;[\4N?U5! 82)GW"%HIO=)(,B//FXNSU6'X;0
PWYC,HH#)WO])0W52T0CH$\K]CR?IN_61EK<\A3T9X*:(6 PL_P.?7L79!L NR*[ 
P2!'XV_"D,IJ'4?_R3/LV= J8:0:UN+#E56'[(9B;4L=C)CE+0<KS;@,"DCO7?TI/
PQUZ\=Q&N]\I-8T+T#70N&L\"I]GA #<&8X$EHM1M^@7UM.]"B-FO,%"?".@"2(!U
PQN,!2RA'G\'I"#H^]$7S=A+H* F)&<W ?8.AAK'FT$ 6\97H7RWOD%F<241%$B'N
P5>%< _,QA,W"&5;)Q(;F^A$B+LA+I0HG$>\)9@I8#0.5VPZ*+M% J<IW4JF"IJ_:
P.FD$,/3.&7%O='"P&-.5$-DR^P&>E;D;\11\@)):+]_D)Y3P9&RFX'<]G+(T1NN4
PNZ9IW@:K3BR->P8_:SCJVAEJ"_?X$3L? XB5K=X1((-Y,'DX4XFM"MI)Y'UK@:P"
P(^$7\]-MPKM>&(PWE0FQ=)C@DET^KQ ,C]<0Q)VK6N#0]L__AWE%IQFHH?C:V#5%
P<: &0D YF6_- P8:W^B)V4JZM=!"(&H3GR#X);7BBE--#%X)1UW?28=-C1]>5VGG
PF\<JP=O#FG%[K];P[%LFNPFT\C<W(-,ST<9E%/R ;OD )D)FX@F3D,\7TZC- L=T
P;+A,6-"LER8REP*\;]"PJQE4>@[J40W8F8SZ&^^*DWFB:QT=[]7>DF)?TT-H>A,W
PV_[9<),^'6Z^UK&>7,_&.1* ?!I55[=,8X1?._E<Z8Q9FN,L2J*/KRI.4VQ*@JA>
P,[ G#G>:PD/YZ/=.3'KR9J SZWUW?#ME)]2]?!B30"89&2UQ=Y'RK@D?+#8OUQA<
P"L%Z03!@GR&H>:O(19/11,%8<U<@ND]D\)5 "QJD9/Y7I= ?Z(MW,7B0!83^09C5
PF@2N#S UF!IXE_Y-!(E["TV@$QCT3R HL>R#T,FY&!Z;9#?RYYI*HTL,8X&;TIOD
PV&-76M>[#+OEIDFY5GEW9#;F.D;=,)NOJ1NH,M-PN;2Z ?I0VY6A]!!&@]++,5/#
PC<;?C#D*4E327_ [85Q=-%[;4MBQD)$CD5X8K!0YK:3>2^@P'XU+S&6_@J##*38M
P7)C8W=0XR @E!P5P"'$]872W/0%311SD, 4>VYH [3, 9U2UDUF0:-?D98LAJUMN
PI@)DT(.D/<H 'CV-O:L"J19>*?>LZ>ET5^H1GY=(%-\VV^76@Z1!F]4TF%0![GJQ
P**!XAHS4UZ05#L\N[L?:C9F$A>I'+NUXN#.Q/X::ZHL>J0@M2/- =M.>UK5H<03X
PN)5>O,=;SREAWP9KSA/&3H%"+<(%3K.Q: 6G0+8!:UO(+YY[&Y0-O_OK:!XC\M/G
PRM=>=!K>0@X3'R9'#/$S<+H3AM#[BU>Q/(@I K.M1R^$.2$4<P 6!BW$)-A[%"O0
P;G%6M,2 +U;K3BV8I;VY$\!?JJ^3\="-I:X*5,JI,9-FM-_+-/RYPKK9R$Y;GI@-
P71[6YN1$(>+K5'.PM?D<#DV;Z2N9?Q7'?]>SG*^,^T1IG] 41>9SS_K6?.\W)",7
P(*&;EPSB)+\]RF[ +_4(9X/IFF3]DTU'FONJTV>8'CIH&SOC5D/ ,X.85M GHD0E
P?2&2BHN>7JT9)VLP+MI@Q:Q[JC(;%$Y<<)21-[TM_R86J((@K]4GD_ZY$0\XY4S=
PA<Y=R':7-AYA=,2U& :<H_ _!MU0M5X44/0R"]Z3^PPR72:^=@-FJ;Y?':<9< ]]
PZ>%Z,[_"P*(OGYYDH8;7E==%(;@0&@6!"B1^.4(*#/3$=-_M(] !*LQFJ&^).<]'
PKH06_A@OG.DC_+Q;Q',)[\MO>?A:.HF<Y(*8W>&'_=.U>@Y*@%=*U,4/^=8@\G_Q
P3H+;)&FV'B]XP5::K4/2=P9S Y&9WD:>"V3-&!1'%W5AJAS<E_JYRTT$3&F@,C@L
PI.Y=RX@APP=*T1R\LT9>.B,'3%H2X2(BL5^0:"IBX*OAI-D4,38!XF; >L/OB./=
P$39AO!Y(0X.$9^RBR75VMKD*&M@V$6B/4AKM0T0,AFJ);"2U@.?1=U9DIB;[X2CZ
P8^3[>7%K!9895V@"=Y4832F>2_#";@'.JX^CV)D)\Q!DW[S94<$(#D,AR/CXHS(>
P=W+ V:$/0]H8N@["C.U."BA]T!1ZG>)E.:"B0 (N7FDU6H[U/_L7XG$UJIA;?T@A
P)4RVB07J'TJZ&.?;M,AIJSS*[L]5*P3,Q7O5/"*JXJDBXO@RYNW1\6_T\(^UY<$C
PQ"WTCLF=!&@NM5\25(ST5"2U4ZA\R6^Q_R_[[LLUC%0@Y-=5:@!%A9(Z.#I-2K$_
PPU:TK71?B#E)X3)J=VA>71=-/RD,0AI_0VH;;!0T=-V(\D]YO'6I]U03>5T>LGJK
P!V*QQVF=R0!'K4M<>VK1CU*V^(HY:F'&E%?B1TOUO-UM2Q!=7TX%BF<$V<(4\;Q%
PX1UK$%\4%5O^):5 P@&3?2H2"UF^6L!@.<#Q1U/.)X*N6RV6")WM%GWS21-?A)O^
P?E5#1[,#<B?%TM+M:;!:-O.LW0X50H+Q)8[+^VD29K*;4DL"+]T*T\9<?H#+K/1\
P '5>:8K87E[.2L2:UMWY6C.]1I>+/J&IE-*[&"MA"N@ONMF*"_1 2Z_OWEY1V +>
P\MOHT3%HBR4$V1%! 6"<#]'9J!Q@UFH[;'[QI0_26;UCB5^!#^\(]X#-Y,_P;J^.
P%%-&HQTM7,QQ1,7CP4""2D>EJC+2'E!+ZN'@I)IS_/U>D^-&)YH,<E&EDF(U#I_P
PFRH6,7G5,,Y-O:-;'-[JF]0('&;P,JU%JH,-A11$3BSM@KNZA*9G&@+K=\86;]A\
P/6>O- )C\23]=0Y7&62=>U<ND,\"FL2]N9A3Y?,4O#&?WET1,$9<[60^UM;9*/%\
P3MPA^4$]*WBE_) JAQIF,(/:B2R: TJV3?(NF_$->1QA??+I])DJC7%& XV##E'F
PA-^ED49^UKH76[18T0[0V!"WQ$0W?0-O?2I*J9R2&5!@*?5 0SKE/1\J8.S: ZA<
P221&/BHJ/3.8'Y9=_G]5>\70W]4?NV HR<V6.A@];FYDKW(X,>(]&+G;O='B??DW
PL3*D3R!.N[\K;LFBZL0T=G,/7&AU_B.D*4]!8D*Q>]!O7:%!:6Q*[Q@0^A/IW4ZI
PL)A=EZN5QQ'7-;]\?.;HT:MDTF[C"6>&\LSDR2W<27WY JNLM)@V%0?4RIR:9)3&
PU0>3?18S:)5(C@7.0_<7K;H[NOFP,9JRTO;#$DI*)Q'(FF,3&4PYC3K=$]"#Q=[9
P\ZRC:-7\NXRF[R7RO#>9Q$N?,]^<"/)>1A>U/D)@WEOU ,LP+28Q_B 9ND<I6\FA
P8N0%R[#2%]\7.$C_\YN=3'[D6V.52WP#1_H64 \09SFX<]"8S*<:T\/Z<'R,O,#&
PT<39ZYSHV3.!.:DE4>G&1H%S:I.D?(Z7#SOD8\Z;'KFD6W>,:&X1(]O2'3GX497O
PMAYJ>-A#EAO2E!XG28D>6S$W#"@R]1[K5Q:,<R2CQ0="P(=8C^84[-.DN\?7<]7Z
P3>K[WV;/)R\@./I-?/R=F_MX1H)1R=?Q,V/AU/[!9["? N]GK^00%&=*3^7<JY_-
P= -\9B%!(A-J$PI9]&M9\UN#$P,XEQ"*4 WC3'%7R04=UUTI$^F\]MC2[3XNG"[1
PT811.=7=,#'Y\1.7OEM8QFLB1[)=;AD4];M.%RS:LN^& GYGHBP56@O6FO+__JQ3
P\V";WCU*Q8I4U5+\&/DLGH[E)63+E]H%9YS&CR2S18#YB6QT5:56M]+X:IE(J_5V
PM8-HAY_4D$=*?Q[3R?$;\-ZMLK<?<94HX#0LW(6I$APE-.Z%7*#V;'=1VFKW4EG>
P,=?(IA6WDU#?;3!&D\MR6/W*'Z>.NC:P[*=+/F5TG0$G>C%%#:KOQXI,%F&IOE*<
P4GY.>6(#MJWOL![2M<Z,01IQ9596K+4UEPN0?I35TDIPFV*GYR++F&>P'C708TA/
P"J?=ONZ1Q%[+P8&8,><@%<4T&CN8-%'3*R9&)9R[\>0]AEYD%MUU1=(:B.3JY*B)
P$QNDMM21<J"E<6/+(QL+JV>@8&W@;<%]%]G0(!L),CC[I(S%<MYK"!P PC(?M7R7
P$UZ*AZX5,P-?T2\V(/I:)OTK@H[B9=H<G[:@JR8:I.N*? ]V!#LQ4UH0.^:BL4ZZ
PS:AX+G:XQ> ^-C#CEN9H(&13:-O28N<!OT^V*4#\XWJ_$+OUT0G(QK#GH2KH-8GM
PI=WM.14!JDK(-VZ '^?E0U:9A4T7XDN;I:2-,T*JP("G8/ERK;US2VCB<\[98!GD
P?R3 ]LKYMX)DM++'/8A^!E>HCF<XUW76H95!/Z#00B.T%%D/9*^+ZLC2!"]@HNK4
P]R>H:*X';V<)X^F ]D7E'TQT)3'XW149S%"#*=!CP4;F]G0!F C(G0Y?7TTN])[)
P]$>A3MS,,:HG8(%]"@FXCTV;)ZHR%[,:9E'Y';$MH^L24324$\V(IJS]G]Y/Q( "
PL '4L#/8\EPWD!:3#$;QR-F<7 RAQ@1[!,-.),'C'FD%=SQ;[+18DG6U18.V0_H+
PATJL]:KP6/G"<@A]=D:$PH 4^1D#C@A9N)R90ZU"P*E1 \P"_N)[4#&H;S@N:.4D
PJR#C5=]OJ-Q:)(G']E@H:?%1'0@UE?-GNSA"!B>&118S)/@EVZ];&("('BO7*SP*
PQ,_B=#)%3H[CF7J/96V$(V=+M3_T5'&M:S:4D5%VH4<XIN:^&I%+)EI9O\9/5$B 
P47V_U__$1.UBO)S7F@;&O\/OG.;DU:/9RT6&$!L\OT&=?M7PG]:H+31N8WVI4(P#
PT $7-ZWQ4DZ??K-/C!7.$ U!%;E/YZ1P+QT(_DAR!)5(_ID #\-:;R!5(57!Y=AF
PV+NO&&W[G/ "EII=8*12_6X\0)_9:\PB>09M"1*:@WI<39+KDU3'9C0LT.0%FE1'
P<H;85QAED0>*\)'_/]H%#_NW=_BLUQ.W'_A+AT*+PJ6F-489)+ZN1/@S=A6(2O'2
P?W=&%ZK - \"5XH2EK6F["V2E>9BD!F)P],7?-04@3Y5$1TM-JQO3D"4C8MF1N9Q
P4[\& 2DI@\F1GJ_"P^UG8)2M^"^]SO*#$QL\!>>-SM6- 89_T]I(P)N!LL+!KYLB
P/W?](6?2GF?M@%JR(L,P5=O;WA2\HYIL#P-1V&?HE@@<DMQVVS+-7%C9?P\HT@6N
P*(SUG3'R'M;"OV._G/*9&A/B: 1VTC=\@98M^$]?WI=T9>9)4E6/S*'.:C(,%R90
PM4+PUR2;, V3ED^]A,IDYKWLATP:\_]TWOHP)N4<R-1$A.KM=?.B7+TNV73<'(EU
PT\'UGO4#*1-.?M+ N&9L)&=^+.D@R6&A=U]2Q\"B1C%LZWEQ?$R^.XOS7,VX[LGZ
PN0] D9Z[)&0L*^XQ845393G^0Q&L"$H$;^!9]:7PS&8QCZN\?-G#3.<_0/WR'U2Z
P>6E'GL_8GT.,"AWY#DI(8\&G3O912:?:#JM&2Z(GSE.XKA#UTA"C+%M/X7%Q&2M 
P DM*/^GK*]JCT#QMG1KOFS&_C^QT>!)#V27#/;#X/YGV(Z2->:&\^\5S1!T^XK;=
P%$4=LRR4E&\JD>9>8EOZH2LAYKZO6-/,X+@3*% E-O.4-,\]T'<F&Q+]X<]&]CI7
P5,U?CU=Q/Y<PE>FX.+H6?W[ .MJ]*@NSC][UU9#<LF5*Z64RHVU7G4)UKJT_C^88
P6INJ3:R]@]E1#BCMB0*HSC=UE^S$_4TNDFLO ,W-@&*R?^P)ZR;B9 !XX0Z.I%1_
PHG#\[?/0TK_O9*3&I',I,->)&YG7CI'-2TH8,HA?UT2RL/*S@"7"QTBU]#NM1&H\
P1E\A*!?X50@V"9$A*RZ]JZ]$53TN4[9R=K-F9P'U3WIE79WBP82Y8Q=W8FI E9R9
P=<7[629+E S(P8A6$%NP&N6)X.)F3>L()X+:- 'AZY''&:, L)VFD2W(#D?R?T>"
P*H//S4.?3FF8@_&2*T#SUK'!8GB1726;9>[XS$!OG'_FMF$^#/ .!A;FH-*L!F(^
P=9I'\J,D5MV-4/EX=S:GP';PV>.ZN3Y,=$L?]=J[/BPIR.,U-8_XO,DD2Q:0)PY\
P>@(JOV =++OI(SITR-D;E4BGQG:OR=-STBDE?]ZZ^6?E=4P+P]KI"LJ-3S.4T;2[
P2JT[*'<L>N-D%D/D_Y*JJQ[U<;M[](K(*NOGBYSQ]'8^E_1H4? !NK;L :R(A=)A
P"JV)X);ZR(0H4%XJ]^.05?H5U8<O8:=#1(^1(]$^MA7(A.QU=+8Y!)]WOLTJ:/@1
P_R/76%<&@RS.NI0E$)7IHF:8V00P>R=/U^X03=*]@)%!-3ZM1OX<(J>VB(J-@WVG
P/= ]E#.52A(SP#0:F-PE>]3T?L+;V0<ZE4^DY:<S(#Q_H.D[RMDLJ,1]+#,+)F]+
P?FT*NJ@98)+*D=$UMFN#5LF-QA\TCTUBT?HF.<RRMT_R="ZL#+R@N8<D+@:;?Z,*
P<QHV?%Y0O1?<S!1 ;E7JP(_<^-94J!Q^$LH;$*%>Y3AB1@: 7R&1W3OS" ?* N4%
PDJR'B?Q?W/AT9LC5 4LR^>@L$P4$*VM(0*)>3^D[L?M_+<Z N9)OO=C09R!R-]0O
P"%JQDO\V;N"X@/9?UT#GT-UHZT_[*\RQ+J#MC10T"1W[@$<N,OR/Z%2.. -TV@A>
P(F]B&5D5P#&#U(D\<XDX6>X_VA%@D&N'C^&#D&O=3\%=9OUC_0]Y-)'OZ3YE-=Z"
P#)(0(6H//8;K:>\@ 6RQ/IB.QNA@S;.(XQN1BZA_I0WX?]/VG<+5!!BB7&EW -X)
PM7Z\K5CSC#Z)@ZCU@Q#_"62ZHL/_;,I?^,NOX >L=[^PFS&OE-37+I^C_-$]8YYZ
PROJ9@4-B:J^AOH3D<U#J6EN\RH/GI*:WJ;>B=\4.XU%.^*FSNQ]![;SY0>XFJ7V\
P#[/MW#J6$]Q* 9SGKSV*^,*KEL,/WSZ51TCP&'4UNWCE*X[+&[QE]RE4KW6.1M@7
PY-MP1[B0',8LECZ^>-W(.7EED4$J= LE+!0!5KUV%FM.+L=U@KX8 LZG(:+^\4)[
P])U+;S6B3A0%J7"OO>79/3-JK0%*DWG?5'O^&.C6;#QA_CD.B7Q+@;$MM5)*CO5K
P,702DFJAVB]D9XN**9T8R>-E)"&(^6U:;3DT#2C-7\UUFO"7<:3E>'WRY$DLSL/%
PVR$K^6F;]?G;C:ZI67;G.SET1IWC;>X7-H#"&(V4_097!A?,T.G!Z+U)4AZ!/>PU
PL<T2([6!6^G?1^(S"_6GFHX%TVE9(KQS^1T6+;E$\:UQ>WX@#OR %H";P/Y$88/,
P6J@^^5<?X<^35G ">]<M1JF;O@(E":?O ?4.I.LE=#'ZL>^G/G$</42XFE[V1^*"
P@9*>]5L>+/$=R$939B9[.E'%1>K/[.E;H9W^B'V19EV !UG\Q&=[)HXP\FE[0-8M
PT\A3E6.4:^8ZI]'VK(J92%/M5^\:.J6TQH7V[7HVG+=OS\?&P4D._ ^@]'-#;A1N
PF@4RG)[\9C^(PP0E;B4S X1#U2H;E$0C#/JN3#0(5G;ZD++ZV;&L$C8G&9G7'23/
P_E'<\(*3'QF;]:IM'7<: I#/-$]A4B8TQZP(:23LTHSG7NJ6EPAVM1H:H8"1V>CR
PGJ_E_G8YX%N,MF6SJ8Q0  12,FFDX'_5C".C(P%!/'2@6L]>?J"E"+/R_QFNO$_<
PX.(^_ R"2XRJ'BUL?X7$97;QD.7/)E.K?NA^H/G.L*@T,GXCJ"[8KWM!BT)@FI1)
PWV!7^74H/QB)R;H$:/.TK1*#'K8##W;+V KH40#8>T:.L<[R&@[FEYX%2I4:V-^[
P#0MH^3OGHBS(P(^3Z40-MVGNP[TZ8G3<BQ*UH-CB]I+Z0]+0P<8T 7[&02MXE8.S
PMO#AHF:JW>+Q6>VV9(;Z=:STL^E5;D(U)10LP;@O#E\^<*&='$F52.D0XGK@P:@)
PY4'3KCRDTCEE1+:TT@)#=B9_<'05Y1__!,1%BY1']\)KKIHA@]'V)IDD/TZKN@\:
P.R7N&GR.^?.28C6U0Y6\V*$'P8S+=3UQ[6)_&C,XC601<B_&9US(&CZI99U$>NW8
PY $[92[R^2=[ 51W&)/XL48N*0PKP[K]N_<2[0*KLH2O^LE,[J%N-HP+W26TIR+$
PA]QAH'U8[@BW2)#!8$ (X9<;+0>]!(MQ#&Z+,1 [X4KJ5-])J4&3%?0=28)%^F.Y
PC) 34H9[>RU,95D->AVVZ(<:.UL%MI_>\X>=#"389]PJ6&%&/,_84 QO]0:B8/AB
PR5P2JA2P6R]01?:3/*]U/6)H<BDE=!5BDT0I? G FA ^ZJ_9MOE=J59OPAN,?5:D
PDQ^5D+$O3,C-+Y#5*LQ2&0I)JB[@0BB( 3[C##[*_M)8H)RUSTJY^FNN0"O7$K?J
PZGRWY$S]NYL,<& 7893JW*>YY,U>:C,IF;Y*A@A7DMR]C&TCX\8!+D=_>_5<3-CM
P!2G9JW^N51D\!L"Y/U?5A[3<<9,>H*NRVRX2TO#=>Y(3%.BKVC6481B4G?1:.L4C
P.^:!#S/=,&SCW\Y\Y! BV:K/\/[3SC+!$SFY_+1@+LW(6MA491=4!9*7VZMW6[IB
P J5:?"L>W:-Y([?AK39]T:Y@>D=AW&%L?O@#T5M'],2LE( R/\C1'U(RF"[J;@W^
PLB>]=F6(3<VEAA9#:Z;!-A@G?124TXU[,TJ-H_$: W#[L7"7J'GQLRWR*>)CCXOZ
PB$:Z=-\XG+;2(+SYEHU.7 VQN55G.]^A_J[H%]=WTJ5N%XH;T>OW9=WUO%2EAW?Z
P+ Z5PCS;X>+1 AA@@II6[^UKF5(\EU&_)H+&<(;'9U2*([.U]&9S?RN\D9QM6/1U
PDG/D8/#Z7%0?\-##18C7GD56$8P8,(<'45#=)_RK57\L-K(ZFN0GVU(-/"A$<_2.
PUH!A(24((B%G?"_ S)V^ZP19?]0*:>KR5Y/) Q-/MDN:[A;,0MOF[3;N>F0C4^G%
P2=R'1JA8OHM?-2YKXB"2I1;T&$@QXS*!\ 4!@YZ+W SI)8VC&[$":K5VW-F!,-3A
PG<+"TN.A7A"!\]/B "$W\T.U11_AQG>I(DWJY4?)[RFV2P556MSHU.0B8QR_K:DQ
PMA(>:O9F:!DW:49O#L2"H^-/6JT_DP[@>&E>LB+&U4P<4$S&/^!#>QLV@7.@2.3I
PDW][&",5=XPT4P(.=SU)C%5&)1+$G.EUD>L; #7T,I1M3Y@F*UFD[D()07.]9E8(
PWMZJ0OJ8F9GULFS5"5SI[](SG#&";)A#7)UBR$6.]3%H$<S5;<(&B+&[MT4'_C4K
POP=)C$%?<\ZZ*-%S!G(1J_NH">@<J!STEH3?MTB#TC0/![>J2 EF.)JI?A\U.7 +
P ,)XF;V76Q\F.X?CE1^VQ#ZD7\7^CJ7 D\9;?_2GZ84R[C]1 B]\7]4T=.?T;)-$
PL%/KJ:^L GXF/YUS)'ZS"W:T+&:)AW>3[G&?([<KKD&WF-E?% 54+0(@G+O)5U7V
P!5.6)J $/1'XY_\PTE9OJC@LE1XWGB'Y96;_?7)%9_=#_JB1C)C:.H^P%"RBQ%W?
P%'L[XUV[N!>X\?$?23&JRUT]N8O>4<[,L+04Y1<*=R0J]+=/LR+&554TK'<_)?3?
PX3VV KX%OS8)R%@91Q:TZ"9(P"(GQ?H&['V-,QFWRF4.;N>+&A1E.&2]!(9E$^+)
P)$^\^4S7<#U"*M#DMNWS?J$O^[[.G85^\RWSAD=+O)%_C4Y<[X\3LY*?30%, ]MA
PQ!FV 2$)ON#"A L*?)Z+N5TQ%D'-L,X9F!Y<,OXA(T9JY5\0"T"HTY.'9S&<DF#^
P5?A_WB+B(OSDS@[F[OS+A(4$K?IKX^>IEG@(&\=,T3A4V65!M7P>)+BD/<ZZ%7DV
P@'\AV*V;'OYZM"G=W^X0O$"GB<U%,=+!\.69',!1#+UJ5&;L^B<?@IV')_CV [17
PK^TP"O@K4=N1B1EK%?62'&-T&X^(I @*DL63IK(W+0DS_9/SJ[DZ?$[+"NVW47[]
P>E[('#*(KP64!:)0F552%=S<":BRJ&P.QR%B;T0U>\6+%D')V%^[%VZDHL^#9R-#
PJ!_Y"B)/ZU>G9SK<;>+=ZBJNW6B$O9XRG7U]Y6.&T$9"^YUZ*Q7?0M^:9&E'EO%3
PVU'$-DQ!_W+/I6CZ!4;&Y^.RD0!5W?%&HKQ&JGLPZZ+9JG3B"R/1,\??@BXG#/:.
P('R]F/L,% 86]-[5AX+:NUYR5W#.Q();"6=F&+(-$NR%(J6)%DUQPB;6^B1OW<4!
P.W$IK&@63_"J/.OP\"\W,M61_0=)0*TK69+X!SAF(9LV-];VL?&@(]X5E+@X+T8;
PJXTOQ]@ WBCO-SSJ.IOA6\K_"-\YU.5GAK$G=X"_ >C0I^3AZS;$*51(9B.KJFG<
P$&D'%99T2UDI@W,\"@V;7=L4Q.',SSW1F((,,-OIV6"KOA=CWR*)69WK6?R<8L7Z
P:?YN]$V;&6D(EWZ"L_[=QC!?KS2S(8^$IM=[(@TQ_A+9Z;%>Y-]A>+1(C)4#3NCZ
P,>,1Y9.CB;E44?KFINDBAW-?!7?QIN8HH!4R*.A;E\7A1K8=?IJ(TW[*  6I@#0P
PNVRLN4$\&VK4:!X?TH=CF2"@VQ(]!,7 LGI9>*OVX;&_L9 7DOP-D^H9Z17H*1F+
P73I,8>)"BGS1^H%S@0)#&8%M>+,Y<&A8UTWD6V4P208(@K>SC$."?Q8X _)2JGT)
PEKLR/]?]LB&_=-U8'E0GD--\W].<_'R^Q\=%/(C@Q2W+O$&S$MBR$H_A5/L)\9Q^
P6S0!.\.)QD"MY8)Y78OS_\I>WDOM($IS2B>O-Y:S1,&GV!%HWU>FOH_[,3G@.1S=
P<DV27YKH\4ML KP:43UL,<VZWAD/OZ:%93.>3ZTO_G#V))W.1@*X\D[^>:4$__\5
P9@,&^_;IG^6\O[JO$L.S@ P:<34)GN.HW<)KR877@' IRL&1]1ICS/4*8\>Q[G)_
P<+0Z!HSN!.UZ"Q/SSFM[! [QH&H&Y+&LL^%?9*5+\&;R^^6_;B_1#VBFN?FLX<>"
P+8.%<EJ[/66;S]XH5R ;(RMNY@3H%SPUF.PO'QZK_D.XSQKA0/.6ICX0-@V$>P9I
P9WK$E;8R>.H*90RU>+R8=0+%?Y%?I^ZSW=K ^:,"V_:38 0(C"#2J*S#;J/ZFL-V
P"Q6JA_E58_+O068)17?,*7W43'T8?ME5':P(EM7V$%.!FE>>Y) '5;\CZ'NW5'G?
PZQ X?&,70(.^$W,V]7.T,H]WQ-\=%O_[K/[F'VIF[B- [&GX'$C8DIA:*:\S0;!K
PNKD^="%<HT)!=T..*=]@UXX%K53.H5TXLC7!O,4U!/&\VDGP- TEA#'$KW1P,QB+
PSS0VO)_W9%I(P98C3NO5N=Y)R&M<4BC5*11;@]?#G*I!#FL^5^\DVM<Y9$2BZ)]#
P$'-D(AB*9^<U9]FAK2246V+05+CF'V%C=/BXQ4'$G"3V4(9U@'?$'<6,L^5#,T8=
P-2+QXUU #$._[<4[>RHZ6JS=K].TRX%>D$172)I3V8">,Y[0UN/.%A;]['W'CTD"
P21U7>H'U)[Q Q(N5H^F0<O6IN6 G9VW25 )-T'9((I\B%FNA0*HZ,*?I(400[\:A
P'2S(#%X+CCB77ME4RDN)%B+/[3.  '.NNF>=>R260^$R)K<=]]3Y1"\[HJNWOI^A
P23F[^QX\,26Z7@P:W.VI1]'D&!@TA40O%IW<QZOLY0U/V3FN5C!"#RN,&$4J.:$<
P24[C0LET*%26A+LB*R%^A1>"KK^W3K?-.(:2BJ82$$>7/=<H?1E84S-@OIO[FCM&
PS:RDR0^5!;\VFK6T#V4NC-:E4XV&'O6%;AT'8VH>>Z0EWE*)=*9H-ABO*HXBYY$"
P[F\H%IH*%LN!%MF$,(.NI:.<']AOPXL9BX)X#D!Y]_A$U<@2:5A6(1X_!-1  S*V
P]H@Z>W\NFMEW39C>$Q#$XE96[26&@5SL!0"0R=T0>#U_RQ#J7F^K>YU:$:L^0-28
P/.N7TA&_IU#5(SCDA[5R&MWK,(%W%K+%PJ\Q']DCQKV?3JT"AQ_7D2 Y:96YYLV=
PEV<"YS*-'O6L^%;RJ=]'5^!JY.;JB1.QR*COKF1B\<(9Q 5!/%0IEB.Z(H8$R\97
P/XG4&[ Z_V>,,"2N]@G8T5BDMY)E8C$F_]4JI_V92C/C5WODC]_/DL2VI</4O(??
PXDF&;#(YD)ORM(D>W.2LVEB=:.2\L@T[^>'1P8Z>S:E&ZXLO)^,\)-KW8!N>0T.C
P8HWO[ICARD,VLDXN:$V$1TU!P&/@/>-/N1HZ6H7YX3>=7F&W3HQ)_%(J33_<RKO]
PGK]Z0UO(7JYC&"2__KD3:2D=-D4&A:$8A?PTO@N<_S9AQTW7FDO#_ 3SLS9G(:4S
PDRQWB<:?F+QW[XI,C/EO&GCH;4C0Q?M 9@5>PG;NFT59=FD#U#<#L?T5Q1 N8^0K
P*ZIXS)4][FV)A=9#^4>9.6(<;+D5/5D+G,])5$U1@??K*':9F%)T_9\":\F>62A\
P&;(K7MPIXY8XGB4DDE"4.=,EP>I;D0;P:$OSZ^$+A#C_1,*:$!_5CN[<DD.K9V<=
PGUN&441K!^;%\+^ 9PO9D"&HLB>%:3'@>=@N]]B42HOY4+5=<"?2F6'!#\W84"&C
P=I/I^=!AN<,L&)V!,BAX^T^)BFZH(51EQPSE?5?;1FIR16<<8R+:?2))2Z(6:UK;
P*OG06_QN\DO3M>^DTX]L3OQ L;Q6*M=%]D &3Y.VN<V5> AS.XD:@?):7[D"=KVP
P;6#;V.1ZDB4 :,RC=K1ZL(*^:V1K,XSEUQNRL! E_?7T--7*LG5&G]MMR-?C"VE]
PB0Y$@"0B$U^0'^(@2ML,.-_) \2V6QKWPN2-^IY>1A#X4R6C/52O/D@$F7M3?.$3
P["V)\E 12,"VHVV9M5/P3$.Y. 4_H8XN2_+QW_+?K'G*A0(7TP7N "K&0$&AJ0FC
PYD729E(]!JQC$"F?Q)T:ZP@/<;[P&GU@7];<.#T,T%$BDQM>@4I*W9)V7&74[[5R
P!]#FGKP).'^V/&;"J6L[)<)/=#G*!W)\[34RCGID-+EW'@G*OE>S)@<W_RU\SDGN
P1S21%1L$;#'1 ):-RW$'I0E.+JF=/^4>+N2P7J)#+UG^:!4BA==R5<R8A_=AC_QR
P0>-^NA\8EQ$0E/)7IK$1W$$'I:-D>*RV^D2>V5\BNOGF+;80_XKN:#SR0!<*W=WP
P<7.9L2KB(5J)TPD>=)QR]^2\VM!\I/<(G>/"P'V=*M+;9NY9?!#@K^L"I>&:V,_^
PMK5$U:P2@(&^+GX[*(1MSK))J@8ARO$<NDS3WZG( 18CV>IN$N]NSC;"#VW!Q68G
P78\B9U]?TOG=UX'_YJ94'S%$*/XO! YZ[O!YX\Y>3"B2PZ2LS7X'R+L*RN:&,<V'
P4(Y[0)R.-.U>Z;/?W89&R0U^%-^EW>'T6%_-^])Q#=W\[ZC)O/)]-A\Y+2$D9.Q0
PW:+. 2/XQE_>4CU-2[Q"KC]L:3?6\^!8&KPVMQB6G?L+<H\"I7(F':K21]J*^'NY
P[C0X+DIDNR%TJLC5<Q0^OF<8=!P9?'W$2@<.)# L@GS<"H$Z#A"357)R%O5L[9E]
P,NVQ9+PV,PC6\2$*P,$](RZ@C?R-HZ5!"UM;P^8IX<%/8,K05R78Q-Z':6#5ZV]D
PY>7F<STQS["9CYAJ29WN9UL)6;M8?[L1.QZ[/-U7CMGW>5L4$Q_'PFL+3Y'/[7+J
PB:G8,C.474^'_-@^J1:M-+/K.T3/S4[,J-OH5:V5U4+Y1<&$%:OZWY.1IUZ#F\1E
PW!+]#=$HD(P8B@O9"LXWT#?^+R#%2/-I0'N'HXY$P1^;W9;?'_ED?1!2;0#OYRLY
P;4U&!APH2_1W^+OW*XIK>8,VB"YVR%+"F43=$< #MTR#]?4H6'FPI0W_)Y3;):/5
P:$9.(MZL(9+ZDMS0[NG=;'(S$-.L,N1HR <U3(%<5?MK7<SBR0B!M"97U7..M]-S
P_..#,@XF0_Y1'SF%DV16TKV[\53.MSBR]O&U]EJG)H?NR+\2LY:U4,+/$$9,W =I
P%5%X)ACUW $0<7G2W:GW)!XF%^W /ASZ6_8/DADE1$TK7M"23L-8#3^6]$&#V6N:
P^!)8_#\56Y*0.*. 8+B4%#C7.E9I!XA2C6I%%:^HSYE?;%UR!R^GP0_K=3B_WDZ_
P^S9 \#+N]#G&SV+Q%<%(<,1'C1TB"W'8R><DZ!8.WT"OF/[&^H)B[<<36H"O.#]:
P)1L _88M<&6#C98HVY%)WX14;T_&9&GXQLV12G0[F%2R^Z+3W SU-T:HP=U@IP#F
P<S87!*.-N%!8ZF!+G-I6 2'CDIMJ.8! B7!CZ23FT$SWQH"9^'+I-)T!XUDD?AW9
P]&OLQ0!AJ3BC"'JGVT-VI=2<VJ;H[1D 7[C/V)CT[H9MS!5\X[A;=K#'U#Z_P4<_
P!BBG*6X* 6*1WV\E=!\)]Q*->J!"8PR,-GG1+:[$A%J"(#?<@D_(]IB9/=.@__2=
P]@$;R8%'^D&E _QG"RAU _R1"FPIT:QJU%^6R2$L5$A9AT]X2$ZC.=ZV4@Z)[X?W
P&<. 8I/91QR,C*3XSS;]W@E^XTY\O#F3[6Z"]DMSQ<L.FR)GQG;[D&KB%N[6*8_S
PX>^LT=67>]E9X4>^ZX-^1N(/C<_T-HXQZYRAY_P"6*J#WH]<]T0R5VX0@;YL[%&K
PMM"+S-\N<1VXG[25!OY9Q5.RW[/0_CNS+9(10CV ;6^F2P9S3?L7;>G@C_OY1/;!
PAQ*+_->)=GUI0R(@6)^ 3VHS]OT<P0 N^GK?%Y<Q1\[=L$1JN)1:;KA.%7I05\YC
P'2_NJP .*YO'*(_^$69LYEH1__@(X?\$P-R3RI @Q8^-) U!,3GJO,I;E3Z_<H):
P@\N>!W=P$T$YH."Z W9!^IJJLUF# L38]P"R3+#5IU;-#8Y@<\,==]K!3'H P0-&
P3!+[HG0X^V7S^F)-GG2Q[J?DF8XJ&%9Y_-'U&:V:M&?2= [.F?^R$D3>FIXZ!5JC
P9SLYR7?]DD:ND!-AZN?U\'6&]#X9WLY11MNU&C4Y:)9"P_QB2PTF8("9(8O9 _OZ
PW2N8:]F[,6%MV(J]=+!D^[5WRG'7BX:%C4$%"XP=R&! Y$Y,CNG$Q/5[5(H7FV"8
PO1@4?A49^<J0O1#R,2_W_F2=@A]4W"NG]< I=X%%@A_*CS1%YG;CH"#?RJ94W5H?
P-H2FA]HU:5)3'C( 9YX*IMGBQ^SZ_]X+B=/QDPJC_[Z&!'0@)ULDD8%?EYC$=,_N
PVZ#/0T=2W)2]RW*_\62Q ,]HLC:TXR5WAT^[[)#,V\3#6Q?3E/DX%.&Y2H7]E;_F
PH96?C4/&"0_YI_6VZ*&/.M 98VFUVQ'1DVK%J*AA,S(3Y.LFF*\"I#K% =.&34XN
PLG_ZT[DI,A:N+C1U) JAVY?<V:Y/VV&?S0L=>:T#KO8P\%QS[X;'BZM.51:3=*5W
P-RF&$(TBIY9,SKC0I>O0+U(8Z8P[>%S'[5SK#J()Y5V-AN?\M.5<P0"Y=0:VWC[M
PGM43,69E<4RH4C=D ))0\RA?H4E/_L^ #>=AJ]PF)T[3,@=%:+P@Z<*^X7R$1FGA
P_0^R_V2>PYZ]0#^S(HO7L32"<X6RA=6F)E<[IE0&_DN,Q/_7E&WA0X= UXWTYW'_
P2?J%J&[2O))9TETR.Z\&H^='3)TU,RGGV.ZJ<?9_"I/MGJ.$*@"N+8SAE<4FII?%
P:I&N^LW#NX8,%*X$D5!A0N_NILW$-Q7:G*^HC=6A@MKG''T [ :$67^H04V.FSQZ
PVR5XE]A6<Z2I H&'6O8>X/T<*/W@<Y 9O@(@=R2-,OWTDK0;"A=!Y0Y+TU[:\ZN 
P9G_ZHP5^N'GK.[1'\,@.<G8NU.C394)_WE:)\NA;)Y9,7!V;_O#-C1RN(%%IY7+9
P;0,"0X$#Q1OSE^&'*BX1$F*YH?R!$GG_)*E.4-KR6)[I?N4'"=S5"#TL1?K?-*A)
PXIR%!'ZM4JOZ$IUPC@'0#E&L-4>N-B;6,*;N'^'S?'L)6)V%9[N:W(!N-(N"E1L2
P&0ZOX'B))I+3IJ=1IISU>4+ZCCY:^ ^M1B]1JM7M]'-<,NG!S<K_!M2)\=8767]#
P5!8&:Z+UI")X5:Q6/SQ2P*3*]'H3>$G::3_KTE%L'OU$(#6@GZ8"^LUI%O+]4F8N
P_@9[HQ>N(MDXGM,<98(VDY+)S.GRIGS*/&8?8,NOL#*PWH)PNN"^;AI',T8G\10@
PKLY%^LLP[,'KO8*E%@+<\TME)J2"7%YZ+V?W%V^%^^0U"WJ%L:@1$(1%<<%5PS]U
PVGNJ)7YFQ#'68ZTH0>?#;AT@4!<.ZG68+1ANJ/%I<(;+/-Q_YL65) :\Y-OBZ>XU
PI#!_47Y<0?9>*^( A$71(A=$Q&G)D1Z1KL4_:66=%9%++8&=73LM$,<."X9,+%:C
P(.J8>'5CP;4O4CXX5RB52G%/)K@,O&V;].6\3\]ZT; SU!):SS,^2!XKEEEY8 *:
PURWOIGNN=*Z)Z[<E^XA-/Y&Z^* :QY:WDF:O&DIFGHBXYWZ&(@_O"X46 @Z-<3].
P_ZZJQ5+B5?? > M9K MR^F'.. V COVRB&$!H0Y(>@PP''6.,,/B^BY=0](*V1E6
P] < \SFBG]:Z+]>K#E09F. +H \"!;BW#S(BH9R\Q_5);MWZH;14\:&)'JSSL (G
P#@G'UX+.--774T;/,<<9FDB1L! ?7TX&/4J.T/O-2J>6L[1)77@!]-41-A"I#'JN
PIY!2U2<YIMO=@)&#+I20^?$N6UJ9-J!>&&(O_9"P5!6SC$>S7_>!:T1+=C%9<?"7
P8$&V#O!:A#, -$;T(7L)0IE1?=%[8I\(ZG=/=E9<JZ'B@Q%Q4\%.84HUHG\Z-9\K
P=?*=V$\4(E Z$;UIK4HOWE6 FCY.B*BV+NHA<,;LI[#A1X;&OEV'.P@-;W3\"_"S
PMP!7@W/B[*M#[*4RG:@*'=C ;"GJIEJGLJ8-+L1)3'FY$ .AU9:DT;XO3_V'X,B(
PB'KOQ6L3; +3(VVPM)-?2Q%Z]8"+TJ'B"4=^*(41=E5D_04@ ^UVT+Z/$<GT3NFS
PN<=X'NOP346Z87D*A27W<2W'0+W:K)#^@QK5<3?!@FJ1=BB+66-K9:SYTS1]M<[P
P^ ^3O0#1"-D"-^?%^8:J^FJ,=31&_*!@U1\D-4!*&_,,U2H:#0[(Y*VH LT%!5AJ
PO',W-9JITF&O5=(9G=FY)I  !I<[U]<,LZ@2:6I*V@L^S1[7K9V\%[6ZE:0NG5*9
P=JU.H;['Z MJL+_1_Q6NST.G\K)S.Z&DV9PN43O:E]3H4%FF+C!57*-&;.+906UR
PC+4* H0#Z0/Z^S?T)/U>7K%-Q2,DK 4+A65OS=@3/ X6Q>:KK+K]+8%L6$;'@PA-
P>KIK>)B3$K4N7X+WQ$$0E>3K</:'&E$&38J5^"!Y:LC%>2%E[WW%KEA:#=%DA]6:
P7G-[G#MIPY1$&,N]2IU@U^H7XT]_Q9U=/3^ 96Q_&N9O)9L1Y17:>A5R891G%Y0Q
P@=TOHWYP:D./RHY,%1^L?@H'+Y;O$'PX\@<+IWB*RYD%3U^(% ^:K@%#62^M-#X5
P[<WN8??/AN?K :(YL@Z[;MCPZO&/-LRZ3#'Y'8MLS5G6,Z_L<,8G?A/_=%G3OH5A
PAI<T2"9ID&,D;YAFO52;ZY4XJQ C@=W3VTA%"^E Z9 \:D6;MHI%\WSH!8,3M0BL
PQ29PDG4XG;0A*?L2D"*QS@%LY!\]..1&YP>&J)C2,@;"DDN @KQ6EJ!#U&U #804
PN/OI'^%%-@%DXXSR61)6_0V 9?)#OZ6]#C<TBI9WO6"*B!@X>)@53'Z3'W>B.;JE
P?+4-:3X?#33&J08B+0=AV#X&TL[;B*Q*;)5K4HWN_8\8_+&[:)?T#O2H/3,AG&Q>
P.K"%V0-/=I7?GO-5<^MI>K5$J!O+R;;=DS_IC3O?<OA4F>0BET@#_1OWO>7PG'D(
P_(8Z;-S*G&J'=L*C/<Z=R4>*P>IL?Q8'C^4R1+80*#VX<!)6VQ5JO^3;N[)V4-B1
P8NB#U#3^J ]<2E'/R6G[+;PR9<7QV)OC<J6:EB8Q.IA':UQ?K[">0T56H@,>VWWT
P[($%G \!6Z'&BES;5OIU$E 63*R<W99O1:N)&PPR5B./ B%\C=^T?SC 6Q?YXZBD
P>(_B'+Q89;5!$55FW"5_3GI#60 6;@!R*:VN_>IL=;0,.<8_@TK [DS?15(ATPFV
P:G\Y],[5;,Q)MZKEV72)B(@,E;*X*V4[JOYB<D1L!P_.=MAPQ?LX1$B'C4QT.B<X
PNP",!)T+U;:<[*P5>C%[#N ]=JWMGK@K5K] G&4R=XF)J7-4B[3,=61 ,5H0 8,A
P![Z\5F3M0-'IQ.+EX;W4UF-;JD?] ^&AU9Q4Z5@YX(BI&8P.^K6RDZB/%?#+/*D1
P:XZE@_#A5Y4JX&1%W)QB__FD ^AFPXPEP"XB-Y=<5T=@*%/(1Y+UM<_$X_T!'F43
PP!43A[9)\SY%,X=(PRUX,O'\X..Z?X?&8)*^GX*7&6M _K312S)^D&#JX/DUG2[S
P)Z8HPC_I^^.OK""0%7E;%3BTO%>=YO<A2#MJ3R[3IMB_#U1MXPY5;#%G^+/)=I5 
PW&OFY]C2"8IVY=KX=B/%5X(NA-1VMH4I7"2B5%JEN++<63VQ68!YY.TL898BN""(
P9BRP!/UM,S"+ZLF2GH>M*KLV5OFJ+N9G\6=3GH1YE\(CN)(UC//3K&7CZ55O27Z(
PQ&C4(^"%@3@DY@G&"2E!J.=\^U?R[ #2K03OB_3!1IAH#OYI!;P.,E<F^F>,"Z>=
PB.[<&=,1LN_:'";J6-)/-CNE"TBK&[3UA "H8<>,>_")@,U"4!I'A>+H-,2E?.F^
PZD%IW!'_6\ #B8MRBFWOAAGK&*$/44]@'3"+@[A.I,88PYKBK1LQ$A$"05-<FR25
POEE)AZ^HC 0; @UC^!-V7J=5)QYGE:"IGLR(>FYU)&QW^XCH]A/2>WY7M/I>2(;#
PQ$#TVFZ4-(.A0QT$GH/JQCJM;+(T.-_K>TSBL*E+$_FTJ+<Q,WS ^U+@.5H[GZ,H
PPRNQ\,#7[&01X6*F FV)J##O2!@\D(13L,]S\)1U2(E%37)RQ2[]VH)[T/:;3"*[
P5Q\#%7]6\3?"MR^&K\LAA%T/7<-H=N8K]Y*-ZTD;8;C,TW\-#5M%*/FL/869\C!7
P(G^NQH89+TVP%_4V6,_38RI$FI?M:U(@7;,/=5SKZ!4X&9($0N-FU7<TJ?HBOG1T
P,NI<WIS:5$Y?@5I9>1:(U.&!@F"L0MQFI0#F2P2RDC <?*88*K0U/[/C']ZU'S<-
P%K )O  +8EWY3([Q>)V^IK4-K:>P5):94/&HX$:K1E]WI"D)5GM[R[3/7DU0QPX-
PE-$:-H_7?;>.7PP"&K,-=$M-)C&*)NCE(:"X:()HD2@-Q7!%O["??=N('UTW1@IB
P"FGP<*26-299[9E8%9D_?[R"6$D-- KT?+>T3)S4+\H&.'XP"P^"52#E!:*3I0)/
P'U$/D,/6]'8CH-G]%X@@B,@:RV7Y987L?/2 %7=C?JQ8LW=O\S@DS*:&?U>-PJKU
PN-#50.F7X(3;40,Q52H&'7-28XG%YY_7Y+@_O8 H_YIURP0O&:UQ'Y_]A(MU^W6H
P_(KDN0E(SCR?U7D>HI*3D0DNCA9L")3QG(;!26!K0>NU6JTQQOU0H0I?8#<0=9-B
P<!I^+-D)W<E8WU:U3$V\U<#4$XI'%D2[.QUH:AE3-$IB_9KGGDGK'>:%[W[C"6/:
PP"I)GI*/H,B,OL0E>!F1RM71T>M,R<6: V*+&;%QCSIXET"[)D<KI6S@U+_%CXJO
PAK*S<89#!I\2P@C#F^?X<<_*5*FJ )=JRX@B.$$C >:$G>^>6BIWX)>/H$U3?*K0
PQH3>H\R< Y\:F0,OOPHR1OM*)*2.R/=^B8I$=W%B1E9FB'^W)2EB#[&&Q<3F""OU
PZ4#>K4S::B':&UGPHKJR8=RWK6*TT;'BHD)QI0?N3YZ,<-9<)(#+1%.B(W<FD:? 
P0!KFIRY?7F2D=L UZKG\EFL_)2KBIW^AP,40,@4^R!A0I[J4N.&>]XO[>\HJ+\B_
P'#JR(W^A_GN5':J9\WV6O+ 3+<S^HX9&)_'$%]I%NY<XS,"D5S?ZR@C;\C_-FG,U
PX6\'#@'7@MKNEJ>OJBRO9@A#''CB(BAKL6-6 ?I(+IZ+$MQ5N9(#BL!^^QPRS%6Y
P[V1U;$QGN@Y?_^2OCL XG$E@+71B1?M()!W@Z%XUG$^+,6S(V*\.A,@0P18.#PNA
P\$+):W%W8PYT>DLI?5?GM$9'UL^$D3W'_3;RG'^=6GY'3*QOR2_-IPT26TV;A$.!
P%H/]U61@L!]8UZP6<K3#AURP7-HC3)T/H+SK=9()2\:RJQ=6 ?P]I7A^Q2XQ]D5G
PP@5%&!S1ZB*KZ$:D:T4]%;\54$CC_&T.@(&&0UP&<(1()?&Z!2Y08"K?**5CCJ0M
P!$FW$1?""T:8!)+0H^Y?^I'"CO;=O32#O=MG8.XZ7OE$!C1G: ^_(FA9E/E99MI 
P/U+9H N,DN55''Z0V^$S4^N %7+(2DSD$9+,XA1'\[>9Q)!'8SS/61F&AFJO(BT5
P.MUH,EW*8Y/M<R,E _3Y,?)9N86P9J:!L1RS6V]U8;2 C)I\DRI-8^$948TK1%_+
P1B;6_("%) C4> ="&=_*P).:@,+!'LM.)D@YJ]VPZC8P*2/3RQ>]VV<L<?,(5^6*
P,?2?+ZK)YR!+R>21 &"_K*/6O:]HUYG^C/X_L6K^RF11GPI]>D-/ZVOH]3D=2M\)
P8]3YA-K #=))B#N:9[1D]>C03G'W+)<665=)2=3.<Y(HB;#!?_I'!TA]N1[JCOL^
PX35-B?(U:"5D)!#AD1Y[#LUH]'(!^S]CH\BYU/XUXK&=_7=Z998 ME6\45^-/ IS
PM%S4? RV#?7Z!.)T^?BB0]EBR;R4H2T9I4CE,.AB<C:I"!6^#UD2 *&&.@1C>AAI
P1H\]A:E("(6O'%1VR@$[ ^1 GA9)1,B^#%!HX$"L1TTAORVB*+JE+PHX[6*V 29:
P%RR-5INUG><@WNI9103;Z>, 5]9*&GYU/MV2@I3)6DZD8RVZ<AZ;0?,?7OO_OH0P
P[2*5*KW?W2^]8A8&>LXK@O]63R<E<SEW%8%$=@&$B:'4+R_<\]N"(AL#N';+ Z'8
PZ/:NJ-YRX:I 0J B4\#?O?]ATKG8TT5:,XF6XD/PG0O0:B7FN-HUL3KJ7S17"OJA
P&!%#C<$>?&KJ^")&!3<IY43O\#4MI#DB40@EL'OQ J0YAW"'&+5%W0<[U/1)_1SS
P<K8B#2=12M'URSK%@@H72@@&L_44ES, 'H_*W(6/[ N=IW4OANS(Q"@Z+:YA7%ZG
PB=(\'C-(X_T-U?*Z>_(;NT-XI13?6@NG3M]\KF*N&))!:YC9_G]X:M.L<_S*COF+
PY?(KD$AHVP"BI\D>V)D$Z% 5C*V P547J?3/<BN&S)([P;NZQH]L]=+=(1&W=-&L
P]%L.XNRQAWYVK[U3UD2P-6VW:DC'6?<&[#!<!0X@\QI\KGI4P*:0'>](L1TB"HN1
PCMS,L'@G*JBPL?+K)W!!S-R_ 9'XM'P:/*OY*Y7X1JM*QK:_LLN_D9%5UHFDA"7V
P;$,PM$ELZ2X#7;62:)'Z25S2SN='H!TZM;&^GZRO;20Y8[8AYOO5[>C5:MAJ!8S8
P&FDECIN)$<O1J[R:P3M&-(QG#TAEO]PJ1&WCJIJ>P<&R?VT1E=3( &1&'6RZAC<%
PCJ2L$T8_=NG@?QGH[FT []WN,&6RS#&U_7F$0\._<O5U=CZ>Z?XCOK*ASD%-<H#]
PT9F*Z[FW/RP6H_WB-"*N]8NT\5E-Y"N8YY,+[PZ,=DOJ:3[>7S4BSNRYY+)4L0_K
PHD@HX2+XF09"K1AT9;P]U1$,F_GJ]T ;QW]D_Y^(F1M.^[4P;)P+R=H1DN=I. L\
PZ=JTQWI_XD*);![>@> 7+%R_V)%\C#Q,:'(C1]@V]HU[1-G'<_RX1;31'%X+_!B>
P6@XGP=XQ"OV!DZN:9:L)<QRP;T!7-0\28:Y4^1Q):D$*CW^URR6OEL4BF"]TK/DQ
PK08O,"#).?[;5(R!BF&9_/IB?^>7_"L;\.MVT]W)<*U^KZ8)@;*1_ESFI>V/2J<3
P8>*SQ?!O"XG(U]*!EC B1#&]JES,LS4NJJL#*'F/!\YZG<WFJ79\(XM=4;>P))QC
PCP&R#>Y"='%%9LE7!?S7D$.I1-"IAZT!FCMVH=Y<+>H[!I^)1A"(2Y;Y&(5-0<]R
PW=@";-'V&_$Y1D$A@CS1,5#\@K9'FI1%3<32X]K(I![!"*33/")+R!$<+.G$2.7]
PU+R &.1'5[VZ=4&;\<(KR[FC<A8(LX\W250/O76W$++14R/A -*-?RKLZ93?4[\#
PGRH. #Z0L+QEA5-P6DO@7!['7D%PND_(O5A\CVB_@^[M=6HPJ6=Q_0,,Z)Q2:SAG
PLB:IJ+1G8S,9?9(4Y2HXL+ )HMGRO#)K- PCHQZM07%4725R(D$"(?2D)'<=RP?8
P,&1=@%1/$"0XQ]JI-E=0P(FQ--6 5(:*/D0*LCN[=:@P1T71=GI]Y*2U3KE]'PZE
PDR#BET8$<Q&D84+^&U8*(&H_>4RRI,Z4!'S?]'7IFNS:0 3^$H@51'S? SS#-Z9]
PMYS5_+KJ[MY,[WBE<K/-:=C_6Q8."E::3(XINZ%J!6Y \V4!^P66*Q!K<*2EOA_@
P\)#*"TJSW!"X$T)1I9P@2)#/I'P#C,X@$16J."GSU$DS]:"PZ0H07=1.>R[QFV6U
P0:-UQ$I!1]UE$_EG+.K$3HLV7N<UAX7"=BDO.3J"9;PB2Q<Y,5$B,?#L(TD0DHUB
P<BITD8-\C@_&<<J43/^P$&I</?+""0-:)<@QUXO<1E6/R.G:O&XQ8EK>H[M<.1=L
P"J@LG^147F+E*^I\R!Q/P<2_X?DD^,IHKMX<'=FA0VPG/';M^VX;F'V7J>AW9H98
P>R!UC%:>3+05?3VUF0!_4 :(D]>Q/0<O_RQ>":T^ )J S:HM@E<>3> *'@O,2O4?
P>2?O\LSXFKOO=W+3H"Y**-Z4!0MK3]=]L&S"U"'+LX!!?LRDOG+@_PVK++B%)9?'
PQ]0RPFFP3*^D!*B+>*6X]D+?_!Z04XH)8/,YZ7'+3#H Y%4_PAL])2/^P"7"\\RQ
P[[!*)L^@51'NVY5EYTZP\>&\A.\)8DG*JNB WK;;T#G"^3NEOV4,=*V8<4Z4(P:=
PY%6+"%N:PL0 HF[T?$&5,:[OQR#9A.I!IG6M1$]AE(0!QV+ZJE.%HMAR6&=E0/K<
P"]SU.)AVC8Q#*\I6T!*>D:8E>*Z/>L0U =KX639=+,&T4ZYYSSFRTI$G X[=TH09
PA3;0*Y7I5,'/N'K19X>,Z&6V%X;W4\DMF6US:]GZ\Z=1[HM.ND9/7YJ@CZ>1)%"_
P'GYB^@076UN/Y42/-A2S!GK=2#5%,WV7Y@*17IL9A PND#Q?271N(_XZV2)&^55[
PZL+X.@KM-+B;$>*VG0*I!SB%"W+TX"OT-#H  4'$];GW\PCW.>.S509[7:)G0]/;
P!;N"UUGL8X5+1Q,)\$/,6814#+9&3_,1:>I3G*BA]'5QO-Z[F.6;_UY[$!C/37.U
P)BH^WG0^8$MN6=1F0B+@E9_F"47CD,,D U?FM"[]XP92FOT2D FK]QCYQX.WSP_Q
P68.G@PMDP,F+<NVD-&_Z(Q3%EI@J&1>TIOA8#V%H!4I/"/GV'C0^\]?ZR))&$F=Z
P7]D,8!Y)T2,M38/!ZJ*(PA)4WZ^_^HP?AN1SXYY&A3"X2CN\;.HB>\HFHNX7"E6N
PL^WOX9Q3&<VE4(S)1CD>C@%@A(%8R4.VL2%A?GG0!68P# :R1Y7/%;%(P=_PG#,A
P++\\$NYVG._7B?6E[OIK^TZ54SSR2SAW<DI0OI&.N=&1/RCCJHW/W?-XP7I(8A-^
P$\(G8=X+$F ,TU<1U 5D+W=$N? 0B8B!Z)UP0"10'Y0THVQ0'-V"RSZ+>7Q;NF7,
P$T%17L.^1B'+,7N6Z]]BY(K.#]?].F6!<PF7?>;Z_(W$S@;D=EBL;ZMVY'4H0]L.
P;_T[3JMO#/SX0T][Y<\J8T2>N%-)S.LVEC;>$L*U4T'D$52U<7(C!0OC+U?%:LV3
PZ'SYVTD5L..?&\TIZ@42Z%9.F<E6I\F-]6U%&.JM?RZU8E641\EY"@^AS/S8H>W)
P-$%^$S<O)%O2C)NVHO?.8FBCF.,2Y'U 0X[U$,[N$- ;8Y"8)2T./RIQQT0Q:%S)
PK"-)#$H-6Z(#= V>VPHB_U*8\LGP>DE[C 32=;D!JI$G#Q?JGDLJI>6L9-W?I *5
P'KA<A>RKFA0;H@^CE=E$1D:562*,50><(@+LPPPRH#,M",>R &7-U5@+?%VAJ*6]
P:'G"X4['8WG3_B(^'6H8CF6'03:999I[L#ADH:T&GAU+1$;C8@>4<E%=O6.M1\A^
PM$N/5@BLJ(]!EG>NB^=- &?;H=TT%T$1F[=X00-LL\)WVP\4TBV;D&V@;#:7I4(5
P,L.^:+=7%B?T/!>>5<'X+O&TXK%#Z4%,/SR%[(>2#2)4 W9Q/(XU/JR@4/UU#(\%
P=^",M*/'6"*P::-$5>PBP,ZO5C*<DZ/Z<]5HE:97( <!RV]1=FSV%&ZUH+LH&ER1
PHYEHE5V<]WAKQ62PN)3S")KU1)O%J&7$JK"*^!AP2365K:%5MH?9)?31?3Q4E.E 
PYTVG^-C??"I&._(/OHL0)^-OP#!EO!1*^-FQ_D")P&KN$HGGESX*&ADAC##AZ0_F
PE(W?GHT&+=M9K@&G;=(W%</V5BTD6N-6$>G_)CC*5MT9JT\/C/[L)1-SP+<P(OFH
PX+.]3%6F%$(8E$=D:+"K(ZJ&QQ(#.6>^?R5/&0ZXLE<6]7II!;BEC=Y\^*(" V Q
P^=,;PY:,0JW3O)4?//MNV\[M-A#-9"H(^&N-0:H&FU@%1>7DPL$LEOYY2/IW1VOJ
P-P^.* #YEX[L=6N=/:A17PS>>1=9'(('-?4XYIK1@8@$EB>B)+M>Y'%+=!O$"=*T
P&=Y>(XB;#*U72+/U6W95C[8M3L?&2-PY.QB]FOIB5LHW"GW=L- \G+[A5,L0PS2$
PN&,VAOAW%2:\)[-Y@KA3ND\IW]S>, V!#^JY$427:&J?_@-B;!YQX2RJW2 6/,I@
P\1!XG@,9HN-29BR:G:8.(SA.0WS[;1)=S^ /V,$3GO$;NF[F<I\ZS2E<MP&$?Z1S
P=F-!V54+CL.+%LB+3%4A.YN(?O--Q^%H%V/IXQA"G\=TOT=-C5W,K1W'W;/PDGSF
P:5Q:N#3K+A!]QXLF0@;;[!*0V<A1)O:X(Z.7[^O9>MQ?7/.V8)1 RDLEMCU0OW;\
PBB:H RA DCQ1R%&2F:).EDCJ@ED1X\6-YW) 91X(%JJTJ.JB$+R1P&M-X,]SR1'U
P!)$&;K@'HI<88* U=F/[N^1&$AVN.-2&^,[^NL160K)>P=1-, 9FS&]17C*5%>^]
P8W?+%/EB'G)E?Q+EP )J;YHB+%>TD_"8QT7N(#X!JF.BQ"TZTOLF>M6E#6*E7FIG
PC)X-0@.,@4+$;L!A4C1^T'=7MU2"+*E!,0%D!"%$YZ+V8]6:,S9Z'0_P]J+M=_<]
P+L/-EK@M*SX]Y#.MR<3\DV36C4?? E4X]]4>JQ+G"ZW0)*?I%07^X6M15=[W#*(C
PRE_[VPO^85*:NO"6C68P7IOQYD47C(<1;C3B&3P)Q KB$:RB9,M;<L#';E)ZY4N&
PV?B1YS'0:YC':W[ICB-#X6OH0  8]F"!V79&6'A<4K'$.$#TO7MP[*=$B1ZH&]KC
P$XU5(,4 ::_-=8WFN3)'F1P(31.EZ7!B9"(%.I_+W*2Z<K?XE#32+D>J-^X2V0;3
P'&&GH=<$D7FXD6XZ. 1*++_:PPK.K(B4JO@5'Z+U$-87+ +REI@"8&7J AG#B?83
PX4PF@L6O(RRAD[2F2L?7\9-1%L,$'6H;$;Z]QB6B %4V [%V IVM*?Z;Y@MA5*;5
P5#?V94>^+6+_-2KZ.A045>SCH.P67$.9V2HCBFB<:16@)PU4W]=N+N_B<-K[0),9
PHNV'.;:Q=WIIP19Y_MB,W=$UJ0*L)/_.A_T[9:"])QH$6LF Z1"[F[@14F+*LGZ'
P,*&M*9K/A#-PS.Z!M<U2GSHT*WW\QT<Q)U/B2%1!^DU<8$<ZM*+WW3/N0)ET4&C-
PLD;IAMD\A:NZ?RP)C.KNVHPU0DCN!R5R]_?Q_2$+@-,JN\,1-#V?F][J?XPSPSI:
P][_)9\U@1M&[=Z,O?&34*8PFH)%<U,O>1+<>E.-I'6/A<2_CXR59*+K]D*F5H"U2
PTP'YB)D5=GM:<?Z9UY=T,.:I2*,+4QT755,/L]\E'"@69M]G6TK@P'+#Z=6=Y)H2
P7->NG3B&0#N2605[9'@Y\%TI^%DCT+Z-:3[ :6XZY]V/QTG8MROO^3P;Y9Q9*\%V
P( T<LU8V>I2U/"FI_TW 6K<7A[#&DJHTUDY@.DA2!:)E1-"/@Y>:R\<<U:Y6G3D2
PVQNA]I^QFO;NVQ2L$B@#1!_DZN9<%S^!E'?VW/BN^OO(07BMT$9 ,JVE V^M:Y=:
P69K];7!Y-E1&^?6!/(*L8?'+*=)0ND1'J<I)+LOZF$.&@W^S11)QD_MGJ<(?V]O@
P_H>+PS^V+\<K*T#NAB,'/@EL%D?/A!.N[>H)%^]Y)]KDQV_;;%'[,[,J1VL[L5OA
PNJ< 9ZW;7+7Z]]7'2:'_E;;41=@OK.H0GRDR.J*QQ&;HZ=/4";*I5XJ!Y@E'?SXN
PAE4V1U$?][^NJ^FGJH)J1),0\.O#*[Z*H#D6V16 >!DRBF5=I+..D_';#FPWU$/7
P;H>(?-06G())8B/>*M%W.#V?*'<F27G/)YG3-_Z&2?& VCB>E(G#'?8&;(>,Q-)G
P ()C<%?DO6M*CO&=3#.4N_)'%#KLT8=PX]_K")4OKRJM1%S(7&*(F($T[,U(LT"*
P-(;]$-V?C:Y+O<HA(O'VNI*,4P!J-K=@(<(4C5""4+TM,=]:M*)72Z("'?HLQKCR
P)/R?F2[C.'*/9?H<-/Q]45(!(WD>SSMP_?)4/,7TK%XH?^YH0 P90:LBCX2#:@Z=
P)2'NI0!4$#U+0:WLEFUH,&+W#0MS/?[;<H61$:)QSR[[[5K4':$UMG0BH*R#R++Z
P/:N5L4-*\39ASYI4@J2-ZZ*EME4?DG8R#K=V$^^37HYG0?A$5MYDGBBSB1];C$4%
PV6?IX],'L1U1#C-CX)M)?D#L!&2'.\FY,_<Y=;:]>A7M&8I:VT>M%VVRBZ:3+E18
P55,C.L7'Q=5C5?P?MF,,R!#U)NL!JB[0H?+?HA\S,. W'5@XZBKJ>;?6D5MYW KX
P_Y2];QS^00PH?K(NW4]/X(#.!:2@5J%D2:I4;?%/MA3,5I:KEEAVA.S*&,#9OVI,
P IMB%R8<5IK0D!\M]C=7ZN=^G*4$##M&@ !"7B?"$/;^@%-L+C[/H?U5"K<D[SSD
P,O\XA<<QUY5TT^4[>RW!I(J!6:>B1R3<"8AT->WY_.4JN$_@9GL&@E$L$_H^609+
P>FHHD.ZLS"ZJB7M?_8@? =LV&GD[UCJP>@"[K7,/_A@:?!9S2[KF/]R26"U*-ZG4
PX8^3&DJPU$? 0XH>_X'9]@A(%3?GW/JL?8D_D)# R:L^BT-/.N WQS"P.!DZ2)J4
P:'WB='&_XG3$[;_,^GUHA+#Y@)HAGOL9Z=N]OJBI95](LJK#W[!,3_Z<N$\$ .$G
P!3 [=EZ%&5L*BT8![\[0/.\B7(AT8U?5LGZI*7:]*;4*'$H?' [49Q9B2[S>Q4P-
PP$RJ@1!FI6W\N8(YS[I4'TWM"-=]Q_RHC ]<S:9?J1)D$<\>S:0:ON(RIV$=G!+@
P':3.>X7+4!)2[H0:D4XT=MJ$J2[17A.T=:_! G.&#"FPRJ?_*"L6ODI.-GJV-7WH
PKS[9%:6*,!TNBZ_+;*(T9H! <N"Q;64P1@@.B!HN9]&4,S5WVP.O[[CC3<-Y9GJO
P2;$\+] (V>K1T7_0XG!=_2(C2Q?ZS@ZCVD8#:+J9EN)DX<C77L0> [/7(0]FTV3&
PM* ;V30/" GVK6<:SQ\/'UDHG5-A1'NC_X>6HFQ+-EQ=JRMO3$E;,#IZ4MRDA>37
P3$>0(;/D;^&TP>L.)?$E4M0&6^% Z7W')@ML9ZE^"+S]T-D0.V"?5[?!,U64%NA%
PR^HL@4-W4'&'D:%NE[O!!"_XJXKL*PT4:^0O]<C7B*8V+_E-B##J!N82(QT],/06
P_C<!XI0_<1S ;?(LJ#$-5OINOU.RS+0WMF(W6CI.,4D(_$U_TE@[^S89F,Q1Q49-
P]36]@<X!\%"7.FTC!4?%'6?"(] ?\_CX.9(+ 9I6?4DW@3 9N8/></J4(T?SB@<;
P"$L!E'26=PU_[]11^2O?4#(CZZ'8YTTB]!=?2'9)J%X6 .#OJ**+G$JA(D]HAYH(
P&/]U)CT$G0U(W>E88LD#5,(F+.!O=O?EU2(!'KZI89HO/ALE+^^8EH5&3 9"8Q ]
PZ$F8>WKZLGZ!*$"K)2F7^4Z2Q?_GE&A2VY/;\P@'R&H18^9X(&UV-4H\/:B3T9. 
P@&<Z*&BN5$>H.:Q.OH2?AD&1AK]M!P@?>0:MW"C8%;)JZP;"I)])R89AIN@"7$B]
P]-D% J^I&&37@RVLF[H8/83U.ZN!DJY7+,9W:43ZOQ80,3$S^@KW4%CG'&&_;O51
PO_=?Z(L0REONVGYF4S4XJ!-.YB QNN*BH91VJB=4]0$;' 4O,C.5&V#%9;.9VL&X
P   U*9QA\X:"M2ZX2OMO^WGWP\/HF5"3S(G$J4K-4=Z2YX+!6A*2OSJ#+%<^!X[2
PL,BY]36D& Q\O*64.!+ '")YL*7'&2N $6^2&?BS<=;WGWB&(CQ]:^<6P@6[LA 9
PQ5NO_65I"6*UZN-M#@O3BYO</(5^Y2*7RQ81B\-96WE92Y/X$M,[::603ZMX7T;>
PZ\^VS*Q^B&$>O3/&AHV\U!I'P82@-*Z7^@NMH(OLB?R'2NMFJ-5]AJJS=$G(S9W9
P%KH0*8YL3=?>[D< 0WJ4K7+MC)W/B")P/< <LN( S5U&B> /P"BZ.<F_]3%R.H@?
PE6C:S"1JF=7AW]YI4LDA[D)0#2,4<,'JU0/<_+(!25>*->ET@OE]US#V9'WO7DG)
P23R?=^T*'^U3:@:7]G8WYV0Y#UWWT&32I*$%\]VW]9S_$R)D,:LEZ,A09B?#FMKE
P+DR/HOK5A_@)CTA$P*!=-225C'_L2!F*X%ANV>1*(_Z1E78?"]>P5;X:U[89WYTW
PTOJ9)?^25@$N;RL0/GP9GK0/R.+6^N1'RM8AKLOU<8<*7]>KR//A 8^*S6<1C3/A
PKH+%YIWZ,(7KL.9@? QY-HYY$//.S]_Z>AXRH"%ZO.W?-(MNO#>C4;OTB5P=#5.1
P<#C0T3RAB/3=?FS#_00S61QOJ9?O2O3(_HFMY<^$SP"I+P\<QC (&#%0]9]'FKM[
PTI36.DIF(5(X=G&ACD6LTAN_WVGPBKX?VJ&E VGY*TA\Z[X,W[2MEY-E&"C]T@] 
P]P,\X^=2R<QW[JULZ*/,,2ADHC_;RWDR>ZBC8UWH-I@_":<6*(B\IIJ=G1R:I[=%
PH<X"<PK/=Y*EUEA%%O58;UM&C?L[VT7W'U0LV(]9%2_=:[^%Q@#KNAOTS,*K,BF_
P!D5A(SN6=61 P-&I>VJ:P?Q0ZGP4_FY.-/N%2#Q#[*&C!I%3Q>V1+K[,]M\BW;9N
P5.G?\620_)Q"6'I*U5%UY)4281-QJ+:;BRX/!?M$ X/7'4 K0FU\%264@V,=%HPR
P$84JISN%(G6C;YT6TZ$W^(3 87 OZ_*)K%'TW2,)'YFPU1G'-R[HUR0N9,(?QZ">
P!X CTZ'R7I9[IRK"5LTB5A]C AG\H$%]D:\!I5THN.DZ(U8-F,C(F,3S'!L;J//U
P%*DC,'0W3[<0N4X%*UQB"\Y&M4M2[SG+?,C:_M\NB3&EKI@M/18I-N D.A59<1^'
PV(VL<5J]:L=O(2OIQR6AL5S(/L5\RF ;^ZL,V)_<%#J=-\UGX6RS0:F>)R%V>2AW
PA5^M3ZZ;-8W:,KUX.L51HQUD?9Q%FM6!-RA$N^YP+\BOO[5-<50VU@&]2(5MSH;(
PRMY&W_L?P>SD<<$QVP9AIG85?EYOT*5N(#I1$MN];'S7KP/^=*$YGBA]'[4E&<.7
PWV-) \N"'@VXD/LHFIYKH'48,6>] F6EP)E P+,FC;_KNYX"-)@YN!GUDV3*-G4S
PZ8'UN79"=;-T7Z(+<2,H=U03*.^Z(T)\6 ?3[[9JH\A4C,2>1H#3.8J[TD"L&3N]
P+J^%P63C<,Q6KQS9SWWG.[A4=*?65%9<LLUTJY8<%FUSO*4CN]G!I.+X-Q3$@/$E
P2#$V%9ESR\]*T8=H3&K&73*_O^:U(H,^ZEW6GQG(<2*YT#!2IUZ4J-1@X(E\_$*%
PW\XX4Q=_6/$QWI;O#=L7WR9' 3"AB&YG8_O77O\=JYO+J)2<7,V#! JX$FN;IHQ"
P(4\3 &[B6)H$PO'8D53](A2>M=V&8#V'N(U9A2+5R[MOQC#[GO//#:SO&55*HS(P
P@KC+.6-?*J@/;U#4HX'D(2D=M8@R6CGO^C.T<CFY_*F:>BIXWP!HYH\:KFAZ$^]_
PY>1ETP!"96YMX;3(J#QR& XC2BMA<,N%NV$B(Z);OD2'"@"8">]LY: IV37P@"G:
P;AA?7/ATZ!9_]PYLDB"BQ3B<)-S'B92 U[.@ _B#DW?4JW=TLDL7ZB>SS U<R40^
PT08W\>*YT%[@BRMWN4[EH) M.]H,J%42<OLK#H3I^00RZ2PW!=2(W#CY1RYO#H;3
PJ!T-]*L=2I%L I5.NYBZ<-M#P)G0!VN_6_4F@J8!O5UW1LL!SANIKR-D$?(RSM=;
P//:\+4VQ/GOMUWK2(.)39EMX*\(C)MTFV-^@Y<LW.@F&A[Q1U"]\M@S#7A8SO\#5
P;-G7)1+DPE1*#4T,IMJ<K;7W/\K/A6K:$PP6^$D:HAZ+!89[UVK-;794_F5TA(,H
PQ"J+!0>R=,5%C>^E+LP("PKS%2Y^\-698)'!PJ^VR__AC:+U*9OR22<DO>D-3ZJP
PC''H+'R?RWQRKK3S!S=D4/.2]U)$N0:/M'5:*9?.H^0%EW_N%Y?&B">7A!O/U-#V
PEM^GB+-A>MFU\ULZ:57OE3.RN]YAGP/'OQ0B'PKC:%>I4MJ2A[>9#]7AX3V&1-XL
PG,-A;LZDU>JK=41T%R ]O5#-;[ */57$>;CY+=:&/CSLRF_?&4SS7GZD<E51V@\$
P L8 \,4JMX^I;I.$J4()N_1PMBZA&6VG7,T4P^V57+!7,%QPIG[0;8?:L/FJQUS-
P*R1*]P#/ +44*<7[%4^A4,/A2K].PM24*IKNIJIWL3)+7Y>A;#WUFQ&ZM.JE=A'L
P#?"3V;2F;_$MY.WD!HS5^H;6:'M_4.GYKC@R3]QLSBK_7/!9<*Z8='L?-0G[V2O9
P2M>AWXJ/,9Y89\8XI#0)J?= _P+AX5?JED"P-E@IEJ^I40WV![D-J[M?NXP++YCQ
PZ@K:U]"@DZ=(#QK\LF L(2V$A#]6TJ=+/5>W87>#QAET\)5\0?>!?2:A_>KS?PWV
PX:N&SR,(9EIPLG3:A-NLW/R::W2,DA?,CT.GKUQ-#YZJ>)K X?9^$?9MXC$Q5UA\
PX>S-11]6;*EX"QY'@O,E5* (ZGJ.8*\2"!Q(V/L>%"MX4G:]MH&E+0X!F_2R4@Q#
PMQC05QS[XA31L7HG9':S8&IL-UR41DO?$M2C%3V)GN/#$*>W:P]);C2+SUR3*44J
P6QD-OPN_FO0/*-=ZJ3UJ:PN0B > ;XIJ>9"[5S+.FG+Z4K\*VV0=.IZH)S2L\[F4
P!ID(>J<@3Y45!R$7NOFN!^,+=7*(=M3JF,]]F?*H!=>\*0RWB T3)4V>XA4$T@@D
P^MX4^@1#2-N2P")FIG.[,:MN3LLK-15MEZ(';@W"2';3E<TX"\#\>+Z->161:EY0
PM,\(:P8V&R<&SN"?9Z+Y$NS&6I&,G!!3LD Y*_C(#U;@#I<*3S=B3C[SF +F77.5
P4Q$WN[1B N(&@T:WMF/VTDRE:ZUR:8'D7DZEYKD_!_I)'KQTL VSGR]^\=?$$-QZ
PH8CEH-'$SL!&!AC#"Y2W563P'VSD<R"F]9041M_9.J$K=Y#@SN,D8N@.0/0X\D4O
P6,6Q0RBZ-:D1+7>#D"NN;O+K=+)Y0!?=& X?=< P:)/9;[J;GT9\^6^SA..?XOV]
PCCQA.91XBGHFH3J#=KD:LUS5I*W2_HZH^%?4NC*+2>ZM#P&Q?3U:[U%H46GXP*(5
PK-X:CYRON)1'34UBD3(5[5/%DOK]N9<0MWDQ7K*?<\=F0L0@W4?X\#SJ"C^)JKT%
P AFO*7D\G"5-U[$:_JB><4.5$^P[4U(YW/0W9T<Y@9U*CTHT8:)J!"Q \2/0SB'Y
PK!]K>13+CIGK?7CM<G4+E.:21S1&5F?M'S_4<D2SJ%7TU>I$S&L&G'D-=#38R&[$
P2JGH$6,?$AK2AJ:09;TA1#+^4[0+++:DF^R,!1"A!EQ:,1Z^\K1XM5+<%M!M1[DJ
P\;$M%WY!311A>_"F/N1&T\)PSWSQSPNZ3S"0:, :<"[/EDD3[)I5343NF]^X+CO;
PNIU56%PO5E&-MC<K$2,T<+,,) N$YH/B3^2R)\\U&!/,,W_A_GMW+AH\-W=4:TT@
PL#9[:=6,QT7#AVK5W_$!-'DEVSLGR_?9_?93O0RY&F$,IWNY#B0B#%_A&VO4G]0L
P4U01'J.DJNSV$&,I0J>SKGD,D>GUBX^HZ<MZGX_E))?Z[5&X[$"[S'YE%'Q**&I"
P<@\N/B<"@F$/OA5NSQ>(4G$9Q"X#.H[L-.T[4@;L6C) !>4P'-%!2[/2N( O<(&@
P"*TU +7]@TX0K##H5M;_ ,5(4*$I66W9!&%H",>N@$TM*Z<SI[("Y7.+&#1*[EHL
P71!NGW[8!*$6@<"/$>?>L^%C&5POPM4G=K$0Q#@=Y7DFYM9L("H!_J\_E6$\G$!!
P#F4(;?#"T)N:;>Q'\QKENYKF&.\?L"[2XCP=V3!]6WV&!J&+P?C_P=6&*6]7?;:;
PI0?42&W142>+1#TZPF>]F,>/?6$])HI8G*DF)AF'6XO5/8OFH\SM\!D5)'@$W%-@
PV99"M_I6OP=^K$%6Y8]\WB7<-ML:6>^,UU\O)R<92"%G*M$+@;J5@$#MA $:^Q1-
P'PU\_K_,S@,+];GM1?/;>[N^G7G>8M*:W=HB+(K0XKIH8)R7JE.F 4IVEAS8X@]4
P-K#YH[P)S4<I%V//"8[=B!0E0G)4<7X]7 4VKE>W+=KJ)K!\+6O&XV<^/^:3)%/:
P_^[T$JN^6HV,?T7^SMQ\TZ 3(4*\TC5,8EF?1P,_W]^\$ X^^@B@H8E:92_MX*,/
PL]4_A$2*_<#-O")--O7_&ASZO2C BBMEB]%P(T<B6S<R.W[580[A:T \Z5EK:7B(
P&[Q!(^3 CZVS@]_SOT02!"+K*7G'VN!U5D;.AI4;!?$$"_V3S"&CM[6@&E39(99V
P_,4G;4RI*5V(OI,6&*/L]+K.1)&B#C,YA@)G"'"PSX)>NBW;><U0JDSN>8'<!.%.
P=%_M[\_DJVTTG N:$)BJ(#\"%BGA@^_SC!,L:E:N@<B7J;1FUV>BYQ*:%*@7_S?F
P>COG(_GW'GI?OK^;?W:1X$6&QO4U@I5J)QFV9M[4MTNM+OR5$@\PH5NE!>0WO%TH
PE$"Y:ZRP43<"P7I7983XKQF[,_&JI96Z#5$-Z$W338'+A35[5 +"3KA3D2'$,G;<
P7Y[TL"XK:5RN0M.4CPFVNFNS/47R>&<\,0=T*[F]P%] B#==5<LRT)L:47H]D8D/
P]1HV.<@W #NK:$I#+J8 J<>#7:A?0^WB-)"(5R'"7_'MY3RQ:)E$Q\]L%_%(17G$
PVE(X7<VFL]UB:A_2WJ4-SM\R(+3KZR/P9K>DF*WJP[E6O-TO,6*NM.^FWVT,=4B*
PEB<X4Z\*KCX$7O.?V$VR@C<S<+QEOAIA#^9V@G)K?$R&P7@\F_ZYXOOF'>H9JJ5K
PIM</RH/?!S;6T?QR@-@R)CYHZQE?MC''V[$X$IN5@_#?PR Z,?!!GB:49500Y_5C
P-63UHE2+4[?MZD!@#*"CMT+U4-R=F/Q$7+VQ3Q=M/O/>,LSQ3UZA*P_&60\R42!&
P+%BTGM#^I"5;/+MS]4%J[]R N5,/VLKF=_JQ*71 ?U<S@JQQX&L HO'RA7,%8 &J
PB="9BG$2?=*F+,>#4GEF.@$+^T.#84B6S!,U;FK+3''[0V[4[P"+FJ/A4,;R%.L[
P#Q/DAI)I2137FA7@,4;TI(?7O@WJR2GM"<%GZ1.!Y\)...H\*GMW-(&<',H#PPTF
P530"\O.B?S'O@C+ \GWTU/^J")$01E[L@#!39)*FY>-,2LL;@"'*E>X JY3AS$XT
PB8RPL%UD^AA9P:5#&RI,8, X2EM\/U$YO>=OL<I]?3X0+T^! ]<'AKY3Y6$%9+LM
P/1%)JW<GKG)O<S/Q))7U)AD]QR%PJI=6=Q*)@*.HG\DP24,_T?_ KE=Z-O]VZ?<[
PD^'>*0A;5ZF^L74!#HXXIXP?AJ!,&=J)<@",!_^B65<O+]&4/GZQ^11D#FOJ6[QZ
PLD\X@RHU"[XH!YDHY>&9AAB!<<*UL5GW8U^(OQ'$"*MQ!:&X\0BB>N]0$.;-JX+-
P16,L)*HD7GAW>1I"NYJ$RMFAM17+9B6-A^,6JBN9JR/H5[C(I0*4@*2=X46V< )>
P?Z58]3AK5WS\UVSEV#A:,Y^HE!^6/OT-L'Q>-DR=/3<TB_!)QT8]J:2AC&#L5KR\
PV"=5.8$Y,':8)^&V<[QV^182[8%>&J5!FD&:)F/PL=I7AHF%XZ35Z,3YX\X:%YL<
P 637Q=+#?R981V>#I=^*VNH-+OT355];,_DX<KEC=1%=:^W\5P:+C7O2I*I:]O,P
PI:@Z,X(=;'QN"-%@7PS^6-TENZN1OD;9ER%-]#=--#:A++:TU>FB*;<(2(!!=VNK
PMGNK.%$P,![.F=BB*G-?NKS2C4"!;'4S\5CTO=6D%1>Q\=['FTO"^GP9@( X-@$L
PU^5Y8QXF4%\/>R*Y8CO\E$7\!Y5<4-T&)X1ORD:\CRG@G-04XO@SYL;$Z6P.VKRO
P?1$'^Z:J.U GVT\W>*<7T10KD2G0@#&8DU0:FD YL@=\6CAK@J-39B<"5 XS,LT5
P@=8=X8/0JE"_63C-1 ]PY=!0L!)&0CR&4H G67.L+<#R7BNT:799=9IX\<7TV8'[
P:-%-)L@QRR@/@%YTJ4QM$2[NN08X'KAO,!5="80*/DRXC<#OPFW;L5#D_,S@NB*W
P?B:ZA4EXP\+!8E<)8^4-X'2.>##1%=LNG,S*KR*C6+Z#WU:"#D(3ANK=SLJ<8#AW
PP*=$&:([-*(7:F?;>>5Z$?X&S'C@ S?<XES9MZ739,<V&.6J^,LL<99-<S<_- <F
P%4Z/80B[S\F:^9+?W)UX,M<WQP0T-BM5R-B2HR\E/]U ZX#W_0YP2'(8-B_WX6:S
P)^HNP[9J"G7K($.XQMU V[_J+I]OZ/(*L&?;U<Z)%\FD*%9%)U[]HV$/G;=,4#T,
P.;D'M!\994X]O//,8M:  L$2BZ59@X9SC]YJHEG'01YOIA[S35H\3TJFV"?%U.8,
PX;E4- WKP[+_6YS7<?\H/2BA[S-^8M$@N1Z&<%TF3\A.&1)K6\")FP<VG'S5/DK:
P (I^S>>V.1EP#OI0Y[\ZG ,-P3@S%P&3N4;G]&8P.A>F?08V\8!\D%)0:;@2JM5=
P?!2E^(UJ$RJ9=.'S?&"?#5\??)UP%=D%W=<V;<>:(DT\Y%V@/R,X@P3_%';Q\QC7
P9Z^?8B1BX#FD+4=I2Z!X5Y0-BN( \<?XPNKZ\M(*+D4'8GPDH/1!+8QUVSU2$$[C
P7V:(VO?LT\DWRTKT7?PK[XEF;;6L,73,<V))S.QV4+JI>F0=8.(L7&ESEPP74.>%
PT4Z7PUJQUHBGEL[N6)6"R;2=53$8RG*UYJJV52BGO*M01T=XJ%:JZCGI(*_]K%NC
PXN"R^\XL,0.6Z@'TJR+J$!UJU8P;C%$1NO"D#C()@?B2=GOJS<@9*9G]LCX#.^&F
PBHC_71P'>FPB.[:\MXBK$T,W7JJWUGRA'2:T*/!I@B;I:5Z/:D L9ZE'!-:-= .A
PFTIIS/I5P)1< )U#L*@Y&9_G*74P>R@'"&T=,$&PD+*,Z)I0:]"=W&=<]SAJ%TI=
P;O0B9#]S:H'""4!<9[]9VI!+U@=<!T6Z3D[V0X6I(5A4+"<SV6(O\4X1@T8,4&QT
PB7#J\DS_L^7.G_7H[&G>//GU#A9%71)7Q!CT0?"FZ4:A$D3H(;3ZGW>32Z5%78L;
P"VK(D#I3\_[#*L,;*::<-C0/1^ C*[Z,;([_C+G,IIQH6^:S0[6IA0Y&+#.7718Z
P<AVGS;>E$&_@0X2$*]4N28:0+@QQ>JM&KB/%3T)JI@P%]Q,NQYM"L#%-G>JSCBO<
P4'I#6Y6QN+GS%"&^]751R[WICI&<)8IA_?&U]A[*]*@YI7W\6BQ6*>AD:1AWTN&@
PU^&O;6]:)QWVFJIZRCH0-( J7. !G#6'2_:QX^RW& )9]@7G4<*O/_<'V=;1\7M'
PM-Y""8!0!3(>9R"P/A$D#.1^09A:SK]Y)SC?)^2+> :C%68>CXNW*?*?9$*$3W.G
P%0K]=/116VJYIGZ2W%%')@6@6MJ;QL6/;-1K=EXI+_I)M\;^>E/6Q.LD RY8ML@]
P.BT;TYQU$O.W!X#2^(L\'1-+'7D+R"U,@5(+5)NV?G3%#HWC*C-0K'M[.(\39!H5
P; '&_X^\.O?/# 1?1NBT)[D+%"?NK4O;W225^I>U^?R?8Z[04P0T0U(K9&Q0.X,0
PK>:='X<U]/AI*0WIG;OYYQ0*%7T2JB/*,93O,_E>#8,I14 -OH;>7YA_:N:>TG<[
P<!3%8+=";\[M!S8C1WS+_<+(:3CMF!YI#'%X(\/.BE:0I^'OHDC!K&6QFKYB*%H 
P$>/;*/QBC&X=B@\_)"'(!T$0GQ_8YQVT]CR*$?B..$R >GG.F3&1P'FY>D=EO$5K
P3!W\7IAVVH=0T:2+8"_H(A3M7#=.ZJ@;D8!ET.)NXJ"S;<;O<)4L;#+Q(?%(!>/#
P[RP3<II7FOM&0S4S%-!U6A<2AFD_D/IK2T](9^5AJ>O'!]6\/_R"(T)RDHC4@?OT
P=Z2P@#0CIR:X#H6=S2EJFZ]\4 52?6>MFC)5&_LH"G-)?98?QC0YQG4KH7;XM(?Q
PMW7 ,GWN^5@2K2\@O4<2!JUXBN7_FK;T8FN,])Z>\<BB1X*J-8R8Z9'VD)*T9&VC
P,<4E9[]VJ-_ND'ARP$\SVDR@F0=";(Q=@MRN+[?!'(@+I]Q_P0F5L]0OZ.OHF=4<
PH6!13@:RT3;T/&>Q66OTBL>&Y_S&HSEA5/Y2'-J9OGR%0VXBCT02DF=GAHD7BA?3
P6-6PZX16.^0H2D%93OZ%&-:) )PI4'  ^LP4X]5I%:E';21(.0,@B&KBZ+9F,((W
P@Z))L;(([2 4"\I!!_""MTXR;HU0>1$Z%Z%[\<GLRA 1L%)!]VCB@U,=%/(O=K$*
P44VF;V_95\0M(-W@Y0Y7&W= 'UU+=V(<=4#E+VE:EAV'O:;)S[E28L?E>?P!>X$\
PGG+OA.;H5;83\]+,_-6KOP\:%)Z8?&=3>X"?')1J17Z60? MDK[ZW+>#GICA3T*?
PK]*!.-C:<9=D >&5E\+GNG'-+8\;"MX(M?F#-%I\4\O5=MP\9E=A_C.2I^2QA0YP
P<E!U'F2=HYI.KLC3MRA(("X1G%LT6)+88T4^!.L]=7.J0W^O<%I<0P 'I(*>@+"!
P"]3$]?%!YJT[^;YV[#C$O;SCRMF2PBN;CXJ8,J!G>W[*))L2L4]5+9<PQM0B;NT/
P#8[YG/@H2XP<\%9(OQUT_0=D.5T'/S$(J^MQ[H&ZZMIA=)IVP,M/&G_G3)61):XL
PW1/7_J_)5FL[21YF!P\,H"/^8MU?['71H"V1U4A=-(73P(7NA0Z/^0/"Z4/^"8D^
PD>35 ']"P%K>:5.F0QA?KS>)>)L9[K$M>L%"@C&I)W#BND_RC\,.^,,>)$96/)6_
PJ\G]A@Z*E;%/>26>A-0ELLL7\WUP-J TY.@7#_(@H-&QS-?MVE!=3^!VN"LHL-\,
PKQ /3($=@COWX$[<54__7VMH&GC'ZNZ@BM,/ZHR3&[\<1S>:$\V3AZU8>BI#GR-&
P_R;D<TD;Q/>(+Y&^LB@IX[FYO3W\"(:D/-YIP^G#CX/KI@SG$R"7@2#LM7*P-B1=
P4GC1-X@!P:1A8O-MRSM10WY07_S%=NK"B"BLLD.UO $,G&,HOM<W-Y4Y- NJK%!T
P?BHM)H7BH<6F(V7=?$N.%3U4]JCUM<C&AK8 \:FR8.6.-!7NTF/?&G,QQDM<OAXV
PUTV3X[GP:3K3\/?=AR,]1=-C_E5B[6!TY_KV C^/T8:<H/IF; I<C698W+ZBP0&"
PO2T9&WCKP=7BU?LST<4%*1COA<A[6R*G>B9,P\4K?NG*_/Z1Q:=0"MIWCNZ#0Q=E
P\@67_'&Q)07M\P&FS ([!8HW ONVVD%:,\IC"18=7",S))3K*[?:)E%'2E+UG5K[
P_2D!$^SLP!9'FP5V!D"0%_T3K)']J!KU)0:WT>4U=[F/363R))5_=0-\H(]ZW4(]
P-S)<,L,,^:-(!C#M!=J-W"L(5M;/65A.HE ./8<[VZY*D@H/A3>HQG7E#7%6,LFW
PV[#FYF&#,H]CHM,^*$:_G</@L#IEEDF&@RN!D)-]AR: DI?$%U%FZ5I+731]+(/:
PYC5M 6I8_GNS[7#E1[YKD%5#[\FA9C0:<V/6>U]F4(2/Y7[[?XF*^: DC 2"U2+C
PM<;H_<;K56+QT/&JIX"+TY44WM?>W:^"4@SV45Y=<KB1/-6T.$7,MW5OYZ?*TX*+
PO(UA&V_)'+W#5)F:.]A9E1;^(L_H)U,CHTL^W\Z:!W3[F1 0EWBO9]%1PN"2JAF$
PXSD-]HB7FE[GXTLH_-0[HAD:YJ@0E]BS:0<ULG^BF+B[+P"*KO2()4E#OHDOJ8" 
PT4KSW\U>[,0,^CE*A*EZW<GD$*2^47DG7WF53S+L[O*!8[."]!HT+$NM[]03KU=J
PN6AQQX>ZZN^1<!(D9J.]KN+R0?7W4_#GKWZAB^:=/EC.0+'+N!1*?F_!]X=/1G;4
P(-A=99P;;DV*6>=8I \A*>:[HE3Q<:C:F)!\DOO#0A&2K[D.4J&<GR+18()Z\.A_
PS@DL6'(!;*Z>K&E.-)(=C'PEHH5B,.<L<[PT$\=&-7:_=S#A(\DDY^E*PZ2!"WB[
P:'T"RMRBD42^,.[!U1,AS4DZK-J\#D=\!N/J2IR?@,\%]TAYBSI"<7B^I?(53UDB
PJKG5] *Y12IH!0Y&<E)Y !9V@'[&[>P#@MVH6! K/3NXY?&MFF!;2Q32)AE,"7S)
P\F"7+K]DU0!Y-ZUPA?/Y5W2IU>B&5+L_1/ZDF#WQ*7@'" 2>^*(D1Y^G34,@?G_=
P[<MM>A[4BJC#GFS )O&RJH%:9I,^;;]FJ/TSM/-/X8<C.VBA5L0-W%VK#.^]% '&
P%F?>^3R&>FQBKYJQ<Z/=KV('/)\P ]#(>/,L50N(NA98IZ7ENP_R3'^*=;2>EDSO
PM(XL'7EJEG<)^&UE'3(EH082N"J.VR4E;VJK\0==\ZR B.S+:H(%6YH-'M 'W0)=
P.>'J]-:7#[0@#^Y=YX--D)58T,Z@C %@D-PQRX(Y*]U^,JZC[GT@<6Q/Q#M7.L[E
P&2HAU.IV5B@KL&=??@>@%(UW1D;[1P'8@F?A0YFN]9^X9.*6U/G07%2GW^/#0VIX
P69/\L6,EFG.==T(+>OE48.@>."_^L<Y9&]UEF&HW&XV*VHFQFG+=,23J-:B(J'T;
P'IA!W4+'P\VB2B%"$9#68/E>&98TI7U@?=\1(S;+7Y6_'*Q*.<X_\1M:A9$[17"=
PD6(<3HIY%-PX7<NI.P18/IL(*^^0JXQ\!_JFN[<"*V487N(UJ%'FO,D5D%\B0K]O
P5O)^+HIPS5E.1WLV#5(J%;&JEG@N^H"BZ#QM2T:WIV"93#6L04^O,1SM 1:..93,
PG"7*1(8E;T#/%)ZVF<74=0"DC:$4O[K'2 LF_7'G?[_I(@!3$JA.8\GVZX4C'U'L
PO3L:@;-CNPQ\1%M3AY3R'7I_LZW= $9?,?).TF2YD@*V"Z0T;XM;X?H+3M9G[LMY
PL,L-NB_9PZ=BX;+:ZR_IQ9=='%BG8U*K+3OL<#@>PL_D)+K7U^J7W(!90N$M*E@'
P&$V-E<0W+EBJU:,1$)SD*).93GD^&%)GEJ6?R#(8J$]082!4]*#DHL\?]<,L69JK
P)</9+2@XG,KJN1!*[HNZ%VS/]-N:!ZZH%A:'XTUD;+*JKF8N3 N.G+'0LJ]?\UI9
P[35@RWQ\17_V8NSN=K!6-&YH1LUTWUT)Y62\(6[NV3M =7S1ZW5#CS; LD>602MT
P]7WHRQQDI.-U@*AH35@3H+^D!:_D-\ /BB;S_J;0 A@/U&CM 5@PQ#9EM R*]'I%
P;&!#YG\*H,M]\ADA9>P5*OCI:&89:#X2;YIQG@9/4+6/0;?62G!Q'E4'A $LUUN\
PW$EV/E>H=T^F" R(! J&)9V=/W4#C9'BD[5P4^3X'J'T&4;(K9ONE4"79"MMEZQS
P_+@0OE$PU]/R T%RPP-X!"?%IE8!@6L8 CD4SU8YAQY8RI5A:7Y/>WK'.J7^[-Z0
P-5Q7B%K(7AMZZG1V5C];>9VSRON6-37] ?VJ+UI)G&A-^F-H% 7FU$X"EKYI5A6&
P27.J:364"D,GUBC$(#EWBGH1[GP=B[LOMA)*: F[T\F*^Q1C]4#10Z'\I>!\:>A^
PQ6>?-\".@=VUK9JL(2_W)\YO$H1GR:$??P]^A.U.&1@+Q?A=*@R^+/ZVEP?4R=4W
P'1+ZNWV[!'\9.;\!,3-7WE?'=G(5^D@#Z4UR8B3EM6EZ.[+S]L>DS 9W8]@1^7N6
P<=S6T +%5IH@,S^ F"Q77W0>?NTVIL0RBX+2%54H^>ZRR?JKISBY7.__*8=NR/QU
PI3)N]B[IF&Z%)'!$MGF#<L&^MS=EO\0#0;&6IWN^P6E\0#3Y;PR7[3L+M:?#PS6)
P.*]W4GDL1.DM=$=X-D$T.3%A ),+"* 3V3GN^%TSHR<$]0P WC-L;NKV6JL-$ATY
P&>6U-5AWNMXR3<)ELU47OB$)P"CCL-[(++TC590CXS%S5E)H'H4\&@C]H?*G,T;(
P:8S37O3'_9?UT@_:"J3S48?J/"$<8G%4U>S?@-.9U>DD7X0&_<$$#V[.2 \IQFSY
P8C\?S7RN<_7LVN7A?- _-UN5@@AX<7IU/SQGR0V%F<=4Z(<G?U\"V30PZ[M\]@9F
POL8J 0;8EN1AC>I@BX:DHW#@K+[MAQX;?'4=G*I"5;+0M&84&U.0EK+OK,BG1&Q0
P* 5S8<">OG#ZV2:M2OQ;;EYT>5$$=RIE,[S,5_P:U-".60*[$]Y*M&<JW,2KMF )
P[S#0OJS)YW7I.DI$="5"#&AH\^&[XY%51D%07P28"8+W/CL4]^N?O-=&N]9A7_83
PN$0'7/IXH[.:+B4C."IX-9R0'-1]*4^D:0]?% #6C0ARL5JX*I#%J_M9G3L:2)%0
P^(YP/^D[#-U (/VW]:F<Q[!K6P(/E:7^E C6&[/<B0PT3(ZPR4ORQ;("YVQJEX= 
P56.E!*OJKJL3N5<\U(-67E[LT*< )4U9;K YT:OH[XC3%"5%@+A"J?63@WQ^Y9<K
PU>WK(6TX;#+IT 0!6CD^W#T!3YW2V=I8\'KDF?HB#\DZ/;^76:^.4H]]':^GGMJ&
P#5IV%IUY5.GO>F--LG*YW17:U<JNSO1U4PC;@@^'(^Z2ME^.R;K+'!VJG20Q9S]=
PG;HG7NN[HXX[G.V(5>.=+@R7)KD6"<"!Q_+KF,&BX/F4U-.0\3*9&C';8LA#BL!E
P6TRN'W,UR-^VT15[73..Y"Q.<)![#F7G.JUL/ 22RD$YUFH9'2-R]ILW@@"C@7G!
P--[0+"RR?KMIV3MVYHX10QGMG:0 \5[=_/I.6]=(&\5.8#],QXUSL?WTG03R/#Q0
P:/R_B-B,V>N)<U^Z9Q%-B3N75,]GB;KMSL0GWVE5%&A\35"ES"^].( !FFWZ_?._
PPFY]<EGUVM0F3!A+'[ L?J\Q9^VHSOKA=;Z."?&&H5L]12)OH'X!\P.I;>-U0:9X
P?Q;?<P;([>&A_O7ZJ(RD""PW=KMYB03XPE_:Q 1W'7&INSCM;,%I!&[2M6.8T:0H
PZ9N\6H@'&@N2JS2^G\%YW5=0JT!PV0Y.*CFY6$I-?,(I@0(X]%K[7]9KCN#6#^Q4
PD-M===IA#MU,%2)@<XE6,X$VL7-%9N#_WL^EE=>U$;7H\/OVY5,Q=UYKWMJKE\4L
P"?7DR<VT&YVRI:=;B&' =HU@G77DGN60;+Z#MUAXW91&<*H>H_W= I^W_:BVT,;5
P^E=AY<(ZUG/BD%D]#_Y^-\)_]"$CE_8/6O%B:A!S53%65B/6]B/<3==6ANB9U_K;
P^8UU7_GY'=-&[+Y7I;*#,P%3"W<XGS\ETL?>8J0CO5XV@>6;DL5$&5D$P$8)8!MK
PM1FLS#Z(J^Y*B!81 %>YY5XCC3GM7)LQOJ \Q#%=J>0AOF^E$LC+F ,#Q7\G4,4G
PQ"\>:?19?&^&?NJ4-UU<IURX8P?!SD*7Y;,VC3)WW*6 3>$$9UR;)31:C/4W@5ZF
POJNMFR_30_;52IF1>VW(E%&2JJ"?<*A/YTFCKT9>?;\U2DT6V90P:3YS/\R?\?18
PTOS?VA@S.)^HK78.Q>ZR:Z;=E,&<B@BI,1X2D@,U%<2F@F:0Q;O825([H3K/0N_%
P358DZ6^9QCZB8UT35CRQ@XSLV"3[4U-5: G4K')R[1PW'2P&AH>AB^&A?HYJR6&Q
P/LFH3*4JQ3M28Y/FR[XYMI>AG G?$H0B%FOSL5D8P5J[<;&_F3I8L*4^[>!8@+;B
P4W:IR?SAI]:Z4#H,BDQD[V^$(%+XC%Z/+,!(U@S8^EDSW[TG[&>0;==9O$BXR@<7
P#F04?$5KSY/$V9UYD6:ES(>8Z/IW@#>T5B3V7GYGOMK:OEG7TJ#W5VA@+8&\MM*)
P3T6_@-;T[W/[+R>T$T,8]BJ$\NR)!VSX[6Z]RNW*Q(R$IDZR\9^(RT0F?<MCD0_@
PF#.T/P7G+8$PY*2(37#>PST5VFK.$89/V(>9.4_\S#^&Y)_<HG+X>_)%D7]JD+//
PU8.9VN;2[&PP#C3;/3N#O73QPC>V._Y#8=AFF'Z$EXT:?EHO?>TINX_3S+7N+0@B
P.M6[*F?58ZTX+%XL@[':(Y9@W5F*OJ09]QJG;DRE[;WHH:$N8<U4Z!J&1HW ;GJ 
PTU;8H%SUS[W.;^4JFU(//#V+ZS"RG(\MTL/[.OY-X;OZ&4VP>M4821]LPCTVK5/:
PB+U[*Z20! ^.FZ1-8B+NE/79CUIPT?Y?.D.-@#$LI_7CDQ"L[;I,#<2O)@E:?&G#
P+9"K1^Q6'!1@)_O\*/W-PJ*\185V%X!ZM1*1[G1?IHO4:HVR\?D!OH,V5T/X+8I$
P*4V=H%Q/L9F]LZ:*VXF&@+A^W:H9=YYX@YDB7^!Y6588/HU*,#9I!WPTT5\!Z'08
P#U_ZB-B$@:D[:MT9+7^DA]-)I-JF"<0!8+(^"T6+V7C,4WYNRO%BCW;K>J!*%\:E
P&*.B,;C*_LFO7;G"02II23+,!".:2+K$9\DK5Z80SS1S6=D4:7)85$MQR0W]QXN2
P+J8OF"LOU3- H835M/[:J,?]'L:[U!PM@&#OD20GF3  J1S@Q#+6 46_QL/AMY[9
P>$HK\+OH(PYWI4V_VRN9E)O(D5,H;@NVNB]F>I?GE21K#5&\-BYNEY87N=?I/%DE
P6@TB/?SYYTO"WBZMF#W(,O#P>HJMU"N]#67-M]B5P[G*P1VH!4>H@JELFGY!SEE\
P9/:NY?2F'6RE-!!?\W392B7-0I:!M/:N%4E[ZK%?MA/LM$=U/O#0[B:\#L45$.U[
P;"!=WK+F8T%"='/U;\5(H42TO4NW_11AASVL&W)_.G_=KU H9N.&H. =+@Z(Y1H=
PQY6@X)^FJK+@YY]8CPH5S'T9?NNLO[<LS(<?VA-;W&$F-K+-#.8W$WW/_("A3$;X
P54PDAH]\@8).4X+IPIKN8;WE(R?!J,/"[\^NCK.!!D")<P3'[&M8[@DAF?1JEM@'
PVP@K\&\#(6O,&IY+K#:1> FP4F3T&323*-5,/!%U,G:)ZRVJ3&%(Z)P,K:&"?6V'
PF%_\?&*,C%+'<ZZ+%>OQJ7TT7I79^HC?$ B@%S J1EUO#[W4]'JAJKR4%<;".S6N
P4V1_9 K! "AWSMV<ULB71QJ!0/!@&;U%;\HW!'O.=R5+K,IVZ?'X[ BTILV+?$JC
P/.8\>+A H;5?'AL-%VD-FWA/N1)E>Z!DGBX20+]!8''!P59JWEPHV6MN8?BP9:A)
P,1[B"*N_>48^\81(H4_)2TGS/_LO%P([C6R:]DF7,L 9 "B&G\$]$!M?=H43'?L^
P$\CQ_7>?@S$CMG@,J[62$H&C:ISJ<RY*>^.T["I?EW,0]L6=Q33^OA?\*;_8&0I5
P@\/^-,^/>"+Q^.17=CAZ!BEA,&.$EF<:A5=/W-X.N5(AH</.85SV;>>[A+O: 7C*
PO-2((2I;,B6?&D$4/.^(;K ).[2.H-="78-(?=&WED$HNJA\=L;:423J-K/;<0[-
P?=2RNQ-7 7!9=3]H#S34IPHZ,D>&/E,?+&=D#@<9L]_7-ZM.44;^JHKWB MF!:DD
P7V>P%R^"1P$H<^QOHP@)Q<@FQQX_G34R3Z;IWG&#T33V#E[0L.)<WA5_P+'TQWT9
PUJ"C.[-.(23<($ ,Y0C"7?T#W,VA!-99"2!>I?F:C]#!K,07CLJ<LS!O"\[0S#X=
P097H!%F[O(Z8A.<*)8P6$F CJQK]_WW0^]STORZ9K\[:I6Q%O]21H3;4*%9.=RD(
P?'4$W4&CX\KR&97Q>DE9;RP8=<H.;M/?A[]K<D?@B-PY]!.<<F.S:S>H:($Z^^4Y
P06=.\7LJ)C:9/6RR<YO923>ZC2DY&SBN.WU+4.63"P]< $2E<Z8\""N/QM5^&UT(
P3:<DI"Q@B,(+C6^RJ+#1/<   ,N,G?%N90F\C>DP[PHMZO@GU^BOEV,.=4^9W83L
P_;R\MKGT9B5][MZGS#^6<3/$=)8?F-\M8+F$TH*_KTO=$VUJ%8A=HKG9-"[+-KDM
POV%:+/Y>>:#L4^(5&+&R[5:=]*P7DX\.[*!2@;!5:%/PTMAFF$JCW2CYJOLB<7Q*
PK/N^ZP$Z0X',]QNT2*8G6RO &4 W:LJ1Z@%7Q!;^S['L'GE?OAYBB)1ZZ A<\Q\\
P*Z[3W15IF?'9HI662U+TKO$;H Y4._+)]<&1:9K=YH?WL!@J4(M_!F19L]VL;E+7
PU"N5@CT E.XO$NE)\494AT+4'Z-EZ=RG-2+;S#OO0289:_]9[.=PUN^$BVO!$5.?
PO*Q8QJLUJ<OP=^; =6^"7=5>$4P[2X3C:Y#GI.W28:H=95QDG2Q?HFC&IHA[50)8
PBC<GRG]36JSZ=JL4(9L="[-?U,ABK"A&<%TUY;!60@H@&U4''M)]>I\8][-Z?T7"
P$)YOK6_S0/O--A?P[(HMM!AEOJ5LL69^W='1%^:?6ZQYY8R-H^?S0+D^TY?PCI@_
P #G& Z-,A7L[AV/IRX',N#)3:*>,5N9[F&7U_1SVBY,M@P^$Q2(52@S&.P]2,Y7F
P(U?4K6S#P.=K:]?/ODNH6(U:.M__513\JJI%G)XE'LQ1U5+K:F5P\WWZBGFO,*PE
PBD]MV(@^:X%8Z;'6C#L-%'/9JX?I,PB7#C$K!;!V@GDVN\_\IU)46/E5D6407[9!
PL\DN1%A^N5 &2+J^^C4623J<D)6\#1?$:%'DLB"^)X:FP6V?_KK_^IVL4,U[&.B0
PGK R0-X' WYVQ-J!SX(Q*-:[S7Q<>N*". ZYV(M;;V;EUJXKE3,5!U*]D+2^^&C[
PA&9(V-XV0WOTOP WW%5:Y$0WO$*Q(0/VII<QSCYC*NV#CZ^@H0@=(ZG X>"4H"T,
PF#0<E'8]IB7,-]=<G1)0+4'_2FN2)A$V.#6<Z(>TE0G3([,ISS]U':!>2JRXL1 J
PIK"?'PT1TE0DTAFY&(TR,313/'D)H;A["._:9LO41%I+';9TL<"P>-:SU 0]]EXV
PZIP1F6/CWQN#>Q-4,ZN<^TI!P,#L(_Z]/*BC,WO$?OF3S0$B0-![T//HD[TG']6\
PX1+<SZ5,JU;[Y5]45X 19Z+E6GZTAG>042&+EZ'2_J5M7"5!!$[3Z&$3=N@=N>9B
P:<3ZI:WL6 KFQ>8P2 2E3I[W<$D'$4O\*+G;3 &9DD>!NA,*?K>[_F  6&S]\+3'
P2]5J4O3XM6,@ME9(R6ERX!&?I'(<B;LQ4Z6 8)H@I"%VW]XRNJF;5UZ\Z5<[7,M*
PA!C=PAZHY P9\]FJ:=-O*1CRUHL?DS"IOEDS>=V&[^:1L:!],W4K7&*U/&!/$EU)
P)GYUTR2HM"</_+3GP=+L$S<2=GEZC1=)@2<H,MTX0".G*G2(;[C1\@VHSKBJ\83Q
PIA=?S>H%!4)8 *;7-SBDE5^^6Q^YK3A!?A^2Q_P[WY$W8N10+,ZKI9NW\&I41QT?
PLLU%$)/U9R']>_Z8B0!%0H6SQY5GF^[>GF/8J1(J3#R 6T"R\E"67D+9,:.![=9V
PZZ*+>IWJ/0 (<-/ YGWG30S44QE<"NAWAG_2<5$"0T_F&J:TXL&TD*OC(]"C+$2"
P7_O:7J $-1L_0-=ELDG+[6P KM?I-VE#(?43>DI=Y%HAOID0"(<!O%"P[R<N^5[-
PC.Y?J3R\)\T;?X^-3G8"AQYE1URTLP&H0@)5"*FS:9@&HL&6EO%ZDKV'L1?1 L/<
PE(CP*?U+OK#X^G#JXF:+V/JB\'<WZ-"H"@]8-]-;+<KYJ%"3W+=L98$)RV@VYL!;
PEU=G]7F<RVZA:H&/CLQYSUVPKA;WUE (0(7NN]G0:)]A%:HZ;0X2_]$,#%U/A7]2
P;(,\^_5?Y:(765.V4 M@/D12B4/#!II"K90P1,[74A6M+A^[L6PO8>L586D^GM*L
P17&YWCBL)'$UM Y<Z)K@23T0$4+ X>S"&%LIE(-L]FYD>7Q/%Q]KXZL?;KA[%E5:
PGJNJXO(T5E"NR[2MU]+&YOU"6CI9]7U48AY85(PF'%-8,B/#M9 BBN9)399&/:X 
P/C?HE-((3;1[*NFKG"PW1S&48>CM]&WW#VMUOK7A\F(!8I:*#@ )U@MX!T25<^._
PM2'%D]NJ1)Q6?W)V7=TGWQJY7@C/QAEDT3KWVP:J?ODOW9<&=_UPH*K"!E64W\[U
PQD>\Q3$8[P(7S<D0XRR-7/_M=5G SX:?(IP^P7'_FZ)9Z\[U<J%GE>@&\P"JQP-7
P3K?*_6G0($7HB@^'W7I<^)*DZ=8NJ78EW8AK'0]$KB)G'YZO>4RH@.]#/I-:;GH*
P_P$SEXCA1AZGVPT]I%PF+-&T:E495L;*!RTN0E<[D<GONL<Q7Y=XH>FN^#1'2H\<
PYHO<2KG\&?^+GD?WECJ:H'7*[/)PK,![9'U>'<G7RX=:;24_979P\+[3JO1Q,K;@
P8S-:?]<]0$!IE0-^$;-8=G*M)#ME(K>9!=JN=,DXD&P>ZU;,6=.,$ (/(554!\&N
PAB(!I>QF6G<2\[W.N7J=NZZN,ON\Z/):IV>G#:S'>F\"E^(0BG!.[61)IMB1\)0]
PQ@;KU*4!*R?UF_A'B"FKEU?L^];(\6%V]40VE]7HY/T]C7IF0TS\)[ADDO10?W^.
PP3+-VOI_G?UA.4'^69<_% Y9S[JSXOH=JE\@=D;>(WI&08+^+C'W4(#%B8._VXJ?
PV2:.L2$?K 'HP%*&;9<O8E<5 Z_X/.^*4.SDW5S!MR:2B_'SS<HY7S+"^(5>Q,6G
PZ^P#7ASB.O)3^LR+VJ4\I2,:Y9IJVA=J]3$[JX'64W<8N/$F.P/)!73.Z10LIO?9
PR%S7GGI7=C<P%^B/P3X[P/05 #D/2\+IW$&YC!?0>S-FL2+9'H3Z@+#M8HAG>:77
P^I&6/!>,!(:1P3>=@@_L3&FCMQ3LFG;\(KL&=M2 S7EB5W+G57)TA=/(<023/:3:
P;8LPMTVP1W-!7CX<_ZBVFL?E,!^"QS0-;@&HR2X>*>!AVT)S#^5XGJNXSI7IK>".
P<HR)TGK'[D^<X9O%ML4J;K".@X7HB2^6$\\NW88@W5!V;04"RUA^OQ23BX-LAY1C
P 9"%M+P0PO#U"60J4"EP/' =)@*=5A@K[REPO-X=3W?.&V0V(M>;T7BE1"^XZ1'K
P7>U+MWQW9_ZP/J>,E56[\Z'Y:?@(]5N"<-91,*$C9=:O9G@OA%NPI<2D&[Y4"_TG
PL!E =8S+ =4SN!E^S,6*_9\STUA\:I ZLPT-LF91QV!#"5_Z^52D)?Y'1>GJR#* 
PB"C)B^OGP8"0[4CETZNQ3XGT (\VSVT)!.8F3<2M]:B#T@<+(<DZ.Z%?(+RU3/\5
P8,\=NXQ:6')0I60KD9T5RF25^I@7:^;+!_6JJGC/',E59)DKZ #"XG"<#GC@+5M&
P$B&Q['#ID;YZ;_K\+S-ZWH1_(^H\BT_IP/5F^@5I4O:LCK(IKQBKQ%F)#*-_]Y7-
PZD@_5S_JWJ4)+/2:8@CX7L%^-9K>.Z4U\ #%:$G7$,I:&*_9X3-5VG*X5GMR))5;
P^V\4'H,ES.VC!/@R!1AX6D%&Q$@T8I@L;WW9G)Z>1G90_EN!Y)15^!45,8^9S?U8
PC;[%C]([,NUZ LZ!$G$=HL2:>T(2=BV>2GFKN5!\&K-/N4P1P5(SZL.JK*6;Y N,
PL*-BNA6NTB6PI+)TV#2*F!=C)2A^MD["9PU$,;B39GQ':72N.1-/QH'1B4IR&@-R
PYI1ILD)QIEWNN50V6%-"A?X8#H _Q3Y$[VYV[83]<-#\O:G8@DZHN4.^30X7ZAMK
P+0591$NYWZ67O[UF:81!UHS$[BAH&VAQ2N=F1*@;3X,X&YU@%\OHEAT4X92KG@Z"
P30D@Q6!3:89DMJ* CUWR[Y)[3MT7#3+OOED#A)HZ6-2@'/LCHQ%&]YHJTE>_\./H
PE=6A]Y7<+2I(U$5J@^4%WEGU]GXEY*/<%H00)P)A?&LW>=P<.BE@/+I_89L^3ER9
P*[>\%;FV:NC="(%&%:_JI42>171@<E8I"K''UJB@0+(>>LRZ<012@*KA1N,V=UK8
P0I',P'"]-",Z@"!GQS*B!?,3-M-F#!'1$Y,-1)-%[SD/ IR/U =6,&<P&UGA[I-/
PL,,#0@:5[^4(]248 #X=4$PFV.>.M;M!OQS7\9^Z=4L7D1E-8.)VO-$XM$#S#$9;
PJK*]%XTZK_N_]Y\!W?N>'WT&DOD>8M Q*MHY]:#!/"I*A%V(>K/0*2#E^.>NP)/E
P3DK!9>40&0>4!B* LZ/@.4V"N&6<?YYJ[A8=WE6IQ30]O_32 0:=9&0Z/[1S5"CW
PD$&KG69UG@F_+._J<"]J5BFUM)P\_4-/]];Y.01"%'T\^ EZ$60*;<H6^<<96_)P
PXQL\>-Z-+K1*:$G;S>O10?N_"K(L3-'_HN6G8NN0%^J>J5\8VVO0WO%G)POO5HH.
P@]!:4(NW#)'FC1-1Q@#)/73F:!#JE";(\I0^-LIA;.'(U)OF?T(]9\0HZM_9;K)O
P HD _!:,]WE%]-/JN_ SD60G-[,OC*BAB_//CH\2R2+$D ,J?JZU<JHN604 7AL6
P<[]!1U30A1Y^5 QY--MW2P9].G]R"DQ)-4A6U%31,Y4 =-Q;A5<IR-3 8,?=S#UI
PFXXL'_+ XYE13#/XP%",:G:34HFP?Q[\T%[?*.N$[H=M8@(VJ) Z)FE(YRRTD7I\
P,+.1D@S' K4'83F)8M:PJG!M CN&,](K#?-WO*-2(K_(D1;L[TI&TW?1'GF=B0:0
P]EK"5"+3E_^V',ZTH*>,BX%QJVAB:=?SJF*PPM-!A4IO@EK+G OYCB9N#IRGHOJ$
PP/[EOFQW;JD-@[J@"='-ZCTR&++\XTN#16\KL1;>B:\-?=1["R?N5FMJRD^93D1W
PJO?:A=.RJS*Z1J'H15,W"@PR=V%<Z>^3[68TW$'0N$5?U<=I6Z7#T>_<!=A;RQ^I
PJ+^#C/!LJQ)4$<-TMVA63L+]AEJBO\ZX]?SU9SZ#F4JLFB2/L] T)4P^C8F&X7M)
PP&7Y4E_>ED?#6_]CW!8L5D/]9MY^D';9;4 SJ;,XF;'U)7S-$JB79\$WLRV?&ZE6
P<6IKDJNVZ4D3IB?!AJUA>Z'(Z&J&)'0SMIRF,'KH"".^Q^,1&3@/IJMSPL!'M:Z-
PVJS8_CB&PC9TKE,>TEN.#^FUCMO#DJ5\SS+4P&H)T6 /[T&\F[F$YO5]4V/HD/B@
PVS0#&6'(Z^&Z%YI*X0>V[2D^IE,.S*DZ*Z8/QBPG6^G_5TODU6EL9/JNV,H=$YZK
P&ORG(- %#E >V:U&-*EL:<^H"6(T1AWF6PQ!C"9_$9<L7'!Y4O;%K?ET731YV!C:
PE,Q<=#'EK(&FO:W( (\>%%*/RU1)>.ZD^Z9ONA/V.\1N28]CKARY9/8M.3-V5C ;
P'^(?5);(5M5G,+A&"1X. @&0H0<+:6SB0V2)4J>^^<B1B>#(H(UWK!ARTI3^Y87W
PG(;K$'F4Z2GN'FB"X1+E8=E@*^N!ETP)M:?WT)"DB;@_MVNB$W) @\]=,QL*7')\
P4JK9FP+!@C][PY.\F,PH+\% #VT=%3_Y5ZC9?&NU5K3,<_:H0)$C&1@:W6N_(VK9
PZ9M_M/,>#T*W2AW:+9ZF"78#4+A7*^P_$3\*W@\]SVZ9>AOUEO"G_]AKK:&_,Q)8
P%LL#Z@7D.M:M5/=+,87\\>_?$C$N?N>U(N:->[3=!FQOYGWV0YD_ZR0F RTN)*]!
PCH4ZVB09:ELR5%9%S?*I9<%VJ39[#^-GBPN[X&LKE?L5>43JJ4L2>/T$[<2D/X.6
P_*\\9&5$JDT[_;?-G-RDG\*=%A7(6[]C32_O+-0L'(P%E4;D99$L<V,,M\-8PKE-
PR-A7&<O-;Y8V01YV*+D[.^C?W*A#8O@/GJ,9O:\ZI? GE(<<]=%*]E$[;E]>8^;"
P-A^  N5614 =_:T49I_WK'[Z<(GN<G3L]+$WQN=SQ6*>&)"Z2?_]+3M(AM;49*\'
P,B=*Q[1 .C:PSRY->HC])RT(X/[=Q'K\DJE@W@E]2\+\0^L]C&@@J!WEF]^AL9!H
PV4?_INM1&DS06R6Z <-LR(?)M6+]]1>'06&-T"GE,_[O<J049'LW%,61PK\'6%6C
P>-KLJH5V]E.'E$A?X@? JZ3,E/!9U_A697.LRQ13GQSW"<(N919B)5Y]?!>"U^4_
PQD+=WY%/V1T@"<"5!_'CA&*/A@64F;2"51*&J#>=A3L^H9RDLK40&7@TG\QQG^SL
P#)0:^%&4LL;(PW^=W..%S[]ZS\/),5F7S\H;]$IW!Q@(6MC?_D>9Z@8'@7()WVYW
PC /W@NT*+<(R Z,N0Z<<.4_A'3RPT3Y4F*A.T%JQPXS4AE(4GF(F2;GL8CFE\K[>
P8,5)6C9!%\1PX, 0^8T;Z+L32DQ-<]<E/#"Q9_(S"/N_6WGN2;C2Z3?//S7+S=UA
P 8!_&YABB<8WRY;!;3[-#__LTNJQTZ<3XRX0HKY65?1L9NZ<%K*V3)@#(2,S1H%>
PXG-Q@A'VU[9895I8H^&G=X5THMH[K<$&0GT1G-VM)0$61:\M=>.0;@P1!]C/9_+D
PH<<;QH1E@0VB*\_>>= -AW&E;25$R$==Y8]0P<[7-\V-T* $K3P3=&D00/H?P@M%
PP2TYMM>4NI@YIT4I49'! O>/FMQG@=%GJMJ'+,EJC#CL2"V?;[:Y]GBW8H:O'$N=
PA$J=.-(]A"^D%LL%#A0,9;R4,X^2Q]Z'=<*&B9*VQZQ"0(=E4.-JH@.YZ/#Y('^<
P#)>U#XG:;*A'Q\&:V!. X.:_=48OV71*JF%*IX_GHFI:$P<%HFD0)6&_F*:FG'V&
P:0JX&5;DYO*W$C."ALB%+TCJ:P(AY(R(/^88X/2?*G<^7=J$LLM ]7.;.1@(^/9-
P);\(N]BJAE!Z-930F44>%K_\D[MIC#+;!U^A/\Y_;X0U-F![=3Q P)FZS*>9:.[N
P=XIM)2QIR$J]0C68=FFJ-,=5);IL7MJ3:)M3O 3RTS<K17=:LF?3F+[ZGUFQ>!82
P!((UU.^HNBCUS2Y[S1;C+=B='H/@I4"UA[IAUN.#/Z8IJ+HG9'WS+/"(51=]X>T,
P8*YO#A!+@1Y]^T"4%^ \4TO#V9UJLENZX?.<'VD08Z*<S888,3+>ZMNY8I\()^.E
P[E1@B"^)_5=L"Q^FR9-F$UW']%I6L$KS\97I4U8#V?0@G4%RL?8>4NPL*8*G55X)
P2ZK QP['J<.61O?T KV/,3MN1<$IS% .Z.I>&_1HE'*KYV@BS'^BAX%Z#</;4_+&
P&9R")OJ7.U7(N7&S=6BKWQ'0;0Y+&U@?"C&58_F,UDED[+ZNR)6\9LAQ!Q.$@^M7
P C0QU"73-T@H/?%7U.GAZQ$M:K<+JL!#X+?Z3&J?6SR)M@\ZK(7"B$-A 8E9:<5T
P_FD9(E0H_6"T05HT.R%+4P'RN EN7S0=Y&MQ+-!3%HHEBN$WVB9COKGZ2>W ^ I2
P6'TJO_SBWLB$F*SSRA55]X5 C\SHIMBS#@!K*X5LS7N0S1G=[H"8NK[D^YV%/5XY
P*$^_ <9(*))]%8Y"#--'J>1U9Q0K!,_G[E=AB#1W_0@KWV(-'=![:)C#9B1XP4VK
P;6S(G>R*O)3E3$5[NGF#Z]LE,0=G/FT;%^%L1&K\,HV9<U]76KR\I&C-QA88"8O-
PE[9(@0>&V5?E@:@]=)FI]NS53>FWBF-C2VHE,8Z;BRQ'QE3[BCN,K%BY=BR]&U.E
P9(AP#G'RF=V>O"&%>N./07Z&[\(1&PFH-QS9]&! VJ;LXD4BL'V!U+T%K\FDY'8I
P2_E@7@8!)&CH\>!U)E<T&9<6X.?(=GD>[2O_[1GQX7<B$KXO*..P_VO8JIWH>G;'
P,Q^*)T0.A \Y1.Q_ZG!T6GW3+C.%"_@D-W9KJ<_Y+$8_<?_4J]&".'0UQ4+;EA2>
P4Q,\R<_NSB;>]$2H#N&P.#*W?V6;.:H4S;O/%^.H$TV\)SB+_KTRF91F5=SMXC^.
P$0+9H[?WS=E/G1O3S!M6OS1\\NP!\.GV66V#!TM_R2U,3K"%E-[:DO0D+Z63YY'T
P<,JI9N;=[I!3GEG;(7E&%G0YL/=*-]\7Y68H5B6246.3^-$V*BQ!$T(DA2_A3$P 
P)@M^8M_QD0T)SX'=[GFA.33M(WEZ:ZN!SLI1AW0S-D1+&/3^)Z^Y"]R.[JX F6C^
P7^7;8+GUDG@\!3QL,("C-267[1&\EH*+!A0J-NYI8?4("CJJXRKP*%4EWT.<0578
P3OMTK.BCWV&*CW7ZEN:X*UZW#.^JE!2?3]J:%R%UQ% :8%[A=+4E4_-P1>N41!CN
PLWGT(\T>,Y_ LN7(W]HT JG^#JR63-?9[:5JLX^?T4\H,-0Z8?=H&="6?>A:>]&V
PY[*X?6'=7C:MX 0S*\B->N-$='KLD@=I8I>V0 G8"<ZSZZH%T(=INJFZ<2RGT;=C
P9&;O ;D0K%@=<6@/BL/-+%9-Z(WP'FP &NMZRE:W"E@:XGT("+0C20C5!4%'/5Z2
P@@AIGYI,Z1\A[Y6UD2-D,BK.Y![C4:2KDT-@?Q^;X_RVD+RS*%/VF0[!DO5>VJTX
PXUP58WP\,=,+'2F5* GK6W\[T<1578D..7=MX%_,T&/#TC+0&(E3MR.X%SGI#YF<
P03>P^] SF2<H YTFM(PHE>SO/1FP.%) ;X?=+L(Q7=K+DWK6L]^EW@O"%,%J<# B
P4$I*=A3J[UU;PK?E[[#W&ETT6,49@# DO$M6@^B@KZC<58/Z@]O4XM,NL\H>3+IN
PSEF:'. !;&C?G^M^A=L5O_]2LZ8N(L/I&KE4-\P^V 0Z>[.9"];P!%J2=ZIMKM04
P"R^8<\M$03FZB^%50V;QV9776?BA)6W/ROZV<!X<6+ZXHG5YLT@PDVIGSK^/U"BJ
PW*0C H6+D$<41?SN;*) R4G3:'>L;<-PY:V(V3NP,*0J(?/(>^UPUP!-XB;Z<I-N
PY0F U..IK@#)=S!7@J-I]>"?Q^[VRGKHU?O^2T2!@O*TZ.XX,6VDH%KJ18A1, E?
P 6;/B&>2<?K*M)LQ*8R\V2;RA)(\>EC?6N(&>1$:XB:@VY5K[V.2Z/VG*:"T_T+&
PA5+BIJ3#C75JO<$5^D'SPZQL]?5^"1NJ3TE*?<">#DRATXI3I;T33]09L+QW*RA*
P:]!P(JG4<_ 4I4"*W>M=:M?D/''T<,+0RT,),](P,#<)!H=5NO1C0#08'^59IWH!
PX=Y*"I'ZC6>-_>MWPCS+-=U1*WG<-."R#G-X])]"VBFKL"#E.Z 63"+CEU_<NMBF
P<4!#2$4),W-?TD3C0VZ((B@>V0C7-9*NP29:QR:6<4B<;"-BHBM\@%@'!4$^XQ%6
PREW_6>"TFJL$S7^_ T<=5L@.Y>ES]Q^&;FEI(OM%U C@Q[*Q=12%H'MU!8TV3)S2
P-XUIA$YS(0N=]#T0Y<#8@DY)#8 WP9$#&3(T5.'GG/V:-T>\[Y?.BBD?V4::M-\!
P"#OS0#U-COFPZ\PMF&@P+E'H-?#MF/1_$70T8"%"AXQRX2^QAM[W%;M'#:STPIG'
PNRY&B<+S%&S0WF>"E/9V<$95KD5/R-#%H.5:S?G7ZZ?12[LCSJ5#6*IA<RK/^6Z(
PW/7CV+<\%G0-GI_[-?Z':?Y=/QB*VK>#@",OC]/L6I5K[#1\#>9%3@;"]L)TGW^4
PK48&'8;-B(<XRF<X9+.V6T3+.D;%;^!?(P2(4DA\5E>';'R5DK\!XBGS_0-=V'=$
PR42,2H:-!_3Y2SH9_S0Z/I#@W, &KR\/M%P&(][;OYM+-M^[5,K;*U&@V)S8N^_ 
PYB55^JQ8>$68O/&2IQ=_B'WM1TSP!U-?4+JN!63^+I0Z=*A5R+ZKVWG;:U(]KUNE
P<^E^U2Y**A;45Y'JD4_!^8T*NID;N8=5"3IDT:J !;YBQS#W-*B?IF$#3*->6D?O
PN1&!\C/74FBE,U*43?=7N5A)^*J2B*K%8AS4*[N6;>?>;T<1$F5ASU([#S"'7*BV
P@+2KJ+4U8@=4=D>R:G/D9RA"]%Y'E<:01F<5*S2ND?AB!3>B(((=G],?0GK4E)0@
PF(HYD>YBKLM&K4[1<\CL5<WZZ;2!\3R;JUD1D^ -Q+1^2L#0.42:6[^M2/@0\SUL
P%<E%/ @>HBN#6NF,3XLM_M(,#"LFW,O$\"LL+I4,Z4HMSP.N9 6-*AGS@&]Q=K;6
P ^7O,'%KT_48JES_+R5W:=APJ7A3ZF ^EH+!ZB _,EC(1MN0IH[<$7G,BB*;#7=V
P MKL?TW$]DFAM.Q1[9'4N,E 5/(07P!%%8#*G[NY,QK_YEM%M<*[L*QNU!0#[N]H
PN815ZN9_SD,!5,DX:F#M6H,H#"'&LI+MCL=J5APP1#&4ID8+9F5S4[O*H["7J J>
PJ++MX5DU T1H0ACL$B4N^5O^+<*V6 L5K<TT2BR.=DY,6,#[IP$=[_$_=STS1Q(_
P&NH:8W\))>-ZZ-?<&"ICPQJ(<'Z8K[]GO?T#A.O+2Q=>&IR<01.^5+/W=',5>C.D
PKT !>M3^ZQJ7(B4=;D\;5"T!+OSU"[Y_9H7%-*(HG^YG9G4^G5%A.88QQBO)J#S-
PZMD&0,:B_@1PZO(@P.8Z9!3+]P9CNLP%)C7?(SW2R9YL7K37H;6T7QU "OD[UO);
PO00RS_.PS9BY&@HAK 9YF\'X--A"T:4L)TN%V!U27XK:L*V#H$+["/^V[.#KBSN1
P11_]%]0&8KKDJ/$'!2$F<#B:_Y>D#\[/8"1>:S.@/HX*?9IBH>X"7Y]N</AWZCP?
P\L!V@&.)5?A%/;WJY#C_L)=0S''7\](YV7GQMH\G/(T;)"WI ^9#1L$IJZBMI(9,
P/(EO$T M-*/V&'';\=G+!;?^S;A@GTP"<\Q=-*F]*@I@MQ>V@X= ;Q!8.0N567>1
PD!:2-@W#] W%:?+%FHJRZ,X1B*BF\;N&8*QO,VU<;<4^1S+B>.Z*)+FUHIV71RAN
PF28 6Q*%!2(B!6_F!"]-TG<M/^#(9]3'JX-XA<J]1RQZEC<A]GN(I0_T0]H]_^-[
PG<9OLMG(0FYW=CA#!\3PY([YA2L&<=/YW"/0[);^[<1TX09/;#MP:D1,3SJI$.@#
P+=LVU+-PS!'YG!3N'\V+VWOM2>)D2G8B1JS%"'J)\,7]+_0.[+N6AILFS3PAJZ#=
PBN,^"6X\X.D7W-([,2/;LDKMHA\GD;+05PEHJ)0QPEPOG8UZOOG\RQT2=?QN^IIC
P29ZI"V NI<G.9D17UC= R*1UV$BK#@V(]Y&BQGS!E:HQM"<H!C"6EL9<MM*8**BS
P64/W#H-538N?(YLA97D@Q"WB'89>LB->7WI*R>BKP_H1?=2SOW)8:JRHK_XU&TS%
PJ\S]FXUZK/, $#R(W)!LBO@W39\.W[^ 0BU*%@)%R"4SQU**)=E GFQX)5,#'$5\
P/8E<O>0LOXRXQAIB-B<B;/KS%9,N&BXYMC6)V==[:?9*999_0'A.MJI)1(+2;(%,
PFT6?W+]_S?1?JB'Y@D7BN.TXA:#RXHVI$GMB&G</H+Y/A.52M 7OR^/SU!\1E=UV
P/<W\G@";&JL@V<@@C5I<OF+D#7AB6B-S#_GWHVP6@&!S/E7L^2B0+6#GD52UULOT
PQYR40WV0[MDTV,#3U<3R3@[\DO6./:H@*GT$\WL)'&>P96N(BPY9V%>'+4EY>&0'
P5N72J'KSTV?2&>>]EC"%Q)N<1Z!=!YUY]O<*=JG>!!%J&H3(:D71Q=!:A8CJ-;F1
P"@(=B9N7< 2\+O<-D.9]L;B\%-+KL9=X-YE2.,3*R1Q<HCS)L9#VZO8GW=YK.:$-
PPOBG"HXQQYY^$TTB";X6[\PF5Y^L)Q!F6D!W\<)&&PG@$0LR="+CYVM(R27;/9^3
PK>-NM&A0[MLUE;LU ;.U74TAR[MG@7]>B[FP$6_5&^$UK N@#S-WBGO7[GDOS">2
PV%R!<U?,9A9Y (A?&;PVL!YZ*]C"MX&'1W?Y?ICKWEM8#+ RP1@ '4XVZWAHGD2Q
P8>7U=ZH!E"LD8M1 1EF9KT!1R<0FMGX0;]H/WL1USR?4" ><5+I"&?6JQ04)B3$F
PT['4B\OCT*9KC/0SHGC:TWWUHT.O14F+*1_MWD[?M9";L'A"D_T(\29F9B;P:C+;
P4;<L%VI(.;[;)/QW7?*+OK]7,A^!* \FE?+KLQ1[;9,Q$!D:U2RRH,,4.(+-FGY%
P%4>\8U\^P]',@%JXPL+E?%J#G@=F2+H&&M ELN[/S]HX0O3[^Q\1<0T0!8?O&_PY
PL#%KQ,T\\9A-(6#XO>VD?PR*V>.9Q(X@T7F$[ >TTM,>9M:MO;8'K1W'LDI'%QZ4
P.?B6B08WT]&_Z^] 2OPF#=W.X+>KL@K+$7/$WB6/D(C: 6RM80_:45E,_) +L>+I
P$W1:@O>SEL+9LTFDD&M-^.><E;VZ#VU-Z82CC_;-B]-<O,88J+$O/=!Q4F A=T$*
P&7E:0+DS0E_:#6?6;J*E=$DBWG-W+O22(TLXB !\X>#NO)AYV1TFUI,3)<5.KN*$
P(4GL"#+/3%J!'W2M3SN#.M_JK8;:CA;HJY@Q5)@;(7":!<J"D4&\EHGID?V '2F^
P;HE0^OKA2FKEB=LEE-9:I]?BN8#P4XL9=P?$BX8E2"4Z;HO&TII#>M=J*)4H.0'E
PZ9.MA'9G&<>*YDZ@S)>]EP(R2 #\YZ >HB,# ^*N,T%J4P"?-D]!4FP5PL,2#?X4
P]+R<GNU"W%B1=R,A8T)2GA4UONFKZX_NCT:1IFS]_NKRKOQ$@XS)D+7+#EK2[D4$
P,;9L"W]/D4YS$A@\0P<JFS01?7%/V;(R)CSFXV8^,PMNT.-(94J>8$!;WX$IN=-&
P2E!^;M0BQU,EK=IM;S[8/7\,IT$>E=@:?55VJ<".V:'."($D)(T4/E]'[ZP/,?%X
PU,.CJF.J-6:A/0B,QR9K/D&$F^?SJ#%-"+Y5;_WA.M< $%?<PKJ8WV9+?^?:QC5*
P_Z';RH"8,_$9$Q./&"OVHW%\\J=M)QGORV='.#E[Q%G*@PLH^>[(HA:0Q.&J*I3.
P?.,HEQ=GU\WN9#JPO'0(M^GP@.B9<0E\H>\"R)'PH*//ZRUW<;?@2>F0Z8AAU7F=
PX8"ES<B^P;PV#5IDRWA0XU&Z5@GU!SO+6"H9P/3R0*=+96H!PC9'KJ(22_3!!FA5
PJT8?B"*R5U7B!>C-:I=-H##59(:>=?)\8I;*^3G\XD2_#^'QDX>XBL* Y*-WR!]O
P(W="!8JH>Q.=4RD+G1JSSNL&9[E>PL,O@B*R1+O(/^)AZ=<-]6Y;T[E#M#1Y%T#=
P)'6#:#+LS9$!:GO_YNO(:38""XMN(.=]J/VW400Q'"B;M3U,=/++EB>"$2P&#A0 
PUX%_&(O>'2*V<8B7[M-3,'A@]D#YG1#0^L7Z8@KI>(\M.C@:/^T"DKL-" =!3/&V
P[\_?EMWQN #%O@3:(9O'RI'W +J:9]EDRT3/7YAEO\>W!=IK_H<*G:%OZI<!V%Z:
PQT]U?PO3T&4<MH4FGC"Q"PM1D@81WR70BCN W8D<[!EW JP<&;%8(T),.Z#61X-4
P69?0A>'07"6,@UJ%11HXNVF(6PYGF>HKM"NQT46AVYG'T+&/&_ OBANYD5IGH-'*
PQ]5.$NJJ.GWD4;^ @\-*],/*,E6_Z5RDL&V,EW,JIMKLK36U']8DZ4VF%_OFX7HO
PG4_T= 4XPJJ/Z: ,_(K\9K=_C=J@F*-LAMX )"AI]L%39E$1$&0Y4TT$4+/0\A^Z
P56P-EZY+3-DP5\R\;DF*T%=T-$ ]!X15L$.DT:;N8TL'U#/ ;W0>2T]"KDL+R;>>
PMVH&*$I]S27'IK@)8%#F*W,#2K+T%K[&5P0GKVC:7C/$#S7/9:0;.F+*B$1,7C >
P_@*Y7O233QDC/*][2M>0SU4_ T$VGR'Q9TG<GZ^Q8Z#N"NH2X#W&:[.@&553PV07
P3$]6)FS]O0H1_\PEW\>]G=/F%WY6L_W!0V9*<ZR?]PM%;<C9#ST=P#G%D[L<V*C6
PS;\/%@,FGX9))YV+UMX>HL9(*) _+/\9R#J2!C@7DV.&-!^'T*,=$ZN(WG8:.^VR
P $KP:>LN@+MUN83QZOPFW2]/\5C*ZL7S'AU9>POF,6P;GS:[.-C67QJE0C"@AV?Q
P<H):)B9 +CJV>B%$(0FX[@6*\!8"NKJL':$E,NC'+D6RO2*>QYOZR8PNC!WZ#4ZP
P$I&_&LJ7_IA5&(+UWX:KB" .L7H66FPIC949(1S+;6&>0J<5:F&#)G088M>S+KX1
PRWH "+,F*6*KW6K:92>A(@$Q>W1@FFQMJYZG=K<R\ESH'2O5D9!?KN1\L)@]=+34
P?8?_7B[N!NP$-J0^91++2?0RW J=.OJ7X#;1AK7Z?8.Y[V_F^#A(&EV),*2LOK:S
P@L]=!OU[R3\.X85%XJ]L_HVAT_,:L(.='3A,4CFU/;"-*?9F<.TG)VGI22[UXH_8
PV0U.?4_8Q])FZH5,\6Z^R#H+H=/9H3'>H,*>AU?$7Q9([5&QW#7NR]$%9M_HN.49
P7?8B!"!1%8/P;"W93D?F[\WDM)QT;8+?S[RI7"D%.PX1SI8N[VMA?K!5F<<!"[!N
PLF4FC.T*K/<C,78\((_E#9M$]#-!?^IU,<\H(U.54-HW>J%U5H):PU?5Q7I)P.#G
P6W<>6^NWR]#6>T1WBKDA^$,-6%2N6  MFIK"#O(R$4)Y/=F9>5/[6*1N9M*@,JYW
PXS;KLE11O0YZR)B7U@BYV4 W)F%01 <^.VJ[I)2+X!6*?Z155T:R:W>$'U24BI@1
PX]1E_Z4DVSL6.8\#32-@$G9[G1;PAK;8XPZMFX@]'OZ+<O9[=BN&6%'7S.64M[*[
P/YN7L(GI*!\U-&&2,GSB\.IHTNVM=EM=9U9MOO<J*+++)@_/9#L?'B"B:E(!;*SM
PR-%^&='[0%K9;70"D5!&N_FS9'2!_\1;4_W"G)Y5V$9<6&!%W_V9U:10@^&L]D/X
P]1JX>HYR0[>7X5+I3-@B(DRB-<5="CBJ/A&VOUJM*!@/Z^%]B<,N/''GX##_2DN@
PGR8&.6"QY/(4C*'NZB$;BQ#EQV@9%50(S6PF3%&95XM@J/*\V(',T\])@JW7J\\X
PPF)7^N 4W =DE1*52G1F3 ,$$/B')L=7@A. L9R6-75;8IUUHM=S/18$WR3>*Y2'
PAG9)?4 *'<NBI$Q!%\E5.^K@E=M"!E>7E:GB8YI-]VZAUNH9H ,,PM:]_.F*@U;%
PPJ>,D/H8R2;%4NGDQ4 A)Q9V54"-BP8H%Q_8K$9^  ?EGM#\M@\7+@:B@7RH* E!
PM4;.*?W\TY9BDH9W+V%:BPNUTY#I+6-<@49(V/SWB>CHL_$<JIN>)<L%$4^WM,ZW
PV._MGR5A;7!B>R2X8DV()9,<$-#/N/[_B1SB\-\$ ERVTD\;K.D%8[KH3)1"E+:R
P%@.O-,.S3=VO[I;O%2<4B_M1E4DFF)%?(*R TT_#JLK+J#1;'KHX>F21NR,'Q?BX
P#+MCU7ZS:0H'-;D#8_;^ LFE'2W" ;$KT^&&%<UE>_4Q'MA4=&+6XDDP&+0038D<
P@LPFE#*R,ZH!HOS052$\:'<,5^A3,G2<M^6 Z"$3N]4;8,#W<#"BE.;.LUW4S8XY
P&Q0S[":([&>H_-,FPX]S*@Q6+_X Q>P*18JTQ$5!^=I[X4ZTHKH41%^U7;A;><VN
PJG,#@GNK=H%C# //VU_*M,^>/HG/J!Q,3B1@ !#,?)6\BE)3]L5<.I[L1P]FMP=Q
PJC98@W\#%O>._PZ-T47@F&U]OTLSD4H=8IZ:J60HZ&H2FF<*U%I7,"30F& M/+%A
P>PK1,;8"2X1></9Q#;&V38UC+)ZK.#D+(=08L;F$(N/F6W+UB&E5D=2?1T#L -JJ
PNP$7/5^*D<Z\=J"UX\H,>,;=KJN-+!*-=%BH.(6\H6Z*9^6YT#EA;0Q3F17X.C4A
PM;^FD9:9K?-35WP@M,4]N[.[MEY@'H=:X L2/F5P18#6>NN4T5%;RK9@?(/J?+'O
P=.ZF[@&Y7V'9LU?JL%\5XJPL3*SA:UN.11IQ5U6GASBM)HT;F?WH5R-HE?VS.NKF
P1]/*LWR=_W@>?GK@NNAUNVD\Z+@90_E13Z;S&E)^]DD @9L39LN7E:$#34,<Q4SS
PE5)S>>C%A% #;@"#KKZ,DGF,:LE\I&N_EMWF@\K!,^W=;J@3*XYCB\&Z)(;<,]\L
P5:R4H7 ]157@\!B DBSF7O38I\XOM>?;[SF>YN\R9ARJ0\RX,KS&GT^9X]3!J<AP
P_ZVZ;$/-B>7:]>GU #("*B:FPRM"%')N-&XTFE#&2H1"I^X@RI_7UN]W'-(=NPN_
PGZ?(R*FU%2D2G)&A,UMA1[MCDB+FGHPYD%/^@7T7"*OX\R30!859F@ZA%SN*Z>'M
P@9Y?7[YS=#X-0A9_)M7E(7SK_.95&AXS0V;<K;9>LK\JBY,RF\3]^,"P=BG27 ]:
P1HK=)!Y?A?@V;N8>341@D)NI:LT84N\<30""5L%-/(?4"O9$GW67H@\"F*K)29,Z
PPGO*Z?QD #T[Y9^7\MHI3^XKI85:DS,?3]MLZG M<D)4NY@_W8W/7C/EQ-:%^8G2
P9+8Q!V %9]0 @12OR:MVL1+_?.H[/2.)(#LGP6D6EFOATN)^90Y!GW3-";4[, ]P
P3"7HL-F;<EX)7]'0*T#[3(E]/PT.2F$H./N=K(%>NQVRS0 @*%PZ>?G8 W(F^W=I
P]<=IYPS[)V*MP/;C('*^S,^@JY"5*J8X0UUX^ #%=51 %]ZIM81=="R8/XW6[9)5
PN@Y;A<\(8&YRMI X?;?Z 4<@F$F+&HU_J^I5]I/ @FM-!J0OO.JOO 3RMH7S(VM?
PO"01UCRXGNOG=<V$\%>E0^OEF;EV PJ&:^-9-$!VPZ[ZUI*.]DMC7I@Z$.D)&_#3
PJ],J[T1$P")5O[[FE^!<7DZ&+,<D$OT%[22N@9B[&B@DD:!(%7*(?-8'!Y56X7'*
P8IQ_5ST [B"SI/ QBM;TK\PV8%<_<Q-Y6OU5T")  );! !B8R&2@;H:[!1OK&9,O
P=YK$%U5=SJ>^VV+GBCAX;>>HK$J_%77[)S26YT*#81&>Z]I#E5)HKR]Z/^BHQC$W
P5U,Y#RXNRV.(2^';DT* ,5^HT_Y)U;RL2,E-OQD\=LN!]I*\6_+A?/L/4.X/CF]Q
P3Z&'B6$X7_+DR_TZQ.-L+38LAM0"W:UJOKV[Z.+/7 W]HL';]VVVC#'>.0;\1+K@
P?$<X\EG_^T>-IC24]*U74?&AQ1N@.1DLL/ .  G5F1662MHGL-5Z/X;@R#F?U$Y4
P( MW/[JY&SZ9N6'&J+B#]W.[=4M=?<9*W],FB0N-ZDR\E8HCA%%$K6B0AF"LCR]%
PKN=+B*\4(Y5UM3WVAE<4V?/!6S,%@+3@S;F.[HR[(AV+E$'LS1A=;EA-K4&<)O2,
P(;(\DOOQ7%\E2/9<VN_<9[])08*Y5JNV/** ,[.,<CB1,;)MJ]C*1+\/_\!S*U3>
P$9YD'A/MLU?[)AKZ(TF^0QX\:KW3RBJMA#J9;?3WC<8T5.PB:07;AOMKGNTW#Z)8
P#Q8[D9Z-=T7E+3?+,3DCUA3ITI7H)3%JS#4Q%*FQ- @Q9.XY*QA*!R4M.00+Q2]T
P@!0=U_9CB^++>/E6-Q>MH%?^=1)43C@ZGFB>-M,Q!P\=5V^J(+5N3J>[AX!/[U:2
P6S3B!> !O(^4F?5WZ?VIZ"T, PIO@U=X_NX;(=KT;C^!MV^XP2^.+*E*8R G>1,'
P[ER7?;+0^$!G6PQ"QO0Z6W^G@)ST4-%T@!QM(H$EPVZ]])0 8HWTUQ5EMTUC$HFE
PG-F8#5\MR/(VQQSU)1>&+5K&H@T;#)_K(T!NMV&$.E*P(3G^KK)%V@ILXG!L>WA'
PS#\8=6%2&LKJ*(H@'Z YTYFS7NSU6*U+@9*)\\DX6#[],#9R9VDM<+LW^3F*$6"P
P9-^3:&!/6Y,QHJ&ESA]E#->.BMN3K!H=ST< 1VO<9\P#7?L2/O%?QK-TBD:#5['D
P%R)^)&-$9FX^[C_Z"OEZRWT"\%0+V5QRC+E-0']XB?N+TS.@Q(!FHM#(CS(O_@4C
P)5:01[']MC*2*9,K FG+'IVC44]2]]#Q9]+Q;#Z>:"F,4^5V$Q1V/VHI68-5;KT4
PRTB-3'#U"9LS<SWU&;-"@8?@O',BY65+ZQK%!\0_RG'+BDH(AAZK5D38ZD7T.O&=
PW'&:S&0S!JL]&HS/3J0STKO"&I08YAYTDB,.FL6M4X%C#-/'X9DG=$_']+1N%M8=
P:MU<58W!6DR5,J5-B)\ED\70#O4%[K:._NY(HRR%4)]GL(]^2NI=T511]DF5+KZ5
PPOO>%E'_C]49[Q)IJT</FS[T=;F-8IX#2FXHE7]Q:XYN]55W=Q/7LW]1EBU7 DV?
PBFC(Z=R'XP'J.P5V]%=^"MJ.*K><(N5O,*4JB^G#,+.C<P^FO=7FG7_&@V[#$T"$
PI<YWR(^93%K6,)\]$E"'+,Y&*)PCUP_-9=CHJOXN<7TO3W8S9]@[HZOSBG89P)48
P[>M )[&^9Y=8Z7ZK8[:G-(5ROPG3E%(W(2ZDJ\[00#9=2)SAL;' )-ARWA+<R$?3
P6!:7]KUH^]^D':^"+6.%P&S=:,\86-Z(<C_B@_34$.RVIM$(OQ<G#8'?C0MP[5M>
P[O7+3-@$EU+&4_OZ'8@FZA;BDI^8$LR78=&UU\Q P=] T >RHY&5X(N))T5:!=K2
P/E093P)KWN]ZW&0N2T2/-FCRC;]R2YG86)VY%(%:P)Y!C^H_=DO,D_:KN9[<)W_H
PN](8C:,34"R  Z163V"HMD+I34<3AI+8)#*2YDY >#E_B5&.@S53K5V'0+0E%C#R
P3RWZ _7(U6K=''Q@ ^V3^ID^AADL&^QN3?ZF0)D*3JZ+6"X7EH\59F4_FY4II="X
P5XF"7Y!@?QAU33]Q:TP/]OGM)>.GH+<!Y+,/X2Q=4V&JXI^:E$$CDDR.%_Q%EB"I
P.1?=GQA-@[.T\9DDHH R?0YHP+%:27:4)HPVC!%8N+F0#G2LZ 9*6\0)2/C@Z^.<
PPD&-N//62Q8PNE=Z0%<-#0,<!8JD;#_/P%O1_$?_V]0M[#>0]!@&-*N<SSP3(Y5(
P<^(WJH43%7Z$7R#HJ)]%''UL%$PS+#K\?&H?SD/;L6797\4S%MVB[LQ!%IUN,1FB
P["'TL*8"4Y92N+F;4'@&WWN,B+<&H+:S]J L"\<!9%3$=6"DZCH[!5/]IU)I%E-G
P&>:ZMQUY?+'[LOJJ/GE+J*59?C4'MN'8'DFI#Z"GRG\*#"K)/LRC.0>\)B#N\QQ1
PO$]<A=O F[>]U>:]LMD6'YT=>,)RPQ(4J)J3!##::G.MM!*^M'Y?@XVW)X^*\07,
PW#%]+P=PB1YP[:1>@Z^DR1_[%^;]B2S9RQ:P"P T@3 ^.#_:&_ W@=19;KSV*.0Z
PT[L6)&F>L^[+S@/Q4J6/?#DBGN6;STA!R8FW3P$]USII!29FC*J4D[LH*4>!#(7C
P5-8(=,[LOCLE(;6= WK8!II^>0?Q^N4-I>.Y)AK XV+8>J6F9<"VP+?$!;ZI0:$I
PC!6OD\79+9*5:Y]?HJZOL:TQM3O-42A 4E>0-_\(DN$;[M*=>9L9M-=?D@(ETZ7S
P%TDQLIX2(S:OF(JR2W_9P)BJ/.>OK9#']TK+Q\&\'H$Y8H0)HX+9A _FWK"KQ%*G
P5[I$*LKQXD. 00RHO]+Q6L9Z\O":]DVSH,V ?\0WT/;QY4>-=4GF(')\C%Z59/1B
P@C]U!T<]-91HP]:S\D@S&Y_PDUP.YLZ9=N:2);@]M_S3)]390XW1TX1^'CQ3&#/(
P@+I)8K6G!MX3M>E?FG 0U9R]OYXA0U%H,&1N/0[##0I=M/>)SO KR24C2:0XQAB_
P'Y_"?K3*>![=66[B7U!CV\&IW,%Z.0I[F5)2+M':\QI@YB<^<[28P^$[NL_>\1#.
P #QC9JUZDVH@$6.P_:H>$ "TGSX]'="0Q9"2#2A7WXR[@?CIBT'%Y^=4."YWZY@;
P,<$9X1H;$@KJ>]@1?P>TF%V%B%2XY&T#@U[TRI$ 7KR<$ U:DCSQD9.&L*Z*2OPG
P[#W[ Y;45+80+8H(<TT0GN8.1SZ;KSV]:A^$0/8\ &I7IGZNYC@_G2QNEV(T4 ?]
PF@ !E2AR2YL??'[.9/ '^.3^<JK*?D]&0X_R 9K:G3%@8HM3:K_P70+MT*:;X#<F
P9ST1^ )H6_W:9OJ)05:?9..*@.RL5)C?SAM_Q\8TWW />]PVX=T>QH#7Z PM4.(#
P$J07\8_":V#K*ZLI<2L=9!21VPGEE(+1\,\<I_\-,Z/=L%8*R\O&^P/?7/3<Y T+
PGR^ZCZFVLX,6(\B9888##4=,F9<:<O'45<BQHS0C)MF5-L:&G7'_\QZ-<Q%\J%S$
P1#D6IZYU(-6*;*M]<(PZVG>DF[IRRI=UIX^0)Y^CX5>&-%5LGPMR5?\A!X>+10W=
PTZOF1"-K>CE?.5FSC4RA38=3,(=44R[<QD .W[NTPS-:]ML7=8:ZE!6)-,(<QUV'
P?!R='::P'FT B<PE1Z-UF\6O \X3D7:8?/M%VH?J:$3@O3NMMX4Z[?J\-.>VG+%V
P#[;'K.7%W0:>81+[5/L*.^\.']8F?,QI<*9?:_/\RYKIQUP^QS^9P5%%#Z6$G1%$
PRHN8(%RHF[S#0*429*$9"&.,W_#CG#QU+RW+GV\C\!"3!JC!L>AM,6]@.9,($S0<
PYS-4EY<*%H;HXMZ*I:$?#Z3.V][!B!C6X98M;)[0;Y5_&4U1XQT^BROY3O.%G3)R
PQO^E <I2UA'3C9F93:=JK]#_$W1A/!VR(%^F.I+!CZ*UBJ-6GT%(9->7QVDQZ#B^
P*7\^(1URFP4%$-B,_CK[C$RA2IY84DRL',F*81;>$0CZNF8V(U9NO0"9>!),  0^
PE31SX#E?=P7X$:T7[P:M6[FZ(;?B(9*J_P.E5L+7')!*UGYKJ-72\19)H3U6P_R<
PV8>)B5Y:0^N?I:(XD#-LU 0KX?1;67TWT.O@NAT_8"UA(M_;B8KHVL3F7R.&&T!+
P;#=WXQP"0J\52](8 N#WI8B:NAUY3$F?$"ZCW;NO-=WD6J.$4K^!UY9,9^H*/.E4
P?2=DRSG@S/)OH1SZ\=(@*'4F19\QFLA<:*E5\/24L>&#%F8'-4!NY*0+ADRLU:W4
P[)SR'5CG[@;K&U>9129!,B6"PLY=;,B2I">BYD!E^VMM!)[>6= UJ'S73V%3@;E?
P\.HE5ZJV%MFZ)*'@"!9BOB VU4MU N03?QGM24Y43HG[S5$E+Q$FQXMY%.0(I_HV
P)I(<]/+7,T6!L&@N.Y83NP,T;[P:5Y'2'ZP^4N]#]Q6TE&LKTJSYX \">KK=NEP9
P]!R[CT7SGUT#N_($"HEAGGZ?6$]18(COQF6B0[H%)5<VZQT'W&"T5L;P6,SO(_0A
PJ@1'Z?^@A&-A%JRU[I<?A.67#<Z-T>"#9+A.S -><4TL\390B9)(6UR['L88H&X2
P:9/:Q251N!BHA?]V=\)_OITHA)\=$ENU_))]I#*6HP#PYD.[Y1PSVF0Q&!'D-98R
PK+6SSU7ASYT[78@'1*>LHV?![*#_][X7K>3T6%=I%'P.= V,!^0%!59]7DI1 6*)
PB0]IM*^I;2H;&+:K/[*TWB]6=6CH4&1R/;C\[L)4N+WBPJ77_WLS<B#( K!/86[Z
P;^7EOYI+9.>M. L'M!8S-](LFB:+NE?BZ_:W9#^L(\[&ML3\1D"#<$/9%9=!4"UM
PWN2X(?IQ$U\ [;_C]K!3X^O82V.V1B#OF%M]NP(VHCLCE'C33R7GI G+BE,Q>SIL
P'0#YM69@G0</]<FW1R1U'NYEGRT@;S9J8;6'[M(4M))Q"'8*7)C\'%_X =$\$?9W
P(Y5475^UH5'=XOH,@1HG#4I1#MN%;R]7A:RG*YK'+(B/BBUK?RGK#1'GUN:<D:4"
P#+\Y",UVM2ASQ:!E"R2<$D2H60UD=2FR"7&?*-E?*Q\^'0+N<&^DE!KF[+ DHY'A
P72_IXAN2'!XV98IK0T5,SS5^T/3W$HMP26NLUSFXL33*7-XHV@_A216@&>P"3\Y=
PP0UNLAH<90U=Z2]45=MKL@S$)T:Z2_BC5.TU5-OJDSNA=<C%]@BQ@4BLZ0O#4\D:
PR =</1D:.[' SMB^HON?R2C':Z#$%7QOM(SPAW5?\0>*\X2(&Z[0.[[Q_'U'4SK5
P(A-4P4:I&'_@8VH_IUGZ<LIYW;-KY39A;IA&,;O*9"'<@$.T>YG^. IXH+?$]28;
PQ=UXK,6AY;DBF6-9T?+Q2R3SP*:%NI:S;34QP[0*G#NI>O4@J=)B+Q1-+<SITJM^
P3&/L[URO]SG8DZ-OS#_E*^;.C:R; </DNDE8;-V2KL4W0_,V]<'#^Y5H;#*"25A/
PP7G\:R^J%K(DTGSIA*/#'")=5@RZ;;U868WG\5Z;M/+Y12E(W!.A4-%_*V_:N0W4
PT11"AQ9^!(49M@+AK,N# ;EW\E6YDK8)B;8,5@6N8!(F9%:;/F'Z9EVX?=9^B@9<
P#"[5W<AG<2L;YILSE2LJNM+I0WV(%NE[#N$K^;FP08DJ0*",#Q$+]W]55L,T <?^
P(@9&[.+F_O2Y@A 030?K-XQ+,3Y?;NB,G1&3)9JV2 H3Y#_#/03V@XX<WZPL2JN^
P(8',W0AK#AGA#.!*-6)+SIN\X4;JR.D(@X^'$OA]P)%%>PJ7N\>1R^7X!M5O9JON
P?A;9?V >=BI7H8>B)WC@'(V%L.P1;L)\IWT:(_89RA08L+0=9-HK?TZ"@W,"PV.]
P[$>?U,^Z2,Y0L4#WXN(B(+SIDS5H[KQ9=<(E_R#6MK8(N?$*&4H@,+UAQN0Z6\,*
P$DA:?[PA"EM4A<%:<+7H#SN84@:&.R>/ K1E]T5P/G-K4(ET\A0'N2PY*;J:7F=/
PV%7F^,6]-JP<6+07DE"I#&>^;64">U=$2?+%Z%U*A\4RN?#_^8 "PSOIT+>,S!5H
PI_K9*@.1A.DWE5SQCUVWH$DDGH4V 2BQ@8UY@OVXI/M"K0>QA<TC>B>(#IVU)0U5
PS0Y0[]D8>9S%G7885WEO@6/FQR\Y4=:YIW+4'GZ0#KP%.\0VP<@8%4-<2RJI"X?A
PO0<T0/\55#3QR 03"N15(%J%5)/JKY_@\'NX?:<U@##5)5:BB-4$(G%K&&'RT2.[
P#_'>AU"DT)X(2/9G'8;Q=M(-9.VQ-Y71/2J=;C91,QE[,PBR/E!&,.POUI8M:[!6
P)!;/Y<,H5+'8PT:*AET@M%TZ?T/2@\1A+7@:3GO "E9<6IOR]KE]VV+M;R9L4)2)
PJE("A#@L7OTA"0355@RCM41>NM!+XK5D./2#&2M>B&[?:U8X!]G_:UMCR.O,;Y;\
P6T+,#IC=U"T$,(B!A",[KV]9QPU[7DK!.Y$@PW<NE@YL V+H2Y=<7F1:S*KU++N<
PW&#HF;E_(>?GW7;'X6YP@CT$W@MY@-6Z1#=@#Z&;79KQR0J68#?"\,6ER:/R<QP0
PF0??.>/J P"E+%W/,SI/ASQ3S8.$8E(&>F9X[?8:)W$"GR!!H961KW)@*10NQ@=/
P%O;2+.Z'V2%J>C*=^E1Z,01"6$9W![I4' #Y^,L]VP0YSA_H?>%?JHL<(;%L/XV?
P;'X%),9%("R!<CVAK*:R8B)MQJE@H"?V2R3)\]^(#X1ED_\A5N(8Y"$CYX/9SNBH
P/HKVQNUJN0F*TO!O-6:S;V;2737VYQ5<[G?6 +N-3AGNR>8G-P45,N <[/.Q"5I-
P\@70 P17,Y(8NH[Q;V'F"SB4."O R2/"$?$212%49-P!,Y6S";VT)'07@W;JG4UI
P7B>\7$V>9C>BV;%2X8:479M%HZSM]2O@T25DW;7[041$^$C,'R5R\>Y+G^!(-(-R
P4T<3)3CV=/'-U7G#>PV_\Y92O"AXKR8GF+^S/N@\5C9,8JQ8AQ:,;(6!G@"?.^"D
PN?F I=].UMN][P[KB(X"RN%TGAG=NS*5]ISW[!,X(?C4X?_)7P]0^B-(^VY?"BVX
PSVH"N!.RCZ,CJEC35K%:94P]<!&@9K/3P+0K@L1D$RU8LI#3<-XXJA$V-A&C UGH
P_!)Q\%IH*DK?YXI\7W03[YYH-%80@5"&'\1G) -NI,>)DHK$LV6!!V\>^S%65]B@
PYH@8CE>K,),OA@SO-E;:ML?UDJ6N_S$9OH/H23_]A'W15$=%4Y,VHG'!_QTKHZ#Q
PS6L*7)#-1[F6+9,DYK42LP 9'CLPVVL'7>F/]@$=<W[\6C_FUWR;KT& :#=:](*G
PX3B6N>$C[C*"N&6X]]\^4HR/#$@HH!^J]3ECI\W9]-GH;'9%-J#[>N!B*'(KHWAD
P&4AW08VGF)P^P^A;_KA %HH6G\MO#QQ]EP!!B5"K;6G(.(%V#2N_+TTML&-^_#".
P/;[<OAQMGW\8NFC3A0V/[J6K0=XZY![T+!I@VHAK&C#O_3V!DS/^A%?6Q*WD52F?
PJ# L_$2F?3J9<R-+Z!1[Z"@_.6U0C&(<AKVOKW=W52EO@>2'&U<D>A<7J+"11B()
P6V1:HS5+<* %\26</:-EHQEBX8LD"?/:Z(A5_)A<P=4*+BB1C%07WHD"?_]D^'Y^
P2"(F=B@;,9+%T,C=G<X\R9;^WK!@U^$63DE_*78 ,.IVD-\,C331>&N4(-?L[K$6
PC8I6.*6M*3":C;,Z]:>W_2O^:E.+!MD'I<"LA4^.'^S-M:"R$ KH[S[1=+VI%KK(
P]5,2AAC>MEU[>&F[3M%.0"6WZQPTMD.X=AR/6E/3 4/*3BV,F2&N((!^X';*T%?M
P[9F'TR!Q7/H&9 &50,"W)$Z77453;UCW-F.$)_ 7'1RD5W>'+GZ:[[0Q/[0^8*A)
PRH049@\D8GQUUU5Z:E>/=]4A_*%H:,3&%(5"EN07PR6 3@CU:!=;O]14_7YI7K9E
P'TH.J42ONU=6_^(M*;+^@"1$Q1U_3X^IVE300#D1//Q0]11,A8"ET+_G"2#Y(R0=
P6N7\.>+;#XB+ <*\^-0)=;>+PVKU&'' !HJ.0LCV[<(:H1V1RY\"NV;_,%<LIVM:
P(Q;?$9_,SUVZ70/[4&& 7A\4VUMY0;X.0<Z0PDEURF)BRA3<KEHA7CJ75.E^%<(4
P<Z!>(/==2T66(L8QZJ["[[%Z</^==5JP\P]Q;J<N7AW&T/7L]2ZG_@2_ASSGC4Y 
P#T0@X3DA6B9.O)1@9F$(D5%_K3(/5#G<S.%^:(-]Y6(?_N@,H,\MAYZ-)K@**#^\
PJ)%6@;B0^ .*=^_8$$[\G6C0XYY8#,V)=;9:ME%RS_$2E!.>.WVB1:5UV]4:29+#
P\EB 96&EI_;]88PY,K%9L]#'-CRX$:3W JUHN70Q,F'S6&KRE P,;Q5JCK36_W]+
PVRT*E="*@ON3 [207"9+L74W#(;".5TU AH'Z?J$SV05M.*D4O:"RAJK*AH2N?%H
PKOOYP+<?SA+*W1Y=Z5B*<E@T"[T[I\!B(Z1X3HQQTGRU0&X8>BF)^ZN,]),,5DDI
P\B H2VQJ'[@ZDOJ',?1G$[!8NAJHMGBDN&E)=/SK?JA57'^B.CX"O76T:E% SQ"E
P?%-L#2K<G-JFI@0A;9M $GX9)N7-8T7R18P8I2&V](*)G_IN='*([,ET4)BBTUC8
PD<.>3Q&TD>[\,F 4EP]&W_H>,+Y5!@LI"NK$&+YDAFR"72_4UQ'%X3Z'7KM/1>&1
PPC5H? / )4I H%#4*5;)Z_F0'E2M"-!((05UN:8.8<D$SOX&9]H$MWTQHB/NE0QL
P\)KT_ 7U G7!T.4LXXX70ON)B_]_3_0?>5M(4&D_EA$MZ!C:# 85(_G :F9,,[]A
PRS=(UHQ',?MT14.!1\'')Y_CB0OIUO@EGG&M7-H\47I\/ $C[7TYM8?6F/+H43,J
PEK*])^NMIS#!7QTNJRJ8\&SINZVY8)_#XVU1E=Z-S$U,.._%/U"-$/"#>K,++M=1
PL"3:WCV4R8!3H%O,<DPC[S8R8>=O1Z7'#YNR-X#$\P]AD[L5.OLV(@U(MN>')E?!
P*R).OO:0V)%O>)*H#V"\NB:97/Q@:A>=S^RZ2;C5SV=IS#%A%*U8NIO%TC2U;'Z<
P3DT^6OL!^I<E!"A/QQSA"^2]*;)'4/A?(P%V(EZ,5]#1?2#T9J<QN8:\,6BI<?M^
P%&%HAM\&,A$.*&12+)HP'J%T_]+OT5X3 K3'LKMA%-* 7B6G%" V%7G4)0R'_SRL
P,(\L5>=9!*!QK&$"WZ3G -OG,4U\X-#37U:) %'S69M)[I\3WF@T_DH2'U?MN?\4
P6G++.,TL*!.D 25']N3UZQ-<AN'"-BD^IYH96A1-'HU<GP&[XJ),=BF*71NN+M')
PV20+M'MI>A(C\(_G<"!X9;[X6(5"L$\C]KFO<F25;K^E#B]=!@"6-HKA'4K*+A&V
PL+"C/)02( HRA1?GGH>HDMK/2RX7+8/!Y;$!><S#V4U%4R-^I<GVQ1[UU2*C(%.-
PYWMV,[3!'S)5.2%IWQ[% 1IC+0F&I HV/+VC@(\HLO%[@8'5]='8\%*2\:P4"Q*-
P2M@&YQ/+BN,&L2S&B+Q>;ST.(-6<(WW-!"+1:\R#\N+:]MYSZE!%5[,-.A>0!'\,
P8QG0DEB0>)BBU=C>,RP(^ON"" W9/7[/I#5*/H<6\%.&OKRJ3AE#WAQ%1GE(C ;%
PC[]<=D&YG6U?/L"*[@)[QYF\KE+).))6@'DC2(%=E G!@.F$4!:D<Q!<E\&1/]P&
P]'+B!>P,T(Z6+PLHCI$YU 'MM'P1'4Q]JMW$7!K/05HNKV54F<UK+^& X51/ *:B
P;#2!'PHI>GF 35FA!K1/T6^^0G!4@JV:T1#BC],9WRT9XPR*F_UO$7L!+G.S9J:\
PRL)HD?Y83P[EP?JXN:GN8;]%=:#?>+ZGG!>=_%BZ[=2"+AI;>VUC(!_=M4DCF9Q"
P?G&1=B;/&H')S<?)<R&;'P3&ABY]X8)Z@U)_PWL>[V;DRH +R@$YV3R.!8/]@.7N
P[ZP36]A2Y#MK<>-%FY6",QV#C-1WDY_]M\V!$UHZZRL]YF4'-J):!GE39^B.)UAD
PRJILC*>%3T_PH8]AUDIU7+LSZD4+3AL7,1J53I6N="$]X@$9^QM8BC+^JS1C7]\N
PF+$Q!UF&3U'Y&,="8F,?@:/ O<.T1WD#WR--$AU ;H" @7HEFHD[#>$7QA&:5E>_
P*\4"R/L>']5,-^1.#!5EAZ6SVS5IXH%+QC0K7-H.5A\H&X4<F]V# VW@ 0NHE&T=
P>-47UL;,W>7]*TE!TK*8%8)>D;3%0LRTDB^SIF5AA9IL0G-,/+'*10TG-ZTP>_@1
P>HG!/XQK_#T%8M&Z\T+<$AC  ZZ(QT.;&FD-P3^[(^BJRCRCHE>0 %Y)DL?KY9XS
PP0DQ7P<BJ78721?;3\4HZ2TJ!C;6D\O@?NFOG<'+FFG?./\D?Z&1+4'2Q4X1*,I#
P<_,E0DG=] >*K3HS\.C^[2O80RRFW$!*=,K!+EJ9/#)RW[-)KIP$T-KN6"_T::&;
PM"8T SZ1!79*H#D71\:5<C[_9+*A]S,P<L,)&\0).9H[8X_N4\8=SIY;V53F[;IJ
PTEH41_FVSGFDZD@U8+135FH.N5JI<Y@;C+YMODW.(DWPUQE^[ D)C8(2FCR7V\Z=
P4F(X2_;QG'  T!\2Z==(%IU>><>9\O?*DVW>!.?AD8E!Q\U5W@"#I 2#;_.[XY*1
P5\GA4ZU'@QGR0UH]LC(;"Y_BE8-I(3"\:]D40_-OV[&J4UL.K;QIEV[&/;@P4=:Q
P[\YI384,)&HN9*\#8I8(A!D-OM8V20X:?EC&^2.8\)D-Y$G*F4-,+DNX/Z39J0R9
P&(%5%C14X9QKHYK,XC,[ $(T[M2C^;^0 H6QYN=&#]L)U>_5@2K@A7)KBM /(N=#
PMXOE( G@Y3>]S+41T[9K8:,\X-A,U0*N82]$DVCL<#I?_D\C""=(%O]</[X57K<D
P*!'__@#N3<YO!1?/E#?34_<U60[B2O 8J+\:;&#?73#%_20D,452"PP-\ 211:>R
P: 1O>:\>.<D,[,H)&55'IT#G=DI*/'((,@N: OYV!S7@=G*@%3SQM-]6*-L9LC\0
PZ7 \GSQBYON0H%RNZC4^HNH@D#;MH'F?>:7=W8JIVH]EQ?M9UI/U73F4.CTUO(XP
PTK^HJ,WC_51O^BC["AKGC"*<')4.SDQ>[UR,WRWKY77N(XBA;\ZE+K0F4#[VFJ!U
P(];"_1BV<>VJJ2-(UWWB%>KTSI]Y<"CD!VZOPH2%\X_60W%.G&CN02A^WA* +]'P
P7IYVZZ72>0XJ%1&.;_$4U7#*-)-9X3ASA!K&X#!,IXAQR4>]QX;!<[W$U5\:N0*;
P+K,OH\$=$ TG;#!S5UQ^)AIS7"Q&SS<R;I(K:]0,:7%9/A5>[W(U?,H/-VM]+*WT
PQKIH?R!6.?,1@%TGJFY^_%QI9"=;*DX0Z3'!Z%#S.D-#^2/6!)'JFXH"M-/706?3
PLFFQ3J+U'X'0_=-V5J+43.U,SW3<907]]7C[2QZK5>,N<^K!*0_O-,=3=T*-CQ5K
P&_J3)ST).4ELR3MT$WA2X-WF.!L$Q2608<JNN<WT8,C=!J4?99^6HI8-?#-02V!-
PT"S<ZM4;GG5>R>VAMQB(&G"[;8FM$D'UUJF.#6I8BS=\L\'THP,;9V6"-.?X3/M&
P'?0MC^.Y7A"=0%Y!]^_C8W+)-F>QV?R3,@3/'+XX>H</TZBL-K/4??P> R>0K\"9
P'Q]FFDQZ<CI*C,P#=:J,A4VZ5):&P]=Z.2]3D]5N@5?;0(7MS177[JTO&P1:2NF=
PZDS%I)B<XFQ"UE"I;SZ^GAK=!WSM<2D=&"VZ6S#03.81T#.SS$RDP]E%12?Q\G\6
PU45YV>Y 1X2GPOT-IZD[)90FI;<=GJ6F$. "BX6[EX#U2TCTJ:*%@D+  52+[].*
P D(#Y$Z$W8'U=]F%@&>4)N"VT(48@Z[T\YA6X/.H8XE Z -:>VD:;]#;&7<1LI2.
P!O22"3>7];0]?1M,%2TAB:XVH$3:*X)( P CJ/-2Z"+ CD!1<X5<A\]!8K+JPTPO
PM06W9ZGC91!V$O]"696G?5=%V#O2 6EZ9G.IKFFO*O)<';4I25[*V&"7-BQ[NS!5
P]60\7F.>?].HTS+J1&QO,Z"&;NE.ED/76[]9?;#O>"BT=1#A7KNKH!\TA>#L&G$2
PRDOVP&QQA7:/FPQ-%AU->$L),/.(+]"" E'?$HBZ*B0J%]-V)O+0/DHJ'E@NPS]T
PN[=<L:HP-.S3^5*?GVJ(3(<2 L8D9&!U%AUB&?F[AZ;'0<4:3!F"YI8."ATPM3J;
P5H>]KJY'F3)$11O'\"YJ-F(TEJN--J**NHAYCW!7F^_U8,GNQ=R[UN.^"7AQ>ETO
P0\2(%1R\2^D@'>V;:Z=5=1K7W[BR07\E<R&.F9#US4[C^V82SREFQ&8[($N^!.Z7
P+BFW[ZNTP/IHGE@_I_I*+(%D2% 2V(#:3Y;]"%H! FR<I9GO<;N :)9^1.-N6E,6
PM!NRL[0 D(^_YPR"Q.*/#%?P-VT]KF8@)BF?Y\Q OL6@L+VD7,A$>:LV^4&](LW2
P!(A/4&&IJ2)0$<&X6*GW@2K!W=SL"S6<^UQ2Q2&+$]% SA5R=#4-B:.0K.7HM3X-
P=B;RM-%M=?DXS8V^N#>?(D\^E/461#T;;6@XRL@/0X1?%)&M"\Y#9CQ=A]3'$W*\
P:L0\O8K3(>(]83SH\A9ML(Z03680GB;!?9;:LVETXF;Q[75UH<9&&VENC8?X^@VS
PHJ6*"WMSIKF\57'=N!YH='WYH8D)WQ_UTFJ8<+A#P_W78TU];EV'F/=X(8]?RKHW
PY]6\V$?/95N<(QO,%Z/FI\D4T\LN'!=/CP5$")D\5X&R_6[#$87.!R>>_Q%,A-T7
PP6=IGVH3+<C6<>P%GQP=ESQG&56-##HG>%+;0.C#G+.]%5I$,RMW^U"!?U6J?7:2
PLK_+8YRLRZFGDJK=B5W0M$5O^X.]8!7;BX>>9$?2 5.@5O*Z-A*:&O'7PQB=Z61Q
PDF H&,?36_+%H')"*_;[NQEEE2#G=R\8J:;,<P<*1NKC<%XSPB.H(T$ B9/7X?EA
PJ,NQ;8G>N5$S,C@38PT6/G5J>O3W7@R=A3'GMF0L1&])<NZ0;?:6L><+;"-->[GH
POM9B/U6Z&",L!%T3NG;NY($M]#- >?^?!/!"62)"G\@YI/> =GAD-;*=4]+B^#UJ
P?DY[+VED1-AR5BRACJC0Q[[822$/G@?ZGY3U<U0O.0VWXYK+% **TO;QT*33D7H.
PW1HY1N!80DVBUIO] E8F-\2+P/G0-@QO.7.^4T-H87WG$O10?,&1 N941B"X<(L2
PLLL^^RFMM*DH$A>P@GW0R:O!"2RH$@P0PL4"0^_]M410#K077*>6IIG"+^)\)>OC
PRT*= 9<*J; 9I'HKP#,6BX%DMDMJ4 ^.'8O+P6Y3P'@O5<WI)\QAUP.H;E8^9LZ[
P$RP:F61>2<3>3DY==G(:5*3#&X&%L_2#9[I#;/]9B'7 _LWKIM7!Y#V "#2RV(>"
PN?J[GPN2^MW;8"1P')@@5)?ZX0^SO<@19DB#;),GC6^8?*$/'6XJ$@,@@LAZ#_><
P70XM]STPU96#YD[''-V[9>2%C/5CUKN"@$[PQKL!/GXABO.E7?7S#5U$Q><LZ.WB
PP+R1V7YOP+PU9NJ3Y5;T,*I-H1:1/CM;O/#G?+$]1'^!O.J#\H/:2O"^4>_DO!A<
P.00$FASD1,Z;PHY,O_BP"D]%[6+]AZ^(Y%=6%O+Z9$B BRR[AS9^SXE>Z/N=HZ0$
P ^1N>Z<,I@'WBR5.>YWKDL8@C0FA/1^B(:)8/7E.*$+Y_V<D8Q:ITC[/+Y.;H]!Z
P5Y9&+!/R2F;O8@"1C(_R..\7B%#VA#.0==-;](\)$&3%6U@2$]CN^6GEPX-)G\K.
P7'^!AV =S*/\ DA4=2 >4KQ%DPF%OM],FEZ8R@X62B"I)1U5;)D!EGAUG?,JJ%OB
PH=03F-YW<\%=5"O)C.]DQRFG7%+;2EZQ?WYM<)FIKG2@L#!,L:&^-\53"EQ@227O
P:4!L"6TE2;%CRCV=\)\X8DDA2GS@->9$<0[SB6_")#G;++,U16.F8)+B)C >S,S=
P_BGB3D1@N8'#MWQU\L-G*TP>X>P+7<-?M94N>-?,J!O4+/('D.(>9MX)Y#&"EE-$
P_#24R/YS)>M;8Q9@CM_>=^LDOBDTU31A$Q#^S+$WDX?/ITLSAO8'+$F_Y8S:G<8*
PNF3.EU _<)G'>LX8@HT:[.$US)-;'M&M!M).7-LA,54W]J/>(T/78@"HUG!T,B:O
PO1MC5XP8$PN/$-/<1AT2.'WV>M;BHA7E7$308ZKB:Z*BP-9C8SOF55"-&[+LX+[T
P4+O >+W@Y*/Q+M;./*J4YYQPF54SSZV!KTVP$!F_L7T$M'L5B1X&O>"YEE6]>)FO
PM#SI&>'0:!^"Q-WEM-7&=\AX$U>A@TL$%&3.%!K3;[ZOK;5YV8#)X_QM0#".*J*?
P+[1I@]]7QAQ9*HU[3#"0PTAJR-NZ&VC_,MD,1$)(C+4)=T;MK>=MU,"X^F^K5]S'
P3?^_EWZZ!T/M:A91?BFA<@XT.,!_F]0);9?&V:>3H8QG]"T^>6V''=]59!X,K*.@
PUU;\G'<B.Q_K>4=#I!Z3'L?PP>_4A4;W7$[S^K]8 7M([QREY6H=VTB(-\83?:L:
PA96<D&H3YO7S>B++T<7(-[+DPST.T)?6*462EWDA3%Q@C"UJ-1Q'2RSS'X^OHK__
P6_31[5__N:I3_UEU=*_!,SWT=Z)UA. HI?$"YA0PRZPC-254:8?4IE!!6<!CPORE
P@ DTRJN. UU:YXWG-IR[XD)DB2V8RV" /N6M=+:TGJ^R(_XKU%,'](]X96+8 HCK
P^:,5J&$C 9BR,3&)%OX"M%+JC,.+J@K-!<O;^U&N+D*:2'7"8[I$P6B93<D&-.%(
P"'M$? ?L"<;'#)7@[Q*.L %0.S$.S!#\B*;+.[1)VK1HQC58*+D^8 (M>#W#6A=2
PVK0R\^UOAZP VCE,CYQB)D.5%55=3T-2&W=%%\<H5%(CO1U-O\9QC_@H9O,=B.Z>
P[DL'K@Y5BHKY:7PY2SBN+RU&:H+]TYC_CY46B*<>N.,O74\*JF3J?Y,5L3G61-[8
PE'B-8JJ7HN)81D=K0@3*?>KR Q[KZ'NVNBQU+>@UE9M*=]L6\5("+T97IG%<TNNO
PGI;N'!ULD%,,YU-@&8#X"6L8;UGF@8"=>X =PGN"#Z[OWX#BQ"+WQ":X:>2D!A.Q
PE&3R70'OV+$4R=DDC"F##[,2>:?9IE3S+G%VO$K([O-;D4WMQG\[BDT2S8SI69(H
PWIWNX@*1V>0H"VC(ZP5Y[.E>+A)LJFJ;1@T6VM.7LX=\B4T.('+>6$C2(@&:3/EC
PYF:.I'#QD)^([W\A2"(<"3XYQUH\GT/%J+R[1/H5FK]X[.F'MC^^'H6(,07'AZ>0
P1RSD5;GAL@-Y;;(PP0-W09JU$*XC54&WB!ZN-$[@.*DD4D:I?:PK8^DV$:S_$%@L
PB1?-DGI0U!(?Q1'9.[!=BH*V[I!]8?K#5IFCV:'.X^;J ),9=2U!\[=.7>@^$8\9
PGI)=/8BM\>(M_P;:=TO!F*G*'I-7L;O9DS!$IX:*@LF91,U76=IIJ*/VL6QR]O\,
PX"SL;-SWWI9/#?^*XQ\:+A]=NX$[V $J2:\12,^7YUZ_M=V?.('<J.^RA/&!2V!W
PIB EX)]2<;'+KE2!(K8^W9Q;F<1DKP9(NW*=N)=O7D#*=YD;RIHZ%"V 8_A<W)6Q
P,@F7K><<>Y1<6BL X ,62S^<EW.$H9A;C\6\2Q;54+)@>$B%%^8]K'-UKU@8\@N:
PT 9PX"H%#,I$R[=;K&WY*!6TERW?1^[=38E/O4]8MR<XU0T$_P4JGD&2$P0VQWP!
PU9]%1LB<HX_[/E9-MMYKD7Y0*DR<V*&[1$ +F%?[=*Z^5:8A9.&Z:$#,-#X_<V"V
PT%IYJUE1!%HDT".?MAKH>+K2^ZV"-J2^1S:F>(/W!L[+J.G)S4/0?GQP@,(2H>F;
P!#+-^:\>B3AGGN\F;>N;#SQ/7X0[=AKB&T? #6G&S+/6(+$U_YM6S41&%Y&U)[B)
P$K*@QV40"MT4FV!#G.Y3( (QW8)/O=0:+N!EK 'VVZZTD@["[:2C]&8_R?52<7Q'
PFSR==T&3SY\]I(/9FAZC7$!+1BA@\0RT)+[LJ9D3O/?N,L\H/AV T(^\=,?T89ED
P"4J#604X&FKZ[5*CK]-@1DWS1/*SKL,&I-J)A4?^9PL!8M[>N+LM#73Y)[1E] !*
PJT'L'-1RG@-,2<VG\=Q0>$E6&1B>YNV$2T\H\9UU#]OJAQ IAI;E1MZ/%:HE\XV4
PD(4[]%,\#1@*68N#<:,$?GEHYB.SN:\VF0N74OB1Q!:?(=_I*JYJ^:7%+ ;X39%G
P#(9],59'O]0 B?O>4NR[A*#)M%%A5!V[R0"5E;]UYW0OU9JOBX=9WS<RH'MJ8 T[
P>UJJLAR*N^^ +[TLA93% G3>!A_GHZY($\4>,)3-Z$ XB]>M*;Z?AC/[X)3UM/?;
PEB1;T:/=$#1<B.S1Q1H#P4%U"K6VPD:Y?8M,)1PX 6[W*%#WPH?R)K_$.<@I_&#Y
PKV^QCW'CLP ?=:UYBD>?:4"?/&3PP%I]7,Q_#"H]?"VMPYMT,'N)W<KG3@[0TU&V
PV:^!9Z;O(1H&:[[O+#B:B>S#K40?H]Y_OG_!AE@^1K2LT7$F5ME0W+[<@A_P@^85
POTQ([*I(>EZMMJGKF#XX6%B^W[NQ%!>?XI#\3_HT3^F:^OZTE"[;^3$=SIB^A@X%
PLUK78E6"Z*BO(\72-O6!7I<"K%G +@+:]DP-I.H-N$FW9U?KSX%K#A<G=M";"A-0
PBMCA*BI(L(CGL("R-"]N4.D1,0N8*=LV21-'1J+98]X5*5I'&/Y,#L38[TLOL^L@
P/1GZ4Z&.87L1XZ"0-(:!%G,VET>:,%[<J1"UP?X0<6R:/44(?.BQ0+?XGK0W,-*^
PI1B2CN4+(O)VOV]/</U+RZ9^[DOOJ6:NG,P=\70HK"K.*85IPZ(QT+E))QQDW+X-
PC^I\!6#C0.-:,1,,/KVAZ'N^]O-Z;>O#5V'%+39J*+)+VW#Q[FN"!S[?MC5I3< :
PE*:Q%@5H03G[A,W>__SI!#XS?%F;Q".JI$[MD_F06F=>"WH?=N&B[H)O/&;Z=WO2
P$<!B.%V9+2 !.W#STMT$#1Z;YD5]&6QDF&P:%@I'ZEIKI\;+1(^9"_%WS=Z:_R9A
PR-,>$BBNUJT  !VL_5@4.+@0FZX6<[*H8*PQQ9.3#HUAEU);_U@Q(! 8^_]$'BA[
P9@T1'U!81T(/>@:WYX?!*3M[OK!V_[?IJ#,3LE8XHQ#0QMYA:!_B_>*F_SO%R&9T
P!00[$:1 V([I?IWH U9G]^F41GWW^1J@RU7O;O_B+@@:O_YA9(++)!1S!]_#<'\0
PD:9-<%Z-ZNG*^(-D8;D9I!4T13^=V_YM[K2?=J"AOEDB2:9:;-*.'8$!CRP &-%J
PV$ @TL_R,HI--ZA](,_6)U._+M9U1_:#*3?R9W NU92?SI"1B[;;*[Z6<PF<01QK
PK$48-IR;X"RVE=H4FR@/*P(ID(<G(#0&*3_]DZK]X(%K-BV@3U='K'WT/@2$,/>=
PVBH W_$/")):9,>2 EH:,?_UO91I;0.%3 7T7R#9C OMNG10';1F6PK/M;VT3L8:
P<I/"!=_9=,]U%[-7,7:0RU9+#B:,X/79LPLI]X>J7A<IS<>/)^>B69NAIU1C5'B&
P2OEY250^%L&BA[")E_>O#3P0A2]SS.U*MKV'SV_]@[X-QVCY-NR[O#,23=D?N^S/
P?^929S7A:/97PH)-@_;2Y$EK,I6\5IN!2<UP6W9U?N9C(X8+4P/F3%EXKVZ85?P/
P>'<$4V$MT.0HW9]3C,G+CQB:;,XD</R-HSC80+E\M<07@-<AB+M&$'SP%Z'9(=4K
P\2D9O4^S#&:?OJ$!'5)O95WXW6:A)?%4- .EK@B%7Q#Z[ (!C^+R-^GUZ)08"1;1
P\"!]*&T4C0OAV%\<.D/DI]\^-7;#H^;.-ADOXMJI+OY)5:5&54/5]ZR-$U,4I7\0
PZR'KW4T\:I&.8ATVM1:%$Q/Y(PA8IHI*)W0&*GK9<;:LWDXR>4)Z;(RT\%FKTV-6
P]VQ#VLI\-NC>.G.-W$$11GZ;HP]8=Q/LX"W$4@CKA5I/-*94Y,:[>P[HY@^D>?D(
PU6& PCJN5]-.&#Z,Z^F%J$F.')%=EM?G/(%>Z1S0G5 ]R0NQ,-E#X=1\0%V?/K[1
P[?E'U5=F67ZA<?L@RB4'_Y[&F,\Y7"@QS1[A00PSI29T9KD*9HP\E&F8UP*WC(82
P0?C<!'BO/PI:X?F(S\@3!GUKSN;<S%#(2<SH#]Z&)">9,8=W1M2ZUO/96'N*%SR]
P^>PJRV:P1@N@TFD.]F\@\8X'014/$4=EW:%S !30$Y\+O84P5'%TMAN@G?.R?7I;
P<[6Z(=E\MR,:0&:LGXM6.MHWYS53; ?CEM#U"V%;=K]1"6: =Z&]A-= Q@/DD2S0
P1=HK[M2;;TX5]QN2(9:O5#XJK?\95L%O]-A^(HE+JPC="569+6B@/C3I V./H)WE
PC?7WBT59_DM,[&[?2PZ!X+1ZB*K(7B$>H30++;36NMK5W^S38HTWW=V>)(876.SF
PH"%$@(SEL-:[Z+X4]:BI'0F[8A7*'YNMXQW)8? @#V809Z%(J:H?YE6C/F+,T$GM
P([#E7]MF9@*?STFR-J'M <[]P6^+P>YNSFAH[X'\T\!7-E#>[5;2[3Q_UHQ-X7K9
PB\31OF.I(2TV<L9>+#"29XF,IUR5D!0'7GR 6.*HF2(3@+:[2ES+8GFWVGQG[A&$
PKR42I&]"VV*!!9=S*"O#?@EA M!P<6X$230-RB('.@]NR!-<Z?TLIA-PM.Y8NL9M
PV9O69/0"3)6*#E1IF%/)(FU9^ *%""DZ,;/QTK?SQ:4=&CH]6ZS?2XC=NC%LWS_2
PH<OJ_';? :"Q+,$2-,$M]%5Z# -F4_#132RSH[>> YN4TO-]ZB8LR+27%.CJRK3^
P4T!'3O_HUM!0,,0W2XE'E3WY)=<2,(B4*KFPN&=9A'ONO.Z!3!=_"]1-9F?"FU^7
P]H3^VFF"-;#34,_L<]5^TKY_*#_I)_F$GAZ_1RWM2'REL!9?*H46/4.(E<.>NML9
P^J5I[AY-:Z ,NRAN+A*9MF;O'CN:00ZB]Z F IF0QPO<<9^L!.&!=2ZL;OVQ[;#;
PE#%7IG#0(@RHT-I(T6G=]+G[*1T2ZC=$D%.5=;J:>+*CJPO25%[5.X-B^PR;L-H_
PHJ*ICSFH?L2:=-P(K:\IRQEJ("\ I>@Z@;GVV/D.SLVJW54H<DH]5':Y0/9V@]:A
P R^?V\6W+5'%<9>6:JT$3 6_4%'V(T\4+H_9MH8"5B5C9$(P M?[HPF 93!@1T<J
P"D-Z_3]:0&3Q!W"HQS'XC/EY,._JM7W+5W#+\;8GXN^7 0?-J4-XB#2;/HHX$$F6
P"3HY8B@GR;X= -#%/MI\NL=I)9J<9LSN0=W&C(\W[6%;JA.:-)<H]"+"F#W[XXA_
PF&W69*<I^A UH:4:RF50K&53:9@G )NCL23/R,+( AX"J2;NT-\#%=T=2C:,)L1.
PD>T(FA*PUNOEL/A"QT ?QMD+S%T4%JD9,\A,(EX1GY$A[+,+T %-V7Z+])38P;XA
P$6[H/9NU3.BQ-X@14<:9LE1MMGD-*]>X>Z7]2PF8Q'TNCM,ONOQZB+XUSSZG53R]
P?%=-?!1H@$Z)PQ3E*WT1_9H!!D>V&#<):;%>;\_"1?N*,&NKD>@)W;)8K#?2%@T&
PNI?]'OB%?H UYIC/;<$-,DDOT+U6J!.5:TRV<$ZM"S5E7[:#JF>C6+&9RXOQ_7J#
PG23Z!$Q0=Y6"^?3&=13=0L1]>\##O)>,LJ2!D$LCZ*DXEE*EL^-?58XDJ-+N/EJ=
PJ*8MH&7\GYY%$%RZ/&U]UO73=X1T0MJ<D#4+!E7.IQ4 J.[GN5X8[)M3_&^,N7-6
P>?WK:1^XS^);L(#Z"2@ZR;YE&LM+O6CLMZ3N8(5%0$/6.F_=O]]VZL*N)>K:7Y56
P#XQ@::@92P&Z* ]<?7+S"LN)Z^?O-$>%88!\4GG_EX =SR9$-2$VQTJ#@_;)W/&Y
PR+ (U@Z_<ZB45A'9[U>$IZU@"UV$,'C-D,ILW;4Z$.[[6Y1NYFM2)T;Z*CHIZ%@E
PO4>(=S!*:4 @\WEU= &FQ2<)?N2A7SXPKES8#RP-$CGG+]*>&*EM/%AH@Y)(#-;J
PV3%.AX+W1 ;K]_% 4K6<#SC::68]P.2A\75D%IA4=H^).E-U1$]=&1@/>?];',CP
P-$P1^\6X>9,!ED(N!;@OM,45MQ-+=WVXNN(Q(8Z00>:>?@E!5 K!E_>L#=[+QZ1,
P5AIUXQQX7UZJY6GA1[O4T3=)<Z8!_U0< ^&%&& _7,<&XAZ-O(W[];SZHM07J"O'
PQ/PN>ES'GES+NC1,%.Z!W)J68%CN-LOMYX=@5O$,VSJR5N@LE3SU]V%T'\H^X3I8
P_;W""=&5F/1)86MQ#4\W!7,M1\;(_MWN?[WCS*:8/RYJN&J]%88Q1DN+%\).P>T_
P4/8C,C8M2P %S:81'6%8N9+0;BKDO(SJSG2-'>-E)9"OM_)81@H"TW(( 9[F.$=<
P,!='VPU[=(5&&Y]Y37VZ<B$K)J8D"2.S02\?#C?B=V-75HM/*-L<M,G/5T/1NW5&
P][OLL=POLB>&*2> #AFR3A>!*3%+4+9L/\.C^$%KN*BDY:F2V1TL9S>S<&Y[L8R)
P'<N],1D3NC+ITE^>E%AU"OZK5!QS8-T-V"Q*"KB*QC[[^]*9C77K^XI!<---(SGE
P_7C5 CX<;J"QG8AZ(.D!+ED4,PE=I9BD;]ZRQ8%0=")N?0YX:;IDO,QH+9P$ A5)
P/BQ-$((Z"0U$2:3S=0TD&EURQWLN_>N%'J17!\,3E.ZE',9Y9 0&9Z?]@M^/!A4X
P%FBV$H$K.98I,ACO!>C>>5\"P2 2T$>GZ=G?V0K;K&;/01?Q_J8.[WWW%L:[:*)[
P7(CC*=D8=5238+XKQ9+DS\,ZMH'*9,!7@"70_8#,S76;K,0XF M"X!?6L,GU:^<"
PR.\SO!:15T7Y15\D5>XCCE)F_0,E/T4 K)LWK%<()-K'/34%8)EILWLE9W3G.^M:
P/,^Z%=[A_-#+X\.X(VKN?ZV1,!H)OC5QM??A"^EWY3"\@(^6]5$:U"F1EL*[TE9<
P)^9AD8YX>4IS9EF-H3FAZ$V&"(O4KE&F9%!#W(- _!0)1'*5],;>W$ ^D6 YO(9 
P/ZN@UF+);90^)=)P*<K]G47WQ0+$O?[!^XL%-=CH!? AGP27?=+S8*U>4 YKO:T(
PK248P]V6Z8N3LMRR)JICPW93^TXL&6/(^CT7F7X;/45IV3SQ0)K0)(%(81^9 ?XT
PHUP=V-[+Z S3?19:L!!&S" 80-;,#R7FP,/UFRYM'8& 91_<V[S@D5O9X+UD7!&\
PKP=A=L:GQ^+2;Y7_9G#ZN EQ#1-)Z.$6P0BVU"BV<<@2(4?/CM/_O5D:&;^6<MF@
P:"Z@/P!IC]%#VD-#UP9CR^.<4>H,%(46/5B9/OM.%7VP2A+FT $PFLR(J,&R?@T&
P[;M&^X[> #0\+\GIDH"KA9#MOA 71L.9,9R=/MNA7R#5=!:OIN3Q/#W+?0TL^:Q:
PDNC%DV%I8;Q?')Z'4C43Q@V\QBY9CRJ*@S 'UU!>4EM#Q=O?V -Z^<M5SC+)-X&0
PM6HX>HB8MWIIESUP/UUV T6IZ@1775ISJ%@+GO]&5B\&]!(T'5>L[#XVDI*J=07Y
PQ1D@0X)B$MU9L6YF;'"+T!Q7Q68O\1576F;SI "3W05TQHA!ARB#1V,FO!TW](YV
PZT=N]N[*[!J<#]SO03UQ[5U&)3W(T/Z3(/:M+0+HK5:.?(SL U79A6E#WW<#J!@ 
PI=T2GX% 6)[?<=4ESR WAT8.CM2ZA-V K&6#1PWAK3#SA*<D)0I,MN0WVR&VQ&OG
PVU@/1:WGY7>A$-=@/^Z3S&D,!/,*RR45)D>TU$![E<@2Z/9M=U,=V&BL+GJ9.Y64
PSMC:M@0C2K5<??YH4!L+I3SR!3]3&F;"\Q0@/;9!G2\E]'@$L3X*^$W/=C&\$(M?
P1G/ZNQY4ZJZXN9H:EZ8OL*R.W0SD&!3H<"HGVHOT=N64:6 E$,(5SAXW.C[:[2>O
P+CO$)VZH)7#V)K0=INCL/K=,Y=#[A,).2F$)B9!'](SR=,>_'GM*^Z+#K>%F9WHU
PYKV\>1L[7?'7$-#1IH*MI?YD94L(&BOA($PP(VC+8[NQ@;9B( +U]&&5F_6B)Q7W
P:5N_(^265U9EEO:.J512[/WQT[V0J26LH\6[W"<LP&9VD7+W?Q')6 R&<V85?8&"
PPR6])W;I0]6%7*N,]I$MA%TZ*CYL80>J7%I$)M07_.2<[(E)[1RYY9=D$=[[:7 E
PI5F*R,.:Z/:C2JB-@'AI::7<#B%'5R0RCV0.0G__XW1"2C<LWG#OAD-=58LL[31L
PX2P@N)C6^;^$;#6HU'Z5X6S:W2O7V*Q ,\Z)$T#RI\'=^(6,#,&I@)"V*)(?.NL1
P*PFB!L1YHL9^91]/U*905FX:#K@J_(+D2&K?AXIZB2M%Y6AN7%_8YA2LA!@/H&PH
PE>_@YBIEU!_+GC,L7D3VL^5LE\N44\H)V30&V :_Y'N9S_%K;CBA19.A"[S &>PI
PTZR&AH_MD;Z]= N6#][G8R,)@=BZX*$1( BI^D+E6KE"/?&6T0])%4_HC<%$2$0G
P!OX.9_889!^>$(2\(O"G3IA+<ZIE'NGUD&F\<B9NL\8U]C<Z1LNZ&ZEJB%@]^^-+
P_FC! -$K"W3K)]Z(%NH?3U=?( ]DP$1E*+()9J^U$Y&^]=%"VC@^P'D/^:)6GY:K
P1>J3PZF..GB 8-7Z(N1?&\^6O#NK*S;TP30)9 &<NZ A1[^P?+_7Q'P-P^%]!G7O
P+HTD4)^Y*[.LF]TYR^0Z2\DL1%93A+O#)I)/";..=FL/A.F;O_66I"%+Q IAEK^W
P&8+1Y(*^K"N>5FB:GMR'PVBPA[::)0C'(?I'G5NDI3^I-7,'A^38G@\$V_)+?Z:I
P?/CI,>M$"?T*P&TQW<?IT*]F(A1^3DZ6]_1M1)/G'8.[4./D*UN221*P$;QA<K-X
POKPGUA5X)+ [UJBVO?]B9ZN5]5X3S9C*,')1[!3%&SV8W\@[1!J03^Q&?+-AXU-"
PN%"9VE;PCP@FCU$3=9WXTAL(W/(F'1ZAI\P#[88',:"")BTW]3GJ)>SO:DE4T<HM
PYPO:8]Z)*4ORQ[EX#JDL<^MTCF#$9<.5%MJH>YN4_.-!KJ6GPCYW2QS3#3,-4E#J
P++YAGFB#*[C85YQ=&?5VC<]HKBJ"BVI':B]'33L#Z]0ALB.Z4CMB<%Q3*+&+80A9
P9[(DQ,1P2M*9)B95$WNE(F8"<O6I_CEE&!X;3H,I60MO"OT_D/6_DE*&#7LJ [1[
PF=$38N@A%/JX:(T/SOA"8YE6"PEM9AOZMD!-*V>J7=;(DG0\(!^7H)>>B';K/;1Q
PT9G.O@K604=V8-'L'XU(SDKY#,UEGJ0 8Y+\N6DJSJ!&F98MPEJ2*(>VS*U\R@+I
P-_X6^SP5]J2ML2G_&2LH4K$A>_2"?)[7O"5/Z"%NZ1"6U=>H!?NIF.A)LU:8#\V9
PD,T "6*0WU/CKQI_2+\<T?I&D-,K;A[%+-IW*5I!5Y*#NL%2.5R86#576NX$'E%P
P^!)2['+BU^C[;DAH[_[^2C;#!G\33&K^ _C=+#1W#?_TXD7C-?W>*QR2L5Y\T@["
P%QJ[H78'WR:(Z^=*(O0[%LMH"H4:G@C\>I(E3U#I-W"B'-2,MFC"("E':KWU#2C&
PB)%>*2L-[PX82+GJ6"\HWSZP/'LUS0"#N[J%[/NH[A^HQ"].QW6??XT/ZAUPIZ/?
P,\H&C_5B2(71($/2]O.JSYZY9- :SIVD8>%@F/5AU-"VA7\\XCDCF4K>&::9M@RD
P4,;(WK8L%_&^E;R0J%RFB-1G+/Q"YU.+ RYE\T4Q<&Q.:XZYT/)[O!O'&)[4E.NE
P-L?7&3HU\SKQS>W6]U_=R_W)0'>;+,*18/QY?=87 $TZ8\]PYWF<R!9CST5/@YR,
PDS*X=.G1Y?Y=KU+/]/;P[?<"-+ Y97R2HGC**KW=2IUXB*0Z9(J_&BK^B;Z;4++:
PWZCQ; KY-B RX*/' &7>_<:Z[S*LV?A=:4!^*(3L;Q2)X&W9VYV[2'/R$&D8HD55
P4;2I5=&+&0C'9VJ 8J#3T%B[XA]A);J]8.]CL=4)'R,F"GA,@RN:7D]XE5)-"SE=
P,20O1CVI<(4* $:H[,:P6D$J\4"D1/) 7%:G\4RE>L<#W\>E7S-HQ_R_#:A\T"+?
P1HY4QZWTEP9/G/@Z;?B&Z%QI7%;/V#P_9/=;U,@(G2:J]F<_Y*$7_2'B+:WBR)>&
P4LF;-?J$VY(NQ.-&0-OR;*BQ#Y=-^J(_1A-RV^NY5D)(X<2/2@AL:>&+<N?^R$TA
PLQ](U*;*PO)GI5BTKUZ,:,UKLLZ^.VDLHXZ(/8IIO^AO681$WE1<=X-9Y.<V:N*_
P' >VUU%*,H4=@;%<1*?G(@A4R0W$4YS&7"V%@V,Y=[;X7-LJ=4LP/>; 'DGY8^Y/
P8K3Y3:U+F),EZ;$6'*$" CL:YR'E>4:XE42Q,HYG34Q?1("4(C3;82G*24)ID$9+
P5/%;'LIOF=0N$9*BZW0Z]413H5KU#<K>UYL6#;EBA*:ZS+(S&UISO_%>$=85JWC&
P4'5&/Q,8Y/MJ!\H%G F771O@^U@"U2+9H8J>]:*.UM!G$HB'SF"Q4[1VFISG;KM*
P"Z"/%:4U>:'TXG[@<<@::4!_DA4'+S(C=7DJZ)W7J5V34KQ8GP<Z4^%499_SJ<:)
PCT52&J'U!3.6"OL]\[M-DGT/U[8C1E4PR37/.SRS]&GTH4&]9?NL\@ZNE[)8\DUG
PH$_1W3B]$\$7G0L^FL22 #Q+N1=YG:!V1NP&:<2ITEN]-;"@Z5_48K]-\4-5RUXD
PW?^ [CE3C,)NNV0PP3\<$J10V2#E%B),#@(M!('H#4'C.X>@K-Q;S5NN8X]&^.Q$
P!;SYU*3Z?B-C<JO+)=H5]TX<<:I%I*P;91$;8>KPRG>/":AK61:L)8K(:*JK&][]
P'H7:C8D(QQF5[W_%7[9QG^VT[N5KV5:)W"%YP6ION5(_4 \?K:HCWIUBI0TYM&<W
PD]2"VC>0T88"<G=6?L?P$>QS$=0L,_0Z3B^PIM:PTJ98# QPQ6?%F=NIW1DC;1L&
P/DF%:]6\I-.]U'P #W;VMD[.I.1<B3BQ"$?R]K&0+'ZWA2XQB$!YWM 84&WMY'[ 
PTY'!T$W6)@A  AF,^<Q=6R=I(-/*<V<QS&PCA0../!C+5;IK^-<U;H1J+Z0;NR R
PR ;M6(^^7P>]6(<9OQL@/<*Q_=A#S>LG=D^"8':*][O#',XGY,7U'M(L3<#74G0F
P"3K:FV(*DDLYQ&U+U;,D"*KL!@L[TPN;!:*1!%H,AEJ8G]FYJ3Q.Q.5JF@Y/M\LJ
PAV.YE;_E*I >/TL9(<]T6JHT2II^+=&D,.%*E*X%8J3VL.42$L'\ \4@A6>TNQ9M
PLO?=B0 K/_?*O^ @CPN^AA[*>^"%:X1<,1O]7B15ULX'RZ;P/*AZM;\0Q%%/NY#N
P:)[\VU7723<#23Q9PSC>AR<?E)#= \H@=%MM_Q,8%,RE5G*=[)2Q[5<JCT0\@=(_
PO-^59M0ZCI\7:RJ4/R$)NP[=$X\H)+UQE;EJ9NSG T@ =0-^H'6($SUA[ID3BH30
P ]1YY2HV2Z( [CL5T-.!#$5'Q]C9!G._<^8PLUG/#W1R,=G!%4D18X7OI]-E7=1O
PP?3R!+ES\A_/,GO0>B]G2H*93"\,^23S<6*7APM+NL6HV$^\%Z[- 5Q%(B?[CDQ=
P1Y0;BPF!E,'A>$XG:6PUSUF#)]'9I;BG-'\%MR10(3J5D4BNIX>#CE7DFZIH-<JK
P-G4UJN8+MV]6TINFY\&V5[J:BUG]5-#E&F[;&E"_W9.3<KBI3)X4695\P5.!IC41
PZENF--4+DX76^0EO;E6*22)OQ$SH_S^9LQ<=(&(>2A>_];&!R;,I9RD,H_+OAY\D
PY/NERC$\3;-TAP+9<(U,/!GM";<[VN[.%%W(>90Y28F=1>;DRG::;"</3\UD-LK=
PML)CJC8; J_,E -U&G 5QOYR/?@4DL_GM$(7*:S@4U(N H.TY$S86*.P76#!?S<6
P,@F4[CHE#X&E-+NAJPRW2NCW#=KOF[,0G-G=IR0LM=C\B-@;(>'G8X#'W_F H&\_
P!F*C@09V3N/-K.\(D6..F;3@PG^'AGL^HYU-&BBOR(@Q;-\?)*\)K"]>#RN]6R"[
P3K V .9;K!/@_1:O;_V+Y;] T93^@"_K^S5@1;N,:ICQ2^16P "]!ZZ11.7&;J^C
PLLEK7CC$H?ML=^FU6WYWT8BK?C;P?1P=H1>M=H[)F6]_(8QHC!^* )68X2_SD>M>
P+4]&!J>)/82"I209)--U,H,QA^I:Z7ZNN.UU@JC&\??60#W0VOA?Q"-&+]W%SIIU
P%=0.I<2?9GWJ)&33>MOK%\R +&A;]RE13$.;=?)RS"=)[^L+)<I\E_ ;^K#$<*(Z
P2].*HS8N?25>I1M5*9COCP@?M=-.REJK#368(_JV[YQ(#CK,]19(1H6E8PEV7N G
PTP2,^)TY].B&5Y](SH"B)&^[M5M[ 8POJ[YDZ>=L  P'>G)2?/7*GI_I/(F=W=K>
PV"-O5-!)',L;T9DF@W/E=)/&%5>'[6PFON5DH>J7XVBU-[]YT!N>*>EUP'ONQ!R(
P(@RM$&CYD+0^'LPM(*XE%=%P>@$)&(++DY"?9YZ,=F87,I+D>;U;/UJ.*WU&\@\J
PN6HRT-'HVQLW%AK?=S J[H$IW" R<:N'9>33[R78:7]@)A0H'=B$-B"98SW4O(4*
P;K0BKW]//_17,VVU4!-A-!'/V%B+A"3T2CDK/VY8@2 $\G)58^(RN[J=HHOU2Q.>
P.TL[.STBXA.=_C(H/Z#T(IJ1O5IE-B _YUE$7E.SZ2M;7#29!2,U\HM2)2"LF]/$
P]2CPN=;K^RRUAS$;T+2/_+V9WP&!0CC2//\D;P4ERCCV5?2C6D+V/6N1=YG(1SL=
P^SJ$HOV#\:HIZ=W\U@XAYO\$NY3[Z+I09TQ(@;J^22,/=@K7P=Q#:#ZR=.%FQ-'3
PTG=U#1A0Y)OMJ/R-N4I>JL3J7M<21/E*U?WLH(U;10 1C]M>DRTO1*VH]\O_'--Z
P)B'Z"=NSQW@/XQBI4TQT+*: 65O[60>BJDDRTC=IZC G7GY_)-G\\9M ?K-#HGB*
P'B5L#-R7.0^HGJ\66+%EAFT+EH,.'CT]YTX'%#[MQ;/@]GW[)2-L/<6&@0$.ZKP+
PO0^!B"C#?I-+SW'+ZNY#8J=$"]2K>^,Z0&Q_:@4>2E$#=C2C)4SO@Q!\L46I1A8A
PPVZ+[R.@J&N5XX?4^+M&NT>NAP4GHG@2+8SHBS+Q:G;.1GJ< M"S4YIP]T E%-T6
P.43X.BA=GHR]CO\DQ[:XWMN:=A538)<SPM%.$Z<?2AK()*.H+#4+\1K+Q 4Q-7$D
P .GO&=X=(#YH23<CK>>LOL9VJG*8!&Y^@AZ"&LB:WRO"*2RT;MOJ6^*#+"G#.@QI
P9[K5W@*/G#[B.P1Z1+<&3\G*J:+12\/G,-[Q-F!7.A:HS-R#W/K65GKJ_&-(\"5@
P)[UQ_T_.XR]L<=LZXP3[?@>H&!L:%SML]XB5]H=@$LU5**?>;';Y@U$9<\'O/-1-
PR TM#<D-!ZO1#7(I/$)=93/9(T4ZX%F>PBGV.0Z(QT.(UHT3AH ASJ_9\@L+91KS
PK>YT/WXZ=MVH+J""$C@$-3]K%:+I@(W1<\DTL?,,N3G'+3YO'A*4R$ZNB=VWU,3Y
P>!F&1A'_;\ 8ELWJ0]I,NN:V8JHA ]%,*SBIJ"U^!K3T)=E,]:SR=<KT_3A6':M?
P^M=WN.=U)EVG!;@HC'%F5E.%]TO"@M[C*H?!GY)CNG%  LGT&?1- N\0'!U0\>9-
P)>?Y+S<L.,H!9J0J\V"+;HB3T+S%7054G].3YF]<S5F-,YOLJV7]::V4SLYJ1KH;
PS^O#*$4AQ:@5#1%:&<K4R;1>)-2W5C;1':\DRVIUAY%=+[)[##3NBK=7,C8!MYMA
P;F&W":/^(<'":LLD=<K)?1I[&;^P+_V]G[^9X4=Y/HT%P*!0X@YQ^85CE:LC3AJN
P.915@=BP(<8</#YSP S5_PM24QJ>!37QV'PS:A'^4\M]_DDKTW!240J_DQ2ZIM/I
P33^<B;#V/I4H.*K]? 0.R*YYOZ\<E<-KY72(Q+4+K<O<13LA^7=EJQ=85'9?>RU_
P)TNJ"Z\+Q6X'8:FQL<477WF.AAG1'04H!Q"WZ_?ZGN'L*,$:H'=  M&'X DOQ^5\
P[X-W+_)"M@4/&AJ\7AWA<DL0\D8 N]K14U=#?:<T%:LN(V_(XAELSV2:*X?N;71U
P9&A%=^9GXOA041)00:XLXX)\?;P#?:)FG4E:@:/-]/TN2J1E\-%E[_AJOJP04#7=
PAXZ[A;FK16B#>3=_<^]T&UERK'SR[_&8+$+IB"YX?L:C;K]]$1<"%&"(A9<MG$ZT
PBMTW%W95:*PUHR-'B-46&REQL6Q<0^\0;=EG-D,_?"7R+7Q0UCA)D$!_O3T3LHX2
PU9_"/+69D/I+6RUN??>_3_)P_88F%='E'9*GG$KSJ7!"^UGGNO?.RLA6Z4Z=S(;"
PH\J^H- PT K_J-0?Z5\@6AWS:Z"T-DPJ/Y68;1%@W-G@M[XLZ&,8K*4=F-A]N2>A
P7J);X2 !_G1C9BM2VF@K'=[H'3L@7IZS%"5UL9]13+ESFZL0Y:#HO@?(H.>G<A0@
P/FG<"6$Q5I UF,V+>^#+[%*J^ ]:R=#1X'?[\T<#RMYEIIFW&_S;+<>WQG 3?T0"
PTE8:*O$11I/Z8M&RKH2LM_KMQ&>8\BOB 4J5[3&4_IU<<V!$0>.V.^!2'"2-)%Y$
P"5:D#2W\FC=X2B,4:6#NWK 1AZUE];T\*:%X-TIK*R-)O ,:J!ZNZL;\D,@'OSGP
PYV+(13P!\A*,JG3ZW %A9U?H,L"E-GF,@3JBKCE@9?R.H3'CTT2U#$_3D,B_^J'$
P+"[(+H":/4=9[Q1TP^-*$X#& 8<C%49+K#AZ!ZN2273[\^;>E19^[GO]<)3ET!VA
P\4(=*3 ,<.^G&:>9>E/KFA.(TR(WT$!<(6:S$6?Y*7A]E9"'@95TN2YJPGX'1#,J
P2-3-<'*&FT36E)DTU0!3I#S*D(2"AG-)J,'\#L)GED<EY(]V/T&NJ>]WM&K!?=68
PM,_TLK(=KXM)&/5,0@VMB=?&E#7P4J\5^V1>XYN.TQ[ <GGIT9I LV)CP+GE1/ F
PFOE=(5/.^/&>X^OSQP7(RX"Q$%FP[VT(5][0"PRX$Q^*V)7*)+@&0?*M#M=>%LR1
P#P%%D(_$K5?>XM+"14,(^LG!?ZC=Y3&VIRIO(-.;FG/-X,PUBWOUXX8.E !Q8+X>
P A#ZW3,G$&;I)4BM;AO P<HPE=6A#0] -5]:Q!5 =(N-;EC$1XM6O45#T?Y-#>:.
PQ]R&Q2'IT.7!:2^C'07_B+U"&<&&O3V&754=<&.#4;P/[GV&?9-AC?:D<#:E$XG/
P6 R?-2CZ1%D -\DB.A!TCY-7EI R?>Q5_4Q&3VEL"H45LF$!#+.EWFCHHYU=Y]%7
P5*T0Z:+;"=(!^P4MROLNJ('-RZ8^-MA/6:C;VK7\5RW46I2<1-]NWRASYN.AWMP4
P)_4%/I":=A33V-]UKLTJ:H'P#0>%I@Z1TS\T9Y>;.(+C-&7V1S,]RBV(-!2D),#+
PPP\"JB11GQ;]"#>>[0]VHNR8W53P:KX-/^2>ZE$C7';I!KMT97;ZETO10V3D+D.\
P!FFP(6U?5]-B?6_('3I.JMC6I6&(1,Z\MJQY>\;SBH5$9GL[_+9X &" C&QKT[!1
PG[P>59L6M]0;5@K)S:G*9UL.0Q'E"-M9ZVM&W;#T'[6%,O-'>'I4*8-T#3H\)TE,
P3;V\O,5U=^5.\VIP.^,7,5X'.=,O_!!3UVI@>LP0OC4E6W6Z44B%^#BYUY,Y0DPU
PYFLOH/.!E9'][%5HQ>:Y7"FK&,J06F+USZ+7AD:YOOY*'H$/-,P&X>QMVG<3U-]3
PJ' *<M"^9YG^VX?E(A3I-I@8\KN'336 VB9)QXU&A;]^(H(>&F]TB'%V0B;A[P)D
P&BX(W:+24T_O\2WF+-: KTW4P+*,0 V#)IN_]N2F %Y"B8>A)1EU1IE951KF%=R3
P%DY2G$IMOQVOO010_^[]3&Y?@X7*-UA3[]4R,S1 K_>.5["3[IR3A'#FT=\,8*3!
P!IR(A%AF_G'N%+,9KS?R_11_Q#=-NJ<)53"#\0R_LSCHZL/]AE8C4OZ5&7\&&"'A
P\BJ2G'_4G?<-U@1N$Q)GDW8W7X=_:.0)O/YG!R<# )<I9P&7/.:4TLB]UV)HO(H>
PORYUM%ZR!M$X=.@L+4<<RL[S!9?PN2Q;I5DNCJ$6:*7W6:BK\I\'4LW,AG=7]S$E
P)5[5R%0GVBN&=X)V$V)67Y(%4!NH'X44)+B6RPRW[K&#A;.A- M2_+V:KWM*_AU*
P#[T*B6"9H)PJ:$A]8-IY<T_I$CPD_E-192:OKO.4FB9GJO)MDP\#RYIYB!3QZ#C<
PY\Z1J=&,Q-'ZYXP<1MZ7T'B!A!UIQY1MP3#9'X89XA:*7S$[/0F]8L%B2@E^YGZ$
P/ZR?(?_IM="^&,3*3O?G$(6L#1P*E"Z3U!\VC7TB8P\ G9G0,5BIU1U4=A6_7*L0
P&KZ$Z1D$P6Z@(;Z2LO12Q+5[:^(.>I<F")ZO1X+G6&RM%VY4N=/Q$[E@:]^8E7#F
P%,URLP/K?'MU,]_ I_,.W&][B(G-8'B!-<_&N>I:9EDJ0@^6S?9\I14JX1&O#]B:
P2_+>KLBZU8Q,H7W^^U7;4Q# 'AQ'!8;.J7\7-3&*SL(-Y"X2P!.:\>)2W<Y>?L$2
P!3Q+\@%1*'0Y6&^O*ZT;A$R=G'TU(<2APM$JD=<U'@0+X)K,;(F%V@!?M90P7Q+(
P D>!4*=.L[.M<M_;O3;('M\CANOM@3=ACJ^#)]:_7J^%BPN <[V5QVTS><92Z*+/
P77BSTTF'M/,68U[:V>A=UC.+!!T_9DH'6[UL^!'HPA557UY>)21VGR6JY@F4S747
PCWQQ<O8RNQ-&@!/03A6AE*AS8#EU5[W&RQ\ :M%)9)IFKY9R$\D<*00'(W!G))RQ
PIS5CW)')49_!$/?RLOWK'#DK2\C-[^'C(7EA<7#_&P58UR96H!;T]>A%PE99]*>#
PU5_N8F%MLX?9.1HWW\40ZH9:T6AH$"PI$$I.?T20?T,\_:+\39WE/\CG=A(0'TDK
P$?.;TDR*0Q"TOSMOBROLYM/P^Q@6>F.7X,WUWE#/7@ [--^WAO_@!?!SPN6LE\!F
P;30A\N;7S)MI>?7!.)9&PE F-EHSQ]U@,RB6#>._(JCP(B?4..,%KYF8RY[B*:%7
P-\]@'.#?AK7%*#$UH):2_B)J3*/+"O6WL$;KOL7AU;;F*VU Y-,E2VL\.)'>-(;H
P(M[F;U,8M,<*)&PN)%L/\>Q04<C&88[A5+FE4GN^H(6<0;K'%(F>+F,U6O08<.:G
P/"&K;B*MN" :D<=_E;N<EE8HYK#;=_<7>U,W+LTG[N$9)%*Z;:-:W__@ND^X>=X9
P[T:M:J0+7P_0192+$C13B7V2-U<0,=\G)Z0,_RX2P$@3RS/'*F # I$$.I9BO8:/
P@$Q7?70K3)Y3\U-_KOP\S-SLR#-\$G4OKBD0W)SB4R -8U/_VJCAQ>E!\TW1NR(,
PL(-L[Q *IY=B=^XY:NT*;#K'(X)XZW*$L"1M>N-H1&::'NVUR,Z%Z/CCY X8R3-J
PUWDP>ZL5V0-Z$/$L.YP!)K[BR-:VC."V 1TS[\BYBT4CZ5RKBT[AL9=9;WO1 1S5
P!<VI?R>>=OF?%5RW->M"D^V"4L[K**;5ZT6D#%4[[W.#<JJG;[+FN?PX0=FS J<"
PYTY:J#9=>YV)HB!HTX=A3;49#G.H*H2%2]QN%Y?DT@A?:WSNB6G')NB! ,_9JJE.
P0)U*EJ4]K6I*RKDR/"XB%,RAO/ZPR(N"-PR/-3H:[ J.]FDT37" XK8[F0'Q+D!?
PF/+XBY>M.8Y,Y>EI[-TJ"&:YV30KQ&^S+RK]BDFYY4UAW<^JJE%,4P,;*@DH:(&T
P 6B5U=QA3U25\ V>YVX>>ZK%^V@7YU R-:=#?_A>MK%;!T=R#_"9#C=^((7%5:9S
PBFESX+Q!M5B$4K5+RB,SP3-Q$20(/[LN/K=N,[O'"98HI'<@B[!P_K :N-"O!%C?
P>,LW:%UC(,/@:C/'$ J3A^;T!5<<ZA)[.3&;V4G86[K4:$F=):7H 4IJ\6-,LU:(
P?!;O<4.D?<CXEM"=_'Z [M4" D.D?F1)W4\+?[JO>@I*>LC5O?!,\R3>?OKE06.%
P9=&U%9K+*8,V$,F-%^F^Z$-<JNUZZ(IWO!"1,R*>721+V:2H)3\2)9/5WX'N0IGV
P=A^'-RXP-C"CO_ZUM:"BT0;5IPM2C'+]_4<6'[8V^_+.Z4I8W%'D"S;AU,=>P8=7
P>2>HV+O%<^ _TIMV[&:4_>"Z]DRDDN8J4J)HQ]=CG*PJC]K8+P34]HBHD@:,C'CW
P)9?RT++:7E;7."O;=,>(F;$PR]0-7CX$#W4I]#K74LIBKQ64JJ;FL-C!9W+02C_@
PQT<!EG*G1ZL_4HY<MR^M41\MSG.?=$C-HCQ6?U)ZF4&_6ZQDI3!KU*0ZYJ57DN0F
P^1*:8ME<&=C%A<IDW<EQ0T/<OZX'&%R"(B6.4'MF20[JY/GWO10CX$<W5.@B:J&'
PU+F*9*IJK WZ5EP#<L6 2SKAI49&#@!>:"M?R7WA[-NDL3*_>3:!&#;+:U&"'.1!
PX1F43$*C1<#Y-Y;*P51W5;WNQ,V_"*_,??OY9J^#[-*'E>>F9+?^U6(T*E*K$4WN
PRSIJ(E-1L/.\SUA_O',APA\"9 /Q<1RMB;M<'9KT_=3DE:#B& L/V*HAQR]1<N14
P<HX5*P@/UB_]U3G)RP,Y%J(Q;41BFAP^>7=6*B[Q%55=^8;AMU-WE$^JE2."WUVI
PJK;-6>APCW3*JKV.'1!G9[\MG(YKF7@INLGQ^ZA48E_?.1]Q.O?QF4<,/\%04N/6
P<0M@,VMN@M^);T,68Q*K,DY:#QO=8EA?)WG5GO#GTA7^&@YT(=AH#02]S:>'&4Q-
P#&9I!FP9,W)7Z\SE$JY',7&QZ_T9\I+VF6 0SABUZ*6"L_.?QP%6G/S?Z$ ^=8*O
PBP:)SEAV;&_LG)V;[V??'0+3$%K:>(IZ8M#/7S4H! <T48:PS9@7;6XKH5^-[$CB
P5_]6B>%\DZ>>%BZ@%D0^;S$')"RJ0IS4YZ]?]SA-^9Y5NT-5LG;WB2$9;$N; #>7
PM+7:O[NTEF(=S8/_+_PZ;)@V58!$Y#F2G-594VW;W0S@YJ&*NB>RQ':H&\M:-Z%O
P/ 2BC\?%MB=8<')?U:3[C0YH&J2QMB;,V+K9SP&^\Y6O2&<N_><2#350V7?E+[)W
PAY1R*"4O:J-0TD>LAN>3M3CZ.<7__8&P&;/S:O# Z>KM4:"+AB+OY1% I-J  !/D
P->((-8 -)V\DG"\BAN/P&Q@I+AJ5Y1O7+!-ZA5T>E$]=DQ(S.#>]'>_""QP@PBY)
PY\R33'(^2?Y@E1)UE0I7M,KM9[.D*"!4O<<40S^AS^8\":"S!NQLV=""F$H%;W\Y
PXSZ\, O1CUB6F;Y,0\ >:5>D;B&MCG"X_PW4+V<A!J@:?!)'MVA4:T02N?PZ_;-_
P([.ZRK48O4#OP!?RQ;S"1\3SBP I<8FK.6( V UI+7^FAT,'D<*VR>AH;\HE2]S:
P<53%/N^5YCJ:K(TY0@8:<?YD//A60>(QBBP<LZ5VL(Z>3A$(X]Y-;@E8R7Q+KFC+
PO\J(!I+M2*(=$,(#(3@#,!BOCNME.@[Z*H?'.4=IU+1'S]"Q!A[1T7"/O>6!I4BD
P+].TK-U^@:CX@5+95U\H$)G[1?@4 F&6H,>%D_AK0VVUGKK;,,N?0+[@3>*]PJ5A
PPBIIB\!/"\:<M3&!&'^0@9C7<1!S-,@")KK_SU'*&7 _-%$CFV#T<TE4P/A)N]H 
PHUS[Z*%_2G0*7X$(##7#%'0K\S]/6[=,UB_9VHW'"IQF.VT"D;&_VC_HP*Q>2ZKP
P;TE:/]G*H0\BW%3>ZKHZXRH'<3SB'T=3VUS0/41DXLQ@9IQI+5<FY(?^ZY$,X?),
PY[-/^YQ] 8"F433'4[B#"_&5GAH^6%8Y<KA5LL'^X0_45]_0&M,T5@1H&68!,B_$
PAY3*V/O1'GB(<[(:UN6"F;V"D"FRE[]VH5DT$(T9+"!JM A$;WBO;4#*=,E41>%C
P+S-.@T+Z1DY29 5L-.MHD'+/B0$'O73&9\'J;'\=\.AP&0<0.F"*0AI/)I8D!L&@
PDO-Q/A'3_3K*=)1C=\J?G<.TSX6@OOWYPH\53O$W5TU\0MN10E]K%[=I $S>^H+S
P:<"E)SZCS^0C1\]^GD;YT3RW[@WCAQ&F7(U*,^Z%_IT1H[5%I<*S]%8D?.NXYWM(
PY\X-N[.%ASQ)!CL!&P:1<1B@!$_M,^VYU.U.<D7.-P?S?;:/A\>,8\665ZT0&XIA
P4,LMD5 XF/FFR[..M5R&U5/-8H!FX;UW9BWN,T GT;DYR:-EV?W^(#O83#/FLE",
P;'.9[CWN^ZNR']*XM^$76A#TULX]]BFW#/I\IM:2?E2J$:1EL!,#3N:W'7BS)0'A
PGDG "0S Z[/$.B-QI?D"<1+S>[>7]HE-N$2$/\U\^K%B208644D-V<]&A^BE:B;,
PYQ/[I#E\(5'L,+Q-6FW%P6D]37NJ1UTE!MBG?K$/3W&&U+)H@B:ZH]4\FXZGJ=Y$
P2]H+X[%YX\3,P(-6HL,3;K>8IFFI_LQT2@8QIWZ?( ) R,KRO';7%'"N>; H_[[=
P3V5M7RV*,]YQS;-B?_$0G,N.0/-%_+[OY4+K_"YKW;^+T1&RE":-I+TLCPV=/<=&
PO+78'U+":G>J6F;H7 +G-&>9]E)40.IW?2,F9NEO)XR6@@(A)(3Q?:R"6UQ<1<@@
PH4"=)5PJ*L2$N\(EY$2U)BG( Z7NUVN+7N-B\-FAZKC(MO,PG<[<NG-=(V>)(U"7
P"-VX\(HYR7(;Z]U_8@RD+F;W)(P_X@/:,4/(RRB+(*[6#EL\$]5AFVA:"$9QR\_S
P0XKQAT4L+AB+KD)6M7QI-E6-42["Y^Y7L%K/J?U-HREGD_<#>%L]H1J[*0Q;#1YE
PE6!ZNC:J[Y2+N8P[^WDQ(1[SH!^<\Y1,1K/(7W)O*EM!B.;=\DMO6H7"4^9Z4W1_
P'KPER2H-(6MK)QTZ()%P3F@:RO]:-BX?S117EED+/$LAH]^^(3'?685+TE14CM7@
PH*M@1V,%$RU,6KB/Q%S)&KW06J:]8\(NJ@W/I]8^%]43C0;$G7^LOV=!-,7U_>QZ
P3$K[DQ<VCBL=->E)5)G.VZGP16$Z[]V)J=P?J0QNIKT'M0U[@9V3K,\ ^K^>&)3T
PB8=W'WC2H5^"_N36RQ>FI-H<!RPH0)L_DBUQ<\.3HBQ+DH<+[#]1'/"'AD#,\YA=
PO?HV*&HEX($#(0LN(PUT;K;HT78.U86A.?N#/K+W+#O'M@"[>'0'PXX$B=LNEV&'
PC=@7MX\D?I0>,7C_KXIEY&!N';X.FJ_!-*;]*CU*K3;-@ 3GUXC&B"_5+/7[DQAB
P3C5PSYD=^?B"#U\\*&15:=VP:?CKCO!C,!_?$F!E=L>"L-/DAT8-Z0Z8X0_!=?6'
PO%[_4B<:6<KCZ!72 @!:R1)@4,@2M2#RB@1;8MP#9\*C:)WMO40T2E8^)DODOJQH
P?9!>CZ([FN2\.$UY5"P(,! 9D7V8;&(KE\A$SYPN,]/*4GM\IHR:)=1E(I;)1-+A
PN@\CL!DTKN6-+56?,<$9Q<V,\?7QTUA.Q<147?Z;-_?MDTFIT8.SU*V_629@V#R3
P6OV@:A=/-$OYI_(!Y7:#8X1HJ!FD-ZF52MJ04#:;A<;MPG@!%;T^>PCEL4NT;H\\
P7R,/+7J>] ##\U^FA:"VF%7FZQY]T7H)=<0KYF*6@'D\N:-$> +3!'/2_K*.FK09
P9#@9T/X_PM"@* M"[_2/18SW.D4J=Y$=2#GQZ)"VH54:7J]?%6\%P XZ\ZPI%GBE
P0'/7P]]^CU7BWCF!6F!\Q3:$4Z;FULT#>I>$R/98 Q_=:4,\T-0JYA(IY&3W&E9P
PLY>!W/\54D\SBFKX3?GN<LS7'E+89L\Y_MLC#&]Q!M=#[6BLQ7[<^8=HHAGQ)<L6
P?.>+ PC]T)/$AD\6I+N*/XTY#):GIM2Q8J2'-S!"AWLV8ME.!\B\,B@TWGO'7IE'
P.P(@J\04D]'\^!5]:W![N/PB#C '(1L\;:5^K $#O'GBA5WO\ ]*(97LG0A,RBF,
P#^;Z+:9T"[]B(/N<NSHH,*')R1JFB<#:KV8%,U3 ;SE[ 4)5MAI4NK+FH<*0 \GC
P,"5SA#':E:EK24G(&&-OD94,X\#-D)TW&B,[&BOK2,XYH*2+!Z_L\M5P_@4GR!: 
P-FVP*EO9=43I$Y"6VG++U?M:D;_4Z CR,7.\1,Q?#MICA&*$QRNUI05W&887=SSJ
P'AK'DV^<7R_<IH:[6NS&\?TA_K6&,;Y9LM@#6?_N0(\QDQ2S(66M3&\3G[#-#]RO
PU"PC(?/>!+LF<-]ZWWWYM!-T6UYUV>TD#>&.-E3=P'Z:CH(9Y4E@3K3Y[%WNL0 3
P*>_20Q@"M/5D;'"::0??SR-2[GO"K^9?]-%NYBS3BD[(61;2R:*TA&IBWG!Y>COM
P_) WP.5*L)[A]K(]?OKF?Q3QY0KMH(0XM]\]4+2_Y7[Z!4\_D^$5V*)N'(T]\AZ.
PI E;'4J5G<]96V;N!"JWT /00#^&! @]D),.:%1:FI1+64R.5W"VB2*PC+CC#'6\
P:QESESS$@/?+@R<0JKP])RFK;GOUP;888Z&HM(-BZI%2X/^,$=ZZ+NQ/%AR.%"'A
PS$^)3]KGK+D_ D#2:T0GE#D5Y0*W4$4R)2#^S]$:*7%2B3H6E[\-[ )XG$@W@GG)
PV-EV_@_I>. (X_3]$)90PV\24)/1KBM1'3@&K\5IIL+R?@RT^O2DQH:Q IT[B 6]
P".#KW4);D&>(S440.-G]CW2X^F^H>-)S0Z3K'!?JS1AHGA0?\U8A;;H#E$FO+IS+
P)BJ<]V^Z@!?QUMM?7G-&A1[,7$GKL+S5R]]R,0_XQQS+^O]4?V<K0E1*PCNJ#A@G
P#\P@GNA 7"29CZPW0/$<P?E=Z=+<27SR^/*<"SAU!$60V_;] ^R"E&-9AW!<$U"1
P+6^+W<]8F'7'%N[,%)S A61^NSC<$N[QD; MGSX[5\NWB76IR%"\J@C9*(X\-7H<
P145.)U,A?8.36LQ)QD&ILMN4K)$,@[5#C@7W LU=%,HRZ*VB'6N]V#SO+JSXO?S*
PY'!:''R3D%8N<<SYA=9F=(?;/-YKA1+I^7Y+!(YU\P T<U3(8'A1IOE8$0_'1I0U
P==N-5Y6/J-=#.;(MV,>Z,'IE;D(.[\VT])C5+I2<U83@^2'\8KQ*$W?J<_FR <,G
P4#E!J3#1*,%^@JD6HR4Y1?P"PDX$3PW34"TDY94G"UQ]^R1.OO>.P+6'/%_]L>D=
PO$0+#]?WKT9N07$I("5_ E<!\9BUI6SRX^<577G\Z.O7-VJ8DN-%EV1] DQVALBZ
PU*R-M8<(\1)RA #U \WVGY;B6SFK'1F9\A^1YA_X(]9>Z&5;P79AI&<8;B,)O>&T
P2]7 G"T8X!*E_ML)6="#]$!#\^!$8F0'*1E-XR\=^<P?Y=5[(-$TB843;U@TE5>1
P8.?[8QP?);6DUUD(?9"OY)QES*GP&?NED+M&3 6*DC9[:ND5N/3+5M2L$_PL=0!,
P9R/CIP;O":L IQ^O!*<H@4[R&^7I#7C*2C,17WO>6/-1P[SG29+W-06>AH+ ZZMA
P;/QI#M)44,OR+'*E164!-KIAY9MFAYOA_Z=F.HQ\Z2T[M,9]F&54=BT"/>T(9M6.
PO)W[065AV%Q^A9/"_ML\SBZX_-4-!Q%3ID3V"73BSXS:^$+,EVVUY_>%/5TS[ 'D
P(K@16X'MXA&CLD9%KSDB-?%3U'3JJ24*I6K&2S["3A$,L/"-0+H(=4%V3IQ[>!7<
PH5^X"31+I)MBPU=B\;H_SB6YU"Z4U2_##Z 684/ F"R3>2?3?$EIX!#G#]T[/)UD
P&6^>\GY"=:!-CJ1FHAFQ@Z<,*@ :5G[:?,V1'Y/6.'@5)?DPN/813ZAND!D-B<:E
P23\IU-Z:ELPDYTI+]C57;JLC4#WG@..WI@8LQ0#48A6@)VB5"[JG!\>K(.YBS)7)
P4/GD%*DN82\N_UY;WE\?@A'S:P]RYX9-+I$T"950!F^A^*Y@(*"2?,7RUAQDI/-!
P,,M!M:#G=.?9=G6VXX"IE2^R80=6XHNDT)%'K;50E@=!'8=7P(!R 0+T'[+"B$^\
PKZQ"][D)&<@EW_/Q*I!EA$.IA)-0>8W@A XM*KSR4>7,,B:QEI0_>8HV#)^5ZN<<
PRV=78X2[0K3D)JJ/R>BJ\"U<M-IN..++Q3Z>UN05QJCR";7Y28BWC9ZJDQA0BSZO
P ?>REM%0:(7L*V2YT0?.\].80 !W>71^/_AO&,#N*$N^T1P HWI,*(_DN+<WL']R
P@/WWPJASCF#2SK>,FH!(\!E3[6]_6DE1>[R):JA17O/BKK.#5+/?#Q-1^* X6N&J
P_]G-*9YUK/T@9UI/UT7'6KF13>2^ Q$?O03DR? ,^\P01 R U3U^_8J./ M;6FLY
P7PM@?!".)((4/3K$R*%(Q]&9:(SYMUI__H#6Y^"U*63,T.;>4WB<+.S8'T//\N02
P+"-"WQG)A-64H]1JFHJ_-@.FZP1[U!UMTFZ8C@YB'VCP!CY&_S).I?(IH^6E&5H2
PC*<=<,6!LI1[A>IT>TQ_/E5&V+5GZ)RS5@2M%J<FVM&)#3(HR&W7 VEKFWPM?H*\
PPNGCT;<JG<P ;BXM/S2T8L6AB@>6P3<0.(TX\@^]=R=%]Y0PM^*:K49^61H??P-M
P*XYRGES-1W7EZ"!XQ35/NVFSC8<\8T2%SGJX2TDJH01R]B2QQ9)=Z#YM=^.XK+=Y
P%@D(T9&8'LP)T%.1=]3(Z6ZZ ,;L.!ZW+9P+65)5,K>A/=FBIK]$H>AU ZGRSP5!
P1,DIAY2?)93>[<!=KI"B33F.AS['E=M]&(?@RE0DV2B-V*.Y6_S</G&G>N5 VW_G
P2;JW.;^?8)?60*>.#RZ\<2%(QJ[[6X1<&*,\SF#U%"#7FD^(X$+'\U9Y'^4<LVW>
P>Q9'+$O %1%!3_:IH%QQ82&@VL3X.2YLR6//33(=\M+,2V-,]4\DV35^87G;G3K?
P<R=4Z-/4;'\/= Y%['<O7/#M551_H]PPD-LQ+@WF4*F$[%J%@Z.O1WM5JHI-876[
P?E9'O!2M$B@@M :EK4M?<Q2:)3G6")$!@L;K<(-E,>3[U:EJ1?BY9NMH&FS,D(0$
P-EA;NE,U= RO_OFO)M*JB[B!DUPTZ,,"8G:\ Q#_A&Y3"CII>+H'&G=(YCH]4B1?
P<(DIGXVG()GD0<M1#S*Y/Q#V<E4F4S+IU>J;X"5I\E4X^,>CD^P>,8.TOY+*/\R:
P0U-]H<.J#YY!?5F =LO2DX$%:>S&R@MQUK/\Y\+*X/\F=J++\^)G?1[^N>PH[A52
P>1UDND@1SBFYJ3WE@4HNZ%E]0I$9[*)KS%B]^945 8Y74Q9L_ )4%G9&R<3\HOFC
P].]Q"G=:WI3XK_+$&.P''#L0N'%FUBL_Y&*U0P MW1N\90:@#BEQ,-9H86;/I[XE
P[G]\52I# $UR>T8-QK GVP+[_BDM;+R-;_;;='>_Q!Y[T[6.=1M'KN+GY@D$ONN4
P'2JN)*>^""CZ?/T*TZXQQYM;8^3N=4 JNEHYD.UE>7<$N-,N%LL3"CW6WOV)N-)6
PP;(^;8G) )8%*@2%UO#@5 ,993NS)'=D'&+SZ+6G;*QU1+"W^C;O"Z51KOO_]W".
PQ>5><+&;B"Y+V;S_E (O7P4O?BRJVH@DFSUD@TCIEA4-ZF"K&ZJ4>!N4EX6;2CY1
PF'RXJ>LV.LCCXTQJNI:GZS("05_FDE5?H0C>Q"*M64G^'C?._QQ+Q=>!6_)\M>[P
PU=$4U9[*GMO=S[H%JHS!?UR7ZZ,6>"#JB!;!>_L'T]*3A>C#:"\<08U!6!'$E0D6
P%$=L6PX0U2;H^C<$+G[0%>]RHU'O >Q#:;DLV2Y;?U5!Q?FY^")WRH0EW#+5\MT3
P"K#1'<UG4TLA"'D0'"L]VV4HWWDU/%>N6VP@4I:OAC&K*#G$ZC2))**2)%+P>$Q/
P+LNX:N1B+C?OG.S@PN>EQX%8H9,R2TWH:CT:-3HGT2)^[8@:3.=HJ=-VCP?/NT;$
P*P'Y'VB6"HTC#BWMB+U>T+/.=+G[A-IPI&B19MEZJ4FB[<1"$B/=3*E,B_-^PH3H
PNL&2GW?B"(ZU(L7"AU^LK2&+./ J$F*VDB'H5FVUC_BGRF!($+N-(WD3QN$TP3#U
P(2?L)@Q^=9_#\ JO,L5KYK^@EB589K!JM#[)\YK-2(VIXX!&!?FMV 'XA0XJ$UR8
P&P(?M(??1RD'QF,^BT"9CM/8F#[R;34Z1:8)'WGU,<*P&!V)-];D?E5!+DL$&P"S
P3@HP8.,J.DMD)<XJ>:5DRZLGU;7+IL\W5/PDVI3^_;H=7Q->IK YB-X\S@E<I47_
P_8L+@>Z7+".-;E>]<" 3R7838U?Z=A+/RWJ3K'(AWP,);[:"$7VHTN-$NO,AW92O
P8EAQ<[08CBW-3;S>=E4C@@Y9.9Z[?9>XF2#.\2M#OOX[2[5G_K[9K+TK-&@7_X[[
PN,66'#XOR&$%T29RV%QU!HX1VU%:?2F8?M2".9+6E2<R:LT)8"B@+1,K5X" Z8JN
P$&&+<#B]I!*_ ;(MV#:8^_2#_H<_6VM%]?COA88+F^/ &IZHP:E'9\ O!"0\1F6<
P#'G5>ND=7$(? N C"SUG5(0 @$7@!1JO"#L[2;[Q*#?.MJW'?.)A\UQ!P9"_CZ>#
PSM^TQ-4D09VSQ??M4;\21TLT'6XN+(689+V-DB4974XC432)+-4*#5^8VH;9W?IJ
PO\I0TPFUQ)Z@/U($P KX*GSN-:F@#*TD1C&#$6FG&Q/V1IM+'L/MX0 9*73-^E7L
P /%TGT96HT-)M4PNGW\7 LV'+-7W>_'$Q<D7\'QS%[G?&.RAN,NA=8^Q.^[5].!T
P&04J[5YR=HI4,6EY:0E%)XFY.(<G9SM,@UP6NO_$# (_SSN'(/ HL966IYQRSW(]
PA>M',!^8B.\QZ:3R0&\JL5&)PH]3IU-^<L 25-?K\1O2+^%04Y#W\Q+"HCF$R*;>
POL\BE&^BQ9(6?]*#"8%ZZPLGNL!0']*Q/V3("V1KHB9KJEP[K17TC!/& $RXQ++Q
PCJUUF>B"D,HB$(54W5,CEB4)+*$AEYF>QJ<P=>H$)LJ(L")WTX*<)9/0&)]OWPU)
P'W2:67QFWF0LIR8802[173]+Y!7B:VUN%^83E0"/?M 8\V24UA@N$>EB%M,;2#;(
P]ODPH&2?E:W^_N2Z_6V=K<';?=!88NV!8;CQK+('"UW99KL#"YVXQCNSQY_V#/V8
PJ4M[G0I[%1?/[OL7\O5&D'EM/'$?1*[!B<% /0=Z[G0KSU?=GAJ;F[+GB>'O]=3_
P9Z +</70,;OMR(:-3V_$V]7KZC0JD^DA.Z6J31PY5Q\_V_/D;VW*4Y*#^D.R&=P'
P',)N^](@/C%G</9P\%-GI6N0%^=UQGJ<D6M:2P_*VSQ[-==W91N*K7L?S$+BG (2
PS05\";(7Z&I8#&0H41H,AYA<)'SW_CR5YN9V]R]+2%<D=524*LM)W[3WZ=,%&(:H
P5:KL8%K."*\7[XW/R8 BUQ47"Z5#A#3T>6&;E50"*SL145X.'/N(-B=A7YW["Z-N
P9-(F-.'4KO0GU9S&\^G[ETOVW)G?$I=A;\GS67K*-<E!J8OE;-V*76EJ8RYM9TE[
P,.V:P41Q!4Z/R8">P3MK;'!-RAF;BN/CSI9$'BF<-6E "M*J1,*<YL!;\PN>(G+5
PR- K+@V)RN(A72D0"!!K.;2<F,!*:!].@LIJ/#EL7Y 0!6(>X!+O_C)<O6*'1>5T
PM9_#F>6DDW&VYA#<1:M^-3>UW]>C#K/&[7>^]_I2XBR-^GZ,UR V^P1<=9CQ!ECM
P&]S>X,L+]==>NG)0UX.=KEP_"*$2#'%Z7)!JI,_<M.+S0RBBP'<:!-0BZ/G/':VP
PD!!"JFS-WZ>=G$#)XH^0T@->N3E?5(:AGD6E87,1$\%AJ\6MY#)^%:&[^Q4S7APC
PD!J^QT%V,A.?[=HB 7N>A\^K%A*_@'R*[)H=AGN"!@-06G#"9B@F];M$:!UBG_;>
P&&+8M(%1;D\!]W]VRON#5T3I R ),"UR6^;O_U,K(\4NQ+C?QOHU#T*DW,)%?"VN
PN9-KZL14A=H9LEUDCL0WN8H5&/SP,U+"PW#_\J11/2O-[(W%#KCLVB5,1@Y]KSS;
PECEZ%Y'.(WVT<>Z)2<5@4^.K;?+04J5BC#=RV+5F$W6Z?&DWP+2^U8=4KA%Q0A:@
PJRG@:P\(!#Y=^M[3<8Y1,3W4#>D1!15DR^2;5:;7E5=;O7O_QHW"FY8^IX_.=0!$
P'2G, /9LVB"?Y,-7'M"E6A['_W8UWSW.KS8E5C.E@\(BSB_AZ%(K3W,W8,HD;2>U
P97@VOB0!-Q,M,?@F+\@S@/(PVS:O)N)-AKV!17!+T17]]/S[QR._LFZ6MP//$Y $
P'A)4+K^#L@N3S<-=E,-5B?OTM#,8JQ3>S\ZO,R)F_D1<_VHM24?BH,@X8JAT0S+:
PI\)</R9@<?>,[)[$Z^X_G*\;>'+0+IV5]ARF)O'\0RQ37]%Q.&\10>KU)_@4MD91
PB9BANZ]>JIO".FO3[BWXAFHB>OO_AX6UZ!%V!T"V,C!YE"O?-A5A-#DR-V4L]),Q
P.*'J\DSF7D@61(]#!($Q'GU=\:??4=^&6)@KS0GW%[>CJ:-JE?-HHD+]"M$QOJU+
PU+U9A#>DZ( M@2DR+PGBVN*. W"\DO $M4,82-L9V-:U+?U=Q8ZED/#@>DB.W<5!
P_'T!].SM\<+I-Y0"I##*I->4M'>Y#O'1]KCI4U D-^_*@'"RXB2R]A 65L?LJ?&:
P^ZD[T+)-J/]#]'?KQW9,G!BH=N^!/O4Y.7_26QVL6;:Z'$]\=CYO86(J+W?4Y=+3
PJ=*M]Y09@4AD%Q3\6K%(1^3_Z?&85C1VBG^R/0T3J:$B+27\5-.52- @S23LJG([
PB:1^L:)A&"8*(.LW0 =.-6-F!V*"U)X&W2;>:G'"$/7H3E=56R[%=3*R_8L?=5JR
P(AR[$-PV^#>Q231&1Y)/-8;&9<]7&NQWAOM%UYDB30PSBSJ*X7QUD+J2D*RGL4]V
PBMFLT;(M8 @S?1.Y&^9-[SZ8GF-)@%_;WH6"K)1U3]J5M2N BU6QV"%(FZTHBVBV
PP[1] RT'>@HRW:1'[_0^4N$HA=7<-,[N8#)  -;A+>,S/K"N-G1!H,'*Y!JZRBO4
PR< (&HUVT.)5?:F\GI6'>6DXX(E0EM@R)+RZ%'-I]6H=?8JU>+!3^TVIC*C[:-WO
P,7I5.*3\CXUMRU,\H6X-X6=MW_NW2M!IMJY7^_5WR$1U[1+1.EWWR4P[VII)[[DW
P4Q3W/-DU!/ R $X!>MAQ?*85OH1%8+G4 #EJFUNC%O+3_>R"='T\ALPJ1&W;6*-Z
PRDQ<'R&Q)D,.&A1NW,.?^5YD(WM<-<KB&:VCN,4F(G&@,6<'#U7 *XAYICW:+MK2
P.,VC4IUJWS4;O99=9M-GR('^U%\F\B,8752K$$\2[.5,5])]DDN[%(T5 4'+=\]3
PPH6%MC 3+:QD-Z9_6SK(/PR/00K[MY6]9HHGEI!(U()?L8LS&1900PAZ<S\SPY*U
PI>O7>#6$'GNV4BY/NZO)#!V$$ #A<D *SE?86$.:*HRG(;U_:TGL8AY]7<R*EHH[
PXUSG3"]:(,4EJI(5U9#:LNYXLMAH4'"4F;;HG<;&3!4(-!6Q )NF.%7*[J5UW"+Q
PA-MRW&'_/]YS8-=XS(4DS?1JW]ILU'":G<3(6C\@:)SS1BLNTUHDY]HG6ASI5;ED
PTR/'T -3CO=(6@HW]]S[Q\:QW;LZ<XTDP4K60&I-X'HXIV/[FE+3[E](@S%)1O.;
P!2FT !WN%\*)?8>7D/-)._+KBEI;&C@3['UYZY]K<_; Y8P.D?%=MB$.#F R[L$M
P\1;_IT!^J/'N)X91CLR]L*S67XDJ^ 2V**%$M*C]AKSA1,/+U0W?KKL-P9]W<\G.
PU2([\W"WO @COI"R1!@TD82I0[NG-3('IR<6%T;7,YE#10O$/W^(CM[%!1-5])C@
P$CQG*Q?>4L6KZS&>3-:VZQ^I\Y(!IF%L'R4#Q0;==LQ_OJ@2JLQ 7OP;=+-O<I>Z
PCJ3^*,YK'X'^9% N'ZV /$QI@L0T"@5JF&Y,?[^&]T='SH""[=?=,9M(!-;[IK=>
PU@0\?U,H#,$T*A%R.4J_2X#0!FK_)@7VHD)(UBD#CC*4M"&,+-_I/Q/YP;PQ9(2\
PI792C6/1>7FHNMIC]4SLQCZ]WVWP=V_M:@=3D)KU6WP@F#V=HR!A8O6DA.W)[H38
P\-+>5L&R1#XDS6C@_CY($ETV9G-WRVPE:+V@E_N9724^K9T8:C-GLD8;88?X@ZRO
PDC*TNJ"CTWD&M;7NKK#>0QI<1"5>L5[_[.[K=>\G^@.86J@8DG&FAE+M)1YJQ["E
P+;P8O(6!>@XF'UM?.&?T>$I%.BL67K[.B8A?W:51' *O/38JIYHI_\?DY$,,OR:R
PQ=#+?2V_<L74XAZ@5B5>N5HU\U9W*$72U$56-0\[98BT4R3 AJ^5?CLR*O!";Z[4
P::Z*.8)/5E\6>&Y!AWP9 ::SR2&@3GU8HJ<#.X5H>LP[ 33[0;3Y!#F>O5H2YTM&
P!A["7%^T)A)PT0KZ/!)QU<Q5L$ O!NF\T?-YUZ\\^A%8Q0</IC5\MPETVD!^';UL
P*B1![;Y^R,1"I='9R! ]^>H-V,!8(2CPT&F-)8W,5A!:<-6.(Z 5N=3C"6G4,9!G
PHY@N'3,&'W#78_+*C<&3<L<;;N:WC%+_XFDIC\.K;2DH+NZ+DV15%ALZD*[ 4^!)
PA66O>]U>S:1\8"8FJ;T35\]+_]N[6M8+_%6EOAZ $XC99W+(%'<G.R#_]B6?R4V(
PP*85.R(+ W3J 4/W,H4_4GQ$23F@D.M&T]I#R!A'>ZQB-!OC(I$7^PZ_DDCKDC M
PQJU:5UQOF[AA#H2PUR!PGV7)$*:X5YQ3E)CB*?N2@>LHQ2T$M>Z3RK6#0C@WBJ!0
PX,YC W107ZFM)?6"SJ@@Z[)@0GX+Y981!WAFF5GC]?)0K.LTDKA:P-IZYP!9GJ3>
P,S^U2M^X!T)1.9T@X[ ['D'UB+O4KWE;((3^*1[EGR.U<7;_./<1[_4J@G?6Z3T#
P+2E$A[/_6B6J]A-.G$AI54#KZ2W8!OP<D<@?Z1IB4TC*=50$QEEWUEVB6)3R[MU^
PW8G4&;_8HB#(&Z,1DII36YZ.6;F'0WALU$I.\=OM0,P5S N0SC7X2';^VKLTK:+H
PYFTQ7_!'>]$#]MG"5=X8HN#/U7$5:5_&2FH.=>;FT1<>,_C^MVNF1I%C'@,'R<?C
PO+T:#@=TVT4M(9K- T=#GK3]+:Z!"4/4[*:J]Y>WNIMA9$@)]VLI<<Y^MG<B3*N3
PQ'VX@=<)VHNR=)Y_5<@;?IBOA-O+6A@$&#'X>C</SKP<#]JBUR0#=E+Q+JP8Y_\[
P1ARC,AL,F/P!?_5J28<ABRR&%.<P+)O@8=N+/U%JC=^S.X/F-MR, SHSUW@FL'#4
P1\@V>KAV1.3,W/'HETJ7\U!CR?8PG#9HUG\,7IFS&LN'P.=3RWW+./ZW_!&^\:#\
PYFH2[2@(81V:$-58?[01E.>^T\ )CWD&8_AA$WSIN_S(-6W$T(5N=[K5!=!$8"65
P;4CYPMSTM*"2X1^?^#%0P7J.Q][4Q/\I+%&,7V<9O1CFQAP+-R:+%H?_>VT!Y[9H
P^R*VXZGI69W%S?-+KF(C [![@2+V45+C$A6_K*,5S3RR)AF5H JJ0]AS4RU!TN'$
P&L>37P'WP[JP  -8K-.O^([QWIRE2H"K;5AR^B)LWG>:X NEVIS'.O]4(R*GQ3"2
P')CBE'51=5CN?BX]F560BQ+3-$E*J?>'6+RJM6 6Z'N>,0)M3)C2F17ALSA^13+1
P093X1MC\1Y8@@;;?W'%YF3B;D$.+R/=="G&<6%H+[N&L4;D;$("\?DSETN,=(1TN
P7O\&YGB'(4)9#(115E?VO.!S.-[X%N=7E"3S$4@H40L.3E<.5;]\WVW$ECF>]XQF
P<VD,F&I:TK,Z6'D;IH79%%;,PY"L6<<"&J;GV@#.K\NG..9Q0_.-4R"RD/*76*Q8
P+ XA7.ZM !N=&.&T;Y\?U>_DU.8.V]<U=A&6\K)0QGWM$GW4SV$4N!E"PK/NU[^*
PE%FXS@F0X1G&476P)<_4S^?BGC.[O0?7O_C=-E?\ZROS(32;P"[,@NF(3$-M(4R%
PK6(5LMW 52@O(K<K9A9?BSY)G0$\@PWA),O7+52#/L!X_.%-(7V-4X]"MTW[HDHO
PGN9U3KW:D>GR0N4[YO? K"^AV3.ITRX0B'%4-=HX*_S]%J>."KC^%_'2U)\/3<"V
P=@_T?L+Z&C30""OS<F@[R7M;F1$.Z.X?>%TT:MNIZCL-=Q\\!703,2E1 86.S$.3
P8QP)#_N'1@<WIP'RNAZ;9[NR<J5-D'B'$G,#W(@H%=<BZRPP5)S6H04'3*?Y!MZ&
P(N_1-X#M+0!9(52O'E7WLJ<_Z:U6X-3<U!-9_$#S'G[N]+JS/,?V5_7>TZCT[+A1
PK3-EKJB"T&N:9N1K02ZMFIPX*RY'L*5((U[S;)X8S!PRU5F\8?:C7(G*$*+(^9_R
PXC*?(R3,C$"?M!SE(G3;/G*]\EBXI%N8MCD)!CZ,="DC]KO W+'[WTUPKK68?=X?
PBO-5]?.36L*@XE=?LE2-K%.V.7$7Z$N%1RX!Y$]Y<2((S18%/Q*6$=.'HELYH6YJ
P:W[PW(KT3L]3+16CVDI'2(+Y4+"Y$7+,8?U-]YT59W?M'NPH=[; 8-H.%C0FFU+A
P+,02P_5T)4$"@#_V+^\KPG\<7ZV:7A7,0V,4=@H.29"EI!'#/Q7/8)K2SQN]TL2[
PV[?8?\E /$I#@^G;#SL&@Q'+)),IBV:]A+"=FY22;$-)K:[Q1FEIQP?!_%:JXAD@
PC DD(O?9?"R7W+^3:7W@_]KQ+PP!9)?QP# &SP+Z,'@_I@WA61]WWUS'$RN<0T<\
P07I[G'PPH8Q&5(N3RV%T**CS)S @2M5.5:E]K-KH1"UFV$4'-?GP86%LTJ/N$LJ=
P1T >TGEM1369LH*CUN"\._,-S*@VJT4L40HB$Z1PD#1@Z'7%#AOI@WS,\OJXS49Z
P0O-""J?JZVQ5G ^;SR5+B\9*]_*9")H-III.4(&N#Q)$J0%SH%4R9H)75N+>SER)
PB:=# OZ[HT+GB="_=^&6(]F".1V\=ERA2SX&)W:?Q8+!N03 9,#-F;8ZIU)_!<8J
PR/"^U#3*N@*M7-&$)DQ$F4Q=)&6?60"WS?%X^7,UTQ9"NI"+#(II?HY4!>!9"O; 
P*7L7=SI)V,##K*1*KC.LG^5=CAFFU_(8/>9*\$86HOB(ZJ'P3+IA%[VBLDV5A_TE
P5U<FF+4G!4Z **TNG'/ !Q.JKH2:[#2 P+P?,_0#.F"B@JET'GHRNH.8#6'8\M1S
P=)!U%*#=#;_,]HF*Z";\\@(B^BDO_LPI()F/\0P< #EYDFPOZT(PV^1]"1,$89"(
P>'/[=K;!CM-?^*FKBP>ZPKI^>H[C9[YXIQR_2-X[ ?YM0U9'OBB4AA44>33CKV[9
P3@C!]#F9*IKLX0(Z9;8SV4!4+0^\/';*7B(!VM$Q'IV_M]13LO>:7KR#Y,)LBAZ 
P0'EW\F:-\3V=JS?CUZ'X )4$O!VOUG=N%.%O!::2^J$V1</O!?-X51=4>)(DNC'C
P;GQS+?1S>G!9_KP=D'::R>EC0K\8+_X+QQ%>VS]&E&X[DXT*+B;GUWC5'[+,\&2T
P@>6(Y;OZ$![OP:R)SB[AC/3,*.=DVVS3XV@KX(1 K\W&\I0+80P^N/0^CGL][$U*
PK1^C#KTOZ%4\GGD!W;T"F+^0-V8 +V)OY5I<%596]O+%Q%(5.SN$C=8N:28%S6@J
PS0)'X.I]G "(=H)#AXE1V!#>BG:&-H0:UY#;@/ KMS?0]/LZ>$ZA^G]7>&$_<B23
P@?<N=$6+&5W!$MS9G5:VSWFLQT00%BJ5K6%UP3-X3/4X*CHCI;_EJ]J6&--!<7)K
P+TPY3[ELFTZ[.L[S =]2O[]>UIT2)_!R4D)QF6_7?NG"IFOM)<,NW=#;<_0UR-,_
PED=(::JJ;"1W/U&SE%3F"UE3""<@&B>H :_B'#]4D!6%TS)P[,FJ[APGW;5\#VKP
P#.QM4;2%?(J=TPS&U3X;U%^!PAJ"JCI:KR*I)YJZ>^!C.:_GQ5K2["G)5SZO\G0)
P]R_):0!<Z$K.Z1"F!4/>T4]UJ)$'OSN"&Y1%WHF\(J&UB-BC$FYM4\$?QQ$*28!I
P^# FJ=Z=-MURCT;L0J[OF2>;-E5'1FLRE_)VDJQV#:'H:E>6Q>,R $7X35:<XR<"
P;D_Q1HL4GBIQLN+5"OR1H5Z">P+'DDA2&7+9@QIG1A-[>S]1HH /@55D;5.PFEK%
P,')8@?$&V'78F:GKMM[I>!C0D]=-G24L'1U6V"W"6+*E.M4QJ!R+4RN#W;-0W?;P
P \FCR#/\(VJADSM"##37HODA/9;N2:KH1JD^U*%F2J/)X',\20(5 YS(>VP)J18M
P/5+W2-B E4J9U6:B*!5G"G"A!-M2YT\3Q)/7NR\HSF; 7D6<F'D:M&W2LJ_[AX_E
P+!LH;YS;=F8M'SK>2,^ _IA.O@O\&2)1=#)H?"8!A+4%9/R ;:[M8&Q(><_P; .4
P-I.JM=XWU;XK0-&B X*8!+,F[RT)>]*E<&U-BW7'$')N&]TGE:4.Q0I)C$OO6J4M
PFMPG_7%8X\B_5;Y1 0_9W#!*8G-0CFU K2+]RR]G79=12SB<2#W:J5WV6?']5V>B
P\C7Y,&)B/$S4_HGS7WGR_-Z%WXNDDI@)GMLW5\@8^]\0 353^AR8UJMS:[D+9(!5
PXY^X66 02E:S">E 49RO'9N_B<BK(^W/&H*#-B=N4A+S\K;5BK*IO0.&HO[PY/8E
PA#XO[V'@;I\40=ZNHA!&RR!NQ4=F+@C@"G'39.AKG_UKI]Z<FE$L>PQ1;4>_3GTG
PQ6C9HCGBH-T;$=:ESU1F\4UV5EJ]T_N,1RY2PV4SP* ITS]^K52([H*V'IYJ;VLN
P;QLU.K6<J2F9.3'7&0LL1EJVBSC#57+XTF\>FWYL9D2@9B:,/5E4EB_KV;2"?%K5
P3CYH0I1/D\X1"F R1AJ,.\<(#Z#/S]"#'NM;L]DC4J\(K@6102FP"(;U&BF*RQV'
P%1>1WU#_#@N0,:!Z&AL?6:40=E^$+50L /-/7IJ(?FNXF^/A!E<L=!YI]\/)6N"L
PV@]="5S2Q(J?,:9;/'EQL-&A$AG:]!WEUI)38JFOD)"K4)A =,@[X+>?@51F(4XD
PYGU<=.[2IR UI?\?">6F>P2TX!TU]0W#I<]C)07^I$V+.^&TL<N,8%01]3;O.\K\
P\V8L=%;>]A20"(JM+7U7B2$H_^RCW;FA$G/BKH6MY_A?LK+-<N/<T7G0N(4.8]))
P*B#IHT&"#P48_HXAVFWAYJ6'B5D8"*/!<YAUP5@&*_2^G BI",Y_PP.8?RUYKVE-
PK##I^O=DM7R7Y5=O=Q%HLU^OP?O4C>GCVLL0C&W]HO9K+253]/[F [-!-YLYQ7L?
PK"@F=RYC?2F$=XPL3Y'A=MF((O&T );Y+>1SAR:BM&Z!J?1L4BH^]2$P/R^ ^GR1
PR6P0KR!Q^INZC:.X:=^UT[:>22!%R:>LV(I^#@"1K[=)+%_L/]Z01Q$=:TO\_GS7
PZ-ZO',#GFH]K<,4UU^X,!\3 .\X13V&BI 09?"']??,B@CP/>R>A;9QEUZ;4_(>X
PT.I*!,&O%3",7F?1U%?Z#PBETI@8<%/(B;CK8=CZ!W'D=VR??2F._US@U;4EIC,=
P'3?>M0 5_D4AB>BNI?HXX!#T1W5CM5W*C2V+O2=4[RQ<#.B1N8 C?[6CYS01!PBB
P!Z=CQZR1690M)?@^XYIK4HCY#PI4(N@Y;==V1\HHT.]]877 0O<MTUW"?PAKB[;$
PW@9T(.IUI,U)ZA1YJGF:MQZ?!'5%L:T6J,,KXEGT79>,7CS\V5"DXW%>Z%45/[3!
PN4%5?W$"+:_"!@JH 13NE+H-15IA^I!&V1;#%*IO:,G*&'GTBZQFLFHU/FZ?3ALC
PB4FU %0;#8*(IJ":3'T,T6$WI692)]"]-Q1EIK<A-7P2,8,OSZ8PF/(1XIT2J580
P26R[NYS83$SXWT& L=W*_L!J.=F\KF7G1D,Q%,<UG;=,:4YY/N+89?&$LYIKYAQ.
P5)NPM#OJ5C=R@F)18A*_ECLJ%5\;XH%*B_?" $N\9; X"_"ED+L",*1%IA:V:CE9
PA<DX2K)/>Z54[YPB4(BPW?UT)"(N3Q'B ])D5K9XU08#4O^CS4LEZ7 M*QGF=/G4
P"$4@ZNORZ%(LVGY]8=";$CP64 @5FQ1'+H8!SW3M97WL2R$[W@N5!Y<,D8@CWJL!
PA/?A6:,4E.J.?)FMU6F(I90L*FM/R N:#NG$0PI;'^K;!,+/R@9""HZ7J6[%>JF.
P@+Z'B,XQU=J3) .17R]3'+ILT@UY5AZ/E-N;,3'.N.CZW'_>^9Q.04 O/F39H)S;
P%[M0F?S&7H-VGG!_LQPW<@[94=0D#7;KA/ -U>E^#C"MR),;\T& ,7$H_9!@7#+_
PPC+'1+@%MP&>6NL?$37]DP8$&S#*6)@D<:S'8ELO?C5#S6ED&;1AT!VK#C0E,X+W
P_!5<ASI#I!D#A!24JCRJ;8:!X??-B7AZZ5 <>)P/2YLY]DU(,?3A)E!QTKM29.#L
PW&A6+7&[K&F<?E-D<2\8AZ(<?W66E)R?5@5SB;_[#[.C66&*Y*<.:0VA>1(/:@XI
P]DXS&M(AXV9^0#=*75O6!N,V#@(N:GU^HCPF<2W8*F1SU1F.$-[+LI6W-Q 4Q;$$
P>BGG= 1>)6\"%Y(Y,%:D&9HF5P+D<72@"\LU>F_0B5(1&9;W):94,H2AOA?-5D%S
PLQTQQ@1EL9:$V"Z\DSPBO[!\94Q5-BP@_S39F*H41K!:78LKQM53>-SF*Q]I5*IF
P6MTV9G+W#S%@18 \M_MXD.1/44YX-#-^NNU?0FY^HZK[6/+J;9!5N7EU=/2"&.6"
P3+$(IBOT73ZE/UKU:VM'JQ\:H P"P$NPWWL-F@O6DSL"" $L#W0\1QYI&7O88UCD
P,?PI\#;D^4"'8INU0&AMZRE"Q=ZQPEKO?<#$#ET 317"06;GCR$S7@ZKPCTKC"Q$
PIFP+]LC<(P+Z+C* K^R!"F%F9/G/J/DE@T0B.1:0"O%_7&8(/PZT(O=OMCH$?F!?
P9NH*+N5?QV0D^1?XT!PT8J&I9'3.#,82?Y>AT<P5/JR%N>VE.$^')P"V=M?CY!/G
PH;/$)=18S':LKF'!YM\I$.8<,]KX)\:N3FD)B5O]^M8Y/'O.(AI1(7/\QV :G=&M
P;W?7-XA"9C>,+-I4PUT( /JJ\^/01BRI6.*I&$BR>V7I0:N()[BB!<$65Z\7&-)I
PN97P<3";3^@;9EI,X&/,I!9N&[:)J).9*\!!Y4X0E$$"FTP/']V2V9^]\I/J 60+
P:_0KOVB!FC7?01EF& _P96#]-.GQL-YDTGNJST0Y^\YX= @4>?:2YK.89XREC=A>
PEWV]0XNS(!.*-,I[*8C,-#%E1:^Z!DR1EHVCB_W*]B;A9/R$YLVD4H424'KLZH/7
P;WI8>LKW&M!-&Q=BRQV88#I()!71#Z>V_57<5Q%<_!SP 6F]_!.63.U0-4RS*D]\
P34@EJ*F5!'\/G>H_0E6$W>W98#W2G":RXGV:#S5H;;[6O<H(CS64]S[J:_L*4>PB
P._[]3L!]V5E#QJ9%8NJRSX%&:->%TJCO@'S:?4FM#5]@A+##V9Y 6QW0QY'(Z8YE
PMQBH;R@/?5ZU%7DDO1;%EM!/QKX5!FX.L\A&%E,=&[*+38:=%TRD7=4GO))?Q_>"
P8;AJUV6/C(AOVZ"GMVBR\GE$D2"_C/\AON#,-JT@I^_+_\__7T9[)XZ'O."0TOXW
PC<\+V^2[J%*+=/FR#(TKHO%<L%PG:FSPJW9R$_<;94HX.0UNY\Z;.(3L3L9J#:6;
PF:?;DTN7$,K#/!*0<O^)@Z;L&SF?9E,<H(&=ZC<^IA6!'U$YCD >G@LX5]AF,Y+"
PF,81 2*.S/+1ZJQF,59!1M366C[\D]F[KHL:W&>9I&SZ[E^$3C3-\\?ZTG/I01>A
P#.ALK3!:J"CS-RAJ_-B^F*6=P%A,6*JG*D:@;*+_Y)P@@'*]TV5+CW7Z'Y#BA6(*
P,5$]$%O#Q(=ZX5Y^ZD>MYF._B*K>6'X7P)ZZ# QK#0J/HK(1U"H29!#):SZC%P1<
P#U'N&$4[8;L:_P@R7M7(C B$HR\W_W3KU#;?H"ECG?QMOA..\ZR6.$K0>82VI"4M
POA(6HU(7K9SNQ-EXSI)26U6>9._/ *>5G361:\@MZZHD;R\:"*,J^.>@;4P:JJAK
PZ=B@KD)0&N5Y70@.6*F=:9@O:T&GXX,NR6 ENALP^<"@524"7F+T4@<3)HMU.9R-
P4K8!14V"^HH&85.4&-+5*Z>*4D@3;]5\\<AY<$WN7P@8L3MV7X% -G!],T"L,19P
PWG:P%N7BT*T3>IPQ2D1B\_>;RE4U>>;AE#D)>BT]SD\J:<X;@X14(!@2B,/$!OQ,
PEG^]B@B7]?F$'1U$1MB+MGO $5-3W'YV8#)H03KU?9I-AYKD*!2]BNM$1/9[?D7M
P7G>1/NCRC.OH&UPH,3720(J=K 4%")A2(#^*0L&;TASH^<#"/;Q8R-&H+B<JE-.1
P6<C.,_O<$W^GN$@/.WTM#/#P5(('>C8Y_1:T=V?80 LIM07RBV.,@76L ($!%R5S
PI!.)/YE4 DV+_CY#5C:!D%LZ!J[YD3+\-T,PS*G+1$@W5[_"N\J,^X!L <UU26X8
P4Y.I 3A+")'<,*\5;,CKIT %S(Q^[MQU9V"U 4O*-H^X0YF?Y N6Y5E1@0$,/[ #
P\%"$N"TTDIQ[D*RNHH];X_-3*%55N>%EMMNZ8IH K;VFVKKMO*!+&!IJT$M"1V!S
P'[S4-Z?KT)?929+?0ZA=07N'*?1_V<[Z%HCV;KJYP3ENS!/2OJZ#S]/DZ&MTY0;8
P)^): XM(0#3@C6[2FS]Q]8[$7?JNB J/CB:7BG)2;M91XQB4+5-F[O%;8VE%@&HF
P)I2> 2 $6Q-V)]8 73H[&M:[C$K.EZ]*R1.1+DF89U6Z_HJ004L4R2T&QY([7]^!
PA3CWPB @P[S7W^O$I/#FJT/:_8#B 5,EBKZQG&DD(5P=[VQ#JQ.^?_% ,RBNTN]4
PU%.\HT<5>:JN^-D9SA-HU9@J#92O(D2==")LM3-#/1>US%'ZO9$7=ZL_GZ3019\!
P%C'SX'L93^!)$/P2 V_P0FFF1&RNE@3AE1CZB?U">;NVK=6QLOK,+1]4.%Y(4WUE
PLPX4+K$2Z4"+F L<#FB(E#T/*9W<<5E!S(ET%/]J;>^#R]ZW5E!;P;FX#PT  LH'
P;B[X0@HNNZ3O-LO8-&$<T7XPJ,A'&&(%J2P71SZ.I_^TV3V291=#9351. [(F'&!
P9HNS)EN$*:L],-?JG0Z*DP:WIF AN&7+P-\]T16/OJGY[!DS+W3V\>?,W87.X+JJ
PR.S >15F>BS*O"XB.!F9";X9'Z%CZ=9XCR)QC=L1SRU'F_AP,6 ?>E/$L]EY4V/'
P*MZJ.P8$8)FOG+KHH>;3B^0W["&1/"_9@I#K\X=M1">'3LL1!CS_'3 AD$22APB;
PSYB">D0ORY.%CB.!8^<.&<U0 HVI1\QP[+"F^%7XY/*LU_BY!&?TGQ<V(MK= R$U
PY++WZ&C1,@.O(UN?.2@UZ-P#FGN039N5 :2/FCX5[?(L#-BFW?"QBS/XTL $YYP8
PWI:%1Y_Q!_B[BP,=ZN5D! ))4- L3G.?+O?KT^Z:+.MKI!/'@?OS_I=1S&BK89<:
P$Q%UP,9]\/B QP:^/XQG,P+"N(G_'#!:T?KH1;AFZUSIRP,G;D6U1%87W.UIZ%\*
P*Z!I=>2.UAZME0UP8N9;#_ASM^GE3^4\?>YFUU/$5<PD<,7'#>KWE0;:9F="%.<=
PH,;DEDKN2\O462WO!^)G4U>G"SY315+!43JN#@X5UKVE)G%F%?". ?BR.X3RK0-R
P^8X+//*1]UK%=>0O0;RZ5',C*'B%.(H>#4&37&GQF'L#LB \7:BOYDNFY*:<UF?;
P)8/C)*:LS6A1P=:ZL)]>TS=*<!?PMU57>C:TQZWQ_ "%=S]7+AX&_*8P)H]M:NQ&
P>H)ZHL%<'42>5"']_9@5"PF!;<G;YO$5.1X]7B1Z0U[>L[:.IF[^9>Y2F_PG65A^
PR&F-SMD]ZY+5DLL'WJD0=?$S;(>)O^050.Z C7.8.@&4Y=R&CJM7%M@NO)H  %2,
P*'2<9/O$ZUVLBBT?GME[R:VFO2*,8*2.\C_]9]._<NS%S[+*/D2+0NX7@33FJ]@*
P$!GUY!4YYQL3*N,K^E9VVHDX[1G' ::3;"CN&X4;:U$^DW]F;(F;AQ+>]"C=-0<)
P9.#!K8W7 JG^8>2CYR\*A2?@OFS'9"W9- HP.XB#WGQ>_"+<<X#$"D &]Q 4_H02
P@$'0EG"E]@'?KH1LP,SSOL=/A7E]WMH..SPKB-EBN6-V.ZH*H,81B<8(!RDA2'O\
P_,]@!0X-%_*DDLM'0>>P1 ;[ADP7Z:9/&LUO%X3<UMZ[L1/>#'0D@I):Y)$NWB.L
PH-F=%06_IA_M%NM10UJZ$O%#1#LR OUGO=Y?4#F&@]1E(W2"+A!E@!.6KX>2@1V0
PV.]-I7DX*S;V?K]L(>8:-_BC3.KU#=UN"Y03VI9)V412[G1J O42HFDGI6XNW6OB
P5 GLITS*SFC)T,DH*);9*_$4BH4\S(0_NN]\LZ,T# ?69>K"32><.^S*(*3_<RG 
P2-/ %&&EFRH8#]DJ5]I8K;3:'RA@-OY'526-,4<!'YI@L'SXR,N5TAVX69#^>8N-
P_*=W.U%(75%Z:ST>FLD72W6^%W\!EWC"091%G4)[Q)1KX9/A NXRO(JE[M\Z/#$^
P%A;\PY="MN\UM8#F\A*HC6( 5T1(\<"8EZ,8;8%; PSD0UJZK0!=IR*:4 ?TW+<[
P0&76$IWN?!I$;AR\&U%W)?Z=AX&TV\&02VR:Q)"7$6-5D3W=-@A$7=4XJ"%] ,_@
P/N!K=Y,O[3O2)6YV?@ZL0J3TB486V JN13)CVG!<%/]NNZNV8LEFG\IW(DFM/V\^
P"/)_(,R<.4%/G?->;;$)G1*-\4G0ASPIL4)WU6>(( G3$X&>_#R%<-A[9JK#SYQQ
P\U'H*=H7C\CD\7K$-YV]%X1U9[.><AV/?S'NL8^Y_VX ?.'H^A\%=_V&MS>#W@M(
P.P5%4!0=6L@?BI,8+ /G2>V:(RR:HWVCVWE3?6U%6K;*"W%-XBBX@" 3Y_#6S&6(
P/N]T[6%'AS"^"Z^:$MS39QR8"C/AC=]?B6\]P.7C=-6(#?=!--,&.@1J.^S_RK4%
PWD;J8):4IQ%B-8$S)!66N\:@1?;EOE0MDR$H-)KAX==:%C8]O$&L7BJE>JZJ1TE3
PADQJ(R#C,LJE_"]5S&A_>HC04';Z&30[7_)3*9_?JQ+.X]:=&P\] ?FP4'%/T;S@
POB(2I^6HF A!K*/M<%J8:_X.+)#M1CD?C[<10]L"\@Z<P*;L8;<^1S_7G1^CR9T>
P!G62S$F:Q-0B"7U17=!+;+:;5^G=H/*#Q7X"&:M1$/$916_$:/ I4O[0UH]Q>W_(
PCO*+=.RR4&X89(L(B_,,)%*(KI6HR>_H2#NTZ _I,,PRJ?*P"P:</Q .9N,6.\!L
PSYGAU$)G?JN$0&)0?JLE(-_R;&0B6]9+UHCT*&J/%\W9F9J+?7Y#4M]Z&*%[$7O@
PRR^"P!SQ$<W.>0J*2)@O(Y$4!^773@HER-J(.&VJ^H\@4:1N;N%B,,=V!._A4J1G
PR*:Y!LI0\>X_$PO8R@V+(9GUE.Y<*##J.?J*=]<>X\.OGJLC!\9C1A$G6B>WHOKJ
P7P"O5^5Q*0K?<\2$F8KS5Z!3XE&]B%J*YMFVQJ.I:)&PI=D4X3^[4NY&K7U=:Y3]
P'=FW6%@P3C'%ORT@'2[PG<CZ2@*#6=B^K3VD7/IHW<\S&Z=:[Z*0O:;<#B%D_XRX
PD\Z,(@]%>7.4NMM4PP"?'Y;5^I66VCYD4ZWL@')*JIS*@&S@S<5^:2RGLB2-\_0 
P6WS.LE)05HH5>F/<5MY9!.O !))]-._IK9*TQ:\$W'RB^B0A"_\2Y5'9<*!]P](#
P?@^O L WC^R(,B9K-;"MJZD$H$#]W2NIGDY6&EV!?5P3-SH:LE\D.X#5>X#^,C^[
PTGIT#IK.+:I)Q1S7MP+\,]8Q U.AG<MES@M,MT&,4FO)R%9B7%"GL>1J+2>UV%=*
P?[A\?9P-RT'\NX#UDD$G?6^Y^+^^(S/0KBU3(H:4(+XJ"O#?;,+"].8SM\6<J3:0
PBTO7U@O40\?*,.8I-6C=STW^E=URIJ:TN;D=5(1%N5@"0XN.H+6"%FGSAKM?H=5+
P4MDR8"TX^6_F'.-#H#G?&RP*UT<KH?Y?3)+*M4VG ]W)7&=*>]C#*22JMT/"TO5_
P8S74VI;I9?5%=X5 &-/_/G<NBKABMK6JD'187/.;0F/NBK4*9^]@^]1U[=@3WMA)
P4HWC-*Y9B]&51QZI72OW-W!15X[T(DS&V@]9*2VKONG*2I83YQMY$Q+V"D7D![KH
P6C#.^OL\.\GW!5(&?]][VW?!ZFQ0<;4W$^9&7=>L#L^O,R<I2@JA9>N,ULBBF- ;
P0:'2QQ<X> LM,'AN.A;138H=S&C^ /^1G"D)BY]!I G3B4W;>5%N,%O8F!,XD&W:
P<*S.O!F5C?^L?1!'$J8S]V*%?E\0B%""'I]NDM;MYQ@A /\R$B>,V&L!Z=AA&]=X
P92FB7-7/:R0ZT<!3\',L3>#WY _8 H:(?;# "%-8Y>,[I7>O6O"B6Z3]$O:AJ#G)
P.4[82JE/[4VR<O,CDO 0;:Q/+\6TEY(LWO[@%C8$HSU8  'G[_I5;;UG6H7V"5<5
PJ**0Z]/KN2\0)E4DL,45V'%&E/_\>R<\D^%P$3__S >"$Y3_)MB2(D-O-!^;9J8N
PQ-KH4X':/#[-@6FDJGE4Q8L)5'\[]/#)'7BUZ1:1@]5;%\&S?>1__(01>[R<4K/N
P0A=+"'&**",DA5<'*P"QLFO7&U4L!EOP@[_1+U<P-.@GX%C+&K>GE767>Y:R*N=F
P@7N';HD3 AH.8;L)&<7%GP#[*49 A8'P*^/'2"JT[B'SP57H*K:#/.7Y_)#K+(]P
P&WX*4%#RPPZ&K51ZS\B<?<MS-NO5A .Y,0G#$V$@?>LF(W'.++8*]G2HPC3!\L\,
PQN=OTJ8EJ\XDBM^BXPKWR0%9-3@C; ?8P$(3STS %R]$JF14C4BH$QU: Z/Z52\M
P1I_,HH>_._YBEY@V,7M0=!2\'S-MF]%"/DE9Q8!!5YKU.=)0ISFRN'!Z'!*6@EX;
PNXS/-"12-CH''Q-]3=GT/(8#!RO[U.3BGD/J!IVPKSRER<\L@HL_Y\MDB+%L)ZZ2
P3QOXGZM^5Y>)-9*O]IU(/LX,XB4]-W,NY@P?=MI=@Y_A_DUB['UBTIAG/65$>^9>
P GI#+MFF&2I6G9GK81-(:[Q(3N4H%0[$&3+HD$'!CO&34A&9(EF<[M7CG]G<4LL7
P[/G5$]%/MQ\LG?>N(T(M]J)3-UK'ER9%5'2'9;6Y(=8Q,W-*$VN8CRE1^R XIG&V
PHL YEPF4>T<+4HVPJ"S_O*2701JTO7K.&_2_D88)*N58)\6.:$40WOY[<"!9E6-C
PSB9F=!_Y4=$YXU:$F5<F7TX;5#EKJG327F^389,8!S\!TEK_(^A3^NQ__D/8<T/.
P,$KLZL<WU.BY\NL=,EPH7DM+ >IVLW%]>*MR301'^QW"1@E4Q"$X:G* "MTZ7 O2
PJT7T03XI<F3'_4+TSVV_NJA=EYD%4<>YD@7E_530V[?:4G^V.M.^F#7*@D&DEG",
PLCJV^PGO>SHK*GXIFKEUESM9?A_M0P]F[D_<C,I=?YRE5BR+EF<\CM650>MD9P[\
P"/<G<8<"W\:<"9!%]F=!88WDX>HR"LD&9[*_LQ+NEX0?;HZ5P$I(9H[S)7\,Q$D^
P9;=7EPVP@98\%^2OH*X(#+PTV-D^.AL:2VV=DJRJ1N9L&-HW25:")<YLYSO^Q97.
PU2:"D 9O\8ICX#FI92Y\5OSAPGE;8B)>I0'S@-=+H+&_[@%@#IZ),1IA)*]*! FI
P328VDD0FNK7$[/"J^7+J601/GK>029?W6+4G_G (C"#6M7.Y\8/C\E/-U&B_2UH9
P. F#"%_>Q^A&-S TPA--<&$S:64.]8 #L'HI_WD>0/OB 0D'<X\P1==+DW*@S4"Z
PV4$\?@U6 $AHOI)<LOR3;!+VC$!DW#C(UAB"/.AI5K\O5,,B5^ >>&!TR#)9+X0Y
P)YYX_JQT+C"'A+]05N4&RVW_8_8J4F;4_'Y (;I@59XZ4^5G@X--HDG^ZNWKO_#1
PY49SW>1AI2>[+2DJ7+KI$4R>-[=_84Q0)J^H,);3CBMOA?HX00!D& Z+1_*KSU>(
P$&GB>./)+($""2]ZN?,SWM3%BQ'<U&9*'XA92PIZ5<*P;J\@CZ-S16U!86X.BKQ+
PB4F?<=A_X[9NX\9XRX1"%*8/BQ$E"%U.L8BIVYL+%-T_IJ]&)" (5E.N#3[Q"DSV
P$\VC3NJL'*T*%CP@?.\3O.C8 $-S^T?$=[:P(->[->KJQB0Q38/^SC#X[>8 =U7]
P0EU+UZ!7E AS\V[[S/]'6"<W SZ9^:KT57?]0(A.>IV+8/THO#JR%#ETV<WDN>U6
P!/)"M&=19$EE!!]HWK=JBEXEI>FI9L'WT,8S*%V "F;-#:-,)J;>?)=1B3WCN>ZW
P0!-_%)[#X]R'/#]1KX =D5Z-31F66K,_C;KM;79PN@E$3CMAN&EK)JWQ;4/RCJ)&
PRUA;3H @7WB$?/"Z\C>1-;@[P?O6\?NF_N]IQAT$++%.=2\JTIHD6W @*\]5Y)?&
P+W/&N-"_0)@*NNIW=!*F<IX&*+% 7^1X?9GEX(SL&#AY&W>K"&3KV8H;CL\S2(J.
PVZ,,5, )U31W S=:1&"E=9D;K[OMOQIH[G$*;JWJ/,<-'>3FR0KX9D++QAX_S\1,
P@9G!.<1#>]Q*<9UVK'\[8.B._ IVU]%A"2%"O\@#,(1MHS7<=:X<'FBSLY=*/E>.
PKIX 5#0N5B:6OR?22$X2YCZP[<SFNIA2Q524)BNG$742AV()*_5T\CD6>#6(G\J]
P+":0X(=^*0E2S!$SN0L=[*L573;$S_>GHTNF3JPGT%CEW<WH%0=(W4($13: _;EF
PBIC_HY1E)R_ZJ<I6-]=&?L*H!0?02%8N%Q?E'_["E_V1G,;@V;.\^Y4>S+\ -UO<
P9Y+B!N\@#RRZ"=UJ)M ;(]<*\#L? BGOJ;#*--B7]18##4M.=J/EF)Z6%\/_BQA)
P.MVF=0_779S#N=]"H,@T<#A8^H//OTY3;1-H,C5]1!R4ZX"O&KX<)3SJ5CH,=]B#
P-57_?=/))/]*';V::!,HPKR$Z%X BM 1> [W;\'KFU%5B&/9X[S &08T1#5MW$PJ
PAP6IPP@Q%WSU.8U%QABJYAU5-: *0:7FN0 [7KW%4LNHT=P0:"G)4Y,%,,(_1H9W
P10:3,#P52(G#WZW<*\=?W-YI6L3C7038/EW84S2H0^QZI@8FEPU/U$R-93ST^<?V
P+P4>_^VA!,KEQ'[$W)'Q,4M6Y:Z .XV:4HK+ M9J3F:><Q(,!T\/U1S9!\=?:.DQ
PXS(Z]7#J1!%: P^3<V?[Z9 8R *. ,X&IPSI#1=*P&[6QTQO66G]%%EI&^?7EQ@7
P"UX^"^F?<2K)4TN&!C@IAX2&&KR[K%&S?+[>E%*G:BK-O+?Y=WF#H20OT@1_68K,
PIH%CP5E!>FK0]]GHZ "TB\ : RZ/;1WBED)H8P(!^@KLL$EH^]!HJ?:T=13@H4$<
P4/$SH(-8%J %,BK&1"O$)"MLJ)?8R[VE'0FK'[AY1I8;7KX8W2X"OWQ^$%2"B4-#
P&;>6%U"(_^I=N[I\4?O4@R2":L+ PF/<^&8VWHJ @O5F:?UMD<FK4I*^#)_FG&X]
PO\*6E@QK(@ 4PHRUY]W:=CIB$ 3A,T"L%]4U];7:GQ"_NGIN8F1!Q.%B4Y60A[_@
P4C3//L]57DD!,4KX]"P5:.A/X-4[MW-&AE%BSU(4KP<W%M1,$!TK_PIE63J8]M:V
P!<F;5/]YJW>;AE3/X8[&/6HY[/(ZFI*F!+4'H#)_8Y,)Z_0GD]<0]E.M[\/OX4E.
PHOSD^&-6-9L"4%1,VO@O#*LN79C\)Z&BI!XX%00":;7O3!#TN]M,KT4YD&L_LOXH
P.=D\W5ZQ)?*@ET"?J/"RYM&[-^S)3)ZP(6[JP[7V2%^M8$ ./%Z[YL@S$=S"K22]
P4"ZT4<LC*[]77%T(*^H0T.T?PS!C20\@!CGJ_Q7"Y=7O;I=,?9QO@&D'B>"F $QT
P/Q?&, #@4!2V"8GK0 Q\$5JDCVK%9W/V%[1X+_X6J!/1(#6(UZ#?-\RZT?.3+^4M
P@=SUAZ'V*?G9BOJ\9]#$^J)G;E,:8>9K4HSXSEIOH9#<MH5X0=5ZNZ&L'40;QK5J
PI2H\)S%X@.$G)0RF&>XBR%EYP*9I&K,UF,.7+D4,*AB<WJ1;U=XW.-ZS$"@4"$PE
P0^\C=8)UEI'I(,[^0 >'HQ+?E6&2,,)Z'K@Y:O98H69DJ;,7*E!MV+7"HFL2G2$J
P<+NWH#"K%)SV/+2)+V5)#"% '\@!A2I-T82']!DMN0B6YEH* [7F].T; [2P:?VL
P_HJ9PU/>_&D*VU%%P>B[-NP&7-(>P'3_+1^'4I<$_3G>$]W$+C+%4L3VLMWB^0>I
P\0Q!.D25L 4:13Z- +]D<' !CWP->V%)GG,+V8]%:L-"UIX8F_J6-1T[=/K]\VT<
P.Y@5!Z_MSKFU4*[VJ;!5;?9MXL@ZC6?J$E UTFOJ/-07F#WLU9:]+/TA@K"&V(%R
PN$085#-X4BT7P,5>U!<WG\C'@;(Y8@EM@<1^J?<'*>*.ERVMGG==A\R]A(0<@L#3
P!BG8.$;BY9:2,V)TEJFM._U9[DZ22TB ?"O(-]F%!*F"]*E&<!HJ'>>"QPGU,Q,M
P(Z2/>4Q^'1VL/J0:8-9,3%2\;7\SQ?QPI-Q'B6S9M&K#IS%4)!X"&U%94!&95?JP
PJWT[(4L7KE]#UIB4#&PMM\Z$06@_C9PB-BDP,M!'BJ^O:!$28[\>-O);;&O7VKOY
PH.<11,;9@X.Q$1GK/W#C1G;UVBR#I1LO/-NM[RI:!GAK8BJ\EX\,A. _E&B34GG*
P%H:G[)HZC[)Y$S$[DG68W]!TK=RIGUY1+6H=>8I*OU\2*?2'W4_AYD11X?,!04K/
PS8(CKDJ*9EI F#*'F&)( <FC'_J@<E1_)K\%]B._#".?)RO7?'9'"R9Q'=]BVS]8
P%T*9@)+&?P.<O/(C_JA]9#DE?!!B\B6Q0^-.H7M@#$^AR6R'EN?L^@7#.9='MLYV
PN^3D=["C\L?/)^7YK2TWE/54YCN*D/7=W1EH.I ^EN<B'?:Y),4M\4W=V22*&[#X
P>3@E>3)X["]6].>?[9PX3^>2ER@PZ5K\3F1N4^?0(+@6?^&',[,\1B/<FS$YC\K9
PIM;CL(1,"6E[D0:M*%Z#U:< 21=>,%VCT?@I-W<-/(OD_"S;\;C29E,&^-"KWB<R
P+>&M?&'W869JLJ=\ MF7C$]C3$$_&DKG.VW$:/NR?^^<RV@MGG)HLA?728Y/T7G\
PJFXT3@'5RK>MQ5DX>(V1HW;H9TN6Y+A1%+2I;PW#0P+5"QF8':"3!K(*N.D\HZB.
P5C+\_Q'M9.6TTJKPL4:-59%;#P.GZ\F_.!,:04CG&GL"+%?(H74N02;$TK-_5UFG
PXV3@6T!SRYUD +PLBD)@*NSOKP[E')EWHRX>D F\=M?R.EKYG$2][K:\?3W.+:H3
P+T&.X3A5^LNY)IIA*DKYBR< F::ZA(6$^#K%8UO1+3,%]YX. ,40,231=63+C/7#
P#/_@"NU-,*\2(&':3\3K=:K,; DRQ[0$>,2#X=SF=WVDAFCXG/IS4_C1@F=R\895
P33/;*3*>#/_GI=:JBP=>^C[J"0[8P^*\1:F'P>47OO7.7.)D*7JBT?F2VQN-TBSS
PJLK!U)&PNWD!JUD;8TL+-8O7+M9MI)R91TF)*Y^^;*.U1C93*5H84UL^9-\7+:W@
P7_PA5W.YHX0B.NT[K@=MWR.CEP]B.05XT:TMQ.WJM:@:L>05.BDJ+D:MO).#W-<P
P^6UKE%56ER]-WP!!2A;Z0815,R(\@]M]UOT7IN<=9>%(SN3S]78)YJVW>A/]+JGI
P>=PBF!NKW()?1H%HIP-7;5Y39B<P&"9E)KI-]<M>HP.-HZ;LOZ5_(:R,U,<-O]W!
P!Y9O %HS( 7VU>9-<;S/2T*UY0$1%6KV^Z\=&^H6QJY(0'K):'M1FJRRV!F&SH=4
P'?]_DBE_^$_G:0-5LC>Y/4;$V'3H7(&UB>:KXA*,Z2P<VF5>3P.\\!U'>.Q0=6Z?
PK73,[JXJO0>7,'[(TCG?V1KE=8.H@Z$0ZXZ(,ZL,3T\UV:$=2_=).=ZVM_3MH0M;
PLMD@@B8;8M22P&W#OD6F)?4Q#TE&"7I ^6TNUCP!9V;[KA@%V_ K<D:$&"'(! 91
PR@X1&Q?E7\N!:'DN<1*"]*;(0#^4N./6S#A8EE; +N1)Z$"51.2=QT7/'9^89_"4
POD3_S+Z? <@M#FFU,0EG=.5NF45?H>;8>SRT"[AWZ8F(8@?N*BE:Q_*/9VW7OX '
P8;)V=2!ELJP$T>#\7>5"1W'>ARV$HN*FQ$9M[HC:/7Q7+D(GX1G="AL;%R_/Y2]%
P<+<F1_JFWLCKGS<J44NS(:<:$N,&K\S9T2A&-L3T8:1L@,G2D$]PJ7TO,%SI6:]@
P=M@R86&O,3N+CX6TGA58$F:8=KV0@1\R<=H]N>@8L[?%\#3J%S/%HWB8^%^!P0@2
P4(]X9H,:#B-^2[/46[=4H,>FWL]/'42N,T'^5]E),2SBH8-.W"F;UK7W&([4W#B-
P&S!1U2F:RZ^I&*P !&AM HQB!\03J1C7L1HU>*$BV&+IO [+CDXZ S$@D^\A/@H;
P/H9*D1GO@_Z(PH4/?7O7\Y?'E**L0A-4KB9ZT3&H(.Q>]2]8=&W-UA>J?F*_TWP:
PF[.5L"_D6CE9K$/5SAA>_O)F.^>.VT#L7&XT[/HMF)L#>+4[*=')7''^DQ"2E$^*
P."X9,<;T@>6N6>Z][6?JS[#V@0?[1K>ZM!"$5Y;:F!!I(-N7);F0"8;@\48+:SBS
P^6X5H/!(Z 2QE5.9N5R/ 8N+ ?TI?4Q$MIA3 2/*F83AJGMA9SBG1&\2.+W4]'/4
PV,$Q=QDMUK@LGQF3?99T;0O]%&@0&=FF>MP:PQ@<'&.1 U+60C'X6S#L31<5:E*1
P_Z1$HR<:\,QG.&DKQ3HPP0B[+ASF-FFU7^SI*5F<ZJFTP5=%L]U:'DY/0\9@'_Z4
P9FR:%H-J6;KQBV:)AD95\ZHU?,?G.84JMJ *O[( 44^#,PY[>8L/0/:QK^E"%J_8
P'N\Z@7N-D E>30N5?WQ1D!2C*";<L0,EXY 3K\\O%>(4!3TA2L]X@D5$22T3R_3/
P^LTM#5^QC1SF"\(QF<&E-V]W#D"E[E2+&,5)6BH$JZ;;C$;22UU@<*<6DF[B9'Q0
PI:.NI?^ ]>7^<=PELG+&!X>9F%:N7KT#2!+M[:,5?K?F8EI7[Q1)3?P_I(Z>/S/4
P-J<)L&#[M 6=6]W5]X_FRII0<K):\M;([.I^JV0P<)D' NS1[5:DJZ>59'8.# K4
PTOZ[]FM&AZWZ_B>C.(G(CQHA$TLUOM0+_XG@)5'$-WIA26+[%V#)#.!.>8D27##Q
P?DM]]M57(O&*C9J"E:B@%4V(>CD9DG*+NSF!N=ZBSL7:-V;OHY:V7 R ) QE\9",
P#WBMDQ0GL9^A9<+&+&)\AKN7RZE2[2CH=EI:L><DV'Q4#Q/_;IT4B]-W%FV/8W8+
P%UBP:Z:.M1<@$$ %P,C^#7P]^N,R8C(G8,@77%C]4CG0A]6,@H?BDHW[2ZV\7C:T
PSWG5F#I90$%9V+W%%VR&'4,ITR4*B8]O\D)W7:V4OG[OE^0%5HE+8S>I3K)Z05F2
PKH!FHU+_F,AY->DC#;R5,N4;):1&&&!2R\S.K06!$H7R?&&01'1],2Y1EPW04KCE
P8=$5\O)G^PX)OB#XK8.B^:N&T+7JO6&F#D&C^\(!%0>W[0)%M=<8&$Q/M4^X>7YE
P7*YTW8)>!6F+Y03]3LE@6C5M/:^<L<EYZHG;W*ZMB+V7=12]&3?0W?U)1?TN$<:"
P@^<M3]6VT>&HDL09'!\JMSX$%BE/AL^H;]PLKU@>"DR:4JYBMLXK?PWJZBY*.M1P
PV9U9&B$S4?P6PJ<U Y+<3]K[B>6];C*9Z3X#+S5@J**T3T%EV)VV/_5MP_SY\63]
P&X1I"D:\0MNQBQ_UZ;V77T\,S_@69W%3\YU4(\1A=&U68^K;9;:J,$R&A6X'GN0C
PG=AJ@C1+R!Z]M\#O80ELHAY<P*JY !!%,YE5Q4G6UWUI2XBF;6VE<O., @9AX+6$
P1LIH85S&FM\NEZ%,EV;9#I[N=3(T*2^C5?\NXGI-PMT *%TZ<7*HK^9[KQ8T-L:0
PX\>?R7C@F8.&/1\'#Y_ED21/1#,D@=_)KDQ0^KI4?/S?L9G]L)/_P8@!#E5;TI9\
P>N1RB%5Y:^O*X?]1B [W9,\,G_QA*$LYD>EK93[3(1.%$\OP2)_4_A ,K+);:M9G
P[SM1P?+_3R?C(>Z<NP81^T+B:=?([9D &G9S-[^9GN#/[$Y*FA%$_!U<Y<4TST[#
P79[5"TRL$],7NWP3AWL,0Q:-)J=<EP0S>LHN@TA$6&8#5^>[TM8,?Z2$Z5&$K25I
P],_!RS5Y7V@PV/;?5^5PTCL.E_8I8_:CXK;B'&,ZM#<.'&CV6@TL"=*U=GQLG[@&
PB&#[W=5K4KY/:'W O;>3Z2^.S[F>YMSBUNQ-::C'$GU:]1AB"RX-Q^SV!4W$,ZIG
PRNL3MB_#;JB\F6'3).Z1?C&($2%.QXN[US4]/*3:?1VKX H+EKHLDN&<FMDG[8V=
PDK],!(9%F^62*V:-PKT@A)*Q7N_9%97GM4M#9WL.[',9"X7'>$90 6NA3*=IX/:Q
P]5;YC@MX B'UC9DG)68?RA"MZY#:DC2LVPA.C,*&>B+?P;6!2:X](:UIIW?4]D7]
PU) &F82OVHM&3(^>0*%LDTN9IZX1$.4)*00W88_B/GQ+V@-=CGT&6%3BB;:9[N+Y
P<!8_HINY]R/4<N4UK<12"ON_&)//L+?DW<ZC5LI<BSZ"41LB#S3%]UJ=[E1T88<@
PF-88/_X\UE Q0$'R- JRTEE"*9!^U\0,0$-!H=<I)SQ[?W.%1Z1Z#&JBT+6UB!3&
P!:8 >5V6I\"WG^5]PD:C9GO.Y%#]Y"Y=E$>QM[IAI\2],Z$]P]+0=QHE4C1^#?TO
P!DW^A-YHH6MS,H,68)"V5B*# @"44Q8X/'3ID<:I0?A?BL", *6 @8OADL7*CGZ7
PT )<TI3(3C^L3Z0"?;5$:6U!+A920RY?UES=HW4=S_3,PN[=FDZ5BI;;^@99P.L5
PF4QK7L*:( :R"71N%X&2*XFF 3@X_M)E]2&R;XQF-S_0S +<['D+$E&E<;?Q[_8A
PUCTKQU.M-&_+(8S4DN$ZM"0X/K#"B6O7S*#>W%X\@)I4U?HWA.4=QS'W747# X'_
P<=5$MXBI2]-/%.03?=C_.PA6OR41Z"1[(WO^::B[D+:8#QYY8U0Y2$V=T[_91W!Y
P0&-6;?GK;@*JF+/R)N@OP#1-S_UUS@. .&#>>C8_\R=.B">7W!2V4;:UJVX%*( N
P*B[&\6)A"3TJ[Y?/8%45K^FAN\D)+BZTBE%$-X.WA=6<-FVTEMY[<\G=E5>%E5@/
PJ!IJ.^H,YS%JS,[H,JM=&3/_<8H.BZVV?M05V:LZE&LD')DFN.T*Q'MS6H:%]:!?
P7-* SE[(<;@V+9T 9?KDCZ U&,9_$2*I;+C-R;RW?9&F]);[_R=[/E'3KZJS.L6Q
P3$H5PE@-M@-V1Z5,ID]=X[ZJ5QCQ$]S;JXA@9WIL0+-7WHMD0X ;9/&=;FD47U,V
PX0%T(2!S@L !60V4&/?#<?7QZ3I,G!.JX:L0L^^<ZH" +8SI/Z1'3M6DMB!ASKG@
P::MVJ66/1<H*K+,-E<$J]0R_Q1KC+&2I TLY8Y,SRJTUS0,+:@C<<)YF+\F)W3JV
PK,$QO3E'3<+*S4\Y&154D+[P2/C%C*\T>!7LZ15UC!/'#,8Y+Y:D,O0MZF%S26" 
PTQ'TYB7AQEDJSMAP<G7QLQ/ /RUXPN"O6:G_2MIVM^/(ZT$V?H L1R9NO]XL%9$5
PI1@RJ!M=:T]":R&'0/ND87LOE=F[>:A+V9Y"U4"B1R TO"%N%1W=<\#'54U;;LWS
P9NM+XKU1;J*#4B(UX7\D1CB5$*K8D> ;9<D=*!XL^F?,Q?"/R!!Y*]WLW'40/4(*
P 1G1^\V"38?)&'-$A&QE$O/_Y"<0. ?T!EA(UR_1,"XE+=2FQA-^B%K&JV9#>ZZB
PZI8CT>O%!XES'JKG;3G*OS4Q;O$1#T IJYFNR"K@ELQY5PL@=K*N)5 K/.W06I/N
PXH0V$+,CDKR/+>+W'K8%<J?\X^7M;]HT5?^"M.;8U1VX:(]T^ HW;7U^6M<ZM/(W
PQ*YD;0F,N^H&"<>DM.N=%K)FAEZ!(=XWS6U+II6,)XL]HSHP)*W-PSHJ/=I_&0ED
P;OXC(?$Z8GA,P\^N>K+,B*@/\P,=E4]G5IC]MPNTG/?<A';#=Q<XE-ELNCEXS^3G
P P!7RDG;-$&TMB<Z>/==W#VD,('O\ 0N]=E!B58<)2CRLT8K/ Y3\\_Z0SS*-C0A
PC1HU#HV/#H< RK[:V-ZTRR-WJXIMB<YSD;6-P'</?!F-\ DD<]3@VC0:S5X"+(+?
P.1VOX^=-20/8P4??7OR\Y$WX^GIZT+=P%>)^GMA;AV8@JTML(#P"(&KJXRDL3D6R
P78)U_5)W,FC3ME+M&<!+?M*7:\N,Z9(DTV916>,\;>C*TPI>4[DZ<?5?.K[6D1 &
P=;CN\N/YPN.?28KS$N'02J@?Y5] 6!A9S*0*7-=*NA"SH+'SR-[ELP75K )795!?
PL?7(X"Y.&OF-$=2Y5%JBXKD?[P B3=_81OXVSR66W'"0T<B AN9IR"39"95HO"^)
P0,'K7[W'[J8-GD>RTXH=.T6B.G)AJ%FJS)8,(/@Y:!@QO>3UP :%@*B9!82B1>@H
PMC/M="&>6M0$5RSOX^2W>"2U$FNR MG&4U_M>O:2ML?P:-6M=U!,.)&>=K<BLDK(
P)OME"B)8.RY(*&[E^\C86F*MM]R-:(JX3H*OV'CBGW"IPZ)/P\*N8">U--)"'*YB
P$VR&WN"Z_<"EZPZ=EQSWYO-(_6P>YK*H.A9\9RB-]@Q3_!F!'%Z-3)1;U+7^#/R]
P)H<C(T;]O($8V@>D*[ND*R^FQ#!G3I_]J76BK@OS6%U%.ZAQ4 Y'.[!W"H 4B(ND
P2 %%V=ZGR>!O/F'41E14.#Q+'?+O5[<9W?OF5V5AEM9J8VFF&B$Y_H;!Q0\-GN*F
PI@.FPI17>E.C?B.1:5@%DL72(1K,V_@&H,YOD2OJ'/V3=FKHX%VQ(-U13)'VI%0\
P_B1*5RE]7;H<F(S5O"+?JU:4&L%>QV,>@_%_JW)YC5!UBMIYOYK4R^L^Y6%_HQHO
PVF)*ZY--^J(EC3=<#WBL(,.7ABF:M),LTT'S MU3K3^J)?M: ''WSBN<ND$D6E-R
P1J:""V[!S(V:F&0WWZ -!UM'= "0QRS6-_0UX5RWXF3"MB&+7DW ,#=5J8C_]0X3
P%\FB3S2.)3\'AV7:;SDVIB/UOEM)<.$S#EG#)WF8L+-M\5-WCJ&/!HC+A4L'*.[2
PYV!-/B6AX36Z8NBYCI$-5#9DE?5#+/%Y][8N?!0G_DVGDCJZJ!C"%UTAM?X.UE)C
PU;JV@VBVD*1:*II*2= MB[Y:WP8>-WEHG#X (-DEG?8*698GOO\-&*U6SFMZ:1V#
P+*S[?[VV9*956(H<)?LV(7&/\=.FLP^5J4IN>$KK'AE@52-I!&Q:_#V[!?F+>7]1
P/'V;21 B=XAT]F#&3*'C_C(K&E=.8W&H*U+8^_?H([Y/)=VI,MUY9PL25=+L@P R
P*Y!;O96<\="C?"@(X.S.Z=ZI$3%8P.PC.:/4^7I$ ,_LK^C#?$!Y4[U^/?T%-8W7
P=S$ZNYYULDYM:;O-)!4#-8^I0E3$RF,^[+@X-WA[9">M I+M/4@EK*&E] 'L_L4!
P5&Q*);Y(5AZS%KP=\6)2 D!+L;1>6VMU.X:#TY1'+]BH%'@1]#WZ,GLORZX^K)>\
PIO";3Y[":X,N2HZEN8N^339JG<>AJ_N0^-38$4K0R8@9)=&UN5<1SV,IGX#\P1G?
PA&2[U3I&+V+4H-NDL^JXWG:@4U_[A);3(/-V=X^,29"L9I]38!T5P'=?;[,=UA V
PZWD8S4DAYWG&9C(I1,RC_GQ?QWW-X,@-2+R-E.W$2 *!I- "-"T!:0D?T*#$$"!4
PTE=DF9A;@L_2H023]:L^TZV;A,F(0SSGW+_0&CX^<,W#85KS8/6X"O#?2+)WV'4[
PJ29F0"T#YS7P6Q(=SCYYL) +?YS8QJE][HW-'^QP=/5&_(6C]MU3*')W#1I+I*\X
PD'9HU5T>< RH\5SK=-AA6KTP9K9C$_64[WOVER&:L#E?PI@0BKY!&Z_,#ND]HYQ8
PG;5G%9"/I]?W\E#OPTFDUU#E2Q;HE$E>*\WAAQY_LPM8&&"VE7RMDT_!> )%(;E!
P5#%(&/&7P2;H+EQ6W&+P:QFW-,!(/EWQR._S QJ><.=ZRX:$FL- ,AYLA@7U_P::
P,#:S#'AB;+*0Z]U@0/>0 "-;QF>1E8=O_KP'5AV-Z8>LQAXYTU38GO]V30M<<H,8
P<M'6]_<CW4L0W:GP@*\(RQ,RB?GZ1:V=57#BOUBLOEU,EG\'J&5$2"8LPD>+0K+$
P*_]1!3$'69%I/E9XBIJZ#$)1!LS;PIP&U$/<2>0/?F@8EN&,W=PH%W/BLVI@$%;0
P=B E/8! F$1A'#(*Q*WZ-8<\M'P($(4^L]/^*@NB:"DFTL*.Q[5K)?V+5%F:]VN1
P+_5=TEP8'! Z5?VB^I)^O2GL$ ]W5N"$E^3DW_$"]3AOL!C#(!P\):K*PI#5M[(>
PSL#QC<?Y9=;A"2C\F^CV/ I5$"? M5^6+4YP(8FSAR*P4?5AK45-\D-.E[!),%1Q
P(%R(XKRD.97O7]G^,WD*C%$JWK7:VOY%,9YSP8!/$XRL-SAYZ;+L3YA-[,F$R,\;
PW0$]Z=V^11@!RK?TM2U<7:*?SJ<2QEVVG[ZDI-;X>+$.X3*6D6#XFK2>G,9J>#E=
P;^>ZI48T0H9MBLK5;]RB9>H[V#B(L^^=3=!MS$X0E]Y$ 5CW+!C,+_;ZKKW9C_Q"
P<ZG+XO. M2HX@_;+F2Z+YR(..P\KSE4$7!Y'B.7LL3V/5,52)BIL?JH>O\]A=>1@
P5 !+AUK6/DPU0E):Q3805*@$F:U&(#'YJ!1.7C?TLRK<R]O&A,;NLCF^2H5JO$K2
P/*4?H@2T.%=:3&=>Z3@((KJU4S*8+Z%3A0%]:H-,_[*@&;#W'^"%#ZRUL;5:,^I 
P%O?RD W1BW "GG+A!8LQ2Q@SKPV$LP[H[\'OYFQT+X=IAU!XZ8V0#/8[.:[_,]OE
PYM1<OX], 6=5>H92\5 =Y\[W$/#L6)E]4ZSL88=-)<E+D2/YK!B!F"W0+##P)DBT
P@NSR<M0_EJWBZQBW0O'R0FPHKY&TVB][3I"<J[ONU)9IRM<_+F&ELZ&#X@5 -(T6
PY#;@+($!\YZ[4LS,T]O"J9(6NXV%MEF4+#Q</&@H\<K#-=+S6/IH'/X@H#_758&)
PGDC)ML%C).,/QGARZ>+IX"4!:N1%]$(/[5KG4N]7-DYT?):&CX([$$Q/;V O8B5!
PMO!N>&T<M/U__?G$*.[$GOY4E0'E6=MS#!3B&>;#$Y5*8$XD\^6&?X)96HLF' N#
PQ'\T'N+%'9]\>HR?ETM*-N*I/DL@^!E@T(2VI%TS"V! W[Y0TIY]#/T%^5!2&FB'
P1\;N!H8]  ^_OZLG^6V'%AR@)DR6@4*8]IR38E#.C.^JWMSR'<00D%[RSHQYPF%!
P:8H-,-Y>2M^C8;]_5R6A_6HWHT %=<U-;,8@/TI43:^0\FUU%)+ GQ7M'U9?--4R
PN"9LJ;E>4C7?XL0S<-*;O/B<,I0(S7,K*B--EC"Z%&N;X>G?4HUC-I8$O805YM=D
PKMX#,]293$%H\('N'?RXIPD<&J*2Q=8UZ9<N9*X)D]T<UR_?P'BM@#8V0D!()(2$
P_K*!+$5U#SV02V(C:NT*$]\8!G=3!^,X#:S>IM919VNC[9K*] M'@^VPB)LXO/F0
PM(W'UJ8ZJBZ?=_%G;>*\DJ^KD]5?F$V+)FV?K[LG!9+KUXMOP_T&"J+NHJXJ60-!
P*,! +L%?L7;BS89=TM[D2Z5;3@1;AK49G/^@&GPX@>K4)6]0-*O44+^PB@.=**AQ
P)^J*=T4%<<6!$Z#8NB?)3I7K_A@X%#X72MRN=_,'@+N1R9$(U1R&BA&<>2S72S69
P[7=S9I)0(&E,,VV4D)2.5,GYS$12?18S'\5^'[.XSW!]%:*FO&PT=Q7JML703+F#
P2U]".Z8*-WM%=I76-B]&/_+=JF/!_M7WRX,\\R2B\&6R+6YU?>V=(OMFOZQ\)P<L
P-6@NPW->8NHT>>1LQ"S$.WIRE(.I]<OQ>9]POWC+]^'=V.@8%ED)>L0&;ML8F!Z%
P1!>8G_EQ6T.?WL M/\M,)EX"$)/9E/!C[2/# 1O<1J<TJJ[8$4'"(&F]+YO'$YT 
P9X<)[69#\LK1\9W^"E5/>*MS( Z>&*0"H7KO;D T_OO^7^Y16N*ZFIUFYORYA5#)
PX^ 59H#72?11J]!:,*'+\H5=M%SFZ6&UX&K"4<H& #.N\HY:.P)R0>C+)KBR&M$7
P/K-E>JHQO(Z\SU\&S!2N$GB#XJ_>K^,#O!?VE=6U@_.Q0?_%O'C3O0*_72/":ID.
P?")N5MH0. V"X$+RY19X3+NE_.RQ;4HLW#@<5\N;<!FI?=VK^03;-O_6^D%9)@8"
P>[$BR'K?=%YM:D/=14?W3T^ Q+ ="2=/NB8W43VXU<_W2AO]%0Q+XKI?#@<Z.[5B
P$RD0# L9Y=_DPHHABD/C/@2&&O?/+S.S-5(EYES=XS7ZW [-8]Z?)TY8:30 BNO2
PI^5*T_MVW8? VD\ %-7^@2D+E)_WQ&I25%JN>VDTH)7(9E+10#IXECM_%^3;RP^?
PXL<#!Y.__9B/Q-!3Q%.9L1>=\[OW;)J5^N.PS>17V_-.'\%Q&[5ZG$DODL+P5(]<
PL#D]6'%(7 $\ <J-:9"N/5<CK-#'A?Z]_3?=%IN@ 4*))X;"<H?[/?=BIWH@9@A$
P8 (J8?3<VS\6LA,_P25[BE+/3HO1N+1GQ<;,7JC=6Y0H693E.63Q9;#> '_.(28U
P_I(\1TV#S\Y6%V9+A5?0X$EPL.1-D WT_L1EFNJV+[@4M8F6>6%$HQIC4QGU47H+
PZ07H8NQ)X21%M_$RVKVB2Y_Z> @^*^:F7'7%7'H4R93QC\41TE[L.>;-3T^7"R!V
P)RI,R4ZWX_ENCX;[@WL(=H][LBMU1;(C;0W[TDV">H&._:N_A+I **RLUHW55LC1
PQ5,>/OLN2;P]Y$<,1?&SV(0^6 Q=8*,I=-.M26>8-#D[@Q,[/3U=GI0\(RP/]PJU
PMFV+9 $;'?3<AAAW=0!!'Z/$)ZG3401_Q>4*^_C%N06K$>G+SE@2IZ>7FB;%;(BP
P<OUC_X=W70^R+[&J%+B_RX+1ZD3I=J4F[8PD6['J5P(.&_,K6*%XL_3JHUV;&3<Z
P%\OJ&TW0#?9!D(07O1-%XB=%]^ ?-Z,Y]*4F$FG'-<D%YP0TQ#F,\)CM[5N-LW(I
P8I6'R(ZI'"43Y:#J;E7!8?X%RD?K&QCCO9]3>\5:K,517Y"!/YY[W."7MMT^3J#I
P^. JN-%9\%GX78YE*DK(P^..L5)30TP#T @(+RP+F1%6>;YPQNK.GUC-;J(]- O/
P<_AR"5]$R8U'(]51-QI@GOT'Z@RP%E'Y&3$]V&9Z<C\F00LUV-#NP&<X<4V^G]Z8
P3?)S&FUW 5>]=(ZP6@=*E*ERLI"5[3PAEGV&2G]N&GX4<YQ8AT9>:4VS2HS%17I;
PEW(MJ.5!E9YPL_C$4T4V*)OX[N*"*TQ>,?2+O*F829\#)1#^"]*5@9$=F$N=&ALY
P.NXI.Y#VLGR;!(8)<#H1XA1Y0O;=_>K(<.I#IEP=+FK0(SV\Y&U2F=YUZREAM=X8
P;71..@<&M>H3"3]^=UU;6[#>2X^IK>R @CJNI:!G78Y+?Q&8C-NF>YU?;[>_&$><
P2I*#WP U'_<[[?J/ER1:K>R??:<Y#'4]<I^P<2UU-)F.C!GB\$S0I)VL19I(\8_$
PC+4>FNM4B906]L81)QHRLIGCMLZN;/,]7[+$V&9UTYWAEX%3.BE&OYC4PS+G29O9
PL$'&F- FF&;C\7RUB?[AH'@O:@!I!&V:7+S@",N/8!LS%N.0TA:)<XWRXBIJSWU?
PCEP\.G+2>X'3?9>DCS'"E+R*"[4P/XU@=$BI22@>^!>8T/U)7@O .D)S_[+NX)62
P7)4C\_=$=3K-ZH-:-+$90?1"P$7@OW2]K8P:H'"Y5WD7L3G\2EKN[JE2$=["SN31
P,L6)J=L9J<?E=K"R89Q-/8,<X?.L@?C-XW94F_^Y'5UZ+E'HH4U;T)#3<$W%[?H/
P%H;O7K\(S1(4Y?:"@(4C[C6]2)58F*JF*5]2$."_.;/"9/[:?E5S<Z,)%X#E&&9B
PE+.7T77?^[YK*0NS:*C:4?&9?@%2U4_%8O$'2XJQ^8^QK$NRDQ4.@;0,Y[,Z=;Z7
P7MZ*SX@6& V2OF<M1_[R4?&_\F=$!>ZU0L7;GC$6YR&33B^$S#<G?_:.3(,>P%D=
P+B4/T#,"[B:IWGURS)W#LKH#+6GHLDR8T(H%(X%?, I]I(("%?0!EK0]#L1Q_,%I
P4CUOP"YIV('1]!0UP#0!"&GD%3[\B]\.';H/C,NC=\@4(283!&B3L4ZT(#5!!O''
P;]E&,V0>UKO^.ZS=)"2,NG/7BR2#=;>A\.$1O(XS#>.)5H0HD([X:7ANC6!FL%4[
P(0]:R=F9MHQ8:Z8FR/I/N<$/]V4A_^"U:CRW)S*2L.NI9<XY(N>2]GTSVWWI%/$$
P:_A+GR-7&K0J=-^_S!=S$]/@8'#P8L2-+W23]QQ]WC(\+@9$R1&-2;O0CV/KL_:M
PU1S?X7LD?F(F'D\TO%&ELR(V(8]9S_A6^(QX!,FJQP:5LA_V=(JHG6-%F4!]H+8P
PHSV+$TV5<L<ER+<2W A<^(&[4 XXT>.YM_#2>:03S;R"'E<>0);@2IL^&#^S&UW!
PB835>U=.3)\99T;%^RZDHUYXT?ZL0A(A^VSLM4O9XBK+R;&LGHD*KCU.ZXG2U&1"
P_ 0&>=3%RAU%^ C@':.0H^<$J>JP?K4?V?684XFF&RV@K&XU,O>E\ERZ6*SPX'C1
PNVKD"*<QX3*2.CLGU%'[)M_L*OD\_?.-NF_V@N97]M*1"?KRFI&/5<B>#(:.M Y=
P3T[4R=^O%IO&O)/Z4\'LP!IID_G7[:W<MP[7Q5\D2?J@:>!7=03+<"X;_YQI&K.)
P5C.U$J.AE]8LD_Y\_@B5GV$U/W[8;S&- Z $MO?_]UC[I\/Z4 N,E'"T=K:NI^B!
P!MFP.&:[>2D[P2<?9JIEZRM![U3,L\X*,C #AW[V/.L/&%39P9L2Z!U1\PTH5 &+
P!:;V9WTQP]X+\*%FE.7?KXEKQIJR&'P]_W5".U<L10:J"\!+3[PA<%#(*W]>R7UT
PB=7M0E0QNY0"K%? %[_^;$[S53)6/\KYFA$L&T1B80_Z_ZN@_B>5R)YPRR./T^'Y
P0Y:,'Y;F!J5AROYX%5]2)C_\#FGRQ3@.+0.#D"5WH*35,,'G^#E!AR?T46="9T8(
PAR+)8D6_Z_\6&,GA8?EUVQ#-,JZ#'BPP  O"Z;<T^DC^[DOQ>=?&!7EG)<UT]]D@
PFX-[[_'#"H$D#'1OJY*;$'K0XON;-;&Y;$KBF';O++<B_<V=MP%AR?M)O$.(S)RQ
P$L^HCH0R^T_=>]_8('J-,L:[CT18#^M4LG@^0G-?(%.EJ8?3/[F%?P_*]][^5UC[
P\/^.^+S>3 3X=ZZQ1=&G/.P=G!I.ICT5"+U?LKG&"34G*8$,L!M*C4%0C0E\!\75
P ZGI,Q%K'KCN!Y*N4YB-N*P47X,< #S+9%UZ[?22;CCA.<K$6HEI%CL&;*.\>Z<2
P*T$O5Y/@TRRY";V60"(C#0/KCSD\(V8$T+.AKYDS+\=&2>K\E?\ /0#+@'T<9V.T
P9UI>7@X&KF39N1(^>T%-I)8@8S/ B;S1UU<'5NU-3PY-$W&'KR""*;D:.3NPT8X\
P1&8N$PK[I)+EPNJX+[5FV;>@-[SJ#_XB<4$Y-YF7P>Z$Z\9_-^>NF"/Q IX^YG2&
PRZV0$T8V7R\LMG#T%!>([&S0Q+I19Y=:W&*L@L')).0VV7!@5=U^XG!1)OSUWX >
P4Z<+,R;NP!KWNL'+$V)WIXE8TCF1:<S+>C_Z47"C4PY84X=7!:+<\Z2IRSDNB)]3
P%+KI$NFBR(3($AF!7T4MV[__$Q .CP-XJO87CWU_?47G .!\[*&(1F]9C(\!M"Y]
P].$QWS*/.5KX71[KUPDU*'*BR(HE#MSI>U5D!0OB_L-#I8R29D Z7D.EQ*5N>F0O
PSW!'9>6UP=[/R6"Q/%%[-Q-U%6?:F4Q4-(Q?>S_:87J"<.J(E!;S(E;I1L;LI&TD
P%TRLU,XCB:5HM??K]WC;8E>:+.AGL2CN1,N086:[#'.;D7_R\7* #]X?%X'&@_ -
P\8P/B+.=P0(%V:FHCR>HD:"9^N[%RD>4[0\EBM3.)KLQL:D LYZP][JWZ107)1/N
PFN45@ &<+@O+,X6W#T.G^K8_B=$Z9^)1M3KI--NQW0V .&S*PT;YI G=#9#D*5SY
PS'T]SH'M=$!T# /AGPKKQ?G34RGXM6.6;.Z\O_*HS'/,QIV"=V#T,L;TSNR9H4F\
P+5$D+GK.:W2DX>%;*_^ADNZK*]ZGR=Y.8C1'*$BS"7Y=FE/V3B:_7<S@=_TPEL#%
P./H%0-R2&$CH5S]V35Z)PZ,W; 5I)&*]R;Q:R+"PFK)1*-$S[_50(&\_S'TL7_%@
P=/3"%INV22FKLJ(R-TDNE#<E6C'\[_'L..TA"#0RUXJ'X8^4P'JU4C@KM(T M8"2
P*YM"EYC!XF#[F1QA^Q:J>@VI0^VUY94HOH:FV3:9JLB:"BW)-1'#.[0SUC&P\&?T
P\$C_G??2^+W\)FDI9H&M#75X2-H'+.!N:,N(GGT6\&R/76KGU0[>:LMPQ_0!@ 7Z
PI>,G^,\Y=(T5,2?>:[J.D?=5-OFZ8>_Z O,9^)O@T^?>F+1,TDYCBXH')67@[CY;
P%)ZWZSP@:K>4WP1S>*7<G"X><7-7L&X18#AM=]"91ZQM^(\/&/F[?BRYUV,%MPFK
P_(C@2:-&H/Z\SPC,;#%IN:RNF^2FI!IF/<5H;X:M$!D)G"9).'8 +/C(B!:=S/G@
PXS?N)T0\/7_[X,?XWB8)7\8U;P[\V'2MO*) :2VMA[[/O>BK2K6/ACI0V_$Q_T+J
P\0)7N;/U"&RX&NO[A"]A1SK\G=3C1K[%\+X])$=IOO-$0"UDS&]CB')9!0N;&K8\
PY$*5#?X&91F35 ;"$2_26AL)\XYVQ$(>W37,1=1YLRJSUC+I6.&+!550TI4HF9F:
PB#6[EJVE3K!CH5*K[5)'#D%:+5F,?MJB^OX )18+Q*#)/$\!@^EOT%J<;<XZ723;
P!]6C[>1<^#52E-LY2.<T^-,9*)O6ZQ VOU;DD3 Z>V?U:X)0]%5'Q=PF_<,@-BGO
PR=" '$Q%.2.61XL*S#8\LI/P(-*HLNQJ^]ET.2ZN-HUM\.04Q9-E_NM=<ET6+1%2
P+[.R9]BB77@%,!0W4R =9 @S2I>#- T_IIXLY*'J<9'^E8I?=7AV'_V98J<^<K3[
P'F5M>M>/-FQGAM'X/!G&0AFA_V*P Y,53BXFUE4Z?+:+FRV+K"HE]V^XF*A^942I
P>\)VT&[LQ KWK[@_*8'ZR4J>ADJQ?(Y8O(^E2G+F@_WO9$7]E=S5'Z+$8JE0 HI*
P,_\P="I;O:3\X)9;+!T9$MR&+Z042N1)NK$7EIL"WKE.KDF-V$\FQ*._C3]J+Y__
P$V\6Z18C -^>[[W($+XKN4M 3(!N!-1"NXP7_CV&^)O-#.51?OPQ'Z^5I'A!=1$=
P,@$Y8"@EEWT>%JI<AF_RS!/ZSI-/5=U*\@>/,H00:47@-HVN17!M#$G10"'&Y-&X
PH(%*1V?CZ2F#WX;8]XDFK!I1Y,1+I;G('T@5Q;*-EX=<7TIEP\-*?=.3I %12=S'
PZO];3*<V!0<71SM;NX)!LH]G)>*Y<;Z],DE[7N1"T^S_4X G\Z$+HM"V(QMW1##<
P[@=+5E!Q:Y\@!T?.2 [@\:#YTP$^]Q7-9/7R(JY$:<;*X<H"%7;I$(4-G# V8K]<
P_]7L_X3^#5IKD1>T^!R3Q[''FXBO?\7X-\;+_0IZ%,'I!WF&LP1SU->O#+,QM$9Z
PH@(P8-Z3W@$[;=P5KSG<^W W(J4U>M@R(XZM6KW2?T/-&WB492ME#!@B!68S)'M3
PKI.0@H*RB_\Q#I-JL;&>LI&/M@XLUO<GIN;T5W4TC:DZ^,GWJ>NP0W")R"+19T8E
PJ_ =03+Q&+1^L>'R #RIV'T1$D>VN17<E>J9&O-Q943FC+R$PS9<J;CWNU0P+U G
PX9?=FNPO^$;9(T8P:&XK*&2W)N?FVRM6"'PV_KNKO(F%6\KQQRYTT%#_.SUTQBP$
PN=6<C\@U"_=1Q><P/.MWH-"^DD9'=)BAVEG&#92$**,U(K\//T#?=&X#U'X@I9AQ
P15.R>2;'F 9*00:'%EI6MN%JK;WF62#2KBQ80MGDWKDH>!7>(C[5PJ@"HS?A=QU&
PB;!#2JO=07%FI]-9*6Q_XE."+ME3!/>K,9>6C[)/,M5GQF !_D3CI'#>3Y)!CH/#
P\?M+M8O11<$.N)(]V>O%CBR=G 0:FFB=V_!Z\>\[9BET9+*E%?4Z=&..#?6BV?$5
PIC[&)V,;\PM8 N8(\Z[:3&B- ,/<.+%D&+9HCCZ#.M79)LNFM_E,)QQU#T#L9)#W
P".MS9,:<5BO)HB*9",D513MKM7I]AL;>F0C4 &%)@.(OV-?#LYC<!A:]C_#%6:*=
P,#122S]0$1'CPNCUZ)U^W(=[DG*85H?\,?8_&OC>6(B6U0[S<D/9:\>:=K=#'/H]
P[)[-$N8AJ^*L\N"1]\T )ATR14=XR9=Q@0(]?&RP2"R5:'CK33<E,SLW>[;(>\+"
P!\CBS$S?E"?02A4(=U!BS!S8^??NOZX@81+>)#AZ3VSOG1MYHHGW-RPN"(2Q$T]+
PSIWUW$;!B?GL5QGAFY@H>GQ_[76P15L([!YE>/>(\\B*@A)* NAR 5)F.E*GOC)S
PY\$*\H\W9YYBPLB6/OM6=B+PG#A71@>$_-(VDM@K%J[);#=OJJR;F6K9S@81S*I7
PN,,GR*OG*#!SQT8>;<>FR&2^8(LO$TV59R"RP1&9*=PGGN?;["ME(?%3)BC.>#6^
PV%=!S=&^H'8@<5%OLQ>X(F86OU18@ TOO'54LF]<,]=ZTXC%892MK];'H("P5<;V
P5\2A47+2U (19B NH)N7J;_J79H2",88O_^UN7&NNDW?.5]4?OJK)7U^#'B"3<?<
P36YVHD#+O;D+YOPXE;CV.V(%>U1T0NM\;>"/5(:D1B_+AZF5B>*Q/602ZZRM@!W?
PS>OIJ!*S.-1;YXNNU&=#OCO%]1[1%1Q<A\5F!BA$^/[)06+#KFHIT^3Y(I-S'36P
P,Y(S,!)I2Z1R/)2 =WO<%F2AU6-(P/\$CIAE5);&N\*5JIO7])[]%N:E:H#$7X/F
P"<@WKM9KGJ'J'PWB[AG@/4M\*Y?.%EBWW3<TC.!"SX>QJ5@S',49][#/\/)/^\=P
P/^%KD1H%_AO !X[8HV",5V FB]HB7SM*@[?+A^$WY(L*LZO-EG%:*S.,]^KO9/;B
P\I9^:A9R(Q__95D <(6=RB*^,18T+,2DA+&/Q$Z)<&]W9J(UN1F]+B(>]VH'!' F
PD9G'E\S:=9OR8M*=+V!DPQ%\/3)E/%G.L@9Q 1,MA+ I2;4B^!EJ_"S&:2+#MI4:
PI@&F&'7$;\-U@?;?=*T#[773:WGTW\:8R(D,M7Y5*\5$KS!KB5N78[.J?_*$W7!Q
P298P@'*OJ%KL$3']THA>EXK&"8[()GNSI)A\.WC>-NK@6&0B8Z27CV5!G#;L6.2=
P6E=ZZ'KI9MZOB"),)8WE2L#]/R^37(PTW72_DIW>5#WO1:3^OPD+K5Y %/F#/3IZ
P!@R6A.GJH(AE[-PS617+IL!K)/#+)5];5*SI2P7+%1B=P#EA<@^'/-P.BDB-A4Q'
P*'GU:RPIHH/5XQ2[-/&7-^%W(WD6:P-0LP;KL,0$!X#\:7E!*X9%JSY"0*/@I@IQ
P2\^3,W\3%6.\-.6NZK^5)E$301%B&_")07#%=9*UL]BV/%.D^/4?@K$@VZ<+"L4X
PL&^)&/="L.<.N6 T*/PZ']#B/?/]^+'Z1(%QK'DT/&[)_'[]GZ3?MUPIP#<ZG#>N
P6NFUNK,W?[4!+@/4%4.&)<GZ^:5-&=/>("="%9OHRLQ5 1[JP96;GU"SPXX_=+$(
P[#0T::=(9&.%@%%J\5UM'\5P'OL]A(87S)3G</7OFL8RYR9_831M%F_1G,S$5\#Q
PK).G9]-CS$ZG,EGSC"A80+A74;&3+[AYHUDL<,GF?_66F7\@.5/+W.Q/G_SX(;ST
P2?'.0XWP,T(J;Z[J]MRKMU.C8& &D/_%XN_Q<:92QV@7)A,XBD3&_%F]YT%-*V7$
P(="X<,7K:>)@2?*O,ZAO3>>D0,QZX5E,G#Z6;S!%/B9VAWN5=+Q""+F]CDZ30!K\
PN2-V-26V93QKAIOJC_+<LV*-K2F9X@?H+,>)L&.3#0D6I/ME#,,_1<E.EQT$.TAZ
P6#YY&H8&58:"IP[^49B P>+_1"CA=+^=L$?CIRM#=M)21'G)^4HE;&A_N]/PU!6'
PJLHW1P@N[(QS _2T]9F'FI4>A2OV /G,Y=<U@UXW]11R<T#N_0$0ZM>JX7\VQ=I"
P&Y=2VFQ5KQN:_"<K6J#"DLGU!AM(GVY]Y=Y="8B=4JEZ%58MI!<R.&&=]?(C$\]9
P5_C"C" J]V@JY "!Q%*)"(@7QSH.^]E$TB3(X"*3IK 1?W;DQ7(!03,'/M=2WSD&
P?S]>W&$,0#$[U"(E&PMX1@=!-.@%UZ$8GBU>6WO:>[_Q>H_52'**#N @8%U*V.',
PF6[O4=UR5M8$\I)*EZJ9D:2OQ+Y3>02WPW.9PBBE5#)?X1"5A(&A>WR,.GM*S/90
P'Z@4@!W((3>X^M6*'#V.+'UX?VM'_S76AG=$07CE=KOG++::M2+$9K7J9U2Y:$R]
P.>XN!=(G/#X81YQHA,3F?6"QS'9*&150+,3TIKHQ];@J%^'XJ%^IEBZ##__=2+L[
PFA(?U=90=,]I]&7+:T5<.%B1SF>Z01@-85RQ1Y.Q@\;^YE_;86VJU[FUPCE"<2<#
P#HSKXA6S@S1_07/?#HOW#N3S. [#5'ZL1,#/QI_(M.FG>="Y]CA8%NIAV5*;DR _
PD-EI@0ET6Q[7UCO#(7TL#3'"7@/8+QH$0]@6GQPN*7]M>HVE* <J2"9N,>^9<1]D
P5OHOI']D!)_@M7>FM>F>_?085T@A[Y,\!<6UCX)Y,8HR8@8ZO95GPAB1B63PS3NX
PJ!-#GCW9*H%']\IQCX5__?X#*H]#RB>U^(]L/$,L<T#X)XM7I'@+2RW[%'V+/!'J
P?J)PJFB\K;?MT!1^.-Z!Y"/%?]CORU_=W8='G^$10\1K4O09+FM'4VI.[/D#)-?X
PG<C8_KN/_'KROQ;SY/_H>X4> <=%DCW5UZ=EO?(+UL'C1@H""O_0.]TXZ5Y;7K-D
P*I6&[GD X(9U$1/P-/.M1(];XUYWW-L&-;.M)7'U?AS,.QRB%NWC$6S)"U-JG$C^
PBER&S+>D!Z3.,^L[(_=%N*(5!M]R/T'<_QTRY^F0K=B;38?)N99R%ORMV/0X6;TN
PHHWKB):XOP.$F0@GJ3EX1C(RWS)B$J#QF54$+1,R><"#[J7QV^!:K.4G!Y8=AU?F
P9\@ZG+%IY@@+%0[E>/]W4A2JD5<G]>/0768BXPBYCTH(]";#\ZAZEU>IZ+<XJZ/@
PB^ EX5D.C&>9S&S'Y+H4N^C*LI5S)1O-*XG/M912HVL]'<&4#8\C'0'F@,D'VC1&
PQ>#UW'\0133Z=17'3]!>TJB'.@"_Q8U8V<<O"YSWDT:VWL7I7;&P?C40_8X*WT"N
P *B^0+7,QE9=?UO]4G-RC"3>J0[&65_W]Z8RL8K$C\8[U)&=ZTORF8RBFSLRL*W/
P$2KG8&H-BW4*M_39.5.T/>K1@OE=D@>[?VV>K=<)*_T>D#LV-H[E)22_VBXJOHLJ
PPOY53O20--^%[QR+^2B8B;V-HFMMRW$_>)*A6RYNAA-F0 W;R\#5EJ3U3[Z.JL&>
P:9"<U'?)FCQD^@:8+N+^H8?/'/%I@CYRZRI4LI5[;I';([1^EG%-&W?@DONJ..Y>
PTG .#R?BJV4.35TM+/B3Z'\2%8X(@T?D11A:T\9A\-.C1$  ?+R(+((F9'WEDQ%*
P&BO%,*5WV;XQ6(12-%;JU(^@/B\L5[#\=?6M5 O&,Y-;+L@\$EAC3_^U_]KQY +5
PT\B X:64N&Z8!]2Z4@KQ%BN^4%ZY^&WGGP(<%IYBR<;[2U!O57-'%@K_>J5&RD",
P0V\]KH'C?PL$A"[C\<D:DH%/@07:)4?/$]CSR=8%M^92N:M4Y$P-S4P-JU&D7,5R
P'^_6\J,PK)$$&R:XRYD;9<NJHYE<I5H7RVE$#=_Y@.V2F:9APZID6*,LOJ/(Q=9!
P("'*;:QF_;@U!*']%(=@PK"Q!+F(?WS]MXUTIDE% ,>@ 3/\KN@W+SODJ7*:4-M]
P>Q@ASO(61,NJ,8ET7]ZZ!,CY R^>X;_*2$('6[/2;)]3.,9T\Y\MI^7P=E919](M
P;42HJ-,7"PK8-_<RA"V-'$KOLE+PSK\O)"31>58O+*13 YXM9!T#?,XDI89GZL$_
PSG/$=+86\]"ZV:*3J=RD  0;YA&V+Z^6XR^S[8!9QQ*SE_&+J?W0LCG=HX0Z)2$ 
PK&I,6,0QY8#N!X_/@3ER2 SC'N' 5VOWP3A]9PMVZ149X"$"C/$\< S1>ON,\^N4
PGRS5B^>7%#7]@*D$=MWG"G  ^B:92RZJ>PJSA,)L9^6@N"YI16!!2X#%PK_>ZVT9
P:<4;:CGCXCL;KUC@4U0Q(7O:?0B@(N?0!IE1T&&RJ&2_P*\6]//<ED2)GIMH-V&!
PJID/JX(9_1X_X8&=NS8I_L-C$ ,*W+,)-U-[>$+13'V;V(A_%"_1:1*O^8UWK?%;
PX<L*?;K72:*(&LD@3#*8ES" F>-4"=97L26B,&\D9$YC%OJ2A/ZT2CY!L1/%,5&Z
P2.]*^\_/'CNVOK@!-F<9FK!@+S8 ([<[Q3**E_3';ZPWS(*M3IM@P_>RJ&L6TLCI
PG/\2"YZ+R\!.Y!FN?*4_*D1_WG-&B)K]'PEZY.E+G%/LN+A1'E!.;I\1'TEH3NJ>
PF"3^Q5?1OR+"2-*LEN3&M^/4. R 8\15,FDI\;^NN>!Z0*22<H3.-?3N/T&Y\%9H
P.YF%42Z@ERF>>;^K>"TDI833FB5(%*)I1H!"&"Q,V]N[63N)&AW1,%FCCF9;= ?6
PTRH R6)E.:!*-Z@L(/-NA*((Z1)YG3#<_OH]<<9\W8SB&]J6*P!;D/=M_[K1+GL-
P XO!)+=L!ENX#F[XG6%<2BB<"+TO74A+,@8C6.,P]R5>1V=$IQP0IG"DAUY22'6/
P,?Q!U>CU@,V\G EWY[)9RZ#D!3MMS^NLD)1 9,VA.Q)Q"Q+\RF.KN."RZ4<:,^-.
PDM%B8C=GK6N+E^!;<V)$U2>2QA=;1_DO$2M.SF=/4[O([B=R9J<&$I>9'Y40J)*1
PGF%,4,RK#4+CO0:RM3&P+ @KL=&=SF@H^,/NR'0XQ?XOG59N\_*P[BLL'//&/M14
P^GRF:MAILZI<U8 RJ9<(66'W>C8K_T5S ++;X]R?.+<PC_:A,Y6L^<P]+9"Z$KVU
P<0E7X-[J%M[PF$F4M8F/$=M2$H_2V<<W:Q/N9H/>/S:W0P?Z.1=U#NP7L?;!]>K%
P!KR,66$,.\X.4=D:G:HMU15?(B\&31OM 1W"JF5\NYI[OMD&&)H@&RI/E);'55>\
P=,,JXM/6]4;_KT =1\46U9!2DQ!^6/=SB#P/-9@,DKIML!! '8WJ.E#9N?N2U6&$
P(J-60RV#*U\;W=3KQZ:O64)"TX)60A:!!?44"?2&)R^>?]5A;-W:/W%K%P3 LRX"
P*@Z-$0P)M,;CU#XX?*FX_F0-#XJ'9+Q(HOX:UP&D;L/3/F&?X_%DU$GH!%NQHGIO
PD;,!@CFUI)OT^3[OV_W2K"ZYBK.Q+=&>P>/*.9WAGJ\0$M0E:(Q@EIJ(.UX5L+%Q
PDNV@6=JA4!72B2]3V737713[9&TU17']V [Q;Z1KF/FE$FC'&QED\/V(H/-$U@Y5
P>]K%DU^*>L3VT]7.O2#^@E:FW%#2R*-X<>^X#=J391X"EU!20<,_3"U+G5KR YO]
P0$9-C)Q6 ZRG$H6H8J,-][L99U:R%HS.Y_!]1B!E"Q#))-D-!B,UHL3#0>8*EF(J
PJ_75RE^#<0Y6&*G=/PO.,O1_$)/PU%#,9T0J$=4])(Y[T#6E*T"72 %; ?*E9GFD
PV?GT*G:OBKE],>=GLHD+-7&&7NLAW-K2=*H#=_"^TI#^U]74N']$([V]33P/#O/-
PTAP5#_D CF?TI/2.YH,UXW X-F4$,Q9_N7B$:EK3D<K1!00H>(W5%^.R[E@^&6WJ
P2G'R:J6:IG9H(Y)S]'V0;/HVNEG\PWTO!"P!.P4%,V_+RJ #J0(-8NOCUUR*,C*)
P>6;CB:P4O'O)8+IS(AK.7/YD@+]B_B;[(2,_']IQE?E[!Q;V"=$1S5C,>%8&[[0=
P-D9'3$"RC6?746'572![3K[U.<_AC=EL!#L6G"8)"?W!J<4;XGZB)S>]"4W948,X
PE]P4!^U@7V#,%*'_R]>?-9A;S"2@/97]#UR#9S<6"4I# I',9&XL-'.N,HN3WN=?
P<P2\4:&Q-8WL>+.+J >(*?5/'*I_Z/?Z7QD2]<1[X^[FHZB:[I56+[@-9O$PC>F\
PC>8$DQ^F]<Y5W3S97O,51.'U;[I:?OZQVO2U<#9$;GGV"E4?1BY&NM*_BT")"NY6
P+G1O.3X"3RT8T0;*[IKL!-!=3Y%[0D\_<_L39 Y '&M4DR+%KKL7X"N:.+TBX7=/
P>N.2<MB;$*.8J/W*5_9G9K(+F58^WJ,)TIFU4KG#U!$/#6B@ER#_CF+RPBMT(LM@
PK%6OC6CC2+81Z;^Z).W:9PI!-/FV7L.-HVZ@.[(SR"Z)O[NX]GLI$%+6(;2KAG<R
P<5 IQ 31Z7U*UBXT@4-Z_<5E][_Z]O+.^Q0(T,FHK:% \;\VGI1,KMT4%]T"*N!.
PKO:EIA6U5L0)X?Y"MCGW_5;/MFZ^P")'7],R'X3ZJ5N.9!- ,5,',VG?GWX^#'C1
P8J-?:_XHRLO<LAUG=N[CF2K/=1CNPU\X !'".J_8S<5J5;,>S!>-O#[IND(D2@Y6
PH<\$"L8/^=4<CBN2J<V9I.Y#\\SP8HL\,&R= )AN5<WK*G3\(VW!HE&<\5VAQO^Y
P.J*KIWQO*_8)-7GQ%7C#SJ$QBM&JY\_#:-'!Q4Y?;\FR5C4GYV$8JP20.C4@@77-
P?.%MR[IP[>\V_Y7+\S%'J$%\F"(:;_%K4_1 /DN>GQ:-(GL$DAKYGE/3#-(F4-[9
PH<=XH+CSS!;P0+_+RF3D-&JKZFR;UX<9Q[,X3YTSMY*._(99KG;2VC=O"+,^)P['
P"YL8?^AKFI0;"> 2\HEJR\O\Z$/^ND:8P3<,T9+_</F0"+OL);41;AS7BB^?.;8/
PN_K"^!X0XX_?=CED1PQ<3 _B=PH"(NZ<#R;WE,;@,7_'Q<\+_^Z).E4X93"LHEQ1
PO93$/7L@;#B%Y6EL0U6C&8X:476=*0VXJ0"3TS2ZJ!&]'GP"0,!(.RH<N)\2SUG2
PL18^"TB\*]?&RT^9 ?4 7%XJ+#"Z9$:!7ET43]WW4.!HB=.,KO':FFH7:(;-/=0.
P(%.]PGH)5ZND? >64(^026A5T"RAW;WLVO^0#OLNM3[$_7L7/>2" X-D8(4/8N\%
P%(;&RD//D=3+8I*5JE21$;\<!@#!@I\5!A-V>3S15SV]!R4!H6(S#X_:7=<MIHTE
P7#0Q0:6[P+8$ISJ%I1%?DM%)-V!AO9#(5@>J R;ECYN.8.\^>5"=PR</W=,!RS]+
P0/6456BK9&DU-XR(N'$BL2LML.!6@^D@#NO:$\0_PIL"&^++\?=U<?B=.Q =..A"
PA8-U 1%597:N*#M3$:I^.;40&89.[J+.O6LD&RLTA)XXB^_8/8")>[&%[&G4,6_&
P17DC%*2'+SSI*7!)!^%:*JWP-$;IE+S#T?1J\3=X\').+#)R[+ZE[HL-!RH6#C<\
PI;3WV"^29G[GR?MK-@R*27]K[J);.!6"-S+1Z1@F7%I-+7)[U(2"(1.1X8;G,"A9
P3LYG*4A3\(.6JSI5M;GW+PP (^J.C%[U-\_.3&+\UXWYF[R%33#7"SXPC%;J,,GO
PA7YA1K<G?& '-$_T/I YZ(>(,()CB, A8=6/9V'T.)3)^@^Q#6E6 9H+ @LY;Y W
P[1BW*4Z@DJL^@G*DEG^!6C'!G'(8KF_$41VUJ=AQ&>X1\A?90/>\>+\\D>M#]M^6
P/1W$]M?2BI=$48>*ZT@,^PA,6Q;4F<S7]@^!X_OD50K/T!16U7;N8?0Z!:/(D.!;
PT(AZ\5EXB)/&/\&5@GW2>@"0K)7J.>M6]$^@^DFB8I9ETT25X=N)?S%74TF@_ #^
PR1UNT'^XP6[*4P6-@AW&<340N#_;A"[S#+,:+Y\<RUZ[GLB9Z)7GCNS+D4[*\?EP
P//="P:5L34E=YXB3#?4U$_[DX02?ZP@LDN8+]>06+/D((H1_*-VPJ_B6MX_4W U0
P"8 CQ \RS1=4/)D-+=YR;]NMJG%?L'W1PBU>>!9OK\=NEP'B$X?<@+J97&A[H0X7
PYS'(%CEC5[=DO=A)MUQ>$XS1TG0&;2U&5^A^EU"#WB1[)37J0F3R%9*4L>CD>_Q2
PPNZ9GVD!>A>#NZ?@MB&<"J-HCB] $-Z]^LRA+!_'T*BUGE$(-H;52.TLT@8\5^NQ
PZ\3!0JE2RW+'U\VP]G?XH<CG<<(#:1^D>*DGAUDQXN(&NL]DQ/ZC79%%B$#6PB*F
PC C^YTIJ(BU6%RM##)Y7.]PU_??.QFE>+A"@.VGM@%IOT9Z.5"+'ZNNF17U2EM&V
P7P(FKI,HPUGW@77:'Y@J)X&8"'X%0 ,PN">AX!M6NE:@J4;L%C9*V=*(O_&WCD1G
PCJG!BT>&X-E2'-B3 K#2/IXZ!#=],((\G^[:!>>E3)1][9JSK)/YI^=$C>"K[4V^
PI*-R=QD!Z1MZ!(:\U)CX/V@VNK_TCN*@E:BV" _ZD8<TK\!F,KMN:.CS9:DQKKK6
P6@%.P-M5S[D\-_]AA;<9:C9G2AR'GAX>VTP^_!E42/$D@U!Y<O0/08AB$L9OS7X*
PUAWGM\&C=QB9/PBCU'MBFR'$I-L;I>_8%A[S35Y5J5E.@FI*8V21;OY)35MT33A?
PH,N]/B-8=]M,L?(*7*=JVS[Y)7[G2"5W93@KU!AS):IRWWGE 2"*W:2)IK00N,V"
P!SZ6YFFK5H"+N,2T\PN9!+W:@!=B:$QF@D?7!H&ABN=55BSA'.A*7S[I[06 H6+^
P'Q$&A/K0WV)%V?&U=Q%L#,G@KT ;]X%SN67B0=RN&_"V[NW=44S=.^Q=!!>P3QJ"
P3+*Y,5UWM_4ZB><CF,M<'7I-Z&])Q=>'V._=80Z(4TB*./S]#+=TZ IFY'TA!]%L
P%ON?W@.S<;D83T^:10=$P',MC5O1,GY@+#)^HM>X'[_ Y("H&VZGF1?C_K7["H$^
P+8]2%/#_F6LY:-.0GE2$>6H?#0Q?K91)J+ZJ0_!YH->U&Q&LHL3\.L8.Q]C((H5D
P!K ^^-)J]$PDRH9\U4X TJ0P"( '_'Z7!_5K46:M%V^MI6KH,:DDP;_FP#&QR4W6
PGN05)/T7;7$#6^;HYH 2P,N9*'F4B_U/ ^MCL0/,(L4](HF=C[P]_I?V?I%<3KE$
P\[W[*"ZIN0>S8*E?9,9[MAG1).\DWW!J[C1-TD39GC-*36+\KL5P-U.";K#M>9G2
PPQJ3HZF%7]>' -H4.T!)'?I*;*2T^>$#H38_XE+\SB.HMFLB!]<W)+GBX-*8)@8\
P#W221G!&2P<]W ROMBUS*5,K]R/')-/$BL7FHZ<P+<)GX<>QII'W63DUE<!X*/NH
PL3F3U]@A^Y_R_^I>HT*<9#>*E67IYQ$J\R\$Z;VPU76$Y>%+^F7,&WA@<'.9<%;4
P)XE48LR-Q%OT,TX ^Q4>FM?R5W7]/)*H!=HX]/4Y*\CZYI#F?_A[_I?P)D"N*<RT
PR3>$;Q>#)EN>2IJKR^Z!:,:YH!1"MR6-Y.HP;F-=>:;)69//8 JCJKN2D7T[TETQ
P&8O3$R_\Y$(A4^QK")CJ06XJ0%SR#4M"B3ZR<[;@*.1N;,=,"ZW;)[+6&<B7ME^=
P975+%XX_ZL2K9?%\Y.:$PBBA57L8176EK491*>!MGHY%2@<>),G$@,W]R8QQE,T6
P$(TCMA\RE(ZR3((G/)EAY>M;XY.CQ/.D38NI35'U6*+&3&8RG:39C%1V)5RIB(-X
P2O-A9CLMV$SM:E,X)7I/T=N\/!)3GOJCY?F6@0"]/J:M[1/ K;M$@$WX#,)>^N8W
PON=]%>*3WYO3V1^IWKVXG:GWD(D.N5BYV!<9P71G0:1C$F\D"%"E\!M+N'7P>"$#
P#X'<F8*U[G(BV_J9-:N1"FK\R+B9>C\/EX*2D-=[8TK")/V\'%2O;XRJ JUMY%GC
PFA46<4+ ,\5IKJXWO*FP:,U51W'\N+,#O^2#?2?=). P(-?)%*R$&ZF#]*C1W_)Z
PW <FV_%%ZEDE_[B;'F@"X-RSFO&-I$QB8%LXS%BF)OFRDB.2^KQNQ$M64K'#<P '
P+R^R6GKM[R\>:39)I3+'@PIC7D$,7USD783DU3U/'(/H/I\2E>H#4(W1Q"Z:$M5(
PBI%_^RQ((]@T(^F5PB4$.B?"78+GI0]HR4P/7TYV3Y75P44%BR,?X4^:YLM:W/WV
P_C<_#A0:L>IW%I50##<,J_^[CNZ]82\""C?GCY&G1GE0X-NDSY(Z1E'5APK(N8PR
P0(?(,^1FK; # Q%FNV@>6Y3M)U5+X<V^B&?'HD<7&53IO(88+!R,7Y3X)@;B^2+H
P<:PN[,7%&H>W&3=ACH=4]P;7<1K+A1V(.L=6O:PVZ:>\XG0#A438/AE$T:[T%P]G
P+R8.N>QX3*\G#KI2+&MEP5=34_AJ:6E: RG]L- _@ __7C/[N40PFH(A"N%"ZSR3
P%:HS?V6O;1>SHV\.K/:C8 0A*@YSP1K3>JQOD@V6J4G=(7>Z#\;*6@B=F7.,8K5N
PR) 3JL=B]!4?2\KYVMOWB+X1_A6Q;WS>(^B23D;6.%H?VIO VE5N.^<N7G'/RTXW
P5,R!^+BQ!"E+_%PR?VYU\N0X^+'';ZCV<U_:\W]\\O5M[[$5J'K %-SOP*;M*T,"
PKJGMI:.H\@C(C0D:&([!,>-8;'!:2-5,^[.Q<EMS2FDA5"TE;69WM0+P D[-1$ Z
PS]%A8!7M]9/&6'%2>KV7A>[LA3)AK:$QLC)S<'-P F;C(S Q@E/Z$6EKW@84ML^H
P2/!3E&*[;^EX<(3)K)^)/L"A^_]9:'U80>L9_'B/+,!,S/^K8# 1$N=X; .S$2LL
P[EM]2$Y:=>\(GO!E>Y_!6I>P1W!L8#Y733P+;D4^:8=5>*,5'UK&&7;Z6"II3IGV
P4L/-:3);4M?'U.X'^;L> M(A 9-.]5?PB8:P&H7]L3N:#2*23/G4[FD"RB7/>DVO
P59HHR$E=*R"O*&2/UJ(<_88WAKKCQ*S1^9F Y9S#0(KX/Y81^'6X#D<W2U4*=$4$
PDB<*L"N9)C&(Y7L&O'?O0=Q',5PQ^IM@][C1_(I!,I^]L_WK<3E5EE@L.I,%GTFF
P*!/R!4SX&Q@/J=@AZH31U.USO$FB:N0K=V-2NF+#1<1Z]57_ ="N%N?^Z$\52\JF
PAUTYB5(/S#'[5JP695,1P9C,;?^?!,_Y5\<+08+I4Q</HR>8PLS.!\0 + G^VWQ6
PQ!V!0@N6"==0#I[XGC2A['$)DV3JUXNZ*X7#DW7]D;&OQO=^KD:<:Q\OV^II\@*A
P)9 G1.4N#TK"GN4J_1 (%TI0O%D%>L9L\SK[#$:SAWSK;K,H3ZV%6,-.C'=F.;^+
PG W3]391XS7[; _:S(N(@#I(G^.^210J3] ]%TKX\WN&7?EXP\01L0?7$[.;\]1&
PD)QP.&3#2W?#BZ0XM6EK/4$!_A]?#"H8O:L0Q^21"**^+V:,5% TEKT7PUP(&CQ:
P1L$2H\58+_UF4)ZK71-S=.V(46Z)WV]0R#7'S$(&S\=OVF9)Q3YB/EA-X:/(^5#T
PK%%6E@:PG8+G=+K?A^\NI'J+O"!A?ZIA1<IQ\ZEYUPY/)H3;H\M[2"#Y>Y]O"2V>
PW4$=XB"R39GF>_=] S'PF2JH#!+[O25*N+'L.-83B'$Y$$YA*'HVT[$\?H\)3026
PA4VPW_V-OKD!5V5C!F;J_NY<P&:9. LG-(. F+H-RX+;K2^?2J"Z8"*R*^]V\%!1
PAZ?*91KI=^L[O\[F$)ECUP<CRMFC&TG!]\,TU GR>>E*)Z+:_9\\%_35!YLK+G[M
PG!Q<':H;@HRBP"DAM"PV,U%($:;-#>!,W7Z[C4.6#**PT@Q//<H54I/70 TNFF[C
P4,-Q8(]/71!L/MC#_ZR[E9S)"9296H;7$[[#6D2INIG(<C.KJ\Q6/EKR%;\R0"1#
PT'7Y<!HME6!5Z+I!8,\;35E&(HEWQGI3,2]?'L!E=>T%(-IS)-WN/@EQ'8EN++5P
P10I*5/?%C^)XW#CX\D6IH+6C^\K\Q8*.BNHW<';4K_4D,)H3$:\TF'XS?;!!8(>7
PHW81] 0-.G97:.ER<"2ZV<UN:L.F"8X)2=K2N5[.=Q[&_<V?WW#JX0,EODO%T#02
PM"T..VTBUT,;_N%\D$IX(?K*^F>"#K3&3Y/N?K3LHBK07WL1&D+F"R5-'-&"<L3S
P;>/L B=T&.T/U5,^'52."/T75FB&S(UK+HK];(Q\=R?X@6OC($OO,Y$TY@._9SK5
P6#0ZQ7U02MW]/*CX0[TD<]")$0Q:?58IWJ%<!PGR M'WOMLV&B_&RG,.V/'@)BXP
P[0&_8Q+O1!V='W<18$?@D[X#54Q>1F&<0(7 XT5VI4<2[3"$FM?64;D.ZW3_B/*J
PY6*9Q,_M#9(?-SBTK+#PIXZ&"=M:=);7$,#+,Q'G>RAY2&(-R16!^G_]5HCM>+-!
PVH/2[MQ-7D^L3$T+5[(!;?X"[SF$+-*32WG;+)7;DXQ>7%\I'&>5?4Q[TMX6>7%*
P(RRN\?AKK-SZ R&I+&H TF?NNR3ITWF8,4 U*,-&Y2JW-GS9-_2UM3P\WR:LK+_0
PN5/8</)FG2R"A%8,1H;$C-22\8C9)YYHK^D=Z\-)AN\+.)/6-Y#$UW]1?FDU3OD(
PSERENWK,M<((?$1K\3J/__^%?TBR:ENU9G_!=)3N$]>%)-V:6.4.*B5M]\8)Q;"7
PS2W2Q=E0>+:1G"\FPKR][5$:0SYW%(5G-060Y-HW 8QV<6[P"%V[0U5OTY6(0ZZ@
PZ3 J0D!WN3][\&$"#.E,N.4SCB@JID$NT()8USKE9IG$*K=],&;)2-5Z7KG #<AK
PMY,8[Q(R, 6FUI\Z^7S'6HTYUS*,!P;"NF@;&B/H$Y=2K?/Q8)3_X.XW7(4IL(E(
P>"_W9-&OJ/4@.IDAG("HX_"B,)E) %PK#4F!UN$=&HA^LU MW8_0JTK.,":+I]N2
P%;$)]O%LRF1)<ZI@@<%/ZNL+7D8%KD.]*,,(&U+HUGMKM%<2ZK32DH-W%7,- RY 
P]=X-'76UK1J8A6*3$SWLM*5!>ZVAU:#7N@)+K+'CR&"%+@A?#OPV5\LGZXG:"0]S
P062D)OA(8)8J&A2%WFZ]1;7:J%N?)PE:LW)LSMACC\O0Y2:RR=/?!3-$PBG@8E12
PGN[L;.L7R$66.-"'L^=NF H#.2U-DCVS.-W4ZFMPO'SY6V]US?69C!5V^'Q-H*A8
P4KD-"(":W*LY22TR39%'('T9[KKQI)4V7GF(!<W ST71+ '&!XP'=8/".37QD X.
P2.+-J\LT+8M[ ADUB0Z)S_WF4?PQ?E?(FM%K^#7AW\*+1QX@7V" !1&$T78CRX+_
P'JW1_#>/FT!5;X8P^(M6RZU@@I?;N_:6KU.5NUM?VC'+P,)C?>4];H"R863S[,B?
P39\#J?N_O%%#<)%0V(/A[U L@O\4;3)BW^9'! ;R"-6^F3HF+- P-E=R"CYL#-X?
P5WQ&9_/0DFF"=9_2L7FRK#V;\G06%39_ALS/C!6OJ=[<4Y^"?=EF -RFTP0_K4QD
P^GY&<M;^/@,4$MD^I4 H#=FN+),H9V#*YQ4IC R/8*/AW+\GGD4_L$&8>Y:EI^Y^
P1+WTIAS@;.K)NV =O.0'8_!Y2]!(S%GS?Q"DVCHAA+N:'V9G=N+3QFA\,FFXZ)CU
P9J=F9]5VF;<^HR'E\[5V@E&6$?J;0F\KB2R>3\_<WUBK1M*2NI'7AZMSS^5$#WBN
PRY. '%,?T_GVT>A.5SK3=24&VQ6'_JJMO4<XC+M><T([7/.%3'L31H?LX7E]FAA1
P<[H&@6N/\_B3 %D@V!_V!D?-TL93*L!6WO7FTL?:71PK/ BA?,4=0&R3&4Y7M 0A
P$@!R'L3QTMZ\V02H)EY'6\ ^3Q.Q36-S.ZP-4VB7%J:5,W+CQG;UW;->_9BC( '?
PP[RCE)M?<-M"6SFWX&K4[/S/B48L8I*7&D6$!3P^JF"LP7I:=/JH)@T30<@ .^U:
P2BI ?FOY"BH:+--\*&*,S79<3.@I2B,^K$G$C(A4[[M4\%PM26-+5%=6XWHF2/E1
P.=.$]+S)_]$:PA6"@^',B@<E;\I#5\21>DB)R>\9UV&];CMXJ>CJ*K4ELZ8?=,)=
PFZ1&J_Q['*SPFL^R3$*R]0OXES,IKS._0+OIN[GLD@R4D!H%]O,BJ -NQFP"" &V
PF/P.1AL@)/D4[G6;^!<5P!J#Q$ZQ%JOA_9NC$V"3!%E+25@FZEXJ>TI8PZWFG2=Q
PUB"Q3,@#+6%6>/RVED/BWNK=D+E)6D)#L^^[<I*Q +8CJ.L+8&61Y1QV-TH42:R0
P'1$#G#MBF.LAL/.WPK$YP4<&1@\$0KV%!QH$?;NZ<P S5]S="*.L4SB[P_5*R0?&
P=+Q/^I,#RO]ZDCS!]EIAEESMU*FX7;7RR%-@M[QN-=[#(H#WAAW'V TX(@V+Z*_F
PX[D:C0T4RAS!TW\W.O::_GW9$]S;!5E.Z"61L(P]H#^3&3+7 M9>[A]:A:$+@GJM
P_*%!Y?4M%][+UDXETREX,3CWM38K,KB/L>*!=O8OBDN&T?^ZDE05BNO#_#)NG:##
P"/Z%%$]I@ 22D;V%;=AJJO#>9_6+>JWU0WVOU R%;_!][L,J/DIO-$!]^_&VZ' )
PPD00U9,:\>*S5%F94<<G13<E2ZMJJ3MJCYIC7_Q0D/'VZ"GGM].SZ7K/@#T5XW%R
P9,NJGAM8TD^'O-G ZQB"KHX)3H=#@A027ZNM!VC%0P/Z^\P+LP2:-?>&2_E'(6E=
PLR)<VAUKX!9LZ<J;SPK/I9B'B["&B"0Q&%4T#Y9]Y:"S/-N+/J3ERL]@%L/WOCY,
PL.\=VS4!%))8 :^P]1'EM"MB(@X257%L0CZWA$8[L:(""_HF:6+V\^:O@LT),:%Z
P&I ,Q=N'*'-7\OMP<YHQ$<@B6//&O-/NHPJ$YDY=KB];7--I.UF'"DL'NW9C,(AS
P;P,+'PG[?0$HCCJ7PV"*XSL@[Y(HCPZ >3Z,.]P;W0%E&!EE3U3V>TA" B6\%<__
PX]Y*TIR*O*8U$H9./X#K+>!X'EJW;BYN1G^\L8W[R$'TUGNN,IYR* 2$5))=&]/N
P"\MX)W <S=BU:LEQ+#DH7_,B(>6JTX4*&&\G'B!F$S6<L!H1,IKM&O]SD/$%PB'!
PF@XW$8B/M. 7+)SVWCDVDM%*<LH(514L5(0A[=T*+*MXF/XZI.?0?DWG=/3&S=>F
P4T)[V='MN[8/B[6O_A:19/DQF7 (.UM8( B:Y:3CR\D@W;&79@NMR@;&CNE_Z6Z<
P +(,<P83""@;JLV6K+!";-O#\R)F:B:LQDQZ+T1X$+#';<R83J9YT)"'FX<QKD:B
P1\RUG_?P&R;V"T1,84MF[OA\O3D):%!DES(S)KI! #U 5]X#1N]=*V29#/TJ$+B8
P+6;6CD8KFQ]B#<E9W!#"*(?HZ&M@BKC3'2Y-FT.'^3FUP%1LT>@+T7%06CZ%8Q7P
P3\'6+F_J<+C<J'>W_,##5PD;VT>&J>W%ZQ%>N:&9%)@-'"$L=%'PVC@.3'U*?ALE
P\G@PRBJ(-=9L(,T*4^O/7=4^=[0DK:Y<>AIQY,]0:3)7*_@)EHAAQME;[O<GNDW#
PX75;)::8&__"#$&WB+KT7B/:9KIB:_X?U)4P?EYH"8_[&XO$TBD+_<!??#AZ$H,T
P8;G;/O\08_X>8)S5\BSK01VI5B$MM\J5NB^5NZ/L'&'D#88HURK6JXY2F6N$T1WT
P7GQ/LPF%8;8V[C9M5T.!9QB3?V2K2@,@)T@LN.4.):UX[(IX.'02<#_--/**V26&
P;*>61\OKOC:&7ZP#W$8F7?;,.[@/*QDP.6Z6)PJXRP$9[6&@)M :Q,\*ZEX&N]<G
P:WS23\8SP"785NL]8_.4LF:O[$P%6B>[>\'4OU $!6A6/(6,)F YG="KP6^^UH3(
P\4H%<9[46&+;$%*U.C)I\ ;-_?('[5,0Q2&CP%F0>$5BUAC:JR!_090OK>DGOI# 
P8&RPA?:U30H"'!N^I(48Q0-B'L;1<=Z.^&'/N\_=@K8T&_G[_MISW#.$%$L6TJ1U
P__'M>07+I>L-<2S2B:O+$8??J161XD23X'3%-7U,6C;8TU\]_G3K\> +.5P "BRA
P!%8CPSN95@%G)YY3RHI'NRF=/>E%-\#>JL]\2JA#^NW;9++W@*"A0&IS"BN2;8OB
PHER3?HE:(RUK(A%QQ3@#+.69Z$ *]);X_BPOM$S*"33L'KNWDOY38B:.L!D^+;61
PT<]U:/5/^;&HO/*:!B-"KE1?5MVX!X!T6Z'H!7#2[V\F$E(V7*KC4M_M>_[FSOG%
PZI_1^WTP:D3ZJ@D/=SV!&?S K#?SV "P2XV"U?F!&%TC;-2':Y.G#W,I#UP.5UV7
PMJ7D(^+EX:U063M#F -;VC["K_RM&^<7W%\<)?2"@1[CAK<+AQFE1M0XS P2+JG8
P CK)J+D0;J#P%544EDGBW'W-<FG34\<JC.4OG1C&DQMA .D+F><?DW_K&MUY$=2U
P<<\*:T;$M!1*"J)_4L"/=,+G]GRGHE4[]*H@5/B4[WOLB_SX4!%!'33&X496!X*K
PD*O%/4W!^6VZ #D$"E47O3/]L3R^?ILN+JW7Q;J.?+L$S,U!),-F<6BOY]*WYH18
P0/Q51GM*NB-5*T+WD$-7K$@XH!08-6J"9IF;:' C.'Z(P;F-U\E=H<A7M#X?I5?U
P"#&A8U.4/G^"7H]S; ?Z^6@IL>-,1++V@'AU^A];VL[4-I.']?&//RD.OFF*,'0B
P;;5'[&%=MGOQYV;I",T/R<PQ)E#8]3J>^ D]*K7O>U>4!N.\]$J_<Y&B7]EN/(\+
PU8BWZ*M1')#TM'&;*9D! 9XE;=4*D%(T$VY-BL.0]K#_!C#:<+VO1DT<F*!:FP,_
P]JXKK-23&?9D_,2A>;P&W%BO<]B=]\";B]+ U<C "X>JV$DBUPV,?UU+;5.8^/M=
P900;W8F$^!$,J[<<WWAU%TW#Z% B^@5<YX)_1XM+MDA1+@VBL1=+BEP=FC],PX4B
P?M(B])MZ'UP("_QOX#K$UM+S,TL@E='VLZWE79!W)P&99X#K2CM2R&Y"XIQDHB; 
P*P-QA7/L[2"^7L["A,7@W!:ZQ;5L&X,G[==?_0X%I48+^BI@V&-GB?A&#JM-1.>J
P/C%@],J/^RU&,$0K/,+2ODC&68;/_;E-^<V5??=)1/4BV1R/,S#:6XFY:UM??01O
P#.2C /2ZF$Y@%YZ/X.QY2WIR"AQ\!\,1"5\^Y9 6N1@"^C4%4-#11VHO,'>#%%C9
P^.T&*[-'1EV^\LH$'M;R6G=LCAT8;K! -QK82K ^ N?4GYW\1.+?2:LZ@?1!"W*4
PG"X-;QSTU)0=<Z@]0HA3N!+U:B7X\KV_J=YU]WH;"C[UVI)4O 38EH/D6PDZYR&(
P,6=_'O3<9_]57*5>6<KH=;+WH;W!$1FZN/_\45702TK*MXI KI0SC53CS8@'I:K/
P G;"M<<3')GR I3 $,GCJS^G=N'E)]*3TL8,!U"B1;.Z<E1?!@A_AVE"ZD\#5.A7
PJJZ?"B<#P0_T#JGL9O"26T>X$]I)69"=6W/8_E:HD@?U08XNNE5=\C(F%+52-MP-
PTPJ!%PMXV!%D3%?/((1"D-VU=4<]=HB4,I.[+Z<5^[I4M13?(":O S\@)U/>/ OP
P%/S$N<-FY!<E@L((!<Q2E*;SC6E$M)_[IZ+WE[@C])MV#XGU%T9:IEHDR1D@.H5$
PV#$Z%D[N!:D?Q1X@1FYFF*ETF_2)V&?IR-9>6;\P/@I8XXMRRB#S8Z\A+>7@RO_=
P&](VD1H" RY:T"<(.21:7E/X[/5R6QJ:#X6WQ!P-U#T4*-.X^-MB;L&.*H>O]+CY
PM_.7@#FDPJ2#^=Y+<+*!UET#3ENF1]?[V*LT'^75CNI>U(?TN?V9!=& ;B-YZ52C
P6;-Q4MQ+$8#<GO/:N:+-V\_;OW0<6RC$XFPW].-V7:-#[C?9EFR*RB&$XCIV^:A:
PH4H&L/Q5N+)H\@/EC3.+7\/48M\L<(9-%K\U]Z,N:6"OXTT(L-^@MW!8(EZL[ZAF
PY(#XWZ\W![8MLKN)I-1<O,)1&VCVBTTJ(/"<LK8WCI7E_U#2L>FPXPA,ATQ8'W!H
P=Y]'*#"7OUNF&[LC\Q!_QD_",]G#,7E=IR.1=VWYNN8-V8S@N\6WN'@KG^V?0WKS
P!_,JGMMA/@LBS)^S</XY\#H\M!9_3L!**V'=*&Z-4EUAHZOV 3$1Q0TWE_D!F1LU
PC6&SV5QJ3KVTEU%0;7B0'/7C(3^^I9R!H$I$5<H_C%^JY=;7\6R>Z*0G_:NE6$ (
P^Y"3COZTCR^0Q9$H(R8&\542EKBATZ>)+(N=ZG%+$;SG](]HL]/OEV7)=[;I^]&H
PS)UTOM\"#X<Z DY)Q"LQI'0&&._TAL'0RI19Q9NU^^4TK6FOOO.T*<BSTH5^;>R?
P^'BHHH\1'_NCR0^B#QM =NM%*IQX 14C9X)Q?>Q)\<K'*V]I;>)Y9YRP,P\])1K!
PTXQ\9&8:7',W(6MJ"%UUAFZI*YTS+108V0!FGSDBL*VO(%?&5 %P' )[ M3'Q*?6
P3X_,6/F^?A90%9;BF;L2S,0)(9D&F'0Q^X\6;8F(,Q*3QT&G$'0K\5=Y1A1]&<;]
P[[R<P[SGPR?B?!D=CM&:0@:7FHZ##RS]%,Z]\Q9U%9@&TLY9MZT\03#46GW@N,_M
PJ9E,PD802\0--5YN'"9OUAB\1E%MM!KJ#E%(_ZR$PY5 8E&<50 \<TN7][PRCRDO
PX]N*<-%K2Y;I]Q4QRBF]FPL NXX&+69[C=F%)[[Z0H9&<O&)H$HFC?H=+$&FD9PY
P&L=L&_"/K%K:=?#H)GW*D420N5]6]SY61"OB)>.*HP!$FS34*'?3'95X7 Q:I$<+
PQ3Z$2]WR#56^A>OGLOQV1RD4\(3H(O>&49S12966*.X$7W"I['P72<G'!33(;Y3 
PY:X@W=[7*!>%)P=B3\=.RY)XVU_]71WJ6UGO 6N4%7YMLL5-;>EXED/8<IX:B#Q_
P34NF7NU*RR\F,#%/_!>+Q&[3A$'R>T- TCSL%:[K6]F44 TE=ZS_;;L*9PUNQESQ
PEL$_BA,?H]]VB=^O@ZY@A]$YC:[/^\?MRTC,GNUS=^H9($ADM7F\'@P,(6 /7 ()
PP.(*:1:$3$00 >A\OH8J;$]O;(DL74.[=[%1)]*M#J;Q4Y.%#2S^@O&\,,VQ8,FC
PJ5@A@NFN>5M3L+26<YLO.C(HUC03@/@I %/'&CA^2@.#!7:>F_UP!8,7'B.KV\[.
P31'BR7K46,WDIF<1@+1^[?)N/.HMP5EI2-1\@!=%QNS6M4LJFTX79&>:S_[_=:W)
P5L@#D\"&0:$LAD4)'6Q(&A@6JXU'(YN*<&<591IHNN.TE]=<%&L,.WCS9EF&>/6?
P%?H6,^T*J\X.186\"O3C*=!$C+V'5'$5K ,%=7QH%'_]^EM55$01[*',S[?^6."?
PA6Q8CJ.6+N@'<'&.E*T&F&MIAFTN*2^Q('Q% '&G=88W VRJ45UUYFY8#JC_A54+
PQLDB@7EK07@R9"B=P]/0>[&)^+K$'?A)Q]RA.DEH_B:'3C/M&@_"JY5Y \XK'*-E
P:?4^?MMB64 \@W3D21G,PLV2&XY: 8PN]UELC4;-*(FY8)"%)^:F><=U\'(HI901
P(@O&X,0#A8H1LB?&EEW^6#7?ME=TPAL9(7( R_AMNC=>*&*.YU,RED@=(0!9)5L>
P_3NZ<C9VXP%B@QB9'L_J!P[MV1_A][S#@/E5^^X!YB7YG\3;A^)9- ZBX#XI0=S4
P/9.)RSM-P4^5X%R_"RT*"#TT2I,\P5+AJV]Q0R>4[ULI#:TBZMZ(X.%$EJH6-\^<
P5M#"56F_1\K'QX]0K#MZ)!G=ID&4@W=LDRW@DQ8'/6(?.MD+\XM;I4/,^JG,;2O/
PU8T$2?QJC#@N7%#GUS],1_(V#.L"%+NJODZ&L)EZ?)N4?I]20^\SB45)VZ#<"[' 
P!556"5-T.L4W[CLJQMJ-U@^!.8#6$N_H!OQ(/1+O1EC3.@;WKF%[(204>?<-0THH
P6!IEGF^WO5V:%:<1C*7-+42P?>;16  +I%@A+M/:^SA4ONR=R"8G'ZDJHO6!]NOG
PA80;''FQ74XR>K>OOLL5,Z$*%!1,W%$F?KGZI%S'2-4+YG4&HO8>F<-)CZF*E\0:
P$)M<2ZZC?LH9091^03>J<YM0 R*E@L3YQ5+3BF;I@__GT=1^AG[@IG]IB,H0PTUG
PR[V>:<^.H+=4@5Y,$Q\KWC=V 4%3_?7=']-(YKGFHHBL5R]PK4"<GL2O&#O>ZC_(
PNXTRV]WJ[:KV>4=ET8AK\]J9-IU\W!V >S2 B#L+KAP:3QXICZ2I3TA.7<]=6>&-
PG= <^VHR:; L$ 8*$Z]ZZ8*6$Z  AEBHB?!+OITY30#[0!B(4H8^Q>R;5+!JL/M:
P"QAVK7\(WM+M"?$S-RTZL#OBR\DY6\\#[>A\T\6<%"N:=\X0@HK)=HIU"<F_&H_6
P35X2Q!F"KW^9V[Z>EK_UK&:B]NV69O(P /)A]RHW*\2H4R;$T6ZKZ(APOJ5O_+LT
P-V91Q+I XEYWK6FJ&6JR;?;46&&G7?V JO  &O?>O'7=-%\6!DH&PX'#>*;(^V[Z
P42^;IIS)<RSLT@6B7WUSZ:^!9V"L[;;/3S$%!V#TN !'F5M%#: P+&(KD!T-\1#R
P(V252S1*C44J^,7&Y_'J18)FG08R3X&R,?SA=_VY[1$7RGW>-O$/'"ZH;8.20_2>
PDR^T'T''/-7S!#QMJP<./5X!I977#?NP2O6M*0:%YA(86[2TFO?D5H/H:H!\J]IK
P&4_1R40\Y1 $NLU0J7S!?GJ&V!PC31Q,1L\#AQCT::MW8C'$);3;8TH'[XEJ?W])
P$*QG"FS^3\IL0DAU\@\-W>K4Z[N08"XG%@06%--RU5]*$09)07,Q.,>& R=3Q]7R
PY7DYDXNEB5'!+CR8"5[>PA2+_D>XZ8%Y+-H,U.B!+X=BN^]:T-XQKPQ,"?=)#M <
P-*:H.6V0C$6._5FLJ9-[T(.SZ160_)(%21H/Q<UX<1K2ZE1RR<+NEES3MR]1;Y4O
P!RI" 80LHO9ZF4'-E8'J+B13Q5NO'D)UIFA8@9K1UK3V=J>\_+I<&)T\2JB )0*H
P/R5'Q#A\;:76>I*ADMIO?E)+#13T>8*BC[.D!<"BOV]_/ UKG)]DQ=]PIFO09BF5
P4?%)F8-BAZ0<RY+_>BA3!SZMA@;!DVD973]SOS<=4AY2G"[G,RKZ*IC[)CLM H72
PMW8->2Q0T=RBHSR2*$3)5CM]SA2EG@EBU0Z5-Z5*:P%KEZA=VE:OE/EZJ+X120+D
P)7EPIXX?;3MU3*%NM!(9##,8E@PW$.WWZL]01'E2VV) 3_^ED3\;"-X"GQU*4U>B
P.UM3PKM&HMW-GA;*RW8\JBT%K>4?(C 9>-\KKL+.53D%#<7Q"?#$6T%?"Z ?*LJ&
P8[F&9J2L)%P5&]Q\M9Y#S_,T5Q$BXQ,0T+A>1)78&VUD9PN9GP2Z8W@F.G X(>MF
P+W&6 ( O\T+DZ05L#I3691:%=8+F[OT?U?1RZRD8@,@4];T Q2&W7^?I9N?PS[!#
P7^^,8>Q9_V1NOTVMEK]W*C@KZ"UQIH5K&5+[:G12'K(&#A@K4/$H'A$"4Y-PS&@O
PMWZ.@C3I\]V.Q(.I^>5.7>QC)9*0<IQBR^ 3EA[?,VE:7=ZIDI]($A?J^QU0QSA>
P:D7.]]]<(6Q^A5ET1[_V1EK9_(263861#=(&7U:PH.(&%3YT5I[.B5J5)T#9W2:\
PXAB][!#D75^$KC,8O[J@W%:1T1O.^[->M#A',P3DGLAT?2<^RJ]AB38AK5[5 O!9
P"DHU>JFPO"4:MG1;'=_&!@9 #09I&)=I^[RC3P 12.Y^"CN[/U6(W\:[/QC#/7$8
P'/\A.!?;BE!8$:3RQ@$3MP\<$8JG3D%V_P.9%.A97&V]/V@/;GV#"-%,;+YUIS)I
PT-!>6$S%)6)A);C'8C0F"!%_=R@U;'"8.0JZHL"3.<9WK96#5K*!4-\>0SKS?GW5
P09\@!>T'3:[GM[^T6?8RFE5=>LB!>=_'A_'C))\ZA.!]I$=I$G83,^_J=<256]!5
P6D^'SEC<4=8\*B 154XWOEG)^V(FXVW^L D,?!V0#L2H:D FZYO"Y4W5>W?(NJ_F
PK0XM$GL6VU"2D @E&, U47ZSYU'86WXD ^%SM<"1(JS.JSR9P-P=1R<)3O;6'YH?
P/TB<^]U*[&A%(=_QP4JGV)#Y')/^&<1TJX)]>6Q@,T%C+XE4]/IEV+VC/[_7JXQ2
PT[/")I%!T1+^VH3,@1Q;Z!J)]PY=+76T[3]IM5N:,E8@1;A/N1.*[Z-:0RJXQ;__
P"U#^#XN4R65H[7 (X!D]%083O<VGG/-CX$J[TCR:+30_^\XOGO1&W>3&VZ6^8O54
P# OSER-Q9%UEX.K-* ]91T.UE5^B^95P^6R\GATSPRD#9-&=#J?))"9C6SU3RTL 
PK,'30$2\A8@Q-E8GEZVC1XXR'J+=?&3.QG=7;/EP(2N]=H.O]\[M%G!B(D8/SS\F
PR,S:8G@6M[5"<X5&T6KCT5/'/*UT<B@D#MJS13O=/ (_=\U%L6_P=O8T)9^["DE@
PH0GP2MP<%P>0D@Z00LUPI9:.8NU0-A42]!;<'\+C$IZ(2]N.#!;0<EN&0+F.##4Q
P72Q.)8\^CL3)IJ*I EJ"DVG#MY.TX7UK@)]OJ')#Q?@DG!'46S_=2[JFTO!YX[=F
P!B[J;>ANP7*](F]U;%WHIJ #0!>5HH8\FX0 [L-Y$-MR<Q]]]!G+&5JJNN??BZ2'
P)<2BS9C;\;>3[6-\V*A3=J8DR;4IKL'X+8H0NB9"XUUT%DQV&O'OT-Q-.I>2$NRP
P2OG>DWJQ1OC]=@!LAH?;AC"J'EROS21 R$9NK(S[TKU]\"LZ&G7W2\Y?ELG"6</V
P+/=J1P/^OOW: 19W)VH^+T/RVAZ0 [?H%][B,=MMGFSJ>UX'!MIGBRF8UZ4[B$<C
PXA_%>@U_]PRE!/F,(4>>I>,Y8VP $_L!C;.6I'>ANIUG-K,W!NZVJ2:\%\)_=^/,
PU$T@&)%8=%HZ3;@KB'X6G;6Y^'+G7+9FR$=_RKXF;@DI%B&/?7ES=K-E*[U,4N%R
P+7A3UBI>W^L985G 06.%&(E.0O)<+^L1H.FXY\E&\V^<G08^I_U&QAHT#*F/,MRW
PHG)^W 9ZN&JB>U"_K7P'EYSICRFOY4H"R#=(&25.&'P[I2.[1I9!T^.S[AVE&LGK
P4_$<3Y?(.<_2%_[5+?/KD3]EJFC;WVH=R\GW030U'1:?-Y1"CV#CPL G#E%G$XHM
P9.@84:A_0U%'QS\U\6E%EI.!Q_S6A,=:PB-2R2 =T6$AT%K),TT[P3ZH;78Q=VXS
P3XQ.WPH*(;\Q7S\EF20>;B\[7$?G%9@3Y5;PWD0SKAC:0"&?B,^P"WV+L-)QC:>>
P]E4VYE_X-:O/^!8NUV!=L*GBD#K_( E'EART(_D])WL^U\""TS9VOVU#%T5*"$7'
P'D=L4PI=;6(0<$?5C<"XBBQ+V1EC4RPG1BT\(#91E9DG=#MD^%T7*NNID-PEM^HM
P;QB)- $R%2#U=\FF<7G8+6OYZX&3YV..>2I1II?'N_VLW6^DY8@*^!AN-@A)F?O%
P$J")G)A&&*]A+#DWF.<83%;-:50/S3OFZ3MS911[LI6@_JD :&HE!5'%-SB1];K8
POM^S53Z4+D[76)33LSM5[2[[YM;(?^-/IWDH08.>AZQ3&0MR3^XGYLMY$7YZ>*<O
PSCA6'>E9$L>C"'4-/\/)*4D*O^]6[0FV]GL&5R+HNE"*VF.2 ;@RJ2_JV>J N^P!
P;?(!&'&_Z!W#/VY(\(%N,<$2(&YN_@2$?EIR_Z%#W" !$?!_7&2F[7.;.?CZ:%08
P0O]"T+JE?RKV[/6S"L?R_+':L5/8-=/H(#EW?8*-$QR"&JN@!P*DA'PL21K-E62S
P]CPCI$<F%><[;Y",B]-?9Y_1IW RJ(SDW2(K6?Z?O[W@&F@C^B_H@&7(,63@3)_:
PU$U9;.9EF5WT2_];RM"#*:IBC; ;X[8GQ]/%XDB8JP,T120PHE8R3"(&QKNII;GJ
PM5X+2CR9-O>:G)QX<@$C[YW^*\),-15OV)&,I;U;9E/;_>O5,/+$ZQY7;I=R/=A$
P@J&4I7==%8+O/?)J+4DF'Z$BY5&#;(2'O&]>]N2!PG SG1VTLOX\_^O%L9T5W+1V
P'CB]P3U.%60& ]CMQ-NEJM=-YM6<;)N@C3\LW)U/AVB,JVU#\]W?(W$;%E3*IF["
PDDDCP%MU8K\5WL%Z(!TN1NLHE!J;V'A1LS%U8X%93,E&2>JUM+N3##(*#C=6S78"
PU4$E1?$OUQ$N./(QW/A\R3Y3? \^4=2NI9APLRN=#5/<%("$/H8RA9\9TDBKO<O(
P,':1ZUCC?E))";FZ12J)OL?C%I;%W(VDD\3&<Y<M3;37XN3S%'2YU9\0JH7?$ .C
P7^_JNRRJ0NJ:L#4 ^!K^P&/-"=K"H;T^0G2, UOW@0;X*639-\%B$G0XCYLOQ#V%
PY=;>5*/CD2[@)%4SL+@WW"K4M5ZF:,BG&&)\I 6"ER3983,]OVTP3O87;662_1"-
PJJ&%CC3_T.ATS DN^;=9@R5\C]Z//.0A=[<B^#=O'E*);(9OMJ5+]8PZ7<NKT,"D
PXDX3V"='8@6%Y5R\85?2[[SIU)I&2 ;"Z)L9MJQN->@]/21$AS-8+L,/[&KH<>K3
P#G8^JN?J'5SA3TK9ILF?=%+;5Z6+V'B,51CC?*MG>4-[#_OF>KM7EO>/6$SWM@99
PE@%*\U0H=O@=OSP[-O['>+PPB$,:3EQ(WJ?H%W/T=8]LET:(];[ 6#A:=[_,M]@M
PP-2ZYOH7ZHGQOX(>**'#S!@'":U;^4ER!V^^3V[8I2#&1\-Y'QFG,M(4(1G><U4K
PKQ/SQ240N2S+<OUA/ML=(PLYL.T2FA*:\Q-7*"(CGR6G$X4Y+G.*6Z3P:OQ75I+_
P+B/S!Q$N88L7[7V5A7^R6'KM_W5;79R.--5"3*P\FTD4^JLZ'3_\8[WQH6KUCJ?L
PG9XNQL9(@JHV()=6!RZ>6T:!#-Y$@^1/,IC*C)4GJ=A\+$SVMQ,>FDBCJ 1I(DPO
PF@H+CIKL0UH_CJO#AS?9VSU=C^N5$!&9[AF(/ @2/(D*T_VU O/(I%6T95_D>GXS
P2_T5XB I[P-4%-6*_NJ9$IKB@A7#W%X-$B50ZHL9%MM@?!+I0A07^@;#S(KV!B]Q
P:T$W\!_?8-[6(ZLE' )<J_?8=9!Z(L8G_J#12@*[MRA=YP[ZL7ZQ:4JFGNJS;QD7
PUS#Z*:IKHM 1.51 647NO],/;(6S<U>ZTMQ6C'+#C%<$=K0,.RT0X%QJ"<')(S,?
PLBFNZ$(PSOUZ:5+OAG^ !6]<.A?=^39-?5%H3H9\;$HL)<D+RH.77DA.T%#5SE_A
P9(>XNU[TU";HPR]62$,TA,+OM533Z#!^>_#M!P.- NC$6F=$G+EM=L,\.!6%H(>$
P!GQF)JF^,L"GG*'"HY8OR=+5P^:ZT7J4EJ^L;E,4K5+N>OC@3IDI7N_=W)\%@IE+
PU2@/B(N,2G^]PQ]5WBF1L8R3/QU:/HSQX-A^RT(SABA-)Q)=X*#<7JN[0#?U+G"9
P$1QUM?Z=VI2/9V#H<XSWJRQ)<2\7 J*/&(7Z'/]VSA.1(&R^KV&D,+A>A".^HM=K
PHBY&5I:X!!,04_,I]8;(L9N3[]M_.]&=5G]CLLF6GB$[(?]/=(8TE\]6=\W"&I9W
P.F?4I2 J+A9?.$*)0K&AA-IYAF>6T;/ GGB"7#_[<B&,2D>.AWWC4LOL#=(:KZ)G
P\_*5LZ]S>2Q]_SST#7WAM[//=6ZU8)"(;(BP_G=%<P,>6;P^^#$&JSE2^MH!U!?\
P2>'/9,-'UKC/"&7L)<R%E_Y' \-1BVYS#M"7O.)YT&7;IV\;D)85)IO82W-EA=R=
PFVSJG,\XU2T)\9]XQZS>FRZ)!^X1U%.)STE;S)7G07XR[Q'M?<!@(XED.$%<4V7(
P%Q&Z\H/ZR;U#%8S[,.F!WORQ&.E<O("@Q22%<7]C'%QA4_[N&A_:6W])+LX] 0QW
P!2'5= -#;BLR*]YD&JE]MHPQY,YWJ>YK$KWL :8UYO6,\9^ER0O+MG<F29RT&B./
P)IEC\_!E5BZPYB5>L -F;8;.-+Y?7C CP//MHTZ*]!R!?#*\1B"*..-J&F9,B&Z+
PEXS<N4*!C\1!VBW%ZS+$U><3=>.]U(I.Y-BJE947$.>FZR&)EA.NR)9SJI_O9V2-
PW<%LA6#$O#K@_57=$;5;;YB&M%V<O2,0R==U33[L5SV7U)/ F+O64A]S)9EE*3MF
PH"%#0^KUV83]Q*3Z^&YSK8XJGQ'"0'+Z"MSZWC6]DTS*57YF/V70H%J; (0:S: >
PW"/&U:O[T#%Q0_^.]?.BU)HA,0S\>(7\81,J(0-^&_& WX=0']"JSGR0=WS?L-R/
P\6MD\7 8D),"M%2\.,.0H*E".M,6>=SB\9.&IRLBLM3.+<>IS3JF#ZL@TD)\S)/U
P7!#\@D]$46, ZH2LE+6;U(G9?ADC+H&,.D\1:>LGFQTJQ[1[[M,-B$3:&FTU%-BV
PCCN$UR@#<4*;;;54*O,Z,U.@!(PS;^M]-&X$R"I\XOQ(KF7BZ;EU*+WW_OUGZEF-
PG/[,=UZG!.^20G!KTC<^MB@4R6S(A_ FQTHC  G9P)R+!D9<S)'Z-5'7](FL8]0M
PCQCHFE8@Y\+YP %,"]]ISKSR5'?O4!5*F-R79<I6S#+E=SA]< U&1I*--HQ4/7H0
P5+2,]_4LKXGCW81C5&UCM;SG"O2_8DRN!M:BL2CQ/A]<)Q.#L.H3"U,QV6;>'%W]
P])"S%FN:4PLY*KO=+U]9KTY;K[]_S:.;B94/8@)D;X!S.U]:@048<MIE4&9U$(8.
P55OX(A<YB@9D,K8S_Z'<D37-F05\,S*=+6NK=U@])U=,7.:5&&S3)4VHUSB\WG"Z
P$5GA=W.0QT ?JO)X6I%9\IB$KTRMDV41@ <:;MS$_P2T9.$#I?, EPK\A:4_H['O
P3!V_]JL/$V@:WA4X^E+:Q[U]1V!7G)GB(QZETP1T!;+N^UIFI2MZ*LFBO:<<@_N5
P.[L7_&343NX: B"TD&84\FK(BX\&_.:E"[4=3;&<3:#WLW2+SRTLS-#KBB)5(8K=
PF8O=JF[+UE^T9J&.+HR,:>R\6PR-#^^;H4H95J((B!KC3RQ;ZK(GOAH%D2#"3%4:
P(1(1A'_\WY%BBJCRKL)4\-]<!ACK@2Y^@$%11Z==7NEU?/^,778W_L&"K<$.+)#-
PLW@@04+D-R+: <>:[<0J T^%U1:E9V<OPS&B@^[7!R1=+-/6N,C Z2G#>Q>5'O_]
P-U?&C>P-+CMXR[@BAN'T,&2%9T$:^7A;$/RXY[NJ^"W2H0'KJ!NC=="PLK#*(=\Y
PT4BKG^"JCF,#F:T1^,Q ',SGM_MM=M9E1RM)UYQ>,37#TB!O=6[%8$PU!0\N"0)W
PHMG61UHB'9 SA?K3*'.N<YQ.Z%\\:LFW,$BH8\^10%+O= +XGF20?F$Y.F6%07_/
P)YKC45B8.SY48=1*IP)39?N:[#3T/6C!]464WNI1<-[7EQ;C]^2B^3_)"H%W$63@
P*,&?3VP.:?E*T*6GG84,FNP$D(3.\UYD.+XI5&F!QLB709!G._ L^!-NMT(')H#$
P1%LP_C"*H/*[JQL&")2?<_K#2:P"(B%.DM^W&.Z+6\EV&19MXT&C-4]#\#$-\.59
P43FR<>$'>V=>TYSKICE#,^4KZP_]PAUN=4U?-QM*R,3_) G6\.9SO=03&"H"-^C9
P=R]!;^DU#-R5+7R"JXN8\8C3"TD=,Z0*WMY+$*YA;+!\M<"G#H7Z5MEI)&VE^@4%
P"QE*#'T_EN_\?Z >XLR85UI@1VD:^$)E5T&Y?P^U8LD^%$J1E]4#K2S@/.),;6C.
P 'W>""IQCW,1Y\M:#.*=C.)%!% C!U'- K*?E2V$:L!"5C _'>+!%M7:GRYX9?=+
P!6O+=_$UE(UPJC;;@A]Y\Z=P^&NIBIX Z!>M5U8S5,M03T='SSY3!!96B@K!]>I 
P7\YF(?';I9OC4ER]@/HHX1\F3#M,COM8[=OPFFAF,-<Y]*MGI0HT,[?9M/+@YX\_
PJ[JD.D.C%NTT$KP3^B$R$#@+ZMNS[;@A+RN\&*2L"MX/^I/WTG!5-'M"[.S_O!-O
PI%MJ)M*QDA>9F898';K?9.$/!;(&:E:T^X%.9TOE^*3/TV<KB4_,?VF&L3NW?C:+
P>J<&S@W0"FQ[Q@WLU833\!Q3WE:P-,.98$6/[9)# )&>5$(+$B*YN=F7R!N>;_<A
P"@O29+,A?B*Q+G:\GV9,XA<JE9+<C$(ZX(UD<8!).B:+(@DC,)M" ),2X-K<O#S;
PDTXSO-=R3.LZY;_HLDBU+BC;WD6L^<12C/2IY[]-9UJ$;N?;SLG_X<A#<P\?&Q<W
P$0L\$612DB; QGG!0QPWW(,9>@1:'C'G33UC/$1+?(C]_B9BK7++9[GO(A*N-<K+
P3#;Y3J<>X?5-2M^SD%Y&EML$P"!5.B^I8GIH<<K)WU\TT// &;21,G=+WB9',G/'
P[<16XN4OD$38=L=K68G#9W?GKW]96./*8AC]%MJOT0CX)JEN@(M!I<K%,6AZT8] 
PKK5'*/$'72AS(B.PAZN&/&L&"5I3&%R-LKJMXAQ,\K@]!<3 WR#LWSX-LUQD*R9=
P]-A$F[&,5) B;L0T^,D$1WL>83VL<'. !8)0VYPU$P+(IZ$7<]KD1M[4RRP)\(KN
P\HYJ;13,NM6N&;AXV7/Z<[P,G9/RNQX$A?+TO/ABA F0(O/WV?3H+8^$H!/6DT^U
P,@XU976OVBV5'_*QE55)UZ[*B!@YV)AMI5PX[,VQ'"3M%:ZKP.8+]D6>2&'YI0-\
PV(-T";ND7ZE59V@T1N<P%[E&)5;0<0V6V*7K!TS0)0SY777;0(P)5M]PT"B>Q980
P0*:!T%ALH.NH-/4 %/C?-5R6T,H  JM[QS:G$G2,V;9[GV%$Y,UBGX$U7.&*ABS3
P/,2*I'X;@XU.C@7OL%.L60_XZX'0PY]'>#+]:.+21]G*+N!?OS9U&&N0A?X#Q"F]
P_NI)NR,?L5V[1?J'Z9JLM2<S?,S;-F4XP?3@=/[%'>@:>TL].J+,._>O4PQ*#Z K
PY08I@;(9&!LYJZ* %O,\F4R6)B,X?Y0<BK$;/)I\@ZH/SB29I4N='9IPOYARNB4^
PGMU4D/@X?*I"%S:VL'W*97CU:DT^D2G6OE3'>1 7NQ2 "XM+V)1L#7"^GX+B%@?U
PRV(&JXH'Z\G!%8UK<7[=0N"YM=NN.]X\HCA7=-QM>=?F74ON8/P?*+=OX&>+^*'(
PZ?KENQ@$L]$!.N#ML;&TH79H13R3A!G^ZNT[D=Z+9GS@I7P#_U1"/8A0NW ][?K\
PF2B@N.^QR(E+M'Z/:@7UUE_R0%N^%EP7-,2GPO&AYY4$_FF;SK\C327L<;^6CWSY
P]H5O%JAG)_<$M%L'O=+W$G#^/H+(@/?07CA<H'2O[34BFRJXLHFWNR8@Z_ XQO+,
P>'!E:BD"S G3BFP@EADR,"N(M=&*-D52-*LI9QA\$WSG\/'U!URM3%H6<LK1:KIW
P1)ZHEQZ70"UH. 9<.BL5IE#H+>%C0^AD$V\6/\N>F_7U5%W/[\N#8#YW&4QO+9O_
P+Q]"[V/:1Q1+6H\#DE+T'_B+W85-C*4^BV9[$UN#XOZ>I>'04D(P$',.6=JFUK:%
PLUMQW6WY%]/%EW-A"+R5A8 M?P.U9-)/PPMS4W:1*T8FQ&O].79ZAIXP3P(ZW1HX
P= &4D) 4II6CQOQQA*'FYO8H/2' J"-"H/,V$D<MUC.;$,7\CI5_=(<5+AOK<&8G
PA2 'GZ5;3,#<,_;C:'M#T%/@<\:9N@>-"+H-^=5I.C>H3L\_%V'B31E/;-Z^23?A
P ^;>V+&L.4;9SQ>'TZ3E4XZ]-KLK+Y"_) (HLN)3/2R<UE=K/W+3ASF2P38<D1HP
P;$^]N28NV/>ID  **(NQ8S36YCNEK6+LQ'!"%5A$RN:0W'SR^6H9CG8)[[P39@3,
PLW[2M.V"#D[!^7"IHHDS3=5M@O9C5L3-EDJBVTV*RY3SWOSO$#&K(Y$08]0XC]VD
PL7Q%&>7T"B;X,"RA1!'XU]2QX.<YO5YF:.RI?E;3E!VV\@S5O<R MC+2T@#;-#WN
PMD<$L6%:,4^MF6\VH\D9.0@B3:VI^1HP]"77ZG:^46P8I>KYB.IZRR8VK-O:LZ+$
PP+N./J>-[^W^3Q[H5#.,T/,M,]U*G-FG.E2$=SQ1Q+;/[=DN.R!/]XPK',5+UZZ0
P6\$Z]!H%\ZJFL9DW];CO>L1FJF0DYXA]O$'4E&H[.:^^V(+!#J2E9!]TD^#VO5 ,
P<CUO$J&Y=_P0S;!O1[.E&B\1"*ZL/]8*H]([BT/#E%6K7$M1.-"$EDB;28%K!I A
PFU5OA@YP)8YE((B3W_)N.X8AH#KP)1-T#1L9>H/V[8\U1DNB\)F64%DD5&/P?K8V
PRT9<YRE92:C[1B[W2*>9MX+$WHQK"3B+Q(.HO20N#\A::9-,I:%_[S^<24-B84HB
P=#CZ>80K@T-I/I,,8V>RCY9#P(.$65&U,OV0%#0:(9XS%8=W&#B^3OX*T?YH6<A/
PNUTF?<@8+,&W(2DW^/[3V+<FWG;*)36'-4[G9CUZ1#$9WI/+24FN'D#)T>X)V+&@
PI*CUT\#D@^R!*DGTOOM4:S=_":KI)@"+L^TH>2=*R9=X0R_=)5QSY')LAH?42%$^
P]7^+(BXMWU-F!6GT*;>6#Z:PK%FG/+6OMBT"?Q#+1B1QJM^UYH(D7D#L8$GH>L;S
PC>!C5HJQW$KP<!K;4\6!BP/%6[-]LB[YDT:J4[Z$=!OFM?7)U< @RAS.T-WN%K!<
P0<BXCD _PH.$/BZG=[^,%)4X+E<BO,[=7=%V@9S<EXK0,0@K#/L'+2BAQOUKS$G<
P28N8<V[( (]$(%AI1]81^SPXBD1![57;<^1UI*$Z<L3JK#M+N62+T7_7]B&7M-J&
P9P=-5Y^0/6+V1.G4FHSZ#(,,61,\)OHH52J2;(CJ0"T6O/<ILN/)01[%_7TW*6DO
P7?SL0E1UJH]@S#&KPB:I+=1X^C+]RKEQ2F1@H-?9-E^JP0!/P!6;U57"4BDCZPV8
P.ZCDK?C+LJ 59/%<FR61DXWD5@--^C^Y\/,#"10#BEU=<$'JG00UNXG7#*.,HYIS
P,W%>%S%D8631VF+*A&?>-+>8"-O/\]0("ND*M*)EI@LT&>50]%H=5GK?C='0V'0/
PK=&TQICR1=L!6CVKR<LQ='\42HA=Q&A>, +8VMRC+8(LLQQU7J>V.!([$OUPDCB6
PBXN7RQC4Z.=$K3-.6:*'.R!)A#PK!EL59;Z"[M)V& H?D/>"Y(0;S(0YDPJQ9V'O
P"ITOU48%H$*BQ"H!F!<_H;(&9[L9< Y;NG* (X/"1NVQ&:GJTEWE%G)K"B^XB8=>
PU0F)5==&M5[U#>$R4EW@F<ZOPR 9S^HMR Y % NF0 =E\VCG=LY4T!P$7&'5!&G-
P&?ZT:+NMGT46#%7@%RG<0](G.+7*9DQCMVUOCL%#KVW>YQFX&S?;6/_*"D"X[E9]
PZ03:"&I?9S!"]@]RM3LNG7J$8KKZ$@D\Y':O?FHW].D_6<8 JN$0VQ>2-Q22W;]7
P8YTJ"OVU "L\&1T8\.:H;DV0@0$O'9I$[7! *ZO(J=A_ D2X&[KN;RJ3.YN&A2O5
P:I/ 8N\NH1!D/Z Y W]MHI6PEXU E'\O[QVM&UN,@!&,(NAR?JPU-P3#^2,)G"@)
P/I P_DU9\5[7S]"5T$<&AZ?TY%GB/=&_,=R]=O:\HX:'+H/7I ]6Y]DJ^D 0CH,@
PG7G#<,<I'F3\TV?&L($@J52]3)@TKG@@0]3Q$_U]5<T9$>^IVH_.HTL_31Z!<7AW
P^L,S,CM%6K4=D +M4:&R[Z]TOSDY38'VEQH6K2RGB FB;O:CS5X,3;Y#!#KQAX6A
PCXE>]T7,SF1%/7,XDU%Z'OEKP7<8&4%<_'AP?=T!V5Z4MSKBW$\D2-7=BK7(ZW%;
P]FB(@'5N)*T%W;1'1W."#$^%(U$?:O)G/.'OIV?D!:,4"=7FFT1P=@KQ\PD!;7BI
PJ!Q+0':\+GI8& #TO?=:/5,/"HA2D8"=)L:$L8UC\#8$;<R8:?K99-TFD4ET:L$S
P$AZQ6?;'V==UUOOCO) ]&5'!59L QS0&A_,2-=NS>)% FTT=N 6*?<G&:\*L9; ^
PL6VO   1V>;&:O1T84S,+7=E8R"W!%U%'+&\N@,OS#:-ND(1SR,+/;$6#9P[H@$-
PG(IZ%J3HG3CV"FI:<Z0O+C%9+/E'[>?MPBP-/PUD4N\8 M(1=^?Q/  X-2;">_.1
PB9W?%=MR:+=/6 /HO^R_T:Y&]B<9\%R,<'KR(,#D-P'PAB??^N(3-FSR"+MJ!I]9
PE- FC[7.&\4_7L4WJ=(X#UM'OEF-$C&UT4'G1NC:'90JK( <N%F2]+_I+&YA4%4\
P_G26<6\_\Z1K4+A')5CG6]!QB>'BYH8]L<)1/[HF7%??2(KL5JN\MG5J5*BYO434
PGU93MR+JG;X"<9023$;8BJ1=EG#9==JQ%R/)"HU&Z'"GS21\Q\=%I]?$5S9H/S2O
P2Z&"=F%/*<-:.\E]Q2>Z4%C*RA]?CGJURU9Z=)8Y)/S1=G>1<RC$9LPLO,;^-X_6
P(40+^E348B15JZ EA(*X""@N%7LLB ;_JN%4+WMHH8#HY S A$DO!E(8O68N*0S<
P<T[P3,+#B^P"2-T@0O%A3HGUF&]29O)U4AB(?"7T<B&!=5G4/M>6'+ID?0F.5D5+
P,(R3E5H"&,'=[GBDU-N!FH<K2N <+;;;+81>OJ=_))W??+HY<HZST?]'?BQS,=FI
P!2]$G[K"5#KDS=R0;F&8$;IO %@O1Y<P<]2"P^-2>L/L1/=Y<]\QPUBZ624!/%L)
P<P4OGZ4"+>-1I>O:#[^J?((LT\_4C\VO#$]'[EM^6<&12/I@5IG0">&C>-WDAEAX
P3LXOW(N0$NY&POB)=K15KHXR9<%\FN<B(=U:C2##0%+7R3(]B->82T<$_.!7D46\
PFT7_=-%ED@[",<;+*9DA+PH9(4P57BPRP-0VH,_C=G'GT@YM%4""?@+1B)^@/UGA
P?7/Y(C(07QWUX;X&OYU6X+>YP.N"PU<@#/\%EKCLM[WW#7%E3;'K2]EVD =^!>^<
PTW0H*:ZW%3<8D9;SZ552[0<0]>!]H)FBAFF<6BJ;OM)5@A#^*A$*KLV"^GS:4"02
P>:Z-<S>)S'0*/R7Z:?.E<J@9*U2K^'*9D6:'XH"*PQC$D6')[]W*AR/XH@!P-W";
P@T+T#PWQ%8*)>/)&%ADFX<[2NUV\4F?D2)S21SE])J(&.1?OSJFY65].M@OHK213
PT5#H *3N?T8T+OW4I./\((CSGZ?7Z^W>E(G[N>C*0W7&_[ZL_3-&.F*9BDM;-\]1
P CDY^8;\,7@+;1#R=#66&AC!D;([6$-8BK;^X'Q#?:IDW\GEUK8L_P/S&57C<.N8
P59>XMI?]?;34J-<S473U^.1\<M2*=ZLCS)[Q7KW_9]+,E;F<M;EJ]AD@:/VR3%U[
P(FF]6G&\WCC.!F >B:_970>1S:U=4()EE;#2$1A%E)-H<)J<0Y6T;-7KP;NZ+_TF
PF"Y(-"2%WTR3K^VV"=&YM8H&ER:P>49E?BR$Z9H=^:AQ0HJEM*!=6"K@=+ZL)<JY
P7&%YN?]?@IB_S(LP4&J@&X98^8_=X/E1KA&[$;S)81P(^%IUQG5E7WL1*Z1Q9N5.
PZ8R\ L8S7 "C8Z9R@5P&4U/Z>=J+^NIZXC<"7)93@9X8T>[F^M9%CZ6,'GS/4CR<
P>'R9$UE4:&2I&C6"UR8"N(PWI"EK$ZLL/&?**27WD0[[B/#H/N1/'UO,-I3*W?T"
P**KD=*UARB>B-7\EOA=JL;H"H<U+8.ZG#$"15X\HO,U_SX!<4TO2IK\+\XO:O3V<
P0.E%3<9!-(Y7/]0V4F:[ZT)'-B=4)00)WDM_S!G)ZYECB-$]\+LU8*?!KH^A-016
P,K[<,24#/%!]Q.7+F1]WS?6YI10*KYKJ%0;F].L#$6(A\1R\L_'@DLP?,RW/ +>Q
P3C,R\X]I@+9EC.F_GCUA+]9BYO<1W\6<M6VG<VI4V#\A%Q'(Y@8>WP0_[#Y@-,ST
PFRD2E: @1JT-?D=FZ?(X@0F U1>%?:[ D97M-R<31!Q'OIZ*$$;*_3::Q&S3RZI.
P@#V:Y*TKHR@Q.!S*PP:X1D;]C>^Y1GO90$+.BM-P463+K813!CW7N*\03XYAS&@1
PX7+H(@IC(39>%LKR.\BS\?B8WDB)D-M4_1C@P,9K'%\1AXR&*RM$8="_2)R2]:]O
PEM7*7QG.HI;3Z3,[ZZVB%QM]R]!II%6]H;>S,(B04<?J:"&*I -%C&H15\$ZC%5_
PMLXAZC?/002#Z@"/G.OX3<U/.WI@&CDFCZ\ W $&APKW_AC-'4Q>?N)A&>8>\Q)^
PAB-\+ARX.8MJTO+Y,2Z%7 Z.;VQ5)8_[+C2DQJ'DF"CRWHE[-LES!W2[?&9?"DK2
P9O;73ST>E)1;_IR]QB!BPVG^;)(3(+M-X42=&H[^Q $&PO4IPJ&1#2Y^7D:[:TMD
PE1F/OMM?)S/G#+%) O@;\['#6?WF1"XG_9=5&.:0BFZ=B;LD("X0"X&/Q71)W(><
P@^L1\NET\Q7=4P#QC2>0?Q/"6>FE3:E5K2N/3,*,*@#:$P>&#Q*/V'AO&=ALDIP<
PSR'W/%H$A>3+Q?$P:J(2C]S"A$G$964#^-!AZZG'SW_P"7)P<&T7WP@(!7!JZV'&
PHFRI"=:O&@<.9592Z#AE^#@52= ^U'\J$$1;K-A611HD(N.^4+>8#.E@.^ND6<&^
PY"5S+1"=;E*CDK%+GHG!]\\I(<ZMN<KN0@>=8$%2'N\(6UWE[D&3)*'70433HUK"
P3NPLPR\#^UI/OU$T\92R!'-V740U6=& Q6'B4<\$!4$'2>^IC$HX]6\YCR.X>5/T
PEQ93(532HXFAO2<./:[;?Q0)3.W45=YGC2B$#WHTP/>LP6$D/5"B!7-8!_+PC/S(
P P[;9('U!G6>V*0>(&A<^E8]BM1Q2PWHFA11_;JO7S(*=[Q^AZH!SES*_\QN) I,
P\+02:Z#Z&<HS6.+_\U_,F6EM!(CRK<]"#3,J4]]E;DY4#=C.Y:69^:XE=GG\ 5P 
P4^?-$&/X&C"ZRA_N!;GMS0C\YK59N0L/&?@: VOV*.1L2Z^"RQ=_2=MH1A:5T:EJ
P#]6I%,K5G)M <2?'!%(CJGR1.^A("+7[7Q#@/ZI?A92T'1=?(N80N.H/#W03LJ+K
P;TT5"$5V!.^4GZ) 'G?V1-30K]+O7R :HTP?JB)8+YTZ0R/F9ALHU'&=_7U&K5?W
P/FR?\).%TB= R9\J&W\T%VUY_@NGWC.N[_%!H!D*NZ"C^D#=1;2G[@L%UWL%Y%F*
P,68%P@/6OXVK+F&JB,KWD^F%%D&/@P!E#*!V([JIGQ.SUM,$^?[/'DT^.+!=(:0!
PBVB$G7VE40*FA87D!;*Y\Y=F3:*!Z(DJ;W=V6\0J7*+5!-QS;4*X^?)J$5>98UUE
PTU9G%!9D?5?M58EMNN+4AUMNR4%X)K"TLH>S+XA_X2V\K$P@)@T^O&TEU][\X*=.
PW*9<\V"9O$ ?D@OR973Z_?$R7?;"&V9L*J$E!6<4,EA=0C,I3QG+B("=6CL+2ZHS
PQO#8!9(XPV0-[_.B/@[HD3XYY*^E+))IG?!$.6VUO1\UV*BJF,Y\?JHM!TA7 _1I
PD;?SQX@M--B%V^JG[9GM.QP45H_/7T9.MS0FFJ_ZN=EC?W>PYW<H1L[NQW!/0H*(
P?*=/89YG'WLPZ%B30VRNX]F?%C&(YM+%7/R?O618AK)S$1J.5('EZ1;!-%,G!IPY
P,LOSA;U)VM<L91C7G+5X]TD]9'BSZW$5'<&SO*P,IF<J@IUI'ZUG7-_4)$9F FU]
P$'R2;GC.Y=2-%MHG5)XP&\JVE>>>P5P^,NUYT5F(QHS"+/9G3/O_B%DITM7[A[M,
P]#8"A(BK9/:88K:?M. &W]B6^%7443I?0\O9<BR28O.O"7T$I)-$ PT9?"&=_H6 
P%L8J<@B.@MEZVVU>'YZO3-';^,T"",2?P8\6*?EV!\9G^=N B%9KO%.1VO&9]YZ=
P?RYL^B\"T5!3@$WND_>M9*:,6- B@&:UBL#;W# 0DTQ@-<K:0:UL]XER8SA:2N"Q
PL;I6D)-8#K6$P3,)@4-%K1*C",CMH/-#RZ?MQA D"]+(12[H"-= OX2PQ I97_81
PRTS':09??<Q"G9E^<E0W>AAW%2<)C@I)"&#]F2 I/,7=24$1><@.//+8!H[W[5.Y
P1@_#+_R!+_6$<R,UWQ$HY9AIR\D,(MQ'>96B/OR*'.L(IQ-[%XI4-Z)^__<I]'S5
P>D8'>'=+F6H"9 !T6KY]HKN)T,?#BY2>>I1@Y HD9_J2Q%?[K[E<[>O+T^OWZ"HL
P%R=><$8O2QLV .BZ!3%N'R/\<MY-::C71%1*K:ISG!QE,YO'R;IY0CN_!M;ONG&*
P'VQ:U2DKVG2I0WMV#B*:LS_VN)?G[%>:6#L%IZV6&\H^C"QV"+YIYYF9&X<B9)*M
P0I<?6H-):-15A[2EODQRNUY"E6$>QI"8JG%D$LNL?,"=EH"5T4R&M&^YMY*<# R7
PTO2T:G>X&2_8A8\9E<ME^:YY5!Q.C705/J4CG8XN,W#=,?I]N&H4S2P-86)@1TH#
PU")G/GW:&[>9(Z1">#GTV3Q8=NXP!P1F$!1.6@&*K+PZHQ\0H+-!6!/VX&S33CL9
P148?W)@W3%Z<2S3MEU^,64O'1X)+1MY5P.UQAX?NSGO2&%]\8/] 4JB9V4>)">$/
P@\[<?(H(E9ZA1K?GUFJ^^2@X"I,TEBZ_>*1U!+-0@/21!/3B0!K!)O&^=$Z;.PX 
PH*^.VB/.\F:%1A9#G6D>T^%$%AV]G.-Q6T$1SP ;]><MM:3'2)VQ@$#<LV*:(5GD
P\"5D)F\=TZ(&X\+L-TNCCYVNT4.*COYMPOU"C^KF62_/U:-?YKK OI:+H'!-'.M)
PQKW88J?[G_R:-\G65O *JUE0Q:PAP-BFR-SMBMS5"*L!@IGZ>X?#470(KI  N)"^
P%0D#L81X-N5]QJ-9F?HZWX=Q7W.%>#7(U]3O"+@3X3#8Q+UXS1P&NHR@$F9,!9AD
PF>_(.^>$,[\.3RA9N.I=-$I/%30HVX860:4:LL+>2=E,EI> 40+NP!I+.I[1F8+ 
PU?:/^FP4!':\ELJU](:<%U;[NB(-^[84B.E! ZQ"*+[7XBD4BYHTPS63/YZ@:2VP
P-P*Y]%.&Z^AX5[31%)#QK_<XGI'4T*[=1T,Z8*]/&+>+3UZ<4'P7^3LRD3CCZMS=
P8M\*VM&49O,3W4D#08@B\78Z([('QJ Z!LRY2EDQ%@DR6D9MF%"EGKM$K9[^4&;A
PF\\66<<$ IA)>*>#+?2A7-(90P*Q%)K QR:M3K,#%Y_6A-\,W(VTOR0QDA^!#G2I
P'(S2'=TP3)SQ52YVQ:+Z)@ B5SI*!@^%:S(TB4]6E,@<9F,FTJ>;05R@UXLOK]/^
PMF?MB[:IU45$O*SE5?B@@)6IDPKMZYVKY!DXC=@H+14:=3M6P1CD7X=OLG*1SY7)
P%FZ.W.U8=[D_1S?QBU"+#8\DMS^CJC,-:A7R)W2]#C+_T7&4LR3WA[9>GN8S<!(/
PU/M-05/_N1ZW;N'3><^ #RUPV78:16$4;T;\*T96)=NB]P@?I)PE&5/JN:F@RBQQ
P.]$G?B9&&8W5A[C'T AV6"5.YKD^^J)I7!ZSID8B*Z(DL>2$5KU;^9UT-@'?;6BU
P6R30J+K$[%.RV:)#/V_B)!06 /((OHE#&#,@TM $49$"8!)=$3>,P7)+]PN G<]]
PC8EDY !$WF6!PJ*,(Z$['4(9=Q+CRY662M $_H!?LV4!@]<CSWG2#2<N_6/,* I,
P%PE3YOK/52(0L#O7D;\L7E\ZN1<@9,**A)50MJW<F,992'+XQ\J.!\BWH:0SI,1_
PD\0(2]?C9&Q;DWS+G9[I.BW' >#O"MG;.M0)Y-QO0_*PMC9$M8[ !$#T='9OD 1&
P%WI@>O@=,@9)A1;[Z& ++,U+K1)L5. L#0-+2K.8'(JZE L?3;D2+N#?\L/B,M?(
P0]B4/<9N)ZU@MSP^*; IL[3W!^YM$LPS0!4["JHR9,O=83TU**R6ZD+>JL!#<DD6
P'UKZX)>'7O5_2(*\=SLK[IB#.(J*9 PAJ9M80]BO7^^)D%C,Y-8)$X#ULT>\WT!!
P>'%$A\;8/19HOO:EN80<T&X2\%$.XD5W>NR(>9_&18&\)\Q[&%W'>U(*+R;!8/ID
P;XF5P6H'X:R45.@=XLB:]CG!P^D:^IY]P\WS(/4,T[HD[ "N!$^)8D*G'ROCJ'TX
P7.^D_ TY"G=I:73\%+2F\MX)T0[KAWK4V8PU]N4YLI7/Q[7#Z\Q((*X>DH(4JF5=
PW%/,5I\P3+PM>@\V(M,7+I>*.9G[PVRD19@'<]G/ME1ZSF:7Z0D^B55=J9AR8CO)
PMX&(4?B0%)T>@320$^V@(E%^N&FU8P"OB=Q^@D>YY<"H6G1GK#^/>C(9H+U,T9M$
P)6HBOT! J1N^ VN3N=>*^U/#&_:*E ^MLG6-1BD<\#!PH&P$K 7?_GR[.;BSV5'(
P\1=6Q,N>VN;30#$'[XG Z% :O%*VL9,5!J?JKH:2I3B*H0)[CVHL1@8;;/'@6,E[
P2PD[NFP7X6^R*7WJURUDMQSS16B#Y$:)WQ?AV"SUT8NI+8,JJP"3(RQL)G<^H]$=
P= EZRYO)6:?GE#0$/U6VE$(X&6G0+'5 EH_OY^9V44:B!)!Q!O]%@>RH\]QGTP>_
PU\(Z[&5..<H:;]#@W]PXG;QC! M0>:#BZA+H2=R(=Q5%V1F+,MST Y@H[\A7A&(:
PQ: 2*'_4H(4G<)$94FESWI;.#]U0S$X#W$Q%4]H7,E.C)K-SE$HP2%P171XA'T;]
P'80N+VH,%*.[R1_@ =B-9 ;39VQ,& K[4/UCIRQ&#Q8BK$9_12H1>@ZA6+P1)(1@
PNS:GAJW:7;=#B0IJ\2%\I3#I_(\-2<,Z2KYGLCER@5KG28$&NHVGL=5QH(/--GTE
P-&H=!,XEY=Z^,-L:"CDY'!='#53,\PI5L=>34,'T44RM=]/TU-%EF!+^CZS9TOIS
P66\!$8.0 "0<T[N3^;L'M?0B;FYF/7\#&1 YEJ$;RIK,PHA *&$_FP:+:93SI:?L
P**Z@&*$UE6MB^K!NW5)"A(Q/(5(P]_1N_(R7E#\2ZZ'\=#]0O]Y_O)L]T2'LQUNM
PB^DQ9%:OF+3*@>A^7A.9(DQJ/653$]L)<M7+WR_E( :&@:YC\H+%U&<)B?Q0@Y9F
P_M0@'U7#YD#BKW!=K:^UQH1\SKH%^7\=3!"6!3783NT\,T7-@UDV<OTT'RU=2^0O
P(&:!0FH':&QUSF?URN\7AY;(4YJCLK6 &4YTLE:)2[276P5$34]LY 1GV5S>-Q K
P5&;//+M=7P"G\?A^C(RRL--,@2 8A\I4%VG7"[#4=V@-L_C$RT*00@/M>&>R]VG&
P7)9^T. \I> "FT2=5<M#/V[]#R]&%X6'^YECWJ:Q"A >0 ;CQ+TJHXQHO3*>R.][
PKUQVETG_<]"&<OXWJW:O'OI]L[PCN=8>)EM@&C;(?:.QN%F8@R#-N3=#-A U.2_(
P=WO^9?SP\;2 /ZII.0Q=<[6[-4GI2/&MT;F)Q9Q3%V-ERFVT[ >MR17(<E;A-BU0
PG0X<A<ME:H.F>>6D:[%CQZ!!ZRG=D9DAD#0Q,[*"'XB)Z0,OIM]23FI(2YPR0W]-
PB/3Q57=W&5]G="??L=I\3-4E;R(WL2C42_&5AFKIP,R5G<AG@QI:&I:X7W'U&Y,^
P6'@A\?1ZT':3N^)TEF%J[J=#0('L'"K5)GO-6L!1'+*4<T@K-<2P98(M*)P$T(A#
P*AZ&9M"&?<\^E9MK<EZN+* .[[-C(%T>(.<"356@\E'@27\2D*TE@6F:?I^'WRCK
PM'0JT!^QF=EWK+,JKOOL@)SK[91]I520)PA/D:>8[Y+NH'$C>$XHC\P8VN8J<L7 
P@%P?(3OI!W,=8:G8E9R0W_#]SZGIKVAYH-^TDKE,*O;280OJ=1<<4=I:7Z]-*S;L
PP;!'()J&EAUERUQLRAZ;()RF.RA1IU")<@GMDYYX/0L;R,QTYO,<8-H_B&/;W(OL
PVLY_+/*!.+X @YL_VZ2>MCH'VFO?*S?,CA*4-6&C^L9RYVK98/]EY1B AT,-*#X%
PNR7]/KSBU'O60!ZX)XB/>$]DUB@H4.:B@)PET\;<IB6WHW@MUCQ:4"RA+2$3VB;]
P^+ZN'<YD=.KV-)DZX''MM0E;L>"*9^*W?\T%0CE-DW%1#U;9NS.,<PA933.N^#NJ
P=BN.]+!6@/034W@ ^>P0,4^B'"& *.YL8@$B;--! FCIS7*[XQ!]TS7,:^YZBZ5;
PHQA4%/_O5QV\U130XH:^%R]:TWJQH: V#)J2R@E.I&!1Q(@R< FXQ@\[2#MVD,Z)
PFYI+(/V\ Y0WMRM0-![)"<LUZA?=_%UG!QZ[91/\,B1MK3.-8L9:N4>UO'M!2YP?
P7Q]B'\<!7'D-7T(QDFS-9&)(47$8Q5WS/^3<-8Z"F,9]F1S:9#:.EX[&/ACX[.GD
P$//G4=RL):"!,"X0&T7"[OJ!8TQ;Q5'S*]X4/N4N[(4M1686-/P"=%Y@(AARBE=Y
PA%?6Z;L;!!'F-W)BKD,C A^%@!43JK9:(-YN1E@_GR;YYZD-2ZVXB2D$U+JPK6%8
P L\];BE20P(N<2D =M33N N@F(\A=/44UTIUFZ#XJ'N<6?FP_4[_J45OY$W0CPM*
PM$W+!%THLJQ@/C<4#UN"SE+\,EZ@@YRN]I-TT#?)1'XUQW&;2[ E"*7 HDGB/=90
P2[5551EH ;B8-0?9A<4 10&1RS@Y:8M7?L(?;\0M,,>0/$17(6U5>0P#WJ=WA.GB
PF_$:36R&.8CMT"1 JJ(2L@H&SU#S*PW:L7/DW>1RE;V\MG<.">0S7A^Q0:BS![@6
P4.)'Z"BB0!JF_B\5B)A)GYJ=BP;3XV5B $B01?ITX)$XP]QLGUC!U.F8-$=>!<8I
PUGL:>:$HD0Z+6OGZOY;UJBAJX,;DP%$R,OY3],##DI,+!!LZS\:$6AY]TS?V-EGX
P18- W! (48@4#XB%2<SAX",^+974L^*[MQJ)N\*_&7L0Z"W.OHYVH]?BN<UIIV#Y
P6O;YIQ34Z/WIV_+T[*5\/,I4(;(CV,:&R$K"+219<'&6'. $%Y()QP\W)9D*Y0_M
PJ!N$AC$D/-S!-C,O4!:G(?B?$"R23[JE)@5D91BC.+BN>O:?%?MWKH@INA'R7@=5
P.%I!YH?K*'4^X6=UC/)'A2S/'RD,IH7.'>Y4'[/4PP'*WNA9"N[;4(5:85\T1O#_
P,O[13+&@R1DIC^IWS :;"+05XG3]NTT/99$9H2-;:H!&<1,LGOJ41CA6>[3YU6*;
PW\[>-]W9%#U6"\B\=W YH6KN]FK]3Q<.#G$8,*'^I-8\U:LJ_$PXIE='2)-ZR3K8
P,UKPM6!:+O]VIH?>"UDO+=%L#INBF:)I<&=6N/O3^88<F_IJ"_O2E)!2Z'>DQK'\
P&9G9?JAP]TD73&9[@9FJ(\:-EI>OS?EE^<SOH!D@P+%$='M"_CK)HO!@"Y)I98_L
P),4Q3[>U]]6\$X];.(:?)G$.!FMGSJ/PHXG2I#@6Q"A)%Q-*T75_38$TGY?LTK#1
P3E,@)TIVVC\7!W,0783!^VTR>#8L9!XYV7I!P_HN,DZ&=#R6RM T#:4H*7>P!3M"
P2>'N0;:N7WB8V'Z80[XK[BY*'WVIH<AGQ\!82#R[>&?B8D[APM+#N>":%47!Q ;[
P_5RT-88HK_:_O<W4H]'Q>H>ZL=E2IUOZ7ZWQ&E]7].U5X\K>ZU>GH4QR?'<%%LS'
P;Y4*+^:VW^BWUE-+ML!?+C.9$2=3P9OS,]D2E!KU1C#"D'@:XJ.Y[]_E[%SEH'::
P;ET90B-T\OUUBK12*H6JW+?=FWK86Z=! W)Q[77WY/'FT9"PE0M,H0I;GQ S%9IV
PJF3OG&;C4R0-2QM[8DNAQSPA#?<& /32.L2PX*X95OS^UZ-X3C,AJS2 41+)*]>,
P;&EZ*):@4+MY41,/1V:7R[P#6<_92A8EHM"7]]C7&ZSM"P60:XR ZHE0V!O?)):N
P,0OE+IM-\Y2@]#U*W#*]0 T"CU$7S#+"35C_O3@'8%0/Y!V]1'O-VCXPWEQ:GE1+
P(4;=RA@DI+?M)043C3FK/6=Q^-5F:#)^505%-0I<N&Z"K=GOP2<?&1HSNH)!=LK>
PS99,3R^.S!BO&Q0/ []WO2BQJ<$K-9:6)_A/F&R+P0,@Y3(ZG?]<J>.=:11>%50!
P4I)<C=CE&+)$E*AR>TH");3J<-X>I=!S:4RM630HW<6#_4;%I))0YY[%6BK1 R7P
P?P?.$!20-D7TQ/>! [M\,\B2T*%$TH3BY7Q=NK .$:IK_0KM:\\7D:+D!Y^/^G\C
P#-S>B(V()\6C$A3QLPAI=/BNX^U'!CV;%WXL^A<83=(?3P!P2 4-SD/6*0K >4N\
PRZ7$-&S8__-3&DEK4L76\8"2P_P@KAZ#"_.'RD0= ]Y+W!C#8M_C@1M0*BOFCC_-
PKBWOR4-.:[^PCD\]2KHDFK?L63I^PWTM&T(B2H*A\(G+].\/@,XS>[%0Y4)Z'-Y+
P52<N'U/6)UC!M<G^$%&%OYKX/%*PG9"5S"'E'X.(+,UJ<SM63!MU[@S3J0BV>+(K
P7."I$(.W,>^PQI$0W:Q/1,J+VT.:\;/G'U;&4N?__1]L"QL%'^!]D UVX''5$J9$
P<^D!T[,SBE%<I]<;]NM[<24+^'CAE**7C?187@CHR'1NK#6"CB<3K1"C=>^,<C)N
PX@L!-K+P[^K1A(]@"$_&ZK2EZ&)? VOQ >*M(S2X3$\:]1N.=+;<9U:BUS4'+%SS
P78K9'EQ$7CV$!4A,$)$:DA9VU4^5NZ1%#(D"P;)6X?N"ZQF-OE)$U:PRX.0@?2PZ
P.ML8YH=<XD<N*9O=5RZPG[SRA<+4(_;E%0\5(^;JG4!.2!&30=GYF&SW0%[>QTOV
PX+%049V!R$L;D^HHI;IOB0.X^V*"!VPA$"(7:A##,A%SU0'/1E !TBJEV:2.E>M-
P^&]-A,,<XE*@8J2\A-1SS8$NF2!T6C<\1/[)X!-]W0=3^X7O1&P+>4FK0JII4-5%
PH6 ["@!^8#MIY252(*RR=;QM;394[KM;$@+C@].\)->J5@#+)]@P:<PW?>U<EL S
P_(O*46Y3?W0(#Z=]63^HXKK'LI31/++GD@3^41WN7!&GX65#?:$GO'WBO\5C+!MD
PZCI.UBH;.HX^!(EM_7%@Y+T25G,F'Q)6RID)>H1?HS6"*V3W7<_DA%Q1EOAL51T,
P#8Y<*"^MS/,.,II/># WR]\P-#?F)77;\$@89/SP]BQ&)WQ":O76XWS;4.)1(=).
PSZE"<\TND_@WMD1C>3=#"<3KEO_!/,4)$HF.$R!Z,N@/D=]9$,+3.R(:@[$LL0]Z
PRM60N"^B4J"%T6H)FL--3VH2F4<#RG,VZ".'/-39RO$X:-VIR*O/FBXD13Z -I^K
P\$::$NE\QF,"ZNDGL7T96!730%STVL9R2-P](3^3-ES(38;LJW2D(E[XHK+X#\R;
PB]KK6G+0*%,.#CY$T?MXRW*6Q@<IA9BN[7QY"'"851R=-T;F,'R3XD]IM2W;"O^4
P270['Y>Q-[F-^TQHH/%V0HM&29IELYCF1F$SWCXN&5+_M5R V>G\_LAM)L$@+P64
P'57!H'/EEP;#\8G/GY([0^/F^L19WY9[3TWQO%N:4AXLD#4"K* >AVT 5FENY[>F
P9':IQ*: _\B=Z4(^I%TW.B=R^J#@(PMI1Z9DU>@ T[N+/0=@+2=#G7T=,W8W8,@!
P/$FSS?_ A))2P"]3 O6* (.PPH6#Q)FR)Q0Y<HB6.$U34NQ=IN/K/J#)UWDOL@:4
P/T<S,M*6@ZW83IIAZ;]9/C=Z8UBG5T1L!MUPA+<]J1/Q"X+C)IU^A8ONM_:55I@:
P1>'+&F-C^&\HK)0!+ZN#9:[*GJS;G49FY/6Q'U77K\P/E%![_I(A5SBZ>@ Z0]VY
P^GJJ8-(I3O9 T(M_6TQS&!AL<&254P.3H#\TC/WC$7@8_Q*>B'Y(&P"W PA%J[KO
P@;HQ*.(XX1MGS\/>X\%0R='!1/D*A[>T=F>TBT\WH7&.QVK>^OD[20GC^5FG%JYK
P;#?CT_T% _A*I)1(DX/,'4^'B%K%"9ZN@FJX9N3:F5ZQ.G@$R<G9G)XY!SDTYO J
P_3-.C!%U1.A7<V0?:),\F./1!# /RC5!@GXG;9.HOEY0"1\E\3YCJB2,(/9'YGO%
PZO2@^);9M<@]$D[<OHJTK,[N;EXGP+?L]+$G/EJ=ZV9"OQG<2S(&,D8YS$MG.? R
P#^T4'(H(W31"Q:$K\X-OQX0U&:?N4EXXV:WM2( &]O3JD5S&?8$T!)+N^&DGSI8*
P:-8A(%X<EBVI&F_ ]/&T(?$UD_#Z(A9!(L=;93"<2L"A*->?<[;^$B8--_8NL[E1
PX-7C"9/R_O]IKL)@8FE"R'ASC/E6%.S"U !M/8.\Z=%#,7%SDFI_6;E_&DMKE:SZ
P6ZT*O>D7X)"'P?AZTQ:&!ILZRC_3E>YD"AOS<YPV(JDC3&O9+ER'H@-+2$SP_<7X
P*ZAXMA#(S09][._S&/:!8/-F^4V1;HM&[7.^5_9EE@.H/CVHST?PJYJ[%<[:X(3/
P#$'GWDF^_7/6%J):6V*6?&ZKKVS&\CI.F KT9EUR642.^)5T\=#317RK0W#U-/B+
P!":%@@:PR#X!JU&2UXJE@.>G>Z"8_BMGRB%V4 7SF&9/-'!Z#1H)<FB(SLO"Y70R
P_>.=6487=+@V?$.%"&C8O:27W8OB, (0@J-,)QHP@=+'!3,0CA]**5"N'5=O*$"/
P,J+K&F[?P#7NIM>]<&$K+U&&KS)ZWM?"H)M(3!"LO)^L?U]6RL[.U;#!M'DMF# G
P0AGJZ<(OPYS]1\'6]9R]EM$O&(,L5+!^'22*Z_^S _-85S.U%<]RY:J(E:9N-(@B
PU CC5$1&\(8UD?N>9RN#M3-R$6> =_9X@V,:TOD=8-^3(=!R*TC78"8%)A^%0U$S
PPW"9(86WN/KI+CG*1W>CV>"F2DOWO6O$GYU[R*GI"B]C%K?"H-3S0DD\9GZ4TH*5
P>(Z](_;-/RR@AU,L+J_@(EX&+5@3#?Q1A@? +;9FZ(+F"J3"4>7ZK"1CE!54ND=R
P^#TZ;N2+P$/K5SYJI*Y]%OD2H;))EL?5KMU7F@AFL3_S(^4P+^"<_-Z B#WN6=;X
P*QY?B%:LUN)(QQF-3SG)X"-K%-T>G>\ICQ3L-'2K3O]I3X!AZ8F[(B1:&GZTZ@50
PD3TLI69J5:%[W/W4^ <T=6?E@PE=2:$)N77-7I!KPT.:V_,C3F;8O8\!]T<+*"R)
PH7%"' YK.WD(_'M2.S.M4S<3M41,87<CEFWDRF0"M[X)7NW]=33(HUZ5ETL2?;-Z
P393_:[$VHREP3[^8WP(^H=$"U;JGK$>7GS+=" N$D?(JX!K'X!5Q:?>=6>59&>&O
P4Q/01@A)45GBY6\?)C]QE1+->!:[$THL%D1&34&N+Z*24KL?6"[*+Q PB1O@ "83
P!9X^-7,(BO3M=+%S&EVXB3S@JYGE<@K60P<R*X))X/#9@,^0='J0E5S$]<>D!*'6
PILDKT:VN2>[^Y9 *B+%C9;[A_\XSC2%+H7L)4]WMD)<F+-2$X%?%M;,@@1OI&G:M
P7B?>,2[@N(!5[5'GXFZYDZ:AR=K<5P+@+_1L_GFE8G"@H,7M' 0&&;5,&9,GZE4>
PL:+ ;[G;JW#,HN>6^<AEQ=.6QJ7+H?/B6N[68>T=:""EQCGVMV<F=A9NKG3MT0A,
P-,$[HKC"T=@MH%*],$@A/F%)%-]F/EH4SP$.@4H1(Y98MY/JP&3:Z"&9EP*T*[*3
P05<<#'N(R_J_-I\(%E"0 P!C,EH!#"W_ >'*LB^MU1+*C%W:<[IKU)D5-@LYEE=[
PH;G<E[QKR/<FA.'LQ.G_5PK,,0LMWD1&<VZUG\A=1UQ82U1K)?Z6M<D GWW2>QK1
P],011@_J%CZ 2P9$Z#2,#W>>N@L^=E_YLF]M(%!@D?=\HK_ ?OOL+;G4JTL6$_>.
PBG6T$X1>-B@ C_RLX.+&"TN336P65WK[,ZPWM!O$WVM"[R&U-Q-8'"*M6B5$0=)R
P)__G*!@B[]<=W-8$2#J4=1[M,073.KUZSC(.#.1J<CKRI$O%X]8J;G"5_, 2%3@@
P4<"D]@*:<ZR+V_.PAA 'V+$!///3YM<-%_(8:^7!I0EC2!Y4O22C@C[/^PKPRTA1
PH S@S=M$!H6;\.>?T)_"6SA./T*"%E0!7C<)-X.%$XKK& \42#Z8FB'U^M?&GK-5
P@X(QBI,[,Z+%:YZR*,FT5@AO4)$5QB7Y[, Y.<DP0,#]PUX>''/*H0JFBR5LW2%%
PK(_1G\&>VQKILJ%V:?R%%3<+@C=KN.56<#Q"2+^37B4H(TP-(8Z)E69 .E*[W$W;
P$(X$XWZJ2)7$ -<GUXVI"Y+B$52GS?O371KK_CG";$55<0;4!"EK&G/<3ESIG]DB
P !F4ZOI^ES;G#5+4J-DTN+O^\-' 0<7#A4*<][5M="T]:(&NIP:9$I@@3(5P.];%
P?=42!C=I".4IFV$$ +K4U<LB_[1R( >UBKJ>$XLW\O7UI9\KH?]#Q6DDF(9RT6S+
P@B#;+1--3"@=Q2'7#R":36_ZHD@7M9"IGH-L#AZ<,:H&<D/^E4X;8O1K'!(,C[N9
P,0]EL,1C"#G;J9J,;(;NET]!F+Q@Q:S?I^2WYM#!V?:,D@?]EK<1*MA?/07^\[0:
P*_6#:UL"PW=@081U\%$4ZXFB<7'H\$L9_P.Q (^,(?)XWI/'BD:&7.D @U@EX)C*
P0<4^!0&! V(K@Q*\.TAO9,R4?78LX1H7\CG((?ERP1X_VM0*W((*M6>,QG32?/^W
PH(Q>KSU4:U!K\06[O[I%IV2^I^6 D<)I=ICR#NN5H9JN#=*(L4N]VZSYU>Y-2SQ;
P?.G \J$3UD?4E6WKP132 K:HLX7^$5F[H'KW0:JV.7T)4.YO+T)DH%\6S2;INZEN
P,K8M2R*W\(%"RY@:-#&^:[[O@7,@!/D(OD,P!JR,<-UWGYS6F_;L>>CUKK'M\VWG
PZ*R?68'PQ/D@8OT=1L96R4J6(<X_",JT!7IM<8T/$!MU[0 M80U81;%[R73989:G
PDI5X?FR#7[G5H'XED?W6K8GIRV[^?;M NL6\^QZOQ^T8*L%6#Y4A%%=5CFK^TNN_
P0V$>EL-V =,"C*Y5U9()J.?UCL9,=7,+(?85?[I<!,LAU;F]]WQTFG.L:'AA*^?#
PDN)F\>RVVIEW*;''!\[<?$_KIR"C3/Q<);@51B&^L]C*^>Y>AU?+;,8EC[,!<!=0
PV>1YP\97UYX"B1F"OM$'VZNC$)[KHVXSCN^?=F,'H[S!):4&3D55)BCW/35,*$8?
PM>RC<57+H6*F_$]$=%HOZ+T<,ZJ7T731<09/DZCD#;<K&01T8@9F/?ASB!)FIPK.
PE-<T@S- V8VO"VEEYX]]L8@G7)+MP+;[5$2PV5K.B7N^:%L/9E)\M$L7()DP<A/(
PSR[:L 5%M6=2']46R._>^!J,0HU):<FN4*83??O##YPP'7?3%RRRZG=84L9QS/0T
P%=]T(;W+RDC[C^4^5Z5EB?6K@M)TBI+:.TV#]7H8G!V*X_NO %"!_%P,6R;>P_S0
P)8U _\YV9&R7V_XA7MVA#TD$JF-T)S2RG"BK4YL> $Z1WA (J-QHZ]?R^-%YT1KZ
PE+@5M7]['_MB(M.-D5H44(!4BAC-2F4O7,0&_(E!&[G> N*X%)=$\6FUA<#.7E$=
PP.AR\E905!]Y_5;[8?*[<K"3HC?5?F.T('DV9H0/V9(6H)SG]2%,[08HJG_JI64%
P(FVWI#%+\H 6/&DL-Q("I5]T($1JI$!92)H<E$ %+4??%#A]\&+G,^@7W,;*VJ\T
PM\@!<CE$<LRCAP!NZ>1^@#+Q"W[!9K\/PQ?U1"ZO13-OI6'E03D)2^K/[];D3Z.?
P$0@O.@)TGW"%;&"45@W&AJ_R\I(HI$Q^K-8"_QW,0'NF =-)6Z3>2)[+Y*.RU6WK
P3$N,5DC<7%!<:RM0<G4L".?I?R43H7&&7PF..SYR4099.=R""2=4G"II:_HS^NSO
PY1O3,]*U8$@NWI0F4\#DR&VRT_IY'U45\0W"67)Y*C*&K:@D94U%$8T>J;5B-KTR
PWO_Y;EP?OC\\%?;#C4DX]@0$0P9OQ^5^AKT3N>VLQ],Y]=UZ6F_=G?O_''(WDKRS
PSJ'S7])<W**9/9XJZ&_)TY%7?"_FV+6HA2$ZD&AO4&1G7"QO0+,N!X9/8,0!B(F\
P##_\A82#4FT:Q!;\\ZN,]Z;,E@0&Q#L?#,34DV&BE@XJB138VP9GG0S,' +B-@<B
P&&@29(@-*/M>=F\\X%;JVN"UJI.LL7]CF3#2F AG'HC\3*@4X>$8&(T&;%KWN>4:
P^;91-35L4BKC&(5WSM$2V*?1I0Z@73\MY$\X04[:?RGW);FI\Y*X54F_YOK6%$&=
P6@43U@+5&5 4^^1D[>J"NM2*%O&M@R0K H%V9<N"S(7& =DOS&/Y]AK_9S*JP'(<
PY^R<)O7,DVGQ8-/C>/,[G1ZZ[\#%Z#&W!)^S0/;CL_M82AR) "?\7$CDA6 OG%']
PV@2J<RZ[>8>AVXT^S]:PSVZJH"H[L3W- $[%\#.3"3E/7O)V[A9=8Y!M3Y3%DZ)A
P-Z_Q03F^Y#)V5-WX+T7JF%Q?B=#[W :&_X,'&\,8!@7\X8K3(XR2]'A=>(' C+ZU
P*MGQG83H6%<R87 ^]$^(+VQ('\1 ,$Q3<B!+Q(Y0#",,AD2E6OBZ@[[L+=1I RVW
P4$PSDQ,7Q0 ZS3QM0X-!:>T?<&K+/K_DF]$*HJR%0K$*\JZK6D0\GI;0R 7>_65A
P$:EZ!E  ?XLI!':]C]6Z&#6W% Z,:H*VHX<S%/D?6**D53>-0K17:3GI"^+49+'G
P^I-WJA#E2RSUK4S>DH]4\SO0)B1SO/FYQ/WN7PZ+WPIGV<7/P@OA<;V9C5L=$K#7
PP;0U'1!(CV::QT[L%83MT'5C8221*85'#'-Y'LI3"65,N2&#DTX^__E6(@3)>S-Y
P=T8K=JIW8!"/UGSWD _$OK-][<%^43P-6HRCF^)OI-KTDU5BJ_SRTL1TV(4;=:-:
P\K77H/GG#2W?5N-F0I=:/%=).=6LR/<9T<@_$.0R4%,%2K[JD NX\:FPERAZ-%!_
PL)JJ);;=#C-0RP!<%5@VVRSX.DW96[Z^H^&(=<$D6I-;[@N77<[60'OMJ9PBFI-[
P>\R*]U6.(NTC8,^N;<!MWGP"3'K)_#9CEWIZ4F, W4/;A06I=7B-EEGCX%])7VZY
PD[%Y]%QO;@Q%$<;_^/U4U0&9&.[;1DW(TR&;!D6$!4_>D:J5);TYI<ZW2_.R$ALI
P)SI]&FP)ZMQ/Q@80"X.X<3SKC'->KQ$*B;;)\/J) +_9G#QL3P[ &:E>P7-!4VW3
PP$G64S(: ]?<4<.'>J*2,5+6F3WSZR/XYOT<-Q2'!D^^T!(P:5'>KBP^DWB81!%P
PIYU$PCJ(9H4$&C*QYYN5G[79][NL/@5WRW>D%1H:9UAR:AASW5SV)#F:U%)%/W07
P(XI$-.1B_PK3M1$O4L?0  8/$-)4)PRBVU7,]4N#G3P:CV>1NOFM!<%^F<Z_]!P<
P2D!.0C@C#V%8<44>*:":?6P4!.0 /E?DC#!3D'34HT]/4\:(8I@F3G9YW.!UAOUL
PI\O;4GF>4-3*^7G1(LF637"U;R8 +,SH.,\F;[UXKEBHQ4(PFO^X;JPLO,2T0$>'
PD3XCW+.7_/8XAWG 'JNACP?U'QAN$:2X,?' F8YOP&2F>YT'@HYYD)X5;$I1;UA6
P !3,7I\!;EXK/#./,5%]4]><[I>=119K375=RD.C %U(H(5-=XH3Z!.7:CGH)/GD
P0,[])(:@7-8.+8B4X97T*;-]?T==X+Q>AX6DA,XMO>1KIT\ =<L>Z?\I^Q)]$,#.
PH40\H5^CPU5\84&107-=X[D^Z-Q9Z#$M)A+L#[K1#D.(",%#^U&LM98.=I3G'XHF
PMD<SU/IG'AN;"$#RB"* EVD%0%W5JL&(,?_R-E^TDM;H*Q< 32;.C,7KGF3Z?:,[
P;47 7SO,P9E(]]%XS(O!IXR=E]+>$C)LV\93V(/5I*C%PU7XT-ST1,ZY_HM$:9+(
PT;0Y)X50Q_D(#,,'>,I8R(E$6AW%P&QS=AV]!>K).Z5INL/S2[$+C7;]WZ FT44B
P$3C9Y =-6_F,TZHJH)OZ>MN-HO>)D4M4%ZQ(Q3FQ)I=XDC(885P:L=[V'SJUD\17
PKTQZ=0%!;A33(4X2MT-I3\^/BQ?5[^=2.H(HP;E6>-[J1?G!]2?/0(C^N)+XB=,B
P\7,+]VWDDS*^6#["C;:-4569^VV$XJ4-W.I97!Y^4/YS_+R'"2(6#1QQH'C]C*M(
P.XF5I+$]9;O9@JNR;AEI8;@Y0*T:<T?1\B.V1D4S^2X((T9_/IN@PPFML(39&&F4
P=:X/L"UU=QFG8@3R%O [(KF%@"[6R"7N3P8*$N N8EAD7*]R*\O#BOVO=-M&CJT#
PI<Q!@K3FNSF#0%FWU4=*4>!C#[!'26Z@Y@I?I[Q9R%U8(BUC6&*$C6"J@$^(YB4]
P8,P0]$A/2D3'V -0F<1(=NV%G2&!'<=SO3CTS ^F[V$DF3?X!H#D-%JM)6H?38%@
P; '!:OT,MJ-R+1Z:>;S44T_N_/$:PY%=U63&O:G6O"J(Y;K#W3[J,A7EJ!RK:3F?
PH@;0Z%4J5R'5;38N7+\U0.X.@S9;,<.RTOS[1TVNTL8SR&Z6;XTA ,MCEM:<2-66
PMMVH Q(JKF8T2^\I?0,> 2DB8"R1@-)&"#$H:P*S3R[ZB.+MX5B L%RUBI_UX2*B
P;),"!ZW*@Z*Q\[78;37)!]J(TH@C$9"<DB0:<*@A%?X]G2&.0\%V])2&9.1AXPL2
PB%HG?YE#23=KT:80UP5]X?<, +LB-/I]Q")^+O>-$ZONW2Q%%_=!2UQ:=[#&??J*
PE'Z@G"VCKMIFHZ1]M;L,5:9W0_J>"[AR]0B.@,2?G!9 IS_*JCYO0L#%@2;@TCD[
PB.WY B\+@@<F]R)35UMA[_@$QS[TGB!LBCF8G>,B0_Z+W0>)U*.Z\0#I5_9/!^5[
P[:P/1]?@?HEC<ZF=[JLWU] F/0&UN2VQZ:F@L"]JR8 %"S&#]$A\$ %]>>AB.V,,
PC'5F!Q34&Y@0@R(&V&>)L7Y<\=/QZL9W%3]?ZFMK8W7!%'/W-4C?28]?#[R!SFA@
PS7/<2CFBFS$F&P!F$!*-[RCNJ.G8U?*Z+MEN CM";RE"P[IMX0N(T/[*<.F<6!-M
PD.1.3:HTF(",BDKJ-S_ZXQ+%;M5 8+)C0;D"E!L%$[FQ7PMGJ=_JNT!.Q.OVE*LO
P/8)T77+XN&^/0ML=1I7+?L?_7U ;>Z'>@G]&.4\+$/EA!S%IM5% /]U[L3B5\N)?
PPRR0X>H-V:M4O8N\S%9;;>0( JWY5>&.8[?^C<2\BL%WF3F;!#3ZB4#P-M6:4%-K
POTXE_]S'72C? 1[016JO8X"@;V=3R8O@15#H_)<IX"=&8\8%_.P[ _770EJWHR'P
PYBEG@Z>J46I>BK)T)"OW@W<P-_>AL4O$.=8XL*GVM_];@[B <6G'-7JW<^,5<F0 
P)P[]U<@9W( 10V7;+G E<G#*N4#Q00W:H8 ?S=#HQM3A;V,26+L)*B][Y.,7B0:-
PATV&KK@KA,+Z-.F)_IJ]4NR3[QTW'6)$13W&G4%M;!N.X_@_K!U]X 6^K9LKDQX@
P6,<G+-V$?ON-1]D(4::'C)S9 '!&;OM\:12MRY1; 105S,)+YMHM25SAQ(@H6!Z5
P_G'92!6@AY9<N@W?.YA7ME/8[J/"(. ]Z8:U6CP[?=_PAR@:A6=X2EVOI$R2DA-M
P:G(K&T9 E)T3=G?1>E-4SI N$_,@FJ7.,SM\#P??+VL=3TEINW7!SNNLGTC9U4IE
P.R>+#,TRG$A=JH% 6^&/M4G[M2O09J5<\;N8<@3F_>8WJ?ABJ,V$@M9 /,)?36B5
PA]C0\XVHL@B[_^HSJ_ 3!3V6M03Y+.Z^W""U[@)7X)U\#O*C+]T((NC.$'#U(S"!
P@S$Z>6!AEW_;T-^)Q^M;@_-)+'3R<#V3S)W3PE'E-K[.!/=X[1:GEU]IS "$:]9V
P1U?(/,IO2YX>/GWVK_I%'0-MQPW3V%(_9+J_>GXT2U,R07FA?0ZAW%]"X3\U#BD&
PX.*J^P!8A1O++=)M J8W'DUMSLSK9:PEJ<Z)F;9JCWM?SN "=&AP *3.ZFL7(F,4
P4[+5IA(JV"I)(V%3"4?9P1WKYZT]#9/.MWRNMK6T&\A'[LCL4L+AKMFNAC*W?/.'
P&+20L8P#D/S5\\TI>Y6O+U/Q;=AX<.E: 4L-(#O1"C]US.:G8S779$&MA;1Y/@'(
PH8L.)O?R*BU3#4:GPQYT\K1^^O>T,P!Z#N6C3#](:*I&_1#NDZN1P6";3_WIU#E"
P- T;-[)XR1[N6%/5IM*J.$)U1+)8+U<..L<:);S5UM>P:(J0%%4.K$?@>.LGBXFB
P%G>09%L]E^A<6/CP>?IDNSO?LB[URM+HUT[,]OLC>4[/V:T@[\7OEPW)00FL.;SD
P!"+**+YQSO?BEBK&<(9#?+&X)$0F5Q$KE'"_=-H)E1!"6^_H7A3ML=0HO1+7ZT[<
PIU1$#HUL:"Y7K_Y%]98P.#>O=ZXN%,[$0J=@ W\_CI-"@Q0>ZRZCU;8E7L#+H(P@
P;Z.!NN9WGX>)[*6RC.<I2/C^\2,W,DM$OY!MN2GWEA'+1-MF64I8@=XF$^D9>\(Z
P2#1_9.QBZN:6)F9%Q(0^ =*!LFN<PR7_]*ERZ(*JU35=)JW1,QEN0.J6$AYQA31G
P"@$\N(*LZ>L92!I5G/]F=X8ZRT[+.RW+G"%L(,Z:%2U,1'Y+@U@)9O=2\O26J(O?
P>2\=3]NT=.JD<5OFA2-Q]H:DG4D]D_<K8:_2TEHOE\#*QK?3F\FN PT?;ODJ48;!
PC*/)'\['2$W% !WR%J?9WJ=]J&^:Y"L&:UGC.$AY;0,(Z;8]11KS\P'A0!@WP2HW
PX\QP>:Y:)27O5RJ$S-G4N:XS/@^(1GTO"O+2+E;(319C=I9G#)K7\<PVT>2\ X7<
PPI6D,M.B=7(1)H1=+@@B\0&:\E3!)(. ?V/US"46KPCH>@>]QW9(?FOP"4.SDJO;
P*(M\Z"A(C#/WX^!G63[2K(]JU*DN 9S[W[O("2S"G,:\_7J8@C\;WUJQ^#QR0$+ 
P,@LB;L!._0&A2\&,GXC*]4L8$C]3,$,*Y>XX/3RMT\9[-Z"D&>XC&(W-(AT%>VR3
P5G/!0<!9$Z-8<OQR^!Y60P$X3/ 1.X);WJH($U#?I@;$ 31'[F)84*6>^#@T09!#
PDFE2.IM\AT+Z-A/W6CE1 Q@FOQG;V6=LQ$,>2]3)V?4:/+*D1QUC YTY#FFT%^O)
PLWJ!A =^;OL5G:LGLI7Q+,;,=:_CV%)DL!]8LJ>VVE=+62];M0R=B0W+*",%L:7=
P2A5U$\ F:^<7Z<5Z%I2GA_V,QV)*6[#7$Z6<7#/KJ7D:4B15RYN*GX6-/5(PHCY/
P5!WXXA/R 6Q>WAR?9&=WI6G%!-^W_(E=M:U%D#=(:U5$ R*&(:25@J6OS'CK.[XJ
P*0B5[$M.8/>Y4\(A![G.U@>%RK@@:!S4%=P#4)A:!U [<*QC0,I.^:KY(8; BVBX
P@O0F?=PB6MBIX,'A;G;;3I,I4-07K/:HQ@6%@HQCJ77WX" \!+1QAT D=@WK/@84
PSOGL0G1LV4*R/5_W7LCP @XL4W52^I[E,_C:C@8"= 7"W+_&]E[QZ,D)^?/U,MV3
P3!Y(PN\ZD^X^(0\FDQ_\QK[=ORPHU1(@ OR0R'3#.U^0 ;P7CU'UC$?^X6-PZ6S0
PA^'<;<UVA'V^@%[^T@O)W[K'I?OJ.CA" ETKPP_W<8Y[0WEWMP;]M:6BN+;ATDDJ
PQ*6>G!/$V&Y'ZT,TRFK-I ;\B>N+_R&=I).QVZ:NBSK XG5X^K)@4LF??JIM.?>3
PRI;!D\@)?\%1'I5Q=7P:49.0X<W375XYZ&708JSI!CBB[[U.41UK&KP6'1LEH-+"
PYU6VP^HJ\+"I(E3HJXH^>MXF*W?2]W- /Q. OBHGHN?/)8?%T+7/NNY?@3MQP[_"
PR^YRCN6V *>_0B#;30UOLM"->#TS!<+1WR^7$"Y^M19T\RHOP'B'Q,5G,$^<LS&X
P97^1T^QV2\5:[QM4F"K'/27DOSXLR24ZQ(N![P?"U]\+V+OU(*B[0.:3W!V_E@RS
PD)G%QL6N +G5RH?">';<\,,3?+]6 (OD)E9,8I6\:;&S[*&K"1+^*W/-:]:-N?TB
P?*#H*$;JCV%!#EXF!FUVQGAJKF+KD\>P:;CV9*Z'N^]Z4<Y5A5'%U@&_# X[2V$5
P:CM# S9QG1@"LE7,VG*IZ.\.X<!X4)?0&#=&/;5=ME@I,QX#9T',0&!U4(LO#D3#
P)9&AMBQ0(%^2!5PK$V9]L3E-2@%N4AU(>5J[(K",S+2Z./17T5XI"^)+7;@V2S3O
P'J.K/^[R0N9>T(GQFKD-/<G3#RWPZQPZZ MBVFXH*FL%1!>&@)NBBDJMQ\92[+WQ
P;P+%EBQ^NR,Y)1-1=F"V@=?Z0NZR-J] J D %F9>_'N&,4>["O5)#X.>PPLVM6Z;
PJJ=YD<C]RIAX\ML1W!/^6'(5D&;8&?\#N[[3)X,?ON5MGE:QU3%)N:X)X5:,G[;P
P;22*)G&9 _!)])6R7)_!F'LVB4OBTTKH-7DA;$M?>]-^ TG)IN9W<<$QW7-M(H#H
P=KE?_S]J^<%I.KH'\DLXD*]I=>:.EZ]A>5WE:LV9T5P31XK*3V;K$OJY=B_<5BEU
PJI;.<G#%QH.NG&6EH[(V\$@=GZJ!3!5;ZA8$7Q,>6!WS-H2S&&4D2O92\8,]HI]6
P1B!PDNQK]RCL\DOS-(U%![Y$M8=-78?T,V49R?#(LF)P0!&<ZP&SI3((N(<Z%SD:
P&E-V?BX%"S3$&5!"YHN,9\P1U)^3EA'&MP,S]2X%)R6OVI%Z$6YOYL#$@*Q<H^9.
PEX00W4W-BC+X[V87T,Q.HR<SVY>%E5DCXSQ#:#J=0*#&;E0;.*LO_(!K*U'C-)LX
P"K&:]K.QP%,CF6>72S3&-?NNK8)!0,[9>@!8\0ZJEA1\!=LZQ*!AVC1UV /T-&$/
PY6D?CPLC:.RP^2Y5 Z,78]<SKH1U,?/G,E?NZU$R(_A*T#,#%BW^_=?RQ7&M-G'V
P!5.U]]H-U6LKF^5O"6M;PL59):MPP-.$D#A=DE@J3)]17(F+_450# )$\+TW2"Y&
PENUX,PV?L_<UI+@6D ;DW;4!BM@I$C$S N&'*&?S*WZQ"&7 ,]2G(:PQU*8[AD8D
P,>[;&C_'_S$5@!00W@$;!.@D3EGU(!S 9(LBC<#L3,'F<C:&P@'=W?_$M]=C@0J>
P?<0*$*/ASUX<# #>$L^@VUJ'($PL>9JK1&U$K)@76*4<1UVS?S8*J6HJCT;KD<0>
P$0OV]HDS4V,TCZX=HEU(9+C.7F-^,9E !YXG[)C>@\O;D;5)<A?KOYH4Y)5-C53<
P+>^-%IV 5*HI@+_>*N5RX<AF,!A!%G3%+I5EWC_T[P0P2UE6>CG4N5B6JR'E8W^#
P-86)QTU>UP&@(?,+W8[D6@.NS09)6CAVEJ%DX\,X$;=9%V1UF(#%F9:KY8W9C#D@
P!!PH\\YL^R*P$RL>!7>@M..1'%M0=#.NL2L@\>UPN;^'<?BUM2VX0E:MG_'L%_Q 
P0P*@@&T,AKQ"FK1%""H2$C\>,'!:9ID*HO[*9HK',G,Y'5]:E>W]\?5,-EO9MMZ%
P?RP.1^'15=@)N ,G^!)N2A(NCHY@2[,,J "@4$PK(/Y-+ROE$=C(?C23PL?K'YTB
P+_!W4.XV,E>"WA6#3S_O-'O>AY$;;,_J.9M':4-V2JJ-X_T54C6/:_#DNH@F! 2C
PH1H]KOTY@Z;.T-F2./5<_5$HK<Q=61Q;H#N@V@0WW7%@^OZFH4)N!%:>$H0%QR"&
PPR,^J^RIMATF9]_ (/DUXNKXI*(U-CS&(MHJ!*JZ@XZ#M/U^;ID[C?7OG /@+;.R
P*;U08MM7:02MRD<$;82WKG%9KR[:,."K2;-(2@[C,9+7D@A> Z,=$H#OQ,L];Y[L
P/-'<UG"4F.VED1R<T:KHP2.BP38T<XO7WM@FZ<CW3@5%:W@:D"_ 5U0Y@]$04DO_
PJ'I@G<B,WM30P>E0O9"-]@>8JW>\*K# )CLS<;NB'I,#VQY6#,-Q@5$_FRCD!D='
PF!*04R_?,K AU<:M/K8,I#02U>O A#7GB=EXE#NIF?&Y0".ESP$@)_GU[3K,:D8T
PGLZQ,J6P2?H"HK$R-2;;1APL$<UHV9%JFE>A58QZ;Q#=\6/2-^'_F'6H?LNMT&%>
PR"<52PLO@8-?"G%;0=R/GA;]9N<G9++6[CS5-%85?)U)Q*&F*R !5G!M$H97#\U1
P_EQB<,VWDMZ.I+@>-YAWC/AB2<&G=(OM: %=C*]ZOT)W#DLB\<(,G?#AR''Z4<0<
P)5C3TVD3<B3G_C;JF:<(/52O8N^PL^P4-4$J$_#C=O4!_W7O5#?YB)<<C,21P..I
PA7+3=HQXLW+?$6V>M'%,?!>$>:VL4<[5OGO_*CZ&VF;\]#N(8CL_;C?<OVB6H>GK
PR:0MXA62A[6>ET#TYV$G_;,$UXTY1.&&H8*O623RK]B%*A/99LX4%6.@$"^T0:22
PO2S ;.65-ZB,(RMB(.*=QNXP1UL07LK^=KXIG.22)HZFX5;Q9;4:R5:?SL52<-H#
PD0(<9M<+1!U* UL)6\P@,6;W' ON(=7H _GPQX#Y=C_.L4SS\>-.'?>=2E1GTK@9
P!O$L[7$9<EQLR.CTHOO2WJ2#94>E:J,8V8V'A"=]?T878=F5=JK2SRBSKFHC2OX=
P"6L1BKGM5AR;W:>C>D$"/$$X9#H?)]<UHZ_>)Y#^7$XLF=X#ZZN5ULI^I884M;=2
PSS0OL.S*^=O"74N0VCDLX6S6HKG2>N\;*$+G->VO?ZVK,RY) \(<AFXTG1&F:/@'
P^IN_OTJ<+!F. R\O=.:O@?LD(VATO#72]D?= L,QSR'AF24PK=>@VY%8%A$S<##!
P$ENYF3MMCZ)QLX0!,* ;+LQ7DI$;)9&ES!>&D7*HD4_\F#L/>P97?ME>;HXWG@2-
P#*2]5?Q[V)55=<4$N:NN$SP_BNF 5!/1+JP[QN<@RN(J!2+H,A5.,XC@)@3UC4[J
PU(J#"\ND6A!--^WS4Q#R+Y[![A^P##A\8.'J/?5CY<(2"0:D%&_J/IX,M!(])@^&
PI:EUEOJ7FGZPA)!^MYEY98T4#:K<&K1C.JGGR.5%3Y"?4$U:*WG!^A#5ZC_P1C36
P]YIW-R'FB6E+<E]J6K>2L9R<=!Q[0;4,',^CNNQ>R\XNFSP1O]2W69&OJK.E'%52
P=TU KTXH,V_\1J#D2\\5!N*Y4(Z%V*B&4][_BQKGMB&''74QY*::<1)PK%\LVS-D
P]+? *OH3_L0<L_B.7VJ UV4PS2QTX5"O<[T(=,?T_&-K13BF;H K<F( =V;HE(X/
P9J<3/2]#D%&1C6]_^B3JC2UG,ZE)CWK5VVUQ2FI':FON*HZ2CNGR$N$<"C S";^$
P!&JN!J/SF#(NA@ODOTU3STI(ZW!TI[U:**_#3D\*ZGTEA3$YGPAN[G/'NPT\(L51
P>=S ETNEJ%\!)IJK7F=D;(S #E_I@JAZ4%$Y;-V(V(E2-?'^&4-L%5JBDI6S#0>@
PPH#A^ <_-[BG>V8<5W^<36>08DJ3ON79X#&ONW^K8^!"^W^2W:\5]S0NA<8YQW:N
P5R7+M2H>I\4X'Y'_8)W)T\,_7-\P@1K6M9U8EPV6] I;\O:SDI_02#C2T\%N+0*Y
PV6F;?U\J\=KY"E@G,7K.)V?11I^Y+1$#PP4IFA3J2,L!\DCCOAT_:>HH2\MR$"[/
P^=@)VS."YDI#(0:4>2:'O&2O.^/W0=9E0$E3"7=J[%ZR_^@Y\=X-[3@96GUVVJ?%
PR:4&1V?#_V@CTN%O1Z845+_#Z,GR;^*R"/:-9^O!V"S2TTSH\!SPG> ,>Q60A%1B
P'$@/(44J3FXQU^K:9K G7*^-CS&+8:E[ _X@#%+%W3+4<ABP%M-]"+"O6?3J[V(%
PJV-0. X<"3=RO"V)8L4XN4?91CJYP11*(FEN9K#E/T8V_)L W<P.[X>.<@?%5TR,
PGVC8?GN4(K>V3S.].ONU(,G2#,=OPI NI2:5;"\+#S9\%GJ+XF.\RSU^8%6MV 4:
P*CK6,2O7$1^B,V:7I3D3= OR.;-"W. /$YQT-Z[0(M8/+L??/L=QNDP\XN*L<ML%
P'W:(U7]1 [4/X4__"I]TSGIX)X6J6SXR[ ;3^X?UO(^^"* V-< KSSN@9"S0*SHY
PG_V"2=0(<Q3U;$4W.)6MQ"S\0N)#)4'<XC=3:5UE.C?D3=;A$]3C1CBPWE-5MPXV
P&EPSA4[13+P/4RC7,HH/8'VQW1%4:"(;*">/S*?H[I8SZLL-W@Y+@#AY^"&_=[ZN
P$\3X"%@J+-N ^>8);$\WQ96PV,]/;=.P'9[-$E_B/T03*">>\W:T80M;IQ7)28+L
P_F[7*!G%B)$J\?T.RWV^N@*N^L%7F 6*$T%Q1H*EH1C--GIV7+Q2/30-@O^SF2V8
P63'63D/6?<1PC$6.5VIPDDCN(7.$ZT+N09!UR^ZA23RV*W.$IMS\Z1B8.NI_BX/=
P%%;HIG%('6,"%:"\V+JHFRCZPUSF)@5%ED":P'?8X%3SCP$)5&Q^2"[_I>6F58BL
PQE(V_T8-$/PN^QXY VOSI7#?ZB[#J$)&V/>+1B?!/AV[OA$H7BYOB67G]/%9(A<N
P/,@H#'L*R"?R[9>>M4C6<>RY<50H']8B,?9RL>V/;@0#-4?/;?%5(^IA#JY]3N5M
PXYFOS(\#7&7>0J*N4_@3HVLTDBQW.L^Y5F.>$2F/B%IY"2XQ4O%&MY@B4-\[A:4_
P5')3L334)&7@E1T<RYHF1^B8(FV1V#Z.L?"_#HY6VRW -D92MU$@TW*_GBD@8+, 
PS"+C]))J9PV%YX-8ZTPTO/?%]6QY&2 N%?-X=*F0CW:36C_WR=E?'3M]+E:XWT9Z
PEU5L*;Q"^>AAW!PZ BAJ'=<P/3TT\*R@BY31Y9Q0?\*290WE/'.$?MGFE D1K0P4
P^;&G^G2.0C=AFEWS@AF:SM CKR:$.TC*Z<#3-41,(?@40I^F?\V$O64BH>NYR_4'
P0$?W#6S4L:T!VMJN#M;IV52[,,FJV[9ZIL(CH"^C0:].Y0Y9'\(+%GY:Y9<WI9O:
P*<D;ZOY-3]! H91CRW[;LYRY^,]ZR3-_&\+L,F=1GK](!'7RR48"Y(4!*QG^S[#F
P'*.[9X]8/[(:'X(>U?CJRK.E;ZF592HP>4+D\WD#QY>J@&?_0$1?JF',U)I>+?7V
P>"Y 7[2BI7_RRLM8#KA$8?SMFY^:'NI"' 8/"I$!7B6J!B&@,6=GER:J]OPL?M +
PF;DA;]\_)8\" 7B#C!\:_\,0NI\=<4FF?.5UG_:@?B-8TT RSII-YYP\(CAH22V*
P=1"2_S=Z^J27]@&#Q7FZGPIF9F0LZ.P.A9G@K<@=5W_BKG9QF+'DCM2G$_<:7&;\
P8#8MQ_Z=T[L3LM;B*YJ%721O\\(UO/9HK$#V;M UTQ:EJ\#SB*-8P7<_@*9Y&Q^2
P;42_\Y8W*BO,B(K=P]MDY;#!I_XKY!^$'9O7>&SJJ1.D&7U/T$OFKUKS1J'N6,*'
P-/98-2'0X8G3@/@9(-R3$&!<TG#7Y/@_H_T[GR?Z=#58#Z),,F\39_K:.;#YF<8"
PX@.%(#!BY0TC83>_!_MVDX?L/?CA,V7X;MJ:DREOWX\/6ND8#X+Z30OA) *<QV$F
P7Z<$JJ+?_U)NGIUC93/%?83UUZ9;?3T@I;-V;A(OE<M1=QF57RS'YS%TZ0T!GW2?
PK,0&9M&WC'A92H8-EO[2<UZMI:8&'?,45$[X+&2E;RZ+G+I]]T*TH=2)<$JK?6PY
P4N1N&4*G+TNX5N/O<:X<JX0B\TW(F6#+/EHCRQJ\=H96#J9*)NT'TUPU6+U/0VS)
P.LD[@94$9J<<2U+LKM)EAY%6O0NX--Z^IB$C;H2:O?<^X+\NCI'KR?)HTTS\"<; 
PB@B'<\IC5DR;B)H64/OGTK8OVQC!HYEL&D$6^&&Y^E^1@3:%._B3&E#I:-]Y8RQ,
P%<+H1^#2G=J7YN1@,6GB]I=$<C;/MEP#$+1'S1P^AB1OK9I-@[<H1K:>_E5S,&<Z
PIZ95*_)(Y;H!F(:^].@3<^!SB[-^UQQJ_2<]"9Y07=2_CT)K&D,._V[G1>^SLP/W
P&.O&5]?FACEXLG+0\:P;VN[VK=LS&(R*D&2D77GP8=,J';IQ?+CTB6=#TNI+EZ^D
PSRG"V:!OCD+I)FKS*.P8.[7/ &>6\GI33.'D[:XQG3&>_);--1'T.='O?>:-J0*"
P9R/#&*$6&P;A?WGIM8>Y( JD\-;7(HD>AO*3<)6D&+Y,5..L^>)--=(9/NH[P!*'
P6\9D.W#M)[&F;G46PH^+P=9B&#UCG\7(7!A4+PT>G:T!+7F/J<Q-J@O,_^T>3*0@
P:$M;976+<CJ=1=B0AJ>S!*6_@E=C5B5J\N0%^Q3=9&3$H.N%XB:KEJ9 )@>_YT!-
PC'S?'=ITHE0[8,E"SJ,\V4.US7LDL*$@9BH:![UYF^C?LR*?WMP)?/-\E]0(T[</
PB8%[K&NOF'SM%V!7Q6V&L4GQ*@QQ%PZ'[H2"-+"FMR90V6JE] *[]8G-P-29C/ O
P>[G<40L2T+4^1BHM('-C'(U $@4:DB(HR^PV2!]61%1^=6LGG?;2MD8"IK:HQ'AO
PD>WSEUI0,TV8WL?\.DMY"\2P*X"-0Z;<FI.ZMIGWH)FV&A3N&E)'NX1QTXM_8.^"
PUL= GUKI#%<5^(H:=.TAV3JK4JZ-=)T$A_V^4<BW00T]<7T,7UXI(BR.K\UY8DD-
P9;DG/UF![[3Z2PI[_*T *SQ%L?$*!P*HM5678=*G,*Q#X%IP=!ZCHV&#>.H ._9]
P XX JC\80[B3^O+(!Y+RAAHJ)I_DL7]/KL7Z;'+Y:11DZM4?ISQ@ZHW+#O2[ BKJ
PFMQJD->C,N+.7$8^?10+P*HZ SO6R,(,+[%]@M'1\HRT[C:]B_J9E$GX^^@LKT-=
PSFV-#13/*&B2>DW_4U2HD7%R>#C +1B,6M1J(>CP,CRJ$=/)CRBQ0:5KTQNQ]PCK
P>Q=XT.0\<_/LCD!J\T>'O\W97/Q.KJMDC]ICQ+P_6!$>&GC&E:HL6^8]_6PU3H).
P\5RL95(H4M%H"S2%5[^3_VZVLT?)N>@CF#HOSXHJ#;#,ME??D_#'*?M:WWA@I-NB
P",#"TJYZ28^H;@DJ2W[(2ZJ^.)=KQM GT5Z.K"!SU>!Q([* #]?)FFEV6#M$HO?8
PYJ/YRUY[<5*@3O=DQ! SL7-4^(^)]/G[?5P>P9_:9>9B"4@2Z+2JNI=JQ,CFG%M$
PMGBP ^*/K$S3V'ME'1H5X[-4ORU:P3J.,WLZ9H<CR96K;61YM]:O-M%7CV:&D;+H
PNO O7C,';1IY]'LC5"]N<9<H?1_%'4!4.UQ5Q:GLTE>E=4X<=ME2B ),<:5%_0) 
PNFE57Z%!_06<HDZ#'8@#<)EK%E!9I:F7OZ0$A"_;B.[F;X6F)5',(RSJR;/16QVA
PS"7]1X+W!IV0$0<@-M&P7<'&Y+CR7YW!&-M52JPP=\9#]@6<;*MTJ=X^M>FM3.O-
PA/MOO[G=BWWCO0!I:_S&75R,YZB1)?(U+R@[QYI/K#2V&2H;.DLT/579[U@AM*39
PE26L/7S1MO]>_LCWXGN] [3%G[;%Q(=V22DWL<K/[@G/$;*G\X %^L3N .J5- $%
P' '$AR6('R!P"NVU3=>W-P29TG4[;ELGI%S1^IUL"OH,P59^"8[ W&=<OS?B]J64
P74O(3A9^LY/4,=>,G.B"QI:*#WNT_:A/!Y"%VW[11@@I\_PR?8(:=\_@ZEL0?@R/
PU7)K[!I%]3LJF,V/>&+V]S%#[]_RI"TRG5:UY*R!O-,$>F/<5CG!7R'UBV$LH(K?
PSH'SF30Z#F5@P-'W0%^_?!\2]/EB$,_%F2.9<!)F.J G%%$)=*7F_X/SOSR60'?4
PNLG3BB%#LAO4Z'YA&S)"%GA9+'9O#&L!)Y0OMA$5P*7KI 8O7BCL $)N-.<O[GG_
PQDI>G"/I8@F'!]&?;L7Z),YO"(2P^'$>]A$<)'V]6)$8@;+E_,D<^?3Z4'IX>S1T
P7U*.79L'9:GN;$S3M][@B-2YB+9;\=)!S(YU: FW!5'[<SC3^U=R- *#M?6,3$UV
PJZ<6LDPXQB+8<3L"HN_LNLVJQ@5E#D@*_GBX:T:@P0Y6D(L8M7?WJLH/8Y%YB?28
PC"=X)?[Z;D+D4"H?3 6%C(B![BF_99"E*G-E-Q-$F8(+8*,%Z+*>KD=TK$+-4SVT
PHE(F(496:7_1E2"9"2QI&H?2;4GLR";8A6(^'Z%N8'F-R!7?7*A81IC&U' %)X(4
P&K]%@?L5_&XSPP](L2-0"%&;59_%D?(_W9?K:>V>:18;NLGY*<GX2W5@NF%%UM%7
PB?" '>F&9+CI6M4&%O--EQ/YZNTPC+G'Y^L)(,1HGD^K.C1GGBYF]G(7K I*)4R'
PB[>,JGK9!+$2A7F:P0O\U!3_Q8L0,.:*?N U&$XR&@PJT#;J$(_+3/(.G\_.Z:3#
P]4"I2H\#(D.AJ,A<3G*P;/Q%M'B/G2VX;;QT;H4E!?V :=:/_"L>=&_+G)>H.G33
P3#S&E))=TOB1'27\7^'.&J?<IS=I,"]SL<7?@H@UY=HD$Z\8N=.A,G!H?TV/VX[O
PZIE%N#:<M38#P>5OAP846N$%\)[H>8K!!;YR&C7A]AS%D<O58K'+]J%*?X0Y0+0S
P6<)E1;XBK_W_JW"U)&=& #OF#RA V?I?,"(MKGT,1F@?&HLEDCG[45YR?T' %,99
P0Q9^'E@1[]A*F]55A&1B;5\?/8KCX+8?U))2*MJ/*/6)8ZW8*VZ_"6P<5PMANA S
PB"<'K#JZLKSB\Q\;*'M<2\C-A(9%]1<8Z:F/1E+T,0?-CVZ]D6ZH7, -GGWMX-->
PZY?L+W7YD]::[FTO><^+[/$1/5/QD1V+?FU51)OI/0=4\?=*3?_FYEQ*2DFWHNU8
PEW@:N-[7Z<F5-?<B#3SUS4$/64=6AZ3Z)VJ,@ =C<@M%3XA4Q7(KFE]%A5HPF3/[
PMM%RJC'GU75LMWS<<>! M"9R\ZI1&@QCL8U**E(0ZRZ0W8%W^&OFPIW=NA+:$B7Y
P]DKD)>JKEXTJ;<@.3(4U:PWEU#$DNG )-X<6?W7CX4Z(A] B"JQB=,( 8R=NQ$'^
PE35:=IF->;&1PVT"::M[5=*@;K)8<\'EXFA5);08G2K>LX6_<'>[Z66+X"TV=P3/
PQTK+1GY#<3+%T<U#'O3:BL'."2@5)JVT#.'9+^1;-HC$G$""K&1A]'_QO!2G,A%;
PF\12CXV^3(:FN%(&%3TG>"?FSS#1*>_YK[GSH?1%/R]DJU=A+:U%],C];AV@^!O*
P2T=*DD;UG2]]_V\JI5MK4:P6G[7W'')M?3U^5PH WQV :YF(16#B#6\QS%FK@.QS
P@XU'WW"*[\8%):7U;B%@(L,G4L 4^!;Z$I)ZIL_58E=6%B/W!F#FJ!YY_\Q(?>/A
P7/(1#A94- :W@0&5LHRZEFO@G]QT=0I//IW*'E_C+UCIJ9R^<MX"_+!="-80M5E:
P8#+VWU^[)^%$_VUESAEMT)XHC*P%Q0)J_?_%V.J*/>K3L7QU?Q0XG(MC38T#K+MY
P$X_Q'P4& 3"X9=-PES0%'7+L14.R)M@$!K]6"+QW78-_#:'VZCE8281O!73O^%5 
P3WQ$.V%1Q8P3<T!EF] &3G\PT9>4X*"/=X^6V1,*!K0(#0$5D(3$T=,'D8KWP7\?
P_I#KBD62B^E-$_?4/A@:7U;-T+WLWG798U:'+)BT<_GR4G-V8QIIN:-QW:FNVM0+
PAM?$U4>:O@V8)?3M2;9S<EO>;Q9CKW:[MQ)?8%<:88"#HZAK8TC12X1Z^JCM@J:3
PZUBW[)G:V_UU.Y+^*&&:IS:#<[X7*3"X,J.W^0+"7#0T\8H@<);K'NM[IL[V%1NX
PC\281>)H$Y5QS=%T,AR= Y<[ZNO96KP1WLO9D?V\TV%>@HU8$[6^,0*C-.;];-"*
P%_2*E\K1@.A94PF0WJU2BKU8))ID&TF4/DNGXSN'<X;8"Y8%U74GJ'Y^DZMVKNW"
PQ6,BQ>B"+1*4SQHB;,F!UA1H-5ZU_:5=4O[.)+KT%"^I"6?Q;/"$V>@0JIM(\[>4
P>D#^JO&WX[P#LQZAZ'U\3-\^Y?IC%OHQJ"EEZ'V4R:<8"-+"1=KCT$\VX:H9E-A6
P*1F,')XHOG=^SZ(C@+MGMJ\M% LE(/W9A02$2I_8W[&]&<.Z<NV]>3.)P:S$HCX+
P0/PK0%'-%.V[S_ED_E>/^/BE;O<>]A'W>)<*$=R^8G\>P)T_NWB1Q$DGN#VWF%?(
P&0AREZIWU,H,WM"LDOXSE(E]G[,,P^VR7(R11W)+H<+E].IEY,I":,JH385$0O3G
P+IB+TS4!5EI&RFPOYPXJA!/V8[,#@5%1PW2-KQY"9P,'^)'T^=CJ"EVQ)"+Q'C)"
P:<CL]'52Y.1&=WIV?U>OP*K.6IXL#Y,B(DFY5*L%0@]DKK&[JWS6@WB?BAG.#<3"
P0(06KD"5:WY-FBJ$G$SG-7+A/8\@6-@7?@-B-_OKN8&'M$S8IB<^T6'/)A2 ^4"#
PTXO$X[F>)/N0DXJ>3>=EG[!Y]I%[RN,Q$>'(6 1(@+?;F[>$F5!94ZHY0SJU![C0
PT['G/_7\/?RU;W@"Y$T)O-4E,GCAA>\ %'XL&CT7Y5#Q-&BBU*]SQ@P'17R!/\D'
P>4?4<VE9Q=*"-*5-9UH+MP4KM[A=E,BYV:E-("1#I<RC$2%_Y.'P)"^( '/A" DY
P<[A1HK,NHV6-\Y],X?QL5T+OBA7W:Q$1D,,OMZFLN($[$G_^-TR?G).89:(5@]H+
P!M@" ,LVM9N,D)UG. =>9R_Z4&ZSN7T\AW<2,GM:6,>-"18ZG2%K7?K !QI4)L6I
PF8@NYD?0*6D<"=JR@1)!]^O6-V!A%]O(2=-]?U<YR#D-.^VP,SFB9E%VM*'7VBJO
P+@1/%M8:TA=*?ZR,]KQ=N4P@.DDUM,>-<WP+^$OHQAVZ/Y"<RZI N5_] XO.LIJO
P/1AN"^L7PLC0G[[-$+K9M<H+4T>9!X_\N_%ZE4_+> :HK+)D0ZI%7K=CX%:OYFMO
P'""Q$P PKR;)Q-D@K GK!8<W)0+4K&OL>>2811]VP->>-I(MTG-%#X)>@7[^ZZY)
P!0:+.MK N)Y8ZX>9BAZ ZP9MO]&__"L\6U<X5_O6-QX^.>JL&["PWL3-C8LJ/T=S
PNL)^$JJ_]%'Y('-?]PE[4?E.(M1>B4'<?5'D/H&+%)+=CQ5_!=$59-%:)T.:%@W4
P!V)!,JUR=W3KC3W WF;U/TLZ#'L,K?V8\F!:=L' )?I&BFY[@(5:J,4I(NF/H?*$
P%SKJN*I7/A&";F*6:0](EZ:K'E/*I ;I(+XRCHGSN;(4B6S9EN$L_@OU!_R.W)];
P/'[X9'%U&< ZP90>\X:S+-?3MCYIRUODBC 1RL/Y.(**M=[\RP+,^&HR5$PQD=^C
P/JK6A(E)E<,N$:5Z(U)F2T>TT*[/:,ZL%QC,=@%WV#2:9^%AHEOP,45[P-;"N IS
PGRM\W&K#GLTKJ<8FJ_FFDU-+SJ2Z]PP<!03-*CKJ73$3"1K5&W2?,,NRR_=?F@&<
P*E 28#'#:> Q?(%F5N]VNIZE=$;-J;LN[W4P!A!P>HPV X(0,4AQ$C^.07/;,+RF
PASO!4]2W5Y)^4QU9&2][U;VMN- Q8$?%J_+8( 8AU2=KLTH8'\,$X-CA.81D4E$6
PN[C6^R4#8,P^+$,0,*09T&^1M\E:_CB#$">:,LCLVW#(N 1(_';C/.P>E!EJ7_2^
PGF2B3<5.4#7P34^5+%C8,4$RJ/JU10SO2:[FBJ+4;R_I,DS"+#D^AQGEU@C1:WLY
P?V\.8*0%BT!%Y;&K-GL232V=F_A69"ZSYI2I-P0BO-$,TY_3AZ&ZTVW*\:J4GP ,
P74.G&)N$O"YG0]-T(Y9P/ZN<_64T46E?3X$N\-8;A@'0Q!R".0+5),TKWO-7# (?
PAS(?R4>;IF-@3_VY0F!<BT8EJ@61QB.)!1A"?@Y, .<A]Y&PQQ> U%F$(.0@\AOH
P!7N*_399LMIC_Y[98;C>@%OSXQR^U=R8.<\!&.CW(%H/N*-!/WY(!<AI&C:I5$Q 
P?0J)(0##D7_SUN!*D$QOK,X")4V]M%?1/U[9AW&?O5B4$*>$7#V[%2>:P*?%'MQ8
PLH4I7*@E>I"?-%UQ>!F6P(&V+^\2IG:BKQ,XKUW#4./'&YW!+3\FRKJC?ML5>8+9
PU)71S'[%_P!OLH:2>0L&GD$LG*S#[6ZIB!U<+VVS*2;W6#I/^-R #\ =7,L)<QMM
PLT,7UC.=/L64@<JLG+D],2.Y+( R[GR&=XCOI'1&W0:-?GP =B.+P:,]35R=![<K
P+5L$5''30?'H<:.^6*9[/ZDZ7%ZUAN.CQ*QB][9]*X%GG&$6C,JU<T% 330/V>"N
P.2,X,(!%@D?BFM0LZ:2WJ'TRBXO7M$]9+**C\CMB:^+<*<SA^[IA_+.<A(,&X!0Q
P9/-O4WK7V7\V;F$5Z(/2"(>>+PQ>A$=^3XU9Q)Y+"(\)>/.B'OC<=XAXTDN)SUL/
PZ^EQ%?X*^1I\$+Q$-'WR4((B'I[U&0O\]9JBRDP/(#N(/\/"'(9P^:7-5+".)5SV
P,03DVI>KUZ%D>B=;7V+T4=)_![51>I<'%&*&*5ND_O^B^]E<V\P3N1&=I0NC)*N&
PIT5+=^*ZJS87^!,"?"#3>W=8GF D=!P1Q,+RY^^S5NP/3!S,VC(W/L=X3P#B3<AI
P0O(Y2,.F?$@\@D+7R7Y$0S%L_Y[HGM16[AR,%&O(.*.()=W3M]*\/1U\OBY0YJEW
P[^U'66JJ]AU)3S=AZO75 LQ(\:+F3>Z)*KA0'$-U-W02V63< -5&KR0+LF%QV8HJ
P;G6CZJ[^&Z?,% /)?3M//PUVZ45<ZA5R/?'.D0]N1,N'7+1-*JU:+R?,5M$$J&']
P%C*498IBS^(2'R)QVOIJ8@6 ?Y3N0M861:<\]?U#V)-05G_\=B8X'MO&#T53;[+'
PSJ!A"<NR#G*"^7M*YYP]/-+M4>F[LM^\V7FXK 03[@=R^I )#$))!((\'<6C6;"Z
PV4@>LJ+;0U2C1 ERIV0LK3HQ8UK][]0DQAJ@T>VWJ)/WUJATD:<:DGFVY"K1AA[)
PGE#/HWZ7(A2" PE;&E!7+(1NO1L'ZW]Y^T6UKR2W#T&[;J"A8YX12/-:1)M5RU=@
P+(2H<.3J PW2&]84ZUQ-U-VU(Z*2W/M2X8(:9EB53VD!3R]7)R0.RLY+:T<2^S?V
P!542$5[,?@);I,H-)#&7D>AF:7 )+UQ&=<_/YE4SF<S3Q],$ZIN7'>U,D=Q[!T>?
P$<&J(5.QO>& Z"?-7E8E4C0B'=2090!W-_E#Q/YH(F/>EU2^R):FA!NC;X\#1U\A
PH98^TAU;B@]E&DH8L-L-#4+5B])"5?R51>/^<@O6_=PINU%>=,$9\L[+1D:!6;@)
P%>)Z@AVY>T!4BP%X8@3?C/E/0Y)H^G2NJ\@?. 20G2B\XNMUT*HQU20PC<INYG_?
P]?J'V_;]R(8#CU@:B<S?!@@1$SL_5C@:"7;G/.[3.C[A,[\PF8JUX1]3KAAJ4EP*
P\E=E5FQC%[KOE_P&KBBF0O5#H32,&U4:@K(O4+QM^>0JF(16)>KCI81I!A1%5,)V
PS.\BN._0<_2\5V4S8?BL^?0?\E[2*=D+*JGS44K&UJ= 1L+E<HZ%VS?2AW2#_8C2
P3M3%/P7C=VP]='VC$I4!5^F6^F1Q23<2;R@+OR"9YMX\DX-MS/.(Q]H+QXIRI^K?
P$)YUYW/KQ*CFIL.JN&5'0WX:5G%2>*0X :D$!\FSMF.O1R^/>Y-*9VQZE;E3X)2;
P8?0N 68$]%NWH!].E0?"EN.FS<0C]7"YS!-3;8[Z\9U_M*"33Z"?90GD8W(_>WN:
P%"UJ$HWT/4*5)+;A(JNU^L.<>77PR<B)7:"67?+-J_3NVB#268S.#B]PZ\1RR'@0
PR5JT ?@N3_">T,;;GI;!7X,.ZZ=+W*/;J<M_I*D6FI.L#RQSFSU#6Y;S!E^)]Q-G
P2(1I2R\97+*)3>T)R74:VN\AT' [&>@O5(J1\D[>[/_<]ZLJW1W22:MD=OG83(8S
P#\9QVPGVO-?P81"D9< ;0<_V[+H5F.B0"8=16<H+?UY^O[L^\;@NE'CU\1&8SDL:
PU_8B+I,J2MAJ&I]R!1WI*9E_"S!JY:GX-0D?#'H+L<PYELSV-DK$MD.$CV,U4,&G
PUG Z3XQP"#*B3:8SWF75SC1063.9H81&KQSMU/(=+MF4&8S0!RG]E"^(;S@/^\M)
P!0[?VQAD-)9A4T7EC4;.&-WMHDVP<) C4D&%VF19:9V.-'?_(=O=0W.C?P!U*A"7
P;9R:J?<T+A]SC6WE>W./=]U58HS!,MAXF-JL/BRH\OY=[S*[R;@D53E$ !*9$UQA
PO7&?[)94_NSU-/H).S\@W-Z2_9@,2JFP<EAU]K&TU$4I]:;1X<X3^ B-S67555$4
P#]F+@/[<=UB[D.<"R$#>CR5M >Q_["ZSI#5Q!=*' I_.+7YJJ6?*AX%+>^5&<,^.
P<=?'-D1N+LG%95AR/=PXRGW?4:A4KTT!YYL+"SH\R$1EQ@ =^#PA+BF+T(TG9.;/
P!IB>:3WHT=G-2.$\6EBZMBR C>/(O23OL&R74"EJXBHU6#DA>"N#)V]4AN!XW^!R
P$"_%6\:P!CS81I-)7GFTZ%PF.:Z[NI7V=D6632(!Y)8N>Z2HPO].][Q) AFU.1BB
PZM-?M;JDOW@G^![/AZK.R^V*V1HPB@81AM,M%>7R5(MJZ#+0A>P8GE#9ZA$]6E"I
PB7;_H; D!6K[9SY X0XV-&%#^GZ_<:IO_]^1*(B3;DP;X:6,A>W"O3].:%6:>/SP
P VZ\K8[).@N>OYX_*G,IO.-PAS\?IXIA.F@-LC_+-#/>A^>(4?RTY2,:!YOA(%-Y
P?K]O:LKV>R1%QC0<0T(!_9B\KT#S+K+X4)/'-_.U$;@/,-1?A)LM1SV77E,84+RU
P$/TX<$)!C=M^'X&&PI,E@_3G)V+4F$3],/^M!=O[P1%Y6NEJM85^23\V-<[+.U,&
PJ:"-:_O>VU?H6H)Y-,"BII4-<>VEGR_$OCD9&U4]4:-=39PG9"RXPBOH+UDTO[O?
PF2 GMR-'36WY@Y P)*)JXR:#7'ZJOEE+\XJC4)=V!#B0<@C>B=3MX0G>_ P@/_J9
PMXS&/J7:?K.Y*HB](+.U3+ZX BCZE7UN>,H=[_M(%E/,-@< .VBY+E%)NN=9<*_M
P-<(-@4-_U;?\\];8J#XK62[YC<]R<C&;D8TY=YC^XUIIV]%9)D!V7N6T$2_XUA7C
P@B>#JDJ)PV*(V^]R3ERY%'3F.AB_C_PLD)-DUA]BZ_6I5[V] D A%K+7AZUOO [W
P!1V6::V:0$9W8+ZR^WV8%^<K*X!5+T]P2#,\Z7W6-;1J>VU$/%T<WO9]69[.@>RQ
P!03DR+#S@83OV;N7R*2_/-D'$,Q/3 <<OP&K>3U99[LPW'K":>_^*=J^S/60?C#]
PS($Z)XI.M >T+J-S1<3HRR5IE1*B0$N&4'0<%$#\/BQU8E+&-A[4>T=[M2KQ68]9
PQ6?U>(/;8(CKH*=9&MH%Z$Z [-V^L&ZZ+1^%3(DW_<:DKL=O(Y4>1$_J#_R$U'7&
P</V5Z!C,^XMZIQAA(MJ"X69C7YVN=$!.\IM2L>LD,+>P\Z'^-0]]B^#ND_ASEC)D
PYJ89]5'B.B)$+B<9!@/J!1(?7]J01E9$V8;Z'?="ZU] (%:P!Z#<B$OZO&!+S;NZ
P(K8PIHB"Q+%SUW@ %"I6V0(P!]CC636\)N3*KW[E, ,([:H6=@D4(=>ED4%S7 '>
PB]KJ(L./!MEHD$-#YQJ"!^=2:!6>R$]FV2T-HM,IH7UC&T6=Q@ .$0G?MGJ1$C(*
P!WBTP,?@.2:[KD=AVL].Q@9S\)L5S%[KL9HUD]TIIV30Y3_G2=X+-D@_%3R31^4O
P^_,+X]'Y9&1!&AN>'CY)/##;@5JPJ9B\7,.6J4+/#-0$_\$S]BQ$J/=%?_B"6;:%
PBL#AV,GX%I7087A\&9_-Z3P_SIQ]: M7"4J640?&I98Z*MJ++LSZT6]$S\?;^3O"
PQ +HF^Z+;>SX<^CR",[SXLDZ3(#!X"/G<Q%24$8I?=WV^=W7LWQ%\%WWG$1:X6RI
PN^Z2[B*3S+/Q91L.W\56;7C,)ZG6>:BXN7._E&9S2>Z2.?^JA(->##< ?M(@D1P[
P $UU O>92,YI/D1OD$L5P$G%!3Z%5;8N:B:<\V^QV3,U!W$A(_;WA%_GP;JD1,Q>
P 43,UKCZKYLRQ%<+*HG'KBFQ[/]_$'*F1_E&ZI5DA6BYP=@NX6.(1X9%\WQ'G:&?
P5%'TY87&O*Y;&95KUV"E@4*<R14#+8$$0\PEI)E6:%J'F$6^ N!$J&T[M2?B-X5Y
P[:QAUK>4M"))[<^["E(YSZ(35X3D-^P?W3H 1.S% JAE*@,8WL,"743%#QU/0C$/
P"/LO=$V?L@BW;:$3)*0TT,@L!^/>JJ\O-W.IKNH\&'^Z#;&0I("0$*6H6B]>3V3E
PQCA,7N/PQ7#5DR/:^.-(.W9%ZT59G#<??->BJMX-+O#/9QY+766M'&R?T.YU5<=^
P\/.P(3=^B<1;7\>(-A*S=S4KSH!\[#/G]>/) \N9#;][B11/(LPK78#;/1&J5HIA
PZ'/U:6L'?UI/U<CCC92I(4>1*,I;%-C4JU+!1Y)K#[_[  :S$(.NEV*GH(.8]5W+
P[[== C"M,5"!2L%495YJ/1O8-%!?IRC.?9V 7L6?R104$B$]38[&EH<_TW!%@^X]
P@V1V_CM"CE[BP[UWJ8A7[JFHKR'PJ.GJB0UQ1G?Q=@E '/77;+'$VGK$\U[3AY3N
P0!^RTR\]V6CH.K )4=Z7I0'KH<N5!UD<T_<#9-W%MU_T]1SE2YSFPB-@[4[GG.9K
PT$/)NI?J /Q4=E8F+ 5&R.W&N,A\$'C?MVCCJD/NQH4?$.FSD8*E,F5$JN$X)&=)
P]AU;1FXPJTG 6?TQFV;=%"E'['<XV7QYL>T@D3L"C/-8APVCP_"K3:**MI:-GXU0
PE3EVAMP9-V FURB6\'30>?ABRWK9DC*P-FI9LK=['EI;DS/=>&0Z)B?1RX+68RQU
PB#*\Q((_:=_%&(59DWVI?OK=9KB>&.'[ &W%1!(*8VE5KY+T=A![P7)'('M -LH>
PK2X#E*YQ.DK[V4,VM6MSCB:0HSS)A&SI !J9>6B)G9SCMXL1S4;^$(B]81B!HQXO
P>SZLOV5<T@-WHGC>MU:S;MC!5+)O\RLNK#R8EQJ75@6!%[F2$7\?L7,V+[TOHZT#
PQ!:!)2PTP*VS)FY.0UZ2)R[=\P@]*M=9MG4FZFTB@YAQB;DU\MSX_V"@ +>?%KI]
P5 G2KV; @]C9^(;^3',UV5Q.Q:</$,KQ++$48"?;HRJA85OQ5$U$\06F\7?.=3 2
PIJY=$%MO3SW$]@7L0A"I/RZ0,<XC;L# G[F1!H!?? 52WU8,H)1:#PVW1W/8!"D9
P)$?_B<+'(4SGW:+0XFDM[?]?X [<3'J6"[[.%IRE>(^V #S9_["\.(H8L]EA+SAV
P,>]A7E,JWT!Q%X:6O+[SO'[RX16R[UA\,.!@I1&>OZU,>.6X<ET%AJ]#HG+:8HA(
PR1:;56'Z\C(P+G-G^47H\7G,[>T_YPZO*NQC1=F2;8#.]98YB1ZG$T,OO.$C98^V
PROAQ@.\.1?+"=%!>]PUF+>D=8)1XGL L>@^5!P#*+<&[T"YUFR'\QJT<B'L RD*U
PC>L;PT5WJ'B"<[,=!?+0FSF@Z59,-<#HD7J-_.VEYME'LZ=7C;W5'[*%$ED,YIUN
P[.[I=@,).,9%/6E>=W'^ ^<5<;61"KSX1?<RB3"U ;+!NYLN[3LOD@?OBAT/$]P"
PUHF]'T@^22^B(B,EMD=+=ZAFVCRSHQ>L#\[1HLU[\=)X&;3O#@7NL_97!1[3V@%F
P)0*C4V$3!N!#/3<&6"0-@Y@I8U$GH&,D[$[^;/'LMX1#Y-18>L0!LIL@V>Q MYM8
PO8"F5RLO-S[01\;&I50LSE/++ EEC$102D>\<8ZKY:>X3*'>]ZOUH&(OZ<_&!.&#
P&=R!PYLPC*;XLA)&8*GI9#WZ^,FW/"^;%R39Q>T%&<:G/RO1>FHM!B0\K(!I!J[E
P_/"G$F>QD[F!V]'1U5W>-O.,4&'2'-8NH'GCEKA\_NH(BS;0@OR[8BY[_NUY4XH#
P6LN&JZ#<N00.V=^FM;@VYSH ]#Q[*B13)1,_S.76\OS@_^-/#Z6U/RA8#A(&=F:L
PXJ<6]G7RBFNE2K!^-9:?>&>4.8ZZU<]<&S/_T^0RS:D!]";\SC 'GW4%<,W>&[@V
P][?*YII9-QTJ2D82-.8,A;=C2F+1L^3S_$M'^QSN^(CPTW<Z-'+SC#5Q[',Z,]@:
P63$5:E"'P*@86Q]UM-]:+QAU)"[V189U#ANAQCXW^;8GEJ\%1R9OG]CP/OF1))VQ
PRZON5:-(OK21JEJ'+1V-G9D.A\-)\A!I=(^Y<]>3'9XGT_7='^#K^P!VE'=,TW5#
P'T:JJXCMZT))0M^Q@:H<H.&BV2 ])^U_?,S?#!:XWN^S\!UAMYWYC'+$.2;ER%/!
P;PI;W4W;TJ1'TWY_LA&KU1B5^+YF D=V+MP6VJVYC\G:A(.S\[GP?3$XEF^7OZ=$
PR.8YD9R^79+8BV=CEH,ZSS!H'2 ?.',O9@2561G'UOA(6O\PVN:KJ3SEEM%H$Z\^
P7>DC/U%:QNHD8E..I:5M,5JI?7+NN5'C[G4>_5H'9'*TT4!H(?_O\Y+T=+F^@'( 
P0P5N[-C9]SBI^;1**0UF2JDF:%1@II'WZ_:;FPO0GO7_D-$\TC'/39RZDZ!G_')3
P-Z/A#2XO<-D.-O=%(FONH)RY7-!RJX'00PAK<,UMM.9SS%[JNKMLH42W7K>_,=JV
P?53<#-F .N*T8$601P'SU&-T\YGG/>W%?<3]Y?#9AK-IBZ!;=?3W2G.10/SX_#*'
P;&TD*MEZ.I_R1Q<[OATZK0M5DE0(:]IW0=D)TE;3=-SHI@2<GH9X\(6Z>*)@]8#V
P8[9X[KYV.(/4;TB =A"_&]0N70J;NHO9SG!F^ ]]QZ*8@?.HN(DHP!^%$8UDJ34.
P]23X7S]!/Q<QIOG70@?2K4AO2^6N5#3.N5I[GPAHG3_,D;=FX;ZNS]0BS%="OSFZ
PZ1V85>*LF>$O]M^CWKLN&J'7*28=XI7R9E3'! L\]F'L=F4/EBY-[<?GE:WR[+D*
P!_5* H2I!]LV)<V6#0(X(@!UI8S2BM=EM #KYZH]0Y^ \)'JL2;G#YUH63@2AY:N
PP7!.VE+7)C<B>4<X_C0\HGSTWB]N0W@+-8VOAN@^XB6DB<8H0=36BAFM>&FE3FV.
P02LH#^(_*P5N)7TH$FP!K.F>;^W(.!]TSK$2$F9AI2;7[]/';BL@+&@+<W<OEP<1
PM18:AJU@3;#"+YP-='8(B?4G/O[#^Z817W45B)@6KU5D2,H<!, <0]9/R-A85-DS
P ,B]8=>,^ZSA[M1C(]J\+]"-FRI,]R$6[J@'=N$$\@[<Q2O/%H?(P;[MM>)IUU 8
PF, %/_UD>+V+USQ;G*'.:JG1H176;Q74'64^ZDA$):9Q1*4M^[EJ5.@$6%!R'@4B
PK1'1FP;, *8VTDK+ ETL7FGS^O('M(@P_2'3YA,-QVS?G!\R1_+[]T/GH4([)P<S
P:G4EP"4D(F?^+E_>]6,*VRTGQX2_LWHJQ7?AH@0>8&"PNO8)?]SPM%S;@2S[/$'%
P<##U'5#/TT5GUQFD4N1!T5@<,[W;AV@O]8RU#V-X6$I([!0,U;5=DWS;%IUC26%)
PV&2X1U!#L_E?_:TXG-N%H68MI_] )>Z?/,K,:KMB>-4U='9UL6/#Z@_DV)_5/>FG
P'".)TQ3E7;X=F+.%YV(?LVUM[GM7RD\_N'34E]0S0>M;)_!C_LT\R.DELM=@-D 5
P=''21/PQ@K[8CQA2LA3]YEA&7%P843XHWH\:4(OQ6M6=NPG^83:D?',<"C+]\W6W
P:;Q[L^DXI[<D> [>7OY2MWL@^L06MLZ5%OX>' 42A%N\7MVGA']9JQ+X%"RN5@JU
P(H O,C7+//6GW>B!12,J),A6@87.SJU_ ? H^JYT=Y3[_+0TBE"^J,2 *2-JK8-:
P7GS\I&'0+QIV -M*I''(PO"5!JF&G@,)'42-P9RDYZV.@GXV^5$DW$Y1N2FL1LKJ
PER]^2YS[<U:0F"D'?_REEBV\_.2FFIR>)VLMT#XJ:AK/8N>179NPJ$!]R%Y\*O\<
PK*&W5$]O //O<W>S/I=NX;[3V+%]4"O6,]M+7"#(;#3QGOH@?Q.>%-P"_W@L4+J/
PHV7Y;RACE9[<'+(V 8_*<TZ72=/CP>4BH$;"<C/DQ9E2B7K&\SAFBO&1,E6_.$L^
P3;/0)&R6-YVTA3Q@I)?LA"S!DU5[2J)HOS-F%47/@](Y7\?79L5M7:T2W'-@$T.K
PGABBB-MI'[UC&/X48*L+ZN-9RAK>2I*XK=[.SV>_$,H2%#*5R]*%]GX1IFFYT<IF
PTZ/=11ASIDAUD2,*ZLM"0(!8@W.+%-^Z;$W+X\S&Q"*5W%UKB4L=SN3@T^Z4<@%)
P]5_PM!IKS4>%O5M!M-T51.&/IX$OR)3KU:O.$IE_K_=[)**,G73'(O5,H@J'HRDY
P0@#&6%FXF [3Q@472OP&I70KZ L&:+TN,>II&(C)^8I^(7<E@%XWZC/,IR[7.JM:
PU9.G4SN'MJY!<SWI&^!/Z,B4"14 )"2YN+''/C9A;I<4>BAC<1"SNL0BQ X<#\ZA
PZ0=T;*TZF7DGPZTJKB8Q'QT 0P<A?&YQ +HZ;Y+!XL6M^SJ$T=J4WN7--H!9'KI#
P;CD)A9L 4*)V,+AY:$ZDZ'+=4#K+MXL; LLON^79YKWM%OO Y1] (XM^N# <@GR[
PKN<N%I&U419<O\2Z<J7&%4L44MYC@V:2Q;?FP'"V1?"Y>1)VP)32#Y4V,9/@%?2M
PVGD(6+'CC%GR,AKPH;+X"LC9N>VN'5/L=,@-D!^7PC!$Z'P.HVHLGE'F97JG4R]?
PDSU FH)9T-T49@#]Q!+G>S.I=5J=;L3:!FE%!S%//4+AQO2?V@F:1'Z!)\^@C3T/
P[6S  $A?<FVZ9ICE*Z-O[2NIR&FD[2&XT2D)@MGO$$HD_2K3'#HYX*<XR:O>6&9,
PUK3V_:YFN/8S[4TE+\)_ :YEUQGTEA!V?"1@Y19*VPS!-(X=N37BNH3*VE-@L;0G
P!33+XCOR+!2*$[V*O U1)-4YM2-,!\ A&\X-BVJAH7&M:2]43?:Z)V )4%SH6;'J
P5Y&;'S: "@]A0++7_3[?R+R;4;6@TXL$5E.42]7;!Z=1'?IUZOPY8?OAH4]I,[!F
P+.$"%SP\!*,J>D%RZ9H1K)R+/5!5;?$+HGTUKN/+'64>,O&GU>\#UD6^<.H'*4E(
P/*X^@>:*]<\?N:35TT1FX;)T+RD&9[): ?W[@OWD)]%0=V<#%+NAM+F%0UGZ/485
P"N'!D9-M98?.EU_7J9Q(D0O=W6F3Z*=I9^75BH+1;E2(J4X5P79][R'B=&._[Z>I
PA-%5?A*'/"]0N\M:)P&XFF:U_S)3(I*F7_ 0F8U#-(> I3/W%J1RH>B?]LX.:G=V
P()V"O*\"QIW2Z\2,U@=Y-C\9TS!"G[/K%^]ULXQ\LEIS#EJH+PCZ&!8@_2R;8>DV
PU.J2X/?9)#T)=W^)GH@:P!([?H13J_ <F"T[J!GN.R/QT_*WR^.OI'6O?X, ><?/
P^IT&G.3##8UP!BQ*$@>ZI;HSN-N2<AX,/S8LL.(PC0TOUM:*]$E#.L;5#Z\%M4(%
PAC5^7#52/ [,X#XR1TDX/L.OT(&$,;L7GH5*NT7BSC<19+.W0RY:JJ27H?*Q$\E9
PA)O5,&>4:_[.$K2 A+LFDC_139VW$7SZE7B0$-I&C(^;BX,TI?6+ IJ!J$I1A26=
P+<6[+*]_#UTCA+ZHB4"D6%.D'Z)(GH0&%#E#ZBR 7/8["T6=NI9CV$Y(4PU4J??!
P$L%LB"L<2)P1V5$J5G3GFOR!OW4PI9#.<MW;B2OW7 T]6/#W$G?_! -CGIMAIBT@
PUZ>$ERY0;I5U6S<9NPKNRB'8@0 FZW1U1VOA2T)V%0&@A>!Z9@ DVB&$F/Q)!<Z4
P%^E R\,J$"VR#2GA@TT<>P';Z<PFG4'K0[I<S/"FOO50!82^L/2W@8^U=A7@O?P(
PE?,%S<M AY#JMRF.=*4Y@PK+NJ[>)0=B@I"2U$LDL=0E4A5;_AU_W[8YR4YD L#!
PZEUW$;=%4*2!1D%U<(7WK*;F+/B!JA[O'6SO[*3X)8,1\V)53#6H%XH/%9Q2I=)M
P &]'1YXE?YL[75E?4:@*:CI$Q=0;!ED('3JZ!PJG?YN.$&V3FO>SK!:;S!=[H(7P
PM9+F.J76*.2'C<S SS&P77676QR"B+ES<%R"L/"5K4X5U8<9&E#!*-"TKDG>S)@5
P>IPO%*U?(*VZ3)'Z'$KS1\SX0]IQ9DS<IHG-)YA/K52GNA'9/%\"[-"\5<9VQ<9F
PA"N-/&*P;&M;1:<Q?D]H9M^@DH"&3W\9L8&L@%WN"FH5*IB&)IY+U7A(0J^P6&7)
PT/YO-]S',7?37JCV> N0R(TI2H)7%0-T+H\^&NIV2(4,MXK\S65/L2FGK X?&U^$
PT"7A#'"J_W806JA^>0S?5MM)NE^]7Q;$$9M:!&QIN#GYK2GIU&1;M8@-'ARKT5!2
P==X!';V1]+G%8'RZZB?_0K>8BM\$\%M9S%8OU-S\[ECZ21?S3C+P BI0"N*!W]%G
P 3U5!YC;>7PB:LL\_O>2DP;'X2&,!-8,KBX%BU'6YV([1+65E0N-6HSBH%5_5"P+
P_+]^\12/;&H>#DMYW:0QT%XYGNH@N,PFTK(+JP0R82Q-9)J@_N=#!J(%C4[@3:9G
PT/Z 9PPNIWD$JJEYL\VP)UK7OWH"YZQP('I+!'QEFOTKZ.Y[8&?K95MNC8Y"=:FU
PM/.EG FHSV;ZQC_Y[](84!GT> 0*XB.H94%=;15PHJD"NK(4 TMHKZVBJJ@5-3 /
P^#.6-FY\]:?B+_+?R,0NW:?XK/P\MUI\\"&B*%)2MVU"#< %@0(B^!;%I7A\S:#W
P4:5(PTX^'7E_?:!P#:M\W.VIM.R/J,I#V_-:2UM]PX'*B_VOA>CF*0PV3$L-XBZ)
P<K)6PFCJ*S*A/F_;!6"\9#]HZDTI&@=!WQ+0LTLNBQYHWG&.Q)K-@\<^X5NEI"/8
PH"*04E]Q ]1]/76H/5.$<\[ _)0;C1FA-9B4,'E80RUZL(PT-2A].D$X'LQ5C8K^
P];IJ,Y3S#EW/*U)]$G;2PIF<)/NO=FV4X99_5VGHW@#_VC/$%]].^LA\A/.WH1KK
PVE9O2X=K7<F5+QJ?.L/_@CL,^3PQ+IR;QM^+X\0"Y,7!$I(\>Y%C!NKT:'C0U3B(
P 7F=?CG%)<[*;A4NP*#5"(,6?*CDI.)U!^8L<]DJ)QPO??;TFG$"#^;!2W(J-A%-
P^&&)9>5"AGJ^:U7G)5,3DP;4H%MA6AMF6C(1Z@T>%/"S?[95<HAX7?.]P/W'-H@#
PD:Y^$NZD0EWL;9!R="NKY8:/5/E#9+VC'9JCG5JN4E#H@NBF>ATGGH [G"EYJV!5
PUXJCJ/M\D]'#MW\VP'+$2%:=RQKI]'T'"QZ)XJ_](L"!#MK77;W!) &\-_R1E49J
PKS5IKH2N6:&N,PN]TGRJU/9]R5/COPS J9)]YD*?FE+\SC\DZX"Y4!W9KY>>QNU;
P5C)3RP?V% (/?K_>)$NMKOQ8C8F@-=#ZQT4UCJ0C[W!A6J91.6/_YIU/-94,]U6H
P2X6O?J/1O<W*[-+-K %@*XL+X[6,ZB9SDW'F0IPE=;>H"?;L@/GFBV6JDGS3P*+_
P9/"GIP!BDE\K3XU0G"6DC?PT=&'P;]/9WT5%?#:TN%@A_S>K''G0=E QD($FG;:^
P(?G"['!LZL"2)1?[=F;[6V:TK'+.&#_I E 3TLT^N.OL'Y8=)G;'H5F_;;W2;'HN
P53Z@O9HRRRLWB3NN39G$?9I/O27 H.ZE[&HN&?4"-G(\<*&WU<H?OBJF8SYD"ON)
P UEYC/4K"269#T%0QVYY8LTL,EHJ3ZA*7'L+.+_+[;R[:]\-D_,B;&"4Z@JP_Y?L
P"MAFDG_[3/*Q_:S#S<-HV$&+_?J6A6K1,#I#\-YA9^98 S6B5Y/#N1&,YR1%4"]7
P9'+\K!JD](X\;&N.2+Q3;:C8" )JK'GL=N*\S4<V#KR[?KKIWQ,!!!.2,<Q,40MF
P/]QN+5SAU0H)W#/ K*F@2CB-V.Y28??';P[/*&4$2KX) 6!^>'Q<RA<]<=6MVV>\
PBO7KT3J_Z%R#C"ZA.7[\16MV ,6Q5K]4UMJ2PCS:SZH,\Q@Y"RDQ 3^P<7.>R^\W
P"Y?/\KF!8UW]T!.8SU3HU&386)NR!L]U])C/B3[KUS_Z+1PS=(Q?(C^M:]UH@Y<\
PKS.#DM! X*.GXJ"0H^IOSY7>EU$,.@1GQ933P<NHO"=&_^FRI0M^I"HC>WZ(L@R)
P.&4F-&J/VWV?MUM8-G.^@"_2FF.JGR$HB1'6;;3JY>B* 0L1T.W9,*-]!M0DU07+
PW\?P/W5A[PY;]18"WP.#3KGN^@V&<S3E#VK$B3+%D+!Z:.$C[].;8AI90KQ)TS^%
P]Z\;/U7DD7BJ2G?HJ9&NP6LIF^2V-D,ZQ@2)!LW%FC+_DQ$@OI(3OP" F,$6E3VB
PK%M'=,1.63/J%MF=&$%@(C#E UU-E.5/<\Z3NQ[N^M%;&2(*;*!PUG63#FJXPK7Q
P;L(T6I&J^H7FD^71_7\#$0AGR7C,U%/$87.=:"B:[N"]"P17.W?V6\/@F/*UXGK3
P>(RJ)^>L4%-I(4K*;1],"0S'THTG2)N_%=:F.^4#-!4$/:<,K68":'JE>)* <=OL
P84<CC; ^&\@A80UYEI,8;G""M*XQOG$>7]I@6J',5#]VW)C_)"AR ;W:O/VJ7-_D
PBPA%VU-T)??K[.^:LX94RZ>")+,3\37!+G'@(A<:4.5[9^.D@&"C!X_E"G@WS@=D
P,]J[%@!7NCSKS)3QZLG,*-<U%CLY!<K5^F%8"-)570KC PWC@;C9LS 2:T1%LZ8,
PER,%.>971GRORIWWJC%DH0!\00"H^)=);*"2E5.C6S<6!!KIA "ALA;;U-ETZK^>
P,2&W'LT3P6T'^(K45Y@Q!.<Q@NZ&,U,W"=/KR-Q"^YAG+L'G_\O3H==!B/G$#S_L
P73JQI6(-VS^A?5'+/K3+;I+DL9.HA!KJ:>G0E<\3-UVH]+UR"X/N.7>4V/H?R2>0
P[2Q"C@()61YTE7S=0AEH:$N<_ 5J-51#WNCC+<TB)I2+'^VP\.OQL6F(](C:0C._
PL?OEF[Y#UN1L.J)XV81@5.![/FS6.$0&A>JJ0#;E'+[[Q:N]GP/%HK@,_>A!L>UG
PY^?_GE1FH_Y:YN<%WTJ-DTPO? \%&$(SP;ATE#BK^*'BG=^UC3/JL_=@0/7:<O[N
P9."$SWY#;O1P%TBV@3__4C8G7DO2BZ5M%:T,!J1R(TI:#8OI>4=;_6:Q,UD$L[[A
P(59[@R2KO-$BAQ\J4!_S'1X&^WLOE^(T9-P0#\$3.&<1*O;L8 J]/LT&X\S1"-7>
P7QI915L!* QQ^'V3___U/.-;0T29%P4.D1^XVG- V+9?>6^)Q*[1\ /[47[ ";? 
P95Z':([P'YMV>S7'/QT;EU1]N$X@.(^9CH35)<I7+7E9%\L^BJVT>=N-^/ 95Q ]
PS.AWALJ+HUCJE0GGX#T&*%G51S#ML%]?^1G9'T0Z"KS>5#G.;R_"%1;DGU*9%&*P
PM9U?TSM[G%CZE9+2.M8N!%MS=BK-CC9*I=;I[(%A&1]!"^K6J:8T&V>Z[^J3UJ[T
PXL?NB$F #";++/ \53_^:38A.LX/V5<O)Z7GLV*J<8G'C<35HCPE,C0]:3R1*<??
PX1..-B;7L;DYXWQ@\37PFJ<HP#T&TJN-.G=-DZO;8];UL0^OT+IMOD&2UYXNTR)Q
PD'U9Z2/FC2-D%,:#-?9-,>1OXIB4_D&>-N])CV%&T):$Y_)Z^]AVF':*VIT0%A]^
P!U:Q6?QTYQZ!ZLW[?'2J-7<UNV5>;K#;_:_PAWV[[SJH@<9\V[])WF7Q[UND?H0L
P:@DNN+;X6+6TXYFCS]\9//A6<!H+I>R A?F<BMJ]]OLM8S:E@1QW8RQ_J\%$[T',
P+4:WB+?7_AA:AVE@]FMM)NJR:A"/DGPO7)6OEO+_#[2)81E,_CKW@*Q$\-Y#_BVM
P^H:(3F%X!WF6X06]1=_LO%!5Q)/C*-#R1&\'TF=6/(T[*@W*>3J4IPCCR5'6 S2.
PB]WB$O.T::<JJ3^<,5R2]V7D5VW!9NA&D2!9_G);YAH"F+_IC )%)08!S2)P_DC@
P56:>@KG VN7F3N^)=\ CNH_R8MP^6K?-*DA['O21@%>2"KBM"4<M$I=IAR(A-<.-
PL*X/ELNGB.R[3 V">KD,*<4&ZK/*;%&I "GH!#\I*(*X1#)'<0(WPQA*0]!0\A(Z
P6F!F:'^((RR"TI*? K4^0+N!B8ON4JX^^>FM)U#W[3#U>>XS[NRLN]/I+WUE$6K0
PE+;RP6"TE'F^ J+$>09DO/<H#70071XY/9V+^K]/KJ7(I)1,*EO=DI+)I%PA<X%#
PYN_U*5$/>CX;Z);#O8XY\)EK'@;5T)%Y\ _3[RZ#.&/:OJ K/94 7^ W[$T$C50_
P5=?%<7-?+#RWFK;/HW_U4IB<809"\LB=N'#;M&6HJ'UY[C>9Q1FL@UO8[6?[,JX8
P[&Q:5 7YK9C^QJ15(KHAZ;T]MR;?>?3]R#V&#!JVV0[MC(!ETX"ZH#8PV&B0C$"*
PJT\$# 8I<(=4G4S^<6Q8' 8-D#(UY7/AF4+6<)<@3]!N56"\.JH[RJ%/OT7=:QTL
PIB'\TRHRT&FE<4]N7UE%5/J7."H7/ GU#%TF,1%>DGBYXIZB+5$)1^7V@ZZ,@$=6
P]?G+"\Y9_*Z::&NE'R%6T/O<]\?X8F Z$,J?F[A$\=0"N2;TCWG=\UTHQ1,IH.JB
PY[T+^&ZUSE?YCSIN8IP>YS+,&J>^O"/-9%D M(4>O32KGR!2!3>L"RD=G+?GCS[C
PY7H=,E33R9\SKB%U;W4T+B%6X_%4&R;],(LIK$9'<75'%^=T#<JY6@9)&C,/+GB5
P.,C#:E66;-S!=.T$NO,%SKCE6E-'&7D9R1H(U>G>6!]Q/+J3[\;#J1QN9%TTGW8*
PG/I$_,M.MN;_"K=NHZ>P$Z'C\5D2G-7)B_%]+C;W%E$!L12:&R,K?5@U<3"O, R'
P$7PL9.J"':F [HJQFM?BI(UVX1WB'@:YVE&WP*[J&+4XQ9)S)A<!C+B),$XC@#3@
P\;_@E7H:U0!.<1TB=\^;1U!,J00Y_B9P\"*R?LR,$WG1PU9%(GE/6X3%][_Y@RRQ
PS?LKM7"!>[X<+UJ_"86ARH3 XFZ;ZEQT4K/1G'1+Y* *-)F$6MRYN5/LS$U#0_AJ
PE5-4)L@ICUUIE5JSQ<JB.KRINB\TVAK%YEU26^6HS'((B'1%D-[PE2N J6W@<1N$
PQA6%5GE4673N1F_V+DUBIT!7Q];% X(SOXL (&<*!:E::"5M):Z6/?G%\##MKTTE
P4GRF["B.JOJ(FD8^[R81_+M$_C)AA.]RMH $$\!:3CH6/E^$.)-W#KD2L-.FV8(E
P.0EH_FAL<V\0*Q 6)'.NK('NI@GH,:P"+/#ENU=194N3K-O^4SI 9]892<*Q Z^8
PU1^[R?"/9QPLIM_I<$%EJ$\V+KVJ:\"'%?4)P TW-7S4LDJ-7(%Y-]Q2/&@M\O/P
POJQ]="XE?WP!%B]%+LNMDF"'7F/@AL,;?2*:H[$'K/V:\ S4O !78Q!>Y:=FQ[1W
P!(VA(_66C=COT9+ QF8Z; JFSV?<W2G[!)*&89/SPUW9B0GU&TBQ@\-?GOW>3&B#
P#(ZIP? N%00=B_,MZ\?Z^A:F$X3]C*B,N6FV(/.M^WH:Z4Q49F\0A#5U?4QS4VV?
P^)D:LW9DSQ@_^0;FNT!43Y^Z2KG,G<K3::,E2M_7L L3;DD_:X>D1$F/$[>H(Q&>
P]!(Z=R=63 :7ZT1'_]@ELI,K5RQ/<CYI(9GI.PRQ.HVR]NI\4DC")RS%*9-:N-EG
P:;CN]!\MQY"%N=_$G];^ZD,E]9W[8'H>_(V'F&9SN:^Y6<3V#S4SKNXQVB10_2SX
P!,1:X;V<1 )3JNDX/'LGT*JR6YLC.9E!&H>2=)5$A]L09!0D(N[KK!=6XD>#/.V4
PM5N59/A([L_'3D 0'",V28'LYX*0B#02T;J1'7=_!B&$:K8YC;L(^XIE*%<U=,0'
PSGD8X*!+6N_,^))E*VQ34RYT=*JWFP-=#=VP_L#HG=G0X[.P)%:K\VW4'6S1IN3=
P.4R%/-3924%@2H(4#(,KX[(UD?]+;ZX+\+%45>%)P#7?-/YK-%(M?WM\KX2N$^O-
PE2Z=&Q&Z*OX</SZ:I:DO3LT>Q[]A,0ZY;G-\<XSEZU:&7&\0ZB'RVF2 -XH=E\$?
P=.I60COKN=M #N+?2C9P4M_+YEF2&-C8=K8AHJ0Z8XHA+E:ATZVJPL=SK!"2 <A%
P(-[-(O;MKGJB"?6X'U9Q__- ,*;FX0L#N^DB?E%LV6=)C)7^,?,(&']V.J9Y?"5@
PB>[KI:(E4MD,B 5L;S8A9 S/\2$H.=V+U0U\X<C=BMS1UU:!IF2B.,$OIW+>](HC
P^MSE(.8C*\V+*F+2,I<E?QB%R\H> D8L>+1E@S6?I'/%]SF0<6)\Q4<+%1!(/<$+
PP\ '=_7$K>QCNY=(W4LKG9;*8$%*AVM 3E8LQ;K$OMEKF#<$G[E![(>,B7H)&<2O
PUNA]WV7@\/@"=L&H0Y1P!<OJ!.@/GW22+?-T9&YJSM'("631AX[SQ!S'^G!!##UV
P<AO/9C$_UH3HA8_3,J_ (V]5_=Q7[B0,4IO<(JQJ\*_PF$HMTGFJ]-?GYD9A<7<3
PEW4;U?[)%=0QEH>FMY"H0B?*04Q&W':MXMFI6]CWE-K>8+N[O)9[? S<0H4\_<.-
PFQ<:0P'-B8YYTSLK:?[Y!]2AUVDT6^TKVUWG_O2RC?8XL<%F/(; \L@7YF1'_$>5
P7(L%"S!C"$76$KFAHI<6]C<(R_O^83@])K]][]Q<?.GBZR&83*O&;Z@S)O+"C7$,
PIX#;\MG X)>VTYO;6X6=G-7S'H_H#U0?X@T8/F+VN&A==A']>^YA.V3+@[F;\4K?
P#:YM;B^AIBKH87S^0K,9U_12V>LH,@/IG(H-?MK*I"N@L-DN3#R2# @=,>[#&IKM
P7&[['DQE ;+<Z%KT%TS^]M$[)>!F^OL;(;$U8L?_?\GI^D7ZU6:L*=*0KOYIPS2A
P?K\\9/F-KS50XK='%O^9V\A>\8:%7SN<PDN+V:_#Q)Z>EA$I(_','5VO+LK?3OD%
P]F>62V;'(2G=)O0V\?1F&S*OZ;A9?CT9<VE/)C"52J#<.6T/)U3]^(%?YU&^'4&R
P3BI53AR/X$3&X7#F9,$VX_UF;6[B5<VD=YVS52 ERI;->+G8A&,@S@4\HY 2D+U2
PKCL12S0C0N>%Q4#>RWH6?ONB%_IN$N1R)%/P=[-< $&58,PZ"N<S 9KH@!P;)(@1
PRM3C)HYKD@G9?=%B)!MW$[8=F S$,HS!M+7DA.\# .$M[_$1TRPI:U::$P@EH5("
PG VS:F14>LN' :GJF>_GEYL_J(E,#Y?BAD[BR>:.T^UK]-V(:H4!?C%ZXM?0H0'3
PQ2Q")WDGW@?US),ZVM)G#)U<Y.=82S\//MD5_4:BY'*TT;A0P).5&FAJ]NCR*)5>
PY5K-!M1J/AL6X12E8UN=L"B7ASF?9.-4H(VJ@I 2I;G;A-S'88T;D?GJ8=WT=_#/
PUAX('K!Q1JV@B3(2N_WA>OPXU@5:%[#6@H?Q3$JT*"6$VWD.2W0+:@'^]W+J?@C]
P=0@,XM\]\O<5[N%W0000 HZZ,WHCNRUJ;?;&-C/@P@ZC&['7X("EU7K1"E'(L3&Y
P]=\'.*FDO"QQXE2,6_S3/8F\N)X8"B5C$,MZQWM45BT\2A]ROH6F09D)V]"EPJTW
P,>$1G]DYO3 MZ*NR.U/JKX![\++YS7X@_5\$S]Q$G&:9Y%VGOOPZ%>OY!F;4];FG
P5($[M<),Q\BN3TQ]CQZNH-GVE&1L,FD?K;4E +21'Q<#=_&TJV$$NA\.<U'O&[UN
PA )X&;B>!MA((#%95Q':(#+8*IU,')D[I' ,8O$)S3"^+KV_IB2>?/?%B>XX1&#P
P]X_1XL;$N4YO,5A.3W6^3IBBHH&OE&S%Y_K*S<&(U4-[]5<KC"2)AOT_-N;-CT!&
P5$/V?9I]R+SC;XNNA"+\83,4/RNC1V@]>]=Y$9(QU(*5?XM%5R0/X:,R)%#EV,MB
PVQE!Q#.EH&LGB2H<,& 9D);5L$AMG56X:S4'%=H,]>[2PH@.34T3,"\$D?Q1K#C*
PB$0A!_*H73R]!G*=>&D*3I#3\ IC(=]\SK!^.Q(QO[-(NK61=Y+LF9(AR'%-T)*?
PI(W<Z>:2REO&LE";F/D=ZI0QB#BVX).719CS-]M.*SJ/;X]4 62P\J Y*&6^.-O)
P6A=-\J?@(+0I6@"%-J\@[HS;5L1W;^=) 4J^XNYE=X9\R"<-_8NH?MNR7834-*,:
P[Y2#:@NB4K,Y">P$;-S+F:P\H*,LPD!']\BHXKA<*L_X[(1N4R/VCUX1.:[67.^-
P&RA@77FN"SU'?X'+R?7VLF@Y"OAS:QT[LED^7]%AXO+,$9R\FQ;JA"QD7;_=WUK/
P.'L5=_(E"&)A12N;)CN^7S76;!&9Q6/&G^86=*+$=JRU+-VZ)\')M3TX 55SB<HH
P8GK8)+B?'QT+$$'6#!$"&HHNXCG>BZ_2EHM&^R97J!&86%&C]8&^E(($@+K9JI6L
P%FNA&%&KF ,EF%@ZX-]9ZSU6Y"< )",'2\NI"$JUC##]LTW?[,^ OK8Z&/WP=."&
P$-MK@*:VML 0B')%U]M_:-;=X;C]DT#V+H"CS"E?:+3D&G9*>NTI(*$UI\8/]1VT
PL%=,YEE3S?-&H83U/IC.<S5TI]67H8RF3M8K9!2>LKKD$'@!I4*82<)MBR;H#/,I
P@$I] <05?]7634'\:W9CK3CE58>J]%FUH']M&AP$ (E^\L=0!3>T4MA%A:NEX5=?
PZG)P0%???IJCFQA?"V(%\K<&^*.ZD$82N\V6+LO03\P\$VOA (M#&( U:67VT^]<
P\^4ZG$:OE.5#T-^X92X\\/TUD84BM,<=%_KI\L0R8"X;/&O1(HNC<6S!(R1*2N_T
P,MX]0$%605#)'0</0F8]2?I\0]9@BU:L#RY)%;N6BV?"CHI'%:,<KK,XB]FT)M<=
P.<X]$^-;GA?#+?C0_P'CX.!=^9^4([?SXOQ>V9M98*@F5$DKAE'X4WI0\H&<:P_A
PDWLW/%%L-2>:'ZJY18^/1E(2!9DK=[SM_@E$P;>2.R^R@#8O&\*RD"@).4&+#@9V
PCLMN)ZOGH/NSZP\A:+PKCK)?/R-\N*Z#$JE*Y=0TDBCX*L*%*C17ICR[5+<!-"(B
P[_M$JMR32@$K:?=D_'1L!0J_8GXWN^=;5JPX40 \H*FJQTL=54LG1@M-$1?Y,J5*
PUR^P_KQ0 S';2C*@(Q;*(5T&S@8=@:1 .3X\#I5>>YAA%W4 :-+0R4_<@S32SK$:
P]&^(LI/'-UD9'Z/DQX9F10[=@T.LV:Q'4]\AEGA36E)M 9:9(/"I;WAIZ/A?'$N(
P-GIT($UFXFD9E+4'<OX'L $LH\U63XQ+K+8-0*X<3NFD"27++NYU&!#<;2'F81U$
P^ F?;"#W:\+X/:L<^0T6UL-CL4K""5G5TO6=4#7OT)_02&O1:7-PBKUL%1M_CNFH
PVM=.Q>WK)>T8F&[R38^D(3J&/'%<,3JP4K1LV><+NR=XW_VG.MHE/#>H-E6-;C"F
P"!( R6DU4@UOA4IB#"7_HBX6%2B[5AQC *K\WSO[(DH5W&ZBF_+YU]=G /1W21@P
P5*Q"*H+H/310133)@9-*8+W?L2C75)O"]>=WL*!H??.AF8<V"!,LF,6='JR#A/#<
P&K1G^,^=9=6B456N\),S^$N^JBH3H5V KN06L2\7+56]PR*]Q^JU.Q121<?2!=F.
PL9J&*-H"Z6GP\L%-TR)P2Z0O-8K0//!59$M%0XO_B@%=[=ZM C));.9*WKZDX***
PBNM[)0P/5+$!M9UPZ1Q@M4UO6)EC6NF.(IKVDTRPJG\AII,(8C;)WW-;ONZ!A[Z@
P?#4H?3"Z.XT:4/M-B*8WG-NR_R#2J1"([P:@S;I![-Y-B VA!GX9+Z[6D8HMI N<
P84 ]_S:.%K?:V3B".9&4PAJ:?QY5E"(!:W*'CFDX"Q@"YK]T\H'W)&R716-4%3A"
PJ%!IE)=<W/9("-P^*+"TPGSY5')7;MKYVW5R5L=>929]I6+_L;4_-NOH?+=%=HR)
P>@"],F?>2U**_0I9_!!68\H2?H=6U6:#"53/Y0Z?NK:VL(51X7FV$PE8JF8O)GK"
PRY+6-Y6>B%024C\3CS:4]9VUBML]V]Q9#XS5$NGW\P-\Q<!':.1T)'(B0O$0N239
P_]A&GW<(RIUG'+$$7OS[[RMR@N"(O0M*9V7)$?^3EIKPK*M65@@R%A0 REZ/A+@R
P]]G1447^-^5^,R.)1TOIO!^*V?T]99R'I!/&V5TB<ISUN'#V@2/C$49I1"QIJFKJ
P>$YQV5\,N!K7FI%=D(9GZ,9?_#&).12_&QJ:37IQB754-Q_M[FMXE^W!K-I8"TM,
PQ;WD,,Q&ZF$8T)D)V/='SU5&<$3Z)%]I,'&QP X;Z3#%;D 3.7VU5F*4('9U_Q0F
PPA4FO1HECJ&N>@;@/RM%O!DY1+?Y?)]X1]^Z$$/SV+NS"U#N?X)?U;T^H,A>(M$#
P6-MV1?5C%TU6$,62EGB^8N&\;AUJH2/:BEM%ZPUF>CY\F(J;!XEP"'?5_ +E_E'F
P:MQHS>7+QUZ"Y73VPWY<B1>5-8-Q)'=GM;V(SPI2^ZOFJ]\":ZW243NC99?S^UKJ
PHQW:U:#'5U:-!,9U]\2+QH*+ASK4H;..E,):&TBQ]-6B1V#"=R1N<^"-%0(.L-^G
P>N5+BFSSK [+A6R3(2K]\T0ZA?GCR]B.<X=Y1-L^?,%\ZIY&O(WF',<9^CKU,,6U
PA>=''\T&<W:'8;LO#84EW6YW@P<,"/L"N+!IF4WQ\J,U>%X0[ 3L,J=ND9/,$)@S
PDJ8GDIC+C+M,VR5_.I,!#7)F>& \UW,D3P]6]RWKDO V/PIUHLC)-GP'?88E+ L/
PD8E[S:4P"&,@F3LQF9_ZUY]L-*:#L:MY05%[JUL04F$(T34B17G\MQ\-AJP?SEI<
P\W['X,@IIIP',Z;]'3J^[^53F$;#99KK_!S6-831[L"J1DO ]97U6N[2C\] Y9G6
P2Y)4$ DM?S!INRH\GH$[2R[SV+M@' *5T.N:L/0>4ZF,.SGI,W$>=-,J%D"4(\J]
P@,DM(5,-Q8^[X@3D\4GN$!=I_<Y:VO8./=&Q%\2]2#MXWIP:/."ZII:O,O'^2;NF
P]"]8<_$VU/#N;'N(!H(@V_/+U@8W.DMUSLYQ?P?KT722!;H1SH%[\(N6"\Z*RIIA
P%:UH:,H.*&6#HR7_J&7,T-?LU>0X&7@*'_^MDHU[['$(NQ& ?I7Z!=VJ@]Q9ZIT0
P$NXA;8#]X-V9T@RBB!E7EKYW^KKC$$]>1B.35ROSLS'>!E#CG5)Q3+KI\MIX"@@.
PVND@U@<6L3V/%H>T\Q!6X+,'7OBVH<!R4FBOL-8%@XEAW5J(R02M&2\E0K4R1NK 
P<XV;*YU;6T+\75P$];U4;?Q^J=+>LV#?HR;DQSQL&2,+"4Y=2_:^Q1+Z,2]C]:W:
P@:SN'\Q9\O.$G5,E(2'"YFUL&(W"O[UIU"X-!'X1,J!-?D^9<7.C>>H"%^T_PA4&
P+,W/Y40PC%KS.5QIHK\P'ND+,C<8)/N$Z. A&[=MZ9ZRF"EAN80O>&"Q!7H2**5+
P 9A;E</5[('XLS]?A(  Q'73YY.9HN@P?,EFUI]60*GHCNV2/CQ)G!^KF&,35+WI
PFF37W5;OP#GC/ #!MV78 G#O$L (.)JKC2JL^6\.X7UD9!BD#R$3FXPS;&(8H O_
PR2[,6ID"U[71C%P^VP;9V%0$=Q(8?O+3-@E4^?7]N=H0_Q6M#.N=9A4Y05MW?J@2
PH,9=1Y8TP-HIKT"#\'YD8ATKU[$69]4[;2=]M-,QU<=:2ME+U'+T"YG9 ;8Z-U@ 
P(!GK.[BLT$6(G600)$(=@!@59XGNAP$T_OG=E-[,OYM?B-JS];0SU GC?-47PKPX
PT$$1:& 3+@ESRQ<43:G'OG&9==K"[1W6_J<#(Q92X6YJO4CC-2GUT^W+!Q_]BFT$
P>F@^QF"R^G.Q<3VWB-N]J\:-V9411]1K#/1M\)H4 6S+:BDRP%T<:!VJ2HI5K_P0
P07:IA[16%'#(\'$6;C,&K6SJZ88+PH/4V\C]R;'ZD@)N>L ,,/K=R]PU1O=54*+R
PPJ7IYPDJUBRI4$Z?%IW'ULI:!'(GS*<X?54TNSV%5^*-P6G32HR6WT7B;!BQA35[
PW>*TBLEC7<6H3A*CFG+:4&33;"("RZ53/R=V!''#8'5*?^X"8,@X-3+/A7<_]>4-
PO'K@U=Z3K!S*?W%+?$M:_L4[J5!_&F&$L!>SZ+J*9:J&WYBQ"4L HM==*]6%0J'@
P9<O3G+3I.-&#NW  T/&FB.GNVM"FV=$9^<5C"89NM.G],5U"6>SH#S(HYG'C%3")
PL;'C02%!"]'/MZR2:3O(^79H+6XVP45 K\S'2QY8OP60S(/Q#9("ONZ56YTKJ"E#
PG0+[O3)EE']53$8O0@U(2[U#Z0KH26I24:<J56(\OQF$"%W??8!W\)B_B05[P!7F
P-^#NPM(E*NO-;=97/0?6/Y3T1C;\H/)7ZIDX 8)TS99C8$\8+_[7C55*^PB@V)Y2
P-MW$N,-:O1RL%L;LVV:L_28]V%$*B57F7$U\?G'#X7U,J /8(=]:%6DWF;)K4D!V
P^XKY3NF-M":+!1+<PJ)6D7-ZB<*34".&,QP=33.'69]',;*X/@8?*X,*'O2^5K5V
PNX3\A^P:CAJO>VY6F*OPC/S\X"<!G_CCMO!C%2 OCN5O%MA49+60!+'&+$DH$?3Y
PYI.^R8[,+B\+UO#?NC\.Q#B BSB*N&5LKLH3&11L@;^LN>.O-!/QKXVLN!!SY0UO
PH'5J]F%*6@]-.^WLURHEJJIFL/J,-99VP58BQ\);" 7_OZ5GMI^@S(UB%2''8>K5
P&Q2+EO&-&EK$S>'>W@G&7#HXK:$PQ5R;)>(1KXQ97V@^['TYMFWGY"Y<PLI5U^PR
PFQ* 5@/?Y=]268:K$:(DD6&5H_%+\<<"-'/K".FQ&F#R[X*I*=&KL@L85FW'/B4=
P]<TX)%]/=;>]O!S[?<0YOE0\0@L25)I>KAG*G,X6/B1X@OUNKD7.^C?\N=MU!7D=
P-@MH4,^$ PPF(+)1(X1IDD?\A*S8J)32APWP)W<+:$G.4ZYE?VT+'P3[R7=1&T[V
P3%$ !N^O,5C<5%>PNQ3H]=*ZKJDR>K'AS'.TTVSHY-Z;_TB22^9,@$-&PR3FPJF9
PKO*\"":.=D:J@4S3$Y)U+MZ.4=AQJ8V*T)XUSGA8W&Z.:M]C="080Q>L>1F'[U<V
PKE0-^ZQ[]%&=O>/__H.1Y=SY8@W52GOT5FNTWKZ80,BHSK>F4W:U X"FG@?O?QP+
P/E_/D3=VM563<\'%2^B>P09 K=(+"PA.N5<32JAQV^<(/F(CN0I\OQ:Y'_&H%]4H
P;>TVE-0!!M>CF"SDO<X93V'5$AUOL K&(#B(;0!8%K&8(-UBHX1I4(X<^?8-.],0
P'=6F$!R<J%AK/_&+:V@!OI_J8CM*:C( P&'[5M*H0!CI;K?P=@LV\1- 4KW"J &+
P_XTA,/S^3G.X_$.T-D@W15!F70$$IH;/EO/>X\@YG-O5!U*G]-MR\'=34A%,KHCQ
P_0ERB\%X;^BJR J__J TMS'+Z17<R;Q]4QC99R4:/UO[E)+G]@2DGB.: I%8FT% 
PU+*DCNH!AM#%+G^;E"0UJT)F>-9DJ)</$>-A ^:&?H1]#:Y$1;UT#C-/288*Z_SN
P)XSA&['D?[+,Y'UV+V3O >6$[O&\R1M1([QNP;9?LC,9OHIC86AP^YJCS"P9FDCL
PT BUQO^L:.'S%3_O &J75.E)O?QU5+\ 9'I.3/5G-V&];!:CA)8$X-=+V.$0"38*
P81E3B4(#@^F8@O$-36+S/"+9W-&FNW4Y8E5B<P6_EQ^_E_ER*"OX<4.?EAC>991,
PR @%$W6(*05Y]:FH:5?*8(-.;*4 SP17X>V*P*:$<\\/Z QZ6HWF&TN(KK&L(.>;
PT<O,W$>N)\KL\*9%7)V6;Q"K:*/)D9+T8V3K3ILAL9=J13WG6":.U@/YN7928H((
PQC[7F_=$_OZKJ?#CZ,QER(O'1RXT^8OCPH&2"8H!__W_ *\F>FI5.>"BURB&,XA,
PX-IN=K^\ FCQGX0IWWXPYKA>I7K40:MIH@UVJ$6UE'Z*?\.$Z/PFF[P>)0 68Q'4
P  \R-/BT3^(SZ>DXK>!^:IG3;+)T_ZO#9"&D@ ?7[G\5::?Y1>J/-K[OWA1(E#/H
PZNX:9HNJ%6&Q?G@+T4[0XE,L)393URZHM3_!\& 9WMP_O#3PNZU[;CD'ZT),5$Y-
PX=%<ANR4>W.&O5RKT0#%\ZHVB'!_O963=6#KI.$@M3FW9[KX"4BT^8>G/B$>[8 3
PQ*,9N1>Z=XOJ32([O.;*%N'_,)]QWIIRW<HJM'N%L8+C=#'1K/KTT4TBS(H_67OV
P[3[6GUC:-N4;_4]B>F"8I)F$!%!\3PA.#MDV6&!N#I#&HO7?RU8+G"FZHFROQB$(
PC$'UE!*?PAV#M=T8VM@[8+O#*\(N1*0\L5RKB4!(RE-OXWC^DQ5@U!)A@T+X<6;4
P1+46ZT]3R'@K:':)U782_70DFX\H%H5-]](@B\W)9/;W>U;F;%\'W<RYG$8P!XQE
P1.$(S"..*Y@+4IK>SK-;9J7KO+6"SK2\,/3[O:_,+?O="U@8V"4GAEW)@UWMT0S>
PF6'1/8&LH#R;OTLD<AP:7;!H2U3?\$5160J57^:Q)*U .-5PR?3J%:D;?N$/6.SB
P(8J^',7[C,&Q1WE4E[?04$W.P[,@<\2ZL'I/F@0AA?=K;KFC BEW&XI?.WA_ZGP"
P$?$\GZ+]%0 0CF'%7?-T[6PKNZM'<QCM8G;3KN1Y:ULL@ Z*OD.#5>*!%Q0H&QS<
P;/WW-ESL31& 7>)1ZVCVK44RKALX"""T_;G5#7:>^RL7PNB[;OEASL&SK>%_ZDO;
P^G]R=G@W E0S#Z^7U-:%:ECZ6"#M&1?]//JW@XG&DU8#A!9M7[+0*/9<8:F>)31_
P_F3S,PB@Q&8RP<@#.YM?/@3A#NZ;>2*<Y)S1]G7OABQ&Q>R^P!"#'HK4Y'1/F/!#
P&OB,+1-V'W>):Q.AT0<UOURTQ/B\A(YL]Q:-<[I )+[;"6+^K='UTT+UH\QTI]CG
P8WO_4\9I==S(.H+8UH]MQJ+;G7]'D:J C^HI2-S><2N(L2/%1#(X1^J-O'SY]8Z+
PLEXV[;\(TZ,O[BML$U\GJ%@CC X7?5AO23\P/.DC2V:.$;HXHJJ414AN>!VV&:)S
PIA+8VJU""W:17M:4B[2GMEX5'XGE5GM^VCO>X+,XJ-0W5$N(TO40+F3I&I\.C%;H
P[XVX4'_H.4TR<HSQ_B-(V1Z%=@QO:Y?QT>RI+LGP6^9#F[9(.Y(+4@'HG%=7@8X@
P08G.4(A5YR5>_%/APPYX<IIP'PG=G=?-Q'=C5#'MP'GA3>0G<><>9 /\*_*^>19.
P(DJX1G<D1(LD1O&GS_*V'81$YP?M>.M#G]Q[=+1 M>+;#)?*%DZWXW,D>(8 /HH+
P"?.J993@55E#HRBTKB:44F?4+C6G6[=^QY]U<-Q AW8-B2^JD6YJE3V48YYI<X/P
PZ*VZ>2NZ.<L6$;:FN&J7QBSC2F)9LG,ET^^;F#I7 <1@?K=#QM\# V+N(UX?Y]02
PT()&#2W^*)+XCJ+:JE>;'@%HP9;B.Q2?I1G9'X%.YB3(;-$=^'RI-H_9H WVK-YZ
P1CG5T1=/I81YGQ<>'H0LF\LF,$Y5FPLL5!#?"0@:)L,XR SR^DM=8Z19LU&D$ZG*
P].#J:E\A)>:UBT1<7.>29-_Z$YEY!DEB4G4\>\E.?CE2A[TB<1YU20CD:H<?6,:[
P^WL/0SE#%_Q^=EP[7NM73B&/2*2QD$@ U+FX:Z3"#E;P.H-GEZ)+'&+ID1'F9D2-
P, $^!*.:"^K98:Z&]3+0$!L-0$8*Z?@9G0=@\_QCZBBI,HQBQ(GO<^1GX^G+*B&D
P#00]-&744('.5<GZ &.#XX@W/R^? @^THQU_TLF>C:C>5 49KZC$R?P#]6KL/8?7
PI!XYOCP=O0WBWJLI$+ZUH7-ER0E;+4?/UIHZ:U=1V6H[QAWX1:%='-=J6A:=A$9O
P(0+UF\7.BH;R+ 2\[1Q*XTCC9%):&%Z0+4\C@8Z3^6J?BJ*X:96GKBP%]Y)V^ R8
P%V[58K22>IP-=NLPA#:>!7G++M%I@BZ:%K"+H:D[E?U!M'(-?XY/_]M$;V3W<QX]
PB0\MR!FV)-J:$UWH-K4OT2WKZ-Y>4V5U)VX' )!^86]8<L8$W@R,#Z5F1 TRK2/W
PU-*KF2$[(,NN4*7;F7RE$L]A*[O#MH>:I'1H*DC%'-*OY%:UQP4((&/IUH8V6R;^
P3 *QAI"=]]__-(NA.+2)I_6.:,^U$';KI,"[%51($2\7.U)FBS=A2:&T+4!H'L3-
P;(OBQ66^P0NX(1N:&RCBH]Q)Z:A26EA(5ADV90Z 8[_ T#TSP5HV@-=S];;O)QGX
P*PE%2\LEN2A\(FS5O@B]]S[M-R^XKD'%V$<F04)"W!!R2DY[^!)KVZAMO%<J&0+9
P%)-UMUKB+M$3@/:2W*\U(L59:HDRS ^6$5;>U%1T]5; ='[T+B8''<F\);%N?$1(
P]Y2&;5MA)3O#5,^IG?JK&+ [67B5C]SZ1,TV?,0RX0:\8PKHE9392-+:S1""KI\S
PH:$9E)$(BA#JX-1X558KZ:5Z3[$]U%=7:T&8 1R!!>AEYI1<;\%;7[BEB3%&LT8'
P_J5%X*O_BDG2CUYA*B9-CG3U.G! ?7,. [(-?^IZP8Y+58<D.^J##'E]I(#IF1F0
P?:CT%)( ##M-?O[T&,&6%INK[2F@O.Y<;)R<V70>E:NRH\MUZYE%.T#)<)71B":N
PE(\NQ!AUA6E\_L_#-L?&FF!\[[3Y"X+HI1<6_*;:)F1OU<KE_!!@ U!=B+T;AQMF
PN/YQE. %&:7#J]CF"_%#/CBR0;>N7%#YGSRPK$K2/. $0@.V[HE8_0,?<?N@R:3?
PGL0&M^^!#8"Y,8<9*CHXCCR-YS HEUIR2E$D"M3GJL/;*OK0!/#G6J8 "L(5N*TD
P!;BN"-ZW6W-<H&ZG<('^&:A ( LKQU$O%*Z2J8,9-!_JB^BQA+&.<08706\2,8WE
PE6U1Q-6"<5A%/JIVV+W#X7/7)1(X2X\))SJO+\,!S;B8SVJAHY@J7TO%0'&1-Q%8
PC4<BYY@?'5;#T4_C1=*EVUT_5>KWWV:40&9[EP8TE!_%.P8/+[+E:S1:23A0#//I
P"(02N)>U::/ B[S>@<MM?<F&VBYADW)TXZT!/CP4#74?'*<\_CM/H>)13J+=@*%$
PBS;CT+;[T\K5/V2)&(X^4WTM!N7_82<()-V,C0$M@SBLY:/(;ZP9[['&D]4:>,Y!
PT?QLXQ7@@WY_,YU&>1:E.S$[SOE;=U[[LSUP;JS=<[IR6_U )AT2KZV[W-N5W8 L
P="'RC?7W+!PUI./P=3=X*WXB@OJP#]>QG3X$'\*A7#=XY:/:EM)G!=EVZIT^W*LN
P,*L,;)J6*OYLXY>X%<K](L%8PX\1I=HA8*?":/6C !3"YL1 "91UL\S\QC>2&1,Y
P:*J($S?':*:\FJ78NI+G\8"@QS+&@6.8B4/TT+':'%&9_T"&UIVG)&U4G/[XVSXP
PT(*,X!%@<@W,PBE)G'AI[]IW=WOF:<--,DY1M]"48,4LW0*J8)UIWR'C-O\5N*2@
P!$0QCKL4[,058&*BOW>\GG-*R",PYCR0&JWIQP7=Y'$]Y4X7PL>L!8\_?EMXK<!I
P78F:PD[_"3O8;_/51-@VQV7<.EH[&;LA.$0J!;V]G_;PV4_TW1S!:S"?_C%>G;]-
P%'.IZ$IFQW I=%*IL(=2]7K=4<7$WCSI-,]( H+T/9!D.E'__@2@HG!!D:R$B5M1
P1<5<7V&4?<8_D_(@J8-(ZIT#)R*^$F#VAO*H>)&?!6\;G>@4R94( CR45K2_H1_Y
PGX\7*GSF0_]V$4F\B7C*'F'2)Z  ;%L2UHC:V@SF<O5RH5T@>^)R+6ZLF!E_>9G2
PYUH:)B"W((URH]8YA^ ATBMY_Z&.?&_\^G-'$,#/-T=1HNK"@#C3(&,%K[!,1$?U
P-JK@=:$RW4Y;+\-!8$\!Q,!338/_?!4Z7*S#75&LWW]'@9Q'P[GQR1F]Y7;Q+7_@
PK1R@3VZ-A2SFEH+>#3!.U$;VD<]V8%,9OB+O@="H:3ZM%^7/QY;HZ .=UFCA8.VP
PDT+5:S1/,)B>:\.1#S_GH8'J-]TLL> A/]IAA-#*J'XCO?/Q8W6_)\T(@2]:Z<X!
P+;02L\V68@QN[!CR1N"&SCMS!(GRD.E#I=O>3A*&10 KQ#6IJX?EE+.S2 QE>/EQ
PJ>U+(BEVL!HBM]@%Z#@^ 1E>HW:=!VR!=)DWIT!L/)]SMWX<.?8'+O;FG_*T<30<
P@H$W8I>0DQ@8GJDM+<DET2/0C38MM^4P-]@*DAJ]/$W;S7[G7\#S#<VHCCB,C5Q*
P*2(VAUU6<'L2Q4*O?G!HZ@0Z4,'#BIK<M,7&8-. KUQD'3LQOEU[5![EA^E>*^F=
PXDD,IWQHS[;]6,D+L==X!$17GO>*T X/3 DFN?2WRC^N2@&ZOOL1\JHJ(<8B&R[%
PP..!? O'>:7;WMO>R>I-T-MT5U2Y.,W&H<LFK5E?BF>+LM3#EH$W<T*842':;)T,
P/1:JY8],^KG;D9@PEC77P;>:I8,U4NZ>$'? ^Z&:<;M:JH,+#X4&=/^,(>H1G95X
PJ/WXS(2':>K\MP@PI\>T@\4/RXQ2A/E*;<PYN"1&@,&Q[L[WUPC&R8F&&KH$(1O+
P'CLQK;;Z/=M81"//W2IOIHE3!WSLH((C69%0N@2 ,PJPXDOTZDOV7K2+UW^M&%Z2
P-B^*=.9#JY0Q?+*TA:Q2,_->A875!*6UZW (U4\O3%J]>NG7C7IZR.='1A]+GF!F
P/$T"HAE]M<B.[TX:C#/IWHC#U/\=^/+Z$DQ*Y4>W9X^4GS'8>/9M-?X57-O-0>@-
P_\Y-"B3^BD$A4)*)^OPSYB+8X(3 [0H&N8$-7*941)\U"%EI'8*/F:"A15)WW"J@
P(-D(-&)+3$S<K1#B1<JD^SUX:=3N9QSX_QLJM5"!O[S<'N(ZD9$"H,G9_FDD)NIV
P>M5#'P<4G,O3ND;*C2L[DQUV("#N!V \P9EDH5+@TZBR*56LX:S@YCI%=8_G',^K
P(NNQ/52">S^O%K/05.N?5\S@#-#5(;"G?3B'7[\ VW,9B3#TT=]"6'X<H25JM,ZS
P,BFN;[Q$2?X$01,##7"[ S(VG/2TRUN+\7R\50YZZP)B+D! FAWZ*-;8%"=7HTBJ
P=\U$Q L!F031%L<,L:A$!I9FIDD*T?FE'4BI?[VLE+^:\@Q8<"=W:.5=#1>MK&HW
PCVS&^9&F1@A#!3(29NWT_F(3O+M"C:V=?#%-)<R>BSTU7&*BZ:H< /@$8?2)3B&C
PY2UV4^2?X@0LS'!Z<AB[C =^]LN>,/=G:]B'[!P5855I_*%41/+WG=/AJ#-G\7O5
P,CNTR1:3*O-VB6U"$3GM.X&O2)O1EU_<X16''OWU.?"07ES7\WZ7WK5P28@XA/L,
PK&:XK3EGD*6,+!K\%%+WJ-7ZVFJ7-+<"H'$0)D. !(J2Y[EE/ !X>C%)W3 _G%W*
PPD30&F'>9N274>R_.<]O$!U<F@#*]^I57(G,@*%%0#&X_)Z17HKYAC<0\QPV1/WT
P$CLA<7R1J6T['] )62"R@:641'-4$%,.%S0Z(!9KL9T;SH7NMRVS.5$8Y/I T8.F
PM/.P4T<.:H*K:8+)0Q2I?LJ6CFK.CCRM^+5B_G/M.&I"HV"4>Y8*/CNF1M4V]1/]
P7!AM=V#P!1/T$V#GH(Y8DFL=2 < 14S8(.^8U:%'UWFL4;K]>9E3\QL7_/+NJ4Q#
PDYV97G"@ISE-/)!_$. _79]GAM:PQS6XG'4&3"X*@D!,7!ZUKB2WHQ\=J)*#.;!U
P@/22X#:#L=,PQWO/V26HTJK_C2FM@G]B">A$J 6_HU]()5L0^+_\16+>-_O_$0VY
P&<G^V1M=DMN7YX8N4BP)\-]D1<WUD+U_AB"0VM)MOAHS]%Q,]%;H0!V!564!*-G=
P(U]V@2158U5#N<$)% E70PXGS>*TN\??9U1!/&5E82&AYK92J.#>J'[S#MPBKM,-
P9<YBWOU0MPI<?F^0H-7ON0'(L0_D7,ORL"6>GDD.=F67E)3VG[=WBENR\U3:#'+R
PKW,*MF!/9[$UF&Y$12C:RMC <,\;BSL&"<K8%='T7 LJ 4;P[!0J)S\I#_/.S,\7
P*$H+[:\[20J]<I!K/&MRG1"O>Q%)??$$TB#AA@OWZDE[C9F#BW? !$YGV!8*8PP,
P@D FG#1Q?VCW!ZE9V<N\ F_0*L'Q2:R>%]$K2MF[2$QJ=</V%NQ"R@*OD4OW+/7M
PB0'CRAJ2WI'X><1QH2@Y3&EI';Z>82!W,R64-F^@GWUS:/)!R^T9H-Q Q+34V3ED
PGX]<1_:[!JIMR[K23#V9\VML-@*=_1-90;ACH 9ISW0HQ.N$&"BSGG#-3@"(+W,B
P'/Q1R<+8*$+:V.V./%__;F:]+%R^9P>LJ7WRDX7K4Q13M).&TM/95TW>@ >7^SSG
P%5CM:$=-X )!S]C/!K> 4=*QCQ>RN4FQ4W']$;/VIW6<[FXGKB9K.=';6;SD3X@&
P5G^D#6.:@I&? ^ 9>K?2R0M<AW3+==T,O/]9*D.2YV[@<''*J/N-Q"2X,K682I43
P;-[BG9F2ZVU_3)9B6.Q=*L>)G1/=C]"SG8NE66J6MU,P:,FXFH.(&?>H=R>JF25^
PZ'WLS'^Z:B=U"2J5FJD%2H@=4[_,LB[N<]4XRZ<*QOM'66@7)+C;JEEZQX,^> 5 
PK/)W+?@U\5D]33&0L'D=W321Y;VSR]/<<4I)O0"/6 A;<>J$RTZ\#M_>$TFK_:56
PTB3I; C.\>?B!XV2.>/'Y:F!V%!2*TM_#YGB1]JR>+QW?@L?NJ,( %^T4&?P@AX)
P0X=;><[GDO9NP+Z(X$F"9*1<IB*S@:YUI-:C:9P5"^@.\CXL-;S0FD(/^64)$LYG
P7NB;^#MD":.N</04Q<MBOX_"?TB8< 0[%F;KZP"BW^J ,8-I<<Q^6&7:=$0)0!=H
PG2P;Z0?8+]O+1JVE.U&BY#U;292, D?BAQLBF-\L"$BPP?\H2MH?N,)3_HE>"1 3
P09W= )/ZA'H=#],[N*8JRF/BH)?:7H[:\[%A5 .N1A3-AK_X<4NE0L!A+]%HV@0\
P$7/N/,_B%0$9 3S]*:Z.'4RF83>>NCO;)I&+>F<181L<T:52UA")!-7C/#L:2-\.
P-@X5MQ!X!P!#YFNS%*;A!5'ICR0?W15=LAKU+G.XTHX>9F"-(V'NM_7C%"(;_P">
P5EP+S!\B+MUPJBYR&("E[NP=\(E;H@(Q"%( F./!@B';J@-$%G: KX[L%.3UW[G_
PW>G0!/QO& :HQ>P6#0<JYO5^7M9'>&1SL]D-H-8D4!8CW"==H"=GOK>L:\+&7$N?
P.+B<UG@S+%>#]>>$L&1^+TNA<BDM>I^I;E9P]E>QQ) E$"1$6'3Q/*HYX;8.KY2T
P$BI$4E)9M7_(-J =+C/;G&?4\ZSJ/B$"!:"AFF;-JELJ!D-!;A1X)%,: :I.YQ 7
P T,J-)H2AYN@2'(_D3=#84,+*%(?XYA]0*ZAK-N9J:Y"\.=?&:*T0"]9J" ZV*V[
P<VBV&A:9838_< Y:^&%*=_!FF9NPP/GN6L0HSZG2=R6!!G#4K7$&)PA/>4I__KE.
P@@67EK2QC3XT5,6/;1$0@Q&R$@S!XG[EF(^0"TBG [(0>$=3M@'1D>9-<C81:]8K
P=?T>CJ33?4[B,8FQZDA_,BWV[-\_Q1G;5\3 <(=)'C,X.WLJ.N]1OU9:RID!BC T
PVURP;/A$HQJD;G BRIJMI&V7]U(- )W9.X6&<-W&N12=]L+S]FN^+JR&:*9[ZF&D
PT<$2[-@AG@<B4OVJ/;<,J(NB^SY39!Y3:FX[#)!@\P3=;.I2_J$?VEFD&9ENE[!P
P4O?$']$+6:*#4^G'UD)\)]AY!"-"PC:Z;K/5+>J>E0,VO4]^*8DR/3=*'.,>AT$S
P2V"IQB<(/*9JS2?@J O 1%(4] L>7-RR%)<QQ'G P#I^$(^6[)[43V#!Y3:R/K6'
P]6$;HP:%2A%$:$*( \0D(905LT[]XQY?]"HS)S0=27S6QJ2ID8$)HQ[79C1F GNJ
PDB[ZXFPEG:?^.S,SM&86, Y[U;B(KBH1MPML(U],(_&6,2Z?].F]_%@(>HB"%IS=
PP<-\,__&QJ#HM:D5U);-#(MBQOG?T\J_U ;A7ZT*3CM\ZPW#C!=YB35MPP@QNMI_
P<B"EB8X,21$4GKMICZ-'[L5^)6 S<1F, *XOD'_/(9BX=245S"BGRZ0+CT%<;UH.
P1>LYX(&(8$CX7'=ICQ?B862",F@8]P?[A2H'5#"]*_(D#-2'.& T\U.[4(OK$8@U
P"AXS6&G L7LA*X7%WKL/;.$\;0%S'_$-:H%U$ ?G%"I:JO_+5 2YC'!(BKIIG]&N
PRMBB3B*H*D(7<Y_:WX_>8_ZD=@$2)UZP6];!ZIDG/!V*)_]^AY0(-D3,D; . VYG
P([UQH*8G)+<RR=9LAVEY<&S0U/&&YVX%MM0Z!YXP9-<LQ79=\O>70T,P3,4M8; Z
P<<:8R(A' :%;@A0"/RC)4:$I*($)ZH,*P[N^/1O:\Q6?) 9LH\=%@F/Y9LI5+=L%
PJJQT@=CQ!1UFS%[MZE_/#2P3N. ?R1%T"2D>I<O=U?,LKU[H$;,?RU\V9H"T)Y,)
P4^0Q7]4M//3[1P8 SF^E#-&2-BH;_\$O*6!:\@V!D\ 3FNM\D* *[17@YB'[_9',
P'NVSYLZX7QO:'POA&$/:E$DX$I3>G%YNXGH1I?;ZR;&SLD57BM/Q87.2B[#YD:E.
PK8^E4%<#(2*&6\_[EU>F'[]8UG%J])>FI[_ /U!L@!56/N,YSN1T8,OQ7FS _ADK
P(UL>LB@D64.[Q:&_6#-5341K:.+81)IR3..>1+^^C?VU^, XS8#TLB(3@</JP.-^
PGB&?:]UAV"M]O7.N^(4?2X"M4IT]]0C9&>_!O,QIF_0*)2/&#W_?7 4^+@(!)@9P
P3)Q9M\E#=4;[C?]B]NN]XYAIU#9[Z'@DI_>27=HTFUZ_/2AV1QA;, "=SL0P.[;D
P/TS48^8.=BR;/\".^Y:T#4)D17#)(,BW=1V,$470(%_;L<@/XX7[L%$@N>!BWQ71
P&PL_;P/TOK3]/*N2P/B2??U<&OY6'02"DJ'F+U,B,JZ/LUQDV$+77E/NX5E)&!O[
PY5O7N$1V4TL*X*Z0OVS42!2%U?$H-(4'^>/X31UI.$;K^OD\V3#!L\P95VS8&,[:
P.(\N.TT%!\1V>N)=28J"<=2&$;CSLY0NURS&2U=RUG+N6LU0\I8!(9:H]%QTVH.J
P@'4]SO?*B0MIFTV$,V#AGS2+7E@?&T]21(OH(0D),XI[2HD 3U0HYVNT9M)$@5#,
PKJ'/]3:W]O67R?,Z!RNSYM=]0WC"9*535B(VJ/W'9IZMG U/%(O[K_#BN&AE7@?Q
P(<XZ5T!(%I6"$*OBW)6W"$X2@)/0YK;GU^I], AZ7RS3IWVOD@BA<M"=;IE^E/H<
PJ;HP4$_'0E0VMTT?%=I^Y^,,KT;9FNUU7VB:_2!?^,IE)EG'&>/$$.5.RJ4\@353
P8+(ZQ3,[D$+LCDGBB?(3"VZYN)#)D:L0D(P.FVF3YC04LI])/28^5*HMG$9:\UCE
PPJPXO.4['>MD.9(6[IJ4GETOO'4ZJ"+>Q$2M?04LU)ZSXO%.A!83E)1P^%Z_'D"=
PN&NK\FND1R7/\0V.\S>@K^LN#<=WQ"<D@.Q7<)KHZ7F_6P4H=S\,II5ML4]:DL04
P"LXK(43P! \'MA&K[;0+5![:*S;2U,3B_C:5E-7:Y#4>[Y%Q;C)2KNRM50;=LA"0
PSH5.$2_3OERM%N6\CLU9[G9J+SX\YJI/) U(@EQ4S:W5'X_38FS>-9FA&]BCDWV;
P"_6Q+/5770_<7G:>D"_K?) *3]R\;7BQ=@:H1F"-<JI0]K01U'VE]J_3MO@T4.-5
P::^FK&A:F SK)DRH@"W7$&NMK6@*:IECWG_7Q_:+NMF.-^8]_@AY!'GQM@M0V4?+
PI3FC-3@0?',T3*!3HPY5F[;\?)1QUG6'@38#8,T68VR\XCN(&YR X>Q&I^5#KPVD
P1&CK+043IL$: *"BG+'^S6&-*;K9_RW08\JCL\S)H,4_M-E?4RYRHPDJ GV]"*Z3
P:\TQG1>8L:M*;^)]VS.=0 <_.@P^,_&1FJV9T'@+5->JEJ;U'T_0*P2>N8GMX 4&
P'U_;V$*/U435$S!-3]N?J@.%TB-,#"7M__FD[EC>129U(GPE*$*T!S101$AH_RV=
PQ&I%]YAW\!2P N$L'1WM?2ZMV:WIUP58#4*3=D9494GI"^-S>J%!KX=>6Y>OG+8L
P3?U1N@[=3'*D/HT4$^KZ3F8TT5QL0P")Y^&':MJ+0EPBD";95K!&^R!G@>S/R-H#
P^6TYZC1G'BP8\)GRD*U/Y] :[?ZP>\V:4#K9U0/76A86URBIYONDAD+T;<6.8 (0
PWC*;!W4S:3,MR*-J\*QB\:E/C$1U9<_A_!SFAHM#HS$.20H9 "D@WCE3F9ST$8,M
P8RH0^4XX1^/XI2^O$&7QD^+&YO&E'E])EF0I]3."1E,)6/[[+THZ$,4T\"FIFSF>
PP!**1OHSTT\&KJ5TY^;4&+P?!W]Q[7TL#H.K(=@I@\#B(Y.7_$')-H&-WG;TD3)^
P6@!+UWN^\XW/<W=HMND=(#\0D5R_CZ>O7@ %C"*);+;HAXM:+*"6#>@K3 V=U 1U
P1Q^'54\M2Q#J=3:>)SL?W(_PHF/OJ)3$S98,^V%RVT8$??11=:.UOS$JHGZHKVZ2
P"@^'O<\//1.\]L]C&*'+I%1A])M'I9$G!"FU9M;5?K!DO,,[=&T(4+YSSP7H9KTH
P2474D.$/F&D2KB75VT-RJ;5'C^D_WVB5SV;3WEA72CU<>)#'MA22LZD[L4#;E'$3
P40^.!+T\VFS*GU]\BNR1O[0 4W*W'1P!*]+HML'F0[+^5:.UZ4K?I?:%CZVJRCX_
P,9]Z7-_9>#/[5(9B1(/D1'(W@U;4R(*7,H=A5I-[++62VIIC6%W7!H,ZW]YVBC42
P;=AWLM@3TCU$>':L9]J29BJ 28>[(YGO'ZEN'N!6A_,?YPF3\&'D%BBZI+^JR*3Y
P^B(<313A#!+4Q7Z]UE T6A=1Q[(VE[,.Z@CJ15&Q:?7!:-T":)/"A-.?*?<Z<1CC
P^3;BJY]8FS5D)0X,>\7F;;(+E6X@2&IS_!VE1#O4XD0:D% 86C[**]K3C6F0]0(7
P(A# M[&])FY1_"Y2;UTQ\"DB22EKON3VF0D3)JUCVU9)!!UU,$L*&#NZO"RPKG-Z
PTUW<=$[ 3QBZQ?N08%O,BC>:M&_&,Q^X/ O\<(].M$5&K)?&^P?F3Z7SDPDATUC4
P+["\#L2_\!OSB3N8D%:'\ S4*#-GW%LL;DY3^B<=K_L7VRNN$H'&E2-RP]F9XF)4
PP>_@**9[X9:A \8U@7JPET ((FH\-=AZ*8NVKS8_?U\%]#&%#M85$:6'4Q;TK<:A
P@E-Y'QY[DYH;*?*$ <:H9&V%M'",)O'(XO.R-V4$ET4VBFF8/<F-@GQ(DF&UQK.^
P.^Z*,,P,:LG^12A61,^R#FF[BJJ-_?<$&O^O*/6>DU**"2=XIC3#E40RV6Z?#-;!
PPXA$:B(E[+-_8C=I;Y>F-&TJM.2U^=-!PUEN QA(H7P*O>Q>PXW!=\<LG7\_.'.W
PR# @B#]KG9]<TK9:MGBB%W*9_[>_'[6RFETAP*0$#Q$=6K1:^4='^BWDL/P?W%#>
P<%+GE5/]64W=T+WTY?=YH$4;K1STZESHC:@+QS_T=:\A*V&*T?,Z?._U85*-E;<'
P1-8IR)[*$X54!N0Z"E'WP=IL-BR[-,&3'S/]\H##61Q7NF&KU(()O  9-R6 !K#$
PO6Q%URBXXU20Q"OR0,5=F]M.$=@*VO"@TW1^:]%EO^PTQ11Y'[1DU(_&CX;LBK [
PP<T#0UCD^Q<$MZ&W#C>Q/%@8?%]WAC@:B%X>CH9+&'A@..M@NQ87ABZ^1N6WL;G7
PL&/2;=((7\@*>@#EZOL7Y?4Y&!$^'DN7$P:+WB40WN_KVCMIM^<!6"56&W.S8_UL
PJ?0']/\5.Z<5*LVR^#N$\Q I$D_<VH:DM[<1GJ]-O+3'P&;]#*/2'O:\ 6,X(7MV
P.3J9!E&SA749# J+?5[F(=F;-[_JN]*Z8U&1ZABNU8L1YIF%6>W1X0"X!YBW_*"K
PWDSSNS1O',_%L,KL"KU2G11]@&K)HU+ Z[1A<-;:081N)K)E90:X& RXS9,AM$ I
PIU\VK_A7<I+97R>"CYW_T4V$)4]]W=K3*I08!/E"3[SXK\-AMVQ-Y[,(G?W%39XO
POC@[K$7B>W'8%,1%H0]JWVJ-N$^A3M%J[D#L;"J=D<LUHTIPVWWE4$[JQ&R7?WIF
P3RWVS_WT\1*;=3I>S=0]X^5UJ_=M/$P90=N88:]$H;HR3+_7[;QLW#!2<_YK!?8#
P.FT5/J_[@E,/O\F<DKM5N%[KL?,LRJ:AS<5O;2"H>_W97_,>LJ)H^JQORK9]JNY,
P!+-+5,@[Z*QB)*?,K&,!H=\DUKQAI"H]"K_2B.I_=R1"PVU-8 4 _%=N<8F4KUX>
P5;UQ>XPQ4VQ'F"<F\U>0*20;/;47_B)&=1$J#^]I0>] <MOOXT^[0IMQ1+FGPGH[
P*Z1'J V&!))HM4M:#D)8($RX0PO(A?*]CEYHJ#HR,3.[YMZA!&N\H@_FH]@NP_(I
P)>VL"=A#_FUDATV8E8B1890HFC?7M[!<)&).)B5HD9:21MO5UXW9=P6P%,W8DM7]
PM=?/M?K'PL&H]^ =^QYYK"SM*4=M(--#IV+/57%Z^>2+'@3T6EA7"J.6<._CKZZ^
PYM/A"79_,M"6! ;NJ\Z)\'ES\_.X\,K<?U^I+)]XLVNA$2!8T/KBMF@TL62ZVFGB
P]4;Z24HS38;;I)%"/-#,;Y2$S5C)C2,H[8..OC_I50A_I <U"'IV(EJUO 1?:Q3*
PC%V&X+LG(CG3QH]X 0KY7SP.[!:V);7Y*!E^XSG>5_'_&(N]^;A47![,;X:8L^O0
P]?4#K!D:-\7C$70"-KPA="C#ZR1CD<%O<>J2&??/#%V++8Z\ 9,O&%;@VR>[X!Z1
PI]6#&M?,2G'DAE5QUYAAFU@V<L5YV3-9RH]TVP_LQ:RG/;1>JN-)-_XE;)@/(R0>
P6H//7U'.1"Y7S D=U?#>O/&ZI/GC>.4B%E8][4#E:FZ&ZEK>BF2QT K<'NU;;1AB
PNIE,DLTN7@XA\%96QO/XL]/6/H1R6"+04B&BA[6JPC5$6B&P+%X#KB)B/6CS$(Q#
PSW4WW5 I/E9%:(T_B("#/S:0/=3(HQN)0+IW]*7_9(=%W+^J517C$8^V)),5MN)3
P]((!A=^2-+!+(C+#R/[.RI1;2.3W!:IQQJ'^(P>Y3H:.%4/V=-.!ZS& H-1,HA5H
PEHZ;; &+FZ=X!\0GPCK='5-%4=PF*I'?0%IN8E"Y0_<+Y[\3Z\N\=.!8<2+#D_I(
P8=>D2@48CLTCPUDK((XJC8^,>B2O?](J)L6FN_;<]V)W7.*67YKNI_LQ$]&)^; M
PWPO,=WO:I<;43?_/4%UV<$@/'-F-\(-N#PS^'D]#IL[=HG7O&0=L[#)6?0IV-9D&
P:2I[/TF$!L4,IMT?B8HR0<!<TQEQ0$GSVK[#KX^H_Q(P('G@B4!FSBR?.2;7HDGY
PMLM#]C&E<5CDLP!W]A'?5<C)-P@,Q68AGD/<*0!:GS @444;8EC>N>P/9[YAQBR=
P_TIJ171O@I=9H2O%_WK,!$?%LD1VE!IL:'+MA/81!G5PWHNEH:;[HJ* S\'R-H-Z
P\4LI> _^.2 BEJ*;7UBS+1X?#C&:]@)E"S&)F_$E2B1KT?CT7K&)T(&E&\0V#KXF
PZ&E#=)Q8KT'BV]7&?<457J2[FOV(Q !"#\ZM,8$?LNA2XH9Z!F.>^G]B[8\,Z9#[
PP3X&?2"O8A!AD+!.#/\J"ABR4U@R"[V)0"S[>!1WX-N#B1%L+1-^OCD_H9N%).;_
PQ)E-_^E;6+Z\T,BB/%_]IJ+ON]X# 0U\%-,.@90XK@6C)SE6P?<A!F&51F^:12\!
PV;P(JN?8B+NF'EC-H7=9< @((%R;_*6.12((9!$0>?@W+HP%X1S]6'NO#:#B4S--
P;3VKAJ)5/;W0&\5MB1-[V13\9N2V%8_FM0\FL?28K@X%E<=BO>,!W^KRGWLNA'PX
PW3BX&FBQ521ZPQ#/^3<)2(S.!D#2LW@?7QW=BH5+=)"HB-D6CM&OO)/(:O=Z>DKD
PD:&^$7)Q552BT]ACN1 AM];$KSLZ U@6)C#7M#YC93=.6:&PW27SK6HR!,?,[[(%
P.I86;ETTSE)IT-WFUE$*I+0,03BMK.WVT9SV@N(3G;Y%.J96W#"!))4;/!>N9NOB
P+Q."3R,3=N)GUA/XJMR)F943<1L[P,BN"1X>S>);B<F-\BQWD^!>SU\! F;.U9B6
P,BVQI,H(J&2_KF\LMX_X,QUN?!OOY4#)7C 79":YKFOMLIVS 4=X!E4RW5QT2(*"
P_<]9K#YAZZZWI'E7/+NDII_1MV2G885C!Z_,B^K\XU6;YR.90E$?&0^UZ_^X&0CF
P0]8%#VQZ[Z.PHY.@^D5$W2+C4KH^FT.%<@U>MC\M$:5RI/.J\&R0]_L[LUOA/LM*
P2*,CQ]NA?!<["+N-,P*FFSU?Y&-91">78_HN$2GRWVIDJ5%<BNBV@Z5GM]'G>]6W
P/K;@B8CB*F_$C*NBS7S!Z8AMR!$=.[5)WI-XM//[&%MYY?Z!BH_+1UC8#@9K/T8+
P@6YX6:J__X9%65V<!(7UJL^?8NWPY-.',T15SP@(>?(#BV;GZ$?S"PCH9X6>/:RK
P6@'7I*=27M'W$_W_QV,82Q'B&9.W5IOJ*(]!D*P- HUSQGO%=8I7)2.S"0TO\RL[
P)P\/Z[>DV59QY#'DKZD##4MQTKNQL*QJ'U!5E<K4T"7KR38:[-)8KU9=.#ZRI]4K
P)#3LS]/>G 41HC:3$=#'A^=LKK;U4,OIUC-CC5>!_Q];.A8H -M^A$O\58SQP%8%
P@R*H->;N[1ZFR.8*(*/P./QNDC2?^6/WGQYBFRGM7=RW["17XE6C@4[P'$)V)RC1
P(5-'.QB??KA9DP#$8>XN5"%XI?1#K5JM#8W_OYAF,[4ZN=#)I181[1LKW-9BF:HI
P/D0MD3IRJ%;;FB;@7+(,;!W56:_U7T>[3]Z-52#]7O$0[LK-(9J8\\M\3,/NLAB\
P8Y@!UR<37%!SJW5N"Q_'!IH\N^JMP?/ 0%6.7S;*D:XMD9)ZPGL9P8$C/C !@'K 
P(".47_1KU"T4$UL'_LN?M!7I& G&0-]-P?> ,#?=P:AR[(8T<-0<A-!A*?NG5-JK
P;V\!7M9.[OX%S@=<J4C7G,.:]U+$RPQ..4>KR,I)2N&58T J10407P;^7%6TD';(
P4F_OT.PK;FQYY5I%E).=, 94!CWVP9;2Y&/?7WD$E.Y]G:O#<?06JU*$<G[_>/(S
PAAJ(;[\ 284]#2%#7UX.,Q\B'5=])$]W[YM+).!CI=KU8GY=$ H 4+H,6R](]S5N
P-K(K^P)=IC1N3-*"])>G190UY/XY;C.HWN.%I[@-NB#M3$ )\-'"D@OH7J :@RG4
P9N=6;EAD[CQE?A\8Z(/]N"D=;T9'H\-(N >%87C3QAA:;:/Q]!"#IXU.])+>=7X]
P"ESWK*U ^H-AEFNTJTF%2G4OMA6+#J.A["#ZT(P9)'5OC)\4M#$B@VGW$8UW;<-\
P(VH+4SY=PQZ0>LU51L7B39&QX_1;P=2LC:WPKN-<"AH5HA]S\QP96$7]RUAGFLZE
P4[!GX&A PWP9O><0\_1)"\-3@6,<Q?A(RT;KZ8_/33(U%)70=\SBEZS!NPU\^QO@
P<E (X[M^6K!%1E&\5P8!"[6=0]E!WJ@0I5%O2&2&?&GMXD.XCQM1_U2\,(Z+/'E;
P<Y$_[PA;$F</+GT$NL"7S5*#BUS%#2U2MR)@G2+TE_C4_<)DDA__$2;WE39:8!I8
P-J- 0FIZ$T1F72.X3TL/9A_6T$E&CH5S6RC&&Z/H*2R_V22/'AGRXJCAGJ+ G M[
P[UW$#XPVD[R,E1+WTDSR'3E!#RJH'O6&EW=CU-![DEZ9=A[:&\4]2-T7O==V,HF&
PYKMC%!MT&S7+,W,U3RQIU_B,V='F5>?PDBP9M&+>624W2UL@/Q2[Z ?:.7MM7NES
P-0=99R/KY2*+).;V36!N"5;"Q:;U3''\S7+.(1WZ#F2&4A=+ A:XV]JP8B9OWP3#
PI9C4U[=S W#YE<K\)0AKW.HF&BWTTA7EYLU;"/#S.'+UH;=@X_@$^E8JEOELH7B1
P-\ET#$27R7'',[D&>N5JR)6SAAI#6(1U2JDJ\F*=A.R'26@>B  $@"EY1JH- ??<
PW@=)CIR4<?0>D>DMB6:PM: $>0+(D]F ZQ1$.OWOTSA@6LSY'\L5[E?#;>*+U#EK
P<<*@-6M,S];3($SO=/2Q%B5RKT=%_7R- &8*HZ_IN'JG<.S1M0!CBMVRFZ&Q :\H
P[Y-=X#-3PHT<7@C3N1YZ-P+ *"=A476SO9=6^VN3,%$B(4FFL+,0/0<C89_LZ5)O
PMS!/]X7'RED$9E,%-NUFDXX\]'P^B!]T0;PAQCJ9"Q%55TF@CV\>TTOL?SW0%DL?
P3-14M&P,]))SDG*#^<%;P)M64/GU9;'VR2,9/S2PBUP=[P/P6RMI@<@H(Z&Q[PXL
P((8YFJ+B#/R:H"K4*)^L,1^R5U93D\!GK%$UDXK^W#F@<)OQ7*%D">';R +R+ 13
PDD+B\AJXC:9.'3_N[V?Z-,X#@">1QIAH\3P+E;9 &L>V&P8="VJI$JD9-4$ZMRR<
P*4T2?6%5-A"HS#NVR5"G;.]='0AHI2<+210_N!LI0+OZLB^2^N3ILPJ]TGB!1%8C
P,DDJ2 \;!^^G=JR B%;;K633=.7W6(,X\<,.=@B)MV;RSZPY;A5CEA+,%MNR!PQO
P \UV,0$,UA%1FX3"SB^S)'JL@A/AY>Z?+]D0AJ%2A X. S-\O&)1>IH:J!Y.HA0O
P_U;\DM0&"I9HP:J0@<'DN= 9NSIT.$&8_I,O89">+^#0W@J^7JJB)8<I=NP5KR*-
P.HNUM8^=:,>5ZAX"]?CB0DAYBZ?5D4-HX $;5TWE9Y@HM]&HB04G1ML/S9V"(,3:
PBY4*V;4A,_#M'"@'*S!-)>](_(/.\#T;,YDN-K^5M^5^^SYRW6G*CA$?31?Q)5I6
P6?>B1$^IO"A7P4"N+BC@&VD<#<1PQ0^ N;"(-*:4#=(-\@.)3?$5B"I.M(:6[P4,
P_3W$;9F8B=L1\_OTHJ30BAQ6,["9N.P0NHVDMX;VS#<4#,=2 =F0'5W@)8E#Q^;/
P,(6&JE"!ZZ%3KKSYFX%C:L<[U1X5R/-1-JRD!BW+PUM!HU%^S](Q_*%!=Q3MVIA*
P9B0$KXU%,66#W@R".V)W^&XC_ POP%JIH!=%O7:J3%HG@J+:CWL>._XL,R013F?O
PEQDW6G83DGBN=$2EG6Q'O9%'(">-?^]H^M;>EG YZF9C=4R,5=YG=<^6&VD\$70)
P39;M[3 H-9#_(OLN-2SSP+)QZ# $FV!EB>X".'KQ(<%VC6)NP]C6UN\E3W=PW^7\
P0E>LHLSZ'-'\FBIFE/YQQIT<-&5@+4@P"]13NO+2&>\D658N:"X2Z'[(VO6EFIWD
P,W';]Z\J5)L&_NE4UAN*TLNG@V7AP[#FW)W^)MAN#:^Q?0.5V\Z=\+9WOSF@-52Z
P2O#['K86Z"038STNJ"-=M3HW5$,"LIOUA\0"EM%<(HN[W7$E6%GH9N$TW#2L?N)0
P2=KGK!E+LF#%LY7-R!5<4S2$U+#'2U6%IJK])'4OQPYIC*=S@7J.J0T"L'=))946
P%79A^>^?<+()=-S)^=C25N)R&?T=N;Y.:^M_1\%GT4W@-*6[UVF=I522I/&T#O/I
PZI!_0CP#GLM+,0B%D7KN-<Z3@ZL(,*7@2A,Z4=%$DIVWGSL.KOR*(&AV]GKQOOD$
P/:[Y[[<'\)N' 5FVJ-"$(HVPI+_1R-PP9+_PG7M,_XU^-X@HV3!=MCX4*D6X.OB!
P3<Q[U0@O'-X*9:+T$"N!9 HC;)\4%MZ#U\$E8<K@2C;01&7W-U$7;8*')BTCE<%\
PY^L3(E7\KUG/DK!M..ZK!F_YM^'VF%Z\!&X.6"!:*TAAV 4]8*3=MPJ@]$PM[6EK
P=6N9;)P<^:2^4J@OG/Y>%Z,&\W6O6>[8R(>/W&_R&3^,H*& 4>4@R0<S6CG%!$#S
PUV#A"4^_D87'PTLP.-/*>DN"')3+DF"$)\9ZTDB3>Z)V8R_*3A8*VD .+L+? K5P
PL$/*I:6F7!<:5UOL#S3;T M/:-NFOF4*'$9E =*7!'9PB]70U A.IW1LA3->_<0R
P; )I6/P"U9QP.^GTNR>B3I#ML?Q61MQ>)9CC\_L2G9>>3$#7^]@42RO1GL>W-;LU
PL0/ZZ&/!\"IU@2G:_T.^ZB1*P.+9HDB 01N8_+DZ /^%P3,J2S!T);-'5 H>4U]E
PFK#\AK?YX]=AZ^4D$MWJBQU_(?U_<4<UF=4X/DV0QUQB_!H&=\PX+)S,R$Z@XI:'
P[/P&91Y"7B44+3\J;=8[,$V41U"J ,GUK!+SM:L(M7V8IMNADOM:W8SWQ_"52P,%
P[1_H:;RW9R\OM9>X\LG4:6(85G"^F#>!<@*6E-%6>A DT[P(CFX*-HV>^)GH2,JP
PE"8.$^K9-"S&12'TS9_.JYAQ97&WKY5W-<%2RX>3MWN3N_W%P3SL(8%,SCJ<BM*C
P^$T*\+5&W@00U]B8(:G7[E<8!K&CYG$0>%#M)CK?W/LN+;XP+0'3,:%MW43&TB6$
PL.?4LQ;.K9OB^@&3GGM!4U1P]:+D63*EJ0EI.V!3>L)S4;'Y=/\)T7:LQ*0=^>6L
P!%"2D.QZ#KO,Y2&_D0*VDAZ7!6%_!+.8\<XRG?:F$U6J7K^[*EX4?4[6W6>F[:="
PIAG?DY>7MOQ5UUXQP]ZU[=\O*/(&O >ITGCF,IBW5"I0LS6W;45J@B\:@N.9Q*?:
P04CD[;/?FC47,U1YKCYT(>1W-: >L8@4,#E8XZ4_*=FH;!=:[O2O@KMMV8IP3X-O
P_<H/WQK+_@UWJ4>PLRL3T>&1:6!!I'.#RKYNCI&: Y60J2H/QKKVP[#"6<OTZBQ&
P\Z7P<X1K>201",$8)KT$TP\G3OLK[$<7B?Q75S-N!R6:?\[4/547G4]> AKV!WI=
PM<SM_+?G 9OA8&%[4.?=^_;.4HM^]F_<;J  = ;R4ZHY!,AI5%:0D+T60%:-G3.2
P"-%=9GL2W&/SB9?D8>()+(5U90T8/RX0+Q:E,-&/%XKCW8Y6K$MU.HVE>?B&K> H
PM<JV-_79%]]^') #M'#^!;!YB^)^9*KT [U0K*[^32:+_N:S6<E=P\4]^0D=#FB.
PL;'(NP /[/5W.I[+_[1I2F=@R /C27$9^#CW.9; T-;8:4/;.=,1M_+5M.[B6<9]
PCYU.TU\U7MX@QUL*25>%%[\I>AP@Z3=@A3'  2_!3@^YE6]FHM71=2A$P^C];&@@
PZ)-%_6\_$!F#(K'ZPUW<D<''#=\NHB3^'CU/'^XFE=C+[>8)090"Y\O0+:O6:I";
PJU%8VOLH2T&>01QSK^85CI=N='-/X_0) .(&TA[#'O1BB,P@")L<L.>/NA36WM)1
P.&L&KRZ>:;2W5'XT'A";$E>1)4(VW>PZ(>71G<%=R4@,54^27H-K,ME24+^(Y%I*
P 4EP?:IP3DUH+\8=A839%02LS0*C&$<LX0X\_XX4%DNPK0?DF('H$%"=";U<D,S<
P9).Q][R!Q%'#"SY.VBJF!8LZS:/W.#]_"'@<4]XC_9/GU\D(*_(-5K;.FH1:5I%N
P04YW/29%+W?SL(I[OC4/\CV?;T$JK3IJU=R8#!<S KUF/$CC]!%,15/J(' _M>B*
P5*F)>P2)E*'VWXJD/>:"R=?R)3IBNG;W X@T3?R]BGQZZ>1Y)G>LZ5_QQ-^^]')X
PESN8F$AV@8=&>9^2"KT,<[F9<KO!5/22LJK?(E#]RW,(1'OHUI!-^?^.A8X<H!*H
P$ S%+%C++'S$5(J*:25C?#2*V "9B:\OZR*C3 H8[+]/#[;?@-]5?BX$J%)DD/-]
P")6Z@[;I)=+GUISVSQTB',A2Q[EI^^0^Y;4VG!=<P.\'ND4O6*-47<[<J'0*X-V^
PU.2'E=0AU,PSLN<7I5]"=X9B= B_O(LB$'D1B?0(JJDJZ1$#4H^2"2<['!V G@]K
PPB(,:@E"V^8B^1-5J-/2_.(F?E31=/ ?1@TXK*:]$-'74>\>J* 9W9$D5+2TDX<O
P<D?E:Q=5XR@1E^V):K35SM9 CX)0D"REZM[5F8R=25JR\MCW"*D:R&Q&-K=EYA/%
P<:RRH%-"7;H '^,CLK)Y&W;^?D%D*1P*&%_A@+KZ)_JF'L.8[HP-5A+#[$4#N,V@
P/1A?'\V/1I3>:/BQ0]W,Y+DV8)/@521U.K&["J-W"_NO;_'%4ZHY)>MFS#N5]K*A
P#-%G2NYG^!T!Z'5(C_\ KULV1T*R;ZZ<@=( R_#!0M.ILJQ$.-'2TDH_:\J_NG@A
PIK8A0Z5J\*@5:R;X#*[8O\A&YNFD^F$)'#_K;. MCT:>Y;7^K]_U]YD2T'&.14(;
P:>Z;*L::5S"A9'=X\,WA8Z>&LHI7C"NL#F\F3#P)H^'2RT<A+LR*4#UNMRCK#*^8
P*V;>XQ*8U$5R/A/L.$*ZNY,V*>PB4/U&5>>W\J]7CO2>FU_QBN3FE1;23#LNGC\%
P0:[%*E"*WIGTC%\^[N;P1GKFQD+O$+_;-$.M@AS6LP"9],05(][8IN2WRP<U"Z6(
PO0$.7CS9Q @D4X.EYCTKZR/?#:/O]Y-Z^F*0S1>0_K\XO0)DRR:OB1-U0)N C6U-
PS\S4YM#N,O-$ 8)LQ13ZMK.U!HS8'Z\;N-CZ?C"<[^!@UG!_G\(&QHO^37K$6+L'
P[ISD94S1BP,PGI.P.?P?9NC5"4(GSTK/2![F)Y/QJB9-&X>2-Y@-]O&<?'J9ROQE
P^$3?SR2)141#9AGY%_9YS'3;K2:V0Y_#4KC'[GBZU=037L^Z(P",)F$64R)CI=/?
P!C?"1_+5]TKPI@;1C3<FBB[!88!P7(]U%,M5N)D6G7$X*YZCPB$Y?,<L6,0).P^#
PE.A"\6>32Z_Y2BI'W'[GF*HR2( $!4_\Q3H62R0S%%0$AWC>F[<?L#D0,>:Z6/[N
P=-$$O5IT3?Q/=YCFPO[TE@S']3P" S I8$H$;P(EU.PP':F,W$*X<IQ@\76?JOIG
P@='4-*3$7ENCX+R_S7^XAX5]R[FA=:E4_R(V\1*0%CN&9 &Z;T8%%64:[G1&Q[!J
PY6[KY&I@*#FU!T'&B$\("=WAY$QC\U98^HW.K=6S,31G#HD&1H-Y%CY =U)4M\AK
P*C=P0M7<(Q@$S(1F2RB$;791JW@QF^2&\<*';)R=]*CNCF@I"@].0/T_J;.B;'1E
PFT].^HM_IO,>9,&3H285*<)&E+;TOK#QV#HNBJZ]'8USBI6S625>>9'S04Y6(!.>
PC-^HR!^E'[?.U,/9ZCPTM4L$M>QL]>(E@5+\8/CN3H:627F[SHUZ_MS1A)R_7.QA
P4T2 51 ;^_!;1[P@A5!)=G.6%Y7?F-\)N2[OV)7(N1Y[58(9S'!8CT(F%7V<I/G$
P4NS-CMOY-IDBHDC2"!V9M8HNRS]<!WE!3'/=(Z4'SXC6A\.H8#'5Z Z<R$0K=B66
P048?FYP_(J....V8^^;T+S)39E,6EFIKC[R^S^M*2CL#$]>Y"T!'LDT8H)5 TC>&
P.;BY38.A@5J<]F07$30VYK77/Z+%%:-*.\+F^9:7^N\*]?_L9-3HO8^PALIH8Z]F
P"I4P853*4:88D140X5>TUU>E!5L*7!%G>&B8'$',T^,4,5 AX(@*6%2#V 4_@."4
PML-)]> 1@:LRRM9)D^N[:Q\7%T5IUA37JJN%4X$:P<(1-Z4\-239I#(MDZ4[VQ<^
P_*NE+(4UZ$;#IE;'G/8\:A"-Z"^ES4H4059WGU)].J+F>*YN%URR%J;'A@U:;>@-
P_>#S+%,WQF P@&84G%?%!A86,#8^Q&N?=ZSGJJ&)N+(T/DYN NA0RIDI/.,-$!TN
P)1]]UKGL@L^(_UNMNP1W@.-K?T)=4;[QD0Q?W7M.1L)^AKV$K;^-1_J)6@UQZ8DK
PQ5<$3UWXVG"H.ITKX>Y]^"TIX@8K@-^1DA]=VK_*#F<U_!D:340UM0)2TA-9J($!
PIE.V&\P_GE38]S1N9<:>@_[I%KF8ZQL2SE^%(=+39C-_I7^EE!:TZ^1!&0;^OA\K
PZ )ET2QK*\NJMP5V7:)Q!V%UM?'2+OX2N^<7!0CX';;>E<:VJ*RMG6:BKW2ZE1^K
P/-SY-G3F?>>M7.%7H5K;+6:K=[#Z+GOQ\SJVXKT KRI&G^><G\'L0PI)ZO!^848%
PD_!:/?AP</G^S9<'?$2+D4TG:ZH'<DL+L&I/Q#5IO/:4_KHR,^G3W)J6?NV/-E7!
PX^7V=G-DAU@WOB6S\2W$#T*8E9\YPZK\Z2I?B0"J"4#\26SI\4=+6+A5[>9UFU-'
PU_A=1V7?_,B):=1<5L)ES3!&(;5$)0UDV>E?/Q^'^X3G&[A]6PX7*&3DTBZ0+WV2
P4WX@%!)*H#5'@H3<@'UO$2&_ ]BFC?PQM9MTOK-._*J$ILPS'>[T5,7JK>>5+SI)
P#FN_M71LD946J=26KA%#*W2]]J,0!JV.L,P*:E[N@N&!4@/MH$35TW;7[;4A9F]_
P#R-WHH"9Y=6=(EZSO505 EF-;=/IUSC*NF:=[19FL)4%M]_#IM6A]!!!='<M>1E<
P5SZ/"K(@P+-3']MA_?8"YMA<BEN0<%EJTH?02X.JA)$L(PG]](-FK )'W!@3%;GG
P!=7OED/KMJ NO[WG8QQ!?[&$V/HUW]A?UW]<[/F)&#69B"F 9JT8K"2[IU3>-)H\
PVQ&&.;[@L2$QZHZ.CSLHYX$R1<&%-HG6VAF).=;ZTS;X?9=.21!8SB9L%JY$RMA%
P*8*6CNX\2F1?[Y7&3Q"YS6$V)]Z B1$G3UKBP%Q,<K<J#-7<,K"RW!P<88BS7<6E
PX 6)@8:OH\B$/$*M/@4.3<OF-=CTC"?-"(H*75*QGD[\G F5Z4E=!.L@^3P4;2U0
PK)76G"^A=T/\A*930Z7XX9,C3::ZA1]H.5X*BFW/*XX8DUYU\G_U+9I7R$WB&D47
P9L-8!)A>UE^5>UI]/C"-U+DJ>:HLL-G7YI],_4[U&6W@[6G!1B;EO<SIS47J P0+
P9S<??!=5UOQ60I,W4Q$A6&<<-IWW<-_TFQJNPE$##M$1&VF$.5PF Y-LP2K[.??3
P,9T+10];J,"%[H7GFHL5W93:79%TP?;/V=(K]-,'FZ5YN ;A*NA(5@EGTE[QOI+Z
PY&"?N8G'NWD7_)_ VM!2WN*U6C:RYWDN)C<]<^RI#-47[#D/ATU!V=PH8D!,A'E9
PW\9\Y---PA'\])A3M7$R.I%SC\N) 6;2#.4MK:FD\;[\O%!OEAEGFR2)3&OT(CX&
P,G1@4:= ;/MHQ/0R(2B+PCYCZWO*7A^F<,5G/P5:? !\&@PCWK=[X=:IPK&!FISG
P/YZ;.HC&]AA9OGT3R!ALB$D#T+V74BF&.+LYJQY;=>0'3_AI?*/YE;3KDBJ%Y.G1
P=0@?W=YADLHA^U<XD"MRG=F80&6@(D4:TCU[&&="?\=_GOZJM,O3='^NI^5E*X%!
P?L"LKA66\J4;3S::).$MGQ7PH[46JVO1),\^&QRZI;660UOKX=[=KS5'R]+I-P?7
P-9(EVW$Q"<MSIHA!BW1G9>6,M(-#6[I@F,QQ V]C4Y+U)6L0 7.@7 !,U'535PK8
P='YG>E.5HJLIA<//;3;F4ZEX\CE"K%R[N4 AC1=U\65WWCV )PY2**RN$C^Z^6?!
P;#\,A''*^F1ND[81K03SU]KBM(5K;JOP\;XV,$?;HAM/U:!,@\9LFVIO>ACV02?>
P&<38^N=H)])R(FD!P<I/>Y*3=J/U]JV62>RL9V>8*"LL6,V-1H^ R8TVB4 <3G[V
P5&5V[V_^:B/C'>TO2<SU8 X9.4\*)#&A\0%9A1F\JEX9 .EULP5?PZ!F;>,!$(-'
P(B\_':,/JR&G?:#T5>BM56EN#]M.$!>_L1+1:0'ID5F9QBDW[?TP]<*$%7[5*,WL
PPSCMKU:=<+ A%XEZ:%J=/%F<&^?D*-I #7,+UGFY 4F1.NE,<R<H3O,0DA<_HR4W
P )A1;9 (K(4!T^!M_AT3L'$$3DQ*^)T-CRM8-8^/QLGD07UJD<H[^2_WSG?.O(I;
P3*:DD8]G6/WO@J^"UKJ!E(D$"/G3CB SN%,&)08W"-V(97T_X-N:0[$8GY3#T\KN
P:T+4] ".YD.>L?B4\CIYY2">%$@OQC+SG4=B#?^X]@G3:0WYXGG&0;'4Y@;A-/T9
P^I(Y6P+25T8Z%-$NQ-/4@/Q=I+V:IQ0XZ9$^/2.#%KX G%LL4B68?5C=1"%]8/D@
PY='W,8CQ#0F;4:R=5K4 97(S;8%R0HOY(AT0[]M"$E=AY$^V/EM502NA<X=F%Y(B
PZ#F\4@7(S"7@">Y?1A:W+VJR#=F9+K*H11*P!0=9EP.FWDN^6 4 6N&*N3S:1J^J
P<6-I](G.^N<>A^^H,"^E:L&;CLYTPO#WU8DWX*1 +R-YL[M*YR"E:(."P86A4"5B
PMXF1#+Z)^.KYK@S!'"'7$X=:J["YW%%RT5AF#MD3OHSES0>W^XAZIWD M\+JO0="
PHFCH#M6BPY+:E1X$!O?E,626(\JS5=:NTH8J&Y2_/7 _Z:D7^DW@^CZZ8*=J)8;$
P@.H&71I]19Y?2@NK66GI ]OB=]P.$9[:]3WZ(4?^I)7(3QYR3<^.'VROG(3S-N;5
P2T<I,A RT2*V?0V 0J%"Z5E_WXC01O[_VD"-N]!^OEJ@%7;2#+F!P^KK'D_LJZJ[
P]S/+*FZZRFL*#B'>Y*)!Q;R@50*L?)>90)@.THK]Q$^F.BI;=GI, V+5]TW = *.
PZK_#F;^()AF@0!3=#M5'7YXMI2G4[<R6Q!NAQ<NH:1ZZP^].$%ZP+*0F-C F/R)J
P9>L= "EI\6H6EA'!I_K[P,&4"0Z,>JRU%;!NYU$XZJ]P91KS;N150J."00%@JA+"
P(\'QSLHC09>XJCB67Y]IX9'&&:(J"G^U''DBXH/5X"B-UL'(\T4>8F6G[&H5"PT/
P9I-@;%>7D7,DL+B;I@,F\:3)J6!\Y\%8<O""):#-<]4=W/ZL=TCJG^"(2Q$5*-W;
PBCQDY_"%XMG^S;6.TD6_[GF=Z/LT]D9BN$SCN&E7FO\='X0);L6ON&YA4-- 7TP4
P,S<_O_+\Y8FGL^I]%_+;0T_):]PRVTIF,)K3JU>&/6<L(\Y2/CU[<^,T'H%<;IR!
PZ%].[?/[25>9MR:JFUJSBH%QY>:HDT;1*S09=HOJ)9\MCBVR=":.0<AH0.=KJLZO
P<#U86T)*'>](?MLQ3BH?%IVIEP???*-76E78_1=BE1RGT^>;7$U[\925K)"9HDU6
P7KO G?26R(5.:';(=.Y#OCJG-:^]J@]E#2N'GPK]M[7%9OQ9?]!11I,UZ#(Z3VI$
PZ/U13-6"VF'46<<H']#56X4Q&8$AVDO3??EHT9>J.EULIY1SH@!:<S4UVHT@>C\\
P-_"L@B\](3L1TN:GS./I-_9_!9LJT@,3 JEJQ\!*+-2BN=1(%WTO'(^@'O5H56Y8
PY"$/$9%8S(LBX0!WS>2X/T#AQ'M'FU]WF-Q/,("!Q^#L>JO(XU3-/*_(D.DN9M((
P)S\8'OT8\(CUQKAQ?[JQG0I@M" #YZC1SDVM39_\J5J$38P:G\M 6[@&0>TZ878M
P^+D'+).JYD5"VZHVR?W5:X$,8&;T0OD>.9_ZW!7-:-1?/O":Z<X!PHQRUA-!75[X
PZ-??^GQIMG+RATBS*UUN_8C=4/*&S^4Z4RKIZ!$4()HH4&?G/U9282J?RWES7E;)
P[%N _/%8(XQ2O/1JP>X/Y2^9N:/.,KZA\52AU6FN N:1V!&E IYR0NCP+-/*> "'
PFQ"5]PU"TG^@<V2;:J*K_K^;&E%PVNG7U:T.B:M(J8*0"1Q[&9#TDS$]&(G6 F[-
P11MR;CP#DN>SV+L',0BQ;+OXPB2:-?S!I.NP')U@L]@VL9&I'"ITVKKOK.BP\G'C
P8I+Q5A+W+ONAYML$WM&1 #RMNW"]L1K!PZF3@-689-^$F_FAM;!8E1Y0Z+)7R!XZ
P&F/[/"IIH<;C>C(_1@ SM4 V,]>J4VW([:OFQ.=$#K4V/&,'&5!!?G@"U7S%L-+*
PJ$0@Y:< SX$T('.,M.(1)W%*63Y.)1BT[ZXU!:_>9:]_O&!4[:YOTVTECS=C@>M^
P^8L3HLOVL8X;_E,C/)=4P$'\1(Z5-QN@,@X%_.NB"XK+"EA1_K#^=Y*F=MP:'_T/
P-P6R#6KZ\5>4,)'UI]UZN0B!B%K;A1BFZKV&H:N:6%+K7CLP$F-,BTA9@4A^:2JX
P(F$1JI3>D#"2!9I/SUJ*:TWUL];B1B1_E054<Q^'0A[ULYNDW[=820][Y)?9A1BY
P"69E JQ3_?8^&83 J_TF2%+%4U >+VO#,VU0]\)AK\OC_#_P5NN4M53,'[2O70UD
P4#Q-6@#4>RQ9U@B%#."AOL;_* OJ5G.F90T01.+0;@0]J?8-Y&8ZW%9-F&@PGN/(
P;NQ=D6V:P1M7+$]HMEWBS7'<<[:O:I/NMFKZ5F%%:$4VEB+"S36!J!O<!7I+3=&3
PUR@S4"#?PNET<'V(1&]7N6HRGJ!_/@@Y6;*PW$V='],EKVY%[E-P(2ZKE+W Q_O7
P?DLV7%(T9%RFP 39;I_Y%!FMO=B41@[,[MWZ"!SGJ).D1,M"J#BYD$5IFOHATE,M
P!U/ZQCE;;K->)[44:P\^;J+[;BA1 L"N%-17H9)E\PC; 5(Y?"-][ELKCK!/+RQ-
P<QH,901T2-4"$4J#0S+>_CTF)]U)/_GSHYQX=GP$S]R(_/1*O(9J2=D-QPY?7(:I
PA:=Q7"P"R5R'/<.N3D]RUN*K:E DQ/T2Y9&63XK[0*#,L-R( \1,!_B7Y&1Y)J<$
P%3,L"?O=/$K?A&*>_O$M',G3:E:V]/#!@&:PWP3N8A6KJ-2JEDSV8XHW],_@+M1?
P%!1KFQO<"HR5KELB (-M<3PKM/5>82NA78 U2LR\3R;;SM)@TI>14R50J]KQK1>5
P=]6QU%2/?9*#]Z5@W9$RJ6B>A]@^TB9P\,BL\**D<^/O]Z(\;8"OO&U!"4$ )O;E
PL25.+*:?Z[0$J%P<04\F=J2\V98AWAR21 W&E_'B\FKZ3#WT3CE-ZQMXZR1(,$8[
P:#V98BP$7C1MC2:&(C@IQ ']@T3;@HT[W5'CA#Z'7CR+U3<I@R*Y!J-P'5^TO0_5
PGI<Z/NM=]KBVH]H2*7$G#W:6TFF9]QSN"L._N^/]THVP6P!MZ!ZQ2GT6J#>1G)K$
P>L;*S5S9NV(&0R;\$&*MX5D(LQFZ2<0NNT 5=(KG4K_)(>*9DR+N2F2UT6GW'F^2
PXI0^ TYA;RBP(*MO!T:8,X+:H]QAB":E;O:S?^MZ)MFV:(M/U]>"++KO'5JP>4?@
P1#]L5#'7P.%>A9G%&/*@B[>+0UNY8LTU7]@Q7)"G$TZH4?=(7Y/\'B<]!2A[OW?B
P2K7RM,F*YH%(/$;C[GM-)B> [".6BP,7<>@>!G9];:]!4#BM?0E][Q&$P""VN LO
PIM/@#7DD0;'H 7B4>]Y$NBZ(*>_W2HIZO0)[BUAU&S$1T"'5(8(KYK<.-C[O:ZZC
PYX+FE*\U98EQ%/:5!C*<,":5T@[O^$TQ*6OBX!DJB0>7K/C6SCY7R8+0N-\(3" 6
PY7AXLG_PF& B.Z4PB/C-&GP[9* -)\H&KP2_/$@$R%ZGN 6"#J^UWHYM%G*/Z!D^
P);S(R^,,^&1\#IR2IA#G+J<RX!UJ>J(Q5SFZ?Z(5TZ1>G<I/U9DKH298$7C4RCME
P\S9TWN%NN,=EQP B#620\[J8:>'W,P:K[E#EK3^Q-Z>3F2?L@07K*>7W,H@GE(GI
P^<HV4R-^ZV)IV?=D/0_;Q=Q*"A6276(5IC.E<X.E+TQ+XG@94[S=KDK6FY>N41[K
P)ZI;0&N,L5#I!HGC?<H>E2[M.;TLNPY2WOFU:DXPUA9F&(BYU'?Z,OEQJ(.7Q'8$
P@3]F(+:,HBFVJLB<,('=5#W]<6HCP! ?#^ PB!D"/KEHHL6_4&! K]\E>RL;YJC]
PZ:[\&"Z_O5T5OT@9F BUM'TUR, ZO9:)&T+ND?+]L-08D,1X;SBPP3= NZE1RO7I
P& N>D;O]+"(10]_4;K>ZQ&9@ FU[ZW J,^S\,(YRB;G$.U"-$*/HL.4&!<45DK%K
P1&JI1\!K< >YS=F"!@1#L3*F7$9@W&]< A;XBQA\DHN2$EYP 372"/*NEU'CY%JM
PW0'TF.<ZEL[!PZC^.F]BQ4.AFRO1[)8%%@J(]:F$QSJ'?*NA[N16!R%HR6+HA]-V
P)$WWS'CT5<]4(TGVK T2XK#Y@W-O_/\HR4)2^$T'_OQ;%2,WU^!PZ>'O)WS3J=FI
P+#OG0.45.N[D.M'+VW&_VTSM9@N]*]RO 0(C7EXP*D10T5S7'PMZVRYIWUEGXW/#
P)X#,<(F;X"X JO!*;'13\SCWJD%N6)SH9\"%FWNXP[2C18#'Z&K4,G*IWU,4WJ@V
PGNP/%^89/;K]F.U;?'"#(VA%[&8'!(%I2IA0K@=$Z^T8U +@PS+%60/#4@X&QM'.
PE_DX4#^ZBYKI 0_H845G>0^]6R5P0.>6&C)B-I88K2[(+'F^<4E"B?'[WR./.@KL
PVDXX7[7J *'.]3A8_.@3IQL9P5&TT*<-D'K-K-' .<1-O'DI)LO0H7QWTW?J9!0M
P)'8@8@UI [3WQVVM1-;W&N)AM[N2WME5]C*$-V*#6NR7CPZ7 U:(2((9?1J*A58%
PVQY:)UX1OZI5*W 4[]%ET('X;KM05]58)?(6/KO<6TJ3RVFK_E>5M]5CV$X?<@F'
PL;AB1]C,?=LP*(OFM_;52WD$BHK4B#Q8BDQ/Y_;+A?GP-?D0UA[H3EC+(%9?:_-U
PH>MR#'TG;*.?G^?D^R(U NR/%=?JB>;K40@7EJ*-/GR#'CGD)PEN(8F12 D1I6#0
PGF(;+*O?,/R1.!TC79.RY@41T9Z6XADM*V[O;96]F 45,)C";2WF#97-#2Y/U#LB
P]&["/5TS=FC-GR@F]Z+6M.R^866:6ZTN9WF8]Y >P@ 0PU632#X_APP9'^&3M:"2
PIZZY]I&T+%#1D(W;UHU>P[O]UB)MWM_^*XY,U@(A5%";::]7R3-Z%495]^V SFB1
P$E;#V5*>LA;3N==50:.0\G0!/H-)XM>J)?<:X6ESBF<,2GMB51U4SDHH-@C@U74E
P82@23.K^&(@*YE9\!16L&:AHI)=![;U5;F"+'';GGV3Y <F@^K3^H!1OAI2(Y\,W
P3OA,5MN#P<WZS9'J;Q])$V@/96]MQ.PWM_\KH:)UE4:V2!$2_L#S[A23R9L\Z/D_
PD@,::($.+(,NL:@D_DT^".BFFH ^@I?,5U1Q>]X"YV.(SL;FO2*OK6H-2_#^&BM(
P(.:%:$01=MEQ2RK'(:5_+O4,L:[EHN28(#G55 *CC*%2W=[Q'OS0;<I3^VO1F0&K
PO@9.SV@UEV+GD.FM2ON.*7;P08<=_\RAO7 L-ZX"F:)\!?T:K&B<&$$H\-N'EX(8
PBS\W#H6P>AI,!-02EI$<3\0[/"H?4\9W6.F]DY49!D;G"X3?;7(=<>@3ZF.+.)NU
P1?P9X+'[-#:M%I*X2M%?%2#'R#&^':T$:;YRC3 BL=G,3*T;70&G&N%@<@<%L=*&
PP3U()P[P'+LVQ6>NRU'K*1BOBVF:\^D55*9D6:"8;4<RBET/J$K_2TCMDVMU>=W@
PGJ'1FH!X.K)@"T($-V!#%\^;!7[<V[++(E?GCTP16M1D!B5PGSFWEJ8<JQ0D(9>9
P*1-^RU]&O54FO.CA^2K$;UQ_<+'[N9]< (986^344+VW6_N*8S+)S0%UE,VG0!![
P>B.*_=PX^!&9$]F).[>?0=D0\%^6K"]NTX49KXFDKH-1^(5B(A.6Y[YL'=WI>)I;
PRL#6RST>1746M4X4%VG2T$5<)&BND<X@US/(N\L.:Z3.(0SK7*LTZMJ1;MYY!@LT
PP)Y1\0N!?2LUQ%!_2,8JKG$U('OOFH'S#35(!]H/3H'E+TG2884F"$(=J>AB#,\"
P)#374<8%ST!>.U<I_@WS--,F(30:I,Q LC5P-JLU4CGG'Q(IRU-^\C'_=CJR]? &
P*).JZ6P(NVB1B2JZ]&<J_:2!4A1>:2Z]$L+Z*6UO$4,DK?^8+1(62^I.VQ+OYJ%H
P<K8?=8KD""9N!@.R*9DW<>S9\E_ZLN9)H'!U4U_3%I*70TOH'SJ@_HD %[@SKW"S
P/0\YD+&_23WO-SFEB0'<HB,RCH\8L^=SZVZ;\B&)<TMJ\3)3B4=[L[B&7YR3M\D.
PHWOK7D$-.3(8!":XM#_^#&2UU VOD$ZJDN/G]JX\;I TQ;,&-2DF1DY)43\8G/GE
P7E2VWP ]>DRBC9Q3?9ITG-A H]EZ^Q9:>J6,\L)]ZQEQ]8#484=[PT=9 QTK1&5\
PUCQIB*1X7N4X6-SL_297.#%3%!G4 D*79K;'M8;++Y6S9)PNZ+Y8Z5+ $KI9WQH(
P:/<2T*_$I-]F/\5UBUS,X)EW0SU5Y<5V9)38OOYOO@J.&@J3%C*%'Q0]F?D_&R9)
P,X:#.;T_C![C'4@>BU>7PM/K,E*DOBA)D<?G 09'K4?CY/=K&6"LA%'I_A]94AJ&
P.C\H?)?_^-#G_"A;%WJMJZQJ(++@@&\&JLJ/5HF4;L5<<BH2^H&*KCEJ@]&Q3POU
PIJC$#;T\Q;?WD0JCMJW68[AF3/"297.FK0C2]-)= LU&4J9P"Y,#.T1 YW7/FI\I
P<\\CNVDE5*,LRU&$NHHJEBN#V!F1J&W5VK->E!+6*.^H<^8$S!F&2@5L7SDZN4H1
P>XAHG4S4*E.=TV4_VQ&5JUOB25/(5RX^EM10N,^",IJ,[_J">WO?(I=$LY'9309N
P=;K!2B@(7\/,,A,3B87=XE$G"X8"I]!$9AC;3A.2(>:8/8,^D8Q/[[$%:V$0FB)F
P#:)(_LTDT#(3*'O(;PVQY6=E0W*DY+ M,+ K)?!V!(\&']\A1IGO2"\G_<!*+:Q<
P*>NR%E8I>S8R241/SUZ(.G<5,+)2Y>PE3M]VNOLORX[>(/&2&K)8!0F)]15;+(""
P/(Y)]26OYL"JSZ796I<O4,[%\"@*80?L_=*WY5[]I[,M8'V;GY]%*BT XB8!27*=
PYD_VEY!ZC*1468+:<Q-5$1K(JS(-%4CP+<)"VX(;W-PZCX+RC?O>N18[O2^NQ)7>
PI5N(F#(K1(V("M$N)A5A?)Z6]$U?D"4UU*.R&YU(YF[<,CLNW9.E)#Q ;+M9PPKB
P.%/:_K>V0.. =X]R_9=(_&G*V\(\_MG6)K5QX5*,+ [2?!6)F95WCVEL;/A*?J;'
PSS> JO ^'(LUA;M).@L6B,\Y,P)>BED&^>PU&'KC.,?]<Z_S>+,,1W2(8E5CA,]M
PO568-"S2@(3%:!]:4G F+_P*A_GIUWE3!#6G&H6/Y.<=6-,LPD 7;G.R.-7V5=[)
P]H&U[$<=_7MRS<NY)2*\RK<H0-%_+!KR>E$-/I-RT66 RQOFJ>_?&1*\"D.QU*.7
P6D.+\33;GGYF;?P_EDMRQSO=!C9IO."C2YV%FUS!P0JVKT[Q-@.$#-8F=-TA^INW
PLVWL"?ABQ*J#_M8A/&Q*&1M;_(0V76(H*&#?]V!<_6#G(73DL&W9%O MS6<<^3J:
PO1.^TB \#&U]<.O77"VBS<E'=8&KD'@]6F2['ORKS0/H;AC/S!P&9!>/\HNS7Z-Q
P0M[[OV U^]5#^(G(XR-TK_D2$N(#W*FM+RN46V^*+?<@LHX=1#3!./!K\Q[(,WX8
P%P0U#&Z^ F%??B5K4/SFW-.-;XB(-:^S[NS:G6)9HWMXL@D J)&X^7VG'/]:LA(4
P.R8-KP51YU&4ZWXT, PJXQ3!@#^_0HN6QFYD*$-J([8/K9V\A5YO>)75I")^K>%6
P@ZT2G%M2G@3/GHF:!NHB)Q.12D=(B>D0O2A6'=3&)2!&FZ_(8WR1:6<\@$V+>56M
P=Z6"#<M2Z;VZ$1?P9D1&/+YY91,+H#93_XY$0=?OURZH;X/+4SU7;"<D9Y94B=;6
P7A"IQ[-@[)?D-XJN]'CIOB&<7_3N2/,?P.E:DW1>5F:Q3PU@"1147L8=#E:.D>CO
P^XN"U]J>+.V-KJG:PD>^OJ&&Y()JM-G"WM*37S%O$991:8MKT@AA]$=T0>CI1Y*\
P7G<H!W8*NO1![X7L#HS9 .$+/ZC,Q=20V8O98<'3AFEN1Q:4N>H/QCL/H'@]D/I-
PB\@@M\._H_N74B4UD6_C'L;I7OGGZDO%?06N5\)F\+U0+J-NDG@HLRGSW:Q,DL/$
PJ.: ]:7:D0AP8S]V*S <!A?U\[?A:Q32SV*GFKY3HX;*"OTDK(TQRG_5H 6 [57[
POPAKC9Z.^%-*IXAV/YH')%I^="JEZBBPL2_'CDCL8J]5/;OH)"!/UX1;1$G*0,,[
PG]T:N+[>1U$TM\0A'B"Y\@0$9.!HT>0>-<5-*J!'583"!^73]&Q+K+-[>D2%$X.'
P?]=<JV1F7<VB305'M^WQL,@F R;6'EUBOA>QFZ5F0>FB(#C0OQR-)@S'Q_MFK_;9
PN#VIK_ &X8NFDDM,<OC-(!E 71ZY9X?.?)\^-MJ >9O'7*27@ Y\;SM/!&G"IPS;
P!J#P'MF^<ZC2RP@/U777/Y!JU:Z#@PF0ZL)+&T2NSKKJ:#Q=_XQPW<Q.QTESS4NQ
P+#2''UGL?(LY.18ZIH(WKERN@MU #B%G"3JWW4-< 27W($3GJR:'R;%,:D;=AUJ8
PXM-)F<A/S32HA12I,Z(T! 7(5%]8IRX*1Q'!'5Y#AQH6UZS<2+HF%!@W^W4E3Z"B
P/Q:CANP3\^#%)AN$Z?WA&IG/JS"0'2"7T#<:U)99G0;>DFTXF,D?76U4])2$VF I
P=XGS(U1P#5!34R='%[2A"[R.$1[RIW^>U,-;8W(\6%QO1%L3]I$16YI+R:Q .Y)^
PG4 IZC#W*^F"I?18P3+-+&E3 )ED]<6AR@9U5@+$G5)02A*+]PB$<"P:E*:WA<4S
PO,;U@BTL$IF0[6M_D1?SS]T4^UWPS%P@UEFKR'6OPJ+Y5S $"57L[&FYN'K^%@A#
P./=@]*YPA"=2!(88:K9HP6Y\(A*MX85LJX68XHKQO/YK$UP!OIIP8 -Y!P*(EAT*
PBQW"F4/;;>P%NN'1"=H?QSJ^@E$B,=MPGC\'O?O-YO#\>9BM.E3N9B@G6'35UTS.
P\[+:_-Y7(J'YH<8$4\==2'F1^T_%%YP8SFT"5=_55))L]T.UA]@F"QVI== FV*FP
P6'T#7_-]Q?J=H;Y&7LSLHP5:0(:U$4!8[]B/001)L!&^?SSJ;].X]!U#H8J9O^<G
P6D -/(^0D\E1WFA4S3B;H-C:;VX$XH/60H^#AEZ:?NBI-5%S6?#Z+YZRU=G!8]3F
P,U5;<5!#V?64UQ]^*B;AS[)K6W9E77]9>6 -Z4S+V90F*<B]J#\2#_KGC#OH=FQ$
P]W(&%EA-I8[NB6W7.]9CRAL**D+!V&[C:2\OU9)">."\NR?Z$==ED>[XOC:E8942
PUYD@NZ?14*%E%W:O<O:;]PF4AMWD%^ )BW:CX(>9((FK9GK^V C8*;5H(?5G)4#\
PTT()E"H>%/!=5"_?0DUYP*5@]D/!1^K+$CL&G>+K?#:1,R5E5=^(8ZA=*K#7@0H7
P?J]TCJ[%)0M.34LYGV3YRQ>6I=7S5+>RHHFBQ6:[1.VPP]Q$Q6 Z?UO-7R[]?CWU
PA6/P=92!#A%K+@$5!)HDQL9@(&4N.W<Q&QZ.%:V+JQ+'1>:C=WNP@C$"]G+N%/<G
PC2#$Q*V[;$=8A#(L^5X)CO7XVZ"]03H*]-.$FJ_NLM0SL6WB(X?PO^JV&V6C;'I!
P>8=[+X8(\*+(Z>2WP+A.SS:X4S) [3^ _T@*N_!9KDK-.O)GTL0U*7MP^8P8/G("
P':4^52JZ ?6/>#+H%>>?S^'HWFT]]:*YM[.?U\-ACP+J%4(W1QV)?OW]0H.L5+[E
P=2=O*HB?1[R!@X,R\;KBW1R^>_N@\_HH>Y(FO(YPF5RYD.#FH%GK"RU^O("&.TD=
PR<4)SP?SBHQGK$OCYM!, #>WA\_9]U%5=#BNHB7"%CA(U^7DX_9?<$:D"Z^SIGBT
PG+D;M-2U?H,H-.VP"=D*'WHNKHZ!12&V,\N&V,#'O62PFH;O+DQ4K[!^2D$,5<? 
PA\?_C5TW;@B6Z4=BP]B'275 *@:82-[K.0,B75@7'-PDNNKC96$IJBE^4RI>)8H3
P+N%V6&A^O$E$2KP%UE9%?Q\7G"-=A BM]H=;'+% J40T^,NYD<,U[6GU)$<B=/\O
PQ"*K##A8??N#Q8C7;BY>X[J0W%A!,,[;FA7<IM$)KO["3POWS#V_<T^]E73R  P 
PKNR.B"27ZH*0U#3 :  &L2 6/-;<<.Y1#=-L0[N*REA,#?L.9[B?=Y8K6*>Q!TN*
P0CR?*Y2< :9;@W0IH"]A*W %P!1UHFV50KT8YT[7,\3+_8T[@1$HY_H@R5\ <'H7
PZC8_*Z);ZEF\M?1J!!JIH7?/WKA#O>3KP>5RW@^W2=RHZ,$<A0<D(V/!\)V/8&QD
P.(L]%M]QUZG\7^D&)_QC%)NP1HU$LUJ7-2@+G19M1/NT(OHJ(KT(SW[;33PK?R#I
P-+$&5Q1EEX7E?L?H6^,S8&WKU(ZG(BO/X!7R?J]?/32-T"10F?8DX>A;6\D/H:(0
P;]!B>-RN2KXMQ%](3[Y?F-@X%O@.T@IYRXVT<R13M6 3C]9O"S8]/?L#:N-#2"-!
PH.;)%B@-.4]N@\!$9=Q?[\RBT1 )'\;G\K]PC3DSZTC::!F1EC080O]&A*:580$>
P5$:ZO!' JSK?^@3<_NR]3J0X<9_S"X":FP!PB%4#\U]WD.*=&?@6=?*_MOD_<)KB
PXKC=U%#U6H;$+J@BY^/E;;=@1WJNZ-^)<A@'7)& AF.4Z)LM,I=^H9P-F9F&$_/@
P[KO((8L<PA!CL_A%F@<+_HRZ\S)<O7B[@'*6P^<NSQXP23A&112^/=-@/;7:/3& 
PC\R4T:G7*6U[S'H0O;XC/\J//K.3N$-EDFJ5KTFD4 4N K6*%J#F[EM@%AES &&#
PR?5E.B'=?\$8J>X]$!)@88"QSLOD3<.<9V]?3V#DW]3['0M/"SPA%T./B$>@-.\5
P@G "]!8!:Z*ZEG6=4Z(V N@G#)ZKP_-^@T7V*MG7)'E*649KDWE<5C3=^SN0$]:*
PC,RP#U#+F.3Z6[I\^6B-383=E8?CA[M*1H1GH7@4'_@6[:!CCNH@SC.9-TR=(RIH
P+J02Y]HL9#O TIHS9IOFZ/&@;]O58/>_%..E1"W FCZQN=U?7+M$=XP4NJ[;Y.>5
PIXJ)H(#N9)J6H%<+?SO,L<#GIY<KBBV@'TRFH;^H4KG4I!DM4<]PZ#J;61$4&?';
PA$%@M%8<!TL.S0J1[]*N/L/V3[O6%<Z$4K9L)+F:5R'CRI[X+=BI 3W489\WTEPQ
PXEZ6=B5*S Y/AF<LH%63<5B'FR2!VR-'BD]372'VQJR%T;[EDM<F-1ZP,&E68>4_
PI\6GK<.N.5! YU6(<=$1/\W)#%5:?&E1:_CD54JK<SHT9,/.6S,&&C+:S%$YQ['(
P*[]-<<?71S*0'^P^<%S8CCCK7_Q]:*02/O7_OO'R%PPK/>HJ+W4NOVG<;1,ZBTWT
PAG2R;Z>H1<M?S^0PNCH+Y-%(=\,_";?2E5"3FG"!&:1H!P>"G7%23>R\UXG _PX\
P=4^F[7+/.^P::<0$/-#*,-I0HBMB?!R$>%>(?DM:'_0VF9N/&$I7781RM3GW(MCW
P?OXA%GWCH$S3D.]..9HK&S-"F+?-X45<E+#U0)]QS<2=27&'$5YDX,3YPEQ(!*6<
PXMBN%6-=N\7? H0$3#WBU6;,;Z1D8!..MF]"%V"*1[0O/0!E%.21I@_26/TW?IB[
PKT%[==)CMRHRA 6PL%Z%MPE:=D^M,"D)>>D-!G*:K8#N)XJ9?Z I%+[U2I+A>X&B
PY/&"B5RJH",3)Y%6>?2/S,.!J@KZZ/^MZ7I*>/^6Z+N9-#L+VAFD&#!\6^2!9B5 
P.4%DT$NP3)$^MQ1@!W$XXNE@];]P:Y,BDUYE\8?F^_#Q/.9 ECHI<%DNT;E]B\51
P^J^E'=5!6C-*.'KR,A)0U-*4)/L)*32NWY7> ,YGFEV[B &5WBAL(FLGKO5-)Z4[
P(@JIN/IPOS*($#S.ZP^#>1%K(F8,")(9!IG[S&:4?,WOG+"1IOR7./T>:JW#F8U]
PAJL=><(EXJ8KP96M"3R?[A^BRQU8?5R!:TFL;DG%LL= ^9!_/GM)XWXROY^."V6K
PSKRM[7,]Q%9W0<6Y72Y:;_9)4DC!L>ND-&F8!$($XYK4[TWRF&6C#K9B.%\!ZB3)
P:\X(W>"597&^T=G[C+G\)"MGJEAF(LQN4X3\QY'/$42ZVI\4FUEV^'N>L+;1[^C,
PQM"ES)AV.7 +,]T<!9,[/DX"XS%W3)R;O^HK^'QSUZG44B<BL+0]%+1N*PA.63X)
PQ/D%,E"F=)6G%.XIYX49(7NGKL:R^I3G2YM;" HS4PH/.Q8,]'O-BI9_VN0'CN?/
PS9>W$OG[>O<JI /7Q_$^WRJ"+@A,N\["KPU8)^( PPC[MOW%RV,D %DG?]C@&&IP
P#-ON+DOO\+*=1R].C.N=9?QVM&=>=A7$2OEVS8_TQ*>U:OQS;EEYA)I)JV-.\ZFG
PN,SI#.1)^PHKZ\N$-D140LO@3ASD>39Y 9(6I&(\T@,Q8B<B<$J_>&9A6F\GWOC-
P.30NZ2[9=4_C-LA+P;DN*GI^MIX1FH&=3Y!CFP8Q5L77\J(;BQ,SA-,W"06=96XP
P/!BR2WRMW-T7L1"FT3(ER>ASKCK$/?W!O&288Y!7\<Z?1&)0_RYT_.S5$P?F3Q-V
P89-J;LKIFS>YVI=/9R/5ZJ^B["0BOTUZQK-]=R];:]LGN-8>$YP:@IQD!+#UVE_Z
P,U\ST=@E1U^A*7>-MBCK[<%M0G%! 9ACAQ+,.]6WW#H4'NCP9N)C,!=^ZE38J6G(
P\;@^61]N0"29'&/UZP[5TZ/Q4 &/K26<N-2RI$6U+P LDUA\[<V"@-8_B>\J]+9_
PS3,U2,I%";_KS\PO!X1IDO RN&7YNU2YLZ IEC@X'(5FDR:U;QSA?/Z2;Z/, N9K
PH1H,>1<]!CFCJO"S^IX1=S:F;*Q$?@[MHFYSN^XV=\V)9#E!G7TX#32"M7S0%63"
PUU@M*QK#1JDOP%V5V_,>*&ZO\)X< [8%YPA@;=965:)W5WR76'_*QDT,WZS%<H6?
P5L1\8OX/0DC"S#V^2]QW3*5C1LM:(^26PF^V0@*(_)?) 4:Q,H4&HO!BBEW\L2;;
P="4FAP>F6?K,FG\'-5;#\FD()-1-^_.Q,W4(L+^1*!A)L5.%G6+T\TVVV^KF4/>&
PNJ^LZY: 11V2R,OY)#[ B?8YU\ XG$_IWS+8<Q9]UB?&(Z+JI#--]<N(.5@JB(=]
PK*])EQT]=52].J,* V@+$[KG!5K(2*.,4*M[5^/G PX>X#7Z0X4X,]9;>![//,*/
P, +E7Z%$X*+P)AB2RB<;)[F233Z*D=/)B/<*V\IW=YY?T&&*O(W4+'JR<\GX)QS$
P^T/RQ*+8*X)XP=OI^BG<G,(($K[+^'?JGEUR*=,PQO8_D?U#V")STX9X\^9KDZHS
P 5=#EHJS<1N'B<=GM$J-E1" ]'9!21+S/,RVYM[GS,T-% J-<7G 2RO+5<[*-<XI
P7E$/%W48G63#I&K?I*C@/1(U.L\]U)1GKIFABA4=9.;M&IO1FTC']22A8N6WFYT2
PD-['TW;KUM(78)B\?:^KMXGFGA=)[U^UQ=1"Q)]+B->MU'XYL"_?2S5_=]ZEO3MA
P] D!VO8^1_1:::4>I:[?^]7<'!9QHV5;B6A>)DH]H$I$;H!QX$T/M9'FE8"^X*M5
P7/%J#+% (M?L]QM+ZG+UX;D9B[@H#=@T!$[3)RN(S4TX,Z2<6<J+.E\G\[^ 'FJ'
PM*T\1_)@5R(9Z_=8/$BK>U#[L-?+:4N4,].J6/*_X ;2;G8#J:#4M>K>'IW=;4EL
PEJ"('&+]%/4GFN3P\6_FBGP3Q&3!6$U<6VRHQ_I\9C7UW?S[M=6FALV*!#?-<8BH
PZ-"O#+HF.X)GA@6)J'V1?@9[@L_LC3W3$:TWW"WQ)IN&@:*/LC*C:#,Q5H=I;YIP
P&$]'I"?.]?#K8AY5$4_MLJ.&H(;?<^#V\AD!:J4D8(/+%SG0,PD_T!T'-F?FA'6F
P;5!!6TV0+FV&:>MOS*4Q)L/!:L GY.)!1("JOT>6C+V53ON"T*.0_LJPZ:>MB*1S
P'7_*M;#I4P= )7I?A(XK=.6=41*@/):]G8OJG6U]UKON=96:3C?/ =;H4@@ ;85D
P^'_]QT$D^(C\-N2M;1]4EVT^*SF7'"'?311Z><-X.U$LB>4N2,0(\AOQJU23G!V_
P3#\ "4+6(1'<87PU-?;K;0"P-C3.4A=CMN[<"FG.96HHEIU)N.-LULMR0$O>,>*Z
PVUH5X8$%_CLC05D-7&%QX3$$WE_TH"+^Y-1=I,[+H9%-_PB@U4A:B:J!VJ&_JXR)
PL83%B]+DQI/]R""=$(1"06;1H0X."FEAI)X!@#EB@IUO,E;YOV(ODD6$,->7:,NK
P@ S>BR]\:'&WWO_TLO90#M!2-+:79: C,!I+,;[XA<CX-/45/RR<H;*/D_<W_T=G
P$9*)V0KTDLNL_/@UCZEIHR:/UU^7PL;[D[/2E^.!-$SF[D-S 70JU7!:.. '^#_#
P8O:$WCA3VIT^= K$7W)VDWG! [!^K!O]@1SR\E2#G$'D%F5_HTC2STT134M--S*S
P9LNJS+U6OHE?[4Q^8MWIB4F69,$.%^^1&"'"-HI!-2L]W4#F:XQV*M$(E+H.ALJ-
P>R.]0!W3/R@,T/$*M3^BO45"(%@I#]54^%-FT44M" .:VHSSD^$2]\%8<1: :X)@
PHQFROH]?@@X4"$8JTAUHK$KL.FH^SO<Z5$5;A-L&A8<=Z8X1<9RC%L%N0B(,MD&#
P$.4\ML7%.5MHV#!]X9H=B/%DOI?*4M V,B;])6 &#+-5^FR/O_.A_,EZ'M8AV_&T
PH.O]@Q<>*%0>ZW/0F8<E[>6<<^RPOX.]F3N &0'S1'ED  J\O[JR&'/(B]Q-_4!(
PF+8PW:=)UAC:4,<TPCH2[G]"?7$&#3-=QLB=N?4\.?5N3&:.\-9[5/'5Y<(\G>\M
PD]O+*5KX J)9Q_F^2(O\&[VGO,AV4F!0ZCI%*NNHJRZ]^.-T6Q7Z*PD.0\]+>\+P
P6*>L?2+.(<+TO@HB:Y4WA*9@Y+B/0:,2%4X?T22+6O[J@.\&92 ?>#2H"W"3_L$:
PT  %F9%E)"T4_D+A*1&;F>A4N_S?]01:O0U;>=E, L"<4['Z@F^6E[/'X PU$="M
P#RY%7!W[.]Z[H_TX7NFDR QK=J=E]/T3P5X/I4H1[ZD6J?U>L6Q;3J&@E*F[\^7W
PKGYB>D !9ZKSN/?=S-+ )I':LJ])5JQ.F2:-1VCVI\>Q!V#U4N)*X/F[PY>[]J)S
P951]'3=/[D%K5%TYV5&W>@(K4-P_272O" ?FM(&,74O;[RS 5-K@GI!:%L/ DT<?
P-O$B-.\^7%MFT1\UE;I)V@XXBC;S))WW&?,$1S^<D;H&C/U!6D&\A6;4]1ZO-2Y,
P'8(K-[0G;KM-G56V_@N%B&:;T--'LR4$V9"NLVIQ>:!L^S%2N\I9CMVH'XRHYS40
P[TRCHJ^\)Z7_7(=9-_L1I3LSN9=PO6W1V' RNDS;^AVG%><7S3M[=_DPE:W_*"'V
P*LU_F_*NQT^0];.7R^XO63D<*5<A+Z2=IJ&@BE%NL2QQ28OIA_XLJS\.48J,A_Q?
P'U95V)TZ'\E+_UJ W:_05ML:Y5O$YQ#9[B3GD+.&X#QK@B62LY$-AAMFE<I09D9<
P!&JV;-,Q&BH!T.[C!5V&?J.?^3V8SC-@L)#PMX/!$"2^C@Q[V*.;\<7Y913RO;4B
P4F-1BZ/< \97,T7&L"P8LU2?<G5_(L:P^+"CG-,';9Q_'E#.YI%WIC ;4>ZRAU-L
PL1^N!!K#4*Y_+,0QD:JGNYB985+6-HHQ<?.-Y*C.5A=$QG4409U*859'M;I+[ZX$
PK4Z<RR(_ETI41C.:W/:89[(Y;W1'24ZQ'/;(RT>T:N\[T*U>^CN>"(5OF\9L3=21
PV\G>-HPGL*##2JV:V*(&$O18GSLSK!B*%*N[E4 GT1@,O7$YN&YJC2G\$!'2;/ #
POYF[LZEN4:"-4\$#=UGFM^IW1YW-T=N'VPC2TQ+8C5+R;[E>8$_Q]D.[*=0G$?C"
PA6E*=KU ^<4'T0CP-YZ0:*Y-9M'9HG2Z0OV75'UVD'OJ&U_@8]=V:9J^6[Z>N9P9
PP$JJ(X/'3C];Y9$ATT*Z O=G<1K7ONC;GV=&XSH_L=AIV69SJ*(Z0C6)VD'%(E&X
P^RXB4I@#7[!9-CJ9J:[<^ K3%SSH'_ (!(EW#1 829+(WX<&ANDL12:9=9"1A9'G
PC JU%;,7@&RV-IPSK3^+Q68W<YDCZG:0HU%^WAS\O:$07PN%];0^!\U 6SA'3^UJ
PRX911HQ"ZK-1W;UJJ-%RB&YI FU8'7[=YQFT>'NRXQ/>^3PE-P>7;S<1]%?9I.7N
P\5!\M;&#]ZTR\!V3#8P1091,=)]"P( K;$Z8>(A.M$JD@Z+-NY:X1B&S(6W8#,Y"
P:>6=#KS9NAWCH-%5-614A%5>]%<C'G<2&A,-WBTD=PP%P,M)/CPW>GVU3Q_ U4<P
P=AUAE1< GXK0'3N*?4,P <=0G^L&I@N;K\?'*I82%6'F+5.%D.30X@WS?IWCOE7C
P/=.$";SYNQP?,LBLCC3RG"#$/:;CSOMXX%I@SDYA+>$1969Q8, V56\X\_:+3PB'
PWDI&: B2Y504;S7] &DF!T@C1OM5#:QC[Q>>K6$%?<'_@QW8-!WTW\.PD,8=Y68!
P4^87O<T+RD9U9O^+[>9YJH?:Q%7.+5U!;'4.YG[#O=+MGS'P\>/ ^#*QY0CJ)OC+
PME7G/I>^3<#'4E<)RVN,.V;Z]%/,_7_9BK<Z1VLH\OB4L$]O]6< ZSJL&HO%;5-A
P6Y-4Q>[P4<5,95[X <RR+@+E_G9B3'-9T<D$3&!KP\'_@-Y,9#2"K&97,RRXBYD9
P::5D. /0I4VK^C,85()S5']A/ 3 -R"'9-; FL^DG!JR_9H*\?N&=O1[^I,XOM(B
P0PM9=4H2/H)?MU;#M0.=%OY#RI*B^I02;)6@]S#,O:J[1NN&O@@=.'0\B_+[+Q]$
PY>*'?)N^=("F1NM5="3P<?&::@W'95HU1>A7F/55\WKE]M<4T/E^Q$@+7V6Y4AG5
P6Y4XS'">^ZW^!)!RXL$YZGPE=X/9JHM@3*-!$2!T'/;<XX3"F(=&*#F@0 AP(3JT
P\?G1:_HOY*N/Q;=]IK>H< U&-(W6^\G#&,/J"_4CEZFUS5W7:?%V<Z!D^4Y3]NN]
P7J?P\!42B$BW\XB#RBGR\?:6;6)OP>/WE)^-- NGE6(WEMQ0SEK7<Z^D?, HJS0,
P>O4U*]M!+P _* A/(.T$%,.R;]7_^72A$_&V=?B[!(SD/HM(H\Q?.<V?VBB/5OCP
P692.YB,>].@%!;"KG6%M\CZ?N_CN+;'J(Y&PK%CR '#-:,'RWS :402!BSEU:]B'
PM6!ZL)\A.)(&^(;^"?IHF %5T5:.H9)V>^:NK>R%%0)/%]T55WK:V+NC-"$ZD0*J
P^5HDKGT4*YGKI0=K_NSA7'P:I VT_[\TP#2D9J08U;^Z9\U[86C'#DCM)#UK'2(W
P3/3$-%BX<:,H<[FR; -MR1E'Y_\'ZV A\7(.D#Q+IP,L("X: 8FZ>$J!Z#J<)??8
PNGWH^:]RAFGH8DD:9P0%<-E]"S^(:2%0L=&ZI P" C?X6C9)5 $<&;^IANNSP9FY
P=$D>R@O'8A9-EL3>^PH2WB:I*=N?]BEA8:4,7$@9@!>XTG+1<(3[R+;I0]\IUA->
P%Y)+MX(]QI2RA#YO2M?6L6#^UR#5U_NBH'/S&XC<F-5\L-U"LG#;8[8G!N.^9=]H
P"^E<Z83FJ;>F.?=E.&UOGBR_C9:66FHP8V&[;_UT\.5*Y.4D2+X:,K %?%ZYT3F/
P*2O)@'WBC+QS-SL'@Q[J"=M3EVH10Z5;Z?(]Z.$_/6DC. )9%%FH'7U#(,R0SE@W
P?!8/L2WR5'\V)J'+=;V:CNP*1K1V_"!S0)<GE#LH#&C!: &!8J_B)QU<QF@X.<C(
PO;2_AUJ62:,-%I@1^#Y]1:J8]&_PHC+]-M*S;R7&_+\II$[>-QG(Y?  >,0\V=E1
P4(. 01L.XP+]7O$$^CH/XKN\R(1;!'K\7@#^2NM[4\%;[/<AW>FA&*QI$OW;W?@D
PTK<J/L @3CM4#L%TH%8C'%I<I/K8YOC7<SQ@)I(\/8C26_H< 8YA-",TA!<>_#/3
PQHBL]SYDA('LN*X]C-^!%_T5D"W&O[&+N:IL?_RSU"O>O!2<"]M<NR^UX=B6GR;T
P!H"['L]A+#P?*THI]5OX$:SE2 =>R[SQ#O;9L7ZL[).M>K=UQ?N87TTEF/>/[SR7
P!WEK0A:+WI7,R8M/]]::H2JF("ZNU3UX4GWL<@NP&2QQT%/M2E]6%CTD1)G/FC2P
P1HON;V[$!Y;/P[9V:FVJ35*\#2XMJ?:N6?8P$S!W^.>NHRI$W6?M&]O7PNU@>T@D
PY,36NI"-QU3].R"VBEGN4B('MD/",!]\POQ-_VP:DN*R<RPI'DI6Z^#"*C*ZC7:A
P94G*X,B1QL,#(ESHMZHR!'B "4M%9JB37P3!T<;?4;&T\M!-<;X6I<CNR:9B'XL6
PZY^E63#NQP%.F52E3]JJ\5 OZ>\1^001/+-37O.TAQ;YS'HS>_:KT:QKW86QZYC_
P$O2/J'C-Q6A%^BET5,]6V\Z#=KI,C #X#>GI)I*7>%F@C70RD,UQPLOO7^2H#<Y$
P7<0DFZ9%-HJS#:>O?4*^DP;JEBRUGK^;7:JWP,I^J36 )CKU: 4^R,RJV=4QX8&C
PJQ2\V8]FZ\;!WF09C#NZE*'LG3P"80:]2,6_T#PR425\X9KAFP;FBI90]?FQ!QHT
PRFM\2CL7V::Q.P:I0Z=[NIY>3#0^5UV47E.N&CLX$(KDH#X/40MBB7]I%0)RR9MT
PH&N!L3/&GK!H/AF \TD/<CO+R&%;+H$R1OV] "8W"-N,1GZ4M)D*S S5D%G/"@1L
PD(7WWF+L)ADRPZ?A(H3D-HH^Y[1+'0"\MQ6N)^O3"&K%BX-M/,0MF!DO$GA]O,H@
P,MM]?XOX ;+J3!G.TC$]5&=\'%QW&5;TB<0:IXI"_V S9%4R$5R1$=WR7V,FKC!=
P;+QGK;6$_.D)3_N)#I2.X1G]K]]H3QH*LQ:Q @'F JE/?*>K?OQ:<+EY!&+=:V/K
P VVE4*C1,;)9*)<J!IP>P)XCB0_T:55=HWP.CE7Q=;+LNAA4&0?D!RSV5/XF= &_
P5N'ILS#B;%05!Y9!L/RU5B,B\9N]GT0/)HX-^+'!*9DA@CRYZ(U]T8$C$1*WLZP5
PEW#]M"?,XY==UA6_8G^L[: H>!$8(F)L ^<S5I'I;+'\=LGNAL7MOK)40/2,NMXB
P ;>I<\PHYX%.Y%/(3]VIJ&VC5#ZIC9Q,;:JV@?@\W%>V"G"N*D58AVQ.N7PNV@QL
P?>MJ10RD$^.*X^4C3_ZK"V-E*/F2ZK#E(\#D2X1J4E3AV.FL6VT'0BJNGC^/*7B]
P[)PYL=,1\"$:1 B'N^W>ILO?M,49@682CW*.5&M;]Q#4$)<K>X<GX<8^:R!]#<LK
PS5/S5AT9#WKM!(^K8_,[G4TD;W@FD4+B'&;;/[MW9$@6=W<^=+$-TP8KV,,LZ3QR
PZR4R96B=$2*3A+[>#P0@\+R^4,\:C\'TX(0H/1VK_-KG,O4I4D6=A'WC2AWZ'-IB
P0'8!MC&%P<%SZR9:VN)OM9^MR?EVGZ), L67&=MT#ABL"Y&T&7)A\NU=G_EV_Z6F
P(1[DC 4/S\!2J*I68(.[8O" 76T*N^D\I+#C*X;Q3BG^<+3;Q$: C@4-Q>QX2(]1
P;=EUO>Z_[$<\/WDXAPG?63*H:,&\'"W=Q-JKIJ*N$U\<S3O@<;YHQ@4$6BOF6U,V
P^YO3!+U!5*9.]D)R/.+W'915ILFKM!KLQ33MHP1O[.N^7,I)G$AMR1FGP#=(^J"6
PQPTA%L# IAPU6KV) -!EXU*Z49!QN,3G1?D$NF[O_MB"Q90IS(^C_!(6V84:W]/-
P="5:J=ERUENIK0YBI/4_.Q2>7[>U!:8!0B[QJM'D;"H*--UI*2=;)**'['IV%!'Q
P8$@6N?Y/W-^JL'2)4+>8XSK\!OFU3[^Z V)9U"Q"CG<(3<ZNJ&F\(<6A_,K!2'?X
PZ\_8M$4GK=V+PD25JO3#X07]S;\R,D;$LPH%C E$1&2>95RV@AZ-%^S+"3LM*Q!E
P3&%?/_&VJP5LG?8D>8 8XT*>.3<__%?>"H"S-;>/[9!-WPL$[M7@;7I/LG1MN)L 
P5*7$"&W3DA5(!VY?]?M8I0E\Y-T3(F3]BA_ZJT)][;(Z*%61'SUK-).9<5<D39]+
P\TD2O8);;]04/;DDVO>O\:645<EOEGA_\Y0?DNC5+7UM0AAO@ZTY-,-QI7!:$YRU
PMN3-S[RXJJH8B'[B-E+*ITBR'QZ9Q]GF8@GOX=7A\?3T@-QZA:V1!6F>,0?.JO,-
PM&!9#\#"5^ZQN!W6X\*=CZ#/=*/+T@B.E%H$JGS3C#S.3Y!VY>29+JK[8OG=9'F7
P4*D(3/&=X?'6W!LQ-J?"([0*8._DEIL/*L,\ZI8Y0W9,-;+ZU;?XQ1U?N6@B+:W)
P 2FT/!7QZK5%J8AB/=[:1!#MHD3N.21D(R1VB+6.WB;V_>D$.M@RO:K6RJ0Q6%MS
PC8"CZ9"4R5Q<>/Z8%DK^K_#/K=#HATKXOA.TS65JA.GPD^X,!AWBP-JT)K@%H4CK
PO 5[(Z(;W>_"MD47P*Q8AJL$+=Y16K4%-V%LEX?2"^7[@8+5;XU6%\U_F7B%NQ*8
PCS));V1UPM$<H:)I/E'T<.2ZTW:[%?Z1UP3.JR?8<NZ&2I#O#Q;*;5RTTV*G#T?I
P/_1Q\24;J/J^%4K6!7,AZ)J&N(#K/9I3%3%K<@(FER<5^B)KW\/^U;&2?X[2KC4C
P0[?H]5_TRE8\'@+<:1TVD4S.24$D.NCU&?6:F9=%TRQA],@9E2(:ZM!&]E@(G$"-
PN+2.WJIODX#TW?$+,CEFM-=@3W$E#-O1,6_TJ53_N(<M@#SF<S&TZ[M%0/-"7701
P3XH+!@U*2@_L?V=QENZ;5=U8!YMJ#5R<IOEV]N_ZX_69ZN'S"D%=T5!&HC>-\D=/
P^9C_;9D"&_CRBY7&!#C?T^#(&G/>)G2AO3T]U<#6P820_]DJ6T,T5;1T2_1[I+O0
P'M.3$;438\C8#;8O<BC22-O.K%FDWHIBN/.'\^I&@WWX6RJ2S)T,!"?BARWVWUHJ
PSX4.E0F55S,9@IV1EU-%&PN>Q6 =GH4W5@;YD8%['ER"@QL<ZL_PYG5+_-2MN@(?
PFQV+- 1K_4(*6,&'<\A4-^-?&R&24ZH:=#Q8L3FX.T'JSY;HK[EPT=J4X\,3T_1L
PC1U-S-[$GTPT5])<\5M^H6.62"].0+P=?=$K2="W'4LS]FC3)OOZH.Z$JL"0#8=]
PD0:G$1TVP YEK&!#1_O&BG3'LYUQFZ-1;812X?[=]#_IQ8.>46Z[L=-1_ZU(]!%6
PR#@N:L\OJBO^JG[_=J\2H!]%'!-;=/]HCD >_[_CK].2BZ),1][M1CAG'3$+[^_$
PTP86*@77!7-;?$;7.-E]:/.=**T-Y1T,%]LFY'"8O ;C$@<@QC/7KFXF 1%EH53M
P0O<0,_/PBC ^:MGT/'_&4T(4^]4YLK9^#,F =>!WXO]Z+.6G*(/ PYY.-!VWI%%O
PC4UV$?")I*PJNRY]G:3HG,,I="NSSOY4<M"K.&"7EB.@</-,V.5R0:5&AY@IT1HM
P$6>;*23+@ZLBPT8P%"[=P#47H8S%M7?!/X440*@++!(IJNW)X%WC7L)K1\@Y2U55
PWZ7L%'RW382*W]]_@-.5V?XE=>T9(Z!LEYVZ;5*C?RLH<=].'N _?P1AGSE]V-7B
P4JB*()?9[761:'8ASY?%!5=(''\*VG*4<S\.C%)\IF5)@<*AZO]U5>GZE'L3D-@G
P2/O[-,%!Z^?7JJ%N("1A-LJ/=3RF\[U:\:VRG2A<>QNK>'5?61%M)S%85T=X1TDB
P4%<W](PM<3:7ZBV!OE6-,B8^F(KJ2A[+N_5?*TI)W%CL:!#-[V6Q 4\*F:+9:Y-Y
P4]W7.(6\+&7+;NFB=YN(R230I*:YT$_SK)+<AI';^BKXO59)=#ZV<8R"CH8R'8('
PQZ<7DKLUFP>U#865!Z66:E6Y/<HFR_-%27*[4-5YG(W-'&MF3"!7P,A]L%O>+SRO
P;(]*BR>4IK 9\&'&+Z0XA'IF-:0A/^)\&[AQTOBE/PIRA#LI0DU1/O"C>78+AC^H
P/K@32-@#NGD'B3^5%E)OZ!&[_Q?+KZ*YOFIUT-Y^=[E-8P@=">N'1M?*3+R6\%>3
P:Z@?YY/T0]E:W'5X\>=11!'Z5##5I=.-EJ.@)8-"*OB @;6+,&XLQ-!@H?X)(U:R
P>%%O;R=15]US &.]S%?PTA&5L8Z(EDS'@'!J*Z44^M:#'%2"*>4V;2;1?"Z$FH6G
P8$?ZU,9/Y+._4=Y8:OXI3P\$_^I20I+E)'#18#L,O_,8^%E_)E3V6&'D\>ZZ?>?L
P>F_&/MUDH@R2G@[5<L@1(+R6NWD<QUCN_(8N28O9M%]2J-3FH#LA&9\V^-NV[?"$
PR!2<N2%?#@[X"P]13)0[\W)3NGB^=SC.#8(U\"2D:9!.ZI/][7IIQH'2FM?1!M/)
PIO/.S SG_]/B,(G%[<):(YE=<N%*$%BDTO]M)C\TAU7>."2%S/@%CDVHB>.KQ;L5
P.)*1QNCTBLE)J)MD.2Y8/1%516/[LX6A,DO>:/%&E+7Z4/[%9"&"ZES]HJBYNF>@
PJ+;@WAMFIY>X_F"+A!R:?M'BJL28:W:A8*M5$7SV$ (S4?=(6/A M1-8+\]D.FG_
P--I$N5*15,B.W;)+SL;$1N@ 4!OKZ5ZIMK52^D40[=GU)1T)=?4:;X+TYK82R T-
P@:Q*;5C+SJ\%SDW?#I#]N ,5B7VG=:IMT R#7V1M7V8*6LA^#=A/@$RV?14<)A9*
PT$V"TJ>_9_,I7]\/D(:H^D(24520I(?=OCDM@Y6GX.1Q3 5I)S$3/AQV!FP?O>L$
P0=,B>]9/4R0X_8T7C?XZ/I&_$5S:%9AQZN2OBS;?8MW2.3^&8&,6)$L#Z#B E3\K
P< :MZ/8Z5'%U@R8'EQ[S$WD:75W-DVUHT4O:9>6_<)J(!MG$0RV5ZYRD*GR?RF_A
P#1(8GW5;@>84AE[ES[N2:1,0E;%<Q[$R.Y3'FFO,:);6H=&UPUP2N^,=<)>11/&R
P<:*>%CU0A=9W.]EJ:V!Q-<#=U"41W_$:=B8/Y,<+4;ZLGI/^QJT]H"1VJ6H'LC>I
PX$OPWVRT"Z^1_[)[8/V)GHK>?D_%0#!$PS#JS?M$?>5IJXIXVH"Q0C-!2J=65^E\
PF12!OVBD2CYD/[E#CP<*Y'VA6'9!7U]R5:*%@G/D5)@MNS+B;Q2JV19PA.#0VF$3
P4?QUZZB)X,P*'DMF\F6O[CW)LRR:2@PS(Q]W>EE:L[:RQZJ0MH1'$JC3!M(&@=L-
PAUHY#>1<^(72GV6D_#& Q,/]&N:BG&\^\7)5RA\%8?!CBU^BV5)")$1V*S)/FJB.
P-(3C_8O6>D9/NQ<I=P5I!;R@WY&99OZOQS?@>-D>>3.H<0AR(6-:"<_MQQZ((OQW
P9_Z_4Y<LVP;=W4?"9)C<BQ54FDK^^6;#KZ4L9]!E\KT>6V+ZM>(TS05'GEE4YK6M
P_P98<A[;15#RFU(T< I9]E0T3<+C37D1S*;^\,Z9,4V-MT?9[QVL:R.:8BSW_:=0
PU4CBG9 GMU7[CBDBZ3[5*2^3@'8M-+T-H/FAPA5)D1P;-<E[+*+HY>M8?*>N),Y\
PP@D.W34XZ&&'AV^@VX[9KJ1^NRQX6 #,/.(B]OB5_8,X93R2(KIVXQVR)NK.6/#E
PFU=WMN@C:Y>J80536UA.A:4UOI9CTE_;=_A%2DG=:4_((A]!84C_Q&_LFB!!ALG2
PF*=O?-\TE5A-VW%R3 H55D@[:^B4Y6R@;N_PD"U8*8_+&/OZV=(CD:E1\4H;(5>Y
PS"/F]/):NCWGX**+3[_]\^*3,1&4*5A"=.B41!R<#=SL^3.(]2[VXF#/9^[>0D3)
P=VQXMY]/^!T_Z9RV.=RC5.?54N+X"V7 Q<":Q2A5NE..2XHY(7;YK_#/-GX5!.DO
PMM[D&$CB^'][.\W:G *4$7SOA(RT%*A32FAV0UO2<ND< V(\R[&_0$S$;GFKZVH"
POAUK&M1M=*YG\Y6NN. 2? 6=!&%V&>443OQZ</2^ITR7"=W!\VZ_82(:^4.LZ[;5
P*BH+I(D0B!T"'YQUB*8%PLZT#D[GH@?0&9&R"^1EO"I#.)1?U%?K>.X%1L//+VZ]
P>87R2BIL5#%YB1OI%@OFFH@DC^C/)8Z?"ED"P:_#F6'>SM=:B3SCHAIMJ&UQBVU:
P+>B+S:\W1!O3SACJ>];61$!S/= )/R_$)59-4JQ&XUX]CZMG4?<NC.^<I1S][^)9
P0.Z,C(SHM)!;:M<KMC'SS +=2&\O R!V)C(%Q=@30!!^C2^2F-R6M-R,E93E OQ4
P+<R6U(J@\%6>DF5:UUBRQ^,DER7\<@J^3&:\@K;+>F)SM3 @"TQ.B'FC]F.9[U]7
POQ$0>#T6081R*=HC]49M0]-<>DUKG*5&?$VU?] APZNJ0$S+_%4-M:<QO8G1N[SS
P?<M19[LPY$RK  \MC(HH>SZ5CQRK%1,-7!5-H0T0T#4?I_JTNR0)S^=W/0B]G2!<
PG/S!.CF96IIO&!&#0^T9GS1T+!RA5GA9?=^XAOD' S(3LFF$-Z#'8Y7<EO Y52?:
PK;:\4[89%E5O$6;AP+FGFTE?6E.%?I@<&]*(=G@[F?"W4Y8P"@X67#?*7=>O^$6)
PNP48B'&C45[X6I+N@ROR\*?>[2!Q?8]K4IY8PS4U*Q]G'/-E\ @A1N6&J\40C\&T
PZPJE_LUJB95@G+$M^IEC6@ND9=Q NTQ%\ISZ5/:[4>1MR;QM>TOO.Z;=E(H*H,V/
P7*$M@6FRZ D\)LXP<$"8YP][2D7 :]N?+I(=^.W2O(.=7%CSE%))1'9[/5"S(H?"
P4SSO4&>V7 04>' Z%0>IFCFM.U0B*],TRNN?I\"P&]\3+B GO CMYO!).QLF?"(*
P^V2JFB^Y+:K<@Q(#9>(8/NQMMUH2HUN2@Q87\O?F<23A)W,)@6:'8T$S[U=',7N^
PLO"T5A>&0Q:\?#X10F*-]-I'W5[ E%3^7U3:NQ&61PET9W)U'^#1@LY)LLPKR3DN
PQ/#L,@BX_5Y<*/F^G8:+0*'OI_54)1780C4VI#Z36[7V ?>\Z] -Q;Z@=(BC'9_@
P<_A"G]7_KO0Z-;1+[3IK4YY)HH1PZ6KL_3A_4 B5Q]_@K_W@+OG[/UJ)\-7)"G+R
P]3[9 SF(D0]&:IIK>#A-*<;89MSA.S&Q6-[ 8D B#V/&2-B"<PX+\TJ04EDU:4.<
PR:'."HQV @7T.QKV"_0)HT;1$ $W%NDO,1&B,(^DEM<U U;V\V[=9,L-%_OEAEH*
P9X[8>;>E@EEQF_04 V5US>;L.9$U;LVS'ZY.!^<JX;"0ZZ1DKF6(L,"GYPWIS4"7
P0M\=I>-W/#'H?MFEYK:A0C+G18C38%$L9)L2X^R+M >NI:?5WW,GSQ8)7FL(8GP2
P2-:CB5O6FL2%*.VNC;K$#$MNZ:56D$^#T,NR&%]FU5\6=C-=OI$- ?'6"';X8V<U
P2O,6#;P>->;#C"%_OF+Z@R*B)/TV,](K8DAAZ< X4._FO1I$D[&-?5=(QZZRVSU/
PV3\1S#Y2Y3\^G:@@)K'5!CXC"6!&""+?D10W,+0@?3^Q4H@<LD:4.278%@5>.ZV5
PXBP_93M+]RXZ=(3"-HW A4E:U^PB%>DKC "&,IG,LM:*X@4B:DW$- !)+GQ..SJI
P@<M2-_A>P2&J*T:M.2_!E.)%^-Z341)16Z^40WC#(DFS>ZI4AO]E6>3+FS+R1-1G
P3?=2W)%W4L&M  $9/DEGL9.56*-[D(TK? _B%A)UPH6ATJ$/5O9Z@8L(.ZB-U^9*
PW\7EH%I(D9&2G,[K#!CE[.'QD=6J42Z)2$B]O\(KH%QII+>T7M1HDQX]BE(F4!D%
PQ6X20U,[Q);WMST%AE2X&R*KY,R\;%S5Z"M]O(<'IG7]1*Q["+:UXD9,LX[H"''S
P/HXPBQ%#\]N4+A_%609TV<ZR(U7SBA1PH?[E/X:KV'2,"*N1X]!1.42X6\I#UIW7
PG7UFN3LNQ&D\%77)/IHYV:HOS?A='EO.W4JD0:,\9M47]'-*^9H+R5E"NKP(.L21
P(1'JK@W]11W:B7Y(<E)86(9^-?B60-*G;6 UZIY'(,>!?P8=V00IE,>1-,\EA!JP
P.W2=;V;>;.\#Z#'=H0*NT=$.ND$]*?E.[]\_VJ>$SH*X'JGH,;<'H.IW]VQ$4=N2
P CUKAR75['Z@%ARX3*$I!MI3-E!&;1="W#1J75@[*3[X2D';LQGT1W^%&NI%$33]
P8FTX"RB (?X=\B8$X1?H^.?778F Z8OU$<[E/7Q5ON(;7\^SOO7:&$('(W$P<,DR
P<,JC,]$$X1H=#1C/5JG 8'HUQ/VK%8$11P_,.'V([ZWF<4:]@TU&B!)Z R23OF5D
P."QC?@KQHQ<V;/C.& 0EQH5WU>*,,V:WJ4!^ZY/2 S?>:;-B%9NTW3TP**F_$++N
P3L;@<"O5;N_BSU-%035032<]-U1$6T?0BO_B\9>(WG(,WCSKB:G?8RL&Z->G;9')
P>F*<[GTE^7JK>E<!T-0DAH+^^:0$"&?NS?-\J!VU\[6"E$'I,1.%7R54\+U&7)IC
PM."E*7B_^-2+K=;4J--YKCE7];H?BNLEZ-@S7:J2^%]>(G".C&+GAD$.N7P3XB=L
P0-E?@*%^EZE)N<4D'A.UUUXGR:S.*-D7RDY^PEHDRBGG+TQWWF>3.<.3"?K2E&8H
PP>J\GI]E(B_L3QX'U0Q9(8//:<UP=NN34.1FV'6NH1[HMN+O0Z>!\%,\2L3K(*TN
P2!Z=*,A7"+%T5&*RLZ\2$_943,C=O[CE4%X ^P1TQQ<<8D7B(Q[T@\R\QF$#;QR"
PU9+'532?M9I;],<4@57D8FRO]D!G_]KAF2#)XH=-F>9M="A)^,>X,A Q2T+T!0_+
P9"M%\GIG;B.,"7.7QOX$_EM9%B0QH.^\]YM;6.,8>AG+$;JD<T'; K#)I!JN\D[9
P,_=1]S_K=7=KZ#XWP;.TMPK/MO=2#6U)_ [$^WWC;UH[QS:Y5+'%!PI_=UO#/""6
P4ND(:FCBS6TP+#J=\EZIV,M^ZZ%Y9["O73N6=OT;DYE352V!@YP/. RU/5NR\C]T
P0APYV_W/C!!/%2Y;"6WBX39%U7WAMZ6LZQT$#?K2#?Z3_4EP_$:P1]H%)8%*])CI
P\4G6=LWYH!WQF?&[GXL>[HK;F]XF(IE(.1Y0+5LC8?RR76#1.HR5[@9.3* 1Q5.!
P>@Z/^P.UP-]9<"N"XP&VD\7P0!GN:%K\ 2!E86P'?'T6.G%B(!-HKZ<R$9',5P/'
P6)JX)$.'8AB,-> W>]K[(@^Q/71G%GH7\0=,L\P47D.D;"I?9N($7CX8$[[8"[7P
P@PKM-P) <A5F65T\C9J<8H6-;%"L2)*]FH'D9$QF<*"LWGP<#*!^SU6(/O,[K OL
P4HF,5'S?>C'P*[&5_4B,8E! ?@=\*BRXW4BF+<ZV(9@R[5+_1>$>/F ;A.]<7],!
PK.-HM4^QWN8'(KN$!>.6 ;$U9-O@MY<"K#,4'4?"2SI"^K_[<?:X)DXR,<%545/?
PF1:T R&]<G "59J7U+Z<KCL51I,DE"#Y>4S$B3)3-$RN%7(-^]5^Q:IQ7,P!8]++
P'./%1IR@8=*0%OH_'2(KX2)11AIB($D#IP'N3WJ'=3V\)K]NJIHT',J9+#',P6[K
P8L,@'4W%[?D**;!D<O6@ =$_:GZE >?S+\/[$7,Z 91K8Y8OBR1!IK">L[8R$UH#
P@"&>2A('],0J/(F& :_+97-?;[=^>O@#F.Y\/T=[)RN<;;5/'(!PJJA&NLVXK%"V
PG9O3-P/P%,^4-1*-5&FS/#H\[VEYRP'9-$^E3;H@P $7?$!?BP?5[;!YU1)(TJ\Z
P_XY6.'E$M%UO&25V?6,'VTE]O!2?MJI+ZL*>+,IJ@7BF('K"7W OT1_DE(!(E0T!
P[UH73S5A>N48(+L><]A>2+-XJ1X8&AJD^F=O)PE^ZYMCY@MI;P/_\MW6[K9(4/. 
P$K ?/K>_A,!">J*6N\P9JTR@$3_2<X5.F]HUS"27(FEU*JVV)X<;OU2G\H>+-%ET
POF+!'#".?:Q4(72!0N]Y-C%3$FO/L?(/F?E>T"1R?&]EYZC3(P,EJS?(^P@OQ!W[
PIN$N%AOS?@/WX<HVF1,'1,_@(>;5?+>(N639?4JFP+DJ$<,J%,#4?9YL"3ECC?AB
P,A.1\,2J,U;)HZ.0_:5((%T .\M&RW67#6<HBE(B[Z5L]WD[=(':8V5A27BQ;!3Y
P_@(A&VO: S:!F#;_]C_TA:U$$L-C^&XL>C]"2Z!A$DHX D4Z=UO:8<75CDR@X!RO
PAQ%-OXH6B9995X.[P8EP8B \^9L5' *#]\%^>A//)/-!?^#;/FU9A/5)7A>[9![4
PI'%6::*/&X5_$F-DLO70EFR4-WY6T?,D::LNR6*\K.?565CY7YS<ZR&=5,=;4KK'
P_II+?'66!K<AS% 3/S]G==W&W)IU(SY4/%98CPIUR09Q03G +7M?>="][>F6 ]3J
P/9W[FVEZ0T3FGIC*6DZE"[#/;TIBP")V4'G((X0?>M^Y%4UUXYKA8'9[ME"[^X]H
P:N:.-.>^O7B<DP. Y%^U0M&.GU3R.-(#LD_#S7I-V%1D,(Y@184D,RL;@I6BV>1V
PEV06OP7EC0L;#U)W9EA1@@:PDB.612$HU- L#L7C$</U\AQ8#2U Q:%ZL\9L4+X%
PC:.#- ,S.">">$4:X4_=J3438;D@R%GLMFN,JS\+V302[LS&=L)4E^+ -?_9T7T\
P /;Y'UWN/[HZHN^)P>A[B.JM1[\EAH$,6J#9;.M%LP RJD>&D3^$/U/P#"$JI ON
P9J:EHSJ>;=YPEC+KJ!+[_\]3W\MK86.UI?2V6(RQO.>&J>HG5,&M^TH/FG4[@[3N
P:DP6R":A"Q\^- )!B5OP;4FJ*-<,!4DIL0X$L87]=<)>XB)6ECOPWWH0S;-?&HYQ
P.7M5-J4C*8\[1(6W\)>5P< A012AS:<JJY:)':#\_SS-0>==38;4:YVSPC"KJU-!
P;.@M6'/(APW_08>F8%FLDV=0UA/_D$]#^P=BWL8IIT]#WA8]"&4@<9==KH$Y?M_&
PD4^D_"=:^$)A>E^P[;D0.A,K*?0K3J"K86GK5R_%X/7'PZF%(\RX<Q/]2?'!"WK<
P084ST,N8)RT6DFBF$61FK*B%/,<%V$XSUX)?#&S\9".=>; J"?H4>2L=(:LKL79J
PCFZIYGZO_28#^(Y$;+R)1.1%3\..#*(6DLJ&=2+/LZ$1/ZXMH'^ZP[_,0Y3G,SW5
PH']*?9I/2A+,>.+D66+ZQ9M\3*1))\TE^^=W/@:L?0%WHUWPZIVP'_MP:!A[]MK5
PF%Q3.2F-/5R:9;8&Y;>8"Z9(WQ3,LGFM0<VFI>_]'QC^X]KUY[$+N2_D!3PG]+ML
P(JW0YJT&AC]>*^H9Z%=S$/HPCA9$5O93\?,YKF^NLEW+*P6#]Q[%^MS'ET58M:1P
P [?V/,GMEL0(J5UE#5ZESH_PSF<TC>#$HOZ\G/\F1=+"KF0J_0W4;M>[=)7N]M1&
PC4&+Q-:1"\%Q\![Q6D''6*YD>F.F_[U\LO6#F=S36JV2^B_WS[[O?NPQ^IXNNY!Z
P74=/*PDO8(XH)<U H)\D_PF3*4_*?"7]8Q<+O*P0WVSP=(W\JJM%0'0@=(RS=S.<
P:&D.J=3@\9#E ;PRA2KXAH@=,9E=DLG[5$+I&HCVZ<6A05DYAXA[K/\?_<OXA&M:
PQ_>H2P9*5R&R%DY)'FJVKCBGU+I32P]/!;\I[_E1[C-QLH%USBSD;6-C2 %9&3P_
P^U83JHS_8R.V5J-$7&>K [>'?<VCV-U.'#553%6M:,:=+6W+:UJ; ?O?X$0&RQZJ
PYT]O+6\FYX)V4;Q$:O.]QX#E<EIXN6:3$.Z\CD7]>U"X#X+36\QXA$7QK7T=>=_W
PP,[A6(03SV^]ODJJ*/:+7X,_()^E7%9)?!KE]X90=K<#UF4$^B44%6%N[+4@Q*.;
PL.M5XT21 O3VDZ-1 ]?@0Y36[44@3R&LE1K_A4^.=: "#W."'K=O8 !^":J1+; G
P-4Y\:6=IW&GGW?CZ"+UY0/<9A?DJYR3F'\?>.]]TP+,RMXX?CI#5BJPV!3$'U@0"
PRCZI)>4\%AQL&#:EUPR?4KTE*(_%&17 B,0I+I* ,VG'H\S2MH_ 6Y30.?9SWP/2
P@O7NW_-AA/[<H>5#_;+^U<Y14S(^!08G%YHY?JQ/-+M==G+26;IQQ4D=9-K5 P!)
P(SEUDWH4P3KLD_RJP4AQ!S5(K9&?\8E(1EK&N [[OB#^4<,.7\8WO=*$OWVVQF?8
P98-*U7'9#T>F\&4V90\R]\ =)!B(NU13T$,DF)HD?E$;3UR=+$C!.CGL0?92T%-V
P>]V] J,\\4]%VCSS):\K3LZ-X,@_BZ8J0/!^DS*N6O@74<; G/A,B<(2$",X\'VH
P@INLS,%N0+L7=<TZ<D$B $?,%;;=Z8?"G@%O6N/ZCD*@RZKN2E5!#>$DCJWH(PV(
P4$$\EM$B]YZMGDZ% EJ8RXLW1;VBIQ3:)SR$_GN1D$\P2'8C__,H>'EZ>6B!R/V:
P*FXD7'&76C$3X#=RI=3"YD!Y6>;/0=6I[1&>4V3F5 :O)WADD_!G\U(ADC2HGW,2
PTEO""R^^8N*<F$9$%QXB:2N.;DMN46_^#2&/'VE.;7@MLY.X'$-.Q 1TNFK/F=HW
PL+D3^&YK4EZ975/V*H\ ]X7W'(F&J6B'0I*2QEEF W6_VAZ9'9N&6G[-BNRQWY>!
P:WAL^>\"+KA%CWL!'.BT$[M8:&/;$)K<YN89(;_BH$+%T@D*:$R]IAC5,!'_M2<S
P*3L/E 36M&HRV_?'5W0< /XQ[SB7\/.XUNP>"2<9NQ<K1X32*F*(5]0T*"Q:M[QW
P^=N\O5N:!Y9-JBVL.#X$8W9)W:Z%UUBGR"UDU<.6TB<]B>_Y+Z!'&,=["\K]V=P0
PDV8\(5;D;//C,N0\"#!]O1A'6E]\/^2)(-7H>PG_OHQ=U,XF>&!+MQ.0D,1^BEM;
P;/#_JD%FI+,VVO&022$TS6H))CV^^ *N;I&8)?J5>E#X>Q!9/G^ ^=) <QZ&+V(@
P?E^H*)>\%7<8"=ZT67!P\Z[?1&.:.SE!DQ1"X\XU?UI6J&SME@?1/VG8ZB!;Y$2Q
PWV1[424=D$C:!QE)UN-)YW!!R=Q#'M5HD^="XK4S[QF&]/VG\<<VMZ&&O2CI6&,;
PJ%QJ9<1^W*$LG)8U1YAVCTJ\@4[2<^KY%^ .)Q]0I9>;J^0&IUV;D?<0JV*CHD\2
P.-GV29%4"]%8H5 $1B[VT1P]#3V4<?!QXSQ7=Q+,=!EOV?]S8,U9+WT@=,,6/$NW
PI,R]-P!!1?_6O0JZIX>[ZSTFM%019PJB/;SYLT-O9?C"8@=ADUTU:D/&^&=I,;H#
P+ESQUL,7/ZMY>2C-C[&R4S+Q,%G$=;/ZZTKE#3I6W@R!+ E+DSCS)0D.N,:/,EZ2
PE["X;;_\6'-R_9=96X)#_W0/PB[+&C_@&0(-G',=9NV:6[Z[L>ZI_RM+DUM"]TT:
PI+>CUBID!&(PS2 4BL3*$GRBZJ:Z[<@8;8_*S_9 FD/ND^T%-._K1S!5]%'0%W^N
P^MCUL3K&)D@\7^7(7A0"$!E96DA:J\S!-^C3)1BG(R_.[.?<;'Q_I$_4?12;H7'Z
P(9A/1\;=8E&_Z:)^?G.>\V86P=RRQ +/Z4<1<'0^B*NV82=M4SON=:5DH\AQ[_20
PG,51J&6!NR>SB4\/=(DW ZGH>(GO_I#N7^\93H6^X& I>.;#Z*E@;SA[R?8O-$' 
P[/>7".O4R^4P,ODL%ZV+'CXTS="JH#NC_\];A*R7.TQNRJ/'8V !IC'94"^FZ?J3
P=V\A_8><I3X+0--U.1Z,,]Z1T2(5K.LQU4MNMZ'A_JMOP_/C#OP?<%_MA&99UT'+
P<]Y<&UU3\0!I6:RHY48A^%QE3>8Z=CF3<]38Z?Q7[R[G=- >WU.H@$WK^%;J-PH>
P9(RI.CJE_N?\-L\V\A.X^T\3PWA=TQ^UX[;0\,+"C56\R4!K7.Q*3?)!*,*NGFR@
PM?_'+C;[<#:>.<#_"_Q'#7FUS7O='Z=G=,#8!?S9J],'.J";U"T.)C+C7<P1JKA5
PY%N^5OLX5SGRD@*5*E(*.M6*/]ZU+0/I=R*-';L )H"QMS2)T83#3G$7<3&:_RD<
P4$@\SV@SBJKOJ&UJE!A[_MO_S4J,CW5S.!DM%[D4Y_JJ,X\HX=BCES+?;2YKLSY0
PWL)'Y>>0,+0!**([+B'X$IV(,541#ZT,,)?,/CB>3-G2PY1BT4+2RQ:B\9-8SF\O
PX!>>)B<+.FBO;%IZZ>V0&[]O]12)M&+0V@U,UQR[F\E8Y'"=7!BH*?3YT]ZD"TNA
PN'R; *KB!+NT<S>3YY\W_L8D?H"YZ@!]T[VAM[>"5'$B^@,!KF2@7=MA8$/X-"66
P-:N;X+\RUQJ:LG5BD#X)M>W?)WIM0JK8MKU""#YRH%W%]GA()?V5[9D8<-3PC<\W
P8986_N7# I)(C]O,7SK'=CH%-["DBCOG?P% 6OS8Q*1MZ.W5#L5+X*M 4RJ\7\:N
P5<R2].C3QG-R/$E$8NE'0#(R$N<]4'!L4FP%M-X1%<_1F>9(#X-.[%K &5K\#E/6
PN0+<FZ/%^"J?LGSQL?R'NL#$$-5J%S,<LAJQQ[(\KL\H:36.VMUN!.(/-WD] W/S
P^#1:,$ F.8?_W2ZC]2>Q6K.7?RR!0![>8KA10U*5=FLE8 DI-*#3ZPE&TY.>$#HX
P+E'_J@RAQVS-[9_)I4?3>=/.<ZDP;J2E:RZ2%$8.>[3 IO!OXCAX7O?"LRIO""!R
PUO0-,T)WS@T6LLL.IOUQQ-IR?>UKCB6JTLT-$9&U^VCQ3:=VC4]LGDOM2#;LF91T
P"9F1DM!^X?%_EGUE_7;,F/G^44%(6=8Z^7I(2*6-RZ_1Z&M=1O4H8%^K#K1/:-#&
PAQDS#)Y9)1M%M7"P1REFZYJ3NE1+B;LJE/NE"@3LS.QDP.PR$_>L7)8Z]=BAIZ2"
P?3-=N-JQ.5S24L;$A*^.]4X.-:)(/43]X41"OGM;A'/GY7&/7;1[;HC/$"7C<5<4
PEC0X!FGS6:+2V.R&)KE0@%]^S]G<RV\3]<TCG#>C3=I6Y;H<14@.E*.C4T4;0Q/H
PO6NV,WCJZ)E6XO0!KXD# Y'(YG8VA+N26)E_B04N%52I/CABD^B7'2^HHN#,T*XD
P*/\;]AAZ)@^=]6< /KEZ)HWL/\5N)""991JQSABP_]DP:=@'P<!VG-&:\4/P253?
P*$?K: R2HV&AH/WQT%1_$XR.N@,.2OR)4YTLH<=YNW;0">76% 01/5@;0TX,4>*M
P5EYQKU.Q'VY<K>:RK(--8'3QWLX9 0((!U(=D)T?#W58V]$M=BF6B5/RWHB]W/0C
P.Z[AH7&;Z(:),"W)!&PNZS62AKRO0&(S*SIZUJ)G!;$P\\S"SK*CJ-;<;X+J'9GY
P[(-^ZL.3BO\-\#I@H- GIQ'6(N:N)\Z;39V'3>".E4FX8TQSK-03(C?AJ)!K.C[!
P<HH![!L+?NHOP^ TA#(G)YDXGS#;MDCX ZMF7_]1!M*E8SQ?X+E9<#3N/@QA3)H&
PF"0AZJ=5!FA.3"1N.DZ/(@:=X3Q#2A(8LW4H 6BKA73G@O9U D0[2_SW<4<R$*AJ
PK6YI+U+<MPB(/)(%2]A[$0_/L ,UE$M/B9]'=?JD;91L3J1U<;LKZ^VI$*X+&K22
PQ0@9(XPHA$V7/CDCH]P O#G/V0+\U0=K@V+&1?"Z6AD7!V)SNL7G_T=31TSRR8-B
P:@-PKB% @,(M:!9FQ^:RN&+!:@$8NI=C2;$UUA%2NB+)D&@97&QE2\/7CVXQ6XL]
P;DH/* D'("RF9!=9I 8O:JKEL6CDXJ\A\)UIP@[NB."_XC(Y#^>&6%X9+I]:7<#-
P # @ 3O^-BFZ6<O:U+#3CU_'7+]I[>U^+^'E"(XGX7S/<(#*%+/NZ6O)=4#GYV[+
P9OUV,:FHE2L1*L4\(_@OS;@A?"=/2/;?YF$\]6"E$?VPPKP2U+@X?)855,3(UHI?
P"NT$4T3H6>^4LH^VD.XG@QT3X-PYC) ;!P2T4O1&HQ]4]G#61<\'TC>C8@O[A^_Q
P"1,67 71A5JUFKA,L<'FA&^C?Z1EDA#8(%L/DN!AVPQIBDA.)I7@@#&N8C?X T4Q
PM8>?S2']J?Q["ZONS$[YP$T>X#/09J"8?'A".Z]N POAD%JQYA3/X4U5(=6?1-7L
P@%"L=%.B_BYL%1M1#=&<K['[V6"[VS4P><:,QM]$+1W\C_G,EXGV':>7BK $!LQN
P'&(>A=QRL"&6R+"'I-^N"P=J%JL8!Q5ZW_6X@JRX]6N+O4K'"4#)&4K)JGQ-RV]'
P6<UN;>N)I^4KS8\.N/EH$CJ-=CK%E]_]K^J@\R\#.BM3AMH#Y)B#]>.J$1_VT8V#
PH+LP'URVOMN7Y#AA=[#V=*50(@J5?%NTHSP8-(2=P82&T#]]"&#'GW Y^>6K0PKT
PES';\1%ST*FRF&QH4K-(0(HK"3T?E*5^MRQHCQ\*U)M-/O^VH^O(O97PY,/U!3'+
P.D;7'P@4LE@Y# LZ?T4*52*B?%E*QXQ7IYZ][H*6YA=1&+4*2E?F9GE+_;!X-.4[
PS] 5W6]HS?(A485$K?B,+:O7>-RT%OG.J+IQ7CS+Y:,*O2/-NSF&FV@\_><!VHK(
PT.IIH?NU:$\UW4<^6%.JB$GQ:-T._G08[\+MN*^JZ7P4=59BGO&M@=B8?1LD:L4K
PYCL!-2Y8!>:W!UB9H"H\/2*$+4UE?_[E!7)/M/0ZK A3!05(B=>HMPZ]WB&VC;M:
P QJC4;XHM\&;$PVYV]#=9Q@";0RU6+W;DCS_\3("<TX%VS?1G( D?05 UC;JX!/N
PVI=-YNH,E>$#14"IELF.:;V4=BX^ N+1=.,+L4WYMS:"T"1CF8.73\-KA[HH"]+F
P5R3ZD$%W]$4.P;4>)Y3!(JT'(BR[N&+*:^7 C?E>[U8[U<RD&:3>BAN)(X_ML[-T
PF$GF BIU<]PME@LA&&:W\\QT;X_Y9P=P1AXC\M9^:^>7$*UP5-*,KVJ]9SJL5>(U
P-,PYWRL>K^/,7_:3;37YF3SR<,P(>+=W26Y"JBBGO3R?FI$W0O2%JU5O7I8@I!?$
PQAQRR45_Y1E5S?8G0J%KB>"B$NZ#.5"L+M,UA9[:FLO9,<P4D?$[BV5$@Z4?\1[L
P.T/=W/;E^DW';E@V1\U8=96K!]2D<7\HD@58,VN2;*G_+,9@QGO\I^.\.BX1PNRE
PV@7@-JO')/7)HI=JJ4,4QFQ>!CU7F":3O[7,^*O\]=[83@RR5NC^Y<15&WLQ:E_N
P7*I'D/S!N!?_ N&]/5<?I&S]C/I+&$G34H3!&AAX$"DQ4OY(UQ/2A +7*:[&6@! 
P(UY_:7J:\,NF#ZX+ZWAIZP,[O2818=78XR2-J7%/1[-WM"=*[S?F)$NNG_^#IGB[
P1<!#4;:;<J4#+>C!5Q,%C,5=X2M)C1!@)P".) (6V":/3'O[>MZ<RS;F"&;:KH4#
P_9G#L(M?L&.(<-#G^2D^T&:X!>,#H!O%^T[9Y#D-<))RA[TR/3XD?!N>HU"G([1)
P5R!9 5):*;SC0:T!.ZL8Y])11.GS])%GP/PU_5EICD44B6H2:U_N_AU J&[W%!("
P3T;=E!WM=A60GS%T_$]4 \:S^DW1'2^24UL_ EI/_':5K(9LR* 'ZT#!PELS!XU&
PC"F8;_FQJ920:8GXF1@_%%88H]P+AE''@O#_3);L)+'/:,OWG[075I/IVZ&Z'F#H
PN$TL W8>= J T)9#]VY%]-%:?D=B\>'5\\QC-G3S&'BEE7*2G0Z)IQA<%&(#O598
P]VC1]WQ[C@CME+PLJCW_G4S3W$G"?80,X7*O6=SX-@@E]A'7$X\A^G>&$S64"EMZ
P^3L<0<D];-_/P<#MF^\#&<20&PYQ"UF-KHJ/(57Z\/=O,"^*=$-3)LI=M?8\6W\J
P($Q.)C/NL2T[TIHT&,;^.?H,]U84AB>=U$GX]-I([.H"GL@L>!^;)V0Z_!S+/NMQ
PFC)%RM,L_,/7WO)&^SZ0)59GQJ*"\V'VHI;9$JF:L!5:AGJXV4T%/K1=41/^ ZN%
PAV/0QV/IP$2/[>Z9AUCJX\Y?(J:<'JZ)G730G4_='SI2K+N^VUC\_^)\6362WH.*
PDYF0 N8[),8P#D]K6>4+:F*#VWDD[%L9:!R4C^YZK?Q,K51?;)6?/X&U5VKT_L E
P^4PS&=73^ECXNJO<;NM Z@]E+#/K];^&DZ93HT E-%)I?UOB2K3LT2;ZR7]&3WXB
PZ1+D""V%(%$=QA[4D,7=>$RL)U#N\7 !\S6[?-PM')XT 3,K$57_1>1,-%^J)+3Y
P+/_RM1M@>7'M^OF!H!ZNU3R"1(253/Q62M@*+5G%:!. 'SB7>/20/S%D*,S92H;X
PREE7P-!EJ7:4I KKQN7'<"EO/7%) S-[2!0;\KZ-%4"G*;&<3LK;<?/A"&8(0V6;
P#6;W&[DLN#?@ P#4;Q$L7<SEINRZ<1%MTFPN5 WPHH))/A61O"8VQ2=6I=CK)"XL
PIK-,TF,<)5=H#"(-I/')8.SSKUXH [ [XF0@P#S$,X+[@?LID?HGML R)U:\0'#6
P.6_!+9N3>P0_>H@!O[G@(=U*<#=5;;N2Z H<_'1: _I/PZ;G=+N?$QKQ(;YM]<NL
P^^1$$%RZF ZFV'-7J_ 9#O>.E2:!QE$6K9%M<6JMU2(*^?#9?0E'YC/[.O\Y&>*H
PJADK)6LV[[E-K I6JD'BUQHJAHMAMIHD:X:[-FU[K#7QTRSDI\OM>O+O,#^CE;@W
PB$JA9SB"U.6\^1[+Y?)PB9&6BR<SLW6Q6YGU&^\V_?W#(,P<1P9'N%E&O2DWZ2?6
P''U.RVZB"I)?$D'<K1K=Q__:]K"1:A@@1IB?_DQ_JN[Y-B!NV6U+\UI1I2EYV$)6
P':)W*\ KR8-Y76=8-@8DFNG\>;]&8W<35BON0G;PAG!WEO<!6+=$+"4B>P9SO8D5
P:JLPNL!1_L3UAC*P0\S90)'X6\H=Y AHK5.8L@TE/9]06B'5>S5)J#?D2"P?\541
PT-NRWC<9(\M,^!*,,.QWWF9G+!9S-5JN_8G5?U4-;\9/^2&5L<,(P*RH(Q*J3,U=
P1: 0YP*^F3V]G63;MZ>]8 DMU/:;U[P%& ].XQ5RBO?N,98EJ"C&3Q)L;!LR"22^
PZV D3O6.QNU^HDE8G&(-+"#K5V6?O$$1MR0IS%B:^$8TP-7AP9,S"^B^.-H3H1\.
PU.@NLM".;X6-OZKI_F,M.@+7R$2V]0V"(.">D9FU :,^N!6_I/..AIO#\O!&9/*6
P]RXT<>0F%E.&N0 ,S($K(9%=$ZW1DPSDXH?N1# _[3SI#GW:L-0)>VVYXF @$(IB
P*T.MON&#Z]1S[<+,"8X6@T)-$9+S\(Y4C46Y94F%_$A&Q_:@(7?Y73%^UO+VOS&O
P 0AN_#'2>QB$'O5>7^OO.G%',F/[U=!J_F4;3=KE_5"Q\0QQBTC]ECV+NLE00X4U
P"',L>(C.Z+%'G>CXQ5E;SM0>U6R!U_TK(VD9>43!J(: 7V-/_]LZTH"/2?>A>6"S
P??:K\"LW^SY8)0E?O0 H7]4V#MEZPU\_MYTO6'868JT#N9*V>W.<8F%\[SG*+1).
P5HP9KV<=!!_.2M!R2,_^;R>8P*98I7DMFN5SA@];_)1VRJ/G.6\HIG\F:.T1$<9-
P'V7^TY^4XQ4FQK!?5+"*7"E;?QIQ#>"VIS(Z5+_#H7N<G11=FCX4*1'[E^(KYZ\6
P!QLRY$<<W0KT7E[;<!41]>1,6_\XA-9F*HB#4@@&7_@^O'A'"CP&SN=!W?)+/#OU
PC<O_O-D+1X"B]4EAX_#+GH(?+<L"PM@+TUI8T-R&*',^2H(XG!=(UA7V !EC;D)Z
P5=Q7XE_:GFG,-C]@B<Q:-$J0D"CU_&;%CR=.N'^J+8=+_<PL9%,A]:(F[PK8V%CO
P7M.O20GIZA4#IA/U;"EO.;SXQ9O*[^7@Z<BZQ/]A#T)E]N,F=K3FQB1MIE<_+SWL
PB++Y=' ZIYSV^C#,Q>)_HKDF]4==<[(8L;:QC/(4P^8@/<G815FRKH<R66>(MYD^
PG:Y07F1BY>$8WFDU@I>?#:8_@P,!M*7; =SXS;30""P#S5)!D38S8W9[?41%?,-@
P:LI^ \R.$]J\C*K>G(N/Q4ZNGYWN$=8SO<0<Y5;3V+[VF&8<:PK8-9R!=.ZP$O-8
P=_Y330#I3:<E *_S0CO8-<QQ$7JK3T#.Z2=]7!9Y+K=O(-3,%L\DAQV?(X\8+4XS
PC4VPM\14;*^59M]10(L)[JK$.:]S^8T$:XZ+]GHV.O,4'TPMI"<W(BJ6(O:*95R5
PR3 :+-O5L:27[2MIVJ"D7=I;$P>9K'ORFM/PUV!"J2QK_8R&E7>S^"&;#L-[/;Z]
P  .6T5)K#OUTBF,_4"GX^X7:DQOS0VYL,=3SD9]PS><2>1 -#7LL9(2(R0]S<20U
PX\-!]@;"[\:9X"_BX:[5'D;EJR9(G\/QUF/80$E!S8DS>+N68NX81K6_SO],<G.P
PPF)3,H'+^)%:^1:'-*H5":(L>8BFFGO'$BV1[GG*,!-#?[#N4<RJ[M>*#"GF-KA0
PZ08_R%"K:"LTIA(C$M;>,@;LY^L'5 A7<&3 .* /8<O?F4V>BC:>7Z/DO+GJJ9<M
PH,^%&[CXZR#I9Z'.//+=;)M7@("QXN*?_9+M$SI(X D>G/\B]>ZT3"Y/T/+3[]?F
P/%#HC0VR7!AG3EVM8G\K7H)E<_7?A-.W'4Q.6Q*TEV?T\)3OF<B]Y*GY'TR!NE/W
PM'V1R>\U=":@%,N\GEM,^*=)1E/$E)F4LK/-(EZWEC88;;H0UBD@U3T=NW&[;M0U
PKG&5RXC<3,"HW$<M43A <!I9!-PS 9OGZG;1!:L*WP8=N:9O2SUH=.P;*+:8OVIB
P,FQ'FB!"A@?C9(W/S 2Y!B$1Y9-J925F(3R<D5&0&Y7=]]XK?(MAOJ)2"*D"4QS7
P@U _0X&XBG0!=ABP%(R6KVWJ"G-\9-YMBB!)EC7PTU$%_6A(_+<L"#^>9:J;U-=&
P-'XPTH$JV@"A-X69K$@FZ!^S0G[B7)F<S9K2*W(DG&A27<9>O],R*&!".N#U]V9U
P3LPT@D7C M+TI>TJM.LO<+UPF,='=+I)D5=?)'$.%$2 V[H"7(VR4';^;^7MUV?6
PT%IS_+Q=R#_VC8/R5YJCZK(#TA\8F^]8#P2ZLHR,B/87)!_A.)>OB<^*?=H+H056
PEU(<9+>?'_%>>2(;4>+&<[R8.0US,6*A8S/G2Y.X%L%"/7+0Y.;1#6QI^R*J#+(,
P17<QGC+$?GN%_.,:I#%N':+H5+GUGSJ14F^ %MH#XKSA:>HUN?+( ]T'*W7320O@
P@IO\'Y6H=[H4S>[2"[L-O_>+':S[TW7K> XJ1*9#5NV@#S6C.PQ?-JVT76&[GB1R
PB&F>E*<OGT.B*Y?6VA]#Y2>P.MYV=@4OER18K_I-=TH;.#,2+)PMHXP?E2O2B4';
P>N&W>2=9<3\O]SVBVBR3D'<] <U(VH.(8'4*9(9D;S^:;8B1-%Q%KD6P".ZKRZVZ
P^&C+A#<C8] ,'KAY"Z[3=C:-W885%-C#$EFL4?J.WUC*87 G3X2R;Y. FJGT"$WA
PQ*H,C6!_T<L?-&P]+/J%GIC;[[$"(A-M5*0-(,,RE'3P!<9$6Y)-/JQ9H>J62K?1
PJ(<(;I^7MP_RT/14F&'<-C'T3S.)V]>W6,:O0Q2SF1QNXXBWTG4CT@#PA>9KYT/U
P;+3/#KTK?I?5WB7_GC6>GXZQ5!:S-(#: @^@K-H]6=1KVHC5IBB1:.7[Z98W[R><
P7:)5MICDK&?&\NDH%,DJ:I;"\W]K!*8RIP[(>Z4+467Q48J 4Z:<HYXA"!_(LVXD
P J&!^0)=2UZ6<K ]12D\=K<?N'3QAS:\!WD"GH;0H=AI?AAXG1A"N3S63CQ>1=8I
P];@IM:/3HY7;4'*.\&!$=1WB<>@0?Q<X:(E-S22=-$U_<3,AM^("[9)?@.2VS5VP
P!$IF^G*"#;"#]-+M?AE:%;D?O[Q-X5#3E6@LO@OA#,2M*;/N ZB-, V."TKW^CJ"
PH]]3F-_]SC#[85"NO/]-5I?[\G*2D/]NB#@<G/^'-CPF2CU3#;+Q[46-97[DUN6<
PVS9& BRSX=:D;]"FH[L:CAZB!K-5J22\V8 U,%/G(GT5&#Q%X(2(2FR1'JCWE-P^
PXRY39!8)*UU,>K5]@SH3XG1P2VDAWV,50%9K0K+(4Y]MM!A_NK/*)#D10@>4&R9?
P%N\\F (G%6)*5#M0XLK18IQ-(+*R01&GV+7S:2<?*'(;78(B&65\MN^,("]W2J_Y
P:P(K2Z%.%<7A.URCR%#(=9B6M 3_S$Z:1+#: @2P0I<D3^]PMZ_H#<U_ 6.CB;.N
PQT6QP-!N4Q>FX<EJ/MX60M\5I2<HXOG^#N,&G:T<K*1[R%:X7L@04?GKE:WR;QJE
P9#Y\NN@&1SRZ-V 0;(8/8-TW'&$\$/'\EDR8V2\M/>*%QHRN :;TO?/,Y(*-H^M/
PY<++#2_:?5$>+&UW+"!0"6+0]193D&*=O56CEG>Y-?PJ<,<K/Y"$>A X.V++9^1(
P<N+6;P2@0^])O32BF#!&0S=JPH._,5"N3A;'.P\$F0)P!<S!2BK'3C&H_*:?[$CB
P73L2^2X40?)N\%WH166YXR'&B.H[JSH#1_TN< YA6L <]#5;S&(M@XM?TC$T@\G^
P,:<+79EM!.L_ H\H9-].!3]'G(\858&N$&<=( 4M$Y>#.=D%*I+Q_"$_M2:,%G6"
P;B3]YD4?IL5MP##<;3D_YW(/57 I&S2W??$1VXZ[8-28ADVJM_9OB&<AM+86GA@6
PBV'D=-*HQZ6#701)TJ.C/"SP^9 ?X!BO@ 3=CG?Q@P%["E9C <5C9XV_!>S<X$YF
PJ($Z$LZ,98D20'7C0&#K6HW<?9+]]F3S+%I+<NREA759#1%<!'OU9!OM;F2?503)
P.ZFH_U*%: &6CJ.)BIT/FI<1(D_+S\H'X.WQ3#*R$20J2U!\B$;3KPBK8UV4"$TI
P15]L"UJ.V8Y,8W7)3)E/"3IE&\#'=QYVL8>[+#O6JU=[:F+'39;542U\N=QPIJF.
PIEYH*(5#>7V3M+W,7H$:-3OV/YQLTV,F&-D2?2GNKD(QS'!=)[E>JPGAL0W>G9C]
P5KHQ$%KWV@G4[5W:/$2Y+)OOC8LNUU[=J&<,16A,,B,1WA&P.C;4EJEQLJ=JLE68
PK"M*L2X+OJVR"7R;[?*#-L*B+E-=CKG\VY2K="L#60^)6A$8W4+<HR#,>T8S[KVT
P55J<MIKK%0AZL_Q1Q'VRX/9LS30@RA*E %]U@F*M*&Q11%@U84[SRMJ3US9+N&7L
P^9+[0O^B].PTT%.[X;0UO6O""Y%Q,^,<U;%!.];\K/L577JWQ+R%_MHHW;*! VE5
PRP NMBOH)<YK]5W"Y9_5E;81 :,O\LFDGGX ++P3WG>=^7<:CZ;]T"\;BKLJN7P5
P_%%"'*0,-MV5IO??*L'C)\EWJ$=W>@5WC,=U4\".[)C^ /M# I/;5<+%6G);DFT)
P3=/9*$?V3.Q4X<E#N'YRPZ4<C:N^KS76#/Q5?E@U0T1:F!VOBC4U KI/&CR# EG1
P$N3A,7OG*L@>_4[BFP@V.A5?"C#ED1>;TZ4J2K]6VJ5Z\:B [;'K+HT:_#*OC(]7
PS$(&DL6#)#3.PBAFT,J#G GS* C.0 Q-@U8U1)LGDBCS%7L?6>I_*K2PF7Y%0 %@
P%F ::JM-N%$HZQV64?;X'@Q]P5*6YU3!^:#WY!IMO9OJ)NB;-MGN6^\,!S2 6'-0
P\ &OIU^X\W?C1X5>I+UXI_S;35V9%^$H=[=9!XN(:@9&L"E-O[4>DV7X0=8NI7? 
P]69([*KO7C"ED</.MC4RSEH?;-SG]3S4V:$(T.GD" R9QIOB]Q%("3[^: <2I_+&
PPBN4((.VVO)BVS,Q4BTI20D&O$A_W(%)P]?2[WCH^QDT\0 EO5<6@>] W/OJ"QO$
PB0M+4+P!V]:LH?GNLHDLZ6CX+TC;.T(*M'^'+C#8.T5VH@,R-#AK@](01^<-,KT0
P-4@@OX+%H+=OGS^RTE,WG-[1-+VH97!QP'\AY[\K#59 P+";%9D$\WM-&J,\+:HZ
PMA@O'IZ-(;?K@Y&\<:*XW#G<COA[<C!305H32QH_3Q,VPBG_Y09/H;3/401*&8VZ
PO6V54*M[!_B80K^\/(X:YV;P& YB.EQ.[-_YS_;TIO/!JF&-Q,<ZGH>>K07N>[MO
P&P132NS:@8X]:*.LM7F#3YP:DRX]2X;1 I8/'DX1D$L%1YCK%Q#;Y<ES@'@^L-!]
P6%D*S>/U=](]!Q-ZI_]VGF+< *[CR7("C69*/-^]+T_":/%ARD7X,=T*USM[B?HM
PMMC*+,&)=-43O6BD.-LN269\#D= G[-/8UXKP?3_]5&D(>CK3B-H101_5-U0G$0R
PWBU,@[6E9Q@%0D6B:J-=X(Q$X9L(5KO'Q[(;DS;NW="2S,)JA0ZAX1/YW53C.[2T
P\KRHT0UII:'[F$WHZWIZ-43_:1(16><T7'"RW@=XSVM!4$P15]_<3!BM:D\"2@;!
PLL)L&V C& ^ 1DTPT%Z'W)_:4)UL1'>Y%%N[[N;4OY\I"T4@=I3F\4J-%#"B#^-/
P(!US-X,!($'ZL!G-\@+$Y L2\0.VEUJ!_E52]: .Y. #E5+<_$J=2<6[$X*?/-V"
P(NV> #EL0K9OV9O04(7HYW8%%0KR,C!&<#18X+D5,!Y'[XE?AG&OEWO@V^B+>'=4
P\*Z0F0>YB#0J(PB+#1T\W40&B.S7YCA#%:>/@IO\81OIGO<_,R=+P9,,,&HHTJ+;
P\!\/,&YY8*FMDC[%KY&@-H/7,-(A^+4-25,#@N^T8RK6W\GLR)WIFVFN=_!S!IQN
P1(-GF$-<GI_?/8X^.8>_V8Z%7MEU+=/WL!YA#.@U^[YBHQ4DP3CBP%B'<?>S0&[U
PGWFQ9H/+Z:D^OUEX90QM#/Z] 4=MQ4;9T)!1,$N[=$;$%YCZW5-+:6F!-4@QKI]E
P;3A7I/JP;@N@(\>6--,H=4T"AF\-Q:&N;C41>QQ@L469N8>3"M/B)AWL0O0HONF;
PKZ$J@6"7F=HW;#]2"U'AS!<86X_]JO*=HSEZ< Y<2>: T(;&#_NX*;<M3,EX2U1_
PK<]4*O].TFXR4C/<_K>5VSK.7F$3-R<URG'L>UHG?V7Z"J/#.]^:M98_B+.44-3^
PO:KP;((KL"G&QJ5>1M0!JN9X#'<N/99("%;5!T<""G>9T8<LZ2FL_6D>-I?P3*8G
P0OMO35/<[MC:289=J*1A$DCFO&9,L&ML/8_\I2)4>=9G:Z1Q1OL9=0>FZU!8-)S_
PZBN6G:.Y4%\+%#6NCKBO_+'I.XW#(\;A8G36:Y,_#.P)MQB%V%YC54INSPD+6,9$
P!D<BR7 (Y:_ZYJ0>:!T\2603"_KE=B:<7^&5>9N##:6'8,F(8LT7AU,ON _SZ>+B
P^N-8;C9I1,FQ6.U ]%MAC%LXIX3TH"[;1-[7@F.JQD)M_::GD\?%R;##K[C'VQE>
P>S=<>1,J7[1GC.9X'G^1%*6S?'PQ+$X3K/(?]0+1B&>,.UQ ,OBN6NW;@ ."/)BF
PDE@93FREY7E\WH0LHX%F!^3^W$\]*Z)@U57W%P2;40OW9"#/;IGZDX-UH;D1NB 1
P&2YM#L T<BS_(2^XV":86WMXA<G.,1 9FOY(>T"KVY+EM>B ;*C@:LA*?>O9Y'V6
PQ(Q7U,ITZ1JQ .>$=NP++-TI3.OAD*'=:,086-#X.R8>T8DX>>E(TY 4C@@*(M^<
P5EU I:-H/E7"JUT<)]<L[+@74*5!KC?6N]JOZO1TT5R^950ZE8"-YI-ZH.J1 FP*
PI:;<S!$A=C]33F!PVTH44^Z4GZU,B[^%P&@3;)+1>D93+%NG#*95U2AQ%N,G+$O1
PK;'1A'??KLMY0[AVL6G\7I9,,;!BWX_D*O2F)OF+;)OJJT<<H]#(LP-Y7POG-:B>
P310&<T(_\=BKV@WDDM94H",#09HB<@L9900&RBX]VXXJE//0%L*5#"7%9 +>BN,[
P8VSP0H-\FA[XTGXU:<B=#=&HNNC1%X9LJ2U, UJ*5$?W?>3=O\'^ 6B@DZ<7VUMY
P2U.V^F3QC2O#B"?9>S\$</@N6A&P9QX"[ 9GLE)V\OS"<6/+KW+]CK?K[NS"']X 
PD7_1ST'RN4^G[2L:OW.2'*5HUG*6-8#>(4QBAU@A!%NO;WY<G9KZJ)6Z;]ABTSPX
P#$O/2T>&3RNI&HJI$==<4=#?L!O;?!11[U"[?D=:I *<!\6B%&>DA:Z*(RO3*Q]J
P-IRCR]#="\.MON:<2\YNAY+\QDUZ\]-V2$6?11K?,ZKX[5%$2++[7,N7]5@1;?XW
P64>,@V""%II.9N8AAD4YZ 1VAMM$\ Q('+Z?)+9; )HO;,Z;/ZQWR"!F*CX )E2[
P7E(I,L!810 KY7)V:&*+@XV]0.S+H.[K\"19?.^?O="S^'>)@JCE%0G656GZG I,
PBO861]!H:FZ<%W=G(>O/V5-/GJ@^$4=D+VNV'!QN%*X79)LI+,AVLR[3XH-EM6-U
PG1=XS/E*3;('0RCQ_KTV&)G4F^R^3P\_.A5%)J5PBBD9N\*1B<)JHSSZ9GN)0J69
P0@1-7I*#5A$A6%\N&]>G+^^1)FG"KT08.IW"^<43>L%F.EB#3:-T>]&R**/+5:8S
P>!L.4@+O&^,CASJ<JQ.B9MAO8,>ZQ9WJE_#* &E** BPY+YX#N1N6:7E1=Z>W0I"
P_712CTQ((J+O.@&T;AD)>V2.;FE[?UG"?HDY/"G[$<5]2OMMA^)4MS\+N<Y;B*S[
P<*_" I_BR[B'U!TH1=Q$86,'[Q'A\&!C<#6=X P>01-W^PK#F,49/]^"]04NFI!#
P]$F?X?Q"?TJ(HTJ53IN4]!*%X]!2K-R-%,D]!8^9)$E=/ZNP(B55@O1"'5\%B"9_
PTX[AV@BZDPA5YU.5#AA0M^0X24)*%P*YU75D#(\@41H08"JK**Z3/W?DEJ?J;J U
PO0KW6' TXXD$-QJ>U(U-J"P@#[A@4*%UPU?:@M<#!6]F [Z ]H!E1&U6#FY;C2G*
P)BH$W"I>'$;]-C>./>36=<L;)+'3$2(F\5.Q9L&?_ EXL'V<H)0M*;3#UB6 FC5T
P@5VV_9JPQB,W;G3_U!8)HJB*#"3.2VZ&2X_=4+[@*_<;VU3\K;-!+34IZZ^1.P,A
P4N7GAI]!XU:>(^F<(4TW)=+YLZDM:V Y3&RQ$YP=O*=B^SC)H '4_K&$(<Z@:-E?
P@Y-^S#.\<0V"7Q=GLF;A7'=Z'F'?7$N*^^:GO&T):?,/OXC9L.V*8^/)>6#9LIUN
P/M]=+/?!_#@6KB#:5#7F%+W]OXD.6&\K!6(_*5YY1EW(#C2,?+\S:.\,P<I3Y=<[
PI5=40;]]'DA(;B3#I@,&7#Y&G#Z@X&TME]4%3O=XU2/T@"?[WUS2E\Z@96)5QKF*
PM&1H"\3T'8+5:0T1WHDG3+M]"Q[\SJG,GF!I#]G&$=Q5>.0;P<4P+-7D94U#)G'U
P8ORD\!M?CPL7;GWON WN-X]Q"8 L0N ;M1DAOMS>&XUTI;_+/[AN=&9 UN@OY1HA
PF5GDR0C18=XL!C\JF<A1&D U#/5])3S#Q5W>ANW/0M-Q, 9W1/.Q<7[G\ Z&P'[A
P]'Z5OQUS8XL<;P.@*AY_YY&V:T%'.NI*:S?C>M5=N'V5<\SFD*RK1IS+5=O7G7Q5
P5QUS"L8&F7N,]IMMI=9B/\)-\L'70\:+7L3L1,=_M4%[UA7DI Y@C"API0,,W^SJ
P]AK#RAW9^E8 JD9P-;4D2"?L6!VW&@7J>H ). $6]R8=*UY#@+ZH.@EX'Z  )GBJ
PSFFF)K+5[FUJT8J3D)LU(N0/YD^^K->I39ZD]B,NYM]P/;;[;D<;1?"A7YWNP,? 
PD7H(ZV[/+08T62_I WLHO7;5/<-U78?(4LBROPL<]F"OD*@3WD<-(M<D*90\.46W
PK\4Y*6E[]W:[%<D[\^"WI";,7R3:["'$PT?KYO?'"U3#?EH9 +VER\%3-)L#(>A%
P9&I&INYM"QP[1DJ1$]'I#0P6(4B%U,^QV DU4.V,61DI<U_A69"C180](JT"^(Z*
P5BG4A.HYNT^H$ZE7M7]$D;=?Z>EZR$OT90TJZQCQY*#5ARZ5+ER\@JBJ;@8_=^H_
PR!^H54>O\D#\54_.[JLR#>Z_M.(FM0&K4M1#^<)[]V:F3V4$'",*@FR:./7,65'E
P22(IR3P@:@<UA7OV^H3(%CE=2[TR$6O(J+NT!(<F%CXCY^5D?4$4N99!'G!-(^!2
PIND9^ QQ40\:L,H8OJ*$:]C;U/3B%"3<I+97R(8]@[(=R$MC+%(RX !$_*S(Y'[H
P]QCT=\/?&A'V*J0E]8_=8"L9R.Y2&F]<?&U_2A1N_CU%3:T .*@^5_T]RK/*_B4"
PM22^QV3#A$O=JG.9S&/.M^ Z7G6)$M6V#LT[[V@S[RX'S^!H<\# $CSP9-9F%S!_
PZ%A)GIDG)JKIP0&T"Y>T-L.D+[MWCOUPK"QY2*DE*0#/#'@_\RT?8-IAD5?"UK7J
PC-SR$/]>&7SB?#:G]"2<V'OHW0?<)9OO,8*3V"=:;IKLF+"R"]$WO.)(V'IO J6U
P%DS\A F"C)[;!:_UC[WJ>]L8/28WMO%^/I5!>.F/A%$L<,'WXV\CY6T@+%"FLZ4C
PX9]5:DSH;U0JK2)WREOY9G?CMS=/F<% ?-7L7SUI:\'9!U_(<^\_U@_C%?8DAB:S
P"&HT27"E3.ENI$E^$_Z3(!K'Q(C12#)DKJM!U3WGX1SB"^Z?V+ .O1\8YFUJ&B^&
PO$ICW,JFKR'(IA0WA"_9_('"$ ,S:*!X>!;D#@GE!>\ME&\GT4,N!FKBT74\"BXM
P-8KI !VPHJ5_@J:@MR:-;GKNGR)#/R>5@]<: Z*V+=W<,QT#_E#<R.M\WKAOJPM@
P[">$2QAD@ON6;3&=C'6HE*H*@I>[?C68V3 8)5U3^O$<5?^0T!=J&.=G87/2RC6[
PKSQ[$@[$O&S/&$L$,M00];JT1$UIF)XD4.DU1]L!)+#_TZ&=#1 )RN^ :SN@&[Y(
P,$/(>2JV13XRH%4>^&/HA[A>2UP$L+P-0;#CT)="!NNFCYJI%&&B?&UF[ 7\#E3R
P^OG6M"E/0,NSK2Z,PC"$LO8--2/IA&$8S@P N@U',4TQ)"W5T?1^T1U*_C9TPX+;
PM*2L7\*9S.?6I6;N'PL>$Z#=JZ)3*MA?; 2"(XC;*[Z,\##T2TEO$@P+WU8DM& O
P"!C[7]V-B*ZV"[%G5VZO(FZG(R]@M-&$,(#X?7S(?]0&';:9P[4N^_TX%UY56)Y>
P5+7+!T:#TDT!P9$9P3GI1_Q*/#;OT$%4XBGST?>H"N2)$Q75S;SIUZ^_/,=*V=,-
P?LLCG&HK^2SG ;DY9*FQ9#-$>43+PO7N)7(S4X<AOHQIRT;F,,&HEV7348,^_INF
P_X??? VOWJ4[IYW0Z$V-%'B74NX^!^-8_Y&G@?<D=WOZ\GK&[-T^&UK]H %8"G=7
P><1]L8-JW:[U>4/?<-/4N%'W/KW!2<C__EF'FAJ>4X.X@#@^ _ZY\6XL1U7X,A7(
P]AAE+0]V-MP&?=XUG-B$_^/W&WL,%#J=5:4/#]'10WPI)5V8J9L"_=P[,H0\N"_N
P=S(><0<,AAC.X-U'3N&7.BJG@"@LL2HW1$@*!Z]NB/35B18!@&&A%/?\2U'T *+]
P?X>\E",1IPY6Z>=+!M9EY/.<*>CB) -.4/UU<ZXZ+4LDKZ&?XX1@6)=]NSB,0+AW
PF]$N\5Z<H8<"!_91)U4\+*02SM18H1;5%Y/>M0V#VGJUY(X.5)=94M8K)XTHYZ+=
PT(-+,O>9@DOYOEF[1((B7)?MBH[YY2(%NK2B_B=N$^'*,0#2;(5C]GC[Z#*ISTVG
PE7[=/F,CB/<YV)A73)P(M .BS6V$?Y6E8>SNB*1%Y<O.RF4H#''F @N$&=3:1<C3
P9+7S#?I(T=I(%8-E^!#E G1,K!B;WJ"H>9K\ACK&QB/52(BT5F4+/;U*DFH65#S;
P2, \VV97I#0WIA#[RMV !P3Z_./B2^W>)1_BI:_C$"N2S?$P"A#S'[F_A8"T"&HT
PLI;4>N+I78>__+=B8PS9;W^#(=K,G)E>(#]B.2RQZ(CU%&>QSF@>?D7I;XVR=+?"
P)CV+<.,.*[8FQ5W%L"8V:=C0[M0@^IG6SVOJ3&0@"4*.&4G4"=<OK+&D?7#_;T?S
P8O8KG-0J(/]W 7SF;^.8F"#%@#0C1+J*).;F4E+V9>R-]. (,N),B)(-:+N]X7<C
PW5T6)@I63(6!+6+ +M8]%N+4HKQ<D_20URA2=&#^BJ;;^.UQ2>B11>E<FD>5@4($
P53R60J0G2UQVS.UR4#,DJ4 ,!O^"YK<\O/N0SQ5*< 5O,R*RU-=0#;W,'(B$+H3\
P^UQ4+XLT>2R\>G\I>L2H>FHM\3")I[4HA934#98EQ]$;2>P0+=Z-'KM@[O5975N*
P2[G ;0%0CLC8,R$,9.&]@;*DJWJKQ_PS:(R6]>$UY<<>4=N6PW3B=KHP-Q^P:U<7
P7VMHA,$@F*XEAK7" 8+Q[Q^#L13GOR*Y]N##\7!%/RA5/^I?9>E\\4_NP?<J4\9W
P$P^78_F'DN.6)^4U'9+QM2@0B;\S7IS0D0635!#6@0P4F\'4!;9RE!4CWW'N/+'^
P8).P(3V)L2LV7CFOK>LBM_ 7GWBN7U-,PBQ9I5&[RRCT._OW-R./:1, @PD,NH!1
PK?3S.+6G[V!TV BXJ3N[P;&\+">P,WH1(-9+3NC;RO5XO*S+5P>Q!%E.;-^C4!!Z
P '@<4VDQ)_Y3S\?3U#4Y0 ;'9#XYR/TF&!5P)Q+XM8]!D6*WB =#&2+YD% *;B6+
PHFQQ@?X+O]$)H4O0I)XFG!9Z,=,)GB(:-C85S3.<OL.Q+:19@95Z5;4ZY_HX1Y$R
P>II7B$4X^:_E5=!S).L^79%:V!;CT \/5<.ZXB*Q5Q'GE(-!"6T5X[9M_)77VV:3
PL0M_C\HEYYXO9<W ',W9LM>TY)QN!I:6&.Q*WW(X!2TQ2*H%F66FFCLQQ3QOU;F7
PM4,[< ;KZ9'9'MPU]E<J9J^"H>0I)%"_S_5TY]7!%8S 454/0 +J\YCP*8O/KK/(
P*KD 6XCP6T[?I/*/1_QJ8=S8_UD='3)D5J7#])VC7W?%3<:SA;>]9;J7')Y#>C%V
P5 N0P[7(<HN".AQM-1730=O@,C69I$J19>!P7/N>T2<Q!5!LV*;!' 56>'S' .+J
PQS )&FE[(/B]IZKRM/.31EO?W&G2T_/O3;ALDN;P2.HJOI6</I">\H?W&C^6L-S=
P3P>#(5$;!C8U5D&-S_F>ZIV@3+TPGPZP\*E6W\UGJ8B, S!F*:[<T)NRS1.]^1.)
P@S8!0K$.C,MV?2M]_M0\<60)Z5Y\'7HIR?]HSJ:LA/F <L&A^6.8M0Y$]?IW 1<;
P*I$UPG#S%[^21:;3.0,6$U)[TOHD9$LLK' ;_'2+8CKG9'/HN3F#JK/[\,+\-' =
P*;;6[>IUR_B!R5U)"G!)(RCHI570HG&%1W;OPYG(T04\4CT*MCS"!9R9Z[]:R2R*
PH@NGJ?K?P*+WS&SIN/L1='_V3UL'Y-N@$"SRR00]88"#"HGCR>'9D09NJ+\B0-MV
P^8M?AS\_%?1+>%],O/@MVRF4QRPOE-MZ;G;I>.>I 7+6)DYT'MU=C>&#R]D"L:;1
PC@EW<6/.P&_]-6U.T'$6:<Z:1')(5+G2X&^LHE.M_?'5^LYJAWR 'ULX7/C0\1-O
PB@P-#?>SOCFD+4EL ICJ.XT6N1M)#"]".DL72+AA&/9,6\*M,"J!A/X5P-'I49\T
PY[Y>>U HO3:+E_OWNW?$\E.!J=:I!1UH>_M"3"PILONI>6)U">:72O-K. 26.+8^
PV$?Z:IDS9LQHQZ0"Y'%MLPV44TG"F3?WT@9OG!,R>L=*DNG[@^ =13Q"[P=_F&4*
PU_5UKWLFK[ )N'2&# 9:9D%H4$)_L6UAG"VG3M1_'SW1<I1N"L;#0VCX_P_^(O'\
PL*RXS.IUEK+GBH/A9<B)A7D/)EO2$^^/CC6FZI"M0NY[+1LXL]"J^2;R.UHJ 7[$
P=U%K:"D^/ XFB$<O#!C",F3*-Y:O:S5<'73P6#!\BMS=&;@C<$(!M1U::LWQYT97
PE@IT7]"]%)%[(R>8YC012+]^W-,:7@-Z9 P9LU67]SZ*5'C+T^/&%A%^]X7+1>*[
PJDKB8^IUC\W+SOFJ');EO^A6H>?ZF$IDK7>,5=X7,+8M@)T)8*TMUS[6^T"GVWEQ
P^%'D%<Z+2N:G!J$R"HL]@CE:K'C!6H?M3E@S4Q?UOS(2#S^%,4JPSWMG)5M:6!6-
PRAO/>KH"1'R;5S>RU8M6D1;F8NO!+.7QB@*7.)?"!GX7O-HT\3QY*GI8IX6CGV]N
PQXH[)+S5RL?;R/CY>\M3B'25^=- RE']H.3IW")S<G7_AWTRQTG:F)#B1][B%6U=
P[;U0=IL91Q"2(AYF\ ]#\K/&?BPF;P8-K$2I,B+>&O[9U'.NJ<8B]<X?.[S,T@%B
P^.W$B_ BUB #'^[C36?U?(I9T"&9? 'JVT#3\2O@T2$/3YX<C)$%JVZLM9P*%Q!'
P)E6<Y7&?@Q /R<\FX0KX+ R3'+"M!8M8>+71G-=8]_G2KM.N P; 1VQ41I:WQBX^
P3GR](OPY@\0L2-U0KQ7]"0GJ/7"@1O60D/9.P4:';Y=+TUJ2'% + %\H*'L6=3&4
P=#Z7$ABA2B*/]7-D 9U*S-R@*[:F[+FH? -#M7]7SQ.<X(%H9))ZZ+PFW#.#TFZT
PK,-BL-0+<?JX2;,]8Y[;7RA;6?)ZGSI,Z:B07GW[.).!<YPP -? (V:*XCP':R1<
PAP6D,$F_ZU3W;0=)O.L++:P>+7++D-X"^K-M[*-2*9;.I)MD;.RLB#D2R'0]CMC:
P!3IORCW\NG!*(J1!+L=;R4(^QD./V-::! P).KI&, 92O-,4=,[AVV"#1/&V_"A(
P9M\FL:F6 \2P*2I=5WQ@ZT>0K##K3 ,4':1HLM!Y0\78V2T.;H^XC)3C\O9%='\B
PY@;\\6!R-[C/^&$K;>CRU;Z*A9X:-R]3@*1 5;D-\6T'+@LG=AKB#IS+8E.$T;#9
PCY3>?44Z)4CCNKR?M/^911W81-5&%\']LSH^ _ZGS<KH477_1P,-5\*+>IP (S?,
PQ]EE\3T\2F)&.I CPX.[0^SZAD"2O.KWR)0Q99I(FV!R447=)NSIA8&R*#,^."E6
P&D26E:I\?F.1Q,U2P1C<KY-/\*!C+3UMWZ45,HUIO !V(5Q;8V6^B*@$,6)>,<-Y
P>4GZ#W0&U77Z3TC#A;,$.*CZ.&$5R&&ZQ29=IT6@KO>2AJ6>*:7UX'ZBOH ZP![I
PZ2A5B*=Q7UUDM03MPY-FT@<Q5GOVI A&*"=6B&=JH$@T2\E5=[\/T3TN%R'+]\JE
PA?E%XBE,_CQ]2=L\T^Q?30S1_I<'CO3))BP FNA5 [>4$J]\)?P4@/\%PK/N,Y#L
P'8#+PBZ[\%JQFBQ2P(5&>MUQ733@XZ>1NC\L+E?6K]!V9>Y3J"/\\F&!3H\.)R E
P$;1N&%\XSJLEJ7:S*8Z#>8;?KR.3K"5.PL'E0A3L*9O5ZV;%B5=K: E,,Q"/IJTC
P3]GTD72CLRGA4#\\=V%J6(=;L#D.UQ*CO??WQ1E$#PK>^WQK;#+G(1(-AJYT6CB.
PK>W_P[M"1<,_^>KFFSM79?W3!;,*C_,0@/A!TZ%!8<9Y1KK7P4>NC2-% A1.REYR
PE-NSP07X41&=V+:V4[K4"L6DX46%Q+ U:/0'+;@]9$2:V=D0FYMF8^*FJ<?!A>\F
P;79L6>5A3R*X6@+<*#3\\*>W*;<!@FF:O[WP(>)-<,B]7$32B?%0!\9D%D(]$O?I
P@JK8B\H2>BD-;MJ_CST<J'FU J)#E6A1CA40YOP#*+"R(>4WP/GK5DD4;N>J$*%Y
P-RA_[I<"G<S)8>"\IC$U98"HR+%]%(BVG0NZG-)XG$YT3NU;'ZF5,EH^\:J9L\PA
P.T2M<9RIY CL@4<4P 18_)39!A)\',!$KV^9U$_?DS,G<!KNDN449-I:"K^0)H'E
PZ0#0V)3@]'Q&3;&Q[3'J B[&6)>WN0XC;=G+-';9$ +:28'%T4&=7M.7</F W_(3
PG7DRPX*"CJ%R6_V>&M@Y7LWF.-"AU8Q4V1R\HHY&D;Y;)9F7*8*I+^!S&DV065JM
PX:)*CNU9'7/_L$*?SG1N.0;-\,H05N92X3S?DS9!U 0&>'C4;5"#[--Z"<>0NX:$
P=QOSOGQQ:(:'Y4HIN7D)#-D)<,PQ!YH%P[RS>=C7=?5HW^3 (1FSNNXTXC?EY^14
P+I$]]P93D2H-?.BH^E4-]S/HMC>N>,V8X [Z^@#FB"YI<7E?5Y,SL "W=1+79U2K
PCHT-]QCJRD]WE):.'X\FRLLUS('[X"?#9HF])?1#LNS )B0CK3G;I3X(+)<:(<N1
PQ;)ER@(6HPXNMXEI%CA1W34P_9W8AY($6'A%>8Y*\..J# !II]9A5<:-PE4(7E30
P!'1VE.;/<@59X&G\"P00IYLY(;%!YT&S7H5&0D1N"_G%3:._A&E"L'VI\37X5I$:
P&^;5\W%_YYQ_T)=T"!G+I-$PB(N6WM\8Y#&A3^\0 .%DLJBJ9A\_']<-/..A>RY^
PCZK1#,I;]8,,^Q/4I\B'2I\OZVG1IX?<E2=5]GU(W;&[;Y5T/MNR2^^J>?\29.L0
PBQ5Y"9_(E:;!%PJ<=E!F:(]]@DL+96BQ'+=XJ/$"=Y=J>2&=OX7F5MWWWUA5(0[W
P'2$$93M"I2,MM;F2DS*-T<3>ITU2#'>C[& _P^0MARJM'2583',A6SKEOP,<0F6Z
PT$=X/UK'LW7YM(M*2UUQL7OT]%?)P&5C*4W.F$Q+BK=2>;?$<._2>8G9&G&H/Z$[
P(_9X+2^K:!-XE\O)3MV\>VC#(SG6'>%*/^C.&^\MQ'_E9[8^]5BM61CG:G)(\>,*
P>\,PANO1?]WJ2MU<<W20L&&#;S;6\"/&K4O>+XJF0@7S8V^\N6D,$]%?MG[HXCUJ
PTK1C1AI&K!7M!<9XBIH8=#'Z^H9\5C20FZW"79&^<VLDR;G*EG!D$-M'2K5T>/^Q
PVK6./DP-;>$2XQ[I'PM/R&T^O&A3=,RYPB5G#9L(FSTO+SV .E0=F+VB,\P_E9"P
P[(\:_^K08M2I[P!S0,RI/R(L[/$%][XB!(5H<H9[TQMC.ZO(S"IC 36&O$1;XB18
P<=7<QR!?735MZ[:5;F6WQD9 $96Y_0];JQOAG; 4PT\129JI5,JB3FE<DYTB@$%_
PTRI!)1S5-)=^'Z-RX?#_PNWFYFP*,_6<_<^9F"'DKC]1PJ,>Y=4BNF1<)@J 4I50
P'$8^$+9R#!?L3WMQB^Z*%^.%LE 78>F^M!3J?XU*WA0C.LR_5$1KI:!=.:-*VXN[
P">:53F9<$S23?FA>8" UHH?JE5QR\,\3S[0#J)4+N56'X_@1TI/_0@J@5W$^BG-)
P@H3TGX3[;:&"[E\)9?@!QKD]I'-^<0X^89\*-0Q&>%\ERP<+[XO/"AD!:Q6<)C"E
PZ[K^EQROR6)KH<9$)CNOOH\)^?*WIO<-)O\AFEKA-O-M/)))<ZS\&M/SBMHG3=_K
PM&:-(E#:?GDCY%F"IKP,!?$:$/I5%(A3%C&J]22)R5'AT29*R)I:4"HF29"O0YQ.
P&%65,EJ\)='C-,R<LO8(](I1QN1$DMGUN\._LXO4DN:+>MDF=DPMQKJ;G@O U,N&
P@20A(RWAP7L]PCEPLQV""$F.FYL; *IOF,^ES_PUDHC*!;5K!A6R0SNC\]II=$K+
P7S](&P$RG""[UFJU2*A*-ZWT2"D.819=AWT'5_.4Y!OWZ 2KGG6B2U[&B'X>380\
P7->)D'2/)+<A@C@%Z<.G$4-X(!$$AMF4!K'&W@WSGV&^K56=M(=KEBY\:W6O+DPG
P?-WV)]&D:',U\6=$QIHA<> ]Z'VRH5J=2XM5IB?EZ$0<@-<+)/BLG8;%((+9*>&7
PEDLQ",SK<N;U@?\8:(9+*8"J6<Z:CQ,?5>D$IR7>J7-SD,6Y=B3HQM_)S7#;7A-Z
P+&P3;=];0,J$R<"01>"5D/HG%D[.'N[M>'5/?]<K]GAM^Y?;0*H#53?LK/(AQ/-6
P59&4#U6Z3OU)@[Q9XF@A-B>HEX?(/W2R#7OGL>$49@M]>]S@W(G\]]3#ED/Z]2:Y
PM#+ L5^/)U)+(M )2"=CYK./[).'IN5^$8MYN?0NL]BZKH7RD^N\L8+?24NJJKR]
P\G.R1.;\%[NDWHO/VAH?D(@'UM0B<EO]BL@YO.L6S<%^;C99M 7:@>,9 G[D[K#F
PA9M?Y35W=/Q(W/H%%1=-7D#<N^U0Z5<VB[W@"'@7D'?(Y2T2F-7S8I;L&,4WH<G2
P,?!GOK+ZO\,;+'49WR&ZZ<0N(K(;D3C7"?2&N=AS:]9_<G8Z13!;0QY/J2)L?X\^
PM>&P%M)DQ]#DE9?=C'4*:]']Z^ YO<6Q.LBD>"N5+@JRH<X*-W,0+E@3CQ1NO,7>
P)5.DWZ:7G9HZ990OIG,;)NS-S+']=M$Q+'2\C1;&X$0#BML2X7.G,O20IIG=7TX%
P9D]4BG+5@;K42X+#KRM2I\F;;7HZO$8I>:T#B /M([^VA;H"O6W],(6'T2L]J5=M
PS;B63<5<6B80&V'<<=?F6XVO3[I\'!;6[DK(]4;[6G.),%\QT[C.,E<]7?F0OB?T
PR,-/C.XTV"8)5GB&JJ-1D6(N$4BA^H7A3LZR]9D-GF<7!(FFTMWKC]&T-U\^, [9
P/Z^0HV@T4SQX-:CIOQ]E7D1[I2W?N6<2LW_IS9PHXIH]'CB5W)@$&2X,2;F6D!0H
PG&66%^KT:;C4MWKR4BN,T#W*@,HW-?ZB_^P4YGZ;MJT2"H3M] +/>SV#QL^WB-$Q
P/7MDD_ )*0T^XR;A'G/+<Y)AZ]K7[16P'V(-@P9@%0MWO=%%/_M6=?(W=] UJF1C
P'A24.??2$+,8@_,PAHH@E>V.F+6MQ'1T+$P(#)I!&.V)0<1&,]T)F5I1IT6QLF[P
P\\ZX?PDEYW W)Y:SH)TEWD3*FR2FJ\AM(VP+IOE?FB! @:F5[+%O%)50 N4<3%U@
P3>S?Y_>\3RM!N\@2H.;H^4CJ."3(PUF;82$K46]N>*(_*%'2P;Q4GJG!HK!K]53J
P0TY,U-.^D".4^O#R _.<^LIL\HQ UIQT02>*O>3T4RNF5[@7)?-YD+I(3QZ9Z6(I
PC-FE,5]%3M."$/J>FU@8D$O]L1XXS?AMJ P>@@X*=T>J\(_QU<^.D,2KALW$>86H
PV"YO=]/1^]D+>62\EXI9<X37[/-,BL0*T8\K&QB&E(*,4F9=PGX*NF+W__HU*+W%
P#?'Q%:*;[8!OT@>K28D85/4A^O 2)['<UDP@K\W6B(DT7)^[Q$74PZ(Y)!9BB^)I
P(66A_C3ED6<&$Z@OI.@R\,;^X&+URNU-%F(K@X$&DWS4QLF;9$_9>QI&(N[,W%$F
P?Y-XZ%K*(,RU25H1K)6X26JWS?1V$T]TV$:G$J;,QW/N5!\J2&P+'-<S6*XGJ%V3
P.J&:!0OUF=C%@)PK;^B["I*NC:G@$,._<7'U(4Q6FH*\A*3JSM)QP.R>?P^Z901;
P(4JVN28GIA)CK\-!+6Y:)_F7-,GU([#&$6)O@D&SOK2<IT.3P;1,[^5=["J.)D9H
P+]7JYIHLOWUPH1,XE)K\0+4'D L2?K::N%(=I$*QYP1HR,WG+:QK!Y#Z01.["9O'
P&;:NL+BVPBANO J2N&*7$)-]"J8/.*GV#Q$U(:KPSB?6$$6B4Y);D<"@PX\&QU"*
P.\.SCQ0][-Z;Q(&'\,5[/CKF2["H!")O$2[%9J[$;P1.R L?B*4<^;NY>$->L5OB
P9 <*XG!#>-WP&E]I?\T:@9_L#/K: A6]%5T(A1<)UZCY2\_83>P>SQOR<T'3*_7F
P.8;<L<! U&M<\*O],"FVJ_\0IWR]"=<3H]UST%=#)]A,-/!AT#:>38J]$.J/WB+K
PINF8-?GGM*"IRB,0K0NLV;_;K9J/!9-?_2=,P.4Q6_V/8(%*MK/?6!@)R-9MV_FJ
P)NT 8!S=98)V(/+OCT17F#W#*)V[.-YUPFR0]V/:%P'1ORK&: RM@.5T@%57VW<#
P"%(:X!%QSD+53?A;1'NEMDF55P*N%SQI*E>6_/,JNS'%EKV/[EUMUJT1\VD@NHFO
PKA%OR*T#^Q7T@?KJRVD3)M-L$JM9*J>NDVAX!\) H29#>"=>I,WEBWIID*J?<0/C
P**%E\ AEG,JTZN5X[ P# !Q=W A#L:_"=%)(6O@^3@-47*$SW:I+TQFW$51X1PLQ
PI?;2!!OVY%[2T3DRND8%P-50,<3#D5PX/G -S,07\=2KG\>>.L^.#IDGDR]B5WNY
P+WYZLZ/(KF.]BQTS>PT^V>,']2@VFXQ8;_H:"OWY>#>V#[&WUCKG67MF1M%$-/2D
P"_!\0H/J;F)=>]V;D*&[5*WDV(T\>./9V8/GY\A$9=UPR,WRV;KYDJS@6?4&L@-T
PM"OF$8WJYQ2/50;69-A\NFW);\DW=S3']OK(5EGR9?7,J 2P,\_V>*7\]2+6AI@Y
PM!#"7*<[2GM"Z2^]AK+G>\:KZ19<]6_S;I8ODB@)^JDKW-RACZ1@K\-_!O2ME$% 
P)7L0Z>,V5DVQ<#)JU[JVY\PX\CARM.+QA(U7529BW! %G9()69F,YI=[Q7F*W_*M
P5WT@PT8S]# R>9%O58!G^."]_-E</S'ZH2O@G/'-H0;T:P@>K%)"P#8==G3?WV I
P!MGN.A>&(TT&"&L5(])0"^@*C]<J5F0FQT?L(H?-:7'^=ZX*OHL5UW<4E7G30)O;
P/L)@L,K(+MBL-V,QV&GU%RG=<@;2/>75!VWRI&]"TQXEL"2AV0%7K+J86*#'WBXU
PD8CT( 1G-_)FRZ-[L;RUY/U 7^&HUL0TDVFE1N (J% 4-H8@:10>!_;-^J(TR4A1
PH10&:8HE3U9'M)RC6/Z>2,;R_M]-R"1/IUPA7ST#$-I37D9N@72NBX/#X2<LWB9_
PNLG#6!=^F=5>F0J',S'X:(4;I.0PJ#EAWZY/@JX;BO$?>VGVPC.'2;G#CUMIL;E_
PL^*='E>XF9=,2Z@7]HFU2(_(XJR',8+ ?].1I*TF[#P"9IR$8:C!$)C7*#QXFSLW
P=%;YU:-[/8HW"4\YA=)&Q8.*B+,75X&*1SF>G*D%QPQ#V;775T8Q)+":N<? K-\K
P1,!,M.PT5C( ;^F,^QJU#4\!9 \X'"L36'@6'>Y0[TK-Q/P1%,M\-EQ;^#SI@*>K
P;W& HOW)B8MWVV>B!1E/UF6U_S>*J1V,6GQ89"LV?_RY ==,E0,Y4,\BCG8JMVZ8
P>B,70G7Q-03O*E,P[T=Q<P\31LAEN<M/&GYGQLF-:NC_M#_HL&K\@H=[\*$[?#%@
P"1N8@H ZM7UQ_3)O,(RD!WO9JAE_L] =.-9FF;Z+,OCAP.!N?"K9I9I$)?Z^FRVO
PO?+PU[Y]CB$F$(^)>JZMYFXJ2E]-=M@*A@FXP5QZ8AL?03R7.A6 HQJ+K*,*)G6C
P+P+Y)^2XJL[Q=HJ!;(FW$KY9A:,M)6 ;00V%HBH?!*XD\*T4P2B+_G2&Y,=7ALSE
PHBX4ZROKQPR@?<'O!Q2'?@?8%A$[%-((,!=-&,07&U-[HGXQ6Z0QP0"VP-7HW>/W
P6K%>:=[??P&KL"OQ]-'_<1L1X+5HXBUQ7B5V6N<IMJ,B@Y">7[)Z=;;3N3W1UF_.
PO,A+QAS^*75G$9<X13O1X;GGH&/[??!TSN_$MP+/5]!O=_^2.XEGJ[C-O*JSQ?K*
P'V*4Z_ZL/$G ^SS"F(.A=4REML6F9$YK$5RK#GGDZ'729A[HCK?3T]06/TZDU'C*
PEB"--T%.HF.1LH<$W^'2")B*^F$[O_Z85)#''3"/':W6\-O%/!0_@Z3U0N.NXH:/
P];CAA#1WE&&H\$M:<AWJ.NVBS24)4N.#9RO\ME8-V:D20B<O>,HTNN^M4.!OVS]:
PQ>^U> 6Y"=1?>>>'S.C Y?7(&.26*VG]__T/R9^*,1$.L?NB2A_?;=B8@7!KL\R5
PA>KUTH^D[W:8<&YM^M$Z+&8&FRT\<!CJ%9&&BY9#NM>"*RLIRLZ\3[05+45S6VOG
PO2$],J7@[RQ-=-I2/Q[4@6+DX#>7,R34,51U&B+T2H_U%Y,A8"6:/&71^"9X$3<<
PX"B.ZQ1&X]4*,M^0_W8V%;3@?;2?J+\NOL4LP82]'=>]8\/&/QZY[)#9HZ@%.H]9
P=[OS$F21O#OBC.-]BT5Y=',3=E/"INA%^K@3HJ1O,\UL1E[OE3[<O6C!B1I42B=U
P3A[H0/;.1\IFV $YC[ZS@>ZTIISU4V9Q':T0<<-*A9^2M[Y/9.C2','PO,4-?"E+
P6B<U%M=DQ<[! A@Z87XX92:$^5S&6\_@_09[*'U[502WX[=J V6&CE%USVL^GLG2
PKJOR9&^#6W/4VB,D:7@])'Z45$VZ8Z6Q-J(P[73)C#K_(@HPQF:0S_3%LUR$L5:U
P^"7Q08PS:]78K4=$,P_6"]J/17*4]6ED>^EW*E154-+$NF(<2HR<*X<R>,UW)Z5=
P4@H.3%$R(/=Y028U0HK8,;FL]^JDT)S0*<TKPIXC.O;)NY6L6=,,R"!>371%^F8_
PGH=?;-GQYX(/=$@81(M"'K*;L$?]/A.2'?Y5G^%NHP#$NIJ4;<:,CGW=TW<FN!OT
PS?]61("M^T<P5E2G=)LAEXOGG96)*6*T@S,;\X!\0EOXY!]A7.[1E)>7%0'LUQX(
P89V;5'[-$\<W6U@Q.__F[+PD3+P[8!]GDUG]3NKA=+W1Q-;*5'HGU&(WS)PV0D: 
P-\W_A6CC;B1)WWU- 4V8NJG7R>432UF!6#=]%.*ER$WG,+F(?/92I\H7FMAYP6S+
PIE4:AR.YV-S'DF%FX7%0JH:>;<F7:@4A4ZTJD[Q+LH^6OV@),X# "O]?^A/7842?
P%D"2YF8*^^9UZ_UP4FF ;-Y"0U:470(QDR'BQNKI4GI2A+_"YFC'EPR>+.&X,!V4
P%Z-" 8<F>Z>K7G?76,EF(Y&!'5\&$\%;9*W,""MZ-,EVG*ZP0DDT/\MT0,ET^-[D
P&O$8X9U8_:'A=BS#JK5(!5JZ"LR_KUEM+;_(KILF0=[Q[.BTI# ZUZR[5^\XT=87
P95E\)V;ID\Z_%%TRMBU*?'3VZ)2%Y+7^Z8E<IF7%NGEJ$#:\Z^85G]+/694597!M
PA](Y/ A@M%G7?/MT7\N:LN_%?TOQH^IQRSU:/+0#55L(G^G_ Q>:/YS&IZO[Z7C]
PDJ-?WT?JK.!<OFS%\[5:B:]"Q1UB#A5V*]!(LN*TU4,IA<%_70XBQ3(I8$BQOQQ$
PB;?<9&SN)]#@S/K^&\1.:C*(.?^@Y4X,!])'[W=IOX?Z+@;@R=BL']BC/69!Q6-M
P=,Y,V_>5,81LCO#+>[,M8B4B)+XE>*B_?1VSQ1".T)V>-KE'];B*/F^-HJ9U?/+P
P.H])<_I =V[K)DE8SDCC;>$N\QID)J0AO* _^+(YF:JWX,]=QN)7O6Q\A:@YLW<B
P NU=H2+<['HU414T+GM(X0*VITIVE,1:_2&K>.$-07K@AAM;SA2V=KIW67O?1MCG
P8-I[/_S&V9CSW@).OKC^11YEUP1^G04(A1^)MURFL$F]9F)EB>2IN.,41[K$DB$/
P45[ZUA(2.7_?M7.RS5"ZG _X#0%AV:7.<K'.%S&1]\:O<MYDVP)<1.VTZL>B/ 4R
P"N]C*:URX6 7\'7'H7--F9&VQ*_E&^Y;$TPJX5:,Q&*NJL]\-[<W^XO6N!]=V\RD
PV IX_5H1;'Z(S[=MTE:63N,ME^A?(]6<IN+10R_\%*Q#=?<5 3T91P#\HCJ*#CK=
PE/XG*&OVA(/'&.#VT'UK>3B_B*)6Y]8&'<S^H5B<G+LK^=V!Q2VJF^%>15.>]2T[
PF:M'OK_&_P8,NJN\05_'=8;/F*:1C<,*5RNI\ #H0BU'0^J S>RKE\C< RXL8/E<
P!\BR-!U"Z$FT4>#H [QR1%^ I=?1XX84(@O[VI0]'B#(5]R: !RU#>B_0'0/A0D7
P_@]T@ZO_3F01DJ*-A_KH 7T?W*$$&4C5]&-6:B>C.^(7JXFF,&:?-?&W]93?FL0A
P4"D="ZF;N,/=Q7O>8I_33A[@ 4_I* $;53C8ZLU1T2.:4E5OR3DXXQ0B]:K<!*4S
P"&S@RZ]_.5G; H0N;S_%?AV4D@:0 "L]?2(O=UD9]NQ=HBP&\$%I7VPBL4T=?%@F
P?U<M,7'-FJ(#<?5):%8MV"Y(O-7]TM4^UUX^;N@C&'T=NL[O0$UV"94DJ[%'!<+Q
PBF-:3D5?TLSPSJW0\!S<=JC2:XST"JKHR.W.3J:IU3#"!'D_%Q!?[80]Q0@))RO2
P[!JRJ/J$F@\D; 7[M3YT523:CS^$PWK_M%LJX6_T$ZSOR@"A)5NRN:D:1_1ZGT_I
P ^TAN)\_&:%V@ST--98K;:\RZK!ZU6@:8-;>#X'C 2K5A_/51 XW?MC]HI%IJJI;
P#8E.#54'U71O*<=EDWI3!G#WL$0XSUY]!DT\F!VRTS%P/6O-JV]A4#."! 27KBH<
P[5;&E\.,=&7T3KN?* BEO\99,#=&/3&0P4F3CKN5Y*+<JB.X^L!@TRR#M@MH2.N@
PXZJ:U;^J=+GG1?[$)AS+ZK?Q!\.22"(&O\M,'%7-TU#+/OZW>%8G1N:X"4J$.BT_
P[-^#.7(72_(GPOU8H:YQLU#WG//5]@22MRHS+%;%7")V'N\2@E;7L#GTGE\O5-/(
P>SXUPGH0L[RH./;;>.\K;]F.!/E7+H-]$B=GYJ7J\!!.1SX^6-[L#_JN#OD1,'7I
PH1$F#6C0[@J[/QB?RI#57-&%9L>1QCC@D0HP5_NCY.N:[RY4]Y%JJ?(BY6DIZ>O;
PG6<=R\HLQ#>]U&)D/8+"G,QA*?E[&@1(J(1."+C4GL\FMKX6C"_Y\+F2WV\QH-D/
PMYGI,Y&W7JE.3M3$6..RUU;=,2%D" U+4>#@K.^>C.Q^=P+*9.O;?%<[1/-_Y0_U
PG<1TDO=LD_32$E-!_J,+U'>(GC84$0BS58J]R3JHX;LB&# 4-S*<<'^>GXNZAX\W
PR/VES69)D!*.C"???[-E1'WT-Y.1,[Y1,G[\CJ(6?11!_F_]N 5""M%-!FB"S G7
PPW5)(-"D%)4IAF[MI*^_1N Y,(A M3VL<.,@^+-B*/88;;@[89Z1\8SGXE KPLYO
PH7M^,49/NZPK\QE'H59N6@:_V6-2OZQK.N;0K/5)R=F!-24EB"T'FW[-QN5$AK^6
PNJ\(P#\H9$5._,=9=+0VG 5*'W-==\=3'>]'$^$)DM]J38L/&M%N]K['LZ=;:8.4
P>6 *G@$%[L=T:A5Y;&R]O6LZ1*&N]3;I_'^\($;Q5]78X!G$B@[A.U+-2R$2S3D!
P.>"*/VZ,\CD-^TFM/\IW*?F2ZJ@9^,ZZ@]J<2ZK.^>YH71V03T#?9BW>$%:O^ W5
P)<((/7#% > 2OV0+LM*$=(GQ(B=TLB\5E:M*^T")Y90A 8:MLD5C#A@)XK9Q#33_
P&FS49Z8@IKHMG#?3&V4-[Z!O3YT<01C6<'/8%)7&2?8L^31CTR/?,@0AB7R&CNQ+
PMQLTNR]H W6]9>A!490PO%,\)"%JMQ8/F&(8:[R<YP658^P7",:C'+;RMLVS_P<]
PVH3*]M#57!RN&1GR/X(J%J'>:*3C0#B;7J8<9Y/^L9&>K'!_"&5;DU!ZE_ _##/M
P:AL[08+6_ZOADU25&5B,>-3PAILB)4:CG *R7!T0!>;5!W>#:**NM%9]KT=[$YY$
P!KB4/B+H*.+A/T^&E9Z/\&W-[QMX.CTC.J%PO=QS[H DPG@V4G_0(\$L9GO0.VF\
P50\5_2JNEZK?H])&CSG/.3QC"A$*/&2S@>,(=DAD0(1L@0OH!FCGCPB7S22HF8TB
P"&S'T65=JCV/\:6X?P"GXNNZ6K#HW=88TA)'=SVC:GV&JA-]S3$J>U&*:JP QN_U
PX-G!/LYR5?T$SH$_P/ZS<X<JC7T'!4 EB)L1M)J\$[CI!638]M@O!'MGO#URK[?5
P_G)[@6%<"C@,?EYW$;0,TC+55X\-6>QY)<T;(*&EW[_BDO[EMIQQBA;&GY2L6S4Z
POM?B1#_\<-_4PRGV<X1E;82J4SSN:_:,1<$Y$L$8_HQ7PZ5U']'Q)\84S$+M<J,!
PU23'#2Q**S>3 U'P-./-T4YL4ONFY[HN(99%;_KWSSGMMV/9\=1$W";?W-,KI9$5
P']>"1ML=."13C6D*EO.1CW?.Y'%!FOJ/3S0O%R/X)<0PYMC9?MSGDF8 "ZD(JGA[
PQYT G#+F^^BL91$B,$U#KQWROM&VT?W(AAN#,XKP+;Z0?\O"CEH]Y?A=U*/>G$5^
PQ7;I*<O?">7$H]OF5#.=Z6AWWR:I.W4><*JY_CUW4D_\+^UV^\/"DB'1!: PW1.^
PJTR<1S;]S"$\X($W/T[-=S(?-CRN@J*H3+PSY JLJBWTZ*/OP]?P/:H0>%N.8A0(
P_:I]F@5-9LU[@^,835-U$*7&ME5:=?_B@SU+>6Z-AAM/60 MR#?5L%[T2_C*FWA2
PQ"X'929J@&!,Q(QLM(9 5O5:E^<7GP9&L);!A\GL?^)H[F'G6Q '%?S45($=;@1[
PEDQJX;(+>@\81/$%G,A(Y'BGIO";*'R>+#,[#J[NAZZSVE[&$<U9P(%,Z%D2'GTX
P_BA]'[Q@*%LMQU.L&[2CKF/@88P9YN33&WNFVK]]OA+YLE"/5$"@&9DY F1HYU='
P>.UL+X[-QTM/R[#DZM:$$ \J BTCAN!UGCEBCQ8K$D%8=A]T'IG5PO,M4X"ZU1:G
PA*7-\PQB,T/L/B*\LZA^W/MU$45]M0X&OU&M06ME5./?HN!=43;-2V4J=I%T??.Y
P.SQ$R[HE<XTQ](Z5],NO[?*L/G(Z 0H@<S$8:PFW)5/9'%!)!"KM*2Q+JJ]I3EUG
PE" ";NEL76MW9(,]W.6%I"6*\$_$YN>Z8O*GI(%L2=IP^K;S4OO5L]'M-)IW=8WE
P)"'=7>V8FZ/FQEMU=F/DZ\N/8/4WG38>XC^3"\$(WH4,8FQ_M#9 L'8Q.F GK<KN
PXM777KCMW]@C>7]^H3DV%">$_@2]BL=>S!3<-L7'?V"V+G TNY^^S-Y_ROQ5=78E
P6@.(=&@(UU[A464M(+H5/@)N 1?!Y>I@']@B)3!>^VIZ%2SF9F[F!:YDD]T9.^[Q
PGS$3]-GI@C@F^6]D_^;WMM#>:+#U:K,L_#MMCU751KT:"#DQ]+CKFYE"SR+MJN-D
PF%P@2LIY&H'FEV,_)A^DE$AW9+"-#&1,&^:JA=OS#JQ"ND@ 3%,^83 2H:]:ZWPC
P9X[W1/-_NM$?MW%J86DA9<41Z-(6-]<$B!X6-LE>KB M2OIWE,@0BD!G8MQ; F.4
P,(3=W JX(K%U6TI&MEA&GI7]Q]SER?>)6,BF<H2<L'J=CN.8*?R[2(V*7SG1APLU
P-4JZ"!0R-N83?LKCPAU.:P@D7H_=,U/!XZY/"53?^&HRU' ]LH!Y%R+B1^W%53-Y
P,<03U_:!E+')%V^V\H0G2035Z*13" GR;H9C;?(=5<1<&+F^Y"<MPIIC\,A__K8$
P:UU?@+2-=R?I.LM8 T#U$]V".N.["(<5X'MEIHQ8QH(IT;.@/9NQPX+Q05UJIW8N
P0^*5RXM) G_"I.P_N[#<4\IZI00LYA;!X=) !YW(HH0NSSQ#%^C:"L2'9N7#?2)@
POWBDW*S<EM'S9P4PH\0 (ECR%Z0',]J.O<<;Y]P&BOV+Q)5!!1=T[$@UB8 I(X /
PH_6"!\%.-U-VS=&3V( F]"K02Q9K9W'9-XI2._+HPD45/\I#L#IFW-[:_%TZ*<.A
PYO!\P> -^[HBC=THO.DCL_M.!L_ZQLUI?!9<C+[=<*FB12_1EY^@:EA=GFYS)M6.
P6:H&T5IY:D/4%W46[&>4@-LU9?9:,7-$L$'XD^6@/H+0]-8XA\X8&9-=SEK1@7H[
P<KJ(>'G\U_"L=J?\:BJN,H?3J_,+.2DDVA=<OAH:\I+GOMEB,_+*F$TU_5S_>WGT
P+A\8\3K'Y>\C/6:5C#+>XCWDBR"+H%;V=;#\9@L@*+'U?ODX'Q)(B QS6;A$!=-,
P"*/EMK(@PGQ?"*1TV(X>#<<K2OZ0U8E%^XVV*-";J/VDI=)\@UA5=#S!&MS17^ I
PB6*JH<"X)WU>BGP!'C^K9FD^!#]'*HM[\3IBL7V3D]CH-O\,RJ4=MADHE<%NJ7_%
P]MTSDLAWTW*2IKS@4MF'Y17FJ3M8?RSD& @09"^CGS+SM7/=KS$(T(VY$H<O$Y)I
P(S&'/>L01AS#J!I8E^'N(<9.R?1L0;B&WOYB'O<'Q]_U!?\ R3U7$ <CW%^N_@1S
P9R>,LP0HGGPPPRJY?6(@CL#_0F>\[IL&EE)7@][N?T1 MJK[ *T2]:I]B#\QO-%L
P/OI(U7=M1$!H[7S7+G1+I8N[UI"V1:#LDG@;J)?+(DMA_RZ_ ;W<[\"&QC(C.ST\
P=ZYS(L_XZ,OZJ>5$OBA%M-HPJ/G\"2]4SX+)1HCY5?Y4_./Y$<W#E B3Z1GJDSVD
P+?&#I-5BR#G-L&C%LD745BWE)"1^1\XA*7GH"?/V?I064#H08S2W]P$989H'WPD 
P983F PGZJC+JYR)**%-/$NIA5P(ABAQ/#24DSA#0-'TK-*#7DL\@/M#$BN6'6^?V
PN5JN12"K?2+F%O*1SC%E>HC,/A#12]+]"8[+@2S&]1KXT9(49QXCRCF%"AE9#:+?
P\'Q0X\W4T;GAA.2+IL265:2!V)Y*<^VF_]DAW+(1Y ?G\>Y_3/[J:W9._UONK-#:
P6F ]Y05B+-W5H(I =YM1%06D=4])%YET!8,;M1""](O?'[Y3*ZQ6C0=/\R4)64A2
P%W%/3/WO>RRM*;:#?A[GF\8,_J%<="I $[):F(L:)(,*F&L[KXUTVS]8<9%+ @$R
P@^A7=QR)NK5#/L0&,(O,^O(V.+XGV@!$\[77K,=J".5ES4GJ-?V5<MMB@IM*)>BZ
P.^H:36S?W$9B\>-?+EWG-^%0O>IO@@B>/SWP1^RE6,D0;@K02D12FU\]C4^2+PDS
P$O-N-H:T_(>42%<CK>X>3K'BL__I#RA2$$FCRVS953<[8/]*_TP&,[[HZ;=;1)9<
P/YFD.<:VHV_!DY3L>,Y<P>O>#.4=O(S=7SGT8( ZFG#2N$$BHC3T2]HJVT1%:U1D
P8CBSI?QN]D<L-T[$BSR?$M$=<F@X VXBR#.H!_YC,8@P)&PV2M+[CJ<'P"LD6H(.
PZ7?08?.[A/RJAV&4^P-A-K5'!<AJ,9+]LPL1WD@]<M]R*O0W=NB5W_$2@W\QBQ)#
P*!8/!.OF@$[X&:#Z=.BR;C2K*RL%R=MH;T=&WW<QY =NK;J,><%M37E=HT?6C/;'
P!U":4)BDL\/1TD%,%S7OTZG*>3A<E9\L=#%OQTQ*&YVDD_BT76*V5B02P08_A];2
P%V4_(N#SL8;+D3JWGI+0CFZYH-=CRE^2)L(IUGM8*K1[5 /$<;K'CW0&=&D*F/^&
PR_ &DM[-('XKI^'C%"F[6&]D0FJP@2-2SYFJY-O%X,;%C8OP65WWN:%?UHM3VGH:
P $^$;Y+/C C+9(5I"^%_"=S)%"\5?<!7!9V)@V]7JUT;45/]9Z.)H Z6^ #TK% /
P$<4:RY"B&BI45.# :D.$-T:8%MUDB6MKSC]L-+>B=WT$&B'>6\V,7:F@&!&2HR?O
PPL9E!B-/I^;Z7/!V5>D$V%[9 &2-0P&>Q51N4DI3&HJ!?!]X(G.H<AR=EC(H'UO8
P$R^4[KAD9A( F\UXB()T7L@4-/?AFD+S)LOKII<4QWPN$8FVO#AYR_L(@/P3MZZ8
PTK?H%HOEH'0QM[H3S+54% P$,K4M8/\"(+E3#?8LE#G/:[?31CUO9H;_ODU?IW,,
P "T^!+K\F[8-0 /@]".2&'@,L-4%#8/.IM"'+)]7BY8/ 56+<//SG#4KOJV-R:&8
PK8ASDM=Y'O> FR6OW#$1NT@K-I//)<5Y9$:_7E9EN1]@CBC<;>.2^<X?5.I%:4><
P1R)Q*SV4=Y4ZD%V>#+'2NLQ"=P6ICTOV^-3]Y#OY%)C353)(*G<W'_1IO6SM@U/;
P>B<C(IBF6'%#L* \'/0VL<>^;P&WV&H6-NX$QF2J:7V>N";Q*"A@$S6_J&BH![>,
PJ/H[C3FP]%=X+)K:_(S/V>BC="'S2P/-H#V.;V!QKF#EF.Z1UQW.>[]( VXZA0RA
P$]/?4 P>A0 "P28RNG$@[*TKS9L$?-SO UAI?P<]>1^D HDY2(NX$-Q?.ZMFC*[X
P%%7>H9X&4']>'3'Q$R22S,APYG'F\I8$FGXW.%H?=V*"NF'31XU"J7 (M#ZJF=<X
P&$AE?1H2"D./6++7W9)?EGN2L*H0L[NKQL- =-ZV=4M]@[I8R(F6J"%4OZS*)3-7
P07X-G!>=?)+,9<M#PVN-OLA\^61=D99J]U;WBNX>2>*FSGN-Y7R(7=M_.MY?_=-C
PK+I,C"!OYN<$H=H0Q.2=53!;P8,Y4O^U6%2!BI-65$C) _C)"#;+P-H;Q&$5DLC^
PPI7KW!BP=^K$#0#;1 T$AB+1ZG?F.]U+-C-D)QHAM5Z>EOB+D!/3W3 0U$)08'$G
P];,OVT60C#"9N:<W7W4C=: B476 P^7FYC=GD_^JW7,1R=<A^A+](>^DJ;0SO8I:
P.PIR4*9^NK;,4PY,=Y AD@%L^'+#WVK+Z)/_76)1*QXUN]L[,X2ON;8TC\BCFC5X
P(N<4R["RDKE"/<(=-^[AT1<FX/K]=,&NN^*2XM8ZXAA4H_'=YJ+='691"MR(NZA=
P.\?E0#[J]79[5W1N&]P^Y-0_.2C;,4/!G2C[[\M XJ^Q,K&Y9NOY!2L1O'O/%GG'
PK!M';)AN[AAN6 25E#X\+R&95<SJ66Y<KXJK3;FKN.NEA86-5QG, 4Z!)G;8'H,H
PQ^+QZZ71C9HPE=;-\)70<F9?.4X^NJ7;[KX2.8N&"#<W#0N<1Q 6N$_V:&HL:ES 
P9%:Y\8)T-B22I/22XQ*#M+'F)B,\)0,M;2+3M7F\U+>2E>,><@70GQT9$^6 U8PQ
PAFJ3L/>?.X&L<[YX"@S-\DOA%%:&" :*HPID.W3!T4-;IO*O&?[YKF<^9J5@;N:/
P?(A:X=5#S%]*AYP[6QA['(;&X-IV,FO9=HO9)BQ)$E:H1EX'U90C#*HPZ%ITI[Z)
PG*4#.V)NOWQY<V%9'FQO'ALMBOBR',OZCDQ\]B^<<J9A9X%&I38?@WU58]YKX:?U
P%P;=6NE#"7%"45[+OE@"_1S8__%DS"^2G2NJ,1O8BA<M4D>;\"9P&(0J;)<RTWB?
P"(6>&;T8N8CNCL]\8)AB60V;\,'=Q6-<!#SS;:LV3PP80NSFOH]QT1,S)'9. O:[
PYSK4M/*\97&%T,B;5[KE40Q(,6"MOLB(-SG(" SQQQ4,"0.$4>&&:[W$#J_NQCTY
P:^<XJ7)A U]7^UQ15&7_I23<P8>8X?%='D%%X04S30+NT5<(>&NR!0R4.*B'<?, 
P7) 8MSJJP**W]=I;S2<'!&#G#].S1P#5=UA:KSO@N]Q+">%?<XC&T)R8$K?K=J&=
P8ID"<ZMJ;HV@/ K,3!=%:M?7'5&\KV5\1:8XW!J Y)K)[,T#8]-^.(8IDOH$@H\>
PB['5<39J(T?9\.9!<N>FX&NL@_CN1:6/D]MI@'^$N?1 QGMBRFL3?^/$@:(MY60!
PN64-#M&D<79^5FV,/M8#MNE<*'SZ!^HJ >:^@E"3RN1RMK2!]H%0:I4"* 8Z8-(9
PWW&KV=-2 MK"]!YN$)$KEV?Q*$%J7/XL7I!I[8:)RF9_+!S]@DY# PK5P>H1#STU
PG?P2M*GPAT/Q-=R1)7./\(2ME4.*:MBO (: %HBZ[92X&QL5,&Z9)1]RRSCT-B;_
P<;4]:_.HN'L+U4V+I"Q-)PMTH>F;[&.--WD>^<?"<.:\.0G9"F?=3]R"EYD5=5KU
P<0\S=13@'CM9."#9#H?&0QSKRSNTXF8;:\3#;T:M3N">-)EP>H.G/2J;+U>0G=WX
PR5*\3_#.B&!;1BZU*MBNKDZ(XN0E"ZPP=%)=2#@POQ,+2USG6,5)K!'Z8M94PM<E
PY>Y(V*..WULLDL4R1V?GGU&\4WS[J' :Q)]Y2<>W8B+6$5[SUVIU-@/"='/@*7FN
PK-68<,I0;#=^K^\E]ZB<(%=6/JFJC_1DO]L9[KSGYX>8>T$8\PAQC^$WU;[>\?6.
P3%H "_W7WPAKZ/ICN^?WN-^X7 > *5>[DM6DN1AY&\?*E@B7JX8;/M;.$F<HY,&&
P\U.+R:WL![,MCX>ND*&WKR:X04/V?X)\$8L/X7EP@\?R9QVD_LXV5?<,A7Q=)Z\,
P/9WPMWL74P@_78>EE.%N,ZFP&O:NZ2/DQV0*UZ\/FI)FBZ7L9P'TR0D'HYS!,K7[
P U#3"/;[HA3EC_A6F)N(X>\856R:I0KK,E2HO#(/Q@BC2>\AJI!/^;[OE$8R)4[<
PX*<__T3Y83J=)P+?HX%FC.YT2Y$,L[8_)1IV =P?[!906NL1#"_/"LV%UUNE??;.
P%>EBH^\0YA];IU@EC*<@Q)AEWL9 0'-G7M=S ^?8^G^G?X%D>K.L* 4_&(0O^)S%
P!13F[PG^*N'D4,M.9YXHHX1*@]BR3EVT['S"6N?ML;$-T9 Y)W4!]Z6H,!'MNK]#
P4'/K%S^P",'!W)07!R*61GL"9A>WBLN<Q@1AX$=HGLPP!"RV2_W(P9$!L'/>K*2S
PM\],Q>I0PSXL1N*WH+$PF7/WAY'[YV31E1GWBO$_4=U&#*H>";A%WJO24T4/D>8;
PP"%XGL^Y*/WK/=?*V%6>Y749[-E9-,0H&+I[!G@$)2.WHAJ,%H<#P75D(D'GE@%A
PV5^T1M@QG.P;);5VTVG8_!^C-)Q*H]@ +352]/&JN0B81*\F0(T3'GP=1R7<9J37
PCN@=[A]];PN..UO@V$A\R&FMGKM'7\V;'C"I5JV<'E*,FT20\(-5QK3HC+ZSC&99
P0F;R^[/CC9?)/%*%"[*.@SH#N-< F^NB[%.C] EK[4MQ(2<5E:J['\5Y)C7"8.EH
PQ2K$4)D\^AT Y\9_:P0%$9ZIVOE :!A7KHXDQ^\6MV7.8])9:5:21BJGK7@0#4HW
P\-_<R7_K0XI__W_!W=X['L@.^?)\D59U]L6X_1RYTH?2S>Y42"(]SWA0:_;]U_N@
P8@ZGCS]K5U%%+"$#FT IZ3#\W^?=#.<TJ"U_JTVYW5J'VZ$*1PI26T-@-!ZH+<E"
PQD\8X:&.A)^S\S7OX0.=%W)8_^;%8E]X=%(;[A8DIB/Z("ZW_ =@6^,!6>,*?!1Y
P7Q% 660E[!I%TF*9PTI,.QJX_:%2>3''&V9DK^FQA_DW.ZO)HKIJ96P6P,:]:PUC
PV=4:_[GE3=1,LF0=_\6,=.5G3!,\P*Y&[4-:SC;TB4E317D#< 4!WY[.*"_V9ZBD
PDH,'DOAE@.M(%>N+3"'I3 'BH8H9&L[78>;U=E/Y=(T>X!%1P2/F.#NE=Y6@"::4
PF'LKB Q:\==<'N#3!G#4:.'EVH]8)<&[+C,$6.%PW2CNB.-.+RU^5T#DGKN9KX-W
P-]2BF[&<&V*[FAGOLK:BRYCK3MIB_3Y4Y,5B5SCE?_/TAZ!OY4Q6X 86>5P,IJ&$
P%24U%_A3@;F&@6/OY2&$U$0>QU4BM. VKUP%CB_ ]71SF#":U%D'9+1%70(0;[S1
PA-F2_"(9!T.OXV%^/-6;[^!^RYB:.LU. IOO,V7_[9@Q<\[NW47M"XA";G"(\R=.
P!1AE2@*_?58S(F&3'(B)VHZ^0VWDGG;210GR^6V2[R%L3@EM\LWF5GP5^?#D7-MM
P33@!>C&9_520:,#[P"H-"=3_/ZF.5UP:JR"#<"SNY@?AKZ'<V26H,T'*H8R'L!GH
PB06X^Q+:V$Y-N[DW(?%6M27J)4+X\<0R::$OL(1HMHJ 3X[*/8,9;J-2-^],'F@ 
PP!S6 TQ!K=TL*.3*H$;I!2^*66Z,[E_$MM) )42&D#5UGQXE;I A_SKM8E\W^"_:
P5<\-JFD^&1?TA-*A:8=\[ @'EPO-22EWFA P=9#HJ3]T;#DZ2T.SD=EOOF1RAN!F
P+U/3".R1KR7=+? GF)^SFTRD,4*0;2[*B$.3FJ2>VI8UEW[I2*F/26F ,+UY?QI[
PS>0EU8&&W8-SP6^EF^/7W\K\'</[N!'>3*L>,#Q[-T =KBAO>>DHBI:]FA]<W.T+
P9E[V(E_$OLLA1-<"U2>//#MX_WP9.S\PHCW^6<REBVQ2%K;\-5\9D F^G7BU]7? 
P7JEP3U?F:O5I$>/F597P>6!*%T\> Y,F0)IPG5!?CW(XQ\L30D$0BY=@1[I._7;B
P+![UB)LZ9L6C5Z_)RX= :W[O$"68(Q)IUI"'D+(\?K>;\UTST%VR&GC(2WPV9_$(
P(Q7YA/U.NW2R-T1H;C,-![?.A@OBT3\UYA "IU_@&=)TP;O8R0(GQ?2CP$'LW,"R
P%5ET'K--TX:'8BST0"]280RI&M0Y&Y<$)9A:Z33^LMCI<<GH,%#=3=H/%0^"I[R$
P49<\!7D]6X-VPHKKK0,9%#0" ':>VO2X6:REL.A7)2L"3EB]4Z;\=!/5?8MO9#9I
P2U83>L*TV['IIXZL(V:_)_IYKG-^81?RQK3\:E=.T3FK)7C6LNZ *Q^589R#S3@&
P+]D6,\&!I&!7.8OQS7.6[B]<O:U2<R@26*BB$W13GVH$<!'E"LB_/SO,F].G$]07
PJ;PDW^TX33M/!H!3(8=S]U)I71F/=V?^C^EOB-G@%Y%NL%&&D5-"EIBGC2CC"PS\
P836V\.V)\A1Q+2;(>WRZYHG@O:[LK+)]$D%DKJKRO3U^.O_,9,!P(!95)91Y?_-]
P[LH [)$DOR>TPKJO+^M<G+L< OH>6@4D6S6[7(FY,W=A6G6GSW7+[B0KWA__L!:J
PAME-=%HRXNBK<6W"MITZSDP>1DT9*HZW\G"LE)2V"WG<*[X;Z2U9<DI1+P.M2)IH
PCHFDU?:^_#)$$6FI#SGM&QASSUZ&"U.#D&.V%@'>,'^/9SA'2\\B)$0I7!);SM.:
P;;6#"O>XU>EC=RU0]CUE:1@*3\UNU7O7"G=E[;UP#J:SB)\3SG)NX<?,P!T<Q;_W
P3,ZI(T )]1+U*.[^S1X2T>%B-LLL.OH;4<2/6/=;\,;I(%T=R9<6SA4+O4KL?[$[
P\?K;5 ]=!^B+"\1U;=ZBQ[N1,\OI%KJU:FI]LED*+V4<-&6J?"V1I#3S,;;3F*1\
PT5Q5=0ZB@*SH4.WPOHLBH@+B+^.Z4@:;!@4A[:S07'W 2.]4XX3-:\@%M(A96N5'
P$IX>G?$)B,#^7_ *"&^=-P!J#5S//_,3*SE(E&J3/P:OH4[< SL(H*@ 9!&9'X?'
PH/+[?WAK;C;1F*2T$7J1I2Y1<VK7+!" 5X29D@9$IL1I@?^@HJ.V2A4W0VRF(EIK
PK@(&D97UA*[M:8+-AISB@-7&H4R(XRIN0WW4QC4G 9@G+14$9Y#T;*.\?<HA]+1/
PEMCJ52%8=Q,2OS#O:P>VSU69(5?KZ66A3TX9+GLIB;,@G;%D;*NRIJIY1[N\D(; 
P'I3VM.O#7(G!G[^_%]&;_B5HEO$*SDMY<3TN5*QK=8.=/N^U]-</\],?3MR!;['<
P]Y_P4,I(*.QG&AA FT6H!&%\G)\@DH.R,R*A[);"F!9VT^3%N3C2RQ/!J,W*+(*9
PE:]3IE:<8JWZK2TC'E&0+5 3A%55RX"GDA$,AX(YGTHVWQA9:>WJ9KQ,, (+?M##
P",AMFMV1 <%403QB'OD-:%O6 O:JJ-=C'+K'\3*ZNP/2]WV:D9ZN-/8I'UM@=)LK
P"-01NXRL3\E8GN&R41\@&SG/*VE+HR[G2Z6ZC<_$?1B1ZZ5UF/)^E19BJY1,<EAF
PKRQ5/:PX8?B',S"Z\+DW !/F44H(W#2.%9D3[*,8-.2"RBDH/7&@$(4" XL%P6+G
PV-U?G0;K.KD/65;86I+8=(<%+T#\#LK9D9HFY&1:QF@0&OJEA@^R377,(R\.DP(\
P1>$I51R%\TTF;/'C<<60HQI1XTH;0V2%/>AVE!%/N&[& 5GP RB.*;4C,<OH)4H3
P,R^7_+7)$-U8W+BN7<\FL74F:;$9)\;U9Y>4QW9;L\3UDEWRB<5HP\E_A)7#H%=)
PC0W5;VWV"R'9"7-9"".+1I+.\5KN:D#;'2?;[KO$E&TA;SZ/J!4[\T.$A,+HM@=Y
PH31[U7>_I$)(6.UB]#F\^G'!*9'_]0:5\4#LACK3L4"V7>L^/.O!\3->DI%^@-H:
P!#8%9$@:S"+9::Q$/ &3UZ59:$B7H<DSN\*OEJC2H8; A0TJ PI8HPDAU_4H_MV5
P%P3_?#9?4'P.)J!'6I?,@07?H%I5+P^DQQX/3AG9$<WON.T,;:WJ3V'U")2^_(5!
P"+I5J%()PA"-P.A$LVA,@VJ4?,R)):1')H:?7>/$W:=^ ;$!>W1"_&Q/U;KAYNJ5
PHG%NVIY@,!"%@\IDY"$3]'40$+XZV#BD />BU-#B<TN,?#1%E)<5U\ZF^+82O6TB
PED"I1,+5-Y%K8'4B]Y73DWNWQ&)0IJ8:D79QU)$P-=Z^?'OR=\PSO^"K-<E9\<( 
PV)XWLC7?_CS-V6\\NJ Z"9'0C7,X:I6(4ONVMK-VVC ;Q #,JK)!<]L.&S6+=9HK
P1 B+_P%0^88(:+.E>>;BZ='R%0[)S.D848^!AL\C_4JTR#^ ,,8O^;B4/J8(';K:
P5@6"9^L%YSZ9S:/>LQ\:Y0))"6$S^&B$2_'2:+=>Q@/SY]N(R?.GV%[)2FC\OEOP
PT[3A,F<2;FKX_\3H"_1F^<$H2K>!9#V"+'9=3APC^J>H$ZQ.).O .R))O\L]J!61
P8B^VSE[M(<H3V^2B5<#\O082&Y'NE%*D0>10L!^?N [>.Z_*9C#N.3V*KOCUJMKW
P61>G7(X^D&R1>!P> $%$(F^&&5M7Q9KY"CX6-8X(#Y":^9F<!#L718;/'Y?<;88#
P6C0A#C$GN2WP1-AX<^4+@],+Y*[\Q%:*#OEP=BV?X:BT-0< %RP#QZ,OL\R+U(0%
P7,- @:E=:(I]8$M.A,.*=B$R4907]!YDWS+:=D[V=^KZ?MD=>=%#.C\YOJ[?5KD)
P;T'3]B])UF%!P/E]S9RFK6M.T"!,HQRQZ'QSP F-HRRPFBY7$8VTJ&['9QB5&+<>
PU0'E"R%4I?.@F%]5%_$90MFA55/'GU];"4ZEQ )@TTVO]RZ-;<):'(YNHOEX(3X$
PR$S=W4=]/2%AHRF*S [<G41VZ44JB/3.;K=HK2:6QSN(@?5=%+^083=-]H#C1M*$
PK4?_P(]>+VF*?5/4K9YX^56M)[/ 5KAYN_ QF,MJJ[+.''C&U" #NNZ'5MQ!V5UH
PWOR#)1EA0]>!%\VAC2WX;9S2 W:?>6\ 0A3>-+AX939<(R1MRP<VR1P@VV?KRI6S
P3T92W_QDU/-#8N;T3CG5W'U<,)DH2$71W.21\)QCH#HM=E-^]N)XYT$/V65A]ST%
PT3MU$^3GY^];92F $\!^;\QU[$,^<;#AH(E$ :"/0)Z?Z+V.*;@C5F9Y[):B'WEO
PRGP:+\V(+_-1D*RP(?D4:8X$[!V+H#6J)0WO $=(EU!!8XZ\(,PRH<LI8UJM"[J5
P( )A49O275?PJHEJLVUCYY/JYH5IL\Z6!O:>BZX2KUKK/"&AZ.L[AI^3Z85R#,Q-
PK.X.[% SE'&EU^'-:6VB#J6,!1D1J#]V&WZ?X63_0PH7@!%MKV]O3*PB:#*7^M2E
P2X'CS5JG%%!U#U\<O%>^^[Y( XWL?44/HJO5?5E^\V;)'F(2A]*#(QA<ZZ_(H>KU
P1=%]C/LR(GMPK05N-)[Q/9%$^N783W'W\.,KQM!*?1^K+X-1&S@#3"R[=,=Q"&(G
P.&\M4P/2,WZH$=8.)P5K)C2S6S HY\=W%07BBOV8'FL3S"&?*VBZH]I[GINM7:R?
P(N, O!%Y4C;$''[CS2P1G& W1[*L%G=M<0CMB&93&QU6L#A_<*O6#7D!S+D9'O9X
P\C\9"X\B_+<5X,V;C'\"&8#[TSEB8Q:8!V'+72<$>I4^ICE0&?F>"O3/984;G4,E
P>P#VW"+P-2G9CLY#[>ST*-J D*\*PV&NPQZEYE/[S>W]@?@0@5.O^HB]8=^J3)K/
P6_I$!G>>H!\.;C3S+)VL^%G)$-"[M($J9*&+=V@]OR=IG>@+28<HL5VZF(:>!U>;
P7AB_&OW2JA6A714W]1F^\QALH^4NV8X@1Y7-V/JV6]O>3AO.._;3-A*O-QB+14/)
POT-9:K-V3&<GX"_2QAY@Q'A.U<<GS:S1W $5Z=O<\WP&.<H3)K0$&)+]5'2F:V<_
PJ@0TT\0*=YUJ@3=[!?5"0BI6O,'T["F$Y[.^'R.RB73O0JX#_(+#*:TQ>'<6IXMP
P>,=]>CX_E#Q4OA4L-ETSPJ$']BSG]$!^PS?0*TVSV?A#;=6BA_2*=AMO]6FP@;;H
P@_B_%_:6+7WCBOM[!?[PK@%![ 6,+7-11P5X.BS]+HM.)';_LO&7)F(%J2M!;>=]
P9^/#,I]5P>6DFO@?UD22WHCKH811DZ*KP#/M;YK?1+'=6Z?=&-%2T[(@/[E0;B;-
P#04T\0[6-)(PIPU)[:A'.UVV"@%_/F$)7-"^H;FNR1Z)B:Q%;LC8Q"OTP(>RGS:/
P]+HM,T[L(_,VQZB$Z=G&5CW#@I/G@)[FER%\5L'P<% K?9*8I$R2T>B\P5M$ DJ"
P)KLV)R"D!-!]T+4<2_:*V'-N#1196N(-+%PWAN%Z;]M?2QC[?HB!RZV]UVKR^3?<
P=Y)L"Z;R*IZ)><3:'C-E\I41?/HR:[4/7HN;*5,.PK^?!9_6#;;L_QAI[NGYSWEY
PH^Z 'D<U'ZE<;LE]Y%6TO1W?<Q3\^6=='=H8M,Y:C5M;Y*M-,?F+6N2C59<"DOFM
PO>ZP,3'.::1V(-_$(=T#"?AE#?V#UX^9HMV@ AW3ZK(#>QK0(2#B.%<8;I,-30$+
PB>&Q,;>PP22CYB>-BJK.AYSNKE%%C,%S!2#0&0J&IK9K>$W*U?$TLOB],!'0Q= <
PP\?CE]/>,\XJF$JD>A9V>IB7.*44NW*7DR;52LKQ#TJ)BM).5<H-.U 5,J#:K.,)
PW'G6\H&B"=Z5_ZD/%>SW#-0R&#[TR8?7ZX(P,X /4Z],XI\YB2,O2E^O>7RBWF[V
P\#?JTW=^*X[WDI#O8WN<I@@B-ZVH0!5W*<M#I4UTZ'2WJEJY.X[JZ4_GWV])/V;>
P!^O3^W[G2'*^CF"VE)_XS7=^GQ4E ]+0:ZBE\.0@VEA6#-6!^:="Z46*X%?)8B8D
PK@N!/&AA*&MX3_-I[=8">%SUO[5'8Q?6K?TP*$IS_.;90SMU[#_G^HTMHT$I&E9D
PD%V/-IA&! X*.63'&)R K\4G7F[ZD!+-\GS0Z']+@Z1(UJAYD^M%;W%E1&]53'(I
P2+M<_L=FRW3?Q_KDO9.)'CEG?E1GN"OT9<.]J3&7^UK.HIO*&\CSV9T\T"R;_",J
PHB"@E^)."D>\L(J!)J)TK8!.++O7N0I-%88W1?,^R^_5^)+S;1E)B$V>L63>LJK@
PF,@8,W\XYTBWP+70;\$5+GD3M5@=V#E3!,E%FT6,_E4\EZ>^$:BQ%[L1/IO6EG*"
P &__TH-WE??1DFOPT41+3U?H.GF1DXV-NNX/*R13+%#C8X?.I(4.R9F:WB:- S_+
P@Y:IT3)WCR(^B*M47O40#+,5+.5W!)C\L"Z@7GF@,QA.(; _1U!Z#7K2Q$*5+8U.
P\#B_[#+K&R*W3BP@X,OB1P(ENVE$N?R+S-"BP29_S  $)%->H% 4*Q*]'"9SUO3=
P?&8Q2J#E?%E/+HOI3V@Y;_&)5LH>AN$5+PUP[C#:?&8']$JL,K3GZJ!=-9,9O^R7
P3C'5%)U?;Y.Z";L6 BT4JS]E'((W_Q";:OHO?""B'07RC(\-C]CP,SL>QR;>T4&7
P8M+*Q3A=RVR/ 555Q*$)6NT1?-K8,_T!T>>8^=DR7;7Y/-:OE_8NV*D1-ENC\]TI
PH;N<?L9B=:$CT:HS1.AF%4Z HC0W1NFNCCD9O#.U7=MT72ZEDQ*2L%,)*6P V).,
PCW.5?7,X("3!4?E4ERTXH-7HC]5ZD 6.(OP58*WG<GS:L%1=A@Y,;F+>LGSRT1,_
P[C?J1Y,^R *-DH'7M4GB5;+4<C9X:8:QMXY&#WK:K2.>-OLFL%$BE2=C/??6MD?L
P[[%CD^ ?U%' E)*DW>W"&Y#^P4T*1,^.>P"!GP90XS,XL6V<8P.:]/47KFGV<:L)
PAU1\3OG^Z0(G@&=UW3.5$_C5,]EL=(3DJI :7U:O)XE'OUQ2=5./@1E=DF)^H]'$
PD:G1A&3,0Q6!C<GO7H@DL(@\24AWJRJ<'Z;/W'G-I7,HF\_V!#-:GRJ&[7UV4MFQ
P4[NCO\2N3"9;D2<-D684ZT]/#R%_$ZAQ6RQ>]S*FM$++V;RYN#<SW]8U7OC3!KJJ
P'HA2H0K)!Q.%H+?<_X4Q2+!OF/[UKH:BZ<HIGOUJ=&C1$/TX5,22U=UE'X:%38+A
P#]H!,:"#&$]$\M.!H55'#@"8%P^2)RVYYD]+T!*PT<?(\\X7#U43#58>B4T!N,MG
P&]COFX_A'F[H_GRGSRQ$O]#MT*?;_PYBHT% -06?E5EYFSU+*G@6A+QQKR@R-1P:
P(I+*=&O$R@(Y$OQ0HQ_\/Z:M!PIMS*Y(]^=H@8(L2O\D6#=G)JEH2 )G&XU,B2':
PL9@F%E-P3$*@XJ $"V@^R@J]R.Z'3*O@ELK.VQKG$.[DG,#;J]FA0#Y.[T;UNSE4
P?@?A,=#BD0Y1BP)M2YNV\7<F30UX,T/7!N,6CZ#!:< AXY1<8OFS\?3H?[B8?"$>
PP&=VB,5%E37H_T0NJ@$Q[,FS\=,_I5JEQ00%?_42(8 -VG<0ZRB>VL <W'+D9>F 
P\. 6N-*YRE", ,(R1K>$<@NDVF'; /A!TX=*BW!/'U#V=9_R%8OW*]V+4*$[]RUO
P<@CV9A$T4H>: 5J ?AL:\DK-_?FD?K&M4=4@4;A,@0 "M'EYY)+CZ*Z<;\YE L!4
PW,6TOC50+9%M2^:KR&%E>OLD:0P8X#6-..@6(L:\A+/GZM^7E6HR1"C^ULI6W::^
P>1O MM%;[&HQ!]#ZTH&G37')"5/*X!9G_GY%"MC.KO)J!)<LH-)#JB5FC^8"M3-0
PKB]+Y'_\8B6,S>J=?!PV6;WCC<000N$DYXMZU>2DOLKM)6!BX>:5O1L!&C[-IX=Q
PO.8+&!R5(DEDJ301WAZH>?;+$-Q"#@5J,02%W5CP28?^A%5#;TU.>!EBNA9P;U@@
PWO<I'?U^GI8U._\T-G+0^_FK<X070\N<$=%7_TM -'109C7TR3S3ZQEEX5[MVCM3
PM+5HD)2$C:Z],0Z<N?2/PV\),<XG_2A.36.9HE(E7*0B\NQ/;I!N@U-L\LB^TRI]
PDW.^E^ZEBL%!&*?W??*4PEK@0UPM?O]<AZ>,S:Y$X5F(RIH'8KQ?5&\KP>B-1PGW
P,EW_P,O-'JLHL_5.61 YNN\06\@KT$@,A=1G)6J0O$IAI&6NZD@7F;F%-6B_  -F
P)ZAFBR'>DSYH'@:I0^KMWU?RLO"+JE(>T@QN$WGCS?*BUJ]M1<CDLN0C8/3L[Q;W
P/G1J]14S+$B13^88[J4\9O$O<)BL* WVL(+MZ2!NZ!9<X=O,+2>$83+A"(6>K4'9
P#E>H,6[_JEZ#M%8! ^T7!,T#LA!>DVV*/-3Y]S.SEX \UNC9R:IJ;XUF:J6<3*I!
P(Y#':D@B0S?@OA;M3WR9YC  ._%_K\\S(%;G@A+PHSV\5:W],] *&;A51/\B-^P3
P0%(W,CF"W2J^\$>9LQT'*9[KG40PQL2$36R&_!0O\J';7]R1#@=5 OL&?ZSH3?F$
P[S!)>T3UG=:UNR<<N]G5P<*Y-_B:&3K[UM! 11DKM,,AL14?BXXJ0S*/.1\[=M\P
PC4BLK7_1)_VK N(D9,[M(0DH[&3,GWSMV&\]VX>C<^7D3_B\3T7#],X=D4M#3++*
P%)NY'9=./=^'RY&7(7(E2&:UE5G//WV5!V%JWEV,V8A1P)D3EDX9\K".X*$@P3IY
P3\:0-B\?W#EI";F;!*(#]:QKA.Y95$UMJE700RDI@"K+&97L[=;@(?#&14(CR2_B
P51-!B!E-@Q1&<>1&Q1+2::V%OFHK@II_\$&GU[#:-3T2[2T*7=/>N)BLI#DT%\2>
PY V!>_59K)O->C0Q(%;<HQ*NQWYCMXL;NIRZ2RBRLBX"4WQ=B&MH['<A(4[NW BD
PRP=V[<DK.2I>YY6V-WD@Y3#[[T5@EK5]H<&O6W#/@^\LJDT-&Q-3]_+^ @:S)PHX
P&76:<SV9\GZ50^-Y:P\)UL5VT5LDE61#?N;S,9]VK:QBCQ3GQ),O"WKJ3UE/9?U5
P!T+_&:]^Y9M(N"M4G(;18@YH28&CG[2GRD,P7A-R_%E[B<"XM:35B!S][K4(^U3O
P[U\(5]73'U@H/N/Q+Q?!WIEPB>[OX- W?B,,)J"V^GPB#+I7^V<@@0FZ8T1A^*3I
P.GZ[%YQ< YPBP"\X_C"P1H=F[67=5@D_#0FL<Z1E34_.FX*H0#4PBL[:W;_1XEOI
P&U8=-FCH"^DK4[4]3-BFMS )?SNM6#YY$S(L$B;4_T22R<8]^- X+6C4XHGZS@&-
P/?EFY;(>/1.F9M31 3TIHKZQ,1SSLT<8$&J;"S:SIJ$#C&>%*/T*^,H21N5_0IEH
PO%J=6I+>]-+96<Z0&>>&3,8G[[S^2!9M'U:]HJ*E1."NV@*>Q!1=FT]EC!Y&AHW&
PWN"6M/:Z %] %>_F8J,#8$V;VF\QA';PLR<<>%FZ5J#!C9U: 03*>@BXYY\I@@6R
P!YJ7%N65-0>$AE/?8,'.'T?& J7^/UO&Y>V+ \6/]>7D?4;?(C>>LFTTP842M0VY
PDU78E674 -S#U.KC<E\.,,]<_#FZ"1A, V>?. !Z,*SY*)ZSTB)2^GHGVPI(ETOH
P]$.R//!J1*US*%*?C/)5;V?$,0@9IE>-B;ED:_F'+"$K5PW$.6":8;SM;!0W"OU#
P9:C17/!7V6&9SYH++6B$6H7DH$?T_2PUH\$"UZWEYK%/!4'H'/VLIQJ\D/Z51^^?
P&Y0XU')D[5?08)3J]Y.<XVM*H,C="$^;CZYV<FCY.O*[!=LZX)?*'"I>@>[FA2YD
PTT#::]QQ-CH&\X\@S/E(ZP?<3$9IW\1M?T8'(@466**K9G[J9\S10-O'$YEY^)O,
PL0NL73V1;F!'8W]9K9\'T!ST> ABA_'E,+MIWW=J+X_;..Z]/"PK:!,LPQ]T%;M=
P&#BA][S;OP4J4BU$IO2QILU:!$5R6?^:JTFSY$'X9V]GA Q!]3W+X"#BB10%30Q?
P*&42= \IM0D1!Q#2,!:==G+$3@7JJYE&,VME5@\EN#TD)D*'I%+!\CQD9(=)-;CF
PPQ=$ZQS-Y(68>QC]NH8BWW\EN<(-\F.LE7.[N3(S$[[UD,,];%^0'[A'22L><:?W
P;+9W/W=?:E?UD)'WNYQX[J[A!^BM%:K05SS*O<.F8*^4N1\QT.DP+/U_42F)<[MZ
PUTZ:I(FO@NA-7GL!2I<>V P_FS,D,!OL"$K_ ?R,(*^5;?-E17Y3*$6WEU X7N%%
P@1-H%.[4U6MN0R'G&8<-C:?)[2X)T#6=#1F=RL]#,1D"QU1'*7?1A;=,34"".97@
PIY7@=5</\*<8M#L_=8?M)J72I?^K=%5_574RZN^I"=#E0Q( 8\T\TA?6C0__-!Z.
P_,?]C7+8W@&O[?NIMQ!LDKH5F$#\BX=T ^IN*"]Q<YF(7RW2-"'VB>(1']PJI6.?
P.%*;I0P%X+*>:_>!U4NI,E>8O2S8SC!(7BABD_X0)Y8+#@,FOXH10,"I3RW\)/JL
PGE$G6;\]_[1J%H_O-_' @IG(KDN@UDT]>GC^E(Q>'.23=N55\^!PS47M[)W#_O!M
P#9I:X2U6KX0T$GGZ?%-UU+1NM; )&G7#_YVSS>Q+\_07ZH?[N.U/6X&'H+-)3&SR
PA4"QX'5N["40AMQKR[*XK_G<#/=6%/'<U"[D,FJ!G_:233HUL$ NQ_MGC%.9V*'=
P%M/<WMI/+%[B9/+FH^-"F-ZDD7<U!C31\A5])O;7K00\TZ0V0G4F$D'6B-U<FZ4+
PI-.0!]08F(&-&3D1&H^'6V'I\ZTJH3!>"E[8'FM=NA0A!PL:S$3%OC!B:@^[^<,W
PXYWZJT\9T*Y0Z_,4W3>1!8K6I?3J2XV\5[09:;3JC7Z'U\15#9] EN#ELSUKHBJ-
PBH?UH'RRV:#)//8.["=N!TX9*<FX"W2;^'X&<1NZ9D#HSWL)EL1-(]LMFC8*YP9W
P\LVK0>["A. =UP86=TXJ5!BABW4?OTD<5>MED6KFU:J.*<]+N2@[<X@]SDD;>,P7
PJ=2ML&O!N00F$T:'/HI@AUN[K,K2KIJ@Y>CW*+E]EVW,DS5_%Q;%1N=58W-'A>-@
P\-;IZL#EZ]*21&SEGV8.<^6$F3.<O'ZY3)2@.<<A(DNZ?C*Z!_$&$JKF*)P,'][P
PRQ5LMLM'S:O_R2=/S:"85\&XT\/\]TFI<:=)\%'ZC5KXW*Y8B8=WG</NW,SF?]BV
P*<*[[$!WW"B9IE2^H=/28E3K +I>J@0IDN8K^<*#4,U,.AFM"+?H?9.XZ7=!R0?H
P+,$8NC&<VGP-1XG29W])@*$3*X+,!/P/.U"X!SI&S41,+09]-F(!RIX'O41US/9 
P5B$(O)(YS6!#4-:F-"\3V/8IGN]? IQ#'-T_+QM!$6/95^C5U#S'GJY]Q7OJ%8&$
PMQK78(?TGXE!E*3 [#+]WBEY-0@.]7-\2-OJ''Y7B:3PH46T>B#7*3,K-Z>P!O/+
P0 ()"E'[?B,R0U2J3>_MK(H6ZG[7)8320+;[PT%9HC$BF%JZQN87]]_U Q2I>4H=
PZ]:VT=G?$7=6]'/,!8+4JVA)!-]3%+F/N!TM=JQSH''RJ;=TSCV"UQ3Z8"V>OMWP
PJJ.>(!WPA \[>MS<MM8@[=N#+T*/@/$;*RZ3U"'LS"XW8/+,K8*H5=L"(7ACV++!
P98H[U:TV1#WA4@UV%IG >/:<XT!6,Z;+K>\!RX)'W#A>0R8 U[.W9Y"$)-^@3\A"
P!%"V+4&J1%#9@;#.Z!IY,:W^[_]HVC\(KX#Z<,=;8W1*,J">I\Z^/%5='E]S$3'/
P;&10S';B^%WGCSOC%RL>ZZN;,4SK ;%%9/1&=^7$%5*E.KT.MV@*=(OJ.V1?^.&=
PBM&-8?DZLI>!<PV<8@R^BY(:&5NN%\=.<0M;RF6G5IT0<6GDXOEV4<W5J-O"JK>M
P+QH%#W>].V293' 8CN$07KH*IPQ< '[[(QQC+ETX."$5Q-&7>IF@BO)GK#NB'^,M
P)3"8<?\<\3.T0^Q<3@/_7FCKJKL6!)[-RXM;M>R&TNE?TY<O!E#AD-9E>,P5U@R<
PDPP&H&0M0"'X+S'N_O$[/?7L+_M'BF18C7D0;*H\?<9\O6F,>D*[$0U&5!#"P#4%
P0T,)CN[/F_SE#XV=CH5=-<[^[URN+9T0D/?9.X%DO=X/[*6>1!"%U+2+#HHCSWC3
P7D)3S=.C5L\/ZS]\H]60!S(Q!=V4H R%[7BB;D3H._I)S3L%K^XR:.%HTVXYD0X9
PLR1C44\LT^*2_,2\T[_!QO')QP.:RB[XD2?"3S$^\_!>KZ]*)S&"6)"=\S0+#A!H
PM4'(/3]T4FR[K\Z2=,X/="&TO@H,%8XP2NS^DZ6NQT*&N+<3X7OM@^S6ET1![5S.
P(.TD&HI>8UA1!CBG!]!DI_=Y^.DH_=<]&ZE]H!;T@BSSRF#9\9Y:]DZO7O!MW6XF
PM19!+'O+"WIP,TQ3G1PB4Z7J:/CE!PB&X^XT/&[*0^RY[E#7MN 1F!["5*Z6=2O8
P9'RQ5BJ!G<@FP.4YAP6%#1#;C7YIC!T.LC95\L0O[!65=5-J7]&G\Q?=#:$;59"E
P/YD?C'L /8$X0>@Z#2B%P7A8;H(%UV"\6P C82>W ,86*5'-DZ''=J7K!3:\ #:2
P77&>E1J#!7#\U7H#N\IT."9(*YEZ$\==)<P"?[  Q#@@/)8_4*]+LG.*0&!UCPY,
P/PARQR2K]XQ30='0SF+U\Q-(3U:/E?X8>M:[:7^'MA6\QN#;0F =ZJ3)X8K/K[^-
P54^ =YVMP^<Y9_J/.SH$$8!H%''9ZN@J]?YLQC3T=A,A&+ 21GK$6U?I4@T# F^$
P'<[N6516AP'S);C:CC 5,^T!=D7 8(X@[X4HGVA)84>A0U*RI +<_O_!JH"ZSQ(_
P-K22J9P"+M3UKPL>H!MQ%<LA??GE'<A^(2^F)M$:K9+>'TFP==?8[FB";(!KPQ'B
P-<6R@N[XT<%ZQHU=3A9X;^AXO!'BG%%G8W6(0#(=3Q#"?G39G)78ZN\Y,H$<-I# 
P*>&H6EJDGK_%1XI=<BT'#VD^FA$&%RD$K5ETQ:\&-\Q4&= BR2#:VS^K["WHI$IZ
P#@)O$:Y TUBA_Y<<03#MW&/>2M/K^7RVC+!D?NKM?MM_X,BG@A]S"#XBMV^Z_PK1
P03;2:T!*N&$,(>:$Y(V50=,_QW=NKZ_X^NTP-M6PP2]K?95U0"\> YG9QP6>-$.X
P]7Q--.-R^.T*CFDWGEO#G8GESHKW*?"=Y<_FMQC9^K#3I2A"L^RX9@&VY(BY Y!<
PJCVI_;1=0/]:GVK^_7;JK%5-FB6=7& ?QY8D&>^P!_*?SR<@A, 8VV6[2._(^P"0
PZU(14>**/U7$;U*FGT>6,* )'!KC(:-^D&@I^X&4C59 9!YW/M[;>7,09]!0)D9_
PM$#2,-$!>!ZTS\FWB4J%<XF:)Q#L\ZT\E$YC0U[+/*Y.*2E;WC< NKK>D]K_ @6"
PASEA0!7&75+OH\Q]%IL)DHX&623 B2-Q"1E=A)(PL3POF8$80CC15OY&P^!GDU.#
P'A@'V40#+P;*]A_A_-=^JP!6>6\-YSM(D=^;LSAU@8G&BUTK]$=JVM=$<GHNQ/&*
PX1[HA9Z'<TIOD=./4$;WJ?</*-..Y?+S*PNK2,:BQ<H[J$]$P])GCW@^H4$7/B$*
P3)@$7.%)ZRY8YQ[?S2UD-?F*53#ZOBT@QRNIULJ=2M>V<VS98G@)!P.QB$5VE+++
P0*#JWP7&3R4,,-4NY'/-+L9 L^(3QU$L"L@3I"0B!Y,#^PI(P>G/^U7+R%U'57#0
P0F#_.._U2&WKC0N5&D:]KP<L%7* B@Z\N/6D@7?-A>]5D4>K<.,:BOB'Y[B"Y4#3
P4*B@ZRQ(G5V)6_25IMK/$.%UT-U?KE(Y8].BN.YA-OJ2^ TE>.MT)#D7B4Y$GO-9
PJN<)D%F:]'X;\IRH;4 BG;FPPGC3F693'IQ;@KL/)=$9!9.R?C0)V=89VWJ@#\1#
P7C:GMV3SX?*[&[D7&M8N<["O6/D.TZ1Y?K'MFC\8<:L8$$J&OYX)OK;:C6DRM! 4
P^<QP3*X/^;A(EIRO)3KIP;15%.AR._E&:"GFJ '"J@\@H;(Q1FH>U72J&!$E+XQ+
P@7HB+3E($*;9S^ K^H17%VSGN]@B?L9+L UHW,JX).3N]F8B#(B&Y(C'HN<A&5/@
PI8VN"*_LQMD%VX\-?4K!&93])6<+Y.VOGP=:!&'#O3/K.Q9)^E(;"4E.6*I/S0 >
P'OZF(U+K$"6JUR@T;*G&W7#&#'$* V-XCEL)SGT%BA"(;(X1U*=7[NLEU9YS<6P4
P?H*F0:>.CMST#UW07;?S2L<T$[+C]K%,L@%S-9$M-E%J<8>G&R2(IQ0DYP;W]9=S
P@R&<E$M@B9BO6O*T66)@:W/?K'GA=5;X;*!*XICM!Y<S[J2TC?;Y[0^MYXS!RR.H
PL/S>'RO/BU*UI:;Q2:G3,OZ[2G19C9(92$X)%#UU?WFF591EYD$U?[D6+[TV#UK:
P!&-NJ@"<4,"@/P%Q<]8$RON2]/H)IQZ9"11.XB\$H9=DQ:PR0JTDPD@,S0HM<EPM
PU;#1O?),,-4L'N 8U "5;H$.&B,CG[O[[FE5HH3W9EGX*Z# SO^'<D5^>CVOQ7=F
P*Z%0B13W\4[G_.;PV7\Z?9D&#-8+VGF7('2);=C]?;@PBD=SU9N:]DU-&9-0.4((
PHONVKJ:$J6?DE[O234Q+AI \"[B S%"2*_:PM*$Z5 "F$?'6]5G"+KCG>N=LO$+_
PC\Y6-_9FP;Z@-7S\]:2'E_=/C,N=LC8%A+%Q6D5PZ9(7\![G\R<B84*+_/@VS_0I
P4.72FPMFYT<'IX4P!HXWLFFB8IENU^^8O-;6EXE5$&P(+JI'RA:/'JM?+O0^UOY8
P53_^?QU,+GF(;_HW)0^B=@\1KS>V>FN@"LE>)K7Y8D,@UG ;+99%I\)2]8644S 8
P!T3)]O\9<C3>5[+2B]R33CS0G#"Y91HEVV#QQI(#@3@HJ!Z&Y?Q1@RJB#NB;<U8Z
PB>2\#QM(2-7EJ'9\6C+]XOZN9;F$?-O"M4;M+MJ;T6D]IVKZ?(BETX!+!")MD*33
P8I+><=_(%_V&)  ES]#-J\>UQXM@9E53&=@?V%U0.6>OV)-"G<#O]000@IN8V3B6
P-4=^I:%&YM*]S7R(;J(['O$1 0':T_F%O>@;K<EBW3_2@QUK4MBZPU%@[?TBSON/
P<KW4Q+B;?P(1X)!L,S&.]&[J"E32=N#B4. DJP5)S923$HD^V1B^F-.:'SPVG2JJ
P 6-K3FI49G<Y*ZUP-U1Y9O+ _Y)_DZ*)O]V6KS+EKA9_M[3PD4)[A9=ZVUM&;78#
P:LB@[[7_2.#S<^CR(;\GQNY3JMH2APX9 IPQTQ@X 6KB\=!-@[:2PAJS\?UC),&B
P-OC/GJR"J3:GTGJ5KW*?\EP1L>1&&!_[#FS["OG+Y+>>(@)RE?=,\7 #!SL'M+L"
P81(KI5 X,V0%R*-[K\-JOL",;<?DR ;2LW#-)7!=^%O7@ ZFF:/X^&F#F1-V),$$
PNRWPS3F5.$FG49S<YM0G3T*C2SH/2 U^]N^@P8]5W#^<)1QH<LK78' ';*Q\-L7U
P%CH[H\O]_CN[>BJ5@HAJCF?3QXEL4+C@]<*P-MN5\P1&/N.[<MFN$9COHTC'+SS]
P; ,6/P]6@2^)8,UBU'HA\I9%&@UQ'6+5YA'0BE]S8\$;O!'1E<[G)4AYW\B>7X$]
P-8G4YPC"G-U393&1SL-@A^8!7;\3,=]N=ZEZ8F>108QDG,%$+7]K(Q9-(HC?$%>R
P4W7Q;CNE$)V4E_17,6%A^YY($.-DABI?+#+'H-S-TF+$GC=VQJ>."$8;_)DT)\04
P2"F1N3?;4\Q1KAB])!N2"+<O@BH+4RF"'[0R%TB>H]=+,,%LU4ZW$=SVW7]MV-&-
PPB1>K2Y]OS]X,OR.AJ,W(_)]AHU&0E^ %"N:;1Q]2RULN$D4VYP= D[Y!730H')$
PYZ"O#@>J56Y+/%5Z862SCT.;/U[T/4R9QULA+>GO^?F5,_2J6Q_W[[Y@,D1R"%YB
PO]3!LR$*&4O?LCNB#EV@+'$O=1AD0L4TGIR%13+]ERKT@FS8NID[CTT&U$FI]AV*
P/GOK"*.>,9]$ CI$RI*JY6D.<XWRO)R;*;"3CBVGIA_.:)@"SE#G69V_/5XC8HEM
P&E!H-Q(6X!]< 7"@<,2NN"O(./^7)LX)CASF37(\&?LC+(]Z93?%>&Y1H00QH9>X
P;D:#B88.RWTIELZ<)+KT\4ZWPYE ^YY7'K<>/<?*6*T_U[DDY.E[MSR(YRP9>VV'
PGL[-8E0_W8UG"S.^4O-'4LSA.5'R_N67QULP]98U4 1/TMH9K^7PPQE[U'0,C'S@
P/+@"#C*^BFW#*NUH,UA0K3Z/6X7=\R0 "S.Z;)*49K)B",F3Q%!0T^LMYFA.8"M&
P X@YM:&TQS=USL&@+VO,\5-8!T?L(&V?$_1K.M@33O[6VQL;:O<L@#G$$"'F@)ZT
PM6<M]-#AAE1O5W4.8R"GRU"71!)4%3FAN5C-[0GV-V.<A6E-R!=].Y/*2 %-["0@
P!+PL.R/0WT *)-'2)8*D"%*EE$5AWF<A:*BBPGW[489L:M!189I('[I$J'V"0%?,
P9C"S#G!F>4/4'N#1&&G$Q[ YKW5"^ZTS <\).!PR5>71^"_7)3B&43CD,SIC^N%0
P>TH 59F-_E2IP5>6OGBYX,," %/3_IA'[X' B<_QPYKG#!\8]!2'1\EZ-ZVC42R?
P?\0K%LM)9ZPFJTWM+JD'6(;V\K(<P:<&-JL4(UT"A95OF!V,#2^R&'5JV?Y,F_E_
P'6.KN"JB2)R(8[I&PWPB@-OM&=\4Q_]*+S4T3?5Z7PN4;RE2^PG2,N\1]#()_W5I
P9&]:6I0DS(5@HZ>%@84*GSPUILS%E?79P]JMO>G&)&TZ>4!8'[0OC";2Z3%1BT.X
P010#')CC2RC\(;2#F82\^6?Z,R8*GE]1Q0%J8<NTYZ20>UN!\^*;*I_Y);*98?;#
P>:($G,"8T*0S7D2I=E*^V=0_I?E\*U_IE78XBQG.!(\5)K$/IHO!8&*?L9GN/B%!
P9)01)(NVI W &TNLM+S!MS,ZK&X&45\X[J.9^[PWX_Y7A'X6$7?UWI+(<GA.R@@;
P>T$$QN;%H>@_MQRF>5PPQI@Y@PQ0-&:]JJB91CU2+"[&^*^HA-9 !$1G_EY"U7<1
P;?)=#*].(\RI($#_PH1UF"D_)972H)"0A ]-\W):(TOK\,L7E_CWO$V0GD;@=A>,
P,Q$@"OU>X % C$"*8A<LU(WY\XF.TVU$G"3=-[\$< E43-],%TG/+/G\KVWE';9^
PEEL<:KA/F!F[X*GL,=;]1=<AY(H9I?@Q+7O:P-&R[318\IV;=/O12ESOXV;Y680M
P :/I^TQ=D6YUA%KM*H>: <V%OIK]L5<1<Z7VE4U*[>1NQ2G*\^38+YYQVPW;T.:2
PJ7ZFCGSD+3+>S1"H%T)P_$GSOM4SYF7(\M\ A6/]3YM,DM_V)"D<88Q=V#5XU7N[
P*K<?HOU*5%G8Y_)M[S=9\.Q' 5O3OFIJ:SD['CNQ*(W8_8^H),"(+3J$SFL!K5]P
P"3\YV/$X0*H;59EL'H!Z'VB^VR)P9\;-$R'*E!VO[AUZ-4WD+MIY1 ]1%3/.W6=B
P.&/[5T/B..%>@J,:7*U_5LCQ;U?9-E(4H;\FP)W?SCMAJB%;MBNJ9/LF$(7KUA4C
P;@1L_*7IO# 2"C6VON\YC(:(J34S-XS+/0(YR1P!LB(DU?Q9M<(-I]O)BO(/EP $
P1>ELU ;*M846UM8KXL+O9U90VJ1ZEZ#;R<W63#<?GZ?,$:G?HJ*3?A_LC 1G@BU_
P ]]V7N\F?9"91'' JKK.X 57#A54>4 BMVN9=L0*/7ZRR;SK)FB)F^K0;C83H V)
P<EXNCYP2"+!5HW8?F3"!@9PM>)M:M8YER;>"P%F 5WR04EJLVLQ-VN81=O%*:TVZ
P)U=1?(92 ]7E#0O?]ZGEG?UFJV (08I6%%C]"3-7<;<U#P' T)^P9J?_Q@CD24@C
POC3&_2WR6)X)8>=F3!5LMZ&O(<A$66NN>.P?/:XN([ CR[WC^C[+N9W[ERD"HDI6
PC.A<3#*Y[."9VB.W[G,54/2GOYXZ(FHS>!^M7]2?4'0&8H89^V;O 7WHC9;Y$1Z,
PR2QW[SC]#\P?5ZK9L7%'QPOEL-6I'%4]>"A<-J7A*->7?YN[YIGK&H&$:MVV$_+\
PW\#&<M]R=3[1ZT\;!^G*<)HY)=51SK[BC_]6GK='2L.K=,1EVQ! I;LU&6@TA/Q9
PEB3"%XSU-2<D[6Z';)2Y+)Y>,-I[SNI1+I!K'U*#IG&U2H@GX4MD!4?+S]9+1?78
PO=!82]4EW"<Y/C)3-32JX#T"H^1^-=2/-JG"3D(!V'>\>--&?=35;P^( CHUOTO*
PXE_[W Y)4[#L\<RH_$_DY]?EC33V8JS5(:JZ'Y<[':>W[5K@FY'E%RNU3Q1]G/B@
P+O:M6GT-[PX)]N68.47(I6'M[BN)+RACPQS7'[GZ.2D7$F)!T1+?8I)T^8G)W&SZ
P?UD#F#>+VM&I>EHFU*39OBOS7V. =__XA/?A9>8WN_R,#)(4PG5).B$O\F4](8FU
PHRR($7OGQ+7)[6J Y=6CPTV7A<(MU\JD1(\WBAO!'1M&C9?F=]KI3?Q[9DEMDPJB
POV/@3 O6I\1'*F&&EF252DZ!/&=O0(7<QW-\/OQ^=T;PPZN$%R(EO ^FV\\HW^?!
PZ.LI+8!!Q=CYHM'0*R3E1RE!$H>7[VSFC8A-"OAF=Y2?PZ.&_1;2IH.5CW/C+I=)
PV4B#;TRD1RONB47\SD&)8(H)YGS4<GRH)\1O#*#%WSLAS:4),!"5HLJ$)F$&J1SM
P:+>L&%AG#$B% !)-5MM&%+&=!LVII M]J16%+$M]\^OC:!%C$X*(E&\Z7,D&^3'<
P,;I31ZND\ZX;H"@>-42F^\F,50XDZ9-VS[-:^Y7]Z"M2XC80<GD(.1G)%2V_KB\9
PYIB!&>7RPT&TWT=6@KZ>%M)J.';-;^S).+43^QF:%1<C7CG?#5DT>FKMY% L&2ID
PCBL(&K'L#>0V>%4_2;A>O'#%'KI:J]M$RQ,.9#%-LHB%5=3TIATQK7"-#IGM(K_[
P .+/_5LRQJ=T7Z2+[*?00ZUX ;CW=?I:O_1"J$5_Q^?OI.R5&3EC:R3-B10:2V>U
PAU/Q<R5ZA(T\L-+4S\[3_2RFF!N::<B:8/LC"(.1W*NNG9\4P($&97?;]:^]112Q
PQBSO0T[QTPY<<PMPXR68^U99DK235IM%"KU(%.,#B0.1B6L+[Q/.X$8%AE<5"-,C
PP7T&0G\I:W.3_E(GFCS%[AWM$,0?>\I#<7$7!,5\(FTTU56$K\("&&/'!3+I+4ML
P-,8O5<3R<(&$FT)19$QETM_&R>N:&ICOBMS5,*F_G-!6E(JXWUNBQG57?HYU_',A
P3M :F[:LUJ)S9*-4&D X'CM(H6+M0=A0WC!=Q33 @NTP#SAE,)(U$TE</.V7)"P=
PQXGV9L]X$3"E2[33B]1@O8#ZFP1,_(.=S&'IDMX6\)_<03ZA&"#R;2*I0'LZ\3AW
P3DRY/\Y'C]Y1WZ9%#@#QQ$3DU^V 6&65-S+.X*28R5LH1QS;@"$J>&YWQADJ'U:N
PPQCNQMTFU<7F'VF:.$1$JD"BBZE\-)4L,#]?4>P&PC]<K_$U$&1DVL@10-9R*5N'
P5>J0)L@#&/IKC8-0,&YXFOBVZU*:'\A#:)YSJJ&F!($?_F*OKM11FBG:=\MFG$7E
P\HHT[P;YL5&^VZPF%A+?*.K88.9+)O&>0^.3P$Z2>)$IHE^GM7X>='@2KQ]>2[PK
P*'1C5\:%-*=$NP^?6P$N.@!2W':&([V@5<X "NSPWN5X&E0CK_K69^-L%SSK61/G
P++20,A08EU;F@L>!A._GUA,P:Y*+HE.'G6\ N\D@"AW+1LW>Z#>R69)!O]-Q5EX3
PX"RC8"GM]G:JLZ3W "#6(3Q47@?UJ6<:B2W.L6'Z,*,?#D/E(GH,!?7RU:F,&2H-
P\RY%3@[B4<O4R/0K9&R_Z@?]6K#)<B4X='T%%;=STC5=.FT5W!\>X-J*G]8#"2-?
P6;S/M1X]P5L#5CGPJ7$CAI#6^\.P=(&DN(E(PUX*T'B)HU?KS][O2LGJ]&Z=&98^
P_YD1E29>^Y/AY!#PPQ>+YGYSG$_$?H9BM>4;!+Z1\EI2"",#?P(63;,4/VB2+Z9)
PJ-;,:P*XV"00D='.BYX44CBTEP\BTZB >3RH5_%(R":JK^7=&L%1.*98@HFRA:1K
PA%.X]-[,U7T>_0A>'N_NFXBGSAY-*#-1I(K$V>C[_XF\$_ OWS10O'NEEO4DOS;>
PRJ$@=1&F])ZDM.H/A@[Y##H[5#=F\ W$"XE_:3S,C.UO=K]#3/YWFC*,TA6N$U:M
P&%-=9PB2HOGE")TE)*L"61 +\G,+;4;E&+$,-G _Q8W0]-B7,?3%4E5_=>C+MIGD
P2"'HAQ7VN?G-2*089" E0<1]O0(-L!!\43XQDP9?W:HA;I3U=>MTD[)04S.4YD4O
PN@?.=P7*BGGYXT>#WSHASPE2X%$F!9G$ 1.E*7<1-QO-XSTY4W$SB&W)\B]R#KZH
P&E_=K+PEK4*2.Q@= !1"O]4>1'_:P_$ [.T7*$XR^>,,1#^HGZG\S9"IM-0]P0UQ
P"LX*0<TJ,U*".T&9"B_\7K09:_FG]?DIY/PL[OPV]AQ517#)]3)U$,RHCF/P,CQR
P-(3\A_AXF7TE:1+9,0K:'$",%/6:E=I_REJANO=\34BS'SO@JQ#9*^TW(M"':/GA
PVCFK5LSBA4J&FX>5I*(N6-#,WB"[9QV/(<P'0WFMEDQ%OHR+P04%SR."+] ?_^-'
P)4M,F\="Y?O%LW=LOGCXA*#F4M- 'L-BJ'.R'_^5Y(]+2#CQ#'P4;#^PL5R)U4!A
PR=/".-?1HKF(6I(KJQO^*?B1X'0=LOJ')NG^9@':%S;I'(EN+&Z;E0QRM=L"R,_&
PD_Q*?MLC9)G7-EO3=!*11;;H;*CQ)/K]% -1[Z>V$/<> "VA:#+F<PWO^^EBQ(Y@
P^TG\AEE@\DAW^!%]V"1EMP+"YYNH/M$+56*!@[P2+@9[.':5_MUZN,L#5D!I5RS/
PQ[6^!5HW)3^@/[32&Q^FQJ\VQE9)#_@1$&C]*<U;09R-RFTBP0]V%@RPHR%[R6)B
P &X^/50DE6S"%.RBLF(./:%SG5G]XUD',9T;'TT&.5%8\.P\7BK<!5X+T ^><?%<
P5/V"QUNJFH0[W2#"9Q07C@13#WOK-L #L;#4XXY9;2[Z0=Z93:BD_A3I@1W1(&YP
P6"_H:!MGD+G \QU/\:J4607;/IC6)I"7NA2,>L$ HOV>;.?HO'(7+EU:2]TR9"='
PZ">3/=Y-7C10Q)'@:N/PQ',/J_75O1<[ >7,B15)B%^B9WREQ;Q 'Q??FYAY/Q.,
P4D4M38Y6^@[PQ@Q]"=BGTO7&;(Q04_M85>T(=&.9ECFVJG_H=RI+RIA95)<^"D=?
PH,6&#1H($A,.L-5\/_<H(BDA__NMEB\PZ112A$Z'!I\AOY45<&&JJN%%5.BJL!7<
PVH]51[RVI_XCX%>DEC-9PWW=)UDD#,&\*J"EPK-S3&,?,WTB1 U+EM8FF'?O_0FY
P;X H*&L0D8?M%@CN2'E'?VB.;U/4^'Y:1_U1@IHHN4<20WL&@A(2T74/Y<(YH_RO
PJU00V&\>P9(T"MOUZH@_&]*^8!LP"R]%:13VEY1J\T)UDHM5Q(:*-.TBX)NM8(U,
PL+%^7,I8,=2+63#M!1CB8J$UU]HI==06S,Y)?-1C_6A2RY.J^U6 G1=>>2R_SUQA
PHPZJ24PNL<UZ7A [1?F8R)_-X,TC&Z^0#=QF_?7&K2Y=@E%(X74OPZA-9^FXB+4>
P07=YB65*IN?M;OPL6H54UK V\D?Q(-21BQ9LR]A_5,?4OS=]6D*HK)9%;7^#MS (
P.<#@YB@Y'(%LQ-R4T[BB/T,%+^A2.W!?/WH[1'&P3_3PE\%9OA$*7)0RS4(^&6SR
P2-@XRX2*'S/UPTAGU-T5HRF94PLH7F@=L/8,++[D^\/1G4 /B[!K*CW:$-&N\^69
P*G52%+6ZE.EO598T7]B5JW1D8QDP'D3<@1:JT+E*+>9HKH^,7U@J96T<NU#O]G3B
P@NR7_ @#^ZCTE#-2FZ_H<1Y1HU:PZ\&1Q]+ 8;(0RW6KPJ[9[HWOC*#"SE"ZL U?
P!THRQ.D,2^:(+@('Z!O%1EZX4>B[)R6NP?5>6,$S5<0K!PNU8\VK_07508U 8%N&
P',X<4Z5PQR6W#7_[O?DJ8K@F@)-T6]]/R@JF*UQ&)7_23'W&R,1]%V)OS@8SVRG4
PNGF*$#^\+F"%M"^W7B)J7PI>=E!,9\G]JS =$!N4#3A6C$"W8[^BA(,D+'+HPJ'*
P5]UCZ>,5<@/E_'9&R<<!OJIQ?\#;CF'ENR9SPSU10^#$$CJID^AN]_X;WI_'D3]D
PL5Y@]X,I!8UC5K\?$&K[<68K2JH8W)K@7FIB\ZSWT@/F#5[XC1@IU3)9UN@503%*
PY7O$(#\'[ S%'#IP;]NVL?T3];EEQXA&GRVB09Y=I1 \LZD:T_/S%>%O/MG7%N_<
PU)O%(RN!EW)H-^<ITQ C,!HD.2'8Y65E5[=*;YQXB%#<G]LISNK059J_3M-<,O!-
P'YTDECA%V3K9Q4$F8,<#E\H%T5;7'PC.&QD!C#[M+PT97HM2C>:_6Z7,H)9LO";I
P"<-87G&D6RF,HK/(/* 2A8/K"5YT/YZA_RG(MM(#&OSB";AQ*"Q?VI[N0X\"A(J?
PW2#S*H$Q]);NJ\/YA$-5_#H/ZC9VK6D?&:9-DY= &7GJA=AS:7V6=YW:S?=TBS2U
PZ+#ES800>9D_7-9*2\8EP?*1W2GM6_GVFB-2J5'8@+^OCA*#>NC'=0>Y8M)$D?%Z
P6QZV]T5*;9I?M@1W_3F&]DJ*5W4S%!92+J!8QN5-8UOIK*SE89L1>3YK';I*T_HC
PV!3D_M2D:8,:- ,0:I#^R<MI"!K4Y\C45]VP [?JHT[B%#"C8*!(7I+4ZY2+][[<
P0UQP9]8"K8(D 0Z(4H?\*L6A3"V6BYO7^RL'VYEA=\EP>"#Q^?A$X4ET%41<!N*=
PY6:9HT?] >0**/1VD$C,9OBF!*:[2>J;+%'WY75JZ)YI9/UN/4P4C;QZV?25A_/V
P/#^%QRN %(+"VNW:^.&%57%9U*W"ZP$#O5A)'<UEB$?+&3P*(OPVDC2)JG.?FK_D
P-$+V< CZ8BE%H?.5%-WQGQ #8""(4^%B =ZS&G+$'9_YT%7R$:ZYH;P,)+)#>:;!
PB+:(_%36[DRL_V8A/#7(ALZ;@TXK[@ITX'%>('4?>G,RX!=W!F8Y2(5SI._ID[]U
PV8 YK6%3E7O0G"+XL;"^-;UB35OP8/JF-[J%0T@IBT4[Y$U2;X^/ ESK-PG2C),L
PUXGWGA3X#5\?0X!+:*.3F.1E+_$LN>7-$$"SDK5"?HB>> ,G?VT3=ZBIBNK6#M48
PY.-1X%]R!*3.[ZT]0T<A>LSO/<J_RWN(_ $\:WSW, GMP.)JB5THHTO+7)=X(=V#
P_P\(=S%A0H6(=1./1R+F(U&BJNSLEG^Q_/M)"<]2<1WPY&<EI-@F08?0CYPY[FD%
PPK7Q 6K5X5@BYP%&^3^:&,:ZG4B5;L/?\?/W5"TTAD"+Q;/<,K^1*D":="!#'!]J
PKY9@+:00S]WUUCC^F<?9@*!Z-I<R9/#\CU:>0MU]Z? .N^):GJVU/6.>ZWW;VYO@
PZ4BIKI?JL.1((EC/.[8[-N/[T3!I$;TH5XQV%G_*J#HALC)5'.P!L/)D9\5<NK&O
P%W#P7"2*XR-5GE@J'?,W@+/CL=+G49_S48>4*J'\;*512/XV.-2G<##[3=9NS"Z]
PU&MNQ]^M4V@E+@CR7ORI<UF9_=\I)!U"1?C>ZZ=KE%WE=Q:PP+W@&ED>ML.KBXVP
PW6.3N?L<=P-[^M@J>5MA"CZ0NMYI1+P!\@IKL/QG>_[+Q_<<<W@]6^;=J$5>YX(T
P=^;GDT(!Z*7#*<T(AD=5 UL"/MH8M]'F\#%,GU#4>&$E(ZJ-,4Z&%6BU9#&:#8IE
P3FJ3H\^WP9<;WK"K@E>0;@%R!)$BX]I1<!*)X\AWTZ\)48,0/#FZLR=P6X[%2X6[
P)\F=L=1,O!*!)OVQM]R::6R4?$2<UL%<6PLQ>+7CK!"C0>7#$B+#1V)[-?'%OK9%
P^N8DV,-;33@AG IW1^K-Q+1;-Z6"6C_*(:NU@I\ O9/8X=#3PE?D:<X%I^24"BT>
P181.K:K%NQ-[O"U$V#%$VHQC=Y]9Y.QOOL&QVM-6+J76"7G!@.'#E>O?<=XUP(8%
P^VZ%D/SR(2/- HSDGY =*/7!'"Y3(?%L)!NCU0Z&R Q^AL.8^;9AC9O.<QJ5<<$?
PVDB)'5\X6P-1@8F0\,/O$H)])]%Y*15 IHJA+ !%)BA'G=%U-H?=M5 ]W>'+S!#5
P4-#OIC_]OM_Z:>M2TV)F3I$RE[A="1QJ&M)UV'C/!:UO*$I_73\8N]LA6)PK%[_9
PKK 81?X'L<$>'N!VK/G "P%G"ZC9/N#[6MVP?0%N;N)%J0U<"Q[4!8?KJLR^"Z($
P"KO' ..C+GL/8.X%C:L&9IG4AOI.!C0 _DF9/DST(Z/VEH,A?G&MYJX="_PF##M;
P\4<__:\GT")J55!1;<_7:YNGK^IE)-Z%1!@0KHA95P$G 9&;I@?>T6T =U25*'S=
P3-2T%KL#BDMMEX^0Q7WF4MTJU+\34Y/A5S,W,';-BBLS[^TIX?TZDQ\,O!;Z0),Z
PT8+M R3?U_O !'8J?JN2CZ>V+43"'Y_TOE^L0=SOVO%' /6X:0_NT@8_^[2Y='[_
PC'CP/D#L"8+GFX&(=+ 70G#K;P#]Q2G)X0$!V#@'_]!83MXKFJB0Q?:_W7_G:$/K
P\Q8A18/TE)4Y+-3ZN+'/)#;K @6+JRR=S5JL ?#(N4[5WH%2Q"VB1+==PT]S78<-
PI7HX-JJLHHU&Z<WK<#?V9?]__M$&J,DK!=V'#.S=,NT2/7B"3__1MA@A_,,">8$^
P"+6Z8[S>] ;7[A>*T;9LV(,J8Z]+X$7;8U=-^CJW:OA@=ADN&/@9K[STX3<F?;<B
P-JN+S^16TGXV%I7O+1S(U6_-*Q"SDJ3E#9Y<T>>=^(E[M&">93>7#L6^ *CAANS'
P\/]08U/S>$<0JCZO/7,-(CSCR>:K&E"8Q(=#3M;0GJ011*HUMMCEZ3)85#MX_C) 
PYZDRF!'W+C^D:YDW>JIL,'+9#(')#8RNJR7N&IB]\. O62IL:9J?Y$XR(HOO^HKD
PL^J?"DJTU+E2[1IL7FACDA!5+E9E E*976"*VGO4HTD+6\G6BN ^NG@:V,4:_%!:
P&;+VV!QD^7<(V?++[G@.#]<D7XQX,E,[C-0EK0;-7EV,A:39H>J5T7[P]3PW,NH'
PIM!UH;(V;0PD[P7KX/UCMN5:KQ?=D)TQ^(';49@0[B] -!5[=MZXE_0(X9Q! &0G
P4:M7F*BJG7AIA0$Q_C8Z$8VM&\T!-HD&UM/$Z)_<#X"YR&>W<(?:V"2F.D[Q/W>8
P)WB  X$]?'=/OUFH#G<V5WU28V&T_LM8;9 :S@M^M"/0L+D8"$N&-IPB86JOXY4W
PJX8[)U29_H%$Q2NJGQJEJ<$G<RA92R:S-2X'-:/PO5DQ/#*Z65%^U[F[>C(?/LX9
P1@(9<0$ G;">PON05A_))\I9H8N0&GBZ^N&@DZX3>;BJ]+S( XXK5UM!S*^'B<>Y
PGI7SA@GKFBTFCIV#,IHPOI1,?X&_K=56\58 P#_PK?ISI%69A"^=*W$*?H1F$YV=
PWS,MR#8EPLGSAD^V;SBY+;-@V6GY@:@QIJ6%$+&6(UJT9'0L@$YG]2[(8O;0FU1I
P YY!L#+6ZYKY6[O9H+DZ2RI7 'AX;'"?*^F&B)AS5\C..+0 X-AD/]E?:H.W!N<:
P>F(8)A>F+(?OCOAA?4=)*(5#HYS@K89-F7J-'(+RU,WS*Q*18BA![[[*_8X>.Y/K
P))SP+^AL'"?U"I1K9[*6S:G+1/1QE0-G-YCN[FE:$RK_[JO;%,\N4\D&]XK7E3V 
P>]B],TR4$.:0B .D9VJ8Y"PCMIINS%3V!&\S4_)K]5 8*BMVQBVG-&1):,?!=/K;
PBA4CBHE[5F+E#]G5M< =+"VQ(S) \B59R1WA(97)(2BRJ\ZT:)<'^&5LI_:YW.P+
P\LFVML]M$<.[UQ\0N\)=VZPZ^Q$F28HI8LAMNQFSKE:=%!/Y!G160<W<*4_/C?#&
P=>O;H"JVF5VG B3=#>_^AL[.FI:=\Q,5.2KP,/J1?"4*<**$6.A=O<D^$H032CI 
PK=)E!H/96FE7"5--!2=DH:S@B/XQ,X*F$^R<<:E=LDW;)F*(%>C2 XM5<;8XA#,"
PP[+C@@.%9=[(GK 6K1W)\)&7<551 @+@*C73FV=451VEZ;DVKT5Z&"TJDT6PLT(4
P*1[J ]5&,3N[LN#T0"R@5K(W>&V4:T"-JM2!XH79PGA/1FYXPB(MHH0 .(7A&9?;
P4PFM_M:=0)\%8 8<-!AAPIO3,I*MFXU-=%SMNU>NQ/M 1[ +0FM>@\!6'C$R#05\
P^8I\KG>>"(!ZY2U1]N'U=!#C&3C<)\!W/1N[$O%)HY=TY7!B?[&FOL#!<Y !Q"B[
P4O,X'9QU@!D=%'R "S/TAVMRPFI>UZYHX:C$$,Y!V=4Q.028FHAQ1TFYC\3O#0W8
PG=OSDE?W.#$0P[()Q&.&%N),L^)Z>N*]]Q[D<TE&(%.#:B>O6&S$(3O:/&O>C1S2
P(=:V )VN;M=A>I_>EB"SS#>U[^FQ:0AO;HZ<J0\,1<3F4U#X(6?0K 28ELWO"R(R
P$F&$,,_N51@BX,AH8)@D1R7]2XE(<L(QV8JBQLKEFF\7>4J[R^!QR#87YX]0MQMG
P0<JZN7<@SN!13=$HHAKTR]\3NWEEDJNCB@.M2>B$;%K#.L9&Z'"Y?/@B<8N68E88
PRB=<;R?IKVVA_Q:OFEN&I@Z@#;IG"73@P;J/U<.RF>U5YB%;"<>)T<?]K.L@T]U5
PW?K#,S8<?\1](Y.>79N5%9@GL;.D],XFL^/R:-/B:R0)&OI/CIN3P&B5&BD1>D,\
P.CA!)85M7Y+QXY6MKL-&#_XL 4;\<$(:YG(@R'-(?BF\BKI&?WJJYYT"F5XR'F'[
P^!B(R<Z\NZ'\4BG63X(2T/D^UQ#:36##6(O'^I1GFP!'Y!^E4FQ1T*:@>(CF6P(X
PN$3_&4_XDL4.V6:Z!_EE8.!SG.D]H%!!ZQ+.(,PEY>-TRL <W72VJN%Y2QFD1] )
P,@>-B!?,3T:("P>6S!3V;4ME;MJO.D<E,\L+C+P-2F61,Q+8TZK)%KF.7II)A23-
P0 $M @X?M0#'2?>0@MTODC]_-U8Z(8\HPL=WKT>BTD@%>#IM%%.9S=U+F;DR;JAG
P6^+L>4,>X5E"[PO)V+Z!BS0W[: B")N#UQUPOODI AXH@3*H?V?B$N$-LC!(24-L
PC=Z 9M ]]D\L].+  )Z%45V)2OK>] WB!H5<-%]<\BETW7#,R1O\<['*#EYV-J,F
P?-R5CB= '&M9-RJ'&#$H<$=^'?*Z ()%WA? UA8BI4[V))%'X]8D#[F^4TGI8\1Q
PF>+'E:;J"K@://'&.+O94KW!\OQB7]5AI%&M;,2(K&A)YJP24#]NG[G.ON5[\!7T
PBUKGE\ULA:KF%-+3/NFX95F(1]Q.?G/L,+J'N(,UBTQS,_K#\A@^IQP&7?)39>&2
P]]=_=P30U6Y_:N.KM>/>SAO#1TO=O0TYVM(J>O-X6K,O"5'9>^,%1K'?1_X(.5BY
P?%^=#;/E7H[52IWD6K?!_>M&F1J+I'Z&DR9L&T:KT^JO4HW1P0FN=) 9@XMTO  C
P$QAY[BN_'2&13E<,T_/R5GZ,"?57[/.W),^D/<;,&>H.Q20];4I3G6/WF(-DP" +
PW9!BXL'7=OH)TKKUN %*/G$BUV!LY.WH\[57,5+F< <7P:_D+P$9FPMXDSI.J9H8
PY /)Q& ,<V>O852HMRNKPJ^(XM>7ZSB<1 _YY\)G7+ C952:Y<86R1&S%[)#QM-C
P%7+6R-9@PC8RM!*5UAC\% CN_UB!!0]RV0>+-S],$)F)DE/.XW\ Z+,YX$X0#1HG
P-7/Q""RLZA! '_J=9)_^65;C[FV$BZOYXG[0]MH"=JO!U6[K+$G'C@L02 '@^TF?
P06_X6*B [%^_;^K%_3VD-#Z%605[<D\QJ*HR.,T6SSW.,1 G_3W_,\O/_DI.5#H4
P;P_/RD(OI/T/:PZ/@>C.*#"6BFS!@E SIJ, Z*FF1%8H(A[[9!"HX9T7 WQ'0@ _
P\(45)BYJ#@4C3'@[:N%%7:6/]']:Z>P9WZ'^]PP3]WV;T"MD7!E%VK=/36B]A(R9
PLNN%W3JRE(8:2Z7NH\=]O+)]1*0X[8-1B+DFRQB[Y"R;YU%+"*\O1P^>;=25<#R-
PBUK.M2E?.K^-4A>+ @]5UO1%=,%I='*_0CPR^2$TN)VLIK6YZHE\@^_&=F%267L>
PT)4OR-S<6Y_?"94,6SFU(']FZ<U[KZ81T0%:COI*A>\LP_:)\[ZM/%]0D/,L+F'Q
PX&F((;T&WC-U$HU0R(Q>D,.\SQ'GRMZ!41!0^^FG9%Y& T=\#;'E20_=7WA"L-M&
P&"7SLS\0#4]KH:$C0A10R&#>2%V2IO%W2P*"A9)^X52[/GKX\FR?OX"23;84J(P$
P*J9TK[ &VT>_C1NY+\[O0])>'AX%4]2\%UP'KN2M9@<+8''68\IJAZ[P;2\&/^%/
POX$ #HQPXB,BM481&><8A<GJ+CB\B;:+IU4%>IF!'Q?WDTU/]-OA6E-$*L-[MQ9;
PS?;(:O 10$9RD38I>L=2X^KWD8T<KAC>_BNJZ&NILWVCF'L/Y/5K)-WZP@5H&])<
P#G34U+7H!U A>&Z8-(8;8Y^^6+S9P*_UOY3/3=1CGZQ$Q Z3H9W/C[>7Q?Q=[8Y2
P@$M(K5<] ]/BROS\'4<T-:.+5_T#YW5B#O[?HP'%_#>2"SCAQJ2%@58[!&ZG3^LK
PJJM<"R A5GRS]=RJZ+-DY(TO2$\@GLXD!OJTK7L=24-SP/^-L>Y0;7 DYW2L7V&Y
P :+!=E"A-_ 4TNF^@Y(>G$#,?F<]0?LPSJJK!0&G%$0R411$A<![VK3H@#RH #DW
PA467SQB1BV^L9#NWPL'3I[)%4.)$*ZB'/,T<E/9E.A) M%7 8^NYFP:DJ+\1WO;B
P\@LS8O,XXSK$,B_8$FONUV8_=<[U]=-47,P"G>.[T*XR5?'<[9,3[L4R77]#B:BK
PG2"262@&ONL&P3J;_GL,BU :P(-2+!YNWY(A;_M-KGM@+2LF9Q#S#N&Z?#&8I*CG
PU=^NR-Q]%R1ZJ_F[TH?&SX'\9KG;V%$*<EM#@3-ZYEW4>8:HJ8=WX_PD:&GV42D@
PQ;$KQE24\#B5I1,BRUA2RCVZ'M14DLN#I>PRV7TEME[]63!8)RU6^&$! *[&>/'@
PAON/;YNQBETR/SRGD!,O^I&0-_R%)!RNZ/=)C?B&2>435S'KR ZWL1[5F',>/+-H
PUUK!"%P [GI@8-4A<0[<(Y.E+#[@P@O&TIEF"=*?9(']NT^>(@8CC8#GHXB38KP]
PVO%B$MI%!4V$IEM<',2T^OP&^Y[?XR?/A..%-Q4K+O 8WX?NN:NRJ!MD9[:/<+#T
P3E@286T+Z,E]-^S*<IZ[8V.)62=>$N>+,;#E>YJM;76M"#13_L"VC]]Z;_6D7QY-
P.;+0H'C'^3!]'2J;>,R.3QI0CGLUJ>]^F?S6!$5R'@M#3-9T;SI"0$5 [X4"OFZ\
P6N3KL?Y] [_FKHB)_'G>UW;YC<JE_;! O8DGT[6*67M$$#R4!>D^R)-CCD.Q:JXZ
P4NU\$SC>[EB"!\#U-,8$!Z[><L]7;34TVW\^.MF5XTD;M&$A4@<-R IA!MKRL_:0
P 7B7-_6(MT*%YY]5-_[H>N4HX9)5OR=@+ILA8)HY%:BW8PYG%X#X0ZUTVA[OG2!]
P!LGX#/\'\(D%#VAM"E7'HY$VINP#H3OV3\>5:JB:K-K?.VJ %[M@M':&%D(#6(EM
P$Z5RLN-4BL"@25D2=%8EY;J7KBI&B(TXI 980WT@XA^MA B0>3 ?&FZ;WMGF.:=H
PYM9%T@KGCMLQGJJYMRULG.3P4(,N&W7[PI3F$S26/XV.\(.44GA*HC/K>D W6(L<
PBPL2Y18^&GRV.9)N2<;SAU: )[F%9RM*BX'#%Y2R:VA@5$]V@:M!D?.2_EYB^BH"
PH'@WKRY5R/S/90[/;Z^P[#/V5K\N'9'$-;9*H4,G0U(R5G,9=:FD%.UFRF\[@&7N
PU94[H$@3M"(3@VQA3+UYH@*[^V_S/E,N %IB^NAA@5'=O>I$I^&K^M^*W1'N<K=<
P%T>.29J*/;'16A9KLPT7O5?TFCOBA<#95>?T[VWL,O)W-@^P;WCY;&0I*0/>LG Q
P5,,QR@ [:RCFA??U;%6F53Z);$U$:*=48AHV "L0;S:2]H[OZ_#BV?5_J@/ZAS"7
P^"VPJU>TA9[M8RJ*88/V]1N<_< ,YT-HUHWCQ2Y^<RL"NCC)49_77UG*_3X8/%J/
P"@VNC>.E*:N3O>+?4O6#R$3IC_, G8(/.T]%:M3,:&S@LR34-34HMMC*<:PXA*"P
P#P2HW:BGD1I>9'S?I'8HV-#O;'&V1FB>9N6G5L:T#5K8.8OC3&P55"6[-8@G+_O-
P< &VW;)7TC]?*SM5"ZDQ8_ A=Y!_;<QKZ"[' 0Q97P:W K8V')3AGIG2H[6F2)-'
PIJU/=V%BZTQ7YWLI-A=N*0A62\+5+N$Q20'@9!)2/6 ,G' Z*-4M0Z-TDSR3>Z)H
P_7-="7[./#SS+83EQ\F<!RH-2Y&?M$7[4.^D*/H(OOY,C;2:F%4N]XX>>Q>F*9PJ
PX4CKCFD$J=JU ,?<RE23=\QM]ZC\R241C^*#3']9QS+ @)2U2 Y#[P&.PN\C"5UY
P!XEC!L^!M0:.27< SF0 RXO,/O/4O:"##8T'=9_T64S0:'6^";MWCV+A-,=;24U:
P_0#4Y0=$3]MFFC997D6CSI9P)L[X,O>,TA5BN]DI9K71=E'5JA.0"N[5)&>&;"\9
P'96)=Y+9J_5(N(%2)BUB)7SBX>)@Q-O'?G67&'^KM8,$1_:TT5<#F0(&]3'&H]QX
PF"2YIM8@-%*\0IG#;](1,. X&[V>$ KAD8%0T9;FAPF^F*92IL=G?&@[K%68]S3H
PIK^%Y:-*XZ3#4/G4MT3PK\94 )01 ]+,4:UDKJ4&4@\4HCR7RZ+;E7=]M +/(A>.
PRCQQL2]%(,#%/_[2Y71 H9M#I7B%:MNNU GSP2"V@@GU$71IGHLFKOK"U%O]RU>R
P08%!!4W"\?D4-68_9( 6 W.T4;IX-@!SQUY=7RVY)=]V@R)V:<1"B-#@0#28^3(#
POO^O)\EVS7<&L,?8C/\IJBW^-PS'3"7:4,OCV1[]V%HY\3<G762"5OU'&I3*S4Y2
PY)>&%QTK+[73EPYTAB[-@ '0)Z^'MNZ&<A^HYHP^P:Q")98&HZ3-[V4N)A8+@\D=
P['_211-&:3$/"*T5 ,FC:6U5<UO2T45,J1.M>?W^_/H4M-3[,OR$" B::*]B@0(W
PKQN(Z_I$OI079]IY =?<$7>>N=SM!^KN9\2$1]7_:B[90*[B] SJ(^2"[03+S<SB
P7/7)FA4#Z+9 G),*9CF.:@)Q!K<CHSFG"LNNQI#,XV(+$XQ;UX9S@A[]^8-Q[$AZ
PLI>HG/E1F-#TL1"<8>W+,"*4!G_],H68Q@ T0S@<:5+&O]>\?OX:38.9K99&&4L'
P3>.@Q<#HDO;X-*>?P=.(3.KN@6[F2NVGKG+6;OF;BLYL)% +Y^72S)1R!Y9"\L <
P73&E'AE(SH0M@)\\"B(/1ZKV-C)Y>V<@[;@/C80P#$&V_\9H,?+'30M!S\G-Z)H_
PJL'.0G'F$HU\-=Z9?\L9WV8/ZSDR4VV/K,,0AV>E)@W3W3Q@4+THB9E,6$JL6@.6
PNW0?DG!+.N62'A?FT<7%*@ZYXC"PN)8IH(W&[B;R!T5:2/HM665S"U"B*53J:%)"
PCR-!'!9^Y9EFT"Y<7+WX&X62&W%/2G<64Y=XC6?H*]MFEE<88JU(M=D3SZ>ZI-O(
P%1/@&FRF&NG&/K[G!^C\,.H&".M7ZCNQCQYB>'3&E1KX2^=WM>S=[1XF_">S2NZE
P>_ C;6Z4QR?^-<"VN9:/L)*TXR52CW>"8A^F5?JL![3GEE\W D<]6F[KL_I/H:E#
P+AFZBF30EA_,!1+\&\@#4D&=Q+Q\PJR*;#(L"*84E5*4,LV\ICD&7U64@@+PT)QF
PW PL@Q9[\I*]"]P"4@XX8_WS?<_=X#LW_VI H&%RG\:NY@.K,%MJ/^EY&Y4R26B+
P/(=%T\6OVL"1/N5G>UB&RRR8>)W,+)!$N44-#*8G.TYN<%<A[UQDG""R.T=_V@S,
P07CN+@I\EV%/DNE0K>0:L1[I1K%52L<-#H?$T EKZI76N"9!EV0<!^J)+!<W/LQ*
P'B_<IU^![3Z\<?=J$UO/@,]T&H$M!E^!'.OS@M6LW-D2>$RBAV)>JC,,H/*!R+C0
P?V>*C+%?E0*L/&MC^9."_2?KCNBN1K"<\:RU<2I$NUP,2&JT\'%QC4&M$9N<-G1[
P99G]8<X4.%.LT%\(WO6T\C^]LFVI@@]N&%$"9GU](A!-.R?PI99!+T.5 VX#$G5K
PAL-WC7'0R?HG#_/\0*?'Y_'N+5!QSD &BS/ZDKRY434,#E@T8=1$(6?BU#794YQU
P]Q#VWD00GGODWOX*3+_$TVLG>J',.F65-6['Q&((44ES>)1T3/:1)Z%F;KU6%.N5
PEC-:+2C96&2LP?.5:#\2D6H3DU5$NZE0'I7X%$0:0<<5^%+.2"HQ:S?>ONDVLTMW
PX3KVZC[::'3@W6'"/]!I'HK:Q#AHW@JB@OC&-HM-F$%RD9E8=HFS]6T&$0H7M33H
PL'J_YM_#N--Q(<QN&WZ%.SP)JF,Z?FYPBYI)P,A_LZ7&"V#Y+BC/0QW64#2;4ZCB
PW=&F/WY--\H[U=N/ESO>#)!&#!C:3,BXR79.0T_FNEO0]?%'%7RK)K#%LNE"PFDK
P,],'&B/.),7-D[&1S[['Q59+L-XN*G#GCS1NG>B[FF-M*7;[I%6%I;Y?+%D)6JXH
P@*\_Z87HO @ .R056J_DW 2MVFJ9),7N4S=>_@QS]*W]\E.]+)==.2G@)DR7LOU]
PQIP"@*G7*H_CO'!A A+#Z-]8:+9); NXS;1_;_R_.FA9E>CY7@0F7)RK1L0/(QLX
PT&3CW@0JG?7ER0VB,:Z^O!R)C% /&3 :U42T>"@(X62$B]X1@:P'1$^P*&N#*6I(
PO\BX>;]@S<!8,!;ZU!]2G8N$8N:*C',@>*E%V_P<+7KM:E\#XOS?@JZCWM$C,RN[
P,/C4;KJ$Y0>FJJ"H^*> O/PHMO_GZAO&,](++,7[4I[..$,;81#WQ8:R1*90:@ %
P6_ KC68L@3-.&.UZ6J=Z/MN[$D-L\X =FO 5O=BD?+&W:';)RIJY^!>41:"")[(B
POU-R- JN->E!8$4".OEOKJFFF,*M'-GHN:AUJHCO7IO98R*%Y3XM;+T3C\%'7?/^
P_RLMJ.>0=1,]V3LZMECNH$69L$G@9;TI1O(0J-5%RDB0;>S6?L+%;P,$#L^)BG9A
PCU/[O>1L]& KF.NA #52MN:$"S"G(^A@:B'S)O) P9.I#>6LBM.=AD;"1S-*;,S^
P5N@',SK\BS&"R;4U!]!;HEK=)K$%E8!S2;URISF&8PD?QP4V_6^?=I(LM-L)%E2_
PEX,ZA17'-QF3R\,K@1MA@HS_T#6@OPY6T^M:+5=:R@A>P7WO:^AL!/Z>W8W0K<^S
P:(_RT<K#<L<?=#239$JN)@'HRE:&>1)-?978T&3"5*]L#Z%NVJ&@9$='AFDH*N-K
P-[1U?.+Q;-R;/-""'7@GK/4]BMLY,"9.MC-6T@&FOT=,9YWF1N19:43-9,J7227J
PZN1*_3V;_]R7M,7T:!^(N<YV(H.QLHH'&74E39?%IQTVED_[NF.1X'FM#KXER[$R
P:P3Q0H=YMKM5Z(5T3LWENV\D.=CV3/S(YDUV).[7* $=[T$W#TYA9\0^T:.2\;]'
P^JALC@"A4)"->@5I^LMT)2V2YFI3C'Y#*/9UCI);/9\U-I]&L, L>6(/M NN:6Z3
P@A<KPBV2CY(V0?<A),N6;4 1CZ]931# W]U[G?AX$)C'AG6(W>@=J@@0,!K@$X<2
P 6[ W2]Z!&6N DV5"[#J5(%MQ&>7H$1V1([._Y]CTR6 F%?R+XRO4HH/H[8=Z)\M
PT-[$*6(-)]*^_YH#N,?"4$3$T8:A;2[Z%CGR244846;KQ5B "]PGGE21U/+\)10T
P S^P5Q5^J:W$Q$-(LU":>WK:'!;:&0@@_LZPW5)P\-_H ,:7K'W37[1"QQJ5"HYQ
P\O<6L%J]UHZ_7RCX(BG>')A)G&9KAV>ZOH9ALO&5U)H5=*LW#/>3=7^X465IQ#(X
PJ\K,$G^68<?<,M]H9G98C+3YM8K_2#<;TU&=X-%M11'ALRE;#T\I=ZF-* 2SNP"$
P[8 I\"<.:&<\'$F"17YB[L"$!9$D-_V*R[-?"55+-86&D1C>@9V_(9:>]@B*7![)
P@R;Z^6O,@MG8(R$"@.%PM_\\I*G\E'-_-C7$ 0*'5V)M_DKK:Y7@O+M7DOBG<VY<
P#3+I49ABG;NX[#@%X ^<PEU"#91)XN"M:R\_L[=\_P1>.:,E52;!U:YA0829?HV]
P%(K4$6[:^-M[R40(^AMG1CCZ&<?VB+8@_QYV\ZLWQ\;'WJY'E\<Y!%""(E7HG@R9
PAJ+4,4<^/:Z*3K5&F(;K2-W=BM;D/"%!@YQ5"RT 9V3>79E\9\)K@7OD@?)03C>'
PT(1 7YG488]TX;@T-.H,>?6VAX1%?ZZ@UM0'+,\(*1[QVJXY<YS,CX \.3S2S._W
PV0:X=[MG\P:>&&"CM^8JHPRZ"EYS4OE X= TC*=D[RH8&E7E*DYU(JSE6Q0,\B+W
PYZ47T?&8')O4'\Z"1I-9,%(.$O%5^2DNG1#">UA6V)SR*$7-JD/7$ C\3YQD^&TQ
PR30-Q!$^CJEVPE!N6^,'K\.-)G$0A\8&QHJ7OW"N;>$4=&G#D:%1!IA2H%@"P#<U
P]RP3.6R%%VSO0'CO^YZ,)PAEA_5GUSMQS48J<'6BXUK7T1'.7SERS46UI3<N_),#
PCG7L=" WQ:,)XF3':J^MW=UWN+)=T-OF#@%V# MKR4\]*LJWS]-W8OY7Y0I_W/HT
P=8O2YJ]X#Q,Y/9W<H)'&"R+>'MVAV"?NB.H%B."/&_:1SQEUD=XM_KEY2OZ1@J%V
PF#CL_%6C)8_]&/JD?91!1A\H+6CSH\!,9<&8Z$''%]H#JOSG]6E&":+!W'3AL+(T
P#^%F;[Y3#I_.]EWE6]4D&TEJ_ AID_#L))%G:/H42;';1;$TLZ5CAWW6<LDRH61/
P@HQ_+PY0(Q 0%JN8!Z1>7"DDM302!7*IT'(?C*C,6E?34+%A,+K67F7^I"C<]RL6
P$;48 3$IE(4XHAP)7K<7<CS($I&]B)$\Y/_4*4:D<24T?*E'N5,[L6?M+#)I]FHN
PVJ'V6@!_% UPE#7Y$%<,02W3_\;D*/3-Y_G;O*97M!)'WU-MZPL%<N<-D4G/ KRO
P9P6U!DPP;A; T4U_#/RA[Z6S=7CV[)*;II07[@7$!+]>Q_WE(R80CG9=PH9&TQH(
P[$<ZGM-.MM!WA6E+&-_/+XLL$I"@6BD8[DW3#>.@<HJ:'>"M.-B4VBYED;OFV2QR
P,_W?"M(M\8E8WPQDV%4"B!1*2B8S.6"3,$61L<S#B:+,:VE0J+-J#.*%7CFW-B?P
P" ]#('][83W^ED2Y;SAO*+ XZZP2)[.:'[/JM?#Q77RBA/R)@#8U6>#O>_VG74QQ
P1MPQVYZ5!R30 -+C+%TSDL*W8ZO<<R^P[?.FI](5;.?G^C#J$K=+ZY1.]U82>O-D
PZDN\"?]A,,@@!BS'6=!FPR],M])15%[B2P[""B6HAX(W\C TGS<Z7ER91RU=]?-O
PM?@]L?Y7 -U<R<+AH]1:.B\HF3FIBFTNH9UZ;MRRM'^P9M8G^>D.I]O,S/B>;U-N
P *EF8GE0&.@"^< ,Q]W?. +E).5NJ/!4+1*UWX&7C0A7XZ0@JC $2-+#&G_N[A.5
P9B:"EF4?N<Z9_](WQAB'ZSM^><6Q ;ME<10*X.N9SC/R_8XF3FB<>2$B/8RNN/9B
PZ"&QHZ)'EBA=+,X!2%Z0P2#M"_2^0G,!3U=#Y\DAM[#W2A=CRVLBH-!?X\ZR5%_[
PSV,D$:,%RX.H=K$2,BKG"I2_LEB<O*U@N)P1T:W3?EWC2;V#J*WEN2WHT*_T%Q7)
PNK(P$.]7^M;ICR)&C8BB NN:/-^# -.C[4-.$YGZEG$]J)*B/+Z^RY?0W+K"LOY=
PAT<'8X[GIS025S5*K+[QL0 J-+OVZ6JS@']HUBQX^5_T%-.!>VZ= G$?CW=W8A/'
PUG<%SNV1D&V=-!T1\ -GY5QFES-+XJHD2]#VG /6N(J$6B@IDE%+Y#EFC0M&57H@
P,XZ3H"OUX-*G6PJ096#/4D#'H D5.*792?0S-"'QG26J)52YH"_W-FX))B1-VA:5
PVHQ#WL*Q/2EG$0<7U^Z\IUKKXF]?*Z-R-C!<XI9@B0XVTZG4AG&AO*7D3X!#S, ^
P[@/C=$C4N%T-A*+NSO2X/)(G+PRQ!H+D%QH?UNPD,A#IY21N8=U?T%2H(.,:>&1D
P-7#.]V 97=\,UG6E66H\D<M9!T94.D#9@2862U+KJJEL&8._Z,J,TZN$-$1[,I2H
PUFP\'.G4&B/PEG3-9DQ^ZA5#=[%>P)A-E@O,*'6]=YE[?AJQ7/!K*$@@3S\W6'*T
P:E%6'X:[87Q90G*Z!Y;>>^F0TV6KGQ5!$%^;P]BM!3DL)$:=CA8)+!26Y?MQ@/.G
P=MB)TQ/;"<T\O2_+>L4#C'4#5[\VD5D!WY5=C5M>KA_0'KDTZ-BS8BVFVOMV71,8
PX4B7 <^ MF?7B=K-)]^'W"IC<U7 :<3XTDZ&,O1A[(0-CQU/%+@/ 6$X@&DOU,1.
P'AB@W.8%)B<T:+>"!";7,"]SSV*G?C'5 \& <](Y6[>"5,PV2UWTA=$:\7;I@>(I
PPI$=0@-':>I$VX4769Q#6-7T@GHA:0AR&( .[M73:VT&,#M:T;X2 C7P\^N!3B/0
P7;!8?:=P*;0:T(I3@_UG 7^P@H8/]6\)I3J^"3$G&$PA?/:?C=3R*P,Z&EPO[] M
PM.>Y&5Z6SJ5VE#OJ027BVT32- B+= 0HR!IW4X0<,:"S60+MX!GNTL][SZX?- ;Y
P1$,6/9H4$-^V+?_X#0#B72_#UJT0')D$)E10OY/<XKP8^%$S>9;ZM=E[:>EP[07A
P/NK9RW.*Q2E>O[)\WP^MLKP7^ TSA[-Q)8 QB&MV)R$57G-,7*/F V@=C%I3PRXG
P?C38O[8J0P_5RGG-,.%RZ.>D>_"H3Y4HYC+O\W1\.[R:8$W:8D-T,.S0KE]9+2P/
PRD(J'KME11[MT) &0OK\9G-[N.LQY&=QBG&B[&<0RDW_>B"L.=+<M+EN)?0K@A<#
PF?MXZTK<='=(RE)@EP&JN([EV.WC.D^[#M%B^L=:T'*JBHFYS-CWH)>HBD8E+%0=
PA"%"7HE;DH*YJWY?QV?\RL4VZ4/RN"93HJSJ81/+BG^S)M]"T:1/.A\CE.=$?0HV
PKHM#J06D",=/$LA0-DSO:\OQG9C#K2 &!R.Q!1/#JP2 !22A*5S@FP(E[Y4;]G:P
P.RU^65AT3,B4\]1OKMGO=98?N9$V?0#+Y"R-^-;(#\@42]D<X6Z6%V-TT$6:L.8C
PW>L_29NDQ,B28G$,[8<)IG9(CY]L! ]O/U/''86=T"IB&_S"=]"J$XGW\VD'9O]I
PDJE^LF\D'/AM(9_'47.SI=T:B\\BS,]K50@O0UX^Q%7>;D1P!LQ"ZB^NSQ8&&"G9
P$3^:^3Q4/47G88R_N;*)FG/UXX_JCH)=#2&H?HQ9@V0"ANZW\G*[]D0J/!0NKZ2N
PQ..:A$+UI:E?&)6)[!3 VN<W(3!$B\]$L(:LX?9\JP.7#=X16(-W&F<-^B%+!NNK
P<RN3'69CA$7RP<R/A+;Y0X)KP#4=<M#'+R1&]^,5:4MM;YC>#%4 A:#:"T@0DI!8
PN%NU-C0KG=M]-$:7JYRL_@*K(4]RU!96J!NP6:WVH?ANL33S^L3(3W-NFM2LJB5J
PBFY:&]23^\\S ;H)S0XVM#%]!-SIY2\W^I<?1SM 7>.%],_O$1L\VN[!*D7^C%/Q
PI$,:R?V=_;NNL^;5)FJE;"'I1D22/I@G 8R(V0V$"!:^+[XI(['<MQZ>L+]X/I8<
P54?+O:E:Z&73%-4+6CU19=%KAY7D(HF\'_, #<0M61#BKK)3$:&E]W3RV?>70EI*
P -I.4Z@PXC-]\5OE&B[B@AZAD]\U'YGG=5>FPN=.#2E"%GNS#QA"&KSF>\R]&X!2
PBWWI*B$B(T^ _[G2%)4)XRO(<+7*Z0]LU61BI8Y&N@<U=/VAQU!L83<-:25@6W='
P+QWF>,BP(J'/\H7O<VQ<KG\D)=^]H9<W?S-)-+0II)4V#5R::V\@P3 K=U8(6E4N
P.$87L:R]63S&8;/].Y(<F=87P+>4J<# )>W@-SK96.&0BM09%ESS<L6^H)AE**<:
PL1PW8B%J\97SA39!/T<6D!R$G#.F0YF"O!O'>RRM0CH]4E@Y8D9R^$!$CTD;#K[%
PB- @^!"<QPP.6.P2!KZM>^L*WOZ^BD2GDA=G3])4+GR6AHI:[LOC$B:- ;H/]T7H
P\B7@-[I,5Y2:5X0FHNY'9X@FPD+W@2XB-EJ'EX;#.#29-BP;7T8BJ'6;N']#9\<9
P&(Q)3(+\63_3,1+>-62Q(UDHKRH-9XP(CQY$#V0TM&K@$V=I;0'7@_2%=/*3F/*4
PCLT:%#/$ L$20J<!J@O^4,KWHY\N1 * D9K$E96).6LCE6A?K'P)VC+J>_&3$N"5
PX$3-VU/(T#@J+73N66J< )]'W4LJ/,"#.! LPW9U*DX-X9;20@<,-7CV0T3CIX4:
P@7*I,<G[?[HJ,9VCX^4Z.F_<:H9K=F(<S;*:]7KE/ZX=]#+*YMIHH<TSY3FWF2AH
P#E+'$:$$&_-B*?TJ?O,)3PQ.=N@:/G>@PL)H8"]M&8ODC6%L J(5O4?-:94.<0%U
P#H*HT7)W^4P+RX,&F3%_FL )*DFL<OK3\+%VYD%W89,I;O?O*5=[NSE0<)1RF?IT
P*C7FV-,D(*;,'C72I]K)-YA\0PF<N7G@YW#_-%X"I-G&4!18_U!PR%FS3+@3P(ER
P"B?ON_!._AX^;K,^6PR/QY. Z=]E?B@E&="MS&&E6EG=B'51Z*H5PQ+E>0.X(;SO
P7^?8P26D,3W$LLQ8@8IX=K:XB.+\(!+N+#IZFPCANLJ_H0/86]()16RJK],D3 U[
PMNT"X^^6"/4+0$J[T*$-CV%^_7L@E?+!>M#_WG(OL>MB^!(N11D-^QA:$K'TUU@F
PO&<])L,_+:,C9 "B8[-@7E]20MCX0]W5,90$P5 =7[.G=:D"R8N1['Y)@$VOR8:\
P0#X_Y&<\;)J#MF#>M*'PZ ,FM)E,45!R]Q)#>T87S2R@)^NI>/T?;G;[S%!IYK>K
P I%L_,>'<MK\^JD5*WFF40?Q''+8^PZ S#.II>ARR@^=<A#Z$,[RLBJ?Y81/G" V
PP0)N"((0G]_*T( SM0AGBP@AV("!P?*/J%?7(NN)!Q$2U]K16+$RLRL6[DM,T 8Z
P960=*S$K.GQE;GL(:,0!1&FU%+?,V2>U<,-28\@41P6)JK-F.H(XODPY:<S8B""#
PH3!7&_WZM+'!VRAK94]@8P3&!%I%O$D<"=;8),WSF'7Y-C\)+H% C<<^=AK-Y]N!
P(FR3>WRY5VKF-R/4*C%]MG% TMZ7,BPJK(%+RDL([OJ#99/%P4M49>:NY0NSEI?S
PO!- .POB**P38X"=-O4(,GN<\$<V&J"%80=!I7(EX=K/0?N2.WU]C/'SA+ZEVM0Y
P!BLIAP64S!Y%+2\ 4V_%M@\>$O!S^7RV]NZF:5871:7R=2?P+@>VRLCEUS*X$8ND
P%BZI1[_+2BJC]75_P3F9YQV!S>_=X<L&2_5(L?2J'!F7I6W@NG]B&#U!224?E/DK
P\!Z'IG/!:=*_<TK:8;S3,#W?'0*?7;Y&@S0EW@GQ68_QD#A+$2;5#4/0%HRX,PN1
PLMI&\3,X\!=8UC[&@;:-\8_/?;U^.D\P$/SOH.Y?%?;C+LJ\"NXLHBY=PV?E1X/Q
PCM<5)@(-HI8YMOC<D-!I%$O#6FCWTWOYZ!,]S9[EH#2E*V-B<)QN6FNQ(T6+2RQ'
PX6]<N4:(>Q%(,IHVDN;:;>$X',_8C5N_#/-":<<=<"^O7.7@5*(.Z2ZN.P"A[_BG
P)@(U<*XM)G@Y ->CE,*>GVJ6%)M8R#18(>^%;J :]S+Y+%29L.E%'#GZ32?NY@7#
PUI044Q7"-X1K2@?[1<)?$2Y5/X'CZN#8V@2#+#/@O.A)0:7V]W':^%U\Y-2"":)C
P5GI1NV[7-G)LY8ZF'QY;5/#5>;= :H4'Q6&\R-#7H*(QNOZ3-L?=\T<T]R*M"I(G
P :*V)DK([@'=.AM=$.9&E>9\_V&(1%TL8HKTB*4(B&GO)QMBED=CMY ?.MWL?<&[
PI:SUYN@-4>XW>48AQZW) >CJ)9H;;<56 -$ZCP!!";?#ZXYFM+W?6VM[AHD?6(2H
PD5SNP[Q =;'J@\63\!L<QTE#1*XX?6<:9.5Z] @E-F(J%RHWKJS_IX0XI+SP^FY"
PO >WH"404I":_#HVM-@7 A6E)9NB[/^K3E[&G)KLXF*,_D*E'!TS?1O^)*C=&DX8
P"WS)%QWOZGQQK4PSE:81B?P\ZM=XI#1;+W6I?C(O\>[01BNIE%%#'P3? 2RD !:\
P0,1'QA45Z0)_S?7U0D<G[NB4UXILT<?L0$!!SS4OB88G&_%UZ&32&JPO_@\26WRA
P7G*TC10^1, J'?]  P/NX6E8IJ#5+8T=KD@;P?E@1O[!KBXXC:K>B#5TTY>0PN2]
P#_Y#88YU!55R" 3[6VAAXL$(Z>\.,OC>B8X 5?\;&E5N,&#1DPN:T1U"Z9?22TQ+
P!3'PXA:5R.DM+7O/-"H88]TC9H8+UEJ30)G6L9=7FUDVHC*?.Y:CD!$$E\T2UC(Q
PJ<,-"IR[Z22O3M5RG>PS'NL%06[3);999?-4C14 XTZ;B]ND0[6[FFB<!OH:,4Z 
P+NKJQ)RBTLGPLE;2N0.R@TIQ!!4ZTH](XX__AU0!J(E&HBI-*IKO]'CYV*4@M>@M
PD_K^0J%90UJ-8AX::/_9B2CWL&(L1Z&-J!7(J?IPC#/Y$]#W==T<^(Z8>&773S$:
P)J/RM[$]N:VQ+I9'_!<>Y"3_$_**]QLI+-X0/>7S?<#QM^W8O!B@(4MC(?T"PZBE
P"HV"O)50$1Q7%;2>F/79YO"L*4.>]HQTF1(*A3810"^KL?B)R"=\G<+]<_?%?415
PB0Q8F:</R'AC;%$L:H@<:J58:4=LK M%JXU[[OZ26.=_'<#!KG#@T#?D!$QU.0(7
P@$:2#A<D"\4((4EIJO.Y5[P)*8(>OI @"L*3KA_4"%$4V=;_).DN7[-[2.R/+=03
P62?+17!Q;_:$F%D8M54N&Q67R AUN9S_HM?Y .6!@ON4Y(<'C)9& YU[Q'M7S*3J
PH7;T1%8NXIS7_HNGU 'YF[C,2P4KF"*:'.!GX2HW7\<8O!T<M2]@"?#O1T]ENYEA
P"I_LD9(6?P,;E5*#_,%U&Y2YR(:&_;;]]+"I/7VK=8I%]%![&5_Z)?]ID",J\K(7
P*G+9+S=^@(368*6SR-N>;:(!.5&94<^%RNI)]9U4C;WPX7"2?CY8\95,8/0%ARN,
P:\N1-2N%I1UQG"4^#F_/B;5]TU2L;8B\!AX!]$9V#?P"C>:U9MGZZDH9S??U,&@]
P*3:ORN-$1X!$S-(HO$R'H<#7\O!P4-./!J(GQXK;&]?1+7 .:%9JKAG24_Y"">;7
P?7+#P^'1E8)[1YIB4+Z. ;J&C=?Z[]WZ_(*P&$.I[_I:*.9;;Y=>XAC#^G1TZ6!N
P.B98EXKO"$#JNP%&Y\P2(_X$-PE=L_A'7..+/3,MJY]/'X<X$)D#F:1;*D>_W@0B
P8$^>S<=T)%)_0\N7P'P'O\NEN>B^DC+/]-7P38/=2S)E9 ^I/2Z(-_((A^M;.DU8
PCCK.Y@ A1J/KKU/N_4QM\X5DC!G0'D,1 H/D[R 7X9?# 3BTLON8W_GS.+D+$+M_
P95&?O&0+ 9J/J8WY'P]1Y8YKFKVEOWF8.K4U!_QTJGTE[Q?FN(<U2WYK6$I=WO&:
PX,.HB^7&ZW9!JJG#"(C1W# YYMJDG>7.&_4'--E?^0<OP#BT+4W?,AO9*VQ1__@_
P&]%#145"EKW2DMY$V1[E-J+^1(YX.N3D!<P8#8VH,LP.6=4T%<QR 9$C!!$VV?L(
P%F\5 N6H0C<=.^O2Z9SV4CCMPL9Q7K&[[9]+\;9S#O0;[72X1?03L-Y7BC&F6?A&
P1"I+')KYP<+R*;[0-.,%+W4V"%8   E!JI*?.3@O$Q9*735^I=6 @4X#;ZG>F;U)
PR!QX:[WEB_F()BQ(K-<KCYGGLQ6.DC4.OIW2,_\U.'?&(63%7FM@GVQ[1[/;]^7>
P#;^PP[<&$SYY&.S5= VET5K_P-0!SY=.9AHH:QEI_G9)'H58BG-O".&<%@-,I"B_
P.#DVP^.KLM0R-($_5J-NG\05+MZLM("0'R<\G4^I-!86G<]' U_70*KJ.+X*I?'Y
PDS<6Q E"_.7 ALP <?!E0TIF!\@AW\[A>%@.N^>#VF\O19,Z3W W?F)F;1.>^ZEE
P"]QCY$:6Z,G[D0E\'+"1S-5XF[R#&8P!-;[9WU!Q6.\SZ<RVP?K_+>RD!L_-'\]+
PQHS*?3\.A@+@(A[6"U"7,1J7D1AO(4[AZ>,[!QAMN$NITR[\ ^/2@U9==$SG]'16
P 8,<&E\7YC+*@7.NGT8%N&S#T(X5O1@_XCW,7X2@H=(#M?T,BY' EC!R!>=M+6+P
PC@)B\8!!QKDY084=Y3>+-2*ARQ0M-UV=E5AZ+E;M(0_00H8&8PB5T :_2(1L[.]^
PA R&Y^I$X\U)U+\R/4 [J=LT',9$,)D1HRTYU_SOAJC+-];K15<@EZSC>(/BCSF5
P_:'[\, SA>J>$LN>99W[-Q(@5[4V"ZKB2@:._H=]@< _P"!BX(M>F!HZP_PYOH[=
P?=B"5=*+ 3T?J[K<3I</)/IAH^(-2;UV@#%5<;F(<$>O9TTO(LK+[P,I 5W7$D]:
P@% !T(H$^GI%H\MB>:3',A(?< >NW3 [S"G+FN?U<0B(*B4CWTJB7\=MOZ?3G#Z&
P3A_NM7M8]_#FK V5E@7$SVF_?4,3&]A1_R=KG^T5#VZF6/N7*-H??F9,,Z9M'33+
P"@S9C,LN&4)RQ@1UH-O0Z$T9G2?LG2K2HO]0D!G0T#-VQQILQL5*]NL!YFSB--+)
PF+3%Z'!PQ_T58_D&XGR^/_PK/LRAI5[)._Y)%F()! '/<-X8F^T7&@#A3B/6UA<N
PH2$,>>]_0N#BC348L ) H+^7QMA[0=<6&3V$YE.;O#[<U':-J4#[O/U1>8=VWPI$
P[[[;J:NF!X;D/'=>ENR?Z)3>8II[^YP_.**=T6/0<C./4NMSZWUA2K-&+57J#[-@
PL!3O"A<)7D%#$AT>@4%8Y-4, LC[3G)K%N)6!]-D2IFAPY9H?H0ZD]TA^MH5,&EI
P:)9,ZHM;58PR=Q=%IBP(_4S$@TWR*5^TEO,@>;^4L@7 M=Z@(&</-Y]W. M&7T;8
PNR72!=YHJ^P@: E>ZYCI(^N3RG\KJV>WIUTG=)7E"N?$ZXO Y%)NGM)\T^\$*-(Y
PO= HW+Q_/K XR5[[IRH4Z@+=0/+Q5"*;$MN&S%'+4BSNDX-^L!_33. A$+$_DQ,L
P\O6B,FVVX&[VS-AH.;;GHR8['QH_Q.T!5*(^>(!!8BY ^*OFI(1E5/=3*?W[P;]]
P,:O% 3M[1;&(EQ!\-#_@9Y4@-;:TWE9)P3<8/0\WRTTV/!8IWZ@YNB;GT#@I+7XI
PN>FCW]QVPH&VY8[(JE)7U'.*L2F4X&@B0RFN58\\*JLV"MU.\ZKB]IE(YA[(&_V,
P.:$&1#-I"XH<>.4L0:@8[R0#;K7T R:JAA8JN=\+1J=_?+])4S2BN@75B.G:=&^(
PQFT[^W3O6U:96@'[F<1HOF)>=+.\KAEB&V6)Q:'E7BTP+K51W] L2I.EZUZU#Z6Z
PW!B([8(YF!=UX'!PD[X)$.EI\BHH>U!D!?*X*CIT^"'-!?8>I#=%W4Z,^70 K,T5
PZP&_,@)[)&PI.U):AY=;/FQ(=J>@1-Z8P8)#0D 8PM1XW4H5!_5F2H/7_$ J !^I
P-==33(#K%AP]$<)/,>+2#?TNPMCS5P5WMXMI&<BTBNNCUU+8(P/".KK/Y=L#TND_
P0R&F!^STM 0(O)NO7[<O?AP?Y(D-"<-) U;M9:Y$6.5)*R&)EEI9-2FU]9S>P/X6
P:$T4MB>K8MKEOBZ/-XMT5*.-*;DU-%"U*.B.].73<23N? X8::\ZT@&!RW:0<2CW
P/1%D8$(?@G(R+SPA%>E$NY8SX$V]P0QNOQ=EMHCTLW.@)<W8U>+1N=M?SR/(D!,Z
PWNN4"K*8QB:/C](PD$)P\?AF #H",-3C2-G=CKU2T1A8"-G:E[U3Q%E@@P99$(@9
P>'!EC!C/RD&(>DT!VA)\P_L%01'FA0P299FD(68)1FP%)VEG^LX_+VNQV%>FV ].
PU*\JQ(\T[5V-_=IETEZ&XF8DVAQ8'!% Q6?L=WU*Q"TDQS>1IOCM,:(F@+BCM?3\
PTH6<9:>CYDO&QC>;13W(I3Z<K5O?1.(AC?2P:(J)7+;X/^XZ7['7WCF\$@Z &;0Q
P]YMAI86MRSG?QP*L25OT[29BA(Z,]R<BW=21/L@PTX +5*"6&Q="SP9\;I4&8JZ1
P!@""]+H*DK?\4.7RGC#4]Z^^YV(OQK)C%'1G!O&2>CY1P-C Z (/0%R*L+_1:2&9
P:A#<B=U6/M!QW^5*IL&$SC0?4$!Q_:^JQ)&L'P&IRZ8<$+^T8"X=->S0T?:UXJB,
P/'I'CTD^Y;GQ7\&2TL[ _RBT]])>MV/@-9<T)'B/3)F0-JD.HTYN:28@<X3173;&
PM1CN[$&3K.96%)_GE95ENF%!,S D%"V+I:5M?B_*8T-*# UT"9$;0$.!"7:;>]P(
PJ%&*;/RT(9:"]":K8G,D^M9? D'FDJYNN!Z$W0XNE?0&&]]9BP+)<6"#EM1%]N93
P8N .W8RMM1I0W18_B;Y0XR;6YDKLK59P9(*&<N(<4D3-FRYJ0PX6]G(DZ,AH,>>,
PPPV',$%! >7A5LZJSZ)I+3RM"05"PYQ< "2.VB$N[%3>I:30PO]L%U@ATM'#;$=0
P>PFU]1IK/>T:\K )'+>2P_4BP7P1W\8G(9ENL%^,SX=DA%LD]S_N!O=J^Y.HO#6;
P@,CE(P=&V/OYWF=P MC6R^C/Y7KEJC^;&BRQ+ S.G@9;PA^M?7]U%B'2RQW,AG#-
P;QZ(AW]]]<CZFC7,A=S%SHWT>*;,+ SVY(])>['2]&-&1S0-[Y M"ZS2U$6^MR*6
P)_6@ W(D58P8 ?UP?(D7?)BOIAC=4S^M&E_6)B[*V4JM9ZWYS? 0'4&FC1RQ"EDL
P50*^6I8K8,BW$M]DO]\,4C 3DHFLE?4'2%Z)$G]&2-C>G@>BX5!H-$Q?+U42S5$U
PLIR,P%VBR%@@/B%C\E"4L/R8I^/8&92P+,>(\:JYH9UOAD?:</YEF>T+S>=05"F[
P;#PMPE$&A0U&&Q>/(35VS71/$.WRAA*&:C,'9+R9U_I2_"Q?:V1ZU[14GI(*CZ/G
PF+!%'Z7@A$1+J@1$MM7!4=6&MU_KT+*7&4'GDK38+>8CJ20X2I'WTB8STAJ?G]X0
P@70#!D8#)IVX.<+F0]5322=CQHB'@:*[C,IAMT]OY4^R7M:*%ULU47E+=/"QW@ZE
PS]D_3J.F!450L859\M/BQ4S!!<L5C*WLFN!;XJSQ_71(:,N,-C/P,,0M?_6O*F7B
PS.V[8GJHR4LGF4=T0)J%-#$D[LA4Y' V\SB(+ESBIH[$2>R^C51;P7KJZNT.-U'6
P_E#!5[?+#K/OX@(=>4I6"D@IFC[X8CDA=/<D+K/E^3 LH4^+DJ1,;D$FPZA$!2>!
P=C_EN:B1K:?([A4)D@PNUO]F6")K53KI*U/UOX_ W&W[I0^=S2MS>O.DO6C[=\+]
P*@[!%&X4V-74;<;SZ<C.L1A4W7BGLR%!=:WV*M3 A.C]PAF6Q8F3=\RCN*E3@7"L
PM,C^!'W%AOYL9*+F1++N9LGUL>5DJKPG"3W+!?SI)H9#^M$AB[C-P?Q[']4S1A#*
PRLZN1AF,O!B<F =(=[9,@"3";000"[YT.&IPCW<I>,:.['7\]\[,ZN]/^>\6QV6;
P2XBAEQK%XI<%6\@!_OR 2H-!S85.(BY4C2A=R'IAXY#\*_6"1 D61-G4\5)[*/#C
P!<^"T$A=,HD#DS+V**1Z%+K9:MIA](=7/\XC<*\_B$M#_&E8=+8EWN>1.]%2<]Q@
P/R(S8'U&I247+]WM,9:5+_:1 L*!,1:R^3QZH0+!:),-EY'R]E8H*N=*$.CR\,U=
PL$^8*#?B?'3^=3C181(\=]I$*%>TMT0]X+=4>3LO#;E_R7D3*.5/U@_]/&$*QH]2
P,NBN<$+XS0?&VFN\Z$1S3R'?\BCR'# C^&! C:#'KF542..$G,8R=5K[\!9;PA:=
P<MB+;2S?$&E\!/&Q6PS3]G084-2Z_^)OM\C"JP(-)*?;GC4&\G!+;Y?M>Y2-IAS8
P#G^:EU:)$LES9R3FQ+*3I$5SHF90!LA&\9>?.HUX$VJ,(*(N8<S6L!STRI[U,.AV
P\N[/!0PS=/J>#077-UBM->+=0Y*/!Y)K]^9.)Y99% [09_K.*@?]U2U-!9D[*\Q;
P<PY?JXAI7O]:9Y*884B%2'QKW[:]#5UKU#FM-HZJ#B88VRCQMT[E8+N&MDB&OI\F
PF[DZ#D[2;9!9PNDF5*#8]\1FUCHG.Y"6]H4>3=M$)?/$!SMP@(,M%3H39DG1TE";
PM[Z1"A\,-ONQ">IP<'::N.86.=MEIZ$,,I/A*Q-RGJ0(\CAK>0F-REL,[C7Z<7W\
P?Q)E< %JZ&]<VII-*KYGZ'6&D+? G;_"J5S!"\7'[(>Y+=<=R&[G\_H,S.8T=U>(
PP8<R;0Q*6:(D-%VIF#C\]2-[3BET<69(&AV0<,HAA /)CM9/]^H+:%)JZF1U)H-'
PJ/TO1+\#]^O*A(UOY%/F4T+R$_H")BXQ*07S:K9%MKM%':UDGWU@$;8JH^?Q((K,
PAC8P0YVU01G@27= Y]U:DP:F=5[HV6/Z.>\,/ '#C'[ZBJ@Z6Y1[L#.ZXR %%UV*
P9N:>$GGD8O9?):+?<_^8RZ$$(QILN,P:UDZ]#_;[R3C/0\XU &(_W@ RPF1YIUU1
P+'%Q(M$=++ZZ=5C!W[)%4G3A$ E2A&U)GP:7!&8G9]99H=XL!B_[=M^Y:3JLI"F^
PS;D2WG$-/%EYWJ1YT]^D9S8=:%P4[^7?CBG+T/_Z=V/Y-.2+.0R33-O?HC1 =4^K
P/C,^G308 Z1$-;4/884P7:(E/*Z21K<_@X_IJ)^+QQ:HDCLX9":U^8)P=VASLO/2
P#X2[FI5J<I#%.<5>KO2J_T>;;\IN/HH+575)']EH"'T]45MV?D74JZEMLM_^E<N?
PI[?HT#I2A8<< (=^FC?!KH3O13&\4B(CRTWCI5@HGFJ;(=DLNG2Q=U)EDY&K=H3X
PF4;/"9 6R_W31@/'P;@JYO'FD*.6<;.]I.)DJ(7TK!$U="YKK=[:E0YHEO3>":%E
P1[>):;T^CR\WMD1HV].X3;':.Y@"!UL=TY'526[%TBEI@"6XI/4*KH1< ",29.4G
P*6N&\OS($>LLU&92_HI8,4%D0H/F4=O*38GO%J$>-+O=,VT/KE^<.T;)-63FP"WF
P!8/B0 UXSNPUL[^C21_XCZA&=X=]VS0N\Z*H]#SCYU7MJZ_3 Q?9,E,'S:4=]8&]
P3Y+HRA\;KW"/4J)T+D9<R(X+RQQ9?^Z3=MO;DXF&==PGFNU?M::^U$>C.I=OE^ZE
PGE0(N8LF7QE$!O?:5D0GJ,"Q[5<;=N!II0N*>#]2!U7/&%*!R"RFVK-98+WQ_WX:
P7LIAH>UIFH@0?KXQE3+CG*,1G5K!\"GZMB@(DZY(YZ9:Y"[JE8NEZMSZ(M !MIX2
P'74R(ZX"*!)1.*4S[[R&I:PLS!\KVZS;SI4ES=+?R7-_SX^B\C&)3!%HK*V%XC^'
P"'R[-A4[3T<BY?2<!:7J0&L8&?HU!(&WNPMHU[?2'KF]>S6,N=N*&1!;.C6=,ACB
PZ*STWBR<6W$X@84^SXOH/09/=6$VZJ%C7 MP7, [C)0Q(*[6]GE*T4\F 2M0E2_/
P0[VG.XP-;B?GXT2F$"&?R(%5] ^) SC1I//CIWZ]+)@05I[5S!U,6[^&5S"#UM,&
PZ1I%<*9& XZR,#*]ZE,W(OQ&J"39L.VI:_OH&UR.<TX-"DD['HILOG2.XP;9T#QX
PUVS1Z;^*O-@ZP[$";YXB/FE%T$2#YCK\2'_N&!8(H/:[%^1=.I59YX$"S^#*E&"X
P26RPN/=[K%X#20^)A-HWBG#;!J(HLH=C37.XJ$]7E% 0O\$%K'82@0(SO(G;ZM4@
PF1:(GU3ZT6GA2//O"3)=\8'2:B/G36#C8HDO4U5:W#>\H , &X"9$62J329&]FKX
P-SSA1>%E(%DC[F\=.5-&,V)M1/7&$IXU.9T/$0CLO55^R)= BDVCPXTU90C8LP\)
P=(!)0?H"[@;70/4/X+(71?D9/:Q.74N1R&"0509@4/B/K\Y5?N?%5KO+\F33"J1-
P<WR!'1]%A).6^/:O#J]85*RN<EYZ[699%/;_^Q P-U_EQ/"'\R]" $>F).BGL'7:
P0A._.YHP1>:K?1*!\E-Y#:R5XML<:!;"R>9._4YXMOW7!PU_.\P35'J_-GA0=Y(&
P/8*06.SK->QMK1*H&E6GD-MF;<AV7T4>-$R]9YHTI#E8^3C< <!\X*K:HLB&?XU1
PGCT +3\^5<TAEC^<5B>LO9(I$$4MFFWX\J6YQ -W')R@):&7+9+\*ON0.0B^C!#9
PCX%H7='$4\F,Q&]^',EU9H!=3'6T>Y&J3=;O#B,I/7K*=>%@P"I?6M47J2 L0O3&
P7,4<.YPT[VW2\]3.,%@'7]UPJ_"E8\#.+@DS1&GC+ <1X&U!-^K?YU"S)T=AZK_E
PT>YF)O20!L='4R217U7,DXQ:U4)K6YL#KOK[HA)YS1#-JX%__4-XM1UL6;)>?E$>
PL/>5$:QPEZ:BAQ14%Q-;*_QM:Q#_[9W77@YS3,W)@SLMJ9>C% F:O=IV<4875X83
PPH<F(@^DE8Q\#MFN:LC,2L9"[8DRR 9?K"UV?->%/.,,EK%\.SL8/1BD"C'W[3D%
P]FKE)@FYWHCHD D5?JUK G<*?G'1I&X\XN0P8N9C1L%Q('_!?H,J0BE.T32=M==^
P,G_->S*/'5HAQ7?4;:F*Y>R)+[,[(KX;B?4^B0*V\D$"'087B67K[&^5:.4 HI("
P'2#@ZJJW]WR?6.GA9!H[V280_Z \,Z$W^WW#H<8\3'3>I#XS[9X-]>\6'PT'%0NX
PZ+3I<U?1$*PD-2B\HUPC2=VLR-":3K.$6?=45@D53YCRL:M:&>J_-'?(K?_;=0'M
PL[$1OOM$;R4C56&#*WL>?P#A3#:'O62YD2==^3[YL%8,4+12 C3L&8TTE1R,_EPT
PC+=:0XU_(#_9QFHJTGSN*SSRE>49(^KDF_5),6)C2*<@:3(2T%^,AAIWQ=-CPGI3
P.QR$@TC&LA4+VA$MOP'C_TK#I-%Z+*1HWI;W_S1^E.42'\<RB#Q,72D$0<_=D!FR
P#.6(#N+LE8E?X%(ILM2$ZA^/V]<\-15D!+*DC)"HLUJDRZ;,#&11#GW'_"O$YI0B
PHS4%8^[UM)R%GL-3O1/-?L4H*8^ W*^^307M.=TW]B-=F/XV.2^W\:ZUUTT=QN43
PN&BZ751C !,2F#A/[3I_$1Q'+74@5<QX1](9^H'V(XMBZ"MHYX+RVW=ESF"$AR/+
P!822DY^%-Y.@G]"I822<B_W2;WYE<.:K1'ZE]*>D#"(4X30%06%,3!MX<^Z;\I^O
P;=3K$B ""$HO[514%11O\;6$UD,A?P6%==1"CBQV!K;,0M9\%.N0-IE$>"<QMQMW
P&5/F/S=7AT0'T+J.6.DX/@C6#M,(-;@>@1@>0,%E#V+(O8AX^5TK;%:+-AMJ@L,C
P9&)?Z;):.N1D52A62]G<!X99OO EV2]15(0UO7J/Y!A)E-?Q)6&X\+5!L*Q5^S\V
PB_=FV^&%7Y-B1T(  ;WZ@(]-&9]3'9UY1X.BY5NPF"#AUS@5=8J#WX*X?O!"?>B(
PQ$3^*+$4] &CF9$&*_U@3'B^=](C_N'D9>X#<KG>?S[S\M&0NP#]>>@&>-&.!3.\
P: W<#_:H^M;9OKS>8<+ 4=0Y1/@]O(YYX,N/"C-^,>FC=^F!A20.IV7" 60B:86J
P4K;: D92VB]QC;  <XL;^%2=4265OFOIDC-KI=5GFFOO.#"]I$),@G^[#:.+P0YP
PZ5^ZI,K/\M[;:'Y[D R/^1M0)T;76L!?T(.$B9\BYIO_1^>JMA>\V$*.><%(.IF]
P-$&+"0Y\<FG^5@A-!=OH08ORYK6AA,JP3R\XC<9Y AI"LB0-PG]Y/A\4 V5KZH^(
PF<@L3-S<_=T*F%%AX[5Q3ZFGJ26TYL307,GJ[X&X=!PC;J/(Y,:5E!+@$)0Y;I'[
PLH#& OFWMVG<9XP6GY=Y]O)2!Z; W0Y7AQ2Y1MQPT%$H*<LA"UJ<@SU%5KT7I&\=
P(M6E>??E2U,*4#E)H*8KB\"25V/WY"G?E>KXS2R6AJ3#4"'M/YR[%FC+'R>",Z,L
P:VR%7"'[_89:#/+,TD</YAH]UMP'9U'^FP"9E2A.7QC/$.?+U( L(LB+^XDQM,S7
PB(6;=TNZMP8HP8BB$VC(0<]/1BFLGC''=CV9T@F*8T';YV>N+;T^A :!!E/FH.S<
P6V*SEJ/Y4P:#<=Z+3H@/F\;\2[=,R;K> 0_'UD??E+" ZX5<4V!P?TT/%'\XF&O/
PT/MJR[RU?L#A%>U0ROC\T[9H.::;GVO8_NGB@,'RR=K=G[>9A$^VZU6RLE)>#H'F
PS('^)8%^<LX!L?*($>X8+<1K91X*L#^[]+9$P->\@:4,H5LUY$XR%S&=JZ>8*/G2
P6872R*\?3Z[L%]5V5!>5= \P!(GG>;!GW+N/;@M>Y2#++P@/GEI+]Z"RHKM=EW$J
P! B^(/%N>E9T$?D+6.+/_OH^T+C@*L"O3^>.$[#C(\(+7O3NT(I%HLF)/D&/</EB
P4QDSG6&J.UF9YC*KNZGM(6&LD\%^3#-N6C,/P[DSH<E[/Q)M/N)LN[L7>S#7'/EX
P,H =*_Z3B@(S21S/;R=D<)0S\U+Y[V(8D"_9E(@+6G%*0&C1=CC75H$[!'0.B0A1
PJ0&G0-[$P,S]6.CH;R"J'4M D\BI[=Q"^VC0MR9_@2;YH6O+./U/>@X?7=YA)U04
PPDC7+%SXQ6%KD/##-M08I\MTOX(]>@:N-^YI'6$DU<<$O/J;FHSQW.Q<2?UZ)B?C
P$5U!DR:B[@*NM.K#7>.D.2-(P*6$PLE4E81$9IJN@@GY+UT"-E?:[.77.><O6\YA
P$E%1>;W0&M^0]0X;)P]L:8TX4D^)-+M,.0JV\KQ(];;I'6@T];,M,0^4I[=W,/O"
PD;F"R(2XK%4.6N]\H*+LM9S2%=*:(DL*)*P6JMD+N">6CST;[B>QOF'%Q'B>P7[D
PC+'WN\\]("&JVT3>O#\\<CD5-A)G^>8Y4P:#@[_,+2TS[AV^(3CA19B96SD93M<N
P)'^!&R2E'GXU]I);7%<O1-#\JC:0_Z##Q\&8_9HM"^!A1*1$37P1XK. "[$L?AN2
P_2=@18-+,=EN<+)"4!%30ND:':?"L(>T$\[+C'Q45_91B-O=BM1"4C+L3>#5!VD,
P3T(FYMXCF@%L>VO;)KX;.XTW$I%+P0*D*FZ,4BJ3CSI<L3YJH<HAJK1!F1YNEBVF
P=+C,N?*8ZC9%K6-M3R8,"MAQ^_^3+YQ&_-:TR+YLNI4YFJC9$A@)EE6HJ3&?<H<(
P@[O)UT7JD(P5FG0=DZP,:XY?5"+"B'>#7^!UKW9S7.Z^J9B6R2T[I)IFG[E\_!)T
P :2KL]LY2GY$N/FA^A4CC6RN)^6 6KYGWT3Q3%/.KN#=S9%TG/+*>'B5.R#36+Y>
P-;<U8-U$''Z\3O?9H8]E>-CMZ2GOC.5P24'XD!GL,N^8#[\*L]FYU<)J,:SZ)P2F
P_I-S7G;C0R#7F%?X,$%C;_7X8+!$^_F"]MGO'.0/>+.47[@7A[%.DNCA(3P'0B'M
P5R0W$U[C.>TE+)(\E:&%![@&QGEW:IE*!"DVD\0SM%=.5<]5"C(&GZ![0N '\IU$
P(RVE1^3"1E\Y>2N OXP^MV=CFSK9YI=<QUZ#5JQA_:W[6P]W2-<M@*!8+6B O=L2
PQ!]"/;=Q.VH! ^(>8V=?J]R,0EP;9?5^C4;MB\:Z#&[HXON(K;FSPO[JZO I,GH>
PYN]B0#8C-*V!'3P5 UO?RE1SH^^NQU+L<FSX6V?DQFK:$LA T <^]3!G!(V<A:$X
P<*_;1F*,:+.8SS4FN#)],7)@7'<_D:QCNV)?9S3\\@DE/@>#AFG[FS%17@Q<&-U*
P'X(OC/!BP=H09>WGV9D<1XAF\+L^_*,E](7>Y_^&X5N I95O?FM)/9JXC )J.N>$
PAU-G,'8( 8B(PQ(XC5&(7I8G_2#'F+&N*'*L>RVN"5[<(77OFL&0K3DJ*:*J2_V@
P,@U=Y6^W^X0WXYFE#:M3ER<X^?:#_C5N4>-*W1!WFJF+G ,;BH^SG&?WMTR"9\&\
P/)=_AZ80V<4V/$;G*^67#1I02V;TT6*8TJ_EYDFYKB@2C#@.DE+DQ*J=6^;BSA.[
P:2 6D]M@0*/MHZ^)6P+S?Q6^.0#2[::P,_3-:_;:,X9'2]RXX_\;-ZR0/[CW (G7
P3&YD+QCK"2C1Y! F85<U^FSHLSP$I8#6C]HV86]-#:A69PE<.A-^@]_LEDAR5H)S
P=J$HTJ_EP9ZG^V,5G775*BDFWFKK0NY;!RV'Y$VDC9;$%P8(V+-SB7V_S,9(N3<4
P="C>GYW9%O(J=":T_]Q-!"H;1?^ *0MD?Q#EH+[NL?WV<:+\8RIN0_7.3%67YF1N
P3SYK,?X;#9U4:W!32-<J]8J!;X>5(QD9:/F#3:3S0<5>U!/7^,]&*Y=E8#+%&@-S
P7=V))%J>^LTX4RZ<4CJ*T?B+?RN[M_JQBEJ]3/>PM$HP:Y^^$O&.O@;O]4DY]J*+
P'?WC"'P,^P2K^>T,(@_NL%3^3\9O(GAEIEVNA!V9Y.HL=@)!ZBINQ"4F$*;]DNBE
PY^KXF$+=TG*15T18FPW':JATF(ES@.I8 V:+VM,M::RT8?C#=//+#IRR:$2^0L/5
P_W_4)T)XW,V6J/0<4$OU>X8_Y';M$]9\,F(F,\?.NAFZIT^KS B#<I;A2%39JW+,
P]XBKR$*VD;F0C3PD.66;^T)F=#;??<*/2E\.^7.$?+6C+D UAN=C;5V$D6ZXE$A4
PB.4)_JU6^Y@&G)K/#6=8 ZA=U!#80D$XB!0^@#5$^I:$^KW0V]GX7U4*OL>B6//8
P+3<*V*EZ\>76; X6SHJC*DF7M<:)E)U.;J>M/RD0TC#7+,A9X?!UV^TJU4$H%E_(
PG'64P@_?]9Q7HZG$-Q NS8K5]#9B@J%Z^V+#G0LI:G!CMZ,/=(G$7]IK4; T)3/?
P7:7P*;+3M.=DT;;NY!LM:AJ_(;ND0IYR2-$<8V2P_D+0PTDC>Y,ZGZ2#G+'P1:I5
P?%@#',#(KTW?VC(7VPA><Z)H*?=NVV11V!"[/B!XB/]@>P%=F&DP2,M4Z5R(T4A@
P&4&=W*.Y.T3'?$(X6('>:YBRHI<*6K*^\8V"8J3H>,6E 7,O>DVPT*TY;^^CM.<]
P&,F^H,[I])+QL!E:3E,HO-8FKVEJ$@/ZZ#.KO]0LZ[-@Z5EVE(@JD9ZL)H'2TF3F
P,3_GET>L4LG]_YNS.GI#C[68\E#X@4ZU=627,TM^\>D+V6OW)% ^5=F-2%N_?VS1
P2VL4NZ!J36_:[KB]E3..8G.D9[81<*-4OU"W%=H?<'JOPC$]19#TG"3IM0<9S;\%
P*M08.>&LVE.H5-H'E6R!T<9Y"<+[&(((>NIN6$FC%\*X[3Z*S;*MUWWII\B$C3(@
P F,Y !WV/BJ'@>,&_=5F-HX&$2K;1"IUKCA[C0'CHT]SE81DJNST2A$M,8'SDJI7
PK ]$6)3<EDP-[W]UM?8;K]#6O:F\W;X<1#O?.=Q7\OTCXIC%)Q==N"-@2JG]5$K 
P,>!P33G$TX;G)^2BT*G;ZB,5\,@_C)''XNG]"!DRNJ.$ G%62!-2/TT9.FA2NLAF
P*-^O[6+"8>A'!TH:4U!.?,EJ!:V*6,3U2<WA&_*LQ4]XVO%DD2PJ'L:CYIO#)WAA
P<IBN=3:M5*AEK*Z)#,%M"#XR!-KUT[^_*0L(JK\\C"?>]VAN*JX_^H:C4LAD-M0N
P)896R'\QNV._!;[&]:EBSP)-20,%?')!'(;HFF8QG ,=L6-[]+:C?4?9(IG(@:6I
PY]M)>\?LBX5Z%U6197&-V1*NE]4)2^D*Y C*HLLG \D5%Q&PR(@RDNS9/TVW(1WY
P$8T XR!*HY?_H\ILKP9F/.O0C.GZ[0UFJZ!V7S-"?MJ&+6JB?GCBO]ME[@F537XG
P+I?U^7:#:KT55B"G)Y<*<5.."2'H8ASXOB\"IM!D)-"V8T#/*E_V62BT+U3[7XZ;
PA38I1;?YI8PB%PR[CGZBH]0="UI@;3G.JENC](/H))G+\*E+R,PG1+<W%,PHR:,1
P=-Y,0H +&0Q97Y#YM>S"A!5EN6'<CA0W]?[[$8R<XF?V;R%[!$FD=XWR&H)LJBK:
P:(C][>M\<X\$B-@%6,0XM@;T"1^3V%T#J^P;$I:YY R,)6X0CA8YA>5:3. @(9T7
PHOLHNY2-@D2G7^$*YF0!O^G>U&2<+$_I.,LB-,CP*M]E;=BDV]O2\H]PW?5 P*N 
POT-"@%$9$)T10899?ZG8$X ^YU_ZNWK9.I&0U[70(FZR>_.6[Z/@E=8B+R&:D&P#
PM"KT.@Z[FK(-]X.0T@2;CM$WD_=$QJG5:6<N%Z'C]3<4WP2!KOI S3Y#.L$_P>N:
PWUV*8^7:4%15'8^3%'0::/NQ?I1,,&:9N )./Y.VLR1N)G$$K8D:7G/QS(D\K^91
PJ'H 6'Y7J-$#>';#ZA)L_K+W#FA%"Z8QFQ@41XC.*5.\@5: )FOM?S.&CV2^N>;(
P+7R%H=:.,_S95.JA<C7/10KHOG(E48Q^F9'NW!+=Y,*H!2,(P(9FR<ERJ#3^KQ/D
PU'AP:*BVL\@AA!N9*"CPP%6! U+<28@-7\ 3O"MELPBCR4X5T!R, _H&C/-!J9NP
P=U3C]*/ 9"4]?_(7]CN)%KEVMQ(F%];<JM!K*]6A\O4[0PJ-JG@%BQXKO<1%$:/W
P[,!V_O"G<NV\=8*R%L.;Y5E2?=>@[R/;A[M@I,\)9Y0L 4R)I>4-P/P-<[H++#TU
PMB(%2+>='VJ_0D8LV.+/(WA1Z9EDFDK^FBZ=$ +<O7TCC],=\E8*:6.1Y*J!34-/
P=,?I_=@8@0A) Q$/38;K!ST&81K%P;)O6?8Y;MMK0^TK%>>9J/F!5_Z18^D'3:E$
P"<+UYX:Q71CJ9HIH5%&*9E-$T?_A-;F1AT.X<6#@)3@;7>O-6SV.;HG#4Z0M8 S$
P8)7ERC2XE9<IP.V.<[(NEIPSP.=BH1M1'1]),@#C4R7BOB+!OK-XR756GB&N\0Y'
PB!&$(:QS.!;(XJ*WQ> .2_88;GPJ;):7G 9)D;3@W>1Q)J[KF0W6!)5F8<-G'AT[
PNN86@H5;IO"S'<)VNM#+SX6:PN.YU*N\((.*2%>GS "W@]IRY0JV ZFWC*,^CS-4
P]SVMS]V1SUGWJM&1> -[4O;YO6%=4YR'0'?:MW<"E\I:O=K93Q2_PF^K)(D]E3:X
PP<2J5LU1^/L#9P@\N2/'$)5)&_&V$C2#T]*X(*H<K=ZW=V$8<YZS93]$H0N)([(9
PY3UMPAX[-@0@14S<>RI^/XP GVK]%KYK#CW5 3M5N0+LWOLN<-0P.5"WX1LKX&+X
P?'H@6.*4;S!7';(YG4,+R=( +D/J8:MF4-?%[65;>Z>X*G+8-A^&!(HRO%7(L#5O
P(&"*J"9&9SP#8 A?ES.JW(F?RL\WS;\;2QEOD(PX1>OC*%[UWVAC^/]6IZR%]4OY
P''%0F4NPV?I<T%FC495JH+705W#H5.ZFDVH.1M$"@U5JT/B&)-^R#1^W8GJ3&05K
PR03HF%9Q.L>NN\#:]W1[@7IYL R&NT-7*[\,%($80V:#;Q"-;JL\24Q4$R$:0XQA
P7O)SFC-3F/KSYM'_0=:66215TPWA>F$Y/&_N3XK#LNJW<M@9EM9L*?FUS:H1?\E7
PW)>[FG(UC&[%(%CZW%5'Z]C3.!,E:\+5$G!Q]#0))['/J'R521^+^]/' ])S-M'D
P7H4]/_:GEC_?#O;H;&V'J<K.Z_/UDFQA9P;Y=718XL(F9];.RF:<@IVU>FIT=N@#
PC]C(C5- QK5D40MFR:EB;9:M7B8QCW6GLK5/Y7[R3N .5V'^QE+C7FI-PUZDI'<:
P>6KK_898".Y.!!%<,0IL]%,/-;&_RG&3?&]DQ,7RV\T=.6"/.'J(Q=*G_:]ZC<3[
PUN=GDZT=-@A;B"=3=B60J*R2T6\KW=U3[VC2WH6(Y-WLQ\#'Y-+OG(U6X5>T*@0-
PD;>-:V^OMT6:IRY?5'S.C"(@[]*?WMVHNW=>NIJK^2>\AYERH<Y3.V-5^69(HK0E
PV ZGYR55*Q2&1LXZE-U2QGL&7VLP#=&VS'M4MEW\.IRC;,>^-8\&NN(_(0SOV-,H
P%T,?!_?A;F%7UV.%_]H;' N%ISYK"#D'&?CUAU&\WE-V^#BR6KAA=]96G5G.-WG+
P9><051ZS* RIR!23;TEO.. ])USD/7FC*W/9D4@LA-7\+JE@=8N[ISW\%C_$("P]
P(^X]2Y))#IG .8,SA?KGN8!++0U25 Q7T@_9&M(?-P22+DZ[ZW6YZ)__4J#8DF]R
P#GF?(RI?XJO:Z-6W(7_KG[,$'LLJ_0^AKB34FU8HQE*SA?(V.O"S8EZT8>(_,@-+
PN<55G\1O*EL7,B7T[H]%7<5&F(\Y4\(%TY?V^[YIV"-$>$ 6O"H(Q_=O5!4TWU#R
PI%?0=:XN8NC05]H&SFM(+ *V(C.*&:;U@F_RD_O[VA)@:N6 1.&^80%'GU1WA!.3
P =P34-KMF0VE2M<#\A$N*>(ZF0[ K(51?QWZJX15UD5@5JB._GGT%;PG^=@N[_1<
PN>F*E1S8LSJ*@'O5A6AA!T;(.#XZ[T;FS'PD978.E[L!XO@&C NJ5ULOR7WN@Y G
P!<W%>S"=)[D\9\T @\JDVO-[,3<KH(GTZ/QN84%T7D#S]]O.XQ2UA^#79Y_+4!UP
P:),>*5V1.6A]A;>#^JJ;8K0H"#96G!STS3IO/T06=Z-J0W[EE"=+7,I6;!^0,@%F
P8E,<8;?7Y$V[2))-9U$P#V1=42R (LN4L4AE7%=R<+2K B*=Q"B8>QH@MIV<(F_U
P+U5E T(0=W7%RMU>B'+\.F,H#W%\2!C*F7#NZ/]!A-3>L+9@P_O_GM"*,?+B.<[]
PA5S0#<TWG>Q<?+W(\1GDP9V1#)ZWL$"HZ" 4?X-C42?DV5M=IR&DXP]$G M"<BC-
P)48Z[.%8FCO(#@ H?6VZ>"2<B7C !@R*Y=\(\[PIEQBBRR.@FF&4^ U97\(UF_S2
PFN@F<0):T%^C9WCTDF+;">_TE7X'C4,@11J$YN9$&)NC[CXH4CIA/:UO8 OCPA)N
PB_O;DUP>$_T?1\,F*"^HS\Z 1&"ISX1%AEFGT76@C^CCZS?U0NA*>(57<.Y+786J
P[F1T0\\*-9D^5S&:J,@#4P%'H8'X:6VO1SJ<C()2#=.4I=.$!XQ"<?C!ZE1PDP12
PYQSG#Z5)97N6A,_AJ(<:RR9RYQ"9S%IF5]7"NM8+Z[A(;XJ38)!2K[C:9H!\5P4+
PF2VD+V*N@KQP<IL)G\P3'#DT+!Z>Y<:<5\G$<B,W^!-4FBF-7I^2A[>;_*.1FG0Z
PR_O*1B3)$0*W1-^'_44$3KG5(U#+'2I[Z>_O3L^;I4+A&C?<+%^'(H<05!>^3O:H
P?]74F+)Q/,T/#MFMN!:HCU<T-,:F=:]YF>=7,5[=#:H*B0S@#46)P7CN#48!=8@B
P@R#"1HT@V2PFJ]N.=66(QH6F?X@S#L8[MURS#"L\G- :?;G;*&>.''\^P6PIZS8S
P8A'^<^IJ%*J_A.%?.NG Y!8?6R$<Y*Z&/=I TF/S;3'OKV@@FF_0&"8G_?=N/F*[
PNU8IA>L1Y,K3X2VLIYS7L'A59R!'HYMIOI<2T+B#$.A6R+K(<=NZMY6#X%%IOV,5
P?Z'!]D)C^:YM>VK<S$&]=JV0 GHTH/JY2Q6&[BN3VL++ G?; Z",,</M@I;$9TK]
PT8]SOXA./EP@1!>C!63=489!-_1UA/R=F"E7_\Y?:FB^#_!U#$?/W74'5:L;D>N$
P)P<+D3)JN[PC&]NV0I<1$&$IF ^<Y&TDRYV=6OWW6K@+W@8VF\R+X+DR.32G0CN/
PJUM[\9GEBPN@G96#$=&$<K<N#FH9'TX9L!!59J_:VM/\J9!LJ-@^[/"^_!"3PQHQ
PS.(^D*2SQ;._JC]TDWQ@?6LL;@T-'HJ8CO]>WU*8[Q$-ONM$/RIQ;X%:Z=;MB<LM
P)Q_NM:5;\OU! $#G\AQX7!+'JKQS2SR'<4Y![\:Y5,+9"_^F8I<.Z0UPD@]7\F^O
P2894Z;EK9WRH2;N#(9)Y?HF3.X"<1@T+X*=X^#=_$(O,'*W>C?8[WS?5G$J)2%:0
P7LB\OQ5*F83._1.C9OS2;LX?'D=>'6%BDU:RK\_<13-0W.@4JO1G(&8_ RR9(6YP
PLO- 5??ALAH!(2WLB& PENX\7/F00LFT_0"<*9W&&>'YK9%!$5G .:X@UW=LK1$/
PO,9Z@ 2*_8TB]JC')LJ&]O1&F:%,%]B!A7KJ[& /75-F-003GZA]R+VJ#D""E$@_
PE'[ ?$M&2ZY1VAR5*;O!&OAY9W+,NU9X2' &')4>S@:6O(L?I*Y .6M7N^Z8/H,3
PHDY=$W&#T7>[^]^:3$FRP^M1WF#Y?)P[#AVP)ZH#341C0]/BQ.NT[N:_\YP'@:>\
PT*>KL<HU"N62<.L"YQ! @?E'/I(HL!0_%L6(Y_:4:.CX"8!+K_]ZZ$%<&X?!O[G4
P#JO1]&@<0\!-$];#<IPN1%=I6= XHB+#M:J)<3HLI6 9SDND#UX>H"?.M[9YVD1[
P?D\:%PH%,CTH^Q'Y&:(1^VO5P-SW)AY#OZ:(I%FEO7)QYYGB0I^NF/;'C/ZAL_P;
P1"."U__!Y)TCOJU(G'ON4@NCPG2:/.:JCGL\1U9BJL##-U<[ZBCP&7_(5DM"AA&[
PJZ7ZZ9GMH221U#_094.H4SU[Q3DOWIJPN,&ULQ>Z90PYGK P[A</Y3PP%C0ANL#T
P<==X)NBX6_/I(]7^4>)@4^4 Y!R+M6JG^.@\]@D^^]^TNSY%] [QJ7@_;=X[*/1>
P(5I;^2,L$KTJFT$54POSZ/1=^'+,.2K&)A;,M*AS!;'KW=46Z'Y^V A]DCFHF:(P
PIW!A=HR23S[!U;'&>MIG&/:YX_.[BLGJ%A2)#WYVP5AB-1:N2WQ:W#:H/U:W/NCA
P#'N::CP<GZ+4G'Q[!YED\7,H7>U)=+0Q5U=BI1^TW#-[9NB*&?;W*K <Z$=)! N>
PHA-AFW>&[N"9- 3A;19)TI&!?EGRJ]@#'_[_7FB:IBJ_1/H!Q$R<)L"/K7;1/;J4
P1.*HT\QF-N0IRH9*X;:=&!:2ZL]:L!<V8 K[;K F'00E'!V[#4Y8D"@-%T,[LR*P
P;78&J6B"-0^2' TW 4A"7*]V[4(F&CD].<9&*/?J11H[;+"0P=7F1P<"V^A"XV!9
PCU+@[X\'7NZ2F]X4);XAE1"YBON0=\W0Q79B2/Y3^9;YCVAPDIBD'B1SPI_=!9(1
PP, F^_C5JG)4N\X5&G^:9^@ A;TMI-3W\_V";EB(8 ,-,&K9@A]5'T4.0>[6X@RX
P*ID#R^R&+1G^['(2TJZO.E/HH\51ZH,NPVYG[B.8#WYT)+3?6& /52  2#P*IM=>
P#_^!BO[A*RM(P@R\@;Z.R7X,FR6B5?3Y_)[="?W$)_].,,RX!>%@OLZ%#:)Z#H!Y
P, GY-D*M3=SP=_$7:1Q20,L O$8K*(0Y-..(#G+GANG+5BME>W]3J_#JZZ!9N&.$
P-*E4/[.JYPS.XU#O4KY$6!!@I%4]?M/#SUH;.69"N1=ST5]'K6234HH"5?EH%.8X
PQD @5EV :I&X6$FV:\' W !,4H,G%BUCETT$;HAR(^T;*^[\E(1QBPP60*Y?#GJL
P[0BG@?/U#V%#\*HTC_9O;R9H^RME*FN9XWO>P_MA;@_/CF#=5*)?_N0+GAT%*CT?
PM*HT]N](B2?AZ/=]/JP5>F")'UPXM+4BTK%G#4;X-,J-AL;& +0$!J#N<367^B=$
PD\E&':/367Q49?*@5LUEO[\17&T>[ZEXO9"%<_T%6S^LWT^'&#/,W.B#L*/@[T,2
P0'K2B)?Q^3-,32M.]NK"__?J(,H+&YF)Y\EZ8K&YJBV+S]?5K\AB6!97FS@D1CQG
PKM^=5VNZZ\J,KRLQ2?0\2XC3R FGHP/L=6<!M-LX8O&R.M-I@T6/33SDT\^C."4K
P_[DBBJ5=GJ4#WPXY5^[+QIV1^,0K*249'6EWD30TJ5%9HP>@W/,I N6F4XU_YP_!
P_8J5;2<TK=+W6BZ9V:W?CNC_)(2JTJ+(T!(E$6KT9;=SC%[!D@'L@_L(S$)^^=%B
P_MS\X%  >>&AW6;&[#A70H:A^5]--L]$ 868_^1<1,9Y(8]</,;V;;1C!H@P 2^W
P1+ERB96-^K#G#$MO#YW@;W^]20$\)KY5 JEZG,HAMM.A6^Z K)P@JC>* S=+6ERF
P^9GMS3'9@Y2=+IP2+@T"S$\(BX[#3'B%9]3]QF*^6C;52+>T;4.+B^4+XNR%$2E?
P GV?"&4W#TA''S5E(F!K;"L)&S<]*G:-&!5=;I9,C.^ &<GI:)X_V';O8&<X@W'8
PM@)0(Q$9UNF..9J"XLC/?/I?IQ3X?C8=LHH1!-?>+O11@"JP\_3;7,%O5':J2)LP
P*,*VP^?:-^GFC]=?RAN=BB"T)AF!]KG?UTVTO_$L0*YC[FH.0;MZA\!P!K0GHCU1
PYGG"L.!^+#_W*S*\D(6J?Q,-G17VY ?OZ,_P VY+J?S8L6HU,>&)LWO4U3"7!,(U
P)'=2/,IQITU&*NM!QLW$HE^>U,<]@ALI\Y2?&SHLD/Z%.OJ4P@8R:$7A_2-TMZ9\
PNH4B7K&8HXW:J$-WUXW?X/R_M17*;%.+<NOROAPJ'T3+P_NOU7&>((%B7%C]+&-=
P&F)<.U,I<^*4 G=_^>W<FTF<7K2N11 >0-Y;QQ'JXM/&MOGE .S.$FZ8E -,%M6J
P$9)-V#</H-X(D*_/8C Z8@.$_RYQY/_G@G_=)*'@B1R] !?F$OJYM3^7A@+0O$61
PKQ7QR:).('XV=>X!/YTQL>_HCYM2R5,A"T(ATY6LT<'($W/JS:>>Q?&C<R=O[;:>
PMH!TK/MD_I!#S46[;$/GQ)?Q7+US!LW5$@'CU_:[%'LVVYR@FW)@:ZU?;JV<WL_*
P")R"[#.\ !7W_^1ILTL1@<Z @Z6)NFT;:5Y0[G0U>F]N\ U^L5@:(&>[#W0@M==[
PF6EHW[<_(-4_6_XO >:KE6*X"XV7[T6[#K"G59.&S3WIG%0$W?]5A4T=M9]:T 2Q
PL;WDD\@KL>F\I=\1B9%:8&5%WBNGZ9IK\AVP(85\T/Y%\;N%.W*%-QG&6<,-NWN)
PLQ4N01*/_L[L>,6H4-V8Q6S"!D1YPU*^UO !!'TDT]\H?I C:4#"J@\OCN:GA[B9
P[GS'7JK&S:-%P,&1ZK#$3<?1P(<&1SBWPW.(C_=9>\@%^0?>!_JPVGS)'@@KX)#'
PD']E/5AF:8=7R,X>-BRUQH(FMP7N+"J;8Q7B2,E67 OEF$>!OH;Y?7MDG/%4%$DX
P=JSP7^DAG  >V9&0.(#[+F]C]FRO3[I.3@'.9_F:9%XO0>;K_E:[IZ2- .)T;9$:
PNV Y2$!B/I&.& N"67N1H0JW<X-"1_-E=<IBT/U2$PZ+'3JJ-#KKG=J+R6"D OD6
P"[RMEI3X5373!NCGN5&L'?]L$Z)$@X21=EI.Y-D^0U,:$!^**#7XI=M]\?@?TJ>S
P[583J2$^?B=[:6_(KWP;9> =^I,ZTQCU*DO>Z(7>/W-'=$9K^6:R^>:F5FI:O5$7
PF?6N:01]=2D!'BN+D-(?LC[D1#3 6:W*YVM4;+.D*O;UUQMS!V$ K0!'?]8P/?6D
PM_L5$)Q6%!&,=Y,%/G^YHEU,-<8HP;P*0(I'ZZ*"U)6.%(F6^X=N4),]X'TDB)=Q
P:%GY, [ZNTS7S+$[3(O5%^=+==9P9(,YF4@;$6G&UL"7U'2B$]II2Q7;(8IYL586
P;O)N%S9+WUL5\-6C3_=]/@D&)?))>A;B:#L%"L.WSHQFUA\/8C8K_%Z[023ZVTIU
PM\QI/.YNM%RI^*S;QU6Y4W^;U*/H[!U0$I'?Z82!7M.VM=@?SPH&6*C<O>_K3/&S
PT,1P6D@U[5!( "PWYQ8$4$A+/NN.PB+^)P'<:X D/;1(T5,?F2I0#"T>H. N&!J;
PT2>(?7_'$OPZ_I/XCP)$_ITQ&O_/H'3L'@C(485_K059,^/0WSVC_HJUI0S$!K'P
PSD2M[75F0AU50>C=+S6YQ.QR%O"\^W/?PE12:1;#28)QC*LZ[A-)6\F@[25)\.# 
P [W5?6AQJ?30;U'*<<V51[2R*5 6]L7YM"0_S//,4]M@)45.WZQN0I]Z4<(*F@[K
PG>PL5D_^V;HRI]>SQOC_9\\I#T$4!/CF:<)%A'R1FI21,T_DI>8&1,+)LXXKL5Y;
P'&;<M3O0;)\7>N1*5RACE>_1(%MA5U','$A\+Z/S"?7M+OV((P:'#3A9YC'!CXQ7
P'S32[@W),=I :H-&_*.'XJ+HQPV9"3SJJQS&)B?3K[ ]J*831\='SL_)I1I?Z:B4
P-=/\=HX#8H:<!YZ*(0V 8F37#MB1Q!/57L$G"%@!TZAL*A8U;OZ6W9RB]!/&FSD'
P9\FE^9,Q-DRR?-]N>Z*>JGQ:'N@^N3@!<_M03_M=VV1R(F*%_^2C#832X7T7-M2P
PP0>>A H9^Q7'*J0&JRF)^9Y.HECACQ='6W*?><#U!&4DP%O,."RFQ=%XCK6F6ZKU
PWN+^FOT1:5-H(J/.GD?WNL22LUV6H3P-L!:"DB^*2%IXNMP3SB7 5%]"N?/V98[E
PR\_=&TOGS>L]E@PD88X4-9?OU)+"F>8],EC)DDXR3\$1P68_WX9=_$\/SE1\J[IN
PYNF7R/ERNS&*.?C@:9M$8Z[[.=4@3LXZ'$EP^/IN60 W/X^>U"6YR5096JI<%#]V
PZF%'SEQ_I@6H@BKJ7!&IJ;C<\EU/U7/7K02,H 2.O] K$YOPC7^ 5>\Y$(%A.ZWH
P_$2EK<8"\L8OE%Y?F"\!DROV3)_QN9!@>M&OA@HP9PXU8&\[>B[:)YPN!4PN2@"A
P9+_G=L9V_.XJR=:AM1JG%XLILLA;=W==S"FMJ$,ZFK0G8!(CEI5R?6E7BZ/4[ ??
P/*D9Q <AN0!.(>-G9+S"_[W2*7C5K8QYNY E-_M9M%H)/SZI*QBV7=L&#,E#69F5
P]NYPF@YT^ %T*!9]N7Z4MN)\:R9*54>EO]3L#<4OO2PVPP!6YH2PR3R:O4:_U%E%
P,L%MTR<4'! ]P<(C5QB=!;LV>A42+N=?A937[*?Z%V6.H[\5-ZIYBP.G9GI<OB\-
P"N7_R\=54S'F+>4'OCWJ6G6 _0=<=EN',G$P'7I95VPI.4:']_.=\]"@FZ"I[+3.
PE0#K$(@1P")GV > [-!I3&0;P#0C*VI@L)WVK\F?@2@<\F:A*]O _/-V(O0Q^P7I
PAZ9=#1W\JP!=R%Y)NJ:=9!/73Y8V71?$<*I#ZG">N>>O[$BY/?0DKWX$=,:.%SK 
P\">6@?)J#J$8XRI.=DG]&,TBQO!Y7$-@P_ZG_Q /$&>:_S*1'ON%5(:B6"V+IF_C
P!GBXT\QC.#= M&G2L!HGC1ULM<2/T ?2](C1ZB]>QFY4N=-R92GC*4W]]?L 5=(/
PKE.*MDB"%W*J]&@CE\MK2/K-R#A'/NC1(4&<?M2(O5A+ZOK)GZW 50)1_1A4<88D
P7V#A1G27\DQ5EOTX5,.WAU6>,/.!S K/J6[JC4WP46) <@])_ /-Z;EV^2>DW<X]
P?WUW2\OY?B87>/H??0PE!@OK?7O@"V:U$M2XD XV1DL$2%I@%M^6*6P1#:'TAK#0
PZIO,FNL^0;-@\M6B8^;F&>1EL^LND@'2]8#IN7Y[UM1M*PJA&>XPPYY$D;_,8H (
P?,OE=[]H7U#+YF#MZEH/JWWEO-L./EEX<O"0;])KLO$DD>-0>@NA8 '15B3+4%J9
P+7(47G&'PTY9T>=U5#KLM#'+>?SK]U-I\O0!'+PP]C337!20?X/N9->>IR %N1$M
PSCRN:?YML?-RWA49DCWOX.6EV)+>4-N\G99$;IE3BYH]W 5P#$X5^L]K\NLDZ(7_
P%H6W,X-">I.VP:EW[J:ILR*3:<C%7&3*+CGCR/(P*U 00D86$B:WS 0PH0CZ65LZ
P "GC1KJK%(0W,(TPEF@+T4HN)O1"+J3.C^>+CO571A0F:-:VJ^8%EVWXM1,#LN'?
P23D+VI(MCT@6?W6B"XA)'G1^GOG'@(D]HW-)P%!!97EE&5T9)S-8M!][S/&SYO*;
P"@]2KH09K;;ZDO%>[^FYO"W^799S,>:%E</'&12J3=9[+OSYDK3_<>>VS<6^?.IR
P0'QX-FG2V-DOI5L=LT"C/N0%820R0RP5LB&8,WU^6Q8J=C:7M*'$N)W''>@-O!P&
P/[^88D7%5P!A1=(7$=C_>C@RQ 0IU7&@[BQ%W(@FNP_ D,]6'C@%5F(KN%HHU8B*
P08>2\2R$$ V&^_.Y^7^ ZQ9Y+T1(F3 M)"57_3Z>Q#6?,1\:,A_ @_9'TGLH6C &
P=:Y5",GU>EA8$_YU+'M:TL<\!A1F*H64L)A\GWBJ>O,6W'&BA;["%$/$8*R67]]:
P=P/;](X-2E9@@+?D;ZI.8DS5B^,__;(E\122E3<O^O4;KRI=1B&S+HCQ]]9![->_
P=/O"L.YR]M!3A7P!=BBN.(V*E <BIIP^_JS<</;_2.K6[XC'"I7$E'$%1X$@YS6'
P/GBA0CA#K61WYW(W4'@0L3H5,^P-29^-A$!3%W,M47P[Q&-_G='G? 2M=CD?,H@B
P=,?7#1Q[%81@EMT'+HRMPGGMI89LJW7=AXY#;^>CCKPU8B<#%)_X3XH)-V>V6YBY
P[B7(_K^8_3O 8Z=^/LD%_ FKDE_*H75ZUENA'PEC%@W7+]1T[&2!5.8JU8F>P7'3
P+UEOP^W.I-B9.);I9;,!Q\9@,C\GQ"IW9QW=D;-FS\#C85QPOIC\6NENH.ZLE]31
P.&OINS=#CGFZ++% 6IS5+;R A-@-X!T3G.V0)8-W(YJ*P+AB"8@I0X0?!2X6E,Y5
P/GH!KE,!U%7^E]XZ1E+;]ZEX>Z7+B^J_-.2H=FS+E%6VQS91*9(=S/&?G#0SG]H]
PGV[$<HL ^]^$>H'SO+;L\F164*>9-PBH&8][LQ,?P33;DWKF/W4-<3HQ^[C!N^X_
PRRMI]E)N#EK2/Q@-$D;7@?WR4[:!0$Z,92\"J,D%:Z$(UP/8:I) RX!Y\<(0M9GL
P[3_P#LT9\-!$%S =VEDLC<=/A]IYB0X:C#SRO%VD=7G*G4M(A/=W 4\@JE[<];_*
PZ(^H8R>M<0:063LOG'DJN6#M(&3?#!(B^>E3%LT(2MU&&5RH=',$ /C->GC36--V
PY5L'ZHSVZ[JN@B5\7[\)'QID*Z8B*G<A$W$D?"T)![YJ2J-TA3K(W#F\^T[G:DP3
PB9A3<6?KZ_Y/0'0\P!-5GA83LVQ NB;!$&I/58C\=R"#]:I';Z1H)UTVS[!D<X&K
PWAAV+CKN(4_JLBVW#$]?A6:>-7CVM]8-JNZ7CNEB\E0]MZV:FT&#N%\(1\G[$C-+
P<P0D.@B8R&3FNAL1!\[R79;OWN_,O<7D]D'[1ZA6S=_'1=2T"H<Z9@V#9)OM3&2?
P*F8LQB]B6/CH(-X)$##?3RL^^D<Z[(J/$Z^56(2Y1<#:T<QX7W2%XCR[X\RM]!OO
PZF%\&9EQ.!MOV$@UV;.,H#\^1#W88?D/(3_QQJ&PT,\!H08(7ZSND(*8N*(MKB^?
PI0!UQA75767HUNJL8XSV+7$A\CVHB6]20"SX@ED)>^9A=_?V80C$S)&+>=+?4V?F
P4B?Y264K"9(T6>5IHCJ7ZL<=-4XND81"U7/= ZL@F0MI[AC:6T8(9'7)$D-6C,SV
PGOOJ-CV"! 70C0Q G&K?/9;E?EI2NJ JG'(R'! H6F-:L)7A.KU<%F+KFRU@0B'7
PZ%^. X-M +/]@W\'C'4N7N#!1DZG6XP9IA2^$QJ?QK_U6=3X0QUX-FP-E'DW')TR
P(!A"^#\%)$G14S:6SXK,Z9ON.1)/.VVR 6C[V\401=#P!0P6C('CP3)$S*QN!P6O
P5.7Q"WA3D!69WYH1DD [QTE).7+67ZLO#2B_)[R7'X,B1@(E/-6TINH#TYL_LK6Y
P6\1G_ESE"A+:;,CDYXXX'X9*/T#<-]HQ@%X&'VX,XS<6E\YK5.NBL.3GP(04 GX]
PQ>B8,HM3Z QT7WAUX8Q6L2?Z.J;_21*30GJZ^<B%NAA4^V1_LK_87*+8N)ZW.$58
PI8)Z<5(B.&GO^ F['(B,V(KN3V?%HU)"UQ*Q<'&4V+57$&)\!56/D5M-3-IM))RZ
P-D=D"9@UME&69R*F^(-(8!:OJ;S8$X0397^A[J8Y\7]>16O^='Y?';Z/V1>@W2AQ
P#!)-8%KMED8I /-O)ZF(X?6R\HHIXJ%D]?\$F JB? RSO2N@%>BW#%,>;-INEL3C
P%U=>-ZP1[XLH)J6[](S)K0ZQM?;)-\5S.J#75V)^:9T7MW=D;V _XJZ]4ZR8K7>\
P-#@_%)P;9)?*)&!.)8>2XV#83FLKW6U9QR^6L"9_+U<G)?Z\'[K3D %.C0RNZ1GI
P%%&7W;)>OL^$O%IM$9$X.L-0?<\C(>J7?7)WXW]#(6A.M]/"_VLQ,MG++W<YB&56
PXKC12<O[D3.>&KX*4CF6[QTE5O 5Y%V\5M[:_GTV4$4OOURZS0?9+;^<XA= >PHO
P5A9H"=P1U';]_5C%5]=)0BXI#] U>0+U$E!/AAG/NEE"HXP]Q6A/HUB;*TJL+W;9
P;X2AIEK>:*T+)#:34D4;Y'K\9( ]QH0U,+-(V8H-ENCXZ:WHOP[U) O6K5R&TW<M
P&/Y(RH?Z\LE*@^3BN+1M?<M[\\:P3 \:4)TPI5E[P(P.F$JD6R*?XNF]._D+2=>$
P(8USJ<_?0OS0_=#18BQM\UCSCZAN(8!T$._3U"+@UU'Z/U>]5R# ::P::[1IEAB6
P$_8V C2Y0^S!W8'&U%F*11[E05CM4E*:*&^WI^L+5W=PW2N/BKC)CF5!"IHM>;ZZ
PNFIRP3A''3HGOE"K%,*F/N*@1@"3NWMP*S=W>:0^0HS.BQQ/MNQ02^Y&-N<UDDSB
PL>Z'37D=8@O&O&U2HHZ>&S)'T__%;SSEPK)( U'5 0;&E01.DF#G!<FUPA/.!K<X
PT5NR6QX/J6@N"I0G?LE2W[2(:5T_ @M2&7MA+NN10TO;EC+>/\/&G";AK(92?8H<
PXPXR6&ZA^ Q*VBVV BD>'++*SG)K@ZNY^ B[J_)]JFY^"CFX(YC)DY.[;_UP_(Q\
PD 98%O51PO7G_JDSO$62S9O(K?][MA5S#(UU0U,#5Y\B".:90MUSK4G5 >Z5CI9Z
P40>:M9?@O_HF'I["5TL/^B7^>7].,TZ5GU4PR*N/^GS6T^V*LZ +J<;B=62&+C7$
P-=*"X^?C2!;<8Y)F[J8L[&'&Z]3"J--Z?S>0# ZI2/] PU3(NMW_?DD91[5&%C<%
PWY'WBG6SW82]_$RZTV:)VVA>6C3PRJC_S #CS9?%H!K=WJ4Q ;Q$CK[@]^S\*!]=
P,/@.I]491#;%+&:4BUQ,T19=GWYCRM(Z(/5RI"3?M9+)&AL)I(4-I[^Z/XN:LGKW
P#2.>56#'\W#;1H[H#VFH=([S,8 TD;SK97\Y;N;ESSR O6%S&F/7=/@'B?RM:R$>
PS=C9^R 'Y*3TV$&YM#;ENZ*:LHOW:0\@"KU3!Q17X&5/I=H&ET_+$]V]%ZM]BERS
P^N?V_W@.EY[;]\F[I"9T)MGD5'02$*G>H?MY,*0S# "Y!+!^;%JM*V,\JB!'4&UB
PF[9XB&O>K!X4)7^Y=D17[$I@R-4,L ,!^\"2'#QF/LV.GA7WS\:(B4A!Z=)9;+HR
P7IW;V)/60C 8*=GJ^T3Q[,;:WTZ2[/23K2Q0EBA8"BP*ZNZ/@!'=97]+%&&FKMK2
P(G)-V@&9M@F$M4Y9<[Q#;7+_JYL$]AL7E?>:27-_^6K%CJA1N;]  4$#!:BV-G/Y
P$8FLJ>47"EP': [F9<DQ=!#LB_XB,0Q0AC.//]8V,8_CU4O]*E4 N3#4WN%/]EU\
PW'5K9U@KU1D!091)7)].(J)'H4;//R._3XY$$EQXIQAD@_AXB824ESY9MC.8(R ^
P[[5 ]P%0'6TZX@M>(+?I>G.??->^@6FH9$:5L0'$;&*PALJ'+\#E6';@E:DHS)@%
P1_#CUX],[DE2*4(H%DC\,(LFG_)$:7"0C%F,"7W%%V!<)Z@9"_RI)F-6ST6.,NB:
PM:8":A_/(1?*#$^%(\=OD,;^PZ<QPT\IC=$KVC_;Y%[KMFM=W>Z+M\.Q+WGP1)7N
P">/?ZP\(WX2[5@"XUL>913 @.6,]EDS5=I>T/+AX5V-/9]9+('M,+:=ZL]C8ZC[/
PQT&&R5T?DL_EC E3,JB\4:I,<"842UT?I((B\0>IE ;F93Y<6@,/DX45G>+8HD!V
P=!08?8P)@S=)N!^*Y.3,JNR-798 "&!$Y-X:6.-%U@P..1.)?ZE&*F>OIH#"WQ@ 
PB]QM>ST$_I4V'3 CSOQ$33!"Z#/V"QEG+_*3L*5V,M*I+YPJ!*CL,K$F)<FTQ$$N
PBD.B6=?<?,.J1J7=C (9<A9@$=&XTEBF^ZF1(BC8K_%UYF!H-31N-&WG7OE.BHM_
P=LNK B57>M?IEPX"1-[67KSP 19^P-L#)2KB?R>EWX#"MR09/CRE!68 $5)&Q@5>
P9'4L")3VHZVA.K>_4VG?A&2U&>:D[;A7:N%R:@VCIQDE^'O=],:29+PL!8?X6\&,
P:,7$@)76QFX8"Y_):2*270<X4*5@!=_06S2AQZ!+\9<M#%6^*M/TGJA6^-+H,#5@
P6AO8LABWF<W/OB*K]']PM24N$# B,%KFWK^#BF<,R^^&>YX<D^.\Q>!L>9"JUXZ,
P,[CR6W$<F@9F[]!'>$X-P7E(3\J) *O]C/KVJ(2[IV9/6NTB)]PEN5^-("P\H0ZU
P[GV/#+Y7!MB].5^/'A'H29\?76G>PR[NQ:.;?"P;17R0HCQK!KN4X9T:;Z#\L^EC
P%TS *BIIZ0;<M6<A&6YK*!'$P^Q)KQ^V&+,R!9D%L\5,\;(3>F2'>!52\76D "&1
P(\J>).B:@59,M07/DE^%.PB;P)X)@;<H$OU7GIQ%*OL@!,6-7H!N\B:.G4Z4=_Q7
PL4<5]*_P_C)_K&B#K;@3'! ?M[<H_"*( !I$ C)"6;YNCUI_YI2>\C)R_/;,OMN!
P)"Z:_?6D9V@S>!I<8M4K[E198\/YFQ.=*#8?CT5&5$(5-MF7[@R@GF<G-<;H>4-]
PDW=$U.&=JF?_/$=T$D$MK5GCCZWO(%^NQ8])CF;J?/X->P.)C-?!D;'I3+OKO5LN
P1G74=3H0[&<?@/:.MS@D47&,#> @%.^QP*R9^)02=$M&I>8@(LQ[GT;'X$(ABVCM
PWQ6:[AAB1WZT\'6XU0 R_XV_<SHM@Y0<$B*]Y8(-H7_+!GR16:6N(%S^8U_C.SFG
P/*0HV#(?5#."=RW!CR'7]90O#N<Z"&F1QLI.T."R+(MI8*8Q>]&>G=+-^A+T(1O:
PVE)?;-$(R+5]T;LAO?C'KDG+.);2?/PK,+BVL4T7)%.,NH1QQHP-MAJR/@WG2+&R
P8UY[&=Z&8R9,]:MI?0+I:1Y+:B^K$IJQ"&/71]/DYZO_>L3?(D' M8#=8*Q8T63R
P%.[91.0*VQ9_PHAZ4Q<0H\SY*3@YUM,=8(DG<82$GX#SPZB\< XWJC.7\8SGDJ"1
P@=I-*L*@8LR%)$CP8_4XG'"#B33@1MPGB'I8#SP-NO]!7/X?RJ2F\(%D6*F-7A\0
P\2*QU[V4&/D:,3P T"%&OG]C#WALS8SPGRS%L;-.3_+=5/-ZHI'N;%>_P62LFS[M
PRCZ6JE^=[^Z&WS;O-&I#U_*!-/(J*!7_:!3U_ENNV+BC'? 4R=NEX B$H<>SI[E>
PD%R.YNJ[PN$Y;QQ IQ"UNR,IQ!&VDTV0$KXE+%N?S!)3MC:82MW,M[6OSK>_KJ6B
PEZ"GWF"2VO!0[I4A*V4.55^7UPF#,DU=+^YA-TO5MV1QP&8V_8L-5@<[ LC3]0<7
P0I03TU&[6PP1=NGR)19BK\Y$ M*(9X?VY,]YK?H+P[BNK?&.\3<I1?BT-N^L&B0;
PZIR QHY!AV=9)TC;K]QYTHWU2B=,7J#\Y5P_%Q:Y7)21W*WFF2,W)^0Q4]OZ7BP,
P#\W8XG)JS]$97;IXXT46_-J!%E*GFT%3-5OTY^/:AMK,QQ%_M8XXRTOA,?P]G#&1
PT*H,*?@R>:(A,BW2)4U/P)'6II<,5DQAYW;?A@.="X!1$<RX79OVXX\?WD6;D[G>
P5H*3OEMAQ\'X"8[NJ_A?P*?BCF]/^-R%C':TRWEY7N>O"SY$X;8<>X?M.@2D80."
PPI(&LXA?#*T?_W<Q %'\2IGX65S1@=E-=5#3^LE\%)_Y=/*/,^4:^ E>;3,3D,8W
P>YAA9%T.D?^1PTCVVX'K$"9$<[C.Z'^]*?!".5V;9^&0PX@E-WURWVIU8QDP<'N<
PS(Y_D=1^T<=B3"T,OL50MLWEHDJ5%EA.(^R]> NF1)G@Z6V*6F,^"*W+.K6'+DP+
PZ@D'=:/ \J-'WWL:M"U?4YUL;3T7.3PXU&T3;* =-R];JFD>MOU+=W.&VD;$#5L%
P&J!HS>>2[J=V1QU)OS=BZ9?9ET2X/4JN,KOP-(0X<YZL_^45J_,IL$BF?MDGS&;F
PQN]7+*W+RA.%V1X&!L5N$+Q)DCP(Z6+<)Y5%^Z]T+U0DA"H\V5K")DMCHY!7VN3?
PJ?)EQEMH.A!$I?1L[YWN]AR?J@\B=08!-E9J)#D=\"X*00NC"&A#T0((5>J0E!X]
P.G.1A1FBQ!8YO0K9EVPBILFNF6-7SS=^2O 4NC2=_URQ^<[^\QI(6+#L D.8Y/&/
P"FIRWX$VZFK["74QLI53EL%"-TF?P;M9@->!F'0@*=:!+]WHA8KL>'[Q0R$6MS$<
PR[1!6G"3D3-T)1QHG<7"FR1>4_8@\)(;\--* -6@N22N'S;_$[T !_BNF;'BY/(Y
P[GU12==$Y/VRJH1F?C]56]*Z$&GEUU8(#T@(MJ<V0EZJKI%KQBZ+')K3O0H]"NC%
P4I!9(CK-6"&DW;"@\J@%/-J??$7EZ9W02P>/?!=#A-#) [C8.J>P-?D_20T,89^X
PY.Q;LG?43!/# \@OZ6Z0ASTU?/RVHS8 :%]L9A@;P/I]^K_E7>'ZO*&*(,#0,(\F
PP>+6##T7S.W5LA9;55&3^F8'TU7.I#",Q5'@RN7PN:QE]J'U'J!K3W!\"?J?,2GJ
P2H(I!F.:+!'*[S7E'' ZW?H"/7^FLO?C3134P?^9E74A:(1V+)^H \U)B*,[5SA+
P!P4_?"8J'<;YP#TF#]:9N'WY$E]R(J&BOR8AP(?,E,J37HZ5>=DD6\^,,'R1_^>#
PK!Q\\K$.,?8)_$IRE>8@B7J5./L^G_O7>FY0-,P/YU/I_B+WJ>(V@RTOE#K+W&.J
P/OB644U6HK^P40(M&QDK57?I4;BYC32,LZ$I'3!/[JDJK4@L]4.&<>R'HNE_6_I9
PU@Y*6Y%VUL&W[G3$BIT?T*\ZU9XUK42-?[D$[/_MM?!1>L\<5@^=T* YX/*CF$P;
PK)5=V+2G5W_+W$35 TMWU_D"3+4_-#L31D1)N@[A6)#O CE63H)S&>X \6ZNF9S#
PD-:OH^G<&[6<(!MCSTX]%'-%P2J>L8DJ)$/.(DV/6*?%,YM$E+9DW<3$F]-=\+?L
P9X9J=*Y<0,]@2^"HDS G4N@"'X5*.%S;P7Z0,@^I1DSMI)A6.N_'!^T,M4381YWH
PP:](>K@*"K>0#(>X#FI)]OCQ\WVT%W[K&+\7[*"QN/Q#(7F]C8>-2JT5W$1RNZ:F
P]"[]TX6S>OAM4N@T6DD23RUTJ+\BF/8D"YU%O-9DT4E66C@H <B8"+-6]8\C(1/$
P"-?#2%-,X?)\Q6\((XO6*Z17\0$Q<B'@--^_L:1=EY_DG,4>ZS!0KH64C*V,R@ Y
P=$*YH"6<@*3F9R:9GL8+-=K\<H_#)_$LF4BO]"5:''CZFNN6% < 0G=_[JSN@<@#
P;5)=A#$"6]?FB<0N=O5S>L@E&RH%.XADH>,S#;J5OB <J(H.&\;J4*L7=(SDMV@@
PWR7[-!'O>QJ26NOW5Y_B9N]:6A[W=?'HSW\59!1FE'FFTGG1&I)7_@V4,?FCN[H>
P0KC)TV#XY0NB,71:XQ_*[B[*3NL*$OBX-U0C9U1+UVW\BU;BLP0BD\H)A 0@.[[G
P71?BCB,K%K16N-35U]XD88J,AC)P:C/7*I*G,8R@E#^6'_Q_!>_P*L4"M0D'0?RL
PM.U'S@![XR09IJRLABB7MA)[/67$Z='N%OTG5FCY8($-6,.5<GN!XLKRA'%R<8QN
P0@LM1H4K@%C==M+"%[/SW)R\>!>J[?.T;)Y8&6Y2SN?T6E";H<EGL[=!S_?RL:5T
P@>*VGM6J_@+B*/FB2]7Z*MB#D;ZR/(*7;1#<>A5I_A0<_V+8\G>O'YZI7Q,[%N_^
P/=I)9$2V]01@!5N(IJFM4DISK[3Y2/4$ZO&\C<$3HHHH0=0BE39O[F>PA-'L$\NT
PS?H8@U4#YVA_4JG)2 2JN7F-'01\T.(FWI=E%Q%J-K91.!".Z=KR_P[_[PO"+/<)
PTY4E%E=MUD!_>U4J$VK3#8KK:RH?AA;ZH$_A&^$VFWNU+60.A&TOH"KX P+)><4-
P+-P0W2_')V%S(>;H&FC0(:OF 9^YEOM9XD96/ ]M=Y(/L5"T(46Y(5(0P5PQ6[OQ
P'$*6Q-.*H0HR4.,_=^Y23KPQ&P-67Z\"EB3WAGXR*6K)T'@R[\X<)S]NI\VP6\^A
P!O?A*,S;+F*>4]]GE+ZXPY(4@,#,]^M:XT$IJR<'*BKI)'MI1/'QDT;QQ@R#%XBO
P@1\U1SZW;8[O1"[W>E$\G1H>XJ@AGL=_XAIN^70K%&?V(G>Q%L&'DN:=6=_BC44H
P@;-***FG<"8Q#M8_!Z.@6BQWTLZ@Y+J/4Y],>):NJ3BYI)^>'],3@2T*_5G*'I]"
P]%5.&O\);^F4)II CY5S5U?6C3P\8O'7.EHWTZA-^8):VY%XG):UU# :'42M%4>/
P]KD=-49$F$2_:HDVV^H"4\8KG^OL"B13@'(3&I4R!0WBUH7CA/Z,5EY'D2E,N'+K
P.C0-_-4#\K3R1]VSJC[!Q0& E9&]"C%BC!Y5QQ16R1/0@!?&Q&Y=NV[6<$W[L5'T
P*%/IV*6UVQFR@SUO2PF<+#KD&,7JSQ4MV0Y@+E?-3(<-KW+SLOFT)&+"PN5@':?\
PR*J0.T0G,%U4DQBWCUY^)*[*47^;-B8\.%YXC]5%+?0V=]&2?I?;1(>3L-/X9.2Q
PH>NK# (;DMN?4/8-#CT7-'F")LFATD$Q(?6$)$ ?8'AQ;\"9&.\M\A[>X4Z(!NG:
P['Z>BCGM!^7W--VH@I68JC CR;M6!RX0'PJGL'W3(%TC!QG,([MB)E''P,X*L!F&
P2NOWY'Q0?9 "!"3HTNG3/40-)0]-/BYT\$+&_=K@.']_0K3$N;U^O[!54H^&1V53
P?KJ'?SS:X.458G@Q9K\\*VUU%T6+A#ZT)8Q=GM(XDZMUL.:6S6#Y"@WM$4\B)LB5
PRP(>IF)@T(5_/*V@)[7["I"U?7!9Y$83P19Q<T-J/IA"2P:/E20=GLFK,&QG/3O^
P2_%Y56/B.AXH\UELT!FJY+/22L3L*BQ[;VL)"Q,!.*M@[%'J;;]IQX5!0O,0W_;'
P'VHT.I-7&JW6Q$3H58:^4AO%V+&^1Q>LU3$[83YBV[9Y4Q'J5%&[]7V#(!SA^&F;
P-OZ!GJ"=+0%D',K5W&2?RKH*<D"GY<9S3.]A=8H!(TU@:>'=K>9L5%TRH/+NMYWQ
P(9?P?*]PK+PK'<)O101IV'B ^-8'MTLT[R\ID8V"YN4(7W,*@K;C_!<(>WK5##,U
P0>8REAB3WGBQ4#,%2UMB_*@*.&$35S<R@)"&4AV"ML&RPS ;[>;6/E#-!BZXOR I
P9#]TORQ=5=:%/Y)X^BLK<,! 'V;B#/:@S?9L+'AK#PO?)0QH!=%_<H^I.2U%&IA=
P/3PG?)O;X\W<1,VLW5 O.FM@*&24#5%DFO!;QP0O*API!]7=B2L0,OBGA/-1@A@"
P@OJ8N$#T)V1SER YV:;LL,)O+T)$Q). ZHEML-5'I9&:7HNLQ-EA]^UM/WM7>XKG
P3(TJ .G]U[.%FSVK@GE'=WRXOE7[RS)^F$7&%0[O)&7QR*4JR!>+F$1N8(?/##_\
P>#$CD^?\=;S=2]CV1'_YJBI!0SIV4\)AVW</7^, Y35<6V4/ ;[\U]V30@XAXAD"
P!\EF7HX0T6U1!&[Z@2[)M5E&HWBV:$R@EB'8ZQ*)-.4PP9*8&^5I$M-C=?1 ;K?!
P,XU590,@R3,8;\%_5<QKW&W;R32.6#[X4E596=,%6$@%U G6+F,[*S<GLFM)Q!2:
P-ON&"^JTL!A)<,(_C&-_E?<LEC2,W*]M+EF536UO36L\PZC<?&0!9H#\3[O1A3C>
P]T9(V^T3H.E]*@)WWX[<4)M?@*5&Z%1O*3LN6-I@)1D%.8*LC]*CX(?2/'8PN 2<
PRF-B([P&"#;%EZD=Y@\]WPP]#IK3NX.2@K]5:3(L$.@VNSUM9/_( 5YYGECN]I78
P2W):S]TOQ1;QN?39T.7N-=!ER8L5:;?'*-II2&.VWH X=J^(X_)*!>CO@?5\Q-3 
P&[3%AA7SX1TJSTE('1"%8H'A" (%F0'7G3D!V_ D120W7V5MT&+SS@->H5] ;KI\
P#>L/1:S;+IH&<TIB,&)N=TLBHBS:CHL0U]O-%#Y!7]7;A B)4'IWJL*VS+YQ8=:&
PS^!G!@*XL32"#.7,F&#L,3W,V>BP:5J:)ND+RB#90=<5WQZO,L(P*<H-Z2[ $5J@
P,,BQR%>4\T=+'C#[$:J)[;;R*T2B9^@2<,U-1@K+JP"/57D#^O)J.]I()NFT;)A#
P&[SP#:G:KLFAA&Y=M9;"6L*861"\H';GW-!R+P#_AU8$R5U_O"&^*+ 3VNX:C+ )
PH/X80*FAFYC<7?"NR5)K$XNE!PM<5FY24 \N$!H,7T"/P1#5/-9A$.S_2!W]QUFI
P<J.5 AFB#7$8KJM[4#A%:4#LV\1N*FZ7O0^X]17G,_RKL],L%;NR0/)'X"9;6=*I
PIF7!>N8J7"& JR-$81P=9[SB6_4U["F2%F#49@911T_>F/^=D!-OT./-X5BYXLUG
P&-!R>$S,B-WU7)-E!;I M\LWZ5Y<Z<V#+H7Y1Z(R''N9/\-<,N]\>4M<*F<9%;B^
P1"XB$D[ Z(5R\P(P./$V#2:Z[P$F$:, (JUL9(I G5%C<,L06[<!)DY&MGT=,6,@
P[$BG5)*F23\&LW[ 7W^\5[%YBKT2WBQLA>M()HGJ,U>"<9,86LO53@A2R$^%@<<Z
PHF8UJ$$2)5*>70MF3&7>VNRH^F?9#_.BWK%Y%TJ<-?'VT]=0Z/#%%$'Y:@*-D-84
PJD<Q7J1YU_]30WQ(JI=(0$\Y6W8=@/VO+,4.H3 0!K%O_U7\JC89@),;)IZ2''0C
PV@ OI'&0:<7BHVN D<)S-U'3]I[=>0--SGST%##F%T)P8,EU*X;M#-:PMF=YMMC\
P?P!46D1L_"/[YIXOS*3OXCR3#41MK_)YZ]@5Q:B'A2-:]%^=D&"*NDL\C.2Y/*<"
P6.N6'APCXI@U1OX_+ <DM$CK%?Y+7+3B;:%J2;4T+-5+T 0EH>^2,6L$Z(MO\@_^
P2B-!J<V="\X %2)]4DYHIH^PH+6A%O7,8$<MD*TPKW$_@LGTAQ*7YB\";=6V_+E]
PL@-N+W @*Z=^AN #G6_SW0<W8)<\&%NB);X]Z@EZV*OY?'DO"\-Q4Z1.[TN71<QP
PW7>2[K4,J^($[M,-!8&FPHI9_:9*(U;+6LTMLP,O"FH >!710ADP"%P_5IK3Q[QU
P;B"9N8\IMK7<45D5_BIDL_O='94.%]JJ.4%N\Q[4]N[%O&I^;(7$7;5X&%?42>E<
PV,AOX54T\=,21[>O&BH-RO7'>\E]7"<2AQNE"*V]^<V-_!(\4+2!.?Y!DX+OJ[HE
PS18-4O5!JOWYRWI\JSWM&75\NZ]?%R<RJ5,T\O?\O#1^BJF"0&41+1[?B-"CP]MY
P#X;-WJ;DC$* B1[/W4FSK@:-OE_R/1QO;W[1_0K"84D\K;XFE!4(^+=MK^5/%"Z+
P^+&*)F&#7:Q:1SE[*7/+J\.5D91K/[(=+E*LG%39GP B,"$[$2TU6<'&AQP<7*!)
PM(R"(&=R3<3:X:$V1_,^^]EX1E]PWR8?GL5G25!O:@7EBRYG\RW>=1XCMTT<1,3Y
P<7@;/FT..+3IH&(0:>?+V%,I5]"KE;9\RL!CD!J*8 0?(DH__"E7F?JUP?6=D,B[
P9+6=>HX9X<!FS)" '%4".V"AD@R7'@_.,;GQA3*7:&C?6_D2FLV=QV^4Q<D9);@K
P0P.TW1".KX04LGQ8S4WY@66#;V=!<)M(*XHR^"OSDP2<(91 &^?I@@AU?[YL2'L*
P.A=^&..\U1A81505<*&@;V3U4T+QB+XS#"=R3S38K9?,1\CH_E[;Q[AX3(Z=*U%/
P5(/F_V)^RLT)$-("SD?E7<%1GN>\:<O+<=4FU<S@($U5[Z@;>TG(^T;A$LZ).=]6
PJH"J<X_ '@#=NJ1/#US/_D:)UWOG7-4QG3RT2OGVP@.)ILP4BS>9>I<0Q;ZI2)9$
PT#;4P2D(S&6O:AEN/I(\5.=7X.3R\Y3CJ&JJ$\ZX$8N,IHHU3C8I9 ?U]^V!0RN@
PLIM#ZQ;Z\C<Q^1+>V;,,(T59:WS9RZ_:<B3V^EKL]Y-B@] VA[GGA]P,<@GHONS%
P/$3S]&[YH[?&U.*\+Q!RWW.@>:[8];%.($HA4P!?9M:B )J1)*OP_[>-XO+_V"9Z
P5COW->U?+&_:IU# .W!*M,Z I@$17!#9R_G/TT-JQ@SW,Q 5COV<UPWG16U57?P1
P0S17]4)^[,&TC@A@3U&/*79ZK3)64]QOX;'D<Z*ZY)(< &QW7[2_7"TL+3DT6JPJ
PA;PP &M6B8(_9[?Y$WP5P=E?.)A?3^&=]!_ZEFVSZ$*H=UYU!SF2U+W%P&+M=X7Q
PNTKIP6JA1NB'3VRROPY7M'.PU)?_K[D+SF4G[B JZH)G/K8JHO=#?:Y=)I=+Z@?S
PT"Y,K[$"K*^Y \L ]>@LVPN\/3 CGZ6'@%:D':XE^*RC#!7CH4]];V5_;-%G934D
P+Y!M,,!:W]%N7#Y ZM$1TZO.$RI0:>_$M(K41TZ)T!7:*,JN#!-<U6)V#FLPAH%V
PV+]35A3I CON:Q4^O%I"O[/"P%TJ<WHNU&F<0AG\WXY*IN5\UA0G_0A?S_(=EQM*
P[8E<CSK^J#HW=$=6=!O>TDZ8,:PS]D%J3G6-*Y-+[4B,%[;!/60_<VN(6P<G@?HR
P'GD!W#HTZ)J[K-&E4SRD:HL,PSA*_^0/H@4%%)9&P"_UCI)G6@^\?FXJ/8%\GY"7
PD PS7!SU1<!NRI7%L]7;T: 1;&!SN51&K=$$V-6Q'4BBV_)YR$5CU!@7.O\RH6H>
P.8Z$",;@4TNY>W1MX2I9.&'&\,$@TF'3M)ORMW-S3Z5\K?/,./;*N%*QLRMW*-/K
P]3I!,7X38MT<K6W*L8E+N[),$WE/M,BH[K(2T)_[,@L$IR@I9"G+KVA.HYSG!@^#
P[O'ZQX,+6$OM$U"X2>$'0,ZMBIFE/9K8(Z5\^-89VQ\Q*%\O:!-I4&8$)MVWO=NL
P B-&O<X&%RVEQ%6F,SC:SQ5>L)*2'WPM)\^8]G0BOIZ>7?%F6RM\'*-6'&D-BFA^
P*.!'@]+237]ID":BJ1[0(E^6DE,9+OR.:./,!F&3"NX"\1H4P;[R,D2=EJ107-WH
P=J9.U24;T-1\J*()];;F^6\OZ%$*P[D9D47FH'(\WNG /&%/6B>GI8^=$5*S&XCG
P@2F!8#;R$Q0HSB?>Z$["549<>;ZJL7^$_R)H64 \U/"90F(#1 "U@N N?6I^4K?,
P4'XGL^T4D4G>6^MX\\0O7J$/+)N5:7L/]=29'>-["U634-F]_T#NCR\7[.;CDD6]
PU=R9!-6P/3U:,"AJ()Z:U'ZBT>3W3&B3\BB,4;ON:H;Q33)T"T&%B(R0$B_ '%VR
PW0__.@M.6!"#Z("T!6LO<LC.IMC K+[MY%MB%G#8?W-314R0V=\IRT2]W8PE*]WL
PT5*8:/"RO'8SQ9@M>P.O7]BK1^]H(^]97$[]T BDIEI1]!!*3,JP531\DT5B@Q.7
P/4OZR#('(0_3VOC^NI\K9.;Q2.LF!50AY4*,=Y(7Y#>IH*.ICMF"&1!@3\#OJL*U
PS+E:3@7I:0E"+__)%':G!"LJSKBN48ZU2QK(SXG'+*!U>Y&[;P[Y 3ILQ#%#*$[U
P*AA$K ]C?R=,%C1()G6K<&Z_#1'H,9WGL'VSS",5YDMB,E[-;3"_6S!I94]36I#:
P8U/9?6ILOZ103NB2^(YTQ.34H,ROAZ*\:);7^E,:R#1\:]WSK+\@Y"8"F@!#62O#
P'HC=?\V_^#F>$%@@DW7F03D[Z W?YERV1: T.&$@'D:IMVL&^*OJZ_I_JE7H+<^+
P57:">6J"=3JK3%U!0C1T+70DA3++@$!^/;D2_)HI)>@#:S-'E AQ04H_V 3#/F$5
PHQ9J8=X=<[VJ^P]&(&(][8DJTP!,J1QQ3H\"T0SO]EFU9;AC(R/*+#URJC7+D7(,
P1SG[")E&AOM#\6T=*>4ZQ@[8[#MO(>'G7OV]<#T ;!F(*HI)$RC!%>%/\;X<LYE-
PW!S)37 +@/^U968+X[$X)8CD**NN>S0H49AF*<&YA!_)\U;<SCIA]\G8Y3"J#@M@
P4:OI2EN.F:X8IE*/J03?Y%([./R+5<I:F:*4KLKKEMIK/+$-$JW4EV$6 %&:XT0G
P"$^^R*:US$'2#G9"YL/$U=-@%,8V'I&\&NFNT,8-O]_.%"Y)# .'7R5(VL5*G,Y_
PZ^)F\_EB\?E79F2V^"69KU*!J$'6YQ#OR7M8 4 UB8^R5+J./9):'0'F,7B:=\%*
PS1KAAW3<.7<2#]0^=[BZO_\B;4_R'07P*/=NU;T;\OW)6H%*-?1!+T;8C[;CK'97
PS'N7=/%Z\&>TV'RP!85S*A*?!?\V 9(MO9UIJUN2Y%9NHEB$-LRCA+@T"OCX(6"C
PCWV+=7F/,^B0JL._:*=?JFHFD<$S4)W_!E?L8*<97=D?QSK*-B<V6:>K4PCZS26C
P+!2?K$6S,6:@?,>(L!HT=,,ZHOO?+MC0_KJ_;>AIG'&0[;>N-*<X6?;1WY=H$#&[
P(0XTB-,JUCITY9R[J;=5=5^F0%I.>YRDKFQ06=M$C()!9?()SO\K:*44-JA[!,<8
P<J(PCF<] &\SDT5=T!J:-D>+9O:F?TBO;\6UX=XQE]6PWQ\?R2?CMNV>?%#<P?"_
PKYYK&VUU!_H]T>E9*<)V+4&] =$,".KK[8^-FN811,@PTSY$6O5FUHW5@"G:]".X
P=3S@U9)*"VW_"$;!A"*+CL>:ST5+Q*:YM&,>51T'PLZM+_. ]:.HH$BRWA:CT62=
PU4W>P,M/([L=0@;&3&LD?8F:S+H1?O/06X/RN>2<M%]) \CF,VQ_>S9%)1\?&C_4
P@BF 4QL_C+S;N"0'DKOB.@%88^*K?O8OJ09@7!&HF"C0!!\4KVS#UUF'TW$)RTT#
P)AT1-,J)[7!/0\&J'F@&!>&0 7PD*YWNG'. 7HZJ$Y*G\#2L)>2WP,]3CJJ89^2L
P5^_-X>N2GW]ZU2J'W ]<D!=IBU-:,3$ 6478@[.#:M<,&+C%;*A<VR"M<:,;B@&:
PT%U%FX)" 2FF#<:G1((+<$KFE2UD'"XZPED,UR,7E[*YO<#F<N8T>#;'KG*8[%;(
PFW+2.(;ZR.7F4E&I$<E.C.H5[9BJO]N)178]80IIMUN!-?&GQ:47IRW>6=Q*LH)I
PPP3W>(A054F7+N9>EGZ[B6 OE+!,)/9K9\I $X3]@U3KAK&$2HH'.7"#$Y-?_B<^
P %YR/)L[_T#_AA!8#*]TYC)LMC%<!D:J)RZY7;I)_\C)4UKM\F/0VX!+UO-9>3*0
P3D#40$J-DN@V"D+F4@!Y#DS3"/,<%RD.@A/Q=WXS-P5"858=Z<UWP CLZ-X&^ZR5
PT[]^IQO%"ZJ0'0]UV"N"EQ\QU3[@,SNC"40/]NX7.<;K'/Q:&Z%_!/U-TIZ#6VT$
PKX*<<(Q>Z0^#4'W#EQ0MO8ZD/]N])D[VE4Z8V-7@G"F"[L27E_M8'-HH'?6(4\IF
P:4(Z!B"TB,$TQ_%?C:L(H'@E2[TVV\Y(TZB%\Z5F,:*W8M7Z34)TY"K'C"B#33V^
P$H9/]P +X$2@0QWE?U?T8\6'0^T97#AK5*(XX%9XA&SBNU'"AZH5L]N=A)DMQ<-+
PB!'@^HO4[SDO,X$+OJZ3-Q $:.?NK\.?+(A':R2),WX8_.YI?^S9+@'*:!UM95<:
P)1A'YL"W(DW9S]J:_U@8 .=N8KV>PW/2"1/,6,!?(YXC3G(U;19D"O4$0P9G'V;1
P=I!LQ1J!5.IA[V /%.6-[)B)M']UE[M75Z 10U_&=!+5^"X,C-*'K3-C%^9$D0;A
PGLY7!HD0G 3+1TTZQS]G0%,&J,06HT9U Z*_YZ/N0<(L'3[N(7[@@BT/&A6>ZV1"
PN'J+C]Q7%Y7=Y)!IW $U(RGNJ$KZ7K![\/S:\D5;X]=4<'0/^F7=K&O=D%S!N7.P
PT0TL<NNE%S[CZ,SZFALM[Q7QW"\I.HQ.B0D&W81P/42(MHM(.#?3B<]"\^(&D>;"
P(?IZ2<1OC",I6"M@E1A5] !MOT=ZU[]4B75P?C7M;/#&=2<:$3+4$T4^0:-WJ8M 
P%V3'QOR%Z[19=J-X9E&/T+%PK+=MB0F?>2J9&A4.&,5S!]?CK@RGTRF?\WX?Y5OR
PW9  W;UZS(@^RQ2L/5"TV2HT&!D%9(UD;%,2:U8^TAX06.S#\^Y(175$.@? .T.[
P:\''0<+(60E^21XJ[#B3T_]U. /_VAB4*9 KMG S*6<I,MJ-_I#/XU'Y0^*?+\37
P*7.TJVGS')<V>B@(T[YK?H7_FF>XI"7+?R)"@9B<382/6KJ5EY<L62.R4BZA</X1
P=<(D<FKE@$U#R_#G>^SY*!2I?'D N"V4ZM.L?Y/Z5&^[<KRG9)T3]789+[<YQ=.]
P>[[V6ZO@+JR0$$LDIBENB89*)2HT"/9+'0'Q?69?W]D[TR+CDE4GGYI0TVN7E+2"
PNY;TTU>AP5LJPJ4CN(& %^F8@E!=W>?I_O&T$F$RO[K*!%-;@'?* >L-=DI".\- 
P*6= S>D6Z MWP6KR#LY"A ^X_B"B,HF23RQ2+B9"*6[S4)E0D$,YBGLCR;VSQO$4
P=N3A:X8YL>0V?6RD[\=[6++>I(=#GH$R_J/^[BU5U\8(C_,^SC!!&(ZQ'%7(1("K
P"U3J8+#AI(4P7/+OD Y-1+!_R!]BHXVC'[B3Q<3QET,#<XSJNGMX@5Q^-$E@'.SQ
P66>PI<"__R'G!RR;* AE.XI@/7G+B$CJ-3VY\\U[2R[BU$X:IQ1]7D!Q?!Y<NI+D
P*JA5(Q_;*KQ(MWZ&#7$"DI/NA]U!LF=(+JW<Q>F8!08U?'$DI"RP%7A[_;/?U*_V
PZ3)D@,*3ONLMT0SO4E/(^>\9L.WH'Y((_4PT@/5[QG%S;OT&'%)'*8.<3+EX*C*&
PVR/-A;<,E]@48O$G>+5GM%'3N;QV12J* @\X-8D+!"NJR#<-UN*8\^F'/L+>$3!+
P3$4*KQY!#.N9XHW+_V@ 8Z"#O?#S5 1=;3=5(QM5RA%DP(2')_FH+H.*@U*Y7$('
P)(([6B%.3\M@Z6]2J@KM0]_Z57^V<N#9Q#;!;:G57.E(K0:1>Q]E\(C.I4_'4"#8
PRW"V$&-TKZ</(Z#5<#MQ@MYWKM3*Q<C1.7(-E6$!G4+&>S'EJ)'8DV+9,ZX,)AE#
P*(R2#?[NA*"D^E%9)##S14F<:+<!OX&?I88QN@P*9FT ;EH +/[V>MF!(&K,IB1Y
P'4'777U,% > 6UF#H?%P=;K\LUC)V-ST[.,P\]"X"QBE84"MR(70XII0:G*S02^1
P3^VW[J99="HJ=6 ;Y 4'ANL Q/3U[7M 1Y5!>)3#=*PP2.^]!+^@()I>?R5QV#A\
PY3M;?N8LZ6^[GJF=(70S)5P.'+Y*@/&449:Z2E:>H0")ES\YW/D0>Y2099<@?E8P
PLQ(I[)XETX8O[4XS/ (X^OUV!"I89Y<B%1C(+BIN::>3'N@1O4[]XJ C\?."'>TC
P<AF5YFU]TO3E$;= 6Y<E8(P*+MU9C/#*^BPCU5BT@MTQ%UZ7Y^:]#2>"JSMTM8'%
P.<F< &NYUI"(*K;*][K9LK5<^%1?BD[^\5Y(\[W?8_?%5OH9"SEX/D.;TNX=*$D1
P#']Q)@/LNGD>9E0W/D=(^_'=:5NN;GZ2EOI6W'^BHB))/HSPR9#CWF%Q; [?71<D
P+NZ'5HLA$K$F59ZGHM_7P*F-?7.[+5<T "_F #P& CP8 /N !1*U!F=L1XN2)W>8
PC;<?X;QU:_.RX O*0W2S,D0?60R8T2+9U7GYX D9DJH,*UC#Y"2T)7/>(0;5[KR&
PCGP<GMLQSHLHFW\NH9W(U<V%?X9JZ3]F;4*>6@U]U8>;B8=QM+EW7QXC(-I$+=JC
PX(-Q!$NN%QE>#9;PE^HRR5@1<P),&NZMDS:15Y1I!(]%*A#(5Q&/X16EU:@<0MCZ
P\> 93)(1$F!0RHYE$WI;,R;S:*BV^^_S8R%;$2/NE\K<_]K?0IR?ZJ(3$;E@,KCZ
P1('TM)Q4-"+LZ;-J:@3+1,#%[[<<HQVZ)350 1F">/;E)U/4KYE=)7@(2A1[_1#M
PC<PCK-OW6\T[ZJUP!KRY3.T$)4*[EO6W;?H'/[E*!J6IR>7*8@5".-2@NX']*C(+
P:BOOZ7T1G=6=>.*T980B78]<&_K;;DK6%^#G,Z]QH&D?S,5*>^G%!F11LRTM)[5:
P/E- .O-AY^6[8%EV_[ULW#!GY,?,DQN;I*.Y9B4#QFKY]\^S"KENG+C*49UO,7<*
PP.ZV&-HM5B$U6PW?X<\,3Z^#B)3P5IH(,>M8TV$/_;CG298;V/P\8A_)KM*6AP(F
P?K1]5F3%PVY_"H.W$393 _UNAS!<?=F$\_(W]:M;P<UNTCKESV\9*_JZ1Y6#WA8<
PH$1>V[;TXYZ>+JC$V9^T1?3NCCR)Z!U-1:)@O^T$]20.93//9IWULB5>F*F/LC@\
PZFW3&/X/#W_#(C=RF*';U%.(*'3A0KE/(5)992VDD?%N>=FFV]-<E99@9$9\F48"
PW<%KS, 3^_1@.ZQ48H2HC;"4S;Y#3+X6X5)*2YYAON4_A_>=TA]'!P8Q%/+XNX3?
PO2)'KYU$TNH$)AWE[KX&K0,=BIZ4W: -V/%?6R]L%TS2F>!_UJA5<^?2352G)06.
PT@@E^TQ3U0^00"QZ"[KB0JT<YJO)"?]U-8"0Q&, 6W!SV8!I#H!@4B^O6BZYPM>N
PQLO$<HJ@V0=U2[%DCO8#>#-6SVH/D93P=8IB*U_3W\R5NN[Z5"QJ,HB/RO76"67@
PBQ!X8=:HG=,>A&P\PKWOF)E>$3/R>-M532#D#"7,138F*-48TR20Y<7@,9AP4%SD
P[^_$W3QY'N@%E5+LDI6"'S?K3.WPJN?)R%T;/J0+#D!C?NA%)TJ7L#CU$ESS6K\0
P9B25'V*C8.UJ/*GSF +(*'E3U!OP:( 2K_:;?1+P$'&HL]QF='N6[SE1;I(\C>9#
P%8$>F8PX40>S8A+W&%;LS5E[7.)$A@Y0KK1^*2^:VBF[@=6@\-*'"?0J-QV1,,_$
P>].>,R+Q:(H&O&C2=:3 ;D#&.[$3>6+'U1:$ KA^GNFD!N H+:[5O(U8K<5*A_Y&
P<L-U=M(+!(I8SL;N,P']C2O-A&4ACY#PQ:!.IZM6PA6-S&0*.]G.)',?GL^:Q1;V
P+?A^_O9V9XKKW]_N@L2H/-.B?T!];AVIN>$\LX0Z:O;L>89 ] X/E&';S1#!1-_W
P#U%A?<._]OB/8 %A,Q^C^4&98O?>C &XB>%BULUV7R,+_ WO>7-S]D0[\.DR9PZ<
P8DX#FNVA^NDQ;J,XYD?VHX6:DJ6DW2J3X]H];. =4K/P*#H$X<8>I/W:O$/_0#3D
P45#0$H/7HNAA]-(UR+ALH?]7:V@JTO#IOGYDW__NMH[A $[M.KI8&,D7"C$7"] &
PNE!68,\G<(Q)$]9GM#IC6J5MC'43G;NJ346_M,-(=9_E8]0-=>X",SM1R&^#/GR9
P^(U1N:G'.U7+@0INKXD>P7HNJU/IN8:_>Q&6_S8\CT3YP8NWTE<LG+LK65UZK8'9
P2VC4=O. /VL'F8S-!88HNLE27\,Z#QUX'5<P&&67/W+(5Y>^[[KKX4#P*FO???6G
P Y %CR;+J*&H=@9YLOWVV;RPSTL7TA6>8Y/4*\?TGL?$:_8Q@;Q:A%?Z=J6FV \Y
P3HZ6?UFQO4^OKG]N07[!2G]L0=7?AE)Q[^T^YD\\N^F[\-YH--#  &8;)7GPL%:C
PA/T]\W)Z 45)_X T6=PW!D-9+48U9:B1"^1M;!R<^];93_-@:89[I<MRO"7#7QH1
P)%EL>%M\1XW>7J8*.)EUXG^6_H_,Y_/-T0-U+N\,^,3-".'7X_EG.4!J!6)TH4UW
P0E%*OQ^3CHQ<)]9J'&A CB?"JZHQX%3-2=HQ.V&9T*]R1'(GTIXGJVB.=*I:(YO"
PV78#:;4.O9+0Y'G=YW6RDK78[5.=8_<?&\H;PV?#8<9BZSB3]KEG=LWS"#P\B;8R
P&/<!].M3_=,O-_@?G+@,B0^!&^+;39K3HD.H/&4Y/C)2KIMF.L9KXTH)'=S! SBE
P [JQL)/;/(\+ZISXPIQ,^2GS!YYO_>AFG<\[_M4*!B1>4G^VR77!8+DMT\UY/5XW
P6G+:-4M'UT[D^#A9P$>+IV'$U2]8:*&&NC,\RWUJSE%R$C=KPT;C4Q^ ZGW:1#2K
P^<4^H'?)-\%@5!^63")Q"K89]Y.9F)R>=MX13/EEF?!EMBXMUSK2!UZE?47[>W1;
P<7W^RO4/XS'%QWGR,3 /U@LY2TG)'W,V7,:;':O:&_W.]/PGB<;] 9I@+FH(5N$N
PU$IB!>BSRUGHRE'@T'-F[E_,)ZV&,#5E#.3?=X"8%MS(36 _VG7/TT"PL+H5\>8.
P?!Y#5N#J]F@((W-I+T+3+-@4C+UEE&RO?5I[R7Z?;'$++*]6#YZ\3!8>M14/?U*_
PM;+Z09)>1ZONQNU)I7SYT9]W?2J65(>3#$0*VAP%QXBJS*@.!#(.R]BZ'*SO$U9C
P66-4@.%Z@HT!\N?O.,;(NC_(>\"Q-4(>X6>]Z],\-TY2#F(YLF'Q">[EO:RPXJMA
P_RA(@0W4JF-#MJ MUC-OUA&@AZC58=^8@)VXC\U![AW45KBIE$9X+F,S'"X#TN)A
PP8W946<)S8"K*H2/_IP8.(UPJ!-J>2$M.'T$.\C>+_WQV@%.*0+]6?T#;D@I^=:Y
P5FV9VP3MZF2^3?3]4]4"M SU)@:3?8MKMNX."R-GO4<-&T-UOL'6.E>[XWJFBRZ:
PZ;9K$Z.5S-3E@50/!MKUKN!\P[S.G1[H>MU;4HC.?S%L;U(?3P;HMHL4(.-44>)U
PQ,82)2UC(I1*,(L207H5R6+EP9/T8']V1#L4:7=A&&F0N#&JTV>&0HD%\PUV=B7U
P4&UG6XN@4?A^5Q7%E7)>D0$S$P H-CX-"%_*.J>X%C2K "!-74&F2_R"I(CS]KK<
PSRO8!JS$379DS'/FV%:]"1E5?TI8BJ1%FS;<G#JM9-G1DZ00RTN]9'L3 E=Y'(?U
P^>P?'==V:--I*#I;9OF;_T:>0S4:^T]"44^GGDSEKRSRSX@.5?872&ND6+*7KQNO
P8IWDWA ''Q!K2??#56,6VZ8.^J"0=OK9^7LD(1PK%]CYJ]D[$719=$JV7@1=*;""
PA*)M=58(G%"(0B0W@+ [:'KYJ"PTSP%#4PNO!OHC=')GR9W\!E# '@O6F4T8&I@M
PI2/5/QE"_Z>H">V+=6&4EP!DE,#SDC>NW'IUT+56"-!R,>"?Z7Q'S@/D1AM5]"=F
PEN\)K\J6J5V4-DL:,/KHH&4I)\C1M<AA, />QV#4IO13,,+-<$%Z13^C69S>W(G2
P^)+T@G_'S[A(2)NUEXGAWDP')_  >A//EBW#1>6/\>0+!*.-R#7PSRQ6]W 'I^A\
PT&^_^>C?V/K$EH./%0=@3\I:X$K12"O#,+MA8K/XD(&X%*7<XF+KMP'EN@D%)A+:
P",@YE*/?NM1JP>&L]=?OO\*;_ ^5]&M\D KDH F=;"+1U6!YP)C_&$G_D=VBW.JI
PP]>"S5)@$H1%1X,+'FCEZC@:?V> .7;OUW#>#U0BY^GV.(SZI:LS4IA.9$<-^^CE
PB2DPHWM(TV+7<CF7MW Z#'EXE+:UVSGGC S=MND>&'!3OY@DE'(OSS-GD:QUJRH8
P,8)GB./%#E&&&2#POQ&.Z$7 *%'=:\LP'8]](I%MF.,Q*EKG7USNLXLP]7XH$E=%
P\OK2B\\TW56C^=<BVV6W:V&(/GH[G;E0+Q:6^"_MLYK?7-]O:0JAK= 9DH_) H_$
PW1PG'%'\H9^:2WW\A,]?V(7Q*SI/-\-2M)]!H?]"]Y<$\-VD0_WZ<ZF'R2.+TF?C
P@P"AZQ4QE1;CI.7P+;<-]?&#+F-0Z99#F+9"^[3#)8@"0$_?0579/LAC^^^4OC-.
PMQ[@T!=#9P>XU# [73VXY,B_PD6R: V.DVE:D'/,G-^.EE)%5"^(C"(M27B;=\<T
P<PQ8;C>MSFIOP=(6 <&%K+&-E_Q,.J%02OH DSQ2[<'6($JL2B7O)QV+GRPRSO9H
P@T(.8(ULI;WGKLZ8YI0F;1 $C'9RJ[NR,S8*VD]0PC.>L.<QMLMO.;R:#J-,FC=@
P6\QBU"CL'KHRYNEBO^%S(;%O. &=XTD=M1L=3<P)I"3%I8OB@3.';M,IYA?$]#QX
P8'2!3J].][H\HY-F!GM$=I6ZU/2F.>@&*[5B'W<0SA+@WIV@]C[M;8:9?*-J^\?.
PXOY09JA@%0#>VO/_=-U:4O/EX<JK+&KTNQ5=IY9M""I []3H4Z5CUNY_:9CGW3(D
P^6>_"'<CFZ?^&>^*@2?G0'EFCFIHFEH(G[9$R7;A?R.[?@&/J48O$\!2<R+#$S*>
P7E"2N##ES$0^-3Y[]=S@$LC53/BTG.63\7P+O_=M#+?X1E8 /?_9Z:/+O&$+O#B,
P]$(*>EO'\\2OY1YW5IE89W,_*G/BN&^(ZUV1W.Y/P$.%=B.3*%/1>-7%MN?!JI_*
P4#F_$#G7, W".D36LJJNO"(W,;TFP#8.M49@[;/#(P[>7I="\1XZ1KDK3->]M;!?
PN8I:$'A %"_7F/&%LP(VG'(3^K+;R(*@$8 B;ZV1';K0*W/!^:D+;#WW=U43^ Z'
P,E%S7,I]TN%I;*00#R]/G[D$6,Y*7VF-,%@ YH;FM1%(1X[15-AIR/L7&B/> SCB
PY(%]269A3N>Q<?DSD*6RGS^B%#'21H:*U)7&T8_'O6Z$M&D!/(RT%6Z+9KX[T'U-
PVM-TZW*S/ 9F/#$(G?F7JM@9?Y^]TN0WMIG'C31<,<-76ZU]TMP.DS+F@3_9DGS*
PM. [F@:&7>!1_R)>5(O6/"JDHS?TGR +]0<"[*K,M-B0_Q'U2L"U)G>#YUU?%XDF
PHB^AF;U/&I=M@)JG1J3WC0VYP!IQO 5D]W/NS[OR:#5MTA,1\;(\*7%/*O3/A M6
P3'U+;1#-=3_)X(NH(F'OX1="86+[G7;"QGY6\W>TVY0>3C*F6F(61$[)DK"IX>6J
P61Y/6R!/V2^"^;<2>2\U[Z+VQNI"&Y9RPPF8)XP,N'V\O_EV'/0!7"]WH'>S0:JJ
PV0%83>*3R*INRP^CR/<#&6/\CF(@"Z"B05;3K6]O@HX 6F<@1V6R=44;C 94IZ6=
P>OGGX4?$A_()5MU^D-=>$-HZ: Y3![+1VK[I-6+KNJ"!F7(HD:I60)["U;PZCQ<-
PAMA?G( ?<O$P=_FNL+_.MP9!=)2S8/6J&&=]];_YY/CD0''..^/J:PD!M]D]WG::
P2S'(XWP>NCXZ.0QY*/IKW!*;@C2$X07X%(H&WGC+5!:C$U'5=;N4D4[4#%$Q2+YK
P2 ".E*GZ]""FKU$T3Z:5H#JS#1\&@GES6&1]^#3;=G-C$BGU=1J=1!$HAO*<JXC_
P*0N\&K?GODH@DRNKQ74/.&^NCXDCC0]ZSC8Q:82SNZAK!'.+J]X*ZH7 C_'2N$2)
PK:KKB$M&8BHP? O! =GVT[X4M ]4]% AOP]Z0$EP]:G?C5@A@44NV#(2B0\D5QN4
PY$G^9_1DC0H7X\DT&G?G3_"6F4GP0[IG(B[59@Y<'ODEU.'$FDG6-MA9*/L:RHK:
PP2'6\JL:BH^X=4.N?( 2@#G4T%"\UU^Q%9/SEVW )/$+8+:[8(;BC]2?=3FUJ/T!
PX< E8+"$K"EC4:4*8'LS R)F^EU:S'I>,K2$1%23W"T_30J4G:+$RZH>L;.RYY'T
P47>L5-PPOG%Z/^GQWD,(ZSR<6&:L#@1&/*P>*:Q%QQQ4V<+-Y?@\_63*V-RH$79$
P!5'AE1M*8$!MEP\0& XE^_:Z-*69!:1D'@,)32/IF(0WRW>[+MZERJW^&J@U:I7;
PJD>)E\UAM6-XL38U;(F)7* HH"BD-(LQA@K MNG[L3J4VGDKJMFJ, H62U68IB[Q
P;]ZADPMS^;0VDBD>0\X IR#\,B^J?UA#/;!8!]>&N/1&(@V<#1G!<6K@=/KU!>KH
PP"V%KNK6QZ^E+H.@^-L-9.HF*KS%.V<)>\F"4O8$2"Q^39=H$TLHX' W))37CB1[
P#Y<3,, =MM(98SG'VQQX<')P1/ZCI8A?Z6'.5GT<J\DHPK@\*%D6'?R?Q')J**) 
PT,$+?2U$#G;GVLJ>5GVMWU+' 5@P+)M;SX\.>S@(]G %(XXWV$?/]L=QR8RCZEWV
PMD#S+B^MXN'+:W\W9V\FF4VQ0!L2#7(GI8\0?0^*MZWC,4)U7CX;<2)I,)LDOUZK
PI=W*W[[LL3>L"5X97=GF)AZ$+ 20YL)/2*%WD%,T4F+3)R&V8J^M1PJ,1%P]/3@+
PI69?.1=@>LES$)]'Y3<V7!+5\"!YV^$&C)[+GH+W=A@MD^UXVI3S+]"_,[B8R;2F
P+4YI6W=S3B<LQC'_[R @Z%B=N1>!&T3Z'1)=I:3&.C]?@UC\#D2*(4UJLE60_]>Q
PYAA^RA(ADIT['<^"@LU][S&R8.)C.C*K_QU^I;:FCE;$8X>IQB!#<T*=)=M8$:QR
P*+"&E^#/-*U3?;)WP-!L,E R,"DUS>TRJCP:F4#><6LR&'MOCODE[TD7,5V"!_GQ
P2O02Y?#GO#QRGW+F.O&U40<H0.?7J.[5[4L9"RH3!#$J*!E^_J5[ >J[(]218?*=
P:9,7:D=BW>"E(^,&0XGQR8J.SQ3)67JOM,&]^42F0A;L0^Y_P/08^Z^P&\62AIW7
PA[9:08U'F(<GN6*> @%FRLWE4IW;GM9U?9?6#2'&S_@(L\I*=8?+(CNFD#DX;*NO
P[6CZN?18U0!RMF -B\QIEC5&P2;H$P( 8]7BHH76S%BTE-)7(J(KSHHT#'H-*2PS
P!(8-4,IG]L->,Y44//-S/\27]]Y10%S,Q8:9@)2\;YFYY.(H8+JU%;IT1K8@,0#W
P>Q+L$D[OY@.=C$@#L(%PY&[YF6:E2][^VB\X(%YWZBO#>DXV9FF*7P<[RIY[KT5%
PY:?MDE_R2=!^04]\V')#Q"K7V.06/3O(CF&>O9#C(\)W__6[P00TW[)PD[*LX[UG
P6(J+ ;[3!D7]Y2TL2A3J6I,*Z#P*P%'%!%93074I'00YFB%7/G:(JA1Y\[]L"#J/
P+JHT@:XI^N,/E=830TTMJ9<5!\L&6#QOYO!(F&:3[<HT(C](_*YD-<RKGSD,:&5/
P=6 RE5U=R,B,BU),6-TNJI" VZ4)MS6 ??TGK0?.AH_14"4C#!GT>=@-[;*B</X6
P&0:R3[!>E^Z@TTA+]_[$-M&HE!IY_B:)7PSAC$@DOK=XWUTZ+SE-G=MJ?[.+8\P?
P\# 07ON1CA2G ]UW$8\T(8HJM"?E=U9O3_1CL^J9&58UH<>;3X$HA&W8>97[@64J
PPG9C@GN0_R>4Z:6^>OC'[]]+T3:H-S;J@TQ'+&.L4,S/[)SZ]Q^M/KJ#-8SKT]Z^
P<#/S!)+&\T85# '[-W]V;Z/HOXCW+_MW4[>S>(2IUX,"T91RB!>O+UWD$O:C*750
P>7TQ2CP*$6=A%G;$> T9K=!$^\4XOM8--1U%SM>4C@WKOAVF$-6B>1NI!_<.(!;%
PU[YQ)S%\*M*(U?554,2:U^*(@V'+4!^=Q-O9VZ&8B%/K\RW66.,'IJ)L-#F.(N5T
PRYP#6X2TD#IRL/MB(&C)NRE[K-3SX5FJ.\A',^& ?-Z8Y90;JL(X+F7?82"-U%H+
P\[E_ 4:AEXBYP]\G6$!JWVW8Q\PWM@&JB4_9W)9P/=0COUR _(=9A1X2>K';1OJ-
P8PQY>:Q8=R";($;;EG\YS) E\94EZ)W0CN1)CL*IZF*T/!JJ9I]0H<)'/I^\,!)>
P$F^+K@OR(+WIHT^6 NL-?32GH[!+26P04]U;MD4:;T#EQ1P/4?(&LDF@VQGB+@!2
PVR3KI$=[,&J)HPN%9"'C0SNP'PECX]@'+^<G,NT^5ZH[*--Z$S@Y#-0"(!%1XW+Q
PTG] I?HBR6@-1.VB:R']'FC<'\:I.8? <%>P9L%20/DOE/X5*Y/Y<P!"_VVU:Q\;
P4N+"92JQ>DC3[=U*EL($^YBT.OK+4,7,P\]'4I5;['=8@0C<AM:%*2[J)2FU]<K"
P#S:9^/Z"?W W-N)O*QG6U"!X[+C_;_7R5['"S<_Y++.?[[2>56OQ>%Q*%P@J$2PV
P5Q7$-T"SZ/L)4:$62W>E^]4*BL+@PSO'RQ9T[U479&PN# ]1)MIKY;FDS 28\'H6
P$2C>NI]/K=XM8=']K79.!'!C?=J7B8Z"=%7OALEPVW)IAQ=A/=1=S.L]YFOU6,$7
P2(XSRS!O^I%W0J7BK4*426JQGC%'*[LM_H9&J&M['SPEKT/ZD/2LP&1[Q"6AP52H
P..-N33,G<D2%E'R<952\L(!T2!:(8VC/XU?CK&ZW+AR^(J--O2_6P9_;ES,+I%\5
PV)IXF@6&F.W/3S*ES">+NL=4D.;9Z$9O9'3BENY>)V0R.2N61X55M@T8U%;?YO-(
PODF;&2H<N'CZ3P.U&4@D\O+55+5A)/8 /.;FX%;L-H<XDMFET0A !0B1[9/==W6Y
PZ^,-K32H?Q5ZPKH+DA:O]00'J[?-+E>OZ@^9;$ZZV/Q_ZI&=Y9B$F86B![CJ?+[<
P<,86<BS]EZ1C='.+*8H')UWV&THF7!6)/]*E-4S\=^VS8'M!286&]DY*[SMH[!YK
P'JA^@<@@TQ8J]00G8@0C-Y%ZD]\Z*RU=7\3EZ!@:Y4*>5^RF.[#@N -X#1^BJ(7M
PZ;1,GJX[N-M))K_6#L(SY6( 5M7_URO8BE2AY!+H@9LU!"RL1=9WY*YQG^VC>\;/
P8IJN 76X1<DHR2Q.Y*89.A@'"@Z/JO25.?,.J9<\90'PW)&+7=Q1=53[KI0^N?M#
PB.=&7^DF/+>MS!UJ(Y'%&,[Z<8!"!!?#)8)/NFL(:-3MP#P'=HQV\3 ?>A".93]5
P9VX5M1S@ O.BA2"3].^YQG!$<7L%0!JN@C"<BET6[9L#'3>O!0]LU12H5[[OISM%
P0#B>D+T0#CM9!\S(@SPY@#<=Z)E%NJTZY79E(]SMKJ';]"<!X&>>V!UV0+T<(AI>
P35W95%39X4I,@;/>!1Y#':?N<,K8^BR.618*5-ORYT\KXGR@7.2D-(@T?Y@@+/&F
PS"3.L'E\6C([YWQ859]C=$(?.=+MBJT^ER:?MZ SU!'^8N'A*)V<372!Q@7LE+6A
PO%DZE=C<**/K@DO(CAK6R-LYT!/(IRW4+"B/]2%:QQWQ"M2?_9*X4$(.>11\D8V8
P"1RRU0CRC(S>N<X[=]E2SXLG:.D%$UP50]O,> ERF2GOW&MO&YN_$Q"5&NF#LKEV
P1[-9AP%,PF'=18!M4 6SSPK'2J/J#KQ/4\E!2/*;GC/SYTK"]=7PA^#JB\]RYDY@
P'N)M@5"4S0?CL-NY+61/[<@"OT1@LJS42@!^A&"V=Y=!_AUM;".7;ABS:68"XKV*
P29K3UWA)A0:A?@TE@/3?:"&Y MFBX!$FW*'?U;168GWCEN#-'0H2D_P=#UJV)6Q%
PD\&OD??RD3O#&W4@L:4#%Y[F$;$\=F+R&4++ J]SMB^ *J<<00#[1#4(X]^<>J0&
P(->R!><,.W @/UA+FQ8:-M*W@,1[!0V9 */]L\ UF]/'^Q0HDPR^$KBP-.L3 /-'
P9]MGA#V]18, %%6(DB6FI5!WX)N)"O;3/5V<D*[TK!O\]<26W&<K7-IQ3HIT568=
PJ!?/']\ \<M9OW\7]!W!"VH>.^(N[C>M%'N@V4.3F?GP-:.%YW_P8/!E4.'[S6!;
P^-HL0\WK^6C&C79I_RE:O"G"^BVRP,8[=B[=QQ:'$C#HK0:M]N6JP^WL<4_X.Q+F
P\$99JG36 W?!5L:%J[DB@'=I*QHGH$TQA8TTJ]<#4_4U$NT"52HQV*>\G_MSJ9)U
P-U+)VAEP+]--HZ_]0-E80Q5Z!6('"IE%C[2T-<<R>>]8EQM7%:C-M^=HO/)FFFC9
P1SLR/#NX\+X0FSEJO\%MNL!/2<O4#C4L001?$^8NF[$>H!A"];.X.%;BX]$!_&P/
PC)U3Y3I@@*VJQ%&\:O' ]-C9@:67B)H:((-F+'>%1WO4*$-1'B:HH7?J?KY'4O8A
P_&@41%&V ?GL9>BT-$Y%?$T_FB7LY5IA&<YIU4S#S&P7T*SN9=<+0]$&,]"X8/B&
PH"I0"49FM"0O.K!$OX=R0-4':Q7PK4:15"!]V#]9/3KM]M]T_];[Q4M"*I&7_F#5
PJQ!"D)W(]1+Z1!_6.CR]I[HH&FR^LX\;+I802,-&TH9^7;RQ#1X;"E,GDW\1JSX'
PP+3C.3',D<-1OW#D#"E=&C'QNBMA4X<%X$5MUO8TPM4>%E_I:F3F20O*K,/JAX!F
P/5;9806X3W1<G$0WJ-Q/!)#_:#9I_:3_-P-J9S1N'S[%1%CD=RN[5Y%>FMG5B'QK
PD@=?/DW%)_O+4%R JQ_-C['^GIWN.L(CW3>Y*V1TZML<#NYZQYNG+2'!>(.>LE&9
P-K):4=]SJE]@%[0HVUOZ@$0)D-W:;YRS;?RRY#,\4"#6LJ[EL1A7JID))(;=I-%(
PE:$4A;+7Z$*-CU"Q],38%$3"#HCXN.Q""%6ZUA(>?$>S61U=FA!<0BCWB%%_GF.5
PI>1WAWV&1"V?H]AL)!&S+D<,8!=V*D'GG_$#7TJ[O,D8-6=.+M>.O&&@F8;BWPQ(
P7:D_.__5RJAF; [>?:U<7V^UZTQI_1F?=@OGQK]([8LBT8>Y);N6&?PP(&P2OIT]
P=TK[ ,R1T7PFDV'0#,;=A;5!(TFD-"Q1:ZE574?L57W#+!U![V=9Q$R@7I9%TF*J
PC9[C0D03GKKC]]M3&>T@1^CR1F'X=9^&JB.@)@]734F@E]O;&=MTI:DGVALUWTK'
P%TTT[\5>)B_"EYE&T")0^XWI0?1!NSR/3&-<>GC*X+NG6G*)D=I[(DKCP=-.P8-,
P(>I%D.8'@-IJ$,C4*VJ4F%!.\5IN>7I<O)G"N@5CMJ%E&T';W=$X.^[-+TY*%A,^
PG1)TGG+G]:WDU-'7LDWE#:2-&IW%=P64M3WMX&:K(@UV",LI05IFY!"T#'8L/0M.
PM+'(N3'NGFDXMF ^(*NLIY^?&!XX$LSN@Q6*T;9!Y!F'>QN,"*;0A&WOY]==!Z F
PT@%LA;X@6OB[6)-Y@/*6'-1H2&&-@*B0[FS\&[B([!T"'9:,>9%H^=0DG0U@O9^Q
PDXERCI1V2E9%=MVME2Q^$:X8[$7).G'^K[ERJ+5>VDM)M&VCR5]1?\@,[%7UEX1)
P.8BP-B:>+.OQ&(QF)?#>?R?_#5>/L(,Y&"T !_*2,_A>.)0P62^0'+W(Q_!-T1%H
P^QS&TA:[4/^6F>$?_X&/A77(2$S!['-,%LR2!O,/SB7/J\ZX"HX2EBPO[<Q>< (:
P#*R.2F6\2874OJ4/_+5Q ZRP79/,,FIT%^0()^1-<8'17<;8IAE\$CBVVXL!>:F#
P1O1UCBF/63BOY9FW_O< ':OL:V8N#F$K/>=8ME0!F_8G>+5<,AQN!4BT+X>S ZM1
PJ,?3^"I>?/0(3')0JJ._S%O=/,RU>J8]V)V*'FN8AA5B^)( \N.T:8V,[J>.'RLK
P&G#_]]TC_9Z9[_10O#98+B#\.7.X%J&(QU=+/VPZ5'>]?.4?8>+A0KX6W9_N2ZT_
P$L0IH,.-7TN D7@@1$E#5Q'[20L)' R0L6L<0$1#K=29HWR%#KLZMC(MV;RG\=,[
PH[BAXO[E=!HG#GQK3#]/%[BT"WCN@=_3L ZK=,#5_6X[RX75OT0.1WE:5ZJ5QJ^S
P_W*3-+]!!ZWV!-J^$FW\B0V]IK864%^3)3:-QQ&.J?>-CX_Y9>L\N:G._!4R+7K(
PLV!\J(#FP&)29ZW5?<@KR3C/.;2,,K*5#>KXOS/*LPX')V"3&#-9$SBY7_OQ4S-C
P6KOFF+_#M=3>$Y+;2U(CT.RI]5"<W'7JN3&*#_4L)Y?$7[*O#$RU/LW+A4%/XOG&
P\U3@49:!;:^!=,&PD,@MHRX!T/3)=)S<JL"(WPSJQ&2NBY^ A5C(@XB<]K:?H7<Z
P[OO*^JC^ HSD44#^?AB/<+)J7PA@ IQ.J7M =% -O_?>C%1R76&BT'ENM'F!FC<8
PH<=[$[7KY0';O4)[F(PG\>A<G8,/P[&1K<3-)E191PT?\/:\846PUM"1'B^)@VL-
PTL$=FYL\'  Y545Z PO5894ZWT5(,E!6\Z>.R#.W^HU 1]K5BR: E5@4L'=AACQ_
P'S%CI8QL]$TS!(Q*S!:Y^-8T+6-X+VIYQ.=@-\)O1WIU_/] A_3C4O5UR\%39S;A
PQCUK'15F%Y]^Y5;2'O5DU!<.M+UF3>*OQVMGRE[V&GQ]O?6-@O-U;T?N76*C>]]2
P(=VTB=,)7W';. J +GII>64&N;QF\6Z&M;L3=?K/*?CZ]NK.8FM384%B8W%27\!'
PI?$L!W75L"5&<1I4YNU>4CSRAB9Q@%<!_KO,)R&^833?;5-9M]NRD),'^MN,K5^O
P+=;&3Y)6#(!+J'W<>FR#%[O#O\/7N;HG'X<[ !,&0T^PQ][T&\<_B"(NO1+3VIX(
PCDP#.+X!1:B( U=HW@$+7HX8FLB*'Q^EV=*A1G>KN\BSFB]P# ]#\MN0$)+>=AT*
P*97X/!K9UL?%$\OXI0;++IZ-<\.@P (#B+PEA]F,EJ^$_8_HE#L%PC!^>XK8%_4H
P#M6&CW?SH@]35NULP0?P?C3?^&VU@0#]"7?@'9'Y7724_F%Q/A7Z<K78=-[\IQ&?
P"O49@\),#>SRK8]:EJ7M7734_.8_(=X>@)6@>41$Y?IR<R:_EU1\&L!IZ8<UQPC<
P]4"]"?*#45>2U>K!8N5U%MP%E'8PC 0P E?V%Y0!#%O##$CWCCGRWZ-/XLXRZG"L
PU-V*L U@FT;@2UORZ'33L2>:V(V2/N$)F7@8[J5!P@4[.,B2H$ T"BPJBO<4)U_N
P*BT9[&004E96*,<'SE3C!WR%S ,YKEBY+KG>*# 8\G-\0-G31053DJZT B^D=[!I
P7.#L/ZKSKH*N/6$#C,^BG!3N"1Y"$M)'XZ,UF;[Z>(IMTXYU.\C^'P );! IW.E(
P6(;<JK/OQ )E]-:P^V-Y6R,][DU[\5[52?ETZ1V^P/]ZX>\@$R4<CXA!O.C5&N4A
PECS?$.\@?.Z/9QV8":<UF\SN@8!5QL2N8:2FP$T^NLI@JAGFK6. HH:52Y')+;!4
P_QF=L %<\%JH)-J,C%MWZ^ZATZR-?G\Y5&0D8C%TETX9B)NP>P= XYH-@>-WB'ER
P'G'H\G$["-:&0,XK%S\!D3 VW9C[5!'C1A;LN[;]+ #&L%"H)&FI,N((0EQTZ0LB
PGWO^.PC?E&#M3K#4Y8&7=P2P[V R!\%97Q>(U%^]#(*AKV#[R!C3ICD5-36VN7=0
PN(8@K.*Y:1^AIW-)PPUU<?U/,AO4Q.*!:^FJ)$I 7^QXH 2;,#9?[=^/"Q#C5/DK
P>PIC&4S(<%17:8;# $4UFPCXPW4*SO6JE7];D!36AUH&>*_6EQAP1[\0P[!5N:<=
P%HHVM<W4NL.B\>XM*+1*P_?G@9Q\-'&C3Y_IH4T]#-KQ*:AB74'EHE]UUX\6/VI7
P@>?9XBAN>S;A>J!J.\D!9]E7UN92/>8^!L<X'JD <1#S53B(*28RE)T\Z4$1E-..
P; /H9!8;"1)]-EPVE,S1X(FH;VI 1BK,71?==LWMM:-7V$!/BJK8@^KXN&\+QJ8(
PU_,J[_!0DCK7AY?PS2*G>@@U<435.OYCW%0]+?1K70N?9@+]V)Y2H<.<920<;L"R
P/M8#KO]6OOJ&V?+A.W.M&^I+G-!R?C$6"G"10])UCN+8WKV1\G=3Y-$9X@BPPQ;)
PA\@GNG5O@U#V#!H<)M%^$&*T@_U*F;8/IR'SI]GJ][!:CC'G<C;JV+I[]B/L40?U
P8I:/''M%\VP%2,OV(N&8"-P*W!Y -2!FP8%B5;UATA&XM: .U8AED!H^8YJ;& =R
PT*+?R(Y!* $JT%%L;GVNF5O<A?VQT\"74R"0-V['>74FA,%@/F*./>KF'@\;WC/>
PQ_M?YO[/-V=M;VNQ_NP26-L$!VN0;4\KO?AL 2> >NO#:J,=?<NG.'Q?F!MZ(+P2
P /$HS\$L'A?W5VJD6@#&<;8W4'(YJH:5+&@T02_6//9]U91BQ1@<<FF@^$Z&59EL
P)R?RS>N%2&1VJ N7>VMIZ"*-!?V/>.!QM.__[ @12N6A4XF*$$QL1DTB1UMDD9-$
P[ISUYM'_&2313"6J0. /]ZCE&%O,&V?3WRQ/%]T^YF>0%(XY-?# 2I=$CK0*2F^K
P'3<F;<TJF<):E(P>WPB^)W2.S+8R.70D?"9^B.W=T]5T^6EL'YJ5!QBM2<AG& =\
P?9>)?*J<4>3<%\VOT.-J0XX*P598'HZ8UZ>8M-11G)\RK97$X:>E,#0P9\&-=:=4
P>G+%R!<\)G"&V:FM=D^EW^T&D"=?[70#W3)>L$<BB=<C.9TN];QW,.=I3[STWN#-
PYLGLE=RK3I<"W?3>]@<7X,D(Y4_\F"*YI([E@HE)#A(K$F,C(4%D&<.YRD>FQLY*
PU!^0H$T./9FA8>I UWS)E@9N!D;]XU7Q.EM[H$V._V]E)M,60^IT YV45MVT?^$;
PEZ/7ZKWA65J6'.1A2@YA*]\ER @4_1E1H(HM">V@.TZ-Q44Y($ \RH?AST0 R'@@
P;1$!F';S&P W=?+ 5*PULB!O#M,D<RE=:PN2CW-*>_>=MX!?=(!Y(''4:/*W\ER@
P-8JO&^R4C;<0:*1M[[@XN"55JJ-V.)KVCB.-#?P]/@F/14*<EFP:60+ZJ'%#/W1#
P'$I2=M"^\]9R&,Q,<"3(E7TCH)@_]Y.,RC?@%5B6'7W7.4U)>^AXQ8:QMP2=K5Z$
P@%5M@POCI5IV8-M@)8XODH_5&/MES601G'Q,O0?B6[W9FJ\0/L\DU;!3+=_>BIF<
P9OG,K\5<M;# OU'>:9&4QC<5X6:ZSP]9G#25GIQ^,3D>S??H')[8$=L8KCFG?1H 
PT *A;DC?]>SI2F\:D,U?_GA-(::3(#FP^,]?%T:7*;.X4>"ZBVXV<SK*PC"KO0&:
PZ@A$9'/[S5*N22R"*'50:1N(P@HUWI&D?)]/O_[I6[#/,9.78_Q&NAX8E1K<OB1X
P:[8"?TA3SVRS32DV6<+;+K>?6DQ%%(U9^Z_O-):\Z-A5<1_U/>PRZ[ @KLZP;JSD
P.J0F:AZ_])XF-8:"='5XWYP[<<!D0Y%3_CK:/$9C8!KNR,;WA"__UEW5$>VJ&IH3
P(.4.$\(0!?NQ:@.@3CR+#)8STK&YFV^GN<5]I^[,P-!L-4UNN#<]N6X#R-,I+->[
PG2RKJDRS$>;!=E7K3 JEL_>QY1Y\.F4A@:9IDIHQ91V!G*$78D_+W>*TFML\?0AK
P-ENQ<P:C^5_QJ, >%?@?,X851;#-Q1IH]2VXO,MQ:W(R^'<J+I'**_?,O4Y\ 3G(
P/VA&M5@4NW6%$LA*3%!3]@*E/-7*L:6<;OFEK%:U=IT89)7[<)7MMKE4G(YN4_Q#
P+)U-+<P[HBG?67/85'NY0*8ZGBS._EC(-74).4*TE&53@!1T'<#YLF?Q32!,V\W-
PD24L_! \8&ZIR9I_#:*RTQ;"]RM'R:5(7M8E_&:V'L<=2M#N$JX5G:>)W?LOO!+7
PP/C,43FUNR=Q4PXU3BK=$6V\:#5RD)XKX2A]W<*I7$+F8I)BI6SW)=5/0JQM?,6Q
P7HE"S]R8[[4#L-&$2+RI^A$K;+KJG_Y\S+7YTGL0'VCV2[-1XZ/@FONGQ<$'=LK(
P;5OHS619U<6._2V(K3(C+RW07%76FY1H8!);7"0Z#1L0"!T761OLPYZGZL@3U4ZQ
P+L--0:S5V8]$4UG$7^C8G=9'#MMV=)1,X)DL\EO1,M5G)=_!,C:7'YM36!17?B2U
P29:GFM8^Q3%5@G^@;+JJM[R/46<RQ$+A$]#G11V B0=9@XSA6.'4+E,-PN0/PRTY
PXFN28E94E(0ZZ?<.]V6- H"Y#N.A%7,>:"&84\LP"L47+T>'8Z].0=DBV*DAL@GV
PT7N1F\JY2NO[3:;[C>QUEJ!!7<4.*Z/=RW"I_)UPF4&!)ZL$. RSN*0:K@_HZCU3
PR&@0^N6:Q>O1O'GGF9&/%J2+D\N4HM.PK>G <KT-M=Z_$Z,_.U(M5C?W>]O TJR=
P3KKOQCX7];ZCJQ%-?!7(+!-6V)3QJMR:-K_#/@"^=-A:C8PWJ+?HLJ)!Y?4"$HQD
PL$(A[*@/SE-TIN8N\AF[J^JX9'8!"]B?,K;SROI49:NR!#UF'E<+<9MNQX>F!0,?
P)N:B/H_OL1 2G_6E>1[Q/]L+MV](LIYYNE.=^"^+"N#E<+'%>M&0VQ^$O$%,:PT;
PE()NUP\I[:\0[JJ$J]>=Y'A45B: IZY!D.T@7RK^N+8I8KHH-&?G!+;O]T7MF)&J
PC.O\%(@WJZQ[S:O\@5J_?-!&QASDG7M$K*X8=+5&'<?X,6_?A4N]N.O3Y;_#H\$!
PCAXR.^,!&WXL.:F,H^5'8&>1E)?RLA1_G,T@]^.K^!0U#6N_SBC1VBU5G=L:=YE4
P\2;2%3M0P_S@!U1ZUM>-&9W;JH5Q$W.@&-\I@K_L_U*TXTC8K3M\9!>$H7^D96??
P3@W-.!^:(:Y$FY1MHS? ?J=I\X]T=/G:9CSEIC/+C#M;L2L/@,'A;##B$GE5<*!K
P#)_H66?!5VN]ZH41P![\RK@5_Y+>-]09K31KUC>F+U]4:QJ2&U\2!V4]<X>A[W,'
P,Q2S>9._1:;05=J_1W>D7(F =$@$;A3J4^>O:>D] SU7.1H!2[':M^V]JXET-VTQ
P#2>RZ4&592"0?!GH82"WM(&V-11 I'2UJ^G?=GS[6+F6?'-9=%L''BEWO+TMVJ,-
P8L?"FY['E2=O^GYFE#[W!%"HH3(R.-Z) OZ_OO*$<1WPW.I+:;)A#"LI3+3=(T^[
P)M2>I;%2T^;7RC5"@=+69^OF_\C]4E8!F-PFF>VOO:34W3FK&*G/(7X# LR@4]SY
P[H8,Q8D*((^")'%*'YY"[]$[[-L JE:]VO-NSX?59QZ_:D@V^FHATP@Q :+MEOFK
PIR1?_Q J._:/%>0"B$1<8J@1I3Y(..9TWQR&I7BEP1FS%P.1Z@&_.]Q6PV6I#U-G
PW31A\>*U35S]U[)MPP;K0>%H7@Y$R*#MSS@N;3L*2X=B8C(]7=6E%(;?G1Y=G@PZ
PV\/;03@O[(6VGU0.;(W<TWV<#K)6\<BHB@W.0%/TPA"S7<@P?Z?*FU0F]1RUE$!?
P\*.*NZYLAQ6DB'2S"^C0P/-YS_PAT"LN<T[I)W>R6Y6@> ( 2'WA_H^6M!% Q;5J
PSR3.+&E#3V.,*.X:8!)Z.CP$U#2PM\"!IFET?F]C2$RLL[S 3R'3@6<X^.W,5H:R
P1?K4GGS(![N$V5E+CF#T[),>Z)5\C84RYJ4&[#'JM]O RWJ&&2^G8WQ1)S4JT4J-
PA)8*ZNR@"GTY_<CI5K5OFJR:LR)ZP*O\#]<%OK?37\<+;-N&=@#4]I(L>(<DJ\))
P@V'_MV:5FD=;4(\ ^YB2,!AT($Y)'$ZJ"F0;5K9029,-K6%A035$:F$IM=+V(IJE
P_A63%]8_Y^HSIZK3JW I-;@Q[* <4^S#\TZ/K1\K%\.^<O4*ZF=TA".T:-!LLSM6
PKE6.'5C@]J+MAZ_!R$=QG37(\9E^"$-SGQ\PZ\UI)[.BG#:MV),8*$2[(5W56388
P!RCD%*7L[)XP%1?8Z?0^.2)V0 N^)X.' [EMVY2M+68BE"PAP 6S_E+"J$G/U@4?
PM,R*299O(WL-0+P<S+K.1Q4FL0K_\].EEN;3!UJ7;\^)/QY3[:J"[]HOV11&V9US
P *>57.GAS$349U8[]S&DUD@:(3&3"AE%"V4H:A!Z<L&;GP/]#B@:IBX_Q?.@VS-X
P$QQ;O@)M30'K4D!?RV\@N\/%LG436_;/8FC'4Q/U2+8:\VPS*$M28_;C)Z=;05\<
P'QTO19 )_TI6J/'KP5<<%B+6RIO(*L B9R?GHHX\7)9N6NCFF8[/W3W5T; BVY8=
P#",L<R"^Y177_D>8'*;ER(KVF\Q'A%)B&[5EHL)UE?<+7^B(R?9)I.?H\=G9P?8A
PBO3#A K#B=H<\";D(1 SB7;U23(+:W<C4S/9X6Z#.C]HVV!?APO5+<[X'S'F[0]8
P;>2)0@;LR4@%6%0JCKN8J..C2H#6<L*&9=$H3 -&7QNIR\,#7DZKM6]1N\].%Y[#
P\H#?^;C+8_46V@UIZ2=^(L)R,:GI*6RUE%;.BI?B$G4SA!+?G<[GJF<=:LY>O 5 
P!9RP"7&I]7F:*&22N[%T?7#S?4LEK\BRSA4T>:'CPO%[,7XU$=?B[PDRH;"FEB*>
PT\Y>$=WJ .Q+AKW<C-N2%Z@_60KBZLH#\X&!]OO)@.\;K&P?<)%F*4+""=Y(:2(5
P22_!GP$%O!<?3UU\1"7;H0$=H0>F&#S59*)^=K7XM'H#) 83'&_##0H\*B@AM^KL
P+K[5*6GA>YZ*NH>W6)PL,7*@;(X4B%(X"DI\K-W$%\-J=H+-S,5E Q0DZ/9?!:Y:
P(Z/.!2!(@UPI+1) EV1%%,&?S-;8&EMIZ6[[QR8%A*\*)9HEJ9&*Z^N'EAH<TN5!
P+T%Q^^ 9K=R9.30_.>X@DXR0=BY7%%E[J,T!.+K%LN4S7AQ,7[</;8>.;MW_P,_'
PD=?Y5/FH5AZ&P\?^0Q)JU<!#A=6>]_G-E&G%?,QDA80Y1E?R)[X<X_AO#OQZWONO
PK5S0@AOMA1$>21[W(-](2$([U?19B?6^Z0^%;R^-0 2A#5L#06:HA-H&Z8"2LI7"
P([R;K,Z+X<CCK'NVV Q-A9/68(QJ:82:)6]PR5!5E\YQQN,Z(_9W(BJ (D#^&^K;
PIAP3X@TXABL)LE*GR]B<-'$>M?K]^ (PO0G3.!P>Z //5\&FX_Z^SIU+K=DNT+G-
PK_'_/UDZT#(-$Z=+K\JKA -.4&5IZW8& M$V_!"G%U+.0:NG>5SR@6,<M)/F0 RX
P&;DK9E$#UA+ZKQU.%!&K"<6FU_#Z5A'<O>;$<A$3IOJSL!52FJ.C 0. S )5]0=Z
PH(6Q0WM?'.2](JM<Z$K]9#.)$O)3+GOKOD?OD#>4%:2!%'"B-2-^B.BN=XG\7'XJ
PB#,GHOH'!_BBKLQG7X</)XLL8A $G6LE1(($AV$%TJY!-H?AGJ4H791DSCI.4KF-
P]--NFE'8$1B$I:[* B-M]<-8\(L))RVA1+7#L+OXW<M"5\"]\*/__XBZ)2ZO%'IA
P.'J#]T8 -C+('S4<:]1*5WGZ$ 2-'*D>+26AO%%^G(?,69X9N*!S]MQS5J-TV.Q<
P<M;A%$.FFF(/2/GJ_!-O!LMB!4@**D^UZTI,\26<))5ZTZ[\F/(V4DE4-Z9 'O]1
P0O400OB6\98'8N93MNU\90WUP'F.FVH2W#]I YF!P^P-#HWDH//"*Q%U^$S$VXCE
PB<Y M7C*KVL3W9T.SPEBM96/9#@^%(0,@,4\B""E]>\*56SO"=)]A6IT#N>PW<)H
PKO[B0FQM&=6I9%P=5[GJ&3J-C;?%:6]PP*N8[M^ (7^HV39]F6Z9&^X#"1<9^(D7
PL6"@2$*1GA4-;S[X6EH,Z !)[/LL,R=5<9\4_L'\92$@+(=GI-\><MO5B^9)[4S,
P@.=1&B3PS]3PX70%4WJ"7*4IA"@$1]BH; \WUYJ0>G([?V1#!"PLG9[V>ML5IFV:
PAR7Y21)H:!P$^UCAP"FK2O"R]00:9&05K%7I;U8X.N(12<%E>9$"JDM%H*7&5&BG
PK!:0>HEU7D83L4./Q_TT:IZL]=X)S,>VFV.9:+XX$=<TN_585X!):+J5ZH["W <-
P->K65E,NPM6]2,Y>A7SJD\'UM6P_A1\1.SL<R>\IM$887V<%Y5OEJH.JO,5C9WZ@
P2O(?<!_#CR070;MZ8[2<PFH0-2/,N>.HYOB]W>Z'$_K1*H> ^9.N_0/B3E9J8Z2&
PL397L9?:G2]YMJK!K71F HK4#S+E7X5+85@I:IE>*YLV,U,LF,L4^^$Z]@Q)MSHT
P&+C3O_UB>61KUC <(Y^M^I S.QA(&IW\%6KXYQ$F+2L4)]QX4\RUCM"Z6Y1Y2;H 
P9CR QO,T5?1]636- 8S2_R2TYO89.OVA@H=7>^)IA6D[E;X+<NR+NC(6+G7'D2%N
PBS1)^Z=?*O5)_A!]=*IOK=+[CYYG;MD2JKT-P1LD;(IA$!&'+"W)&*NR-&[07K !
P.EZO@"?9IDY@"/Y[YNZ7QXF3_2;>TZ<5 W8[4+->>4HFIM$P*FH*AEI$BG. T./-
PP@FQ=RB[0LB]2F=7)/#$W\_5 #GRS<[Q2S3&=AL9<]Q3Z R3-SFYX&&-0"2REV9/
P\V$F![_26,]3PH!=#=QC1-9[?K0^T__\QQW<PKF;3"E_MI>RDP(^N;AA^(G'0S2-
PDBC>#%]-G311!C_XT_UY +M48D0<QSY-40G5RDMKR.:S7R)\Z6Z$)'8D6DQ*="!P
P'BL=V1LAI<-0\W9D9>;+02(V38L7"D%,&SRZ!Z42Y_)?G[?QE;9:;<=+'%K[%F[$
P* @"%9+7+(+DI.1CP>WTG"7R.*2660GQXC<#*YB78C1-??!OQ[_(NP]%V[+J Q">
PC\;-]P7'\[EI$9E-I!_R)1%$A)%ASS[)VZR)&PC:JB@094"IM5ML5C:D_A&N#Q'!
P]FHVPVK:1L)W"KKH5S23)" \U61N2-F+B;_<X726I>?G'3\8YQ1.>J,U5'72!,VY
P)X^CF>;UCY=Q:&9A:7X"]Z4.H>#Y'EU ]PK*EYMN6; <>'&6_RIP^.+K*2O7BJOL
P'WQ-)1LM8WQ?,I_)+G!C^.7 E3$Z&3K.Z+TMZ@E<D!<\0!6+==]A@'+IRE9M).\]
P$TN?$[[6Q2<=1U2^ Z]!99\,::B_SZK )2UH;=BU5&I4,XW<7MDC@:(1F*.N'XCM
P-JK.KR9]LR=%0WYH$K#?V%;?T516 @:?E",ISV@Q[]\!&77=^3%0Z\,SD/I%)?7A
P;("%U%.V<IL78?A?W.N$R%4,L.F[EI"&TQ$H KP-RE;@7]XI)M$4^YA2E2BE@H2T
P4$7[NX-YRA+D0FMPN.H/8/Q*C8@F;JP6Z9*_P0ND(G)8*UVEICP2Y^I)S\+8/.KY
P-@#B"__T>J"+COX<FM4<1.QR%0YZ[#F'_7H!X<2*.24;6:FL5@&#3#@E<%W RBI)
PJM86M]6*J_0G:^D:W=$):Z&U8#,5.J2$<PD@KP!*A3FHC?$BFMA\:@A#.+ZF22T 
P$R[U!7RQ%!7+UP_:2D-W<?K$JB,),62Z/-DWX:CDA!O:G20[,,ZF'SQM3HY1%6X1
PU:=SP@M8*;Z/Q+^9!\&HW];.FAY&:V.=]1U<_ * F[Q0A1U1$C=70'G-'+&#_B H
PN@D*9W(3GG;S*24^)L3:&B*%:_L9Y^1(6#;.5_<UBYDE":<@P![/U:6 N@=>BH]:
P'6@"Q:@ V++7N1#46A263Y=57(1)O#OTN:V!!8,0PX8@M=G-*]->CZD+T%TD=C4'
PQ8H6;^'E-Q'Z^/ULI6#;KR_^N6JY7%TQ\\F<NPF#&UN$ 612;K"Y[2".. UF$YB>
P^_YF3@H XY&\?_B?\()!1*VT>0WB\,DB2KF!IKNB/4=$7&L]?# 9/AP^;'7GSQ3,
PY"CR56G_7'_P,KS)[0$<RHKDXO:-.Y2"K%SD![T,$<+[.B'*>KC<)DA#G+ EB9UP
PM5+B $VW/>NK1\*$E3J$(GVKHH)N9(>/?F ::G1B<NHI7H#"UIX:"[\9F>&V)HB,
P])L?.A;:A&[HWZ_32'6M*J=WPKPY%A(7@"R="1T?28-"LO; H7VF,K>#J6+BZ!-A
PQ1+LH.-%Z&?6/.\M_J'D54OD(V>UXD:!A<=\C22&HU*Z$<DHNE'+[\4<.+C[I=+I
P/P;X'?M$L8>M0FMU&DC=BDO]-3Z;&($6Q"4-J-7T=QJT 2\'7] [FI&K/P]_=\(1
PVA H_D>P"M \ !@QMH2O"5%H9R>T&:OS&R>&"?$0 =6;#1"QM'HPO<03(]'9:IMS
P;UY8R:!YX_<:Z+4^5X1K%&$=%=A#F'S9NI;BUWOK:QO#@)8/B[GKH;A8R:D9VD!/
PVX\CR;8=*7$\PY15M 4)W:I3WQW;$9$UF>LTXQA2^@QT8RB9 31Q5I9!6PS:W?<3
PXQ9VEY#C97N';,M"TFX:HH]ET JQR,05_>%X>T1KA<:C)B,1&>!K$/9V3_-.@VH1
P^EBWX[,B:EYVK_54-1NUG/IWW7_/+L>@$FRO2_ZJ$K8X'4QHC]GPM]#[]=/&D$KC
PQER_LML-/#24SJ_ WZW(2UT0+)<Z+B86-^<8U+;"]11DIV(S$D8$<W7[LM6%P$QO
P[ZG:O @/R;@3I68:4RV,*[84- B>3(-*8-J7P:J"W BYH\EQR,; :7ZDR1$$G3%-
P0DO;XT.1JOMW>-5$*%[7#(6#KX+K4/K"2JQ_W3TGK@W,#O=>AE?+YN5QK4ZK-4'Q
PT#UFNB29-_!"6Y!M?ZXLF"L@!?"37[&@$VIG'1BH& <_&D*/[^J*E!*]/@1Q2<G7
P03[QU28,.8UANL*4/"153@Y#(?\>P1QB6&;7TIJAV!>UZQO+(O"+J"2\7#)B,OUT
P"(Y3HUT2IEH8-T'90L+,:)IYK7XP4S#FM-:,:>HK)CT9"[=(YOE3C\@VU8]Y)O=W
PS3_EJ0YJ=8FX[4#/AU"I_Z*? _+=G^WOS*9DH[_5>F1MCLG028!YK@UR\<^56DWM
P%I*XF(\S"CY0G/24!K^:;.6Y[T)_*X[KD^83<.&$S>-%OG9=_QRU@\QP.!Z"@]F;
P7.:Q-4>HB&&'V;4L4VT_)_MW,K9V$(-#:*ZILCO=WP_-'_0=?E Y\G 2S$C+P[DN
PS8CCY-2W+FZ]T-7FP;C^6US_)_)7FVO& 8X#Q1_VVC^F4VX_.I*Z!A88V$2DAB[R
PON)K*/ V- Y3X^\MU<$ 6 ^KUK[+*!9\7IASC5R9,U_LY'3 "^:4.[DQ@$UQF=L_
PJ0Z<"+3-E"] MX#TS+I@+#JV]81OJ^QQO[2)EW+X)43B3KWCPYNZS/X$P6Y9'Y(I
PR\FS!XW5B)3QGM%.5"?CI*_A>#5E?VV:$3E&G&(KQ;GYHQPOW0-C9];*MZN,MFVY
P/M688.ZYJZ8"O+<)5!U=BIGV2>8?CWZ_8#FW=J918'0ZY7YJ7H=MB[#02V_VW!&:
P.O;.0D5]I)N%NIPJ&&Y6-[/P M.(&4B?$-^7N1]#ST[=5W0MR%/L,LQWB[DDDW]^
P>\%-_,E$7INF,:)YH%WIGG"7ZG$C9H-+9\.$_+,;-^M/AJ:Z)8%XAA84##? >SP 
P;^5JO^T[*,<$ R$"2@JV8UAZ0#8!=/SZCY-'IX^X=I50YN85 SLP/O/"WSO9X3ET
P/"[CKKL!J,%MN?&DKQ]@?^S!"<<B%6]MOU4V(A55-QGO=3WN+4\(L1/NLZ3!KTJ(
P!9JAR:"'78$MJ]DA<TDQ*\BE4AI8 ^E_C+LR8AW[!/$.#30#HJU!(;3T/@*2:Y$&
P0?WV51#[ /*S.6>F_/"K<'$!BS=1!C7C4G%:*[UHU DZA?GQ89,-3O9%E?=K1$E6
P KB,<:[@[\PLL$F45L2_*A)D_?)-$SOGZ%!:$AH1\S>01B8!AP8#]\+]2S%,!%0-
PZ"L48995 ZU3;&K@[[>"1EG4FRN7"RK%S&U_L86'\P_E(I /<86@=*XXY#QLK*<J
P6$ARM6X480W9MI#0!31?_QF;BY&;V74(\X_'$*W$(<T-ST[--=$>%!;.9< HK2$:
PIUUO_'=C0@PY"\1K$3RH8O3M!\#J,AOP%#/>M5MF4QRM0-\J<4&0FWFR_*WP[Q1_
PAVC7D-L+FNEX#670_7J.0@,D-/N:%]H6:GG,URG1N]7G54QWN_X@6X6@U<4*>VB,
PWJ5-S,+7%MW[MG@$71]DLF?+8CF52S=KN@8!H/L<8C,TF=Y,(*YL_IR1".OT6AWD
P]BT@"E'QSNB1J#E(+@7=1.V ((3XZ;KS:@Y$^.+XZB$0&&% U?<EXG13WB.Y *NH
PQ$L.%*<\X,SIP%E;6!ALC/>6?*OUI/-.] JC 4P@C]V4 +S)W 69GL :T54[N"\J
P.,JV;M&LH2YL^8B([!20*]J'^?O0X7R'<M^D^V97*%Y+E8.X)('V[G:C?5S\\YFJ
PC*+G3*/NNM-W_^A'YK1])L" 3)MV$9>_ILT\I>KFH8NZ7!,% * Q:GK0M^\>H8!'
PWJ"H+F#%]4KOQ%A0PS)%71UY4V,0M4MWQ_+/8TRY3*?^ :3L5Q[9:['>\#-(G7:8
P;N>8\!UXIQ< >P7EN\:7WASN0E_!IJ"%*CF[[ZSCE&#Y2ER:<5WX7T\J3?]J1*^6
PXP4U3M7Y$8"K7O^<, KJ(RK+/ 8@HIY+?YE#/EGKF6-$I6?3@!2/)[UV:I#;Z3&&
PTD$."YROD9^C WNX%]7-V[#.<!RH@:3ZUP W-#T*K4@W!UOM0]N'$R*3U]T*I2R:
PJZ\R?R4>;]=&-3[,_X *)=X[V>8<I8[H4GTXI_0Q(&L@R![2+3YD<ANC@-78E;01
P;^+:63]1SHH .S KA/^1=Y=+D [H*CK18B1@J$J#Q;K9^L@T4VU0;D@TI\W?+Z4R
P4G1<8D]7\-W7./-#+FB6J207];E]@Q6=A(EJ6)7)RJQ8.$"Z>/&IP!2]>:RF]920
P[@\AW6/84JD%'K&[X1+8T<'4V3<R.&F?J#,OGN?2)K4<8(U9<7N_EQM_Q@:8E@>2
P:L <5^PEUI9/FXI)XD59^G+P);A*<*GE6@:$>I?<==5)G:]7//%^$3_GR'$.'UV9
PM0 VJJI-X\$D8?TPSKV_*/UA"T&R^@N^LFMJ]OG.<=#7O@:^4\' CDJ?;UF8T<V>
P@"#!R\\?D )?:^J5)\8$MQM^FR:XX;I6M D@.J)L"+]28YG-V[#3JZ"@^TZD[^,-
P/^K[EQ#3)^8&I^.(H[1@S#<*B "Z+.5QQPBNJ%QK[S>+G):$=-*FPP?(-[^DYOI-
P*)#O_;HJ\ZR%:^/9N=<X6&L<"=.V"MHI?\&A6%9Y<^3VO(R>=:6.Z&AG\JO&C)1#
PJCF5!9$>J#1)XDZ4E"?WC=_H=!/0.POBY=@ .Y"S>OKKP=&"]/H6IAI5I\D)?/0C
P74S_P]2MD]CU G01'W*.MW$9-'N2.WM1&-RY.$/'DL,W2V6#R40-80/+#01D$>&N
P76JOG Z9K"_VE5<S=;J0%HEJ3)J%3.$9_BZ=OM+ZL^GGJ=4\0G9XU)&E%3EM\93J
P-?&O)<'.^)^W9<L\/0> 6<<?FBVL#U!6@*/F;1NSVO.P<3%[9&[I!?<K]C<<9M2%
P&S"#0:(\=XA#/-%M\:E?M+GSU^!:_M)FKCX)SS<,]"U34+?L-A6%J=%(<2,ZJ.;_
P6I1F")O!B]=Z_N3A7'IT;L'N"XLF$'X#23"Y2K"+P'J 3_#7)-4#->B<.!:3"P[Y
PXT^= "5N/?V4('/IS.6F&[_>U=A_0:X<EX$OBH."*T]Z7TAO+,QD'^Z!9&T_Z2IE
P-=NYO/O\%I$[T>Z13A^N?NV#MOH7*HTKRHU@#ED4D@)4,Z!_\P/Q\W]4-WJ'M*BO
P_EI2\ "KJ$IT/E6\'B\PJ3RJPII7)U@SEKPG)#J?LC/*"T)/'AI>:J-,D<!XR\X.
P\L!=*L7J6_E_O@<:JS1^+KX/%3-W4[HC4:)(.T0]M'DXG"N?V>.Y 8, 1XH1N\I6
P0BD#+\L;E*C23S-3_Y0E#B;HR+P__E&@&T#/3GDCK8YTX>9Y#N5+C2BL=J/ 25(N
PG%!U/VC&WXZ))=RG0DC[A+9M3\;'^-#(%CX!6C;U(<(/<QUZ_35!!%[C-TU+OW,B
PG%NZ#,@%9.'43I\&7'VX\IZ+B,[L@)B9+I Z"9X09K- .>\\9^N[D'4>75)W>ZAD
PP!E%$Y4CHCJ-4',N7)W:>V/F:^T7$F6&T)+9?7'T5W$7C)E2XXC^=ZIRGD.4A<IB
P?B00O/ X"K.U;/%G(78[]67>P=TLXO:YQ1KU ?G&&DCV"E@8F8E33C;Q./P=NE>L
P6CM;U3L5#MI!+5Z@WW$V]EN4MY.^_S1A+=I;$Q/;$5S9V*QZ_EP.(64A'K$B"UD>
PZR\WA" 0S?#L0P&R D6_L8=JJFBRYQ^XN3/43NH7!&>2<.Y N:5]AU"Q9$NL9F_*
P<&*81W5R<FVW!5'E%XX_<#/\ZC-%V&O$%NKC_\GPJ'U^1K?1/#T=)VZCG@[?7VH]
P.' G#X'A-8M_M2<ZY6M<Y4O>(TMP&OI  567_7\4AY=>CEYON%ICQ/1\+,@I'>X8
P?4J Z$]*>*1Q$2K5YQ^Q]/;Y85S_DO0GKT5,TK0(O%N,@+"=%H^+7]6K+W^RU_J_
P%)9;6E*U6AA"S@!NRSI1!^IJ.A^YL&28HE7;-L\P);%UH)QFJJ8K&BX$0:\!I>8S
PT0"";#ME49?>!!$SF6D7KPS<#^&C=+"^NPRQ"Y/HC[KZJI_YE,5 0G^(1+&6H?O^
P2.'@]<]RIW](\E[;GPNS.NN2X>.SW4UEZY"ONQ%J0!;(MVRW/NZ#U='B;P$/S^'-
P"7"/.XRTV/G[-9?8WT[77V!Q;F2D$FPOJ2"0J9(C-W^B7@72WZK4I3X/_U*RM[->
P.N%$*'8_*]Z/FK0 R93,0B*W&)46!A&CV7).AWS<:\.M],0+AO?;8=SZY-+%^BD<
P2OO\Q+%;1252$NJ,HH@0%LU')]K(0J3O@ZA_A,H'%!FKO.HG>"_<+PC'(1JU4OTB
P5G>]YT$D-@-=KNOQ;]$#-P, _?T/5T" 8WV7N'3N>M_)3\M-L@#+YW!>I'[,%/K.
PUJ%?4*;]8)+C&79]H26Y&VUDB9L?WGS4V_?;=:>PR$ISWOM.*'C[WP>4P^_386.<
P6Z'':'?PX-R$A7YHE>0.!2TI7!4>*$>APK^2N4#!+=;0@>([3V)V9E'2\@],<YML
PT;_G%,8="3O*H7<ZL6:]M3:K:WU&6[ UUO*=2*\\\8RKX/9DDQW&LF>.9MZ\TT16
PHR!F\D2;3&TOZ!-:Y>XZ5BC/UB_+)_5M*_'1^[\#_F06&#^2A3Q?$\4N@9RP',\C
P,\=2QP*Y=%C/5NF]>(JR@AZY?AUV>(!O.2Q7\@X&[!J/AR$$^_-17W#]*LP?,>DB
P_'L,-],?VS6C&JNXRB-S-9<<GLDTJ&_3K6);L'J205Y&]2>E_"'4164./I.RQ_'Y
P3]Z^,MJ2_T&V?X6Y!Q)<727#533#L%#0I%W!QG<8N"^ 7KK?/8]K%J>3C@Y\+""8
P^U>DQ5?_;.)3X3OX&138Q'\T.L.V*=![QK]<\#"N<7Y%,*6/4O&%@W(3N(BK7GH:
P037?*M/8#0%M6N'2GPN-+R@!-W0!["&%J$MPP/R/PW#^<6K')88?B<T?I8&< +-K
P'ONROH3WUS$S"UO*V=1VE#'0LCO-&4T^J3)>R*B6,K2])87?NZ7P^%G=9-$!S\RW
P.BYQZ"RL&O_RT&0N>;@U)<\J![MXM4=11Q06M^EE\3+6!$ [JK=SY_W\8N-,,7L=
P55I9=EY#/)%--3-J!)!N2O#SK#/RHL=?QQLU4$E3;T)I!DHMCY0H>?UI<!%/]KP,
P6&>]4:X^_P UF:$3<WI1'(:GX.=RI$RT<?(08!=#(Y*X3@+P[RNLI[E"2)B.X$F.
P6ZE. #@5_M'/\;W>Z3JJQMZ=R4V7BQY83HT&CO8[S#\_++2%XHY*OOH/EK'O,F.C
P5=+6,I%33<"GI)/QY&QRQWJ%WF7_AL/\:>:OUZX2Q1>;1D,S3.5FQR%),0=FO"[=
P#"L\.$OK#T7MGTCR;^V43.>A();=7:4>523M3N& 'Z38?PQ7 G]R:ZZ?5T24,$X5
P\C66.&\(7LVVB>#S1709?S0>:F,)6V?O#A9M3D:\=.E.);0]?,,[D>$";AWLBN[;
P7(5N<:1VH..UEGY<#Q)'C8WGXIV*UXE(+,I,UI4 9=*)I)KL2+RQ2LP!WJHG-*:C
PLK!\+% OO7'97AR:2(^[[381_^Z:^/I6'398*#,\ZA&/K9Y!'O2PCO(D>/LTB)*0
PW3TZTSXEULL# LT#_?T&$-<./1["2@;^LV56<K&9U_:&P_)31] !0:JU=*$RPX3@
P?6609.&*R@R6RG*TJ9^9G#Z4!3*J1AEG?DTHN;JT? EDQB:AD7IE0TXF)6[$C5!8
P F/=>S)%%S2O78))42F1#JYC;0N?96^#LP;<'5@T2U6M&(D#BW3H-@='*V=;_JXI
P7L9MX:6YX>U_C['&P!YB123V"\(A038!YFR>E=-B:F;XW23!X(:Q;GNMI!PU"<1^
PSZZ75#BCIS8!^V)B^1-YZ&I[L@W-\[I.H$> RH_S)I_(1+B!""*D ]4.>'3I7,6[
P@!^6#A3_1(2:%!*E377;EF9"QJD.RW2EEA&PF[^C1;P74R)G<*6D?N4E.7IW5.7U
P4V!_7)FB*!H27/$!";1U[4TN@H,R#FG]XS=?LD<OK .)P!P'MI>&L"VVN8F/UK"4
PD3YO^G4?/=U&M^!D5[N:-0+Y.S:0 DE">Z1&ZB)>>'7LWE%:._Q]5RXA$8[+HA_-
P$JT&75OAX-ZR5#?(!K_W.CK7:7/3$<KCW"2/H:X'?5 S#HYM TI?($7D<Z-15?NQ
P[4CEXD_FO:M\"MGT5A@6W.$)ZH'[6)9/O5F!.E=\74<S'[\)(1NUT)$"%Q'N4:):
PJL24HNE6PH!S##G$Y1^VCZUSY\K%&Y8?<4'5 JKE6P$GI(I,?IK:8:IWMTAK<*KJ
P2X(L"GIJSF(3$C)])PG._<3K>+-74/KJ$&1;>EZLZOW=,;VQ?J20\I8. &6[2DA6
P^)Z*R'HZS3OG@Y1*D0)D($A%<RR(.R, U^18AQ$(KE[?%X_N;$D'-$+LG^&=J#0(
P)XD8WBIW54A:V&X ^)U52!56 W5[_,79GYMFIH>YEP%,&:'.S[QO%(Y_&S]V,)+!
PT"18,^\N$"K[5M-1"H$CI)MYI8,(T\0S1][OD5 ,+R#$_)E.33)]9P3JG" K^=V/
P@/DNY?)@(PE\XH_0%G4$=>M(JI=)'.&0ME#@@>H7VW!]0$:@ZDCUE+T^M'HYQ50\
P!HJ_-ZFD-U:K'ZX1.%*!UDX27>HXK+U4HACAWUNGX.(9M1GA4)(/((.[DG9;R(T9
PUWDRE-15]B+ZX8G -/<34U>K%KI34!A-]C!6G(\]$.94<7G^"=\$"E!_N!4M)]KS
P36EIS[$[@U75( OAKTQ=F%J!UN7N:6X5O*YQD0K(9]/1T'R3F0]&DE2'VI(/UK9@
P6J_BPY1'D1':BS5^&,P_A+*;/9IJEG6H>RRD>IWD(UQ3)>(7>7%.X]0F(758=:!2
PAD'1B"F]+K'D)J_&#/B:$UC32$^C</-X8$I30 DE'EE -(E$Q(%?FC/TAEAPQN*"
PZ$LU?14Y$3X:>[)^9+-T]LPZZ1P@ND]BT*(-ZMIOV=A(.X.BUHYS'>Z%2A58PA2B
PT9U6U0Y@TL18Z3MGVS'_OM6%,X9'+8:HS5##?IXD9%M[UW7,W*3\A!DX42K/I:_T
P9I6?!HO /70ZA$0UM?*"L)M:N8D_6^G*;[6>R$0*B,7Z4=*WID:S(N<A<G_K!\)3
PA7M^PF(ULIJ[6XQ=W^!$I#>4%F;G]@$SJR<X^>N";,OF,=XT%Y9EE['' S7A_(EG
P[&ASMV>%PM52?4N>>U6,%4GO60XY 2?-1EX:U#I[*9U1_C'JT7RG!_#3.@YNUF5"
P=$_]<+ S:K BG%=#4QZ'!]IX/,KSH\IP>);]0Q+Z(8'+L-KQ.!1;W&"QNRGNQ,P+
P"&-@>:#V8X$[TC@?,(NI#F-./PZ"C&6 )P6 L@&E=')(9M&%C8(E(Z=;^$:(/MG%
P%"??XMM-JBW/I19ZL[_.;SBPD_!8G)M=Q3\]YDUA1RIML(Q'3@+:9[H&E> OT'KH
PK_!8!:89(HZUR69M3B)$,"BGEEICH%;=V:X#!]OM=JZ)L<*/QK1*T&W_]^8@ETPK
P;)ZU'7%0=G_]6!UH!>I@3[?B1SD@)5(23CR3.QS,O>GH!F)TK)*WTK$I(J>YW4ST
PMT:JN>AE<-,>/C6@V$5<@W8K&/P(IU'4RX'LP;G2_I -MX#*(.-.H(W03Z=EX:I[
PY;F#16-G8IUJ9SF, -!/ER,@/L\$:+O/,&5IUOB$>QQ1<@V87:'E/ $)2Q/XM#48
PMBLMG/;7K2#A0A /P*E.VW'O'U@+QU:+&63P 03](8)BX3 R:SG,$MLX0B_$B$ZQ
P9?+G3$H6S1?EO?I0$;4OTY55GKW$VB@(">Z9S_K',ZH6G$78O6QM-,* *>/2<U*-
P)0/4*NDE=Y!D4]U&G9BR1HMC$>,]JK;"\]@2$[<BIU:B%T9-@^R*K-5(*\N)>%+$
PV'%\,K18<6R*?CDL8N,5@2W)/=V3#,@I%N!B6+'V[E>&GC!. 6[A=3A?G5;F@X>^
PUNX0OAOUOS_&&=<@Z^VQ0GYUZJN+3U"M0V\4A4SK8;*NSC"V!5?Q-G82+\5JD]LA
P!ACDKEJG9#*3N7$C9 ,2#)L5[]SUVEMUKIJ-0VJ6=._7*5K+CQ[#[VH>CG.5<7J'
P=PLRU,U&TVC?!]CF([K#FKMTK'59!C09&5.NA, ^B/VV,0A/36JV9CI2B5=&,D<&
P9 ',6B.,YO:R/87=*% /L1'Z'C_,)52.E46QN#DX3_D8>H8^DSR;?I4PSAR;7AM"
PO6'OKS?N12SJN.;0R50!DA-P?'8+@8SJ?5.0,9"DI.*39L1TO$_JG]J%+AIKLI(U
P,63&!>AJAQM$A2308F_S.6;*.,7-#;&/MWJG$>D0HLIG^K@R-7)!MTE3X$]WF_74
P/%MZ,-$'Q;3C(B7TG-9&3NJ[514P*9:Y4$[(VQG9H<YU>6)S+*^R?XQEC1@E6K?7
PF<\34^I;X.$<8YV(+A2!-C,8"5_RZZ#9GGK+C!R>ZN3T^\Z:_V@Z2Q)EH&VS\"/E
PX%61:=OV;?6(DBJ=_)W#_,FQ_7!@CI#WJ+W4H\O 5)P5!U,P%Y7J4KVOOEK8BHA(
PN*$'<5DA8B(F]<WGR[*8"CNU1KV"9DPC>9QC2L][?M-X]W4 Z9*#XA(^)O1=QNHF
PHDUO2@U<Z5,O3WMG6GUZ7U(1I]^P*2-5.=M,[=$EO%;-@S_Z#P/3VYUAMX0+&S $
PP!<I?X6;BBFL84.R2Q;;&/O;/7=N0:;YE5-,B9+ABE>(:O%&&IJ8.X&\RFH*\>?A
P52\RX/ISB0S 5!YTI\=17TK.3J2MFB.D.A9 JRV^)'6H-I+P?-254(XZ2?"KMN<]
P:K87.5=>AB.Z7J([*+%J^*!*S%<6$#K 5*(+.E9L8LMD,NO+D/( [X$,D$:PML K
PLF- .\!83'5!F<#[ 2Q4S#%8>5G2B!"GU,(OS/<P^O4B8 <5-# 5"_.=1)F&OI<&
P&UM++_=BY?3)HLC+):H!CR<6\:['A,:LXOPOR\.]=G/PPA4N^%5$@.N/G\\;*Y8-
PD#VK+)#?[#YE_S\_\)-X_Y2:LR\QP=:S;=5O&T@L-P<8SG 2OJ)?&A9.SX,G5Q1>
PN=,J>71SAC19!+#2D2^F(@N'^.,^_(P4MG=CEF$%\A\RXN.MDB.;8M[QL/)&!9?/
P;->NR6#[K53SX+RGYE<I9/+G-^:!F/Q;_D%'*^<EAJV#,,_[S:&566H1(L>D1(; 
PY( SC:!S;8P<@(WVM<2'#+OQNL"90V1>82Y3N*3OW#IF'(E]9_R4_,.>6$(P=C";
PWD3:F&<F <<$P\U\W5+FZC_UV4C^D.T>9JOPHI88_#.:!3W?Z4,5.4?5K51IDDP8
P2/FPZ(I*8.NXA'D9W2H +GX7K,\)N-H._Q/VH\%:E(6:O1D[2-NOLWR]QD]G[-3[
P5<-TD*YR-F.\P"+/$*,GX.1SNG6)^D^R$S>>.,[1 ,C:^XD!!TQJVA'><&/[WW[M
P8/$!_P0K60E7L$J95:R986K&B</14I_@*VQ*M<3*H8,MXR*G?++_%4MEBSZF4$A<
P=IF^'7S%<7-6Z?XUVU#2?]HSDL9R]"[N.A35R:Z[?87L27-M=CMKIW0NK9(JN?$Q
PA%FY26;!:0=6['1:Q-ACFEIS5[DNPWR '$WU+C(4M;EN/:+OV5VZ6TW\K&M 5Y6U
PW.K(QOQ6_]XAQZ]-CG@4UT]0(N!H5_X40JG\W1R9B[C%L82WM*EO2_O?5N$+6%\5
P[IO-_%EE^M[?F467O@6L) '(2C%2\*IH(QMI\!C)T[P,E^-HU46>)QK(:GV&AAEG
P9NE&ANF4L3JB\.TGK5TX\Y^6#RXDS;ZV!_*T[DY +68/T"NZ/[> "-4^ITEKNBJ'
P>R9 .MQEEV #@XG%55W5ND8*G5J: ^DK#6]&MK^S\#>WTB?JP:-' 1Y+PYPO4I_%
P PRK $O"\^:DOTN,EBYR.[#CU)!K?_*)?2T0U</<X9E&K8T%ZW*M8IS<!,YOX)<5
P2O?X-!5(=.49+4%M.K#R5SKF5!LG!WD/(2?^RT4%I4$-;8^*A,,.]8?AMX)I72/D
P5?M1+:V+N.\0DV==Q="&T;%L% P8YA4 H)):"AEIB%>.?&[Y<=_AC->R2]^;V5*<
PI.SH1CV#RCTS+N_O(M6$!TD%FJ\C07Y^#>9F799)4&IGPX^H7.B#_@?1_*BLUG(5
PD$.85,JW,G7,KEL<W8OZV<<^)8R30B4(#N3FN8LL!:+%BNX&EW=OIR+6F3S%!PU@
P^2,E-=-*?.FCH%PE4+"B!H?3-#S%\QOE<$8H9]J "?S\4<P(_P>.V,F>>@<9AM S
PJ<I+#D)F5")C]QL"ZUTE"W$?"\C\[DA CE'RPAGM9BK^-4?#QIS=Q4B3LBBH0")8
P>VLF3NRA,Z9&2XO-K"M<Z!W#HA2+BO"\WR8OF?] ,OBR@J5P?6EFIOP: ^;"IB6/
P T-Y@(*Y_?UET+*PA4,M/2?=3\8BGU3/V@X_;O%_>:_H2 ]:5 @5$<EC:,:4 U?.
P\BI<-345:2T,V.[#WF1P/O^73F=:C^CA :Y !!/A?"%/81O$=\TC*IVD2E1+X$VW
P@0MV_NB>@5<$@)T+8"A-DQJ4_[F8P2#D-^N*3S4=&/FA< >=/FUX,AQ7>4'TC/BX
P"C=<XUQ!DN_S+-Q3N(C>*@@=1V,H!')NZ,TR'9;7T!ST$RMZVY1A2TS3I26[6GWI
P9J/13T]_66OXC? )(L>[Y],[1&G]O164$U<@/_ ^9=.VCH428W-9YN[ENX3C.=TF
P!,K&8^4<<ELWU0([X6(F.8_VJ"(L9KG:;8JY1<9DG, H<KZM5%Q?^,#L",?=R2<?
P?<RF5/26W1"2S6]L)VL#*;O/[2E:=8C:V> \7P^-'5B_!2O[EXK:P&!OM@F@#65D
PXV.Y$WOJK1/VR^]8@$A[9@947G5G6SNDY%^!J::/QV-S&U>FQ]"$IJ)QKF^!.>D1
P.S?*H^[#9:>0YP[XZ/S: >,>LS2OB;5D:Y\:HC)QMQOGSX[WB5)VP]O^+" 3N)JP
P>YJ$W-5EJDMY*:@-R%WAI6=SS&,%(;<U,)JN>2[!8?309##CZ,7DP9KQN9<<: M]
PZ" J#%#Q#EH#\QWC6>SZ!K_837IY5TJ6MQXCX)W%XXJB8.^]?G_K4O!TU /X0YHK
PZ$WU'!YF5)S,3):[CO3)Q RLQOMV]0HP-K@/LG^OF]]-NU0;?"7T' (LE/',I)1K
PD=I%N 7L=)JKM+OKP']IP,D\*=(/9JWKJ6"G=#_+$"31DK6AR0*G;E$A3F%?[_),
PUO$'FU#:CKYKR^?#FM7U;D_3_XX]:ZI\EGANA*Y1BM9T<KN_$R;#KBJJ432O*SHS
PPG7L:7P\B $LZN9KA"!B]=?KT8[NPR'44 @;*9T93 OTZ8HX"OH^QU%*/Y;@U<L$
PD91^/-85"A[[3TZTBUG<JJ-DH[P5:FE.H=N5Z! 'ZN.ZMP1992B%72 "CM?O)YB#
PBEAIX2;5?  &K;!):SO3_DHU<T_=X"ZG]=-^=O.EO"F84KGQ>51M^R_!^[9O.81N
P21R,]V"9CU-+>'LK"[, Z"FC;FNV*4,&X9=L'TB[.1VI9:(YQ5/ER@ "AM[H=]40
P]H)"L./_P(6NE>KY=0Y4F1P_6:MG#L,(+?:I1E,F$^HAY&7#I9/R0>06QR]7]C97
P?2+:!PT*%L8B&FRWY:EEI\2CX3ZZN8JBC!P_$(A#<.0&J7"+HV#?15Y7^YQ)TM0O
P>R8,JS.[+XDD=? JW:NL\  P]E5$SE1C+1@[DJ1B*8ZMJV^;$,#8:B,0-?9T!_(,
PIHU;9_TCJ<==PYIE'"-#F&2DQG09\-)C)&9[)N%H\P:P/W4_>TDWN4WP\@,X!WP"
P6:NB<R@L(:0\*@6O"(;XU1I(J^Q#7 ./9U]L1<<6WOV"P3!3+E%=[]Q\; S(ORD-
P-UD=#"@MT6RF1H0T?2X0$8D]+\"F"I#B3?'.E*52""2=H^SQY'KT2Q,-3^4 %Z,M
P/:+;"-_=EQ[\SUC"!FWR9>+:Y@!<_J>0^:6$MOMJS,BJ<#M^43M=)HI:HO.OGS@3
P"5XK-07X5XLO"Q_!; "R]8/AV7FH8FFM6/A]>9.8?K;.,GEDY!U:<<'>__^F&%WE
PBEI-<"5H!P-$)0WDY1]"K\1P[V;"L\6!@F?G-3GBGW2)"6=PFY<)I]Y?$*Y!![@@
PCW!_.%!/ARSI132_NB(#365?*IA;2YRC:^5C?@;:CI6#]29PO(0\9;[0MLT>:MCN
P(>GX0?-.D]!\!1 <WYDP@;=%5!I6\GDW>[M7U*F6QY>&4DE9Z%7_^GTP>$6&!O[9
PJO2C'-85FH>6:48Z(U%6,*2- $(LY2$%]9.R-U#SI%YA.*^F=!?2:N[/X+AS8+AZ
P[7YO+>;3U*(A!<4O!>U%,\U%OW0X&5>&7<P/<+188\*O&]VNA<CX^-6T?*>_:%,@
PQU*QB$KP51L;R?K$MCR7VJSUTM3B9:1ITL^ZE^!N+=-1YI(7>:PIA_)GXS:\7!@/
P1B>V8I;!/1BA@DFL[D.G<2@U 105HI[9%R^Q]F/@&WILM:(/EX7X6*G*7"_3P: Y
PB$"5;9*(6;J%C]AM[=9] "^U]OF$>GV6,$NVG>.$!:W_$LTS"A0&351PRS'>S;5\
PBI96=U/=;84I"S:W9"(D&;4:HA;+*/9PT%%HC+[Q5(8QA[&MM.S_]FAXS(F>W PX
PUT7^]=JQINJJ*2CJ!_1OA*98#[D?B*"\6]_$'7?0F0]5_DCB+,T%9J(*^H>ZV_$B
PMN[V-TV_D'K\YXI'$$>,4Y3:.D==^B>X!4M,_>J_QNKE)3?BEA;P%='(:-V?I^JO
P9YWN"FM.DW]("8+YSCWSKZ]X!2"80;62R$-L?W_'$ WI]B>/2<#-UN^$AT/V(^IJ
P=>C;NG%3U]:)U2/'V3D/-=2\RQ9Y*3^]4C/*(\*X>P DZ;57"#"G!T]V!2#M-DO,
P,$?234,;B Q]OT>+W_\U2*/ KL.164<0:#J@4P:X,"XQ\_.N*#23)7WU60)&ZRD*
P=&V7Q^T26"&FZ,*G"2$OCA,+CAV0+BHT^BFAY$5]CSX<Q$*3UPS5G/D'P9^"/2R!
PA?K-)_F>(%[CZ5P=H8EZEXN.79:M@U.1))CGY=5$I[<)?&1^,GZT?C%3(M3):5?^
PE4PDUQG[-U*DW/2Z8B&S@':#5*PJ?)_.Y^R/U&R"Q32'*=8^>\26K%98<UF2D@\<
PO,0@KTB0.Y3-KF++9E);[[]-#RS'<YAF)OL+6"<.;X=$%9/J*)"4BC*-G \!?-!;
P<DAWQZH_#O- D-L'_N!MZ?GT9%(3 =:YC&]/+M8 0-S0M7DEE,&$5(<[0N @WE*N
PL/3JTYR_BU5!DE10"LCFJ5OR*,]D7@%)C6W6U#(=3T0*FG6CP&X);\5:U9OPE!SC
P;,[I?D+3['>;RP]8N-72<+&K)\6LY!\< FGII$3=](/,H=PQ$WXC8$QJ,X,D6$?[
P6PLFN*/H]].0)U7YU%ME^+LAC40FU=U-9.GR=BC&=:HYN8$5SVA)83K[=S9/S^'T
P<"OS#(%\GN0^ E[G1QPQ[H#NQF+WH:%+A&,MU[9A7&+=$=C1>&7@FX-\]]JOR\6L
P7=N?Y,935VC#LVA!7B8$B^.J3>P_2JB!9^,G4^.O-JUCAXZM3=G .0NX(<[G.:)"
PJ-_4(?ODPE0/"-->KK#';EB()2J"')Z<8\3#R\V;[281M'IL%%Z//06I7U4M$&N0
P;PIX$B-PLB5:"MW=7<,=-:F$ KA=TJ6 $:7S2A#-4B6U./7/;<AG]7WRZ^;5CKY*
P')JK+[ZQXSNO%KBT14.9L3I \.N,Q24TQD^93.+-0<PN3V@-6!^KGL8WD.9CAR/Q
PE'[16 2?+(_'2,C0+Y6P7+V@TRV9'E8O%#>$!.O1GE;K^L=$NX6_W!TXF_!EI,6R
PI8L-B#-\]B5E7%@R";D.JF^U:D^@IQ$"PMSO]&Q7-.1:K;#I74 K(#5/DLWQ\SN:
PD>]LJ=0!1Z+!Y0RF?9ECG""VY%3E^P3ZW[8)*X=Q"_P%4"4+*1V/"DQ]]K& 9[\B
PR$9F/^1V,D[$F3,[4WW^J<UCE4U^;.2B<8R5E3KIR(2LF+)LDA?198=[W$G;=3._
P1(7:VTH)KRP.;'K5 9">D<"#(!X[:<&SQ'@\@O$@/C\JLX@_EAQ#EZR.FKG8I2\;
PLTK\R5^;S]='&BB^1GS:5,2XVN1)!-0H:L82/*Q\'@ YZBA9)3.?<K,R[! B'4$H
PR3TEE2)85X$P1DDD_E#HX!:1^RB[&T#(^%\\26G3&X&S#US7M3/S*$.$3Q-4+/8?
P7I[>!C@?1 ^1=!B:DZI0TU8)8Y["/ BUY?^W*7,B".7KG$%?,WAF1;B C*==W-9*
P0]B!*].V1'V CRV76?&%D^?$Z>+>!/=1A@MD'Q/('(2&HU@X$T[8>F-"[UUN2?$*
PM)]T4<[G?+]9G$V"K,&4Z%163.&PW\.AE2C4RP( 3_4E!.8D+W;'>3N/<I,"5)_O
P'7(<&5[U?SGCI"EN9!+IT&O:9>G[1C2-3#!=(YGG5#!:CU2HH**_NTE59!/Y@>X1
P4"N@J1;M/%"JT9Q\(R6<[EP5BJL\^+B;[%C3.^2..<(A-N#($/1U%3 FJWN1<M&B
PUC'-&^7@3[C"1-^-V#RQ-U]8.O)0C)5.'X!)T!\\R=V/_*P@P'K32?KR!O9R%UJ)
PX%AI?ZASBL-()L0??9T@( UFG4]KI):R&G6;(7'D^H3ALIF=.YV">B-=:,7/#-F_
P#YUIZC8Z^"_#9HMJ7)K>O;1D^)_@&_R?"@8WN#I+QJZ*V\?JQU3T4VMC!M3D/PMS
PT$MKU'C+ZC2'1<YP 85M#2(8[VA=')0H;TV3+Z:E*A2W0M<TGI6!:7$N2_09QQ$0
PZUI&J34JZO>9>_5XU%7:PV,W&>C\STM-@K!^L8'2IV8OI*R_65T!>Y??D<"V'8@V
P<$7D=X#7)4N&X78F5A'  <"+*_'8]E(UG96X]=">01V?[Y<\WR@_6U\:Q9H;5_E;
P3AK8U8V[GN4P7VP/R7')3^U9-A'&B0E$\JQ$TTQ&H_U#6R#>+*G/YDE$7A-43/;Q
PZCQ^6>] L%U^'#X\^52#&/D&8=U:7Z/%B<2C[8Z@ .I@?*VD5'FLIWDZ'YN(U^$P
P"'<,DB!Q"2&C3Q Z.LT0'ZL=Y4VBM+_=)PKYM.O:8\"$C4)%55!WRH'7G"2>]GL.
PP.MC.AW">3N8;$=3HK_KAU8D;[B?'*0.(IT0JVX.BO6 >*I2]TQX#M7M5%CP:3O@
PA*">7,**1?%HY5H.8E[6\YTHSV[J[,"2P;IV/$AU=X^&4CCK.)2DF;W]DFLG^L<W
P:PT?Y>DV-/!:]1>-? <^( \]9I'*48E8_N6N$WO'_QX=TQVK!KXS='.<YCR0?Q63
P9DCZ#[H'^&"+&BO,S:2I#E+B+WJBN73G[PL=$(L-E&4>LRUIR3>>5.; M*X52'8^
P>K+==S%A+#46O'GJR_WB^JJ"L2CZ0>*?(;FE!]XB5K$/ELHCPB4-3'A7I)XCY50=
P!9:B3"*%HA4?HK)GMEA/MX\YWFY<ZCDIJMS(/0;<NO@[ F/>TZIP(R/FU.YF-DHW
POG*YJ87AGI#;7!*8L#G>-E-92?N,5L_;%A9.K4SIM" &GFH,E5$[+-(J;:W#1EH^
PHJ1UJ.+%SY+W(YH=6TMI/Y=E+U3??D+C;&C49;9_*9)@&[D%2N%!#:.)B-TZOH(H
PR+2LJ%G(.9HEM3DGMZ;ZZ-/<RKO3$=+^57LANT<+73H7@I<3',N<NZBH$9AD&*^0
P<=V(=FF[]  -9^>;J;#D+XW(D:57H/2A> 7\D$+C.2H)FB7RA;J16+I <G+[ K(M
P<1?H[F;SE(#5:S7T8FK03. C7C\F=J6%+.4 #[$TK-.EEKX\&S:Z >Z)NO;E6/WD
P4?V>O .HJS*A\]I"F3 .H+#4]EG]-3[?"WT9V-.]_)/;G&;G'6O._#/F1FD>L>V.
P<_<L7UI$&#"C6'I%UOT?*HQ)+LHVH5*"L(0)%*=>WXL]$$ED"@AO /#GZ79;4SS7
P_G/E=K.K^#GTCY^D<2WZ0?]/'Z5; 9[@-I14X__!UK<?#<5UQ\>X?3FY,;6B,\N 
P0>,>.N[S[.V54+16_YN!_67VQ5HXELUZ[;AQSF)Z/<!<OI<&:.7J'2,2[\%C!](S
PSX;D,E%)A/*)XAQ>KS"0-Y0O>2O0FH;/?0[FADL\4@?-*64%;T,V:/3+>SI22X@%
P?A@&X*4T=Q]3J:@EN[ST_\>(>O__\D]:T5AC 1SD%8*IIA.6J5'.PRTU@<0 ,,IG
PS5;09[[]DHS_1!B[?4K*P#[@YF3N.^?X^X_0P1AW#+5]/G"(2AD7_VGX))=+F:%A
PUR'=7$I9Z<\T!'K V;:MU<0'#5WB=UU!(/ES(2MZC1E&+?<YG=G=RLZ<<>F:W9TF
P["$>(V.??YH:)BB,,"5R(?PH([!_Q$I_8J4>,LOW2EUYO^337SS,A=AS_YSN3V$Z
P+\@CO])8LM$9P_L8 D(==0HA$K%;(VP'+QVOJ0[R<[4+"B2KL[<U=1W-;_S(3J_X
P1G'\64X&I=&OJ-2SO?=\BQ2"D>Y?9I>MD2O;33BK]A$VXDN?B&M4JL]8JL[MP  P
PW;35SGM_#=Q+\UE(';O1RX8NS.9HIIP!'5.U:BANH84.$WJ4 ;6_TF1<@ &HLQ 0
PAKXD9%(O<Q0^N^VO:/>@=-8!7>-Y6Q"YON\%:[G39EZM 6[9!_IQ#V*_#Z?\O?:A
PI:D:CV%'?CTD(_.WB,?/5@663:,53^1@Z]&0LWC?XV.:Q^GDR1HF7HFH0 H5RGU8
PM02GE.TB$^$62TK9LO;^QOAL?5/FW<'?X[M"<=+\("F7] W1%=WT* !D/?NSUKC4
P<'(R]TA_/R?+BTQAN,^;#E9GV_A%?G6M* S\S$V!9"S7FQ+:ZNWTV\1*>WT:=&[1
P^/RCTZ-U[L5$I\T$^*V#BDP^\-H /X=HLEOL5F!)O#"YNA->@R7.>1 $9P;RY,D_
P@])T6+\*FS'U$D>7?M0ET.*58N1G1^4<_A6&*-G/8V2QE[YY3I09J<Y-Y:^X:#N&
PU H@WH<:SJ8^L,*>;96Q^&Q!RM-^0*6]RM%B/>2J:+?N?(O"PJA9BS/GIW%R.R3J
PQ06EZ,J5KMB<.Y^I[:P_"OI#,E'K .@"EDI@#R;<J6^7Z#86WB66J&Q+Q=L7'-[P
PN! T5^N6G!T"]Q* U.&D[_DIQ$\>62R/V)I072F/S1:A^Q-P@^R^WK%W?F+,)E1X
PY;;B;<9O /WMN=F/.#X6]!?JY4$FYZ E\O:=6M$X&\L4>BH$46^EA(NS"EVMYSF-
P%VA0PQ7-/=HTFNK] I(" BYI6W48*E^F.0=X82FL+:&REE"F J2;C1%_@)UCB= D
P=I82<.U0;=!J$\\^U/SMAH$&;'K@J;/C CN:,CI^T+<UZ2TC[I7_KGMV<9V3T*1&
PIW#8RM$Q(P\L,/FG#$>:X#NE0S.,&C<]L0XP['*GV803%5\4XWM,.OY[SVD"9UMK
P<29$5A_>K1 ^D\NE#5N5DOK^LP[MG?P-\NW;A:WN3=\!P\PR<O0Q";(?)E60ZJV%
P@3<_55;71WMS(D.LCW]>)SJ*[]S1RDGZ<WQN+,<+^)W"&PP_4<S$'ZB-?%CL5)H>
P@MBQS$#XU0L;U9 ?7/YV*7Y@Z<+VA?%T]*FE+8^GF(*VJY#;+?5QQ6)!4V@BTU+\
PZCJRVO3_U7ZWU9-OY>:4*NHW&B:0"A'?^O7Q>KH2IK$IUXC%-]?,J1M?CGIS8F'\
PN#A(O"(",<"?TGH<E]Z"Y9#60UORO5-ZPI$8(L&P"A4OLW(<_NE&1%C#P>6*A&V?
P9_AV$SXY.1P9/1%!Q%(^3]?I-X.2!)_Z P';.;+8%0@WN361VU:U_<I:B^Y\)/E;
POG%NLGZ#=&S_B6\E.159/VU>6O%@39&1$$J_,E<1+:+CUDLT,B$TH_B MON%2!0,
PU[RLOU@ MU+?N=FHK6%,]IUK=.Z]8=^+M;XGA/<(/QJ".#VA4TMU#/2#WDFPQ#?Z
PT=ZWJ<X8#-CIY>-GB5M9=;ST4@'['LK9QZ4NZ1B_^ ',%2*6]^BNYS'-W/*>J;'^
PE5PJ@31BFVSNF-65AJN!B<7D[]2%JZ(QZ)FZ8V5[G%NE6S5G]ZB?SD1OAEQ3"J"[
P.="H>&9KGK@('&?ZZ9*O!?AKXF.G0:_)GQ:W8JE(M'BXC(!;BB<'.'][3O!Q+9NR
P,=+X@_]PU10"A;/1%HF\/],AY]DI&11EJ^H*V#?WR>;R!=_9IEZ]@9.B :$5"T2S
PH)!([]KF9SQX! BMN;2MA[S&!&M 6PCC&+0[_)Q,IIHLW<U"5XJ^FB*BF1<7\PV0
PEKWF#Y&U4BII\2R;KDQ"X8O<7C$9JIR&33_PX1NG.9R*Z<3L=7($\&#OF -5CQK/
PB$"F']TE'DB@.JS/W/16]\]A;B)"7N>1$C+&.,T!D)]F!J@Q+(FP^7^,QJ'(="E3
PN&H*KUS2B2]Y>0%U2H>444 \@)!0-[D&_/B.-V?S!<5,G!Y0""Y=?L>0$&U)BOS?
P J.PQ"[+&@&='W]66N"G)7^Z^1'0R>T'"S2EW?,BUG$"I81R51T$T53<)L"#*Z^-
P9?;^>%M<#/PU#N4:RJ*\#U.I$VM4'UM7-=:J3R"_K6Z(EJ?(JUGPZ1.^1? 4*3I_
P 6LRH_SBHJ$ :\)]&&;YR8$ZT?^$[6O]IY5(<7D:!XM<'6-<)UQ_2-"/)JD+DB^U
PU&I_J^KB.(K;CF_A(U9"<LZ)[E'0212OKL: OD*/7K>VBX\%3A8V<>. 8O1B"+=;
P_UT(E=Q_?QU'KWX\^:,Y@DFJ3F#>[ :V\1 +%9$F5]CZ7I_MS-W +4=W;+[N=PD/
P)OB)V"'1G^)6LQ 3LS;M[.TZ19HKBA-*N= TX&R&XSO;"W8J':A&J7)8%NC^HZCN
P56QWO;R[U56//^[?H5HH0_5%CA0'L3T5:(D/N*]S9FI[+6(T= @)F^;D9G$QV.%!
PO6X$]&+\3>^T6UJE2M(EWH..&HGE-\OTD]UBM-1DB4<DP!!C^3?>DC(VW7&'1FQ\
P!-H8\BK29-3L^ A&W/#NPVR/T&T(N?6?B^,ASG#]N.-['U+-Y?8HZ@\^H)N]GC$X
PJ ,:YQ)-36 JO]_5>56;B8\;;%#3:!B/;WB[,=R?+TDZ],(IH]LS;T]V@GY0X*F@
P!9B;N/C_44'7<4/6HQ>2,SB"%G!>4AL[ \]UW]5H_U&<6EI0S*BF1?:(\7M6RJO5
PD!+V1N!(J-NN[W6F9"(+$NF,*4U/F'>^ L;N<0\^80S26[&B[BX9JOEI61\5U-NU
P_:P:-U.YNCU2$ZN &5&JJ-(RH<!1M]E.AM8,OO:T-V6-B8OL&4S-J8]NUI@Z%BUO
PX %SK;/ 40:CD\!'ESP<L3"_1K-6%*MS+GH$N8("Y##G/Z+OJ=TG5EEW%[[^ G5U
PCX[_&[?<9#A"5B!C-UTS<IEJQPX_9G&2[%!I/<!S%5_CL#I$*WEP :/+M)_E7*XC
PQ#!U'9]'7&50Z/,8ZNC\\;+5_;=]_V08*[=1WE+T/'P#JI)"06E'?BVN"Z8OELIB
P.J-L1:&QTZB6H\4)):@5K<9B.@DA)03L7ZE$-&(.'1Z&7'W=9JYBTA6)%. 4R2N,
P.5"CAH$1[M]*/@/O=NGXIWE"$P21L(.-M>>W4A% ]DP"H4-RMV*+BJV+"G$4[VXA
PJBS[W-Z-!YRV1CW)G/</2QZO,TX?L1BBS]^S+!%NDB&%*21983:;ZT+[1<X<454Q
P6%LR)!2\N36 [<%M"R1\H&%TBAN2KQ,HE R3!-C\FY:;NQ'?B4*O.Y4H[,.& .4/
PO2Y1LMY7[@_G57H%9%OIF$&WXMS<X3/G6< @?E8#^J&6R%_W(KTG.:E))IE2I$<A
PP0):1]$R6Z@U5D)$W58A6BXTXJI(3>3WQC@$R4T'6/?C0^C'Z11=&0<NO&/"PRQ 
PPB3'],VQZ1= #*3>I#P^9S*%&/EQYN=O*P!H3DBD:QIMZW4043>43K47Y4'*W1IR
P#)$I:=(X70;V;\H!K@?_)FJ69CV=@+:XTY5^=I,;M24+5'+0#4-MG%Y=V;C[, _,
P8/((:R</.;)PL ]YL;LQEY[]3$U%7//WX?;\7"B8$DC$O)>_U6UBS,8=[.ZFS)7:
P 2L2ZF/8;L[@\3?P7H&0QSPUT@#&73Z4@_@9>GWJ%V!;T@"4NW:[F6?Y>/F _T28
P+9_DZ2S(WD/+D0WVV)CLVO\W"/^F!Y#HV*?T*K+)6""!5+M5O+%/"6HOK$:O$^0=
P.69[13S46:L#%Q5_136IXH9H!T&Q4'(3N39#@>+E<ZBAC(']IO(URVHO0V@21BG>
P)?(Q%D!<5J99G]R*'N):X/XZ!;-DQ!^LV -7RR^(:/1P74_5L*#S?+_82N#-3UA%
PJS+/9QT\&%S0M=>^V^'TOE^:@5\I,9@A[\WT805."HHYIH]TD+0.C>=CUF3D4S0]
P2B53'*9Z@Y*T>][!,27'1/CR0+$L1+/9M$"8\&?Z>+Z"RJE"ZV2"+P>3.?W7IAV"
P@80PNLF3?,HMYUG:-)8,\A3BP4=UJ+*B!HW;UH:"XL9BBY-0%D9)+W&N.L4OR6<+
P(U^BL\@FL1[$5E+RF&(=!>6[HEO]A?YR[("0@;S"UY13TH4][Y3AQ<39AE+NZ15@
P<G\".$CEZ1H',+7=/&2NTG>-ABPN0!#RR][B[R3Q=$(#*Y'3??>-!Q\NY.8IN:>.
P.63 X<<(#U [YJ=0NLR19"9)EI?ZK>*H0O0-<%!>F8"L?7EF8Z UB[#/R^-!I>\R
P")6?DW^,=2?.)_5"Y..++Q&IP;Z\(IU,'])J4E+WP(OH8T<D\S4FO\@%#T%5H%\H
P<NI5-$F2'%(Q:OD\-!>M^>?5AW/0HAH:US)7:H*Y']#?EXTCG49K5^LJWNXJ4MZ;
PM7NK7,<D25B\ U!'&.I,,Y\ +^[SU8U@CAE@&9D?N:F9+D0G;@Y4\A/.  <LKI4K
PG@C"H?JK.PL9,"Y.:#1;S_FG#SXNV"CR:E9('>D312 =1M/N@D+*WWG2(">(Z=Q&
P A/2<\KK.C!U2KL8OE)9E*"JHLU.59Z2XJFW; FZU-)%%W=$D_(FU*F,K,"(_ 47
PI -7/_SH18AA>[%?F=\1H+9_,T817KV"Q'*1(%!OG<&G _#PUE^1+2M1V;"Y)T.-
PQ@] ZTJ7 [T<1K"U]+J(/%!5"H(G3FYY?7\.QV1T<R>8! F1G$6MSK54[<B*A$6\
PE$*U-JUZM)&$J,CM3-<FFD 9>=S2)?Z!8(46>&! B@AC!V@O6("D0"QA0VJ%L8IR
P<UAX;^@?HDMVCG&DHE^&@9C. "%U@>4SSDG$5[Q>R-&S\7RY1A "-TN:<*[0]/A'
PUR78%"(&0G#JT27>\N)58U:/2(:_M-<^#V&LO+@Z+$2;K?HC-BFEV0T;=MDHMHVU
PTE_07A6*G7,G"8B\@1.J;5B+4ZK-ZW[))&<KR%7GT&:GQ6,@0=G)K>3H9_\IRDBI
P+J'G@:_URG4L-?,Q@I2$"K_4Y"Y414I.G3S=-.&'<S@'_HLP1""NA,O<<WH>#>:M
PJ'.J">OD)Q'6Z>T9G@VC^R2F4;L>P5F&2K"K&!Q1WL3X71^$0B09S;70!'Q'P5/:
P3S.:YV;6)7Z28+YC!$[R4?^AEV3='8"U22\F:A<&LE7-O'9AM0SB:\'I6=7$W[);
P$3U=G&FC;*6.8*U,MZ7PX15N4&7/L'>?,!/HG,G4%#DX/,T\#(L/(<K*O*><T"*K
P5X3$ULZS$6D-38N]JMJ>=+Q'?L%IY$?NL.X8@,WXDJ9PO8E@]^6!4P9\IP(CMLBE
P%!= 4]FH-:B.F+2;9^=S0"H#4@M)2/.AE!Q'"VKJ/!0'?;%G'H928QKZ>0:W?F@F
PM"E=LU"'+$L4)IQB]<"$&L.FJW7TI22S9YP(>]FWG-,+[!8&/,\&DY'A0"@&WV@%
PD1<'@^C#11O=QWD:%LL9]67B3"6LRU&@!YQ94I%\0,I?A+7D_X:ZU.R!$]:AHS0V
P^D<&RL=ID=K4X<&D3--&#LU'@5EL>ULJN^_,':XR&&8UL.>.^P:D3OY?Z#]!@TXZ
PLV 8I('(S(9N,9,",27*LFO<S&/.V6?%F-;&7!SBP6Q5_]VF+%Y]*EZ_MCG*DNH$
P).H!DX/9SKA>(G'.FVKL;&R@;[@&]B%@ 5!G1W/K$6-[,]-]FE..D:[G/#&O<\%P
PN/<F(OGQFJO-QMLM&:"CW)%];XL0CS$Q#EMAFZA:(5AO8 1;LXE_,;&F\_<1BLRP
P%='@'U^MR@U'P5CODU4XF+E](HO;8 8D=X-C0@O&\!VZ+ZRJ#K;MBPFH4+BS>Y/?
PF(O:.X"U9+4.;0EVZV*]%83%=A,[]$Q&XPCY^3**L6BP6*5"-F15$=]2.,+#3OFD
P#^. ;60%LR]/K@8!C[:T=O<^5^O=6SRD=4#" ;++(\S6.E#LW.33,9 .]35T%H"=
PO"86*8.9#2'ZA%)!?(5#Z3C@1Q&G+W$7)%,^6D:[1U#2ZG3 RHER@",[;!H;3'[J
P?U41W6'$A^;H0)%;]9 _9FY#5H8R$3PDI6;/5 6 10*#D6\-/3[7[3K;ZR>0R<%D
P0:)VAYF7*6BKG^'+<W0B,'"K %@3_!#0\CM@]#GUZ-BA9 RRBMAJMTV5R]XH )9(
PQ2[E2,6^@HA32&1\&(82&35\K&-M/$/*M>].@VWT\KE9%C<-:+Y@M8LP"] ] "IC
P6S$:)5R@,?S]GYOOZL8!/F!>/^_TZ*,%<UPU)195T)HRH5G-_[1:H'^S(W0+1^H+
P?0<-W+W)G_U:&#/BJ,B2+5=9R*T @P)8D2;8,(/2THBO-AX(:5#L9N4(Z*)70-&8
P^NJUT0T&!>833#W0EB6S;2N!S\RJ3DM:NR"UMN_G09Z72E(A4F2Y$JW>,L==H2+"
P@1E3Z92MEXEVU@5C7^C$!>[?V996I;]$D*)L0;7G#J"9!)@KY_I:I(G.@)L+N)P>
P-O!$1(F7CC>VFWTXG&*534V5%F4*)'&F^L6H?H(G2N[C9EA6.[PYMAK*TOE(U\$9
P*^R(7^32+ ON<YIUDQKXHB<?A*,U<E<,Z3?E6U?G GEGGYJS;O2\8V;RRQ.ISR;R
P36''+PG*GUFN5QB'>I1$[>0A_GRV9RY#I8_;DV3UPD!O6Y@'M@IH-I1Q"P</*X-N
PVL;NMEW:78A;@.?G_6A)\Y),65W92=59"8C>KU\&<GTR9:!['[:I0T-5O^Z]F\6U
P'G1!M%1[$ VB$2^3DPC2;_0AU;O%K])BX9&/7FT6*ZG,V3?WK"2Y.D0OX<-0YXI=
P[ (.G7*<OPD+1BGE8]7&DOK>'FP#>*1@,XNGOC>LO'0$Z=[:98T;=2#I;>[PG<(F
PL]WP9&58BKI [B\?5%%"'10#$L7;_M?7XM94TP:Y8S[@.A<1]$TRQ$K1LU;>915N
PA+M73"1Q67$;XM>J%X!K5:!"O75>$ >K8V/A0+@+&$^;"%FZG \.L+41OD=(:V!U
P_8T3!3G88S/D +6532?=?/<9=U<0:#=9^WBJIN+C*6WJ/V/IHZ9(GED-KG<^U*=G
PW[AF9AMU@4G4^WWV#?#U>R1E'H&D214A5R:6@FL'\$\TYYWKL^LS5QAY=7 B\[*]
P6X/LUH7!,AO205[/*C[>R2A$UX,=%$\0/21#[B87SRG*#R+GDGLT,8%&\H\&P70?
PJBJ<<6\_6P/*UH 56ZIGQKS57\79CU(1(.168)LUJV"WX>_,7OT[09N#FX6W>$Z$
P^*Z-L+@$VC65<!?IR(ZHI7RPR\"3D:Z-ZO]='P,=Y_'1SWLSHN$;+!3"!@QGVA_(
P-3'A@0T%(O;^C+^_F]?H:ZVZZ]B%6UO[)O6"W2D=83MF/N:Y\)>\M?VXJ$"9'N+>
PY!^V\4H4)-4T=;"7Z-62O*._$1ZQDZQ7HV"FI^1K3J=^Z>-5<7MJW,:EI6ECWB-G
P#_:O5_IJ9Z"UE\>TN.:K@3A=>2W=SCC+FA*N$^Q.,@&BG5KZJ?1@QMZF2/_X@\$R
P3EN&+E KUB/VSRN*Q=37)6$SK-&'9KD8Y3])$.I6Z50QF!I]1LH"AHBY9X&".B5'
PFF2AV];5?$=%#0I7LP$4R.C*[DF:_FL38%0!'"G:)@2)]@WX!R/K'2O)D8GZ#8R=
P+5%#(6VX*J"V=)DRI#O#L?]RO&'5R;SB%"5?8G2QY#4I1A+%Y7,GFS&[>11QT*JF
P\(MPTT<#LG^416,Z:UH;55WP+=%@$&!BM\6EW,:DV<D0#\I,3W[$(HO"M'7@CMRG
P_Z^>'7T[$7?)%D\QT818D35->9@[-;B01L%9PXSZ@GCY!(W2AT19]-#<4PJ@A"QB
P,Y&\;RK6Y0,>TT8NV^O7!35 &\.(>MG;$K%SC*HP&#&P]Z@7?WJ: Q>V9@TV(481
P0V"68WXWH:D0D<3089 2EC+ TVV%>-/)*X&96IAM28[&HKD#3O\-RF_X[I@W+]S_
P%7'CA,I^PA%##MQ)Q2AT''/R)HVOP;AT_6C-]4Z&]#(B?\:T-6>$EC=U&M5J&;R=
P4@=GX@IE^OGBX2NJQX=VG86MGS;U(3(=,7'0DHC?"BPV8WLHBOS="?EC W.(=VIO
P7X+EH-:L=14?<FS+PA?D <KFPF%M]"+B<R;S7VYJ%74)&Z<H=$I;'7(Q.G8][)UX
PY=H4JM\78/:C1FG2-9W0@"S.)^ >M1:V96.]OG;/BM=G!OWVV%@2,G%3-9[SZ=?6
P#>,L<?(*&N??4U2'C$OB+<;B4",,(@#::?SR)D9D,J>J_N^KLKKE13-.&M;+)#.F
PI1/\<M T.9DHJ'>YO.;(+;86?@*2Z^R[W4FV4"NV,\JEMXK-=E!2BQOK[\1TDC#+
POJ_7NSL]5OQ\+!J5/)+@6UC.^30_<4MC*=3V7Z)HW/YT$6--)RZ6S=0 _LCDW^]/
PB(<A6EPY2*34 ?I8^=,<H O+U ,%168HGN^30<G!XP24B7P0Q%W; 33GFP^6H"\J
PY!MP,NLBO_1U*('J1=5$&P;2 =,@W'$EN6 URRI.[<FH>S"L7RU]2(OU;L[+=:5+
PJO"-2)R_Y0;GI#4,QFK:22%S*@U, TG;N"XKCUQ.7KPJVD1,:T<0V^SP$%Q_7JP@
PJ>$!Z%7?;._DG%B&%L28^WX:0*OT02D0E7 Y7$Q,ES(\OPG<W_!-;\\%-?I+BP=P
P(YWBD+124H97@AM?(# C.]T=)I'9JI^&@^_[@%A>8*!_4I:40]-V^%)#7303N''V
P.DZUVX>FA,[36SR6X[,FQNYA6K05:]IXGRQ 4=H7PV_3.3J/+"I:VNCFN9/ ;45F
PAPX<3S:M0/Y;F8,*C!YDB7,P)'%; ./CE@**SGV+.3\\3I44"8<1Z$N2K/CQZUX 
P8 TD%E/EI:-VWQ=[J6$H/+_)QQ/]/K@N5VXJP>G6\U7O#S'A?DL]/Z!LX<ER@-KX
P)'W&V;C5[QSC'"K!LT8@]RO6A35E?%Z#5H^"Z4DDQDV37*TI3W#@8Q_GY/+'FK!V
P@/))=UED;3\;-V_T<)T^<K$1^:@:DH9K_-,0!'I(^E#5.,A.9JY+=E?/V?P,;SB&
P2CM/_+S 710+^3V;EN%$12-[4?44ALG":5Z&CRF\JDV?UL)"..Y^S=OPE">UK!9Q
P+$36)$S>WRD*ZVO>@&(I*_KB#PM<]I=%VK(1- '\\HI5M_8T=KGF%VS*,_D"W9"&
P>*@!EX3!"+@$GZ8DE!;5<1L^Z.+@N2G5W(B4PD7H(V(4[< H_-+"/=,3R#1'M:L!
P8PIGOBZY?^Q.[/PR?R=#"75%I=90#"^W=J@:-OZ'/!8-X52L4^"$",J[,G4[;__F
P9,,[* '12<&P C.R,*:_,JZYX39D(%!^+OCAWNA:CA*'O>:F_!SC_+.1EY]YUDAQ
POE5D(#E#P2UFX& [;;3FW2HIQ.V<]=^N(=1A!&@/,DB[T"C0U%0N7FHDYW'W],E 
P-"SMA1$:PP.\.Y-E+^O$#G_'";Z'0,S&6M)GOE.;+&D;Z!GM(S)P5"[NQ#,IRM'V
P+]PK=PFO9Z$C06_!DYZ.V5D?;Q0":% -0.9=<JP/OX:L!.8;S^(@%=NXOS\CYW&E
P^,;27>AW\\W&DKR\WMA;Y1913)DUSZLR[*%LYC(:A\F+VKF<9L"'N(OXUGOO LE3
P^;(Z[N"3UE,+3]\1:H67LI.6O(Z=EU(KO+OO-Q=ZPSBQ!&+9TT:?H'=^292K+QYC
PL%H_\UPW$U\=V+->F^=1+X!P3>?.>, (HM3$1 Z*R;HVCX'9?EC'?FF#U6=O@N-E
P[ES DQF="9@2D#H9PJI3-[JHB?G]4Y#"V7>7N\-"@<]FHG:?0QF14,4P;6HI($0Q
P;?BOX\&4XO".;T^AH!H!N6#G)AS"AA+ Y"%]<4^O/4J@NCCCF,5PH7Z5 </,WB/_
PF3(6&C(E(K9!U>J%.66](8=& .R.Z ?:L4V;^);QO__K4>.32Z4XHJ%J4:@((JWX
P@?1R=ZEE,V]FV:"S.Q:"M43"-9+S%2]+'\7\8-MEB\K?2GU'?0J#>;PG)$1JI(T!
P#,1UDIFMI5@2\]1>R/CI*@#==5LSF]G'U$$CUMDY'#:F.)L3 RH#]W\_ZY?!PV:M
P12SW_9OC9J23BU!;"H2Y[9M2L"%#C/6]I4YJG!G$2/TC[A,?^D85K#Y=P=Y2NC0Y
P$9L5XJ;?W4M_<1CRS 'Q>_14]U*5VRS7:PWE_CCJ^I09G2 &Y7"J/%&A-WM(^LH.
P8,^6X3%I+U&"9J#<&$.O/T)_<'EV_0#=816D:N]/49#$,#E'\Q&#@HM$?K/!"NK<
PVR4^0:_EATD.C^WZHF1UYXDW:E,D)L=*-"S9<,+7H^]*+GG39X?A[?P33,S.^9WH
PTLP+&I1\0C-%T- V_L+R$;*G--$G&]_LVVK5X!*ASGW]Q+?T.R"^.7;R$\;SNYA(
P<?EYD4>&W7M@@#HTH_"%S\5W,$-6=Q()7AD_$F<*W:[E?L,R)^;<NK> -B]3D.22
PC]4^BABW&K]/#7M4?>SFVPVF*C24-A]K-'&F6HKCXMBA:D9(ZTOQ,#(:3%](1LH'
P8F$L%^U+';Y&)'+YR16=XDE9DLM X8950I\]]Q#5^CP;96:/R =L_[^T?JI2MNRN
P4/5!PG/(ZPV&4B.FD4Q/Z(""PL[-6'WC>C+?PP;<!EVJE>)+AFT)-YSX-/R'Z/X4
P9*YWMK[=#3%FWLR CKFYO;V"W5!W&.0<'3+J0N+H.LF5@(3^350-K7V72=8[> AV
P>-9F<(AJ[7!G?MJF@KTDRZ[2$7E#SVE__2(7EXX$6)_O!0*^7?\*NI(5*UWD'Q2@
PY$^@7F ->$QK \B;"<1?IDQ?+D:.XXCJE%.838K%6"ZKH>Y*]MF/K$!R#%HKAS0,
PC@A$<ZT-9#"_1!3HGU3QGBU&S05(4M 1V)FB" 2V!N,S/R.M27$GQ%.07]ZJ<I^?
PV5+P,HB2SVO:D^?:T?TIM:'NK3+8MR;9/O$Y+&KB\TWA$A[XV( _U1!:O')D.^YS
P9X:A3C?M%;<$+4U@Y@2#).>2@"LK&<;'UYB$[#</FRR%-X&V"1-+"]!>NEJ\7P-(
PL"W,'8_/HCU9<2^Y#]2$;Q^ACPH:67?B<&/=$LF5Y?OB19))U7]D=7UY:9B8 LQU
PNE56U08K=3R\ML9!7&)<4@[MO@#0R%<NI33F++1;2/.:XQ[<RYP8YNS GLT2*K,!
P-0<S5ZO*WWM1JW2B$$_:]#/!Y^>D[0];#F8.J %(,K5#JOX2Q$=""^"\M(A ^^NE
P&ENR:)]KN9QATG'1*\#?Y.K%UAB*D943%,HJ,)$7*H&VK^.SVL[%P^9H5H5*4]L8
PC/9J.N['0LS OJLB29,RG1,I/4AZH->>[JJ](K%FI<<Q#)N+K) 2!!))+R\2<G;1
PX)8EY_WOL-#[\Z_.%)"8+\YUV2Z'(8/2G,A4J?%M=446Q$:X%*'A%>QDXX.9BEVT
PPSN;&L0)Z)O]WP64D\Y<I2FAQ6RIL-]C^7U#XX^F@R+!*,NUTY_?N-R\B]GWOMHU
P/_+N8I>8V3&DX]@1?D^7:)![M#JPU)C>PX%D-WO6_:!-^K;)/P;(^/ [V7,1G3.+
P_S)L6N2 [R*"=HKY3]:VM1K&?I ?TF]73?)DY,J+-P#3($D)B1FSN-#/MR$8 8\3
P=YJ8&&F3Y &J6RB)5O><_LYM'YF@G$9 !U^F%-?MJ@'@C264\D<\CV/K='.)_>W2
PQ34U+\!#H:MZJCG4HC0H<,Q:;Q&_LK>#S2(H5(%/!:XX!+SUF]M]=AFA[_G:(FRU
PY'E5B^%PHLZU'V(9:I].Z0%[WV^SO[(:J.11,Z7GVTS!],6D#T&\4+P5H>8AH+#%
PJOB>6A.<HT=5.-B4(1KWW%QQUYI:\[::/6#DW7(>KB]Z=_]3R?=$A&Q*^VI^HEH;
P:9U08<-IR@6B'A5HO\#DK@Z^= [0]3F\\VPD?M+C00"0+7XX@V13G:BA_:S$RH:5
PK]&T3(<SR. _U&2+&A*D2&,2 /0^+GW#8_7\$\30GJX3_(%;!O"(:+$/2?OUL*Q,
PVPO_7-"6*Z.[5.!.P]76\/_I2E %I& M)?8H*_L328&M]:1%8;/YJV#)B,:<\< /
P\I["?ZRB!XB5OF[6DL7E@Z(X<%7(HA!%FZCJ]=_O\<U,7S14%IFD,__O@/_3F&0]
PK:_XN<6B1I(:3(4E<2"TMWT'N=^,<+N8)XFM!1EM__5/SSF/@GI9I$8?4W"1V5ED
P*NS8\7VL:0Z=4U@70)WJFXGFV7GZQ$>Y @OSQA \:B9%O+BUZ5-"5.ZF88HC<Q6[
P3P0,ASF[XIZBF?I.#!3S,,UF8DL['<J5-OIYU!;DR+?\=C%%V:HOW!K JJP0CDN'
P<];*F* @([ .6A3,<K9U-MUM3^UG0"HF,P!8P*!BX9,\SZ!GU:,ZLY9OB41% ^^$
P8&?!^FP2B)?MU8L" Z8CI3X(QO'!$4ZX@S95$6J;\#'CD'OJJZJ!E$;$Z,@4KU?9
P\VDBT=>6F96T_8= .6[5*;XJ4X5(GI_2H,LU.=?@2!4XOE+J'PN>)_E2)/Y24GN;
P7^"8^;>A#LZ,"E[RK9SX%IH[*6SP:9I%^8(;KO61E8">Y#1P7/G;F/)7VO"7]N0*
P)^@VMC<_DLX+E>>OCP262J-( 9 ((+UU:K%.6$A9TAA_#,_,%)2UH\HEN5?,,2?@
P)V:[2Z&546I+% L64[[C!(2.PM]Z?$ ,F%][ZZ7EZ&I1S[ !.6V)&&*9W?:FB!_?
P<U2B\ZUJ7V*T]V'<BF,F O1HHUKPCZ^]$[9$%[N*^3Y+J0&"P<L^MP3ES"E_=E1^
P[J%H&N_Z):Q\8Q5!_JB_ZT:[QGN>=U9*M@3WJL*AD6_H.XL='E5!-Z(CY%4@B2)L
P9,%YG;08:Z0@-@PM^KB#VW:$=THCG!\-+)6S-GAS N[LE8>=Q_7?!&V5;YR\0A0U
PS&ZOZP\VDEQH<OJO#=%:?6H9$/0QG8I)MIN'C!C0S)8@THD0%X%Z'I3^$,$H<'>L
P U,:]')Z.]#;;K&=U/A-P4A9,>'6/OYKX_E8D.#21K1D3!.W"U1!KR4'RO]RY>UM
PACT ZLD,* I$\!;</G)A%S!Z63G2B?3>-T*)3>U#'^63].;JDFX%?4/VOA>HQ-L,
P>N4 [(F>X=QC-WQ;8S(,,6(ZRNQN,!:7FQ>:ABL[IP&(UWU)E.Q@2?KA;\4O[P]X
P#&UG[>\)Z_O02G(>3EH[T(=P0YGKMTAU\A8Q["A";:)6.9\E(-71CN?,;5<@/"(#
PX[T6T8\&YFMA+J@9:?=/1LSM8EG]\OE8&<$]>0.M4H^20M%,7V,ENM!DAELRTMJ8
P5%H9W0[X8]_%XF[L=7/NE"WZ?H<:EB)SY,<,%S)XFPX+?\]&GH5M*'=^5M >+(:A
PY.V0,^JXCT'/JBVC+7D"%E#QZPHY&.X7_<R5\!?DQ1_C5JB"BX1H;4C4E!L&:#$Z
PNUCI8:OM5 IM4LE?=E?4:R"W9,02NA-K@_GF(/5O?>-S2^R1!XK#LH;^L;]7;;-G
PYRF=^26:7*YFSJTGB=IH5J%S39:%WB-P-&">ICA6H/68\]$8F^=M]OFR3,/D.C2<
PRUCK_Y@320)L0QTU<G9UCO&TKA\B+[1,,S\V%T.V^*G(PR%!>[HU.WPLE0 GN]8_
PLD -?V#:ST]QD.TB/5\Z8/M;-^FOKRH2,W74L@:K9U$<B-=HG@?T#D;<K:NQ$96*
P-V@IU1T8=YJORHY$M#W$$7]163G\W[X," [I;"1(>;G<C$:<6JN9]2L")#Y\QC<F
PDLVD66:AX4VY#8V*VD+UB<?R1D:*!IOWGGTIBW^C-3LK< 1OJG5:8'RPDO >%8T*
P18V/I&'J1AGX4WKSXW6>8_O>9Z?=W=J#ZZ+CN9:*)F[ 5!I[,TBT2T;D,:<EN&;9
PUOHEW.*+KWNB.B++JSM&HK*!/&C)9P/4DN=ZKI:J^@_8C)<TX?.6^)_D=N\_5*3)
P$,\*727*;<2AS:Q6^=$2272L0\=[^#16!GA/E'Q9>VK;IUU,>RR ,,#=0. !AA!"
P)*>,:,'9P?AE\>5(_B6P\751.'V&U/CN=,QHCZF'F>+'[-BY(E6ZN@G!^](12*E?
P;6P[=BU8=&!6,8+2:+W5I2<S(85IV\=X<=O,;E0R8N4;;BIW:6 ,M;X540-%\ZQ_
PNA,)+)J@15LB_,^:PY6N5.MW'PVN_)&!RM2@LE_3M</QLKWI1W;KQG'/OB.NS-Y$
PI0Q?'_Q%]S/1[8S7@P/?X,Y^)*LJ6W/LVVS(T5B:*AY&0=W7UT![!ME]Z+&RR@O(
P&CSJ3>W;,%%5>S"$SL,/TK=EI$M.71J8UVCR$O91ZBNHNZI$K4R' J>U<BM:&2*B
P6QS=]%(I4^2L6&F^LSO1Z<X4G!XU)\@!R#R]GI+OC3T$9##^ZQA/LTC15H]FOX<A
P=Z<N SR>2$'CI74?K&"YWL-VG)MU /GKPJ)U1 >ZD0ZP?/6J),".\TH+T7S\]3E^
PF-E5JDZQ'6/??5%FT)7O\38FU$*C>J")> 6>;$TB^"1>"NNSXG/^C@/QKE72$-B%
P70/!G0\H!<>A;W'=RSRSO8)/8[O@Q7AIZ!B&6K7T#<Z'0L9VD^_X8L"!:9QX^CAW
PT-7$*ESV]-)I5UDJ"/^"/8OV(PUH\A3L6(=28KL0\1K5Q60"4%_+LGL"(;]D$(K+
P(',Q?J\RYWX9UV((E? @3C<XY%0_0E"(S-&GX-X@\+L_J85-:694BO&]E?:VQ)KV
P[%_=Y,G&C&A,50#(OIYLWC.&NF5 .4Q"4K$B@S+&DQLM3P4+P<_YLF6:P@BU":5"
PMTKYMW!Q:ZKJQ9&WL#/8&M9RK2T=YKI=3NUL\!Y83<QK>XJGI?-22K_RL7TEK63]
PJ>%#MJBS?P1-8.3]W.\8R$',;N9-I+NY)#'6S/8/AO!PW0Y:[I#W>H_@3O\?M9AC
PR0NQ_.C(3&5;@%Z2:Z"@53,MLE8T_"';M?G6XB;T_%*@U62\Z.XPG;?MEOL[8[$ 
PPQ55 :16J.WB=,GPEAA_@#<ZL[4/4(@0#)GZ/4J 3S-SX8IA'?(3Y6^;[:)AM(9'
POLJQ? ZSN&CX>-DFJ)%$6-#X .'ENRU3$=>RO'7$*JP2]HIZ=U*L<SD+ W1%JMHC
P_A!/GX]O]J :)_&_*J4E;*&$HL'X5<*1%@F1%#/NV##?'@5/4X!V<^-=+)A/0#8A
P^4%N!5(] X[(IQV-.CK4)*,7O7&_8C%[M-;B/5ZE=UW&Z8%M _>:P7;6;&KQBXTH
POW+)Q?A*SW!Z'>+:'O&L>% 8G3(P< :1K_4F5=[]*,;[[?3P;C$JL@5=[15R+5E1
P0*["-D"S#F3,D(B4;-U-[,K;C.L= 1I!, /&[1* &2KGUW:H-PHSC!ODX\\+U/>8
P7 $PMX(C1 -+)EUTB[>$G5@RG/TB,5[OT(K+1PWN]U* I:%/!=RRK]R2RM12Q7X@
P)?KNU[87JU6P/ENMR@X@"9R0Q*I/!V""/+KO5X@.T8A&76')+<0W^J>AO-OG/\<&
P[D6]>8S'5SO(8#@Y5; 1",A%7ZD?S%6->LV&H(VBD:^<&#T2&X2GO!4]-RI9S7#D
P1; /L/&2+#+XS4/#E:RRD<M\/MMA76(,NA+/CW^4"*YT&G*2 C'=XY-<]_#YIL=R
PF)0-7O:Y&!AM9"X)C?<9XZM=^VWVP=>+0K8Z; UAHU.+*-J-BW_&0_U[%CR)[V9Z
P67(X8QMPD3'0_<R#,&_:ONE;4V:9NU)HDA)*T1/5@B(S5.$NG'P_$+/'G</VO[ D
PNDN,MAD8]K-+3!)R6"^B6*9&"("F=$?]/_3YGAGYV?U>UAD.O[U8%+S,4?;!68Q8
PI'@2#L]JISMA4]/CN]=L/8)O!R4^%HZA1_.4F0]J.H2A+R<*G7S^3=;B%"P!Z"!D
P;&L*.?%H-,(-AZZBS)KG(@S-P[:(+!5:M(5T-![TL=73OXI)9"FZ_ES?6U&N6:)D
P&J<-:1H:(&D/&03>N<-CSL;-5I6:Z3PV>4!Q0CGN&\\(Z37[/;5>56ZN."XPV4*(
P#@($.\=V'X2$CCRF/YTRCM$BS1#((-I58TB18CXJQ0DESVC9F8W -\@<O'Z0+^@[
PAT=#"LA002:Q)#1C0^[_:0RNT-BR@!5[!!X.7&;TX.PSJY$BB%31*8;)ECJ9]VS.
P@@64PAI;(K4ZI*M2FC@MPXR43;-.KHVLL+[.\C^:J>$6G->\&+_Z3@J$&24>+DGA
P82><C__.21QH-RB&9^, TEN1&V 3@8O8%LG\; SUXM>+27[UM:( FSF.G=1S>/.R
P.]Y#-A%2N.^5PXP7(24CNM-3O^X/1!C&(%8KKO)(=+^#F:])Y1;<X\&<)V2??'QC
P((-Y.E]QIPB 0_>>:N=VW[K%&PN9&\!W3AAG+M ZM+\(4Y8]NEH=!OF_DAXZ8SL7
PI^D (/.#:H]PLJ*+&=M4M-1H@&XDAED6M0;-*&_(><\9X C#G$7#(6:(YF.57J'M
P!-9X?@"&M0)-$<+0^S79"$9+*P;IMS'89("TXU:(,JXG&6:BW*HOQRO5LCU&^V3C
PQ@-SZL\_L31N)GQ5R/U;K4%Z;W8#)MCI(#/0+9?+4GMA'SNUQE0W.\+ 5E+.8"ZG
P%U:YAC8R&6D\UC*N:)4S>:AD<'RBF*"F1LX-3L74M_P$PM^\&;:$4S)"K[97YXE.
PI  [+1+0F+]S6ILJJ"UTT(>ZDIAI OFZ<">_07'=E^MU9M,-Y!,7<F8!PFR!,_;.
P \'OWJ^\(& \8BA"A)@B\HRK/CLNU>H>V,(?SE$PXWX@T<$^(<%5311R<.I;>,_E
P<\ "SN_5."HX?5 )32B!8JJD97Q?=_^'\!G,4)3W0[K^UYVG"G,*T@FA>)MY(%,V
PB\TL+IG<1(- PD0N/1];U1]':[A)#L6G5@IOB8E:]UKS'V*_!*7X1*'L(:AR[W*1
PK3H7[WL;"=SXZ;F AY1(T*<58<'2G^-@;5AV!";K(*QM*OQ+;=64U.23C5660UI)
P_]*^)VG9WY.UGF?B3N<2S"+;.HF/GN-+%@T-X%6KW+QM6*#/[]I7Z-'5=I!_YH/6
PIFJ#1]<(*ZSYV=$Z H'L^A2,Y3!7?L.<8W-MF:E)?^&X,$I$:W26$[#P_9EHG>D.
P&_L$-1H)$,.Z,SX65P/&=8E;R<3Y9>V];:%6LPEDIL*D<W$NV7^RR2TWN !OP;OI
PX= F1M3%%K 6VUKL5$)_79.(%LS?OIFIX5Z!'8Z?FATJUWA;-K>S19*8!!X(XB;@
P+>F1A<#MQJU#9OZ^X$G*:A,L/!1[^F91/\3+N80>I'U@2AZM-\MT%-I!O4RF]^ZZ
P=7<>V3Y#P8;MKG-GCA4/Q,.4++2=.#38_7YM1AY+<COLUOGJU7[.6.N[3/8)5R\R
P+^20A:)?#]Y&?+-6=0?\C1HXN.37I>]'<0K+7"Y53]&CN1Q8W@288$BG)C ]UCYT
PJO*%#]HC-,P+R*K3$VJEO33K=ZE)V?G:;'XSZ!._NTO5#M DA^S][)Z?1VSE$A+S
PV7Y"MON8*48?L'3BD<"^>BXP9!F4E$!434)EMMZ%M*F.?M[&*9:WE(G#I$9C7/#=
PENW"3LONG@!@$_5TA6M<D'1.^=V0RC3FFSB'GQS[A[>/ TB_MOL@'OO:!$@'2HE'
P&MHT?G9;?H)$KQ/F4TW[+QL&V[C$/+#!3I=VH,OTZA!((:ES=G;M-<SY?S;VL@>[
PK]DI0S4R%^F3R&I_UYT?<&*'!AT@;W%I:)/<_!QFH8J9X54]F?"741\+>5,MEL'/
P,;SM*!5PJ4WV.40B(T9'31&#A2#/J-L8!#OV_W"9V^A$=I]&+C23;C]WQ?+<@$O;
P?QNL7&]ZJ\^;Q('[YEE@/U//A '6HK[^,C=].[_#LJV2V(]//>U*)7L?KN#ZJ*YU
P"Y263GB6'U#KD5)*6QP&Y^5/^'F1W!$'!!62N245;G=%8;Y_W=13''VY*U%?SB=+
PL:N*UCC2U3;'#L\P*ZB\&72;I#M=\[S8^.'Q%3% FH(K?2:2NHD!8Z["!1.NF7Z^
P87@. /D"]*A9YGQV.M@]>G%H[ E\6VK(8F9?IF%>PZS'0,72<KR/(CN\[+R-7L]]
PX?=,CX1'_%QW1$QV<@]389F%AY&=8XB>$ _>@'/&*31>\I)/&LD 9FD2;[F2K41#
P7*HT-\+.\(=1AG;S&@%*FNZ5'B_,69O5ZI4J )0IQR<# 0"?0BBFT"X)6,<Z"/FD
P'_Z1\@H,Y::K$_%1B:@TO#S?;@DR(<&/0YXC8YFK!>OA'8<^C:C]GX^M3\?6>]40
P./RY%;PY?J!6NFJCNX\,_X?4R\8^$W32=2B,\)1MN\U)3!4IF?"LX;]1[T]36KJ3
P;\K1V*1#!8;H#_&GY<P&^2<!9Y30Y)VZ-"4#T-?^Q;]16;DQ=]=6[X['R!Z-^5QC
PMA.YA&W3XGQT>3$\SS8@\Z"X;*:3E282;Q%2F3(%%8&E;M5K>ZB"]I!E_K7@Z5R9
PI_3LQFOB%RVIVTP: _#MI%+[6#KZ'S0O,G,ZZSFKJI+<D9EJ\4OUQ$B?3 E^9'3%
P"D;7N>Q$VOL<B*.)8BN7!*C%99-,F&S)FGS3Y$TW/?K0Y&%EJ84&(4Z!N6D)R7BH
P3/:\Z7<>85$+@3Q*TC%8W8H][$5NM*6MW$L^[6SCMYW^S9\7[*C>P2E5S;%]!WI0
P#R)3TG"$4T1JT5>:LG>CGQ:-?D3<-UEX9PA^D4R.Z+@-X>N]HVK=_4SSXT\7QAR>
P_6' 2V.9::"MC 7NO ^8'>[[0T#-?;VY-^2+2)PN&Z@]>3*G!X@<W7GA-SY+M 9;
PK,'LD9]\2\4 ^N\?P[WM?$/%/=Y$^OE7R-MR^!OA7])J4>1Q?]_;N">MIZ!:C]F3
P&QQJH8N+[N4<$_7,=#]R[02S3GR>FEJF7QM*4I0$&U]_(%UU>@$7JKW<1N _1AOE
PZN?OGSJ?:6(7LY00L)6SQ*20]\A;PDI-KW"1#=++ A 985:O'QWQ  P^T&+5#0^+
PP22.&8GWBJC9E5C/>8UW6F<]61XE%,W\KS[T#TRFR4L6[[#2QLOTJN%(C&AUPZPG
P I4:'\O_QCS/O=N[5</QD21V/52?.S'9K_Z55P$KQXV%K R57HF8.I%)@ !OL.Y.
P!LG[SF0OV4(:DDAGZZYT*UEM4^H&<F919[/CJ/D!Q893\9+G[ )CR'."Q:_H\AJL
PZ,._]N9EHQI)6OG@=WLK]G6-JQEQO*=LC"-2;/89I^47DF9Z#OILCG]\M>BSZ0TS
PZKB&\-I#>UF"OJ-L#.C,7S3-HA@!1#6A[/5ET$9R'(::[3-'E8,99L9ET(B/^H!K
P:N51)R"O.2X'L8P+,%X>X>?Z^'.7XT<9@$A\-GW'7$E?IU+LBF,)%U0TT6<$J!^Z
P,<3>N%EY,9,-/(6C1[8(J-84)D4MWALR=Y[=%!1E@$*0'(=&G5"",Q0Q%JSZ20\:
PJ_0%?JRH4$7:0E_C 7/TK]=T?9R\K\>OI4O<.2@ZW5B#NR1I!4\*:WS+=_N %,G1
P70[PZ2/MOO)0]9^,5,8\K#LZ]\$7O<&8;U15?B$409335#S?-B\OH2\S*Q38O^A[
PQ%CWL7[J==ZL!<[!;D?5T+=[F6WOO72[0L!8R.D?^,C:U[6A^[O3_0;POY**L9KG
PX"$5<=6Q$_2Y]TCR?CP;.>=B(A2>^KT*$V7RAP,?+-]]GT[VKB>J7U?";YF&]VE#
P2]&+H0UA9E[6TY$'$E:'N '+':%/ 3UU]J\4UV9Y[OD"_)CXLC(;PM2%#WN_)YA1
PQ_4V]69X\J^UQ<6&1M"0TR?3 X)@46^)!!&?")6D,L!Z+JS(:3MPH&8,.,OI[HJ2
P8+E<7C])(T"^@[CWVPWA=AZX!/J8TS%0!5II_+PJOXI])BH6=+8U<,ZE\WU&^D0Y
P0>_#KNRA9#] $%.X2A+V@L]B)?$9/ITBMX\_'OA2U03"A@N2>AXDA&0_E][$)GWR
PC)1N04ATJ&3.X$(8-<*YI7UPL7((J=/<_<[Q:X7Q#9.2^"#))=H6;K^UUSTE)4Y;
PTFV_OP*]$[F6@YU7\YGG63J<8-992PY=I]_2BP>[GD!7&HI.RB&>"%6/@MRP;%6D
P+7"U*0-TBA8B=;VT2H+O/(E\)4W%Q=+_W$6-@0:(*L5V0.92FH\2KVP9TBTFW_@&
PIRX(J7=8_$M/6]_T?<5#?U.L0' RDN:O=@>WLG^0_49<<A6>4=G*1I5,,UW]54R]
P3M<<I_<+;G%5L4CQ8U])7'E1O5AUNO]CPBBWE/)$A9.#WBT=:MRHWYZC,L<.R+I,
PG#Z%%.U64A\B1EJ$Z 7V@7*>-+NQEZOLR%!^N5Q6,+_0'8\S_LD*8@649[45KG>.
PH./D]*"'=V"6AL<:JY$<VH+V2G)I"A)0+]SJ9;34\ IP[K-.C?;\@NB2)C0GDQC7
P_,P_8TK/8!X?.$$S1?TS)WPTU 6VC);-D,;V6*_YA&-L8D&LM,L;2H?I0PEJCP^1
PX\,'61R/[K;<M@[+HP*Q?6TI_"^=X-VFA$=5AL6H86M^X=;OZHJX?(-!S!A/\JTF
P;ID.@53XEA1\BMVW.3!6+#5 $>[]G8U)"V9L%N\+FC=.K$5<PKU1.JL LDM77<J4
PF$UB3W9V4*%,$H.!%"$*^$_VEOI%=U?89'GQU2A[G^/K1"!Z.M_FZPZ=O_O*-5;)
PW_P W+=K0%7[08!C45"PWYEQ!\8H"V=/2SW'L%3_S<F,=5 8]WXGEF;@*MC!;+,=
PK ,5TG"/T-%7>?6K:BX%KBN5@+@%Y4ZX4%0."R2SG*DS=S>.'?KI95>]5_!0G+_-
P/:-A@WLD&>:</8WP!= *'RG_% M_#4-!@YHZXYOO(U(]JQQ9[=LD-HT#B%VI&M5B
PN*B@.#(*0X.)OQ-D$&33:7CP.^DN2?60;:Y-QNU@+"O$)2:Y467^U(W4]D5X!YX$
PZ>TCRBL;CR<DY6V=,"C$*73#].B,<Y892DZ9A_%//PVG6>I]12-I$;$UU"$^M=3V
PZ7=3OETEB^G6N2C@2]BS :!0BS5]5HC:_76\QC'=A#Y11-M W>A69%X\$)8<5/++
PESH([4%7-WD8Q4A+,+3[^?20R6-39YZ(T,LOYHG!4%^@HIDH__@\*AD1.ME3YRE3
P5/M3(]"=-W5!**_ 5DISV[S53W5+ML$W"%4S+N;!_"(?ORRZ(C:2.X,/FF1\P!_#
P87SB4.Q@RDV]H@L=%BVB#^QBZPX:5D_<A6"%:UI )]4I2'W2(>4V$:5&#R$S%IZ!
P/.)9RM V(83A4/X]@.B;ZZKGSQQ(4&8=N&H1-OH)*#?5Q-!LDV#'RW@ NJ=:)OT"
P5+K5>0(&W%>58TFXDNZ QX0YOU2Q38ASXQ%'[?]DFQY, "SCB0N5IH$AO*8YX,N_
P5W/:=1[LZ>+TM*TY-98"(/\%I!]']?<;/%E;OH=Q%P/N30$JPQ76W!@/L-2'33P.
PZZKBS;FK%'03Z^06R,4D3%J;3"M+21_I&F#VU<(C34X6QY%9)/[_02\5D5)+:2";
P*W2!KJ;>/^;MV\#?.6L@F-3KM%TX)FHM:C<:J+OHVW#@O:4P#9"\? @HZVR8^MJ>
PK>5$'K$A810QA/6T%BU4GK(M0)G\OE3&1U9O"D?BA?PMV[\_5$?BBBODV0(+!]>8
P0CB/#B,-%X)OVDAG:]J +_(B)E+[%,@7]>*PD8%WC6<V!*E > ?XF@V/T;NW(($]
PF0Y]ZADN.,F84V1=N']X-C5Y]K#+$/N6\@_2!3?3&@Z*0060KJ_>G!^#A$1IWA9B
PZGLB!50_17 I=/B/=G.X'NKK-GU'<KUBI=7K#I9]URL'3]\[J)=N,<1I;B=;VE"A
P'!Q:MH@83/W6:_E6S<Y>SP%H&7@^5;%X(094&VW':[UISX=4J]"Y)4>8Q(7O*3M0
P=<U6(Q3^+>W"A%@&IN)3V@U[+#=H[JT]R=/<F :<&LD3_?+Q71D8H3"=Y9<CVF4O
P4S&!H3U:<F]-]ZU/CGUSYL'F "VX;4L _CZPX9-R2P8<KJ/R&P <M&%2VCL6_Q3<
P\K*N,P[U]4SE</Y5K:)'4)]_C#&P_A.'PMG_-G7U.:.-H'WP/R])LV"H%D/S2XJ/
PO4-)@89ZODV^+M+8<L*]++ZI;+K2A55HBQ<X@$K#U\6$/NV:,+(FI C*HY>%+8;/
PU7_2ZV/'0L1V\M0\F2K@9KVS9U^_M1 -\*XA=7.HS:8\+7AE^R*-07J0XF>:(AUW
PB<5J?#:Z)AI1D4KKJ:J7+==4:$2\UD(Y;W"QXGH<X/$6X[MNZ:AO1\\<4\\WX\B;
P"C-<V[9_4'760*G16IH$2ZX/&9J'^) OJ?).0I$]SG;JY%S0*:UP3+9OI4W2>(R&
P[&ZH+35C@*UZ55J=.B2=&$A=6YP;QQQ<[NTX&U+!%H1*XX-,SU*/^<G\7;@KF4#'
PWNK]XP\8T^CO:B*MD/YXN3,5RZ^V#NSM$-W,T5&_FN)[\XR2%@:F]RLZJ/^SU[Q\
PD%=)H(*5;XW7>D( B\6=WF7]!).;ZT_( @!'_G(//%Y_+S2"H7NU9RF3(PQY.W1"
PKR+8%J1/"1&8H^*<CIBYVOF<$(QN']V:>H,&?R(AG \3)U?@1PPK?45!,@.ZMUGG
P)& HI.Q2-"?^E0G8#=WA5-S5F4?NA@,<*-_WIE@P)Y>!OG-5Q9=?GTE,&(;Z\K8T
PER5- ]:OQMF_7FY!IHUJ7.+F0T%MK8^S#VW-VV9GD9$("'#YQN=73#<1,I'^D_XL
P@EY+AY 37C+UC'E3"6T2W%O/HKZ8#P^; O$?5\=1;KAG+9NL2<V7;4"(U:!@ .4+
P78[D65JL@[N1Y??C(+VO>WDKZ0 60<L.#;' M^'C4V=^5%!R=P=Z,+;Q0*A&@D(Y
PMQN@2S'M&5M]VOH3M70FJ2<__;\R7(:5EK";[F^$WX(U.-JBV:<Y%U6DB?A)#J0H
P7.;)41WG2V<W,"(/.46V"/9-=&$QZ+]9DU]VDP31>RP7+1)IHOT^$P;(2IL[G:?9
PR2BRDB#!VD#D,2]WR$*PT(,<K*'Z8QF.*KG?:5IY?)$7 7U'*H,UEV]F42.U3Y8T
P2:/[H@.,>TMUUWY@[P_&S,FWG/%]DDZG;X"4+H'KL0U^4*/[.FAZQAB0/DB7F?*-
PAA\@B]&%$OM"1KY_RLM+,(D\X8\XYSPQGU$Y";-\QZO97N4];5*3'Z1MAFIPK"F]
PB8Y5OC!*00QUXH'Y$%DP9J'M.+O(/) CU/U._HXEX4SR$[M]+D>;UU]>RV;0S8]9
PH*S1_LJ=;3#\+5M+ *UM@]/&%75B]6''8@F8W?DR[^Z#L9U@5G"^ ^?+E;2=>>+N
PI1=A^XL@\<9E2ZROB_KNAFHOTF$L <3X=KV#QS26#6V=)<I=U+GY  T-FJ :#Z:M
P?/Y5DIV[<_GA.$37_0R-WNKO53T;[ &<?ICM29!^A#-RG 9E7^GU0XJC=W/KA^)]
PD8C[><JI5&FS^NBDC4QF7UABFYY\9<OV&/!?5'[WTIG?'CEH9CV4^1*@6U_WDXO<
P-=G&R*CVBGPX=,U0%@?V%JO[*7HCQ%GL/+CX@$+G;,FMY1;;+CZ:(3TZVNP!S\E 
PF#91!8&(U;_W'[]*4JZ#SL:C?$*,E?B:#'_^CZMHYK^>R-G-O_^NGY[6BS-C+QE6
P?ISO..#_47DIW2_#H A$"]ZV$=$D'1LV]%C=RZJ]@CW^D: R^![?F<%<[K6._##M
PNKN\?*>>QJYK'*3&]75(T+13W/^[FLE29PEXE6U0UN*8H/65!XI>M7[A 7?MYP9+
P*TE=I_]Q[X<-,.7+12]&//$JL;A[)O]N>><?GF'ALG+&AYU7-1/]%WA>'T8L#53J
P=46)1S]",*9QXL';0-&25U.URIUR3*4'>T _'!CVVZHU"@,C>J-;9D.W' ID(V!'
P&X."Q("7[%ANA@"B+@G6PNAA)U4KNF \&H_'P4,!>*^'XH5E<$/AV01:U<F75<0:
PAE/T%-R8\MKJFDQK)#M4B4%MQ L"ZX#JB&+[]RIINVZBK5D ;,(E!QM3I$V1.*:Q
P8JKV9.1V$"C<[0E21_(4S*#Z=.9)/Q?;%-#HL9/#6&7%?+NV6?81>KQG=0GU;>P"
PPWB-N.X1IH;)J(6%" /8'Z'LAY,X 5$]"C97]'R7""=6ZQGPI<1J Z,KV6O,#[T7
PM2#*@)9P&O&+6W*4-@K"2,6](1+UU??XN8!V\H%K_^>FOKG?K0\,+JH.X K#@)3Z
PYE3CE-LZM-&1):N^H%W^!MM3;H3AO;^_=@FMO>F4W%?Y%Y/[B%933Q!;N!3+L"E5
P:W!%;]F=3.GGG$0/XK$[B$F5./^9?8>&6%[3S:$/]GFQ!S(?Z-,,^/BZ Y%#(II@
PSF6</9^7Y,N+$=JWNG PQATB)+2P'R0\%,ITT,:_ &D7:E#//:M5X11'O,X7);';
P4 OZZ 6&;LZ0/<YCPTH&4U85-,MS8","-^^T7F[)RG9'OFE+@I;!1R=;ZJ1N6"GM
PQA4%<\1$\ N 42]/???_9[FG'[- ]OWOAJ!4U(NPE6/:(<-'NY6JY6<UVUB@KIPE
P?SIH@&=OZTB(9CXS3"*[5%1!%;ZI=O),9/AM&JF!<O?W+L #:A,0*./]O,BDD64&
PY1XKM)55487SSO &-;>BTX61DU=BP,[<4!$-VA5< M5I2P#3ZRIARC]/'8'UNZHR
PX))^[/WVO"-V^"8ZU %ZK;"Y?J6X-;BUJ'>=BEE_]HCD05"D 3=AT6-@ 1D<7QL9
P, 9/ (I]>EG%Q?OKOHN>)K:!O)NF\PW>-2O^CAG\=F$&IB#N@&T%PE>L@C)FZQM.
P-=H>1YY?9T"2D'Z69M%U+=ABSS,]0W$QA5]/7_]7%\(#-LAZ*MIYF/["$O4E\_,)
P3PCF<I\:IMRGFB7(;80%\7E_84GA@;U8VS26]:!)ZYP (;VK(@%-Z#3\4FF&5%H.
PH[40%+@7[[J;4+OC5LU&D'CN"3\ +<:J6C/W.ST DBFVAC 8C7@3,U9=V(0[&S%6
PUHQ7]>Q;\$K(1MM!W.-E /1=C-FK0KMZHN&0'$9K@5GOV,%;Q8N#&#39BGZ#9UQ5
PZH*&1>_MM7&&[V6NTPFI^L1 XMC%,K>@^^EZ!*N\_W5,B9X4RJ3X[W?W=G!6JR]R
PRC8-TAK;^0U5ODSCFKL1>]:CV7Q?>1CO%V<K]KB SF[]/B"L^LF;Q3HBNH5"5!BO
P$4?$K!9(,3'-3J:590MH4QX"Z>VZ,;")ZXUW^@W:BX= @[!'^.9(:M !GT^"11FK
P\$IYP?8<3W=<>ZM'8[TTZ6MAE]FVEN%\Z,\5VW5E^-TTM#.!T,I)%&D(/B[A!'Q1
P%BZQ[&,7CPHNZ<VC)=AO,X*IPL="I![..J:N]GT/XF1WY,(NL:U!@<;,D7B/-W'4
P5MC+.,8\%^&+YS;_-WI+.,^EH,@+T2B(A6J0 CV7 %-+DA)O?>1,2SE4-M4VHJAJ
P(IYE1/XJ)TE'@^CK^)G.OG:U&IN(-3JD-%;NGN]4I,VC46 6LK@IO</R_!?$\&MI
P3;\JBL]&=*_LN@4,2504]^<*QZN"1YA>#;$+(D?D!-Y@</#MZX&_:R=L'HC(.Z -
PZT/S*<![->!T\'B6:/XH$P7L2_IVC1@&0)8M@N/C.0U,CEZB=C8RO8FN/@C58ZJ'
PJ86Q&:A+_-5*=96C*XE]9+IQQT'0%:<:3TO+48B"_+5KX:IZI3$Z,II,HIG9"!3K
PW>2\\M<($[A('G.#,5X392\S,$S'MP<>OD$0&@8INTD&:^20);O$Y[F/Z"<18K10
P_?.NO9^,"[Q8[B ^Z@<VY7K"KMWK(N!X65)@=#> 2$BQ8[0^_%LT9"/T^V%%@YA.
PRXGF"*?DH':3%^%8.4^C:N!PGG6>%S!Z'K<? 9,S^:([L!P^!4U8(E=C?,DFN_DN
P+9>AVFN= 8])FUNC4?V1IN%A5V1]UR<W\X!%NLY'Q_)I^()5:#>6 011^\Y.#CX3
PZ]C&)"TC)XK]:#.G:LT36Q>#WNE?!)F&NZT^M7/U-(@'#$"L778*UF&B/_3@DG#H
P.HE1RZSKR(/E_6%G@GOT>*WOU_1(\MBC4F3HN[+OGCS?DGB/^3X*V;KB&WF9U7KY
P(![/>U,G5_SJVS*2WZ3R$8P2D#6:OO*8I56I_IAH;#C\@78^?WI-=(DM#;16K';0
PX#TN!0J&V=*RK<</I@K<>/)(#Z#*?:6H :__ZHX@7HJQ_SKUSPRO&O ]4#F<8Y =
PP46%SN+N1N>EEQ12,A/ [\R8[UG-$?J3K7Q(':F^U5Z\(<NC*^ ]=]2R!M^@B0O$
P1C@'4'7,OYUKV&5YO%]@)BY[M)/%EKFDTNQG$MW,2M3O$6'L$\-H#%,D>(3TT<U8
PN?T]FT5Z33X5L(3-H3PK-6=(^Q>412G*GAN5$J416+DW^NTT)W\8>'3:"C$??)"5
PH"9W5-O<G9M\0V;25824FLT6TK0XZGV5$J-!T[2\OQXTXP']TQ#JD8)+F)6PBU_O
PF82+^=?=*IM;QEL+#O.Y5\PV=*O8C [A9 ]?NM;0I#C%=_6?4+M@E@XO:+3X5ACS
PB\],T-7H?EM(H,!N9[ '9MN1>']M:XG-0YCD:L#)Z1EYD%(39M;8?W([1$L_8^)F
PN5*4&!56\KV[3.4]^L35\+5)<1*T)J%/80\1PJP7L-OI\#<QL!V>-W::N2F @!+U
P)P(TSV8;D#F]01_,)W7W*K<(D7V6+(:KP]/=C3OD <[EX-#'2!;R[XT9SZ7?U&KC
PY,TG+"X;/VJFR,#' ,^@WU_&Z_L++M;F)FD1"]\YH4.X'%DY>)$U72X9\YXGC[G:
P=,*)N(U<2"88'K%9T-2*+$T1UKZV&"'A^JE$@N:4F\Z3?4$.CN[P^'A$P8&U<*,H
PB=YLS)K7. U>FEC<Y"+_D!.X/<L(];%A ?ZY/0097R49%SDR/7^]_+*L12U*HN\_
P^K_KTI/FCM.([_3<%B^<9A"@6#(FK>PLX<(U$22B,AEL#OP1@[J?J!;$L9YL^'S;
P7CHA4MG#WEDN%CLE):MRW\*"4#K@$17B>P'4W%^.7?A (&!PFM(%A4U0NN@6VZTJ
P4G\;B'DNLY$B17L\@B)M<I3Q9(H=4?%GZ$2&_&CRO%<GLWC'0-B#T4U!NL,VS$L^
P_Z([W<BY:LPYK@,-H:K.,FF,'/L?RR1"A\*_G_%?&XP2@M%U0&;=(=LX.0R(3'A9
PGP&TT8H''-+H%7^< GQYCV;EAQ!;YB+@;=-[=[&)"[]\(H.TYV7F#I']$UC;!6?S
P:9LC JI\GO2S%;<Y77:<Z,@=)^;4K\[J1/)>,>=7WM))%Z=)GQ@@7Y@L4.42TY\?
P?Z-SX6P&=="OX.O-7WO=>N"1R""%@-^3-MME95=:I;?6Y5$B6/F46T[&Q#>RZXA@
P$]2 GOZJ6M:T!\EZ(?-%.;!K4(9(B<LXC_QLNBTDP9"85<)P/O>=!C8V6+;2%(@9
PK>RM";5_A>Y;<KKSM.!P'9J-:P,_[AX,N^0N?1@!'$JKV8S2M_%_F7?9XW=!&>./
PM2=-<+.SUMILG$^@$\KT- 7Y3M54DQFZ0;(J(+X@=?;AN%6SUT=BW'M,R_.&ZW5^
P618O-QXZD#F7X^>!YW#QZA](V'M$HT](.2I036Y1I-G!&"MN<EP!UW-94(C#.9W>
PO:WVL/5U!#*  3M,]N4^B9OIH64>#V<D];B0JFZ&#6NJ)YRC@6D4D_TS<GX[)\/0
P8TA\(PSPE<?W B*E3MCIB)WD!1GZ(SK1<S&\<X,74_=209*9^H 1GZ$(-WPC9DAT
PS=1%&QB]I^53_/?S1I#HWO'HT&X6<ZF-Q\PC0_+T\@QQL=N]9WI='V./]8RJ5NDQ
P(-*XI">1$A$J__%X"THH!*@@,-:U"DAV]RQ4K9,-_^V:H+D3Z-]=D,E;+SR%TCP?
P],UDB9$798WVD'Y)[/$?6K;95K"#RBW6N\10Q<N&<2R=V6ZC'N^Q,<D1=HK\Q--9
P!(XG.TC5ZAK?;]+?='6E%WD"6>'&/Q-B+N*YA4Q !^3&X@-9@CW,X#)5)B;[K]NR
PUXEHL%!<XLH+>AP/H#@7]X[^I&A"9*3RQ+NXR-<L!STF"08]*-B3'V&#QBF&QB0D
P+D7J/MO"]5;"\'*A(/+N*=+_\Q6=L_9=(RP'W5)?H:] 6A3K_'$E4Y<S@&9'SF>D
P9-Z3F=66[*3,B @]D7B5*@P6BZM!<'?4A*S%1[GCJ)R\%O8(!"I#=%YOHS40I<=P
PY+9(E+]WH4$B*Q3;1]_*C;GDF9#XPWSEGIK<1E@#,]9/#4-GQOF#BNZS[=X6C'S(
P!+-[8Q*;_QYWHH+=%UPU_V114LM1#NW/,#)P:8L?9F339<ID-.4P?K_-*,>J<-+'
PV8-I*[7CTV6Y2-.KZCGW^*&QHN+X]\+=)6[FBEO[$D+G7"&@>*=^45:#H7@CD>C.
P L/0H[")F/RG&=+D*U6Y^YK=B)>NS5V5%_W?JV%5\T%KN6_64=0R@/.[UK*"1L!:
PDYI_Q4X6IDJD^L?Y9,S9O8I3+'3Y,O.)>!7U7[^UF"9<.VH(=M8W/;Q#Z45B8DIE
P_Z:HDXSA/NT#?0HMZJ*Y^O4PQ[#;12XPGF_ZUUX]@;;I<7D?NP5OO7(\G4TE?&S7
P"AH#8;>YO6(B..I"KB[D:H,+I<)EH+FH+?6/@T:=&'DX025JP&(U1^3>@_.H+# <
PIIA^2R&"ZJN2LSVR&"R-&$."V%"&>G6V<XV7""-A2R7;UT.(O -$8&L]YG2/N$,E
P&:?JU]^R\-ZP=\U3!1'XM//05'[!VRM%&T3A@[D3?3"G+5=M/2_:S5=5#J[1$8%<
P+/7R7N69'<G:G)*L.PH&/#P0-^<C^#<!VAA+#US9^JW/4MA$ MW%$./[!WC*M5.-
P^\_:JDYZ;2^C$X!T XA ..^X\W,KV')&M9A?2D3WP>^FH2%K!V15KR)& K]A[9B'
P]/2K(C5UQ(*^5XU6@'RP>"J:#ZUVI32F-]Q4:AY/@&;'%,J/'CV,"XHMXUW$!H=O
P3M&ZI<\PZ+R(SZ@$L<E+_=CFS_'L13C)1V ^CW)#<PG*>^&Z_1VOX>5N4+%@'HD4
PPI4:Z_FT/.100!TE?@2P#[;D2WZOA&[E9.=<5*9Y=?19+$O_\A_M7H(3>^EV0J(-
PRI4_A<CIC]Y//+BU0/XN4'I$\/%FN%\26RE>B:&)0LAZ-*[=.B%V\#:TR ]ZB)WG
P-Q1P(=OB>(W?P-WA24F9>R6N)6_/+LPZ^Q;0+,?$JUA@][W0XZ\%MLB^*F$,=D:8
P[-5FCTC20D;D^J%4IW4:NT5;6?7B6SVJT0,YJS</1LS"#(Y+; >0!ZXC SBN]$LA
PZT!S4#RG,Q'/^>P>VL>,BW4G-@BC+ON$P/!)#_6THW\>=BDG!S&"JO(0 O6O,B!*
PAR!6L 50;O>L&R(?@F*GG<$+7LU 1SO2,2AOJ<H!'<M+QIU\<8L>"?HVVC/1+1K)
PLYAS4+<^LLLV_V5]N,IVH#"#*BK LYMJ?Y&F[Y6>VLLF;"F/IO0.%"-Y1]V]?08"
P"1B%:;0V_Q&C=&[\R$F840,,0%#J16:>4_7,0,#'=2!3=VQ5SR=N)IB8'%%>FU\9
P<U.I87PP! *W^VX"*E,QS+ZHFH)Z3CUPW#RQ#J-\':!%-02,0:H0.$U\:>G _C+-
PMJN&=.(.-.?1U_"^<C).I_CNW..\=2))C4$V?ZL42%%G])07ON8F?BE-6:L%Z<]\
P?&N@S"[KP]B(R[:)+72*LY&WYW\M9K"U+(M4P L>5JT)M=7FD\+;:2S'B4+L_-*S
PB9"TM>;R@+)T4)/$BKSQT?*'SJXI#>$& N]FJ)??NA'#81 DYS_R>.@-#ZP;;)WM
P?,^:Y2Y1>W'G&R3#&^%MB8I)-7P/-A?H#7>&MCL20+_+Y>./N4C+YQTL\,0Q_1M^
PY6S,X1_AQP6CA65P]UXGCA0XG[<E-;G*'<( -7S8-M[P%4V."F6.L-K C"'WK) E
P>I79B1U \XE'$+?)L%=S3+(UAB8*@HM@(9#Z?R U*L15W!V[MK8?Q5-_ ((#E338
PXQ++F6I;)U?JJ]:0C]PS(J,+5OWFB-W[+$.5F!\XZ-N8"0S[N@:R8WYHTN8(@3E[
POKP8N\)-002,!"Z1H]\/ TYQ'CK,*]#&XDX>FCG.2J]IZ6)LE6+X#UL^$8+:$Q1C
P(Z$NU.2!?D0L-MQV2N PXTL'?.'8^>G,G+ I;-W89JMD9<;4L5Q<'4[G41TR9LEQ
P!EQ?C-5!R719:U!\XSX@L,$/N'*99]/E+PTHBO(@%36$#8(-G_E]]URE13FZ41VP
P=&L3-MYGE^"]?^NS!B\9\F-<M!(S3T@V\NJ%8\[UQ;IUVZKDMN(S6MS6P .XZ/R.
PIX$UBP_I9T/P);_C_RVS!ECO+SSD@WAUND[B*:U7$BCVV:?R@6CFZ^*61_AEW%->
P2%](G,6,$QO:\86VXF;!2->0#PF.AT@NB1@GW-MS@O!/3%S\/DJ4-)9@<QBI+1SE
P=%):*RE57 U5FN%6?3IFQ[P5%$.?]Q.],0CQ"-8X65Z&J'@K=J$UO'^J!_!RRJ?9
P)CJE@&^Y<1Z>=_]C"#4V)I1!MBVJ2X'/*U3^337FC M"3[1U]!:<L($4'J^ D_@X
PO+2,O(SN?S[:2?MW88AU3%5*W6I&&Q%C2NQD-"@-0#F+G8-'>B)N/52WUN6C@I6Y
P[H6%LSR<GC)784.ER!J*\*SK4?*A,8R[P#H&0T,--XNC0Q%D+^/\WL!SH^ZZ$AA;
P;[G[K-A;20I[:4JNB2JRFRJU!V5G17USLC=.)O^"\AW_RZ\76''N(HO$IJFHG%G?
P^0H,HD088LBHRZ4)YZH;_%94JGK%&"=*37#/)V^D<<GN1--L!%?L2D3DCI?%LJ.@
PZ]Q.8VC+F:T<+QOJX75Z:ROI\MF-!!)4158N*"9;VX9[&#R1D;83PF@:)@#!K3"!
P;7&,\L0EB+.],QU'8R?[P,'=,J'Y[>;T(;)S"?V037H5A#.XHDY&*NCECSAN 5?:
P%"+S.7HQOKIRNZCTDYVU DA:J;XPZ#34#JZW !6@"/'WR2'%<,C[_F*]K@-/9R)V
P#EJ@"^+4($[0]<4;<W-=@?F[2+7P\HO8]]F R\1G:' QSZ@:#(L_M6R!/;/DE(21
PCKQYCO- 9@#"^@>93,:.1"_TP-CO4%B@2UF4]\>%VNNE,-N6#TU9S;967G'9 4+5
PYO#EC!G5!B)!I[8=;\L"9/BN3%X/VK%(YP2^HY ,<3R?4;]Y@WK6IX2]]2%=& $R
P0;7EO+Z2TWU9>K%FY"3)2)@%V7YOV-JYT[:*^L9TLM31!X!W8<-\0(DSOEB>(Q Z
P@S$(.@UW1Y>?IN:/2?HD$7TF+U1)(1;S%Y[%T;0_3X5/WNR_]BZEEFP]X=*W&K'#
P6^,F17"(7H;%JM1HDY=2&]7&R'[D(87@1-*=US)8Z6WK@B0WCH*,G [CT6S2V.DB
PI[6V45E()T$;?I6,(% &-7/@19]V:.FV6+K,\#]/:&:W[*U 0'2H?T?,8/971WUP
P^K[\37ZW5 "F>V0)DCVE72XL]?[]IOGI"'^&0AY'5[@,U?VI_;A[1U:60"^%W/*H
P\6/7FA([LB94W%><O_#/%>'*TL =D_5-\;%B-5+&/[:^]O'$XMC=RH61XWUAD<=7
P$B,KUD%S3)W),5^YS)^%@YU/\&EYV?UX]$[\.3O$S+<<E!=B6OE8WS$A2"L<_$+R
PYDOK%,[E"[0Q:27Q=56V3<LG!1">JJ7\0K>MDOW::K- LA<ES6AX!Y+:5O(ZL',V
P0FJ+L<'7$MQ[F<=QQ:Y8,L<]RNPI.IQ@*K3-8W];;)Q3<,!H(5<:>495.%]OR?K9
PZ0DP6J ?>5HAZ2'ZW&[K]@<-5,SARL!/4WPQNQ9*[8YY_+/LF>ASY<?R6H!/P=6B
PN7)[-=WG"DIHRUL@<]OWXO#5+/LNX&7N-<F_0RH@L#.(U+!5*!L^B7,N;N"-BXG1
PACB3::^!;"4[= *[Z]8[X6$' (+W2R@MI*,$+,:G?(?=, $W]PC^6"H/U#BPU%,"
PZ1XANH-,DLIH2C#5"&*_*(6^%(/&E7+_@<SC90.4=S:%P^D6',2(AKC:-\%?2?G]
PBF IKU8;EF";<\SF[0VCV.@_/LK2UHL:C ?F"\'IHQUY:GI=;$7?=PZ^@T<8KOKA
P%(_CZI>_TD-6?J=Q[]<Y.K%'4#!%R'8BP2F<%W70.0AQ00R_+3H]/MF=7'!42%J7
P&69+0=0VI2&=RVUIXM#2%-LX8Z8 &-6P2R-]M9U<35]CYL'*IL@WV<+[MDOZF:LV
PVO\^2018R[6NV/2:/%&LFJBH(=%J&M>5@<DFL,.F\)39TL"L+["]Z9$6M2GQ&A<A
P:GO2,DR)! ZU!52\VH'!&' -@[I2Z,3NJ*>*?SBIH8C\PYYPV_>M-G_C&L"IST@%
PC"Q"TII^0OQ(XZ ;9#]BU)-):UP(*8MR]CI[-Z_3>]VTYCA]Q@FMHQX+DUI[+5LL
PV\_?6$]M7I;3YSI3.GD^K%0:WQJV#>E8.WSD!H5:>/"H3:G@NQ. YNGV@9-^"V-#
P310S6$X( PHIJ& 5Y8(9DF'C;WYH3!N,= \]=@44'6OYXDK+TL87E]0T'"]<[N&K
PHBL$1C>!83E;(!WX+RQ[IZ>7%]9NMME62.5PLTZA,1;[G2(&E?)A84/H-,0!_4WA
PU_!.!S-X=44_+W_V)Z^TP)=U3/OTE0N]JX[?QLS)?VCBZ2A "I-2J\K&K%IPYU)G
P3V8S2HVSJ)K%.']SK<:N'PQ>HK2$SE\\!@,*P0KLI<%FC+DX9N7-'V=[8- 3 /?"
PNN-OZ4X\I(BUX][=95Y)-+#B";P"5BP"P3L4M,/&N.<JH,;"\(.XN1SI9>+_US9?
PFT^-D0I ;>^EW3;D J,:K5M9;/TL2;/Q\QI[@%A39?TU1H$+Q4CN?XS@(1TZI5*J
PE$7/[!J4+SGUTHS,M2[6I<51R<  (3N%P"1H!!4D=F=OA<*HD+]G-/]EOV!<IF$+
P:W2Z[FP2C58LVX8L0G%:NB&Z@>O^*K ]7-]XN'$#DW-7*??=(4"^=U9L!L,\H1<2
PPP,5NWWX^V3CR7-LB7L$ P(X"F1GF^&3'O[$2(Y3V'$RGC29^LH=0OQEG.\@#@^M
P@H;T4^M<+9'TQH&,>$A NMC_#GPF&O*L?(Z6CWL*YWS,B*\L&H ,2%AFRF&MY L6
PQ>PY\G=)=P"JA$[Q&7K8^=IHK+D]*QP[=\4Q!O54GI$05V)-#$^1C: 7UBC]2Z@_
P7\#:*K*R(Z'NOMGR.,T1YYGRLHGI4T L5TADVQAW?6,D#6OJSA<][@/#F$05\U/0
P"X[D6]$U'< AX,L0WX!EAZ*:GG4L=:J(KU4O]+5UJ'KL2W8@1Y_@5\N]+ P&4'G<
PZ]MD+'<'ZN7E9BOUIU/F"EY!_RT B9VF !O\\G&+#^I)"C<DG _!V^BE)*W=4+'V
P1.;;,S%8+QT[&?;A_9TW*O:Z!=?<DIUU,5YL7U5T1J2D2.N.TN#0?\V;C!8KWVE(
PJ[F'OU2+3P01?P6.CL^Y9,)"&@]S^+@!VAN>V$#V^><VFP<,FBC[!0_1R257*>[[
PQAN$=X6:P8;V-@I@V=IM' GD0,/^"%XF5ZEL_J" V0R'O,C&A_, =(ZPT-'T  K$
P9$XS, E1*$=GKO]2;1F&(%-FS;CT+Z_M #R6R+D3(GB-B]39"/T>WH>N]G"-%"XZ
P\ R+.JF(MYA$-!5NP0JL=%<=/DM[*OPFU9?7&+&KG]$1R*C$&JH%9Z\HY$67/KH*
P16H&#M?'OVNEX$!4&F ?QV7NI0 .Y2I:Y_Y9R,4^GQ2H2R)OF=2.W,[3*K"PNIQ^
PA3TON*R'_<;@:J64SZJHL9'<#T!GBDZ8YU(S_W$L6D)WW16.FSP.SCD7TA;V%G*!
P\#,W6I_B]@();C["J3JY'!%%<SL.X8]S_/#GA8R$$2LCJR%[IEA#TZ<G&E^-0$)]
PS75\7IGG1_72FGOJ1.2=:"R<C:8#WL+;Y>V,JRUQ=:Y8C$?].$%/",)K3'NJ)OQ6
PB8XB<)\7S?<M/2]Z24U2(!(LN0-8Y;3Y=H.'K\3"@FL>K,'RZ!P0WW''%QMJ-.&<
PAVCU5*9+-CH9B@H@AQ;'.&MU$/ FC?!@FIK:'^+M%X+!>:2 O)B5[._(MYI9# B(
P%3Z-F3XX#D*M2M=G/&):,7\09-C[4HNAZ4!+E_\7 [OC>>L^H@P/>?L"ZCO0H OL
P2Q5O2HD8K'HA=?R0O!+#1BT*[Q4Z*<\BT0.J TW:1L=!$D$FN?T]!T57GW_= &QR
PR/F<+?!?,;<>7NXU>P8XIW@[!98-\GEHG)>^2[%)(6B!A#]Y_PH.8X&S$H#^6CO0
P'W^&B(1*+'#ZQ"-B=RD6JM12,2Z2@IMD4[R:(<2M8<*S6'J<(TU[RN;W(0&MMCN7
P*27X (T_DWK:-RI#>XGF 8#S8S=4UC1#E(8G%<_-"W6GO]XJ/?%M&[%Z0^:L!2LN
PX\C1FQ=_?30&VHW4Q JD3TRMC.E>>L'@W!1B0H[?^Q,$[J_<;LPAB!:JM8TY@KM+
P"5)HD/^FO<Y>H*6:\?Y,ZS/_JNCZVWEGCQ\0Q;K[UK=W:*V@E#*U]@ZP(<"GM_G]
PM1YXM:432V+/Z!:X-;OY/&(E9?%2)=M5]G"5"71-@H_"V&:DIU'4HK/&1#2W:;KX
P=AW;AI0 J,MCO!D("0I'[ZK5G,?4VA0]<\PMT>=6&4S#7*A:6"R<O4>4T;-Z]<.8
P+P>4XM"2VK0,F J+7&,["*G;]<T0VB*H&:#D=&5/A/YGCE?XLA8" G-/M5?\+<5@
PP(AC) *CXYC.HN10 %I"#K^QP"0"DFM0K.?]<\A:*&O3O3.CA,:=1<WJ_@M]E&#7
P:VK,9F&XY2;"PA4\#9+2GSZ8!).LBGIAAXP!O@U[>\2,\\[?.?O,>%#.(**1Q,^2
P="BF6(\R&Y+(&=TC.SOD@,/^[%[LY*5:-M.;MQMK1N*#7;_*F-LTRPDQK?/%BI/ 
PPEQ-H-H/ /-N;MBY/=?<DY%,2+ [B!:3OEY1R-/-W;W1*Q*\B76],=JKFI-4_G'$
P72A*RPS1 \%:NGB+0I-,DG(?M+X<8ILT&--^]=UC761NZ_WCP<0.U'$_7=R$=CHO
P/>4$? ?5#Q?EO7!WZY\4\V[+FP36EW]$%<@@.OO?3$NE*Y6-R.TQC?)'!];+[_ #
PO0QFUO"F2?EEHG):& WBR@N1K#MHK!0[,!N\X-/-2SG?DL\*"#RFMB0,.<9324O-
P@A^ ('B)KXQ/HV;^&Q85*99D:U%_$PS?^7-4EF4BW84!'BV5[*<S!R56J )8M0XL
PE)2P[3S,.D\+"Z6ILN6*3.#UF*/#%AB)8JS:^+,=(E75-_#D>=@ V*W")XLY,KO3
P""TA"56W3P"S8K!+\.9M%>;*R0/ZGY/ZSI.0&7FP@T36:A$RC2-U*I219Q;>\_W"
P[8*!')T,2J9/U(CP5>:"MK]7Z1B.]+PUVY:1:\]3(@RVK"(U*#KVG=.U.'%R)CM'
P8P^7WW0G>4;WHW&#>@]"BJ^,+#Z;^26HKAF; 7/1.9P)'<[DAT)64=!P\.>U8'LS
PCK7X'^_C '&I#TR\TE&.0Y1(*VRBHTM!B GPF)Y8+$R7 LH/3L*P;I?5%8 BA'^!
P1O00BXW747D%@UAR'?H6XZU_T]XM9[BF.8.:?J8"X] J"*IQ"NF]VH3TMT@JPU!B
P?]G#/CZ.RT*QZP'51/V)>WW7DRNS>U%X,L4/^L+^^2D*8$ 3U^NMV&DO,#Q&**L#
P[TNE]>7O/)]:K1K54P]/[3*J,&% LZ6Z (Q,4?I;P+SE:L1TT5P<Y:,6N)!PF]3!
P:TA"[+#B*ZGX V-=-%E,)M(RL']5Z9*Z"H;ZA%^+YU^_:)^2HL6IW;]CO/F<3PNA
P5_'?X*D2@C7:A\J'KHAL541\ZKFI,)\HD@OD&,5#C^WJRM_8?C7&DSS01!G(#)<V
P) Z3!]'>*Q+70'AOV+&9Y_STC>[_N3.72),%B[JG09WK=RN%S[UO+PK6Y[BC$E#P
PET'WF.S%QFG+V-2XTO:7)(!O]@107"?I7L^C/37(\%D;9=TM<?E28@&1L1C0 )5J
P$$O\ YS;F7]NBKX,DXNFG&3F8_NZ9F# 7J%VN\H7M(L%6ADAV%,-X'42R6B1\ZF)
PU 3Y)G(O6]+UH)W)Q$PS)*(EK/N<GB!"1J-;)X2LC<93;(S>8ME:BS)1.!"-068T
P-&/3VRR7]GQYBX$47<+ :5U;#J@.GK/ZV5%C(!0,[5$VBU-S*3<VF8GQM[M_7".O
P?28XBB_Q?1 0MRVO%O(>&18/]ZL4AQ#7*I2IC!DE(&D2LFWDG%![CRSKLZ+4*,EW
PLN/&CW9&VP_PKU/H 6T^[^YY!L-^7C<=@7*)5ZAT=8>PP[GMO8I$N,!]+C1RX!I,
PM@$0)/F=V[2-8+O66B[DEAXW1[DAI%I9^;9E?J0!E!-LG!(1G60J36+TRNRVH GY
P5/(!FJW^VI7Z7QQ:N$/@&5QH?'5T_OY%SZ/J0&D?V 3/J+&;/LGWM-YCZ0!U/NEJ
P*I>L]4^!-W#9U7QYW1T3X>BL(*H&,.W!W0OY15*!-=/Q/877<05N9/U%QTGJUIBY
P:"P$7UKMJFXKZG<%->O 04/%_&D&+I=<J($Y?)2.W@'4')Z; X)-A&C6D_K4NT-!
P^4</H;(G3V]JX$$PB"K;:IUV\W/8%3A8Q1A".!,0LB?3XYVGR3PVYOUQ[O0IK"B#
PG0%@9 %?[0W4?J+%66G@?ONF@-AZ-7T-6S.3(?/I^(4KO>W[);4^5BXN>-@,\*JE
P.C4#X6*#]YTV%2#@./T*AVD6S8G24CN>X%/O0#JJO!59// //$AD:#D*!!;9C8S0
PFF+CFY&[=F\M)X/2L&6R,]LMB^,0/@;]'$!ICI!'Z/;RICIS$S3>O%:'9BK9,5[-
P7)EM+TY4T>4#R,LXM[G<19PT1*]"YS>;'DRP:-:43-D3U-'RCK%6Z4N8 K3/%1<F
P6M>Q-V"LH-D/4W)O6&]@JK'W/>[G@ 8+PYWE%O;IVO%LZ5'L:W"L^4;E90%7ZO1B
P& 8^3<!GGI^Z$T]3(6])WE8;]V7DH==1&]O7R5?@B4-4WPP=3Q#<O$ECNJX>)^=%
PG;HOOCMT6C1G0+QMZQ-SNY:R[YU6S>_9MLO9-VHRQ%<>"D%&Z/.2P 1 ,%IX?[,T
PH2!,XW]^./>3RNVE2\]$+7#*5M='.&5#F%=I&A&N%'-1F*X/ /AM!6VRLA5+%]OR
P@G!E(M7FP%V+G2IWLYKAZ1(A<^^OA)]*-.OT<*N'TH@@31YP10.@-'0B8G4_A>MC
PBEP&:FN.0:W@?DEXJO6HFW%-.59JI*JO0%)K@:PN$)#N-!&^:K#J"/O"MX4@#:"%
P<+AB/86H_$*2YOICG;[%W\4QB5#<:?OPD.O[]F(-P0CZ_]'%I1PN[9GC*VNQ6$NJ
PHXT'KW*R"P G]'4!<VBFM!D2-J&+:A>[Z/!0/=1+W/DUX'HD\O4>NQD;&6_)E@U$
PY*:+K,;!X2^#"#C!&<))5 ;J[A7SS\<27=+:'B;P"'N?).61BG6HQW*V*J+7Z?I:
PRYGCW+*W95C:Y61[=FPZJB$\ES=+D,;6J0D?;59,T@&<U*:SF#&;5Y+W$G8R* %G
P+ XD3Q>UO(_*-F^VM*0>@;KUXA#H:FTO^E/]6#\TP_/#279U"F'#DT;RGD-U1:2(
P:KU';+EW8QY3.SLP"% MWS^&4;76BN<0V3'Z*+'99+A9"0X[/S^"YE95T*B;(;UF
PN)Q"W=P-# 5?E0H5#K&B,O&P(PTI4+W6=?S14;8BN:J?\Y1TS(=;XFAED$,?7:9%
P0; +DTI,[1,,A\>]2&Q%')\MY@*Y'%F=XI9XO3MNZKW/1%\ZXJK%"N21*<LW^#  
P7II;*/DS^G> M/1^AS.7[WOZW]DSS*C)S:K*&C$C@JW,Z)<M)O#<M+3=65\!\0@=
P=Z/Z%[+TN'6]5#FPNB+D4I/0[!5'UURNSZDLK'B<-Y8(%F9)1]CDB@0?/'2D0B@%
PW):+&QL6<7PT.4$)ECN?<8'%#>8A<:]& BQD;U&@;:@LL!34;)]G+X@+&4J"C0WL
PE/!0VGPR'0>IZ6,+=DJ.%$0P"_\*-/$?G2^K7,@ _8]M>*+:7;;]<G2IVA'#AW($
PQ?E;"5=(8E]]%[[%K (165UI2RUH97MT0P#\W272-DE.DUOX_U[Y9,PX3HF[7C9D
PZQ*GHU$5R\]BI[ !Z8AO38:1?1]58)&>_*%RF="0R'X T_X5@'%^\(B2_U@#[#HL
PL 1A+H.VW_;41.?KE._P8/S8(:1,5,CVE?6!%MWTO2^Q(7U_ZC;:S>7=O<?K7I4*
P**HEP+6*\=")''97I@4C%-GJM%S!1CKE!]" XDX8$C:A?\WNG@=F2^_" 2H_7*EZ
PZ!=P-)R-OVHF%@QPL+D^UEUP,NQ9]=*!9]#0!V]4Y%AIG@=?1WLOHMZN;<G>3Q@J
PI:&SM_74I^H55G3'2*A2^N]3[EG*^$))9%^@!),J<EA:AY!(4@,.IW<(43\IZ$P1
PJQ)^.]L?5?'!0C8B)?XMHBE"^KSL(/,E(3W[B^9@B7/^&6@-$ ^3:+Y$EJ#)NU[;
P=V[FWB98LJ:EU]+#GG"UP/SLEBOJ_QW'J*/88IG(T0JEYB]=/(!BU2G7*>(-7Y'%
P$+?D4;3NS9-5.;35'6*<W<AE'5ERM#0OPS4@1#P1"_3WJ(X]C (V[<KSY*=*C 3R
P);/$HQ6Q!Y*:N^+C>6"O0/$185L\ #S<N[GG\\6*N00"<2&&Q'Q*$5TM@CH6A08C
PSFYFNBYT^7KENF?0K:=4-5HBYK=1VMD$CZ(&RH.:\Z%7@T?+XJ=!+AZ*<NM4Y@7,
PK>/*XP:G/MXOI( 21F/_M1[K<X$#UHO;;?@)<U#_\U^^>6:!Q4T I[5BR5WM7;L/
P-NCM76CKI! ' ;#8V,3P?F1SQA*]JIOU4F59,&SRKT-R'"]\KU1#"QWM<8IK/KDI
PR!4>5BT+\/^(R%9D65KJ#5"8/ZZ/>]MS:UQE"Q*GTO&DI5@^RH.OWC3)9>'F+!/I
PX;: T&L;!%Z?:'M0>%F&6^UU"$S/J(+S+]:&:Z'EDJ3IS2Z@*1I[LGRAP) ]IJQH
P8%1=9=6'9:/8NMF/!\J+.\UB#UW\3$)$DF:NFD60,.+Z_?N!2J13&1 _I#PG6: .
PA96K/[V%_URCSJ_%A%?$7\>:!_"VB)CE5]XNU"%>TW$S0LK?5/)(!0?D6N!H-_H]
P'ALE*S!8U2=W)J5@R=[K,EL=M.#JF3P7Z%,%/-!A(QP]9")VBI&*T\K +98?%IP'
PP0YU/7M\*YDHQ:6[>1OO#(*P$37K+H0#<^#VGG,/?5?:8,KK:\Q5AX!5F!> ,6XD
P9U%%UM &-;9FP,F)BB=C]]Q\Z:N'1-,$>H\?BB/)@[T HU"TC*^(K5-B3\>O3H\+
PQSDNEL\>6^TK+\2"NR+N#LLC)Q9<&7DAT<%T4J$R0UQQ;[C[0.: -<]C_WR]HE$&
P]+NY MO5,-<925> KZLC1#M?UR].UN5<SQ:^GU9DROOW!AL "A(N.P#I@WKU&_WO
PIC+4'%+L/,+2W/@*TA =S)4.0VWP7IS>JFXI>GR84MM_KV1X9>/ET/G^_&<4?4> 
PQCPLF4INVYB6@6CW0;GPQB-)0JL"[VOY "[H;=-+#EI7D[\]">)I;1#Y!DP9@]UB
P]J:UK+5W;4*I*B1OD%&T$K70VJAP,'K)TO(XLF1EK6E>.:DK<L,00A%C&%6==33T
PRXL\Y%2.XX,JU/3BB-I7U9*PK!K4!QQ)!45%S1QU!E5-V#+TWH8X%I:A*D3A6E6H
P(@KEU/:T&4EO6N3GO_U@<2>V%W?B<)YW)+HE]$/L#Y8H6V0Z,%G7-TIGW3IF.O*<
P W;M$36O@WP .MGT3 /1-:K!#JF/!9$/LL6##W>B&SQU-SJ4WHB+OWYYSAS3LV-X
PE+G@8&-\M3]GZ1&/_B!3;8^,H<SS*["]W,(EZ%F"&A2E98X4=\U*+5J.H9<@I D1
P&C--5O' %RO23NL4(7\NR>DW'9[2<]X'<*XVP;:F*\\8NNY"!<2NL0OP84TDX.1A
P@(T,QAV*,7U%=Y@2USDCY16K&#>7FC:Z-JK:'+[I)Y1I)DYL>Y",5X!UCYH E"P?
P WM<9&'2[.\ZJ?*V![0@!N0+ZG4 &48-<[;KVDP?IK5DMWS4Z1W4.*'=RT&W('4L
P46]?YGSC3<EBN;10+45HI%=(H7OY30*.%&*@0ESDR9G6F\+UVJ5,/C!C<7#6206_
PI<-*6Z\AZWS%=<:NE5+\<-$:^_M!U9LR"2@$WOC\"A/<]@5+Z*66/.V 0,4%66MM
P;.7[!_@O^D;7#;HY[,YL_S'\G@$03.1_^)+6&;.@3<W%G4.597Z I(4R5$U+@BTG
PP S]\V+=1<"JB41U^50(E:[Z6Y:0:]"HW)./2E^X23>8I\I9T'2]>QEFOL>]X$C2
PG1@(]T]HE?A0 U]5'K_[_BDY/J$:.,>(:!^_=ZNSWK_U'&*WT 9YE=7=AW-F\+OY
P1*1.FZDL.M+S]8+7Z0J[)$'L8K8AH?RSM \GDF'Y2!4*WP,*!;A('M1"B6<3AHQ]
P'!E46XB/E6/J6U=CFPYCE]ZO?:I#<NN'$=6 RKZ'%4[,5LP!,:\VK207$P=6$XG8
P8/27<<822K \@M$)51S/;GB)P2)PF8X+$W\=P$[%V]L,PJ":P;(?WA'BGQHL#T&U
P+GXTRO;:__^<G2&SR^(- *"(-_@A056>5'5\)J,2'D9T=\#?K^ZG&]=5<Q_LQ5W"
P6I"PGM\>)]NP^#\P-Q2E&C9 &2P'7U3@40BSX4H$EX#DI)4%AH@9@?&F@!AW1U\"
P=%TAC;1_QYGA#@/JG9>*4;:P !.4C+1(Y^3C8/MM91./'SYDE?AW4#>%]M=9S@<X
PSOC S<PC.5E;O_19ZE?P__N>1T*"UHJL^^%N-9]28E_(S=_L<@&=*O%Y!!0>LS3+
P)*22VG.] 9'YJX:T%%N$[X^WB38^%6:H__0@3'XC/E_H+8[PXAG]]!J00R',@[Q.
P$=4P@R-^>+J(-<7=3[Q2%6GZ@K!T)O]+;I)M56WQ;&3505&Y#4Y9.))6?HY3#:G7
P?'(D=JQ$>);#"]/N& U"P4O+:(RA!Z.G2++CI5<8L,F[7'P4H/=QP7]XO3C?N,Z[
PX8@(B%S[NX_O' -*0).)$>RE]#'PC1,O"NBY&3\6 _\*69@FG7E(Y#3\P6^WVZF/
P\7TW#[B(^PMOK>GGA85@6S?&T+;]G ,"?P*&0].H."5%C;JW?XTH RYR1 >1<"<O
PZ!3(--KG3X_W&8#:55D/O&*2!S3XB*G+LC5BY&OH7J#KMTW+X7Y(UT-+U04.T@*@
PUHQCU(5,PN; !1%5!^X1C\D6> -&G]+$_TB83%$+3MFG.XHPI/B2<=] BSWG=IV^
P02QA\V4'>V2T@<T6M.,U+Z(LL%<PUE9G +%;M78,G[DN\#BY,!<B7KGWH$3F2"@$
P<< .8LVD4YQA%QJH",'P25L:AZE9%($Y7303T8\2)E>2?B/R-$Z3!<V^-Y->_O'M
P*S>@'LC[4UV+SB*@\#MK2?[%FN47#-X-#6IUBG>.@+U,I?BZ=('%<\@9$W[K3Y;N
P[$#NG>5>2A5V+]9$213OX4^41UQ @;T9[^3'D?&XH"&),8\?GHU6N@O@Y_\0_F#9
P=K%G%%5<=Y:7S9J1=]G(]<&JS#J7A\XA>BL?I?)R$N>TV=[9[F$SYYPIM_[M2<(\
PX!'H!(G>9=?C[QG([G[-:L#(D:(J>,\[XR*)'SD2-*.ID6!R-JB@*X)3&BD9<0#?
P=S66B=D6J]9=I83X2\R3S$RT/;(7;!U,(_K46AO/EF*CO< %2N1DF0P*3*?]OL)"
P_G\7%[JQO!:EU9N7]Q%&.;F1SN^)&42 W_([K'(VB;;!N@EDT@AQ1"=^1)E4R -^
P%98'=+= 4,*<SY<A7I&2$JG.&A,WW4/!SALKN(<^R]XLCERLF%,B4E,AB).=MGEJ
PC]U60D))C8$&[\5K\T>+' O%VINOU9VMNAP:KUQQ\%"?3K[\XS_]#?([>0RZT^OF
PKY8_H#?T4G;"#:IP_/(Q;H,%=])B5>*]99 A\%K%HA":D6:J2-%$49,;+9RL4LHW
P?S.*\PX-@+@M;MISQ8,R%*7_K7WZK6 &9+HZ,V#=!%#I P\C)7N0.+3P>&&X V)*
P^).W>D:013MZ0[V#(N52LFB!<TT2KU-T+1NEN-,ZR&A[VGS_"9Z&0=!9H_DU)D'_
P]8H#RDXT;\2@-:I8C1,!\__[5D>W\Q;-YYA*56B+^24]VLL @YC+C"@*\7$__EO9
P)WA8N#TCW*#-],Y**]#KZ.-=B$0'?<,0<K%QZJ7P\,G.(]GD;*9+?-PYQVV_@5LV
PRO<&"_<7'Z*5'BIT)Y.^ZM@TL89>!XK::RWKH5[>X4TZ(BI[,A>L7\ 32WOK.?.$
P]=Z;9^W9GSU&L+ DO^2B#TF!B?JV8#?9PT7+29?.1/1C'(((A3[!3#OR?+DV[]3&
PA\J-.A&[P ZIG*A'F0E)_=+?Q&HCHRV4!=UN[.>XBXK=RPS1NA=Q09P9;=4$U\6P
P-Q%1JBR-]G5W@HDI(>O][0MZ2'D3YW.;Z&&![5 197N0Y5Z;Q^=YUDAH7X3'MNN5
PU@PUW[D-0R*\ ?BJ38 )33\51+O[B*1'MBSAG6%IR] QDNOQ(0FHXT8"T \]]YY*
P-](0KXQO+51.V[6/HGK$F5)]&#M_5CH@MI.3(]36K9&7"#4:B>]_"*>K4-*]3]_U
P0CUC&+#'T6C$FA)B1P'M]".V'*>FGJZ2(R4>J5H:%L7LWGBR ,V15_*9TKDNE C*
P(ZI '8J1HC?/ P1K(,LFD<L&F&VF\[!ZE&L.%46"M?) MFF'_9 >QA)=[!8>).$K
PL+[)YI*K:)/9L^F=U]GMG]J7";V3$:V@YR,]0$PK.<R(J6D1J'48=(E6/8X=TJ6U
PQ,R9$?-L7D",#]]3D'P5"GE@0U,UKN2U$!N7$IID4HA!_BSF9M9Z(2>#DD,Z%GI%
P< Y94<,$4H?1F!%)PFNO6]%,G=ST XX2!J3@A>7DAS215:XPQY5L_W3VB"2]1D!8
P6;[(TH:9BMR)Q;/1G9$LT9<7N 8$7XNJ)=QO*C_5@ST*V5"\B7[MH# 4)ZM)<S#S
P4?I_> ZQ44QLETBF>".N!3!:<Q>]1W(/'S#CW</3R@#C1H2CT;[M$C>.EGL(12"=
P+R=S'UU".@-DMK'Y=@2V1>[CCBNSP)S8EU@N V!ZOWPS PDN'2-M!BN1<N=)1J %
P+/3BQ"1ZMB(>%&X$_CM*-^&2.,<OX@L#7.<>:8<92ZSW!RYJYA)?3%HQ-;MB4#]8
PBP5 ,Q1;D(O5$]P><>/?,1TP<$][(BC?1)U+<Q9'O#=(_BPI].^,*'1X?6X&>%DK
PO.+NFVXL>3-$T'':T+!OT0<#\8M<'BQ*X*CL0^\4[=$ JT0 1*4'%]U$Y5I5-X/K
POA&6]1;(N/"&'K@,Z*Y!(N=I\9-M^(CFQ_A9QM^&N0&(\'U*5&8E<G9)+0]V;YO-
P0-X"A!&]0-ZEK;5N4 PI)NZF#AC0=6#;?-^*O1QT9-'-0#'N(/>BR:@)KL]QQSSZ
P.,@[#P(G0HN&,P$LJ!^ _$IN_BC5*XA^&36#Q!OU9<%YV=>(AH^CGFO$3K+Y__ &
PB%<[L?WWG4)!@>5MA\H&0S81]I8:5:":6VP(97;KOC?AOFSXH[.)4/HKCPZ?3Y4!
P_)<SL@=6OY6UUMB2:* 2J.]HKTS&E_^UM8_63,3YQG5>:Z(/$%V7 ;W(H8^8R10H
P9_YP\2B5X5.7 P U#[$%4#[DKG2MJ7:]_#@"02,ERX.N&1)VD#M6V *])^N,VB# 
PV'(^LR#GWXXIX0D_<MU1?4TSIZ #X92MYG\&/RVZ#2+V^B Q&6;)?@$*0J6MNVW>
P6E1[DX [3B6]J_I: ]6X=,JL0M-$N[] W)5_4DNJ"@!ZZAZZ183]G,8QD I;=&^L
PEJ'JZ%;*C()B+W=+SR8RV1B>]ZY6K.(W@H@.!T5O173Z5G<!LHWG[Z5M5+TMYIRU
PO_U\S$,_15Y((V\6^RO_WJRNUFJL-<1ZK:O9>GF4,%O1F1B<_)D^$>T[5V[5+3H'
P,9*G"!FH/\5:Y1L:-.E<2%SU0$Y46.(DU;J_.Q:D2ZX[5;=]!?'8CY_:H<[</E[3
P@G%\;FM[I>?-!PE&()[R[8*Q1J!SRNB1FW[!L&^]BR;LC-GTZXVU.['^;[!%RA)1
P^/ZN;QFN&U)DVU4 ]:Q]UX[L1H.7L';0*,N-)D,5GK,= .60,SIM.ET#$029RVN 
P7X?!D/GLL"G]W&[\/3KU-"\QSAO00AO;EP0+P6O /--!%/]X1FRMZZS,M]*66D82
P7]?0W;X&^"?C<(D9_%.@LR_MS9!I88SZDNYGM8",T9C.WE+0V(NC!.3O8#*7H?MU
PU8-')Q,O*/??*@&0%G$!F::*+JCK4:W^I%%]M\(V"FO[;4KC3R02Z8$+BDF9&_O=
P%\K;U B7)EX7OE6>YT@RVW.Q4IP!6#5"Y><!@C!=A7 YRF@AFW<%1N[]>0^A9*'&
PV7E;4U)0AXS/1U!K=S','C)M(0=169(W'@5* :S?K-6JR'!3)KK)40ZL0"B_/8=M
P<A+&.$-JI:2F[$X<<1441F+V!8-"+%L?_QSED5GKB[5Y[4E0D,S:Z]_95T5SNLA=
P"3*(-1R3$ X:/D)19/L[>]-G/:CS/ZZC[*O#\[)D^)I[O3,!%JY24P,%3*F+93_=
P'P7^PJW3P*.44\ 5I^7EYDY[ XFK"E#'\3J&0CD\+8((B+6CWYU71HBS _G4L*@V
P@!3ZXGA=B*]P;T^ _A6.]']$IK!I!#CWY4[N BF>>I*F7DXN4O33L@5KQG#88^S6
PTO!I5MP$ Q$A_<"\%(S)F5S9&.:I-03LH#5H_#KHNDF=%78\GEB/"OS-BV] S>9(
PHTF1FD+K?)@,>VS!NW;(K90CCV=X$6QI>C+0NB%C;19KB;\![%878:HE&PM3;D-V
P,_>F2E3Q7\PU3^ 1=GXR<O;$O0";KECH18S)IM)12LA=^D%BJS5\O@]@9637T+/H
P<]^SC(/U5+JL9USR"1TP0HI;WDP\./MW.&1,+:\:T$E%3N?SG.XF8C\P6P49W?VI
PC-K4MQ.(F($1:@EN<^>X9*N[S*?Y<.QGM%&(VA@!CJ??N6-ME DCKT:7N[Z^5K81
P1,G;X</VJU#(0+D^V:*L2$>CC=F>/Z-Z,E9RK^UTJW-'\V=E"9^1:_#JPN_ IEOA
P[F&3W<8C<HYV_3]1O4.! KB.<A1BNT,WVR^RQ+4>S#]GMRM5O^N#Q$X*)BHO]JHZ
P4;!EL.EY5D9%M.R=:V<:(OHCVH=, JAMIY#BHY^S_"%%[DJJ3\P3RQK'._O2TQYC
P%J$Y"MVQ@&?(-?P,FN-3"<$,(>*TW66G3F^38S;*K,"L_7U]U/N$0O;3'-;>U\LB
P9"O2X@QJ@S W=_,E;6L\BV G?KF^8&*);A1%T,Y21H!U(4.+; [8''-+4 F-P^JV
PX"B(_E@1<*=139$/\]0C'RMZ/:ZH ULMZKW^D)I?<H3\P]5DMR&',AHGZVA44-=?
PFW:1D+*F 60ARN6\%_=<6&9 Y8$3X=$Z^#3< F9%]_F!8 I@G)4'B0+Z2:N,LOHP
P-6B%]B+5+Y=3/VV3LP][JN^FLU(.&NR!%VVYW6G?+]UXOION&RF@4B"J13^W5DI5
P&U0TH6+SB>JB4O>%7]+!QQY*SOFWFN/6=7"AU9D^X$(WQ<%T%R*'2!XR9-?\I9%8
P1-;UIA250AR.CU*US3+O84$GDMQ5O:7C#-!C2H(Z:.XQA^,$7JY\/Q[+BH8^9!.^
PNGF*.RS:,)DD_&O!X_%@MOL>W.5U.&C4<!0@NJIXA>UO?I+ZIA:[MG,I!QO3C;-Q
P1KE5]R7<]9]'NC4%,#\$DNJHEXX#A??G7912<=XZX#1S__E$PLSO\J P!11W)3AS
P]HOA0PHU)*!K>SN'GC2$GW_M/ODJ=V#SW67?JS2H=9!3*Q95\D_J\W<7<^QG@59:
P&'AO?:/&Q<LSV<46'G0B")_'=1VO+W7(!4VPJ.YX $;57!RK[#F&6Z\RWW8I]L1*
P;*<TKCA\LB+XC6SC^Z5.WU,0SLJ.";- WAK%U\%W:O@QSBIEJ\O'<Q3,E(A. LS<
P>&6<8,^^9/':H_ZF'PZ@<0!YK[U*$:GK6Z0J&G-G4#9!N'Q0Z4&F=E<\-<E/>3+#
P]_K0U%*31"'[W;"V;7CLW7(5EQM-@ X<8_V;6BU'IO\TN(#4>@?Q- UB[)N'P--A
P%080J_*_(V "R\S0<J3*]T;K#<90,H8HDR3ELHNE5WXFQLC%^^DN#9_T@OQPX]8W
PIG"U50ID;S9M%[:P)OQ,.A$WF Y#468B>LV6W N6&]2\H9;"93V+8DO+M;]()C,.
P=*#$E(;?3,K^6&?R"#E[S10DZ2:FM#2YY9L_#E)/\RVQ_H^"J#OHM-ILSV0W%^2V
P!>+Y>4]..3+VN=(\=JK/FS]*R2SK,L;I Y\]Y08FT[6O@#(!2S1:)%,";-TE#]7'
P!2&=M*B+<42-#W?+4P4BK>V*L*; A,XD*FAR:)6O:P%S;L/92AS='TTE"&Q'\7I%
P;FQ3TRE'?,T'^B/Y@,:&4PR=%E/T=(4UC+26 3VQV 3FTTR ]$9P#K!$2G.2''"F
P$*V6EB8,+*[B'"<@B0XDZ5\Q\<?0/O#?BHZ6 D G ?*OQ$,M6$6C;O%@@]$40'E(
PF!@O?SE<TCJ$^##0BDI[]QJQYPM[HZX>#SAE<\U2J>P]<H[XO?1"$%)86\ =;RIZ
PA=O $N:%&6%X")6<-IVMW)#HPB9\[FW]5>DI02CGB-&AK[B![H==DN*(6Q7W0$-^
P7R9PQYFH<YJ<DA.@LC^*P(0)?81Z^0 )[M8-HG^P4>N$?+^B VF*9T,K.YKRO5T5
PUK,*I'4YFH_>V*6!(&";)CR'6Z_XDSJF&S9%KA"5MBM;F*R/?B8L^8?@J8?TX..9
P/FN[> W/. H[ G AW7:_8@Q'$C:PZ$K"D"N221XP,G&B*U?@=96Y;C^R>YSZF7(I
P^SN#];AV;N%_$ J:_</>)@5 9S/_.HF  VY8B10&7>TDU2FPFBV' ;H]EL-7F\%D
P%PI<2&?MF7R X5T)#'[M]-LTO?7T)\+J)P6@L;*-'M$=53JE70%Y^3%)F8P3@X"/
P(86:+DDI" /QS38>3)*]271OA^4VH]?8Z(]OA'0ON$VLP8?_S,9_^KZEYCQISKG=
P:FW7I)Q?F/+_N4S$R5A93G%B;YK'] ! ]?8+Q08EHYB'L%1X/CU68>N%C^?0>-J&
PA:*NK!3PIML[N<K/-6ZA4R(WQF1'>3Z>PUG\' VT2)*+,=WES\0A#%)VYD[VYUHL
P1/:0OE:KI6M$;7+^=>"]^59N5!)R/$2"W0?FF=HSOKBW6KC?LIS5#C7?.J$9H1G@
PF\XY492 !Z[8OXNH[98!/4%'21(-02XV YM_%TBI75 ;@S>I$HIQP'/F<;*^!YV;
P=<*Q3!D;V3B;3!4?#'/ W,=/"@M-<LG]Z,P'?HUH8ANLR8"!]N\P$A<5%SNLE\+"
P(V?'(IE"K_XH]PT1G8%D7*@$!8.+/P_^;%=/L0F0=[@Y?^:J]NU+B=,$Q7<)Q,TF
P=$7">>W $YW&0S_6JQU\-XJX],NEC7@7O>$P(F3+@TX@F(]@,[5M#,4D+ ]^9XU-
P2@DC#T:DA0ST.N62A(ED<2U_3P]U\6R< ]IUO8.E)?LHL"!!]-P#%Y2(F?16 !V6
PT;2YBQ<R3"'G5&46W8P(8AN@^* Z8D7EK.?T@^D#YU P1?=Q[4G_1Z 7'?Z3/[LM
P+T[7PL,4O:\3K,<!#']_X%(,;A<^<7L%#S.WMB><]1DY"O[D_V-M(7V\=PS1FL'V
P5DX2MZNE-26491T;T?(&Y+F/\W^,5B5.#RN9;LI8&1NMI4CO@=Z^[#9*XB7P6>3A
PK@:@JKWS<[;@OB:;W_ ;^LUJU1YS^HK ^6%O6ZB:=/QB4!K*78'*:7AQYS,_'L1M
PQ6A-&<4XCX:;>X[56PK$[33SU:4H_!)'L>>?FYH7BT3DUNAU8S !;UP^!+E8(B=P
P3@LC$)SSNOQ0O<F/8&X<T3W%%G#I;\\W7J^L^YY8>XUD\*__E-"R*C1"1"SBYIQA
P8Q^QZ1L#/=V1-G2"J9F6/QX3JO:T:W%@R'76Z="HPF\59 G<8GP!;K%X-D>G9R*E
PL=H(7231UAFC.V M;&)Q G@9T6MV"6\W.M_Z3*/VC-1I'L"0Q$F5K?.G;"/J0$Z"
P(\>#VK_(P-!)M"]7]D1$!2?5NW>$D4&A=OK<3\C-&^9EN%%SA.)A9J[^\Y>39K.:
P2SWIW*:G,2!;HH NB_LZL%.[^!0;^4<^R0Y1!<DF.MSMU,X$_Q"?"5DZ,B^(\V.C
P"/J=8=E.K7?RH:4T8H918I.OSQV94K [-SJ]&8FSH7T>I$R 0<^0K::EU'8&M3V>
PQ,6UJ2=_#(1M#PE]#$M<YQR]+K:XJ/1AHSUU!X.K E&/<6]NO1)IY>X\VO[SV;3 
PC)E>R0O/\BX Y- S@31[?MMID,03>'5Q5/*;M;5V_S\6<$HO3?S-6QS8$?<;&WMU
PT]90\4-BTG#2/X%'3[',L.-JJ^Q2^#L9EUQL?SLDX!Y_HC*#9IJ0-5F-JPA\.%?O
PI>GZ(:,\\2R1N48&_*9P-!$4+42Y3'9G(PRWZ^=C@$:A\+AU[7KH99"LD[53>+J,
PKX1OQY\H2N&!]2[%'I"$JY;Q>F+>'^O##*WC;N02M3%4I9HR ILTE;%AH;,$+Y#*
P?42*V3+8/)ONCWJ[QZP*.3B243_9ZN!' H93'.4NA661OEE_&T$*3_,X.N$ACF'M
P_[&X'2K% VHQ&&CW/5!M!CY7!3S74@_EGHZJ-UM5V'ZZLGQMVTRHM3:!'B;RP2=9
PG6.S=U3((U^VP*=',^ZL7A(<)G 43OI$ 13'/GER,IBJ0%X=S,+^-K*7"N<YAK>C
PKX%4)A/U+T5OJ1P;M]A;14< 3O*17&^A%^D@+=+V/2U1D,VQB%(0]G:W:PY>^4$P
PYGMH&7^"0:2YV<<RK/3(8ZX<L-=N@C4NCWGBYR>KB'H>F(%S4__99X@8+YPFSMP'
P[II&;:/AND_L.02< 2K874S,Q,?H16HFA8=/G?=+IM!WS[5<TJF]K>M'(^1RE@9E
PB/R/>F'UKAW0BH']="[<F26S";1C+ 8K8.?SW2A^ZD>PV:]1O'&CRJ.A[LK9TGC$
P)>Z43F%"3]E#Z)S[P%G]Y_6%(?,7_]K>961?X8%5<&;0T1N 8_X&@$K"^"8HADC?
P)*<?@JXF&TQX6AU7V0\1'@UG1# OCYJ'(HX!1^-::\@;:B*S *XS1Z<4DCU:/C#G
PX0(+FWIWDB6G$RE+I+VM[D1'_N/D)><N=T>PVTB,#":;]GNV_$VV$MMNWN2(5-_F
P/*(5J"H2Y*8H2-@[SV10J41*IWX%3])O==L1CW0L7>BSES$<[+INV,C0_X=23'U1
PD*!4V,N['>4=+%+4.(4LVRUQU9$9<_?XD0M^"DO*9J!%.%S29KKA#_KKW'33/03G
P"]S8D@,RG;91P(1#>[;;)ZW.PH@4L+9P3-#Q@8$7V<L^VB=](D_,D@GDZR.+"/.Q
P=]DY705(-NCT>"7YM)QKT2Y57^4GK*5-M62OA4SL->ZN'A'B2\3L,1S 9A4.+6=7
P!^K_^F'==V#6D3P^("#(Z5]?>DWP.F5K_B9+_4KXM%:36 GBX8J;LBA[$JUPO<BC
PJYO9#;I;_)-*<3+0&FM'BY[7[A)P#%5">9N+09VTT4I T] <FJTT ^D_S6%$5F#/
P?B92L=&S/;<A3<FKXX$;4F" F9OU%9W10*Z='V]@'.+:O<0OKY#MZ829@D[VCF9!
PL/?/^9P()OJ?)&#Z5T_GXX::W^9AA18UAXS]YB69-ZBZHCL60$;/K#/^Z^-,[#9]
P=,&P]K/95]1&<;(4E[3&X@Y@4&O?V3,WTDTS-X%#MBBS0(X4X8) #A*>B_M^ XC-
PE@]EA+91<;AT,T>^JS=&>->91R]+$R.2]6R#U;-;85,RL%EW\4P,L5A *);6K&C9
P&8-JX!6 %/5R'U"QF5X\PHT,!YP&RJ48Q?-:I8;E@(<-@W^EM&9O29:O8$AJ>HKR
PB+DJ<YNO_)NT!SH$"_T0R6=I=KG5*,;(G]@5,U=J\1P'ZN*,P^=(M^W5EIJX]*T"
PB,*%,![<<[JQE[+N2Z\ZB2 @!4Y6$@Q-ZPDW&DT0DYJ3G,0URX.[4R%M0'.I8D'?
PK$E0J96Q@L8FSFU]]+?*), -1UA *(>6\/IT'OG[]8@4)'7?"Y<C$MC+./=M3GY0
P*K :*_G?I>-!KJ$5?WZD !8LPJ], LK[ -W+:]-OPQ_,L\46OCO?<?ZDF&D!E)W/
P$@N$&A:JJKCN#-S M\>'5.L(XTA,ST")/OO&:ZL 7]'196&WL&P%6KK6S7"= WB#
PYC1.UE(1-%JT[8 CAN> 8%<$1QMB;+J%"$@G%^*/<(K N>5*S6\R@YRY]T;5OT^J
P\1/\5CF&\1P@BMS\%5Y>9SL1Y5>9@!P/6F^/<UC/C)@)G##]=T(T)&'IW.YMX=38
P3Q:<,)=I+DCN:6^/&"K8.45H,FCI<[([D/_[:E[>\0>NW.N<O!/>PG06?Q2G]C5&
P4KHUI:1FT=A0?)V=K(K^SH:_&!.)<K25PB)ML&\!]YSKK/1Z 1]@K=N-[A3?#8,U
P<+:#:U,(@X5"HU]A[S2?EPL++FU?;.[22A<".IQ ZDNAS9$=>- :Q!@6F&X5M&<?
P8EH0HFU^7W[]>-7:GJ#*(!S/ MO0R /B\#X3I 5&,C:JZ8TDUAB5@PYICR.NIU0O
P7B#%<"S&O9ZIA8MZ$FLHD<(T-M>(@=8\DG":M3)6UL..(=W_G$OQ6C=S5>+HU'C0
PX#)/4O9^;N:R3V_*"+P<RL% Z!]M G,W#:4/1U3N'$V>*L:IL:F1?_8'^ZLN1EM@
PR36OH,AFEU"\>9I8V.XK<FX(+N]AXM!P'BL=%@:O\=O>>PZ!$0K?=3RM&:M*5CJ@
PPQ^:B8(FT>G9AYN,RUF>=TTN=52FF!V,BG,_+<8\(:[XQR)3<'08./]-C[?-44@<
PFA2E=,V]PIIM,K%>)->P]BIM'%R_)H6%- W?PFK),Z1JE?=36$Z\:R&@"<":,O)H
P3"5E,*^\T;.!/\IPBRP2*RXR4&+#[IOE!6[,+^[AMUOL7)7=:FDE5N0\+IA#6LW&
P,MC2O=*C,P\K]V@>.]!9ZU6XPFQ'JS-)<"A4"VL*2ZRS00(TCQ#@G+8Q/^;J$LJF
P3RA:,?/;F#S"*I^)(T)]^XO).[/?$\X,9#EPR2!&U3=H-ZY M"P(FB<C >1JI>=/
PD(M88O(.0OCW+V$CA D:1!FJV=37PKF)BM":@#7F\]"!GZ!#/A\A/'#2G-H9]P,2
P9@N\K;@(W=Z?P='AV;8N$IXPWV! IR @"H\DOL2",;.$X=6370B\3<J\P2%J1CZ>
P(OMEQ%UKOIL&,%1==SI?Q/Y@$V7^!,\W33WF6TM33,6)5_Z#-49>N/T<W8T[V@]E
P MBR=O+46R43<+?;) K0W.M&A(HCBF]^",3/_)O!>37T-+T$!,JZ$\">J3$9V!CM
PY,:@(4R>T#V!S+,(:?VP8(=12FXYXA0#H!7+\GB;3ZP'/^..]^QLJJ^,NX7X\AZI
P84(MLXP  =+4R$0Y^TFO_:Y%-!1I[9)CK- >B2)8Q/ ."?MH F?7#+A_OI7_7R)_
P+F,%.'ST'>'C3Z:7O4=]8VV/8>JM&G/VK8AKP07THW,BS7]!SI*9 \%]U-^O"TD$
PTF,*RJEKANW5)C^OD=&W8(?5+QY9<+>'&PG 95C  IO[NR00+P7DSQE1B(,TP%7H
PBRGZN9/D#7?Z$&A#=#G0I *2.CPGLGA#ZU>$U"("VMM6?<3.,_^0';4O*7O6^U--
P$.2#6N\D. \5K5>Q-@)=JWS8W=,L;&O;;UG@7(_1K)'1\<N5G2>XMR19J=787AFC
PYYY@?X6R8Q:OVW#+'&E.=*-A]O>(:Y1]J7LL:8-]4#+TSZER'[?;5?+YOUD:[8S7
PZ$]1UJ:?AN$+K&OO#ZO];5,*DR'1+9UF.E<AE9*22#5]_D]<EIF-=0H1_%89#VRK
P:/6"!%@O@^^XXU;MCMD]B;;NQ\P0EF[69KP'<JV18NG*HUD,/]8]+H=DO[4%#:JG
PZ!H_F]L?"('FM"TS' K@SS/6;$/&B"MKG7J>GFY.O=BDO+>AS#65OB%9/P1BI:A?
PQ(U(T AQA86G(+X6\G>L[(5Q$\$0N*>=YUBMT3Y$;?4,H!EGW;LSZMC" @;?*&UW
PTQR(1I EW54W(U$O$F9=;T*0A!P21GJ!2-DD$3^Y#_V>M(F4%R;6Y*DUA<TT\9<5
P@Z"2$JH$P6TL>[1&B<G/[&6M!SP(?^1A]NZ\6(XWK?8?S>W)^CJ!J$O*H!D?@\QV
P6:TZ:?8FP4@LH/,UN+?B$&G?#?/[RW4URIF_476:A^EQP.PII@EY]J4NL$"4QI;<
P.XWKAKK)X@N&(OJ_U/^?H@KK=2SY05%OLG6<//-L[^5:E1>,A71_LB^R0=475I60
PF_^>WSF$;RMOIB=M(JXP29P41JF< JUV!:A "VX3L,2PP=Y*B]+&69RJ+_.*0G>=
POU$5<C&=-C*0=-DL,XRQ$;Z]DC/@J*9/RU>Z+61B'%0V_BH"RAP8&PVL/$<&'=T7
PZVMM\./*K4*Z>?@0>WG$*\'FUV IX<>X]J;B#-2//+R93N>4 ?GU>)?U"?Q$I<MP
P=*)D Y_%8U";&O5#M:'>]1)\+"^L!U# 8\$DU=1WVS!+M1Y>W$+("-C-,\46P<"?
P!,)[F^&\D=Z508 3%WVB_>?ZEBN-5/SR5^QZ%QQZ_J6+1+E3].,(V0.=#8PB!1U3
P04"(W;Q:OP)3QDZF[]>,Y=/\)Y,*/3F">=@^6;$AN(&0+=O$G@QA8=H#)$AC8J9?
P]Q=!'G +OF40#5<5*O&3^_<6,)SV*.'ZV5F\NI!;I2?-WZ"9&V3RZXZ(3#(>X'ZJ
P\HSC+&8-8LSJ,-)'M?F )@SZ1#!9VV^H&9!'#DLJ!9LN!"-G%M%?O#4(+E^(\9(!
P0*DJ3-4C2@'%_4D7^? HG3;+TIN>)_.Y1;\X7MVKW?()GEFD2DR*BF<;[5DR?C'H
P$T8E#63&IFP$N='3H<%S@MJ.(*QOM^#TN14;3'&6NRO<<'(1GRYO3Q,U"7DSI&AK
P<(&=*>AP\!A=A<[77+B&NY6\:Z(RRKCAWVXJY^1<I]A2 52<SQHDQKY3[R;'E9FV
P"=\[,!1@0+\9! ?!UO]1+I;B96*G6,2 \'A<?(W57E86#?8GSWO"YR\5>M7VNIB#
P%'/,ZGBRXXGAE\2KE J]%B&882E$95*HW2*[A6\ME4A-@?R.]O"Z$18V\N#4VT4[
P(,7M,X0H6^:ZH;&?[+O*8/;.6247(O LVW3&G/< W#9(>3Y ;<Y^=/-C7'/]%)(:
POX.>\1$\N@ ]CJ+;,,=!Z9I'0@1!DXB(QAZLIM[C2&F#;Z/-C4\Q*<YP22&3ICW"
P/JAOC_&2D7Q^0H9VY%4:3Q1?95DU=OM,!$,;.7U *0#-7&:%7^?L)C"92SMG7H[6
P5*FAK%MYST$0G\'ROE."=M+1G2O?C!8&,"E)>!Q]+S*<XF-]*.F?9)L"KS)J4-.H
PA-"*/=GDP[5[V9X[#>XO5W"*!?-Q5W/E:-0O(-64)G@G<#*1K?3\1@JF+>QZK/^5
PZC)'M]]<?3NZ7?A5CRU.;^&C9-H?F 8TL<:9L7MN"T"7@"D)%FP&_O32=B*6$2A+
PG%U^=Y4V<?5$9(5!(BP!_K;V3XEY**H?_:L)+%@RT_@=*M>6'^WZLN?3WI(HZI!+
P=.YW@KVF1WO8",9EN0ECTQXA; 3D)G) ..*P!,5AN!SXIZ6Y.B2_#L9#]K-S.ZJA
PPQFME+7H,YG7G'T@^T'';4]'*%.CJ)3MXS=&SB '3?3M%G*/Z4<?:!;25G 'I_C>
P/\G#K+E-IR?YL@%GG?T]J@E!M4L[$BS<5.BKXY.%P:?/=]>1E(W#OP0M!W_11^8)
PF,8.0WOE./GQD&+N)7%5-T? &]M2[Q3TBN:+N-*UN;+&K],")K^N6\+]!3&\$;^S
P:73V$/$!8Q?2#:R:W@$O=&<EW"N=,Z^+2/CBVU_'9AQZX .&Z0]SU+Q1#(0TJ@M1
PF&;.N-7"49_4]UGX>"?*&9@+AT#Z4#,DS6ITWS2M:2!,J@__=#>C6I>?E^F1#A,8
P"9J<7W.19;\+Q9!S[#-B+MFCV''X>-Q8X#W^!#2O]"1;O?YOFW.&2#_#X-_>U60W
PA*,[O:9+EQ(S?,N,Y7%W -A7#A2P9LQ<K%'G2OL(*?K+NW6F$;/$0'Y3M0Z=3DG3
PB_2YJ7=KD!14&Y3*"ODJWJ)>SC:FB2)JS."Y")&.+J/(S@NV\5\;O7'$>1 J>6LD
P7(21?\90?XB$P[F.%"C21'PREG0+G2>^N7IO2U@YJ<K*"42V,= >>XZT0'/?N3SD
PXHO091&O-A,Z4OPO$>8R#++P><DM+ER%/$<A@^>!] )DRT'T55&!/[9CYZ"IP"8H
P8>_2/E;'Q/U8?7?03_/#!P=-F-Y#=F@-1RH#/5GZAJ61"(P$:[JEU][4CGF$\%ZX
P@@PLH-02HM8$4_QLE^<]RTVDP?LX>UOLA9]AOTN6?VB:.XG\JA=_W,Z7P ]"F5WO
PIG_]JK*WFD/$ YMC:!9N8 I0@*P9BP2BU+@S+*D&E.60;/M6L?]"%GI-8RN40 F#
P<CC:8"VRX3^\9- IN;7$9Q=EIDF93*$S;9?EC@ I,U8"3_#$=,C,9-<*S!A1\[__
P9G/:3G>>1OO333+3H"B0Y#%N*DM'0KGHXITP3*N&R(-YL4=>EKUBOG#%_MTN9RD8
PB4[$&)UKA:!U04+-!BFRBL\3&<Z@FT:7^WQK1V?\B('/T.!Z+%$YW=8_0T4HT9 !
P#]C9[4C$0<6JV'IO83AM,_S_'FG#'_6 "S:BKB=IKX5RMY-Q(3#<K:%W5=[QQHC6
P)F8M]A)D%+K"*T-;5.'2'L()]<Y29!5B^"0<M-_XXZ7D 77_&XJNW,["WEK&4;'_
P/I%VWXI38&QSH),C1\1W).8N4R^)CT./+H30EZ +IH6#,>.4X;]@RD4W77W%N)<8
P$>Y!#'UT*T$J^E#<)6U\N$7@)WOH6U6!3A -7%]?;OK1%/4AVR.$%*.<:UX"!:V?
PG00[U"KCJ(5<4?08H_Y]B_%]LPPD=BHA&2_S@'66[%740@%C!.2W_+HW9H?/74,+
P6&DA;R?VR&M_N6:AR30E*1OSYA=8 @:FFCGSV:.?4.KYCV<H:0\&3/< F?"T__<=
P97E86M*;I-NN^[C@#5:T=U$ G&WP(OCUPV0>G1<+EUP(R <3W\914722/#Y_T.#+
P6$B:$R?QNHVSCLA[P,9_PKQUZC@,4UM\2>< &J6(LY-7Y=O4B<J^(MT!3$\3A%79
PPJ(!WJ!5?Q?)/R9<O]!R* @'M>ER^PY< $E_NKXTY1O<I"[(XP O(S@<.2/-6P3H
PLBB7^CN($)V*]9X.V7T,-"V0.C%W >1\QDY_#(0SI2/+/2 []MNA$>2R@* SX0%O
PHJ\P4+5HUIP6[IIB];WL!2/V%87]&32PTGS"O\#+\*>=0Z$O-F-]K[A!D'3%OI/5
P#DML)=Z^MX$1FYTMP'G.;R;*/YRF].E\/AT#  F;K8,.)WP?J_:[Y%[#VOB!F5F+
P6\G/X:PL/[5FE4YI6E2^\7TK7'7\/3:GX @@$JRI[+Y_BH ]C:L'M@X>/O5S/DS'
P<HI LD#7F)(3E8-Z88ZG!HEWKA/KU &QALKQAP^?ZX-G$=+ @0^[;;O)?ET6-]RY
PF]*T3=4=J&U9!:LZ: F^CD/6F=GO* .IT$X:VCUQNI?33,=%?9C]K!#RA8$:G>FB
P'.(J? I=.A[M:<BANZ@)5Q06-ZO UI/<0;>I0L.]4D=>TKU(,^O]ZD(["?R!M/*T
PJA)90W/CB32J);$ 5ZS0#\ GU:R2>1Q$HH!8,O1'TRE'X<R9LP0RO5&$)LW-.V)3
POL)$9M)GZ%&C6)+6H.CO$W)BL19\;A,X676B$L116'%EX+@A;&#_YF_'.X$R%T\$
P!XZUFHO_+WKO8D3D"A3M#"GW5COQ&(V-R:XA%Z5E#N^8E7GTD5%9>)!;>4]2LUI.
PQA%@S-/6<%* 1ZMJBZ!$U*/\"T99@TO]W$.Q]0@TF:A,.B:=/CN/N)^TV>R6\]A1
P#;+99FD#R-*S.'21?;462ZK)KKUL(/E>EK(BE4]4(H34[7?S9"6A;C>OES_CN&^S
PE6^GR2&K&:5/#I!9SF^MHU^"\B$1F4KRS^5"? )7HQB2IX0 TAWSU,V=[ZAFP:W)
P5B,I#4EA&AO#6Q].CO#&_J\DWK7!_=?:? UY5H]1XS@080H]EC*>N?%X\(V;I]7:
P$X>$KF5X( O<W_5IBV9*,71:KGEWU;8=*].NXFG!+F$R+Z[T/.V>U@970I66X9\#
P-P="GH:=Z3>&5NV9-D@?>F]CH\C\7-62Q/OD=LA$X&DJ1@'1Q]3_/'@1+;#G2_%/
P]/+C".%!<?UQT[S1G22_V62.DB3AJW0$4#:G?I5QAF*IK9M<+B!]R].B.HY<4_5Z
PB5TRBK"XMY3;H9! -(2Y'1EB)@14;Q%#J9;K],8M#UH.5[LZ*[Y,-4:"#]/=,=^C
P0P,KKM(0;PLL#/[=)'=3H%U SN(R^ 2"P"V.(P/X*3)W%O!_WK POUQON0E=*[CQ
P.L:A%57U@DIH9A(;>Q@'%+Y^Q7R/01D 7[W[MM'#4O9.!_9#/5-X_(L0>&B"(IM3
P7=3E0;Z_(?RZB[LAUX[P*-F1AMCA3N]PP<F\NO_YNO#8A5^I-"P!@B@)*A)V@-?[
P_DQ\\PRPIM-,B'=$+B,$O:,$!8+([?^]!^<=PJ\#<TI@8+Q/T);H>-+PWOG>@W^'
P+,I2A?I17G(:G1L)A9$!H<82X]K+,T#:!(J4R5Y]*P87_ZWZCNJ=SK44<RDD%74S
P(V[@M98FP@'L_*RL8:_ I/FH$[!CL[3QZC4?#)/X>< V756%C3@_%'W30*_MLQ& 
PX$QR%W''/7Y<&%B'B.=.B<:<#_2DZ<FZ54)R1--(]F#[/B,(\J(&\C; 3/40?]_\
P-: 7\$["V*_%Q1HO0H#K(2US"-T]F7AS9(W8=US+_"]@2',Q();:'[Y 6Y@0XPM1
P+A2"-SF]0'4Q:$(H@-T>%-+%,%/](6 [JP>89B%3,%)@T9O*'?(TR9JL7&SF0/-F
P2S)1J6AE9.]D4G\80#G$%+0>?[,.<A#<5B8!>?*PPY I"%K <5C23H47JG-&!7^^
PJ+H>8VY8?3-AM9@QL:4_ZQL2#"=_2<\&XP<GB2*$.48D#:ZYK\))E_%WG%+:]X+7
P%N!Q,?50J-$J#YY+>D7A9(Y _9>\#V+,\O<RWJ+!J3[_A/JE#N8FI'J/O@>2[Q0,
P(GRVVE-<$ LA,)*H9[&E7M@Y!,I&XXFLMR!)&5_=)J66J^N5*1@'B^) 60-A@?Q*
P3=>YF ZL0W%Q(8K91+W34WG>5:_6V(A84Y[6$E[WKR0+_LS;J%\>(*'*'S!K%+/X
PQO075%$GX)RK>R3< ;6WBN0HP@S8*7X.?!.X?"2+VI<N]2+0E!UTJ^UV).B1'@,J
P(X'NR/]^"WWC88?3!*)E26^Z1C7-#@WCBG/)(TOP;!C4REG&7L_QEV$R0&_\/I;*
P1#M4\5C)9.;1IL>^^I@4_TVW?K#K1[ZGJ>*O ;<'^LZ0@1W8/NK_*0SY<C\S4J3^
P75="+LL'S_H%&^Q[B<*(US*;E4/\4>ZD0_G.;IT[<&H!Y[]963\Y<]^@,#=$7L%5
PS/H:A_[&:W>@HI JQCJQO7YC7L:& ]*A,"^'/0IQ.IV\C26D"D:]BXV9'>3H%NM2
PY*@XK9=QG FEIOWH =&=#2\^;P5B81WWOBD87M@:1<:M7U^OZE/:A2TXFY6<TE3I
P*'Q,HO Y2%Z>0Q2UR$<^ZA!54C8;[7LX>;/X!U;A\:LNHM6O-?*$I&?-I2/^7.,(
P2S&K=P98D4(_[IG6F3H959[PVST?]<EB@),THP_.7D*+Q[+BU\66,]F:1WA%=5:_
PD*.NWV6)B#ZOP1R;,#52M2P#"#<@_.X/2@$_4;6;K!*'EY5> T7QT.>BX2IL@&GR
P%#ASV)P(K^O(PJ\'\S12$QS46-^Y?5,-7?GG246:T@]N<9ZGMV^S0JF>C6U/,HR$
P-<BDC!".- .IW1V'!Y-,[2JG?FQ#KF/B1@M8\WP]^.(MJ#LU(R]I'A*C8Q?">*@!
P83*FM=&^8IPZ>MJJ_R@P[]GZQ;W@_7'4$VM*R:4^@R@*=0$18IMG=N*UZ?%DV]T?
P!TFF?C0(>\FJ@=LLU$?E"Y/Q[A+[_\"2BG'QS:&!'PWUP33(+MWF711:<E1I_HRX
P9+$Z/6_I)N'*M7?96-5JP1D )JY6R#,7T4?-P*%0K(6BR>&Z%P, &5C103K.6S N
PPG1XK,8(?0VC5@.!>( +-SH:X\[2I5"R=.]6MS>O5&J!U:[!=*\29Z"MF%6=RV7R
PXGA;(@J,F20YSXMIFV#7X]>,B9'1&8LFH7P!/BNT<1S7X=\6[SK*+7 G+R/1^XNS
P:/%V?*^>]W352_C%5"NEY,Q^>X#E:7FULY$^^,3KX@ %U284.0U_(P/!/.7N@47H
P9WL3Z,H_DI<S7\K/RV6+^-,".!D9K[([JV(;L(0?V/*DQV .=^UB$N1V[T*]F9H#
PV$;>N:WQ+-8S730D\2N8AU1I#Q7SVZ;BO=.[WVV&2H_PV[K'Y\R> LK!SZO22&?.
PUGXT/+(W!$B8"GJYO_*GUBH<GF4#$W>I1/)W\#8W/5CA4+_--FLYW8J+?Z[QGZ:J
PI2;7!%4@#8O?[COG,H:>@BG(^CXZ7]!LQJUX-![,8I4[.D[AY>J"[&H93,)Y)^K:
PB5OOK9+7"Q+N1GI$RU%?_]1[VHSQLKU$X@6XV5K-Q@NC Q8TLK_#^T7<-G-HP0?,
P[!1_A$=6_YF]4YP("X:X):+3Q>6N\6H-Z9%5*D>;FG*._$@ 2'^E @+,Z6D $S(8
PPMP5:EJPX_94^IX6;LB6+J;>[6M^(:B\;2S>]5")-R=%EUI 7K<] W)7)-( E,7E
P"]5Z!EL=*% B+RTA=96ZTQ1PK[6X@P*;T)2F#A?JUC&:AES?73O7D*KH^QJO*2 K
P^ TUAE7!_2T#^ZCR2)O]QKW92V6W-:*+-[_DXGRPP7-^UZ@^3/>1 <]#I.&\'ZR7
PDZOW<%11:K-?U>5&JF?H/RPY1#=W4RY5&=W./;L/]@7CC$^EO\S#T@UYR1CM(5'.
P]V1!7+52'0DNWM,.'[)%NS)F<6 Z0YZ1;92RQI183R $]K0'(*(O"X^:.[$ZQDL+
P^5TQ/.=FFZ"6'*=$YAR!8SQA9B$"KJ-M0NV?9%[L;!AZ<+U,9*+F_BM^!"&=KSM,
P\>><_ZY7Y&J=1%9]'$TV IEB7NRZR,*AM^#R2RNKE70]Q9XF@)$1*_7S*B'M@V>/
PQTI>/49&"H:YI9MK$$2R; 7*4MH4L+?3/8Z US/%N=PC25 C/?C1:'U9[SAW]%_#
PO\K,;22Y_!K=I(Z2U!1,>&)R9TOZ6MGS42U*FH_TVY?3F'!(DL-O>_T=<ZZ0[RXR
P:W9,82=GU07L5[@Y"@.A1I7P8+T"H*.B44BI_KK;E_O6YGE!1&7 10'38S1-;B.+
P_-=:#6_''I[PIX'?<U0SK_%\Y=Z1E*W%Q4Q5"-5=48T%&$-D%V#?DTJ=BMP<>JE8
P4QE,_QDZKM(NTD7[)\&H3P^VJY=?>1D8+SSC#QRL ']XN06>0CLYO)JT<J7;4,N-
P#@2Z:X,1><0$B3G7X]=?^>T+D]R9JQ)R_C\F$76Y9206;UJ\C@G*,G_/CFH3"4N$
P(^I(?&R<MV[T7PF/R*$2X>!5V2J#H,+NQ&E\HX%0:DM6A1X*VIM]*<A 8*L*$,:_
PS"3GF>E*P(D1]A+8M6*UJ:7A:-35DFI;ZM]U! -6UQ@K#.X> )W$BPDNDFW&1@U)
P4U 8<3\_:1!+4+!"83!RM?%WZE6UT_X@.Q)FC&H)IFBV(J-_C2X>&7DFA[YC:V$*
PD@)YX?@+T,X-GM0NA:;Y@WQ._0@+FYNY%+@M>&MY09">Q-E0YD'<V'1)8:YSQJOE
PFV$N] E86U1YL)G[^7R5JAH/OYS_N^EG! +,B2O&97L;LHY?HY%+#R\$0T.OK>8@
P0PT^VZ#Y["P7.',21A'5AL'[$.(N 10AES)=QM'?OU,W;3-CDC #S0'_R6@*I-Y\
P^K,W<1$^O@N;6JZX.\]R[,B;?<U.-.!(9>VPS1P:US%60U>NBNILJ/4G^MADFZSQ
P9$2[OGKT:*^X%YXN9&B#LR59)QQHO>A@7]@<&%;6<Y@8SP1DH-R.['!&'5SMPITG
P>XFC1'C"NGI_6QJ@Q$^OG2.ZK9'9!OW1#JK[%')V5!^]T])[WD,?67U-X@:DID\1
P,,XK$FTAN/<&U&46'?2FW.2WZ]3?UJPPX&M=UI!^&\S1H8G.H^"HC$OPGX^=QX<(
P<GY35/.JL2/'1X@"]^E9!V>^TLK4SP39_JB!Q03ESQ=F_Q^.,DO<[#&99ED8X2W,
P09/%0.%M2'%4+ W [R+ZFM-34]BD5EM_6[(;+SRD:0"LS9[UJ=:"!7]ZX,;CA]"]
P(__.HF83<AY<C%X?F3]L0)@^SDEV@/-%+>^\@O/[Q:?V<N*BS*HC#Z%@/WF1WPNM
PY3V2K%;;,?^U6N7JC !KLFTJFT,7EI[:,'55*[WD/^7- +T/_J?II@'LP!YMZ/(B
P*%++ES0J/&]S1S?1@Z,5!CO$H_(CW'$Q8E]+V+AD('SI*U11OIB_*-R/H>FWZ<$F
PM=Z X%;0!?V2QAUNO %LP_D[S&RI>*( T*9^"SJW)C'D5\0^Y)Z-%M!/GAP101B[
PK+&$%@+F2H@6$@WQE>$0C6\1;K>@[CA-'LDV%9^M1':?H4@[)RAZ.5P!^Y_\_OYA
PRXBYM2[JCR_;T^PS+$,R]S.\V K[G3&<CQF,> V!L:"7J2IOL.6FB)C1ZPUAA.^(
PD/&'-P$6Z>"L?W4Z%95=U-Z3J[W+V0[\"[2S"B,<94?*P+?27UL(R.">27^JPQ<7
P=@C>,,W*![D(+!=DF<O9<\@W?B?W@#448W<V2/&)>IN=!RBWLM]=[KN[.#Q/<%7(
PO,DP!^Q75BSJ3Y_2=4UEC+BUA^['8".J8<3B]1B\SI?AP=3OIE5_?A9^".7XV+%2
P).6?>*I\551$/($M7GQ@_')XZS![3+N@[3]X4=_A-'[FX+SB),@M4Y!,6%4KL0X.
P6X_&SZ5GCZ4T-L[N$>EQ$#>[4FDNAV^;;VU#$/XP:@K6]#>)Z#G*B?_)#R?JIGTX
P63(X.) 9FM.XA2OWFJ!D(_DG;;*3:Q;.27\SI[U:02G*O6SL9QEB>> =X&$;3Q+1
P$<AT@2-&T"_V@RO#XM=SQ&[%9$FX&P&W %#;=>U+=P)7+><6!FWWTQ>6T8>H%5!X
P8K7WD]T>&A9X6TU&1*.B@*27EJH/Y\#1F-$0?FJ#H^B(H;;/"M^&C[9J-&MOMHH+
PC'^U4^.9]:].YR;Z\84'$NBM^IH!N"0D/$1M-VL399VN&[]/T8U&Z'^O,0,$MZQ/
P'7W0&?P1\",? F)=.7#0W^"H33THCR_EQA*9^/0D#L;B('^SM!G^G*1UZ&%8^?RT
P%SHU*UM.6;);^AQ[L,U2^-T56UQ:?HOW%S NGX,T@I\I+4Z!X>VW4NVEX F<.VB_
PN%K]9+C)X:#:%^5T;K#@[1+STFR'ZA'O9KS7_G=]XMTGX@V(#$H^>T[/1DT*DKGA
P5T1<(7HEA-1&V*60!T8?-_@6<5ST9##(-')Z0G2-U\(7 O+Z:/O*E9TDZ@?Q,0?H
PS7-GQ7CP3NH ;&0<G>20.'&EU\U'AD9/6K-6KDT=\%F7WOMEC(LC[;^^DP+84_>(
P/YW\]@$)'*O2N[M<IY_1[+W=!:*3LW=A22NRE%I4RO][]#0G[_"[1V!. <+JP*%0
P)G[LSF@] B<??=9R2MLD83I>7\;],T8(OOAAMF!^ QN2^L<.6[_7X2P^VHZ%Q;"*
P)<=M,LO^/+32RL(DJ'(@#WE5YPK-^'^<)(5W\\>Z&QZPM7TS8C'0E.ARC3:,&P6.
P3.R^/2:(]@ZOSS8!M B9#+3>B& .Q0*!!KP6[E?0*409BL7>P-Z_&3GG-K%B+WER
P1Q(881*O<3B>FP,_HMT-)$N]^W_I\O5;.[TT[F DX.,(>H3%E^2'/X/T.$^A+P%$
P;+,D-N*=ZQX;DZVXR,*#(-01^[XN- ^(5W7[>W(\]?+61H$-K4"=!W/BH<3JA,1Q
PB@G6Z8H=)/.>UU@>?ZF*]"0&2 .R+1:K,[(L\D!7^BNRAF6;M)33PWB=N >**#HQ
PT])M?)U\H2LE=A+';[":H4CQWY"'%RX#AS\,KWTH9C_&EO\$35#TQ]+"&G*-G0V_
PD.7=Q4R;\P!U<(1!!>V$"F_:[(<9?&"AWLA:=[%8IT1HK=<J)LD2)7P?PJ2H,:FG
P9GPFD>_N3^PS(N2.![:!KT+@JD#<@!5WJ;Y:'Y$FG15^$3%)[ $$ A76YE14#,#^
P"Z#V52G)RV2)$7 ?? 9'8Z6T?3)_SO7:<?;R/7['VG8A0E*HK*DD:VNK)"&77WS3
P%Z^7/>[8O##!/=MOC\IL=%-2UW.O[)9$&.Z;B%,;<QA#1EQYIHH93DZ_%FA*R7*=
PD4*3@?@).FH*27F%KVD.?<&T^I*U1602]=;5GS3@/-#"%\(: <J7'_/B0#!Y/F27
PFO*#V=Z.6XSC+<_HD)%EDU]18'-*W/61VX.[_.':L-"G8@U*8#EVFP=^"254!9-)
P-LBZKPC&IH,K>.,.?L 5JZ'H0M!003>?3%%F4BPE#ZGK0- V_-3#*M,UW'@=!)M^
P\S>Q09J%SA7R&IO<.IG=(VL:0>-=NZ"#95MP"0- R RK L>K>-968#^%E\<[FA^P
PJ*FQA;\'<_5'S:N.FDE-D;'7#MUX]_1A,[6C%-4\E.KA&<D5'F1RFJ&\*M^% +[;
P7L5L*D*(K<M%11KP@.&KCWE$5PR+Q!$XQDT0LZY:%-$M))U5D5R:49LI<81FG5<M
P50P3LM&L=*J&<*I45;9MKBB@Z$C]*F6WI)/!?Y\-M>XO^5<LD[@ %R>CV,D;47G2
P7KH.0. ^D<X3EA:";1W;Y4:(DO (.+L#!$J>^ZB65^7W1AP*;(P.W.8<@-5V%>!3
P,O;^7OI&!ED+.4U^B8]B9_4D15]/,P32H4IH_<W>ORD1>K,H$_1;LUO/59%@2G;?
P;3^H $)RU%P@&O<'C</^,8S B<[F&:3IT9**5A?@CH1H&70;?+P$OP6$ISEVU */
P,#]F&&_$QBFXBE69-_<. >=/JU0)M;YA,V^4C%Q\E#G]XTNF$/FSD-4C\?KC0)LB
PVS6B:B$Q$:B=<Y]&H4?\.Y7]S:WF-$O<4'3/$C;2X:;SGND$[U*"D^MXCU&>].]=
PJI4ARRV#9^D+[#QVDY^/:2IU35MATGX.\ZR0)1@P9*IL](G:;%;E<!R@?*1SL-I(
P8Z'K#(]2K]O0@>AA#I_1Y6T&4RBQI"2J=<?)&<IFBC4H4(N^_8R7&$VC% 26I3U^
P-J0TSUP#J++6L2?/OLU]A[]Z[AS=]26!>VCJ9H]!\K3\B6/<[1_0!_Q(V#&9:],^
P9C'/AM BQBS\RJ\-%E+?15#+!W M][X))KL7KQ(P<C;&K\5C^U6H2CT4")5FP^H)
P^#O#0>CTANH[U@8-G[%%[?^G3I0'U\RW;O8%_PU[JM0_OW[HPG]:.AVEKYN*?!!"
PORB&\%!\SXT\'AYS(*9^06=:W^K0_43MW"CB,U6AA_+Z&PF.!F).O3."2(^'9H2E
PN (9E<H!=5@H=SB9O#:=L= -.UL$LEUD=(?]U$?1-7" 3N!,]Z_$-14$J,&=Z-U?
POJU:X,U6K&Q!J-<;CW_F;)SGCCFSJW%U+HH' 0UQI?$T7W?+<MW^H.67>NV/=4;)
PG7R;T=/_6Q#R/]IY5/ )7\3\%+1$E=NA$OM*48>F"LCV!R;MECQJ;/;A SBO>DO4
P="0R(!:VZ:QD:\=U_7G_R"3PMQ?)7# KOE=EL @5#X7_=7_A-*M$4-%<=3.4R6:N
P_A>FU7E_"2]SIFFUS.5QB*=Y%ZYAC+!#V L]G*)<E6KA##!H@S0]"G<JF-E2IT9/
P*OH\]M)'S6^#YFDX'HA9K9&0_9X&6%V3Q9WA3-:],?*=H':G ,,[5I-?GXFO^CX6
P7!3OX_F-V>Z@9,KCQ#:N<*>!QV-Y3%R'I?:8'^TZ.Z T1OJ.W3<?(P.D3:G)/+7T
PZ NCN24H;;ZA51<<&KF]N S4^FNY8S.4T![+_)'<DL9H?%MR5I:3CT+-[K47K5M/
PQ;$*8S[^W\-'Z^3"!=E.^C">$."8UD+KAK0V<W-ZL"KO6*K CP/0JQYB^+A9/7>Y
PC[5F>ZW+G1 6=^P7<%7^NEA6C<2%=(T19X>F5![BF=)H+BU#8G#)FR"MBV;_!WO$
P_ID#!<%+SPI8EV I*0PC2$/U&V#Z+H^7>L]Q9?;F$#3*(43MB+H&OPP3ES.]"NWL
P3^>CP/LZ<J -W^"T*@VUS\BYFFY$_(G?7(O%UFS/:85<Y[=:^9*#^%EFJ'>U+4F:
PW+177T!YH2"-;_' ]>R+,"!KR*6,=+$P<! 1$WE<+Z2K95DF&(E6E1WPJV+C_/-3
PCR6CS-3"U/I.NRX6Z\HK?H/A"T(5R)^Q"RVD_"AB3T&$\%(T)].$V<5JDA*OM7.A
P5S*KR5$1+/MIQ X.+1FK^K@<^TW/\V6.\RA*5N?;O,?@"82-SR[%8"D2VM2AKV: 
P]<L^S2J=P!Q.),"A=_9C4!:< WBAQT$7=TO@>4I]:ZM@NBJ*1XK]G48U>#H"Z<>R
P-]$7/Q.=MK2/TP*[;V676&VL$DHEW6%VT/W^)ZR'.@7'%#=L--$I%/,;TH"LJ&&1
PSJNDB8M6A>,H0".)O)4I\M%$)8)K#?U!GU+/N%%"DZ[F*?M4/FS:K=5O2@;0K[X$
P9NNBJ&8&E->!8A7%7C/HP[.0BRD2<:D@'-P*[/S=JYSW.I+$%AR,#@2O*6<DU@+F
P>Z"2YEQ; QWW.(!*M\#*_I?MV8OV!!KT93A8R,$YEL(:X3'PP'.]5UA2<U[CHF%L
P'$DW7(UHBTJ-P9>Q_2M.-5.P?Y+FL';*A#8<U+RH4HV;!4UX!_U./1;4DHH10MI-
P,<R'K49 1\Y=DCO!\^X(?3TLWT(='*=:J;M[.H^HA_V0X-0@ S<2\NR/?1%<#!Y'
P,"'#/<9WO+#"%Z<'/*Z^ /4"]>[ZPZPU*QV@>TK <)U.=)9(SH>",T7NU/KQ^*]@
P7_8%\"/^S:^WW[8<OMIP*':BFJ1H?@QMZDC8+*^YN)8 4K2I*3QW]SD*WVQ;!"F1
P));;3>&]-0LG.EO;^U9:F[?)=+U:[J!1.YY)K*W!'>,FM.9JE*:6/AJ6T+\[D@]4
PF$D#6R.5)Q:UL9,QRO6L2WB5X@R[1 #3R^Z*Y(LP=7GLCRL;W@C_?(Y7^<@/L=OD
PM*5V2EGV8KV.;%2R#%/5WK^$!^,:N<OD.I);GZX^S6Z+?'G)GG??+9U>6?AYD=9%
PE7FF!J:RHWLFI\"CO<S3WJWRSW! ][[T64*?9@YX&&)CGQXBDV)JLQ3;R2%ZC%91
P7/Y]]$=J%G[L;D%%.9/KKTY"!XP1?ET<K&6D BKR0LZ_^U\ VA046,N6?B@5^UD"
PYU.=+ 'Q>HQT Q3<^^_B*+R]QR/(DJ;I;IM&&9CA!@K3E5M$^ZN14F:]8+D-,-E<
P-7D@XPHVO6'U'O$T&5NO9">F\5Z:M)9\?87_8B(]&,(&2K<'BH6&4I8]SKLDCQ<X
P6NCA<^(,"[*M1W&-*[/6[-T SP_*J=4'G>*S\6Y##06$O2##H7VXY*CD,T$F?48T
P^94,AOAI%M_#G;;=NUPJ$R(7"4S#*DEJC7)&(&9,F[+P=4>EZ%_#\@]G!).2:0O5
P3 7ZJQU<:7N)/L1>#?Z"N]17<9:++5UC1: JD5R!"Y6%5X@!BX!U=3BK<$@8**DL
P^+L!26"EMH3;+I'HV/<PX_P@$6IF&&8*UC?^.]2_<G.A:C1Z$=&*L;,O]2^IDM6 
PZ)$,7HLD\.C_.SF]VAY]&NJ^=W(^.QMR \);/8\I"3^A@GBR3$'\DK")';BV>3GY
P]L*6,SF:6575<I&61$R]CPK8%'TT(T,^/]7P!7 BBUU]?XIMYIG.:]FOLO>:K$SS
PT_F5&F 7;8UQOEI9E?YO$L-\3YUT>$F^Q[\M^'9(R?>0E/DE&D\O/MH,,TD6W.6 
P[?3P0^4.4A8 =)_6BY;_I>S1BT6Z_:4DD-X)HLG7%1.HTBUEH45V(<7D?+_.5]:)
PU/[2!W!2?"!:TJ-R?ID0;/8P0/\+?90Y6GS7XX?:*=[4TI57X;I&P6+V>F5[2DY<
P.=,2^FN<S.+U&%Y&NX=N>(F7:G7 ##QO^W^)>[N9QL0[>FIL_> !AP:4K;B4KU5+
P>^&["0X0R+%H[KP!^]:2,*S-^!<W+:F6)_&W-<ZR =>&QOIKTZB"$:S3=HCKAAA?
PX1LP6+/*O_D$&DF!A(0_(S4JOB^@_C;^^5M2>/*IPP6-@)M70LCA1#QKG21\UDU^
P%291U$1A*)PB97OBI^]KQ2 6@60\%P#Y^94!TI7 PC5@^CQ6[^%TK%)N@-7NJG'O
P>E8?&1N:N:/+9-K'ZM69V^C1&!Q;&9FI<.<[]X,KVS(#7D9C$TYDU%JX+^3/<,UM
PGF!Y^.,)IO%QFDL9D7ZU(>.V.\L^25%'J):=4SYE'M^U-1=T7)Q;QQUY&8*-SP_Q
P]'G6P?3$3%@F)?/K^TN@,5*#H8UOCN#0<ZO:<+X=XI0\ X-V^0*%B\\3]J04!P\Q
P =W94/JA,Q1'J.+9(QE2@Z$#;@I@Q ?FBXU!=\_6.L/I]4]52NYS%7#3 40ENDEK
P4(#$3,"$F&FYH^0],<QO%4&:R'P'LWT(=-<C@<R2&3^O!3J1]TPZ,N@R"80JY^+A
P5'XIE^+C]]$'F[!HJO3KC,\?O.LY7$!!=#.]WZ%1UNOA4X&'NZ-<QU"",2.V?C&;
PDH%FFN' &3.C/%F++VWBP+&"0"L8=2@^*!<L^)31#J0SS'K8+4=9#+-Q@>[/JMP\
P*:[<**_<6H 1!37%@T'?KAGVP9I7S)5ONR?,;DLU"?,X3E8+%Q:NM0I@P/0M6X$V
P&R\OV\>QD [W]]-:!TQ9C6:3BO&ZJUS4AB>L)^8O?*H_^N2 :TPH%Q=H'_2;&U+Q
PA^'7]:S1#JVC^&X;(_[^O;[R1]8Q&65.3I#]*U=#2VOERF,RX^.62M5EA5@CBK*A
PY*O.4&; "4%Z,T:U\,;Y#"NRX\F"N6Z=C:-T)Z)!C >%ZB+QVXX40LVH^-, ?&1&
PE;[39S='?$VSI-^YKITD3/=UE(\/D(:=?**^\%G,2"7QX\N'=XQT'U9)+]E?J#A(
PA=_--V%?WM/H"_#ZL1.UCRC=F0_?U\#I?^3Y/_N"'_-C*VJJ(^RJ  5!H[L!UYV,
PPL_9#F72FP/59PPVO/GUPHCF9QC"2WFVL9[99BAA<Y*"/.3B?Z1<DJ0J_53R&T?'
P@2 +!^4KHHQ> 0J#V-*'4F\YT0TSU5:1UI[F#GMSI_-#(%ULAQZ+W\@\DN09P]3H
PD16*)5.&79M($D)(!* $L3) Q,!M?":.LDH%)<C,@2Q:"$SI#BANU5V$@1+L"(J2
P&VM(J?<U03/HIVHKN]L_#RCI/*. %^5T _4J!]_*:WM:?T,V!9DE99((\/[AQ>7!
PV2!J\/-$IKG9%77[;3'@F+IKAO&3\ J#70"6< 8(Z+>'H!2J;^5Y0WMR(SL43,^^
P*T2(.'E)28X/OT=>5R.&9U6L[Z%>%9@K3Y0T( =PX8RNT8=?"4HT@M>J0BSX)H!_
P4W*_2:7%6@3")ZS7-18$^O??S4D^!I+HE 1(R;;$V^GU-R\)>7)RDIR**_.JN0(0
P0-4I8&#&%)&"R#'#A2\1*P ,X7:1UH*3KW2_GB9)^6Q'8;0NH=C*\(V.BUG3-@QV
P\%"N#-\L%$(E&A>XBI\@UFX)B"T/E*K=AH$Y6E7<)U*JGTM3BI5T@PEM_\O->-7/
PKLQ@Q9A8^L<)=8^"]CI1K"I647$-D#O+6RCU6WSG<\UN$\/;I^I^%HD&P>(C:O<Q
P=79WD;+W>3IS=W8R'#_1+(:S%4O %H%R2XFOYHH40I?!FTQ0$V 7^ 4FRR71E?<(
PJ7R\I?OP<EMC ,3%Z)WBG&*=J,H-,O)0&8,)G![56N$AK5FHO7 ?BARJ8X_V0"=2
P^-CV@?TC;%#I0;A-/,4MIPXSR1K@O6%";J-)0YT(4 G5-( DE59):\#Z,S!K$N R
P[.NK6VG\F&4G\?=ZN3[S!2S+*!'5-H=^*/&'5;OF7&$;X ^8Q.;:>*L6/#.A#V";
P%LC"ZT7[ZCW-H#O):MAF:4EO8N(DAC6C2JBQR=)>SN SR0NXF@D-5.,0/RD-SEV;
PZM;&,.8+74[7K9I7G'(U&OMDME;X G](M)4&@;AVF[_>BJW(YAZ!4?L(H7%7N)V.
PL;N13D !P:$Z 3<.@1S0I1B\$FVR"^</(XU;<LN$4&69I0:Q#:[J-_1%,*@%SYS;
P40#C)KIE3UH,8$5' _A*%F+MAEAY5J>?<C;,-$( GIRVB*35ET/1(+#SC\WNDZ6^
PEEXSE#"R&G>H^#6!_#&KZ=R%/+U/=#')C13QZ&R,JHR=8IGD J+#8%$[^S4E5UQ7
PM"HFB_Z^I..&9@;V>'?%I)CZ(NCV0CQ</.7:P,@-XOY%FQF4M/U=0_/T^C@SDLFN
P[\O.=:67NISG9K=ITK6;0^<PS1[\3HAIJY5-F;*KV4,L&%6._(-C"H1&#/ Y%WVH
P)\]-7GAI (4=O2$!IM>8ON.I@6->C;A6!M*Y_ IR78JO=9(YV+Y>%#^X$E^$H4=A
P]O;W!*_?&I^QG0&RKG'74#UJ.$DEL6E[B\;8H?JG<"[[$.CU@<.&QZ';:\>-,7L.
P]1)!LA<HAG <OA;T]5(U$XD HMNN#'^&Y,,7-%"J6VEU#B0W(N]Q  M::6"<R)@[
P0"$^[R%5KI W0 '(&XMW$O ?D!WCRR<=;A <1+5#:1(219$)FM43P<UMYCZ(E'?[
P=$#5!(H'TG(CY?Z .'/H'5TO#,4J%I"LH&-:NM*JF[+W$R'Q_$L9T%[BI'LQ&F[ 
P>+,6:4&N.0% 0,(I<Z")/%^=;%2B7V23O6$XA%HA<\DW.KP6@U5.W 6DT:6FO?E&
P4)"T6H!Y&V%W"(.$2R)+LBM=-%E<J$,+.-DCW'SB<KKKHV C9=*W:X19[?J#C88C
PUZ/;U(U^&6<T"/2D<0A#_R'U"HI%;$2\Z%3O&Z&#YYTNC[IR/T I,$"0:@6*(U2B
P0QTP:E/VG5>.Y !'/[]=<V:EJR>>=4D+]2*%"\2(7)/,U)B!)+XABF)B7%OF+'Q>
P0.NDH)YI! >6HJ?_$9 47MT8V!W15LVOHL,)[@CG_Y^_0[+<HX-_>A]"]=95C[Q!
P,(CA,\I@[*%%/M ,)J$5=KT\CU_50? >6$ D= ]9="_!;3/8NKJHO][P#ST!%74C
PXXAZKU?80!VK=V!U'!LFM,E.UN^4J$>%<6*["A+LKO.<4#X36XXMX4AA2=H)&#J]
PT-&,+BET_XN755 S,NN6FRJ9GO_Y:1G^"!7$<N"FK< 7,YPN:?^UZQ0X;+\U%6AH
P[6K\Z[7WVQW2*6F(T%@D^?*N9Z^15;8=@K" FJ:[$CKK?:JMRG-C#?7'K3JG!/%.
PWX+F%<:#6A\0IY(&.*CY/^B8A(&LK+9##"Y:28#7!H>(NQ3.)]0&O#NMNG*O.D)E
P>V@@:G0WN$H\Z8WC?\D-^C%CP[;7O/M[\]Z;ZBJ'2U8VH86I;@#01*7;D"GT2,M>
PA$21IB*) _OX'@7$H8L>XWT\]7Z3/VR(Y0B=D/6J'M&.R9#2*JS1DMBP8FBH9C1=
PW XLJ:P8_%+\_QRBY&YH?FMN:DIT_X%/XRB,SREHM&EVI!T9(C"8V^#LU67Z_1GW
P\2,%^X!&DZ?[X/&$I7^9MJB,TQW-0/-E7,!9C<OH/:;O/Q8*BQ-SKO:2OMAS'#E\
PSO5-G@4.Y3L3-XQ#*HL)1A\20:V.*ID(?6C&4@N<X/[\E$NRL5-98V#P T[$LQIT
P/TE+:PL9C.KO+W!SE*3%8'>,=H4*$J:,&#.4(GF4=<4""P:8!,P2K<W&#J(M**)%
PJIP6GZ/C_\FKFE0G7THH.K'W>$2@D:*Y0\<Z#W&H= N+\^P>=19X"4O8A>=>/">]
PU)<?9I;7Q5^#\I3_VS@=G1BJ F!\\W5]"WYK'F@<P#",I)?Z1-\C(T _LY$2J 0B
PO2\/:^4Q9\ 12 )A'U [@Y4R!4H4DH[C$( 3IB7HQJ\!&?8B*2H,2OH(7,8G/F+R
PJ>C(&V\7"CM7]!8[0SNK\%R^/B$):9PU'VAY[A6P3]O0:5W,32F(<%9[[G@-0],C
P]F\G&]8!_4 AN?$Y,Q+OU\ND]]  T..;_\9'O'Y270MPZ\ R;5\D/$U)="[Z80U4
P&J5TPBN;J.9J;7K3N'O,7^L="R=JDB"N"^K;S*;)L0^N*IEHJFQDSX(A.\=.[HN(
P)N"CVZ.+]:=,@7Q\Y>M%2E910L@'-^%\D3\]Q[,*NZ?Z)4UA@X](\*/:XK*#ZG)/
P@/Y   FUYF"TMJ!H1S\IGZ":RN#R^V<]7\.2Q\ELR\04M3@K245P+6R/.NH?_$#H
PEH'+ U^:KRV*QP&8VE$3)N?B>F.'"&L_S.F@/RWTB\,WD$4/K:/@1___A5U3&E/A
PC,H<RI84 _6,37&8R\C?*#%]H[8/ S=?+,"\LND^V9H>Q[75H$]'!JT:M)6<DAE?
P2DI9ADS6%\8.\0+U1<4\Z2#%&!!F1,-DA#?2V 0M/7]0BZ()FQ62EU0B1\ (&^I0
PH'V]OC4(P.RV^X/"Y\G-K\*I#!CG7-*CT,*]\&"X6CBO%WNWJGKDB_#E*??"7(QK
P 35-J=H36\^H&%%W.H]UA 9A08&+DT#2)L*+_VA9E;L2='?//XTM =!;]AM=:;Q)
P8&%&KA02QD?WN]*-2.5!(<@M+DGM;#D?'[33 S&]L._K;-94T#< IG9_C\5:VQ4\
P$=-4+Y/H3#%S%.5RYV? &2R>&FT,8+*(*]&N'V71U'%LX3!23BT%IH\,O6DF\FA"
P(N\7#ZU84)R^M=<;)@5TZ:[PU0D8.?#]+P2K_$:3Z95/B!%Q#?VK\2(!54#J]'D*
PZ"CKU0-YU+_R%R=+!;D:3;0"(E5(.P(@Q?K!,:=]S+W8!O,7I35Z_?\V5F\NB@HG
P "B=HYD3*FM +IL QCN)%8 X'.Z_18>A-NA+CRV3<'M),T116K.147-.-N.M"&B%
POD.J@(![B9]U#XBG1#JRZG^HQDA!RB Z.0.]BTO+LWRWT8E'^61;;<X< M2H&$#>
PV<MV@VEJOF"U.!43O<#KU7Z;<LMWR*C4Y=A;W=EUP4I7V[SWCVSQNR'D[VCI?J1;
PNXJQOIC"O?0V<3V"WFP./,%I]0#MQ?.V-5B>6MEF<$1I4B1]1'Y'VYQ<>P<%F6;A
PXF8V$ZUIP.)'EF]D=PMW9Y9I(ZZ]95LL=6)OJBF]S%W?79!"?35!88M5I_N+0ZK.
P6RH:0&,7"LOS)K(#D1E^48Z_C051G+YHLJT'FY710Z^QP!Q)&6X#2U$35FI0!9YQ
P-#<P,2%LC$%F\D_D1#-(>=SXX2$!1A!XJ/S_2^UO.6O9.#DN26R".P7"*PD4<[6V
P^IRXA7O"&^TU:T@I<A/]B45;+*G=6.YM:'1T7F>,Z%D:E=_41%%)0F7[J$6J.OIO
PIQYLGG^8O^49EKG GC%JB"I_GZURB1[%!D_U<(2Z>LGS-WFV;Y"*)NG#W/?W)*?T
P].ZBC*?#*<_4E+D<W2F!V \C.G7LC)'TITQ9.9DMDI;8I2U'CMRLO]J>@7 \ZO-G
P?"7.7&]L*D>^LMP8N0V.-^6QMWL'OYOTI])&9DDA-NCY#)S]_P;)ZSN@$CE$@ZIH
P)OG,76R _6JPS3?E+V:5+K!_ZKUR%OU44P0<]J3%V@VU]FN!'0@YF,2=.-5++EBW
P0U#;M9]RV5F_VM%0G3.&8SU<>"<6!)]@?/K3%%:1Q #42M@#($*B;WRFVD;EAG?8
PC2^/KW7X&CX>*.2;-Z>:M85-3=$2*;V4IR7H N\$=A2\['H+&LI8ZVOQ"JFA1H^^
PTX-!DA\#,1;PM[/=G@(1JRMQQCE9QF*)I*?JQ"M7"2I@.J<$##3, 6O[S,Z'Q61L
P_,3M$08S437JM,3,GM'D&V_';(,YU"R=\4!*93TE?&$]$NRBHLYUE6DK5_H<-FY:
POBI!0GCRJS;=>6H8FP:ALZ2XX!E@=1 TJF&$!TYP7D"8^M]J4 CW@.68EXPM%NH0
P+EC!S8*02#A!B:GQ]NJ;D@31)?MZ RYL[WV)&:5TGTG;6!H0"'*LY*4ZA. XD[U=
P!;6 K>YC,[-3;]21&F$$Q5Y,VNZ0#!!5K^>_W+V5Z)<,FX%0AS^FC7\4S=:%CD#*
P/3 6]8\K;)T00DE,B-0W"!4V!\G[I3Y&"8XQB(L8G_<!V&O:'M'V72)^(-5&R&L=
PHH*E&C6:2J,%)2F.)5O]6NM57B'7!B\\,?]NA- /F/]!)_<*!A?O&/PCNEP!T?->
PV<$D(<[6T/[M!95P !1P3J3)C-^+?T!B<@,&+Z2?KQF@63S/)5PO\\S0)/FMC%^D
P!^"WYG<JUQ(#YD9/WWP4<<UDYXZLG(\O$F>UO[(5MOV\*5::W8D'J7-+QE#C9%U4
P2?,V,LMK<,E7J;L7-72&LGTU>NAH[8)?5I>>T9H19,Y0'. ET=,>LNE]J/Q$+*R?
PW@L?KQOY#7EV/N[HQ&+&*Z<*]'\/)YOKD(LQ'H=3J-H7W][Z:'NEH:?7HOZV.E/W
P:M?C-)%8,XOC*R(='S4Q5-$5/A5T'L9N]\L\>N_]^HQR5RQK0LN9\3U[_:T4[>B)
PV^5&*(IR$>X&-Y[,_AKINH;O71A;4'D8Z%W=0/F3C 1VB!C#)W*-:U]'4!+8J@-C
PNV->)DP^JCU[20T<)O>\-"]-VIJKWDB.S)VLVAS.ME@#0F,)SV265AZ^3BR-_0\C
PYL#^I2I2 =SH/D:CF(TATVY</KSZC?#D JFALMZC?2@<"\ 1+[:24?*S#+1_LSHO
PF%DT(+QSD&NTR\[&UH5^PTZ.V]3_\DOO10.VTII*2X24? ;=;V@U8O:45*;YA^7\
P.FHF<P4 :0UZ*0Z>-D(&><<UP?*L4'G_!$ ]XO1#X"D5'&QU*RDUY\T\ ^CE_.CX
P3376V'\3LCQI!2?<GU_VT%643VT.FTP/&W1VZ#^O._/(8:$[P;5MW@<XHC*S=#C5
P<DYLC*;A&C@=3Q'B_KZ=)\I!A9D[P??0$R"J(V:E?/^HHX!CQ,-9/:UR4</73]0'
PS?PD"-MN)=HGZ^$$&U,M)K2+%>S%4:-$=Z:LN<7J@M9.@:%%P<CXA+\2P)N"TZ(3
P*5M>',RU=U>%G2K2DTOT]NGTVLJW3^)YZ[9-&_E,:397 HK ']I4&_^ZW,^3S(F+
P63=CX7R>$NS=EC!WB?S)>A^0:1&B;>BXM!#1G^?]/2R)8$EX<][Y\IDN$C /5R\O
P8[-=<0,/DP^&Y1()H9;:LC@LG)=':6*%A3U$FUV2>#!=JS)J]-\^\^2?8?JZ^6+%
PEF/ZS_2&L3RM1K+ZN5[:7K#-QMH%Y[BOY]ZDE.1BI@MO;=4OU12":U=*&1TEA/\/
P'(C(W2J1Q[5C4M@(LW]5_D+E&9%%BH7RP =O=(#JU]0+1<M1T]7[:DXH;_35?:$<
PV;12,2CEN_-0> \&*$675R_<*E!J+;O6/Y7RC4S 3/7?E]0-G8@Y=  U.,L]Q5P_
PTC@#W2,0%/Z\1+?[SVB,<LV%1Z/)[!?O1)W$ ]1E9+8>91%*6C)J$:#EUFV?0=I7
PW_APSYX]<HNL!O4I=U=O?1\Z=A_T6N-MTRA#AHNR.=.3Q]]"("]]IY*2:<:A!SQT
P\SO0&,L5B+0O0/+AHYC]*87/M5/$I Z!2K9%[CC4[NV@)L+@EX4ND(8SN0^798%?
P<*]08\G@)0#]S\YF+.<;=M3_)U>R=D4R-%%M  )<AZQW(:'-3]@7P+64S6[0"A5@
PE8$3=]2="E(H>_];2D WA:'A^]PN6GO_<#=_C'<,/HUS27U8#;K'"EI$A/-F?D(!
P:CU/U>'VL+$Z"O(FH@2M5AIWP+0 =RTG#$V2?D,EEV)#X/-_/\>EE^*@DJ_5P%-X
PCG4.D]'!7%OTAU#+R;*=AH@3=B:<@0TN*"E9UZ,9XIHJ'HQ_.F&BXGJV?\5<SW B
PF.CGA?RREKEF^LTN<%,*^@\W.63U[QQ-:BJ/V7^T;D:G=SJQ_+<!!UN%F':'&_+C
P3U:GD<VD-+K6"FXJ2<5).;5'\7]3&KDB#46^Q;@9^D;#I]XK%6ZA.4_106[>XYZ;
PJMUIDB8LEX0_OQM"_2BNVP\JA:3EHC@^S$%*'3BK[3,+YA!L -:Q.AK'[>L5YO<Y
P, KQWI4AI,C2S[WI1EV1WA[*%.B^8U>LQCS\NV#C*=/37IK,?P.L26&N@8(F7:EL
PQG"T<Y \(<;*!(T!.F"0OR/OK#?]4@Y3"=Z1Q@R>^B5 F3K(,.^LE\0JB^VTRF;U
PR([[%& 7U!XB,L#6]DJ.Y_=QD%_VT0A*Y86PC^UG<[5?_H.P $Z>"_H!;A0&*L9*
PQ&W"NTI*7 V42QHO1EIK!T,9Y.'E1UVMM@3\O!H ".*2?*1!$--I1](:P&IVQ-Q0
PF@W!FLCR<:>45\:,/5G*V@36V)4!HAL"3$'EQ%S7'"\TJDT 8A*VPRF,GK*$41]"
PB,5&:.8/O 1.6:;#8.(<?!;4OXT?^[@4P5J1HUC#J^&\?6\@ "JBLV"V\HCP8MN8
P%"2ZE1(SD\;0NL.$^O"/EL?M95>.-12^[K#]-41)"#5,RP&:_O%UPF'[W"-GM%F*
PDID,W1GK7B_KM(N:([H>48.+I/:Q+R6YHM!7VQ*?F>J1O":T-F+I&VL(MT>-YLU;
PAW(^%'2M'%S'<2($,M2$I:W,V,)KA(0Q\CORR^$VTU2G*TS#_J2FC3C,=81'AK=A
P0AG8(0:/R-ICYL%=:,H M-72*[D7G8V!GC)&+[P&C#$.%/AV%_>J@1CDA9\<>DT@
P78W3M",&>IQ)K=C2-*>UKCAON58V19CYC<JI8%KFB&S.CW";A?K2L5KFCHY8X>G[
P@9W,=PP/XV+82J6:RJ-3U 9TS#2H&Y==*[IIFWK:P;5SR?[\/,F)1E9^<5UF^GC!
P.1SNNM!GD4\K.@>['$,CIOG2' 2$4T%\!Q5>$KL+!H3%V>4D*RX%I_5#G?&B\%]E
P+#D2BF+A:K3HK9]=(+O+#T$;]E'%+Z.4O[4*S?!WPW\];K6\*)RQ8!-NPH 7I\RP
P6Y%7.;R/Q?ZD8I].:3!]I$JJ<% :41X9LWI"C.E^[UV'J!$4O]WHM_"!&\H!\!B9
PZ)-&KI#M*P!%,H-WFA*J-'+:+;0_0HB@R!OEP&S,)S,&EG()!;8%;2-,S QV'1*5
P.VVTQ?4&;ZL3Y%[V*7W,'"V1+\G0YXO4RYM4MA3)Z\DLWC8&^+:L"^%ZWZ8T&(.U
PX@D?1%*)RL_$K+Y]W'N&,^8KQ/4E4> B&.3OK-+QRA44[TS/W9V23LPZU-JB;ZAF
P)UQ#:K;&Z,LS YW -"5-S7RJ[MQ+J'M*QK%088N(CM$N5-%CJ^).9R$_?')B"NJP
PU/-7/?;Z7CG"086#9, S,[7:JQY$2NM47;GAG[EPH#A(&,AN)<ZP]8BI=!)CL K^
P>V8VVA8ZY)>)WB1A3S+V,3X\@FJ*H;]?[4/K2-^05BDV:M!Y$+#O%B$["<>*TV3@
P)E"-7;_MA4I/BD]]8:<S#7OH'E?L>G0J;2<J/O-Z.]2BT?9O1-:?Y08 C@/H&E:>
PX:.V3W_SMPVITD)6<'?I=K37I/0- D?_:<W[)5+HW4(> '6\X81I3R/JZ(VP-%0&
PK+@I.<CW$"[JZA3'_:CH% <LPJ\DB9F98K:=R+XKQO32+O 2$^J&8M]'L]DU(=WJ
PC[<MRJ1X@'1WA0[X4O05RCM/.;WV5: $^GY^ 7[8XWX>.@*(1SQZ?DCXWT7>K\PF
PV'XPS F-%&+B.U673(XTVHNOTOYOU*O()\6MS/X,<ES,OT4$'KXB\+#MLA'M&.L1
PFP]S"%?QXF$D=XV!LR:4R= F+FMQW_B<MTO1S(*B?ZH2=0E\\&F* WZ2*GKAB5>8
PH*+*U_^SZ@T::I,S.9Z_E\:26&$73RW]?"XR36>7$"SC9U0OXG2E )PBA*&KS6N]
P?AQVJ,"SL= A.?/&,>$8N>%8M@H+OZ:S ZQH?3(TY7'EZJ]?T5/T]^LW619Y^(0)
P>(P,(6]P3L4>[K<A\Y%Y*^(KG*MQ^.\]FC%N?)D=W3:!S3@@?I VT[4L+WRB3XEE
P6QHQ&D3%JQ5^J>N>E>PYGEW<EQP '8QS.0?P+CN40J,G&&M?362[ ^I<J5*!Q09Z
PB^;0\[AD#I#"DZ*L,8_N36Q0N4$$:25:!SYFGC->@'E]ZF9H!?L"O"/E#WUF&%PQ
P7;\+K3D45I9-L8.O%+O+]6'FJV "8+CE6"HI'6;'TF(4/>K6MM/7C*AACM%FD$UN
PMFK]:6,^R8@9>ECE]U*"'T*Q%C3S'G[U['BMM$J=I96H4BVH@FOB[*X7D\BR4<^S
PWO%90J48W;>_U;(7 $2VH!;;B\WGA]01ZYX=XJF<P:^M!]^ P=2?W4"ZK/"3A%>K
P ^L!4F9'\_I5<B_Y84OF&AB7M316P+&,_"02(.L> #:DA6@"<9R,32/1N\,VA-"/
P:JD#/^%0(Q$BPW%CA5J)&3JT%"_V+M:4U17";S9%\;J;]J"8NF>6QJ$""!K%U/RB
P/XQ:=@X%HH*1E@4XQ1FE(LQWC-!CTL9.*7MA+Z0P:D?\_9JE#XL14LWI=!TRGMY5
P=\B?._RGF*2J"+1KX>!GL,#J-OPR@*:,84]K5%M[4Q\)4I4";S^N2D#[N"(:TQO;
PI@GUG<@.Y:^6:8&+-@UY\RN4N9WE>!8'158R[/\9['!*;!,*;>'&T3<A[C%>ZCRE
PVV#5]3PT?Z$K]&DM]&Y=BABHCRN;[D>8*");FBX080G.X<,%\)+X;F; RDL;0 1!
P_9B9O5]L5\<8GO\3U^;=9Z[!7B3<L&ELL5HHYOSWTJUTRK78L4]#JQ6&$LV@Y+P>
PY<QTPU8%&)J4\ Z,RTI\M#%D1>H3IE%E^+6A4!^G! <%F"D0!8#EY@'.I>(5FO1#
P>6)J?U50!#QW*F6_> 45*;I<>ECH([7Z)42\V!3D3E$OMBGRBL)+W:WOPV$6?=,W
PYZD7(B),_XN!,!"=T@62@DB%60V[@K<:G<%"&UD9"= 7&*[)-8%#"]\H4A^\I^SU
P/KJ7TMYYE6FQ4^<@"J=^MKJ9<XP/F!*@ZHJ82O\^_R]-%B0SU;=BA0]OP)^/H<YF
PI>B5"@X TD\7./N;MUJ)A9TVSK![V0?-9[PU9<K/5;_UC2"=?COXVT48%/#X(:K^
P4WL*C I.]6H+GM.4+\\PW!#V,S=&+O$\<]WR0:;LD&"CO>F=<.OQ!:->,M0@];'X
P<JG!M;^EFO7,N:?ZD#N!RWZDZOZ(J31D[*SB>ZZ2@^'$[U^;B!5F9<%VCI*/@H.Z
PC6P+SZF#8O!)A(> 6-K25Q,,Z%G?H=>K1WTZQS-"803>9 NIB[>WRC )&/F%I'3^
PFY$CE5?<E%TIE372C>.%>>":N(*'P4;F$S,3J5TRT>7E%%POIFOM4QR@'S1F<(VQ
P>GQ%]U[<4QED73P[*EA2_C(BYLTT@3KZ-G)\8S(<!OS JJ<(KW9N0C%<R++N4G]=
P#\&MP0->\U&Q#/7J16,/!)*?.0GX5QRWN=]]NU7&D 2NYW^3;7&+K: EUK.*((^=
POM>0,P-U5,SNVDR#;;E0VJVM^US(NL(ZD$%S'L(1+^UP)(7V;?.AH"U[) #=5//D
P81*92'(S-P;@&! KMZ'#U&:A4C^AE3^(5"VW<Y)HL@L-?E%Y3TQLJ'^-#!].QGDM
PY""C7ELH>U/7?'L#%(,F,H77(&LAHE4\&,!#<3J*W'UW\W%7]OC2U1VE+NCG2J%)
P"5BT$-Q595>\HKH.N-&0'40/H7-]G /J:"%W-+E[_J^.>>&04.,Y=S,,2V5CWV<"
PH:=?^D4+L<XR<I3((W_;LYRY0S#92MPQ&CF0:W6!T/W!VIA.QQL0G,FW26YL$/V$
PYML FOX*<55 ,)PJMO]W:;@X[9-4$(GZU>Y112+>C<'>(9&V#*PLY1 ?VG+!&W7G
P5X4^SI?QIUCPY2,=NRV&;2&2V$IP\\2DA#GQ-6HK'T6I:.TF?,ZY4-'G4ZF<QG'O
P$LV9W;I\\J_J7A/)@)2A3V'XJ]0=Z5X-U-("6X'0>@/%D(Y7"N-]69. N3N[.)-P
P$#*:%]%Y_]9L]H\HY+*B3,MZY[$O3RGF9Y-MB:LE\?I:BQ,[H3])[)0Y^=5U=]4V
P;,KBX/!"\&T:#2L'H1-V2H\&:BQ+D!Z==/OYMV]DB!:W3>U#)@XP(Q9KX:_] O(6
PKSY>%D*3B*G2#E YPY"YSZBGQ-G*U]BSVY >X[DS&JVB)N%KZN<4&;JE$SQ>0Y'*
PL#> '=6JNO]OO-0%>1W@WI ]2&YA?IQD:[[VX,*@(?D]"2NW?X%/XA)?$N0CV_R]
P^F2JH<#J-$AO:#K;_C*A"G5@WF"U.*$!@S7',A6V ?A+M[U  &)ZQGC=$FQ=SO;2
P_-N#Q\?[:NO"V;UE;*D7:FQ8[ N%%.;9'/M;O@'#]"TN+I31+93^CGM&H ]=,8A.
P#N,UU*G+T;)@H5A)<F")YRR8TX;=XY">4(YGF?QRF(T=YW8P+I3/TK$?>0JJ8Y/O
P^[ZS:9-UGFR'E>++YUY8?'#*6#QW!WG%=2%167ATYYE9!EY,"3;@=-F+*C64U\'/
P3!F:>V+Q*MFN46F$':Z4"UWY6)9D)*D472\G9B_F 2!K"L?E6F*X3P*(W\R 0R>^
PL3JGHX':C"XM@U=%RMUC"L>@AUK2)!.(>HW"]6CZ.)A!('>"9K21S[T9_#=P)QD;
P6Y:$)\_!2" 'P +?CN-([G@W5=0PFDUZ5$\14=3J/,!6K"+'%1KP_6B-$Q'!5H1O
P?EI:9UQ(RK5X_QXQY,:V=M9S=W/3-;)"4F51</O'"]&"S3_ OS"'=$V1 PH91#U%
P^/14!E?2ADW")OY5MKC"B"Z=W_+_: 96OP.?K&;7@N.ED$D=?-_X8\,&?.487!;\
P?CE#PN)<?8%GH1ZT' YD*_;F[(X!D'1XDV&ZUU(0!]!/38/D!F2= P,IBA-3VJ_&
PQL5<@&I_60--P<1'TDG/[=?6"7(VY [Z5+WH6T=R*/<'\GW3J$/949,3"(,K;>RC
P-A_V/2,Q!8X:D!_Y[8BRA@#)TL,9>X7C95K51KE1<2F1T*9=Z-GIK)5<J9\-+<MV
PKR1M-2TBDJB./^K#T6& #%_P^2]IS$+*-Z[20*6>+84KFO5UD7UBHP4B:C<QFI'1
P+?CJC,MBJ?]M7NF-  <80*<J"4WK\?:BW.V:W'&7N[<K2=ZV06$%^?O[G,IE_M)P
PU$2&US_^K&#B'^()Z'% I6^>#R*<)H57QM>9@BO017Z WCI@D2L;X15(W;^U&E.U
PIW6^LDU)8:JX\496A#6&M:NS5#APZ9)VOUI5@I=FRB)&<%)?$SZW:RN8/D/2AE_8
P]N2,5"'2JA>G;!LL!1Q,!,%IM&O>O;4TIY* 9[A$LI3B7OX0VV>YLT/>0H%BG_J&
PP=I^X"0/)V9\=<)V@7#KGM#@&C%3"A:B1Y1HZJ5X.*(3;F7?SVP$V*//>5+&(^6=
P?-7HUD/*,E;<ZM1PGAIIB[8,0^9+8][NHY1"2J"#%_,N/*Z$SM[;FOJROL<N/:2J
P,][3[!I1EH;'D5,A*34#1+TGB[W89ZL>Y-W:^?T\B%EWK#OID^?GT4VD&@_:,6/G
PRR<[!4[,D!Q: 6G3P_GJYJ' ,&(CN453$=+I,VEUJK5'[(Z=3+X4/AL^&RJ[9QBP
PN?(>%AYMO^7@!C,H@<>[3^6\NLUQAQ'/"'U$EU_^(A=[]80-.UB37L_:W(WE66O@
PXXU@X'5)KAIOP5K3M@,6F(XI+D]=CK,]#G=16\7X*?]G5IE[(BA^FWSQ!IF[U53:
PA_GDP+^I_<,9(&F2)G5(P*3VZH %4&\**,VV;'QT!,G+Z8" ]U\LYZ&1[%G>I5/'
P_0.Q;UT?J76AQR <DG^Q6QP"Q#J.F3CM;(JQ6F9A7;68%/V+'LNE^)?C/GSS/)\Y
PG:B[R-(1Q,LF[%A>C+C4U#6=TGN6\"D, '#2LS[VOV91!\,W'3S81'A]W)&V]B-H
P(X[?"D_\!4<I_[[0!@[=6V'P942CM_T#9<5K"!W:H=R@R2M]HB+5291.H3U&5TQ]
P8I/O%5[5@E+U7(.8J0U-S',QY#(;\I!GTN> B _>QN9PJHRA<>6O_#XK#N*.(@:E
P>"[6/!)IN7&>DY$RMS]:)B(%QW9DHR&0B:NJWS\GWFOT=+%A86*,SO%-!V12P3FQ
P\/AY1R*@FC7ZDTNNUUMH"SJQ;)!ZRQ-Q #K)1;$&(?'G^$.-^PVC6@4.J=GQ;"BC
P5;I^15"TT=GNPWP!=2Q\JI?9$*5N^>M0O,/,'162KI>J2L+:5$@0!9(?TZQ/UFM,
P4%DUP(NJY++0YT1(1/8\^'M'JNF,V%GH4/Y;*!6)7^$HVNMT^LWR6KA)3,CSL#Z?
PGN<0GWY(S896%R0]VD#VP/^%YE*(AIWL%@881&V$V34?Q3CD':E<1\'?C/?L899J
P2?>6[]L"-K^GH*BJLQ+\V)ML33B%9<9?HOZ:<=AC&Q_F:D'[21\'K62#==7<1KTG
P6P)&M$+/S'>=V,U\;5,7WL4@%#[[9M%!*B_'M.ZWE(0 !>FMH0-;';HN:FO2%/#J
PAVGX..6!E;PZ:F^.9.A7@2T:\@<$LO3'L6PD-=;(F$M<](\LGT8,4'W:*WC57K7.
PN>8ZY2^J-J=<.W>TJ5,,K+2KCTW=,[9Y.GA3-EQY&W9;. VC!F-T!>@$<Y4U!LJ>
P'6V\K9=J[B@YL,'&6-_!VNY^__Q=+\*)Q5&"])UC,D;5=@$% N.;</=S1?.I98)@
P^>K Q(D>EX+PMJLT%9E'.HA8WN$\24W&5$4=GH#T\+9807'D^#UDWMK@@7_]S3 X
PDA;SV7@B4=<'UAO^07'"U65)FHO+O)=ND4=<RX;=BWU *M:L=T3F0VFZJ/@FCE9L
P!<*.UQ$8F#30'ZH^]'[ *3]MY0GD7^&IRP&9$>*((J?K:%W=76966%A9 C<Q[-6"
PIC=<Z\% OGVVCGX'!@;XY<JMIJ*.5"-UBQPX"_4PH,J7Z"^O@9SG.8.J/L@'!ZVB
P*1=QO<S#IR\S'(UZ.V=QB9<<^"PA>N4Q4\_+,#_IE_KHU.D4'G7.6ETWAI%CLA-C
P$+%^KDW 1&<$+<<-L\!,\(H;EC5;'%XPM<Q]0')K>]K]MK?>#!W7E%X X+1"46:5
P<>:JU-AO:==DQ_\236"(E@-F=A8,X/ >L"17O HW3H[,]I?%PHE<1H("ENZFBQLK
PYKWU 0TW!.^YR)HR]PD@$SVF +73EO2WI^0!UP'NHA9!1PTNIU*N4D9X,N<PP&4:
P)JT$P<2;O^.?H-%;_/@=?,5]C>$U5U#5[W5U:-LY<8W\C"<(-5EKLKZ[V;M IPLC
P#7L%D:0KON@^)-!M2LBG/Z9.,6[JFQQQBB=_.K) :&4PY Q8%6F%=ATDP>70$ ,Y
PL#LAMQ *=[$M$Y7<@]NX6W\F4*O'=.ZP2:@=;;("4\DSGUX3AB&1ODA?'J)(WQ?;
P_++@"\@/.Z/PEMO=:7[YRI+Z&ZS]!!(LM6K>3[0.8X[XFQ&QZIR]=6?QL[%@MY9(
P_3TJ0<Y,RTI>6!AYN5'H+\J^##]!@C;3C,+BH"]>P!%X;+I&+@"O&'K>#H2GW:SL
PXG:)97D4 LM(.+_88G3IS]4QG:[*]/(YV\6LZ0DL8+D;H_F:J//06=>! ,4U(.I]
P@?^#=4=H/4>-#^L,X'KT(6H9+*]\SM3AL/=T>D+Q*NA]I8A TCI8\2-8OD[5T7-+
P@%=[SBJ9CN\&#R)JN62$:9:]4_T@?2H)9,8Y:<C<E80M_9;>J8P?3%$UB1R7OXB?
PC38N1UZ2-2]VN-<*LX0!!*[&''ZF617A+/MR@'9SSTJ_K;C;Q3^OD2#!H2:-SP3T
P, APB7"<P6T+\GYAH)"C"_#V[!,9_/"$+07Y,@_^T]2)# 2J9[)Y5(#.-;HF]O3:
P67 RB+BQ"_=VK],A,85H?*QYP4,EMH]XJ+][*B9M2%M#%S+84CONVER8-.I>LP>D
PW=]PT/X&CZEBD5K;LE,RN HH<6O KI4995O+4-@?=T&RRZH!7CV=PQG [YVA63=N
P*19HT3GDV=Z_[JO)H']J,R?TO-212\:HJ5 XH5XJ/T_8Z1I>9$HNO'=_)JK$)(U>
PBPIVD<T?M-U7>2+Z>(H.VTN,Q-@&I']%9?R+'??.$AF1E!0!P;3E!!3F ?U;;H/T
PUC6CT7W\7#"@J'A<TC;%024F[(D^&<BJW(Y. R0PU+X9!!.D-?JNJ(JKPY=,K,G+
PV%TQWGGX .C9N*DY/S];7*AVTGD'5^]"@I4,<O09^DP52 #?J>G8_7:,BF/XF*L5
P3I39XN$2Z7)(UM8K_Z[G+)R+KSK@6A9QXQJJ+\I4N%FO?+(W/-G"F8=*4EG/X\CD
P<)BX?:QE*U9Y:PL[<0R*&LA'H:B7,)U/9<X!\_W/NAKVP%O; _!Q%N.4B6D@*Q4>
PT4C/D<&81-351HA<5[-K@A((,_2KV-G+$DVR T$[@P$9A";49 +@=5 =/ZA0DSS'
PTH A#-!US'N_*I.D[%7R94)CLF\7+.Y-DJ@(D*%0TC[=31/RGG%V[ZWRN[[-6D-B
PR1X9]T 3/IYW6BO%?'0]%)*-NR]ZUE^L&Q]@<JE#MI#/\^^D=KE4G^WM#LW8VW'L
PPS(K\@<^ID FI6HPJQK-[IESZ(05K<5=P6##^V?'LV]'EB43\%&["O:2)ST(]<.+
P\E(N5)SC B_PR ALS/AU  )L]AT1E5VJ7&COOH<Y9MS/:Q6IR/?&N;]<:A#$V7<]
PKBT0<<NM*&9F3U]SO]^+G1I@EM&5:1(3GIY):>N'RB^,KCXCSW7JP!?:_._7%5R_
PB0OHTV=.&YN.@Q+;"-8^__,[UAE0L8Q=_%(L00SKSN:XM9V!0^:;9Z^\?[6/3L.\
P!+C\;!*KW,O\-4;O"VRM5]%?Z'1O,-KHAW\T)\CZ7*(IYJ?"[ $*K?%^G9H!5JV[
PT%:F/KH8#FO$FP;_DF.JDRK-_\,4J^()-BAI#R"AT.X\L&&]H3;TG29!<^B:[FE'
P*&I(@WRD*O3*P7.5LH__G(#HI'.6H>Q<*^, ZK!^W=Z&DW$H.W[I2+R01UEY07Y>
P"0&9_V8;^91BQS3@D@;:\<=8*8.H<V]R>H/(+$*SS#50AMI7![B5K:$*(RV01S&>
PAO*^79P+!R8E)9=.8T<*EWU.=1EB@JI&!?"!#.;R998J\[8/S',^<*V(YC?CY]TY
PVOYY 3(RK;4C5(D&F+S&F=U[QPH(K==-0*_0,8Q4 BWF\$C_0E09_M[T.6HVLL<$
P91F>3]8YKYST<2[5%&S+D'Z)<J7A5\\?)[Q9CO[3Z*H[J!#GPM 6..6.%MH ^$]D
P'5D\KOC5W_%'S](\*QD'(&)(2DDN@TF%N]R/#1!3Y@H$X5'F%UF'K'L)',.QO=F'
P'%E#B'1F8J:.A.AH#P&WR=/ <"YHXF@8VN?>0QH5!4GHT$/YJZQ*B:L.7)]P!]TM
P8'^ VST2WQNP?\M-UQ#32$*(%4X.&R"YY*GD#&G>M(I5G918:8AG:)[X&N=VO W6
P/Q&-7D)R@2"GF]HY&@)7__AA&$BN4L"[8%&'2\PNU2U8TBW>^MWS@_U7$<HEKBWD
P=3&%(['G,PD K0*74*E_YW^%N>BUK[29K0Z@BO]*4CDIN2T5V0%TFY\0" 0:?)K"
P6\?FC)M(1>F,M"V*O%X*!7!)P0G\D#9(#/T5E[Y\*E(#*_B)Z0"YK!!;;-QQF][^
PI5>71-C8S%^C ,FQ)C$B>QKF4 D4X6DE.\ E0=NS9T@M%\O;?E=M)&[$A(0NTU>E
P>@F%-G%T,SW\*0<5FJONP@EO;M)]3 YH,G&Z^2<@+<L,18#'3J#I)FZJ5BBF^QB?
P=P (X]9P97E_K/*(3$51JZ4779@SZLL@Q_+=[DM<^S17':!9A"GUKG[&$D6B=^4]
P:6>9<QR+'F_P-VG6%2A.I/.=R&(?HT%9LG*D!D;(,9SP-=RYQ4[U\63-CWS3QDUM
P;54''116AT9+F,(&RH5IR2SMSR=?!LOD2G6#PVP@_?R T2GBX$ Y29SL=;!BUM"Q
PKF7@'T><6X6 TQ10JFH2_L)D#S$7ITIO) 0KDG^,V>GS:!S)>&MG)$ .88MJ7J=C
P?-_/!IY!-#"?A5"6X,B.G2A^)WB_3!>4V9^?5S],HS"2+Q,,MF_"![#=RL0"#L8'
PR?#=B(ERQK8TZUH;PC_GG>]K1&H!8 O2]Z!/E?;K^2)!#(+/?QKS]1^+_,;K05'O
P6DKYW$9))LGKT28X(3V4MSJY"/O9+H/J)ANP@5LC>0&7U(&&2T?79FG]R'QOAP^M
P+)%?$@CFP+T0UW[JV!4JUU;_4C'?'AE&1 ;5EWI52Y@W 5= =,Y4'RPSSSWX):R*
P 1.N%D@B<@K#3G"VR;%M11?PS(%AWI88WA"S#S!(;T8>\W/I2OJS\Q#U>1.G/10"
PNL"J),$;4P"1@H9P6)<?@RU^NVTQ9'W*M[J?C3+^2XPMWK]_ #:DLVA?!^E@.)P<
P@R&H*(O G24N!!%SK4![P>(1?X\W3O]$ $9L0,%BVZ@^4#CBT62\(?FGGUC17R[H
P(CUO%YRR',C?Z0/G"\6\/ASN"6@673MSJWHML W89N*L%S[>/ZNTZ5>&N5O^H(N9
PY@PF_WZG&$Z?S>EE)_1=Y(/R\'T"VO7 <6VTR.O?F\RPUQ[,NPANFU<1L[VYI]0.
P5L$HWOZQB]BX8Q1E<@T_ Q+H'MC]/'OHI)NJ2@LP6B'R @+Z&SK,F5YP,CV$=#-^
PFE9)2N*19 ?*^@432S ]Q>A,-<=#6,4\-ZLH#^R->G_D@?9,)(LBS*D@9D_%IAX'
P4S_5P?QN;LAQ -HE4(,&):N_2!V*GM;!+#MJP]]2IBYE/3E-[.=,^MTUU*X35#Y!
PASJ6%RQZ-]?_8P47"1_9OP>2Q'KR@]!2K$.UD(N+UD[">;L@/&+/5+0=*Y1F]#6R
P"7K$Q=R0"<!_ 5&3L-'&@7LCIB9JVIF<41-_\*EP;PB;)R..-&.@Q>RUN)EE5HY*
PW/=P'UV@[5<Y46-H1-2?8%^U?#R>O8IY<H1YN$[V/& ,&?EU6I;PS KB4G$,:F9]
P!;N!77XOC8HMNTE'S]$J+3L'8 5EJT-XC:0E0'I^NGNOO$7FC90,!-?[9I"8C2T:
PB_G#2V%V6_L9>IE259@=<=7?@83Z4UX\?ZS9!]ICU3>."&O,[=\#>!!VV9'?ZLI$
P;<-IT/SH\^<<R!^AX-5P;E0:RHR6KQ\Z4).S ZUD4E&VYI1T 37 37XM.P!G [?R
P3IOG^T]-9LBKBV'++#'"IVEXWN[V><)  E5FV-*+ MN1>%BHA*SHT&.;J.LI;N\L
P0(*4HKS'ZFD,AN@/"?F-CU@#F^]&I;?LHWAU7T.%&FG^"T?>M#$I ,D>K;3B3\R6
PTAIE5QD\/OJ9&S>8H";PN;T/M)//:6S;_M#?7\4U\6NKYMX$8"A<0G%9(RK=D%ZY
PJ:(]V:\%>HMFU9F+4U)T>X)(!X\!)EOQS"I'L*H,I-;R9RE5%8K SV_D/%=[5A"E
PK5VE=Z?0O0.\C(Y-L;5._8JM =%0I6&<[9[?OROS3)G,;O#J6<3%&<3]@"GG-V22
P]KB:F!&AW8.G:Y<+SCLTPC;/(]44&Q_E3L\+[?-^_'H>;;X$H</4^-P4(+#8DJ)'
P +/R2&*P _M90"VRK;6IJ:)KX44-_2*NU;H.1W_BU.0"1@F\U&K<="0YU13_*V65
PBF:8^:9O52JW(8E+B''D^V#$8F-&#)+2INYEJ#L,1!*K)4Z8IM4J9,],/#LJG5"D
P![^!RJJ2+_1XQS58,+O 037V@H#)G$:-M8D1RG?^+N U3[KOC9L^<,&V4+:^ &A_
P-P</-?21V=.R2YM(0"93"'L-]4],/>H0B8?%UD#L)RK(/U!L! ]&( SOB(MH>78A
P$.MKM3QU7$GE*D'ZM).7LC5F:GPZ>^-C1N..%T:L<-F"7@N]5Z,V[Q1&3MJM)^R7
P*+FY11MR'=/4*6X4NXK@3!R_P]'63D,9=460=8] 1BX+Y5TN@LZ.@1]*IIFND6F1
PNQR4=0)TLPA7<CB"=K)P[=P""PD:7!^HP8$,>&F#<J3.SE%(7ORD_U$6MQ)C"8'A
P:B%=<S.7$^"E>V.PTD$=!%VA'MJ?$=.7W=L8AY#86C&+G_6VZ7YS%-?T27P%LVLS
PQD"OO;@,C8/3(82YV-3! %:K_*AP$/@RIDY4OX6%'9>GYY>!"+]3V9*<A<,+(Z%!
PBF1TKUQD\*^S?93;#L_T'H/4?KU$&IAMP%_%6XX1( N.#!EF;7KYG/4^4KV3HH=O
P80UJ?/J?"L7KEDU$)(,5"$U4_"3S%YD4^(4T4,!2Z[6=-$TR!PXOHPJ\>5_=I7?1
P%3WOH<Q^^*$"V![)I8;U_J+EG!]9TD@C#+$?H91_<7,LK%V'G,U;,G#]3ILZC82D
PTX"#5[S@L[3$"X)_,-6TV*2\$33*LI%R@P:,_LVF=$4#\_I'II!*F^*<!%#\2IBG
P.8>Q<94PO5ZOW7XOR%=UN&D^G@D@7^(W00"LA9/0(WO_UA72P509X#,9V$ZLWEX 
P%#K_\?J/XO/0%J*PHA(0SJ4MA@<SRS&/5A^>I/J;HMTU%R#P]SR?NV&GL^T>;="S
PD?;X^WE,X9$5/*/M&WAK$%%O+Q*MMB,<NOI^Q:?=[QL\1I+N539' K<8<,NHP?7,
PV8G-MR^NG*SML;&&/ ,HY A;WH@(U+!FK5GD7<_"[U")E89K(4X:*81ES^)0#OZS
P]K!Z$MKF*!+%^VN%)H]<J+7V9RM9F\BLKC&,<PU"69%RA0Q"QL%X>A7;<$\)0 ]/
PJ?5M;;V@G6*<?9$H@%X?/FZ/<*.-3_!FVVT0A3\+NXWPD[#KWC;P8^10=M6N?$\"
PDW-)KLS<-$.E<8>[MNV-":O/4Z;BE"42D<RG,IAZ]9H=S";P8CY< B35UU(40NXC
P*N%O#O:-843.@/%2?B @%[<+ZL ;/-DZND'Y?0T$R5;?ZXK9]T(F"2V_>]M+=U+"
P7B6H*A!PO_V!PHM _1(QUZ)#77P,[#C#7L))J?%T[#:ZWC<1B496RM%+\Q8E[X+G
P!N'/'>69-)GLHPB(#<-:L@,6&$N]/;'_1-T!6[)!L%!M/=8>D^:2<%[Y=HJ%:6GM
P4_,.['?IJ]\-(RI-4L+Q$433!ALR&:ZA'7=)DD.L:LGF&<TJ)9[B7%_-#NJP94>K
P0S 9'V.K3F_J]IO1A-GOQB^P^+ D 6_/T]K_/CP&<]_=VK"S=TRP/1S;1H]TY;F(
PM0D:Q,5$,,WE1>P/]C77<7 QI7JPAB,/^LUD^PGA1$O_20*6\(V-&V0#A)? F=&]
P+D4I&E*U*3F[@?.Q8TA@TJB;V!T(#PRR5:W-W>A.O,(,03.P<+RS]>M 7_['\S.@
P:+@^_6L_&]IA7U8EM&?QA:%&Z9W<!BZ+;>MXUZH]C<KS) "U#T)WQFTJ4L5?)G<;
PMTT?W+J2' (.EBV?%&9+#L9&)MEGZNO/JU8F3^3U5MUD5G][<2<OBN/J!/Q2KVO=
P$)058&;+MI?I'W^XLW(XJ59&G-HS9:EG29Y*DPLJ.=8/JD;"3LC[EY:PY-_"H*U7
P?XY>J6-5E"Q6DXL&BK%AJY+OV-_(AU[!$$YKASI95XZGH,?'?6<W4%/#WWS]KTK'
P9-_"2#B_0!-@4.ZTT(ZYV+:8,K"VW:?3GS"U;E43<PS[W(D'';- @R]9CS.F/XD"
P[5;-+2W%]69VT#V@,+-J]8CS.!$]F[3LK34PJ*@,"HPF#S&OM?ADY-!S<-"'J_(K
P9GG_M2?. GM.3LE0-]TL@#$9RW[1-=R&[V<=1ND[S1S*7^LG"FWJ&OGT7-(BH*W'
P/P_&_J'1?&H:BAS[0%%VS:B@G<,)"RK\8?+%!F#3KN0G#8Q>Z)\LZ9I53&ZM/EZ*
PJ+>_)A=3K[X]YFC;;;A<N2+1O5,0U#T0Z8:&&5E@1$1N?B$:OI"]\<O]E98ATD'/
PK1:=+D^'.#. 29'Z@THT9)8\0E^0)0-.]WZ"5SK40#6\5T# O5:[HN/S<:\\&X>S
PMXU-(5$H;#):,KX;;N1,+$LI@"UEELL]"-DW&4"JY?9!A@RI,XQL&\5R0>"M&1N<
PQS]>9-5;I["V20BM>1Z)[8OHLTBF=>I_:SU?8SOQ>L4><[BMN5%2;O-%1</)&8S0
P/;%_\D6^([!NQSI='<6/T>CS52)8180WJ9)H_X3#91-)V-ENQ6$3__?K8T_Y\,$4
PFPJP&C=GY\. 3(^S[R]$OO:X*V!N6?9PQ#*3>QM&UU>$.3]/1D1B5P).C=2J$UW\
PTC3H54?.3+B8;7),7OLQUI*Y.ATTP-\"#=9NG^7IOYPM=I^F<AAY"!8_5SI?\F-?
P#K^FFH"\!QM( JT766.'2!3.IB%_SJSQ BP))@UW,86ACBTJD=[J<9V):7'.&&T(
P.L)*-T 'P]MGYB*716"3IYM=ZBEY;S_+*CS,N<"4)QQ4!W;!BO&6L)P>,9_E(2R,
PSB)CDNTHQU\GNJC!,MM07MWD7O-+Z1NK5X*3I:8AR>QQ [1_AN#V ,)PWZ:?PTNT
PC^M1>AK#*UZPY\D=T^W6C:'J6B/I]5\NB5TK:3T20RR@*\N"2F95&KAD#2N/ZYK$
PJ:'//#VARU)Y@C/$'"8RC6-RL\7(L :8?W+I;CT_># O?*D-P\U1Z8&38^TX?(=H
PBJ,\Q@VF_4ITTT59:37\?X3S&C*EC"T3:U*BAX@":7'U^KH?X3#WYRW!P)B^^KY)
PUGA7+/11;<\[1;J\Y\3T5?GU$R71W$J51&KPM7IZKRFSOG"-@9VN%312>"(?%%U/
P5D@?H)O_.\IB6_D@'^6G0/<P9+3GIM6QLL6\8P<VRX@AP\3U5Z?VDRT&"(HS(+?:
PQM#FE'YPA5T[?,N'<;T0QK[X2H6$%T-\:.2"Y030,OJ\['*/Z4F-<%RN>\!@O-&9
P'B+S3<+M>]_;%U1T8N%D0>[CA]9"9SAMB:/X+N-KVBBFABH04OZK*5%W!NS8FUYS
PRJFT!$62[&*_+7YCP\276DZ)[!G!3LOKFRE;FU3AXQ<GL54\.:H$PJZV[!6EGMB,
P)OBY,&/T\Y=8(G2PY%S4R4F#N Z1'N!Q^B1""*GM7Z3G?SS:2,VYR^8C=AYOWD[C
P.-V]XR^P%O'0<!PEY);\N*/20H#D-O+KOPDPU&-"\7XP4ZTQW-PX&G9*\D^;@7?F
PTN)9M*\QZIEY$T$=%V]CY3J QB*K5-?*$Y0K,\.LHYD#\$6$G6Q01'G?'#I7F"#3
P(9^V4AT<ET>L5X;T->0P2F#>!H:D1!3D<(#\%\43/ *Z[LMYD$=P]X, ]H-%9]7;
PFQYE/'93U)J\7.M@H!BB H/MI7XG*>^PJ<*OH0WF=<>0;^#>!&_$7JF6"0L'6SD!
P6M3;\:SAM'ME5H*N)70PT,=_<9S5B?.(>V8#E17]\&*K;)AWI9-$;/6<LY\,YB(:
P/7]]M0U'B2#T'*,TM:>CT^>UB]U$9&TX5.PC"Z7O4!PNP22K@!1C0!,X^N C:#8(
PT^L@OBS-[?ZGHAVD8_?@]TALE3=3M O\<97MK/N)+:)9@I(UJD;6I">SYIT."Z!\
P)4F3C#P8Q>A.%\E4V"FBPC<13.+;#3EEM++(^3H,\9W1A[P9*XU:J^P9FP60HPI:
P?JNI%7/%6M;T'T:5"NO.&_^;&P\K"._L0:;^G=TT#%S=)EF/UN\S9A%JW=Q=KY]*
P"L6((W^W!00%KUZKQ+GD?9%'4LJ+?HS:KI04E[!F0%"2<#G4"L>Z).HU,S/]?QN/
P[&M<G$P(ZU.KTH-BKLWL9T,F-]RX8UGO.YU:JT#>R^^/]U=!U(1\=#S(A0G_]D@M
PVC:\C$"A6 IER;@077S.\=!N^K=8S)I?BVMM-E6-N4WP/+;1D"OQ%,<_]12CQ@.X
PE34=:V#-)I.?M9<XU;-1*<26QQE9&B.N,4_-1Z?"2/>Q] "]UOK ?C%-6' F_C)O
P3,:,0-/)3"J[/O_EU-JU<-*<+:TH%0M6X SOJYAR\5Y/#4S;7TFDZNO;C8+%0R)@
PQ RO*R93B?,XFF./I^41]#(KS?=_P;)6$4L*(5RC8,!TEI.-)RU,OC^S,2L(CUJ*
PZ!.,H'EWBN?)!J^"ES.'=UV]NS:\]6UUB+R21Y_(FK^KO +3ZFA)W_'AI$O>W*V6
P> %?\.W8=V1%M!2!S3!88+9?V 5<"D/,]>F _OZVU/0N->YD9=YM]X<G8#/#LB"Y
P?@,LL<R#<0(;UN$$N19U4-SZ?<I[0LV2)4#H^\A65958S=5N4T^^K(=S09%Z4E<7
PU&1"9UA;BN('9!X&H?2DB#H"B#/+6LN^[Z],-1]8T!N'WA93VK$+Q",+/C?$O;MQ
PQP1#I%4'JWT\)#6/RF$),XV@OG_N9X:5:D+632R/B^:[=8U.PP2 ]>%+B'81D2H&
P(B39BR"*A:[=!*QJ=]_;!.MC.2,G;MA0TNSG=Q4*K1'DJS\3LV=RM(.6O%:JV*4,
PF[9$_EG*-[H4F-K_(AD-[9]M0!CP[*K'(L'Q;#\+V[&4WL@H?K4V'85^T\9BGW9\
P:-,OONDW(>0Z MCL'YLX^#M%Q_AJWSS$TP'L#T0BX>Z9C"-I=-.2*T/G[*MQU2E[
PDP2*=G2G:$HY^'LQM]2);]S:TD71<IY+C'E>W%>4*UE"_@,(+%;$GV8!D@]E"@FQ
PQ_W&$[-N-+GZ)R, P*%!O#%>7SR8&0D-VZD+CA P9C8G&\>Q-<#Z>3H3?5$-'F:0
PILL%K":231WKU@S;S4N@&G\0125U@P)X/'3/#0F>VZ9H22V"&H4AST<L197(%BBV
POM(&4+5/2=J4 1?$JQ9-32WP0K2:(&]HR4JV(A>[4&;S7N_9BG>1\P%&#K'6R'K:
PV27+6*QSOJYE[N2W4.>E^@^]"!7MF1UYN)N0NNJ/\88,Z>JV)SM];[,C"O^\G=!<
P\=1;1MQR4YOZ@V,XC=0R$(Q_F?3_M!KA,P6Q6 H(V\<UU6E.PNJI&A:X>;YV86K<
PN@0_K3K@A/OTD,A=_3@$ S2TCK" **P7IMP;!\"'1LZ>2Z0E:LNMV#_8K\:&L?Q+
P2\.;?7[ZG567_?Z3BB*,;ON>8A"S:5#\3'V9T4W53#0''E<_<3J)&].CDMCL24N<
P](*@K27=C2!1\%)3IK\JBKXC50@%5)N%2'G2_GI&VH_@:+WU3'LNW&&33U",$A:'
PZ\=<E&S[IKOR<TBE)Z4>9)W5K*6K:/!)%"L-6C4<^?]M&//WU1WURJ9!?IK6-\,6
PO&/Q6A#,WS;E+404!XVU^=('U .>$^-P))X^VQ[%/0%RR!;*FC@5+97J& J3'UPE
PR("G@59GG7A\CLH_'K3PI0B+)-VJAJS/0FJC4&Q(WZ23)LN(<:WBH&Y3TZ0&,^RI
P_J6?!Z,)(E9N39P?<-:YLF%:47C2\=H(FXN4]E &P9MU%:INP#.<2\][?S@]I?VV
P3JW"/QZEY0W&6QD'W;NR4++?*^])"+!VZSL;\#0IFFO4Z^'_Y^H<D2#@*S&?*9!?
PDT[# .C10HLH>M9UGJ7::C*M-2ZXY'*HS =]FW'J+-Z+E::K>]5=?]\^0 N62J_P
P.'@B 9:/J!9UN $3S5!A6^$M[)YK@"P!U+26KV_J_>5QY[<I<YF7$W@DPYH[OB)$
PLR;F'8M#QOK'02MXO[CGHK#8!E#3]R:G\(&Y%NRNRZ=3,%I?SI0VH,7[D%O)@<#C
PUPU7()P-6.>GIQ70L='9[[6YCU]H/R21P-[Y1M%#"\6?6SKOJYQX#R8T,[UMO+P*
PCV1?<M5>!G^UILV!><OA1>",D6 N@/B!VCQP?QIZ4)07M/4X]!8(_GTHJP-/"6\-
P4Q@0$D9%A\U\"X6D*]&+]I,3>'E=M 9B.4(8%'U1:\A;HN'QI"R8M#KAQ>:, );9
P^D'FJ^NDZQ"5X]M=T7N^*8D_-9FCT3_.HH@\S<S2]0--_#J(YR-F\!%OO?^'2*]W
PXR:?F<)'Q]P"%H&ZX*)P[+#XMO(5<-325O6*EF)YCK$%PT=YUM:+]<PK'5SBIPR4
PU\28@M$Z<[B#[A'_0M8@[7 1ZWG".HIKCWTT,%ZRTT<L<@))*M[4;U4U>='FP@:V
PAMH?UD=LMOPR@!-]$/A="?*>$# Q$/JVXVDNLGJ66KJO'SG*Z?9I&93>IP$@YH3V
P36<5(2-2W??Y+)M,:\=U0&+,KA6OT?<*4"V\$()M7OI.HH!H= *Z2!D3NXJ"0N\]
P1UV'%B.7?"I[2^UDOXE(6?*1&N7.1<?94P<@WM'^-70F>#MIGV&U')3%2V-+\G\*
P-2D'1K!ZD:@I^_#FKN^_GNGLX^F*]TO: Y?.UXS%^?EQF<Q/ /YZ+2$>T!X 8*^*
P:Y2W4N.((AB'ZS^U??IYD_7S@":B@]OW-&I.VO_TF3[V88*;![*0V2^;EV5FO2Z 
P!8XJF19:JZ59]]:>/$1/@"3"GG@_QD^IT@AB9$]]H07U-#W[Y)!4,-0&P&*!V7=7
PN64^K25-BEUL$C0"<9 !2;!&5=&/J4U5;TC>$;P:K&8;_MU9H[)]PSN'ZP7.- OW
P59HP=:?>PGXSBV+K6[1M7VXH3!QAK=.]T*G=G@@V8PIN$6^@6 OMYRR!J?#6X4 F
P1I@47E821M+;?Z9NP)#4P<P30/Z6D[O>!0_LM/X*W5GAO[%O ,@+L$IPS:S T=^:
P\W"I\NC+(9 \/ [X T[NJ5:T8E=@FOL9<U-\.A_#\%#!)2-8!?'LPAIT7XGV7?(V
P@=*G -(:+ &8FU$03W)TXP'6-],![[+R-N7%&WK7SF?ZUA$PXIBJKB$B_"?^)0/6
PO.S;W';IF?6&\AEO&DC/U]"+85]P9RHOVB^:HE)]?<-(\B=;>[1".N^1D"!#@7#C
P]W6XP&'P<F[[9CF[Q%87VA;T<<5TNN_<1YXC8-H\R5W2&.^JQYSV5V1U_;0GUG(\
PMG;[MJ+X0ZY#-)D-J3(3LJ#;PW?!2:+M?F'7#:C)WUF!!%,,^%4>$PF'H2<8]GL=
P#;>=[0+"1;0VD\DCFP@)#@'//U]+J7?)1.O:!-^&3VMGN2I'CBD<#T9@P?=OE/0\
PGBNYY,K T%XEV/963='$D&Z# -T:]W[4!W*25T$I&'._-9UY&Z@N] &/45(^:L_]
P6RG-WPC7XG-%?#!%SVU-5D\/98^&H]TJ)H(#C[8,3S3O&D7/,1/$@%1="7DT##( 
P>4K36S,U89Z@N[N'0%PCZ9'5@HV+X<_&4B9(9*Z,L%JRVX?\A<-+/H! ';\YL G)
P:[OSPE= .UF9"RGL'.8!;#O5<&E%^'(=^ U62VZ$'^Q<MAPPH^K!A83YO$)]]3V*
P7_6)2L3H':Z3;;2QWPA;>1V:31C:NP$KX- /&)T>P*Q.FT8^"WO'+#F&P4TA_)F#
PS B+QA6W0A []='YVJ9XQ(BILSXY:Q>LN-K'/CVO.<4OYAFI^[[FN@ ^>IG*Q7<N
PQ9,T2%H*)BFBM$T!>R2PJG1,#J7U_\28=B$(XYV5WG*_($ZSR[ DOXN'TW+=8 *"
P"*!Z"CXH.1=F3\_>15D,#I.4V'3=XO:PWU/@6%'2B@4_PP;-$&&.AUSE*>K3#*<!
P)*Y:I 0+C#;4]CJG'.B8FZ2^)$,6#5>KM1-9'K]&S^\ZNB^65VMW% 82(A11&=#+
P$'_VOPSM)".28* CZOSWV2%#2 1"HZU#RD(&?/@OBAYK=)WU,CMP:X9KI KIV; ^
PL ,8LIUEX@%8D0C%6<&3#M =M/]3F!6&K=V2I]BJ9B2BIR5U,A<T5L<4/1N@_$]:
PCAGX?XWDH8%*VRO(JNX3$1#@\Q^Q/>]TR[6LTK=I8T6[CMMR6U8;3OY/6&RG]V.6
P+BFL6P2^OVVF /:0;6_=K53+=27D[(MZY?H]V6.T4UFOOD=+]I5R W!6.^F.\=&E
P82S'PT6F=U$C$8%;#I=,5T"?YMVX;:VNW+S?$BRY,/E:O.9USQK\ ?54G.ARQ$DG
P7F@1;%IV\GWY/78/#L/-5F?8/K YF6,U)RP+V?@<$[O06PD&)R@UF:<KI_L;9WES
PMGF O%3)GBV EXE,M\1F];[N@F\T-"NN_2=#:F3'P8S2/=0TZFXB)Y%0:$\1V90E
P,O,]3<Y]S\'W-@Z#AW3!,<&_H\.3+\2F]ZA(+DHYQ]:4[=#&9Y$L&M0BYP90]AW.
PN)! H2Q#;@G_Y]1-'BE:2I0&&[!>Y)V*UC_0>?<79>^FO+]A%).C1C9==#X/>@_Q
P4F8F[:!=X349>DXKGY2D#AS+: YU"EKE(HZ)!_0\1DYI,U-:):,>A;- E!P?GFXC
PUP!J2\YH<.G'TX)>A3/9(N?+T=-<"2^=RC9WV9[=]+\J<Q_J5+YI%B$='\(*X8LR
P A-M0(DUAO'_@)^J72;L-B>Z^@WB&YY4T=/N*X$X)U($A6(KS:_A0E6VXM^X!*HH
P$M6?UA<5&*_S;#LG)IL7[L^.:^>:TJSACJZ> >["J.VJOT-?RO?;*0C+' >6D'.3
PU,U1T5!-4*EOD+NT\>HWV:*XC=U<@B5/.R>W5JUJ0P<+\X%-=2@6H#J402.2UU@U
P9!B8=D^WW3+;2(,\57C3TKRV,\7T1<___&[61WE_N.[FT8:=4^H<*6>4=\$:74.2
P:O Q=^";P\(FK[>*B*?'7\\4[^O%FB,.OJ8@U!LWHG6-H<V9;H0!%?(0CDDV8;59
P9WG1G=#=3A<"V"%%:Q+KENB%BSK$G?;Z)K]34*H-N6:^]4S;S&>L2%5MY0.E*:N;
P>&::$\NG5F:.'X3PO1LU(YWT4&H\_<;.^)2[.\D>&X9$)G6/7*2,W8V85A.CN$Z%
P93":[F#7L"^VO+> S4_N$=[\CJ#V'L$PLQE%?V;/8Q6'ER\&F6$&*W&@E:@_7]:.
PV4]@[#=\P65L/VL-Z1>J9.UZZ>B)#K0XX?] 4<_#(1R4L=?2?B=M/AR,!5MZKS^B
PL39",X!^A/'W6E0I0#]:FSEXS'S@ \7Q].L!TO:@USJ+A#_'"HI@_>-KZ)!QYKM+
PLSU5@LQ[6M_2],YO7+* UR4PPM@*X,FDLZM!5-6Q$6ODD0I^1'K:>)GA3MB-/F'*
P"WA5G-Q)/K OUDYZ]\R XDIH$UV#+*H@>\-&>*:K&^H1WW+ F\;W;AH+8 $MDRVB
P+E+Y/S+P>MV761.SH?W?<MZQ_ :]9.5,=?VD&814\.DEVX.QEU'6N0)M$Q3,.;*)
PA?GM5-V?I-_>>L[./O-'Q<_UVC)3O)8L2T*Y5P/,/86AO%P_<B$RMXC#T2UJZ. [
P>LQV&:;\M^)U=-'-0W=EW& ,.J[KO%]DB2D9^97081[]9VC("^X;,%L-!*.WDROW
P7!"TQ3G8BB7BP3F$F_)%]^MFSE8E,"AFVM0VECK=D^N550VKHJC^1U@'%<7]T\@O
PGBJ;@-+ML2Z2\0:/#23:4Z >3C-(0Q/G9.OLJ)Y@NJEZIST1"("!90,Q19"XVKH8
PC^G8!K C891*.02YGH2U\28)*X -=G='"5)L"O;Z#+_8#&V=X?X6A^B-.Z4 2 ]4
PMWK[5>//-3G8>(@+JK9.! .8 >O 1QH1@C@U9WNH>P\"#O' AAP./:QB2HT?\I3^
PJ.DO2?ZR^U&8UF^7D0H16X""F"QR 7S]:RWP0QL@%(4:QY4*@4Q5_[H>"HA]];OK
PNIU=[([<@BD.+9]N&!88_<ZQ(3LF'_Z*XV>I>@G3,])R-E1>8'0?W2*0J4;B*0EV
P*LM[]!2$DH8IV&N)*NA'[XPN<DC;O0"CTPAN!L=$Q]-(U%J25*R, >&M#P^0A#_0
P  ()9#<_XRBXK(3U='<(;)DDACT5TMI<>[?$9?&,+IH,&&?I@]6:?</@T!8V?(+;
P3N<H_LE<8!G;[=9Z<3>7KTM6THWL'D_B0>+[4,0A ^M+]A9[ 2ET[PKYTPF"VVC6
P")06_;1)41Y; BZL.6BY6'QOX5;VC:AT^64]J8IYW=5.CL@:1K8S60 D<TOLJ9VY
P E8:"_] ?9WMZGT8N2 IT>&;^3(Z&VUYU>]W&3AJ79P$@5)^YN\,)<1^-[UX*((S
P NGDF>4&S&J&+:1?A,D1I"W&3-9AX$<#VKMP-/NH-3I';]E?<7IO5/1\@[;4Y>[Q
P'2&9VQ\GA0R-$<XQ*]D.PC27,N?DH^(99VVFS%H(*R V?!<@X7-_C7$@)@B% N_Q
P7\H^BZ!!<>".(6=088/N41E9\MCGI_/C!7?8WE".V.""6K\1P=Q&YB65UMS 27]6
P.MGLL$5<[PK4I0&2YS'#+IW:PW"K!R\RM[WO\$375<V)[;/^E0=)>',PDF;_/ ^X
PN"6#!G)"0@(L>LX3 ,):_%CAIUD]0JY-1%UN24<CX_7VJ)/-^[-J8 J.!8L:VV9;
PQ[*4UFF?CJI7N+"&=*7:5$MS;XHZF\F0CR]K]#$L?[C?(EE=8I&D#CGU0.WWWMPA
PFI*I,/9[N]Q74X=6"16\;:73F[$VJ?^!-(WBJ68R,-P?MG7:E&P$4V!#U+Z2:2,4
PY3BHX7H.=RG%7)<"UE)HQ6:C H0N!!I+@KX#0,S]!3 7X\9:<V"&6&CY!L:)"-SK
P;C(9-BC)?-.=$8T6I3OYZ&(;1#1W0OBX8?#A[9W2GV/?:ZB75N%7$#UM"M]1Z<?3
PM)>K]GH(7R4$.M!"RHE*U*]N[ZRD-BA1,6;#WC%=+ AVZQWIJ)'.F@8_)G6$M56[
POV1T+;RG0.&F!<1N(RM"O]OZ%G\U^,]W+J.)(.LVXK9/]CNE:/'6_I2.5308#U8,
PHO(%KE0J6W-JS-\UG;4U#+0=OIF]'>Y3R5#Y+?RQL3KT )%:O+VU=C^F!;B+58SQ
PN(XDVZ]4GL&&(?KA&#'P:Q%(@ZMUFG!WH>*_7T1+K.\@\7Y16GX2LP$I84BGD]DU
PFGU<%?5(IZZ OR3-?<8.VULE]W?Z%%%0/!Z+HBL(]KQ:>%]>7A#V^Q=.7%+2Q3*Z
P9Z,_\4(5'E)GU]60')<\U]\+SM4>V8WDZ:T"T?.=,AX3?(]$$E3Z7!<!>BIO5O12
PI]!1C;0 ]?T*; 2SVY<1CE9#C<"$SE5/L$QH;N\ZNX%^^X=# 3M(+#CXV*G[6#,8
PZEYN5@F(G&B"<F<J#9D^%LX<N#%J]2>-I&#^W4^H2_;/$^+UE%@*'/,?,*""*F.A
P!@<YO20X66:]4FE4(&C\HG ?)ZAY^]+7F!Q?GOQ'K"&+"I<H=*G%,[3L.*:@L)2,
P/WDQSY303HW^B9R?$4 P;J0)7W#-FN*$YS)V2_"[;3\;:AHE6KM&@<N#&X2 P$T2
P:@C,"^+R9:M<:5#";G2#&"NV93)NJ+&:U%VFIR17V;]*G(.FY*$XV;S,G3)W9**B
P5=N>;?KXO;Q^<W=118:L:.#+H^UH%X)N(F&'R945K#KL0%7KA&Q7P%)%-:_;N!)0
P,@%&:>I#(V@R.@ ,-WWS,=/*+%=SHE)UC5KBHV9<]3S#K1\[] :-5+5.A[3-UV75
PZ\U')GQ,_*#LAM68A*OK:#MF T6*43F05W%K&MWHV1_(WOE837?D%0U3ISWD][T6
PRGIV9]\P(<FUF X46BRQW5OO;4>J1H?I$1T3_?.K/9R L1/!/KXD<\V9=E]93K-5
P'A;&^JP:TXR'KT(>4+JXJX'TH Q<L-T#AUJT4T7NQ;Y4 SS$S(JW'B?)(LU4C<-1
P9%3'9"51?EL)!C$3:#0%69_88ANC59\O.G/-\\?!1W)>4OL$D[Q+I8I'<O[N+ ,A
PC!\EB\)9C2Z4+C66/D63TQ_NO\HDW\D-KJF'NHR-D_/;'8"Z,"B5UX1U%W"9F>L1
P\)J&DTIX[K=JD4^:@Z;-+JQ\".:%YL'VKAO@#IJS%Z'X2"XAK(1#CH_\)"FD,0UR
PF52H& ?()^&#SPORW@[1?AG86_H0J2=?FU,H"?UJ =8=P'HWW.I:A@U@4HL*=NR;
P#/?DI#=J?+]]DOZ,9L_,Q+Y*P"AA[I_3SD1U0:WKA$P@Z&>*I4F(BF/+C];!0I%X
P*RV.T'/.@ZA>=)SF*?O_%S-([A05LN*3PLG0QE9\[E!7#E%/]3XCH/'-%_&@?*H-
P4&G"?*KO:F4#YSC,WSP0Y+LL/WMI#)4< JG?#!5&GWSYV*"^"S7HZX/GOS+S?H$F
PMYK9Z);L[P^L\_KH3$_'V[2!=W4D* >V)5XUR9U#CK.+66VRZS1QB8U#7X'._0E8
PX5XHU))R08MW.T+'<*/H B_0T1ND(*?_A:]6ZUBJ"C"K!/_0)Q/ K<Y877JQ?EW<
P5K&N3^(U&)]?_ $&A6]K&!A</T!HRT&VV%+HZ;7/W<&!HC?<*X5 =Z?Z2W&I.;G7
P6_9K8K5)-62U\#:0]E^:0N1$L+A[B=9._=<44!X49H\MYUYOP:R^,W!DGJZ%=>4J
PD+WY=5:T&Z$'2J2K/"C7DTH[ Z7,?#>%A/@#'.T5(4$.Y\[^Y-H,3836)ZV-*1*(
PE(/]H5+,[%JCWA2)_VAVFS-+Y&J@:=A@)F+>HN0E"#__:&4=J1\A\J) 6"V#T'D?
PMCX?SN](*DJ<1(9ZBFBD-+L8$UAP!L[7S0W0/]IJ4V$#/(8]?Z[7K1*@60Q'SZB<
P-"YBHP0,V@ _25?K4.IINIZS'(Z+)TD-#8_34QUJB4'BJP[Z&J!(B"EMB,!O8ORN
PAI""P0F<&<!)!V#9#C?3;[QO()E;U;RYEVRA\^-&*60,WRU7D";W/F3)9$G='EJG
PH@ICJ7QL@H6MPR@ +EG^O:=![=TX7"+5J:=%<&&[SHT]U.-]8#-U).E*G'6#\@V[
PC?>R3!UKR-@_"5A+X%GK_N+A=46?D]S1X7WQJSHUUDHIH]033=:O8P=CAN<@XN50
P_( :VAPS=#:X-8S:?G"0M"D(Z&$K:(R/YCLTZ9:+SQ= 6O.C-D#'K<GH7)@7VQ=S
P<B#5PNA562F?+MA9NG>)%+MJ%VANHBBO=]2K/RF\]VY3=SQ?OTGC-0SSQ*$V=+4F
P:A?1#,K*K+TXXPV&K/*;M/4ZGUT1^];Z[$Y,N\30*F'2]4TOS7LA^QH'2J(0;:(Q
P:@3@^.EK#:IG'23O3>J>BEX//_S#R<@)0WNPP20,1%V6AO244#FBJ;N"\%,,5J^W
P4S3)FB3C(9K9>*%>VVR_77G=XE1*9[QI854X?H6EH6WYRT/8?^W95.^\%T[/^+I.
P19['A6%%SGU3<7YW"0"10 '5.Y5J-E<J@Y_[.0OVWAH19CQEIK]X;T_X2;^$3 "&
P4(VD*3S-5A9\SE_KV/L ?>9D^;>N%T/]79@^K"K2/&)8Z(@[R)#8OU#!-D:?@F^^
P=5TSEV#/X3,H+9I:Q_.4 &W8G7W0"O=$V $:?)LV;-XO"'\QLC/BZ$,E75%S&4K+
PL7U=F:3JSXVT\)Z-:*4]\AV/IM5P;=]%DZAZ=:1EJ-_,DS/=<1I*":!*0V>'*'U^
P#E>RU6,.N(-#, D]2[A9D&<J,B<C_U+ZYM2-I+OH>0:HB_ T$:TWKE&)9/0&Q7)D
PN$Y,?B:YN+C"ZG/Z-RLF!DJYY:VA^RR?RW!MZ CW#V@4G-06),:[ =<9G]'(@DZ%
P"0VC7JZV6A-CD)GF:RF]@2EO;0QOD+0K,]H]RW2\2ND'E4DN7 :C.; 2B9YHH[@R
P!0.\3,X17C.3*#H;]JK>?\)*B]U.^O"GERB&E*J"#0A/80J#(0?BE7_F/NF+F9CL
PIY_,26JZU?%#(.#W-PI=1.VVFDDVF*;LN/</#CLD/< )>UB<\NZ15=,<*@Z'B_L#
PX),UG@P:FQX:]95C0)PTOK,+9@<$4TJ6;KO)E)R5VO8MOM+2!/RD*W?&6RF-77=2
PMU+0_R%5BT"+MO6Z^P$,+E%[8[TQ+ :8:/":]=)]ULEW@T>J-YP$Z,.,HBQU+7X]
P R]_K*X>$8("8?"H;XOW)["AH_+[F7\-)SVY0;[Z*-D*/ET,54J<%Q%>.V4TP$60
P7O!:8QCDQ([F"_G0@=:%(Q<+- OQ6I* H<4CW+3;L:K6+T_S(ON]VWW)LR@@@DV6
P#&&W#L)^):Z#N&0S8"FA\<T*8$"(X-K2;%KR^GT#7+9_JN7@HZ;>#-=K<<LFUA-<
PFY^8EVL9H HE-5L>,.QW%3/L5U*=DG\W>9%/IF;F@'(C"E-BY[Z9C# DL,8SM;1C
PGX4Q+,9LIGGNZVJD3NTHQ/;>6WG908$.K>;P3[60TS5F5/8L-CQN^73<E[;-PNDV
PBK"S]()A<+DWRN+!0N^S%0_OEA:5_E3O WBU)N3I:-:&")[)1<+6-LS9W]M=4OB9
P\QB%1VRM.?R?[CCT#OGAO3()L)9NJR\:."$"ENTIB=LWFWFN2TQQ6!YR65MU(W D
PP73L-,GG/R''FBQIIEYA+X2GC1J3R/72M:Z)S=GV!.:'3)AJ4%?>,8VE,]4]N/83
P^MY-:*BV(A5KY&.W<+."-%/Z<I<HNS7;8P3:E;A6:6.*?F=W$]EN&!"P,2M[\?Z0
P;-O[%5 $KJZ+G5Y805<R=>O+L">8B1.KO:NH95.CU],X*2#X%SRN9,A),KEA\&15
PV P5@+&\U^R<(&H+D5G*)5RD3\USLGBGWM%J:*IF"Q #?A\=?1S).3*:0%1^>E G
P.1[Q@"#8P9O7Y/L3EIJG'B#OY%#Y,2K'F0/?!DW/]4%5XCP_+(,WFM.=.B9'Z4&5
PTO0J:J8<;+).GAKB8!_1X('4>.:)'LA$\QR:N@A_[RH;U]7I39PR'-1[/,Q65Z_%
P?9T_Z <V(V<<'4^U"=",5?WJW*91$DH:!^4C]@/VGO?,Q)I:2H2?FC[JA4Z]MS\C
P.R2 L,SM5!;VPJX*N%,(M#30P/?J'Y<04MV?@?&NC))7?<+>>J)\9VV!_7L_8F2P
PAD3A'NY&C[19D+MV1)?L>78Z5^N):H_;H%7!Z#CR0*#F8TW9V6EQ<NW5B4V2P@!&
P1AL?EZT.6$#[[):85]J(R>\&\OTZZ>'LX5UTT%40()-.,C^FT,H)/M^(P.%: MS)
P%."\OAF[F]AP^<K(;?@= (&DL4DDW&1< ="5VC78[/F;UQO00*=C>].Y#WE \$M)
PWF5XH@26BNP'TI0!L7CC&-GG]@>^;XW,H2MD*G00O;=9VI%9-]J"[4H/(2MSL\8U
P4P(3:7[+/:1V4^NSN?P1+.K.N0 @[M=,M#S%$;M;"L1YR7/ML&&B/M%S B^7(S,R
P6$2+H%*VPDC#5 I,CT"069!1N@5$,L&H@^;JA(&^TVS!)H]\,:)$7E ;6TJU6T[N
PX\8IGT[,K3O7_K8]<4]B+YE-)0$SO11%6ZCJ*]O$[P_#6"#@ML0IG@R].+0? J2A
P-R_S_&>SD<ST)13Z4!PKFW.UL"W/_F-=(?<]]H'D?^%Q?8DQP>#QMY#%&_W)3^PE
P6O%VSA9/^,;^PN,Z\-W>VZA+1.=\@%FN] ZKT.CQ/-F@\!=,2Q#T.1.5]YC.2,T4
P363%SNW_I',?>9'#&$5G;1#Q+M^Q6:J=%OP@3LMD8&F$DN(P*W<6J%BXO_)%=.[5
PMWRGQ#;M>AQ/Z5/BCFT#>.V2[JF0ED6Z'!=9I9Y7I4''LBXY&)0 4L%^Y?-#;ROP
PH[\8^8-M3OG,+L4;M)O80PW858@=P]?E3ZBG()C</IL7OB/)&Y@3#YJ)D05+%.0*
PB^Z.RS;?H6J$#511&"5?-I2)8)/]C#<_P,% <73@:GE-] +*G*5 8%HG'N&;H@@]
P5I*$C0P>>,ZMLPTS[O<?\TK4U4@O@6J/Y,\N]$+A$8@?MQ&%"J&T36 >K5L HMVA
P#5@I2&[_8$\3E;& 93C%I9'%;ZE@7M@,?^C^BZN=TFO):;5+$V]W=2;:C$D?OCH@
P%JL!M"\;D=+D@P)\>,)B @X6/<D^E0&G>BPWF=O0\KJ']K3=9TB0>G)QOKK38'"M
PTB1JBPD:67]Y2+;65>#:&@:%P:(CZ87)QWNUIH"O_;J-=A.($O?P=GZF7CLY;N%+
PI!.X=G_M^3UU\#:QGVW6%YF.(^PN:>I9@V?(6V"63,7T*DQP8B70;<':QT)%,OFB
P/#0",P+[Z\ZO+@&.RG!2_P,GZUU#]5,RY&M_U\;B!Z*1SFZO7943:!SQ8=UV/!H,
PX%F"B3 I60%<2-HD\2^8R^7/(./@(>QLR>G)KD[<5OIV"2"NG\RV&0\%)%KRAY2H
PAX>V'YKX>;JT2+QZ=IN>OY"J"M:TUAMC_6X^H<,-)4>U)(X&Y "I@+*><H3_3)30
P8CM<#,<R$8;X=_.Y^.JFO_%)"F<I\*B,MEN >V#CG:@M'\*8A_,&/E) O,B?N0L\
PM/C#"%@&_D&14AV3NX3SZR6WKI:0(;G@3;\5;_92=[F^'@YI+I%#9A+2<W(I[]& 
PG^.O-Y: #,6F4\/8)A.D0\* ZUZ43\ UNTJC>U7CV&NF^#WA36P[=1HD-?22.&XD
P1?)N1@,=KR4SU@9#]2K^.3PP5+(W@>73=%@JHN,+G2[J,Z[0=&9&E\X4!@X4./A#
PA>=C4&HY$E@.KF%PY*I\YTYK3UK5XV+=*[DJ1O!?+)_@M#"A7*[:\L L !AXB'G5
PY9T7H$D^[Z9$CD8-FM*'1;#>"=3'9V51%D":*3?R)V+.3/<0! 8,WBUW/%-B&RWH
P,6IU@33*+TO[V@$!5F9"7=MHC9JNPN%#YMM#E8'N2#X8J;9D5)K.;DFQT/4I=@6^
P0HBG6,3G?&Y !Q6KK6-K^VB=E)F=9P\4!Q'S^"LY_BX->\@J(.W)-579QGA@35XH
P<$!3UN$&9:P:OKWU^IWX4T>6Y[R*S#$;2?8;,5X+$-UQ*;;(O<6OQL+=!O >D]A9
PBXF>EC(36)>HS/VD$6-?F%/F_'2,!=FQW)G(ARRJ '"NQ_+67W EY B=\R")C!!>
P]/0#@QOX[I0M!$I-"SNV&#-[R'2>%3IZ_K]+9'/02Q[#M:2JKX!7\C+VL%]1VCD=
P6EAJ&<9_Z:> /K_)= A60Y.Z7^0P\S65'-K3N3M5M!W1T1&W9GNR-R.Z7_RQZ$SO
P/^\\F0;IE<!C^Q^L'\?"-..80+9CCC.V)X;H&;!,>>*/.<[EA,V0)=(7Y#K&3S:!
PM\)=#\JL1\EEZ-N 6/WDJ[8DEDE.9?D\X]!PH&4Z;YC:N=DBW9'6NDBT,B0NM6W&
P#WV^HY0-7M^6,J['-(:>%#"4G9V-3^,9%@^8"Y[3S>G2 *,UQR9.U?UC5_6"D'A)
PF;*^Y<(J*8+\]<6WYUW-://:ESV6:=&_^Y)&K-AM^9)2#/X^@R->IK/11;(E4?[6
PH>QGO9[6\F#B 11T-$1Q[Q??=?JDFV]8W)@BW,GN="94K<=_#&QRJD#80J?5VI=*
PN,<55D9)&LTZ")\X!P-5>Y9GG+'>M=&5=0/KF0+T]0 *DY'DKLT*Q7Z4URA?$8_N
PWX3?/TT\4*(WP;Q.E\XKD<Y25B_H&>YVU$!=:0)%D4JW6\'M066-_VQD#I==G"\3
PU>#Q(RDD#L*N35EO'#L]"^K;OQ30=%>^4:N3@B>\*C<3)W4ROH2'6/(Z\;\K,7<7
P!!BH!0>55X,X?9=,^KJIL&3'J8$?E5.2Y_4(>,KI^WX!''QCQ1;^W&+D[1S<'ZKM
P?#79$=B,]8DB0>I3;C4G.-JU<F658*M^VFT772X:)1/O@]]!PM=0+A_ &#G+FE@@
P '4SH)?)D]KI0J>/G+.@)!.@155OG-!#R$C?AS#8Y.Q7&F>V6I(X:GFWR$D$UL2]
P.!4FZ4T>;9"X)I]YVQ$G7=3\$932D,54Q,-5/_NLI1(JZ;$7R:2C<[U:%([_7 R!
P49HB@T72>J]=W\1J)NG:M.:JDU?\68L_S(.->X3UO)C'(KG0>79#GPZJRM*"2V"Q
PDJ^P_@J1_(_?ZQGGQ0E6W%6_V/#%X_(*R,1VB)6"CPNXWSZ0.-N#6G!.+'P0\@!F
P">9R4,(9@."VT>S?-O4!$ENI2S7 I"+[!LLZZGG.2_>\PQ"W-2]G=P3<3E!6[S";
PTUI\0>#S?Q*O7QQ-WGQV2PR7UYF.2RP$>\E:N%FY[L[5D&UCATHLJFA25OY7N7,B
P$TN+Z4ZA?)S5;2$_9B0WNN:SWB^<%FDHXK>M38$&['&-)X9/A(G5I1^12-/S&HMF
PYSA$:4B]"0 Q_KV_\*#8Z<Q-<Q&.AX#8=-'OL\QQ'1O/[4MXL L_2T3<F((C=A)J
PU2-](^ZB,3(^?'G[[H6D;5$IK5D@!\N]2353Z$I11>W6T-*.J0/)4[QC1K1'/S35
PB,"K4&CFN%4?"3E]-5E*J$\'O.+-6&E\ F,&V<0YCZH2/=MX,!N0'BH&ISP-L,:T
P6_,PG(09?5DL +V/'P_@V@4E,'(_M/5LNF[#<^4M%?+A.-^\ [Y^]EC7]814"/")
P4G (%##95G3?.E]\J%,8D]6["F^;\70=5OYF%ZJHTNZWWKLTNA18JH&<+'>>1;DK
P)!&-ISI*6X2BUQFX3:\F&%6\-<<<T2>TY*;VASA.R2UP^IIC1*60%!O7W-]83RA5
PAO%0D@Z+V]#)Q["(O]7AF3<)F.*-8?8=",ZI 1/UY\(\0+XN 8R#[U\/SFWI.?K&
P[VAJS4)0P$-%$S7\$QXW?PDSTY>(XXGW\3XX2,%=L<YH"-&[NSF5X?5Q?+I6@D2X
P40XH,LHW%LY3LI1A67]QA98U(X-5??[FK1E>E"I&)-05F+1&.!,-<6WG385'-S_E
PNH?EW@3'F$.Q I"O.GK?7CY5LRT[9M;/LIDX394SJ%7<LMGQE;;3=$/#"/=D?G$T
PH"#O:568C]"]';N.I&B;Q"4M)SWQQ*56N=<NW7%J,Y+'!UUL:K[3:<H$G [9CALJ
P\W]!OPU$RR^0A6;ONI$T#?H15U8VM9M:<C3WZ]T!^MYUNIU%#T:(&3<>'N\8V@AP
P^C0(/J=8!+/E0C\"GJ"XEI$B%0!O=O\5F>TK2^DGA,#;H[Y^6/)C,-^NT?:'#:56
PE;TY+8*@.)A (I^Q>$>7 ?\Q#_:-RO=U]0[@4N\-S0I:-'LN O<=YC&CQ>_N!RIR
PS*>W,JCAD7*\"V.G6/<31</_6<<JIKK^L-_-$E(_P1YU#Z\96M1D+8%B0%8-K*H2
P0!I-<[J36V&1*H _8.#S?:Z(4A%*7]Z^Y#JJIY@Y*-!UP<M;\E=26NC/=7"J#%%P
PQE7@\D.MR4Z5%E >PXF#MS^G8'470X=,7"NNQ="@G],U4#%7/I[PZLE#H84N&+HE
PTK\P]')>37P3Y:I*% 3\=G1"+58J=:M.85J]PF,H)@@/Y-'%(8:@  5]#W8U]YC8
P3'=@X18[:;47GQ%$WEG@=,>R()40M9LF9F,JXOO'(Q"$NUW?FDL89!6B'&NWL4M[
P4=3&6[M(\D3&4<(TGMLWEGZWN;K5/G#XC)MBTG8)^][C-_V3!R@'[Q<*VL8MB&GN
P( G54E=WF=Z*".5R8HIT8;()Y]F]QKOQC6HP)(0DI^VUFR1>,__BTWKK_?M14\#7
P#VA$J(@=!]HR^?_'S*N7!PH1L76'\2=..HL-P- RIUQU+P$\)4=VB="3%DKXLMCX
P_7F1 .V'$?;3N"_1$+8W #O">>>""5T*=Q'KHLR7-* X?63GF3B%W6KOGPB=/#F%
PZ+C[?MV.AM_WY<OXGLQUT-9+(&OZK0O:_&T]JH@N_)47G89F<__/A1)6J39 N$8[
P[> =KB9A6&++DV_6AE;:3P3=!S#'D7P!U_J;#F\/'V-%^7;2GJ( 'L<YIJ-G[<G>
PC&7VL21Z7^5W.6,.!?DFO; )9[X2NGCJKP$<"'\)*L7:&P7A&Q4VO>3?XGLM]/LK
P!X@0\N'O'\]U[>/YG.K5#@@C@28">K8"XHG\H.( ?A^Z?CW_%,4,";S=&Q;5C%+V
PUU=PAJW+D7 QI>LV#D')G59!>'V3+KJ?Q@#,"P8+,K8.S&TG*4[H*576>E#JUT*^
P% *^ ?*/$MQ@TP9^D0Z7'+*>(1.Z)3K.3T6F<H_R(G6R)-M-9C"G;G2RZGC_3H/H
P1\^+I]K0+A[\1)O2&'\!SX?V\(E+ #NNVKX!P3^#)652;2W 0]C?!\T?QU4>\:?)
P;0ZY'-UQ># =8KG+S*8]V#F:@TN?]'=B:T;(JC:W;4A>585=VM0J&&8K?U?R3&E%
P239E"? 3"C@1]8D7U*/9<<+.0Q#H$RN)E:@&8 6+N36UT;KYYH"<3L/NB6\<=1R\
PN$-2N%CB_AA"4*ZNR_V(0=]<J\\^K/ZG8R,F9XA!!'&RBT 7D^R&0H-F>K,?YAM?
P#J8QB!-B)<F62RR/'K5(-F[E3A(Q<0+(.^TFGX4IW2/^[:Z,3WB1L,(1]H+\(FNA
PYR6F(P>W:!$8&$:UX97R>9..G[4R/ZXOC,%'6=OQ&MA)]OWR1<"? *,=^6JA19..
P>*86G'709X3H;#X8*3II=1-4)X#,WE/6@DST'H >Y2N&MJL<X<@,2Q">'^U;1T:'
PA65&ZVU-?F'P?>(+X$9YK%T.C\;9LEO5),GTKV]7=K?5_E-V4'J841Q4<!-=1-_(
P5R\YB:JH_Q;+I\P>L;+=* $2HLG6U],67=(RS_W-HSC%0RJLI)9\UD^>=KS>-A('
P6WJUGA%/\S2"=-)K\ 5C6?;<'9WK"SN/(RVR??LF]/AK*E(X/?B6//</*-2&PZ9F
P_;C.ZZ*A.1Y&[U8XU17'O#,*G'=(B_M.UC %0X7ONM;D]?//,+^G3$>L$G>H0*7_
P"3:XLI,>#C19I?XAR3(H2*7F2KM %F;3\!PI^^.004@'A,<B/+.ZMCOR^0TI> *L
PT4[26!OUZI[/"$;T\?F0Q<FE9?:&2+0Y!AX;SX+ QMRDM<#HH%.+Q\+(A^5.60H%
P.%9];H"2":_G"!CT6"?N"5?US G&IK3GU#4FT8XO:I"!261$JP<H):%%/BJ%.G%M
P79&V-<+_;%.@&W+ND3)#+UW<1,]<JQU+R(0RITT99+:U%EZD*&_?F!AR8]+]0Q,@
P^:J,U)$%UQKJK2]WXJA,D+J2UY;W4!D3E#_C-6GKP+'763<!%P".N#PRF2Y'M>+0
PI9ONC^_TO;*9W*2"E,,=QM-D44R _3KX3=)0V=G E5^_6-3#"W/JL]$1D$GNO'<H
P>$J7T\215"-J9\[^,\B&/Y[6&FE17 6\"]P.F:AGX?FFRCMOKIKWB/&75]RIX$HC
PZ:W4=TL<9?/VDA)6,C\77L0VR<"B_Q26GY>+<A<I_%G?2]3&\R+3SQJQ6H5>K,;/
P;Y-74R#%$?EQ[*>;^4 >%^PT0'KHYF8*JV?.SDDKWZFC@3XO>+QGM@YRVR?R;M-A
P,_!V(D4M$&AKD0EB[3O;-#%"?^&'DMI?WY=2\\28SB1E(LM"PU\&8!>_+O*U(A <
P9X.@"#?7SNDN**D1:U*=413-!L'=#.MJ=M,YW,@F.3#\5M=C#BV<6Z56ZCV]%P )
P=RE2-.>601589?FR)0B1;/]%'.Q-&#].K>$#O%1R?D"FVZ=$U1FFYF('?1'4@8OP
P=J! ><BJ>!7'1EAVH</J8&=P>E^]#AQVGP/W4L>I7HBU1S^DQR88D5WGLGGIP3I/
P=%Z5XB4_DM#A)A"J;39I%Z[0-?/I3/0M0'MI5*DET#^^50'?W8M]GV3LD=FW))8R
P'>#Q5E21!:0NUFQB"OKC>77YU/Y*B*UQ21HJ-1C[J!SDQ?GWY.[^M"GF6-:"'_3#
P>VORANX#"3\F_QFWIO';68GX4];O6L6ZH'3:/WQ9O3FIBZI3LI]H3=%;(P=,_,7#
P3BYRO7;5D2DOY!Z\%RK=IR-A<04V'H-A/ A4<8VUO@#+##X</*CY)L8Q\D2< TO\
P XU\\P,43$;O[J6VRWZ78';/5M)$X*2[7U)I.B:KJ  'I(5%4D:5,GOHX?5P#L,M
P;IQW=47.@M-2XKB&Q?2!:K/:K"T2K'[YMM:1BA/N,L0M;BFZ\5E<Q">.^NV 0^+(
P08AZ>RW*:5 :O%_/(HN/8P?*66V -2G5WY>#P'CS%F9$R?Y=4]1VW21!IG$"%NY2
PRJN#*I!94\(8>'63,\Z\,5&=XG\CE=]^<[)!>N&M\VA\_C?38)27KU%F3K;5F\&"
PWV!WGA38I8=-TI<V$I#Y0OY"6;7@VD4PW9=!,3HU&$N>9RF<.V.$D4O_<32I?;I0
PR:X,%5X1<RJUPKO+QAZV=E(*),4H8[] A9YDJYF"%7*!>Z8XDZ0TG S?!.>;=EGY
P$)L2[G*&T)EZ"+_,N!2Y80.-3C&D94*UJFU"F2\.-7<<#,CLOZM_#XRJH)LZVG!W
PG!8?NE4MMR3!O<7@1[.()MPDY;O[(N\ 7Z<YU7L;9X?BX(!4Q2LVIU!A7(I]?4'M
PX6"4L3]YA#:+8U)OVP?V4*)2ZF&U?U*P:B!!";'9>292'2A&G&DNZ6ZTUJJHWQ_T
P[[RP!WT1C2?/,8>^"$IU?"G"H$JRVH+F9:(4E>QZG[L%V[DMY.V:5A>BOVGD4[F@
P?I*XLY@U5;C>NWE*Z75O?X^F/II=(-3A26B<C<KC1<[?A,F?+7\Y)"%6U;F1< $0
P1_G=Y7H1J# 8*G26CA&\(ANG,.)C(%#[A0'I[N2XPIT8=X$!O^K3?G;LK.MT\&#<
P)']TP1O.>86@VD,^1/Q@4CTGWB0(PKN:/%>I:1IFA\+TNUB@^LK7ZMFIDO2[H)V<
P==#7A90"Q4L9A_()FIU[^^6<-3&[Q_7]XO0NF\7C-B!POL.M()4Y,/BTM5&#%#6D
P$?63II]?B8FH>/3VJDGW!#9[Q5-;/-RF[7E-(HSX)O0.M'<<M* 6QN*XK\;9-K=3
P]-X_0!#-4GW,,U4)L0@/L9^ZO/(DQ^J9 3)O!("/L))9JL/K>S-"_FSDIJ]JJ>H$
P3T"[I)>W)TA'[)8XE(Z.V7[KY$EL8*N@@/1M'P@4V?,T<X&!Y>Z._RLP<F")7T3A
P5%K=-T[9 MKK+H;IN,0;2AN@C@/:2XUR1&14,B+5J&)#[V9W0D_]J:GDP(DEE)27
P^7/7KZB=MC1\N"&R\OY8!F[+ 9&#>\V5,C0'7H'O GZ*HE/_+Q_7")>0G)FAO6^T
P/F3<Q/0<"TZNQ8 ,H5$27]<"2UP,69AR%_YN/K2U.)Y(KD1#^4R?.QEU$>DT*6Z0
P40'D/ +-/([QG8:K*9+=\T*'*">M^=2BCD36-5YJ&3"O9'41J4OLA*0-\QM<IUS)
P$4#3EFW3(/6Y1A,ATB()*/>3LH[1T^A=L=6Y?:__YG721/N?/Q<YH[%].B29)=]A
PXJ3'!Y= WDJ0KH3PT<5)ISY3PG(_<PT:#Z8!;D-\%45";WM0RZF^GEWS89L&":.[
P)CYX6F[RH(\A:KXO)"VJJ85X;"<2H]UMI7XA0)07\H)F@;!&5?Y*(\ZF<,<D;U^.
P>\$<0]N YLA=G1O;:$CC$<CS25](F@</C792X2/E0.M>L.815#)MJ$\%MUG^S>8%
P,;;:U)M5-V,%BYG$WWR42$[U>"?5&/@P5J$JKZQ<Y9>$-)!$Q<2GK#0F%WQ+@9YG
PM67$UDT!(B')@MS3Z LQW(RNP>+].IS3UE7I47*MP'*><&Y?0#"&JY+ME3$&U#IV
P?#QQ"H1%FU@??2<WLDHEF[_(L.&WVUD:ZT=A>IH-N^HC_SW.R!%3C20[E5K($07>
P#<#N $.C6INL3O^$8AN+;@I6W)I#BM-V,/02#@QR8&9:P2CU=U\)$UOF W]:[<16
P,L 31"24N T)^7K<VZ%:X31W79&#58T2D>E/A*6LNQ^6H:\*U1@GP"&:*?KWS%]K
P*+T+M1E_]$>6M&CX:WE/[*)]#@E7 R?(06&A#LBT8:60S,>B*DK0G9(!'_%\#SOU
PTX(T*?&S K'?)30\12YOLBC:J.W[@OX.TO0B,Z@NG*$3,:OF3,:L5BC5#5?E5,;/
PS927V>*3(0AJ#37C\7"\'-YX<&4^;$O"_X\+Y\B0.F<XJ.I+>/G;\EJ+7)SF6KD;
PQ<IC>&HBOKW?M4 =.S(- &B\ODZ,?5(0U$(_#?:('4]<'+5VJ35%7,LU5KFF%<3[
P=X(\Y@R0J2K60K==)IKNRQ-UN!,BM50X#SZ)34;YNU951U0%@J^FEHMYAW>]:SUF
P]A9! 8'K2QCW;W93$*)I\6UZ##&*:H&TU?TXHK@,3+SOZ;1!3[C8F@4-I"&DY]4_
P%R;A<;'3B;D#DRAQF:_'0(@]W/+@ H#!@F6F_<UTIW(;'E4D5_I>F[S*%Y7T" [<
P0Z';>P<RO!D^G^AI\,7&@=^/%5BJS#S*]/X]\V[@!9#P\"A*4S=X+.L!> JS2NR-
P_Z%Q;+&FGQ1A?31H)&96ZD ^ /-7'AH6 [Y(S#^[E26X*X!A^Y$:^H]ZNU9C[<"W
P\2Q$-()DWK\@3:SS1;J&R?W"#_0_=M6E0FZ!6_<L;-6\55+R>J0HFF<:*G*AW9GY
P2AO\?&(:K<9D^A+6/)P'-WP26A2R":4*!EO:P0W<2(?LW^[5GPU:K;YHDM3?F!2'
P<4]UGT7:IX:L([?>0Y&GWPN=QD$V%%>T,VQV2.MK@X'#(4QIO4.LRL6QTI:)J7W,
PTVG67V]/V?T+ #\: *A_##ATHV/O>!XLAK6J[!5C987Q<RII01-=6M2XP>FY@+]"
PB"%(1)W2T3I,O[SE;43"N#B4%#KXC8:YA^&-65RM@53U)H/D'?7&[XE^_S/L!4%Z
P/BVZ=S^!,9U.I([\.#V"MI-N')_Z;?^=U;E.C?1=>]9ANEY;0))C;F.F=J+US[,R
PB]0+WK%N'._=V1\C]H@5F=> $R#0):%2Q'7*,<DW855<P*,9&/H7,&*"P[%$ NQ<
P@^/9C)>'ZWJJ1,/**!_+LH*+U9U(BBHGLEEH2,(H4CR52YVB79Q8)8-_"=6 6/RP
PI%0<6G0_A5S#5!2?FQ G6EEG3<A "=($%(DD&K-B3YN3BN%FE/M-X9J65JR.<48Z
P?_MGKT[MJ?KP8UT**0)*V#9N7CB+VW73U RM.@^L^7!QK5ZE3_FTT[((DXQ8IB'K
PGCDA(SVGNH[&]%O.3EJ)FG0=X73Z"DM&UV4=4Z&&'O7T$NVQ-BOTA+15'4:\/U]+
P*4O>84J@?>Y[,@GZV6&ZJ92%\4)^POBBI7=K!NZ>[#L3>OK-HN"9;"R>4] ^H8O_
P8;E6//3P"+Q-<?;UM(T;W&V?GY6+)<?5@(TBL_Y =.I4N9_AE:5^L6]PK]A>-D9%
PL+8%G!W7>3XL/>&'QJ'/'[5?D(:J!;D(('Y<B$0D:8&4<%QF\)@:78LVW2C'!US.
PKF"&[JND3@OB*<5)E>%L&=G_79B4^30_M.JD--524(KY.]<P;>-,,MKZ4\W:ZI5,
PH]7CS3%CR[4<LCRSP'TPCXM:L@SCNL5\HEX%<MP%V]1W=%NYG)70B.S+LK\E+"_[
P)6 G [%=6:Q5KHJY1T3%^UA>HPSJ>_J(!PSZ^<;?+%,5=,%2-RV_*#_81-S-JPOM
P*O^<ZAD_%PI]9'^IN-GLXQ-XSXU.DD][0G<+@?Y40"_KBJ.][@3MHU[FGLV-?BB 
P@QCU-SO+2/!85:.TH\REJQ_-!D L/3\,%4OJJAT7RC(^#'(9IO#[XXXA:].!B4GA
P2TI-X2QSA?YFJH)M?_G%VCW/];DT"H+I%/R2=95G86;91$HMC4 4#>&RPK%['<8*
PC-F#QIHX--B.RYDG":3H^*](IXZ:E@7]\# 76X5L7@O[":8%GV(,3*)@* PJD0<3
P0ZO6W</KKYF0-_.4D>270GJDV'XC=MA.K:OU\' KK,/!-^!?GJJ.)ZUNM])CP9D(
P.T?=&T_E8;!5VI"2L]+>YM)5V\MR;B\V!E4K_0M&@VZ_ [/D+US@+KZ"FO$5<Z/'
POS::_SHD=;3T\77UP)+<U2^)VPZ9UC-4;\6J*E1&M*J:V'=U<56G@F1K]]].#QN/
P<T6X3/0O:DB#G%9Z@NYJ.9$*C?1G*NL]DL";<&BD<V+/62[-UW:Z:$^<ZPEU*XFJ
PI^*&Z<P>6?0TFF(]H^?_#2H_9KMW/L)BFS%4/Z@#B.'K%8_-S"_4*K'FLK?\U^39
PLB,P.D(OO#7R95+M8%=,.D)_KO$LDSN6ITQ90!R1.<3/IPV**]($<B-G[R^J$=LD
PNU-#I'<QP5%[R*0FE)W/<P]W'-HGB*2 XLENR_)O:M#4CZJROY,<',,=U.0<3(V<
PL!/B/LFJ#@:[:PLIUEMC?-)LQE_Q(JP9IDJEI8=;W<L(A0\-&)N'+L(C8O47W\JP
PK7$U7FYP7A[$64[)4QOVP6SWA*-^R2^46C(EG1BCP0W,S'J2,DVJI/WA[W)\ AT!
PJ2]H:31D8]@K[HE?!%&'A!3 )B7Z2<@VS2H+P^2Q9:#U.@U_$R74QM>5$\PHUR<9
P3B\.H'%3FH"MK',#@%Q.N!"-0-EZV*LG':Z/H-=F#V<(&YX9DPCY.2.D]Q&N*V]'
P]@D-D]T6"S,4.4#^Q F.*O D3<[F!&Q%2<'B.7: H^$U-R6#D;F# $=9I3\=!]5]
PXAB@9(H:MY4K&U@63R!R8[]"1;C2JF^B-^9'?R_GB,Q)V5/9))A.66L9%- G^H^'
PVYR]RX X\N $RI&![2#PT^#T?C]8$ZR_O4+)]O5.+&:KR8;#R V0Y;_M09"H=4K&
P7?X@5=/4#!5P_8XZKM/KY<SOYIX\[FP$B$:+UT6I=HSS3!Z@UI '0XNSGEFZ34"(
P6S$<<^N'&R<RL79W0Q+,5V.N^MQ(WU3V8QO6G"ZENM$^8R(D%N@"R\UK3SSB0G0G
P\ RI*CQ3<6\4]9([#ZE<\#*Q7LS:' 9VF^US%W3U-->3>_KN5F'9B-]U!!U7GQ&J
PG8<>264">%?@ AI+KYV)IZ.:)KB6M:^(4H_7'@(]N2R[^>*8IKA>^!UPMW7"JB,C
PKRYJX5(QXNA6'%;Q93J-[O%=ZMS;HR;/Z9H.PU\&D5%@XKK^3'$PD@@%J&-7,]C4
P$8?GX:H'6>C7PSA-E9I[(G5Y3>_-*+6!=%6!95W0ZRU-E3D/PWZ_F>,_#RXEFZ"R
P4^'=C_;7LGX\]T2%X1Y=P;?=B-$J@Q#CV;VL1JKGH<RM@SC9I@9,=I@GQZ >5CF[
PC8/A[ =6R=@4(A576I40*W69(E167<<Z4B)2[KJ??LX8)->#C0W0L^:CB#A2C,@@
P6,I=*6T-MF2LAPF[=S-;6M/O*F^SY0&@EW).K4L.QGGQ!-::ZR_D'47=6NA$7/[V
P4?]3G Q]4?SR0'>;.G&6YPQX@E9TSJ!T=FE=8XSH8\:P+:Z =<U^UTY.DU=C82'+
P"R9-"!597VMN:W-7%5%TE7Y,,1/$'2./D"7F[ 41@ SPEQ));YCP:AYXNKW6XQ3#
P8S636%4X]+/-=[=[>M'=!(&]UHZ^S&,P =;,Z+C61M6L%FR\2M(F^ YNZDL\EG.>
P5+H6&=17R\LKQK!!&A&.^;%APW<TH*6<XF6.-!\9GWA-#&M!;N#K4;V%Y)Q"D9V>
P(* N5' %JJDL@6986X-O-8UTM;V=["\]6UL-NII.ZF[]Y$5KV5VC3QH59)83_TC<
P+*-+ZDNX!=U[1#MBR3Q_3?M%\DIZKE=8R%VI?8PB_9*] <*VZRPAZV1^8H=B"I!?
P1 5[<QM8D+;[1!J@?P5GH57E]@RQ-I[#]=:8A='>BHK-ZKE3X#@FF48E8W!7K8HF
P-*_U)>S+<T_@Z*J@/VW7-]RZNMZ;*/%^427ZR;AV;4#X C" ?\Q?%;DB5;(7^Q9X
P'DH#APCA?EOP_YJ+S%P)(=.4)S_#)A3:[Q<PV\]6%BG2$!3)$,PD\P=Q'.2O(P$^
P[D46Z]+QFJ,#G]H.ND#L69-P^J_VGXX3B><<H40H9]T7I(RUW#&W9:3UF?XSZB:^
PY8ZU.!+ACRWR@W*'>[1XVO:@/H@B/? 6'3J1C%]I''NH%<<@U7^>2/*[TC[M%'6[
P@U[P=>:-:',52,3QE.F3OOAC)LFF>*;!5Z1+*A^\;;WT-OSD&+PZHB"DJ3\"G< $
P/-'T#;U-2E<1Y<I%:=_+JK94/R15N=@+<'/0*D?*CZOZJ$-SY/ "*D /+EO+N5"=
P,O@[;X/Z[M^ZQFG6$I68,Y\+]6) /.M$ W.IG!I3&_Q/F46QX#0_FA,/^'D^Y;^J
P7@L!NXPW.2(I?.]%**L+\N-DD8!W36Q>_V4FEV9*Q<:*[B&A[:52GLVCV'IZ4L\%
P<%OMD,\.*4UG]3IMUX%$F]4XGIOXBT9SU3RMZ_)MVZU'<59>UF=F/7[69:)(L!J#
P-BBCE8%:QP'9'V,YC?'ISSC"Q44 +2'7[:T<__<@"%!P;IQG#&) ;5G2_PZ&VWHV
P?G#"1JSH6*]/PA7] S.XEV5\Y7>E0:I9>*UZ+H*AXU<C>.YT]_>P:'=OZ$GEO8B)
P(O'>:N5F@D6Z2^]+HP&'=V*SAD1:=O(E@=9.K=.NV!DQ[D0)K&BNG3*=L-PM"]3Z
P,W3Y8W5?L-KL#_OSGX6(_&\TMMSE+53*.]<:Y$+GNL.$-#X"(NG0F$1X%1W;>&2F
P-Z&,N$2;:BX6AC76$XJJB!4?;H52&C$>8*A+V(XIOW7>27WU3J,URP-NKD^$HS7,
P\,DNO,A&,8#OUE.F 8EDO=R63QMFS+-)V@#/1)XBNP_H7CS,_,PYG6)*5]9)CB!,
P6Z8[(4R@"E)%E_ 2TA&WH4HG[35WUY5N&&N\ M@K -:SYQC83S@"&!+3W.:NM-I>
P>K-.WI.]*9FS391B:$RYG9.8Q0H0DB9DAVBBF"$/997>6C/.6[5]S>':$<S4@\\-
PX:A.;5XQE7B:B\=I0^(O4 3)!.BK3R&91UC-N]_UX4;T%*SB4G!,'BF0CKK"R*:Z
P+#RI&$#\?LK4,"H!32SG8*4KXA0=FP"./6+N__A+>$&2G_M6NX 8))RYWE6\&8\K
PJE/_(4Z.R>ZR!6H_=U*IE?7_/2/"IO/:P9X@3QU$MK.F6.W5:>((ORRCS!15!7O"
P]2L:7[ST"(01]683L7PC3$65/Z934]Y<=?N%=J)SPUM)@+]FV+G@9@VP9/UVSQY?
PJ0&2T!^OH5=6V9R:8JR-./W\=[JJV?$N/&4!U:A]\\B\0;HSZ)*W"4\<B.?&!?SS
PY5BVAJ[RC!&9FLON-41S[96F_(%Z#S(DC!?'R<CK34<SO[KD'YQ#R(XXL>\O'SU=
P'^.R,Q:'UCII:-B9$/3]A=LI=*B#>6P4P,XA!L8Z1TD-<CMA*\C*X+"O,[WMO*C>
PH)^>,GQU)QWGHB+:):9ZNU63T41]?S(6+2 +("-&=M&=,MD]FU&< !9!-Q0P=O=W
P89PA,J*V,NE.C5B%/'M[ E 4^*9P6XD/\YASP&J#SD3)B^5_Q/PV+TO**OOO"VIU
P!6T4_"#BN=?X=;_M:(R:5#0^A2@Y ?8HJ]*"6K#V>-L7KL!:>]%+M]3>-TSX-R1^
PAC:6M>"YW4$8-L5 67!1<M3F:"\&CWPO.ZD/V?OZNJVO^ET*VQ=Z/]=)1*L_I$TF
P97#A9_^S4!=(DM$- !Q.QJ9U!N-N8*\G'1;2<J7KP*;W[U8<F<#:N8?'FL<?I*._
PTY^GNMEQU*"QLBFB>#/B,%=R.1QDJM&MW9#GM"-M]\KLK'#>]TWIB%]V$X$=&1P4
P\I!IA_^#-ON@+G]H72LUQ\+F9ZE^TBM;"6[L+&R*$>0W=0MT3*T#2PG'M98Y'+?@
PT39+\]^A-Z:N$/( W)D+ %WIYROT=;'U)F(OK%:]FG'IJ44$ [:&*BJM^M+.4H+0
PT+A>>[52\^TM[D375 &Z)G0^UE>"R*BH9(,4%C7O#9Z6T(DB?9VRV'5]@0RM45[;
P5L;1,N0YIE$Y+?EE5Y:2#0E$62Y"\6$B>!M!6>3.X17^%/B.B!8W+NKC9]=:XVU4
P73OU>XW,^1']$ N.!)G/>JB0WW66A=89C?+M+JYP 31@$>3G;#@NO**8YSWP*T";
PFI$<%-4@,#<WMFN(Y?N<?1@X25.+W%\VS>RPP+@!650Y;Y/^2=FIBAMXCRS<.;'F
P0[\9W6!B^Q020K"TT?=;S[5]UV$ /ER"Z)JC<COIBA@7GU+VTR\YDIR6%K5LMT9%
P-O[SD__61V% (8,/(N>/U4M8VN;9*ODBMP93'=/  9\(L$!_1FGAB*]<-+D9JZJW
P<"\KM?]#M" Y*A2[GTHGZBP_"!N#A"7\[-#@X_<Q MY<5D0:RRIFAL[FP6%=X^HT
P";#C8T!V<AU&0(88:&62==_H/<:TAU.]7FDS;A(@72;ZI.F^<:9\*VFG4<)IL5V$
P.S=XE4_:P+WEB,$S#<%:2 G--999P=8>_I#R(%\5\L']JCLA^%@BZ!F\_*U5D8LH
P]2[R,F5CV"$B3)XAH:8&$_.&$>V]8H%@U=LL+5==56 :/W'LT5\K"H/O?2P+6LG=
PQ+VD0OGW"[B7. XG:#@W,@4XL^=(@ A/!W9,*CN2_P+X%SA@K+2;;IY,_2&A.OI*
P/>%VCU6?!L ?70>]A>UE<2C'CDP#<=D 3>"8#89/WDYL Q0;S19!VCN-X(.U<\3&
P<%V!2/;=6GP/+M6><QTPU&Q7Q]3V$OZ[PH$J LDJ^I?X,\YO6L'\H:?.YQ:,0%_@
PF$-\]MA[4!G&]4XHZA@W.SSSC\E32:M?U_"\\6M=]5=C:V2;"-6R:TJ%F^D9? 7B
PF"+BOD/O<>9.RCT!,<F0)ZQG_B0/JH72EMME PBAYU^SCJKN9DL?@!(^\#@#?,2'
PVF]@P+\-J\ZTY+O_Q#K-7!B&'A1 D@HFF]OB5) 93-B7LJIJ444+*"<@+,/^CV(C
P7=8*O"T\N&,EE>1P%.BCP2/9),1D 6) O,$@2GTIP>RL#0)$+/R4VQZN66Z%##?5
PC8I._,.);"+;TP[$-7N'#^E%R#@S4 9AY>5=-0=31<^,JN+9]P+K[Y@H;ZXA4<ON
P^)2.+<37)HBWC:I!DS5$/7<:]7#]*4J1.J/D=_!'(:&T'=L(B*G6LHB\ZZ>;>/:2
P/[>9'H$0%NOO /Z >2"D3?H=C3%)CBM!XKN=ZR4T\A,0*P*LE@&RJ5HI"1_,'1T"
PU$E5HW6;7 [V>/>3JNI#LGSDHN9:I3A5-:KU?!QNSVS5FCBK:>.^4O+=GRJH$;5@
P3UBG3Y?#YP<'VK/^DK%8:5*1N!K/J*9EZBEV_N-RO:P-F\_8>Q,,!X?Y6GA+VT,A
PCC,</32\"^'  E#:OZ1[.>> ]&Y-[]]L!^+:;IN(XG"5_[IHP9Q020Y>\HHP5#U(
PG,O+Y"C4U+)O;B!92Q)E/=Z)C:C&4/XUC7'7EARX.G(&:O:J_+?8?R(@[4+_EU2%
PZ'<YOGB>-80*2#@*]%;HL7L8U?[5"WX(F\N-V4>P".M:E9#*I530$D,(4 [OA[E$
P5U]S  W11:ZPUN18P;<_JM"Y2RJP]B%:?W\'B/L4>WL"]UX[+9<MS]UKA]6J3#B,
PR/T+W_,4A^Z";F6'O*YOEO!& 6@M[(GA4--4X;!&9)I-:D^9(ZO=5L-[E*^4^9;M
P%9)N^6KQ-N8MR$TM?0*&B,Y=]H-YFPZ37Y@[*D9FA[+H/UQ-U9DYWB,\N!*@&TQ$
PEO'T&E68*RE)6&3HC=$;@=.C2X'N '_($55I8]]8@@/?FZVE3 PO!;0(=E[[,L5$
PU;(S(U434:T63,8=M7@'P$!?:AD=U:#,2 \=)J=)&P+3(N)OTERM<\EU#@45<G19
PC_$ZE'2T^4856S<JJ"T(-VW=^Z@LSM6W+@O?$N<E"D29!VWB78^AA<G-^BB1E\A0
P=)G?6T./V6A=G9U&4&CAE;HKR@8/IB9YJ3/V__AT??D@&T209TL*)U36.M?Z9JIM
P=]ZU?P2@EXEL\% 5I>F[]YR"\?;)%'JKG].; :]V]3)@M(=].1 0RIE)S1VMCV*"
PYT!6!4#<5J+G&E-3^$E"GEYVQ)H.9G>:\D.'';81?E>71-@.JXHG";2K(:Z.:0):
PY&5(U&?<Q!P[+/A^U R^$0JZ@^PBDKLMX %RIZYM&[F*=XFS7PA*9L25$ATFQ?J5
P5=\*.CQBD:_HRU:?@;&2YQZY3*H$V8GQ2%E;(*P[D))6TKC4B!IX&;32[>WO")S_
PF_45'*)A/Q^E.;R4ASWM-T;BY^8$C2>$4BJ'D2.<<LH2-M1U*>U%P>G.$5 L>I&W
PD6EWLWR$,^,_18E;]NZVJ6A,"J_\@;30;9@JFM32F<GE2^&UO4X^V&^@8]@+8$]&
P:+$44J8">HQ0UD'#Z?S5?E%.VW15.-57@U3:OJXI3X#4,3%?[0)9C4]JD3=@BGND
P:RI6+M9JV_.A"080&[$]<&Y9K\=%)KV#05_![X/-=7MW_=7LIO@NX:)?0675M7X0
P5<$/MECV!AL7&PI.\\Z5+FPZQU?Y:!FXXA8)Z6C4_&4QB&*:M:>ES\E:J]6OQN"Q
P59R9[QDSKD(5J>V-(^>I;SJ0@[]\DEWXIG6,E2*;J.A!XXCF8(28R2YA]EA&KY=.
P6A"#%_"-W6:L7%F>LU.M9W5;(-$GRM?7+E[NKDUB3O5M.S#MW VRA7'1RHVP#;2'
P%6-_>5UD,LEFL ULXEF)(*#N]4*7:S8CS.^:W8J GF76Q.<RO3$X]*1PP^_NB=\0
P78EKD_&NE:/)^M#$$)436;G.Y%E,&TRW3H.3CPK=)9_3[#TH8L6\,FZ32.=[M\C[
PV9425F.%EOR%CQV6)_GJGF*^2(PCN9<$'M.UY,3SIR>19\VCINM>;F!)C98J^[?$
P -D)E]#KY'Z:" ENAUV-VHY:7J+>AD.FZTBMB3X2<'IW';Y J556X@=SL17)3\C_
PCDU1_O!I;&N^*^*:S^9M9L?CW5B</6!71 A3.7%IME"?I80NSO6M(*ZT3_MO=7<R
P_J<$1U;-%6Z.K]P=-"D\./,,]F":VW14#CXV8K%+ADF>:2QLS5B_0(1]0: \4 8S
PA0M@HMSBH]PV4'80NOBC', CCU@!LV-^CY]GI.T43JT&9D Y+$1+IQ\+%+!=SA5W
PBT!X=#K:WU3*YOJ:0Y<RF=)%KTR:C)16*"VH-<4SJ3&SVE\TYIH)3"V^[#WD[^OH
PLP+0&B30*X3\)AKCOWJVXX<CW!QX/B#^2268RPRIJ!*QT=))V)XR02(11<>9JO?Y
PP.:Q<W&!KSDVG1&W@]NXV+,(T=2&@$]$?+@A.LX8S3"FK!E^FEL%9!OHCL)E@^PM
P5"W2=?SEPM1%KJG^"4MORYYZRQ"3J_<<3^8_D55GN6E=M>\=XTGB76F&5)XZJL%'
PDPY4/IW]*R!=/QP'L]ZQH7CI;)<^:1(T6I4<J,IA?)4W>S+^!?=1W]'NYMCW"H3P
PL7X"R\#)$@--15Z?YD?><YO=QMA=\4IG,6ID4TLPUP/I6U#-#&?_VE2 ?7%3EBCT
PF#E<;NN;ATQ/T&XK&!$ Y$%""0CVN_(B=6,V@*2I?L?5R]##91DW5Z]&>PU&,+NJ
P.Z29R3;HONHO] S'K\@;WNF[A-L4*I"<N3V)H^IKC?!^>@=7SA97CB9--#* _]L^
P_;X7WLR'?"0B^F^3-3R#Z5&G#7\?WC65M_0&@TZHROL(U1%?:0T:/L/,#RK)8J7J
PQ@QB#<"WBRB84$./WRA#SW3BIUI?NQX@X7/? @X":R5L,H-)XN#AVUD"MPP+LP0Y
PQ.^:O*B<";H$EVQ'[4NI"18I@U2Z17(WB!.HSQI6(8 F<2W]RGY,9]#++-,@'WW 
PMW<7(U0?L7SXW;K#GC=ZD_AH-$SPS._%'+2]W7+ZJ9],*BS(J%##9K5/:PG<E#U[
PK:$A"%JTM!L%VMQ;"_&-X%M?>'$\"X;0O NJV3*PS5RYX??'/](K#CV8YW\A4CMC
PIP"M@D)KK2MP'>XJ\CL'4%H 1$HP4?-O(N(2JIY@ TZ4!'YSX0SVI^ 6/J74P9AS
PPE#XT:B769.W#+:R&%8$CB+SW1DHN:128;%N6,G7 ;)&?//1Q$:V9W$ /&.S(;@$
PZC%IQ-,K&.=VK$R]7LY42D,;1 *RT*^P1^NZ'5[04K)AY$PQA_JYM]3SVUH::%][
P:((9 6*"]5\2:$BGXG8$!<X.IRX':994]_I6P8KL7UID%IV/FC%"5)QES<O0CA.-
P@L<VI!"$L2$45Z_GXY56N3)ZE'?+-"J?]Q_L.;1]?70AA*FDC@DZ<N@; M.9[[B$
PSO!)$#*\9'"8X.*LKJ!)L3^U,ZV33EN8%TK:D.VVV&!X'OPY83/!@-(7;@2-$<78
P:%LZ_!;R(BM'X+3+/U:B:RT//?=G6!\*;@R64O(Q>1]6<-?)([Q_R'HD?>C49- 5
PH5*\RNF)A]"R+X6*3BKP86GE4^QR#):ID&MQK/52SPK3+B]7E((*SY<TOIQ;3X\5
P?3]$+F2]D!8>?(*$?[,$]4SUE#J@@QW@IU\^GV>4Z\$O YE)V0TQ:E:^X"OSGYMV
PI2!' 3-O\<36VHV$^4F_@V [Y6,.S7-3P$2Z17S$2YN!O,F%T(>YR!TW$. \!U[I
P5PUTH0'Y1H9_>;CO[77N*?BA ?Z1.A+X34-5A<21:MUH:VS=0 O:_@%_%?7&I!Q:
P=<../K".IG";<_7/6ZJIX%=)2H"E@2^M!6)S*#FE4;6QS?X8.E6NH\?(8:F_;#WL
P'FF9!R/VS/YI424Q#)2VK,4^EB'.5J>;%A^=E>R0B.B>&LVB>4H0$>JY@T/EUK.J
P*@O/]M/PN8C>,(DX4%QP&2[*Z@!;_5A2!VP#&-WPYO_Z"+XO)!*G0Y:[=MQEQ@RO
P!KR .3007H8'9U7(&;YEU-QZX[@OZRCW650,1)C/WV%QY"0 $A=$R<9P4'63QPY+
PTW ,":A@M_O7OS_-A#O3 6&;!<OOG@Q0T3!J$.LPD?+( %\CEB# 2O*1]9%J.,W#
P3?7?I#"G5\[/2V.C#N>=.I6JRVAKP@Y8'K#,7!*S("KB<S\1_F>W6BE$R_?TGQP:
P0FX#?6H_Y_N[:257%[4RW0.SOTN-,KNVB<%[%%#^N\^@_-X[M;\BQ3+6 =X@3[O;
P5UYR@H?8/_0H-]9W/G,-)J)?UF7'<\V[)!C#NW:LW[A+T?_C-TSAD.B=RE];S_1C
PJQOVI +T)+:HF0NNE'J\%!?'3>ME5V#882N.Y%A/S_4VYU*R<\4\_N>#IATWD6[3
P=)L,:<[1"2M'T*.B1FJ?+8?+30THL.;*O: RVJP*QV5IU]'J9=$*.[1-)IQV(9LY
PO\%!FT4_M^'L\P72SUL-+:F6]2K*IXO%3;Q)&/'7A5W0"CV$=0^ BJ*EW!O67.PS
PT,H&"(W;./J<3QM_SQ#T1*XVT[XX97-< TXEO_8[]</SRS[;!-TC*Q[%P7(Z)T!L
PPOU 3&N#[P8"$XF/XN)2US<5U[V6-@_JPDN5%,$1SZC9O%MG^^"9/L<U?$XQ]?XR
PJNO!O0[]W6-ON1-FC@0<J0-,$7=:,5D,?8IN 7Z=YT>3C0?%G4OYV+9MV 0 0'8>
P#1HL0X;;L<XFF27. 'Y-3]@7,T/0J!;)6$-_[A.[NUQ\#SWKQ)5C/3='=_^C&^_Z
P#-A$7EHDP1)_7<"(JPDQQ<,.K-\ %Y*9&J#6"@3<?$N06( GL/K19XLL5"7_CNZ,
PJ.)?_H;%OB[1I,H@VA1BDDGS@KD[*E:: HY(F>:<7F0A)$Z3X3!#B%_D4"U1ZZH5
P;62,+V>B4!;=-FZ\L)8U5S/O EQF9S%7,!Y#8%6LO*!(6>\%02249PPM:ZY:QA"+
P@/O5N4Y[8CQUMOR+E1 &SV"(>^KSC'+H=K.*GBSF&ORKI)S"D#Z-!2C6PCRP)5M,
P],8FXOG3![F?F#TDSU&AE37\9_X4UPY%[1!&$<S24KB7>RU(^=07$?EH<WS<';(L
P!$&-<_3,_T-6)<@).<(5=K$<%*T)2R@4R;1#T($"29WQ0':6[[.CZB<,RK 9IC"X
PU;@^5F2K#>7LT/?/"O7Y?T/G-"](XM@AJ-DL9.J7,TR7RFU!+?]H0$H+,\?-5P;O
P^=K'/'QR9RAP;M3QLHW-'(UW,E+@!+#)D [MUA "KDC'JX6Z+ZDKTR6*-KNG5PT0
P?JM%97GQ/,_='M<IDU/L.VNER 'JP,$8E) "C)#\."J#Q\<]-J(D/58:W3;)LHC,
P=NT36V2,_J0)Z(SXJ&)1XO<.QL72E1-.$]=!133P[X<O(K7=C\89UT5%Y-TJR<SZ
P2UIN;%2\"@]WY+JE+4&9+S;H#EGL8K)#F^T&%RKS] >(!3*HCR*^G>6^QBW:FB?/
P$@\25=:7TDJ/DJT03*=F0A*T-!OMCO]GE@;:Y'ZVD/G";<"U&O,%!A.FMF(&V1D,
PZ%AZ @A1K5R%1L?15>,EGK0WV]^*H4!P_]?,9O51ZU.TNC&G8M,3.46P7I?+5O]5
P%):R@"_U4N%.?Q=/_L^/4*,VMLT.N%4D03'-E,S#H#$FRT[-T,?7?P;,$9#N+T)P
P30$ V' [S4:'N.'Q7 V>$F-HEDBENB7CO,Q0$)OU!,+O\; ?+B%FHEP3<5_9>&FC
PDJHB'/^VP9M#K@LA?;Q[&N @!B2'9\?[JGG&4X<Q1E>MTX:6*N["93\!2#33A>DI
P_RY'^S<LFHVYN_\3]_@4U$;2EBRB%J-.)G]#[#'R-]9&5E^U>836-<FU>%4U=2!^
PUH73(HKWCEDW(ENH+[?''2(L'>;U1NZD1;0D"[F4[#-)FM>NJ>92"9!R@^XHP?!)
P4*&E[8:L@VS^.URH/PQ1:J,4C%JF]Q;^"-G2@U!QO43>JCAAN3>E+&T5BWQ%@3!5
PXYB._4H[AN)I>M_C&>M;+F]K[;!*WX<YX:N E-*Q6G@^G9K;("2,+:T3V"#>VP2J
P,]2(R-&?^$;;-7B[<E\1,]:\3#G<?C_/13;[KWGP\A(K$ZD\V6I(_C-$'V3BW-MD
PD<10PW S?SYK*R>I7R-W,R\J-:Q&^#SC^(<8**K=511(I+D"8,ZN\:0<5 0Y--M+
PQCW=$+CR83>N:)E^P72.5!21G.W7)55_NC:Z+PMJ% NS0AA\/>T9J+9UW!!28&KS
P5M1=OA7&3&<0_RO:MIK<1[ ?C9#'B"P8GS][#-[3U)T/S!]%6(7: :COC>"N2!X6
PZ6@$=R/!Q><L=RAX,DVR>@V?\C8?89 <C[P8O+=)>Y$6@'4V*WU&IG)R3 8"P6K%
P\2ZH+_S.)&J=R (\)Q!$/ [8&\YO@_^KM:YR]2F8)80$4L;J=-EF\MV,*$[::+Q;
P2?ZSCG"ASNU_?/SD@<&([1%B)J'9!KE>=Z#> JLC!_F%<I,A8\%7.4P%F1LS-5YQ
P*5Q+B UBG^(MZ_<&/,H9N,3 Y3KC@H[<WZK2"KM&64UYA 0P1!X>LS_H9&:-?M,U
P OW[8&7F=5D!LD.Z<*WR$:<57W<S.'.H5NNS-(^&^5EO8SR0"F^-@BLXO:X(QFK7
PVNK'$OV=:10@<6NJJ2;7S^0.TC5W ?)2,;'.\!%N$4+GO/6Q'K.D'K1(XJF76T->
P-_]*CC7*SIS+U9.+##F?$SOKO5V-,5_QM5U1<2J"%!U%Z&S.Q'[3UC+7;D0ISK-\
P%/X1ZO8C]P\24^R\K,GB9KE."MR5''=!G8R2#G&"I=J[F_M.S&Z'QD!X0E)=EDSH
P/>@Q!/._+^/)L6\O2U$1#_FK\Y"Z77O>5*V][<5FL6%E<A,N*K?,BJ8] GUIJUC;
P" 8O$$6_HB4U<QS*;2SN65N50/($R9^M!*L7_PM-%&;^_457HX9A)OM.]\K\A^@T
P9\\/5F\3C'/\Z%7U;@N_0ZZRGDL- 35VY9I4 .&'/"M2D6/<E90!"^_W"L-WY_32
P@6 XB<\[3TPMFJJ4>\U&,7<]K0VF3\PDL&>LJ2_AS6P-ZXB:"?2<6.X@[<PZ(G%J
P1]5Z%#+7=,; ?J=?*LG82@1R-UWTYT!GU2ZZ+!KK$#5O,S]',;07_ZR/A7C$J))M
PHO\8(D\MT*J3]B.VW#V/7W4J?A-;7=].MGZ4(+QJ9/#+?ZYI(E;'$#F&*@\IDNM9
PXKJ=&+J";G.IE]\3CJ[A9P'0^K&?9,F0VJT8Z)55E5&:/9B7:]YJ T$(!DSK_/GK
PF]69S#-)T_T053:C,!9Y!/"0H/=>XV^.MEO6ND//1DQV=!*0MS%1$/:M(B8"&PF_
PC,5Q5>[E*76J$)?ZZ/#$2\>EDHHE)"X_\Q%R<J7<30C+1;\XIS.IY[KI:FCI.1(J
P*[BCY79+]";O$2?[ (T0!A39M433:&>=40_E7PQXCN##BTK1+\3?)HHIIIX+Y,N&
P\FB? U4>HTJ!-XMJ!QZ+E [$NF%:'/H6^45K)/;%MG__]L?%8_6F3[;J(1,5PL>P
P$AZH+SZAM;C8_"<K")7E&E_89P=1:QMN#A1@P6K*4-YUGG56AK(;:T7^=D,[&)R<
P%@'6E'8L=,VFBXD%V.<>(%=7ISW0@<$&E^]8=X=VD/G/8XU*C=H1&5"<!5I0;1=0
P83<.X4C;C$UJ306\73@9IYT+-_Y'H$X;%3XU3C I'(#\P*PO;@O(I*AV/R&)B?PH
P:939T438Z!EK\BMKH[,Q?3:-M:08P?QW7."V?-E$_-7IHB-I#4%OX_N7S[J&:CK0
P4Z,XCI@N$MP&LQ_"C0IUQPV=\\' 7^6$3#& 7?)LSN)A"B,TE6IO<*:<BU/60/P0
P]O> FB0?S  ZAYW:@MA(^722[K#4Z*K>8 VTX'_O;\/#QX/4PQ5[!I9H FD\7Q[6
PS-'<F:EH!0"S. #KTF%A8,R2713S[B?!=WF2PRP2%!-7R>TXTG/@;;CTR.6W-B;(
PA$,@T'[YSU)X3LYR820ES!C*;>:QLK8..Q]S%EN1R2+P!Y>/YZ.[88<C_@M&J@?J
PV4LL _GQ[B_A0Y1\A/*P:$&I"<H-5*.%KX^'O!-:%L3G\K95(&K,5*YVL?H#?B=Y
PR4E7=1["%+V?><6!GI_O'3I[9$OBH+)^6N@=%^?M(K7*8V4$0_Z<%2.9]<%23&RB
PB5>'+LWUFEBQ^0GYJ^E5O$K3?_%U_]&P37BCRGX8.HG]HA*PT+G9D6J#ZKH6QP:U
P<X47"P/T%>U&"#]9W@&EIJF/2Y!TO41H:T!8H+-^]!XIIJ !VM &]V S!+O$IIA!
P^WCRZ3AQ?''^,S;/P&4P$-$82L=0> :Z.%'@1W HB,S(FW[J/=2S@/.<E;M@;DK[
P7B<AR_F<<#'S9_V*HY\.2\Y6/5!15;BE1%.DT"AV]/N(9D =YR9ZU,L%?!D.5^<R
PRN9*<M40&G?X"X'K2CC,.,Y;JK]%J9:[D$JJ,)4C,#KS0"\/T-PTLC]F:U6R_3'B
P;\_W>CER_7>6R,QSYKVYN4W_R8LTNI[=2:FIY*?ICT&A*T23#,,'MQM3?*V5E$>4
PGB";".KH:Z? !&PZ!@TB;BX?3M*D?#'XA&G2314C\;.9Q/CW]8%>,-YQX^KV^$9S
PE:@7OT9&'H*G2PDS+9M9,OV;.3M-JMR<7HLA= [V_?Y:I?<SMK&[GM4.Q.CW"'<+
PNN+6S0"4)M?87"KZ*[$\I;20HIWV.^)[=<E6*PLEX\#?\HRA//(EDJ))8*T.!$6@
PU&B6!TPE!.PD7(?"A'8U$116BDT_Y-"$-%L]Z6O'JB,>@E1)$BC4<KM>Z5W<!RG>
PL9-\QC4&;S4,V:5/,5K8R9;?K[/QOMT'WW2[(\+0IUCM(X4>/I+ZZ<$ZIX+LSSKK
P5JD7C=4 ^ )A3M2&1FHH#3T 0#-K/J!*47P<TD&.J;3.X,E',[^CV<YGJ^9Q.^F]
P*=/-3_99_-:^F;<OD;7Z^ZC5 J<>)EM%!&@'2!&C7$'%>C4)FS23DN(C31S[$&C$
PJTD=$2B9#/!"!/&!8[!.Q33=N,V@0"G[0$^O#=^49!(8NO=I*F0='<FWG+CK\SRG
P<GARV,O*U6A</3#VZF"1D$B.P-SB-CNY@-9 6M:>#Q#Z5]%LZJ_YY?DXU\[FP_UF
PP4FQE?YF9DV%HXG-<O]S$T?MHX(M?^?SWQH5QG/=!0[%.(WJ-R8J[%5\)Z!^WW>J
P1$<QYIN1_* .^>!E,">(N']579R=DT2+!%; 0S KS9JBLW8%]^]\V:61LOV>,8R1
P("'[=ZR8=&"+_I[-V&#=7H6$N>9"$RV>N$DHF'"X>K F(PC4U)$4D79AZG+FQ"Y2
P3AO]H3J$?XMN_,3)>;H7UO ^.N0I+I#K4M1.'$0:%3G^,$U?WS7Z*WX03"B7UJYS
P,=^T@^N,R4LHV8GVA>C;FM[;4@HR$7ONSVEPZB!N*1JZX&RFBM13PFXQ&*TP'7%_
POI=)5U\->.JMT6E(PK"V-BKPM@JR.&>"(G)NUR;]3C:3P%%'_U5HON\&]%;4H/B>
P7'WF'V*=N,6)VBIZ/OH/1-(=!!XQ T@B?#UY\)XE((D5,O@J3:A@8V]=*0W2L$^K
P. <PK<.V .P,JRX#YRP43&\*M"@'$_)>=LM"]6Q1>OBW&IRT'"2MBQ#\[=13=[IT
P?#-=.,&9W)X) 7>:3H*PETZ& <MACA7WX8ES*%#++CGSLSNAZ$>%X5"T^!1F4@!X
PC50YMV29DV6Q-%.H[/)V"A<85H,'N"ES3:W<&&2KAB4\[EPPNYST;S',"P%\*35D
PT<!GF!;8%!*,Z#1F3"4+'#!/&) /4]1LM-](:C3,O'?\8%O+1^/WJPG&:L[<>5C,
PIW #,5K"8DO.GB?:)"XH"RC$FV%:>D%]0A4H-.OY-*,;XM+'9$ CM]B/; JW6S:.
PQKQ0R*M<@2XQ<;C^+HPTEG:<K4#>7&6,(5P[?'GO3LE! <,1=S66F7=NC]_"DCZ=
PTGB^S-17^+:M$C/I-\R9-%.<(PSXIL-X-0<>!WPBQ E5:$?TCS+1A95BXN^1VZTG
PGVSV!<W!#N:U[(/^82-X?XZ^G^ ,2CX=1A.'*F08UB7+V$=E8KIYO2>^^GW8YH2\
PUM8$I]TVNCGE2U9_1O&UDYC1>KU;3.U4*%:&M1XRN4\[2+,[(BM4Z[CUVHQ77F))
PWFI\</@G&S2:A\<Q5/BI_)QWJ9.#]E==91_!)(T>B)SKTK.QPN9BCW,/&"3%/L;#
P=PI3K>1H?<CQLM)^X0_=TJ?U7T* "\!&GJ3)J@4_^6_*C6C4 ,EF/*PVQ?1<.!8^
P!8AL2.*Q/])0HS#J!X.F+5%7U3X>'F(DX(^#Q!\9QT8L*H 6C>WBXBC*-&#LGL7>
P\WO45*2T+/5N1'63LMKY(-Y!:Y13L?YTR,&]Y0) NG@+Z&7.S)ADKS+=<VT()N:?
P&WS"5E>BS7I11TW7Q9P+K0YP1SLV',E#U;JWS(6;0]2WDF$.2\? %";F1#*)\@8Y
P%&/&_4K_O[$;[P!;N\RP!3UD0G,Z_""O<U/YB6_966JDW8)*K*QF;J.<J\MG@"FX
PGE[WCR3J"&:WD>W[<KI]Y,\.0&\6-PT:L)_"GT^]-SL2BQ1*JBU\F W'=G[9XW9Q
PTW)Y1BK3;0(AQBQR.=<7QC,OA'#*SGDCSML'J/9M$ "\17^'PZ4V#TFQ/>Q4G^0F
P'V!<,XR#B/5N]\#PVSC!UCM6H2+(Q:3:70%_J1\UC*7?->,6<X*("!8UPB7P2A%F
P#KBG![2(B%V)>+R;+$:=6NP=O$>BE+I;(Y4 03=4>S@CB)6+>@\%M-ACY_*W)V50
PN*B26SH$'\>QPO7:N$Y7N727#ZL1<_R*Z\[U_UG ]FDI-)6QE+)295H@K0&N;31,
PI.K@R6CPP5J9X!U9'<*:+[YB;6=S4'9#WH=V9J3B4;7U:VZ3J#/>Q1$Q\($-B@VK
P3-)JQLIRA=J!$-I-';!V:V?*\1 :I#N])3F5O[BM]&C+DA!_^4D>8U(,5&+&;44+
P#?T*% )#%90DW0OD<$H\=+&^L?B7, 22QP5*I#^&"L8VA=3 G]""BHORDV=4.4(G
PMU-85V-_LQ6)0%!=WL$O'WQI5W0L1#<L\%W7A,=[X2.<!HU3)X.W!\[L0W?[-WE0
PU=H>#V'PG/$*&'2:TR@CROD)Z8:#F]M:_S:;EO'[C1O@E1KZ B!OCARD;XYC]R!^
P-Y49-:LA)SZ<WJ\K]. )B:.BD1H\B6:)*)T)/4,BP>NVG:@ WZUNWS\FLK11MYRX
P@@(Z,<V"CV;V#,19*,C25(T!6&Y&=9@KZZ)DV/B.:Q8 _H^*0L$7"XHO5#'#6/7F
P@WNY'YC"%A?G5A5$-NJ*7"=49W^-,F.6VV>83BW+98XMD+!.7.1$EFMO?]H16/CU
P 9G5_G250&Y$XO"" L 7%9&+R(MN!9H=",$4V'Z4I,@$>S&"=J *R"@8\2RN@+UU
P3"L"&EM_V0J%IQL<7^)+!%8.%O?%7,&^ 5X9 I(>_R2DUM*BP="!3:>W=@UG=!JQ
PY$+F&:X&)\X3E#^KS2S?J&@LH ".86"\/+ L 6Z*@QQV0; WEAW:TW_94.9%!)B/
PWNIE^EY%.))A$K5*BR'D;6!@H,K#ZNDTENA-%HN\.'<C+"(!SC8U9YP18V;FQ\R_
P9 9SCSMJ]:VOU$^M1U_B<VNTWC .VP4R!'6GPW>4$VL,FB5\0RV.QUDLLE>/[UGW
P6736=$_?E!BYR1O/Q/N6+;&TZ=K72BW2Q<]PNM8\UN\)^500PG8?3[-7L0"PPV_>
PN+H0-S_L$*5)11]8S>#.3NW=Z"((3 &.MPLE_7I#EJJE,NY0W=^$'I<8K3B!E<1W
P/BAQ/M.,JRRL.<"UATR,PF_F,@/9E]0Y0)M+;_X>6)#ONO# 9KBZ:AE2!0N8,<O[
P)"/V9KDB #'?NC#O<.9II!NO/\$N=/?$$2;;:FJ#5 A["9-607Q/<KSPUX*@:!:$
PAZJ:,;5Y^B^M_U#4S"4Y6(H #%5FXV^"R&MQGA4ZR/8IT.[,CQ,Q&6D;D+[;[5UL
PE-&GSJ()D\+ ^X\>,EBX/]9(F,Y,&8)*YMW.'"Z_VYBG_AG"MXE3EA-2$<9PFD.J
PW^%EN526 6%[3!IU33GMP0J2X"]$>5<%B?&&D\:XA0?V<)G+[>>"ZRB^.I&X'OH"
P$6*_='0PZ/_EFT 8&GW[0KS'9*!DV^D/]X9!$3Q464+A$SQ$B*LMNYT7K3=6]W #
P(NFAD\+>AUN>?R'%ZSO ,S)N!4=& 3Q_HC0ZGS: QEO@S?9.AOW!9-TD\1U\SQ'7
P]#4B2.U_*]3C AFFOQ@I O>:K)M$\6INOK75,@5'1'-]L@8^NK\V2<S[;5'\S:%L
P+\O@RIWIKH*QMX+L/<JKSG-3>#2?LGJ8-[)L>^14U6-&Z !MQ(:A8XP$ER$] !ZS
PH8<8ZQ4%>5[_KART''(MCO2CKBO6978& ;#RBU[&G#NGANV/$3<6A::,9[(&9&O_
PR[I[$U7_ZT2ER!LWB!'BNXXHK/2XHNQS#KY$A0NE74M.I'^7 ']TVF3#'?*K:N+A
P"ZI,[WWU>0H5&),:>?PJ5G_.3:689FC>H&F"QZ>.A'U0V-#XF;@<Q4+$S+G;M)"Y
PEN>A_.&/T94.D(P.7;;/ ;)UVBJ@V8CW=9Z)+#"])Y_[K_*S][/UO*,G NBZ@V4*
P%-$&%-V?MTS4'M+"%SW.G"\1 G7>^UC7E04ZVJ9@ %*X$FR5"'RR55-JN:.=;V2%
P#4<\DI@WPR?A/M,.< 6=!ESO4WZ0,@D)P6O)/HE?KW>--1F]E%A Y'B_RVYT$O54
P=PY15B])#6UV^I5==7>4&G4@'T>OK!]BU?3M7CN2.8)[_H7F(=_S1Y=6R.1=,AR;
PQZ7WSIP)R / Q@-@.B\"+XW SYTW>NI^6',+:IE1FAR6[*MZ2X[(?_DJ<VD;_6!]
PC9MUCE[!W6)[G +3$HU9L5:F.WC=+P*?PNH22S0$LG'0^1''BHH<,'(%PL'U4BQ7
PR6\8!V\?R\S]N#/KKG$"%P(RXZRR?K0^]#I!$EN#5[-K$'A\W8<Q(.ZD;YVWV._8
PM.W?W)U[!C8O';%1!BH:%H(82]BD8@FMRZ'SQ#OJ;G[*69W1<[>TU^Q7!NW<_A_&
P2')DB1RE,4-9)Z+'X/Y*)20=>#H1JRV5\H])U^2"8P,M]-9A<K;GM#QK&I$:/ME^
PKRKNN^6]1FK'/0.AZJQ84!P'2"D65!9,60(-XZ"?+43CE*\7EH6@2?AQ.9?$1J<]
PXYRCP(I%N_V9Z+F4+FEM@;*)/Q<X"8=Z!HJ0Y--G\:^T4!<>Q*4UU H_U[_T#[ >
P44)71PW44H8?=YSNP1B6 [U_LL-!2@I=HG1OIMBG(5\VV0#"FT%C,#^7G8P=W_^I
PZ)2J=Q$Q7$BK=[66^XCEJ:.,[W?3%N 51?4-ZU*)<A%Q06WMO.OM*@_ VJL5D93#
P?S\H3/MB$Y+6*%M\;TK79?]"Q<ZE-S2P!#43$>C8DJ#F!HHX-Q^-34QA@>$O?SUN
PDM .8]ZYO^W)/[H1CYSR[">3MR5CU'\7"EU6T#7";V]F:S\QJ?SGY_QT%[9T^,>V
PXMCCG]9'64?"QUA0I3? ;O6%<_3HY*;B6#5HU2!1S>*W/Z:(7DZ=.RQ ]>HR]D"N
PBL"._23UXI]P^^:W-,3BUYXKBI^:LJU<.>/BZ7AA*[IO!3HO[I'FUU3M(   3$OO
PP%36AO2?1#T.I#?,%EK*9<OWD27Q^@+%9&%(:-*U#LB#G%58D%$!/!LL7<-W9U.F
P#UH-WC3GKBSJ8?FG^7?SJM/JG?RBAVZHV!Q2>0G6 X *'$5:.R\!0JHF4JA'PSEW
P#0A8QE("#^-"R[O\X%UP3=JGF]P];M0:V0 Z3@\^(RN_OS-M =.J7W=D0@Y)!2D_
P5J_OW%PP[$>B&]98^_[@43O -*CEC6L_+T3$+;DPC<W-2,E&\N##H'QP9%PTRF</
PN?-3/DKG*%?^+EV+J!WY3V%NT@'EX 87:7#&P+RTGVS_ZJ!YH@WD=PQ6&#8=L= K
PGA(SOO?;7 "L+4(>,,Z]N='-W<L'X1KK3<\]QA+0DQ3S6:130#+J2 XXQOWK:-#M
P&8-I]\QJ.CL\IAFB0BE7U?D*RCRT")@JK?#MHM^*"UK%ULZ_M]$!IB"\)K7-M&TX
P"23O.\?#]DL'M,=.-/B.[J<DNVT)'<.S*G2>=Y#M='L1L[V4Y1BM6;H0RV2/>.$W
PI&,8ET,65]0H:,,K"K.CL#KP0VJ]TN2OJG(U=LEE:2C\RVA)DL49>.';^^=O6IOU
P^;_8!<NZ:ZCSU[+N*;1G'@^M>DMR>43=2GV.2TA)YVNN^<#M><&+%/.5SOW,_ZCN
PL_S7FB&?EX[5ZH7.:N4U%I.9BE?LS*EN0LKRET:79A+5<A_F]9V@A)I5ZE5BZC9%
P@J4B?S%).,?#XF,-+/[ R)^DLP7IP'K"TC;+=)S:+"YJ8;5R,/*ZC3=&BW:(H,6Q
P/(P4G(7QB@!3?D^[2V3Q5=HY_S]C*C_5Y^I[YX!<3%1B*)?/XEGPF\_.GJ>U/A3-
PF]K@AUVI:>3ET:&1?%7Q9IR=QF>&7FJ<'$MATS\@?R)<3 GT"%GX6QO/ZDBI"?] 
P*?@1DKC@@UK$'W:78.ND;N'D%Y(>I/\.L!2%[=+[K5I/%>=/<HWY XC307I WB%!
P)V!X2(*#E4_R)IJE:R=XKJO>X'-M_-M5)Q!C(ZXISPXQ\$^W^*E"[ZO1SCHH]DRD
PP OKMP5'ZK;T;KN-GJ-UM9=TMT#\"@SE$'7ON,FSWB*AIS@2*T>7I:DV>=,V )HN
PI0>!-E_*=ILJ7<K.1[D*\"JDA!K *F(R>OX(#^)T4C-/%SL);=Z5J,Q!=3"U&7G5
P(F[E5XH]NE5,U@Z)3=&/FP #0=0I-(CH;7Z1;HO>;@(T/Y4 WUX;=#?:/W"ZO3%R
P=!D(QVIUO@8]@IP-?(A/=E4URYH/]C 2I28>B>I2I?%<$\N)M XF/Q7/W+PZ)KQ&
PT@SO6N\ 8"?O4Q7#HUD'47 R7P^Y/*K]OD.#PP'ZWE&W!3W)SA%=6W#3<2(E[3[W
P+)SBMN5WV'J55OZ,,'Z)3U==.I8GWI4&+]4)9":E2KV$T-YK WEOU*9J8;L81W>E
P%5()QLU@ZS>R"  D-$!@I1:+Q?7^[01%:(&D8RSELSFBJ[#)*IC (_W)7IG>)0,>
P/%CC!G=:8$[G7S7/@(H'KWN4TP&0Y;UX0]YK!#=$5^14CS"<;RW2Z,Z\';KH#4;J
PJW^H*<F.@PWZD\&7OA\>.UVF(X:%00#/H.D'5)^(H%*([THYF7>7?V%)D 4$/"R4
P^L<$2#P).<>.CKG!8*@*^=/OGW"&9"8#,<&IDOK:K1T[(N,(;7(+NY&[G2OCRI!]
P:]JQ(T!/RN<4SC7C6UPN+M*U8AZ,!OYD)VPOI^B*/EM/*(N\SJX9:0:T;0^=."N 
P\[!7W%,]O+7V/S+A36<=]:(^'Z1415]YW$QJT=^4A)IJ<PI0&V*/BCY*2T^BB+$T
PLFSOZSU?V+YDJ.8--;R#RX"4$VL*9?0,S5H=L'>#Y[?9B^:NZ3JIKXC=V,HD^\23
P\*@H:8K]Y.M!2VV/WS$;A)LZ3<(%3(S.Q<MNYRC?+BH<)([Q#W/@J(V\K8?-/..J
P!/O*3G^F Y9H2M@W,1]JBAF\_4T390W-NSEK3_RIF4@S,Q0$$&2/HN>3I)];%N(-
PHKWD4D'1;=%> Y5XP&_B,9#A<[/\%2L4!G8:P=,-44^.VS?E36#N-O!GH7D1^O7>
P=9(A&]U#?QZZN:K:6K6R0@+85/5B<,K;164XMS)AS+:NU?GRW?25(G;.Z4ROVYUO
PSF^74L?1';S7]@K7(7;*,Q1N)E&C'!WYNSY'D:=9X$O$CQ>I@)$*2?-X(>>^$19,
P@I6EY$.1>V E)5WXYPVZ">7#TZ&3@8'PH!M.U?U+*5JE=?_DXFR]8"P((!J"#]=2
P;!R]H[LKI6H4 'X;1=PL<]![;@>H],D:2JM7;>:/HL80_CCT380!T,W(*KDJYR#*
PGI4[2BM"U[S<*-30-@!A8#(!);L"XP61'F\@D6;!+&N6A@1@L]\ TW2/EVP(AUV,
PD?^6#E6-@;*4B67GML^8,R #<%(\!QS%;4W,3)4OWU81Z5?)]QA=79;A+6X6.$.)
P;9I%B3_T\O^#?/+%?-$/A;M0\$[8).0U)?/X-H#,+D.[J/2;0_+UE07Q2OY>)=I>
PA.O_X_()83$(2NYT]D%R:8X.ZQ52_FD$X>)3COK55H*::YFS%BY'UEBHU(?9KAU'
P9E8,ON.C!X&EB9J-*N@4\VQZE!I]GH"\GZ\/=&\QASEXL.Q)E"%R1<%M(]S/N^BG
PI!*WHP]9FQGV$IZZWOJ;GK/[Z3#INZ'"  ,\%JU^3/0X@4%;3RG44'^=IR5ITVE6
P PU9J3'=+M7%OS+5$CJAT,EU7E6XQGG[@T5"_K,"ZX1KXJ6]>CQY8S7<%[010'M;
PCBJA]C@$R.6'L38 CX@2Q]S!H0-3L'O7(-56SC+]AH[.+I.0Y_=]PJH>,9EZS 98
PQ98*FAZH,L:LE/K6P9''=ZU(327R0QN/0C27567]VX"X'^ !Z]@8O_(-1&<-(EI4
PS>8=O8M/W?^ <8)3?0@+.+M-1PPP)Z1@!XLJ!)Q%Y5^D93&?U65/=LE%F.8N=0G/
P";,!4_:4;'E(0C>-@74Z<BJJL2$.%-[5.UB'IC6E"!D$-3Q?K]*%S$C3,^U+;M_<
P#2A!0=PC^F@TL1!KV^B:9@/B+(B*<$SS>8-096AOJZ/=@U2S;?"28XF&L&89MO3D
P5(3_JU5JKS[@2+A[T-;VD'C;B503-1)@=D-SH ZN&CEQ:ADBYTX.0'=E8*[38!6R
PGQ2/\<PRD7;Q="XNYJCJIU@ '2PM>FTBW?N3T;" #>F->6:X\R<ZUACB7?GQOHYN
PC>O]!I6I T6N?LRRGVSHQ.6_08UAS*G??1R,@%F.I4_R48D#*6@P4_T\WA$RFE",
PB*;NFMC;I<EV."+-$A[[$D%1#%"/ ;OF8^7@$M5OA']AP*D-\*+&_A.T3E&B;?EX
P+(66P;&E\D!AD!*21?^I1+[-27<3'W0RXNJ=Q:?*;]<RHL ,@E;KU,LUG+;I-ZGB
P<@0DB+H9/P/M:31*NP[;S5>]%TKMWQ4"+/,&H!V6GMBC.J12=#E]5/\YWDB'_V'"
P@+4U#A].)P=_<AL9-EE[PTUYJ9<8TI$B/":<V*YSA6Z;FX7L\A*2ZJAIY(!B2>=-
PN(IBTJ7;!UOD6 :0AKW_FY[#HGC*JIX%7XR1%+Z8.>:2D5I1T>T.8.W#,NV"1YHE
P^D$(&XB"JG].V%^KW/>W5.4%+)9IT?K3<<_Q7^G382CS$AZ:7&"_ C9/7A>0C<\T
P,&/-0Z6"K33\O0[J.52$W"U,I(A2L$^0A7;OWU5>7S([I9:ZV38:G.JRUY1<R*JK
P6-EOT"&Z1G#%90.[7,KC6.131C87R9889N YSHT5ZF@R/6#8^L82..H+)&X&O"S0
PA>.3M49RFF*AM Q_*B0&MV^26-?J[^4AA?^,R;S>=P]/X\)G>8)Y[_D_SO<]0D!1
P3GRA?7#,E4J]A@!KL$QAN672=%_VR(X1S8+>\_56FRW>41[V(A/8=*I)*7V0L&P]
P)_$$WB,@T(QUY:S ;;4Y99+SRK[2FA^77.8F;17Z5Z;C9K3(/1I$4R(:?O!5@KQ=
PE:MM,M %$S/[+H8YM+E"0?GL5K?T'P\30N0@M'PJIJ**:"4=P<$:6F8.D>$H'D8(
P7<WY!"T7[E6,BXM\3&)[O^K@/V:OQX%6"XL!/M&IO2A&O1:TY]="CJC>S-7@.C1;
PXT<9@7!=<S>]'?Q9;I.J,*JZ7_X HRP0B%61DPVRI5UM5][7>'2M"F8SF8;GFT]T
PWT--$?L.R#I[%7VU/# 1W-V<CWFI<R7_O6]R36CD(Z>$ (G?5=@OESO''G.D+?C$
P1A&>Y<.BF_@JA^>_#JECS10&BP4^FGAS2K#]LH37KL]PBW^J[78LAU5_&D-7:N"%
P@-:]B0;-M_PT;.O+^DFC0SN#7(IHL]++0_I[N92%VN9G#LD5Y2S3'/?H\[2+( ,8
P$ "5--WKE? G"AR&_I'A1^4YUK"8 \ZD77"JFH_)_Q?6I-K/!7L(6.9U.9 QWN"K
PDIR#4<%M1Z!B4E52-3%/Z1V+I5U38)+%KEB-Z>U.6@J:-]MM]W.Q V#F-<_6*@=H
PF]ZS#M)8G_<9RG^UY@O&A//)!9%$2\VWSOUGQS5ZS1:XN:Q^D#CZDJ':V+N>\#57
P&K/ :+:I6H AT=8>UP)#O"*6>,K\3"1D!143/"KTZI]IK?#?=F?4'M=_ A%0WAA2
PR0.57(=4SIQC*;'>XE7W/C)LO5=]@]QH!C6+B8IMY#>C_ =O+#NZ90#)E?[%:)[_
PM(<6/9<X#^0G?*Q0)MW$-9=K=7VF=!T NM/GMV"P3]OMJ,A0V%,=T,8TW,\*Q)\C
P1WL$8^CKA7:5,I[@](YO^1]6!O/0%*_<')YM(83"<_,\G:_E((SG=1PV#Z*%E$5K
P*E2;]-OQB7D0'B4MYR.KMY(H(VFT3=NQ=L)SU;<!I<;X:*%]#)"ZQ?8@R3!I*/0S
PXH%^'##E+PS1IRIW5'&BW4Z886Q%N&Z?9(A(+$6G2!:KHIW[N?R)>.L^L%[(A0K<
P"O</\E<.28>/!S0YKFD8\2@;I<C],[TQ?1T=)W,RT-!/?U+_%S= A&N!<+5C;ES/
PEA*K/ZWVJRP3C/BR%4D)W5.5%N"!DB2#YD-EG!T#@@;  H?^K_GM#8-.:Z]XLS8Q
P&K%9%!S 7&M5.T>O#(#DS:16C"C.<_1I^CQ*0[4%0<XK!Z0??RJX9K)5I"M=@?QJ
PY6\JP2YIPG[%=#2Y:2])^%;%*].?IY)*VHRI218??HE609VW;>OC!M]/\,S,0[!1
P\8FB=O#P]#Y#J/_5WKY4*AHPQ5U6:>)#38\_D;(3]IWY:EZU,D38+#MQEJT3$CKI
P.;/'8:CV+X!)Y/GOXQJ/)Y0Y\1K^D=FB:JCGI48)7[\= T?8MPT!?)29CEV4-.#%
PVN.'_3$L00?]=&ZVO;X1D>#M5*.$H:F^NDDNM[I*U)=T*"JB>IL1TR*::053F =^
P\Z/O-"\5SVGW).]KLBL(4A[JW8Q0D+?@:CH%)@?%GF2'DW'9F;3H.U(#I00=.;H\
P"-'[77L#E&147D C?:;H-);*@,JQIWARSH3 .G*%:$ZCT)WJ.K75=&IYR1[P>8F.
P)[QCFE[Z1O]6IV%/X%J38O13C!H2C.R'S<M<\K&-H\[0Z9+8%+0T\>_"8]**$ZS0
P&#96ESK#,B%@FJ+>#CY$Q$KVF0J<Q_YM/)$.83"#KA)TA1[XQ%D^ZN:C2288?UTC
P_/)]B^*3,E:-JJJ9NV^/ZBC!H_0-O&))=#3\9@-_$7S':_K*K?"$[PM%/KY"^Z@^
P2#3MWL53D 8MPS[PDV7<-NM*TR!*6['*O1J3<5N\(?^;,T5MC:+L&F(X@I@B6#GY
P>LJ^P(U)K:\;%3!V*HP&&#1EP@&@R8/!U0\$5N"4!VQ->I.-3/^9^WGZ&7'Q\($H
PFX.?(N4=IH=C2+%(@^]8H A?_)U]UE+RVO:TL<M6F<#U7C$6$O+]TD)-8P*=XL=J
P>45!"^SGK?+\@JF!?L<*RA,CJ$N:_H-D7^4P/?A3+)#QZ(&,:[5'2!!]NGJ(E$3L
PNCHOZWJ6YY\_1U*9XL<.-SA/+IGSN]]1MJHUM\3F;N-8:$1][VYLG6!'='WA*,MH
P="81SG](%X*J&BV"C]Q6&LH>5+:IXWNCPJK3V]W@RM15?6^/BA)]HP@KT%Y?)VXX
P?YN?BI%)@+ZJO\A##H+07@W[E)^#45SX3T).&%3*X"SX1$54OYV<FQVA@S]A4CR8
P]PRBK)&68L9[U*W[%B-@SJ=MJ%GO)_% \PS,DIZN(G]M#U/-JD\'./5&.4K@8S=U
PSUK6E?)KDBTF!7JQFH@[F>61?O9!1?DZ"N23";*.>84/G;2;%("X=GZW\B"7L'?-
PD()$[,$9+&8</BJ41.A71G _*F!LDJ6'^+G(KV0M]<<LFJKSC\B[:[2I@CPS\>.*
P\/TZF*OP$43'MT2?YF.V&ST0S;LR!J"KK^'\&$/%>RQ^-[S24"2VX19IM%=^.H%&
P0WW/$<WI/,X*ILWZ7VJ(2%*R0 *W<];/3?7[G"S*A%-*R*3U1KK/^N(-0^)^G\;=
PW<AINZ&5^NUA#Z;@-\2S[T:,939P=OA/[$QA\0;I60"NI@?,@HT2*U ._I7&88.6
PMP66DTS&K>6=BVV&%B%7:$T7 9Y=*W!2D+"Z40F29XOEG#65:TIE@0E+NQJ,+R=C
PV >\/DN9[8!5;:DD,FA5F)!-5E!BD_+!ON#1,5M9* 8/,3L$#.2(;(?Y),BFH;NH
PDWR.Y')(*]1;4'8HW-\)?GCGK=K!B19^>;Q)'PXXD59844 0K>/UC+Q*3R:>.TS:
P'EW(F-8#*U8>(8'P^@^6=AV1\Q+%&]3!$+-LOUM68E("9$)K-B!\R?G-.?7/P1'^
P@$NPM3)9P9YH=UQ(,*2J0HS!CV)B752./(CV=(?CXO4_9'=;2^W$ES'Y>'L/:L[^
PR7')+X\3W'A:]IU#THF_R  AUC>%.O>G02>)?;6G&K'(;IW(+AFP6^R,"LTI>=^&
P)':FZ>I/_$]1WBRB8Q8GP#V+^7ZS>.['1[8].W7':*A@H_P-L@S5/@KX(XWD4L.O
P#-3*F([Z49\4C!6<XS7K-1*XFX3/_JX<HGL2]<?ASO+PJ-#3!%599&-$=#N'C-+[
P2V ]RPJ\FK=^I1D(C^/R%LU!_<C:HX2'BN"BX/-@5>WP\K/UYG74[+L))2]4,3)1
P!F$0>W;1OT;-+(;O<HN# WJ$FV'Z5T]&="".T_W'*6F;=!USH2S_)@PZXQ7!M.&L
PGY@]GJI6O+"BB$;;[Z.(P@!CY[QZPV&0,.F=VX-53^M-OC8<OH:&=O%,87Y\1]G:
P27.Z/PX:A(J>&8:L3F!FY+FKQ,7(#)9_>XFV!5+*H/AF)&8/\CQ[B(+2K(C;47]D
PX<&'&MC2(O%\2L!3&5Z_)K%6-.O#6SOF.MN)3<9OI0O7&HQX =D3VIVJBV_;Z=1V
P^3G/LC>6 &#EC%X>.;DPHT&@C*0CHK>5MJ7%YPIG2 P^\M=\T0_[Q3Q>EHD-M;%G
P%MO!M>@<;[0WJDM=PW4/"VMOF/YRMBF@I7(O5;CH?KL 5<PDAM$$@HQP P 5?D9M
P*]NXLU%G24DL5)@5E<[BZ2E)-0;#L<QM?GU$VTQV:WB_&,)XNUWH"YX;+Q3F=[?4
P+:;.?',*17FEOK8:"#.0O\@8?J-^A;8<[,!,9,'.(=UDO&26+]CZ@0)VB,LV'I@L
PE(A.5W/X3ZTP]$?<Y]KYWP50(X<SUBG'PSL9$'@#C^P,ZZA!7*?%6UM//30U9=R(
P4,\TB)L+:C7^]TIDZV>^%1O#]Y\@-N#Q?D;'ZNK$/NK>,(O'SK-S#(\+0:,'\'(5
PS@\*=\CX^2=H;SM=ONC@SS/1+(:85;#.O;\>R>*D..FJ]OK+SC26<V^X>YL(.D8O
P#WOHE2+W\EIXVZ8P' RI!VV06KPYU$"6I$(>GT,+3X!5QK<RH"X)N5'TC+O'9,WH
PM^,'-&<OJ'&)O1RO_E#8?J18^9U^/&<90;)=,>AE3-# H)B ^GR/N&7/@@D-69<_
PPFE)+#J75Z.9W&E',^\?4 OIWSL%*<JN0&H7RU *^%,@QBL!Y)\BI W3ES?]#3NV
PL7T'O4"D7MPBBJE>?C*CY$PN-/D-WY8RW$HJ[KN4B'A*C>+87[,C<>)>KL]8V$+<
P! P2N$8BTR)J3;<<]1Z@CZ63(E*D'@D*Y2JO7;ZH.X*U)FXXH,RH]&I+@1T#2/I\
PO'Y)E5'5\!*S#X/D],@KR$W9?[#@G U]#>21U-+-#MK?Y,LF)[:/#B9@B\(>_V8D
P3.Y\:*TLU_T<@]K0K+H<!7=!E7DD=2#1Z-434IG(>>/7:/92O-Y4]J]"<].4"Q27
P6GCZG.L!#<*G(I4(3H8K)I6YZI,=&U2O7T)ALA[+[,BU,7]5,-F+?+[?5@;@;_I4
PH-\',!;Y^CC#,O00[,@L^+1MO ]UL<==,CS2@2AG%19A-[7NJ7]7B\C\980&2\+@
PU@<4RRIJ?9W<W^/#E>.GU2'IUIBL_ XH\K@ 0GY:76?2Q6X65736(%9W"9WC&<S;
PN7@;B2#""%(6"=0X0U6:?D=\!U#5?9<0JTI2]Q1.\?S2-];"N9'3S*BSH_H6<A4:
P<("MRY0M_]D1FQI2$5 NGW][,Z0[+6=4F_YUH<LCH:@)$?;J3M\I>M9_&6\IG+L^
P,4M,W_U<:F8S5+*ILNCOH(D1,\^\J0^SC@MZA(P,@YH3#VRT1LCP._P>!1'@S.@_
P?Z^=:\J<C<0%'$4[E[=*B;HBT<BC7N16/=6/>)8)KJ4G;I:=HWU,XX=J9_K%W%:9
PB((HVX:98N^E=^(WYC@" ,.K$!BH)=;R^U-("J> /A3AWJ#%WD'&>85H&S%'R-4"
P!_R,W[(SGJ.OJB7EF'9ZSOWI8KI#*)N$DZ@TE(:F'F,5[WV"GB6R;1Y$;B0O\F5M
PZ+.[N%WCJ\L8LKDS_NGU>F*G:$ 4+:=F8BHYO@9#P -'423%V1Q+4S'=WFE:,74H
PN^W]>U)Q\T:KFW K<'$RX7%33(\A@68X5[2X4\P$W7@^YGJ7Q+5TP#Y0W,+6) SB
P";X5@D?-X!S9S:@]09J2UXRG#!)[M>0)<]J+78+KWPV:,+PK\Q3*=;=0.'KDL(V#
P0>+P/LUT\FQHW83:V=<9&>-A4+.K#7 [F6+Y PB:,IV6*__C89R\"L?&<1EWN+5B
PJ&T[T@4?'J.*)(HAH1A="PY,G5;C'^(+;93>PN,P*#9R<@3POC].<L8)'==M*6;E
P+\POM,37'H9^$8&\OYB^8@^?^H7 DC]8JT@LHW+")%NXF2_VJ51MNT3<I(QX)(Y>
PQ,[Y^=($[.L:+)B>"]]Y\+E-BV*^=N-.,8F:/%I#MWW<*87[C%4G@]P([OK\! *6
P%8#NUO9*>SMSKF:;IW%RY9CT_ABK[@9GK;C-]&H\1B'Q #!D0VV _ I9/$V2G$FJ
P[N*$AIB2I^-/Y8(R E8_8&7/2, Q"Y:8>-P4O1GVC_@+/CR]%TQ> \\5WQ\B_#/)
P@:;2\2=?*I4A'8Z&5'(V*H!].T)=9J*!)U^8_Y06T)MS"JNC]4BWWA\L+F<EXZ,<
PG9+9EVXG-PV+F%8O=(D8>U/SW3)^^2@%GQ!;LY/B74)<TJH 6V6K</_6S:UAI-\M
P)V\&!UCF)<_+>GF>PDZ+YY+FGQW4R8ZT:-J%G O_QVTDL\'J0-AE!1;'$2/>T%08
P@ZHJ1%3M6ZL)W%_8-D/_9R"NM0]:<1GY 9QVTOYS,D2^HI:C=\3E&@W8#3,^$%TQ
PF=J61-=',K',/%VDVM18=/\#C\&1NF%K_H;@W(Z3XEJO;.G(J+U@F_(86)'KK\GK
PYYN%4Q9))4/./ALZFJ!85L/![Z@K[RNZ1@_EX"P*SQ8(3<F-1&I ;41!6MCV%ZF]
PL+T1"H+]@*P7JZN6_6^73>A IS#=L!H\04B<E/Y.+\9ZB(8-XF><X@SVV$:K<*C,
P4(71OZ_^ 2#T#Q!K:1Z23SR>$;FJEB&<:LSGX>3"D%^]/A'ZSL89T;^ ]"8M<SC\
P=19*]9XFQU557B<+LRV,+4GDI(,?$_C1F923?X0'$B+,C/ONML7V+9:9G/>L%))Z
P\%CPI'R4L,!AJO+J9G:N-.O*Z0C>8A;>S&U<F[8EU*R;-H9/,VE%7C+5.L>I\G".
P9Z_8KNLU_GE[B&""CQ\G9,;XZ9U_T=;E4J3#H\!6\;VY)*B&SGT^:_X%5]>8RHS8
PRV(TJ!QK1#B G^ ;(X:,!W7H1UM/[ QGVZ(<U,285A.,W!J ;4F?3Q@AY&OS*=3=
P]#TFW.#\\N:5ZX@Q (;/N@(*I=_*_8$M9?]B[*,P!S&$D]%: ]X4'YH$JS]R-8Z5
PC&O;:^&H\ ,@Z@7RIYRKD%_=NY?7\?8/?<O.$CN)IDV-=)H,XW@#YLC83&-*ZXU>
P)"*Q(=R%-?<?(2OI]A(A;\[Q<B\0P[PWRC*;J2;G1OC5>0O0Y[)*7#<I_TF">Z\F
P'/?D4&XQV3N474UVUX=]H-=>N8 ]1?=-I6Y?(H=7:<6S+PKV%O_YJ";HE[U:,..C
PB5[-LPB\/I#G@J.7T5;\U)+_B(>64J+C0ZN(.J7(=F1]Y,D[&P]PHA0R)DW7Q+#1
PU;T>0^'--M,+PHV4J)^1OMR?^=R=^/Z6X"2"Y3K PRPV[)1#TG2OA)H"_@_GA?Z"
P+ZH8M6'3Y>5)4P2T0 'FZ.36;*$M(ZG']R\_L[3:^'C%2N1/$LH$PAZ7/L12Z/0F
P5.4C8-)L/ UY]CV5 @FBK4==K^-K\D'47MHAR0EG6S?%[(O)L9"X7QUX%^EL:-OE
P)?T@,D^G]7EU@U3T1VHW4FM# P@*<H$/154B@\YW-^)$6*$TCDY$,%K7;=2MB(B#
P TZ#H?>:V)4-5)-(!TL'0+K1-2G7W5G')WWI=-BU+TCYNQ>I$$6G+LX%1HIL7 ];
P%(=K&(:<8E.S&/9)[LYN5#]"QK,:IQ^!?''T"V-KIZ?]+#1L-C+15<%!=/"SLTN#
P=&ZG?0>,O%A<DK;ZD41'2TZIL"T+5_77YR)762$4!4N6"ZZAM'OB.2^<=!.[)TPQ
P5X*DH(K$YMT5TPBO%@$67S"+H#7ON+3N4BKM1SPD/3B[(R9-G$&/'K%.VGK6OJ?R
PQ5I,Q*"?V;(%; (Y%\V-Y3=G"N=,9[C2[=X*A_38+"[Y('E9:XW7'<,,R#950M%V
P'.7.!1 8-HS4A\*5_1PA*K_AK<A@6+=S^OF@8693%4--LOTS40%A,9SO^&H%P?\D
P]),]UL<$U?"R+6SRF]7_K&H&WB?=X,/63.@'-"N0JM4WIC[,-S*ZYE9X)@:D7!B!
P42!I<\^G7H5^^!HO,W"O+>*4<7&D)+A PFQ$WX.C,@R[F^WVPDMYX/CRY]I)7:< 
PD:\MOI-PPQPP+?QJK^D-7V,%V5Y@_J?\FX%K,FX6(.L+?H5^W_?=P2]T8R,QTE,@
PDX]92W7+=YQV,$:Z^O>E?M2XYB#@.?JKXR\V5/P(NB64[A1M29)&PWLI07<^M5<(
PGW$L,")E-FR*?W6!"XD+)V^JJ?O]G-HF:6Z8KW-%& -V#&-G&P[,BQ(!&*(QR'$O
P*9?1Q0N;\0$^JZ!U#:+:2QSF',&MS0&)NGR-0! "=0\,H)>\N-4W'A/]+L"/>#]K
P(L(C.7@Q[X?KOG \A+[]@(@L!IAXJ:'RM_5B!G_K?\)E;Y__S1T8O-^.N#LK.SY8
PL\J>CMO+6C"J2*ZMRW):B23J1+#.HGG5D&,JWO?M3W_F#L *($PEAC)$3<91_YU0
P</EKH'C1+^@?9]7SQ@K>)6#<"D+$EZ(TC4I<A -!0B.NN=R'Q:P<4),;V^4EWHF1
PQ>H:DH\-MZ#F T?2OO8K8Q2X1P(EPM\X3,%W%6^$O:-Z5N_HM@M4*BTJN!7/ ]T&
P73/1RSHLYG*FKOD+&R%(X:MHKGUK6L$#.8A9ZC?-GY?!X"]=O"'CWF?8YTR!S)[5
P_&VM[ZA,5NP]"8#(.Y'Z2T!^?Z>C5Y8#C? A\Q2NX9ITJ#62YY2&PM92=?U611V^
P*5$4"21EJ:3%.<>T%47Q+Q"E+<0(>\B(_W?D!*8N"=2R7"^=:-/U5;VTO5V'_1&>
PS3AVO)97:-!B/S&CSQ1.H@8PUZ.QW4""\FWLMT[\@78D]=)C'BB5UQPRS))T.VI 
PT<*4R;[2;Y?UX8\TS2^4K[+E%@:@KB#U6O(3MJZ!!YD*0!V7J>,4W210FMA@I3D0
P_=-1ZF)+MLI<TJ D,)5&:*P=[VI<WH-;\^08WZ_@[&@I.[DK[8:?L+$!)+&@NO7R
PR->YV#3C$>5F6IO*"9%4A4W5ZE4SD7;B0M*T7$OC&%8/@),N\K/*1&NNU*352C:7
PM83*#'[3).E5^IK9>%K^&?[&)W&CY11H'RY[^VN'>GICYP$6JX5:RC'22LD+[<+3
P[3KH,-Z%?9-1\>(B!XZD:9@SJCQ6O6TC >->08J0Q5 (AV$DNM)YTQ8B/D+F_&2;
PPW[7QFLNG4 O/@3.CP)6S ]&FT0CY#Q.2V?/M+.VCBCD9[!TT[R&P[ 8:N_SYL,P
P64?/!=K:^@^XVT>[S[HLKQ%%8INZ[WK^VKV=N3'^[NS>K!,5XQ0M4(0'!T@W3@8S
PA_MX![4^BEEL7&]3CB^^CO1.8M>.-^MJ+:5LF;6E3T _A8&?1\@*GVZ@2?^/\[EE
P4S6T@FB4CJQ-[NYR0@OJ\LNKFIWE75/J'.A[Q#RE)1.89@8FC.'6U+'IQV44<Y%.
P%H6(<W[[.<;5:!FR M:(5[-3L++"$KIC@_#-2Q5XE0@__L B+@>-HSHWV+R[A3F3
PY!^ES.ACIHXPOES-%B>0B=1LJ:1S>57N7,[!ONA?VLL;L@U"M9V30LR=I&TH1Y&(
P\C/D",WN=(.I090.!'2$<@2L./1GT) GFWOPF&1]%9]]/UE$8D<BKLX[:B4#<$W6
PI^5-.! ]AWO#H7(,=+9S%,/*&&=WU _W_+-I^:<2)?9(L"9:ELG'E)&6[U@?8"6J
PX>[+*GFCW#\5/)E)6B6WP8A.6=I#)T>9TOG>6@H>?!^G;N>6TQH:IJ"OY[YV\K'O
P4O:3<0)^KU 1B:@LG[:8[$N+QPT42CHT,B"?WV# :/[OK)V6'4L-(8FUIP]Z,LZF
PJ%/!L'6/ 9+5XFL.(> O^=OZ@[I# J3F450;QOY^LR+5J1]S$'B=858Q"\=5)X^+
P0'W=ZK8+QFC!$PM8>M@$GZ'J*7DKUU[8)KL*X[:R@)#BFB*7[+)![IN8!/8O-HS:
P,-]<;Y!_-,+-;^HH?!K!LVJ'3U:]V[U8XD%<\V_\V,Q@VD\OWWDSG_W0@[Y?]N:1
P53:.YR&\%^9WRSR"P!^Q=?.2<3.4^1L 8"(\WL@9.&!7FVUTF!@&ERWI6(O>\7<X
P<PG9?<9F8(.ZN-FY[CSW9!>OG9UGI@K'@7@I]2NMU> M&N^Q/ P=36X3[!!\L[RI
PI[!I@<M7OOPHMH779DP(6B0OFMMEV/'ZF_?Y -;=Q:3^*MF\,6@IH/3:YU6<E\R>
P?Z*@L,MMNK6"'8#OT*Z(4-&;R',6VB_!++D6LT@B;?OO4%"CZ2\44SK$3D1IX*%%
P>PPIXZ'J]RNWZ?$W\%G;+L*\&?P2XYY] NE9T(>(<=&K$@Z%5@><,+6VK["@[/D&
P@(W+QPC3=X7^WW9!+36=E_'XKE/&0+1[%[Z*[!X0CE,&7AE1X)Z"#X/MN5"<N M=
PF&X6"4#$[1V:6,H )BFL_/NIPT0Q^*0[-ES-_AO'%$4CCN&S21+F1U&(C<+2YWQL
P[@A1)RX+7$D(%+D>MP,?'#TBQ#&,T8VWI.%IPVM(JT:5(@:&&F#RV<$RJ9?:^D6>
P@:<\P7._V,JT$44A (OP1:K@&HJIUJM:AQ"$4.KI14X]ZU,6.W_VE)X"KMI>^^O?
P>;*$%PT[C>(D]NTE4F=I3ICRDO%A8405M#2&_UD6;Y,?X*Q'4N"T_QKSODZS4[PX
P75A)<44G/>F7.N@QHS@V6+SAY/1X?F[K K+LG+AO$7%>HW5?H6Y-S.8D(QXL2A!0
PKMV?![3) W0X5K&4WFRG* %R8C'96(M]@'9=JH*]- PJ"S[4A9WKW&XFP_...$;F
PH-_"SX39\CS.8-:'F-+1(FYMZ^2T%T'0]!K$-<O =T4;NW:KT5FU"/XO>>63K8MW
P\FQ%*#FL> S,Y\3XR+^I1%8*YLA::Q&3>8% +IFT V<8Y>T<J28=MT3-9LC'YR8B
P1%C>6-AQ7;(^5ZEBIBP@73MTC+>'Y)E825 XPS<7UF<*216R=;NU;/:W/K]W#N.G
P!JJ1:5NG?-EFH]F/2C4BKY4NU.;3S[_%)D&X=KBW.OYW"'P:1^E>9BS< [E.]HNE
PPPE'_QFK@\ KN1!GU!,RRZ@,CM*K WKD;MJG>)2I^3EO/SFK0#S'.)8)(0\!V1_8
P3*8\7VT$==UM493U\,H#GC?E@A/@,Q+J"DA'=$%AHZ4\W,YO)DV:2PX=N1KVXV4&
PM.VVAPDEH(NE%I]J52CE(9Q>6@EJ+4&ZA-:W1&#7D).L06)6^U;)]=6>Q'I64#/I
PB<>5Z["@0T(!INP)3B!\ 1I[HZK#U/#[K<_'!G95Z\Q_]"/[/V?^H&XJ5:(W%0-(
P(1+O:V:=0# H],L(2#L0GHBDRS+_16CJE^8844Z/3QD"'D?>J)=L^]CR:NJ8'X@7
PY"E;7-PUE1>BT%U,-=O!'9!Y=@ G3DG.7C/I4,^C\;.64QLV;4A]\@<--K-Q$ -A
PC4Y6_!0@NS8^3Y#[G 3G.%2_C^XJ+*;P61OPR5IKD+ ",#U_FY:RG!B5<7E-NO C
PQ7Y'B9^82TY@1?.VV68[[T33_C)/B,W2P$E8 ]95K("Z VGCLZ0VJM(%/N?2S8H_
P/"2M7;?8?^7!!&T&Q.%*$\ -6C>X.MO+^'C.4@73(#G+LQ="GT>[UTP @PGQU!?A
P*Y(#]Z MC0V<A[V+W6C.:N1'[W[TN^.=L%==<HX5"PGY@1Y[6)3#.Z"8B$J_$SOC
PUW8_Q9557*_ETM)\+X=\M3^8&==YBDT'ND)K+Q\L9@'N0PX&.S5BTXG%:\GE_U&:
P=#Y*@8<G#M&#([#&&,P\K<@M0TJ#+UW8(\C2/R2"T4A@= 3MN/^G-,EPVJ;RBI26
PKN2K#?(YBY3+YE:;6;&U7EWD:P(.K;D\>4<]F9M]4,31LU'^,-L;J8Q;:L,Z )71
PX.;[VF.)NAU&Q5G_J$W;&3/E6'(!./,)I%,-T;L1+SK=ZKD_9F95GVO+.6-2GLOE
PC7*KYP&UID3L-*TG<;I%[6W^@Y&B)8.F^&O[<<IRFV0"1#(?K<R"<V/B](4<Q1JK
P+*C@QOP5!$,T-@4_X6PQ>>-7F$_T 6=0&E_K+^2Z<MJJDCYE03LU(WJ8Z4,I8UP,
P$E O[!A5(C:J@U?A(,%S8"5*#"0E<KO^X+W9N(6$5&PIYY'U&*-9*F</U:%9Q*R$
P>S@T0\_)3TGWN?#]3[R8BHO>]L9,D'+'WI-V4BAC'R.UD(36ER#?2P@HC3(LM)C 
P1'! +6Y4CZZ&[:3U0J#49#VCR[HL4\BW?=V7Q\VU)0K6#NUH1[/-[Q-=V1$VN&;#
P3+C]+VQ.Z(0AEI7S/2/^#.Q^O4;AE2)S*9YEH@Y52UO,O#B7$R^QI?Y3*:XWG<2P
PIK.KB!>SY8TA,]#\T$"7M<APG$J93LTU;D8X[)B44SR!]"HV#3%SR[@_.=;S<Y![
P]LNI4XWD7KPXT\/<,\#E['7=:; DU3@J=9(59BC?K*,C=<84/BX!FO&&L=&=/R='
P=/&S70),K10KMQI"&4LH5\D5_Y*J>+>D[%G/2XS]>9H1[)U6SN$97SS&4%C(Q<W$
P-*'.;+:C\I3 (_RM+>D;D!:AOV.'8M+%3I'R/&^Q18;@ >1GVONE0>E9QUR/R0<\
P;P20*Z%>':"+2$_N E<D_4&%&MN(GX)R&G3-.'I*C%OI6;X[:9=K^#L(!. ,%[7Y
PH2KFCO&S1X6T9"X,)K_3,:)W-(V4.?"%C%.Y=QM4E^;*H0 B_KQSF!''+DK^#&0<
PA2MD6X? K0ZSA:(RL+=%)9-*["]X>Y5O#@AO1?F H,G\:AFL'!0#JFJHY*0KA5XB
PL@- %S%!9S@8*HK9*%C+PL5;K\1:/31%]>D3ZJO186JP6Q:T.$W"PMOL75V[.OZ$
PB5CZO^. 39=CT\6W4R Z-M0OK6D% ]V+%%WY,9GBLT^YOKS9G>!3)?A96CK>O6(S
PG^TB4RX=,&2G]%(/,2\R(5F7T<FYXGD%C84TFR3 +ZB= 5DD4I);UB=7O,N>N57P
PB>*[_C$UMZ7$/Q'2E6R\$I<6&[/:>5(&*\=]D2-05LCMI+,8#8BMW>8$&,B.3MV)
PD@\@1%A 9H4PAL-ER[[/O.[:A6O?10_]!UST,FS!'9FU_LMY\-ET-2[0'DY&X@6^
PC,,0.Z,EGE%)=L2L)BVXR;TT=991^Y5IJ')*%G[P75> ?$$._[*,%P;NE;0*IJ4X
P6I^TE:*OU1 )WSND@LWZWUAN,1*XC:X123GG!/CHB;*W&DJRT?;9U";;#DN?:NMP
P$Q,U@4HXE@YW4>OX;V_TG@;1$JJ7;]8=OQ<9J(V:16/QUL_E/V_(O=E\?^YPD-/T
P2/U06=P(3R656?^\Z;(0Q/E(!ZCO7IX;=[97$@GK]A=8$2><\%F&H?] %ZLVK<=+
P@/=/V]E=8<ICIJAM^5U(!6XYP?R2&: O\SM6+F _QL2'-=<EQA3&XN ]X?S6R+";
PU%I_I:2$A;.BL7<./1*USM<3-&I(9O(M-7Y9FIQ%9-LF7LU1@PJ?:S/Y%G%+^033
P*PE75<Y_6\G7ASV2>$T@,21(SGOE( N4-?\"A<HO_\'$#5,!>B$Y1;/\1 $C8GG'
PPM$+:/?]=>8O(0,'"!5L4M6$E9B@:T;N:-,AM;\ Y8VHXF[\]R.:Y'MT:92&>+J:
P-^-QY![[CL0@M@&+$!4)_#IS<AK3-B-2I862I3-REU"?DM^1RS%W'RH0057=7S>!
PW87<*X^F%H?;(\Y(^4N&7D6G=#5^6S_:Q/NLQ2C%OP"Z^@=-V0A-5K>WP)J8F,@F
P_.;H](R)LW!F"MY6I<[M#=-PV9U05D>!2WH#7_@=+SNAH\[E/=#%!>RN*SU-Q 3N
P^G>CLX(G'P*/$LB.Q6F=&CS6"/^CY!1\\[VLLD"&ZD.+"II8<89%V.M]Q3]5=4WU
P22T]C\9(>LXH;$$7N\U/PCYU$+_F=GSJ.]%T2K?2,.M-X/^4R)G9*(T1"<+PDT-1
P@I?_KN"V2X:7I.NC-6>$13>U[YI&\OC5_+WPAR0*YAPWFZ'-"_%I&Z.;3?+A5GI+
P?CF!H,AT"#;:2&!SLF1PH#A*'D8<6+LQA]4DNHL=1%+ZR,1UW6'IEY8R8G*F[GT=
P?V)H^WZ\K:6@1!J.-\Q5>7W]FDHW8;NFBH>1#M!V&:#0::IV>Z'.;+= C7!96SSI
PGSC"_S&!ZS2',4EJPPU) $N%*)2:3*4]-<VACZ"T^OLWGHX+CGVZF<_5\[Q ):N=
P<.]Z ;)3'G:P^?HFTFRRCFH(1BH7=L-R/H0$*.K7Y1&'!>BBB7[>\:$&C/8H'2,[
PZ+?'SWB'7?VE)F#<FH)1HC]D+?G+3:;[M#@8?](@'XYGG;N]G[,M54I-!(,F>\)W
PN^7B1I,R(_JE>W%V=/2D+<^:EEK<X#V2\IM9,(S&=^"3P"QF]#$4O,?C/W?]0.\Q
P6MJX^70$-* %#2?Q%#Z,,Q@7(A4VR^T+,N!H^3M$$J0:QDM9:"S4?] RHMQ.^AMJ
P  (Z,-=:"P/EIM9>JO>NH>0N2@CI6FD:D9U#<D&7^8#E(^TPWYR3Q:C9EXM'?;8N
PT7XA#7"D-5-3 R:J^*(>X::?O=V=N"_.P@[=J<D0VR".2)CO7BXNK<E_?%XR^JK^
P7K3!@.#TO?"VA@A326H*K5SGI7KR#9'2' \54%,PF8N>43N]I"_4C'RU)417S_]6
P'\*B]%?N:0EVN_=@_Z?A,]V?0,!!"9LY6^YYYKKWYVUE\^M<KF#S[9;.EWR!].8_
P!*2YDJ)6UVXE%)7F_Z\KO*&K0%2[$TSOEI'FI"9FW0C4K%UU?;DV44"F6_4I*=VA
P4#,7-L0/[G@VG)Y%FC_I3(7'^!21%<1^%0-DX6ET4.VZ>)@5SM-O,_V(]^Y9P.72
PK3\O]$S6X"F4O7J(76<7DV:M.,H4OM6]W!Z(/@3*?Y)(9K2*5,B4G45C=3#Q% AS
P+X9G?UP2J*,S$I6Q:ZKTFXY+;?^Z.J&HIFWXF^$@2.>F)/G9)L1 R.)*2)]=S(.K
PYXA<',"\(AZ=_&C[6W9E#U1WGYH0?6-B9I\)'2@)=T%@4=0K#^+GE=H35@9&WI[-
P01IR941:\40*C#J)+\7,W_8M*K/#J,&N.]_!/=IQ\8%DZO*%ZN\_@QGLS#_K3Q$E
PQ]!=)'IVZ5<?ZTE564Y"F0H#;>2*[A%>^,<) H_O#/_LOV(U5T-WU1A),5%B\*QW
P1Q\513T-3[4'[9RC5E3P,;;8R3/"-<JIP>#UA;A]S8AN&V^,WB$"ICKND)__5-"^
P"=Q&+:2V/ IV@(#Y=.Y9Q'2>&*X25M=J72JV$J\=+F78?=2X^:2/E,3(<0",HKVZ
PRSGRZ&J2XE:4XP$J_&?Y^R?H;0O.'TW3LM8/8_H&_*;JT3IH6"%*3T@MFFEJ!>! 
PLVU3E\Y**+(V[9G&?I-:-+-#PN/%CM(+LD5G^7$?*O\2!-R<+]':@+::+9%81@60
PQO RTX?9BO@G,0(['<\.NR<L( R/C-@48V&W=(9US!YC=!R&Y7S(#'J\R4MWLL3%
P6W@F6.>.92^^FYQX$4VD# T<T4>N:2"0>7/5[P99FV:JQ57IN18"G &!2NM:XK0G
P]S4-@=S! N%;9N#4B'X%:@,177@&7MZ/BN.56C,>+H?P2S!G@.H[F1);-9Z,L"CE
PAGL<;0@&3IBF1B"EAE]S6Z)&%<RY9<SJ6*93P'Y$6ZK3B$S1X#TRR),064S@I\DU
P$^QP!U;<Z)C^GZ.-SCPNY^QTA&G9I&J6_%F;*IUH6P)U;9D>=W?^Z>GG65'Z,$FA
PJ>Q+98L'^[^7 !/#%58KT^V3[WF+H5+^@ T8^A!\[7R(N:[W?B65/7+IC]S(-8H5
P<]X@J$-9>7[)J^\IA:'/OUO*PO2I'1;P^PJ--V7G<#5&RAADJ3%SV'E;_TD =XJI
P+ZUCVYO!6K'8HE(BW1]Z*43RWR%AUF.(D<O<66=M!H]-.9VK4X<HCZ1.W(B#QAX@
PM&$:KO&0D[ _K;R:3'.WE$Y'/'68;]?(R!V2!M"=M,K<R48!%YM,L'CN:$%9X\-$
P_13X74 MA+'QK&<D\)!*TK$1<7T_L]XNTY70@QFMPT#V#7>A1O8; M]HA592KG'C
P K)O2T\=90;,BV3:&L%=QR^;Z;-'O4'@SS9"BG,:51%ED,*'18+*YV1GU=8J49\L
PEVR'P<N4V#"W%8[YS^*O72W[;41DYN6D2R/:V!!KVJCX%'EP"3GTGX^(4#D>L$ON
P5X0"H@VQ<*Z_"6^X6N;'I%J=+!YX]_?%Z'<[.U*B/VBHIN>LFC];K'PU^#VZ6S%A
P5X2"=HGF&BY,N-:WM,X]_'PMPX,^^I57"J*E?.!+R2%O6W@5&JU WZ$ B%*P@H2S
PX,\$N;.NEI!V5[MV"^"_!(V+:"+VD^YNMB!2Q2PKJ'FIGGLE%B6LR);91Q35/A-9
P\GA>45(YU6,0D#_X_X"5&Y@ WV^Y([X+K8S/DY^0OUDI>RR7KZ\W2MC-'I1D33D"
PN91(()":Q OUF_PAV,\8P^_X$T%8RF:<=8IA(R>,+1P[5VV=WWB\IY@VH)YXFW+U
P2'7!#CB8K+PG")RWO1FDE,/SA6?>U^A0;9 12TKU+D^;_HC".^=_MNY! QJ+-X7"
PO8Z?MY6@W0@RI=#%\&K,44>B[\?/Q-+XR*RN[ZITI/]986ZT2?_:%V3 @@2[D(?H
PW OO&@'53/0N,2*GQP!!NOTM$0]ZR9F5+B57T\I4.H>%I]8HT3ML3MUI.&M\,S(?
PI]1256[FXF'DVZF*9=.\AA@WG4V#L&^?>-(-H:?YAH]7YZ MZ@?>NW9;HVE=9*=,
PM-A_/ E2+T8W75NK 4<[ID<# 1E/+4?]1H91-;:'YZR9C N\*E0@N"Y?0&C&3G E
P&5*)F%CFXTXTM527<N"&Z<IG]3GAU6",=QA9HS8-5_G4U\6Y(H/OV936UR((5R+#
PS*SGV17B./.R1 S=7565#SB_1:&]7\5>\--AO/CXT5$6@@IW6M#QAIFS2'DB2C08
P _#'D=NEH::(RRZ)]1A^<N[L5!/8/4103X(*=["EPEH/D0F'=-65J/__BR6T:.'3
PU_N80Y'FQ]3*UJG[ /[L,)C?X",Q@+,<,#VWL\O^2ESP(:]%6DZ/Q9C>D)-3JT$B
PD"RIW\*<J;EY*<?7+!(W_W8FFXT:@G#,+)*BY&U; M$F_.C:(8L4)?>RG8-NO[L-
P/]C[^C:T1-[^RC-4IH@J6SR&D2(W#[B!C(*:PSN+@>:/<UZM:;ARNQ4]F&85N-J.
PHA\,PDNY&?%6G>V:XSLHT>.XXSKFEF*SIT#<8(!H@82SM&VK/(KJ1/NC$+'QV ^P
PAW&J(,7[F[(Q4.+FVBV647SC]'R, PKK&/\+@-6E5MI@Y9R.YR:S.-,*VHA1N0.K
PI&KG.BZETHVJADR@.B97T$-PSX@&9N4;MG0)53F@4D'N-O#'A;)RAZ:(4I'R-]4!
P=Q7DBJ>7<^GB Y[LGU; MHD%'Y9B3;F)%=)D_XUU/#''5HJ"7S,1X); )C5(DC7P
P$;AB3Q(Z HT0H*_1@R*-;ZZL1*B:M4=S"AZ*HAO6KRYCP=#DQ_ ;DTTZ'9;O_0>G
PJL2L@4Q;W7!7GU.@;>*7_5ZGC#]='&%;2DS[X6[_  P+P!+C9>AZ+8T/6L5ROQ60
PFTXTJ!R.20JW<]GP5*.9*]JQ:,BZLTI>D<C?H+(:4OEYV7?X4')FM.PRWY=?9%(Y
P>'!  C=$--/Y$++M2F@=ZG5-68#EI76I(0>R UTQJ:AYX*J?\9+QUT3=,LKNC%1\
P*P9R/)U1.^7TH5)$RR,NV^EUS=9<4?UR=O(I+&A94OP_T %8WOG#L8.,%TPZGE' 
P($@0=-6?N< N\J9@8K2YS-[") N+0RE+B-K_Y_7)DIR=P,B(TJ;0P.%6;(!G8&CE
PU3$4&M]"P^"4Y:9@9STR/K1S M7^[.]>)AE9]/?XI?8CZ7&IU8?(,3RB0E&K/.B-
P@EHN+Q=#%._5!%G.(+QHXQ]RF?U=?<UWF%].HR5PL[X.N@VN'KG^AS$WZ$Y'V4KT
P ]-@-.A"]&PC2R>_]SGE<*66;9PT;L#_37MW((. >OID70_A_":GYKRJNV9V[=G0
P6@.P:7>..@PRD\6NB!D?F.!D,62P,F$]HBSFI%][1:V>52*SO6D19YY)XL^38^W/
P1 /D3=^"!BY LHI_^S$6?G->>GQE',*++O=&@*74.@H< +YM**-'."A549##0Y8-
PR??P\M4CR=&R%9"3.++I7>"*HU2UEE$@)3JKV\%4LPG@E%,4_**>#=]<V3=2A"3'
PYS>PU03"-Z .0F)!(M,&\*?6.&$,F@(A][1S!YIF JGHDJ)79LQPKXL&?!Q@G=B/
P!O*U'6:W($&./6 7@Q%VUS(9M"G11N[Z#B@\^*#++AS]:[5PAQU$+QDZ[$_6=*8R
P]"A@\6OD@Y4Q-85X]QY)HI*T>.+FP=1H'!'PY3=&2PAV;]0=<'\L+:O $ &L9H9+
P2)^KJ6HZ@.G&LQ=].2'XLI2M>]L@!Y8YPEL9P(7GM6XL,27U?_3-5XPKYC+D9G)Q
P'J>.V?'^Q/=Q'6(X;S1]((XZ&!"AM6W*<D16<:Q7ZAZGJ&?T(.KZ#!!Q_1>8;YT@
P]'-*F_A'= C9SRJ!:XM+>)A.XX71>QZ'ESW.OR\BO:EQ\GF2IB/ 6JG/0J]E=!_#
PW/]^+/Y;05V8^NH*'"KM*Q=VS0Q%E=LMMX@3QR\O&CLW=Q4&:$N0MZ)G;<KKC;18
PC].; ,#1R^=>BJW')%!!&)(%Z&R;Z @VVX']TQ>,)M)Z*'-#-:,$+@=@Q9I*HRK+
P(6/?B_KJ?5O0,=$ !C*Y3+Q3W37Z4.7I,#1C(X02*@]APRW[!368%D'<62<#_1)K
P$!BBV#:J.;+((X**I]H$_(OC6:*^1.F8R)ZQV(><1/:4-C((9\V$CA(,X1FROPI 
P9"UAU?81UD$S4 $%C\M$#E2_.W'I.P<!BV9Z#1RP ,YI$SE12*Q#]<WL0M"^)3"L
P?I>#>.Z7[+(FVFMGKH1!(@*T\KT9AT0MQ&ASQ+K#%@ZG?;7=EFS'O4;1F$^6','8
P&Q$63.QU&FV4XA'62  _CM!5#RDU8FTU5QO_IAXC"E%N7/Z@()*LPFBV#!US)6G!
P'PS/7W^(U\MF,DY(X7D(WCSE2GV<SU3EFZD3\YO52M UF<G;SUQ:C9G]R)OM$K(@
PF+)NGLS'Q(OB[4QO5_S,<%&1^%]C/=*!=QL8?CD7+Q1(3Q&M1<L/P^5Q%>S!(N%N
P&?+@R5H9P85HLK;SO8'1?-ID+H#:'T)S@%!C$U9@01J5C*30PL<;A'MD9Q85KL%I
PC_ +VT:MHH "/,@AK'&@@+2%-F%^9YIKF'FFP(T'@;](\^Z.WW+>O?_[D2WCL7&^
P0O<TKUMR6&,?A[2*27+73T',&+L6"0YN6LDY=P+KD(47XQ%P!?_"6ZPQ]V#$:-%H
P/+2J_02IVYM8/=%@1SV@M3.Q?YTL%<3W&HRBC>]]M%J[-K=,/C9TAN'Z'YML-:CA
P6YS)0PGF5/'#!H/!Q1N:[T%H=I&=%)1<X\:-OK2*&T$:M4DFNGNJB'+!Z[G2]0))
PICQ[&*[D "Y4+KGI%[] />2LGLK$/W6O:[/#6](%0Q4P%'U2P?)(*_?LC.+IJ]F-
P3TKVKTN<K%%F<9.'RS8"UVVH(H\0O+S5L]%Z[:T A%9CQ=9O:4"8.+<CMQS;+'KF
PF,:L2Y^A;!2R3^%#?M="-[08L0QO%-08W;"^()>65,=8BH@!ON9*XG"^M&^ZHIW"
P!HX-4![?Z75F 80+]3(10N]NS*NZ1TE+7Z$"-ZD>"9HWDO2D'?OKPI<<T-[GSBU+
P'R>!T57Q'>O/Y(&'#VZOGHZ]# !Y0(,P*Q, LH7:]]D6B*P\TG.5-2ZK#$]R<H@>
P;0@IL,.W47-\M&SZ8D6D?37R25(A ?4CF;SQWM.VK75Y*1+^R)X?I2 UO$2=!.KZ
P?(<86 4X71]V38YKR*,ET8#N78$N)\F=1!76NC<H,$G$,.G?<),-!IFC'B<T8GTX
P .L/MS'Y#THN?2SY8Q)+9+N\N"I#E?NXVC&DN2#*$>7_^CEBXB]/RB3G-$NG12DH
PGMV;%1BRT#GAQ?6SG];)4-&T$,3.S&&9+N@P[DOF?*1M38YBN[A[>A*<53-R0,F3
PWQDI/I\FGWDP6=4+7GX"B,%% I;Y%T8>E+2(7(RW5 M^!V8 9_HD!7HQ98ZD*+8#
PN*$M2A_-W&WY1(L>F\U^D_C$8!=P@E% ($<&# E+F52;7U8Z_F [24*^M#AXW]0G
PK/^^J@]N/6_%=7U RM/\OM5_^R\+"0\_)2UCK*G-%K$];A"OI35/0U.B7_<]HR#7
P?.FUV38MY*%H7!6V1'HY'R/0YHT=27L]X]G7#7C!/1V$9>Z;V$71]$76CR* HAEC
P4_&^+,NT&_/TH *3;-]*DPCQ:PQ@S_\M+".R0PZ%QD3Y2F5^25/0Z:3GW7K[M%I7
P9PLWZ?4L1AD[O0S=QV,STPPDSD3X='*#&7D$2.UD'Z4 )8A@Z=?(UR#8_96R$^_3
PI#[G]PP)6J!;?U_$%RE*P?HU/<&?.),ODY8D\=X\JH0)RVJ%]55\!"%B-'0?/9X3
P]MA+Y -I[!NA7JJQ2AT5M;%T[2U*0H\#,;N0RQ]<J)$  8AK'_J)7"#L&3.^0N6K
P1&8-Z:#'X4/*T WC_@_>^#NJ"JEH?*]%[Z434[PCSV._K^,RMKY^V-<OY0]12(7]
PXI+KFL(R;V[5H2:S#-=^6!S^&5] L\[A8F27OQ0O*VI"5E/Q\C/?WI[F+G1J8UCK
PI'_;VE/UY)W9]SF(N%#M^NYUN91:;-R_5'=RPVM"E^P8DSXV_Y6/846O)85MX*AO
PMKR'9MF,J36N_.3"($ .IME2%.ZJ2>?;3!H"XUC>2BP16QG0V$-?=N 5]DK#0V: 
PU'(I68>OO1";<?MX-W#MVGYK2OA!_O-?F#SW\WR")Y>5:W'^N=83:/*H"/S:[XE?
PV56JK?I<8R!!8MV4QHT3:.WQ(6]D:FWT4BQ6\!I*4>:U^6_4#]%2*I(Y#CB3292=
P4#4+@0<G$7IP,;- G(I/\CJ@NZ^;R8]N \!Y<B6V_>ZG6K5[MY8IW28"[KU'/(-W
PD9G:E64-TW>AHUM$%NEA$94D?+&:2PVVF=.Y<&GO$?ISRDR\]!LI(D7&H\)+IB71
PFZ"J^Q<4!#8UOL-7^\I5R;-CJ=,*.PAP3=!\7B 1B"4CVXK.5SW<#(ATG6TX5T']
PA+*X'WAVOK)?)O[L0 9-'-:>.:1*R (ZD#I"Q6#8-0$YS"Y'QT\DI8F/UV+)8-YS
P5$299VAQO42B')6)Q3ZKOO3,F7?07C7EA98$R-!FV66V"?!KK9*XY;&+-FG2Y0Z0
P$T-#),.]AEI$]6<L[F.Y)O_<:G=?P1@,]J[$%)57<VV:.>,TA?0Q#J>8*70(:Q^U
PD0S<REP[+ TS 8NE7B[40%B(T(<%D'04"C%V[#&E;>UK?#6#W4YPHSR3;W0CONH*
P6O[X)C_:L-=%*N._XHHPUW4A#)A2/6B[&X.AU%?H1+-QX.BWOTU(;?[\S"V)I:"=
P'1\L88"#''1I(_V&>2?F<'H4V0*8^-V)Y,Y^\5WKNGH8T>IBV4O1<TP;.4D6?5C2
P_OMZ!?'I>N5=$22'J,%AF%BPUC@% WBG-3NSX28X75-43H5PZ[(NIDDOL /RE55G
P=4]3M@LZC\ENX/^F+LC-@) G6T&09>9(*O$8PFX-O9^8%QHBMXA @?-!FM=M*%(R
PY'Y3@"U8)EC\M[VA6Y^OJ*:8R#*B(L1N>MQVH:ZQG?DXWE89(YEQ0=0W2G]ZV_5H
PO9+_NBIG&[(D,O_]_1\:C1]K,5IB2N^J_7-,11K#P.;'<$M5\((4J"S>IZN22<(%
PW2\QWC&]Y<I-A8<OHJND<PWL*!N)Z.FO;3HT,HO:Y4OUGJO5AZ8&\4"^)H&2BDF0
P/M>:ZUTYZE*M=]^S+Y"O6_@X?VC>EM\'7J[_PR/JE-BK)+6;TLR3 P47]QODO [(
PLJV?Y7L6:CU9WJ83O,JH?'M.*1-=//:0MKK-M(XG(X+L!6Y%T(*BG_R1M[P\N_:F
P$Z8NS0QF3JI#Q* :!GQFSZQ:/X5N1&N13BT[RD9H^,P2 (S6Y1\K?LI(P!(PEY%G
PI&!E5I6J!8.@WZJ JAZ]X[?TK:^%G2NN$=D>5B28R>'JU%/A9B#@LX*V^+"-@FO>
PTINR#6*W8=U!7I'<XC3JBM]XNC5'RPW>65F!J=7UKC8=78M/*8_;A<7_E4@"V\<=
P/0TM:YG:T1D+I*^7)- J5ALX&MVR:T[%&UWH0@9!$6N%EOZ5)5+]#_6!G1";A;O.
PA"*C+M]PW0 >B"NH6/T*3%(=,G,F%)]'=30L.5HKLR5>P8KZ.5>V=4.DQ &J!@ES
P4? 8<RL0T7,HQ.F7BA_@\XNI+^E<&]]7\?44/BR*HOR_D"X,^8.G4_C@5][KB1":
P74[)N!PK>%-GX31-]H_R:R8>\O915N_RL!Q!LK3$Q!I9U2H)#!'NJ10U,#RF]UH&
PM]"JDAY*/:X(S&UINH]8'48&Y"+L LAEH4<S\[&&$<Z 4;2:*7 +I*[O4]OVP"*Z
P-XN3%OUY#3C23>%,\]/'JUJWLF$P(VMU7C:#OCZWJ*4.ZMF"H.+GCQ]#F_+B6P>!
PCU'>ND90[!PH=B3R$\RIF[!.3"QS6Q[XB'#_&[4+8:+RT(4&%Q43G+=9U7,(M &K
P:]D6J@G0,3;IE1@W/F\L@NJ7TW_ @LE=P=G:H#RQ LNX5,K+#>M2SY9.*ZD+]R,E
PL[:UB:K!VY9-Y11-Z<VB=^EYV-!]4']88PDCA1R/8P6/QV8!Z>]1GC1X7LZ^?3;%
PVG-5Y :&MGCKT)]G$U5F7J4Y-3\'1W5PW[DIV%U2A'!%XA=4D&Z37H5JMM:>%S: 
P!WJ("R6ED*Z0Y3/, ?NOHH&AG.FSE*8 %H%)58::>[.%%.D<<4./F!_]* D@A4^F
PLH'L$C8,L9JGQH;F=:/W/L3%4S0G]50,E7.8CNL\%/QJ%CZ8TUL05 @_\MA]%IXR
PSD$ HN/%;G\2LLS'I?!&Y*MK9:7%3\<?;Q1FBY(^:/Y1)FQDT1F8%$V$-*)][#4.
P"BU_/6=/<M'Y]$>YZ2T(4O*<X=TG(2@#W.W!WO4],<J2[,37K:F<T?V538$S+9:$
P^7EMDZ![>7:CL0D)>B8<Q<!LN$+74S$21NZ_BL-)/-;&(25;A%;PEJ8.(:+L%@:0
PJ:@3<4%TYI0QVQ%.'5]6 1%TS[_C%+>N#5-/QZ3V8?R1BK(FM%C?Y4_5,$B1JYY&
PYY^'%D6CR'#BZCZ'C_2Q^&QHE;4VO!R3^B-\9-= "#A9S)$<[C+]GKGE C7FQ*-[
P>8_5[FR5H7#YFCX+*=;);1VU1U/E._RE-VQC:(NTL;\7<18;#R9XJXTKA.+E/]2F
P8Y5**6B$V+VMJ3&GK6A>A(8XOFRM"GT?3(,#(E^DE'<O2QU4Y7,T&TC1E$W\EW^K
P+N2F/G#C?IX4/NG@XPF=,.[LE':S1]RF&;*CW'V$6JTO8V5*'Z\[WPN[[&Y@(G;$
PJ 7O=%)=21\A4?=-+T\\ZCO*9R, -Y$W*I'9HB3X!\#3,RJ0:F(_*QI^>MN.X,^V
P0+U<[E@08E1/*>I)#9[<.)Q*O76H1&51'<>N6.]N96T'3#_GB0$7K/F259UWI'7-
P*)XR^Q>O(J'9D/"#YP\8@MMZ!@6?F*<@F&$"+.*T[\Y(UE_@544"]*04]A1$/8IT
PWJOQR_#-;*ZK8*@:Y/8^^LR! EHS+*)H"S+CUP@K<(BT^(U;W<QS6'GJ3AB3=GW9
PETR\'N>];LM <5I"\&@;MZ:"X>=B^2R3LT=^J@^A6CAV-Z_Q>?TRXA&<BJKQKQUL
PQXU*+DP"VZX#MK3C0V>V1EQ@1%DBL.B*2U&E=U%D/:?>6[\TR6(E33UF!G? Q>)>
P2=OUY\0^C0_&92N==5:'6<"P5^2+G^&?"BA IHQD]-^-)_J(347G9BX;#1HOG;H8
P?49LX3KOEU[=/6Q<RV93, &5K8_C],;/UF;!$<4BGI:=(Z*+^XXN8I;8:9X993[6
P_X9KU4#,DO#]9I<[V_SKI"L_D9_G3C))UW8;DWZ7('JT&E@KRQ5B&TD$;1[[G5$G
P9"?OE-%U$NM(KOAIF7*A=(Q\,@#D.PCR?#4P5;,SGU/8+ZN%42HT&2\M:3V"#Q4.
PB48\ )+A!^#)H5=Z%NUC;[@Z?ZH#5H":-#AX.:^KY75V-W/3TOHP3NYB-T0?;PT?
P<V>X!Y#[M\V7 %5^\!^(%V^')(<=ZPD'.HV(T"9M*5I6E'E+4'R&#!]SSWV:(;"O
PS7<9OBT&\KNC/XC?MAYKB!F#PHU<EJY (SM4R&<ST(6&B="PX.F?1S%'AV=*<)R^
P/#M:3S;!;6TJ"-*W4@ ^9\;U?-V-# :V."_!+[0*"J67=V%,VJ8HD+CX.$S0&$@8
PQ,*Z$_(#%;7!EA#B6:JG"870UGIY'6; P3]#"4,+C6G\PG\!<85MNJAFR8W9=9CJ
P75F8^^X\^>.#\A-G.1\KW2[8F<2<0]*-]5.@,Z5%285!&]Z&<7^N-;9%8,<#W)8/
PS]+J U("5HSTO@A.(!\)>6/3WACW6N&@S2,C?@=AQ.GN/C_=4I7$-KM9)=R8$[AF
PSP%N1\,M4GXU2Y-#2*IU:7(I6HC(/]7&5DTN;(M'>]E2)=D#IRC%<$9]59<B1<0?
P:^1D!J>@@7-*<;0!-310KQ4EI?9='?/,R*'7,8'U#\]I_NC[]2(H%""_<C/DA*-K
PM55Q8\<0*'KG_-49=<4#DDF^TL47*X$\;BP_4X)&H9UG1&O\[Z_VNP-<[P.X@6US
PV-I*0?AZ"F:Y9_5#6@FI<3OI52-5$^W(QW'"W*=G*$CE&9)@88Q=2J^/@RQ=?+KT
P^/:NB-@:]*V8Q33$FE)_]SQ4O% !!$DF2R'P(&L&Y48N:H0@/*L9QBGLMQ\LC0HT
P8O+]FEQXJ+Q1B;_F?"9@W&)C$]0LL9,I'0J<KOR4P[_ [I'T89S5-\56EH)_JFDW
PA.\W9H #\4H[!?>:'$P/IE^$/SH*,U1V=D)7ZH%H_E7:[E\=6]^]/14@L.8+GO^D
P'.2'<0+FCV6&#4)G,R-T_>I$$!@]_5W$4[ O%&!S -.2M JKDM62"^&V<DZT^I:L
P;/OASQ^Y2]SZ6"0>Y,D)[(KM#U+#;?3@97)MM=K?GQRT-\RG7RIL<\0/XB_KSG,M
P^I0;V& -X@*M/41J6BNVC"ZH'XUW[:S]PR&?VB&KS@ZS&CO^\ )$7(S8]!-_/+,3
P#8&(M1/\$T*,'^FZ7UWB+_,!+/5,>FK WD1KLP<#!_O&/%G+<Y8T  W$P\+>A[?G
P6GL_18EYD*3$J;4Q[F 5=[D(2>^09E)<,A2[K." ^QPX88:GTKLV"PNC(<;!6=9R
PA!_^>X)0GIILD?+AA]AVXB>Q#G#-43F:N!.MJPL'NN3.)KN=*;L<WFA2+B<K1!MI
PXUKAJW(ZO3U-B5E?BH(R5KZ5,5ISM.WA/789LOZTR)Z-YHY:1#PRUS52!<SCI:*3
P35ONQ'\7T510*;OS61\#B$]I/[P;D58YB]@15:>\GC)EH,O=8+6\YKP/#?3=7?IE
P8F/HE$TV?W+;V'7Y?>=U)9V[ZMW@.RY)0&G<=1Y=@+))X:2EW#\@_JQ=S:3X)F8"
P[)64Y0.KSWL&@AGR%G+YV_9ZIBAOC:+L<I'8"*>*-%YH+[FL2=( %W3QCL@C$'\6
PD)SMV?R?A6@2[FE5=$&\&  8WJ"/*D3U^DE]CM*=D]82)Q.0UM=\:@3@S<':GN9>
PFKM/Y=$&?W Z/$UW[\UH27H*?=[:--:!D&O33:6#!)-NTEN# II%1T&]8+7%RN+V
P<Y/#5FB[6K;#V=659F^G; HOXE(\,1/+T"3-:'J^.4\M5>+Q1W*?_>#ZM_+7!DL1
P;&<C3<27RB.8?].Y*;F]-/5!XW43D9]P-K%(XQL:]'.?DF+CC&G&-2@(S<<;,ZU@
PB%D/&&KI0^398K4N5)5JH?H(L9YO^HHL7ZOT8/:'X4\SEHP(-O$_"30APS"&HH1(
P#[2:+J98;NKYE%<$/A=&@($13LZ5@[TO?(AU)_E S^ZJB%3 ^)H&-K_BYIO4$-83
PN]4&RZ!+T!3<^*AF1[0.%.[+4IXG2#ZCH;J ?@30'DN942,0V,% SXRU=L;@S<,4
PG]S2M(*PA"N_Q1]!J/)ZTE?2:_$CBWICD7G:*E^.T" CPK (PPD'[YQ^K1V:[.D]
PJ^ROUM+7D9?;-+00V:R71G-<)]L%&J(;1.8O:CM4,EVO_M+@$*_]LK58S9B ];F0
PD!7'4';]"1&'^DUN5_Y9O>_:%C,O\0\UJ0:?C6P1_2 [ZB['>9Y_(]PHO.8&@'H/
PY-+Q8?3[H5SFW+%NMFJXEL X_N:&7*:=&Z^7GJ[>7+Y8^H_G*"K=Q$,/%K5/4M$)
PJ:K3T0%VC3OM=[*5=$:9(,$GLR1]37_4CL:4E;O7@!U;T$A!JAWEB5:*.3.YT(#0
P.:0BR$6W^.VFD1GP*&G2/Q^164[45PW6+%24199OAJ5L7AT\IF8TZW9MFO7BOCWM
P!4XQ!M3&^8 WD&-!&3?!%"H7J7S W-%,0BS%9%%:E5XVJ9W3AK)L^I05?(Z+)M+L
PW!UI !'39T;(DHG,0"++R:NJ ;M\I_6IOTK?2QQ9VX7T+!.+Y(F''S_"M0VD(#50
P6)]9[#G\R+@"/*9<85B@HLXYA\F_5]JZ 6])%48:6N^\K1'K4=[W.1,=$>&"N<$N
PZ:K5K[+:RQLZ>NA U4RG8"Q7M=M5[>&*0<NK+A=DY963>\5%F]GD4TJS\K9JOW@F
PY52 !$L,7)LZ FV"$06K4?Y-^NW,]1 PV67[F]7D,NNL F^BNZ$=T9\L>=8@&7W5
P*L;)1FTKNFE?@3>.AW(^FC;7Y"/OW-2\S Y]>/NB^!LH6@ F-0/=E5U$H5KJBI$0
P32/$KMF,:M'/QX,!D=0O93#62--73GP8(400E]*1?HZ[)^T54IR60(0 G]DI"R>I
PPX=P/=,K G!5%E>8"?C"_H7PF#2X-:TQ=)BO/O.S_P&]U M)G#>5NFA#$ON<@X6L
P',NC=J.[+CM#3<>JTY JG8%X1*:-<O_#,<<ZM* @.)S*Y%)K!N$1,*R0_U<8L2[K
PQBDCG>'U7&BA&6Q,DY(# "W="W#"7K[ KY;P&6)5EOYB >)*(>8S,5\]/_VV7W6T
P$IAQG;,9@,["F_1N1F=F$<MM?)R7*(WZF]AA'1CIGX\(^;I!=FU:10$2#:V@^B!L
P@=N5:6%-S0W FYLSP*8=A<2EFS4$,,!F&&/3B.;Q?F[_.S1Q&T04(PKE@\AF^;&Q
P>C'&J6NHNB[I9()8K)9R!IO/.!HB[GZ<)<'J@^_O#;>G/%"!H<XI;&\@$D7D[AU*
PFP"^VC6U4A]BCG=PEKGF-(GL.RR&9@AD]UF?:YHP>];O --YFZT#ECN/["'>,+3V
P/6L_K[F_W4"9M6KHK]J1"'!-A;5((-HJ,6K=D-W7MC^7YH.&+4[[[1];  98+U':
P-Y/=UX,1),?M4'!*3"?8&(K.RB:LS'CTX(T-A%#*%LIZ@6+IF7GU7DVAEY\K9)A4
P\WKN656PBQ>05&"R/E>.&4_$K[)21\:85K3*8<PAV0RES#U0OSP+'*?.FR7""*W+
PXC'ZMGMH]28P3$3)XQ=E23!ZAF/>$S>>$DXY/):L=-!?@(E++WA>Z;8\0+GVA-B!
P%=E=PKZR,.VRQ-^!E_<)'>@W(A00I=TUYK:Q]@OF?-2'0R1(ZO"ZKG488Y'_>$P;
PE<%G6LU2/C)MZA2".:3#;;"R'@K$@*JB<H#PL"T@1(9"OEZTA:>Q(]'%7XH45!^0
P#[G6PLQ0=_EP;3.??[7"5_&-322$)-OKDZ\QQF"-03QN@[4D^&KP[CR=CHK?#?#H
PH"0_7<\E?,8!U3LQ&8'W2VB&^7<:@XM7 ^!T]]  !Z.<'%/!18S\1*(R(5)&9$6S
P45O1_3<0B%\0"F Y<UUQT/NJ^'QCG[.G6JE8TCW6KEY2KBKPEETOG.CZ_W=[R</,
PHUAQBFRS8U B\A$HS-S;#4GOP,CXW#5L^&>7ML55;N)LIN"W&#(F!"#+(-Z.A$0%
P5X65;VQE[3&9P?_MAWBWIY/DON.#G= ED"H*<@96<Q^=>7K/99&)';(M@XSDOWP+
P=TP\R/:29#[UJ>M76[]"4S$9"OCH?ZJ7DQHK63](M^K;>3:\Z_R_^'-,C57979DX
PAP(Z"Q:UG5@!B@ TT.E_N9@\FMX5DX-Q1G]\;ETX,]UP.P5KU)>D=[S2/RI,X]W9
P1:%KEQGU3>-2Z&"UL(508!\/8D"4]1.&;HZ<<$!_7HS?*)'K="[%G$BT;P\7A-;=
P*4WF,91WLFN09HAII^V5ALG4KZQJ+U IA^*EJD35MU6+2)QDC)RPYT_$/$N3A,.S
P>1^YCZ#E5$$#A[&W;O%!P2/C6T@D,=$IJ?!F5%DC]0W1YZ#//?%5J2,K>A:!*\YB
PP83S,"D9E$@$:V'37$\KWQ,;T<^2IN;,ZAWPHD$X"C':$A"%883<FU:>N=.^=-K7
P_YEE!27%RN_&W#%6_OD\**JV<EH8P-EP4IHGO4U9^:,GZL"K68++V4!SI51;>[#I
P7SE[%!QX^V&V(SH,I%?)K&O?[H*C=6'7]46_4FPUH1($0K;[[RKO0S\*2VEHA_@<
P\](];@<6$@M%O 2>7T(93&[M_S*?ECR%9'X*85^;H\1'UGI:_NM[1:W,2B/)T3::
P'T=:)=["CY:"UM^%3,O2*?&D#1F"(3+9M6TKU'-TQ/C3>$U^D+,55BD:&+? /+*E
PKB.3M'8?:=?GE-]F+6*K#ZDBF'L&S#HXVP2Z'4M1?@.=?A8960?1<T@7$BZHUSNF
P6[9!I C4=F&"X&_GH])?\B26RL-:FHF_GCL/CJ16A9&HTJEF$IC>_Q:T<\_'E[MT
PO2JQ7C2K*; B"&#P,[I"<#KHO@(KGH=_1DQP?ZJ?DS\3P&WVZINU6_"G]7<5?K>A
PWM'Y2\G-_2!_Q^#M 0*/"ZU_MSBCIS<"9->N^+SY25M;]K_4!LIF!%L4PT/+JJLV
P55YHK03X!21*828UF@/>R0TV,F@$*@<!&ZK-K2 PJ'Z_DWSA9Q I@GB#TY'3<N1T
P_'L^JZ!V#^Q!K&8:'YZN<O"6*2!9-^"P.BKU$T9UG'*658O19E3\/B"]>C3:0 R0
P5OZRU-N-3#NT"11N3SIUVD=CT^;[Z7QZ;&RRJZYN=:6V03T]U_K*"_76^X!!__2)
P8_VC3PSI<K7.!L'[0+ 6"C#;+J4']JK$?'O+9ZPI^7G.D"2F6BAI^=J[U7%VA_3#
P5HH%:Z$9_<=ZZNW7.4C1\Z@/!$PGEJPBV7/C.2"=LZBW&&6AA08H&^K0BG==SG\S
PS6$L'@SD"+9X@WGB5S.PL8415B".3-/1!%$?L2*R+;=C"K05RMVJP!#72<_+M$ +
PCLR31%P5 C>+7EK>?8TY9?#6B/,MU1'#L1DF0 &3DMH!"L,8F#$_:8HRBZJ/.]HG
P\%+ITX.O7TR1)EJ':2 M2FV',&H!3V >I*)?5*HY"2%.?I,8U%S:W;/JG"J16Y:"
P$3D)^[6CG0P&P+-$[O_?5F6XB82Q'4V#_Y_;O043F*'IC#$/8JDPM;>).(_8R,\V
P12KQDNSB')Y#L&03P)5LPS"%);NRSU-YK-ME;Q6EQEC5^GJ'$X5D#*<G NA-KY\P
P3C24@34)G%1L&KX]:OU2/R5*^W9$H\(&9X[:=@&:C<_9:^W+P>E[G= B1N=MG@5%
P7-R'@5,<+';3H9SDGAJAJ>C?_OX(9.M$!U#N5DTR<3_Y4>\6'DQC-_H<R&_6V[ [
PQEHJK\$.<2$<G!&!+ *# Z8R,KA;B7\)7!5\?M:*ZA.L+MOY'][L\'G1 [S6Q#M^
P.I<!EQ<4N=@9J6^DI+<;(\5<DJ$L*S%,:=;#VD&:#5QY).7Q9-3'B5>T#E0*D'YM
P*B7\$F]:<=FS-T'7M&\AH\9_DO7/;-X\!RO2G:0:=YOP3/]=AH<9T\V9)=-BUL(&
P6G]NA<$K=\=<!H?-@!+1?%),IG'--!?R<^Z )K78X7KS!<IZ,:XP"VG/>Z#DO]S?
P^%@Y<L5^VPSI_CIH"C*59I _F-^=Z%P+#(T6W(_Q_78>V=S^BG?<S%[+((ZALK 6
PUUIQ)4A_=@[@HFT00,>H+<@)&>DS4\$-!9T;&\4.ZT&W*-Y-_GU&QAIE2;.B'>+=
P#-HT("EFO]I#!DU-B(4BK(&^\IP7[']B$G-\P5"MIRU@U^1:NMH602>A@+TT<SIQ
PR.>>Z),62O,3!J^<8K2O\W;^ \_:&>5L-8*#9FD1P;KB-.1*-^_:T_03*WG9F#-+
PNCZGWHS6:#)<-";QH GZ%WTI5 Z)DF4'UZYDU&GX.5</V^KB5MO7H"HY3W3JV.=_
P/)IRQ>],ZC\WH>5T/#[</2>I7^_AG)@;=T5)#17FOT@'^^7V+D;\,5_&.7M(EWF]
P%MOBC]RE(8,:,HL16T)S3JL!<QX^>#V=%4WQU@*CN37*+!53<D2C>%^OA??%H,7A
P79A,\8)XL"J/I??[^T_X%/S\NKEC0FN5>PK3'Z"K_(F7G+"X.[@J RAXFZ0CUS$,
PQ+:#'YNE ,GHEIESWN4,F3*BT"FWQ/5$_:0,T$MUK=B<,< 8/)313?FZO)&D[;(I
P]4X]MN7^'+_"W0:5L$>7,MH!131]7_9YMB^0=NS5 ,JZ8)[2]NX*%XU9""/CU%EW
PM #FIPMW ]<_-,[+=]C_Q<WEOO;AY)CE/R]3A%7?JGLMTHA$Q,XW5((/+=7BIAB!
P7AMN+5K-ED2P7@M^]9HX%08BAKI6V^A:&G5PFGPHGO&O;M+/U>A;0 _41JRJO_"/
P#0J\Q8H=8@4\%"OS/PO,.7&D=5H9/ S65"(=]9^,*1?!7=3EDE-.U?J1E1=4FBQ<
PJP_#H(@& L;P2<XRRVL^R09D'G_,$TFG_IS&D6.8#6G?/48'O@)V@S"XBWN#,(?W
P/MTR$U,K7/Q7D8]YIDMJ7:@7*A+W-FH5(\7A50L0L59W8H73IV1.P3=>]SU["Q_P
P-Q@?6G&/G_8H=]%X^2 XS.92:0NDOEFXQ-S]XS1-6RPB@D79O^DAT+220&5Z@2S<
P8ZW61C?\'OQU__KQI88KC8LQZ>US!4%KD0R7=;ZB1!O_"VD24A%;><$>>X04OCOV
PTT.D91P>1@?MX.+,^;V+?AC" @&5]?(>ZYMVFM+.U?09@18Q-#/C+@FA79:Y.LF;
P.E?X6 V*K)="O\;9%9IWKOFXOXXF.N-64:$=*@D7$TI^(:!<1,$#/>2,#1#W>/-&
PI]>W 95GES,3O,#&#.0 S!SOQH];#]J" "$__N0\PS*B*V7TNS\-YZKRX6:UZ++L
PA1FPUX6MF!<N<.WISNCOGL%.=JVS!8LH7"SRK=6XU0FVFK:DL;>0K&K$0OU&EABY
PWU1Q3Q[[1#,@0N(\Q*XM<%R;^::IZ$.31!GB3,UE5LKD1O-3*NH]T]2+1G7==9W,
P*#',^S3W\6=X"U-9L:O9!'LUBO\ELG"C,-#)P.X2278X5^!%#N!])GMU1A2T*C@&
P%CNY096LR''@R)'A7@?6IDS/]BEDJ <H^#EK0JER_.:'.C\J\!<OC7]W9O(JD#XU
PR3[WH9V^<G=D+C2@)<-(1SI>_R'!) G$KI$K7'S(4H9J *&@@Z=*F#*.@K@^"!EX
P272$=\ 2X2B1!P 14K\C32X050(SZ^F"3B]UT9+C+FMGT;"]8_Q<B7'^US55O6<J
P1-[KT(7OBBV*SP\ D0<$*8#UMH/Q*M[1398)F1C/_MN-9-7=LF(:^1Q.0%7O&JT)
PT4I5HG8%]CV^S5%ZA]*RNB)],^+K-7F^VZK,7(0FC0*@5+'O$O9>8F#QM>EV3Q04
P(IA&LWA%_(*A8^K?=C<VJ9A:@=:F!]&K9!A3L4)=?SE8%S+]N!F#"/QB6^_1F":\
PXC;<3-2JJLRHA22FLPGP*D(M?#CNRY54MS\JSM'3H&"J[A&1+ NE7.22_MN=R>2%
PW.#+1*/GI #^DHHG)_$;&W.F^&R]89)"':":R C]))T%SQ5%+)N"7?__H+-SU&;J
PRMIAXKFR5'@&Q9EQ+AV%E7_[M%\/P^MHJ3,7D<7I=I@,Z '@"ADK*H'C1YS%T>MG
P\)RG,5-[.F?+_V*CD]UXA/[Z+C-M,1ZU>;"Q@+4\-$R!]&V:F)'HH,<[9M-H&JVC
PH8_MQ%("H(U<@$D;W%,6X#>26,+"&\C&K-O*O6W9\ZO-2T7>%$MV:RO$P%R]])D*
PYH0=(E@4ON#)DCY\\)\O*,)0,S\$U_P?_:47HM)&V>=*Y&P"".EL204J=["JM'\:
P%OO 2G;B;"X9>QS%MNFB ?7W Y+B4A: 3^^"NHJOT 'M"'M/PC6PO5(>.@-6,*Z7
P.VIM#->SL#C'2S>F,M0.I'Q)*D&+P')1&]1G_#=[$:>VF75TA QMV&GR-EYUGE5G
PN'8?;[N4!+O,Q4N&^BF[_XK!3-YT.7X(W/M?9+><M)I%52;;K%")[;JI ?@79-+-
PW;2=C5M,=3H\GU VQPW6.M%,ZOE.MS3Z[=_J#ZMI3.LR)1\M'8T9[[6,JUWKNM1"
PP\1?Q&;P-]Q8-ENF]T7U6]$CJ\A;8>C($]4W]#?9RV /C:)MFH<(PG?I3&78U4>Q
PA//N!U8YOZ:F<&K '6I31=9/%91:]0Z;.4PH-FG85S2E'-AQ)A07[>5.TLST<;C(
PA3$Z.$Z>2$P(^KL%9.APKKYR:_H-\F+4,WUED)C*/CO5G3\ =!-JKW0V\:)90<1"
P*@<1IX+C0;<'7"860%O$@#6/S$YLZI7$^8QR^20:8)@@?1IE:O#0*_HR$.DR.@&7
PMLO?(1\\RM[C?#C</"7W@=2U-1 AM+FN<].*,JV@F**S#)C0:8F5I#BFT^C,[M N
PD6<NK/T\\EIQ[^S[*;L;YEXNG]7LE1ZKZO*L[AD=K+(H[A+)#S%?8I0M;% +_K;=
PE22N=K,%>'8+L4]$Y\*V-:(G=_WCM%U2W9-_3%+6T',#,B#$QOMG]E7X_H.L[XS9
P3^U\# +66+_!YT$C2\XO@&+][E7;=%F[Q!"O#?TW0#,(M"8BH-]!,AD#C]_ =(9:
PL\D7X<K!/W4(.')G#7Z<>.-18DS,<.&"YG8KF"?79;CMUMICPUP/:W%("%6UN87S
PL$[L1W%6^(M.,NUNI83&YKKTNX,BT-E$\^>!C+>>EXF&LOH*+JF>2@;E.SYW\MUM
P>\/_9B#MR@(KH*=*7:?\8'0HW*!*X:;]DV,;8%Z]*@JV&G!ZK51I:&V>Z&8\]*+1
PIJ#WR_?<W@:4 V\^4Q=^]G D,Z;Y5,4"CT$(VCI 8JASBSZ#8(-/=D5-QJ,EK.VA
P'@]:_9<.((6L:6^-VR*H6C(L,(2SK7<GG21@ :42]R_ YD@L0]O RN#9?G)]$-23
PQX2JZJVYM4K3731G^'<6J'ST1L22:1@-E%VJX?7C*HMA1%55S6"OJT5X&KN"+A/;
PN>\ C=W'C]PEF'DG\9J+?9XS[F.@^LKJO[5VL=?XBXAH&_'?NKZ'@O^S5DW_&&A6
PE(7-]DJLG#X@X=_4_V#?-D\LTZ_YQNG'/:T/)8<_DL]U\P4XNT-_ 9E]SH[T:._Y
PZ=?=:3W/6,=RZ+WQ; _=IC50FZE?H>Q9$[.B"4@NYGE"C<*X%T#,.%)H%SK?&G?7
PY[3,(BK<("I+A5%:B U+TQ(E>=N4D5#A/7MP0M1B(X%^& ]'9M:#-UR^)O?F2S!+
PO]8 ;T\ORO@%%?6B=S6EO;@ K%N($0.0!M^M,:5XA\:9F)&A7/T]:JSBD-E-]#H6
PXQ>GV%W^YF0PKFU>14U54H._M%Y2_\CPT>'T=KVH3AZF5Q=I=V@[JI3G2^3^(K?/
P36L<OEP\*D#\;IL& T[2_P4EMA4M@I)62UG(G-C#;#<(@ZDAV0&F;VK!-6<BA:=-
PLS>F9YF^+L!J,'?_1RX:U(GY?L4R2W8$T$&%7Y!P%<(FP$8GPM8-+/^X[QH^AE)O
PF*C!1B=6E"&F;)?11*?(YO A0.-B<,3$8%!<CZ\K$DUM05\4Y[52]70+8"/SM);9
P?H\%[;=.@0:W%[D6Z\:KM>3;RKFY<FMTVGW=>BQDU+_*4\(B&,B<A9NYF(6IUY"#
P ZRG0@>$R%5M4\^;#K'Y4XAI8K,HD,T/;=6&-Q%!86- ?C<C:U>RY'2DA0>'?WF+
P R5=5B;<BJ@AXVU0\..]6?VYLP<I$\)31>G5!-.,5WT+=V8#J1JEKII)(5=8'K(7
PI.389D,CA.M@R]"/Y>)H]+J<Y2-XL>#-Y_/RLQRM_5LPNZ]G25)N2*J8UB&9D"@(
P*R Q?[W=XOLM+7:3Z7((@^AR6%UGQ]G3/RRGU@1'"@.[UI#Z66(JKGX\"Y:.L/>%
PSI/9P$BT%3620^/VP@!!A$HYBJ4FI++@(7RJ)3VT1OVETJX5_-\L(:S,C#G8X&M@
PUMWI5YX/&6F,BT*./D!C6?Z3 9R=,BD$S\],! (=O>A\]+Z*R:XNU96]OC.Y)!0 
PP[S*=LP0N)!DT"GNQL71O]ZU'/FX7+4RV2B;L[L-C(,$G[L SQP P<.3U%V^,IN;
P]?KP<S*N#>C:]$ZP5@9WW/GP60Q$H-^#BQ!/0N&LY")(O;6&,3;FC X'JQO,H[M/
P.#/0DA*J!]L6U8&E!>"^HBR;W<J@EDX%63/+\28H/4)-ALE_W9.M,Z63>Z@WGV)_
P:<L/-+HA@J9%F:FK [/&"O!\<7D*=[3N@ O;HZTX6&=OO>*@8Q&LN&=0E[LQ+IZ;
PR,,-7$AX]U3&[,G%4X>IFBW6_2E\>OQ2H]]^G#$ZL,M8F6F&!41%*N.1>NV"H*N"
P8SFW3(?DT8.IJATD!#96>&CMLL#=WC$K(6-LBA(.4&-[Q8.XU(ECTX92U%"&QY7D
P39:B.U<G4QS;H&<VD[QX&EZ-JX^C>+X#4UF:'3DD49<:V^,RQ/EO=F>\#]0*0DB,
PW=1+^$Z!C$R"9U*INKD(9)K5X92[7,;B!%7_Y5:E(K&JYTKA&?Y4:V_Z"V6KTH7@
PS(H7C 13*M^+/,*K'G<6GHO1>'#"%)BE7_1&PPZDJGX"GT\2 %R4;]/'$O0)Q<%V
PF&IT/;FPK?FA</T,(CU0C.0+&5 'NBTL32#A(F]-3,(:U:N4,YS &RA(4@^=/^:&
P=6-*"*5/<FA&L\E+&!NH<)]N9-@4%DH#^LG(4>25>05;C:Q"@X?HJWS-+":#[X:Y
P&WJH,M]G,ONN)Q35O3H.7?:V3*KD</M\NQN7)-P ?E5G6I5*Y@L5/ @T W_S(S* 
PVKZV A3NOK1-N\\%O8,@=)?R3N01$XYRO\JKN'HPW<=\B Z03&*FAH3G^ +4O1[9
PX"'Z7I)WJZ*&$BY24WZZN>S-N11'\H:@16:AG(N0LFC6 ,37MOT#7W*C4_AWLM47
P(-8_T$N<"B8;#((%M\#2U4E$G!NE2C?7;H@*%:$@@_5RK)(-FAC+L4G_$XDXNCU7
P#@U"E?-]*\2K1>F!V*8%AL=$K1B_,]*]:1YC)/H5[,JF"6'M?'(D!%<6#[&'O+JR
PZ%QF$COF"-K"%LTAT?-#(A\1W3]:-27:M_=%IMCB90I''F=XP15B^K4>0RJBB(E-
P!J=)A@=D/) X)UC7DV$U #7O';L;][LT, ![]/,:8T /'2.B6UKY<9#IFRD4,N!-
P4H6&QZ;+#L:$^<AT)^.Q%X^N2J2VX)XW5OIP!7C\@VU&AX_J*^G^(<H0C)?=_-JZ
PPLD%5SH*D;C7P;3NT+8WUJH1S_#90]T[OR)/?>:.@W9'*VL51I(^ 2 0AG>7MNCS
PRM FLN?25H99.3-*N*A7*](#\2;&']?E]Q!,C'Q@B2\=KE.C=YG?'ITOE0N5IB6^
P:>EMG#;&'$5UF(7  SD1$MIN\[/OS(09W]&%8GARAHD1V8AU+]E WEP\?>'91+J)
P%*KEJ!8!50*:'<^5U/D8"(,*-O+E!P_21M:=&766'OH>=J?BV1-M%]'MNB:/QTVH
PXP5/:UON7%G!Y@J.&IV$E6PR-FD;021.DKP=N\7S?M;36M).7KVSEM=R1L5$*RLI
PO;:C$ _VQ;2LQ!M\@'^63=MV;F/U;/)UX4'.VNT5V2\#^PKW:W<]OJI+$BI3L AY
P$N8K&PLN_[%I'ECK/C+ :_E_5=;[TB, ?1XC:7?L)[%;= TB\WF<^T8+9[^;VKRG
PY0#![\"861/<!APC92OD>SX&]B)']FN\<R0Y;6;]6FGS^O8@8W^Y$M ST0])[]5B
P<&ID"=L\><T_63U"YV1%].7IT**L4\5<(>@K?43>#I"" :5N%"3. C$31(!]+$-(
P0_8GXS19M_DUJX;N4N$S76(/,D^[,>MWZ+88;;:GA^%6?&16%.KT'W9-+=1]*G5G
P2@_ ",19JFAW$H89O)5744N- 9V[SU>D&0JD-GCPAZU-1^UR_S(2?,%"*ZZH1=NU
P5 4D+>&IM0T4E>W7CJ1K7LJKA!K,&!PL\95T&5[8?0EVM$S% V'2%35$BP]S8O B
PFC@;8GQ7*]X(S38VXB^>Q4L64O41-UQOK8YID>Y82*?M'\SUO]H5&2R4]]^)8E9I
P78Y?>G7IJN0;#I,6[RERZTD67:P,HB!7XA6? ;5@7%(T(W:94[48T!3(+YT,$MRC
P&(47%^V^T#Y\FM17?10F68$D<.#R5Q[M.A3%X56W(X5*RM8*\&K?8-0:Z8Q++G,V
PSCJ#RFV4=_(34HDS=P[EK B\,>_8H:1HU* S^2CZJ8@$4TBA]"199@OC<@E![,FD
P.IPU3W'22O(N+G6%8$L\F_X$0]#"M;SC*/'V0!4C1\MDZ!E$!>R_)\SYAT]$#DWO
P ZHM3KYLK_<!Z .#;@1K8.)5-1</2H #E/:\+%_AP<6 9,L.JP#&ML8PUA1W#[&"
P,<G,:5V)@@WKPAG65(EGVH /X\!88[FH%U-E;>P=)&.N\=P%/&H9+-<,AAJ*HP8D
P*AG/[^^"V<;@6JI\;831?P<:?TE"U78#F%"7*^QM7-94PA7'P(GJMP$2"5<,+Y$C
PQ@+.>S)LO#_-+=_=6G#P^M"5IPV\WK:U);)D*$)X?6U@/DP/KX>2:'&U07IS\CHX
P =V2 <;T;>=\*@^Z5PG4_O>8?"*K_TD!>$*$F,%&LTZ[C;722D30=-ON][@,9/OZ
P_Q(<%(R\-&HAG;- T7<SR4<7J"!RZG(N.^IQ(]WI<@O#1%CEGF'3G!Q9ZE F1^1P
P3Z+5\>9/CVC[CK=)YDQ"6_U =DK2Z6,^0#Y[4_74Y.T<W3UAEZ-0H-$1_24B.TG%
PO%M.R?[&IV%DW7_:[1N0KDSH1!E#]E+5$:-;\H0;5@]YBF 2\3D==S KL?)]=Q)\
P[+Y ]1J8;^_<&H#-G%TH<!5.WCZ&Z^'N ;/J6Y-)WV*92GX+BBJ (?V67Q'54$5Y
PH4O0P/-<_3-&[S)2UXB@H_>'O*%_C\/^"KB<':\9V56 U,#(,%FT[OY^6];:-QZT
PZ*DYGCA1UN0J,-.=V^#P<,8)D0!R6QCFPE2?-ZE>GC!5BW]U"\9,&Y=4!$M;H0ET
P<*M@_"%136983B*Z*?D5&;3;=#,5H%FF<\-..,Z71U V["Q#0XVZ1;EN16":J4JW
PM PF6*OH)Y[\:<\AM%Z@ZIOMD6G:5[ZV?7<XX;,67J,TU$\2,Y%(1Z'!_Y*KPG#\
POLB1GFWU J<4IVN\K7B4TO54MZVB;<,UM =""WI=>'15&](S)F<V-]7BR!3VCA7-
P+!Q[-CIWYM?E=SHEBNXKS' \4G.S0<9@M<LC:2+A,L^&+%>!<L4!A]I#4[[(%;MI
P?\O?:W/H7K (IP5&2"+=B4-];&"?NRI0Y@=#G%97@);"[F7%0[2_'JXS?BZJEJYM
PW0K (UG3M"D1C9YD;VH]QIV>0OL5364/[T8JR+S7DZOKJ99'8/!S842%E"X3MD:7
PF86F).$FDJND%'=$ !.:Z4=;V>4'+I%I4S'E1@I%V#E?LT6.^/4J'"JDH]0P*EAN
P@2/F(FV!C-,5DO;#36O*J-Q^?P# 1"M?1E_2)G_T%Q"$I.*%@QR?J.I?Z"K?E<\P
PUC)H+N.N>Q?>R5(J.XK7@S=NWA3V:9+;.*7)O<?Q,$LY]S!KE[$D0K,\;O$68::H
P:AH%20R\G4WROG8R6I>;;W%:O22VICB\M!I6,/1,5&<Q,(X"W4*P/JB\L)]ZDZG#
P.^65-S%(@8/!:9^XJC=U[/,D7_T'<[@(.1P0187Y=V692=P[F]I!=<]LK#L+V"C]
P,(/VPM$QIT7C)#.^#W*,3MW=28."2)#ZWK4E/S;$>Y*U2#YSN]]$3&&?SQYCWJ52
P+M(ET"!W"^455OL]M5*'AAVX5E-F9 =@;,7HY3AD8]3IR5:,_T)J"+SR]^Q*?.S!
P9'PHYIGJ,_5%FJBX["??Q4&^F%6U@<8HC:T'*3A<2LN)#*:P5<XLW/:SKZFGSRD<
P)3M3_- ,Q*\2B LIK.4\1M.I/O^#"RGMX1::X:+.]YI=PKV96)6_3IGC*3J&'1J6
P+8=D64Z&:IX8QU(IRA$QFF_B"89CE-"M/>,426W:;[P! S1:4>UI00>-P",*3\)E
P"G<J#X+\'#)JU!B6<^\5-$?>5U@4^&O68 A22;Z%_ #'X;*E;+?1#5"3=SHGHCK#
P5B$)QV>'F4DZ4>83/M7@*8/&NA;7F2Q#_,*L=DAY8^RKHE%:4(H^L1LENL3!)^H3
P*Z^N1/V:"$(4%=K!GE\K:@4L+^3/'73&LBJD!#T"=XLW)0&:P'[OY-FKK\.CPA,Q
P2*L[6@UJ1$Y);'6)2GN>V.+@>I^0*$$*ADO\BG];RCY47\>_IWE:+?\D3A9CC#.T
P2DUFB!AW:U2I+K[**D->[$P&#KC7*5-^R;$:]W+;2\\?_N&]G97!^QMRU6O<]T,0
P09NTISS&I)5SPY HI+ A\ZM8>!%?2SL#X(@=9(&H'A!'#T,+?>%$EFL&M# V_Y$(
P(<_ [U:9O?;U0A.GEH.J@6V24&(<S2WDY)>_8N,UX T0O1\B:;RY)O 3F>_#T:> 
P[LW\/W@%<;%H!$KN-\$#'!_5#]\#'0!G L[4I*6+F(\\NA'RGE5E]+4,0WLM)>V;
P+GXJ2@X4;>1Y!&B;&OPF!I-UF*8!$$6NE=A[?EQX/\2#[ B&O<T?'.T1B8:1[0LG
P& W!08U;<!WMVRWVF1:#%PE&\L+R(O#EP#9$\QDO+;?V1:UWA(9H/DV6.Q[,3(]N
PU^8Y/J8DC5@0NKZ>K&.E^KJ\T,60#<3L3D9:.HNI%LV$/F!]77KR%XQ./L)-:%%:
PY\9B&"V:#>-WIX/_%SK +8N>^Z[T9J^5&IW::#F?2 CLKO%TCL"O),;8;P@_X,".
P<50J; G8<1W.P^9Y<S/!RA2O'U?H( \LC9YP[9,OM7^(\)%[IL3/3NWI2<A)4#:]
PZGE" 5,2P]#!FR:JQ8F0<4UR L\QGG:9I@>5Q/I%ON:R6F1CT#"71/I8O*[9$L F
P2/5BST0]N$_XQ/H/\>YJESHWU,H$92F=O"R5>[\]27)0S,CO/KV].Y1'IQF )#FI
PYOZP%?8SJV[W'"C?2*OM]M=B2P0@&8L*S"U*?+ND Q,\P:D9(U(E8G9>#(&BB)V$
P^6LY99?7!@-/_GWUY#$B4%1BXKRW3ND&GJQB6RS-LZ"<TK8S#IWC&H/30>^PH6$E
P9;4KSZA/G$Q.:#MH(NOK \ T>P[@[JL ]25T?\J"O^>?K'HN7!U+LP _;:#UOAJ\
PT8E'7LVT5A7A^W"AO3&>=*4_JO%07^RUW0;J+S?UA@\**R57SWQ6AF65?U38N=G)
PJA<"85 HF [86B'G0>T&3<G8:2=%A?*4:O$@R1X2-S:K#>1QY$3LB$$O 66I?J!B
P7PDC_P=\1^G'0?8O/C@B;N&1<HXVM-07<OY&4J"6RV@B0$NX(@.= ]4!4/'5^[)S
P3=",%O-6SDEEMHS4'[1#4&61>?_P;U*HTO!Q-@R39=Z@QYJSM>(<- (CA8MYDG_X
PUS0OT=&M_0DQFR1OX*^AD"JXPP=S8#G&H!G'^X*@IY/[T2D\+?]N"OO*AWV4,*\*
P)CN^[IES55<(N*\%;DZPTZH.P$_;[6S)Z*"O*^03?-AZ)$:)?%:6;!?9GR06#%>Y
PR$<1WU@:O,SIA0]?M=?43[0%_*##\F)UT_])E"MC/Z;%L&,\\;L/:RMD:;]7,&1>
P&'5T8.#J!LYDU24?4#I2?<DARG:<*[6G8A]6W:G,)0L?L;2XT:\,J[HE?)M?3)M]
PN[%9+HD5+=QY#CL%&:7&;$0]?S$D:@QX!9*:?0E /A0UCGM4,7I D&.C1)>$G^L$
P^5TYA+'G?D+Z7,\PG2L78CM<?_H M@C-D&'CJ'EJX4DS#8551=&TP_R&.LQT69A2
P<)!B[,*"+96>20A)G/)ZX]NB&[8?:D6@&[3,^9SK:)'OV(]F/#NM%>_A"@#,,!F&
P<'$KM#9]QQ$911L-5#IYXGF$D.K>NL2H<^[EGR1B]>"YF</0GOB3"6"TBRH!L]8[
P!>%@]*QIWQABB^!<1&OC/N"Z.H$,$G@%-42 O<WJT\TZ9=LX_I0.I%%-:EGZ8';U
P:PB5I56-A;(DQMY(" "D\8>*.Y-"EI,+<[AYOB?S+;UJ"S_TK),*T;M_+% 3QL=7
PZS"KP 1,\&&*)L/,PA?OFA3NC^@#EAZUCN5*L+E_Q)O2.CS?K\9]S7BC.Q)DL6C$
PO%.B4V^^K-3K&A[.P2\[(5@\ *'BC*EKT2I??XH'P>DNN^IGP+J^U98C!"W;[MY'
PH?7A<QKS"14]M)H9/5S1SH;6;*B5IVL=50E>V(>;-OI$JMXR_Q;LNL<ZRBK\LM1>
PC^=HYV2L6&U ?=$N:'?/Y#<\2#4V5W!2PS&<N-"F>^M8UQY(TY$0N0 CCDBL5%H&
P,O=T+W3;S5^.HF0TY_.9;+<"?&J+"/@WX!G)%'D!H\ABE+L>"GD65%OB!$>"W)[<
P(;J[JP*.+RBD9S FB([L6O4[,437*OM/VF0,+M/SNY\92221\%8?8!F@>M$QQ.F"
PNAU*NP'RZ6B56GK^%!'+%J84?R;CV"Y>N]<,2-'S@!?CYK6)H-!'I!*A +DG >'F
PZIAS.K.?#MN.O,50GHB7S7"\LXX<?P1%FAZ';ASO3N'GUU]R :/Z3L>+[?%Y;-%G
P] X< !+-7QV6Y.<'G8,_>@SC;#K+/X2ZHI8Q:41(71_PU&<KP6XK>Z(UUWTLQY"G
PAPLPDT89(COPVUZHZAO%5@JU?X/J3/:C(^@8?!),JGVE-SF:&545$":L$B) @'4N
P"80:1&&L34 ]M_R#YEI!_% )&F#G<=/O;15"W>:O\"J&9."'S#_40RR"1B+U3W/7
P((D9XGMPH*1N6.<NP1URFH^\_5R61.K5U%O:KSG,2B#_OC!EPAGM /_%LHR[_GK2
PKFL44/I'$#V7,.(NVX1-GJL%EK8S3M8OL_[P";?:,49]IX+)^A/5U+3O+5P-[D)F
PVDX"K5FM'9ZS&*)?Q9P@M$ !LUP@+FT"E5$],#;"&,;-&:BXNZTE3RKFDD"&A]&@
PB?#T<.V_BL6J\I:/("_*OG ?::O H5C]*KD('=W)]^V@IN-N=6%\;.)/T?UNMH<R
P<NOK680S1K&R*5:LU(&JZJ-5L^YW7N"ST Z$PUV5XZ2MG3FU)?N$8G9X)VKB2(,@
P/*SD2M74<^%ZMQGH'9<!^0UR7T2$UB-C&8,C,:P@^%A?PE#B3,<X6?B.I-O%%8%T
PA/"#$1HZW/WA+AVJ'KSH)IQ_"'K>HC@<&GH-81>*5X6SIVD%9]KE:DWFB4.:WE.;
PYOU*D+KK/6:N;>[J;#?;(289%:JK*79SFOB&MI_>FD!+ U$HE$1IF6!>[+H"J;N?
PX\R[$BT\0@0]32\5UL8C7F(,!(C!?;OME)AKQ=ZBGC(WD%#%0@J&1$CT4-I^'!&W
P*__,PK;2E2[L3\W?FREI:)RC>2F4[B"[#9&>EB61^1I9YP!UQ+:SRY;_+B)F[,ZM
P$&W*#^-NDV!))H A!E9< 1;*+O/#GYLL;*OS/Z*+33[,(6<$_8_#J=<%MC=G<(VU
PZ "*%EIB-G+S0LT08-.R&QDG$>^/VDN.PA]-" -W'2Y^D>?&B;"2-QI)"A;YL0"R
P1L;]&CV>GOO?Q*SQ8WL9^9L&5^OD1&R7O!"862LB%*%(:A[:&\4I=<S0 -I_!\TZ
PXRLAA"5/FW0JM=U;W!RS]^#WSP;G3;&6^A 7L2DZ?U@_2<]Y)F_=OO)%I-\A@C44
P7D_> [M+IJ:=D==6O1S=$-;G&FM\'J^ZNYH1X:6HUDSGG%"!E:>,\+#"[_*X["**
P^,@U0AVM?\4BUE[D38$6/'L!3:S"RCB^ELU*;2!U1'CCO.;V3];;)WZHH=@(_E5#
P0[?SB#O12JP(%JS5HGT+F'JD/(*JHYVHC)<JJVC4/+1.E;+;50C%1P_+(:/P:/\E
P])."0FM,F*$7\N)IW7#LF,/R/PU@;?8K04]8\4YN0O5OVG_4[5J[3+-P)THL7O:S
P?J;J!.IVO7LT'VU54\S,_X@11NGX\U;4,:S.27!*%<3<G3J!@3"/E&:&EG39">V9
P":(RU\W95U<WPRLFT)A8;_^$PP"6 (2"P,V2*'827PKT,?#,2TR5M"D5)E76RA>J
P5%.QU5RZ2QEIBY9]V[U31-U;CO$\4^GAFWJYY79"H\5_<(72=T8+EY"=:=<=/HA-
P@-BYOQEC1ZF7 I]S@860;&6?,W,V$T\RC,7W*A61X4HXS[:SD[4#SAA;RUR1H1H3
P&[M#J>YQ+T*F3;.I00H;K8&+SCTVESO]]\#'5O!3;NT&([YM5&2P5*^):4>_NS&D
P$:7/NRK@VX_$\2$JT1Z0@I->/2JGN7-3LI)H:8@OI\F-EN&"I0E#%WPI]2PO0RZ6
P)2Y@1C [11Q8760T(,X(K8>>HCY W>5+NU5I5/ ?,U.D=37$,3:/'H!@!S3K/J$L
P$"Z; +0@3$U0I<\ )J3E,BK3F)WH!]PZ[D#I]NX.V0%.<X'/MT]E-UXRSRD A969
POZ!=] -]11 OOZ@'>"2ZU?Y3@.QY=*K"B; *?"F/RXY0M^X4Z8+8S$369%7,/_C_
P.S6<POW:241Y@].LO30!J2:#*J0L#_'*#SUS*3T5T)^CQQ4ZMA@^293%I!',9I(W
P_"B&S%H/GTT0;=VK8XY],557%PTZ=4U;"G+MI<\4LU#IX$QB$E#PK\GXHEKOP(A 
P,Q>#T]K$&?;9Z8Q+0%S,.G#IY\<(DEJ8M0^VQ$642C_5\\!:I!>*#4YE4MT%4;IK
P%O&HI<[<.%!292O*C9Q)3&)-M-]]M-=][U ;T>.M&<1A 9 QT[[(US"D4T*6'/H$
PKS51_/;:?W(R&82'Z"],VRUQF>\Y4OH5IRDB2,Y4;3X@ DMMX"WN2X0,W:&#20%X
PHQE/D<"WQDHS.O:Y7[T>+'3&:FTS\CXQ(,#[>%>9.LWT!/HUPZ-*5AV_5-U5R;&'
PQMH:Q9"U!S,%9LR*[O&$;XY][,;.N@87-QY=;W>[$*U$KZ[]"L]?Z\&&@8YA5Y;.
P<F.@%9QU765_&TK$SS2YRMVJV9#P$6$:G@*)K#6,Q$<;QKK]J-O?Q"AE>7YA9B!@
PSDH*C<!OUU&S:FA/0G,WEWS-M6&!^$P6T#<MY#Q2<6"05"2QQ!2B2*'U.M5<<4J[
P+T]$#<,U^:=FXFY*3I&OX-C@DSMB4Z1Q,/A-N<&^6*BU]O@?*PU  6#S4W2;E4-D
PTZ<[MS)]W>@CL+#%[Y->C-%_(D_J_.WRT(PU>R'C@O&(KBQ+3PS<2EV+79]3CZ#,
PZH&+Z5J!T/Y6LL*N%6GE!YJ2Q/?.-/.GCZX8\/K=?D.2CU,._2SBVV6@5Z_D/!.L
P>Y"6@_S ?9]>V^/\;"03U1Q6;";,H0:5,K8,:"JMQ6*Q+M9-)9@<!B4-'<-OWC8C
PQBR\]_O<[#(_;T3*9RQ(S8A+>>%-MHPO4A"_J@=3#D51RRF=R,O?.R"=@IQCGE<1
P_V*2D!AAM91?5[Z<NT#!)/W/AJ>]GE5E(_F0TCNCR.A7L8)4"@K@4T4F,1+1EW\!
P+/KK0WC5!I<7=6D2(E%L^;HJ18$R!.M=IRS.-WYTNWV'!/*L&6(WS[\[XM^V#?4D
P?^69_I@-D^OC0G<*$O1N@&;6^>Q:)2S^-.H# &D5'R6<DJ:!\D!D:5D=XJP N,J"
P?\*^8%2:504-4F<:LI$EPM%.K9D@@O+)M.#AJ[/*<]<IY>'F*;$&7/Q?[4W-Z^BF
P7L#A/.&#3\8?QR7(EK&:)AJ*<A-%@?-A7O9+^_&,8<T )H9;[U2J"4=DX!?F5!F0
PDDN-\5'AIBY4VJ8X=\E+28D )D>C%N9_F^&J!<!D:48A4+6;Q7?BSYO**84&!SKZ
P'Z_959*DV[Y5+F+!V)&PO.3WSKPH+Y7^ON# ,\INU<52!Y_P]P#QB^];4@0B_#/C
PTF8Q#6GN,D_'*+0R6$='UB.M\"5W80G88Z>PUCB&Y3P93=HL[+?N*7<V@#U$=,DQ
P/O4.Q-4S-*3U<(;R<G#%+LE3<@;OKG%12NL\+_I,62)6.$533$:WMVTDT>"D34?Z
PN1<8-_?PB2=KX[BGJ2]^Z'>E.4V ]<<$5Q%S 0M4% #H-S>RYC9SC)TDV8Z6-Q@E
P=IPE+F2E^RB+.&D*RW:!B2@QM]U&'ZU/X06/D+"IVTN-A]<?N*,I)SZ4WPDG^Y"F
P-BW=,KZ=%71+7-#^31DS>.N^P2SRCS7[&A34:B31/-]+LLCV'_:S>&&P6!&?L;_ 
PGE^6M3I1WURT"6IEES^A#U4SE$TAA2">W!SQEV:>!.K1[SEL.0W,K?!4J! #69^;
PW?IG$9_'D14MN! =,06M,J*OZY5X/7NC8"I2I 796V\#J@V&Q-*0M9K  AS@ ^Q*
PB(T:'+AV%ERV,MZW]&;HYUD=*:COQ3'9,Y6N<L*0]X,[+JJ^4T0(!HUZZ9D& VWT
PK!U?KHGYF)G #$KUW?J44]'FYPPB;3*,.^>S[JD8*F]N+8V9F0FPZ \[H(/VU7\-
PQ%S9?GM1R)AD/=Y^+F):KABE9(@F+ !N]SSNI[< <6P@/;@DY$5;?<;VS;>'2NL4
P$:>S^_P/B.L1.,N[^=C)/\89#.8<OXZJ8K)LM>L8^.MDMLK=LJ^XC<*$GZ_@J$MH
PPD&QE1JO%F%D)#S;ES"YP*'S+ '=\2V<:*,$]?TSH_IG6R/EUG.]5U>_B8-/KEUH
PII,\>Z$#@Z*? &K HM] HGL2='DK\/1L7&9?3D5-5,?*]R%<9N@$17>,\P+@SD5,
P: X8!KZMIF+@7YK+12$%^2]+'#WW3&@"0TF;?!VUBN53S8[,W /CR1"WR!#31,Y=
P<46\17/9_K%+,:?+2F3NY_@W#4+<4I(C:MKQ2.&G."<[[ N"T=22!NGE2R#YFJ4M
P'Z6J4/0>+03?"_M104%/*J=6+8;^EPUX!&!'7[)JC*.AD9)6]N:'X4=)3 ,8XVW[
P9J]OCK&_\NA"S:5VU:-'_:']:LG%LR#[Z.X*\8(I+19$[@FO[] B76!<.:THSLDF
PRE4Q=8<[CIG1^WM_T-W! )9=(C._'G1#JM*0^_=4N15##K;226SJ5AS(QM#FK6$A
P<]I-IJ,YX.X[@']@L1 ESD*&#[IUULG(([IC(E4?-YE8^*2P38079*7OG0NMTE4"
PI2TT-M4HSQRG$&8VCB0@@@;8GX^NN?5]W5./F-D!7UZ=FS]E'$S:LT')01'3([EP
PD,V[F55(@Y<S_KRKV$<$LMBM(RCT[#R.*,7WL=?A%G'C^J7J8K-I[^T;S94O;3;*
P7^^/FAH/[.2+EPA5>8J!TA1PO6*V0L_;('J%J0.95-OB-L:==4MPLMN(K2!E/*  
PD@(,QL&I\]S];ZFD(?:V%(Q>^&XTH%\TVA2<^.V*>F/%[$?G^D3R_ 2\OVF+91RW
P#(I",X-:#-W58=W+-R]J:((9O4R52;$5V/]=0E1+'OC*Q4^D EQ01E)2!Z>+N8-G
P$H4OX@ R4'CVU'RJ^E2)*TBU&4^//J>P(^+OSGCXM)Q9F9)+&-(((5=@=GO/ZZ!$
P.Y)]!Z$R:1D@:<58T#=%=1=0!-RL+7JMPL4F;O<!4"I=K.XVQZ8GH=Q"'YN!=Q9<
PD^0?>6$\PJU-'OW5B?P.\GD=&]ET('@"B2;@*GXQ??G:HZ+GT8K&\5TZX%&ZR(7W
PBFJFZCO9)T'\I'1N!9ZF7N4,N!P7/%L/1["9($B;=R (^WD>WA"YU]8.>[J?TH8Q
P+\H)7UJOR.WC\T*%/:JZBS54XGI,5*1PGX[4V+(:B,$R_&EBCN@ZN4PF%$HCG08&
PJD+3"/L];&[*2[SJ?0C1=>:?.K \D4MQ*L[9UN<>;HY0* )Z4^G?472=RS,P//$V
PSH F%) <W[S#A%*1N8D"GNQRGOMBGF!<+,&K_.;$HI[1RX2*2P[#-UT>5&Q-P/'Z
P'^,Z0R)*]N4@C.R<59^L/-.0'%%8]^W!)P&>*CEZ*,[B&CTZ77C/V^$FCB)(&^4C
PWV"DL9V%.\9NM"1Z2?'>+!+^ =Q8REV8"^%"J&.D2+54!][ZO(_!(39!$EH@T4TU
P^_WC.V>=3A7[WW0>6L^GY5/\HU.':@'DXTILV &J_JR3R FDI;H[H%K9\]XOH!/<
PV4!FQK)6!Z?@(:F/C?>7I2$O6 (IUV@:=.R_G0%E?\B5#:]MA1$0"@)"M1NKP7/&
P9ZB\7,U4%>-Y)Y_ <^]>X'4/5FBX]%,Q!U!%JJ,OS0:O'LJN>1S]L(;8-(,=N*8S
PYR+8&F!YADA+J^(-Q/82  WO67@LBX0HE;T$0@J6)EV&3(I#"7A<>W[2U4J'2,A-
P=S^JO]-.W4RBRE?T+]_3\?<E$,ERMO=0E#RQ<]8ZN,V9YQ-G;"P-45010."Q1_]>
PC>7S:)HT]6?3L(U\O,$Y'\6J3 @V\;BA64]'+8*82IEVI#?Z48?NE@]S^'1(:BI8
PDZ@A84)[K:;/4PK+9LF&1U),>I>\\\_>4W"%>U]L^IR9Y[P6&^&6?8U_LE2'M.!-
PKU8>4S&*A<@ J2Z:';CC4#<)U0+SJ3E^RH"_A9,LY-[;0&K9^H/*ER,>_'V/*25K
P9%._=LU+F&(76U]?JX@VR[[XK%N,):\KK+LWIYH3';CP'$UKP&[\)C3..OZG2GE7
PU>/D%A:K2&H1TF:LB,'"=:X#*,Z :OQ]C2#?^\-LV7CWUW2$"B7D/US:8C"KK5^,
P^PO[N:W">/$SK*:!'2B6L"X7@5[4!*"F?(HB/+NEB(CX$A=$AXJO;;EFN$PA>TGZ
PBB,9XR#LH+7</@W/V)4[.CVXER^\?L+N-'NLT]BZ>BL'45'('$(?T_?C]7ZF?BRA
P^2S&=,2"43*>- ACK32@1CG]P$BPH=+?^"\N<8"XCX9C[)'YLM5D_4C5-CEK =NX
P$<9&AV^%?_"^^$AG#MFK+#L7&:D2/]*#0CEB(T9'B.1LB>PEN9,P^MTVI\*C; \C
P?K)SJF,^\H^,VDR5;';%7.->W=.&%JJ,?+=D#N[CUIT);W7PDA09 $&TN236J --
P\= 7W\[^P3G>!>YL4[D_=S[UAO34"9X6]7>MX$GSQJMM$J/HX-[W6^F3,E:&?;$A
PNFG (!5#>CQ=A,MW<287M_(!*T(&&'L=C?U=ROY'L+@>0JGMO-9<JDR+OC6KS6RT
P\PY0WE"#T$;N.N1^SXY=#^.D^!J"5/KC;#WDO!RND94M3R^]<E)VP!$T'%XY;/R+
P\<[JUZUKFR1_'3T.]^K+0<TQX]2&VZ?I<%B-![M"T(S7@'?QW=;!O0(9'6,G\CH2
P@,>;)(R/T5[U^.:(0A&<GFQ2HFP\8_/N\/K=/AG(> BC&Q<0UWF8#W]%:6.=A13_
POSHOJC! ;907W<LUK";-HI.C?H%WFN $7.*RWNR#P5#L/TKE8EEH:^>UR>#?[_W-
P(W.IU+[VL2:*6>W@W5ZL:RFULK*Y#19^KUI=[<"FSEU6LQ;;;#GO3I-1OP#S,WLV
PC2W#E-YRY5H^6^A!UY,'(RT<&A>6T"P;^KJX;!O0--7N.]9Q3.-#;GPU?8MC>$,T
P<1UG9O].(XDR=A)IW\CAI01B H(<$HPFB$Y S-'4(VW<S_$1PH7DW,V,NB4^TDB_
PJ6'AH,QR8'0KK@0RIJ83$OAS7UD$@F^Z5DWY*V38:\- 7Y(6@Q@]"SC\(R!.2/7W
P!3S-I1])J!8CMC4:J8?O>1$HP?\^W03$?M"QND6JVD^]&LCVXG4.!PSQ$U_ -,,"
P/MA.!\$:BE+&XE'ELLX+=\N598->@U,.L;^C])D_R#*I4$=O<-J),"KI X $:<SY
P9<IY?TKO'2$JQ(X4HV<;2?K6(_GV/AE?]:9(+^@D=]^ZE06E#Z+51Y2WLB'&GKN'
PA\M3=7%0_'X4#B$M-=MV4I*2_)T,-+Q@3[%\>>[.+)LLYNK;-MA7%L"+W;M[GO]P
P\I R*YW'QESAO@:AA*WWJB)$*H>Q%0#E3L60PR3F_W%/5B,1NYATJ$T7HCGGL'D?
P@2BZQ7'4.:/"X/@/$9P9@SB<9.W\7HN([55_-=94)%#-72]:3VXD5=).IP*],%]3
P\ _L,O*[^]:NA^SVC.S;)7NU'U0K, C9^73"Y5EK,D(ZLPIL7*YC$' 3HM-1/Z^ 
PL)>DCP$DI\8,%K>3Y+8(AB?N=JANTD_L6,+,G.-9I)=X)R+U9"#\@TYQ';?VG:X2
P]#++XNC@>"W"L;W8[JG\;RS*H9=)^U:JM0-/@9]+ZT6BO>_;W=.1AN]E:&_:88@F
P,@,5O_@,>'5[T\^<AYUB#<=.@]X-_02[YS<UAI6_-6%5,<I1=J&LW!UUS)L*#DB9
PMQD%&+8V[\]+*W!:@< TF<X#(LG4!#(4!+.ZJWF=(KRM6XK_NBG4R-/0;QUYF:E@
PI/#)TBB^? J>$/'IFZ<@;7N6Z/>J$T"=:<""$_DZZU1/;(?PZ\C[IN52"KUP\(['
P*)&AV_A8"JWGD(_^Z^K40#YK0#E1LKX/+\<5;K&*_.X^$#[6"2-ON^N:]:,/N!AW
P@=1JJ_L)11CLS-Y- B[;C[[:?W45^D]>I&XE_=G20YBDM%E5CV'C^LL'.$-UTV\J
P?\].=;:^/$C9J0J+E$W_PUSK0- "A-*\E>1*$A+3:7E/EIOE9K?S7%ZA$!2?RWF 
P@> R ;@@48*:0_"<.0XP2"^_JM/$"GYL_D]4J2TTQ'CA"M!HKBQR]DL#7O@%64WJ
P*KZNO^* =3SUN(GLQ;-[IWT8--UIGN4[@=<;5G=2MU8*SXU]"@2^_)ZFKXXNAI2\
PB"N(.TSUZ<$$6N(E^G<]*J(!3=/^J@ M8^-?QP?63 V<A02!FSV)/XGY_^3D2Z/G
PJ!_Z_*CL(.6NOXK;+JHE/:.;?;!2O(:E+]2. *3HV*S0&G1\(2VITS"]@BG#5974
P[)$EAP4M5D4Y;U:PIMY8&=/6Z91'^?\7Y6G.X+.(X+FMAZU8"WFIO[L]+\X[8:#6
P\ECDBQ9BQP] Q,[>=8JK$#)\,3>.FNC*F:U6"=P<P8N%=H#B*ER-$C_!=QZ:4\#)
P9<C$4N%16 ^XN>+0!#))'=9EF/#+36QBU1,!^LS ##18(=P<$_K=>I+3IU9I*SM%
P'8=BN;#BBC'+"ZFAJZ*ZU\;BHM@94GF>(%JRM,I-.D%QI!-J?3"R;US_M/W@AK9Z
PV0*AI+B-B@T\B9(#<%7),NS)N02>"RY-/2X=0\*[&1+L.54W8=;^N&NL]8%KLU$1
PKID-,+L%X^!':>A^1O "Z^X3^-Z,>FPC58^,X\S5L!/IGHK!SL)@36(GT.M)>%I<
P&>JN1JR)6:.)]D.#M74%Z$JP ![O^6G<@*='0LT(&[IKN75"W&1-&PJ[$5=DXHR1
P,<2R%XK//AAL2W@3<Y'%9C(=+AC$QX>B$.3FX$I8U9RA[Z:Z11'[7D,;8,=2=NF/
PU\D%<.\"%&TQ=.M6DS?]+1RUO,0MB V5=\//2&* $U,W@-P7F$LOZY55H+ ISA*$
PG.D H(2S$DWW3G>/9.E/%)/..)K,'X/ "9IDJ$74(+(T2,-O.UJ?7"R8C(=9H5TH
PPTF7N\*D9+C;R<ZER.]8EU\5_19YFW=3)SB4?P-M%GK//TLHQ=1KN2PP5W(<9QS?
P/?!%E]# W7;L8SR2/QARE6J6MQHRKYV,VP.VKM^J+\.K0O0SO#]+DAV4,&&JCO.3
P9?ZG2%H+?ZC=[M<_4 B1=/ 4+KXO?<X5?L_G]9Z1* A._F,JA\#X$K=6!>/_+W>O
PP0$Y)7HRT(+%2:I,YP?/N)%7BY3J<,<#=*N#JH_Q!Q0!L()]+0Q5-?LR^HMCMX1"
P3W/&@>#4CCS"B\1<@LWD6F1=\2B2^\8?V3=:R0_:=2=\$,[4N5"XJ<8NUY1]WYE#
P(PQWU.N-(Y=T,9WT62CYJ+-IL3;I >M\'E0LH-%*32O9Z</T*':,-F/HL.;[T,_H
P4^V':L-OJ7<CO+*RY<$\*0,"4 #GO%!JYFIQ?E0B*G "D<3RFUY;7+=22V?G NXF
P;A7B4(B0Z@)?Z2O" 8FB'T[],'7Z1<3-%$A]@4,<0CH?&LY72PXH?XV 1I.LTFRP
P:T8W+#*LR0 UWTN90IF.KPF2K6;8@IG]'#D+C;C#9RH!K%OGWW-%[6Q6C^("\4NY
P%^LRA>51B*UH=VU;]2O;8WS'1&.3NQXZ=]X9<YI_[P77, ]XAC8' ,^AT0!X!7TI
P(F'E-1G)%;:SESAKL)Q3?0Z2I/YISU4NX-72.X&*0LL31.(DP,ZH&0SS3S-5A-Q%
PIE1&+N2?R]!5WI#U\.LEAKO_)_>L7?(5KB6ZI6\2- H22VS8%E"EQ4D4*;*>P3]]
PU\R1_<"@44G/;X$3G[& P""ZW*BSO=1TT?QLB5W+B3CD#:$.BC29)ZS)1]0Q6[#7
P29ICK;IH+Q.(4Y.;5,3#T!&ZT2%GKT(-I +#O.^47HVXQP]L7B<$*1J2-/!IQACS
P\:$T,\VI5%(X7?"EAIT"2RZ8_CQULYF]QZ7[=^XT.\ZE?YDT'\OIR-0]!X.HYR8Y
PZ$V[JG!FL*$1BDKG#EPNO0"@4@"# ES\$B"L3G6X\/+5#&CCDZE)G4:C_IWPG8 -
P/RHI!2PZ1DK&$,'LJ%T4&Q+_)%JJ;ZO,2Y<L'-(TC.5?8;%U]P'NM"T[W7A>HV*6
P1\7GQE;C&8_7X\K23M&%BXKHGQ/%'0J0O24A;&])88+(IO#%F(F@A5 COG"M2%^=
PY^BJM9KK%)SPBEDQ'):FL5(T9!:XZ.P--A;M_JW^OL%-4LODT1F-2[U[9DPCWSWE
P4'5<ZW%8I'6EI^H[L]E'+E-!B5^*Q.E"VTGCPZB#]6H!;1$X;Q-1R5"1HSHD>E@]
PHU42$$DNN0]KJ/:< @:FI@Y>,*4/8N%"1Q?5"1)WVT(V$\-8$1IBDWIU[[H)BC<3
P6GH(#G%=JL&M^VP"DR2%TTLMY]0]HZVL_1)Q/M<N=Q<JW5-&#@]$!R:)N8^I%.ZW
P?YY&W HES$*XN26F7VK.PW^GKN3_.KBP73MJ0JXD;JB,QFH%&=5UB4KV&-3VJ=@+
P0[R<2R\\G8,7(-1D67]G9!WY=M<EH^!D?1]P^D#4Y,G[\-;Q"!'Q/?%[7)E'N;[J
P90 [3LDAC^G(PC):T&"!'BTXH?VY'Z0U^Q']E=N:6Z(^&W%%\1L&AS4+1&$.[S)I
P'=<";CS3D0S[E BUS:]$(,5K3W=MC)*]WRVMPS_=2&D&0^POBX?]S',W;ED29!NT
PNU=GC9$VJ4@I\R'E&P"*WCQ7_7XHS*T-U=GL^POUR%&UQ $!M2/)\1)M$X@?.R_A
P5;)S5.K=@\7XGZ'WQ>KJ.L3O((+5.1;-@L>0D(NX!OIU&+W#YX"^J]9YSG,#HQT;
PTFQF+3CTGLBW:_1<BCRM),G_KZ[[?-"PB_<:$1/^4$$OT9V&DY0?W7I;;V'7AE+-
P';W#LX\8DFH2)"IE)+H5RG'!/*.NZA]'7HU'CCCUJ2 ?12!7;Z>^Q?)2TPR70$3;
PQ=]2WZ&YAYH72<]+HG= L#!7AK?C0%_-H&%_@<E#4@IKUOTTU@R<@^FCHD_9(AI7
PGV:]N_^Y9@$'#I4&GZ%F*!%RG3P?W=&2S9ARL457^AZLIUIMBI6<X!84QS!8NWEK
P2F@Q']'I9)R^W//G%&VQVP_DH[W,8D!U.'J6+9Y#\#Q@"Q*)[A5!6ZKQB#*==L,5
P$J>HCK'XZ3T,F)W11?%<PW+4E[HCP;082TIGV+DK;=2WV'UTUG;&\\]B;E 'F?AD
POQP3QS.80,]*5QU#_PH$C7JP7Y;S=IRK1SF))PIK7+W8'R>K28I5S!M70U9$AH&R
P+)Y@,SW9L^20;>N=B>=6N4%&>3Z?!2B91ZR'#W/!O[NJJ ^=W4DM6@Y-<JO=O9+0
PB_P.0BO]FZ5:6M;/6O;#,Z^B&T)].-^YPHB!BX4M+K$>KI_-M,3JU_[6<HM((P)L
PAD]:92PBBN:D,71C ^SN-I\AC;QH6U\=;@39;ON%'E)/T1F^%OMYN_>",_*7W&"+
PGF8&3JU<[BKJ(8ZW$3/51W;MT0]-:US".NUB1K>JP0 R8 ;NKC/@T0Q!_[-<?MM$
PL8."%OA[ AFO;0F;;X- FB;JYG+-WPH<S0=]6HA:W>+YC=A1$T7>A*!M80M@PTXT
PH8_B H-*E05G7+";^'';4]F!8M]9[+RT:DC#NOUCZRE^6.*;FV4,K7;=5H+"N9XB
PN$"R"7H4LL-WY:J?[ZJ-SGXX+.]1KUGK'(Q&8A_$+S#[0(_EN2GW&?,DE$^?VE0A
P=H;/SI_'33,5E^PTT<>M 51"DUT391*V8!]U7F5Y:4!'JG=?0&3%B!LHD7PV"[8'
PYE:OV;'[PX*V-Z31S$76Z?T,W5Q,K;5B_<A7ID[:$UVZ?GJ\W>C>I /"/TK#)ITU
P4=R/^(^RQN B,..F\$['VXSL/,F:E2!=_4[[*XP;BWL?S> UT@=8+4DNUB_W&K5B
PWHPY/\[-6;6UHY]6!H^!7P,_,D&[G;%H>9I)#+H1=BFZG^3_GV15?H\V$G53,$_<
P"N%R*4/Q%KT;A(4UF^&$( 9NT8=!2$CZ><,EWO<C(\L<I+*S8M!+/-59<I<&),5E
P^ [Q&.>XJV*%2Q YE1S'_+Q89Y>PN*Q +E5I \;OVSUK@'3B%O+IDF!0^3IJ'Z1)
P35!,O1"J8\ZXWTR#)3\$)Y2[%IUA/E4EY-]@'N'A !N]Q<WU3[ZC(6\JL&,?OPDH
P>+T4$0*>WO/]7+W$Z=0^39\_-^Q2AH[:N/LTB P3^_3R*LM4)9XRVM$S>4$(XY=O
PXF%+G0+G+H8$W\._4D$A,&2K<[(U<,@C'3[I>A6&YS:P (^PK_1HNI(RX>!9=?IS
P&WNY=.UKIN6V>>3A!:!^Q9$I'TC+'X?&;%^<Y$>"U('QU;VHI](B:57<*8CX1+<+
PS9@E? :3%D!)N27;8QSS;_50'AG28U"*^9]!H0T&*;4C>MO8&P5-]69IX*Z2(-"B
P<N6KMFPNB'/Z-OF*#S7/NA;5XG^EF:I_/9BCZ@W0N[(-<R,RAV#1<:CN;^(>N3?P
P!RM11^AS(OXYK'&6AZR>JJY^3VVP7J[#BKL/UD:GEJ,"*]M(V>',)KL<NM[I/[N:
PGMHKY_7ET-=@LO;A9J$F2+2\"7!5JR<# \D3=*=;R%GRZ(-#6R%2#@V9A8IQ!V5G
P[/=3GJJ\I\/*_HRLSFLCXGH&UG(D8$<<5[Z6VD%5/FR6X9/5?'VUNR[AG+.6 *SP
PDX;(G$%-).GZ*+-R_-F>)H^4LSC<#'90X/TFOEP&B->Q#XJ!QCS< BU'GC7=2UO,
PT0:%>'Y>)[J'?OVZ=N<<_BH"%(8^C_BPA4"B+;?>7K]P08>Z;G_8G6]@>%(N1ONR
PK*W3F&&(\ =,/ML@S<V>) 9&RR=H,JB!O%X9!K3%3*CA)<HHZ%-L-:^@NLFUV5KH
P''5M2"V(JZZ8?E'U5;DPTE2-(Z-^NES"#O#DS9>;C1[A8_3@7D3!C#*QP#R6<O+V
P(%$V!6-!AQHK!I;0"?*6[34@*31<OK-B3GA!8EOA'1)L]0=NY"A"3QP:SK[U7%TT
P6Y^ZL21WSAYC$K'VMR=05'BL,#6-JZC(XM1J<1<,Q:$YP%OP<BO!"IRFU@#>[K%2
P6R6UV-?4V"E1^&.4%-F>&M96FU6DB'MS% Z<Z8ITO7DHC&Q&?6WC"B!-IJT+LYCT
P<%JMX]V[RSGON91,M @./H.;G*"&EH>X\U@0_ 8FS[@LS;*0@VX'65BL#,G4<IU_
P%.KCYU/$S12ATP0.C8>J[(%\'3*<Q,:N1U_^6)8"CXSD1?!R;;TH*0/['EHALN*H
P6=;)7$Y@N4[[*:"R2/P%H^]QNBMO^KD5:K/0!'+GYC>]E3\W^<^)NO*+&:X1FBM$
P4Y>2J'<:_H=1?']=CBY#JZ/J:<_<_TCOK(!(UEF>VQ8H/+(U%M N2V^52-U=K5,T
PPX@(H+FQX^V(EAG& A&BQ@+\*:QB)"5I0WN,KYY^PNF$K.(44H+$_QCQJE+=HX5%
PP,+63;;B>TF:0WK'%J3V@SW7JOCE?=0\J-?W7>FX/PAF,1.Z1N"Y:8^_D81(8EWN
PMN;?N6V]Z3W@4/Q'.4 2TI=MF)9U20G8<81 U#-CE.D'E(+N!QZ$.IQ'V&2!*P,\
PLU]9[KSER'D$V7XXTLMKX),$_-=XS0; 845#<!'F(BMN5;>&"E\P1V3QGCV+Q[5,
P<.G$ 8XS+1FRU!Z*@@UG8NW@+M!U%QF&[E@30NSBF.$F=SH!K1M2\2]4"=0 K "(
P.#SI$BD>?Z97-<&<MWXQY%41#X_<UI<YFF-V<I<W_!6#>;&Z_ ?D1/EJY+XEJ1I-
P%%E'4_;HKR8:2[=6F5-*,S)),;*SJ."2R#-Y9J2PB0E[4WW.0MSJY^+Z+1'4^_X)
PHKGE\M8>O0"@+G^;X?=&08B,IGOJ, =!.9Y2/^V]9MO;F"UMR<"TLBF[C;?A-J9D
PW4JVX'\UBB)[SEXOPRS5TU$&-H*/\V\%K9KVM%)P+TR.CT?Y]'?0D&_C_0S@5R3S
P[E\R/$J-?]::%7, @:)NL?"%<$#A?GQ7]6V5QQ( K#D"QZ<O.8?K&QO0\HY.5*QE
PFWI/S6M79P<MP5L[<YKNJ^_WH7-8]'6RP+G9;S'5K;\K<%RCIFZ0%1V9< [I$802
P%XTFXH:'N+6;&^@#MZ7]<.ZMW<0DM'"ET!K'>TF+67N*OY(L.=8(+9A +@1,A3,N
P5D;&O;8G4=;%Y6!7?#L#E@]FWPQS],GCE8$H-@2Y_L[:U>1(MKRE;+1NB6YG5BYL
PQ4ZZ+;0M^Z?)H2AJA)\#RB:1EY!0CVW^[?N+#5=O90L_V$#R6,R%VDE/;[E_=!"=
P!KQVBSV3C']G#$"8&#>\D#@HB1OF-@++]Z?>'A*Y,+A!,3T38)&[B]!#]((_[ L7
PU-CBP4L@F#28/9M57 K!XZ@6+-K#:Q=B5M1WU(1-V(?(L8-0&)9$&NVQ67<SDY*U
P%8WZ]CXT#[G:(&(:/_IR1CQ[]L]A&C_3O-PBM[/-FQV(1U+#77H7:102)'I_UNGT
PJ;8J:2X!KZ(+1?<^YT)P<@BAPL?3R2[6("#EQ>FK:G.> 8K7L=1BZK^Z<] V:-SJ
P?O!P/O;CU:MHOP 4'.:2-V_^WOHSO*<L<W@/1EPJ$=8+B6^19B@GI YMI'#>]7!W
PGYT-2>,@R5J^>#VEEUS^<H'PB5BO?1<V!_'1O ]2W7'R92JX2>+I=H>N&F-.0Y4;
P@JF6C>HPWK_7!!-9DJYW$N]1%#L]3)*;V*<PB)D0M)OANO[AF^-,Y$S"=+#)F@JG
PMAWUYT?$^@6D5N5O@#1#=M8]CW^S5%)0$*$J#BG-PKD!/=?&UO*[&\3Y[N^R:I43
PDWX=0$R4-,HK\M>P7!.A8^OZE,:LJ%212\$OX(5H"$IR@A*?[K]KU12.-S?7PB_6
P#=CP^89TB"SF.8P/RP='V ?K ^#(S/N!U!I^EO '=J+5,HI18FH68+ I_9NDDI) 
P@HR$@(J"@AOH#R(6AQS)CD+Y6437 IG% MPP1+\*J_IH#"MC+,<.AO*SS1X]'X>>
P5YXU2WKQQ_0_6\!]+EGBVUPVN@9,5"DH79TPZ]<;8*+(R,[O(>FY"ZN#B-4_7-X$
P6?EPE2!#14XX)J%NQ>,DH!AP%QXTP%EC1.WO68A$PPGOORQL>ZI'=-H@(J1#)ETR
PI?W^7)+^Q7=J+5]G[DXK;:RVUA$I)Y1CS*L]T%!H)"UB^J2-PZ84H$!?:U:GV#C:
P=OPWKS$:F&NEC8B>I,)C4 2Z7E,=D8W6T4BB8F\Y;E1#$-[BI+3$L1.%%#Z-IFT&
P-8K4_2#]+&>[%JN^ZGIV0YZP_E)Z/V^Y16S!62_)@WFS'%3NL^"+M%+C>;E&0[28
P)GSOLD#^*OX^^9&VM==.KIKJ5UVYQ<Q[!NA' TS50AV:(&5_9)QVKD[_.XXZ0P3;
P1*KNC)]:!92&<=T[],_C H%N;_B',W6Y#)FN#J@#"2TO 5!.%D-T;[6D'R/@\GL#
P0T1#T;(W6NF[;1TWIRC4?B2"A[8ALV^!UWJLHY@A^=)$D;U'#%U.B$:H>$1/ 3U]
PS*75>LRY\$S.Y+<AFP&6D7Q2(,G*Q^^T*K][T6NC0*YWZZ0O_^+76CE\:: <3E;P
P)_*T'#I.V''S$#XHS@[>A)_\"/3/VB'5!>B>-L0FAJCZ$.>5!P!+ND7>EB6;.N,Q
P&8EQSD*F2XXWX6VI$Y;PNZWV=AKSDF<=$\:$\TQ>)=/9[]/"PP]?902AX(,#,2KO
P8-Z]/\1A"$>C+M+#!K]EPU%%80'RNDP;^OFC"B[^2%=@H_7*SJ]Z,D,?QZUM#D%_
P2<&BOJM4G-B$(U\,C;V\P\X";TDK7F&6']P:?WQ<HQH:6U :8ZONC2.MLAGM;W&X
P-[1B(Q6ER0$]I=HUO&,0PO)QUG54692WN+:MF2S \5#PWW9QTW!5H:\06\0QQ(E'
P&R[Z(V7&+@04P,#\TE+"&DJ+.#5L]3%J0M$0%PH]42>C->6TF;=\R+G7QG=K#BV!
P&B3L]L%LW"".EU=G9>GU4VYIUX1&:"%#9:4TDBLB^>.I5MP01$#4$L2J&HD_DG;L
PK=R,8-".\>I*XN2A'@Z "JA;ERJ/*U.C?0.RT%0D9[PR*V,$ERA['MK:-^>[#.;%
PTJ@QXH), ND:%O M+"S.4,M!T:DM>#O#^59:AM7.%YO:SK(!$B%0&BG95)_M&GD$
PPGU,<C2LJ90Y\GH1=,SYZ4AR9QMJV*]) TJ1E8_E@O% >8R7T,.BRN@%RKK3U55$
PT7X-YF?D87SD:,D%6ZI=M?+U5OEQ11SL6$6@!F/R![TS;*(-[V8;RO0,& R;__J@
P'[#')APY*H$/47P29I^.!B<.C^\>(7YJ>9DG0KPW7?91'>CNNX'.*(H+9T #S_%B
PV Z#:L-9$_:./CGK/:1J*4-60O.Z)Q&4]\W>TB?VGU*4*&=,#E4I"SGSK>VTV"H@
P(2,;0_OJZ'(R%-_YAA] )U LM 4->H[V,F)?)58<AC$$BK,!'HWNG"?I%-&EK5,0
P+C9^H;JA!%4=]JD^.@E7A@1!A19 4SY7W/HA8T#A'W48"PF+_FCV[NLXC&OH1;P;
P#9B@?5K!U)NLXA_2<1\_HE%G%REY((, T>1P/+$5?@$"9'>;>OT)LT/$(VR116!O
PXY$CGN?$R(3D1*X3E<%4V F#IYRP<U6,L#&FNB7.H:I$@L&9T(1X25N.3]ZN2-HD
P29N! M8+AZIJHH P(UK52>E2?O.K4]OW+=WA9N[1Y\X[CU#!K5.[\([HG";A)EK'
P+]>=&31AJOY2>06!:Y_-(4T7!:8]]8FR+0K>;<HAC5Q8F0'6I:R?U#.(OB8I,3&0
PY:-K430T;\]_)!*+MO7ABXR'VOE\K71O8[P>:MM3+Y*K1C43*?T_6<'#'*I*&WSP
P@D>;T-YZ(&-@_L;>J=,?#6AK1H";.VS8%..R$O(@K% J",VS;0@ ',V[!_461<ZB
P+07H*"$?M>.+FH@PB:U9=VC?:]F-HG[/>[UEB"95HHD0=$>^?TM&W:^XS[^<I^9D
P_"O)5IH$"8;ZT RSMY</'A&W23WI^@2<ZI6=0W7::E6#1PUN\;)=#>->QZEDW9>L
PG?MR]UB;AIL$81T39(.5>2;\,9B3-X=.=$E2-"&X(=>__Q)[@CCVT/Y5D/U?2PVC
P8D)@S\]JO:WB)H+&MY];L%"YU*;<@SRO069C,8<006V9%BE@DL]VU.[>\6Q#@UUY
PFDO\X2;-((W'!$E'.RO+'$C(*R,/ KF#5$TP?F6/3SA":(A_28&[/$MA<!N6*@YU
P$5:5KN7'(3OE^%<CMHK7PYVI:8Y-6T,1* VZA-RGV[),3/;<T^4*98$>H,8C8; B
PT*M=455F*\  R;4S4N)N?S#_=["\M\'D?Z&XD"\T;^,NT5_)>:".[B6 Y$,WGAJO
PW#?E%?S*K*JRP!_;Y+[4I[^0$PH':>&QD[H4R0Y$!V3*!MD(D49+!>="%4#_-OAF
P1^7_H)C[EQZT:'444JB;#*NZ_ Y;@3=KB-QM!N-MX;8;&_8VH;?.E+550B_+[(NL
P,/[DR H/:K"V1CX;)Z5UBB?^6]3Q_\O3['PT##5M-DVV>QX8WL*2BN.4_>A>:L?\
PRSN5(#=?1,T$]!@=?/6]"S @7+Q_)*7_VG0&#.MI670)D79 =06)U(4P:G&<B2SH
P2U>$%OWX'6N[FV[(ZIO5"5S@J#5I(K;*Y']$U"GR4KA\T(1(C;_UPN*#4T?84(/_
P.N? $'S6B\I9TP$C0OT^]'(>Y=BWN==^*.S)-D6U8=0$,]_&SE8CP4D]L9BS9G=D
P5[3GWG*0XS1<\]!CCT:L  J.R&0FE#TIN.HJ*+MNQ!(*$&^VA?3<Q>_AF8)D\I+8
PI@L+U=C,$R"JAL@KKS9_RWK%RKN$F_JNJNRG2\\OLJT0KLTQ4>-]:\Q20^TF7FF8
P&U)V<KY?4J$O.CI-_D<^GEF*H866"FN5%&_S&AA*@675O9NK*2@0.OJ("15YN2PV
P_UO@+"5 @G>I!'&66$]NMI<QTIN$IF_),8UORA</HMN\UCG($/+OO798Y.:&EAF?
P%-=DE)N:^12R^/9M;A@9*6*I$7>H]3S% %I@E)%!LZ&Z-2)>/H_-A846P8XNN&J7
PO9!J6LA6';J7EP0+XE7C_,$G6>(D::\3E*SQ[WG?H.#H#N!UTK?.< UL/[DKS9M?
P=AA#8@W!0%>-&ZPPE^-JN8F8@-VN55U$;C)LXOU%RB#L4M]! I&^P0W,%4="*R71
PXJGR&;W#U%D#Q+/[N3Q@:1EK).E-NY??G+(C//U/N9ZJ@*ENP17&7$1T\XJQSB#(
PNF1C&[:VL7_SP,;= #-<@&%*8&B;NK!0-768#F+4L9U#.2$@J-IVZ5%R;MYC!\!<
P>' Y5B!QMM&]$SH2XB(ES$A+H1;4X9I>H7I%.$RHE;X'4LIPL1,,IQPJ/)TQ4>Y.
PE^\U,/#R][2<3_K&]96>O$GD;YT,E[>:=KN1L !]C0BY)!H(*#W!H<)^_)$ 5MTG
P @#RD)F])[=[DK&'&E5A_V=2JL>C-U!=:Y'2@'35Y7&-A)O"//R*YOFSJ*2V4S!-
PJ),GS:'GYX)L$!G4]ET<B':Q;C"=.H-H640I%<0#^!8$BV56Z24G?%)#,>I1NH_N
P5=B+/):4(9ZX_]?WH8&X"&*;1XAG9TX4^+J;9L-U5&TTTLQ\GH])H0(^X/"NXPZ 
P6%:!62KSCO"!/UDO2EFN21UYY*^O[)Z&Q(_\@>,C%'(W.GQHW\$ "5 F(R"U8?UZ
P C8^9^SE'?$/.3MCB0=[+V0?SZB"%@6()Y&-#CRN_?-G,ZRO9M<;<P:K!G;@>#&&
PRCS)[S1XIF-R87KJV%^59[:BCM" $,= 8%0IC4G%.;#FO*UAI#%F72:J^2>W?9RI
PZY\T7S?!U]O-9Z<JO_.3>,CC2([R<KPD\"UFUN^@4B,Q1%+AW%L8E4L>C$V=3OD$
PX*37U51X529MC^X$ZYTN?.#=D<D=R;/*\0B5N*?OI#6A:M!X0B-S27NGE4LX'684
PKUE#3=%R\;Q56(*@IE=<VK[?.(%4ZUN$&)LZ%6?(6.4N-8A.3.4"0XVN,4 1%;!6
PN#,15?\"4OI[>[)Q0YJ<^# NVN8?X<]Z2U1J+Y:,%.O=;'"KQQL(BG8:<JU#&)JB
PI3TG]PRE9GZCJC*%WC B3D<423NFBMI5,@1#>O3L/!=[/53N^\#,0=25:OKWBL[E
PFN[?0)HI\JY:APF.TE_\&)1.T1JNCQ$CL;=3IK;7>='GQ'VX+=X13*XIFV)[P_4\
P6RFJSOTN 7L#8;FJ0SWU:NM\##\6.MD3++5QA$CEW?&/&68X[V,Q*=;]A:+&]EX!
P 0HO?^O(*M/>$_<]/?*A@\1 F6$L>3#:%=R7FSKADO1Z(M4$/UM*(G$[<Y0H\5JI
PP:$K+5;05C-Y,#C,E7\"6\]ENMH\JI 8R5*:9F:B!L+<"+Q.7RQSG  \&W.AW51C
P?#7ZE P__[^,TFSJG^.WA.35 "OLGL/&3NKB.1"*P6U2T^TH[0*4E;J+1%UDO#6Z
P4J(3<>NBH\-)\5EGN_Q(8-XV89OUR9H#=L8O=^J> CW_!$4A$D(U#D.&[+<*?WB/
P,LXI"!8:Y9TO5M%/6*#6(0SHZT\J:USX^.6 I',NG_M_W2F%B=.02G'W(XV?"]E3
P*]2XJ/GT^\=%?Y?+O3,ZJ"ZJHV>S.,$WE:H>CM**TJ&5'<$'5 4GR;&!)$["A)LY
PR!4 /=BD>7[7N+G2U6:;B)O:_9D7<2^'_,IGD!!.^)SXT!AO<G759FIPXL]5H2D;
P>H8H!!%# \(:=,"D='?M0?48E9I?+N<55;'JT3,]+3X%^Y,J]]W"L%D4H/<,(L)(
P+* 7,DU6>7D,SQ(OJDVDO\+ RLF7>[=H<8O,F9MAF!.0?&"PSU#UO!.YBH[]2=]-
PEAD;Y:BD\C0G\]4LL72AWB!$:#H&D6OJ<<HN=;_B%9#V8^%Y; )]I%XFD5EMC)56
PG:I4^LWY;FW/#96-9XFD(I5?HT-5:"J5#4CZXFMV78Y%,=<%:%5K/8SC;+Q/(/)0
PWN]R&*^)I"22:=B(=XP'E:Y9Q^]PT[W4G]7@&/0IS)T#FGC>;+_.QM9SQ2=N0I=8
P2.EM@O]K0&N!TG\,0-PT98G%DV47$#7?V(]XB)_!O7A%;55*%Y4+GST5ZXQ^)5^R
P00;S0_L>B0Y]Q+.2%M@R2SWBV*>!^00G42!TR%,)[ANPJV\3GV@KY%"4O@R:O+ZS
P3Y M^BD7("L<../;($&XNKO<[Q/_NU_!AN$05*G]<,).1@#1_("9+7UUZ\[F)N]=
P4D*60;M4)8Q#Y:4@L#*"P+NFX'7CR?J"TY[;"#RV\WT(%"R*(D][3<:KC #SAL<$
P>P8MN'.%67SD !]BH(S-<WRAP=MG$MGTU_=^F\$;I;S>^(HT$:+7U:"%',>J+<P.
P.0@'."R9D93-=SW.D]L<,4X.IK@0"D<K,-.F/GI+=*\)]OXR/*K!.!A"!) R)>0<
PK>*9Y0,3</6]^C]4"1Q L!/-D987T=[PPU-44KOYD2MHZ151@*"P)O7LU=2\Q%W$
P;/.65+;5C7/KTNM^$'UN=NW0:4_QZ.]"66AY=M?P$?QTP_IBDS+WDF;,?B<TK0.9
P'LF=H%).WM=;K=[6(4PD@71JCIPHD4"61!_,[52T]^IAR-H*4- CO7N;Q92A&FS4
P@4]HBZ2&(5IZN9;5CTL=1XDV9.W61-7A/D.=+:\4<>;_3<,-BYN._68P@H "VS^N
PDY$1^"CV"G).BB@AG4&:V_J"3+K!BSQ"H7/^3(M)6@C\U;_YO.93&0:10X:;47%T
P)\8'*&(V(C)G." Z>8@JPFDV($[HK9RR+J$S\;?9*?(JBJ/,@82!A5/[/M]P^MZ$
PZ+#?BFL')SN+7V>*7FK!<CYBJ,->Y@=^.>\,Y[V27CEP&=2R_R1;9'5FM1Z7V&$9
PS@2&/Y\2-7$OW 3R58=DW9),T83NW&  !KP>CY<PYU40H]%27UQRX]P(0\>9O%.+
P+<CYC-PZNI57H1C>.YC.]Q"J:^\]+?15ZH\R*%5D9@&9M@3[K.P!Z!9Q3KK2EAI"
PGJ.LK;XJYJ9!WY['$V&)^;3":XCL3'V;JRB.7N>R%@V+<=\(637.W"D&M1-',=I#
PSK'^EM&V>5F Y;<)_Y3IM$-3T+(C>'V=.;)E<B /.SG/+&X31&W;7!&Y]V]?-])!
P=TE]H:Z.^8*F?D1@D@^:RW/BI3]VFRYZMB!BT9[P"M P4ZZ1/6*7BJ,N&EYS5%13
P]VS;_@K^N[A-B<:QS 0\WG= IG.P-DQ^FL?)(3Q:\Y0\W0E%1K_W*SB8*Z'Q1L(J
PYA3\G[@B7Q1"R#WHUT-+,HVV#;5G\486:<Q>-TO@FX>5'FR]>4NJ0<GO+@.*BC"(
P>16K(&$,/UZ_O8!V&33;<27V\[B T"OG T[M[M?RJZ+@-"Y6S-=PHZUA7,$4C"I^
P EZ0Q3Y;4KQ *A*65C$FI^6X=^LE2$ )L>>;LA)UI6O34\A&IX0*H/PM^45WQ5>>
P("W@Q,@W0KC3,^%\UHGR+M6*4=V*4_J5.FR)JLVD %CRB"2/@^'5XU+4O_GW''/>
PT88/<-+R&\//#T^/(H2&:X;9Q@7_&%KH#O-<'.^\:@I6YA'^E14!\N)+J-.2B=I>
P=+R10;4W6D4T@C.^,9E1CU7B[V2Z,2YGY8=#J=D[+@[3<#0_FLQ1F<&8MC&\=@EP
P_K3#T(KZK\&7?\E,^(C#6CUYXJ$8:_# G7(7P5U?;=%:/HAK$#:L\VX4+C@<^=7@
PVZ-&:K]?/ZX#V^8\K+;((/T1?D6 %^7PVOIU&K3]#,OI_0?=J*HY&B5SF$1(PEB!
PG$0 HYK]$XV2=O2 DRT?LQ\YZJ6*[@G)5;0HQ2U[K*H[:0G/S8-W"(FAY/"AS_HX
PZR"=8R^AX%Y,@+SLWN').GN[%ZQ2W;\T.&OJ&N#[A'VA R)WV<\@=",K]@7R/I5L
P3[OZ9*UM-?5I>G #W<E)A,Y]$_.,-XMW' UGD%P<SQL ?RZQ+/R%,SUPA'1UA9M"
P(I31VD&RE)1Q231K^([@?(+]$QX[??MZT+Z$RK$QE949(Y"5X87MD]J[1KLS^XUA
P-TM$2#<RVX8%2M*]+=RJX ,I'K?6"A<'LFR;L!JOP9VA']#$Y05E>Y<;(6*X%#M8
P%[-<OT3<9$A6U;>(A2?ZH\L<3NV-:8?D(7OB#-.Z241,Z'$H-*&_5=)T9-H!\B1=
P!H(;!>/S;]6.3*ZJ*+P;_^LF:)0;!P2N,VO$IA"(G]W;)FU?8>#4>?X3R>DE+7'M
PV8+<NPW'73/75ZC%T60X$@'@O2^GV-L@\T>4M9F0*U(FO==ER C\-Y.YQ/,D)S3%
PX-$!/*'0V3^I+AX.P\TD=6,O#A!L@YL?#A]I$J=VYPUA+)0JQ:X.#^ZFG1Y/3P%;
P"O3G/I)T'L?55[FDV)$\4BV?$D4"WJT8U/?1RWK)4RG7#E%=:!#3R*K"270K3\OH
P\E@ S89+>V+-4[T/*N$84\<>U),1&*A=Z['?U;HFV58M2^$'42T3Z!_E3A6HMZU<
P14X5L&DE (B\G]R>ATB"R"^J2"#=OQX&6-1Q9G7>:XA*I>J3+O$ 80YQNQ09(6>O
PTW*/U%%.#SD9V\5.E(:RMZW6&&H8>T0:=^)I2L.V([>8^IV<[2 !G$@GBQ8B)(I4
PT_?RR^^B^:AM-B!J>'P94R*4%E!*PNX%:A1-RK!H78KD%Y76[F9.J/T[_EXH1C4T
PJ9/"?RVD;UXZ@PH$XNRC8&&]#!CN_#:VW%)C_*>9KFUKN*/ET6CO_MN&LW#4!_4_
P(T3KW>C_(&W+0H"&5'0H<% $Y)I+TY9*_K(C#\@MK[)Y;^LAIG?I5VZ3!CTL:7;X
PP#O;=DL6J6>>[TPU'@# W:/MX9U>--,PO'H&D65,ZC6>>BV0!(KQ>D%*R<@LL 26
PJ2GV0=>F=  TU5+[N#U] (>H52-_>'=^6X'+?&Z/^3;;$,UG W&*K@-!;<W6&6/!
P.L1#)0D;#I=U]OL6$[1"BN7# MJ1$OP]J4D(NNCAW)^_:^W,\VP41<"S1V&#8(?1
P@35;3T9Q65+(*!PF\Z:B3\6]>4XNO@Q&%L.)Z3NM=HME3*Q(3B[C'<R6M:O:T;N@
P3>_X<$JOKLZPI;*$_1TVDPI85;RGS5X.#ES5K*G^WX#<>M!TKVQ1S><<O?M-69B=
P]?E+6VX./-.G(D%5V67&<Z.N""\2H0SVF2BAZKA^&=S%[)QX,/1RAL.ESBT<77W!
PW>#14>1BA:G,;XF;T8K1.H1W>)['G_'3^/T0><.-W_A$L!D%66_5K@+L9U3;X&1"
P2#H?"TZK();,<XR@WK!H:V\=,"Q8@?[X?<>$H]F@19C^]/9P1C@94WSM\34-E634
P2;XO?LUR2ASNC8]#[I"C%H9MN]+)7$P^0+OZ1X7?%]S3 _:DM7*;341C+EO&<GMV
PO]Q' XHGUJ97+" 91<-,B"G/R+++;W(RL''$!N>1_R9J\>9ZQIR&'>!J,O=YTS<?
P+4=TA GOR!:R_[S*I4XXT6]\L[H R3IEIIDE Y\W-#XYIR;/)#:A*)V G9WBV>2Y
P^Z#"0!'=%-[,KA(G7$AX>5HIV\9+$=9@JK,LF^):5JGDTR\*2V/D6GSI5;G39M>/
PI_/8.] [PG?_]QK+4O//]DK#@Q&IGVKC"T1+?IR#IEL+13(N/\1MMNI;L=AA+I."
P(]HD$EMPK7?^O\WE%XG\]!-TQ607Y"I;43*7(2]"U$?)[FPE-I?8^=!W>^V@@+:0
PL^#%0@H7Y3N02SQ+#FRHNF)6]I$>:.!#J1,@W-,WJ,8E)G_9W?9JJ;L>:A]49U7M
P7EL2W++2V[,4:N/ XG13'E4!1MP=2R3)Q[/1BZ>=)>,3"JZQ??5]WKJ.GB%TRCA 
P1TJK$"Q24J*:KS2X<=B;HL%U@<[P4P)S!Z*^7#C1?U%:PKCR,3.G,YA[+HW_YQ[%
P#P(469:;#!%#6&#4M7^-6&12Z=CY%[F!*9=<@UQ?20E#K*7$'ANC3RYO7/1H,'=4
P(NU-\M7Y1S'4PFO T?@MSAY7#8UFG@VF#B1%3@/XOF1;.E%TCOVM?-(04+Q'[845
P(<HXOG9=YRO92VD,*5?#E:W^DE2FHJJ0D2F_5KAD& 3"$]PT38OOE'.S]'C:2<UH
P;[%HI1]O-#B<(-FDE>YA63JT&%N&#+)18TT"8_[;Q,\H=/L3$E,P[&JZR*M=-?H:
PYJ1%HN%#C@>HPXC\%B+;6MHRPD65F-T&J&*+#$&8LE6>TA'#$.2>:&_ (3#NR0*]
PLBJ$6:)^ED!=$FS[)$ZQV-+6W=N]:Q"-ZJTII\4T.!AE^.7%POD? H:DF=/Q[8(#
P>8<--&J?RM2/:'ZX5FZ.WB^%=<O4QB]A:G[J.V&0(OS1J9DL(/-=WJS[D89FA%.D
P<^^2L/>=8C3H%IV&<=OE?HPW0[5T74Z6?IO#!<+KRH"KMV2UR?HIF=!8/?0'CF-F
P"ZYNL9$]AU]V#UX2-)5_L2%L-:5%H;'.M'D9<"'%R-8J8V_2\>$DS^"+99[-0_<U
P#.B4= 8<C\ORA\X=5^ >S$5D^VEZ<QN^.AE-%!25A6AKP"8X6AZ!;ZM:7?\?<$Y6
PY.[NB1FOQT;3LE6.J0%'M=F$NLYG)B4 !163S%=HU32ZTG2@S,BU784$+((A\G:0
PJI(,IFG'2R/!G-.>YD)HLUXKL<!\=[,V[LGEX'=N9'[2^)J**N3N_-JK!Y#5'9]F
PS2%ADR+\QRJI]@?(<MQUS;-\UU()#$=9C&2L)'I5004F*I&6<M 5G%96=O+PJX+=
P-:+_^ ^E)E]W,#NY$W% 57(LEB6[S#B!];'Z"^$4MCYU?L@I*1D $T5 ^X:#U+0)
P(&!#S_"Z!!JC)Z\2ZAA1;V&* H]\=3V32S\T<<)#FC1,2HJ7T7"Z('HH3LD;39KK
PG-BQ@?%X2#6GL:;RZ N@#;,7'[WMA\;!Z(>=E'$+U:'7W20I!A)5']W'L9;U1B$U
PCS[T-)\DWV41>UC@G1?\YL[C#]A&-V-B+LA7&P"?;ID K_S@.N,FILP>1W;L&IJ7
POQ!M#@\S[GV*+XH<!&\2WCOR[3> 2Z48PMJJ(VQFY P+7BE7VZR/+.2=E4=;.B(:
P[7?*6J#__F@N;?:@S2'*#MF94!Y?^H4R1=&:SYKXQ,,^3=:&HX"?.GI>GH/W6RD<
P@!5!G..AN8*5 OY._9(?+VPBB1R?EN^BP3W+2L"8_CBWB,>;.^M<(;'E*@C_/:Q\
PPWB<1"XI,TDW2IF"'8*8+OR#-USDGC/V;OL.&%^3>BC3K)65U:JY%T\D<G-K0>)[
P4<[W;&OOS'EZ-OG ?R1#6>#Z%.+1)<X*_:K+RBW-'XW!' 4;:8$YNDQ8 ;%7CVE0
P KUG-^#$,QZIU LIZ0SPO^2,K[.,!GP'$/F&6@#-\2YP+ \2=6-:3=0L.<%NB<4 
PBE;@6>,R#.TKS3R>,2&OF-2J_('N7=)@O_WXA0*;F*EJ?S T+S'KOVA .)^+6$,I
P<>S)E^-BP_G#[FQ@(Z1=E27AHQ(#C^CIFP<J$O@HY+^X#^&\/N)C(5FTW]6BYQ3:
PM>,9["KBW;4M/8US.^)CIE)/M9XV4 $I7\H*I(([0_70X[C29\"0':/_>H0RV_MX
P*'P;NFTX'/GFVCF,#MK'EYCL)QF6K70>2&_[?QI=6J\1&]7V 'XS:QZ+-PQ/41WX
PF-N_> ';F<NR&J/X)>>V,JG>DQE#.\_K-9]1MKC@"4%+?88Z1OP5S/<04*4;P]&'
P7:P2T+5_E22-NM"Q!]Y4]!Q#L36V9%6<S-C=@9+>),$3]5=>+>N>PA&FTH6S0XF8
PK07Y=N+N8V.3UW-AF@0 SV^M(*+1:>;U76!%7VLS7V)KA<,H;\H<"\KS;G0A2JX(
P.*^:!/7*F=;@^&8RP_$:9+$M65/^Q,WK4+*J7,DG:&19>1W"@MO$H!RW%*<S.UXY
P4P/AW(',H"Z/^?I< .R>C686Z/<[%@U8^()BE&M^KQW&:VH,I<,%6.(G8JE[K*8 
P0])VA,!'S+9R+%S)F/'/P)2N%+LU['HN39ICE?A##./B)*4D7!*.[((ZW5T\-*^$
P<D,2NH?N*4?9>;P'[._>.HBDD<+M<E$UPM00"HP Y0&UZ^Y9SBL>]YFJ+5X+V03^
P_^0^SL\?R"TW4HG?+@+;2LN[96QH=GI#"-YBBF69W SYXKK^8K(#5S'.U3%YTJ'D
PZ>7V>)PRJ%A4@_&*)J/+:!-61"]MJ6U[^[9OC<&U]XH)5MBTF"W!= C W^O#-V>M
P)C1U!7VKN5XW424SGJ5%WJ8VJ(-BJL>A/N7\Z%.L,MG=\'Z@I<*EJ1LU06>69E% 
P^IP,'AHLI-<"S\T!++T=Y".DSX!GL9J!PX0:7X:IRUO*#Z\]I^TF:# DP/E*!<V?
P$YG<B4@GA\@R32-,\.MAQ# J+?!V*?8;$QW;"$DAY,2],UP5/JM7"8E0]"GGI>!O
P-XQ%!8TW!.XWV4A]"UVO:B?H.'#=H&(P"+*(\E3-PZ(6IED9FL0%_052KYI!XQ/4
P5*;'+MI-BCA]/):1?KD\]O>8^J$'T++9R-$;FATT4L9,+,U]"1-U,HNS'\-08/\$
PL DL#ZF9WC:_PP$G7^(.4+B8PGZ4B'=F;$A=J&@@R$69OXJIHQY<\LRM$N=E][P"
P-!>#2-UB,@.$<Z49%N=H\%AA3C-QC+[CAA@N1E!I: -T2&!Q=KU[9)WCI#"/)2=H
P0>9[:'(==1[D?UW]@O"YPTJEK)BX!D>C.>RC1-\X)EZE5FTKNPM5BBCT(P O(DCC
PE 08,[D?H!,-5[7 ACCT([+78V57U(YYCOG:4'SA22^'B*I(J.LE)O[BG*6ZE$@9
PO2N2/'5HL2-EN)L@JZLXWJ!X+T&\3WA'&++/-R$<M>7[=W10B)3EBUMI'R$I4-X9
PTL:^G@_%2%0M4MQ7HETKF\"6BKG2/ .-0Z6ZID6.J9W2"REX8CJ? IR;^K*EU3@F
P@.&+2O;017NG0V5YTGNQ=Q/T(7--@Z'7OZ4ZF)N6O+E8$APAXMK>QF +CUF=UN>8
P PIN#+SMO4''$*;DH)0)?EM7;%;T/:I@'&)=79\4F^R\G9C!GD9ZEQ0H5&E8F=$2
P?--[_0[V.4=79?1?7QJ3A]'WBM-$@;JR@JV@C%*RCVZ,(M7+M9!4WF@?F+T<.MYE
PCW?!8X7\@[O>G(_>.?O6"T2\0D>LMOS!3QNPVM1E6'L_7 H68"M[?898=XF(]DC\
PF_FR&2D/ NEMQPO?AVQ9)K2J[=C"K"8K.MN_DG?CD$ M=.3WOP5<7R;.$Z"\+5=4
P?Y-E9N*J&[H\MX"0-U:;!'158)-E6SJPVQ_IWLFN2JD UV1GK%Z@QJ'\4IT*/O6W
P7^?'9LF\(-UY]5C]/N%0@^A1B&M<E=$E\W4(%IBD@><]2:!"EE65%64/Q'Z^<6$G
P"3F*QD5.]K'?'<"@)\ZH/&OY.7;TQ+7ZS;Q!APQWA^;X<.%$1";@6Q("!"E%AU9G
PT#J_N)J7Y<=AN&13P48C2 (DX;NK7*L%&DZ(5 S@WF:&6JVD*P 83RR&2_[S"VNF
PJ*V#6GDVJCXD1R0V)AWL)N2>Z7.QI&':4+04HUZ2^C+7<<P1"NM)D@R 05Z(^S-8
P#0MCR-OGM01^2TGHF3%O"07DB:1Z7CWU8EU<VB+6Q>$I37#5(:YMFCX[M@Q@&_/@
P>,VYRAIJ+SCLOBF[.I6\3]'%S.# I]L)'=/<?6@OP )^7X%B]:C6D_/3_K7"+0\:
P2TX"DP6$/5DJ.)Z\!#;%IPRM%=OWA\<-M(7[3R#"*WDYM/"<=S#=I[)"F$;O%CDE
PIAKII"XOCRL=.JQ#WX9@YV;'KD(IQC7)Q9E?@]#H<P+8_Q,FSAI9,"[&2%C;[$$V
PX;X3S9LO\=@&O7"[1ZH]N-R2I)6LD#_?D+.E?X6KXNFU>F,9.; ;31AL"YH*9"1O
P+0]MD/XFW1ZFNL2N*#B72+(]'#R5 2"(D+2F384,FH*A@W1M6Z]?-&@!/F[6A&K3
P)G#<?-K-4ZKN(=']E2S?'D+"1$7*LRKHC*6\[V2>#BJJ7AI9O7QP486/&,(2\Q>5
PX3O<:@&0M2%_$"59GAL6,QQ*ZC."3<!NMU @Y]KHWGU6;Q5X1,CQU_$-=P#_GQJD
PXQV3.6.8III&<M 1%SM=PT60S(A+:Q3%,J!JI,H(^N3R(.&1TJW7'PK@1@TH/'=<
PWXV0/,#T2EUN#)_[;BQ+..\;\)7!QSJLS__7=: 7\EZ^,7,=;% 6D7CGH%&__0*6
P1FR$" I#&A=Q<FZ-YU[_>\E=5"2XPL$;Z=<);A0%F,DH!^R>."M'FY3N_SPX'XGB
P R!*WK3T=-L:R=RK83[&W EU.CV,W5BGH9:HP5=1^DYX)'*O;$< P4]N49Q\3ULU
PF"IK='ZVB7P,CA/M:_92'NC)(4)/]/8DY+@GPUV++(D--6'6X,M@?/2.SD 1/L)&
P9;# XNS>7H^;>J@$ME2,TNJ94\$?;QI,\\CVTX,AHX6G[:.,=L ,O_7NM3EZ/*$E
P:^"L;!%#'(==^:'40?JT@P KOY+IK5;;8BTB6(@EO@=\S&@\"9ZFPQ3[#=9W:'8W
PZ-G >R$\EL@E2WG$?I:L^0/#!^V9)!$<:^Q***&2;'L"T8;3<\! <$:U)G&HXE#4
PN$=8B!*A1QA\<Q>4>-E13O:Y"MJ?J3V8F_BK<4(QGY/Z(^J59"7@G&>_?1\L"^R=
PNX8I4@=3)3(AR+PSH]84M=,F:O+DIQ2YTC$>@VZ81^.FPW,2TOEXUU^MR==7);CS
P&:@&Z469!6IBX;SW](ME*!@CV/C)?+TYBN[!(T#>C.KGP7QQ1]]<K(&$=X=-M]ZX
P=N"[HZX.U<HN<-7)<L =<@XHF\<CWS2"W[R);S6/L=+9_22?D^Y:9J/ZN>ZQ0T-3
P9?";C_A&:H$P:4S&/9J,I_B[N\Q3V8D]I@)\>'*\>*%C]!I=G!@V.K>"G'>LQ,)]
P"==U/_*6IOHR^?J @,:++'];$*Q51;SOG0.FDR<BWDN4@A=;H-7U!Y7DQ#L[Z4\1
PB^T1N0$+!@.\Z:&H0I1\MW[^RA(/!\G["%X$O1L#3!J3X\V@';:B;GE>+6%0N0Q/
P.C1E<^2!G=;CXY>36KX? TYEQ<B^M,4[/2[\&X=U^VWIW7V;F&SR=SJHY0D?UB1G
P_@\X@8P,Z::?H)&("0/U-M2XV ^ILQ-=\*-O-UYMC+IDT?6")>(9-!:^'/[LU31)
PF>-8G2=J8GV]#"<'Q7V*N*^3ZL32M\[D'0:<L35:0X4/7R*_K^-HN+M]HY")YIXP
P#9Z<*,L1FBS-=S\U'785_\3!A&,B#69[].(AF=8'J++ -:PRXFO0;#F@TX?J>U';
PJ8*NWZL]^O;@YO.(=RE*\PV.3)4J,2.^M3*:0X/;MTCE.G6OL04<A:[SWX6J-0=9
P+]J@5V6MF&WV36__-HOV)9LKN#Y(PB70T-EB:_XMI YV:+!HWF]/5CK&N+&4K'0M
PR_G>%(CW>]?&"S:4%R^BUJFVAJF7:)W5LH.[QHZ2CH],KIE7@'\(X_1&EYS[0BY\
PW,MO?\/VS;=4)',JRC6UQ^N 5GN@MU1CKLGNV=I_K6@?DDI;<"E@TP,!]/T9JELG
PEYWL=)M":"1/G)[T =373Y!ZTH*0(H#Y/A'HJ$5.P/)=>K<RPH*.\&,I8QS:'MN2
P#+$2'^B,\6QR9:DE&H.LM]34[DIWAM%9,G^ 'V,K=@*&?GK=NO[]JAW\+3$2F&,W
P*$L3S&J!&: 9B1KL'SN*QSS?.X:UB5)',;.2BP]$]4.V' ]@D@44 @K#>O_VW-IA
P\K,YMYDTO7:'>>'(?-DVJ<4V-%5@&=%/41E1U9!QX*_:^\? TL46E"+D2(B)=YPX
PPHGG;R"VT;/%[8T:^%VYIGN&%X:>>>L8>-^/A3K!(^GT@ ',F![?*]-9SYUREUXY
P/*QQ6RUPXNX!7S*4]\/FM_!A<0-$VN&>JUW09M=;/_!XG0V=<FL2KUE N9.5E9=1
PE[=U M:V1%I7JR;/6Q\JQEW-&'%KD'51F?M>4<F"QE<0QJAZG[MRRPJO*7<?#T:,
PKCF3U]0R!]YK3\AWYKL$7=[>IQ%>I]Y<]NDW6:I0S'"3B^Q ].S>,0CSZ+)4)EY%
PU*M1B0!VV_V59Q,.2]=U^:^ISX4[*%;ZJY=1$+1J0SK37T#8CMB9P#+U\'"^+>MQ
P[%/G+[4NREMR*Z=X0*D#_EWFJ7G!3<JU%>$0[N.N*P3(;V1UHIS0BUZ4%TC]'3^+
P!L< J&?\?9_W] .(&'Z:!;<D3E6Y@_.Z%LJ$ULUM@FH5/3;IT]_%:^K"H] ^&"]U
P4'A[Y.UT'!?P*Y*#N[RYSE&JWL+ (^ ;-BUS=ZU>LEEC=4JI2N#F[(]HQJSN),T%
PVE6.KH/(TK\2/CPHY+-DV3HOF-V[EG2TU]E#HYX:Z<\#VJ?&R)[Q,1C.04Y28B\Y
P+.(^;)P1*<M?E.8H4_PC=#M1]\]3E1,:;C_I#:H\P>6O3^T/?"9Z[9UH']+L.^+V
P1;W#<#A7K%O'NTUGA.!#I.=\+Q+2EYZEV4H= ZF5R'C94O5"/4B_L"<(LF5OFF?R
P/_O Y32KQ7+ QIBBAR9*WA*0$OCQ<I49T>:V*>I .6N?V)3#;1$ :[NT7.[CM+W$
P3C!^, .]23.E;^TF*1ZF\UW$YG.Y-EI8NW-'@V4"@)4W5\/G&&38>4(4I.N]_?]1
P?+5+RHPK99R=6P]"G_V:%,L$G/@!R/Z]12S(C^\#?'_"T',\,I:\*\'VC(2J'@\<
P/<%$W^<N1G:]+K=O7)*47;AZ<6%S?_J3!?810+<3@F^5VZ/;0ZKAAIA1X1*'Y?H!
P31HAXE&5W?=X.$8A28[2G#U:?G_7$/V14.;?&#ST;4<7Z##]4+A!1L^L 3*T.+P4
P^)4A@^QM6G:\< %[;=YG?N3!IQXAW+OKW%$ID/7(&.JUYIY(N)@M6CU7QO\8KL-O
P?PV.-]D\+H]U8^JNWBB%&2Q=]J2#NW\&HYZ?^EOK%T393E)@9<"RN,:#B(@FV2G5
PO(__1X1_R"LIRC-/I.*^XF ZS"=L9=.BU"%%5>UYA#(7HTW%&!^25=UD*0GR?$BG
PVPY17P?&T%'\/;(QW;?H5KDV<]!]BU^DQF_U1Q"6[RK;A,'00)5""8,W-Z2PXZSQ
P-][1[V0.A9:8,!70=RF"\+(_]U;<?($JROSG[_@&R#G1=ZE1-RXN<+?\>H68]!7U
P?[P.]CJ"L8RQ@#RU(+\<OEM+%O^D2 6K*[(/45-J8%'?N( $V/:689QX^MLX:.1=
PCJ>KM%;[E\>GB6WU,.N!VDU;].%-78<"8NB:2$HTF%HB2VS$?C1&/+E 1C1-8R4;
PR:5]D?UG+O7D\/@!K&CI=M"X!<$7>=.%23I3%)']GOPMM=SOM;M3$60*;"P\FQFV
P?#@59WY?-<&0G$ZW-HLEB:$OR5,IDNTIQ![D("7W0'4]<ZZT[[YKX38GV=LN2VZ.
P[" P*9Q)^EY1T)4M%2?-X03 ]B%$C['?!<F]?4H2_50M_4U(\;)';QZ7>( M/.;)
PLPFZYF4/,V\AP'Z.!L#N?BYW SVI#^'Q=V&Q=0>LG[MO#X\R[[O1-5P>(7B=H+81
P4^A6[UWX>!V259'W'.2"G.321[/W3SABR1YL7T ^JV='.6K$22#E%"MX6^?U#BL3
P;3G!W#1IH?O\A5CJSPG2J/33_ $U:&S8K2*(.S1P*G:B/A#W.$@NY#-QC!O1_.U>
PZD["%A0VO()2AV"Y=!=7GOMLK>\57,_Z=MJ)1"#H_O5]I#.0Q+MIUV:@/B3-HI^5
P?8YT5U\O14"WT:H1>\/A7)A;P ]]Y=OEZDDM>,"G]*V+V5$M(N';5WZXGOUIN&WN
PGF>+[?VX9<EQ1P2YXK<5_2ELW0LM%XI2IC:U.PNC-(RX#5NCO\'3TBG(6[T^E!E,
P:8<-I_G(#,^GI (KZQ+EK^1JD3@UJ>]^UQ.GW?:ZY2*Z;#=,<+%Q,'9@RX<[VO'I
PQPY;T,/$4)%P%9FA'A4WMV0Y)HJ^:LZ[V,ZQG#,\VK@4WT&CMVXQ55<_"&J!/O%6
PT:]MMQAHNS8)Q!)!Q*:-Z\DS>T_P%> +9#S+QTK0+B[XY-H3!0Q5LZP54#+>VF@[
PA+K5C;00#,T"Q3CINK4 Z1]$-M>$\*B% 52.UJV%M#,0W2@AK3LR1H3:H 9;5T3;
P@4EV#$Q[%_T@8/"T<$VH<#B""Q?R%+^W!<3Q7@UH[4ID [I&4>$@QS53V#?XV8>C
P4":R\7@:<CE8=C-7?=W+)8<-%A#:%ETNP(D>UZ>(S3K"YR7G2TPX5K$W?NR&HITS
P-]-3_>]0.+F)_1 IT"VL>5#N\/[+<8;4VNHI@M"'CW,5T/O=CLXH'TE\&_R_>6P-
P\YK7$%PNA]RUJ8',L_G5O.FPROT^+'\ B6:XV5$*-RG"*V1*U2U1%B?GR]8(C#,V
P3BMI1Q5(PB]U?WSEY>YG7!?-RT/D-(<;D<D\;0&RGOH?^W4R?I-\BZQ[;*6 /I1O
P7S>\'SI$6%X @M-JR"*],I)^G.FU_&<3,-2!A5<E/ J\385_&XNC*72B.PH1S?X&
P9)G.R3)_1;( D.CX")=/SMGA]!>U,[L&60\HB?$3.II)&&LP9LNJ=C-I'MDK4;)Q
PL.Z'>\1^G^/MO4R>SG)*$. UPDC=5K X$WV)(@#'.@G^KT,)%[\_OMBL#34[P/1A
P:]F\MS%+M\#E+KB#1>;&(&!<?%YP);DRB8HM342(&(76>8'[A+,;'-,,UOWD[3VS
P0#2@[\QG# CR!3I)(S2R$6KNG9?W <_Q6H2'G;C3$D.AES.&Y\V&BRBL"B96A*J>
PE\QB<B@E5L&O\S>)R<<WD"1KBX).-C^]CR9'L\9&O;A&PA)SH0UZ61IQWD]8HGK+
PD$P8\4ID $2[87K+Z2Q,_;\!2!45.&A5:^>\OQJP'#J:6;@QF!H._&@W)H.T!XM5
PFA.L**]5)!X#ZF$]O(@*H*<1U<H2/1&>\G8HD=T.+4[/@$#)@A425*_FSZ'0I"0 
P.J+1]*/-/1X"5E0)QV!)]K[G*'PG&S@I/;45?O4!2ZS7@K'D##W!'K?>H<^J6_==
P)584'/I5@,2@1W/%IVBS53I;^URO_&\8Y[I&/ ?15=V!4QP_>6 FB5H\J6-V+9\D
P>SZ?67*:YFK. <:WV A>S$%+-_CU-PPM:/Q!OV;,#L:WYB:>@'=[_QZ!T1-$5I_$
P:#,8QD*0.%<MN?M&$H2!C@=Q[F<)D13[- AX:\/0HVDNX^RCVKUNC@7UN80/<_(Y
P/_BN.V;<S(I$)0$RX',Z'%S>3_#,?7_K$C3LEGDCYF_EQUHZ_G0;7;5)3EGXP \0
P)H DZ6TV7>\&(YGZ<K 5I4L;K83]K1$]9 K0PYK=#"3+I;PDCC;9;R!.8Q^$, -;
P+VL,3.,)8.S95))">M\P;D,\)5BQI3ADSY>02O7R=+7X98UI+P7V6P(J_!Q9[5;"
P>%X\6]J+6@P5='_84J7E +@VI3KG+?E+#5O'E:U=(O>WV> ;@O07"GU2H7XZW>@9
P+\6H@D-_@;\^=0H+?Q^8QOK%V4-(\1]Z>H<)KV:X%$@;-]M42PI!DO7? F6]\@E!
P09U(SN+I1,H[C/S5BH9/5WYO=[)5P^6CC$OIZ-Z)"X#(K_ HT0# X'-XG#GFEF01
P'*8Z[D!SO' Y#J)6%9P+.RMX?&^?\:65AV;5>LN""ESUN!_U?6H=&*M5 @$CP16G
P'-[$-_\SL3\JM.-"#UO6<XJX60XXL$\\4";G(Y$PQ&SF"I2$)O3#^/"<#6#PY3(N
P.+:AH0D]B'N64IB#$!*!!EH>Y#CI2"JUCDWS6UDU#VSSK %W 1VF;?:,"QR$LNDB
PC0=P"8.JK5E,7=NY:[7,.F\",;<HI'^CDY9R/VT((:EO;=P^V\SQ1HTK_3+&9#R2
PQTI02XDVGM*]#//!B!6BQ\R#UE1'JVD;NWR_ E;Q%*T$H,FX+<U/9;("Q-JYV8-=
PYN4G21&127IE<82Q:-CIE,),)9P8H#N>V9 RK7A3;_(+^UX)C-)V<_[#RH'AW=41
P4DY2X!@UE3C96#'T*EUSI91 JZ-\E1:TWZB3 G0+*!C6*BFAF:;8)->WSY2ZL9D8
P2&3\DR/]*=2C9W'M%&> 93SL9Y'\FY*;116[C8<-0I*WB:';LZWA*5?&?_S9V)J<
P_72:U&$_Q#S+R_8'>):=C,C9+FF9[6 -?^IL=9^/>G= 'XR)!,,"@0BYDF ^45WO
P@54YB!32]S-_^CNF+4(Q+,AI+!'^02ZY?^#,\EQNYO5>*=-_$G=)0(E_>=U2"&82
PPF-)M7W+O* 0< D&FJ"0^*>)%8O"B'83>/_4\"ZQC5*%NE_IO'?X)6N3T&/C3!$V
P/CH:]9(64QV9,64FG3?7U%V5(D%U$<6-D(.AJ^H3HUKB0'[TW$6;\AU$M*'+.CC8
PM9# !.$EIZGQ1]"J<*K72VS6=E51<-P@P&^PG< I?F8RSL22/P-2=W\ F=9LWDC3
P^)A"^ \7'$.H$[0BG'H[HKD$)2>D=V=1:09^&T\DDU-E0OH=]KSBM*"X,W1$@\]F
P6=EXKH[=(&XL_1SJ8+VTIAAG@D80S:QRN^I2SN2CZ:2!Y4!*!XLT*,=$HX=.'(O1
P=;WD,*N(R")% D'!1I:I,R*.M^( ;)JZ8<5B+-MDZ2]ZQ/&UL9FJNW*98YY$RMZJ
PO0:I"-#ZS4@'XO4"$W@**P*=%!DBHKC3]!V53:SKOPE,/ZUM-!\E$5<>.UI.$,,6
PL[H0(-V"!7%(E^\&?PF=\&N-V;%18(8M^G D]@$*4:;KRLZ<"[6AIRFT-;-T/:S^
PJ'EC2M+CS>@1-7I4N1)VM9ZC;W7PE$'/Z:8IP^_+>)U\@Z\YL3(MAMDYA;9#R ^A
P-;.KUV$.RE.SX(=JND@K\+)LS?_T3W1'Q+'5;*#Z>!.K>'2F&NXOYQ#H I9FYSU0
P@DE/59AO"\/YMI9$! ZK5V>8F.9RB<36M1+5KU]J;KK%M41%I>](R_TCO!_3B2+M
PZ!DL8DH&N,A(C.R>QKFR52T!QDY6D]0?_+#L&:<.'N)J-YHCM(P9<>0L+L? 'O+_
P*IGID6N%&56FH,P*0:-G=!9N7*ID]PQ(>Q9@ &_K1ON1_#J-DOT$RMFU:L) PJ]0
P+F21.O&501F1^]=JRVOXR$+->F 4:[D6 X)L+JMQA4;O"JS'Q*?9/U.?$9K5VFA+
P8F49P&I <2C72]1BK&?"L^PE4()"QG%$.NDS5.5C<WG/Q "?\WU WHGI(V^IETF;
P0#.'WQVV5Z*^P-5_<8"Q)]Y&'9%LA#:4OVY7*T/+ R"),3P)5P^9C$8T*SI(-BIV
P2N03U@QO2EH4*_)6:J,YS.+[(%MBZ(]<#CG=63';KQG#/_ O9Z?EF2>4[Y<X[PR&
P301^:;'3^"=%-(:WM&VJ&!D[>E^426']B<D%^A[DN)]S9_$K:J_9^UX<MD0.]5@ 
P^!,)H3WK[LJ\2ZV2_GGV\CKM+ 4J3I6/ _"H/8&,02 )MSF< QOD?(BSTE'@G77.
P&M/8\;\[SF '4RE(MN4%K!VAH;/CX[FUX6<ZE#,;&J.F26X+.OU"PSJWDUO'7(?\
PA2XDO1$-1HE<*^8<>4#6-%8"2L7]G>4-%A3*UNQ=&RXS+]4A()=5.H(GS#=8^A7(
PX^$KS$BC"910-U@:1#.(=3]+\7C8E_2YBU[SH#Y5FH#;JFV_!&21"9%P0,*^UEPQ
P7LUL=K?D9?$A"Z^>6%P&&/O_51;5Q3U@UPHW^IEAX+"\RO2WAL+4LM:(N+W<IDPW
PJ)>MNA[,Q/I142"+O923R80.&+G,E1@@;0^FZ6&7?@M_\4[0@Z!26HTH@E46,PQ+
PU,0,Z5LZ5R24X'7Q4\'.!^H3LTP"+>$.(;*X8UPY8Z<J2/[<1=XJEF8W"JA\<%2!
P[UCV*QHHNU!#M2+H]I&"2=#K>3#)?M)W%6G#Y,:AGT&N'U,?C* 'RW&^\R^L7.G'
P@WHG#*)91G87BO6)LA((PSC8D.1$HRS0X[Z2V9Z-.5!MZ#I;!-G9R+_$UH54GN;(
PD([8IR=<)\YG&P ZQE]ZV)MZ67G-&8&Z63Y/N*W[ \44CN!C6F+]>!=67B<QS.0W
P"H:B^J[I$1M,2:]#<:N7,!K-$3N8Z>+4RFO$MHWAFA]L=!9/$SDB"[Y%6&/G^!9'
P+M'UB6!NF-N(0,%_,:82+/']*UUVWKKP]4,UZ_)>-)<@E^BC[;5F(.-R<CF3PL__
PP:J+K_(!I&D%W5NX!0AQ<JZ!G%*.6G',Z##P]1!COI=W8'\;Y5/RT2MM*HM?P+KC
P([A!_8!MHAPACG@AUZF+B@(6)2G^WK6U0LI5C4D9K-4HH%5RXF%@)4IS6>(6OHFV
P]?K:H5YC6!T!HWYSFNZ9D&^=R>U\HL%3PIBZ,Y[VV=&P.RS.G:A!0N:+5?\-"-[F
PDKR1865:?S:IP^+7.%*V'.44TM1KDSSD[B'(%0%_-8*LR0=;LE.&G O=]^@;;3# 
PC=TA,9$^0?+,\Y!.^DC=AQHZK PKT/M+)R@=&IK8) .RWZI;K5B!%X\S4:OE:[<E
P*R)C2K<G=7Y3 /GWW'53KN:^N#W#3M7<Z+2#!L'O^%. I/UE+ \3/(:%Z?5+M"'C
PB=.HIC+ARR>&X" $RF6C.*!2]HC\A-7;\% _S'FQ%;(/ZMX&KO=,2A7@[O._#PB$
P6MI9#CE!^R2?E:BFCB5>GU]-6JKDE/<4)D]D*%5</R5953P,#BBIQ_XKMZ[CLU-]
PG)LNMUZCE9,6C>+5K8&_I6UX)SD.YUWR3U;'\>-OWJ3*H3^/.Q;-NN+TQ/?FL!'C
PBPY=D!O6B9C:XBO0Q0JE*ML+8+&#\X\]#1BL<Z0&C1&M$MK=#1(ZOT<+]#*L>5:W
PTF9GP>Y08X@HPH(9[4;R>GA=\L]S(,J468\"TRE@/&EY6V)='CU_J\.9P%6J3]^-
PN.,7!ELP>TF33=$BN-ID[O[N=#=]S</)A%_PYL=>5P*$-D.?0VK6>\-=9>)>K."B
P-0'4S<LW5C9<6N<)9?9. J%T?'?UI.:0PE!^,*!/%G;FZ)PK4.;Q7%7L UTRETH1
P :K6*9KAY1E8SL;47:D;LV?C3'F$TTI8?Y*E9O<:RXT&GTV^O9V-&Z@%$P?TK$Y$
PQ$P.5 =O6S8+)<3)/,(ZLA#8Y:&35LG#M)\R+^7L/AHEO2$"C#_:>NA79(]1E01C
PFI"D*(IVF'?4)K=E(]QU=0EOU?,J1!K\;7V'K&(U2S9[E+%,Y9^R"<,GQQETYAIB
P/SBZP/J,F*,EPJQWQ#Q]F6 Z'5\[)L=2^Z@&-2$2B\&:$Z^-2\C^9XS/GQ'LJ-:;
P!)H$ \"JZ^!;/).8=+NX.".A;4)*MHI0WZ0>K/GXKDGMW/<()TSO'T!.=G7_: KQ
PO=B1+Z\4SQ /1GF"EC(<;&!0J=R"*;M7?<4L?C-9*(8BD%XLHX\HW @]V9^CM CW
PORITYZ/=U@IE020"5ATCEU&*OHSZ1Z I^E$V<W,NA-LX$O2 G/OAQ/SI0_1>39$Y
PN0RD+#1K,(8R15!=(Q%!9)[QH]R3V9*PL8^7@(]R:Q[]<I.5SER3_EG=R$/U("):
P$[_OEI@T7CE2RO+3 ;)( ADPV/+W$/$7,3P'+Q5L#[YSJE,^H@-N0-8Q#Q.HJGN8
P/$LXVU(TP7=VC75A>8R.\N;EM:L"]7@./_)H8+;[]>! %I1N[)G&T(]Y2!NLV42T
P)4J*;1R#7LA9>YVU7^4P<.(BQ+2D:9"6'>+8W,&_>%\7%^D>O]!I]%SI>L8%V#YI
PX]=.=0=IEI +?"9&Y<*T"SY.BM$ZL2;AKH1COL5:IU@S/UQ+L5EDEN!W)O,%&BVU
PCV%("V+5V4)F(JZK9(84.M&# V^P]:,V3)/M;SUS#I&D8F4N$-#%;R#6DFP5<9Q9
PVJ0AY:P6##$"H;>A\9<V;-V$@5X1U+ 6JQLYS:NZ;YP^-"X_PJGR783&,3RE%*__
P@ZX)+"?+#\RZV,GXVET,E3POM?+OZP!T.SF@8NB'##H$'IV.W)9G@9Y",QP,C@25
P)K'YWW%A(-K6E>_A9/.G_&5]X84DS^41TZ=MB^SP,Z-">.*F\.>:LX.VA")9HL1'
POJ&VYK 7_2=TZ8:K>JYQ:JH2[RW&/0I+_WNB&/=C;E8.@N^3>O%+?&+2C9JLFE(/
P,WIHFZU#;W1<MJ >5.)CQIR\&:LP8D,]_1U&8:>Y$XE[GBV$0DV4GX\D-!',([AS
P*143T_X'3% HZ#B_3>8HYUN3[M&) U5D!(QX&H&J9UGH3X;J1'BQ3SFKW<L@(E3B
P#=P*1KD_>XM9JD+P85BD-JLB"& [69U:0$"'WLIN-!" T[,HI-\8URE@7)!)$-F7
P4)58EGRG\5*^E6_J'07O&7>7+6:G)G8%\U9."MSKQ>11Y;U-:Z!0@JRQZ\T>#1$T
PH5;Z@AG$>LV*S:-B$7097WH+8L>A%E;^SH>KN1K)^$C -:WM.\_QBX 583\!2E/ 
P_'/LILZB(XBB%[>XA,&A_>[,2VS4D(/SZ)PZ)C1B(3-//:B&N)#LWVV>+DV;+K]G
P9OZK!N,=LJD<V1CTV19$8UF_5E)M%\_//8E^@[5P'G76BD?>,Y94%84D'RJJ5#EO
P^LB!6U_F1 H&=HL/'&Q<F$7@/@0H@OZ7$)EA]/=*A[56M1R9PT#]3@IS>$?#X1I_
P2)A>-'=M%IUB\86A-!$[RX^:*"M@]"1IL2!2#\Z@E)#1_ V4$[^99AF^#&^G!%(W
P2NT?G =CWQGMK2WN&^-,^_C3KQU_WIO$]'_7_[=D3&?G+[\#-XJD?GG?IT.UUW8E
PBL_UR5*RU<*02^MVJ="3R#:5+/'2:B-,R!.FGTR&A@Z]1/UXG);E"AA<X@H/(,(=
P^KY_/<:/62G 2A[XSW#-!.==WC1=OCLU 3;$751Y7L=3$\7/;J"R!_\DAD%5M9-W
PI,[[Z>1$M333DR9K"O.?XY4J%?0LG4&I0R[.Q _255LB]_.1YTE%9QAL'^\_HD?F
PH1;=_[J :@R_N ,@&'(OA\ =%L5+IN>F5U)':F3$'+DK%"''2]\W''UR?1-$J!R<
PA&B5/-2\G[K:CB^%!%1+*%PFAT.F+Y "CHD2F5;*VZJ+'4G[%G+5AW(>9PSSPRVU
PLQTV2YKR_GL?LQO0K_E"^XE\F57;314VDF[\28FR;\V\V/;]M'@0G-\[4;DR#92R
P#JL<1(KM6"FKG#?%D 2609QV+U.C6YD<]RC_95D$03K;@6H8S4]7!@?(*1GAU"[N
PLAG,20,(*&TQ=7(I,=HEJ0F)C1S=I![_JFY4FR&]G-I$$RQB+FJ69"^6\00J:/?V
PRHC<W3X-><CHG#2SHI=+Y8B]JLX5,]#*4(LB&8=QX/R=-FI]/A CB%S?YJ8N=\$W
P^+(*RII*P9J$47/#*0+;,2L"KQ@ ZNM9=/^L%.L8E?0@PUVFX7NBF$XN"*G[3L0D
P>^O1)&,/M+[(T;&87P*.)^!UTZ> 6@]+IR^8@?6 RV$BYWL&:.=0;D3Z6IJ34/(H
P+;R0_W>I$AYM# T)5)JPDAN%[W20<J?=AO_?S5EZH<0'93.Q$1]BAF91)>-$#O6Q
P,1'$# Y2..Z5!RECF?HCG),1Q: @E32F#^!H.GU(0N(&S&PAJNT\=0%3! 6AH:G#
P)5+*.%39.MD]ABF\FS&GY \&F0[.3Z;ID=^]R9.MU R_&< I]*U7,@NF+V2,B%9I
PF$7]<8MS:+#L-)=X%1]\B8_A%\5Y!<7^FM1AL>^ 1!,M.>"V*7HU4ZY0U^FI$0@G
P7H8L RS([;3BAHF:=TM#$).M ;V)&#:B%T3]#A"$J'^]XD]2A@0W;:BF_=6S>#\H
P_'#C</#>UL=X.X;Y4%(\ZXB>PYEI2(]25=8],^ -P<U/1"SAB^&E#I6<N] 6?++M
P6?E@5K29 Z\<(JK ^VJ"F4*->8:'@3]W7D62)6ZQ-[32= ;H$U[7X['C,1VDY6NH
PQB2I\N"=KJUZ8DH)2U]7]?LI?DR,:!>'U.[^L">%'R8(COK1[A= A&@ZYH(;LT7K
P1,_K])'6) #)>O-]WV L/_32A $H#J'#Z[\CK\*'MM'%L_KORG1@!0X+A@ :[WPL
PGM^FVIA&!_.@]5(#DH6+TO4Y#:VNCAF*3%)GLS\P>_QF<8KW "OVT5G59PB175P7
P]+O.MP>2YI.T]#DNQU!YCB!1OV\8]"9XGC&31O5,HLA47.]8X T'M:.#D<.8<ND:
P4K&P9?K)HQ F(JZ&9C8-IP'.!A!T%K;1S\@^R.>\S,ASQZ]L.<@B@[JYI/&3;?(A
P%$E ?)# Z8%4C'4<_B'R(Y]*:#^)!/KL#><#<_YO=R$=<;XZOAR<+1CVWB[O!ZAD
PT9/89/->X8*D/)PI.HM]J$_?U,C?":(4,D.9WR_C:?+D<?2^WU!KBYVP@LF-N>M'
P0WTLSL*-G7OWV *-]O!T-B7IHM,Z[$<6&<L;/R1]HA*4V'Z@YY"1M>X5#7J*V(ET
P&3LY)>8H!S0AS!PW?9:* D=.4&R>PL'BC2)++&M*:K'!7<GF8E]"#U@K4BC,%Z_1
P[>E7Y%&%A']I ZBIU.!! 4U70/2K=++BH,L2BM!A_&'_#4<8E];GS]@<Z.05A:VF
P:,N_D$1=*>VP%:L@0'\5==MY.:;,)!D%*H13K]V]SE;U,<>=2NTQ,XF\\WZT<-9+
P+KW_T./, )B]M7H=:V8P)$YJNO[/!- P"\@_C\J:L-\X8<J9I(;_N1AUG<BNC;W)
PE('5TN.1E[ RM4(UGM_M[M3CW7PP20P(8'?<7I\/_WF!PS4Q&PSEI<(,0SE7FG'4
PUY5<7BE-R[^G .($2%(:HB23V!?0P?$;=3_)Q+(![E AV2TYF9&!TN=U#FT1KS(>
P:G[D;_0]R,?;QNB.TVL1Q#/)+HB.L5(#((;NC/_NW"V PM=]K?W"S*_XS[,@5KD2
PW4DD2N(/7E\FN%FA-/61:,OIDRHC51*(B^LZO;(WK;\K=5F(WYM/#XC-85[/ZXNG
PWDI%XT3\JGZO,:Q_"3EK'U>G:OD8J@ Z[4%7+*?C44#+7I<30&9B>D&TJ:M>>%/:
P"?HLT0))E)^,G<+B)3G>_+5\^.+EK17M<,@ZED-%O!+8&<;.RJ$HHW EH6YFOJ;V
PGX9PH5=V!T*3DY2U)- 2F( U##E]&]O!T?L+3H<P![W>D=-\GR%:OHCC'#R <XAQ
PZ%4-ZE'*%I:*YYT6F?SF099,D1V'T0VX>>\])[95*[N?7?Z36363_U,@1PZ=L%E3
PCW,C&&WMI+6)XW>OO@F=+LP'UG0 ?'\?[\8AI-HKV=-G$=K*'D8999(](2@1@ZUC
P,9M0&^$^G5X0AY45-I:RS]E(3&0:HJ7S90ZHRO1Y*('1!(\ORST0)JM8Z=QU-UZQ
P2JYIN\,/)@(%M;GW#6OT&RI?+[&^9_5CG:#W$F7^.-S0"B"Q@0*+NPPT!+SC"LP=
P^BO4]&0(1X0GB3J=0?[I[DD.VUDI_PYM?*;N"_U6,5+&!7?!7'^FW'Y,VD],71CP
PI"MMD*66.D\9]61Z)W>2;>8OY]YZ8CBF\[]CO=N"'GDI_UX.S]<L]<.I/'+DEVLL
P6*&J[UMA0 I'&NUG')(N49P""7ZO]?[52@P]LJO3'RH?& V$!6BBM1FMBFX1%#]1
PF,*N;3Y:V&KHI&TTB,Y:00&'!,$GB;<D/XED['<))G5"TTU2[A+J-+[5D ,0@O'P
P*S*E"1_EWLMF4M2X$\,+MBSX$FDW!9GS5[4MLY/^!NE!IV)6$MF[!61:3:GP/,VY
P9LHN)M3[/) T,G%,8X20P*D3H?_CYSC7YN];-S9AZ<$7#8WN!9;TV3F#RM.0F, 5
PLC3]2(KZ6G@S@0?NQ>9YQFEP:%/6 %0:<ITXBO4MKAZFQ0RPS$03Z1:CUYR(H>?F
PA*;A(Y/NDQ+I^GHN@3]PVX:H]E[J0R'-#N$2)TC,]A/U#$MTV9]3TZ'O3?L>N12A
P4J2;>45-\6A0874="'7*4Q ]#E/M778^'.^/9Z#T%4"#'_91YNU+!Q!8-^[';X-]
P '13I )CMCV6 \P6'GMVI3Q6R_G.]?;**X[8-'$K_:$^EYPSKV2 ?4)\%\7]5_8(
PJB1B0X]HVSQ_;44.2^Q6$Z>8+5L6KV[P1JESY[='R>:H'Q<37AKUC2O5S]^@M_^/
P[X?B!+"V&JC[,4B\VU+U>"DRO9P2LJ;N9P3$GL[6Q@5[^E=\-M%=AZCI#C(<K EH
P'/<G[[1$ON#=U*MGRPCQ@#G^6J&2O4F?9IA615TO4\'R7=DP"J ES^B.P>$]*PQ$
PH9[P[Q+VP>N2CU/C=&?GP+4:CB+H7+?EJ@/9AF5*5JY*\[[!:NQ)%9,O>.-TS!&Q
PR]DOHGNEUCMRY UY-7GF>\RQ+C,C.+DOMHBT%T]NEHT0LM*^YHAX&%;]W @W$Z-,
P>' ^\^G*O-ZSI14-Y-*LSXO9&TCV*@BU\RT)!\ *&*%\6WFS?.Y\<T(3STTY XVX
PRUZJ;>]%_P0-OR*"8WTCQ*RW/*OZ#I)=E> $NOO)3+JKG!G-U.)1LA>KJ</ZOI!@
PFD.T@5P0P(TLY$AJ!5&5N+U=[?TO@@LHF"5[V9%E+5N03DG;[M-O^\+L$/F!R,*1
P48R,V51?4OK@X,/EI;=0&<A:JYQ1'S?8:%.K0?1W) :Y_L^MFP22DO(WNYO^18EI
P>$9'LX<>RJ.W-*\RZ&!$@?IYV6G)+^!(;%.6QE#!9 'T3>T*I+CJQG++=B!<_,,M
PV@"-&%#":*Q0RG5E)G8+@GC$&[&G5O%'BN),%*2MIW#"F99"*\WE1W\\8XRM%8DK
PRK&^P\+-I*\0DING[ AL&F9/ ['-XGE-GH,=BN0ZVYDL39^@+"42>-@X/U$E\=Q,
PZ"O&)U:]+F2Q*A:K0?K":P?*Q2H-Q]PH;QXS;U+B2G&#)Q8TNRT1VO>J>) JG,[X
P(R0X$9I1S$V*(4/(TU"+VJ?H]ZKG!(D]OMW(Q6R(_> =(=O(V4\'6"THB;7@78WX
P<\/&<-YJ*5E$_-.9Z[HM".G?[@>3)2-:A@Q=5_=@!"ID#6UR!M-H>E&&JE85JA%C
P\ZU]55T&Z4TWD:MPRR4,4E*/XDO1G$/9[\M;\VJ[&IU:5YU(HD23F')J?L+UA,@4
PWH411-><)Q?OG[';K EBD-7# I$:>8?^@+"/HBH@-KWYQ0C0BXTS[G$[7KXI0:V[
PD6)$@(^8+E]+%D'6 ZNS#SGLSD 5BK\&J.TL5#ENB77;/B 9(M.*N-1J>UK%E[NV
P [&66]B2(B\5[U8PD\B=P!"!/>] XFP_*4M8$D$:E')HH<07':0BQ:]1)L7,A3QK
PT2KL[@L8&H 2_S$OD15[OA\')P&^1:]@,,9,-JGX64W%K_AKDAXFBA#?Q^54XE'*
PBFB!+='"CKLF0U%<?Q&5K)996<H4/UA>4GI_$ <)C(D(Q'S:ETJ&!OCH4Z#[2E)+
P*IVZ,5@_TE]&J8R0UM\,XHB'T-,@GVY =*Z$!]'(R.>%X:?QA V%7O1A.S&]3IO8
PZ>WHMK;HVYSG5%4\3;&-:[("5ZRG;_LU!2C43[UGEB[&_@$K8((HQ%FFVB7DP/:7
PPPP-IPWT#O>#",$_ZLT8S\%LC[4)BJD5Q#6-0U%H.:N6&NXO@9J48]'1.YA=7Q@)
P\F]Q1]YR<Y_-F%'_Q=0X\!5$]6[N(H^7/3NM*_C\;_9A/I0V/B\?7+I0,T($L/W&
P#Z>/#P_E(UER:5>C=121U)I\/[JPI*9X\*8U.X[<UNY=Z?"CZ @EP,7C=N#CE,+G
P^WW) ^;FD%8BU[R=\3 ,1>I$S]=^+##JX?+&@#BBFASEH^+C=]!6B CBKUQ&N:K5
P7R(R5N,?&VE"[::..;25]?QH94C](<SK0!YEWEQLQ4;L&CP;KQW(?1D'#^I4ODZ3
PKL6VQR:F"CXT(6:TW\8:KFVY'.1+*.?[H-3,-XI;=Q;) O"MGBD? NC0NQQAU::D
PAGV0L!QB86.>GLV]1IHE?,=!B]2TMT2:]Y?PY(X]K+$03<OQ>L0V)@3"B,6GR4\R
P='1,J4</:(!ITM2IKKE,7>_"_P_+A&LIFL.?FSZNH-V*1&2SOYON([_/TD64>U:8
P:82+8/!),E;&!M#K&T/#LQX+I?GU)1  X_3E_J?R@77HR-Y]V_/-#RW""9]]&O.S
PIK@2X+A@VLYKFOJ<Q8'1M'/;V:S#NX#R5$I8I%\#BN>J\$T5I1-WHR4EJ\<*N=R>
P!%/!.EL1$&R% \_T$KO8*24G6D!*5G+)%? )LJ&4@17DIJT%N$!S-<FE<2$%ED3\
P(\,GMDD\/PC!LQ<66 (N)6M&$[Z;Y:8Y=*IB%4\:FT_Y\![B!R*F$<+>ZT(KGZL6
P4"&+^+DUD@D",ZR,)^T!S!6!=&Y(M%?7L(FYNY25[^805QUWDO!5VP=EARE?L*KE
PY6ZW>@_L8=7C]FA,+:4&+%>B=K-T @^B[\F88><K))$QV3*DD=1A!</5>/'T$1JQ
PX'? !EB5/9NGL].C?#6TIE3S!!CN3RUR KB%Z<#LC;]DC1$=.!W1;?H.-6)/9OWL
P$HLY"N[S:[15M\<F %4&T+T@]A+: W-090=.F<FYJ=%WV9QIO=;H[&=S"L;YB2#T
P8#\<D'-9B/E>Y<Y12IVJUEO[6/<H1]8 ,8LZWYR=+I\#(I]%\ DNR7 )_-/'E_(=
P*LB[_R&.PKKS(U92^)L$3??I'[*36!M/);$'"F-#)JH8[@[I]GZG%#5BB%NR$B]/
PG7E>B=@<KA.?F9FKSDK_[R#+[&VQ*Q/A=#G[WB!BX3_N[KP G3P,ST&U5(U&VI&5
P5!9G>_B;+X 7B]  ^><)_(53SD(Q7'R"'(B\1T\<]&+ICS+.#DA6;8 Q@5Y@2WB5
P)I-HKUP]7T(3+;N<&D_?54-WR.A\<V-$R_'09CA>:SE*&7GG\,VQ=%Y9?+/[0"M%
PSBBC8W9JFRIU(2(Q,)J,Q=CO89 \T9PI3+8K*+>:=HT9/>^[O5Z;S9V/&OB]LRP3
PFXYP?!3.PW_O9ST^>O7I1@+AIYZ U5#BFJJ EZ;XB.K-Y$269).P&SN$IUG9W5\P
P2B?W*U/^L*-CKJR\K"+8;"K?FHK+;/'G-_14U8^Y3<#?K>S5%@N7]T$)(KLHF;* 
PH=A7;DSQ8RA@LL:R&.^L=U<-PDS^##TD1,+OTX% #BT";ORO\%CN /\X:>+]2X=D
P 5GZY5_F +YYV1-\Y^9FWJ&21%G@J+A)5GG\8@<JFH&.J37=S,0],4!/?3[H<TET
P,XQ$3[SOOSGOHW[\8)X<*E8\$7S 7:=0*)GQHD+2YN/5<%WM$ZV<8UZ6,3D0E4!^
PH-;\4#9@S/^/)FZ#LI. V+!/Z :C&#/@"1H@2/=S"_^?O',F4WO*A]LY@()A-X$(
P@D^ASQ;@KQ6(5'US.+]_4<K%/(:(&O5,U2BS9R!@XY3<@9-@E#\$[.7%&#?MOGK/
PY4?B[*28I*\%([V$-[L]XM&SKY)W1Q"<#CU"17@'<CX4BNKZUR'9\2GGEAX9+-  
PDQ[B(^].$+0-GTX5YU%L7W*^>(^Y;QB^YV"175@P%B]Y<,UCK*&1R(YA#0O^UL H
P;<,Y$^*#]%(4%Z0+9+X5D. "5OVE9TN._]%_8KDFVKV,!V5?9&-F2@37TY59,4X,
PQ$;@]3&<->>98@/&&ZL*!6N\W_0^E77&+.=G>1:1-<MK'>)_1U" X'MU[ZD6/#1V
P896=\90/MS8=SO%HW,OP#]"UN>*,-)C]Q#-2TFROTR(JQ_[H1/MKV^30"5IX05Q?
P(R!)H*NHYI"A GZNFE4K2K%WG_&U7P7["1G/MDL9><>>G3,LA!K!?<\) RZD")/U
P,"$HUHC<*4-4)7+K7^W9%  R"^-'FC-\V$861_RA*XPN%!^J18#-*%\>&6G+-.NF
PQ2^3\51T$SA:AC:)Z>H* CX_H&S',SQL*I5Q4\0Q[AV>&2E_4%0'4<O9];7@/">D
P7 D;GJBY.PVIP%9?+[TG+#.178;[98T'I_=;T!L/U3&)\:U[9KP)<1;23G1BM&YJ
PB THDI1$I'WZ*\2>QE%?E4.4=GT1"6KI)Q"!U(39VA+D"V</NC8.ZH:$H6H*@T\U
PYR4"7OA4=8""=U'$QRNG!',O$/F+!M0(N9%*JAU]M.@9"59Q +/9@EV=LKX/T'V0
P*C_G4V(5"PJ5+S"2O'> K>1.C.UDZ)E8R)PRR0")>6S3R4%3_)G(8<Y_YOA_=PQ1
P\C<.T5?]1?*KR_':1?LJ0'@#7VXYP9>8J(HUA$U3)OA$710//XR1!SH7 LSMN+.=
P4&!&=H/D%T<W_ PGKU2*57](0PM()X,A.=, 4]AN=K^!2=R_>O:_[W;SDGLJ$=5/
PA"W:"O6P%JI'^:E@U-1:D7-_0'WD0@8"?S/QT,JMM04%Z+JE%^OBZU7=>SU%A)RW
P1C]RP]/A_A@2V"YXNIW/P)-'*?H,M/.,C"8PFJ1*:#SE"'"DT>L>?/Q7E?!XP";*
PFOP!U#C445!ZO9T\>Q1B!_'8]EB*=_2X,YX13((NG^,S2V.Z=*.!T=7.!(*9J>D*
PEXDQJ;.H1ZD=;J;R!MV0D\'SW,3&('"#=6DS+?1]0T>0O^2@<*IX::C>DT<5>4(I
P7W 9<-ODDP'/11:W,[G%(TP IQ^KVH5\9C9UWZDC:3J!H (4F!.)[GDKH*(-0(O#
P]L5FI1]6$I' 9 +7@B8F[;^A7X1[Q3KP6!F2@F4==!ZH0/W<94\QX]04Q'/4JQI6
P7T<OE9W.0Q$;QE;J>,^@7$%@F-4-<&IS@Q^4^HV*+[RD(1"5F3*/J6&4:_X@T8Z6
P?&Q>8O&QM1_]:]3#+NCC)!?0JE CJZB9\R.&[<\J3#)U.Q9LF4)6>/7W!4@*R2;S
P#?S2?%#8&MLU/-]I-B;E9T%JTPT,9.GF4)BYX/3J\)I_QA "]Y2&];",X#Y4:6JU
PVJ8BFENX^[<EO92S+]M93 )8-NE 5+81Z^X2S?;3&E(V?P5)717SNJ^2$(8D7-@3
P(T^D54)8K%C>8UC$/'NNL.9[Q-<?$Z&@P9]JX:C9SZG^ <D7(Y(XO 58@6TLRB;J
P>][83KUN#<,1OPX'Y<1X/"SFSO@G."/*",MG/$U'#2P>E,8 B42E; ^SQACZ8A,1
P3]UVS(:L(F(<=S3K$ #-CTZ%"A*Z6=4*&/SX\7\(_"<,O="!)>!;"!'C..O;>\%6
P Z2]8^_5&L9":C=ANF6C#U H;<A5)>SQ%R*Y"&\%P9H9U*Z&KO=*I9PAOO; [PT^
P M)%A^B2E+3$8 'G<4:\%*'M,$75>QTJMV2X)=V(C@Q=K/ ;=]8L<7RN@B&1&%\5
PN<%917@.4HE;_T@EYRN'DV6OE]%Y!W!=GR6<]&Y,8NC$DL7@J/MVUO%G;"MSJ@ \
PI2P7>?]L'[]@MK9X:('*CTFLS BA_"[$4>WLQ*%6_1$A_*W_:+1=IX$[/@^->W ^
P9<8671H9I]4K9].YB,6+3S%9R@0@/I=:([0VEHWY>GNZ:3(X8R.4\0(]+[WXIU:3
PW5+Y%5T]F6_M3$2G-$S1O2J@U,0H:.J%[OURC:9PX#3"1Q +,8[K8?(>VO3Z^(='
P!TB7C>/1*G)C9* /3W'4>5 ="V-^'YIJ54@M[RKC,8]$V*H\VDU('6\+LY"?R[16
PQ_N]\ZII5]*V_2/"/M@-U/!K@4(6.6]*$DKM.3R@F+VTT1!1.(QNT.42-VS8INM+
P<GKAQ9>N"4AE+#NF79)&9=+X S(L,"3A8;3+7"9#[ !9*)\#.J7#V<TKR-";F@=N
P@ABY[+HM7@''<8-)O+1,66@, *@1V4_!&=V0\9)J==.8.K)LW1@J\_ULF_/\,H[=
P:=TV-E='VDA !#4Y:D>=^#_SYXY^KX#Z1/G/+..'*,E$\LD"BM,J?'A%59^J*''R
P""A[,Q"KJKW_Z)-[Q1%09&AAAJ^<3(>+ )(0L_?[)[OZAANY):HHWN \LS[5EIEQ
P3XB>@7$H&P11/Y)N2TV^.;#!VBVQV[?["?'+Z?7=>@P728&J[8$J[R'V+$,/#/B\
PP^0E0U2%8D:G?WZ@-0C2N+HRS97ST/VSIXM-A[.<QS1PALG'IU^&0%4W)NB/:*>"
PMDK@H#E(>B_"\>8^S)!G>W;_QY3+0H173JO3R,)$ILL/]2G2G*X/B+S&1IY@F)&(
P*FQ3.J&W1ARB\2;&V( 12;AE(Z:SJT++D"KEQUCRQ<:ZWZ*'8\T]@T6I)@'+6*@H
P,R.>2V\'LR!92;U@^UFEI#5KX\HA'T-T7G4=]87SF0LW5F9&,8V:^<^PEIRYD7UM
PI!,W?27IE3GDGB:UN %PN"9;#0>SNEY]6+0C'1[\UWS4/;)4Q\W^1!,46MXX=E*E
P F+H32GH!\7@]7-6[4'"6[KKQ'UXG!_J5RD2BYN4A%#Q31[18>Z8]9\6+:&]25FP
P=X<HII+1G:,!GCEE=<][.$9]E=/W'$Q1>='%A7P;'5!+$AL?T'8FC@IA-$WA(H:<
P=2"BD$RHZO-;82!XJTS#Q7X'KXO82'3A?9QP^'.N(C#CA46\^_W>DWZNA<[X3]<?
P31:K]XSC;<$R1#0^7(%((VI0GN6X]?RU^/MB' 5-\7HV9Y^O%WW"4B/3N6W/GX5?
P9/RT_BB="AC> FFUC5@4+WTH@&R_2))BPM?^?\0W<,_(5*%O( \TZ W4]R2.3Q M
P8R.Q'-M'E#X(,V8JR7$W(99R!9U$GJ1N#8ZRVAID%V/IE"I7;VP[=&1+7ORI!_K"
P#A!3GQ]0B#&UY>2%:*7+N#KL$T=?0 8&I"OX8O>&?#FO%T?O1+TBE4]FR:LD%7$%
P@[P]NQ9UX\+9SG)15F)U3^T^U'"MX:S,B8Y!/*L^O0_Q1&V @+#\PN()'X].#1B#
P]8HROMEAJROG6M17O? ! X$XP/=<XWA/>81?AK*95166$&Q&NS^P0NU(4@/O^9Q!
PW4R.)3H?O\CW_CL1_*6E5)W='#J[@\>XQ-@G2Y];KR%%-'X30OA)[JFF?*!I?N0]
PIT4M?#O!U2:#=:;>)Y3=&NEG77&#H#"VU<0FV=^1%9F^V,&@X'/RNH'088;#%WLO
P0M?D<+3*H5A9AL")G;C=!.! ]Q-Q'#B-[F*<$T^]FB&Q_1[8"M-P]>?Y48/",248
P94!C.[R,YV%$1M$R?![^+L]5XO'<^Q95_IVUK34!9%%/X;40-<Y:5[JD,'<AF5A0
PA>J280M1VG25+2N&]( BB-O>8R9Q\PA\# -:%5"KI%=8[.&) J/R[>OCKO2<$($X
PXP4HK@,^@-9PR]^LD&"3Y,TK@$2!7!V)>HR2?8]Z9[S]0MM\!A*#+E2+&A#%#RJ:
PN^"SQ 86G]_[C]9R0[TI$?C> @%:R^-U7A2&5F@HFIRD?YPEY//(<%H5NLH!PGK9
P'E;#52PY\"N35A=-7(X;9=DY"X^H!PMR5[D1D2O[86+M[B&?*#05[4*GC"C)E35%
PR&Q\;EZ@FX$+ZY^C/V*1_M[)+V&RS@Y#_>&B03WK8W>7S:8-1^&C;_9(]0/#S/U=
PF@",DRU RQ\5+"S^]2HIP5#=Z[ET$]#5Q:6UHBU1/L<L%_P>/O>;!A&[8"A_-!!0
PG2Q2J'NI\=!Y2C$4]]*H*F^O;"0I<N#ISH< JO6A1SJ>]BW=X<^D3O].;9*I(\GX
P=X@KV-P'$V!;FL81+-(U$,ROZ\:EK"$P27#(0]>^.P.OH)JBG(@]4ZTQ9\=]M6]&
P2KN"$$AJV6\Q9) $0<K& ZL<JXSI,,.2K=?ZJ+?F"_U#_D"#]U5";?NL%"!8E[+Q
PY&&<DYJT6T=>DP%@2ISD_77>. *-4".!GS/$1;,P<=/!O(X_N]JR$74#CE;,9RLJ
P16J77\VZE#]Y,K:!Q0L\[ LX$!!&0UC*,S%;Y#(M]ME(]HCE4[9Y' ;V2AES(MG]
P#=^&FTRJAP?+7GM/$" NY;WWL6_+FH,<]]2-V>GOHQ(++ %,/P7!#C<Y3S$]2H@!
PZ85D)8_W3_D'F,]IOAI7NL\X2=LCVMCB$,N0#NR&9T1FE*K5ESM\@-12(F0NB1]M
PV#:NFPE[C5BLA09NE!WY?L:'PXM0H9@!D)IR.[_&J\W3O#P;,N]R2UX-RC2?R4MN
P!1"\XO^4T\AY#2[ :H!@"CT DV8-]WY-;+$I@=I:_YR&7#SQE/=:N@9\:&G0(8KF
P?)YK'6UK^_9!R2(J=8$\';U>$A=\01HYU#N5-8U,8/.,<>%A^U^='-I[G4,"J9((
P(WCN&I!23AL$KBOR+C+"&?,%9!!Y$HT+.$-^RIIEE0L%;HSF2Y&4E((UU&L:!I6Z
PL%U<,'954)1.Z29DV.XZB)D7KH#PA&SQ%:-R3B15#-NMM2/=O'X_KD<US_^%#YCK
P'!%W$1I(\O.WMW!5$?N-IDE4YZM7G5SP4JD4HY'%:YA(>VX1P %N<*.4H8^.@VSE
PIR"OP;=S@?[>[<2&K3?_S8Q2=E;S1=59D-D+ CD"1%'91N6.BYF#4/3!OMW-Q%(A
PW"["9(;[/J625-Z%U"B8 ^%=2&I8^ >"TC^$U<UI9UU<!:)]?R@6BG+P!=)R]5WC
P=X+*A5HUSV\G_-XV^0EL6Z,&E_$&@@[0O]+K^/P#:R<L(*X4Z9-6/EUR8Z#RO[KU
PV($;JJ-*!NAS]]_(VT7_.\JC#9J\X5P!R)!O*T70JA5,*6XFP87 >=Q/<_^7E"<]
P.GM>&$A1[^%X6*2O"?5<[#E*17M4BXPM,.RVQ=ST:XLSD)<-_(U.L\FW-9/Y##A.
PHBVD(.4U*.#$5UJD>'0ZCXG2&R%@R7@,#'A%W#_)\J'BB*OU GVWCFZIX+GZ0!!@
P89-"&M8[;O^\"L<8(,'.![JA C\?PJ"*F,2.&*5[!* G #RAWYN<A4/*UF$6>9>*
PT.(N<2[Q!^Y:O60?[[26VGDWYFM-B$]O@F'X]8_W!@]02T/)S/6^T0-S&_GH;,G5
PPF6A-IE,V!>?\]_!]@&WE\3DS$#G>2U*BOI?!X@'Y$/P)"176;5/&,0E;8%W!6>;
P0 ODTRTRV.1)=2253FJR_R"*.ZV!O5I<3)5T@HO"  > 34C.H?MP<@O@7*^,_IRU
PL5#XVQ=XL2VJG&V[%P>3KY8RW_#^=#>FVY^XAG'8G_9];O^XKQ%IG1N_/X0RU6U+
PW 3PGJ?WV V0]S4G'NJ,[BX;C\]@OW?CZ18YM<Z5;UAI9J[</..LK,V(8$H"?.+M
P[>,X<8K[?Y_MO00729R0[ Q'AM+?NDDX#(/;07GN\Y8JP? V3L!A9>=2H.4@Y-^R
PHB$LO-/+AX1SIK7=B?&K\Y!XY)F<PB)YN52GK7I1X(A-#>2%[(!]X/PSS9+0JBKG
PW"3M/IE>7EL<V[RPKWMT"XFZZQ"DQ."U%'6="D2#1#9$Y44491D<X-&BXD26#)%7
PM2$'Y7+XP\-#D*!?MCJ&8J2^\O\7_<]5/BD3V35\-X.6B^W<69<YN#BPO_\,J,1,
P""2$F(&Z?&\739E>] MK&A1VD,T&;[WW5*X <9LM*V4@6/WD;%2/A4\U=!OY__^^
PL(Y0+>G"U6\F- EW$NB[#"T07A;+GQ3[^G,<M8GR[%O,\8+'[&I$DRA[' .C:X)W
PPJANO&QY\J1 Q/.ZB CS=='\]#E:^"F:G\(D>M$;'B\- .'&6QZ(+/(8M/]?7;-P
PU5+<30!>)E_7C#1P1_(!9K)-$.9^2V>*BAJ5N]7A%J.VTD![\M?(_H#R@P</+@ES
PF=DM:WSYXC7A-?,%%1ILX2-"-=(Q$$5X*(N#2T23O^ZY+N*%.UE3S;SNHZA<Q\"N
PK!*7[^''-E+J[BS0KXVQS-U5P,WB2B";SSI"3T,P(?/JHF/!LR-X.GZ].C$:["V#
P0B$DGMILI&2B<DFG GML?+$P8>@YD1K:Q(BXQQGZ*".\BB;%$,P,7#Z(U>5L%:"N
PT.1](QDP&?[0!:X)>/NIQ?]!9I$5H$C>8Y:TA,8"X__G-$&DA)3#*_.+GTFYW!I:
PD9#HNOS1L=\?>W*F4K[ C)#T,@+[>UN1%/XI2Q)C%C\S INY9@]X\P^AR7CR8C+4
PU?G/BR_K\$DM "VFH1.7/=$8,8?YW7GRE%LU7M5!PJ,V9V!/E_YN4$[I= F*5))B
PRJ4.GWI5/,2$.3M3W7)KO+5Y<4)[Z9\_2E/VIM1EI8R-62IB3$R3@';@\-%).-O-
P<5Q1@K'!"D"B^NT;V#%O&!>-@[Z+D=GD*=URR-V385^\9E]BE/FR0GN^D=4)[/LY
P_\FQ0V_K?%TK@?/L:JL@^/2\M<669;R>*E..WEBF9@>7N/XEOO=1K$P[;,Q^"X=#
P?Q@R5]=34(G(FT[^\\, NDA=#DF3-SZ*\>J_,"RI;I^.+X6):"#$:0I>XFWZKP=P
PH-785NP!HV'WV>J+FWQCZG*NAA(Z)=" $?.*,Q>/^@'&E:T_VHT8FI#9*F#9<L=I
P8Z!M^]$$N_Z@_C8+4.&C3*&\RJ:6'?LM<@(**V  ,T@8G*R]BE.J459@$_[I4DD/
P[*1_T\0QQDS9,A34@\O&:"24ZN3!B2;P33&_ZO1 A32R%1#XF\2A"TY!W7&14&MC
P%+.#]#MW>,0KPP63L/1A%@L1;WY]Q.W.W#!N9'14QT[:OR;RU7**QX%D^Y?$DH^S
PR;:LN@%4H8V_L&RDW]9"NFHGQ@.6K'TBL7BA\D/_7902P=6B<UI)\T >EYTZZPMQ
PX7D5P*P1=MTTY<:L%^Q27'SB9A[:PVT2D*2:14^]6)KI9J>L'&X^HRA(O8C07;_K
PL@:@ACC4=9?! >J>0O01]X3BA5HG-&A-@5$Y>>)P(_5"3J.@D/G8R:1Q"SHT$1=2
PDO_\@_?A?#.GMU@9504ZBH+I_/G+AO#Z59 3!@[WIRT%'0NZ/;U#P]'Q@9QRMTPP
PKS> \R^QAP\4G/R=WA?1<4P"Q9+$,^*V\YF)/\BYT[#ZBAA^&]=!8@%4V.TA^0S.
PG=]9;GJ=RSC.Z,JZ*:!Q/CX_;S -^CC<*;TX)7-]YIB:*8*"+QX2HJS/$TYJD2M!
P1)\.<^BVG-\OP^9#\B1G&_3>YNP7X/![7HSK@?S"5.6QS6\VD0Z\W.-'<&.]/:Y]
PL&6-.1007?8IQ$+2CH^:9K>#V;*#WRFR" <R=VO..75^2SR1,L$:\JU5O+1!5/GS
PL&33S2O"2!#%X,).EWCU#[3$WET]GIK_VHSCF3:$G-N5Z"XRO/DFGH?N'X2 88-P
P#8N:O82O>X9)VH3ZW:;_7=I5DIA%W^"JA+A"]I>1/@1J8U[='@B.LFVG^@ LYII]
P0\;#.JA&YL+1.)I!Z+9.C<:%MG&888<CY%LT:O"+$V[%F:(_Q3FX0<;4&V%28%N#
P!RY,:-J$,V@(KB IS=*IN*$D*6.KLFA606W^5\#N*HHP<WP2/4"[>2B(!"S-L%;!
P(!E:)>J Z:#)]%^W2!2]QSXY;!77EBO2I7$+!"...5H?NRB?[MF2%SMI.1T$A]MJ
PAEK6(,"]H]<'B6P1# &EDZB=&I_;,%KM__@\-!]:/$? &'[T,)P_2O5@C,6SMV*U
P=?;W.V3(MJ.APM>V@++O9L.[,""?=O%XH_^Q2F7I'0[ZX3G1\!M$OC(Q/$2E1&W2
P+W?)6"W'K6]2+*H6\ST&-TG;]P($)0ZK\QOZ)A(05R*8\ 4IX;.(1K@[D,PZ$ BG
P-@7X""SJB\L.GEK/Q\OPQK!53%4:$2UQX#49CX%HETZAR6RJ/!?.A]<T^3"(8HO[
PP)LQI8N8]*"2-0W&=9V#_H-Z27OK(:HFJ*IT@1THM[?VGPO+$,ZRXJ6Q*IHP.'(8
PQP^S'"A8%[L5I<.Q(X'!C-@?LND#Q0%+R4XED%'A^'L,FTB.? D1<)^5%B4$0W5%
P?V4A] # 4%>(\>E; *8M/@B?HGRB/S^5%8ZC[]D[.S](95U.?!+#_EBMR&L($=F=
P^5YC^7.Y[L,5/)5Q9RE41XE<(=/OA)Q'>TLD;".1A/;@+2N\I"53R,MD3,-#IZ"0
P2(!Q>Z/734-B0Z:E"IK&TJC-,$R Z)TMLL_2_5A+L44S/9GUGPY,B?><>2.O??@O
P23_+J^\.^MR>J_]HWCP 7I0.7+W7 N$J- ]NG*Z"76!L.5HRS>^,T3FU^4K=5^MW
P&/C2HH,9_?[6YS=7*G]]'^'0=/C)WG6!.$3U]ZW6?W4L?79IS>K4?@7B*"8_U@8 
PF3'$WL0OYTOCFI-M.[:L#V8XD8K)MQP*K\Y&R[6B/$D?I"F3'/^I5%-1-_O%.-%"
P6*P4((9-9K!!N_,%*E5[;8MXAG)O$WQDB-#&.;!PH/"?=1=J:00H7WI?<*=!ERPF
PEK;M2%("SCS\B[R2$5)<?=VYAUKHX"P-1[C^2X@#<\.&7DU%<X:F JYO(0)Z"KK 
PRB0[1L$\C2*B3F]:!&CUI P<F>Y@9K)OI[]L;3VL"^_6'RKZ= XP6W3/_"%NKX#:
PT8.1,JVH9!ZX6/SDF8PGFME76MLP)%[7-ODW 7.A+]B(W&)T@'5@O_.@J#T@_A+X
P>4B,/+A"]@3Q%)>FQO7>@AU^=]!BSODP<;,S84>(:<67+EZ[)$_RFG2$^JU>RK2(
PK>:+;6P"F&PDQV;W:EYKL8<*_.(C'*U'</;UBB)CT)E*^,X)5W:$JP7OUBF72]%<
P?TCA^H+ $3A[XHV(B>>7N)[ K)&Z@]5$LJ#7=!_0C@7PYU7O#.@UA1O\#?HOQVP$
P55;+LAS8IZ(PBS0R#2.;^L'I$U%XA[P!LQR$URUD^D6)O[!V9N>FP&<KWG*2(TZ-
PT\+)E )76O?(:,!O"8P;Q?7V!W'2:_@[6('V82HNA)<XT1CRG.IHKHNS=7\;31D8
P" -V,S80$\K7;[A&F:EW9G*N\&W2G%C'/Y30>!@)$STX3]&<!J$(@68J35 ^QW';
P#5>>8,;C)N(#\>"B/1K9/5WI__/_SQ1B@.0!-T^5GEJ;=F& P+_$:)P5"9K[:>U6
P^++XA\ \#^HP"T@>H#.P9*KF^I)G36W$46B6"NBF.6V;8'F"QW()HWB%72^^Q34A
P\P6YV\^_Y%2)C&7[E.=5"M/2]W (>:.(ADTE(<V?PH00-7(M$K"XF;BCN,>P&&Z=
PG&O7IAQ&T!NI\V!4"!5HC$F6W_WECY!8V/:KS^O:LI/9'L2-3$S\,0%S1I^*0E>-
P-#<L>V9LF$DK$ C,\X<[HL0P(Z,;H7!7'\\BU/T+Y1O!_)D-$G=/&&!9F2-55@H"
P%-4;X@<YV:-U,F79VMI/1TNH_S!&,V62/1:XK6\S[T&<A*P>,OO##]AQWYEG%W<I
PTO^6:R]>.UI!%ND$"YJ0 ]SR-<]3 ?D?5+TB>,Q5 Q/U2@#5&&C>)TO!F(T43:@S
PH55%T;ST3B9M&88:/-,-Y.0>[T>(I/V$?:JS]_2B!N=058BG552 &Z6W;V14+=&^
P_=@[>_EM&SC>'?@@]$\;LCY/2@KNP"4,7'493-DJ!6!G%I.Z6O7T<]^>^ZPP16\7
P*TRR<H3V]2#[T%EF%/VM;*V\; !>MXMAC]V>3".[( <P:Z85D \1 )&2C7#I(^A*
P7I'_C!)FI_:%&^&>FBG(4/:E&:=6AQL0G:1+/Y:*Q6!ALYL$WE5V&$_ !&0BG<9M
P<NRU/_JIVS&>-W[Q1!'BC>HQXK939(^)XJRAE!<\)"/LA ^$XT@+SE\7_\)TWI:E
PH'!7#J$49VBD.>0&^,,^GOGJ,(%$IOY7O OQ+(Y?P<,2Z$Q"BR:H1W7BG4*OR,VZ
P=4")_FE%89B8,O,6698 U5N,ZYRJH<1#.3E$$!NX*';VW"2R&O71'DJ)PV<!G:\9
PK@V!+$*9N)J'R&UQT9072+LCN.54W.T&O%IUAA>7IB17>;KV)$CQ&I\I@?]:-(. 
PZ!1][U[LKW$4P,WN^2Z28A[T\F/IW>&8QS8HN4[7 ]Z<[ @FWFLC7!GF]&(!W(0Z
P_=(RP'<5Z;L1';]0!8<2U_ 6+)&C*5MED@2%NKRA%9D0UCK_)]C>]3];!.3M]=C,
P7RD%69EO[4TWSA7!H<D!-O*<SMG''S,@]-Q4,Y%AA@,:+EWWPL/M:F9).GV"4X/N
P3B*,,XLC"6!:+%H$J@P;0_2QJ](S<80<,A<&XQQP3[-#5C#BG$LWMU5%IZ4G1$I;
PLJ&IFAP:[Y+HM$T1[&0P9T8E;#D(?UME0BD0U0<_3^:<I;E ]&5P#L%H_L)(8)K#
P_8_4B[:C< FYTLJ=Y&#.'H/8V9W+61</%48\Q'.?,K'>Z!";_^\OA2N<5U8DV<S/
P:U-][U5D:]B(;W(F&@+*9P\:+11)T=3(Q\"):L1/O]9D:@C5#C9[BD<7]PW"V> 7
PD_J[O"I(+PM<CNAO8;E/S<2K3ST3-YT=Q! ,%2.\*HR"^^T?(ANEUDQ)AU 5^;PS
PNM[1L_>7Y_G6_18)L5 >B%JA"9,"5;+> N"6\O&QFASXV+4('G8)Z_ "8;%]1Y@;
PY$AU3, M<P<B$%8J,L6NE^CSP*RJ:IE4#&%JVB!\ %G(@ *GAV=2V \25&3!Z22L
P\]Z0$"I@9E65D[/ ^4Q5=SX;FA8(T%NQD\GYE#AOL,<5KV3]%=W-='\)-=9Z88AH
P0PS^KI%M$._R[7:I4QT._$Y$G :6^1&B')_<V=F"*$G*D,\!<4:XGU[2?&[7N]=X
P1LSX*!<)*>E#)4E WBI-#Z$N<6N%<_<DR]# J:PFD,%,P,:*4'R8?L1E$8I'\VZ-
PL&3_LVTOJQ7I#JNK2'QRSZ;L?<I.9Y!.?FIWKJEW)FTC?:55HF6?;"9@-^@OV\L\
P<!$L#F*QP1$ARM300!SX]Q9(?WL94+,VXF$&$V/33KP*L5 P/N26<*MZ90; -T,M
P!NV<MR6#ES\2N_GZ.S2 UA3D8(>H]Y[NXAHPZZS_.'K20S2@+!"+=3T-G^D%2Y:B
P(0CD?2MK1:2'XLJ0^4]+E EUJJ:BVX?>P;3Z *]9G[8K]W)_B@LJ*@^Q#-+1J?)4
PXDZN>W73+99X?]^WXX.BXDWY>V%?'1?9/![)Z3RAI,<U@$$<ZFC_G1MZ&-,I=S5!
P )T_H=L_WJO$':=D[J3Y(8GX3199%_KFA="7*V3V2,Z>G[>8!^[XA+SQ+0G(Z#K)
PI"UEV7-M-O)=Y5]>X):\Q(NU#%Z7[GE)GU.%?7D OUF1?L\6)%<R+O?W#HY,9T;1
P9PA2Q6*&:W)**GP,^V7,LH>HMZ<\9X=YA-!WM7/< <JTGK&ZV9<L;(T14PH]MP_K
P?WTA]+#5,6,\4,:_=Y<KZH>N@5UNA%Z?\K6)VJ48YT2OA1'_F-;C);;_'2WF.0Y-
PF!WU8<HP Y((7P.V^ W\IF_X=\E\!/UQZ^5%TLW39NOY1I2:K4^69S<E92A9?M."
P&FUO2B(L,>A!+=ADNH*=T5BK&CUW(1\=M3P[-P@-G:Q[OG25F8Y$DI=:(=7SSZ2&
P#8)&\ES%_L<Q3667%UXK(<)QSQ]93T76&OE=T@/O9W*Z(5"R_3V>.]Q.F7MZ26C1
P/$E( F>:CF?(VM[K^>L:0XW5DD$7\]WVHFD$+^=YU2FZHN&YT-@+?;B"3R>;IK!?
P_J>_S/>QPR*O-/9Y,S#U7_"W+&#[[%GE+D(F8B"Y0(QAH!RFT#@"]VC'3,JM4J%#
P.@80%YB+)''TCT'[?,KZH985SQH?L+U6L&V57B[546%?N^"/Z,%3JIJ(1DWQQ%Q#
P$=KAI=Z'2!]S%Q=(EF:[UIGWY5W7WOM">L";F_# =Y3[.3'!U>UWXOS=Y#6#*CE+
P8'D0BT6+P#5="2.S<,Z7NE$YSJ?J\/WXV[=<2T5U:=MH-<B&UGEF[^'3 )X);PFT
PPT_2K+T/EGZAWOK)J1NMA)X^NOTD\RP[)Y<3MH,'Q+=$J0/)1"Q<) 1%3%J&47BN
P5GN^JE0[XZS#PRJTF%^?9R*7F48%36)[MW1M^.<4?N%M@?8A\0,2"S2SNM4-V.NT
P$>)4+^D@/9*SR 6?,4\79+Z9DB>^AK\SU;[=4)]9.RR5%0AS^'/\;\%&9O'UJUM"
P?S]<)*[$+U+\7[:N#?TQE6'/M@C#68]"[<VV!NGA\\@NY<*E\!026[S*!OAYF#>&
PWA36BJ6J[;KH*@EZB9% G;)?TYG1JA.-$'7IFA?A^JRB<"!F-5B_=E2"2-U<@\<F
P_<50'[L)XV.4.&1;?F>H#DZX/A="6S1D>/>JTEG;G5"W\HYX;#XM# "&(&P?D?XF
P/-%85/SN-;S^>%)IB)3;DIF\+F-/T?=@+DUY)Z?!I,^.3QN3:=(Q9ZP,"][23 !T
PKNJ,\'W= KZ7./N/2U9US^1 M/"W,H%MMI#@64 FL4SG20"MK6SL7@SB+QELY#TT
P-_A8 C:R^\GN_=^=)*Q'DY__K<SJV8V?.\'?.(U6WVP\XH?9(?9 *X A*T3W#@<K
P-3A:JP'2D N-H%BH9ZU@ 5\SO%#MUS_$N?XE -PJZ[_$K',0E!EE4.L\^=%'&?_&
P>1SZNU#X,M[6@BN>S].+.CFWQQ8,LFV-UQY@-N1&6H]%6R2O^Q[\+]0<M8K^60W<
PPRENR4GF*GNWT99KSWAFW3<E%*SEF*GN8\-[_*19H\:3F_]42GR>Y$L0U,D[V\_:
P7,0=[:/_?I+_T&I5#_;'(7RF<9G6A4;K6 KN P(F0#RD\'=%K-N1.=R?)?]3Q' 2
P,Y/:"UUXK,>1":+S^9[#&?4T@UTO)8ISVMX'H(R?W+U\+XW2M7DWRZAH[D!N%.J^
PF_P'\F# K9[1SY4CMF6&X6@903UMWHK-@'<7+G"7X9S@CCOI@G\P8[#')7>G82.)
PN4#K25W%N!^]L1O4+7N3H1)%K[+JD3;$J HJC-5WY!&'3=K8ES*^)%3E!R$5Z_VY
P8FK';"H/G&S'/H/A#=B&Y0)&LQ(D5/4\K;Y@#U%\.!#HOGM%:)EIT%Q"'VB&@5^5
PO5<ID[G,3A*>V(U&PK1G3W16M8=-$G QO=NX,()(I]7(CBD0@'RW+TH4QCH* 2Y]
P5-;8MO>U>81W]\!'($\FM2)D]0-_YL?X+5AI9%$;Y8FV)^3C21(.?4#S<A0&N]S*
P,-2#D&N=T3=QCVH#SM5.Z@N@2:(.;#(: D5!K<&NWI)JW J9?R]AH&[)FF$CH,N!
PK-(0N'-V])=FE]9%$=)EVE''DJQ".J4?KPS^>NU>L,2@AO]:I-@/N$ #K_>)I?(-
PHLKCG1@KO*/:Z''FK)@7'/7MMX@@RF^>NR*,%1K7VF- 9#8MSOM=;J22,J!7>_;V
PU&4P:;N<69"X!"<=UZC"Q>.H;'[MW6='!ZKC2+J;17'8?6SV)_F?N9Y226G>='3U
P-%=DX_\3"8."Z;/2'EN$;8EO*PW&V@7%^7*ESN4O U#7K/3B+F]1=573+O#M"Z$T
P!DBLZHI,9AZP7UC5PO8!6>SP,G&"A/D<D@QRHUHR6V9['-@MR5SY<$!/$5-U<SOB
P595\W<4_X7K9VCP[VY%A2J0B4ZJ1>226,&R!6/].U=&++B*;TB_IM=B!/+1W62G&
PC@6-;*<2+5ENO2X628:L$M<!,=R5,'#^>O\V41%\HZ )M\-M&VNZ"UYE +32 +S=
P *(2JL$>)"+EQL9C8L]YP\4&W7!YO'T3LXK%TSH+HDO!5L/[Y-)2J2/YMWQ,+!HO
PB:7N-2::_N*RRC^".5_BO?$//'Z/95[6=NL;T]!NHWAJ?A24<6#Z,:3O3<C?GZR!
PAB-S,$=HJ,"K9H;&9B[;&C4L#EQW'*<Z7%!2#3WNEQ\^,2R[;&:'MR13X,M\KD5J
PP628;-]<%$A'Y*JPGCY7/U>_F3#%P'\# +'I@<"T'+M!]6"KX]]/:]Z7DG+WP>)4
P>B8)S<+&(KI"D"$IT%G1]"XUL@A\;$H('V;EYQ924EXI>:<9XU%!VKM'LQXJQ3#:
PIZ[B+I+US8S];+5H**1DB%8NI*9UZ^](K4EK[9/PNW+\!GS9:WEJ!>-H:/XW:E 9
P>/19H@S?7;/*O7AP)(C[PX03^@;T#5#6OW86\X';X1\!X_YI B7W_5LF77](AII.
PD"6B."T@>PC4A8I#(WO0C#H:+5Z,,\V8_\RC%":\& ((;';3@/^SLQ?65&><>A<%
PU<S=S@G1]M8;Z3T]7TYI#L;S!0^.H=IISMMS7.UI\$U[GH?=-'.I%@-2JLB'#B$'
P[\;2J5_V%<)XQM JS0<R+5(HN(SV78C=^SY:/O4FHSJE0V)A!,B=&<#*A,.!T=_#
P5. (IV_R!*R;N(CASQD-O?4C2./SWHS\@1VY=JC?%2O[<"D=P[AC5\QY#BM.L#&2
P';XC*\^)MC[]#A\K<YQQ]GKD,.Q2'O.JSOKN0/?WN?"[P5I '.L$FP<9=6Y^!"?O
P  #Q35S=-N-0 %^)FJN155W>B[0(:PPOA1* YH"XCM46GPF(3P$O[X.QRI3CJKP*
P7Z5HB[)L)XQ\68F55P, ZNAH(@>"JPKRO!1"=]B<9=$C[>-G2+%/CM*GK3@-9586
PD'NJ6&'PSKCIYA/N*QTB/O"-F2QZW6HU&!\U2LNV+GG6Q'0(5X/[2DGGP>5W"$]O
P<QQFK[1E5HKRSP4L\9P-M+4:O%]P]4R&!LXR6%%K/=A,A>IQH9*L_&1-Z. +JGA,
PL0G'$.$$4S&(@[*(=Y(<^!^_U>![X] L@&, V*'/HK*F[PY'TXEB .@7*9O.0"  
P5@BP%Q*P^0D!2 'ZHTW?<:$@4\D'^2U\1^1L2B]Z$JDP&F<SXGQ26_$YS=0=0<N3
PQ^3.U^TFKL,,S^FWY5Z68=$ A:Q5M.U7F)2_H_#4S*VE,J^Z?Y(?Z(7A;,RW [RH
P8"(]S/"@4##)P[&#OV_J1+P(VY9J ;--KYV$N]F@I%+F/9U<43+WIN5HSJER^)MI
P[0BQ) PGD3-E0S39R*XDPB$-6+.$-?VLOOM ,.% ;O>K?'>N_BF.$/\5V\]VM#"0
P^1T2A=P]%5YT5]&,GX> +A+]U91(P-7)\ ; 1?@:U;Q7N TI[BPEP:M8J!G=SH@5
P)ZY#]GW>,J#?"K%I"LS7".?8UOS>I=;#SV_72=T-TE[/<%9S9A=0OJ-3G6%^>24U
PWF8<>5$AWI&P6%K>;2<&D40F*.H#GIOSG@S9(,)T'/&9)58?[]M4KVE#9^'Q^@2[
P^AA4(LD8_9&1CA,B9WO_9MQO-L(/+G> -^]NT,]'2L"]_0%;MWY#4'+^(WG2?A\Q
P)R<M8'U0S<JDWS1G*%.]KP/I' /"\-3W_U;YO)T&$@9T"=/SBO7#;#V7B6Q:16Y1
PY,U&9G<'4:G[2JMT/?\2/*5QI<%?P/4,EJG'80&I_&'2O_D82PE&"V]<]9WKM\KT
PT:C'AGBW:Y%Q[T@&'K-*MF4^=E%Y5\J+>N6A*-HD'=BLH=UPG>6LCK B>.-PRT9V
PXK N=@44S$<8.MSZI<ZTM1W&MB(MD[H.X^9F"6CXRU<5LT9\8]=#N1B#!Y=>B:]S
P@M<%6?3@:H,6*I#'J\FG:*F&)='4W9+"UX>OGJ-Z>;HU'9-@)3]AVO Y[E-\AU>U
PNL%G8Q$*$C.ES6&H!']58&DJG/_8N]H8JFEU4\78%^V2I_(/K6"2*+E&VUDD8X*-
P J2/,P[5 2B7=*LO#BQ;/\T#PA7DT6EYX<?I"3IMH.JZT9(Z%6?JO+>=XQ'M@;7]
P"L2CRYII7HFTS/I:X,W,ZBU+05\'5@#DNDZ''J^5@)2'BSG%-X.V6A5Z+49I5P#P
PLZ61Y'$1,N5RH$T>[%0CTV,Y[QW>II?4E6$8&_B,UOPCE%(%!R]E*!P(]PY*OFF]
PH^%)@G=,) P4*:;^%4K8^F!<<&>C,4$&RXR*H3D9?3@Y8GY$?[T\=M1M,049-=,,
P9"N<)T0V;#A\=5Q-4KJY494!&_1FFG4U"B5.;BMA=X(\'1 *C(3 NK5YWT\SXG0;
PZ<_='5#_,).Q."%U0M&WL%8X'K+"B$C8+<0@5 VU\KE.7.,.>A'1#8<L^7;DWR!Y
PQQ13,;'V\&>C265(X*KT@C17[$RQ9E!M8FM.>XLBU\<;$DK%O:H)399Z 4\TK_@T
P3T^8W5/-,T"2^+9BY?\.A2&'&((2ER@\"&^EGI=H]Y8$;)0%SO",FR/.)"+9:+^?
PX+BMHW&]U"/6I[P<P-.]YR2=N=)5)"GY'QK=4C*EH^5 876/AW*4\OY<L$"\+\@F
P.25(HC8<>RMA'F9 F\81F^<+N0G0 $8=05>NLSX'7?-N' <J! =XZHO/0Z9+]J\0
PW].G=]M[6%:YH'> V_!;=#,>N_%L2)%ZKS/L?1!5:^?R9?Q3$@9C;26XIJ1KM!"L
P>YF[^>[7VNLP['$/+V>;!WUU?H3]D@-#7:/RW\7J^AV]L4Q@XA.+-8^"I+P>KU8*
P>$D$>/%IW(*1</N<+IRA-NF!NEED%ST7194YT,3=B1T23$EM1_A47(_85VM@/*?%
PG/4[+.?^H&)&!,IIBR901>)LJ)_<ZZ04!# X>H$-)46<D]'6V_W#4=*=N.2"Q-VZ
P6XK%DIV\I9Z]\<K"FH9W+\G:S:^1@ZG@TI9"#8PV-WR%!]X;0@6JND,G\EN]I8:C
PK Z?GD_1QDDW>OXS>4CB((7\0N(W$]K4NU\HQ$76/7=14RM:<8?OE8B9-$TY78)-
P:[>_'H*TOJ=WPJ\ W@3N"[XF!/F>.+<[/8\H^)(<OU&@OG#X#7ZZ?%YRB,F[39/V
P-_NK8]@_HK?(PEV;;B>2/ZKOP#I_XS<$WO(5 >D8X,?37MS[W Q-.N'E,CA);+A1
P+\+#MA3+R&B)N_\>I+\^4X9 _&IR5XI69&&MT9B*:FY\7O)<;6MDY@B\=:0-,L$S
P.E-0B*HI(^,M13B731D15&8$]D9NR9[DSDV:1Z;(%K[V4/+U8_O_8[HRL7(K^N2U
PX@4FL7<TG?<8S!RF9J2WJ@8AA$B&LF=G95F9%:' .T&\(U/N>L! U[V9D7)3Z,<Z
P<HVOJ$5<@K?0@J<L-'$P]D_0Y<)2%#[;X1CNV-WRS^FA/<.%DUL_=RS,L1FD=H5M
PNXM0[/TOULT)6NP5(PA)OE+.S"U@ 5+.8><$@RV*3K\<G,>+P7'4-6]ZGMP).Q^N
PG6FC/YTEJF=O' I"MA&D,9'> R^IH&]:XWFB@E9W>CTC;;S>OC)1.MB!A%J^N)Q3
PJ:LN!B9C=((KF:;+EL:")[5:0_$Z3SYBT+KF]RG(@Y:D'[:UI_KBE%)<5AFW?!Y#
PFULH8XE7,,_J^!1VN"81F/WO(96-(#")'1 75I&I(4W!]Q&A\',RUZ;S-KWI*ZOO
P1%&4">ZF>HB[E_?D$<:1FD[OR4E4.<0#UJG:'#4$D2I" B(?%*6)MC62,;&,KFRC
P[>\A4+;4LE7#(;VB8#=3CBL^32A.B<::OZD*7[U:8;'"I^;DV,]]!I4G*3''GE$V
P0[L$SI7X\7XN?C'O)?ZTCU+.A2Y6^AMV.%B6!>^4B^]7&5Q4!$Z%B QPFM7@V7FF
P0Q)4]1EXW2I(F>G#,X+Q)[585*:;W7,DUE0)K@/ZXE&W!G'Y[YJ'76N*7BX6W09#
P73TI9B##PB@V&SU^PP2K9PDG4TTH[&"G(L><>7*UX43L\7@-?TV^;E>71J0D.^35
PWGOZL15.6?E,7=)[Z3#!FRZVHL;0^*1=1&>8]@,C9T0:L6D]QGU!)F@CWM?1&MZ"
PT,QU"M4+/C@P%)TST+.E] V%P*( 1Q>UZ[<;YWHW/$0"T8OA.O!@E3G:>I;ASOF+
P&;,)0KW4--8<(:+I@%2).7+LCHG61+#3*:AN -M.K!DRYNWCE7%N-#DP+"]00^MP
P$DQC+#?M,*E\5W_/HZ+T3"]E38-L19!!AK2TW@+CSLH.QQ;K=MFO$@'R12Z3',EW
PB[KS&GXM*_> L%0V=I8S$[\<?[?6]3HBEVO4);-7KOL S=H4CF6G&R@PV$1@KKZA
P2$&Y+!*?(A$*F@,1VY6;8:1Z>6+ J4Z)HDTS#64AU[%9 H%O#*.-K=/!"_(#3!#Y
PT*>%'5JH]' C"W*89%&YF4C?N 9:%SE:J3,0JT[[-;T\*I5<.&I5.:8=T<^#&1Q]
P8B/,JX'U^[WB:&Q"AT-81)JQH+>]">UTDYF1/))(4J8OC++L=^]]IK 4YZ\*CXF0
PI$#COK"/L&,M+WGZ-)/7.76$V7,N14X\X#1*4/JO5AU]^C"U,FLM]"3<S4+'Q"CL
PV^RJ\Q6:Z*1:XA:U4>V2N-2@*8E.-FO5!#BK!R_J_C,K6[TL^$]9MBS+RD..-RNO
PE7UU#WJ('?80?_54ILZKR\ UJ:QS3YDA6.DT?AICPR0=JY->.*")H"B0(R6^&/I'
PP@22XMEB9\9;-ZB&U)C *?KZ#?8_LO=K80FA/]U9E&-<3',7-!]+;^HVEF./&,:0
PG^9 ]0JIMW8 T^T-OB#&S3^:URNBS#J)X3TGUV.\R\@!8O]0@B'%3 4+;S!/0 U=
P(B0%Z7W0FD@(FI"3#]<YUJ#_M&4'RR.&X.;2(-Z/V'T'3LI@)M?HOBK5'MNI7L'H
P>F3&%9IZ09SI$['5 B KMY<:BD;*T<)+0,V0(F)GK9\R5 /ACV-S)96T\YM)7?*D
P_&Z,WWV>N\?02P=D2W.='R-'2^[#Z]57(UJ(T?U'SK^FK';6,3ZABX(0YU-JLUGJ
P+GUE&-X:-BL9;FRT/]'T"#G8@Q3.<4/R9V\/S_UC5 L-<T 4$+3<_@:#3UCB!,3J
P;-!O P40GC_(E(!N-ABG7[#O!RWH]_8X 0;0R"QT]8T/$&.*_&D"=70?NKY(8>S>
P!<T1C)I>C8/E+H@,7F6L"T\8W\+I%@LZZV$B_2P\I$V<&?9%!=:P^1K3SG@]5=LI
PH(8X^HLX?S8?/^.:H&B7;$Q'*DCE(.?#DG3I[E<_';])37#(V(^Y+G<#(2KF042K
P&'%SN6$R.UANJQ=.PPZZQ.R(+LK[%:8/8&:!T3?4$WQKG,"CKU(3SCP+XC&MJ*0#
PC9\1:@??[1=X<!M1C &R0@BX9R-@SR3P+]*^V#+?N-UQDVYFA#E$:J!E0ASVLGCV
P(>(-62#@\>A6FVUE/FL^]DDUI\))O!/BE!ZU7TY6(GS%!BH T&$R>/% #_L$UA46
PS?%K5#P,S_[#2-29[UT3?V\1[[HN0M#L4(3="V@X9L3">Z$L5IY,V?T6&:-F&8(2
P>Y5GK6!ZZSK#00E&/")4PU];>XK UU0\ A/K#S X.Z]%8S_N#W*'RR@A-ONL.UF;
P63U! ,.0 -8$=>T7Z0%!HFK?BK\S+0>T,.9*P ?<0KX0![LC[AI]?_HN;73TJ[6"
PV%J>\]JK[GX];>E2$$<QZJ/*8\!(XE"+=""*_-CC'QWBC<Y=FV2R8ZA(&T')[DI@
P9":@$AE5..BL%R'7WV)!X;-^+=2Q>V_QA>.)2.$>)AH3Y;8V8WA^+/O)Q/)9;>A5
PE+=4H,W#!&5-P/..(?')/(2HTR_7SKAH$-A_ZDO(Z=V LU5%59RB;!PRNI[]L$>]
P"YCA<B":B+!?Y[MSL7K-L".#XB)"AJW7;$T95WNU1*M@==;DYD;S0SEZRB2^+%+U
PI.9*H!/>=&]!%;R?V\*132M9_JD8>5*G\?C7P>IJ5*,A>?..UT"A8+GNA:1!A'_[
PY17,FNE:,3!@Y0>Z>8"RVZ96@:(_=Z\Y.1>>)D \@M#W?H$/T/@HV#ZM_H=EBZYW
P!!J!+'7YV3 [*6-GR!(W=*XY*QAKIH-&X&C,-0]ON_!P=P/GUH'D)NO_@&8>  @V
PT*-EZRIU_M+S">H<("U:"Y,OF5YYHRS;R&9?F_QZ4*U"ZEE)<)_TI*^C J/773WA
P36V)5^:H?"5Z=B@C/([T28,)QQ$-H&=)MK+1Q]M2.^R>/6C61#XN;WSG=$^[XNK1
PG9RI^G[&ASD$*V6[TKX'ETE*C-[7LXQ53U=Z:FE'3J"?E]H@DU1.H[&RRIE';8ZJ
PUYQ_CV0*J%Z0G-(\"?I5)5^:][CTVO-3-UD]P %]"LGJ?GXL&L% GG#/,+)9/%N2
P[AU. K5=(A0Z^&<6'NH\G%1;;6A:YI/0<W;!O) 6M.P\X=^Y;;P#-9*L4N-L,U4)
PO<-F&WO(<D (.O<N\@J<4Z'Z5Z9*CPV4HW>AUW8Y:L9T[K9+!S?@*#PM%8_OS(1J
P.KA<M^)&D !J^=B4.RA*L$EBG*;'1?O?.\,NB:. CI3MZMUR E-*R9():3CG[)P.
P^K3;AH=1__[$\XCC;K]IC-K1<>@792'H DXEZ\*YP[[+M%^JG]MKWDGN.S5]R>^O
P'Y1,W.[TZB>^V:=VM-%%QY5D"-@'ZMK'^B7&MK\G?P"K3I1@8Q0  '-(&:#BU$(Z
PK9/Y<\+-N%,47L; @>YW6*0++:F<9KL&1'8<TZ F=07Z(X\/ 2S)^R+ERH>P(UMH
PA* \]5?\%K7BAWY13-N[/#;$@X+#EF"6Z CAS<]#FG;&^1,"@'$OS5'!"=VFJ"&4
PR&Q'M#"Q?A8](77%?(S*B!PYJ]#HA4W.K]PYG<UM;&,CJ?"]&TA&SPF?^^IWH;-1
PGOVQH-J$!6LR#K"(?<;J2@;O:TCE+2B@M@X34O>-+:%.5EJJ00&HYSKX<"ZK7FRA
P[NKQXT3(%$C+>S*;90"5MIMD+I*$ 3;_N#D'B;NWMCE"HTXZ=E66+LZ1ELDH"O\P
P8GEPS;U]Y4F3 >IAC1SCC"H4MN-'#!G(\TAW$">3]]XN=PN8+R#[/+Y13*GIC3*!
P\%&T?7KE6'[GOO@VH'LI_$.1!4!EWY=EA\.6G <71)HZ/O/XB;D)SC=X@FD3W_-\
PIXK#:^ 1LT:J?BVM$Q3AZ)/EY(\K%KE49 &PND 1S>69#?(.'RF$9+$#FX3A41<3
PFWJO@.5L->SP?GD<C+FHF9:/[YM_B"KR_3T,G?&][IRIXU /!2A"4ZDQL\(U!'B"
PVRKQ,B)I69AZ7W7HVN8*RNY\.Y^X/AAXUK_JPXKN"-A#)I&B[E+UGC5-_#F/]1X 
P-^C&[(C-ZB?;'U"P_BX]N"PF;3U-J[(BK(MS:E<[R/G&RFN&KLH>-!2";H5$23X5
P%(TGLY>C@_T,2R/Y_2+;BW"=ZE8&J9GE/EKNL%*N08T1&K _I.(,@\_0T^^OWQ+'
PCVU ,1RM!DV.?S>NUAVJ V]*F@[C%: =4-&I8"J #FL;POUB;!CA&P/[*.E9/G$W
PQF9ZV]?N@_%,7&XPTM0P7]6I]+#2U(HNH/,C35@-*V*ZQQH?Y%$X+[_;J0I6$7WD
P@ E:LA$+Z8^^O1TC>\+"%/I!V;=,CL=Q9G93%LF#.;EAQ_TO\UD!_<D!T+ NO:#G
PQDO-RBY1^RP94TN'<Y-?6Q^$X3ZC(^ YD@Y_E[^D4(R!7 V$?M 3]GB3%MH_R:*"
P?K'*9R43U:?,FOSU<RV?"=F6R*7^[#-C#1<;EU,*[ARK:YE$000 HGHWOZ514.-0
P#:&"UE9PQQQ^&)TC$-P:K./-JUN4[I-WFH_F@HM-KR1_,@#<DE1FY+3EV\3LN)&@
P?Z%BD4 /KD+3("UCDR83'5S^K]V%Q *<B\H(>&/G)E"C$"[&7QO;,TEMV&$Q;E5\
P!XDVJOBS!WR/'MTI1(03*)K*92Z1"P4=1?3!.'_QR &#\O5R-!ZK4I(8P$V?V>IX
PHR8T;X'$:B%5@@$9,$I4H(B++SQJ -D0SI^OZ6B,VKR/#P;"A#K3Y5'%3IL3^B4*
P"J@K6G.\"E*@='BCXE$4#@S-=V)!_/-J*)_#;;TRN .L%!HB0R6J+#>%4,0H?63^
P:O_&_]MQ!FVT7EHQQFWN__H!]W@U'+GE(0F.8#L&TK523S2];G/ML:CUS$OT4-P6
PCW#F@'V+.=(#W8#RUNHB-YH#^^X+1?2/ASMB]#ZT: @R036AD>?$;@PHL#)^4&[3
P\VSL-L6M1517S "H\ D;VG) J2C)TRH# C&TJJ-M%_KO6LJNX%;(QH#(7&1CB#^&
PDP,T""3@5Q3C9MVZLJ(]D$315#ELZWSCSUX='^\4G^R,-:)V3?1[HCY:8(S)LI2;
P]=5;#,4DA3!5XI(*L[:@:$#$">;H1D]SO?QX?SO"29?/GWL3QZ).$&9LN>-1/9\L
P^6)2V7K/@3W&:;_&Q_-,<&_MY?K=VPVVD.5@1!A[S)(PF^#=X#OMKA\JMQ@X-1!+
PW"HSE;T:M4D0[1_(;3>N^>?10/!%V$%?OR2V4I4'F. !$J2*NO[O3PY>IW[_SE\J
PD1*BM.Z4"@^8C;],:  ,  JZ9RQL@G64^I3"S!,6X7#&GD0G?\,:.I$YYJ4]Y-B)
PS?OQ078T\D8JC(/;O7C#[H._@ $F7#X?4BOU_L$N^PU_V5N2#+)@2K/C,?!<H'TY
PX&,U1T,67D\2<C-8G%#E_B12-HA0E=$,J.G1B5M6+IN?&Q?C"XN#L7IG%.=)ESV!
PH^1Y\7OV32FR[&+05L1'HU%TNY]N<_TBZ7.F1/'U/W$T<H>DJF(,NMRUW=FJIF-#
PZ.QHPS6.9627DZIUYH#V=V_T4Y\Z8OC0#N0&MX=-12P*\!#WL*FLG6%G^.N K=0D
PD!4>NS4TYG]XD(F;TH8Z[@E8"<Q6RA:!ERH)7,HA*,N1;OZ0E25#>-OVA+9FM/FD
PM&0J@+&):ABGGLSQ"(D5BWK_(3N1<90+!/:/V><T/A/WO+QTE]:S1\G3JW7'J6"1
P1I<:A/3%SUNXQ*MTQ,3L GD_*Z0J/,2KJRE/=^35]"".C$R^3I5$8;$DW $:6(,/
PO)3 UJ"7'2ZSNJT>D!X$:FBXP]/5C :Y]#\K%#D?,X?UY8G1*Z6F,C7AWL"3JABK
PBDAHI;A]\^K!WMAS')O WZVVF.7U_OEG!( #+3MZ ( YO2#0!#Q4"(\?'*2%3L%K
P)&X&,=H1FF?8I80$JT0W,P!7E "#)N[QCA #=8E[F%0RQXP $MKD=&'LCP>([1.N
PJ40/CXWC'LU2[X[YT,_^PK.12=@JCC?*ECAC]CQE33"K.:-Q@#O';M:%()X0TA%7
PVJG&]9VYFE%'7LU)ZA$RNJO7>]ZA>>B:T*!B.S91 <<9=_S1D4'<T =$U'ENA2Q9
P8<>:%=U;%'9/*9,!YOO2(1L7I4<TEG(.E_T<O4D!K<]K3VMA!BI;$5F[NIG73CA5
P(5'\,1GYDF :>\^5?4NIF\"(' \<V,KL9B9\:BSXIEQ-X#TL4-_=M/G9FW"A)&UJ
PP1H^7)T_'[I?E)+79ELL_O8L^1RD^(!BP'XEH=,LA,^2AS&&4@%&T1U;*;5H\ 4T
P,+XU8"G01?+N#G@(W601EFV4A::@D??8P8;\UKW/H'<&3JFS:2)TT\S/6,^7&5HZ
P3N>+>T*"IFY^N1W463+XS]-W-[W!1;*$+I%4R5S J]NIR#[ZS48;UHRA/PWW#'>"
P",\UI1\SO7*K,;!J$&6>7>Z:Q4@/',^"0!V<\11JU.S+B[?0G73H[X@G3HX^>HO<
P[C-+SR0SURB2)4Q#984VPN;SZ 4,"R+<$]=%_\'J[EXY_$'<@XVT(&LY:4M)0.M'
P42I$5->=%J/.>4Y76=!.T-9P;BLXS8/5XGZOS5:_;("ZJ9Y^3 VO8#?[AI+_%RE]
PC<$7F!D$QZJ,U7I+C)P^-P$RQH&CNH^WU :!S+X4\UY8XBR"W@35"CK+]Z:9H5[N
PZ4&J[W%CLLJ:A>A?=I54Q=_J0_;IO2,EG1VO4P>15<VK#&[IJC!N?.RCV;BAX !C
P_$._/UT1%'98<F84EJ@_0TDMEHPA=2V]E<GJ00)"4GF%;7&Q-O-S-&$9#%=D2BVU
P- *_\8@1+HD<R( ,V^[,[4O7;(A2/TAU<;A/:8==\]C54!W]CEFJ1SG+3>."98#W
P])WX?DYFE$!2,4JZ2ZHBQX0/SJ5\:G WV9MS])3],Y(?W[ V>/+&GX.W2-P'KO\)
PD PZ"4\VQ7((O%.(!SN\<A<3\"9J$Q/WWB[AD+QV#8T>.FS_%U[V=;]0>%G9?.I5
P3>;[EG7"J&$BM])OFIS;H^,X@QK"3C!8$:.IWF3T[/2(Z/?ZIJ\R=_)$WOM6]^12
P8RA&J$:XD88J$-I*==RZ[?;[&Y.*MESI;0V<4.*<;3KMN*G=P*VHY%#8-K<535SP
P^[$CO.5^.T!EP+/P6/>;V5>$U.BJ@YZ?7<OC/4I_<>[N*BWI.&+DK0^1CE#,UQW3
P0U'8.&;_\0KV8@@1/^Z]S1^<8+>ZR3O3.L2Z_<G16J.C00I !9U =!:_ NK%='TI
P#L2@>036U(71\@S'ME"IM]Y2+P$U"2IS.OML[.)8#86BE-;'">(6CY'='26?MR((
PPH5LA=>CTE"YH.9T8EIGPH#T0\=H?A!_CU(0@5_* N:&0\:4,-;@2\6])3JJ%YEM
P>8V,27[<X1,I]^R%WQ/\:6EN-\W@##;2]\UJ6<-L . =Q!LFI0-OI8T K[?(6!L*
P<L53CL-GA+HGY0 +<TX4H<TCZS.3/EVEZ_+'.BDF5HC[X"Y#8H!7"&\'7_0L5)AQ
PSX8HWX%_0:HO;/NA$R]M 7!3Y:I!R/_E]1GLL%,V5VSA%L4UP@T>-4J8@[XJ-+C(
P&H1;0)J($6N!6XFH+%LZ\<0343_>^V3_%%ELEH;@&;D2(&^ZC:?-TI5YO0MG=PP4
PXII0"N6E,(&?&\),Z A;9ZN\.V)=TQI%1N35U*MI72\;2YEY_C1V0U,WA6!%U.A'
PT15U)[5*YS8N4+9@V .CP1XMN719?=^N<G^)9P]WB3==!2G;CO\X[\(^/9 A,TTF
PG;V(/?=!X#^9P8CVIH]VGH,K^)V4G4![-8Q_I_'9X]N VV2#L],_MVXPX+U,1#]=
P=.\9/-#RK7ZNSXUY2_P< U>1^ %MNDWN @X4Y\":EC5)D^JU_](CM^?\[\%%ZNY/
P5L@9I,X?[I=2=Q+EIIRH%'X+3^&=_?$W=58BZ<LE KYIX86<U.DK=TP2HIZL_<WC
PG)>O&'R$IM[F+P8SFK$#B?\']]N\W+DT'KP'"AE-[2L(*</D1_2L6D'!5?9P"8"Q
P)9G&"]U]&Y.2W+71D4HW0B!.#U['OJG7"-@)/7?&A$POF4(2GK>L(,90,^W6J,K?
PNMS "2?'UMU1X,6Q)2P,6:<+0RVV9:5)A9T7(1]\7W_^&)?2=7.7HH)< XBUX&;/
P_U* #+Y,XYK#Y]JCYI=L1%!D:I1^P-:G<W:S__QJWX!EOD?CPN4Y!]BWNMB3B&LG
P35Q$)+I#?3]88['M7A^!WQ1S+W*RZ=+=?&G4U#T&T!MHT5< Z<L(!@LB=<[)JG[N
PN$86B^L!W;@J*RH@G32Q2M%97K.;N4C@M^3H*G\]D$U;AO.8@SAA!70$:XP)2IQ*
P!KT/6S75]2WQWBRKH&Z<!=+-:^F3OQ?7P&A'D!T75>?U8HX"@PZF&$PK$\TTA=54
PN*-S&Q FH0#<F3G<_S<&(GUA A6O_XB!-FE1Y&(:P<?NFM*.T>ZE/2 9VPH%N)>F
P ,)JCI3J:B#NM6*K/O[T@V?%,&&SU<X.IVD8$[!08PQLZR >M=M#&1[:^FT8K[#.
PE]OOKQ%* 6M@2SA#!P_@2P-LI]7&>=!KIY=G&E],=&D PP0V>?OK@0T&%A5G<MS4
PJDH+>-@&)QU%4$2WVB46/!-Z*)]GMZG8(!#I<[-W$Z'@JB#1<N"X4*%$52=XW;UT
PWC$?11,]X/92\[W^*4%2Z]E\; 0[V%'J&UXAWD!EUCWV-=*1!68@_/N:@Z7G9KFL
P^7#WP9!*I_F#T7LE E@.>-^5)5LK=7)8H6O ;0:4Q8NV7347)$.(XW&S[0M#JU^>
PN2;M62#SW=?656]0OI&'P+3XTTG<F*4U; 2T]"9$;*0^A6XE-[N!M XFMFH(NMJH
PYC*&PAYFM,IKX8@< P#Z+6TSZ_8"/>?JMO<18_AJ-?DUD#&&K&9D-47LE:E]4)J(
PS3^I^Y;STX:/LO$89UVW.1(4!H=2Z-36_X$^V[S)!Y:O@N>DXZ10L%9.DZV/6E>>
P@,8OJ(7E^F?;KNXDW6K?O?_6]^X.I/="/$XH"()?'96?.AN*ZSK,:$)X6^>A='I4
PP:Y $.=OB(6,[;/E-]@?6IU?@BXF50+C.2K=3+TSAM_U%%^@&4L,%Z#RF2A?/L&"
PQ)MDT4QEAVFK85\$\/,_G)2^FWTZ!3 AJ":W\G3T_CF/D2E+15.]&'YL^QU>:\+0
PYEK3OJ$]7FO ':9+#MJD*%=EX#YBI 8.DP_OI3Z=^1DCLRT%HAV\$=8$:*.L\*3C
PM$5VQO/W! RWON]3V$VZ#\AUDMOVB:!-7";HP _3ELH@<G+.R7L\F_L0*0A&F!-8
P6=B,AGF$WK[LN(V9J$Z]6T<Y>N!F%BS)1:-E9GUEM9.,<<>=2N#U0^&Q63+'(M'N
PL[ZB(VY2 3?TOM5'XWK[X'J<R1 =!-^G";AYG05L*76S9,Y:"7E3-@]WA9U,!D0Y
P%9'8[U'4\4!'I6?XT-#?\7O9P_6?@-XY37*#>+1AR+3#+]TS/M.#A29+,4#_-81N
P.;*F(=6X>,[/_R<=ZD/*%<YT?0T(+R&!]4;'M&1/^)O #2/!P;^X.*RSD"GV2'YD
PK<C$F N&A(&10 "+%3?61<8:YR!QGQIKO]:1^):%[][P*Y=<=LPBC2/G K<,J OM
P!OK%0*X31@90YRBPR[?ND$\B&7<! XIVM4H.\<"_[0??HC=3?/T&X+4-VW3-5Q1!
PFZEATJN&Q# +FA%^>M(RR_2'5[?[@3"'%R[?OT5$Q%.@+7RE'-[H,:+3/V8TDC(U
P0M3L'D\F%U0XY.IY15TM1TA<85@D@/('@JPO"_=8VQ=,WW6U>=J-T'/D"I'(G%8S
P56Z;HT.TNX/BK!0J2(BOX 39Z4?3P8/T'8D-J4582U+E+5B[G:WVQ(C>@.O*5(N 
P#Z&P.A*-M\&VB*67B[;S_Q4.QOP DV=6H';%SKAJLI4.9[1^@Y;(JVZBLGXV@3U 
PM/1-Y! 3[)@?G5.S"30@[N0!?TK@3^192R"_,>S-#R'\%(XM2R,GI7M.Q-:EH^R)
PT]D[+HH,'+9;\?$K;9.ULX2_N>KJ6H"^6QNY*NMZ "G9KKBF%2]V?_73.QYM.E(F
P5MCP^S_@8I#P2#D*Q(BKK<#U*.\\O(,D#LQ@_==&,K*C>^#15$MI*Q5HQ5#"3G$"
P."T ?JE!>>[/XJ=\ZCLU*8/]U0P2R(Y=E_KM*9HVWM5\K[+L 6DNIQ6L?;?F7NO:
P.]C%M,)H1HN9Y%D''%C2)O['^,T"CTM=?]^8U34OGJP^L?Y0#H='Q^F"R:;2D1L(
P,'6+-O9-FOPCX_LQ@!H;TU[ 835NH/$:!@;.2 4*/R=N-<)Y/0OCD8OUL&C].= 8
P,2.J&% 9U[F0C[.DU%+5J<37U%3X<U*/:<(5^S>A:A)ZM\9E)J^JRH#J]? B#%U<
PR1VFN_;YYCN!;?LS62*>-LB^F2HL@-:XYWCK1;TK\PMYB)3'GCFAAKMVHVL=(QP+
P$R4H9Z<= "KJ&0TLY4N-)W)5L*3!6&?!+174&>0G@=\HX\3QFKZM>'^1Q]L\D1WX
PP]5VK#P9."E UE2DTU*<9.$31KXP=[$^98C?'*^)]'V=W- [%KPMC\?"[%?T43TJ
P-!!!IX-=GK"6E!0*,K0@&# Y^+T2\J2,L8G%[_<<=B\B@&A%$1TE^(:B-<?]HP%+
PAB7R@-/I*K&VI)*T%9R78,7V,;U,()KM2T2'YR,A1*YZ.=@NH]!1X:YT5,20B/4S
P?:G<\LCXXG_+1#M3(Z!E9#_\L CB\XN-%OA&%L\1!^/^[=O86TUH6L02 )O+[*T_
P!2 .O)DH*#H+6'A'C#&#^_9_H\>O]BP?P#VS9Z3CMT?-#I!K'R"^&W\FS?VMAT?D
P>U,7.1]P"M\+<?U+>?F7P6/! @^HM4-L\.#<@1H9U[=;5L0B#LY[H'V0EY3:1TT"
PR;&F"\6RYJ Q;!"&')Y'ISNWKXK,+7E:95C7ZLC2K@3"(IIR>LYSV(YPXX-+[3*;
PPWU,AR%UU\T""FFG"L%G-%YL%H.QH4R[A*'-UBOP<#L1UZHO_Y0L3-BP/-EM1K0^
PW+6X83J>U^!B8]5##ZAX/@#]:0705 X:_W$&"W<-B*)!LF3_6BN,6T$PMBIF3V,/
P8K9HPXWG6KB9%I E2L%:OH$ONCW% /M.IEM8I=G$6V''*/LF0LI]):2<2$C8X(#S
P(5Z,HC-?RG7%) U"\%9LYM*VRJS]O_Z>/[U@65U/CI3C(E?H#V^BI1$8BF",;+.I
P-4*_1++'%VI6(L0/"WA$HO;'\Q/!O'Y])RA=C\:$UNYHCCZE_\&O?79O]1H?":#Z
PZ%9B $E# X$7+(5S;XE_&9(<(,OAP8+!//&6P1V:XB85<5N^SG]!*6S;2DL^EQR[
PU2-=W*["/)CXX_Z$(]8HQ8R>E.EK.\(/N5L,%+^#T97TK!01?S#R9^G>_X J;= I
P[I(GP$28<'=0%6^\9)SA;8W A5:"R2-L=5];G%/W0$1M"/2\*:5HLV)-4AW_218'
PD^1V@6:FUGZ(KJQANC*/<-1ZS''G7W5,,NB4W:T$&$+$K&*Q Z)\;B[.0K%]H^,G
P=QWEA0FF?'^ZUQ\(@9WX2O#6<YA[\3L<0%SORLI2I80D -326N%<=:];I$4\5.L\
P78$#H->JF0OOLZ ,<W/3!'A/H-'"%0D$O0P$H/C!V73P%97I+]C#?@RPH0%L-H(H
PRT<^<)5*C(T:1))S/@$M9A*G&_ L9X"^%4#H#-<WCQ]Y0E,K33<MA3"?.-0D^HA/
PU0 2:'DJ2+64^CFQ#!J46[ZL6Y/XOXFI]%F0VHA(9G.VQ;PG@V=((91; OV7G7_L
PST0)6%K.PZSMDN3TSFMI+*O\+.^AQ=R26T+1JP7Y1:V$KGVC@ASS0,E.\\&$;W%]
PQ D>K%D"G6FO53"VPJE66,E9(XO^V?AP0YY59U)_,X?-QQ,<L4.XM4D%O8[1=MB)
P55"86FC<F@#2C%%Z!2LV45; ?35_!]R4Y$[BX7?QS,L1F7%3PGFNF8N=NN"2,UHL
P=]1S5> UQN]-V[^#;_I':$PDAIV;LJG.J;:3GPRCNU//I8=>Y*SB3AX'#&EP50.P
PUR!U0Q9PJ7I@(LAV& \0!!QZB^K<JGN.VTP(R%-FEE6GB/RL=V&T>2\1P< .?E.J
PPXY3='W0?934I-=QU>%51I@2I7<$2>A=B@D/_$R<X=O!@]X7GN:A7OWYN=0!\]MH
P2.2W;1)(3U@\/"P)ATW&X=*>)Z?R/$&XD@YA77727BDSF59YR=AW4PQ"'W@3\@:"
P-5DX3[V7@'G2V"GI4/^FV@O'DR/"@*F$5&">GHJ3,'IW6:LT')0MOBCB/W:O%W,>
PU1 0P5IYDOUNM^R#O]$&##5LWPUL+:J3^8:N%#R3"58#T.\/A ?( @(K*IK/H;4<
P#.5C"1@QC6#^8:WJ.*O5_QG[EB)P^&JM:% ?D&'D6B:*"3I272-*'D^WK/4"9^2"
P79[^6O :)4 =0Y>CT"]^\)]_L(K;^*$ \V['_A9CK/+6V!;TPLR$I ,^"B..A\RW
P9,KW23&(H:<RICP*!01]2[O8,MCIK%J"/76XF]18[B^H;_TRI&"ZS7XG(%0 IK<C
PUE!34[7286@3F/U>6'=RO^L%23H;.(UQ7<,%K C!L;Y3RJZEPY_/)QVZ$DS=@L/G
PHXVX>\=U;7BK0TL3P(IS-09XQ% 1S;?W/U(-RZ +:_0M1BE+][+_.NK,+ A&\0AU
P.%ADC) RR'C*"=EY#$,E8 S=GL'D.C'C%#:5_(8QM@@4<T7F(?B,H+[E38<DZ,>@
P/4!5M#*8_'IN,@&0<H<I[TPS+UHI&']FE.68EE)(TTO^&ZF+GB4T'4W(_?L7%E)(
P&-FT(A]P>F>(T_;P&:N[F+ -TT%(D$*2&VAO_3%JR@LNT77C'/Z,6J%\H(>=7$^"
PA_'76M[[JMGY-CQ:-W@A8#?C=6#&S/U-K^V.1UOK'8"QF)?77#Q+8[ 'S"'9[R=F
PRGC2*D,/7'&.$:E\N05S(6]7 24(,DI&G%17.E4V#R4_3UE7SNL"MS;Z9LTPYB)V
PCMQ826K2$5VT>*!(W\,$*X+D*]F>QXK<??M'JANR8NN1,GW3%GV/9J_#0UK-MGYW
P--BF5%C3LA*!;^0B"[^G75>/O73N7#''%-"5(63\ 0\)08,JEM[]P!L9DFF_X47H
P\I[6?X0 X:X[U!,.<C-Z14B+\$EM*6$@E$F5=CY&H;>==,?G\U:]JD6W*L">XK_/
P,8U\L8SK"%:'?6OI-(/22%[Q'>YQ-@#.)HXWJ%FR+(P+]ZB$F4:&3IK"3'M(CL6G
P"2]]U-*'"2-UT6+K[5QM;)D2^FVQ2I9Z-V.@Z^;*L[.^^[/"3[G%<9)L7Y&.)@2.
P\L(:7I<M:=\8VV'E@23:U\H:/1^XMXNI!L>A^DT^LY/'E"4Y_@^<QNI6 LT,"<M*
PH1PG),_L)G:;#DD<]6(1U))MUDI:^\6.)& 6HA&!_X8/ZJ=F)DXW6VBDX+2^@2(;
P%E("B27+IH:G(CJ1%J3(9?9VY:;E)]@X_:3#&=XSH7TW^:P/[9@/"0Q52M4>!DT)
P.?LJ^\YFG)Q.@RSTZE-. S3_%^.X__K_)_U"G\2;]W$[D?H("\@U #92MY1R!+ +
PI4IG;3$^/!BNSLKO&Y[WJ!9$9%>O]A:.>,.V%Z*?68\<E0'?%.0RE!6,:'MJ.B^$
P--L,-2Q557W<S&#/*BDM2IR)7Z3OT%V2*L-;INHPC5UG9BP[HO0Y!60624#WR4<Q
PF[$9>3:%Q< O&IZ1WM;J$1/A5Y/\852;W9]'RE#>B^T'!CY4.&E(Y_"BT)^. NCU
P?U-U^F)<3V)T=BZOC%BXTT2W$G;"^6.*^A)R'2"+C9W@9U_NN[8Y^LRA@AC+YF;$
PR?L;E0Q1GH<2?P,4E58<C4UM^[Z$157=RV,=.>%D3$E&"HGZ*+71)$15HA[D"OCT
P$KV6S<U#%$P!\6*1R ,4SG;LQ=? W\OU?Z!,_J_"[*(&#5'MC+\JP39U4U9]+? ?
PQ_X[CX31F,_.MQQE_4ZU4^+(#]SJLK1.F9,'7.&SP(_T@5QK#V:P%_G]DL+]*A.H
P>6^GG@V]WP/T-I*HMM'&\?($4)8:R=?<:VNBS1T]O.!E$39BXJO/E)%VXSJ8;.52
PL^/PCM*-,X?_"@/9W,(UR+A%>+TR'@IIV@THV](QF[]M+%4K+!+Y8$R_'1ZE?(:U
P'. SM3F9&>@^[ OPQ:[P#F+KRQ4G]TS[4 ?IHYRPH]3RE7C/'D+WF3B?&HZ3=K*E
P<7%-7?S!^<@44^BRTOU83FXO?J92NR"E3=AIJ<%QC/^I'/3;J=A%+6G8](V&%FH/
P[L$P81%SC9X"78T5!Q1.,GO-_C.J\Q0U8PC\BSSE-QSGQK.N<Q6'F#&7)72L"*_(
PBO6@@P0\%BX!;AM:X8B @WZ#-HD-KR11I5C9[.%%VD^NG&(X>+-[E-BE+9(E_=+O
P3KYY&\@[@*T3-ZT(#G_%'^ \MO;BR,G#LL@06,=N$;91;3P2=ZY'L<GTJ;^K\Z51
P>_EKC>O:CT6U6?A&U"E\O*IV"*J]==)8=%[*+M-,Q)0%5X1@I6@W3KHX\+$:&;/L
P>7<(CJ.,MH,BTX@A9*,)W_"Y<.V=(6&DH3IBJ@&B[M$7OBZJ>  N5(\< ZNX%IZY
PN:YA\W%]XMC_>%^HOU"E2%X)&B1:Q#.*2-IEQ-B/GAT_MZ[>S=53)%$<XK"E.K$=
P+RPOZ[55UCQG 7S ZZP%Z$.>AH):@VKA=H6!3ZW5 P-F"U2I$JUUU"I.W'NQC0=7
P7IIF*VU,^@"?7=)H2Y?O,H^I%>?;P/LJ91Q-Z<N,S:F@+M9<&E4 PHE1TU@$@M[L
P_F0;%L&'_$/D_,;1T1R5;>G2<(=WA52N,"-(\>@S4;>KE5W:?7CW)\O0@"^4_<&U
P'SVDS"(WFWG VTA5F)&)'YO :WP,6J!P_3E1(/M0HL($PW'TZ_HM,.Y% ,*M*6,J
P'()'T,10B;UL;SM[^J&')1L?6)X,G_&"X..\\BZ,N? \9)BO"2ZS40$67Y(]KA,L
P$$BUT?;LO\KCTG0FI:4;KJE#.6ZKD7 SG#G:#>M7,242;GP5LQ+=&TK8AOHHHD,W
P2P<[)8XA62U"&+D*/Z[KQ^/) KT6%9P;]883+$!.PWN)9^2'G_N^O83BK"<H.\T?
PB%B"4>]86P6:<11T\!WY3XZMU^SO9CET>H.RV^9"U6;WG3L/61QO/F^V-R0AZHXH
P0%&H%>'>IW J.N[TD?]_GV3AR;Z?M(LKS;D4*EMJP)'P0#,CTM%1^VIO(-65+"RG
P]TTD8KK:\80&'S)3DEW:+9UQ-%3DEPJ(!Q;_0;->T6'T@Y\ZP$(XF>BPC7Q=SJHC
PORKXN5LIO?*;RHB!WLUE4F;HWE)B1^&MPJ?084[JKF?;)#>6^+A6W>LNWS9Q/G 3
P<V10--$?%H],ZA&YB5_]U&I%HA'^W/J1.MA?WRMNQYF01 2Y\W#*J:"LH!-RO+^A
P]>>^I#&@C4M[% 7XY_!^&TH!L(_BQU\HR9Z;%D)G("X3(3^0V])Y$& BZ27J<R$[
P+/%.&74NV%I@4^^VATN+"A]ZD^FQQ;*=AM4&_7(1G78GM'7/1!'9+;[[I)DX-@<4
P62X=VZ(F3%BH[?D.$B$9^38R8B-/AS7T$8YC-2BTYF/3PL>(,C_D)@5?^PRJ+'<;
PP'".36V%+T@[,M<I.35PQ-<>OAWU;RCTCE<%'_@;.A<=@7B__<MZCZ&*J/Z(LUT$
P0@/GUM'^ELW.O;ZG9AU\%\SS/?(V%V8:O3Q140>R6("2G%^\6.".0:(OWU[1*PA&
P/_R3/X@6+OYD,&/07@WJYT(I?]?LS)"78-*.I8OI$*41:A&'UI/*#F"?WV4XUSC)
P.Q\[1BY7NI(ZQ:IM/X;\U@>-E]DMC1.'#$]<\!=N@Q=)W=^2KLX?1B6[S%J</LZ4
P2U*5D IV6J<8L8-;V/T5COUJ3;)E^E.Y@D&O"^!YNN%@?:VCQHK*R#RI^WE]7FPJ
P59.!IG[ X=8VS6UU7)WL?\[]6 4E&U]7>E@2N.%B@E@&J+0A9/7332\Z^TEC+PFL
P*AJY Z/KZ]0/K)1:-=UIJUI(4+!M 33D!"NW&7D'P"!FL\]S6HWWL5K#>DPJZW2$
P87YL><>=)I,<72%G'1)&H],+L4_7-LKB/$]-L=N9/5ADP"I6XNJ^9$KD)(Z71;SB
P6GSFR=$R/I\5:N8SYD.Q3AI-4-!;;AC-_R4B(]97.WM[MA.S>Y=ZPJEKAUF.'"4D
P,=+9P3/"KFH<O'==5-[8(<JL8_DI_NDFS; NJ$1%R >X& ' O@L7R=6R1Y++%6KE
P5N",>,&QT<P6QBF6_!@UVYI!\DGPVZ7"]@LC4\I[W63($85NJ6UN\.?T XBK&*M>
P#^+WB\ASK/ZLPMHJW-;QB%<X'G+T";*[;QBN3%AK&=0F0%2E?KR#'ZR=/"8$$:2S
PT9%LG:2@(6('YN]7Q3>@ANON-QLI_@=XCP<OI::IH?P;,+.V/V(>@T,:!U9HLX>C
P4,0O":,N2)<@S4N@E0(7>3N46[.7\0<OGP'&@$L5XB2J<OAC&#.I/;&SB3Q=%RAO
P^G&\#,%"0$(9KOH97/0G[6?%PP?@D>"K=)<9<.N+/%U^#E'A3ZHNI M5D25KQ M_
P%E4"M[!.5R6.&N$E)?"'3S889I1LNER?'C%]P4'5<":?<!/GP:;O;+ 4I:9QM$;'
P5]/5R+#M0%0TUR;M4_$@,YTW!3NPS!J-R6.K_Q>;N+]+K+Q,0YILO<C7MXGX2=ZB
PTL3\''_8</C^@YU][9$?M0/T^_[V+L.4G5P+^_07K43G_4M\14+?>+I47Q0?+SD#
P&GC4!/8%GHD!9I=%A2AY[P.3U1B&N6#;:;-F88C$9?((1X'F+A+%5LTUW0;2 5D;
P*)NCD6E%VJ<XC6(O  $K-?60'#4*5PO76J+U0:0G"3U(7T:(LWUX5>H@*O,8ALJR
P4%NJMT;ZH_Q2^/7TOW>'M0V:*^=F(KU+.@ ND8.966H_'M&:4>N%197\< W4(W?5
PE[7^""[LF 8VT3$52K4WE_0:N>'M'L2!MCJQ2X0>1"+91:[=[MW;=E#YI 8 U$VM
PUL^\\.I&B/Y9XT)<&2ENWMBH+*WL7KF^6\WD]N$E3,G;(@F.%$XZW:!@%=?HX>C'
P'D&MDM@WLD'#1L^M*ZYAF?G(2HR4#(F)1*E"0M0^;K;Q# %5'[_+(_]93X5:^U97
PT=C!@U+#60Q?'Q,R9F,]+C\/4!XVX2K"-+X%V3*,@%>J=6N>9U-*\F?=$>/_DU6X
P;WGUWQ$ZB:PD.;:I2BPAPIDVY 9:$SUK;^>(%52';R,&N*=Q&97H"Y#A\MUVCKN7
PT(L6K5R%HF5"A# VWIX@]']S%6%##92P^Y(B3P'8,M+ 0#0?_=&>OKM@VU3Y!.GZ
P,MTXIGH:+'Y>4%D9.(LU#H(^J!9W1RZ:#/$=(?1>"T][8T@)(;G.P$E_^%T 4!OV
P!3)=UIT<T+XKQ(O,(00IA&6;TS#)'K.*0P-F.B'SY#'C<\/[\GJ;RU+I I/I@^IY
PG@F)OV@D-@2:"EP^"NG\;\"TF8Z06)!DT4WC^=9>BO1)!^6O]]+CDOGJ@0(+]-5M
PP]@/#UK'W414[4 K\0&O A;F]O-6=B%!C#<#QSY6-C%DTI?2?*8>^LT/.8S6>*;1
PI5>OR&_1XP?V6*-JW> ;*XVJC,)0KPNP-9?4>I.,^D#4"8[=#2=4;C%QW0PB"8_R
P]@KSV;?^EF%?E(@NZ&:'^,(G*!OS-3J)>A7P'Y$A4UZOECS<1P,R='DSBWI:AF/!
PFNM=&"?&GFB1+4:I#A9Z6;1FO-@CZ"M3)P"8Q)C'#R)()A^D G%'XGA-*(GUJ=L"
P-L3'G!2$+>*+,T]BFB$/&A4<Q$A-T"&&E.]RW%^0<#W"Y!328)7GJO(&[K4,=[=V
P$A2'&R$9_^4XC!SEDK6!27TH5*6(4K\OF> +[H'[60,$W,7][*38%P>)>T]\.7:_
P=T\P%4EFNK"UNU?[B<%?;"8EU!3),6WR[-+:(5 ]>6]P4RYZ,F =&$4+>1U-4_.G
PXVE(&(BOFOS]>E,S[L60B/^/JIH09JS]?GKT)K!.3><5F')&]*>LF&AI_^2D.89O
PRG;#W1><@[S9-E?#%Z-UWSFK=GG!)<+@XWCJ@1DF4J*WYGK3CW>D+;)35>FKD@6S
P]*8G3J+ <H;TNW[1/9WXF,!CWJEU]>IW@<]'S#U(Y0!HC"_/-:=R5V6IM$%JI4*2
P+.X!4R$C?0:1/DOW2(?]_EL>T3VKFC%BN36K_WL<.F!5292FH(5WZ0[R<="D[2*W
P?D/41.;?I.^D=JY+'X"FT86ZUF0S<Z)#QNHV<3JRW.GO"P M<BB':B:\-)@BL7@5
P\$B:4I?>JL.&E.G[3LEP;"J4T=<!QK81J336<]2D\?>C6MXOO_ZRGDE>_L%K8;)<
PZ]Q[T[TJ@OP;O3+];/DS06^H=I0@Z4((LG%J^@9Q \5<92^TNO6K#7D7V&P9+VIG
PV<HZAL30 OE-=C]CZ*'G-SQ5#.4'[,:,^I2E&T#A_2W_QHW#Z1LM_D$?A*==!0A8
P5I0MY\D7"63>(06QUNK.-_\ZO.1#F.>-IOG\M8<7\8\](>-47JH+*--1P/8C8>/T
P?-_*TC-N)."LR4##?&F6/4$^GO;\S=6L%Q5+5#4TDDAO0 &CW9''>]\UKJ%>*8JY
P]MN FN'1ZWP19[XX\H/4??9-X Q&9A8=C-(1")+.?9*)7<7,XH2/PN3^26$E&0Y$
P!#3:A4^7(@3:D%S1#]&,<B_W=_7)7@RO&CSV;H,<MBU(PI ,C7375BUO&3A>K<,2
P&)?YMY6I!O-F,U*\'U7Q3J6:,Z?3+77(T_Z!BAK+:*>"F).T6U+><SW\OEE6N"*M
PD>G<>.BKNSXR%+NN$J^ZST6'3-\@\+CSNXVW[Q\[(>4P0DY"/$ZQIIJ"01)CE=>;
P5XG%9_MMU!2!'\GG1T,/3ZI4%?YPC.:)*3>9J]V1^5=]'P]3K/]20C=]#:4FX] =
P0]4BMWJ^EP6UR+2VA:UIYY10@]\.8ZPIU"8>= 8USJ=T"21B7+-9=&YUG2CB2XH]
PJ[](;(U+<$R=?;QG_DO2 JS5=;MNZ8^NA^=N*^IS(KNB>R5A/^V3IR<2^/7[K>)M
PW%C#^3F^;MNGSUQG]_A)\GEP+W0R./V7&T);50^7T'WP>)J]GL*TV6+2"(/"T=^)
PN*O 7'4HG\<)+S2I\ [V91ZM*HI+LNA;6KU:5Y)8!:].PP(:_;!NN^FZG'\[\D06
PPV5<[?L+Q0!6I48>\,6)WJ-;*O(,^#E=KGC&<*>ZD#B@)=],FY;*V #I&"!\?.1G
PI*-1LHCCE^Q;U$);EWAX Q:\/HMIL[\,2J42TP72 9,\>S'UDZ/>CAA\86W.CZ&H
P&*"J4%0H@5@Y^/:;>PS^<C580".?P?=!QGH"J,#Z"7EW$(XN?S.!OI(,P-E$$!RX
P+TCD)%4^=U0M/LXV:>EU2U:W-,WD%6UG:56P7,^5N'@^(@B\[1 IG2*,8RMW&ZR&
P*$;0I,^Q$M#HP<:6;"(DO-1NODK^BM6$KXHVU?][./>+2$*GE-G[?"0<W^8J];G9
PKIF\"/(L00Z01.0%7;$.\C7#ZC',F>EA1MKN2.(2V)KPA3V_;.V-O*NK#IZN^S)2
P4 [40PKY.1\X$?H8TD]5%5E#7Z'T'B2$1.;BDDM;M<70,AZ[WLG= 'CGP.,D,FM[
P !I0[A\H(Y7PCL@DM_&:V+R&:EL^W1AV !J"2XU"45I-'+GEI$_*V)_"M:#_?6I(
P%Q$Q"52;23L_SXG5\S*D]/T.U>J8?2DOH1]!7Z$5.GSOI--_=38,_2@3;?FN[6F$
PPS2R;,^\ QW\IG4_])O$U-P] QSVIDRA2U/??"?+,HI1J%4JK/NFCR<N9_,8QWZ9
PD_64GG A%#:M9,-@JB*U$&3]!QX&+SE 3>_GVP^BJ9E@^R9 @K$Z=BW2?\-U0#CM
P9TK-P.\Y5[HU#-.,Y_-C$ZO,N>1BUG65TQK%?.1BJ@71JS160\K&^44-S90@IK@F
PZ^79\X&_0!*&E+3-'M>OT7(?_RA H+,&!_12[#UE./'F=^X?YW8(C7&N"0H&=_![
P6,3RMN\!?;?IM0%DB5+>$5J!',$D\$55Y1>Z(=1^IHW3T\XO782%C >FI%N]&AJK
PHLVMIO,7CZ%S.]C"DU,(]&'-@JKZ^KCQPE$)JL)=F'\?85/ A"<Z^\W'CE%/ZF,8
PL!AF)WVXK CY@E=W$ 2H#%VQ<-7J_2ZL<IN'YE[C&,\E/U<1W63R)"J8%*7.J%-;
PFA&H[X$%><8:F8?STLF_M+-NC,LB6+Q-'2]IQHO1=Z8E]QUYL^8H2+X!F\8K/7A)
P5U;-.B;25M76EF_P6K<-F"QNO/<BTJ"?<\3[")A(Y$T+SW18+6U#8THBV)&CO0>N
PVKPP@>_O;NCZ2$JTFG>^GW+5]/@K!84NW?5*X50=8XAXS[Z(YP*@G'(3&L"[DPQ/
PC'[Q8 RB<P)6A/2M_UZ^AVCMN#'/KC(Y>@\?@!FOW>5W+ %VKI836*YW59+!ULQ;
PI7S3W4AM-[6D+:4U(M)J$Z)YYD+U^([<"<B^$7<9T8"9SFM#?)S+1!1QT9Q)Y>FK
PJ]_77%GBP\1W\Z6(+'-NW5_/0FV 69KQYI$&8I5NAM@\KQ3R1 03?AK8U2C"=,[Y
P5Z#OI,YVI5('8!E^JHL#BN#[>?=Y%0\IX)>#T0ZG=:MZ-:_\G8XA7E/G[ ;%,CX4
PQU)CRSB/N &.W@W./$Z'<?E8_P11CW;?K@V7W(F$F CI@^GDR:-?L7/9$<]7MR'[
PEK\W^ZSK_+*:?73,&@C:[ZM(.L1(I.T<0U1FE$U/JA%\I6%VQ(Q=OISSDCI#UL+^
PB)'YV#SK,UL5^C,'S1$7D[\SB?>+D3Q>/S!> R\?NZ)NVHB\O=?%#!-'A,*LTPN)
P5]?[AJD23K0L*I!.-Z<_E&*+/Y1[S$$YC RI<7PUI4>BI-R9&?I=0@P4$?MM \XJ
P$%D#< X/W/$K3="1#%JOUJ-MO$K_ I++>D.U>B.DJ#A&-YO//)8;]O-^N+O1Q6.L
P> B[/-].X+'':JP O^Z*)&V[#TNGC_)VU/!PGF"W.4]/YUJPAFZ)P*FV(\R1CQ)#
PM/4@]V<T?@AT>7=HGQ41G-['!_KB'8VRC;.1O$VQUJ5M %UI.\]LV;7Z_LIVOD]N
P9V![^E<ZIP.$BXJVSU35-R@M"V#/:#L-;]K_#49CK1NP]0#'KV4G AJ".9M7UD4L
P\LU4; 6,@D'0J\6BY71@OB 4:0B<T-&^P/ (>'P0&9:M-XL&)$X'\'D.:984L))@
PP5JU"G^,DY1%)/S5"$V)X)S8N/D@9*>2&2'X%)J>V)08JP?554]N2*JS3XZ\DR1$
PK4<R_)<OL\O&54;I-^:)QR7#>'#PF]FHO/4@N>VB16"_;ZGY/_%$*,(EK(4 8]0T
P_Q]$DV-?Q[-*L[%M^^NBHWJGI*V9^%@<G\$5S.%7<&?Y>?N(".AJPV-L/3PR&KTM
PE&^[GP$:2E]94A@(?Z>CU0!/GA82'!C5I)Y&[JM$B 0'#NQA9MBL9._ 71OX@A]=
P4MQXK -0NX[4+H"S'+YF>3M$0];^I#55XL159P GJ.S4X,YVNW2JQ.\6)./NO\+8
PT,=WQ\(V%J%9[(@TF%^Q:CA8'=\^*3C:D;$7$A2?1/2JIHCN'<CXP+E:GUTB:&0W
P\/U+!@4] (OQF7.L4.@5_ ;H?L?%$]]18MPLM/GU:(K,_$\F&LNIY>ASX)I)EUSN
PWZ45MW0Z:T%9D?TZ!)^*W&-@:L$LR:V?LG(@=U+CUT8Z*(,1U<7\UY_ ;T6O)/3B
PG5LI9;\ A,9D-U*,452#P^]?:\V%I3!PY&N+2$,3RLIX)4^:89!00*2 =+38:G*X
PTQEMW;N+K'6'C+'%T'@1-Y??#'2EAL+\V7;%?OOQLY+'4M$B.$S9@0XV#YC(8'YK
PVA^LEUO?0V0/(U"B)<-,K/%0N[(OGGY9&]O3_$C@/]9=#.]D+?3?M4T^A%((X?6V
P)W.D\1, B6")I=;M"!(0<?TT;O<,3:0KZ;4J-K1OP+B 6.L5),-[J;]DK*WL>73 
PSC,6OEJ=<:@)PO$*!(*'"%Q@F.#2/TLWGK.K[$LVX&?8*=Y'5; VB9AS6'#18 _R
P*M:)G5&70WH\$82]RK 1-WYHH4.<=X+4)ALY8]YY^?I\[1..FK8ASIE^RX\0=-^O
P4#]3F2&_8@!M3G->5%@E+B'37BYOS#@(>(UXLV![^:YV$"F)H2'FM%<[R5[S5YJ\
P:Y90"\51?O<)J ^=>?D:4<3AN1TL/V9 ?B!:*&E+_AP<;[]AFGJX'#$F\[52/D(M
P&+A>[:&I2G\ ]\(#L2?4*DIU\#!S?7YX!^[@Q,XYP,=D?K:9)Z87G'JF3ES/IN9L
P!2G#Z6N(H,HOIU1E!2+"XRU=!P_"Z6^D CSW@D-'6#+RQO@_!ENHQ 0R2/;0&?JC
PE?9T?%6A<[\L][Y+$WFM=CGU8;@QO ^!G^CNA\V$@P$0\)<"0;UFI!#".*VO_>0X
PCVY4VB<_BZDEP./V9\16EX;UD.SV%=K&K)])*\WEX?Q+4,7=6*F/%\NB<M'G&G;\
P/O;)X'K(%;&'FW&P0I2\.7,Q!T@@'.D-_ FO^^%&WFHY?!-9A>D&1<:JI<,,+]4E
PB+/"RN'IV:'-T\<AMD3C)!PX-\2@OODRR_$!3L"Q=F7SL^<_QN--9<:>3$N9.9.A
POK1(7KMKU#Z(SS$OI0<J MCB#7QECAYR4!Q^GF48LZ_Q"7<71@B-US+FG9D@7L':
P%C9D63N18L=JY2T>MFCL#IJJD<,N*0+0XICG^P?;*J?C23-L_-50L#C"R$?Z[=G'
P:__XIYX0Z8%R,HR%Q8W'&_N%CG3PC)(G607Q6<-6+$MF?O@R'4K\.L1A+NKQ^@.Q
P <8M#I+:5PYAU\0"A;A-&IR6XZ'<KTM8SJO79W%2OB*.0$2#T%]N:8%=ZC08 ?Y<
P607=R++*]Q;TH!,E0-F$FYH- F10!H Y71=(-]D(60#CKE'[?EII?!Y-FD%&.+\"
P+#0KB8(]_\:*P'N_H\4EA38@OLP0.H!NQ(@1@S.R.!VBG1Y3[C3#@=Y*';9X!)L1
P5S-)A=;26ZIH#9^I67:LB9CIM@%/8Z6"/):9 SG6H(AR+=+<.)B^Y=G[<$6\QTD-
P#WX[O[<V(5<=#ZA[R=!A/7V$ B>C3+@HH"WK:-DT.(,)T3N^8N>#5RKC?N)X':.P
P2E[6".#]30K+Z2G09,.?#3SA?9A7UY!5N8VLNUS[SQ%2[C+MB+=+NX&!=?87SSJ2
PX+>.IGG1 \*V<U #\[Z#KEJM*O5T8S)T*8=.#YIK/T43>]$DF%T3WP\D91(8:"_ 
PR&P_(MOJ8&ML=%<VRPI/#L(&AS3D#A7/G3(0R>;9PR[R:R^.G]OH,@>HC?5'B0YQ
PE4]3&B=9)MA"^+(;5>:B-Y)UXMHBJRNV'F K&&4:$[@,;OA;P*I&_(@8)B5EZ PC
P.'N(S-N+!1?R;:]_Y7Q_LL$;CR\VAW+>IYH@(==R+7\PD)$J7X$[3@5D%DO[Z)LI
P,@3[16HF6U>A8RH8 SR]TR4PG,X%/1O63<.N<V1KWY:\:UH= <#QXHA!GZ]W]Q)D
PU)-6YI2ZGW.&5O\22:4JZXH8!LFI21Q;;D)I5)_9YZ8MU.AW';LJ"[[W=M23YWDI
PAX.6L0REX-O"]KR."=]U#[F*PFW<"09DZ.::YU#')ZO/2[OB93%T<M,^*!( 585,
PHYD9)MM>#0<Y0(X<X'E";5R%(S<*/X&P#RJ(UT0?EU>?N&4L^$]LC8J;'^? $4LW
PVC]L]+!ITR@WZL*?^'EJ9%-2,Y+R">,$O-66>6@O7B'AX_?&EG*JTO_[YY^6+^\1
P@:!A%&6.'2.Y5\-LZ[N8A6U9.>=<XS,L9>^P?/78H*Y29/'7)2><VZA,LDG "G;R
PH\+R4'3S]*<BHO!8BIO+3G_.R16Y",SOU<_^=E+J"$\+(:RUX&@_AN&<)]K\<86+
PR?R>L3%>\@>BT%)YY1*@:*1[@+)31Q@698E%PTJTT@-9)?2Y5#8N@7-38V!G' DB
P7, RDV!6(7@%2Y!EO\1!!Q/1S4'U_F^%TB$DI,DS],+[JF')!@<A+7OFRAS398O)
P(3V9UKJ3$*>:891/R7?&T-/,&+TKYU%!S2JM;I<4=@!UVH"8,+='QTP]'2K,TP:J
PVZK4T<,BXUME\!ZJ!LKO=(A;*ET<_%.;PKB(=TJ<?LNMTZY#?@8P"-O*AP=_Q)T#
P\+;L=T E).RE5O\OT4 8:W/Q220R@>4HVZ82V8;#0)JQ=(]3-J7&JWE9S,S"4NG_
PY0Y+P%J!L*-_N%?;8XRS*V[6;N;0N"YH' LNZ)\K G-PL(?J@Y$$FR=?SM[;#%</
P7+"0V$,EKPCO!L&2U%)($''8R9.2:EV Q0.WJUMQK 6.Y6"?N,<;[=49S)W(K*AJ
PC4?%9"_'6\G[T=BDW%7-8ZO&X?7;<?PH4FHJ$/K]T5$'Z%J=#/[O0+P&@S@YP%J5
PA[<G>3Z @00  Z1K]K3[^U]]%62Z:X00!.U]_QU@(G&ER4TLSVW?+X\$A35!"_5\
P7>VIF=L;+3JH:EFFH_ZMI^ )<-*[TUHI%T0U"1NMST$^V^#4OSRH:#JO-*BBC"Q8
P&+Y7"37 :E-0? R7E[VGA?%CT%E@L0YKR.LVV.7XU_\U^&P_M;B)\Q(>.0N1[X*0
P7'Q$=DDG<>ZJ>A;):_2VQURVWYGR;$P]ZB&$+[KRM3-768C,"_9[3&&>IN-6+*H>
P(.Z\]=YYC;,?+M?-=]?)H:(X\3B2S/QQTJP,-Z@W^B:*VX;H/93S[C%)NFFZL"Y<
P;P$WB#[-J,AM->1.3EL%0E>Z\8KSD71-7GIC2%Z5&VBVLG(/(,-OI-M2.-;JQ!1)
P&=T1D17WW3!9Y #G.BQ4W.8IP6TY?!6_RU;ED7MMSAISYGQ.26(;FEGPD^Z'PM\6
P8)@)/,>L>9CVL](&+\5+![Y:U,X\4%;(L1VTCV(ZRM*:0YW7:EN"&-W7&JU)1FX)
P0?)+L=V6Z,\)",.8T9K&F*_-O$9]QJ.V?K!&H1]?^74KU,OP*6>DBHFN,K&,V)70
PF:9E)!MW/=W%K=4BM&UP)#V@KD<H]+E ;HAN-M:T=-2")VQ4_"1>R# (Y!P*#AU 
PU7YVG'L%OG'$[50D3Z.Q2++)I@$\4+]S_DVJ4&,'R=(*"$*> ,/S4AV2:+;:^I]G
PD!"';N#A,TJA1^QD&$,OF#''9/R1#*^LKX1X"4U?44?E7[GS=3;C2LS2#UX^$-SE
P5 ;1+O"/OXT&6N>+_E+T)X8IH*Z)>OKJC+@'T03O=(?\GTW%I4Y[9^[&24\VGFR<
P<4X#2<2 ^YD/@5PR:^.[";U?@;-K@H_G8TT=<F:G<Z<"?KW*YUF/3K4G==7/-PZ?
P.LV4] .E?%"&B9^!;81-RDT$9<0ZK)>'&A6FH>Z)I'5HO( "RMWTM<WF(Y;PBWM7
PZVFAMZBX%3"?0,S#0GB\-J/PH5(K<S$(TPCNP3.C-PP3(BC&&'A;_(!L- JR/I']
P4@V.^R+02]_.X,/!<WJ;<U345]ZD9,OQRML#HX)KW=R(Q-4.;4/P"@H^DYA80D?5
P>8T #\*=:3;@C,A;015AJYSV.VH+(I1P79XX4/<@O.(SC"W(TV9C9I0]+-A-8!.[
PWH^,W(G5<7'&6<?Y6Y*Z]=)DY_\16P,8Y"<-\7]$ X;J+ K<RJJT,HM>I+@O0V91
PC0)<\+$#?]UH<PU7>:RH,OJ:+LU;KVRMK$%TY.00=B346_OE4BFB_"G[*=1 [?^C
PSHN97F-VB;85Y5@&66XEK]'CWGAUG>M:B9I&*-!91*! 8?N#0Y4!*B5W'6?1E'FH
PJ:4C&8)]D_*2NN#P70H "$*O0O4L,._E9%FQ9-4/B3CI2-D0S@BJ+:(Y(^JY>!OY
PY>EEU:Q%D\(?!E.]28B^EHAAJ52'_ 3B'C03.D,)CWA1,UE1H55X=X.UA<1;QN_I
P#XA>E+98JK:V'!C[]&J/IEII\@,LH&5TNT0(^YB(+A1?#PS(P5+P["ZO\7G=YH9C
PL2$>)3$YCJV&%7EJ?@>,E&&_P,6";$))KO4M1/YQ(E7"YB#D@V8P8-\%A?60B12,
P!HGR2>P-W\@OERP=#Y/I ("W<-NHC5D^^.I4:.7Q1/.0?.#)=E%['\#2)X[EX+O'
P"F$QW-ASE@*@F&)/I4166MK)Y!EBK?(5V)L#8N !X@+1 I=T@RH!&8*D"TT PX]G
P#8-V\4:BGDQ6Y*[*)>/O@5@IU_JISR'(QX8S)9$VW/0<F[;QW[MM((T0KL_JQ,7=
P@EW%M*TO4R]ZEJTHUY)+Q(&"-EPS)MC!P+$L9#;5!5%+Z%$(EKE3KYH#Y)PN'/<$
PMLAM@**&L3C'2DY-ZA&(<7NV9ZICLD4PM6))[GZX0A)D\:"Z$6A^KBA+O?WAHO5@
PB0&&, !Q),:2VH_.!5I_NA-1">OEN#&U#@K3%&:KTPL=!I8L ?E1U.PK\Q[PF.S6
PN]@^3[I7;QN71:Y"$XFZ*R\:=OGC=<R"GM<KQUXI62N,P38&2XDZ,$&WUNL\!I<D
P-9AM3^_'Q;N 9#1L9X),3N"_Z(C#MKT)L4*70+'R=2)'6;&5HX+18 %T/KZ.!D%8
PRR0AHG@'#;-+&;;L]2&B[9F:F1EM=<D1<;<_LO(2L%$W:3,2MS%SZ,;/NK=>P>FD
P@F\H;(+@V_)T\6,(WM9R0Z,ST@LK&PCEC+I/3GD-II%0E?8#C<HWYR)OV5T'"H<L
P2/F,BU9L1]R>F.KEW61Y&NUKL8RPL'+-_51+6*;U5M2LE[Q3:;-K7\\+*YE)A(?B
PJ/,VHFYKZ4Q8]@%>PTO(=%3RAS^$,SG=];5["EL28[C+P1[PPORZS=-GX'*)6?U^
P.TB6R#-=0E;L$I> 8&^#W4@,_MR<>!84&C]<@-4(B^@#?),T0C)KK8- G?8V33 6
PZX)GWV:$\#<!:Q&"]ST&6Z$(+-?M2S)X$')161FRVD&DJ. 3=#-4[5@["R?63J4,
P\F^H;V"+P'D4'!D?5R0 ':3 ^\Z\<T;LD+VUI,?C.Z;8</ZFO%_0@R,=6I.3@Z. 
PPQ1TU> ^:9C\@^MK%27[H-7'M.J>=1V[<[-D!>L"?'VFOB3N[Z_.D7L+3+DRZ]AX
P>*1C8C$;:"EHC@K QBW94H >H$!/'C/?.-D06BL!I?'@:WF$'$CB4"T$K]_-'9I+
P?=/*E_.%S!0,V&*U< ,MHY&BC]D,#,BW'(7WH'U2@MH(%\O;=,H)2(H;4Z@?H@?,
P;-;]S*UEOZ3KPE]XX:A-7^R:,G]!:DYV%SJS72'2<)2!(4\#MPE&A\+S=BQ&0(C7
P[\^[VT?:P$4P/:+=\L/9RJ&.@[[%>HQL[=WD4L"U,6<5G9GS%9N-_U83:IRY VQG
PHV:3(^@$[>3=ZP.V,YUM@#.*X1=-3O44B%"CH:N-GRBD%HI9':6Y>I)/$1[9M;(B
P%])<HOHTQW--QQSZI(FE.=\+!"/Y_[>8@(*Y_N7H['A,O="=PC:^I/8K;&EI>U%K
P9W>.:8C?"7]1:<(84EFU_Z1$F6'-O'J\;56@AS;= 41 4M"F];YM!$>38-D773\U
P%(7.X;HFASIQ KL'!U\C$1*4^3L#7/O,!>YU<_NKGWPSTT&^K/,:LS1Y9WR\T6BD
PEFAV'?PTV@C0B<[WHG\H;T/E8I1GM+#!_=B%/^-OMY"LL>='0R';"PETBE)XAO?R
P_>_8WER1N>SZ<E9,2@N\G1])W*_T[$J*>@)B,Q@^C5[#_MA.8F _ =!;5]XED7',
PBYUH].8M9E(C3.EHE4!N:0NJHN_\5)L0P=B2*4(OY2G\EP1&/F"E9I67'N\!<RK$
P;+!'P#0?>\%;>**I/":PSUHXCM7VHUKF8.O$B\_DFY*549AN'H>-M&(<=KJ&X,,Z
P6@(ZJ4NP8QII3$$K5A&/K&./&PA;2N@G:MF?L'\G::773 ]JTE81?N9,T-YAP:":
PUZ$)[-+(NDP#YD^DS#EA9HV'%CYJH \R4*DZMI*JIC@@M6D>B"0XZU4A7"QX2@8D
P?85?EB8%)T'HR0#XWO=XA<6:2OFX4=#?Z!I^,K5R+/6;JL+@R$Z]V#IC^AN6Z&%L
P23/[GK$>)AD^2GH4;W2^@6YXD%*GVJ;0YDXC*Z/+<=,2JW[Y K\"0L.UJ_V*G4M&
P=[7#I[[4FA4=0I1[S?SUZ<'&./3^+3P])N[9B+L47T!!,E-@M6SY6?"'VUXZL[V4
P;\= &&S'3 SXAC2X4^3;UQW"Z]X^^T)0(,#"ND,/I/9RE +V[N%_VRRDZ^MSEW+>
P!\%@2M*0UG$*L$U!WO'E)>+3R_FL.IBUN3%E#W[&"9[$L)0- *>7<G]6*#2?[AU%
P*!H20'H\6<W&H*-,- )AP5/!A:"NS6D!7Y]@,P?NVJ2L+V/.-1)O9C<;\66Z9<S#
P/F8CI6J!CT#U 63J,+A9'[NVFWMRV?5/VAKO;PX%#B+U=B\3FIYM&XB?WY3RO%'_
PG$M3*&6+XS IN@+7W-L<M E@?<T\_BG+X!U@)J56!^61C5<"_/:;#/W+N;Z2'SJP
P%2:F73-#YE-N5WPL1@!KY<8K^XV^-CC'24ZLL,E0E;>0)>G\Y,-;["C"N!$_.:%.
P,>IF<_J&Q5;$-BO-_\)W-P""V=@ME3<!(WLD.PV%O!JTSTT< R;<6>)M/4:L9@"+
P#"E +;T35R2RFXVW0F0'6'&U_JMZ0VWOD%L5O9!*UGN2+FV]6;> VLVPI;Q65RQ;
P9JF)W<17%W)74PHQ'YVY=:OG*,D>.#A24WQD\8O7JT2BY3QND?]?0%*'!KQBCPG&
PF%[@;V.!)^IWD[O&@H[PU[*+5D9"TQQT@ KR1F1_E+*M=^#<9?#33!-HMAA$!/9!
PQ8JB]K=A.0J&D-GWB'R;:8?L6Z8T7%/W8))1 9LNQM3,5-C///.#:(]78T1=8>*#
POI!A&N'F-6(U7 PY[@-[:@CIGQ ?0*]P<XY4JO'-?X]$10_\,0R)Z:"C(YA2#PY\
PW^-ML^QJA31K%X \<Y)-T&/$[33%@O&'4(09"X9V5^7S_>S%7_Y0/K*# Z9E0B#_
P0021^?%T0W$9T,?C\")]![P4M5N+-1)/7<Y$&\G<LDID,SU'R1:?[71R/BL"'/@&
P=\I-[;R@U[.$)TN.\UB^O(Y['?STVT+UC"HMK[,L_J:3W@SW]2M0[Y8\XOV6J[2_
P7K.T)?S0/RCF^!;W5HL8?$Y>V7R^YO:(^SUWOGR/W)UAK[+&M -B>;*=I$DL.S#]
PH%1N."$ISYFGO5K@I()"+FAMY&7J%C?R@%+:,M%B!:,6E7"+3]P5EZ:?=/*BC'KR
PU6FS()(K8=++RF]\%V3_^$"OZSK'Y!,8GB^/Z:7DK:P>![&[BEBL@TW+C!,?M;H>
P'7^AB83DW=FT!(8C<:/YTN?)-X&A\V.!\^ _1\-A#J_T'?>!?\;6$G^0HM*L?C5>
PE?$-K?6ZUHP@>,DB$, ;-7EJ([<4"J7K/R5KJ1=B)&G4(DK.[9XF4.";Q>H=AWSA
PP;X).GF;'VF_G5C -=\<0F/N',VHS4C4D@EA4[@)W=1"-TB#^G"\?[%3ASR(/F8Y
P8_<'S!2UGKX:B8G0@**8Y:22W86WQ\#,W.>-"!^\*Z(=A/?\KZ@8_%[SV_N$^A:6
P8D1'O 44/R<#=AP@-HEO6OCW"3()P !4 2CF8@+H*,.)V3E$\M%(G'SS9YON<433
PH3$_[1:\AA;2WR+CPV_U"-V>[R]8D)0 R&/( ?JIFWC1HH#O =O5+MO(V#WDI$;S
PVN81O(FEZNQU)Y\;MYWA$%].O48F_0=A__LT>";Q5[\WCLIJ#?$A82C^O16+L.9 
PL[*/Q'^[O4A/+5HPR^N$]<TY:T_.;&;9YY0+,L/$9Y;>*S]R[BT3K4]C(??&.ILK
P$@N+&^;X5"L8>SORKJ1B?R'@5WANR8M >1QJ<"O'.E!'_-TVSKL;60DS]6R5F0YP
PN 0S1A'Q!P+$<FY!7 -)"J5QN7/._P6VXGX\^Q#C4K/82A\&B8DV#9MH$BD/=LUO
P8+^;5DU\JHY4:6+P,N [F2<\PFC#$KU('X,X5:.W*A=;Y33S2HI!^/$63(6U/_3?
P("4Q2FHD'9&!+BAYT-@XK/0K(7X:S(SZV<D/!E7?$)]#O,( N1MF<YIY;8/E)+2_
PZ(  73)RFYE,[C<#V._I6\?[0;O^$;)1MC:N&ZV6N/30MK?D\F:-_/LP)B Y8;R\
PQ)A&%E_NMY0YCM,KX+&'%=<^L[N,.(;4%X_I44CC\VN;3V=!$@5J#<&E#J$F83Q^
P4TCC?[FDI,63]8VD"(D]@CFWI[4R)WN<BDEAC() 6U!F9ZJ#)A)/ &YY>T'][HF4
P)K!"+U)?G(3>*,\#0OYBU.<^O$QG^;.(2=<F5J=^1BQF0(1O\:L*+;HBW!S'EJ!!
P8UBB/#ID/J!NQPT<.SZ&*W):0Q=@/N#"J$23]/N5\6\?VHO^NH8CAZ(A#]H]6UC@
P901\'L]K'QE&L[AW*(0SL!NBX=O8G9&PDF@IT^Q=OLQLP^5Z)?G_L,K62W2J31.>
P&H#UCARE!DPGX"'0-(X4O;L?\.1N<= SQB@#0L_9^!=#A_"LQ:9=&*B2ZWK]:D.I
P;\(]+%(?91-B--EO=^GGT</@*(6)9EYGRD% T;9W$04YH=@.*Q 4P< <G/TOJ5M?
PG>>@P",PBH,NQA7]G]6T^3CIPL6$ $%566KWT]'FX[U08X=J<&A86GR+?C;R%TM%
PARZ""* LC$*<T<1, +#/%V^O=:4,#0F\P^ T[?70YE+1)HFP'%("1:Q;<J!Z!)"^
P^SXABPD:4#?<0_18#3CF@.L%6"K(2/[5 /C66C0R&:NU5V%?>WZ.BRHCYE23CF$2
PXYXP;7!7'WO/>;I!ET*+BE8BCC.Z&%DN<[O? '[^:KG"(6UH6U;WRWTY;W7_O4%N
PG%%'+^^!$= X4K#@U/35 W13Y=J7E=)0]!:U%_CB/\G2*CS#237*A++IZ?&R="'%
PQ9H>]X4-N!=XO_MTB).HV^.JD$"_3I63OS-O_<SD'6Z,3Q_)?KDU^2QOZ!#-$::)
PO6G)1#,/Y%_"C9F1OH61NT0<OH["X* ?J?3+C74]<N[F\N#B]ELOHI7D";I$[5S/
P-<E)IIX,:,[6$H'-;>,:NK5TN.D(:$8U$\]FBG6+JE=Q."W0>\QD<VSWQ4> $^T>
P-_ZOUZB<):_QABNY$-USE&%OFV WWUP=$<JS<IS,'4;P"]"1T:(M0#O:C>WV.$RH
P^-=4?72099JJ)C'>Y\<I WYU5YN;ALQ4[DF@_XSC@NGO#MIE9%,I[IU#E1>*7F".
P,/0=BZ9\XG[)/P-.=4XXW)M'!0FPUF=OTG19>"VW7Y-3#<E0WJ6:]_2-N<:W]=IS
PV^W+71[TF0/?3$/>]J#B.ZF<".XIBGO^A.C)5?D%-;.:N6SBLMD&6I,##P,R%XAH
PPA[_=V8KXJ^K%(5&NR_[&9V!H=S9B.>0-5H+F!@BRFS7(FZ:U?4J.LKRU^F&_L]U
PJ;A=QPK;>=5F[ 7Q,NMJY/58P3" :/O5E*WD]!K,MWW_8E+%UEFP\K#TD2=8M&VO
P9+9^O6<);]8%<>TP3=^46LS'W?N+<CINS"#L*!U%.\!L8H*3QO8W+%F1/A/H$:HR
PH>.TL8/1=O>Q1UH7,NI@%^H<1'/["+=H5\VX'9$A/$VN"6 +EC]['VW_<)341C09
P-H\%S(L 6B%#W>&\?J/,J-(+R74G7U@<@W.A_'G-?<TL"Q.LW#%)0SYY@/@U?L +
PH9_NH1;8)7%JF3P=0SVA X($+);NQ;J%HP?2R@4E:25N8R 3O&1CYO=[AY6VT\/,
P'=..%,'4= J\0X7A*ZR(94:$R@+"3F@F:",R18--,L$98D<_D(5;FL$2;S_U3A^-
PH< _XH*+GPQ5#SJ"6IQ"YH//T(H4^B-19:1B'B6%YQD0KJPI[V_<"VK*B(ZSE\V/
P<*>#%8HKYGH.EQ3_LI:"IL74S3#\A<K>+2-0820"I\HI_A6[-(.%"$9\:S/#K=[X
P!%='%6,"'W6V4@BXS(.5.$C497[T,?FZ<@N;-4Y(!IV\U!>-9V+<RFX02I!W<D-L
PZ>LP_7I;J1]<1PFO/X0J3*=#I&E+VI>UA+0^ &V6.,_Q N."^!T(MC,P[Q'8\_S,
PS+?%[?HX8P=>L1]$&4+O[Y6U#A-HC6V-13I=B#<#INAZ /#"8Q!=\4NF!U^BS&/1
P6A';<:Q 3DQ4USS&(A0>!).)%?K.HR:)/F9:;:R[G!#>DT71-US.XH)OC ?[0LGW
PH1L[N10$I%TH1'>>T'?YUN-%TZ)^03F$LSU!7)T.X?1VV1:FSK]Z:>">.83?%?8%
PCA-IC>QS_5TWVQ?W;5!2'_A*>0ZVS1=7QHDP4V Z8M(&5M="='TM 'XW]SIIB# Q
PR$3$D+]-?QWCV)Q O$*V8^LO5?YTFSKKU>M<ASK4]DW@L/"72E70YC(-9S6MC!'1
P[?%SU!D$!&?P0ZK!*B!)!N%B:-KM,/A@\L;IMW50/"3+L-P*V/L?"E.[>Q4 A,3,
P(?=\^];I6MB38 -HP[,,P:O2@PKX.T@M-7R(-1%P;J7RI;0*&*E:)Z6'!%TOVGNK
P\M4WW5H/L 0T1994HA0QUL5F>Y^&'V,]K&V"Q]%T[&4<X\CA\KAH;P03ZZ*A#J%6
P(-$LUEX0[GNJR_=79P\F)]Y5B_@_5.HKL7SI!BT>Z>@-68-1*->RG2P(&<MK=E]E
P^KF=\O1_(BJF+RLHSM<1=P:9RK7XH@)Z=8A='O9WN,%_P+NOO@YT.K795,';*,W.
P>C%=@UI3!K##.R+\4)OWFCP@[9B_Z78@_TY]S#69P,,Q+0RQ*RV\PU%W3^]K$(.F
P87AL^XB52YM2I?58E"A!6#^I8X,)@AMFCU!>P '* LA&UNJ40P+;?)AD^5 Y!AZ1
P/DS3)<UB13U3E5\0VZ0SGV[Z_OM07FGNZI4L.[*Z"*\:$$C ^C#KN+J13-H*1W5V
P..#]7([+S;P$J>XNX T#%DS(#CZ5&6E7?0(.9-:$0)<?R_(_XSX_)T\A9N\@(+3(
PYPXR-";)D,3TQW^-NCS^C[BXJA7&'6N[M-V3JTKVK?N%<7)GC"X2'DOFXLG=ASD'
PLZM4JL_1,L:MY 8"/$W925,XD&M5BS);22/6]YR=Y>[Q^N)UYQZ<R[3S^=JL9WX\
PA909L(>,+7/OI8:,;,8ZOM]-' UTY7>0M/>N)\,H50^S=4WY]PNA+4@/#8\C*^7:
P >B^C+0,>%R"M0B49UA<>$8E8>+DO;C;W^?\1 <Q3MP=.YUV/^Y1O*;4[(\>&APR
PO8H8W8F=1<5Q%_J/5%[V2+4--SP7D7)'HI^2<F:/]&<$!&(/1N)A*$T<N 8#=? <
PJI;PU9-L6RQ^+MYTEZ3RCV21N._;,OSECR+)O"FLW6W ]/C"47$;J>KO6;E&8-1;
P\@4)>!\VE3&K-EL$)".NJIO<>F;1X:MUQ*4+9:$L>Q^T/;&&_!*#KZ4?_,0*+UI$
PU]>P!(^ Q]P+NY=(7@D<8 :A2J!>?A&4\QPR<*)!(+KM!GM+ND9IQQTO8F=HLU3'
P_2W]7KR%.8S>;5+!=/H/\E_245>+<544#P@,$FE$O%4]<^:.+M]1C21.*ME0<WS2
P .3I]9EQST2GF:@;$U[R\>]F2Q9A$,Y"ODKS;QZZT[=IL2X4/#[DD//PSI$JXWBT
P+J5(35RI)]-Z*\R\V*"3CPRI,K>C@$;H_$A-"472 4#YH4E^\P A"!<64TK8%EAF
P1NA_F<Z\,N_28C 19KXDT/."T#?;@6J?;H$;+I\;20OC#0U:))O%4G*WE<' .* >
P3'6<1&'IG-O0LV[N9G)RG .(FV\:?;RMR6WT,_B 3OVJ=?Q-4SZ(-JRJ_!^S$!2Q
P<7\,!Q<'.+&F?3"C]*2?P<E&F*?_D<3&5K&\BV/\#B*K2*I[J*YPA63HL9^@89?&
P>&1I.4#%WZNE8U<C/K3T=ZXA:+\D-FUOD!?@WI]5VB8.Z>]1/:Y0GSZ7=4J#1)= 
P^=#9O'N@"*UC2@<QVWW!4B^(><"DI65. L=;6:H075&IHYR3%.I:*!Y'!)V\;[B@
PV(FI1OMT;6,H^EW_OE''YYW6,1%3M2?;ED8=^M'WTZSHM$ S94KZP\P*T,V3Q37+
PQDI.:+P_T$#'_^&P_RN]5_ ]=DM"@3<><Q"5S!4C<S.W)'X0IU-21U2[H)4?X%>T
PWB#UY2"UDO_2*B<PJ/-_9.=N_F^TT][D08IH(.R"9I.(V;_YADEJR?.#";#6/JP2
P&RY 3]']C+4\THR+BL8T>+<?H,'G9R'+27:F&%=B,+;U<G: :]=X1RN**T,F5CY!
P.FK-9.O@020:C88_5= VRH/TMP39-NQ!?RH?/M%#>>U6BP/87E5@I1] -!N-&E%?
PDH2/O)F]4KA9';[=ZI=7KD:01Q,4X_VZ[UR"7.0F&+SG8RV[I\ B?&/9>%C8S(KE
P<<[9(L61:@$_TYZ4C&0<!;;YA.\3D7NVYNMV_=,?'DI6O,3_/I^8@\,XB8N3.1Z;
P(B-=BBO4S?0TTP"&>Q[/0317/X XW-M*G@]68/Y%H<Y%IQM1A# /;YS'[%)?.."R
P!?K1J;Q"5*AYEI*GGKG_*G>.&^'.;&YQ[I'/>E.G#Q]A0>*37%VF4,Z22:'@RHK=
PSS9+_;*]7Y6%SXUI,MIP!P4;%EY(2JR]/GX/%S;H,8-T.D.+M?-6),&Q]S];&>5R
P]KOX49H2[:[+]AA#F5KT'^*Q'<\.QU@"-_"[AT)]";<7C<P]7AZAUHKI/^-P&/T6
P[TJ\B5XSELC-"TL@>3BDW$MXB;\6"WB"EDVS/ 9'-8QK7=,!S#9:,W!1D2HX<:PO
P <L,]"1^#P8<($>^V?5?#:]KFGU3/JRZP*H*'HYY>Q])0\/-9!D-%TEE0\V/:QY=
P&J&WPFNFW_?:LT%(38'V70D <5/@AY=M\]M8:!H[@52[;+NLHD9'*80 [J!GRV=P
P$3=<=F@22=BRQP7S5#()(;9#>YQD+D'-@IXP2.$M^B*FYY?V:1\D.?Y\&1)!.=FU
PN/@-=/.O0YU#1Z#/F5CY7%94+2D_-8WCO-@PIEJ>BK>>R@Y8!>>H-1PJ'8OM3,JX
PRV%]T%;U?+J/RWL<TD9J;?R""7Z2W7]ZCH'Q]SN8#;]/3*%4$7![CS#!URQ+H?!T
P:2-^( W1A@8-&;K#XHFJZR1QW9M^9H!803_5_/;VCB(1VS_)K).+'"RA4W,A1+[(
P?,^26O3>?CR);^P^7QH9Y1I++1$[(QOFFCX\ (XVUY,=]/=YP<"_B7SMV6P?JRM?
P(]0[=L:HM)(?Q6K^XR:X!A'S2^M3[*.<VC HSISM3O'57H+_W@SQLG4'*=ZH\3Y>
PPFJJL[:#/@/>J:F<'C'%&G^-.'GV7U1G/,7QY[%Z$#F*4G!P%D,\_I"ZU_HYZY0B
PO)',DQ3E.J XS[=3&G;C[IOS-<79ZB#R.(RNC1&$D* ;J=2(DM.-9T2-4?^5#>HK
PSC*N:) =$;Y-EZ-\EC=ECCX394IQ.*)IV" 37>;@ML$5!>*W F:^DI1 <OW\&SN9
P1M5N^-QJ)&!_C]YR#5HVA-1QBJ!-,T'O92W!7CJ>:WK[G8S_\XW(13<3M1"T,VJ8
PY!QIDA1S[HRX"V;>W/Y:6,7\&#5ZI6K&$L$B(TE$U+PXAW?I85OO\\&%_\(""$AZ
PMX0XY0EAE>GRV!7K@5)C'Q!TX^O+Y1JO= +:Q79YUS)&F!JNS5>L9&1N3$!\ 4%>
PKY@8/L7RC@A#V[SX]=H^5TS<FH"Q^9CI$FL),QUSTM9%B1*Z-EL_ZR<9-N!#C]0*
PR$D:(L#!CEAYM$JT*XP!(=WI-A"0M1,M1]C6[(ZER3_!S_9GV.3YG+(K%[+;ES3<
PEPJLJ^/[23[U=]84-),5++X)T,XL#25TXE^@0DH_:4H'8[RXCGFKN2+YCZ)?^8RJ
PSI#FR' C%*IN0K/:)I^XPE=/N5!2TX&$KM+P5]_MLVN3+>7X'&_H'SS:W^F*?L2W
PV[!$;=I2433A@7R+UEN'%95"7"-(,@RAOM)03B>MNE_4_J4)?W'I!I3&D:P *O[4
PIT8>*8HB_SUUM?>G#1P@C@IDLME5)%"PMQRF#_'UZY^.9]KJP4\N#PDZ3YS:O)6Q
P*6J5CH9-FUK:N@,%2'VGY423W!LIV"P[(V\**L?CUMZ9@/NGBE&\?#-7H>_D->FG
P/KL>V\4/':9A61/2\"+0=I$#XPIA"G;4UK@DIC@QWR#L0' WL>!Y^?+<4_+=TG2]
PI<]&>3+G2<2-+D"[<,_1U$K3P(RQ-DG&E,#G1VII1/DCH$"5$]DE;U**LD7Y--@N
PT]/B3X?<.0[9<K'I\5F'0);K2*DSLQ"EA?3K.&3#2LC-$WG[_  Z 95X3UE?/9=Q
P<D9U_JT0R[L;^&43+S?G7"$%4-U=Z<.VZ"BSP-QAC+I<N![125*)ANT@]*B+D(]7
P,',31B9U7I?8:.402.$*E[E'*H," UYR8&=,Y(;$\9:5$70G4>@] Z*YYHGF6*UN
P,VO@OH25* =PLEA7IA?1N2N1$#(::$9<6)-FY1OMCM<L*>X[<Q7,DKU8OUA(!I-/
P/W-/PX-L_WU[7 *0:1T^%>EU.I=0R^B+O$+0##Q8" J"=ZUD39KS@W1/^5RI*4LM
P6RB&OF"]'#*NA2T5ZU:H[2EDRY.Q-62)[ '&?N8.=290*10[;0*3<^4&B@MI&(^]
P*?KL@TQ5ZZ6EB^6)#86:GR7FR:? S)>^]&U CS42>19M+X0=\%P;J?6DC2;3 =%%
P2/R$&,[&R+0APJR!1.F1271H/4YFEXV=CG$U&F6-?*\D0*7'AQ_1@6"8A4R&&%^W
P_?CZ(2[DKQU]H%ME0N<TR^TW4,U+:Y6&C0RAI9HJ_$E*6*6 /[ 5.66K!$S-F"U_
P3A*T/ _5#'=32\0,#X Q4C]>;KDST$$3^T7XQE=H*%]]X, W!T'%EN:/T8SM9EDC
P\Y 25 /:V+L=>1M_)==$IC *;CI?VM5W6TF/@WQ!^FW-T+$"+XITPBIFJMZ*+C'6
P7#P8"DC3:?S?$O>SL6QY2OGYH W5&AN<BD7C'9[J5#[3AJF GO7?(\@(T<''BD48
P<4S/K!5M^+I#TN2:6SNV47XC0J+0();+?XE4K*9Z7\V4;60*807'[4#22%+(9PG>
PODO,/+2L^VS49;S2&=!O-)*GQ+0X_T "\". >'XE%P7R'4]7DGBZ/13,,2JC/V3;
P5[-/+17',>EKE<N)= =I00:;.L^9S2WK;@=+B@L>);W:IORY;E RI/^CXDH3'.@>
P: "P# &3(I*^P<4V%C$4@G5)\>7QJQ@B[UF-2T9?8<BTR>*\KIO5/7F_%?#0'=+,
P\?>[(MIQ0F9>V "0NX.*W=>,X1SQ8V@.TM68K>-HC5&_MA3UX,BKTK7.AK^VX?"0
PZ0NNLD!X4)JN9"D0^BQ4GAU<!>?T)5\#48O+%Q04,SX-5D9(ODXUF=S&['16-[T/
PP*O.L2GXZ>[TACZH$]PT !@ &6"X58AUU3H7;IXBOABE_JVC'&>"Y9:R7+GSL=8X
PW%D+E7I=D96BF0 A8<2)%#<V_'#,Z3!=\GF,3T5;?N5C:A.GA-;:6-<82.)AOY.Z
P% *OAB#5S:W=?2)* X!WX/:)<-23R!,[2WYSL)VN#RS"7/^(0SV.Y K%#!BB;BN.
P*ZJG_"U:N'V;M-:\Z6/F&]&OO!'7ZQ(+ @OZ!Z#%*?$A)\SXZUB=N@]E(VS(<B> 
PH[< (Q]OGQIM .UG>4K%0'!M>H@ CJH.PH1J=,B8[Y 9-KCDY>P(4=9B^48ROWK9
P5S/FZ-BO"4WR_SP[JI1_S*BK2*"+<N.L2XD7L69!X6 2M$<6UBJAR2JZ3/7SPTM,
P9?EM_&*X@0#3J7G=ICH.;V)/A[!CX^2Y,.I_J#]P_<.D&",*#$T-(U+6JH_3]OG^
P.-\8;(@6D!P6W-,'";REXGM(BT/4HN)']9GTWB(_U:.599P,RMHL6_8.\)?_N@LS
P^ ZC83@B[L< M]K\-F<Q USRZ/PV6XO4^>4]*^&\.NM]Y1X2H [.BO>EFIXK#B74
PWO,0 ,0GC&$#%@.($&=]BR^!\/HIPP^D^8 XNR.H-1R/JUPZF#L<[4O2=W]?,8;C
PEJE60.H/%5LS16F6'_(Y^DO,H.X\W=?(R#<)Q/@5@=:I!*.14.:2&EPR^<X+X\XC
P"&YJ<1HF;+G7..5F)YC0"2##+-RUY"9 AZ%F'@K!3Z[PAN/RPK9(7M;?:*&CB;9O
P!0 ?&\GC_I+%?D]6.A\=B1J1LSTP6[G\YCP)Y(,G/CR[YK&8S O_@LVCO;P+[!A4
PP @)30O:0+DU5&TTZ?SZ#DLKAVQ.E.-8VV2^4AAM>)U3#K1'L$DSU(,O$LIQ+Z G
P0@9N3&J0:QU&3;V<+TC!U!R,?KM\?#1D<C 513A3J[54''MO0+>R-,YS0UUN:K&M
P%%B;BE**N"M=W/*],5OK/P0Y6^(F##ZS!2M,^M9"&OH^_[@/;,%*6M7FSPN1NNL(
PZ?-\2@:C'4"U*]W-#>N70 H=]G,.EY8?XUZY78LA(U3Y+SAOW>3TQD(*%^481,)Z
P%%/W391</VUH>O!'=ZC1V:8U?GB.0W>V.C)5TWFY"'*M(#2"ZF-B71#&A?KZ')^-
P,TS*2 . .5%M94W>MD*]B.5POFY&/KF+-^#+NG[+&T['!?L#IZD3:$=7)WJG\X"+
PL*"$4S>,CUCPP4VDHL><[%8\?(3'!1-K!Z+'<A$1I3[1#"CB"N$EU;?":MI8W]G(
PVQK8OW-1/P"R=QZ//"3;_)5N6:W8[+I>/YS,.I4'GC] 8G(LWY\26^/P^:-[3@F[
PQ]@K)L[!Z1IL6W712?<-!GO:_*NM^SH^$+TJ[0-N((T=='NDY5K:/PJ0<'%D)<#/
PAX=&GU=EJA1J8N %8+=+@<:R&<TE=TGD!2_$;-8:W"Z3K(3ZM=>^\$Q!)\=Q*CQ^
PL_:JJR]0,!N>_])N+O<IW!N[(,G*C*NF4#,\=4;!N,- 3GVT[8$>(H[3:IO7JF=J
PI%/?_VR97!SJ$4RPY<5T3'&(\E40P;9#4\*,MF. J:Y0 WF6Q3X '&L@[<[G85[G
P>@RXV*V)/ RZ7#A\!4;'\9&19%*XY:MWP8>- 3_136[WYOP(9LZG.1=MG=^PR)/-
P^B1=U%-9HV2]8N'.J<!X6J/I7;>A?MV^J+DS6Q-RJ+"H) JB?+Z&F V0357&7N2@
PZ]>S!.FI?#)3YL.1-KY*FU2>:J&*V;A=2!4+V'_=/(OPUFW*'X7)NR1740C!FM3$
PW0I-B<Q1GJSP]V((?KUV"A ,:*U=YJHDRIN[T)NNP+F>$!T38_#)R?R\Y%XRX7@,
PEOSK(1D8K&>!+F1I:2P;6(LUT#<5@VE$<4,X(?%M4(X_4&,PJ*-ZO)U3-?O&HFCX
P!!%&P?%2R+=DI]M-]Q([,E[7(7CJNGLV^?"INO0L$@J4HS0@27(I)77DR1>1@[U<
PQ<6!\::@W[_I23=F'L7)]1J>Z*"9\'T)9<>?WO;5H%=6RTB#C;] NQ"'FY+&6Z';
P?62M.A1P1Z\BX?]9_D1[8T^=S0Y9LDA5>7DH)'M([=M"/0U3X+F8;K)K94#%I7H\
P= \=@=S35W2G1V,9W(4_'*X^GWQYO(>;(MHZ*'*DV'#Z-&(V8? 4D6U!,WR0_G_7
PF8[W>*KCXXPU0(W1H!_\, CK :</H,ZT D"@,'H$1_K/K9]>^%().F244!L/[F>X
P&4MJ=B;)K)=-]>*%/H$ZV[SA\<PSOOVF8$(LIV[;9!B! 3Z+J [%I2Z F895]EGN
P2,B#S$G%>\!5F%L, :W'V:Q&VU"PGLTA3#YR*NVP\* '$H(G;^#VX8^E(WZ*7HH9
P_1H7;]$)IS5-0]5(_M+84@\> 2*"M<_G#RHJ1UY8*9*@)HX!B&\^H+F#:N2AREBA
PF4D$X:XX9IEM(SIEZ*-Q<)U978$>-' 31U5REWRR!1GQ$*RTS#$1L+CI5_@1@T$?
P1[(V?Z<E,;BWXL/[J68CN"&#06Q7 ._142&8EFCE;)BC3YU1G VH>57N:(%UX$%R
PVZY:\O%45"1U(I8X"(:9_A5'9,R3J<C8VJ/[#A:_&RHIQ&P?+$H' BA/I;;'BJD,
PW_%$6=L%A_IO;_7O?K$I\B(WRX\ O^>:];RWYL1)5B2ZE ^0U@KL_Z\LO(\N,Y2<
PGDT]G)M:/(, KS8?2>M&%L,!2@_I^;%H3&R_[/]<()\3-VTZIK^]PO]8-![1G'5G
PL$9HF-L#T((@4'8QFG$ESL";BX?F+)6W!\R)VP67S0_I?<C,4ZB!O#*DWD74*BQL
PAR\*R+@LAS%\&NT%"]H%RM!LYHJ9R3H)Z/]+38WA[X;UMMFB!%YR";$%Q8)#*I)=
PD>SZQM,-R$"O"4PM4ZL[_>?UDU]^5<S",Q$@:HTJ6$ B2,9],#O-NVG)TP%#36I>
P2OP_*@#*^ILVF&1C43%NYPHJ+J*G76QGD$GU9Q.Y1Q5&$0.:_T?$ 9U<[WN'Z^ZU
PT9G#<K!5Z[I3)+GP9+5K!_>W<\@A$&'U"T->=<P5N^$"[,O/A)6)L0_?CK7>Q!<Z
P=I%.@8 8@V'%"O>H;VM7JM9:@W-4"Q3GN 6+2KN$$T(QF..2]/(>VY:N3 Z)G8-.
PH60<(LGUMI%O$)PV,XT[ ?Z9$FI"+?AL::PE&M9-V^L6,14?!!JGBEIJ:61#WS5I
P;#>#KMW?XA OOOM .[I14@##GP#,;CU%'@"Q>'KFZ'QKS48V<9^;)+H?V:FYENX1
PX0P MMH$ CD*EJMZX$- VR103@#6G,:]B<X<3^T).?#WP:#NQGOI,][+0E67D55P
P=OEY\$\Z^026&>*^'XOB<%+%<^O&)-5J\7) O.1[1W;<@1 2DT3,YA,R=SS2441$
P-KN.R]=5T"J42@2.M5Z:=ZY 6JG6FL$V901XIT;9>Q3A0*[[.-)SEZ%QX?PJ*:2-
PD^,]#C'5G;]R BJ(D:?@1Q> DG<^)9K9P$L&*Q$-03SR??F]=G%0<N1>R<BC?"(*
PP6H-\A4G2[-,;-D,,-V$K:J?)# BS!QV0R&@_^U?@:;MB$:YI7QG+8[=7),:OL /
P)OC?R.'>V"0L U7)8X7VGOSO!/8F:JK@%I^C1!,%RF+_XY'A'P1J07)B+)@O0H?R
PSB*J9_&?OT2"AP*%/<L3?IP:LP)1TX0>YAJSY)Y)9"/=%*Q+B,4?R/]5;"O2T]GA
P(>0A@975+*<DT/D1$2X]STC/=E@'B%F^9]00XFF-.MV#K#(6UCZ H@.M_+VQL^$<
PVV>,RWU2CH=']1#ZSO>+?>?L4QHT87VUI7MTGH_@9$.*0$-BC*?R$).,8J_=S5'=
PD*CEW[)0H)YST+W*::;W8&V;5!KE;?9+H=9:RS=OHAU3 ,*J@'NB%+APZMV^J_V=
PDLO@]5Z6-I=']<]<([F4A#- X HIJLSJWL7-0JXEJY>\I];KS):MY:HZRQ.!CK0Z
PK\8^Y8$OP;UD8@8,+PZXF"QL''.G?=>,(BE_O P0STKU?68;OWA1,[!W09PX\@@3
P9P<M0//8^!7O>"5,G3,@[4:BYBY,<J4QO1[N2[@C*]8=3CEV7E?=W6VB+P!K&;(.
P9TF=_XAAR>B;KP8V=S4U9R/==+T'H %Z -R7+C';>T)R3N2N03Y93\JH_(C"_@DO
P#M-R'4Q7C'R/VIZCQD.=326A9R,H.2T'"OP6SW'NSVKRGLB-M+*[\JTWW_'7D?A/
PP;L<.%IG]NZ>&3'27A5-,! #P)+2E#7&[>^;TUY/<Z/D0_39PJ8S<.+Y!G-S%A] 
P28C^&%-B0Q:@VL86UXB/N#=2'AYJ0Y=0Q@DNC[[:^=])5-]:?WA-&ED#<IA0/JW&
PL=/FB-"/^O;]:O?@!E4RMH7[KPC7=H9E5HI^C"C^U*HG\_.8J.]=>.9H3PZ J<&L
PBO+T=*^"WD !N!H.Y% M'*:I,9).U(_&EC'H$P:LIWKE'H]Z(L3%^ Z=-F=2>5,$
P>$&J=$4B&O!O/GWMX&:55L'93)I#K3:9;6YY!#L@A%9>G)S@>66+0?+5PF?G4: (
P^>=SJ2%:>XXZE?Z4LGW'0+Z8MF8U]S6C<P,-6OTY7!/$:Q <GX);FC;H&$5QDO;P
P2Q&^R6)^(0>M0-1]EG8)+<I4*U^2PAL!>';WLN@<7$FL.8T8=!>_?>:4DM0>C/*V
PMIT=A<C4^>9EFWVF B-C+4Y$HESMCZ"@"-IR<=PPP 8>?"_J(=/]Q%KX3T,!>!Q_
PHE"B%%"52K;N<WC05 IXT-_^W%>]D,;0//H@V4WS1Y22.>F$:>"K769_KFY&R;8\
PZJKZM-(.AWR =[VB(/VR3R7R3BL&ID!>;D!6/0H/ :ZD=&(\H1)%8^C]P*U\YDC?
P3J2SQ]S-G^7 9LPQ>,3V>+JBM!O(J41XQ(0F> _8WE>J:<]0QMV;7EYKSEH[ []@
P)(I>!$1Q&V+>( 'V8K+'!YHM-\V5- _Y<;@P'*DG'1U?W"5RJU!]\TIEU8BJ'M)I
P>_4XZ=*1V+KJAGSNH?#NY5\9^G$V']Q @_KOGBNDLMW? V0\8?0D!IS)@N,<%5*2
P-:*Y=L7*N?[I(Y,Y-M*>E,9'Q.1_.>6[F/^$_,QU\;OU80DO]5ED]:,%S10==F3P
P'Q0E =?-+$1*P)K06JP7W^A 2S2X_T_1E,[/,*&)P1_@EZZP<, &EE4%9/EV%UMG
P6'E>\X0S\$.IM^0_%8.[0OT.31;.%$^>?=UZW#24P[O=\<D8!;Z-^[9EVW'.:$YV
P5R1T.30E:?D*$PV!D3/SB@9CCDM86137K\8GE2!%OYBTD!91U ^QPNI_$4)H$%S-
PG5F];Z@8+HU"/_NRQ@?$DEDY5V[T>,S_BL>=Y[PRGY/^]=/E7<40QXJ-8]VP%B<-
P7>?8)*'5 JJ5P[(.!G>N2MKFI8;H/&[]H=>;IT>%7^ FVC=(D!@[*&VU\/"/B\=*
P%'/!7!_]SH+BR9W;KH)V!=9LRU$/BK42A-@#),-G)G/ZX$4YTEJ[DO'[&>D;JR/I
P@<<Y]I_B9\/P8LY?UC-6UGZ"/7[G\1GQ/7J6*PL\306+=N3[=,;(E[IUIP0%QU_R
P\T!TS+]V+9=8JK!;H^A@$Z"5A'TFC"]M3->'%@?A;W-76,QUWCHB+O*(G # \OB 
P1+S>2.O63*X>E/*(&U%<D.UE;<")'\_7@JG.D?G=4W[SE.#*<@,0\>:60ROB(UN 
P?:K-'=:&:\L.V2('.^L_VBMP)#O@#>81SKF?&5NR>-6]KI(%BBW?2Q1RZEQW;757
PU[0>' *EL\G@/E)T*,D,R)<#")-6@SA_38:QC.^BEC:7L+OKZ%\XU3/?H1BVN_/0
PNDH$1B+9"P3@%)(,^2HF9;D$ILXP[PCE7@[V'SFP$_'PLYPZR*7:I@6GTT[7Q0GY
P.QY>J^O(RE"RJY&I<S)JT_D_;':#%IMW:9;?E%67Z<RH=%2"#8NVBX:[-_EZ.R2\
P]K)L?S&?O[H%']N6A)?&@^PS=D(N" A<0EC-LR=X'A%!U4A$Q*:(QUXT+NW)*JK&
PTB \S-* A./WJGX3>/AVP 2,W2*+[+7APK)*<,7*/GY<<?%6)I <M5THR$0[W17X
PE/OIT+T@8D&HC5,!ETDPK4(D,H?4K@D]S#2K+H\RLT;,1TTIDMW^"5L25I']WPIW
P9VC3J 7AW?N@N<?$76(92^V4?>[O?3?;:?N SN)X%^>FD4V9*&WS89R6UUR)I5\#
P#U46K"&FGOKXJ-@S!L&5)>2&CP5IG=&#KN14\RD^A;_N R;NC7N_^MG<=RNH6H]P
P ?MR,$D]Z]'R),B)G,154'H"R28)D5KHN8EJ]C4=+@52U5E?'6:"G@^KW<6FRE5D
P[&D=KU9BU9:60[B-I61$*XX7\$%"BQ<H>/G@KA' W1Y4P<7>6')[?_R[BM@H;&% 
P,8;=(TY+R^7CB@?;,]/PFF&OT2?.QS7[SH:YW5ETAU.Q_ L_5:]#(86A*< F(_>G
PJ237Q8G,4DU!N[66+"CO"1YRF-AW?GH<[RJOCCNY"]9/!::Z2[OO9:G#E"]R#HN+
POX4 _?V\*86)1-'5>&/Q11&EI!)M=7]@"[(P+0>SMQ24.P^>D='.Y<3.#ER_YG#W
P 1*,\-'D]H:TK\UELDV(3'C$3</EE@5Y74+%?^-1DBXK9X>;M-5=Q@&8?3Q;::^,
PHD;%-[=%C,.=[^M5^)H V.+.O(4R#Y@Y;=%7(^DZ4JR.@HXM6GLZYDTP;CL:,E/P
PQ\AFQ(+C+77?<;0K**W'55KG _0^MUGKM)K5'Q_^GEK$\HH$?^I/:@@?IK!I0'KD
P3UOYE5U#)^Q,;5Z>&N_=APY*++Z,8^NG<2@83,>!=/<[PZJ)O<;%KCU0#EPJ9YK*
P.3:&X1+J@GW*6D6ZWA)]1I;@)Y;=70+_6WRFOV)5P]-]<.IJ/L?2%6S27_9"DE3%
PN5P)]2=TM[=R^&:/SH[1TJL79FT(%OHL#FM4!;8#FQW^T39$^GJMH?,+RP-U?[C!
P:$FJEYMD**DRIWOFF4PC.R\\%%^F0F>*,2"&;+3+MIX:6^_!B:WK9@MC5Q41K!+=
PXX*&[KN0]#'+<%\ZQC66I&P>W[CYS7RCQ#,O<BZ 0-HR"Z!(C:SB5I(/.<4JFVSN
P<(C1%8EQ>"L) EC&(D*0(1!EU6VT4X]93)23[G._G5$0&\>%$R?]#VCHG1-WRS5J
PS<!I<&N64I4+R"+;@C#%: <]\UC57B["E2L9?#-R]_4 " <U5]- ;G[F1AZ6>:^^
P&!XP1;XN"M8ED./Q +!KZ2IJAKAV_"6,+8.Q1?A+R:<YU[]EAWH.<A,;:+X'VC'J
PZ9-X7S'?''G33"I#T!>]?5H5C2R009GW%_[KV[B473DG[\ *".T4E'9RG-BB9"D0
PH,/'^[I8C[L246CH@YHMC-92K3N:T=&<*G\2Y0VIM160 P(;"KS*\TEL$(U;$N]=
PQ&9O2.B*D:^$71GO883.O%9+HT]8Y#&PSW>\-S7?L&BPO& [?0-9F!RB5:HIM1, 
P+";&O77=[>=P.+4/QNXCFWK:71_^W2E)EH#F;1<H0D\#+R<YN./U<33W3\+@!S$'
PT/$VY.)P?>>!IXWMQD!SB(1XU@KU1Q_-)W='>FM*X\XQ:[(/84E)RQ%<FPQ=(Z[<
P/,QMH[+E8T0]@^QTYGVU6 5H%0HRPM$^I<54.,DS(>YKQV=,F>;G1/WYLP&#[T_4
P Y_!5*P6"Y^6O2^:*CL<?)ATBI E3(>8L)[FXXWQ$9[ILX,=&VPT8QRR.%T+[Q+0
PI_K94=R"-%WT"2M#KD"LX/2W ']/$)SLRUYTY[EY\QHD]_1C+MR+G_Z6S[ - %,$
PB>IR['M TLK-%'BF*@BSKHO.J!U\8Q5.+DY92_+P0"4>R7VH4W  QJ&*+QVT=0 _
PK"\EK4)C]$,Q,:G9_\W=)8T1A6RIWIK3,"G53",Q .8EFY!5T33+!!DM1ZY$,"I'
PK1_&NX%M+R)A=D$>6>!].-8P"M2F6*6A4WC334R^)P2+X"#MVN_."3;@CCS1.=3>
P3%N=>E#Y30I;83 EG]U IL] JSBIH[5U\9>$Q^4GTCVP,K9,ML"!O'P[P.I,M,=J
PI"PI#7=VNW3\+?2?ZQ_:,,(R"?XG1V.*7F-\F@K^-'GC"PVNET-@]M#T/<C*[X%B
PV^'ENH-\&9)W39^FMEZ1:(!]=. 4B?GAL&CH0&\1L]Y6<WU)!JY&Y]M^].D-CSF^
P(Q/+J7*\"GTTNZ5$Q^OZ0/KHOED>%VTBIFZ!W1?GU,'>Y1-X*;6YL/NJ'3-*:1<@
PL\R#E$NBG[P6\(<<]];*@KM]O=5IR0"&&G6-Q_>2)KH[]N>$SE^+"U-#*7RV/)VT
PHD(:&?C#";I&? V8>L262=8OGSCW[@:C^Z9>M=4EM84C/>?>8U<7;WVSZ$</S*@>
P$/=;@8VS)JH0RL%PAO!^_^R::8V"F7 S %T'T@RPY'^K3[*,BV29;/C"??D9PCD/
P>]1%9'_A5JTH$?6((9I)+;C30JIO'E9;]O$PQFF?5)N&BFT,N:QY2[?9@;.50'=M
PKGO9]M(;=YV/@JIZ(MN4!!6/\R$FQRG-_V"_B6ES(F]KR0NG?F<QZ$<!4/L8XH 6
P.#^R72X^T]W#DDS"YM4\PKN6=05=2Q+>KTY0;XBPL#Y1R+W@>'N!A=_%V#Z!/"BQ
PD:II80<8XW4D"]$&E=4%_A!JT,G+Y=<DZ_1-SS7OS3;:# Z24&/Q(>CR6"MZ^]7+
P9JD9)O1JL"6=,TQ*X'7#Q+O>NY*7]J+(3B7S?>3S:9^B^&5RS8?VD<ZJBW\W9!AP
P9:BUF%3--$E8544I2WE!5KJWW5N^K<;<3MC ,_T](*\'OZSJ)(W47[\0W-F-7+ ;
PF7"HMYJK-J,,-NJ%0)R*XS4LM83."Q"X'FYMWD?"H]\H@D<S6(B-W\L[0HZ6DA\D
P.<>3TF]\X2.8X[\2EGX/+RX_5G0YZ>%#;EA>T2'$GB./I( 6@QQRFJF>IU0Q+ZK]
PM%\O-;0K$&VB>VAG(<7'P9#WNHI7)#PWVH!&]^?YI8Y<G#0ZG):/%]E8O>FB8F66
PI^3[@-9]CNDD')?CC88C9P&BM.\$J*P,M 6;CFFU$\N;DX&E]$"TR%Y".C ([VQ8
PX4<^F,9M>S(^N$O%:' L:[LH^;H%HO*TC(@%A. SRK9LZU468$8V+C.QDE-$LMOC
PI.JPTG:HY"FTT, C?\0P<RMS3T]6=)BDV9!3LC4RUV)A+2^]7VBX(WI*;T-X6U!\
P1DEKZH#3!)VY,2RV/0BY.'1<Q@FKFO-JZ\B4JD4E/B :+VQG8:JP\N&R<1-$L&A(
PE7_" FO=>48,DV>ZR,V,Z@$O,64I'&_2^*;<O9 J'GS7.]GU;UTR4=&725M-ARML
PVW%1V@[*_TJO:%I<=G, HL*3C8YU='2FI^ERV!;&V1ZD3DQ7.\@?&$>?#<E'?FJ/
PO4B0,LX*OQP<GY^OO.V,<G"03I*P5V-2CF]W\[0L\?LZP*)SL0A41EQ$H:N8"U+(
P$U H(IRGEP(3 P;,OXEL/:1CZQ&](>V)^<&#^Q&7D-T(!J/DRN-/WO>C"]]PV[\:
PH9Z_T:4VZ"J.T%./]9^.O-\'O RX"G&%M?T FV81XC*T78I6B9UP:X[6XFN:%!/O
PLA6%K" W\2!F%,0S,=\Y*,;R76=*2E%.+(SPK+,Q8Z*8#(-4$Z;.(7CW"QC)2B>X
P$B_-L6TGATV3CFW]189H"B3.43LKL8GGN,1R&D&N+E2E%],;,)0*72M$"D:]!\Y6
P=6UMD=[R?TK3"]HA/-\%&%0"6IW42!;&*Y(A12[X6[6\;P^9S21FLZ>'Y']TWK9&
P"ZJ[ .JB?SH]TZ.3(,6FI,GQW8& ,%R;*_QWPAB^')2U_+TLQ7"B:Y9N!D0D9."@
P4&*4FZFR >SX Z9$9LC^+XID."]_G@-6;J \#BM/KRU68,X&<6$KDX4T]5&(K)=D
PPW60EK.N3+EF 4(GJI!G=]A\OW;OR>O.4-%(4\&>YB1%EUAF5#_['Y:A9;07OJ6H
P#:<N0X\Z$#><+>C\9GWH?_0%%Q4 =)=Y4G9NKG*9^$GKK\XO"V$PJ/+X*VA7-+&R
P,#XUM26=P_='3:YTWL2]/X!\,TC^R;K>8F+<>_$99[)V;\,3ZA:*1'Y/0H:!"'(.
PU?1,Z]%=85K9;:8&5(K:_K@^;RQWBXS]<\"%'F=:[1F([Q.T#\ZJD24DF8DH$I;K
P*9\32M'F.STC6D7E__=X,? ;!64?D2A!["FG%!L.2#O@C:FYR\'RM./CVLM,&(/0
P:TNI^-Y9(:DEQ?]%DM#X"AD5?[RK/2/:S @8+T0D\@+?XN:OZ3?UC7J-W]1N&ZC]
P0 "I9MPY_O,[D#]4R8Y"+53ESR\@H/R/^'<_]=C.[4HT84'-Z)!N%&'N?. CSJ3>
PH&;U=S^+]9?JI]I\\+30,%/]KJ!*8-$$B+?R\U<8+ </(2]EYUUK<O4GA*GS3-=3
P#1S7OSUYZGW;JA\1:2'?(B)^Q18_OF"AS;:F>5MM= 41S*GW(O;\UWX$YM#BL\G_
P"5?!$^'#O!<G1:??VH[/?H%4KCHM!_KQ1NW7<?M6',^%97PRG4V=(O[77CN#AMAM
PA6;BF\1/;>_0Z\_IW08F?3#_\T-L*NQ!L#TSFC)(:X5::I)T)A-Y=(1*C5H3T8HJ
P2X.)FA_8+U<.O&V)YSTIVI^?6Y9<P#!2AJ$W_+\FH%,R,A67Y@+6Z:A^UO: GAD/
P%$$<30^3VQ@Z5EYEP8Y(/CY<0?>&@#:X>"*F4X_:&-LL1T-S;Q&P.ZA&6*0?_K2 
P8KZF2(T<I)#0P#\31^X&I3HH+5I<+B<I"[27<*JKD!*><Z8YRI<^>+N<I VX"A4F
P<I6ZR'O06H3>&*]]?I&!9LR9<V ]N/>4YL$E6RC.'N*R@TG;HK%H$TG\#=R=)AA+
PFD^^,>SE%R?:G*P8.+S*]0GM?V1'S"K*XM%(056SG?"N:B0<B[^<[MQUO=#'PJ9[
P,@RH^:N^]W;D,B[^>*5YU[<\LKIXT'@UWSW?Y&;]YMQ9>(4->:UM]VMJZL)4]RC=
PW @N3B.8^<_I]I8@J@&HF\53>@"@:1A_)F!BOL\IR:$BJA+(YE)O Y-A'CKU+.=F
PSPD81C!N!&_="IW@):&U0^.EWQFMPHDQ &FDM_8A2%;I\:?JT!>6/B\^$+!+>#X>
P%/\DMNMY+#C+3B79,@0C)9&+.YJAK,5H@2,N*]/@).6Z-1K=F9 +-=8!2)5!^G 1
P&5MQ[VFDV-_1F6B#P2YQ_#_QOT"/K(+[TVS+/[61<O4__R675'E1IZ(JVMMHRRZ7
PI0\3:#$F=\9IO<_1$PM/_O%[$@1GDEG8YJ/LHKYUP&U##"6=BP,5),%FJDU\\&=3
P-;N_OKK&<]W%+1W"WE[VI,XQ.#!AX69\AN4TB0R2W&9\B]7K EJN->%S;(4J(5<N
PNM>)F(XR)\ >PL<AU7=,%(<20V;2Q\O-@!>X/&[X<6D\DGU6H>O"YQ(>%B:L\G/&
P*0Y1,JD-U\I:96C@8WCKS=<9WO5Q6M"3FZ/RF"$WLNHCGG$F@#YK^8-\EB!FX,JD
P@Z.%M*->S'':;M76O]R2C@QP]BY%+$MA8J%%NTP;J"2LJ'4@:E5?1P)YE]:T#@!"
PL^J#-/"7[U26:NEA-0MOT4<LF+$%-:?I73C_/5<+T_T/$UB ?R=#:OJ&S8&,?OIX
P&Z$)^N%B=%Y& ;%RA;^D/U>*1Q3<&&%6 :3!+M+,AQ;Q1L Z]T+@#?E-7-S<>2^R
P.W<TV&=7>TAI <.JOL15SZ068T2TVJI0+NX',*P[IY5_>1).)0_T)WE'".5Y1@.'
PZM+^A(COU*B9A>\;)M#!W8BP7UO<#FUVO,I? C.;B[:HG_#HN*E'BM$<8.D"4>NV
P_9(]&L==[2KK\8\*$^,>1'ZF.Z\D&(@J+ YRLZOCE<Z])J&EW$)(,XDK"]K*X#/S
P)'R-!!X 6U(,AA_Y?LY)5?F??_ =3TOC]=-MM;TE*[%%+TJ='N ,- <1KTY"/*?H
P>C_C2G3%@#HS,\#%E#S#>%06OK3[X,PQH!YM/HZ0_]$U'%J<UVQ-?\X"7J2\<#_5
PJ+%&HO9HV?\UEF7>I.+WSQT^10?4"<?EQF(Z6#T)BN!DYZ=[5#NI);C*E</GA'7?
PBLOD&6'XMTF5&*Y.$0(+[FQI) 1B$BX0!T%GL1"5&=M6TG[(R1)L>%UN)G[M^U,A
PNE*$0[RL7^RM@4 7-+2EL)K*_.)<:NT!;@KDV_LH!Y./N7467]G0:(:X*__%-%(I
PDD(IHL' T.&X@6;/!#$N983:;C_<?V[GUZHYXRDM)G:9?/->J?6M!JD47?8!E"Y'
PFHT-E)?OI-KS#"@9=8)L!!.4GS(H -7C)4WM".IJ;0X2D$,:*^E02S_L@0//9G;3
P!K2_;81 !Y5<[7W,<C@$'AV:,<Y9SE516O80+*P]'M$!.-)D0.'_A_6AQK="NBZX
P(,;W#X3[?=GC9V&7]@[#FN6;1^-\/&;[,W#EY=6=(1.,3G[8X?BSU>!H???Q3G&P
PA-F9O9#1EZ)2X9XE6-YX;D60:7/$SR6)Y<L0;#3CVP]8- Y_<24L<GV#!/UY88W0
P_CYPKDI)F)&G:X),'"?R;7II!OR2:ISKJ!S V4[T*)=O1T!L5=KA.)^!>]-QI1D<
PBH9AOH\W_>/K(,E,;L;Y#4U!W^X?3^13W(=:^YOIC%%>4(^ED+7)Y9#*6&)AKXBS
P9"V&6A%@[Q7*&.-*\=T'7>Z#[:E%H5L1)QQ0B*G<JWB$X)A?*S"N: 5'O"0?.Q$]
P?ZH(_!+'&0,#U8%W6TQ6GECVHA1M0SNL"K%QZ>@CIWN)FIXQ7-L6=5;9F/$;FRE/
PV6:@O34.C-@^,8.*Z$MG=,_=O 5FZ?K>9=]';S;?&.SW-J=9$Z8 X1AZ24W*9'*]
PHC\KT57[)'[2_+O1><([CE:R.=GJFYZ0I(03I5'J_2G<J$3YZVA?&/JX5!I61B.C
PN4B3]9-11P>@GO#!6;W: SIP.H_=7>UM(F!DFO"D&%+<>XM3V'Y<9)^*N="IW+M3
PN.%NTT1I$"#F*-=XX+&B?LJ/L0TQA*1-M.>@@V:"NI-T"L]/X?CX;JA^&><T$J%Y
P%UOF]F3_>:?MTYF#=C1L*:[<M(DCT[P\LL*_WZF1^.P8OJ2A4#=4@V+108N7O[3O
PB0[]WA-G[0N+OQ([^NV M9GPMY9@DNA$.,7C'"CY?9X"IANI5,8V]&"[JCVZ!^:'
PV.D">#F5P_FU6<]0GH!D\ @,3CC1F?+"GVEXEIE<>??9:VN*.7%P#'%"1[I_QX:6
P'>Z:=SQ*I+ZDUO?U*>98C4&R8PL4_2U*\8A2RTBYR-=*VQ(0D1/<\. ?, MI%5CH
P[UQ\GZFVK09.+B$5$XP)C:(GQS]BZ'T<4D*[ *)[\[&:G@F<-Z_O&:LGS80V>Q;:
P0!.;H,?^@7@*9!UA7DG ,@CZ8]*QCIX"'1!JU@)6?V-[I @9+'#/*BC&"#U?1#[Y
P^T/[8)_[0K:_JFYY)N7;#Q. *:(R3$B=A(FG75'+1970DA5'].@8\+FL;[>> RMN
P<F^"[:2ZI ;#_UPG8A+V1*GS7[D@A1-ZN2/*Y'*5M : U.NFM\#LTRC>P^""6D6%
P<E@V8]E!9W' FO,Z?M?SO9?'W0UV34+KBRM7/M(8G4V8T]2FMZ^VEL$3'JNOI1_$
P<?/CNO/>("S,#]*;J\_4T5I/49.N!M#T*R9LG"K7UA&OE&3HU"O$<?,+]D:A>]++
PGRK"9:;',=C08,TBV/9)%ZD/T^R %&=28;>*6=0\I:3(AHW26H5*U@TN=/+RX6TN
P=]XP*P/31GUTF&X0#I 6ZQOU'67$G.* 8E09G2AQ?'Z#PC"ES-D&O(0-)U6TICRM
P*H0JB:V(GXKTSI--QH$M8'<F:<N'>D\*@P-#C(1+\,(9:2.L=6H&WDSZF8A/J[5\
PP"6]\9CM^-!5H*M%L?%5UO54X&K9]XPG+N%EJ'49'\NR)&+]6:@UHL/6N=E,9LY6
P>85TWFIC!R!K*2HM&C7Y>5 C>+@VY%S0=<M1[%+<!;$K)?99-<\L@?<1/)7/6; =
P*1[Q,7^V7D1'-!$B;$O&LB(#'S'T0S3U3= 8;5[&7E[?89#-%WTH_#W)Z#;2U,M/
P8*8P9 SV1H_5FQC])9[[VUYWS"]8Q&2*H_@@(;&6C\?UL,;JCH+)&X75<:6D7;X_
P)UK6#/T1F-<C/.L9A%?)?P1CW\!K5MG9F1.K657\02B_2_U_*#R]#SD_4$"!WFWA
PL'S-,__$:((XZLV$(B+D(%XT<4!R:_U31O9TC 1NXEF=XG-=W!$XI1#(ZNM4=O#%
PXBK2ZN5/.E0(.)"*NCS]! .[M?^":%=1+>-S10\L,1W2J6(P9W1X#5Z,J2:G>N'1
P+TG3><33^S)PH=F6[&0436U'[(O<@7*1H744'>\6G5+E&^X!N8LAK?,][%%B".B 
P)A':L>KKSGN: SE-?-?2=? $G/G;4U-+L+[PYU7AU"3[6JNE?2VABD#><<YHM.<)
PL9;.MFM=I6%7[^LY[O-#T.Z_)KMH>-X*AF2>/]V9/B/W6H.*$ 3(-)IGWU^C!P[D
PW(GF\E:;44)ES8W8I(K)XJYO2J>JP9E\BRL+=U$NY[@LM.&>DDP'B"4Z#++X6>EI
P5[WJUQV3#_Z5$[UO8888"&UD0LNT^<$^!:+OC8YWX]V]R:.Q_AT;EWGXQVKH?;0C
P#RZ)UW$2R$&,#_&@=;=VGCN'0)/PM#03F189NW<^*$*=6%*'[.))K."]B0*G/\]<
P3IKA-0#/<G]<73A@[M@XEE5FJD W#*-F0/^4@JS37_Q?_/L/F5E8  147G6LU5_Q
PUJA*M9P&60+W"7(-+'XAQ#U4,$R^35)6%EX(3DZ:[0>EJS%D[\:"B21@PWJV=6L9
P[#>7TJU+@BNZEN2+T QD"LZ$\Z>'9QU%6&UG]41GG?%*"/\TT/9<#6:EZ:A0)5%+
P]"D*%W8AP5.<<WE1ZFQWAGRDP1@[]3R$'WM+_@0WMJ#\F'?%U/^5*],K#X%PQ.&P
PSK#D,]OJU80I@"T04@X5UH: 46)>_B,R)(1X/62N)T4AO[!'V"0G6-+M< \ Q'Z]
P-(UI.VA76A^XTV$J*:+ S, &I[G[@A012J.07*7<5*AK<":E^D '[(RT:0:/'Y-S
PR>37;_\(:42, 4&7-X:7NP,:1;W&?W^#B3G8IXH2YLNVQYAT^VDE+4O-I'OL5-WX
P';,5&9E\II5G^%P;P"@]',L:_G*!#+:43) >MC,N@S]-72(NP?,4C&*L4V#S_?MH
P]PBG/78E^12)\E?0SEW>CO" J[^W]_)\]:KH+%K$0OK$H;>;?S#CG/<1N1P*D7/0
PD\\K%HFXGX[8<*\K1I>F*N\0_QPXLEYV&<D><SHG!0^&*HF\@O1VK[..I[P1+30K
P>=!?OZ0,=<[JP\-N[X#D?ASSI7GZ*^@YBWSVGKL7;_.*YA_/[$I(K91POJ&K.J%(
PLL,T6$G[9>'#DE"9I:N$/G! ,4M';W\LF-/GW1MRYDV*>!H&FPS(2A=;LJO@=!16
P,+4OZYKXV*0N:#\0>G35)EZ.K0T*04TEMV3()8SNKJL$2 *\K@NO;0'^'Z6^13TD
PQ4)8RO+5G8IA !CV4YG^)NJ<T!4"&&CY$H>K,$WX?GM2/:3E]^%. ?CQ^TW)E+YL
P$\5&>5)/A9R&5(GY03_Q5<M5(&U\) @PDH2$W=;!%9YH<&C0>HW=Y7.]%3Y'G909
PE];@*[=T;T?8,PX5E/7C=3 IL/A;MO)O-2=<G26(:FDGWAJH53Y:,E3E.4V2=ST9
P7QDHV1)XNGU]W0SX+TX/:A6V>LL(_Q%*(WOZQ"SZ"5E!)H7\ !J[;8B4)#QE\7GI
PQ\7YI(3+I"VAK*0!(&Q0)&;%Y,T^2N@U]CU[?'T(.3&^_^T*_O;:?D]HS:7A"+E*
P6$?W?4M@ ]*+-)?>1_GZT>LUROX3\?L_==@TKT]&>&K'30;YQ@3O?=(>&?JPA/1%
PO8=3P'G&>L(L@K29-0^))T3 (IN!2/(A@"EF(J67[&1O=<R%UK0>%=:QLUDBWG$$
PORK+EFA0HV$F#7?S+T8?*>C5@>F13OZ:=X%F1B;$+<3J],0OW3_24P@$?=.;E;XV
PXE\]=]^L1H9"I30NK!?VO9 ("!_\L#(M+'I+@084D7'=>@5]_<H5:O"\9IG3:6,D
PW^UTEF^"^.V/ES;#-AAQ>R?DL2+*"#A#L_]!+"LS??/@7T<WAY,>HH5Y7-64HJ?1
PNB\QM!>?VMCAD6U=@-](M[$B]W/$K$3)7:LHUJV63%4"X-,A60@'C#550OE'_>BL
PU5K/^TM=MP72T)-&$9KXNF_9#TAQ-B7L#B,_MH A2[T3'*6$I'_V3:RR:B$QTAC%
P548*T.%O4X:Q<W(S'(FC#A[XAC]CI(;I@1I),\*38<59M"8C7KP6]70 >W6J/PWT
P+5=;?XS0(QF?5%X\!6$J&R+0&L5KU,]22\:<($R%C @S#&O&!;Z!SNF[X9G\>BQB
PP'GX2CMF-C&D\LA:;T8#:#VF;QR!9_3Y*> J'[*C)!O5YQC\@'CK$K P+[S4WZE1
PV!03H)FX49/N*CMGI07[F5N8T>2IP*V#@#*->5M?@8M*^W/5A\&ANF "WB.<HJRM
P9K0X=DDFJ2X%E@A+:5_$!\D[57#!IUJ-,">4+6$'J7)6)FAOZIN>#C.*W'"TN6EU
PT$VDEQ*_X0%4YHYSY1;! FMQJ'V?6H-.O@+CJW02I$08O)Z(Q(BWLIA4!XB L_C]
PR+:3A79)!'F<@5.,.,TOP08^YNT2CL#^ML&<9]!YVKMAF;>>G5!39*-@*8CC?;1 
P/ZH_J"<(JC!+LY(H)E7:;A_\]<LH[!"8$\D"X3A=?;P/R*[6*E\O@]81^W:6#VO7
P\_K85J)[ZLVC*1#-2Y"&0]E0>T7D6;#J>4LO7>!Z]/*I89)),H<=<'RP7[$)E#H"
PZ-&'Y(R.9,>$X(V02\3\!XBI.WETJTVVZU'U6M&R$&,Y7/Y;TNBA>6:$L%+92;@U
PKT]?9)JD.3\-/4$EW?ZG/B%,216C195Q/3'63XZ* _.;#5E'N14IA:CD(886]7^:
P]H?7IG-@%#S/B@%3:*0LWESZ/TXE>P5,N(&%[NYL3')6M9G>K-# '>2U=^JKNGZZ
PV=[!@0IJ=TV+0,Z<K@&RG)J$P27-('$U/_-QU1K*>2"\I0OXS4+O>?!_^WBIM#%1
P]2&X]7^_+;OJ[@N6O^IEA=;5Z<#;-9@G_/+=O?"WI?090Z)F[0ZQ[\$%E2YR%#G_
P>;>8D?JG*J>"X5^V./E+@\C4D\;43$Q18=BP4\J!408-.&+9F?4@E.L&4L_7!OI&
P+]]MEJLLN4U \DWT>O%VN>LY\^*X$YG[P_:2\Q,_A8I.(XHN):\:"2[GI2,R]ND 
P!BBWE4Q?WLMP9;8WK_;I;(8&A@7%L4B)!/4<?A 9/UF(P+Z N=_092G:!ZI%FOLP
P\=^R_KH8RJ>Z.!4UT*/L%\(;;4R:= 5%Q?$$HN_%GF1E9YI[:R29:=_(4O9A5>P2
P)=5KVD.N;J52QC@U0N4ZX9OWKIM1=Y37]Y&:Q#@9:AUXJ(;G7&"=OJL:L@V0LG/-
PZF@J64NC<BY#C",F5(+YG14@)''[,JWCY/):DK.UGOID[729XI<^B95$T'X",)ME
PA.8,G;PG9=9A!W0ANZKMR(7[$^?8BV;-E@R9$4HLFEK8IG4"&_V_3HD:K,P&AH1D
PLGP8DR7F"=$63X>L1:?OP1VJ.# <(C+30^285QW-A,D4&VAGOG-WZC"*)<K?  /6
P=CD>+?EN>E9"JA$-"O=C@C11G5J4&"DP@DUV=MI>O?P-2!O(B[?=:CAAS3Z8GGOG
PHYJ#^@W+),NY0Z,PU%323N"RI^+@)07*+S(>(F)("6G=1$8&W4GE%ERD*G5'AV)G
PQ#&1Z&)ZL"C]['<]M,<'P.R6P;*I68=RY>YRE0!/=]X#, IH\ >K:7'9JA&II1ML
P-=HG9?BJY'D(9<4<&6%MD=0?%1?%;'UX)I0VQQB_LW5UV/^0=05\YJPME[NM7>'[
PRA-#F3J'<C-BT9\^PVLFXZ$5<(QDPQTH+(R.)B?&AD5?1B<TC5+F.?..*!LV4GV>
P/VHWHC<&4',[I@0/Y=0ASU<VG/ZO:&PE-%WKL?)YW02IQ"U$ ]]^Y-0RR^N3L[YY
PAIM;U_T<VU(]"SYCN,7WKB0D4 U_D&2 /O"D6R31FGFP6IVY/%P 4T-9W]92*Z7V
P>V(V&*"1K!R^W8Y0Y*VC*7JJH [E2X)6T:JB9\SX&;-.6\>VHXT<S2H^,S,<CE^=
PL89G0 ]H#F'\1U34%JBH:\0BT(,M\E!J!S_TG:79(G\HVP_=&YQIA,Y7CVOLTL$F
P -=XCY[DOPCECLPY\V+U@4XI45MW2V;&HW%7.H>;L[/\E91(*ED=/>Q_IM?A1Q=!
PI;^HS>6$BC4*EDPXM2"'PX\_SWPPCX03JZ F(VFD"3F?R*77>"CMC>='#5)IE]BO
P QG!?:^GN.%,>NP'MT^DR0 ^G<(P HT*OC8+6\<PRA%CF&C!W\[G74$*'BJ*U:J+
P:2QK?^6)Q/H5CG)-EN5/%I!.M#[]QA)%L[F)(]_%%MY$M"#X59<,>L6$'Q4$P0#;
PRD(R@' ->$S'WJ@U% G<M&(E(;;7Q:]Z'2:V0=[4-B+/UH?GLW)I7*7=Q&CB:76D
P0SBG5#"?8@AB6G)[&JDT9/T [F%7E6"7#7</ WI(X=I!6P<N,&S12ES+]"7)$FOT
P/LMI&(SWGBS+DR0,><NADZF<4M%!L/&J]?.KV$T>HL]$$"0/6JAZQ(S55Z)4ONAA
P@6ZGA_G515H]Z/U)8Z#\V"&RB)2SW)<6L!2&*8/YBG&9"M=).+;X]I#2WQX:NB2^
P>9#!9I)E"1MT.9VJRT[UXZ'CC:/K&IBG01!GL#0*,RRN$".%<$=O."\VW\.NV/5@
P,!WL9K\7HYC>:O#^/:W0YB3I%1#^B1^DD2Z36I_8!TIKTS0\K@F TH]IGL2H5NB]
PQTA@[((O"?=W@?IRMG0-9HYOK["1T;NG">+9B1;' \<,ATD#=A"F#6"Z)C8N5+#8
PN2IRIUS*N[PBR64%?5$%.:BU&8\H<;^47'7QNS4U!A@BC'P=7@#?<S( %>'I3Z:]
P_4*L,*C2>V#^L#HFUM(.[.^EI;'X@F6L^>(QZ$[%C^>FMH&]N<OU&<.""D:CM %)
P"UQ38'Y::RZ]T.L=ZN!/?I'PQ*V >*-*J" %:]WA>HFC/9GM*]^W ,_6GP=H$# U
PQG>M@/AS)PMU]Q_[UP/=G9KC.L<,I=-)- TRAM_57I&HB4$^0E7:WWC D^/Z?$!G
P2\XC;B!GR(/1CD5-LJI?T31J4J46RZG7;524>N$04Y%S,E"U-=;)&")!D)E5I$3.
PW?7"H<,*H^N)*ZCCBH8IJP[*Q<$M J"!0#2;#+"E5UH*7B$\=M+*!W"JR&9E1)OK
PL*',6=T\W&M],\'R0\%XX1,O:OH6]U\ZU* :2DN(P*P>UC9"85>\XR\4-M8]ZHT9
P?8B"=RUFW_K\.[<,=Y''FMRZ%!>M!)723P>N#11EK+_0)GPRH=R.8/5 S,B[J'\?
P?_MDQ_MO<3](*@-O DA#91+CC&I$54(=(KJR3H),X2:O:MPMEE?W,\J6B1/\L[/?
P!63PDL6T_ "ML0OAP?L(>U-<64>L22[@M4MVM5WIFH3T0ZLK_FH$;:_"UOA*2%[\
PFN/?"[ B(9.%'-TPMVR>1BET<NV*23Q=ETWL(+A.10B3]V#WJD"9,WJ[>$]YX$DX
PLU9H;'=FQXO9S%9F[%23I)2"I,/S"95O/U=8+W]77'[0O,>DT0\RH^!&5;Q.R2_8
P[!-JPC+Q+5H,6Z:-O&7?$IQ;^'5&[G&0S)3I=A8XAG0Y^Q8Y-^>7F P4"S*43OJU
POTLNE?Y3M>("FD>F;(/>X^.9D90[:5:164_;SU"6(N#/PJ<W#!1^3C?G;;U )WG=
PPCTF@,CG/A6WGRJ!\7$L7XWV>4L=78OM_(0GWZ]U6-$3+A;$8Y2SZ;Z@W0!I5MD)
P(79*/.16*+['=09S-CN)JER:[RTA!'"(B(<S)?V&]A'@N3]<FS,+(W!G)R5R!L+I
PTB>JRLVY<1$@@_[;$:#YO.TV,+:YP1%1*LL,!]ODX*'7K4P?@2577;5(R28PJZS8
P?>YSHKTQK12G>>7C?BE$/[_R[<H[I6(@(Q/ZCQNN9 ,@.KZJ ;FO*>82?N=%)SD0
PSQ"UJO69:(@.I]QJJ(< T]6H7XI#YZ,M1V/R6IG,\<+&91+^BLGV\<36,[\= ]%*
P-8=#K>CH*J8:O"&H42^G*#>V,/:V.GT0<ZT$.W!X3_P@AB8>[Y0?^F-9J:T%T@8[
P L0;D73@CKKY3>EEJMY0FMU:5K$0484B!4$TII*A*0 OJ,+*.!X/Y=/JE_XN3^ZH
P[00ZPL=LQ/STGRH>976']+MGF0[#KT=M2K6(OXYFIFL5IQY",^O-'W8ROYGX8/G:
P@/<9P1VL][,5H)C4R7!%=UC197AU: AH*DY$7?_ 6SNT:EU:P;=&ZP(?CFL5<Q#D
P27&G/.^T=]Q(G?W(Q%3G(2ZZ5VV1F9!-L[7TBGK$Q-7ZY^@J#5C4(T-;RGFEC44N
P?7O91V79@_B8PW%>GCB206C9B"+<+EO<F #]6H+'  ?*,R$@^MY666Z7IX:=R7 E
P5D7^=WSG*^@K7P9J= YQX+XK=B2;*%_OZ >LN<\1",^ZZC?;9.))\K"WRC/THR2 
P(:/L@Z<)[ZS36%F0PLU3JUL EMC#D&R]3DBP?XIGJIX6G\@*EHGT4>>R63?R,Y'L
P&FSMCXD[DE4&@P1[MQIQ;-";]_H>>(J@0@,2[7,"[?L 8"E[?U 0WH31=8CVU9#W
PA-3AGGZ N[/M0;F%B$PA$Z+.,OKW"4C\;(V%R<9<4T0RB]<]M/*>GEH[FD*.^$G.
PP)-"ZO ,YJR=E:: #6:#D&8['1D[TU245LHU<*BR<SY"Q42BVITKE8KP/D+1W^%"
PIZB+7LZN8_!-H5VU<J/P_Z9I=R,*#_O4%UM!?!8EK_$/<>;[T'+N#[]7)2SM'<Z>
P9+-;>PP4V$Q('\E.I4.<#SY/P6=?%RGIH4=WLW\NB:VO?MVE-5RS8S%ZGUD@;C30
PG9?\9T;PI_KJ@'.M3'ZU6/F11M((,)9-U8$D  #P(E)7%Y0EF-S'<!([5?N 6,&H
P"A=_,-BCT'&BF"@)%&4YNRB5R4+;_*<"]@HY:6]?(@46,U@I&-_?ZH+T:)VPUQ01
P :D*28[4^=Q952Q+10^^(*I[>HY,-O9_>3I#/TFBZ%G#,6W!.D>!#SF@S(8N>>?N
P>9*K-/(LHV^2A,X^)T4_(&C['ZN&'JQDK$$WB"Z7-L]T;3T?T+46[D("486>/\]$
P@X=_5:12TX71<YI4'D@Q K=QPN% P+>4-$[@="1MFGYIRE6\EX#]IBH6G(LQ- ^[
P^%7<1A,>AW&'"+*L!NE^$M2?Y% VJ;VS &8VTK:N_7 U['HEWN^I_8 J>K/@'ZPW
P0&#7^.$=ZL+D9>>H&FCU%/V3[6(/:O9)LPV'+*#(9*+?S@-R"I-$A4FR>DJDV4'2
P,4 F9A/YY3P_R"$:DH*+8NS/7= +B5P/2S+\U!$@Y<L,'Q).F;!8'T*BG4E&($%4
PWV4'P6Y;$5Q.EKUKGC/ C83,$;&!T5N3-8F<J[S,W<@DH5L1.N03:U-[01EO([R5
P>KVT)M=_628PSIE]HFB 2-$W9  $2-$:%N.R9R2BW![>F[0] -<7"5\J=8R@*:3/
P9K)7S\HI2C],-"C&)"YR S<*5!DU-(KUF\DA)*KV0T%9&ZD(4[**IFJ'^6/2GL/>
PZ)ZK-7LI4&:,@H '0D)V#?\X^; -7$V/GT\M5XS'(ICL,6 29X[..Y)\=/1?H"(J
P*Q!X^9NE1K-(0" @C:YN^%0$47?ZS5Q7.47 HGS>_AI%]&AIK:X-"M31!ZE?<F^#
P-0KTT=/?<;,4^:6CL)*Y41R8JF1H<[/"L0];;BY9O&7LG"2<ZDZ<[+OIU5_'#:O8
P\2[?]Q?T:2%S\DF0S<TU!T]@:"@S WA>R"+53()[#&0TG$YO-.O=7AB&M9G7<Q9?
PTTWH, W=LCJZ, M/[#E**"V22[TYX:4;D03*_-[*.9+Q8U8-L8(?AGX4G='-"(S?
PY:JRW#G(8E=)L-I^-Y0**^IX+OUV]#H+"8!"A;H+Y4SK(]\YL6#,,2*K#:NV6.^<
P=P.$\\QZE/UP&?UQ(#5GI^K^:"9Y],7GXA6N@?W\=P]N?=H<ZKT>L^PGH#47G4T;
P^%5CT&OC,<CT+S9+2WY=9PU441/6E*<:\1R*)'\=LZ?9Z>9SEDD3JS8'B8Y*8_N"
PSA:L5EL'NVJ>*A(:.61D0>?'%JV^B1.B&('@@VAZ!;"3S4TI43"*A6K'NLEY@ PB
P#E2 S[5CKND[!RE+@RT]YHA'JCN#2H$EK(%4#:8E"B5TLH]&9\(Y[FS"<NY_UB'8
P:M!Y]6,11I=J>E!;M:L,K#W0/=+.7PE3?R0J(;'Q#84@GF%9934XCBMT74 W9(WJ
PB5@AD6*H@M)Q45B<UQXSB6G$WVY&4:]%0;K;*G]HBGA3S)"#KQV5KGM3IN:Q\00%
PF0\^>7\GG7_]1IY*,@^:W>]BJ8,XL._]'REP?*3V*HPY#?,,P*SZ'G;X#QBW>A)J
P2QGLB#$)F]%GWDJI;%" A<V"QE8'3 )^D":R6;:-6BQ/U(4KF1@9Z$N0]#JK<*$/
PS#_^C)6 D-\X"@""?A4AZ:UBX71*>0[XJ3(@_).W0<XL$+@M-@V=!X=2(P0AO$0I
PO*Y2K]/B<1]NBJ]M;Z'\N@2FXTD'C+=QY0C-@'00&7\8-/5HKMG:<)\-"*XN2FDR
P:DJ%P>#8SQ+#G"P52!T,_2,,I2:?*[8.::UGRJIM^^)%:L&DA%G"[)0J"QWP \3H
P66OX,Y((1(^*&)4KR@4\4C^Q3NP51=&A X1IT)[_@L_'JEJ0U"N5[K%%BP&N0^,4
PQD15#7K<"7-#[4TES,144E8$S?!ZVCL9Q#YWAR>,F%#J.[8\3=O9]V^\D;VR5 DX
P_MH&UO1,;?C1C$$="NG^UX[ 5(!=^&2#GWV".I;PP',]8I$VLF=CK7Q9H/QA3N?=
PV*D0M89TZ6@VJ3K*H#$()ZB[QMGKT0Z[')?0DYQ!N8?P9=FJH( VOZK_<2!F#XD*
PD&_0-><_)>R>K(U;DH)7K57P/T70MG(#F9+=1I$Z,"K4ZS'%4#CX\L(/J'8(E^F/
PO]FJJ$X@A1*=%0NCYR!41+9EI_P,@$936NR@)/ <)?6R!<<M(*<Z(>DV278LO=:0
P$/:MJ!+QCW^SPAV'G#;!^[1!IH!ELLM/PLV B9/,9'V):<<$D@,',0R#I-KKP,<;
PQ_(H8@N3#)PW4@V#I336G";(GLB4IXBU-MY=5DVY[V__HV*"T'A[,'==)<-:-,QI
P6G-'#+#7#=ZVC\$\=ION%VQAP@?346%R%]^RE4-(AFK!O6A)\Z03Z1>22(-04*8#
P0OQ/\!'Y",S@'4OSG\BGA_+=T6=[CQX.$P_U'E?/0\TQD@GCL^R8^B*I*6;'-0_]
PD.#Z>TS=%'JFCHD<^6!OFO_](_EA2VO.K!9FD/0YX8+N\"F0C-*VW9_IJ"OZ7G^4
P7:.9\)('D-^TWJ!B\K17'2U6K,N=BHZ=OWZFYU]0#4)<6?>7Y&^[="Q#4PL)"CA[
PG1_^Y/3AWOL69Y"<3R38Y1&8PHLO#<LV*H6!#VI5[K(GW9 2T1J]S-HF24?P)_A4
P_4CZD,WT,>A6?/IERA8!B\HN!)FMM?"7%81@/O>]'TUSP"8,4R9QVB%:S,[OQL1K
PNQ,?+(."6]1\2E*ZLI3\$Y1;8_X)3VO1G$J>IIZ8EK=M+97DX,7%5!!=133G<DB"
P4@AJU0+NK79GYREB:N^T>9%\=W-[BS7!K=_=9AWN@-7OX4 :56%AWNJ2*KOX!'D/
PPI@)Z$T^%P)<E[OYVU3(T5L!D]I7^(T?#C= V[9,HF>.843S(QCCNKNJQD+'NR.A
P8K4QUS?.9R"#.00$=3!:,ROZ'%!\Z@3.[;C:[Z97C3<#.)28D9%T2%!AMK?JFND-
PV'7^\_ZG$_)S0/@1.5M(^SF&-BE,+MI+N+@F,U;OG\&$+T$E9[*DZ='2:PD(VI\@
P"RQ2]#7(<])EP(H"KO["S3+5#GY]Q07NMY;(5V?81+V&\GIK2CT=FEI4OKWX Z>"
P/#KF,T(IBKB2TN++>F\7E(LRG7,O$5-:4N>F'59/]N=1 LH@(P1&%.\?E:<HJFBT
P*+_SE/P$A!U<A/AHX_1OZ8;\X%6^D0WK,ZR%H5L1YHH0D :0!E<%$!"E";SS_3J:
P)\E1F#%;L]<;C[S;C>^.^7F9QE)W6"/026A953-X86(4[._'HDX "#TWXY^O)=ME
P) .F9%J;K" 5@1%]'FR5SUS/I\#/C'+I)UC13_=+UQR],_;6&KMF@2'9;+/&O5AI
PH^S:7.X%GBQ/+7[\4^*7^U7:N^;6EAQ@0'$>8ZUB*Y$)MRV*Y=-M,1)VTL=31M^A
PH43CK!&L"0?K(C-;5_H^C8LXU;YF,"9IO1:Z+7=SY<.Z$  Z<&8K6[KZG'[ILUFG
P17K.)=Q A&[SA=,W)!JTZ-YY]+Z)(;@CQ#HB_!2EG^16GP0<=D(H">M,-EGP&D(N
PA!)$CSUNA\K:ANF4O&7)-Y'!>\RNX2NB!?$Y64PE"U6&S?:;Q$GG/;';/(5JHT O
PX)^O1'<QLT\>H-LX*7VIXK+VUNNQ;>91X99TDL2L=M$&9:_C*_,$\(AKLC.;V6PH
P7KM#)-\MM>+JF:7#Q1DHO!?I]@]4;5^9S;6OCVGN/JF'@HKQ!]^8<X:''E(.'T<;
PW9>,!$5X?LVR;Z.,'33^-3_SAB J-966*7'KRBFB2MM:Q1F&^$/D:A[P<L*5J@A;
PH3CS$-%[$;171!R8.(=&X6D2&*OK%EE.&NVQ;7/YEO<G"#-?^,[$IS_]QG3/O2-8
P^AL)2$UZ"/9HB?OM<BC7P^F%WFL;\:_XVMF]\Y4BW%,YR-J(U<(/\0K/7N'O_!O2
PF(+8<M[(DQH+9G='(4$J4,@T!L<7!'^!0[% =(GY]VWZJ9Z@](U95+',;\YTD'>H
P%FG220Q6+2OJV1T>UI/^UE;:&#[_LCV*?B,VVRFQS\) "UX#U@0\[G0U]X&/NFN2
PL10+" >N<[-8V4IP;%/H0OXS2ZU7<TF$7Z/H6S#E#(SAR_U;HE<=[L%(=_#!8"6 
PU,.;<7"ME0GE\UU5HZ8/^WK0$2N'W9R],FEP?+82WQQ_"K]'BF6%D?KA@;'HB3"-
P1DKK6<:I$>50B;J@;IZ* 0Q#O!-(WU:,6?W42G?R:"V&Y%,^Z>.^VP=@_R14#C4K
PSG3';^LOM"]05Z2%A$=U6)!TI0/,Y*:XFNSJMSNQY(Q07(FK(&8C(!+=O&(&[^SF
P$"N^\OT3I*BGS1DKR,N$,$^!J1$=CKF?6N!+W";[_+F(@\KDU0*</03H&?UE"I7'
PT?4%F!X83DG1/N"^J,9WY@0OB:A'NZ/,QX2UDT??T4HX/ 6CZ,42DEX**VQ803H<
P^%7$I E3/U *R3X\ZA6- +L Q%6X?LB,Y)3R:.HGYGB\TJ-(TCNO#,TE]Z#UA.J9
P9FQC_2FA4/TGF[%E8.QU5BJ)K?2U)X[^/1>;<D"\<TIOP+A U9?'?0.(<J.>:53T
P8<C$G 5AD^>&)#E>C>I%'M:W!X=]T/Z=I>8F9O06P9WY1@AB\K<\.U0\"#6Y\5:(
P"&%WR*2R!/^D2'5M=/WG>B7D:9)"**!")[1=CN/SZ-3>#B)C.A27Q0!"'AH2R7O3
P'(TV-$0 \P S=D^I[6?_<Z:1#6Z,<KV1*;>J*AJ#:AV>.,SX;\/H8[C&)=%6\02F
PF%7E6N5D2Q,6WUQ:)$O4%JJ73,+O%5C,D)@X?QF/,*"+G;6_2R,1N2T#@4S<8<<F
P3+>U1PON*LZZ+&S,3,V-KDDD4Y4*]/C823TCC& (AV3@KI_EQB^DGA5EO(C)[!^>
PSY$G7/?K^2.I8!1M7L1=(F'[:<!1AV/M-//Y->0) 4]Q=7."0E>[AL5=$Q&X5)FU
P.AZ%IZNK-I4X+IC&L_03(=]>#-V/6+0%"1NSB]E<3)RF<:1Q!YNZTDP-4N"WF5@2
PPOU!F7L4GERVIQUY:3O'7-X+K(OCYALZ,T!<K6*VO1B%1P]$.X' XJ7:,'6$85BF
P+'XI$B))&=XJ*X04\HYN>G'$*40%,P1C;U_*F")INTD^3P,$6\ OMQ:4NI?C47/N
PNAK+7G9_SKLN1^"QT(^9O_<!(9>JG^ ]KQ@0'BS^&T*2V==YV5CMM(34!+.*O^*F
P^*2Z"IA][9NZ=XC=:+BNH68DUTY,%I :>+@AH ]9M>]=NO@]1-@]R=0F<AJ_6:CQ
PY5*S%V*:#ZG?WDT197T30?&$!CU_8Q$5-=<?G9^RZF5%FKEV=1AM6C84GI86(T@(
PTGT\Q%G+12:#-DAS'-A$POZJ5 NCC!MPBCS#963?^X32$8E4BJ7U.#+8<-N,PHA?
PJUC+>T#R"IO0NY]Y-XGBL_/WTZ"5\_IX C5/ G S>7+K1K"-*BL3GY4R07^\0\I_
PKLE<Y5]2?&:DJ6=U@45IQ*F(&O^%2.G;"\I7AH\L647^Q#Q *9F,"#)&HBL?*2(B
PW->CA4+IM4A:=/ 6)ZDI&%Y%+S>VUW[7+R?GP,7.K36H* =8)U96;D]J:92H_6OY
P[!W9PQJJ=5M+$P_"7ZZ8X9XYU!DZ!!0._G!$R]T:7211 YAG#SU(^?4'X*H!I@WC
PY'_@V1:?)?^?LVCZDTWO]Y!;IKV@G-8RW>G/7H):['K+BV.P* _@X%T?D=AL]IJ8
P1?TEYE9QT9-"J0"@BET+@;?0!8-U3]( <2B"Q\PQG <T[^KS\IWL\<;D?88\RNY_
P$]#,C-51K!C6U^2(.36Y^(NB.06'>_,=7? JF (;L^2JZQ\*KGOH4YSLM -!L=Q;
PG?UP_-TKY?-ENL8)Z-SWN6L76KJH]S.C@8AU^PK];VNO+VW210:/>A;PIH+TT)<$
P=\%N[:(\N=&02[ ::G?KSDXV,6)P3$R^I@L.J>M(YA;U;(BG#3;Z$*+\:(55"_J]
P7JLT$?;K8^\.!VFFLV/O_)<IN"=)EIC4W*CV$>_Z8"+K.%IIO+:\:6"OFCC">+QP
P7("_NJG72C$7--+62]:>Q#FW(E#W_\[NL&?3/YMV;>DFHU,W)?>ALFLC6M(#9?(X
PKBWO!DD"$"%>;KDS@!N4>WF@":N MO_8!"*D^I<=VDDN,^5FO>+;N\;H2JV>W +O
P+\T*&*UJ;)>:4 CDD[UMT7KM75_@T!LR0LFTQ,Q!8V"6HS"CA-,2K;C#*WZ23*H^
PR_224,2R--A4<:9:P7XT$<=/%AQ(',_,=L%<2+3 FG$1O_L?$"$SA$7^O.G71$1R
P\;A?DO(O_+@E[FR>V8X[5Q$4FK>Y,R@RM5B+O".W^960T,R,]#7?R8UG X?#?&VF
P2?<HB8BZPLZP @5EC'V\[_!GN<1+#NA<<B@KZ@ZC O/)KZ[1?Y_50KBSV@3UN7UA
PY26E>D_;G]VL6$L7U&[NR'+2OR_YS("OR0F%U2*DO\&YDE,Q?35&!NBB^#C 0A/B
P]-O?E!Y#:H:P MIL9&AQ3.@XI;8I$/MBMA2Q)._*]2O3J^OBZ'CW> M8D2LN%G,]
P"4*Q M/N\@]18=:!**<32Y=2=GL;NW>SIS/4P )31K7"<.09]!,,2EIX4>=B!R6=
PV5?%M:C]FEN^U,)G[:@?:Q.G0SFLZ\J_XW8UUUS>&'V&P'P9]60FPH#ICAN64<)^
PFF X#1G^9._G.XS%5*$12E"29'<KI3V5]+\2U]>01G3Z^>SP0I)EUGV;<=+2E;^Y
PU3#GG&GQ&FZ^(-WM+IS+946K5TQ )@'O7 F$6(29(P!'#OC^3SJU4# !-L.P2.=<
P/,K JBF8N&)OR$TN_('!3>7AW)!OM5[0X9=?\UVJX8?!K4<E(CB$RP_LH?\P/7E8
P'\%[!:""XDC$G6,=DYZ_4]4G#?A316E"2 Z,ZW(G@)H 'SQ$A_/TK-:A*\D0+MKS
P$J"456X^^P>RRXB]7&#?(@WEX]KH@@$Z97XCOFB$":A2,4,'04Y96#H6-IGU)&?I
P#/VN?U\BOK?#7WO%(D(ST.6L/:'SR7B-5HK=!(_/DQ0:IPR'6(J:6[I0J<@)!P:L
P#*- +B7OV;FZO+X<J,YC]G?'?$)\SAZ[?'Y(S.3,76)*T?A/\)>  MH)D8N<$51!
PDV\Y5C7?\GGK+*^H%33Q !64>$5@7'V#N$CB29:[B"+>Y8\2SLO4V=9O2"N556:)
P)G[V_CI4$Q%N%\*/)TY)*0[MQJ3V&_KEP7IXY_7NF\^[?]Q]:X=#B8KIMDS$]F+W
PX*O@*@,3-V3(C<Q@/RBG&4??&9WD]XF,J#.PCL\Y91HSR"<.4O=MG2:RV8"&*_J$
P@.7)ZVF<,@>2/JLQ5RB1WJK-6\]VF#Y87U9_6>S#D,Q^G=\<[S?:O ,A,%JC5R&D
PV^AMF,:]NB%XB09?Y"5$F*FV'6HQ2[BDG;#=JG:"XRW6LWAH))4-I J@T$//^"R;
P JO!V!)J5\PN:SIN5S/.J-6C0+2Y;817#'5FN46<J:G"LFKW?^L9N0SSAZ1< W%<
P23<:WN,2B?&!]-YO_49;6D8VNP 4<!IE\&TA2"6WD>Q-7<+@"@+&"R6_(;!5-S7T
PUAR*]G/"NF?OFN4>A[,G[>-%BY?7-ESZ[(OZ[1IL/N,;!U+A_O7F["?3%PGIU;<=
PVPI3$?'?4L86GKO10.+4 I1>(,35WQY,((>A O!7*^+8C1N9<LJ+/W_:C:=IHNCF
P4OW!D*MGE,$B?*O6[+//3M'XWU7=;,F7;:[R*>!(@OZY-B&C;"HO\5$= 8NB2=3_
P61\?$T%KS&AAC<^30H[OC;F^#1VK*4YR/F^PG,69T+L5M]-VF)HP-^+7GTT8JL^O
P84AP4BL33B"L5>7];.6*!KQ>^>U C_2'DA#&8_ &\O\P$!J9?/Z*.^3ZI%13X9$^
P\["O8;5F/$A>O3^K1?RG"!8&T)GRW3]E';*:;_Y5_B/55'_ZVZBM4J/1X7'X\2NG
P08K7)\FSM^&=$T?/FR3&<0S.MTN>Z3Y0P4H]V1G <_N4Z8JPIN6:;1F(YZ:RAML4
P]!=%%\3S8L$UV2*+A%?PZN^]B!U#U#LI?<#C &Z9<E88QBW\DNI5&,$]#Y<9,7A 
P5H_J>O;9DR3Q("ZU6(CAUA+! W+Y.NQ'L$+D3R /%E_1D\=YG<B)DKJ<( #C&^_]
PDM\[<3#KDT0N;(.YFX\*H4?9?K!W_Q*W:[FSFHRT!G#5^VG 8_/5 K2FIXXWPU*5
PZ/IE$\KM-K=GVMG'P[0U4I.R=I.'LQOES4R,J7Y[@E-=054LSH8LG_A$ALT5PY<>
PNG&&LT2<?:*5?S7GX?0[VX#/>-!O8R!,A"U32U0C)X5(2LY]7,TRV9;$&DG(B_;N
P+=./YPGO9C='?W[?.HPG:; A:R1>MND^ +:B_KP=FR!'T%NCLOI*IT+2@:^/FA+3
P+J0CE(ZOIK+M3F(B(+I("U N!9SL+W6I#YCYHA]HWO>%6-KP[#CP(3UMT2KC;">S
PH)'2?<\><+)"#=9'S[3W'(-Y_;?/G JK-K2-U-%54,ZKEPC* 5NN<N45X70+,0%'
PAJPQR3$$_S$>7(+(9&OUW]T?)SL#AD^!('?IS2&2]]9(DS0N4"A"L%5&_V+@#$L4
P"J;'=2J),;Y+3+2+)ORH)7L/C4FI;C^)Z0')A["PIJ$HKR$M2*8?)RE(8!\RO!Q@
P\K2]V RX4J.U42CD!KRF9MDW%S6-\?9(>^Y>N5+D$2,.%YRGL8#_W;G U_HDY.=(
P8/!-'?]*H[= T['JSRA0'(_4MIWLG: .!6I)SW";BUP6&I&'9U9"P6_!2@#7#XZR
PJC%%[!'M>LS4\@LFBS0O9_.!LG,@/MO^8@/"IH^H$+X0^9^KU@5Q+YN7V)TUUI9*
P."O")IG/#H>Y7'H$,-5*$/]''%,=AF=C$>Q(HTZ^61=(4J.= #<$)^+%>54(C9%S
PS]).,3D$"E2[)?GV5MZ&\:6J+H?K-[98A6U7MJ)+FL-4E4-JBO,DQ*H+E*7NEC#^
PPE#HY8 #K&%V3YQ\H$LKS:\0+!KBB;:3;!I=T%,[7!R2OQN9T;22B-@3;3_CD:$P
PU::=1H!6YZM069$M47MN#;FD[\9"L7M@<=^.[D0KI%4Z=HP@U0>6NIFEC^Q!3J /
P2A#H7@$U\K']6[_N))E"3C/#:^+>N2GOV>GDZL(.=8ER3?!%$!Q<^@A0'[W,(\*2
PKO(_+OW+9Y*3!!-)O"#C0S-@BH-MH3D-<*4R5JW-)YIGF67[SZM)TL25:YTRZE1J
P^&_E1MASW2]!2VEL_UQUUI*AXD2^CR,QM@9!ARVC/BS4MXK$/T52+<>8&%ZQB?84
PS+\ZXXYI3?KIT'V#>A]B]E3.*J<+3.7?7CM:*.UY$X\W086G+[E"SN$V1Q\YB'@(
P;A-8[3#P9%N/ZUQ5158,R[6*&2'3Z@X,B;7O+^RI0YT\1/51"#"FC,Z\N_LPBO#,
PCLF#T?V(5S6C;JA^PPXQK\+9,AN @%X:,GGS3&DAB+D?D<Q>>K16RK910/SWOMU(
P#FLI%*B0Y!.RPP;,"#^#8GVD1&;9]CB.9,ZPG]+):JRUD7MOPS7)'Z99L3US\5!7
P]N47Q:.$&KX^*9+7=-\!@HPRIO3 KBU/)XY1X6?^/[0F]?)#8QWU'K*P0B;=45)E
PGM2?VO7?4MYRQDE3$63K/N>38'<KGX?4+0J[Z1CQ,\I-+%^I:P6HLN:AT 6L\X;M
PW'^A@;#3B$3H"GF./#SU%DM"%!:@A2@#H(0>%(>>V3-"7XT^!Q8& B#[RI6=O!(*
P_ZE/1L\VN505CG4Y\U"U4JF#I6/+I_J(:?^M76OF-@'"=YERVTBJ7XJ/?^K:T()_
PKR&/?HG6_X5N:(<T/\X.-PE5Y>_WJOA.X?[KM1_<:KGJO1<_GKP(4R5VD$V27H?F
PH=HQ;^_^44N[ V")5DH*82C+TRMT G>U%&ZB/P7&Z@"(Z>'UK[(^Q,I?15XLUMB7
P$R/RN$AH"EXUD@B%_,1P48;0)>N?+^IZRFRL@;@WM\P8%D<QB5D<*Z=P7Y=NTI3?
PCNTD0.^JJQ;1 &<XB0W,(!^B6C2TN7,'ICEURQ?QW"/D2J7C0>9I8^):9:">P\CG
P1M>X_W0,EXYR"[5SY3UPER9>U2ANM;>P5YN"87M<A<OKK:-V$D2]$#B8Z10$,0QZ
P>LF@6/TH!$T,OK_!;1 NMAK;_HHNN[7+-K^)U%<BR?7;H1O&,.%F</P I;6U8\6%
P[SPIS'3BY,B*HYA=6VTJ""(N)X S1A\OEN%2B<&J*HECP@58PG5*SFRV%YS7/*%"
PIKIBRS"3U<TVV<#72&V$N7Q5)&IHK;P\A#Y[R1>XRT:/-QT-A!JF'L%AO^L6Q7.(
P11DK"'Q9, XIY>E-]LR!.8#Z1,6%^6N&3:$2# 5H%TJF=<BO)6'GDF#>:?$)&8;W
PJQ)^C</90:QZ,F@TXHO?_P-[D1[OQX=[W&^YU=5!HPFZ9)EE+;A-(7COX93\T9CU
P5(/1I'868_/,!9,?*0(R;XV6[E3[9NF[\_A!J#WVU^;J/KN>H3XAHZ6R6I,'."=J
PV],M.SV0?QRLWZL/7AUNH_1$4(N):X*^-V:%C-@2FD@ #'?HIK?I[D/<V& 98:FG
P7X$X-C-<;$@J[)5<(?>^ < <Y0E-E GM(9+NH,7L $;-)(X2N6FZ,3C=3M1&O*\X
P!&HD)S&U"_9NK(58.K]'I+7Y\%P$&_[Q##,!]\A&ER.27KP%9;$UQDPR:]\B*>Z;
P,[-!<>I&T5OL:.7A/<#%._DP%TBA'_L6VP1Q,Y\"! 7G#NS8=<3G-J+[0@/,:5<,
P;W7D$W1P4;;&? MA  Z2#%Z75L) =%8+T^URQ*$:-276?P&AJG9@U@L'9+^I<$?5
PMD''+1 9=%/;!HP,D >L0F:WPE#-BL-GFE[#*?#!Q&,ITT3,__2UK5[>9H(5.#W]
P\)?/JTPHC\)/A:C6_M8?-<F&1#E;?;:^P(@,(P=V.$#QF'6W5/**2ADT;SU=[YL/
P,2.QN;0Y>Q]/,0%[!WE%,Q)"]J,QA*+V;.'@"ZD9"+KBHJSB?EI@=U89#KAD.-$E
PA8[P07ECE3SQP=F\LNY?FNP-L 1VPK4CXK!*(@7VH;OV\1-K"/6'NEO /(_STIKN
PC-;+D.XXI&S7"_T_ J1'5QHS:YKI*W6[@C46EIUG8-X#2-$.L/0OE *>KL,&;\1]
P23>A:REBK(&7F.W+ VFZ[!RG%&6C6=T;1P^N[S0V1I86FP#!N#'=2=_SQ)B+ W[E
PX6>7B>S3B=)(@)7U7[<*K%'^XD4\Y]DX:$SF(R# EA HFYB\$OU5^@#QFX.70IDB
PI?!)Z1!"1WQU+(<M-_!XJ&*]"KJ)5LFGOQ>3B6G.^4S:1G\/(/%]6'EB>IJMWU:O
PR&06M*J0'+SD=U!4.E QX2YAZ3N:1!'L)'$&/-/#K=$44[;_= ]\!1T4Z]>C/W/_
PON>["%6>AW79MTM9G^EANE#?6-Y0G8TNA$%!:*D(U.]IH8NA@_FNU%$A<0.MC#$Z
PY)HFI?\V>^[JQ[$?7D5@.H0/',[B'=TG^[MXD#\5EY2X'9-5RX-3L=%C/* @#O@;
PG4WLDYG.Y1WP94%R3UV3!8"L:1X,\%?U:\0'A^+ ) SWL3#PS)3MUDR'(D.65#&G
P$O\[*JFA3[XR7F2HU\;<65'%M*R0$)J,KEO??U'3#@9^2);35QEGV73EP\+A>)TD
P :T!D_N36EQZ/$D'+4Z4UJ;DI1VC91"V</J";[/TRR>-1C^CYXC0H@: G:0.XBSE
P,%[E>\*$+07$MY^P-QW !U'\C$V16J]_89W.[>#3TU.;<B0_=XV3\<["OC"$U:Z6
P,++YA^^DLGDT*USEML(6_C8MZUGJUP"8=@9W%W53?:[1[8\'@Q>Q_E*HV@9'UP1^
P95C*XUYF&Z?R\XS2ZTL?"#\'TE]8LO9K^L,OIS&0A%#R94@=,@ZT0"+ \I]CI!J+
PN&UP1Q8R-9.!XK!ID^1OJB<.T+.9%!B3%?:2RX=<^4!,OKO*A+=F2/OO-ADU1&VB
P9OA5KI=EUTKPT LR<I%SR [-DNO#>V6P_,]/8RSW)DF7Z&RL<^H4+5VUU=JHT/8V
P'ZI=6T['=06:)A>PKSHXHO824]KNP=W%"4WCA+P(EEPW^+2H.Z\]M,[DT28Q3__(
P0J VLN8Y%JPV +$N.V)-@<]Z<CGE/45I8']E=^>(J+2#3&20*0"U2<;9>AJA^H7^
P\&FD[<=5CW"^\>B]M:.DNG9='F"K^=(%*.AH=HC-:8<+!8P)2M1OI@E"H.,?C6*4
P <0!5J_[VUC!X3(TO1QRHO?G@?@H5JNE31ZHN7"O90*@=UI<[>&>N6%_E3KB@N^Y
PS@-UBDIJ:U6OW4!'<)*QVA(@';I&2^0/)$1=>S9./T/D&@D=GHXQEQNH&X]W5'9Z
P^+I*!LIJC9CE\WV7S*D'=PHU9(]P9:@HY68XTL#;])$U^1Y/=2R7RH0\,+[%E'UW
P\.NGYS-=KH;EQ,,(6\^M!V&40/A*N]H.;TD!ZWPB,D'>1O8ZN9WZ/'UE4:R)7DM=
PHD'2 1Z!MM3M&W1JU?+X)KMF*B(A:NG8)D'R(ILP<X0?B?5HQ(D=L]FO.I&P8FCB
PN-AIGO3I)]5L+'P%_V4$3QA$3$R[R>9$QIE SMJB_IS(V:RP41=J4SL0-=S  9?Y
P8G8G]A:4(9M^../TMAFPXEH6IB/<U!8%YDM3J1%5H%+AF[4&\\&OMZ0-A]DS+R+,
PE[T)_N/X76+0QHVRXH\ZJ_/BB.?%TJT&EAQH0C/.$W)GI9;4U@,UZPT7#(T6G5=,
P1H^DX1*C2LM)^B(UX -IWOSD5!$M:KALXJ!WB%9]EZ&>*PS8RAVFIP-$.TI>J7N>
P<;)4BOQ'SX@N$\4PB2V=&ZF]&I=3T3> %*0?/65 ?9G;8&RJZ93;&9*3,#*M3L%V
P%3F3) 2P1BH7A@Z\/,F@'3YJQ6<(D'5>^N8:3(WI;.^@?7B%L3\C 5K/)K_#YB8U
P(G- ZKF@#'(7#$\&5QIFS,#,!4H99UY_B:ZWKVXAX+O"GK-J]#^6Z%;XA!HR._#P
PT))&M0_53O(3F_\!^Y?*5CDMNUVIITL^KY3!%IDFG28>B8-3\&P6=A(HC\W#]9/B
PIT#=D@YV+Z:?&#V*J(U^M;"I^!WL!R7$;AN-SO8$QEETTKVNQP[  7 ?3:HMBSF=
PJ<3+&7)VUS56@VL6,C*PW=_]>8 OG  0,U[$90,ZF(=(CR,8ODMX$*E;=MWPZG=%
P;7T1L6GK5Q?^#8H54$23MRW_YPQJS]P_LI!L7S7-O)MKG/@A<I%FKGJ<3:]P@ZF#
PJY.W>Y"S.U(B].RRR&RB"0IC,U]DW1'$!W%>1/&&"B+0O% Z@VL(0.\:''LLC<CE
PH4N? ?@ZRR:1ZU18=6D(2V#FL?_#/9G#NO)0\>)%1S<?G O2L@N-3DN0"P(G17F_
P7T<8A3AN^'^\P/J*'GFSY4DGTU6BKZ^Q\.V\UIO:4*YQL E0=KH$IN5?=Z%_.L5K
P]!\ZW0I@\6-@'A+#A]^F$%O0J*@0ZK9?6F#9!@S^!?GV=J]G3-I 7K"I"X_^O\01
P%OZH7;V3\BT[&37Y2=4K7UL82#>[IP(WY^@:!N%VSCJ6C@I27&',#TPW#<^G!L2.
PD&WB,;5^GZ1S^]_[HFH!D_#LQ1%=#+VH3-H-OHJCD/ VMIQ](G?U+RTY%!F;Q?*6
P<Y,U4^TJO@"8C)!GJ4_]V"Q]0:\MHMABT/;&*=PAV+G>6QV*C)76197[%"'&U3J#
PA[\P=(T/Z!^KM45,)MUAY6CII#$=K@PV&J'4'K361CBZM>A$JN6SF5Q\W5OK/]$X
P=M] W+\D/^R"&,#;6ZRJR$ Q*+;W$!V$QV-.J1PIL$DR):O_N= 4I.+U QEQI-U_
PJ4:,"9%:;=LBL6'I)0GF74?V17DZGIX%,H___;*LNP*Y-\S4N*HBT1$6WSD=MKV 
P#GLO?<>(!F\,Q;U9Y'KX1E[J<@CH76!GCFP9>SP$\1@GS%_<.CSQ<N2TJ[T,00SD
P&72DT(W4+NJA%A?-1=+[.JFZ9G.@H26<U$/HI=)6CU-A!07!;:NXI/( D,1G_PDE
P\&Q'1UYFVL"9UVT_I5C%[F.YFM,=P%]7%3HY4 >3JT[>B)=L&AQ@43TM$&A]%;<J
PW9;D%:08[-,JQWTPPM'.TD@C=S-@NW[?'=2"!;&K8E$I /5$;*GL7E5C!#(XQK6-
P*?S9C!CF-1\C"^NY'\Q_X06LY=D,)7+QV+8T!D]I20<*6"25>]#?E2M_VI(F(>J4
P]' 1@ *PS&6LB<DQ&<W=.2H^I5YJ':-"GVB\VQV:,[^I;IOUI+P'IUF(<0W$[8*Y
P;H.K*,<SQ?S$\4I_L6BCF05\I]AVF6&J!7D9J;P3![C8N.$OB-=!=NB$M#4620:A
PZ?1[VF?KV<.Q.:;Z+&> YNT/8VHTH>[36=K V/J]N-@(R\8EP:$WV1YE22_=T8<]
PY@P"5O?F.[H'_X;0=3/E:';PXG)=DYA;C1J$S BG1WBZ[G_098'K'(XTI",D#VWM
PBFBKV?;J<-!(>Q:-KO5L,,OE-K FKM^BY;W?G$R*SO-.NPP[B'C;WK703&TY2W^*
PPR@Y1/5#4*"AQ^%BZCZ3=K,"4@SH<3<&K:8J/49 (@QR)Z,EK>Y!65K[>T!S.^-3
P%=$&RY\)7O:*+K%%>Y9@GP&>03JNV,4J\X@]\%0/*(!ZQ7MPA=)^F/8AV445\3'B
P!N5Q'J 0DGR?P:[^+K!0%OWO6S:#?"CGD6/Z!(]KQFCM<KQ._,K/*./]&U$=ZM:1
P7M3USEAE[!#>8.#IY: \IU.,-P1WQ!C-[N/0"BVM]?2QZBEZ7UGS>-]58(R'2A/G
P;NH2@1G\<. "+8MAW"-U#5)[5-G,<LTPB\R>3#5WRJ,<U!H4[W<9U.05^-'=AH$L
P6>KC;$)[FPMN@AO?5:.@:;53_5X\3$CNLIRS.K">.S&!8C[>L;W8H9G/>[(9X LI
P\7@N'FRO$DC5=:3>'94D9-3=9?6>=COO!5O[SPU?B'I)_59N !Q:PZG%*?43'A5K
PC8MOT Z(6O6O9_V)5)WZRO@@6[2C5NZ5?AB9]:YZ1F1 V;73X]AID9IO<:2N8DG?
PIEH(F[H/ \$D.'_$*.JH!W/1_$:/NU<U"M&F[Q)M'EGQ0@4Q+JL08?5NWJRQG8.K
P/NK"U-K_C6).8E!#OEHZ;)SZ8NJJ>-L\:LE*XYJ9NK>*]3P'U;8O.!T23[M"R0!*
P^0^^TID:IB6GOH9=M,G3\BDBFTS1/OT=-6&T5KF<$CFR[TW%&(I%L)5L\TGZ0&4Y
P$WSK3U[$LOQ&/536EGVV>"\OOGSAADD.#M!U'--\[\4),=,# 3LZD]#GE4^IW:[Z
P37K?E(_YBRI2A:] W:3,UY\]H?R*JYP8IKWP\Z]/&AH!?R$#ZSNFTT)P/O>S2Y@Z
PY :(DFJZ_MHVV)A4+)894BS>Y9=1T!WCT)& ?6QHE3Z3AA(S075;)<S\T8PX"NZR
PIVB2Z153'P9T6/"&VRX9*DKV+'$^@QP-D=P^..K27=M$$@_9F (L*GNP&GV?WO$4
PBW##7)\"5/TT<7=E8-A[GGSF'Z0KSIOV7R5^AF?#QO38Y232%CX5Q(-(:H@A6%8Y
PR_0M3-JAWZ3TY[H]H>-%SD%UB.9TJO/&9HMY#GUE4"^Q#H7X(XD,@:JYEL&J1T'T
P!+G\\;\LZ=([]?']2YTB ,R>["L+1QVB_"5EH%\2;#(5HB6RWJ\^2AV?GC:BHP\4
PD#8VW 7YNS>2L:&-$*(J_V[.0GEVN8D7C9,N GYJZ1]C7))!R*OZ#+!7J+-%)<DC
P,%4[HB.\)'/SG8H[CG!1FP]2[S64,#[/0]2\J'AK1%-(:W#2SEGFPA()!O1L>7@T
PO(5[Z[6<3*\16?7<>W($VZT$POD5Q3QZ9U8[DH6/@Y$F6 DET;&FH1ZFAF)-(^#?
PG$V0Z!8ROUIM/4?BFNC$%UB:J@^.G[.2F]E:1!#5Q.CE2\-;>?&G4; -7 4[-Q2_
P:D3&,BT9L1\*ZF!_?<DETSD $84_8-9YRD^,@<V-RZU_4-9VHBTW=E97+L=X-YFI
P >A=3>B=0+^\6LLWEAR#%:N(XWU6Y7Q[]$ITK=G(C>P8/\^M]#)OXK2&+L 7 HGQ
PT9+@13]6WRBGE#"0<KKAO@ M4_!Y5=8X*TF^!$8(XASF9;HKJ*[D9>?K/"NOE6*/
P[0-)^^2=4 *,O 8.2^H&] Z9VAC)XLDN4<D.%"M4M*\<Q-[---W\DB0R4ST^2;,6
PU$48W6I('-^?\@WPL#V.@?FC&8I*S#W[#S[1C3KF"CE6#?KV2QR5YUSBK67,74EN
P!^&U@6M=@')B<C?GW#P]:(E:#TFZ7B: NN%HI_85XT9+0]@V/!P#%&5&SLUVF0@Y
P@!L'$/Z&O_MF::@&2T\H9IG$)XSW80^AQ'!.W ?CF@16SB%0D1B/U6^?[X4,60^[
P=+V.NYD9Q8IZ!LT>7?P9=M""2H,WNYVXX:WJ>%+7!R1L= _<'G]B<6)CP_3ESYYG
P-#'BA"9+U'.CHM T-\=_]]LS!BVP@P2G_=94@S5[U8PS>.KL&5SP3Y7T3N-3?UJY
PN*^LFBPI/X7;R#L;*K^[(NDH86;8,"<I@4CC9TQ.C'C$^Z".HNI0*1@/(+YN(3JY
PR4X8[*B'U/Z@\5D%^Q:70#8+:&V+,Y0A<7PBH3J:;;U)"X\<KK4"F]S6-:<H0R1?
PKMBF1IA_L6K/SR&.%B:2W"3( 46V5RKV81N]<ZHS_\);Y-:.*O^0^&E'D,Z$./\9
PB"D,3O'^7S7_>'L?2^^/'O\5^<?T0&-F_W^M5KY(U,3VM6Z8"E0*PU2)L8(9UY\]
P5T$#G1EXFJX_\%8!FP@N3-E:6;K_MQU+5D\7<WMCY_46H*.G,ACU.Q#XTTRX 73>
PQHDX&>+R0%R)*UZ$[9ZP_H:LVT#J<<?ABC9EY--&>H#5MI++>ZJ'*<Z\5)?%=Q(.
P#MI[P+* ?# R00"#_9,AE<JG9,9V)&14S:C(C+[<>YK=,\:EEI!/S7Q=]LS:B%2A
PLVU#5.?L;+QL*MKVO7A#7?!:2J.M/I?*"SNJ,8*$8@T1RL0UOA,B*QH8F8E7.0;K
PJ:]Q#)X(@S]2\&!+#TE2%0:4LU<=] =T8\_QX-R25?(($(\3J8)E?H4+WBEZ7H]]
P\=U;"=;7R"MP2E3$_ ^I-L AO)2BFHYR>E_:7="N!F+?A=&D^PQ<V6''@-K""(22
PC1L]:BO;*HZ^0^F,:3VW=6>A96 JM,'5,>Y5'ZL_A".-V(7^D:> JUDU?[*8Q!"4
P+QYER2'G*,2RX4XREE@5&(C:R8#UA+;E^/UHF>_F590D!TP#*4[UFN_2<?2FMQQ2
PHP8@GSEX-Q;L.?8GE"GDQ:P2/21@#)Q6:)3/E@8'P(0'Y$WER<NES5!K2VQG'#?L
P!-N,'1+[IKF],;3L8EFJH2MOESWDZ]U\/#7@DTAS1'7@;YDSNAD?O<D;=WA:!E*]
P)M/@"'MD]2,O[HS73P@F8)1^M>ZI:@4])_S0D#VH+ZG590K/;B+?]U:V!L2.[0+8
P?4*3B9C)OG5XK?N@R.%:M3/I5$N#DWGZ !/UE9S"(:(.W"_'B7.&9M0XC165##>,
P)6!^Q>;&OI1>.47R \6414=%+>U+58PU2\KQ$D(WJRN9)O1OIT1^V]@ E@M[D\,8
P,6<GS8MEQVN&Y\?(W*--)!\$&'"PCE>(%B:_ME;_%A:+HX)]QF3'003VKYC;ZGX)
PB J&FQRZ16.P3;?7^&+6=($X_H2TU.+HSN9@WLKR9S7W'NP0]G;-YU08 W>6\G1A
P9QOR^#JZM\Q##^(X+J;"E';?4+E@;D9_@W*$/"L_QB),<6?NI7_)+Y!;?A%RN @Y
PT_$1U2RW.AENAGXK#+ 1=@M@)WE+[7O*Y!I'(_&1JF;A<_W.5SWI+I9KO"FHC_09
P?-KM D-;*K'E-@R_ZW291R4@D2FXM]^?PI)_8G%,#@L:&>M7N@I1BH7\>[@>8O+8
PYA:F!![&=95(EU),8+;0(/=B\K^Y4D,C.#J")L9=G(]$XSJW."<SFDQSF-0C,6^3
PDUR_A]A"@7%X ]?>@1N,)1WZ<[\]5%<X92AZ#BEM[F3-%O0Y[,TS2N\@Q9T!A3N!
P(6^!4V"MFZFY4;^Y]3NN,"!7>F"QI]^SZ\Y1@?0_HW)"V!4 <&?A@\!%,P>Q*3D)
PZ4Y/&@9!(:).F:]=I07#]S6Z/;[G,/"2"*K/C!!,>Y<?\I^*3IR3?PQKSW>+_U$7
P2UV9V1C6CBMY=4SS7'Q]8VH-OW4.,?@&5J)LH?DA6<Z:U$\%<;+=(K#Q=Q4TO!ZI
PP-SQ56%$F'2C3<BB@%^1^[$CP&N?)J#/VFF-]F0E(1U0/U5DKC2?AX;ZHO+_%<:P
P>TX_=R0.!A_)C-39>F!6&G(6C(EHWT7&L5:87=%_F$&J3RV'I SS/6NP$+#(*\_[
PN]-=# _APLH0)XDY7QTMR(:2<@^5Y59DYNY.L$U&BV (BG1>IFIPJ_!PE3 HC4.?
PI48W@WACUCGVRY@YY6_!"H',MUZOCE0Q%[Q&Q8[_\DJ87^:T7VTIMD_S(Y..$A=9
P':;T^,8Z "M6(UW!(W/.T?%_6A1!YR1!:*_]N'\!.]KD8V7GYS>"C8>*@K&ZGVZ7
P>H5/DOAEN:[C1G64;^:#N68HSO@U+D/,5<,.X,JYN>YRK@74*5Q(3A7<><. 6[ <
PAVM<)W?Y4E?ZI;[5T.A3ER&T\98R2_:K:@RMEWJ\$WY<;_^02V']34@+6FZR(J1L
PP.?"']:_IMRW)7E+7$]JQ<$]V=?ZH0F;G]9,?O/CY?S+(L5+PLTXU<K\0M--IE72
PN6I"Q=M^":$(BZ&UXP01:_SNV!L1/G*L"DHS"$5[NL10@O+&$_F; MF@L;-] R2O
PS=8Q200'J;\!-"CY;8@O_U\]RC0AQ5E  C#PKL[=5:J<(@KA%/MVT":\&RQ#FC.:
P--3*/5<O;"><O$XAC)+Q7C[2 B4T6)0]R^,+/G%LJTL?,MZY:^[HL[AV&0 Z7@:>
P]0S\'7B$ R6T6]S<7VJY%0<%IZLBEZK&FQ@;64-QU3AD&#P-)<U"K35[-5V%2*CC
PT]D;M/;KWGN!Y@P")S,>?QCNH.U#M'7C-<V!.IB>G2W ,. 16<ML"P'GY#-1)6&A
PB!^TO62!5O==,5F?Y&P.K-%E.F.0.?Z8%J@U.=CEWXN9':P=GK#!Y95NRA3J^MQA
P=&%-[?B^TO4IFJ.X=5L^6:KS+MX/<4GE*F&&9N&A(ABX78]?K)]C\7- P<'D4Z44
PCD<3 ^UKV#9K.O%!84F0<+ Z5/!1BQ2SFOIF$&$$8BS\**/%I'P[\L/.K)+S "Z=
PN%YT>PBV;,3V_7I*<4B*GUXPD;KT!"K80_:1Y]F2O8-@ ICK'Z)B.%<=B=3%9_K,
PV@H0KE=,AZB.I.("K8Q>\O.->_Z;P[95U0]*U^\(0.ICCQ:"6)Z<EI5N^8+?V1S=
P%*)LD3^#]UP-6+,.O[+H7>Y#_95_,ZB3].>LHU\OX]D3ZC!3W''C0]0G("D-&F(4
PCQ)0"F.CJ=WBK1T!6=D@+(39*_EH;K=[K-G34O3/YYJF:'D8I"4Y;7-\LO/2@J-S
PW$S[E&ALG<=92Y];X3X<>"_C,BZ;&.$[.W_S\2/W<$CVHS=\&YU'%BI0YO?+P5%V
P;T L0>>O_7ZP>G&=?<"XQ?[@'FJV>&U<@)/9NFA4+BH:O9R*, WQPZ]^ L%HA;3=
P)2E"7QF1%-RO1+'#_)$^MW\W@ YSG+LF\>OE@!A#<RI^93;@BYR-NAF(RR5BO+# 
PGS54D6=4-U!-MA=!I@ E&2W"2I/-P6'XQ9EJ]BSKN![=I2B4EK,G-FC%]%?69.;V
P&JT>C4<[Q1T\;\._2,3KL#EW!FK: \1QGZ:S!<3J=/(N0XUX'98NJ?87%2=0T$W#
P5$G^HGV,OFD>J$8,%K))3GH.-TU'V8&=^\1[FRMI&;I']V% (:VA8AE=;3:_0*9\
PIWR4TUJ<UN5!*PQT) 0F=]-N6I7O6=\4-4JO9<LT#.!XGR"J=QL9DQ@;7)X>@H\8
POX\RDU?=? H;*\7%/S;DDJ&S-K<M0NRD?U4?.<_NP&D59P]NM4),FY*)"$M.UW%H
P)J3$L<?=1Z.:FBHZ]G#QU^HP[?<SV?/X42)&5OS1@G ,$<,JWM>XDU_D"#VA' P^
P(B!'TG<:DJQ]JW,*>*?;L)@L7)HMU=WGQ!6A&4EY$DRM]B"$GH5+YD!9FU:R2E_K
P%&)8K@>UZD>SRS(/S9^X^P4,<+"B>_N*Y9*A1QVA\=!Q'G!33IQ2?*Z.K(&2WT$V
P>,(8Y6K*FEN8-_4KTW]JTB4GW.?VZR[?59<WG.UEF3KO=N^KV]R'(8*C?LU,=JH(
PFU\ZB" <PAXH:^\$"&,S\L4()&IXC"Q.7N3[TLZ]%6P88CC,]B#7K+./1PTW/Q6D
PD5*($]5)ZAQON'8N\ +DC;-BXM855V16HAA7 JJ>RZ9Z"KG).S5G2-^)X_$-8OPL
PJR-#;GE_C!D!E- =Y_4UR,!PVIGI^5,1 KUMEU$7 Y^ 9X?/_>)3]:$CBZYD#!+I
P8@P$Q]BG8C.$W'I&#HZ4C@&R1-6E05=9+'+L]+!R5P]T#D+C)M%K);?3[C4MZ6NN
P85X-!&FCM.I5AJP!X>!&R/W3 1D7SIV&P3M.:+._ Y;OJNS"@DH%"8ALW,"?#8OS
PP]"BI%690C;+DZDYQGW24=8<^(:K/+@+AG"OBK,3#O$1.!""7>+AP@O0R *AF -.
PYPK9$5'[@=E&;H;TG/EMUD+S?&D'=BAM;##O,S=HF$S(7.%S<JOB!P?2YF<V*[.3
PS\<$G/43RGOO<R*LH.\349IOCOR/#!EK;W30PN.- 9IJV4Z#SU3F_>,()TY'\^W%
PU_?^/5^M#Q8+K'X/LD!OH6\716Z<#SKM#6NVS\Q(3;C2N)8FLJT2_X3OQ4IU2E@P
PP^6UN\P_$QP)T2&C*F;M_%DO$1E)% \Z72<8HU[63,>%]>44^(UM!MD#\R!;J=\(
PQU@BV*:I?906KF.@&Y,</?]>FKOZGV6&V#"W?K+5%]WJG_J0N#91&=OVY0\^K('0
P-#);&E+LSU)PO5MO^R(?./$$>;@8@_5\L)L?F1 A3%J%D2RW"%A"]@"JB@*$!DV8
P@2XY8ALCE.%<!B8"\6AIJWO[(86(\RKYT;<6.4V,39DHQ?1K@])-IU)6$/+0=-7L
PX@3I].[ Z'_R8-$*)>B;QOC]USWS4S$'6:A3 _8S>OY]( PA04G<43P0&Y5$17H@
P#.]F"5S8*V(%05YL8(FB!A[KJ#1!#OLHB;>^CMW.:,:TJT4,-PO2SW>1WKX@A?P7
PR<'V$"[<8,1BH(ULV9=OG.F_XZG6ZN!!#]FWUUR6HFZT9S*O]T4WP0( UAY4/<I]
P_SDP/B"FNC1^$G+K8SW&B>"E1&-\X'SK"7$)O[]Q)^KK$8\,_YMN23\+AEX,^#O8
P4"\>FIA!:/>5<]Y[;9EWM$%@I727S5=D_P8>.1"6*&9ME/=PW-]A[:?7CB/U"VC.
P$QXA;OS.D4"0@FIJ0? U_,269-_KD*:44[-DGL5+,TN&[DV;1-R90:G QCM.BPAQ
P& \V'K5*PIO^-=T;R)#S6#X!7@;?EKL;[&6(P54+.HFV=;93STD/SZE5/X9[X]O 
PN9TP)L\K"_2I2=P+P<C4?)?45+. YG3S6+'U]=#IDH?9Z_?YO6 9GCYVQD>K1<FJ
PV8Y:)(H7C5F??M<&L7D*[QWO=S:%$WQ->+*L8%]N,1.1/]$^5(2D-?8[A."YIM8$
P'!MC376D"L=J_V+=GL%XC;+HQA>3 ?SVEH6M@J&8$M[*;_]\:[(5X1QX9@NTDW4^
PH])-</DW.9 8(K?+=:K^!CMVE-D'PEOL4$Z;1DUCUWL.SY;@IN^P2,M->Z>U^46.
P33\M.D/VI+18<?OUZ.S=_92];V8*W%]H[V[9R1_M_$5NA&;9/1J^6>P(MO+Z1<UA
P_97 8M/16GZ9J26XVU"+,("2U ""2-D'B27O>M-TZS"9!E;=,<P:6*;4X SO3^VX
P]EGK:F?1/](X#HTFDBS?B[Z!H)T?2$6:X"W+A+0?IA9]=-=9-5;&&@%'KDP]N^!G
P4-)\C0]Z)QEPU>.TL'RXZ(W<43-)< 6A9;6!,U$J@;!#?H<O7C%3U904]JWJZ+?\
P-?]G63_#Q$(#*:^& G=^9"4<T<$+>U#G!<?JFI%)(@U21 XFJD*Q-<XM2Q??!4X*
P^-H'Y[1[LO6+9Y"J="ZA?*JQ"N\B::\;X$-<9%98?JEY+:P3.5+"6 D@Y<'.+N<T
P;NS^'ETQ6TG=ZF^_VZJ=(K>45.W:2U6['JEB@,$G.@M-0KZ"9M3N0>+:]#8SVIE2
PDTL5V^1/C!H"["E/03"\KS4CJ!IIT6\O&]%YR_OG@&J*?)7R@XWBM>,*!LDA7YE>
PNU%.0P6CB7H=Q3>8Z5Q6A?0<6>?%#YK1=&&ID8I*3VW:1.,'L[S")\5XD@*T,:T:
PA+]V4#?.BPUP^BE^O0]JE78H&LYG2W% XCR*HH'D C-! !S3UVD#"\+IG=3;H^XH
PY5(S5&BH+$8.!S?:QM+L7.^3-+]NF6T*V3AE/:9F*MF,3M,RAS(IQ7T*WCG/(I=(
P0AJ/)Z%SZ*LS?;<PJ")D"%%3L1F59$AO1^7Q)]/-XSW#_ZJ@AF73%7!X(;+J$-_O
P<M"\;J)2.S^ 8L-=0A;0&5&-8;PNSKE'MU^>G.0H,LQLRL<J/[E!":LZM>S0$$M*
PX'6@GTQBI^JY_N1PJ(26[PM##CLREA.ESX8^X4_R(_T_7<OJ?4-Z'4U5E'=PW"K&
P4I+/U/"+1PY_? BXQENR^(36:,)2_4Y*E U<CU'[[JT/57BHS\(R**(BT9 =PCQ&
P@R*53@QB2TGN>V=&!@"%FL]\HR&--KW4S:L?Q]?RR^OFE9A64+/HCIG]_=>"&XTT
P"!,8(*N:-=F>#F=GL?F>YJUM*)':#5]MZNE9R.O1[I/J#7)0L8-!Y0;&LP<(?2M3
P6BM9[?$^=; CK2FY6!)\E!QB#1TG%;-NA^(G%%A=;_W"E+H,OFRA8Q!H*\'N<L-G
PQP\19_./9RT#J,[1.KWT:$^)H.Z15G^ON7.1/D"7Z%&AQN8^,-"-_N./MH";UM=M
PX)S/D&:\O8-,Q3!RL$1*L_ZD<+$L2F(Q>]"3:$63LB=@$")66KIUHI>L&IP1 .ZH
PC&ZF.=-UYS"B<U\.>5),-G6!U<*KMZC7J$>J;Q8&;8;O(O7H*M/+V&2-,"\\2<11
P*?M=TL]^9(09TSP&)-B2+X\]H%[K*@)YI&CJ^7<BQ.&E)E0Y\%P_6[R>?OU)FP/_
POE.5'Z=Y+&6B[%W<G65T8 ZJG:-5<C0Y<$_=/F)&NI'E?W+[,-XU  MPZ3G2,3'^
P8;7QRO<":,T/2S,/:_1Z=?Z@J:DT]:VF-EU;1G%'!(YJ MURVF(0TXR*"5?P<!_6
PE[[\D!_#_\,\@D,%$\::2P5!9%X0G=?U]J'(6N[#_LM6_]>"_Z.8G/ 7),Y,6ZF-
PH0HS>=[752SV4Q@5E?43IVU=#(8[OC@ *2 @&F%"=$2M>3S!9HRCSSXY)CFCZ%>Z
P&N-QHT&++WL,Q#4FJQU6*]W)_.$(B87TX=Z$M.-NZ#(O3#70+8V_SKX.W2-*Z^'7
PR#K[&V\;WK<"S@<8VH@B"O[#M+%<^Y=1)4K@)YH*O1)24%M:ITE"%%64G*K5"K(F
P _G4[# 5$Y<TF76XK'0[^CJB</;W+*QL19%802LI3] ;Y52\5*O%FTLHA IDJL0^
PA:1!:'K**EHIW9+*W4BAR&>-2-1ZAHQ\F)"AYE'^N>BXT?/D#7C'**30R;_OAW1G
P*#?WA#@A_AJ[5I&Z1>J2$*=$4'02 J] :&9A\39G>WSPZEK1R8]FA# 6Y2=]+"<)
P9KCYS7_!UNE[=NFD" AB96$ L0<O7PMKPQ&C.4+;#4H'+M8/RG^AAPP018O+1EE/
P+U7?$)5>9AT037M/.&W9\3EHL9."A=F*&+TA!YC/4PE>W=K3K0.L]SPMO19E< 8X
P/)4_PAY']36F>0- .$?'4;JU1K@* K;I<)_2ZZ:W88" L,6&[:NE0#.Y0C9S'L;O
P&C5B/,O Y=O$5.YNQQS]>J=XCH2Q^^B^@TS&#WZK5/IWZO MWM(*V"&JX9X$%:TP
PV9R]JV1- K4Y<F:-E95-T*DPO*2 4U&E$:%83W11MSRH&W2D$%PZYO%]#!_ER:2*
P![5;KXV4@ &[,3,RN#/M?@KQ6BX-D&H;BSB%%X/SBKQ1&J8A&J->S"0#_7)!ROV>
P/0= :75G/Z.L\)$4?P]]KK"EYTM\UD_5\]_47F6[@UX<+L&2D5(@A!C<2=I#R9R+
PT"UX7)2?;Q7YCA4Y:CAJH.2QDJR -JGG%S$$O)$7@]C?OS/;MUBO'J)%W9_B6M2L
PEJ"%+>_OMEL/#V-A1_QR0Z(C7HG%+DL+/?\;^ZS34_R'0)GBYSM$76+2:'WYOT-<
P+9VV1&%MZQ^_JB<X9RM)-+92B9;K7%DB2D^7QX-&,4V66"],QFZ%%LF2$&AN]@GB
P/LM14C$D%HBA3Y/UX/9SE&:(B+=1-P(]+OK FXRW,-X,3 /^.: TP46_XFI6:ZKK
PL/05LYATZE"^>O:MP/-L@;EE0\2@K1L7I'$N[N _!"UGG5;@7$G2=$-^(WA;,V\^
PCH:4[.[H[:L[:4HL'C.:&B7Y=;D?G$U;IGVV1T\0/3 7(<#GVF-$!?AZC.1@BD]J
P)RMB<VEJR"%\+//\R*N&SCDYOZ2#6]]+0,FG!%\3G%:21N-::S>1Y%#=!7DH$VH?
P*I:6ZG%HR@2R7S'SI,7Y+4$>QQ=#SR_YM(X@SH2'UQ>2-ZT<$U=D]7%!9%$Z(9[,
PR>?@W>@H+$X$5;[3N$RMAW7J<SD%%YX 0ZWYFY,\L-2G!.!XIQ @COM@N6!;:_I(
P\-VMZLRWK; 85MR#[XW??FL[O'J>[GF7"N!E]69(2GM+IEU0@-.[6EN]E>P##\W$
P2.YD?ZR[964A]E]JZ]>$( !XS%E]](\749U1Q,DNN?7^B<.0])Q-:HPU!Y!.[5-L
PBDJS"\ZQR(%"T>YO&T@2R2L![4V"WE& Y=:F#FY?V(@ H.@[\8N.<2=-\:OS*0P]
P%'WOTQK$Y/.)8SE_53#J)I&RX%:G*D/?0()%4* 7I)/"\P@K&Q1E^;3_NF;HE^[P
PLAKEG+[T#ZQ,Q/CT&VS30<_S+__YZ[F4_B]]0G8-7:]AJ7S>#!++'D753PK&H]MB
P=31,Q)LQN%:M221:Z^H&W/OT(^V_<QB=FX&[8%VWG)'@DS=4N1QXKGZ0\81.]%EV
P8"9^R8)Y<[PR"8A#WVCWON>@N\OY&4 MYHFC>$/\.^*UH!BV(1M;S'@#A_\Y.JQ&
PZ9]"LVB9BHO)@4YGQ1?Y@ WVP(&/(>"D8AD .GY\U6P)2T57,<9YNQNZ !@R)S$$
P.YV*TFM1;UAVLTZ,$1/KL!X">Z>FJP:%5NH4JDH/^REM&>.<D!!A  +.';-DC>F<
P;AZKPO-=,)%@[5RVG*\J% B]B4E"@QHQP*T0F5J?3#Z$D@:K<#O"PPF1 ;J(W%LD
PBL<X]  J<<G(A>O6?_<@Z.V];"<+SFLY,#U T(D<>XKPMK.*98A&B>X_3FK)RRG:
PRRC,C[8#83<&:32]+^_Z=;:L&^('8QY"+ONP_3[J*5GK8D$7D;<1T>Q([0-YH)T7
PCEL$L@DV^X37U'B97Q;BL\X(YOY@(OQ'NVG[XB+0M1SF_OW@X<GTO."7"KB!/4J6
P4M!SS+:*2W:)00>UT/\[U8;F1"+O"*^;$-4G*CN5J@CD@X-B5PJ11%.3R\R'K_4W
P[3J):X5(KS:(<O=9L!T-<45P*3/MGXO.6.\WT/'1VF6]L1.R/9(A2G?"C:X/\X0O
P$ONDH7Q14;(H"HA:7 GNV!SIB)8T$R=DP[SK94&IL]N-/0@*EJGGH)TXF0HERU0L
P>VR.6W":Q93,=@?Q.H$Z(N78,+[GYOQ:IA7*91,,-?!!F5Y'-TXY;514@9%!'6E&
PYS";5 $U>L66IG,4K+.L(F5)Z.G?^4#KF/Z*T:)IR+P3$3H69*QLGHD8GE+AF[(8
PU>[A:6U(!^GUWOF?<LQE4!IM. 'OH2N$\&N,U9.]TV6E6*_N-,'&6ZT6K3VW_DU/
P#[B(=XJ6ON2E;]N28<$-!P5/ 08_?$\)]QU=3H'09Q*QKWYK:$0\;L %A1&ZR(QZ
P4E;*$)_1BMGR/;HWTYR/_/@ S$O$Q6O? S=)D==]Y*>('*&B0_1TTT'7H% :\FFT
P(&?C[F=G@L^OH7PDBVSINQ<6S',6R_]7A;?NEG18=CM/0]F'*CNIK8H'UM^*]8A\
PW9"U*+9&*);XBERH^- IPL- EM2Z68Y&?)D&?I(ZF*'466S/>V 2\.;*,J>4G?UA
P$I3[)&$T7IE4?[(7W^H1GF08'"-[%'+UQ.9UWT9T4.<@D/I]\,:9!W1R3T(C=?:J
P<O\L\R]SF_0ZZ.O9(Q8'[FH5E 8Y>C]0YJK,F6A-$9)U!))[5@"5:?[^"#"PC\WA
PQ8(")E<&6E[#L&_!QE <C'?Q>'UCA_A>M 4T3\&>JV%TL+.O2@Z#FV=A9T\N)@AC
P?#&F9*E&CE)5P3MR=>YGC-9USY,*U!&R=.$NQO=\XA3=#"1VU49%R9AH#8(ZG2Q,
PRO*7]"UQ,#R@&YBKVTHZ:'G830QT?:ET#T=<I#_F0@Y +0X-XOO/8L.=/\&)08R9
P_E)28^=">.&CO8V#1CA^.DI#".#NKB6#I'_YM%":Z+R9:O0?!].T9"U!:?A$U 3P
P6MO,1=(R@ /Q>PS5'8J::^>D0 FB>JZT9Q$W5^!;A^4N8N54=:J1!J0!-SIC\04:
P7OBKMB;4*?\.[0M]> 2"D<?&T8J9&ZV(/ET?PU,"]O>HTA)SL#&U:*MUUIA_,2J7
PAMC1X9L0/EWI$;S^I@<-*2P XN>^D V\\(Q_,:""E1,Z%7L,?9V&&BF<X98/L7F7
P!30UE7?*,)@+>4D4GUM!K!&OWR!Z!OJPXC<V8UB&N7TZ*- 2P(R*7;NX5.-+/T<V
PVC2C+R+;&96V@FN(2!>V<_H._.+1$X774PL74Z_YB^: #'69HR!.72"U/P!U?X$3
P<#;&)=+/7[I%^K<HCZK%=UMIIS=X?&PF_$X;^'>3-G2Y#]O-W$$Y!68(Y4E7:C2V
P";>$(6U ;B+;6O>7;L-%]I.>%VPV'^G<3_Q$WA% Y<2(<5-7*WZ:6C<L,S_NA%0G
P-:8\HI&53P$_T_,&:]"#9XZP21PMDX2:UW!)ZC!5V$K.-'M9E_OAZR.NZ7=IX37&
P7L"D -<<OI@:^>OA_&B]@&IM]^KGDO,OD[[Z_XF7*]!^L 5+M<FG1#_:["N$.T4E
PAJGOZ^ 4WOOW.KCM=RAP-'#I>Y5=I%Z> N/3"=4M'.U&J$\U^. K;^H=Z)9BR%W>
PVIC6#.,\JHR3&G=FW]W#(WL*1P/>4<YX 3%:C$L1C4!^F!#20B_)$X,WU91$'K10
P,0JU,YGUVC'SEUI@AL)OJ0/?B+9]+?I08)#ZZYI61G+OQMX"O!=ML>[A+I0%"$$B
POO88"NR.1E0'1F"IT(MT.V\%KI9K?:&"$!XZ"$XBIA#(51:&<#I/OUH-29R;DOHZ
PE*2&3%Y#,0XK"LW_Q"0B<(5,AIJ;'(P>2-/KKS!\:BQK"J4KXIGM^%<HLN\?@<VO
P#7ST6EO:>=CC]R(\]!KMN*+:/,,;:LJY-&<:L7;9_1@]N55\&7N]M$-I;4/C&EZ*
P2U*%U9;[8%@,8DIV>+9*"40E8FB>^%>]F\[UT&(J."-C<PE![?$25]\(5?E?K6*'
P]0T&14CIWHA#H>Q1.T5%%3+_MN'YE@!AE0(7MCZ4\9!^MMFAV1%XBT#13 YF2AI;
PR.>6H ^[W2E+R0.&G1V[ZH_?C"MA0;)*I9U7U>^A0';DXC*[T^M0=MP\*T+$[9T5
P_&PV]<]''Z79<2M== SS$>!7L!G#SP90SS^^%#TS8117L0W 7@Z\ ;E3'>(+:JK$
PVW\SD55*]X5)%'?DE:A] MY+E #][C_E@5+C"*$DH,1L)I +)I"SKO*(%EH"SS<B
PL!3-,91!PZWS'=U+?%R+^'R6YRVVXU6/::Y!M4<1AT<6IOCU^6#V8\/VZ6O68X *
P"1@=$O7ZD7Y/)/?8>#) B[8)T/=,S1U6JU\/FB+^XCQ=EJZWC(W ;%@;,8W[^BD#
P$(%\2"2[</PFIM:'G:DC!/Z6XN0L8JJ^[$9*1Y"@5($H\>?17/LS%,/)[V9EM=_:
P:#*_/;&AUH\%Q,C X&W O0K=DD4\?R4#LU9K78 "EGF_F(OQ=D6M$$ZJ_);@Y;]:
PESI[*BN?% Z;O\#EPBY+@Q":"B;ZU.K%J392)--;0B2YW/@C42@C)%U2$N\]'#@W
P>]#J]6BN#7?@=+X$VD5"!;(&!X6''P&2[42KG<1U4;ULLSBF7659%;.%]9!3HF>2
P+?X/Q(:.!@Q<57H0MQK0Q"4]6[MZ0#Q<WW%958?8Z"?$SYQP\-G9<UA$2/@TIZ#4
PV6?PJ\("5<\07:P6EFK^(>P39^7TQX7M:P%[P'WL@0^(QJU>].:VA"935D^UU:9A
PX6[@CB':]\XZSIY\[6@$M!G^%\H%>"0KIU4.>_6(;I7P "2Z^$^?)P'V7(* SESG
P:2.0+3A8C<J!/.FVCPSXU'ES,[Y(LL!3VNQR?D561$^'WG^ ']D-K2UC]-OQ[N(Y
PKCA+8RA#.5X4/_R:*F$3;[$@UU4L[,G<H#UM6MZ(UD4O7]0N7ZJ@XFLF?PQ(I_G#
P;;3M1=7)$T%GF=(\\P>UQ*<AF\WG>V&.T@:;>PF(PQ[E\'N\C:2/S1L^XK;GF5UL
P*D(= 9"$Q^: +[\$Z( >&:0A]_)E7.ADLQLW#GVIS]\<^':2;@A/NQI>769YA#L,
PS.W+)BP^N3\=+\,@3@WNZI=S+ T51K9B,X6J3]IQRS-$7AZ,+0#^!?3)+(LIEPU:
P/Q%20+V\%S=M,YV#$8:.U ?9![?I,U(#V>G.C]5O@0-*([W?@@P31D^3N,"O_5-@
P_5W*'VWV\$[YAQJE3VMYVQ0#^K0G^M4K!3OCQ[.RSWHJF%@#Q.,]RQSJKG.[LK#&
P)79H(//U.RI@S$](""E2*\$:\RU">V7Y0/Z9+OAHMS%/U+]1#]B#>)1?2:0L^(FS
PA!J$D]S&:TL:%6*+\HT"V%OB#^_!?A=9&:V-YIF"XT\M#>[(24S"AH6E3,J9N(;.
PIL*-G@EE!ZGQXD KR-;E1T"*=SZ1C_@>U=X+-,I;A!ZE21<EK:FQ\J-D[,BE;ZK$
P25!KB<OAO@7MLI62Y?:C7JMX7]XD^_M%ZL/.2/8Z\TKLGQ.(&5\?-XIFF?8'@7D<
PYNIW^_Q"#O-@C-5_B3C@8L#E"X"+;R_2Q*6D,/&L0*$%1LD\K6*D"%H:5&",$GMW
P[]ULJ]H)8$(*Q2NIR'38740H5EW- M"1JB:3M^!>CUGD 1CL^6+%3;'Q$9@JXKM^
P^2>"*I:DE0 IX87W7,.2#UK/,[_75_(?HTW P!#^9-ER S:UR*/3!F(6V4\K4YR>
P9^6;UG25-41\@!A;A%IR)2&BH#[3^> *CM.'7 &MV)YR/K$=F.#:!=1M)($I'?$E
PP-9<K=&Y'2.P3T9-.=';]\<,3S!(=H0L=V=H!3T@7T!!\O6&Z-8=#(TU6DWCYC]O
P@GAFG;;90XS&09".F6K*<,$L=]!*3(1S75K,IFF/++N#0&&=U#1S9X3@^<GR]@_<
P3*[M1]K5N3P$0S/;4T[RPP< A =#RO6E-1?<N[&H=-$(RKSTXB@X[3JZ19>T'*#7
P4(H8-?)]/(^MD\PDTW^8!)HR-EU)3:]$4QJ\$\[=FWQB(,G,V^XH%!S\"T!>[_T_
P6/X]]L#LI]R&\7+9ZMYR4E!Q!^"V.26NW[^8D\;3H:\LY7 )^R?OL/2KXX=[_$#5
PC O0)*6$#JY+ZCK&T^R_5G)_B8HAH%3Z<*=(?QY;J@WY5__DJG#1F>3]A4_M$+[O
P HRB;8=RQ>B;D@L-,@U3^$KW;K<0$M=4;:Q ;@YR-!Q762S905,M$Q_L<Q:J>*7.
P&=+M*M,@%& U&ZC>P;=BZX/!=N2NZ.TPK\\B^UNIJ.+;_1E@CD34><>\"V.C,N]L
PXK$V.R7&$VAM9F&S![(2Z4D;*J_IW\Q1Y$'U<4U^0N1L: NG8/^!2<[ZN\3QGPJ0
P^,+ZZ$^;@P/E5XA"T_HV%]EEB,0[ 5'K"#P*+WTP6L#5<TO$<U>>*H4TG$\]GA35
PBD?'D[A=A(^K9:\2F%T)4XCZ?KL%$PZN!/.HQHCC3,+*]#^LIY.:L0Z+VK*OJ"-O
PE.RF7FIMV.F2-=6-SOIN/-CCJSZ%LFDJ[G5]\J1ZI/7=4W>&NS$T%K=2%0DL@Q3T
PZZB+2S=,-:.*<O^>_X6=%UKD=Z)2]#8M_=%*%_(XM3A[%;(1M,#(':.AKF'O#WWQ
PX+]+TPUO/AEN,GB\I%/?/BWU!#Z3_7T=\Q'"&)2.']O8B?UIMZP>;G[1>&P19[;:
PKO?&+I0EM80.>D1-''-#^UM[82IGZ"P2GXVH>D5$N"GCQH?+Q+CNEG->!MN,Y8P9
P8HW, ._5SJXU1M6Q3I^*"H?J5<>?[CI;G]!6G\>E[7<.#I^Y+6.;5'FH#V">>)(2
PJ?YSC[;?%FXQC/+]]%9WEK8/8Y:1F)<*3V,%31GJDQK'GVW=?,5QJB9[04.LUV6,
PYLO!N((N !-=M&.E3&H]&TR# @+"/1"G%9F$Z^3T]K=AEXXZDV0XP2:-'^6RU&?.
P!A6"&EH8:?]QP/P#<SU]Y1 2Y+*1S#0?5\)))]KGO$YT=8EEV*.*<HC_U_A%J'8[
P".8I(.,1@K 0FQT>!G\C3\QCR8DU:_B6XO^MZ!J?,19<$@:SG.I DH]HCBP!V1W@
P,:MH2;0S8]< ;.(/P'FR_18C\*J<]@5U@Z 22R#V);5E+Y*T#94188)-UPGWZI_W
P1<G/,VUN#71-;9<XT[$U?#E"4B]";CS<$WO_Z%_4?F6&":6"()A+)E(_J^A^F<\&
PR>\V"N^=HQ^YMVU9859H]NZ0EOW)F='8,U1 F\R6O7;@TGV8E:O'KY+XJX8G!*'4
PXT_-O(]Y_V<YJ;&.,7!08$Y:BB_!1O)XV@=MM?Z63G[>'_5Z:1"2Y[")+?GT05&C
PS3[B"5T]EHTMUX@)*M[(:D<'YJ_;-S(UR3TLX*^(Q:$:H:=Q"@K-Y1Q Q8J?EG&0
PL,@P8J1C#",;3LY/$W32Y6Q(_V$RK-3+.ZXJ#Q<;I,9H3H?TYJ&;CO UT+W(>HCY
P]33%S[A=M0$C/-6UBPB.5O;"^/(9(>\V?O%-R.FEKN"&3&>!"-Q[SW22T'LQ>#X[
P&LYQRMJ#'^M:(,3$1K7Q?06(MC?GB804/"&DY@;S#9KC\S2GP83SP82Y"V@@PS0W
PK.D##,U:[O3X ,$V]SVI8?XX;8V,3-OJY=!+HX-*J@L(+LK>5G5]LW2*/?Z3B WD
P0>V"D;K@H\BDZ5':)@L+J'[G(KO[*>E%3=X3+XZ"]?GV8*YO*%Q4>N&#RO_C\U[I
PZ_' DJ]WE(+R6:<@/#\X>(&C@SWJLM35MD<%P-1S9\>T-;@^K%GVNV&?CB5O6<G?
PUE-^X *KX9)=I[M*I!SY!;41(#?S51O==XJY5H3?VE^$R]%<P="-P0Y@[TX>NXT-
P1>V,#'=HN0MJO+C];IJN@#CRQIF?=OQ7=^EL=93D65'?!U0P'?1[F^V&:NEP.)(]
P$'&M'-=>=D-N[7I!ODT_Z*U+<I&/?.0N8:I)#TA-[/1WZ^Y7Q!8&0X*(-+V@09:K
P<#A @]I_0I$- %PT]XX $S.5H++[$Q:=M,88:'5)&#GZQ.(VFW"D0D:TP:DK)+^A
PL2XU)#A18C?<-B )A)T4K9QOGH/F+8SU4*>FT_(3I3M0TE!TWJ:)<QJ="B+M&/&)
PYT@QOFE.'(;$V#[;Y=M/P28MKV;V&EL>E @<?LVW%LD5Y2VXTS+9JZ.V@\(0!FXI
P)5-03;?AAEO2L\?-OD&67P.VQQ<R.RZ,V%$H?01D^JCZDN^&WJG-$8$"_]RE8/&F
PO'7D:GW&]C4EUI0[<ABW^/'ZOK!D3,%+DM)"#]%79R6L_K=CH@J714ZQ/NR3RM>/
P@%Y&R5QS*1M_,>[DR80T]5TW&\TC0)(V:U_(4 !MV!CG5/=F6\8.;A D$NK1PM(*
P[)*,.0Q@)RQYANTT7^?:^3 ;ALYK\1>D?]<.JG!+-R]-3J*^;:AS"VTN?.M.3_B.
PYO&2CT0CFX></@:H%SI@OG6<9J/$4W6HLP4DO8EFYDN[VUJKX7*F*BJC27NB\MN\
P=4V>-\V5\BV'IS5F$/KO90^4:?-H92+J-D;(P(F76><LN?Q!\]<4#FWSQ&?C'-A 
P/UTM>Y5N<D^4.R=AA7.689]]+7-+I]_\OQ,NW-_5>\./\\YLOE)=K1[>!S($OOB+
PAV!]HXX1<Z$NYD8P>>@HK2"W/FKLCHJ"*_&5KOI43.JIR++DZA7+>R3]DDLTWH<=
P?5E2#A R.',NI*IN<"(Z./X<I'<-B,0/'LJ@LU=24P=(QXW8*@66VJ/)KY@F#(@E
P'83@HC ?6:*KR[\HD$_L?X HUQ[\C*2\Q9Q8*F%=6$:&8[;ONNK!]29*+,;)S6%:
PSWP[_  Z$9-./CLZI69%K1@CC*[">EE,>_%W:"+D::EK[E,=]L.\(PU JCSG_^=V
P"8[1*-4-L [P(" ZA*@/,4#:_"C<5F)&H'$B3RMN]5=]L\.O[/,;L,+O\0#?J?XO
P6%]9-R]UEU9K:1 "(&E([\E:"=YBP?& 8V$/GLT<A F@F>F>>R4</_8&&8_YU>14
P84DV?S6G#R"DXLTNN@YWM:=^;2..7,_F?T.%<198!Y=59]J<A+G"Z5>:&#D@7Y6N
PLW*N? "J45EL,H?ELV)0U$IT\J71%2&JA[1&!RF0Z"S/BEW=54W@DXLZVY<PF)D*
P\)I<_[=L@T<D4TA%]=E1'Y+=H%EYY/=3@QO8/A]M7B#/L]\ X0J!]<):K%-C\7GB
P4,[)0;$WZ-GU"5-6]4OR%7U,[(9PNZ@5)]=ED' ,HTETF4<C]LR$G)I^N (PPXMR
P(+?,E^RCZB4WUU%2UQ$%[,#33T21CR$,Y#YU83. P<+/M'%%Z0:^\7G1YR0BQPZV
P*]V<SF?!MBPN=X<UZ<ZP&?(124T_WU[!25/MP/E7 :<Y.)/%F1?Q97DE_EG0EFVH
PI^FGI2?"U^JSS=YO&RDM!#0"]M<0292>7FPN2C8H!1>-$;CI?(=+3A";<0Y(7E!#
P:]=Z/V@K5T$-GXK]./G'HMK9ZK_+*J(][$^=S#Q4V@,[XQ5,H9VE 'L #GI,'Z-L
P9JB>]A;6]3#6Y6+_[>=IHVGZ>0N*U!>#?(70 KM8/.E\I).L@0<PLW[P:!T*A\=\
P:E0=3 PO@]$TMT*F.9BI4:Y#K4H3$$9D:K<N89O-/M0ET7V,Z/N3M7*3B/U*5D31
P<'9IYM5<HZ7[8[%(6?!:I!ROD-K>>OU'S$,BOFK5&LD@6P@VN0"2L;-]EM3(4L[?
PJ9Y#!0O >!'G[T[73)LYC_@2X!#V^.J<<&"W/76W*TIUPF4:Y2%#H;)126O[B3K?
P%2+A;$B@<=NF@C%/;RNF6\#*(XQSB %'D%AMY_[R/FPKDHD#&($/)#=VH DX[_9$
PI>2>UOO T+;5?N%_26?D802O,F6OMKCNLJ2U7.;L ?+)F.7E:RV$KG/)"O..7(!!
PNV#Z]QVGU46>ZB0>5NI[$[F)D\6"WGY#W(A0YCN1$?M=B^WP;>8'L;FCYO>MX1+-
PHMX+ -^D*>+J!WFVVXH)N85\TZK/YM+/_&*<AY/Z-6TDP12-?W4!X:19 Q[C(C;J
PPDVJ7 9W/Z3=DU -7)SH,E)Q- RPX00E5I_RM]UF.&&UT(&JR5G%%$0GK1'K,]A5
P'"$L\&[ZB5[R0&E*M&6^?Q3=("E)U0X=+/VM2%:'$G2H^G-^B.BJGACY6!V6^\0R
P!M!F/3K#I%8O-G]U)1.D*.B<PN&2H8\'&>07\62V*^U4IAO%91_>$VU?5JW+@/9"
PVX4$>^,R0<^J./KHQJ !9L@.O?_1:99*H<EI?/W^$VH8/:84>YJK]HL)PA1]^W>>
P(_SF '!IZ-8?.GW2#<N;R@4-T+A5+HPT-G@^RZD7K;(F(UZ]BTJ$8OE-Z>N#*,9L
P#/2JW3>P77$!;9!97&^7?=;V;4]:U#8FHL:488PUJ*B.H,X7X*!.AZUJTY^12CA2
PS(/CCTG)T;7!_DOM*:LK)%J<^(]Q2A^IAG$O>\Z(\*YJTE?O:N@I56.:4.OBSD_ 
P&I7U-"]LX_+TXA>K)_YJZFY^+UCSJP87<$;5G4(P=AOO=MOXM]D#\>Z4E:U_:<U4
PJT<QZLE!R#QUE/851_C@9>C,AY*LI5HBQ6/@EE*AH1[F1/\T4)[/0R0_PWEY&G53
P20(DW;>R?^\4(JU:)9J_3V#K;*B#^J?:J:!F=(:*V#?Z?9N<Q@+XQO?'$8IRG7I$
P3G'*PG]#$3\4M63$P(,/)58E,C8B4T'::V27/TAT";88-G*EB>N.H^R^R 4Q+WJ1
PAR)I'("<"3<"Z+(J!C+__AF$*B01XUOZ,N!QE1_)G!I_?$RLC?4V3:*WDW8\S=X?
PA!TKU^D'BV,U>\Y(H$<&ZAL57@SFC" N:Z/&]OVF P?OW$?^RSI(=4$;_Y)]I9A'
P^.XC*,%_OY>F,RM^\F)?E"KX;0O+QXWHO('EVI[BI-$]:\D_]S!R>0%F*+8D"K?(
P\5M:ZFTGC:H/2Y3^20Q]"<*7^TFE?Y?\F4>Y9X4/('$N[<"JE6*+]X3S<0O/=,2T
P1/4J ST)A$M&1@VM8C8-<D7W3!OZA' ?YY% R"DX58%-0#ZXGT9DGZ>WVWJC+<C^
P8Q6%J/[(<?E"E5&X$Y#QQ#BGU=2 CS-/1)Q&AR7&WX?S[H-\8<H$_2F5]ORC8DL<
P[.B-J_W8"Z-$S"% OO3CG#OY.'5#]A$#&'*F/3#;NU\JU0V]MP6VZ B>_$N9,O^9
POIV:SB_>84$ZX,*09A2')()Y>\3E]M=GF,!P"UK2!P6]P6S8_96&__8I=Y'D+H5&
P&T_S&@"\_[VS&$*+,DU#'_O.LJ[5.>Z6-LOY\-!^42^>$XF.M@CM,E6S>J.%9&'6
PC1@9IS[BGEIN6[E):X$N$ FPX2>@T^IMRY\G@XT@*_1!8:1$$OL^6J)'S9^FA^-B
P[%VPGOE86L*<$JT:>ZF?7P25QE&<9&KBB>)/FJ+M$D @&<@+8!3W9'%07*3@IEDW
P54ZIQK/=5!N'2=,8Z<MF%SO62LN761T\5J/CK>:$31FVQ2?Y+IN=MDH\-!^=[/+D
P=?-:V)'6$&SM,5#J$7^*^")6 =R;+ED&NA@&<"R-=$26!N4.YC!G'5X.<8,.K ,&
P,A;S-7[)^>6 32"T&VYA71<""X]*8AAG26M:HR9"0R6F,D"9L@6B+?HOW)<Q%=JL
PO4.!#*_D*5-W.C9)0!S".;/"J#_AWE<'57):'"947-!2>JQ BJX]0XU=0L\(1XD2
PHXU]2?^JMO@;-QW)%>C?@)BW8+7"/*"XN/?=QBW E>[CK[)4[?/*C8$ZEMH[*L_A
P2UM6L[^I:2+C)VBU5I+*T$Q(M/6\+ ;PS<P<+PA<0\%C%YC8Z4!Y2&GP90^05$<(
PB83A@5T+F"GS6%5.&K+T2!X@Q-B=XA>*QUNO)7XX%% X[DF%$;:88U?+G[<1(\^9
P:TIZ56>@%BSCQ2J<KI3C^DZGOP'XP_=#->'/#1%P/ZNS BR@1+B_L3*E8IY9CGHG
P!UC5A0&^,9W[3*3X4-/UMOMN-B QSL&TS-BN=9H-MVWB.*O08_ 9_1#2DY%IF8]@
P%K'1L>UD)E PBL0QBS^3!3RKDPM32\3PBB 3\V"X%]UC]+=(&)CN;_[8AI>2T"E/
PK!JJ-GL?!,N#*%L)T0FQO6% CL\PSP6B0Q&JI&G0V_'[_$<L3*?Y$?OSOCA?:2H5
PK;-W?H!K^GF0UQ)G9:)*Q="YJ(,2))!2UK* !A(E5L>9_28$@@ $Z3AHL@/E=1V?
PN%&W".JFD*W*KR\M4L)O<XR7*(-^?LYM2J&M%E$*$5'=<RW.LB&$%KZ6M=ORF;!,
P/9Z;:"$^PU<.XF_,H?Z;X309[DN])=K6YG[9X9MICNB,G+GT@))J7J'8%AX+R:5J
P&6/2RF?<D;ZHD>U&Q]BSCFA/>-5/=?^/5B957>@H]R,]B&L6@P 5$&_>'MMK^7,M
P?'\X072\(RC!<"B!:+_?WHD5)@V(6) MOIZH*0?,5_OYF$/I%)QQNR.6:37 HA9@
P48G2/9\QPGR5;ZXXPMJ8QX2:3?%O,/Y"UCCB73B?76JK.>G5=(W*ZQ;VNBOEY#T^
PZQ@NWYU_%5T[&OP](=&3I'8PR_&J__-IZ]/$1&5KA,_;.L$'"G&XE)(9[@DR@ .[
P.V15'%R\.4&Q>_I,\\MD51>])*@K$6>RNMT G>U%,3=V <&I@\:$PC12F<OAEJ<9
P+W>R":[.YKB@@VR;/65\< ;4K%CE+F^@JV.[_Y%Y?</9>O2G_8*.L6XN%Q"4TS:3
PH*K4:A?,?]8-/EVPHUCCS1A/-/E]%4(*QFFZ&G ?]9"HZ] 9OYYPA446?=JJ_$]8
P@0XIF,2>,^-@=#Y&61!NZVR,%(0A,SKB[;^N=V+&A6[2MOVH\ZYU/% _M+89^$R2
P9XY$ZX>AR5)$4(EJUP;HX:K;6GI7F A;^0I8C[$U_SIX:;=W#%"IE>D]EGF,&C!,
PWEN77+"Z-4\!'2K4,!'ON Q&P@9@_J_1VY_L-.!$HC@(R XX3ODO3@M15PWY YD(
P$!]EI;HC[B&H*M!O'[Y9- T^%?.\4%?%BF:C^&?#A_/WXH)5G0M<?C5+DL><5[AP
P?J4'2)CZZEZAY3I#!+IXX+863*7)NZ;0.,$F:>XSIOY[Y!5F*0.SHF06'C1Z $CQ
PU OF7];R+;B[D;Q),\C%@@HHXVI32%DT(D4G2KIU-D#:?+/P&1Q$O/Y)CZFU<+Z9
P,/B?OFKFBJ% -=T.(24Z1Z,XJ512_P4D[/9F%3.A-JF#M.LN$O;5-$XE>\/F!H@^
P.&#27E?:F-+@=X/:E[&CTZ>WY-#_=;KU41#P(3E%5"(@>(]07J%_5WA'YQ.')]H.
PFB\=L&98VA&L''N*<DAU;&5;W_2OY46#G\$K0!6EKM_#E81\6;XCIXN 2<D\# N+
P58.=+&0P#Z-F=[$"]@R%K8W9A<#QDPR)-J=#LW5'G;9^U>QJ>M0W[36ILH=BK5E7
P*9?1;P5:A(EFD1:\Q@'@4TK,+PD*Y,7HN>V])JA1(!F6MZ:@F<B2FMZ(WYHFDL:X
PVV_NT?]'7SNW+-2&D:F'WKR#A+N=*B<'!R!M6RKBS2%Q^(TS^EZ#8L0.)!V0X$F>
P,WQE&(%^#+_B3>GW-8K-VK?I-_9CV\->A("UE%N/\=U/".;-D.#?+;TU *^28)!#
P4@6[,(B6$/-^(L*Q;YY]G,!';==+ -C[GM4 M-BE.IT56'],0.$+,^BR'TZ?7M&7
PQ217ODW._N"UUZ@=$S*SR(YBXA/SVFF9I EO/4S9LC: AS9KYIS.;<<E+)+]5(7F
P;?@"/[I52>ODZK...-1W9+,9 6:%4%WQ/@MF<F?I/SP+9Q?/1;:0*;L4#)YISE7W
PWRY-&":H<P33;"E(FF[<$.1N%'H>+%Y+.Z'B7!Y!L, T- HOX+ (.%4\ZFWI9:9%
PZ\\%-.2,A!_J@X0> =];Z\AI:C(ZXG*-+1P6D#I^E RUFGQ^I<DM9BE_^DMW37OD
P_>%,%X[1A>("JHRN]/O\J$?$BG:WA(]K=1@N$QH\I>M(]H57'?_F6#T)YX_S!5:B
P*/!=-U^N'D;UH@NI[472)' K+[.+*D_G S52<&15RA%M"8R/)4S\2<)[Z%M4E;CA
P(ADICE+Q[O! 10@0G9=P-E:R/PSB*Y7WW26=CSUV4P!POUMCPH>9.IHKB54KO*K'
P(UO6D<\@2C4;#U"I',R_'0;""5"4A!,VQ^J##%YRY^[U=CAW%&5J!:3:O9.AXA0.
P?\+/8B=,^2$@7'470)J5ONVGM@F>:CLS8'N-GS^)^<(Z7&\/3QNW?/0E2C*K= ^4
PU] RVI*[9Z?,]POY2%<H[3Q-TO1-M[ T20!!;FJGD(A>+5"N1W S<8+ND!C?81KZ
P$'HC.#C)Z1K">]3&KL,0'V]"!27>12!&9M8:3GS3 ;_?W:3EREA4U 526H@.=07@
P54V+EY'(6\?EL+@!Q.I%&]7"G(_CPRU*.-^;WQ@YRK9>PHTJE':Y77^KJELS02"7
PA]Z\K//0U$<@VH(+/*$?J!:"+D\+5SQK.B>Z"QG\!,V:3)%IH$S0RPU_U9;<9!W&
P/9IH3J5=T>EDSI090^3>.TD$6?2>^LM<]+&?=';)-*&77KU<4I$[%."M2IMM_O\B
P%2P9;NFQGB)N[DQ$.\Z*+1J=-$K6SGDWQ-Z,(E<JO#.3X_9A++&TR?<>#?&[O*^]
P"<#6%+[&.ZJ-=3*G=GEXCBIH,O6R"$ *M:)KV4^&X!L$M8,SNV2E%ES-R<R%)M8?
PUB2'C%;*QZJ]W,*!R@)T"!>E,2!EUWK(L4D? Z"^3FPV502GH>A1):/('%PLG(#/
PI!4!U.W'A-SMW[^1X<+LRVS;%K#P9M8"U335.9:9SFPFCK1/#'8O?1Z+$7L;&3PQ
PQPTBRVV]Y+X5VNPY@Y7_1'BCO;SIG0P[73P9/ZY$GPE$/K;'7^A:C,8SA/(/AJ4A
P!3)O>E!EI<($!_IL^02$L%08(/OXL+&=@+VGKGWFR/KJ HV;1<K!)Q,L_J#*G&B1
P1'J&L<#)Z9LE.S>QI>C4%MGLL)(3&ZT_#SWFI#U[R-5$Z_Q/*FHAH"SG'+JW5B92
P!XNVM $746M&;]=PAK,0_O>-5J#K11$&U):NNH5GZNT YW]]>H6!1R9A2(P$S,:L
PZ+G$(?OA>6 ]1C@QEZGN%_Y$")MJX;S>R-;6.C#)JV\OHG65M5= %2&-K-=/,MQ(
PXP[_0==U:2^'4$Y8EFY)6SLE 1T!F46/1:N1G%W0,"PPR>'/62%-T1 F8;YX4M2'
P&34\)MI9_PDDF"4 +R"DH\BNM&_V 6[)ED_#+DDE& [N$/9VG*VS_@KP1*@_V2P3
P(DW;[S?+-]I<?:U7[:\W-T$==\YP$?W :E*EVO@F;Y4; M4TE+C5SXI,<F\$<#3.
PKAP2#S-6*#.-H->=TX$K7<CEC.FO$$)#3=QM404-T3[P.KSQ'IX]5HCB >86*&4>
P=W6,$SH7/QQ</WN_QO=U)X^P?WGH<NM-A_ C^Y]44Z?C"N76J'N2]V1S#]Q%^PY>
PE_]44VK-S;W,OFQQKT6#K<Q#(87VV% )>13S1J\?L:9Y<^&@_]G+G]^52%",Z2MF
P<<MO#<# ,(1+!7E27_8/BIP3Z:Y Z"T;1G?%[W\:>R0TJP>?LIVHC*)J&B%FD3*_
PF/0Z?AS$U=C2.(5DX]?G25N 8=V(#K)@-A=&F>S#-$<F E7C'S_[&E7!*,)%@4!_
P7!?"RRG'7IIUD4[=!ZQI&!C20B'L<"ZP8MR0MH0(J\J)4*;R1JT'%'?ZY!<(E]1\
PZ/7K@CIN:";+=++VW]E)>P0.<]50)K4V)$"'@2<9<-ZY;2[#RX]5I2(U4Z.KECY;
PQH1XMCF@2PY8AXQ6>363KS#;+CW-]U^++RDTT%7FHL&/V<0&9W!V3=%I:I:BA<LU
P2RL1>2TL@CA.Y%Q$@R,."*@L.M'JGO#*OP>C212NE]GC=B]Z;7U'IO/<M**YK:_@
P7F#7.FD>]]0KI\$AK!Z]/*A!J:'EAYM/*MA*41'""&=;'J D04TM4PF_)%S8#_WU
P@9"6B) ;I7\=@?[[2<QB9/L_I,FU&0OG)#J7 APE<RD\R6!W,0DCR3NYOF 4?[V1
P$CP.4A#_@> T9"Q9%F<+3;/(5?GAH6H,PH..@R>.^\;2L2"31#\!38(#]%/\IH98
PA&XS0..P8E8?VQS%,S"0<MQX^8V:ILN6'' Z+'VIA/G&:,1UDBNP$-@YJ2LYI'5]
P36;VH%PIBV =E.3GG69]L=.1Z!OT1I,8R4"92"*^WNFMS"Q?QU9D82)"_K>A)SK 
P6U"XN]319N?D&<-\5';VA'P&T=<9=I1\TE H(ZZ:B]R$E"A"DY.*GUQNRR4Q<&9J
P%8RTIL"2(\SP3!]I3;0@)$27! .,%E,:?G4:&[W45\ARD1:J<][ZY>O\(O7%&EIO
PG;\??\/5N"&VJ(Z9\( .VRNH1;B:B*DML)9#L[UI7J3[9*Q]TBM+]*74<A]^(%>-
PMHY^!9%5KUQ\8-I=O]2,&/.+?ZKQC QK5Y&",:B^7^#K9M=QX-?BWJX<%<^-4JZ5
P\?;8447=3O=8GAB/WI#4&PC3LC,I#OFCX<#:SO%VD*8]"'K&L$'O=U5UMOT!U&/X
P0_BB<&(&$#Z X3%6I.?(,EDV^MB:/.^*^]5 .6$RHYDM'1SN<I*R:&6\]V5RMK_.
PN3N_Q:-@$&PBQB^-DX"G^#OZL4;X:&Q,EZ!_ ]XCJS'.P<"KFZ$H3<'N2@_3C"!F
PLQ/>?\@ZO0PE!FIPT^0&05:60#E  DMA1U6M=;?8&4=OYDP&!'KVJ/!,!S^3]H5]
PG2?@!)-A6?9>8@_GHS"FDDN\2T8XG^FD&N<KM])Q(*%W_3_&A!?-*LZW^,<DIE[ 
PW\F52P:&[DI-[=TMJNV!OL#7>7GFO.Q?)76N(8![!&$:7AE#B+OE:(M>A*2WP/^D
P/EC@ZGQCK$L['F/5RG0U0!Z%Y")'AV#.'5P"\RF@A$D!RD-1(QG-R1/QUY_%H F)
P,45DB:YUKLF'PIE\Y#R0O3T"0V M+#E0\4JEBD36O3E"*4TR8^UL/^2,R=&N*2#-
PE/<J69/8H(RJ&,%A*?!"N*S+)*_B. J<EJ%%8BYE1R>K^/1C,\J5 ^= '*W42Y/;
P'*1T-C9)T76"XO5\;7RN6.9MR<N7+L7E <3%3(N[QG"Y<<J)4<>!#0Z+C^L54HTA
P.MZ$Y>J,NQ[(&\7C(JYH9%.>@<?'O2<5G:7=,GOU=:1P(C6I&M8C"L(9!%ZNQUNM
PU0ROWB5\TL[&G3X:F;I/V&T,9/UDC>8'XGE1>)G,.U#/4__MD_K-?6J@:YG]V>[9
PZ!=OZ&P\S)OZ:KTC\?YP)Z492U4, DXC6@Y0]5(T:BZ)X\R,B=?F>*11* UYNZ&[
PX=X-;:E98Q0DQ4/JJEGV;W:;A(+(I?)*^SB_,C^JSN5 ,W/&#LE";5I[J#4723,P
P"&BM G@#6BMNLT_>+Y:N]VA.",LY- ;[ ^MY:P;4'KN),> 8RR(]#KRX6V76\K;J
P=@I) D;S^;FD(;@2OM_"-#\C/G8J%\G8;* (K6,B[.#?J 4Z0\ ,(UK5Q$)9%>ET
P!NFSF-#@G=BIB9/),-&+#OLTMI>D%/E)E@&M#(CH8PB=\T([^=[3FA$: =R#59 A
PI'CRB\$W$.+/^",?L';D4KM:3?)'S"Y2-8Y ;$I/%=<T9BGF=[/E&IW-OKGW/'Z;
P!%/5P\9]X7*M*$\^U!FU 72NI6M6E$PA*!X;6[=?HFD_?QLK-^7T>/GQ;GOYU=Z?
P].K"OA^P@]<\_5SI#C#8E=1W5G7 ,:_]!9WA=XD!+WHCW81 'P,?KH[]5']Q,.O 
P8'[&'3&XBZ>%Y5ZMY0YK9)<<) +=GD0%P3]#/P=C1+*'M9 MKN?*C'AZR[OODHM%
P!/U_(*F G$1'=]#;8QY83=0*UJ4&1 9..@NJ#&<]A*"&."^#7(3021^BHPH^CO2W
PI#GVE6I*(/66J9L>(5@:!AR306$!O1L*)OI"[^#3G4>"Q6Y8_C?@^!54#(B9%CRP
P,1B9D[17MIFTR^(V 3#_-ZJDH? EG_!VXI.%Y;/_<V8"C6?N+?AR/%$I'^T>U@>D
P(9"8C\&DGA*5^T4_:G9*31-^@L'9;2E(=<%Z@A-/=EN0]1V.BL@;]?:W!MF0S>B8
PHA0?"4S2=@(5D(Q->O"YEI@(N5(UC ZR<LP(.:$)09G;TH_1EQH_ENJ2P0AK$DNI
PLAAUA]58'YRV$BAM!9*JR@;F?+*OE0/VF=ON!3&52&"WW@OUC'U>$_-/>020<6HU
P%Y=.HQB3K'=+!^<PF*V;]>9]7!G"9!<)=6AC#K^I)Q_Y66Y_DP_QX+F@U6X-)Q[4
P7*6C3Q=8-=KIV)5V]7W)4I^W'J&>XHNLF_P 4Q09;=*LP+<\8>"D(D5W5#9\O4?G
P-]-A-S^ES>[YC(,#?/3/S^]TL#R3VWS32JT*DYCK2>S#] 00.O@HTJ]:$XJ3Z> R
P8BX$A[]/=-D,7!T8P<#& 8PK&P 3]%E!E.YZVWRT.38(M#FA-J,KW.%VEN56A'?6
P'=?2!UR.W#=F:L0KZ&DDSM.D]H3_!XGLSF"0&WEJ(WCG5IL\QAF1O..$^)@8#UV2
P23]N$$]#'H=AAS"596<,D9Z8!N[VWZ67^AA#HS5]>ONF!*U(T- 1G/%DH),0L*0@
P6NWF#NX5+K43B]AREXKE?+<^HK% #"(.IQ>IQWH"Q8SZ31,E+J)(YL:,O?-!4AXF
PD702<Z:&3G276YZ$S+L6=_O%0XKI)5,[!FK>FK\L,+V,[WD=.7SF);U2PQD4?US%
PT%/#3PZ)GICH5NI'60M=T-SDG!"%'B7[4!1U+6G?PM83V,GM5'=0_PR7,4()&@>U
PW=J0UP/_WD(<,=+?>W?A'=>%[7]TM?O:1"02> ;>MJQ<C"^5FN&"KYDHLWR*NV)=
P57-G3E%=_Z!1@+C0MA;4,K*7FGL"QA25W\'.I\ZT6)OUN+@A(KEA8Y1;'_]CA&'M
PG([8*L!- &D&I(F\6<GGM1_83HOQF7DLK9S9.TT^ET[T3<H'4-3<8(.O#>A=TX]7
P8U[)<S?['7L>LB6@4-DE<(IVYD\PMQ<=B\4[M4$8B==3SLQ7Q4]0D6P]Q47'))\(
P .O0 :\6C]^(\26@Y'8LF?XP/XFF>M*.H-POH?,U/Y2I+_Q\75IV%2R5;;I[2;5L
P;5HD1$B?OK!=.6C&-Q(C\\3+Q":1-3O.P4H7WHZ#J9@RB&O)2--!1C-VZ-!S:T$>
PX6665JMW.OGIMCFK'>P()&)FGO T]9;AKS"FB'<2)B3+#JS>1.N 0T.DPG&OP*I4
PHR6MLI*"1(@&ZS$8G#-'&DIYH5Z@Z4?XBH5TN/B)A0&R$77@8(//PW^YY?45?28'
PS\UUH5Z ;DSAU <*%U*UZ!#\SF I%6GC$KBP1MYGTQ:GW(?"I]GF]ZJ=PGV!JR!9
PT0.=!K4G]B_B2$#O+O]E@C_[Y'.PU C'#W6!^!NR=FZUD*G$.)G_F??P*/LKQMS]
PU8!X"S,M@P!90=7Y_ AR%-7<.%SBW-,3-WEQ9QTU3O,Z_JS3_85)M.#)D_O7@4JH
PL-^QFVLXR:+\GBB/KITC<;'&HCF1?G#AE?OV]I2].17YQK?1H8?)VX$=*&LKF78!
P@)8]58 Q5^ [:M<2(! #SIJ++.-]<F6Y^<D+F'KELV1L4<G5R"-R@GM4'63[_L#4
PS1>79M>V3P:^#6S:AB;CV5. J4@6H6*MK4I.<E<##:M@ ,//L[=NT]^)TCA&@9X+
P@)AX4O?DIX1/*6$I5LTX)>3_[[@R)DFVA.H%^]%_Y @A:^DJR+_G'N-X7WN##[==
P96N\<YXY!JS1-X\D[L L:],E*&P"6$.E%OUM!'#PQQSL-YZQ=U&7X7N",L:U]8#6
P8&I9MH6:6@-6RM<CD0//.Q)T.W%P+AZ?H:-X9N)28U^'50A[U![[](4)N*SJ4MST
PU@.UEIV]P1S?<L65]:>OL]W8)0@Y"!O@&(_\X=<?6%NOQ,LM8<A9@YMP=2FVT8R1
PF D)OALQL+0%3*-D'^C].?+NFO:OW_EJ"0S^5UWTQUT*A0O;O:EZ3-0)/<Z'P;!$
P5\S=^-)LE"QDD+\LVEQG/%?1TM\A=F&DS92?1TJV9>@X:?9*D#E, B1/(FB5(GS]
P_%=>_JS]?-(#C?$)$YQ9P?1;"+D,+?9WT5^6O@4 ]#QPD/( 7WO#3>>X2;QM;B!M
PY%>7,;W9%!MRA]Q](.?Y)6!^/\*E!F@WQ8R?-APKYSV1L]QK";)+MCW;3@ZW!E!.
P)=NLW"K.[Z;3I;1Q96PDX40DPE-UA60[&JZ]C4>#B-%:J2\75,E;])\9FVHNK66I
P[(_B?56PMO%D+]DY4ZX.AG>+52?9#L9_T<FU2^%KF)!-)#4E.6H,\-GMDE(=,QN0
PJL=OVKN*!QV%6AYO1;4K45Z:8X-XDKKQJBBA^TNS!4OO-]7)<)M"SB+L.WZ,HL2A
P^AW'EAG%!UY%2UT&J^H26+S%3GN1:^=N(QG+S?<_H+XCC7J71U[-BFT+_H%FM%="
PIE1\LC$7#?U:!Z"F<4@MA4"W"WC5U%G4Q*'Z-C8Z,!'X,FDBT[7KP7UNW@LIT>'S
P.4!\>^T7!5,SY3$P%$E#>=N Q?KC>K0BAB"M0F/LS+).5,L]RQJ8<$=\*A[(E1>K
P!(S5[[K#G"AM!M3S.SVX@:9@\W3T,?.=WJ(L 2A!YPR-]@I%\U;FQJ -'6M+%=CT
PL47:A%'?G%]$%!97*I8O6">4?27*K*7CJ-$^G"6RD$_GET,,M8U6>&&6?^BYD4;I
P@!T,],@F%61G80! M+=RBG\N*%K5O^YD&) ,4F@(O\R7[EF6$5CN34/81QB;Z;^8
P'RQ8&R[/8J="F,3I)ZNC!0DCZ"7?9/5T+[D,S8<C3K-MEF,R3-^9R*M]7@B)Z#!$
PD[3W0*-L9__N@B@:E6;Z.C5T<MA1VB\<40FD4Y!-O6SVX4@"@,+ V"B,$>O_XF^K
PB16&J%J+\9G\P+"VN8G^>/R!EPE"J?#B60%![&\%$)2DLL&"5/IIA:$]!<8%H\D1
P5(C9$@SYLB5%)L<W;IB9E>YWFY>V8\J3FEF/\*W,SOO>TU( AZ)P%6UR158_M5JM
PL,E@(YMC$@%>!7QF_!#:9A;^2Z, +=Q\I;83)+3([-9-$[V?>=07R;V+#*&NZO[@
PK-=$<I'/M)BLWDF/CZ&OV2^*FK_5!E;W/Q=9:V3K?5I>/V3;FF B)/$\X1>]+,$K
PQ#U<>>_.E!!'K7B'U.U0"+Z&AAL;\-)#) @MV(275\%M,?HCB&1.(@5U:ZVK42["
PP]'\RJ[5[.,J_<K]:FXJW1KB>PGHF6 KPW[JF2K9U2-W+O7Q!$.FDU;V0VUVBM0W
P..*B/LRV&\5FCQG7X5]]'%!T+;,_6P@"9I;"<HCD'<[$!G,W(D%BM)PV70PXZZUG
PYXA"@.LS0 VTDP2EYK)=W'K1D)UTBC@82LB235Z@.>@:&;&M/] *L)9A(,+X,X@O
P@6%I11*V^(P+U$BB65Z:IW\P6B7I5078(#L+;Z!\,3+BB-$R/>U:BU=)ES]YE/Z/
P(?9%?C>+]\+X:06=RGVRE4D/*;"<M:3A+?!V$KE;F[5.<<:O<IP-6?T_V.X:V2I0
PC1'9@B;=#_;=.H$\3_F2=RE_AYO!HLBT Z"A P 0%<OL6<34*YO\_<J*OT.71_K.
P<ANIIP24!:+C\@5IJ,+:1XFOE!4[=.R2@XMIALO>BK=&K(G28(?H5V^,7@@#0D^7
P>$ :6>^*M(I>&//CA*)DQC3+]#:$%O'?MQJZ\W^.1B0(XI"A/]+AV+DG20&+V_FF
P4Z9B '>?61S=$"*[PH(BZAQ%@+O2&9$][I*F^0,,Z+^P1103!URS:T"DE[J+!\-D
P'X(]'IPH=]ZPQB(Q76((,=0M2X!?4%"P-QB&-.>[5N5=%&L9QEK--N1B4V&TF&B3
P<6I!->U4A*QI!<5Q#"R@@C1L]#R*QU$6[V5RF,CDOKPS@04<"8M4,)XU6DD%=^^>
P@\LA(TP[LDRG=&Z"7Z=J&#:(IW;D4/G3)QL3!=SSY]TZU?UV;-K[%KA#GUU>I>!R
PF^(7$IK.O<UI$L6KB*ML_#>@$"A5IK8I_R!"@"1 Q>!^[>-.I+KW6^X%W0"!U=$)
P>]28&V3,+)^;_5K J$ZDAS+)0N_-AB*2GIK U-@P$0DG9VO12ZL19,Q12A(4S;\-
P4Y+EA8U"+@)1L?BLN1-OIFK;U@0CF=9W0SK>;PBCLS,TFWZ&<&C1$JY_8BO2SKZ;
PR+9LOIZVTC63= 1E(O=-#'0$%[1'6@#/M*J0=;G7N1I(]E#W5"I$BT0_')V<WB0T
P\@B2X6JBVH^NN04F*9DC];.WO[7U(Q5(Q9Z,MKB5QC\27-C*,XB:O'7\**JPA].R
P57L*C(60"^;UQ.HZ:R3L=<3&SH2<FZ*E_O2@" +5DS12R,9*)'18XKO $*N?/ 27
PD^%*;O/F3MY/I0:@![E0DO-W2A.NL<7-B)[' =7PFW"4BI5HVT4[)RE-E8S9J\W(
P!84I><B#X!$_\5,O;/\>A/,^3YK6\U[/S)-KK"KC9GC@>BWU2X8*ZI]P>( [(W+-
P&_1!Q53HQ%\+U"?RVPOY?A=>-\]GU'KRPH'F.[6XN)!A1I!QEW=%6^ELU*IM)@=F
P)8P020'#YLN9CN@C<*]E\VN;2$H_-.*H.&'.A+J1NZ^J 1/N3"OI3%,26ZW6EHRM
P93#LE(>:;; DC&ST9[[VH*0%2=.Q/6;%X";)"8;TS&M7K3L,U#N !B6Y#0+9Y1_6
P@C_X"&UA\FK#]IP2ALSDBJ!)2=(_$-/7+NWT8_QYC)=X;BA!2'63]SA>/" ,4;6C
P>P9$<EX_=AZP]SH_%2?N9+*%&D@.,J)U #,KZM+[Y2\L@FOJUDW'HP2[ >2_/Y)^
P0H12C 3]#!#YO( M^1B6@91YJ)EX,?90)OM%*:NDWUOX?8=K-J%DN$B#B$!3H![E
PHE4)2>LJSS7DVQ2'PT'O=!DHU"K'2[B8O@#F]]TYO6R9Y;IKB4!&W834G+<?Y,0Y
PV*M,3^TW/@ "TH>,A-,%'.IJW++#L!#%7VM6HNI$95%>P0KOL2"7+YIGOB)9O%#(
P.JMF)I9F:EL2T?)7\;##ZS<* %L1P=H;KT0$?<U#QE4QJ>%;M2)4GZ]E>2N2>!()
P#]@T% QF"#J0!ATX:MS!73JGR64"N+JM[F4(B5)L*UU &X4%6O?\NGQG[JA2VGV\
PIE\W)/$)SKK>27SU MT5I1B@V4YG:',H\%V+EW''KB@*$\:/>3;'ZB*NN'SRM>W8
P:EZAD500$[F1M;K _W[(=7JQ\ >T0[80KD_SH4_ZO31B_^*_]ZPS9!)-)$S)9])F
PA"LU7Z*NN3AP_9P5F$@84!Q)PB,K&LO;XCIY'.&IWAAD_]R=5M=@7\BN7/5::X^>
PPD/Y?F,2D4(,),>])\I(-[#K;W9+P$>VJ%7VA[(WL7"?Q!K&'\2IK-S!\74,M*KM
P%_+-1 Z[J-C E"6L3;UU8PYX:=4GU_7R0;\8$[];Q\-FB0&O>^Q)?(T.5W;@\]D!
PU.%(>/=%,-QMX]\D? 19;8(D+L=%N.>70CL1JO%W,M$V*N%'\@@ ION>'YUC3QN.
P2\=#R[F,A_5]8"0^H'#.2%"9;@B@"A9\3$)/0Z699RX:Z^+:FG?(8MI*7PV&@[='
P(RQICTNJ-"/X8\J>?=1&<?#O@L_DZFGMTT2 >GI 0NOAOAOFP-V<EH!&ZU*! \K1
PC9]<JP#N EUML,QQ8/Q'QFR%)!K69GU$5J'LOST"\PM]%!V<D:BLT&]#/N(+Q>:.
POUD7!+.3(2[GB:U>;)[Z7P!\'L[/I?980+!Q@>]E)U]N7#^%RU4N**$""G;\HH1J
PSWK618^74EPVQ6N1B+4E5NJ0Q./T?](YTLW!8')#!&>$LUUEK1H4V6^;.&0Y<RKA
P#G\U@MHUBL<! -#,SPT.!\KVP1ES0?ZH1B*P:3;$K0<5"7J.=N0=@Z6L(AGUAQW%
P6:%,?Z3NI/I(L4#;\T@]#83JED0E%+OPM=+P1T[X9!N!QBE(E6C;3H"XOOG#G&\H
P3U0 MJ9>A$Z>(+F$]ETMR7%LK=C[X,7LTRHN-C: '/W25*WN4Z!?])A$T>-8T:WE
P-26>6CYONL;S<YY7GCP?D'$@@'-%&-W3/0Q3<;6X<R'-PP%LNPZ''Y-LM0:U$]YD
P]LU;[I9;"*;8*MM]7HEK/K\F#(\[4R>22.$2-2OHEL4K[%;SXF[T226ZC,9'P+L=
P6NMXM$B&LAY_'X.1&5]R>[P&7[,U85U)&C3K[J_UUK(_I.I]Y=+5K=9'&'ZZFSN1
P,V!:VF]*CO'1D?MQU0K<?<;R;%&NE)BR=&V/+Q?F3$$ Q[^F=JM0E#AUY+@3,<./
P;,5L@)))N>'US889!(7.]5WQ:9FS>>MG3E<7BK"MP]#<L7,\J@('=:1L^CDWOR\%
P/QP5@/&?AWW6R<%.X2*G<M&W<Z!#^EGA:+_FBV)]0V!?LQZS9 W%'H"TU@ERV;'3
P*W;6"[W54M<"[6:EID>EW?R"08:E^^SV@55F)T&)[W_UOA]+^99FP0KOVBH9REQZ
P,A:_36>162^!JQB>J/0D8+NAV$5MQBN&XFJ=4X&[@I//SQ^+_J2]U)/I.#DYF;AN
PR4C;[01KM+7QVQ<7$71"YCEYR:@&3D8WW;ZH9@$VMMJYZ@F]H:A<_?'YZ('&#J&R
P]P,3E_*X\YK.2(-BWNZH(>6@VXOF-&$X,GD]X%CZ_$>D,@M6 ^><:Q# 2D#?@WR7
P=K<UQ>-F-*QT#Q3&:-,.BI*JNBV4<XY 8H*OB6R7IVV3Z#O:5K:[SXHYKIAHZ,5L
PI?Z:3^."/&+$EI+-*D+9^@@#;N:GLW:UR7JIV]!\#S45]/I?18"JMNM(P?JIO)VB
PDE2:C4VUM$?M-[/W1Z?EVE;HAT#6K&+^V&5'=6\OEU^S']I+! DJ-%DMH9]S1LS]
P6942EMI_^!&K'Z,JB0?[:OE*A87B_8)GI*O"MJ"T40MI;W!?[3J%[BM-FBWV(B9@
P@0O2><_+ Y\BO*XO[W@H=5\TK!\/]_\&($R/<P*W0ROQTJU,0&&]8%($?VOA'!H!
P!B7QXT N4LDGR@HQJ>>T33X<*-%G$38W'I\8.ULBDY$ +O)IE[TDV?]Q_BIE9YK"
PJG;KN3H)>T?)?ER1WMN#M45L )G>)LQ:Y2O:$"'D7?[!PF.!,6EIQ64]GW^R^_F2
P@62!_9T$=I'?F'.)%YIF ./OF5R/$5R<;):(;/1XUHFOL&4>\ZK*//C@,F?',V=^
PBTU;91[W-ET=GI3-10ESLZ%;]"_Y-3'F5&!S#3D26-3E*F*D=8@)7*$CZ[3R>PRJ
P/%GP&Q*NDBKI??P,[#74I-?<%?FIIKF3C Z@^IZ:#7D4SZ:]J>E$S=;^( *?SX8*
PG&[J*=HEOL_3"Y4E/@;C7RLLMK4YSRD^AFO\7OJ1=OAMKC*-059BD]PN-O32\[I;
P0BB]\+]:/ZU$ZH&C-3T6#JN[J=@+UM!,Z'>7F75=;!,MV0A=/\W$:VSUG;J'6SFF
P9#C%\^&0GG"V61 A*9T/TH83$C?>N4][RI></H26K&#U-B>2+BD-AX#D4K)C(:(5
P?/XU,IDY[V+:8HLH7X]+7R1WQU1<C$-#3$]MM?K!>-JT"O^$S((<LF\(F20*F,4$
PFYX,R(-(,7-YYI:-%0Y8>H1_O6]V3DGLBZR*'4\V.S_.=V 07<GI-P/H]6*L/I[6
P\S;D[.TL+8KR7^/(R[]WOJ)H9?7-:8IE,C3 >'T+V%T2\XF4>A3ZG)ANM"CA7) 4
P<A[GPX]Z(Z"2]%QGY8S)T^>&/M=J\T]6Q@63 #&ARJ];G[O._!=$EUWY&W=R<WMQ
PB6GCS:9[0>\S5E41+Q4!\C<RA%I96 P5U6I9;7O_^[^\#,F"^^>#H302R=]+,,&#
PWH9'\W/*K(D] #+YZ:-2"*Y,C#9&^2)714MKBT1AJJ+HF63$CMXFBB8?2>-!*2#X
P%6-O:-)B@]RI/$:FOCNG=)PYO@PS,:PB,W@J"D.2E78 7=U%\UCCHVMO[H8I7.LN
PHE1NG -SLX@AN:.R[ ((SBT?4C!(EHTC(^#"U;[LE:%_<U*^A3/CR@R#3*20/9A9
P-)D:_%%!E>)KB].A@W,][26UBG&B[']9%DH@"T;@!C(_PF. ,OME5<+TZ6 V^Q9?
P//6YQ^J!A?.O4PK0[W>"-]S]I%E[=M8B=9-Q-X&CM)3,T:QGCYU?J<,'D0S$?\OM
PD7C1-P\9;@"ZFCD/(BSSHY+P]# D3JHHK8 *-JX1O =Y("CWE4>2W ^,R5".M(YN
P*6)!T5YBOU>6HB]6T>?H5016<7'_<!E]4C,W8$;6A(?.&+L&\HL(]76N=_ZL8+?C
PWH',7<YC6(U9H3T!S,#VW3,NZ?%:5S:V52/QOQ*]>"=35^>L8]A06WX^7O[?-RC'
P%;C,GY5"4R=P760A$C&9G>DF'Z0&@:SJGLA#_.(M<[F0WW=$,B?L\:$ZOUWJ>R=T
PM$M+;_A8].M6[T$1^W19*?!!H?M<&C!Q;661V/KN*[SEK&)'=RT5J@P3>78[W4M/
PO?!X3+2O@"V'2/._8$=VWX'9< /6.T&SSGF330!*RR:HB(92T5/'VUWN^)%-0Z!Q
PAACJ>8Y9T<-"CO_\G;<P&=5)$T""+:(>0HR$V8.XU)W$"]SZ%SIS)P*&RV"S5B(M
PQW)4"['$CSX,I\M_*YH^PD:$TSM(//!I\#F#A [%X3B@!NL)!?G"W<8YU:.]"N:(
P. /G=XI*Y%IR":.'E7=+]X0CC^\+'A#5G4%'5/]^@WU04N*I:[XK(%)Q@:*)H]\6
PB-FY[@S1Q9/_I#VEVW6![LBQ%7 >@BW94U\B_C"Z= V[+PWU#<=V[#=<B8Z>D'$?
P!#;2+488KTUK+HYI)T;?AQ]R+C+;]M:V!:6_F@Y7CZ$;I'7EYAFI;439;\^-GBGD
PM)-)58J["E$4EFIP;1%)++U$CD+LX@2PC-M=Z5,7!U1**X,K#J)QO,GWN/'Q8D ,
P"$A,+('/2Q*RZC$L>ARX76$B\3JP%BF?ISVEMDCK66%]C6HMG!/]39Y(-FT'KD@@
P2!&=&8O1G(3_WF=1Q('-OS&&BVU8;J/X#](KL%?7H3RC"^5_HYMX7BF>[D/\1$-Z
P1@LQ<UGK7C/M"]DS4(3++Y['N05+)17G-26VK6J<'NC6]3"NII*!:R2]^R?&Y'M&
PZ?[JK\8LOJ"QD]+P5S'*38WT*!4\8%(["\*EKLZI$7FFR/7MU*#-ZW9%"(&DX^!2
PLJ.6HOQO8TL5I.JDW \B!M;I_B:V!%%DN-4!L0N\;9?+ASGSKR("'K4M^%:PA6LU
P]"28IXKR"XC$8_*C.-V%SH#'3@WP:UBV[J9(;"N%F$(&C*TE9""1J#&O0&9-%WMK
PT7$690&MM)5$]Q+PD94J;H"R*(LJ@/"&$EBH"7320<>4I_S"2I,H[*9'GI+)M.A:
PX$3F-&($U!*M2+:"W\%2<*[ORW&>>FRF6@?ANO PG@1?.F.CQ/E(H9D<6XP!N'0O
PU1EE+:DL>BIQSVTXK(>1ODVO.\X10,"UV8'5T42+C%U4;YD"%$R!7\W;<NK.L0'>
P;OS\K>V1*F5]Y?ARF#Y2H%ZS39J8@058MW]T)/RE+-_1)IKQ1R3K'+@^.L7OLY2$
PHK(6[[3ZI6L@0M$#W]ZG23$S#8S]'++C?./C''0^8T^HI$A?DV>R!K*5@K(@2!B>
PN:ORXZRT3B]-,Q&\?*)G/_<MP/72(A;DG]9E$_Z\2HXC<$CWYV'/:<S:H0>'=STL
P.U,FV*?Y3V^$F?SO4P%4N-8*#T4GI=,V[\SW]0!#LP3_W$5_S+TIZ)FW-6@"W=G7
PH& @Z[(6%19;[QI8[^NH3&>\87XNPX[J2BK%[K2=T6CB?;'[+8$1Q2%Y23$S4.OE
PN;L(K*0"CUM:X5L1S5=:W^IMV,=9/W:^'/USUIB/XA\0P)9PW-Q@+Q(#B(,C9) P
PG-4"8-(/[]U=I2'EEOK[^$[RZK5TDW65\0XWUFZ_5^XW ?Y9F@,^7M@XX_MV24_=
PM[]IO91LW.9G+"++<?V(\XX4/N9,+BVOX+^LY67Q@:R<-P-U#(AJ_=+50YHUI?A%
P#EX%)4\Y;,"1EJSFE<HI ^-12T)BYUQ%Y!%;+&-M#7F?E)75/L@LV! , 0@!7ZW>
P!^^+[5^3]K]=+QA@T@8019OK*]H&8\CYGHENRN)E5-X_C?R@F]3?3IS*0[\>\S[U
PL%I /A=J@*)@<!Y%(>G#;IC!#=LQK,]3LJ%S4&+-BU> W3#2H_),9^K&*>+(B3QT
P2';88\Z//<79O/AS@H]O #,D-H1L!IAO%4"L"R7(!9=ZD,M4SM=XVF!_!Q2TZR4/
P $WFOS0UFZD!H#OX#:^5>K6*;M)98G#G3D :J[KA- LZ!7B2FY1X+N##2 /F@-CG
P(UYD0&- #);0ZPI9XQ:_#_A*FHX#L<N&2+)"X"Q[&WOB=O">M+G:Z8REC^U\T% *
P(-KK;QS:'_YH9C0QJ2HL+ $%(=9"#DQ7C'?F#=C'_]'SPAC"!3.)R,!)6:\M[RZA
P4W=Z7MQ %'+0G_1)J;";9$$*4\AX?^6SJ=24,?IEG8);5"XS<=&8BP;K70OMUY"3
PX+8_UQE $!$-S7"N-@4/KRM4!ILFVN [K.Y&-&=NB#SFGW1E]5_ $P&*6MTD]#L 
P^*F4CNRDT@R&(E_ TSYKMI\_L^9>;G3D)*1,UJD(PX9VU4U21'AO;?$*Q%B39YI@
PX1<SWH(IN<%XCN_U$,E9SEKPCZKV;RV,D?#XFG:&%WP;0%=?P3R_'/;G#^Y6:WH0
P^O%_#BX.6%4R-N+D]6IIEPD;XBSDGA<:J#6I" 4EJD";4,U3KSH0WKE(Q9AL2+WG
P37"^E"E%9<3GPWN[UC*X E$R]G:QW'ML/ZM5H[<1H4-0Z9V0Y^Y/N>[N+X7$K;VK
PXL;A;J;BP.A/RM:J&+^^9(V)KCDTH!J(3"0P8K(O@%BKRUM#_D81S2JH:@W[/P4_
PWNLGI9UM%LQB23:BL.^V);@@(!03QN)[0?\J&B#BZNT* VHZ:]4S>#U.KXW4H8$1
P$#)BK?&O<1%SR0AR?1Y:=9I2*HFTNN7AA1]-=QS;6V$(Y-\?CKQN-ZQ7(>R&9O_D
P0H!+FR2E@,HWE3S'?;H\692>\N+]%#K':P*-.Y 39FAPKH22.LY,"=* P!K[*T+_
P*(1G7[3-N+5412O7-4IRG._#727*(<:6UDA^KLUY+D0D%!]17+\@/A#LAK%<I? X
P<5S1SKW!)""FMRFZ=?W2I*$.HU?K.+CR_^('EN-"U*8@.J,.-4PG)GA= -NUF+-)
PT^F(?&JYN6<L,O9E);'PGJ!#=E>0XV93Y8EJ>K1X,+4%)(@P:@7/ZR==971ABH\)
P0OS?U#EA0921/D\=%EOQ;= 4B50S.V_XR7M\SP<?X1[%NAV5AF&_6 B[4TS/QKM)
P2L *BRA1JOT3=#))35HT34\S9D70A(3XO=_^>.V"V6@YLONM1'G+0O[@%E&*>MKS
PK(BM^;&!,W>R?$&\V'"F:962Y+YN=U^3QB](@=GL'J'OA91>BVH6H?* GQY_8HE_
P=#@VYTEZ#L)BEO78>J>3%KZP4)5LMD/M[,,?F*>UIY6#L-P7K(Y0+WZ $Z<DIWQM
PE--=C5[[#13/!EJ.:Q0XQ*,!;; >L4^HJ5C'VD8M-21@6IW@SRF6VL8@I"KSJ+8U
PTH%Y QFTU0#1M)3.F70>^TLM>DX;3:+?=2G]+E$03@;1*^#6ZQ]"2("RY62\%RPW
PM:?LJVK;IYV+I /F4H;B/BM"__%_S.Q&H>MMJ&8_9&$[6(M-O)Z:(#F?&, JHGU>
PEX.1TI][Q26CWS119N&<&>JFKMM"W:HQEW1::4;1N2;XU^Y"17QDW#<OA>1?-Y5H
PUKTF3_HU3^<E91(*#F*T6*DE=)C02WGZ;T(I4=J*;6 W=?#3<^RW!VKE^P0L+Q\9
PR0FP8L;(K%BMG%A>)3,_Z8?DVQH<NU*G,Z3GD6KR6'T S+C>\9P:1%\R/D\<NQQ^
P;\9J75=^U&^!<D71?./%ODO8Z1:\#C:%WX$5MC+^1>\?/K8DY]C4B)8\9:SRU9-*
PZ_:6FZ7Y:M3!X7";\+IJ4QN7&CG,J$KKLHGZ@/MBM#\C-J(&74=RFR#UJ/7X8,[H
P%TI6^!Y(??*FB$AJ@X<. 5=\F'SLDN<[B[^J!\Y9603 2J]DOW0+V(MO&'BE%Q!R
P!>]\"CC1$7N)?PFS;M@+IBU#:$U:J>=$_%7/Q^.?#'"-96T7EU%,',7M<*)L$5[Z
P4%K:9@UMONC4]*C>  X#<\*X;@]7SP:G"9,X0"PP,!I%R6..$SL!V-@HYSI#XF\,
P@:KY^KLN.0T^6W+"':=YXG:6PE;>(9]L#^E,?2'%PKS05#O]E1[P'9\F$M*^.M)*
P.38+R9N5Z4!%N[L/2KM:$U^I[0="K/%=3HD@6@LSUL":>?P+@+;Y^P!8-GEKG)U9
P-#T$/9+BHZ>KMEXD\\(0O\"NPZG<@WK.@'.SW)QVYJ <W-M9-#2)?#VF)$(@C/UE
PCN)W\2#J5Q8=82YC=-5O\V,09 H:[$K'Z7<OVMR :[))8OI@<EA79>A)H4W"*SC(
P.B[#<<GE_[?W-\3D*K1+O#K-&)HY#D3%6EL]B5#SC#;98.[E:Y,83Q+GN#3)WA,5
PD:D<IE:3_G5;7OUM2>VZJ$/$S]]=!7C2-\CTA^*A$Z#543\X*%X_W\^3$%XGX *C
PZ%G-9\:4FL@CYRJR9(IZ07RWE0Q%_$4X*BV8$G-( 6/M#5:GH"MYT9Q:V9WX%[.&
PQUQ, N+P*Y1NF$&=?E-,JID3-E45%5)E7*OUN56?YMR8>'!B<.)@+@]YJ"'TG:5<
P3S4MFM\Y;4/_3J:M:J6 D7]V]/ MRUXF74.KQ+4XD?8;;WV8)I N%\ 1INUZ&'A[
PF#5(=.6;XE@,T/DZSU3<?<!& ?,7<!I@J,Q_PEYFC'F@R602:$T"=JNY+:J3AK9<
P_?2 P#>]=T1I7N17<7C[R7 &V:"D2\JE$U/!S,N+TLWI:YUJCL)*^]N2//S7:+H1
P=FC_5K(\K0U?.2K,&CU*ZWWI:%>'AC!SF5.=T)+(5=WXO#>4IF".H#W5FH6!Y@%U
P!"+U<R9>UWJ9O/=%=YCL3A &0'I=W;$&?GWNR?A@HQH)>DI/P0F;BU"]/U4?G?Y5
PXB3NT40Z2HH2$DI4H?_D+^#R]9'(Y54#:G=( .)%>))_;TDX2@<<0&1/FUL\S-U$
PFGX.N<_T>YS^JZ]?CU6,]$.CXJ:!X_ -9^I-=A^E!9L56[=$$\@L<[SDF[TZ7U I
P.8+O<\^YL:\\.X9=['>QKOQY46=F=U\M#\!(,Q=WX"D9A3_&+6T![#H4"DI(S!S?
PV"B)4]7N\8BNLC,?YT?Z83A1GC(;*V0DA :$LW=FG3\H[TQ,1[S)>G(>X+JZI=-]
P5RN[W@H"T^P=]-&&#CNQIP2S'S6B'/IJ"2"QA'$ZMJ^;6QG?"?6RE"_KJ+(NZS%\
P#E()U\$0%:P2K'NB\'8G*U?IS:L[Y1\!"!OH9*ZP@?+WZ(B"M[KY/ZOMJ%$5V^;7
PX\&4[EVYOBL4=,OIT4[$\Z( ,1CAW"$7(D<9"*-8Y=2>8I$K*?+?6H2H.\7.87];
POWI@OBYF)1SKP_6$ OP&A=@,1&/#S5,(7>7?I$51DH/N_R"2%H1U84M!,.XH8S"/
PYI7R OXX;O/G#H94C"8M*OT2BWJP<N,EK#=3X\VS$+AVZSJR>7^<1I8XFVN3\63V
PHD(EE3 TZE&(2I\[(*4F$NZX@>\<]).A46<M7*WGKDU6C%L,L)^.,3=%>Z/^E$]R
P5P=J?(@9Y]/GG).,;)9D+RBF2^7)&Z8!+/OV6)K*L^C<]%4]OSN.BN)KWI2;@-Z6
P?@40F+!:*Z8_IQ96X_9CCLHA\;NH9R4HA?FY;WEG]3#(UUW-4+9KO)A*5T!_T^LE
PWJT[J$]"-G<[AC*YU3A6?-3<VN$./CF](\P5]F-4LFX)?TMF@SH!4)'KFUVCK^3U
PORX$H^LPNV1GVA<J[1,?Z 7O#8I6)$+%K./Q B#'";RIP[SJKT*SX)'"52_B?:RO
PJ)M#L:M5'MVMB&Z--,TK&W8><K00EJG&\L31&>/X;/U.1(# KLI4AD/.*'[K?BPJ
P;)*H<!50PXDL\TFYV.'])M:9V:F@G3*&3Q=RN%\4XD]J6OF'A!+M3/_,/77"K;X#
P2TWFY^E^&:/FUWE0H=FH,?N80S"\H\$Y3_:=']/!X($:I+A[J,B(%&G>S)N[IG<J
P1E3(+,?C&==7:B($1>U9SGR#S@ONNAO@$/3SB'&_*%E\&*C+CC&[MEN\<>=D^.[!
PQ^[0F0;QP9#.(ZEZ7?T;^7\*4PB.Z7Q%6\Q%AU:&TE7<8K6"L0_0?E_JZ@K-U:_=
P1!C#>LTWH X5H_/,]5,?:W%K44'YA,W<*UH7S7 !EX0[KPH@]*3J2R*+"!UO=+TM
P+M' ):=>3;Y!J%.9:/P9^CW!7ZQ H=]QJW>(LDD41:!NGWIO,"FQ <"-]*P+8,X^
P7;&!MM>TW1%T='1[C20NK$!%,,6T8U.I[ASQ4>"<M/17WO.Z*T80WMURA,Q]SN<[
P@"[8,;T/)@MAY'2LQ"4Z>DP;L:Q*54KSM_"GV1!_0XA9_%O3RU-A1Q-O+/]\AEAR
P+Z@''DN$'8616?USU@$;K<X'O$=OUV<IZPGK!42SD TZVQ[HTS2SV5Q:;1=X=.%Q
P=CIN=>B;,RCZG%^4;E\B$H!/GL04T[R.DY2?0=Z/RAF97@WBS?EDF%OK>^916Z&[
P-K;7KHG;Q//YJZMC%%!8E<N(11\3>:G:;WG+/R((S8J)@;>;4T'#Y!00RJ4Q$]T7
PH4C^YS53-M=[@]'OX6Y$=])ZD^A8':VN5QYQW*(_)WP667FG.2JF=Z/@3>FU-VK=
PD5#2MV*SYO1V[Y42V1DTXQ^99S6-SN?Y\!8 >1]^L5R#W-::$NW5 ?]I8AGZEUE(
P,&$[==_( 3KSK-D#_G\VT(9@LC"K3'<@TB-J[+LV"U&M$FET7>1*>&A"X@JM^&RI
P2;$%$M9:^95B?J%F'IA82/.%NY<._4D=@<[50R8,@23]20Z:-Q]L/ K9Y(M-XFA=
P2L+2B@ECA&DL@$N]V%C)RQN@Q*-;V.F(Z!@+LM;H+3L*S+QR@#&_D4L9QE,7%;$L
P#.JC)+!P<-"65LZS=>)4*^E-/:^6!#J(9H?03S;[D^#!F&S$TN*<H$2_II3BA"NK
P2*Y3&34K:L/8%NAZT-T7USK?5(EM6"9[Q[]4PRC*C7GA0/?<OTU;OA*3N,=J;<2.
P9O+Z_>]GZ-,@[]_M5 M^LZKU8YVB &=V/,,OEZ^N+?%UK8>,N9S"WYV>VQA>L=[S
PRN@@SZGSSR]+)<Q@O":+&\_Y9!]_7IV,Y_T*IU*D*U:2^XZS@GL289E'Z>PQ^F*@
P/A;^K,F1K(R_$+7:.P_Q0ECD]QX/ XUS/ 4GN";A*V0J1!'UT2/>\0>FQQ)C\?51
P@S(Y5\1=(N?IA:&\"O4(6*13\/(]S&;%+T;C)T>:[,5< ;2(#SBRE(KN!VEW: <F
P6!EIV*)1(GW<F1HA=Y3C"C;NXC4F;/B7@MI3^URA^NAP20_GE6=%N-!_@,")NYZX
P_+[/A%&Y]DX/8ZB0@R=U*^N_O=1N3F^KZG_M3BLLWB:2???-VU@^@/>-:?_O$6HC
PC0C;P.!?N]\S-2#60<^DA.%0FP-"0E?Y\D?5WU;PRER2)9RC+T3)D4'%)\2&87EF
PW.7/;*]L9^6%</P3OEB^,."0JOJ!LBEP\%:$OVW8."=UBY3>+J/1=@2Y#>88S$:(
P,1IQ$-W@CM$XWW2//@L0L5Z2".&)UIL-&ECIDG9XNDE;<%I#+.?V\=PBWFF.QHL_
PTUZKYI9%T^VGX@[ZRBS!<E68>QM'O!8@8)\O(@#VT5^;4(\554"VDF3:S,U@/BN&
P% RE54S.35%R-.ZE+Z*)N?Y2UM6CRP3TE%'E>$?D34YX<#!SNS>?HKK&4_+3\"\)
PR'O84.87^/($101<S22RW#6/BGSOQ6[B ?9GB"(:PD/@Z%RQ]L?\2R\R'CK5YPI3
P5P):7!/)A+D5_T+>#4X3K 5,O;H3'B?G\QGB&T*7[C]'<---@EMI"3F"]"-_O>+,
PH*1&1_?=W,#FT7\6OKK&*_ O>.)@)@!< T"O^[^ /L >:G+UWOXXZ&[A&]H2!:1V
P:!#*M7J;T'S.PPCNY5O&DBN3:=]/*:^"G8PQGE%-U+/'0A))>B>7N,\.]F$,%5;%
P+?R?/'G$RBCKG-Q:!V6CC#7%K>:(JU<R0K'%"XY]"O/F[$)W&3(<!R$'\]K"\M!#
P3F.=YMSG*-[[+$_'-SM0#*3RK_,Q[*+QM]#9F:G<YV?-+@DJ[4>)YEB%_W367<C@
PEL3]XAWM%0?YR:ZR^!!,JRQJ.C#:_8SPA$,9*@R"7,"#0+\G4*910=URQI2EX^CO
P4VM.\@0RY>GC524RW,SD7[+28AN_CW:#",X=L%=#AD=P2S3Y@A-I^_M&:]>F?#6*
P@6M>55I\(/[I#AM\O?KZS%D:@/?K7B.6#N=5&CQT-^E=_7-9+-,POH-%LK-R;^D;
P>^PRYL917A,\5WBYT1]K]+_3M042&GPKW=?[%7'MWA;I[&R=7Y:+Y<^^3$IT#7@W
PM0N#D':I:KW)6YD3DA [$J06P@+'54A9K/@74;)52"3]9H&()=OT"M$G=I5#GU[+
PQ'S;TOX8>ETM4-;Z_RGI2#K#W4D\EPSX'@@?6IAG"S+/Q?['@E0\06W(?PG:/(\E
PWNK$@L"("HWH46AHS9E-? /$#WD3O^=("XD!_O5L- 1T!05)EO['A&<,7#1\8IHW
P[!)=><"*9"2Z]UF7(^E3_O9E7E1%.Y8J8,B3%;WV4<%/"?RJ:3C4>\=NS\U/3M85
PDU# 1U0=*.8;4IN%;+<?M*"]87J#(S H[FC1G=0)&%2 +021.V7T[)%JPW!3V=OG
P4""/2D5Y;X-^5P)!X.SAN=4U,VM+E(L/]K.-E+$@C)SNC>:(]3M <CBR:TUO",I'
PCT<4A?B,U<(V7SC_(-5@*UIHD=\0^M]?WEQ#H(LW0?^1HS1@@1_#F ,+1#K"WE-%
P9=8>W4FY -RT,4[6<#-(J"P))K@NP-4#2,KV#B;F5O\1S.L1P,64_CS]2J^[]T$E
PAG5MJ55I9H55Q9L5^EV?\AUR].2;: _D9>#MR+0M-L>B0=5/M$MPH%J4K8S3?;7,
PA(EY<GK,4WY,M"!JYGKV7&,8G_CDD7?LD(O%D9;%04[C&1"T$EO+(,J6RGBA-M3+
PK$X*YU2@%A695P53:9JL5]6P*TH$<PQN%=@.G,%X7F[DWJ5V>M<Q0[=+7S$?(U+)
PE:=/^O0$^OE3H(_,0GC;$ PQVZ]V;3PLGKDOV)0.[.50[Z_-/MPOB]G9,GN>#_!E
P92L-"688K"FWZGRYKQ%/$[A11[D"0>"%D>W^6)5$C2SK3/3V3 3,ND*Q[5CKZ:J?
P 8W.7FV+PUH ^4A;2R8=CKB#]#JR4TH_*PPF@0;VC_Q5W\Z\/MU+<$[6]WG62&9F
P9OM4RN4HDB\PBE!XRJEGRI?$TV_^@=/QH,%95KD]VA)),XW")9H" 9<,QV1H68^G
P:\CIUM4-5[=1,3S8/%5>RN3]3%L8W_V$0H=I8//Q%*5\W":*:^.$UN JO>;>Q,OA
PAK]/T57"@R USBW0RXLS;DZ,1E"B$)Y1N#!F2IB(:5-\BT,RQ)H[>G4Q_ 1UL/-B
P'I.XVX^><THJF3=0:%+'&(5FSRJ8D$S6B"5[ <CGLSR2H%"[Y%+P\293=2TI[I_D
PC[K:#/R:6O@8_A'RI#[QFL/^($7L!+)]NC$M6+JOK*M),$,[2>&)E"-@,=^:^JFD
PZ] GNJ:YK12]R":%EJ "?+0.PSFX#L9S#CA3(*4Y'-I?2B;YD$"+_Q$UWM0=&*DT
P&D=NFR9@RN&4P^_IM_(Q$@#@%!S >WGZ@!U\"^J,2J2Y>]![QSD=NWN-WQ29L%LY
PL,]K=3/J$L19S2 *O"L(& L!R[ ;][*O#^17@8MS6 IQU_K']0+C4UZ6\CO4#&5>
PW\D+)^GP]28'Q')4> P/(L>@GN' KL-LDW=BZF#@G3:J@M]GI (LB)Z,KA!U,5NM
P@>+%R88S@;N]%R\1@6[A3B?7&11L];]@SNCE5#91>X/+WL$5'LX4EUH/ 'Y,SNA@
PN-8A(WU\(FI@P^8@\0Q;T&ZNXC)^8\GIAY)2=SVA@0'DO* (\1>F'*SZ68@<;B,-
PJ5>ZW33O)RL35G+/;08P)&X^\\)10Y*>6IH]0^6B;X*>.FF\96+L(;Y-TYI:)W'H
P)T:I7:Z0SU]53@YR,!^5+3*1)@"I5#M/ E&C4>VUCPC)J=Q\<'$Z.K":!E8WB!"B
P_CB\Z6!'IF(##6XJCRO+T$PMC&"J8I@RM1VC\TWG][<R!3FGXZ>&&\I%\^H:2+7D
P6V6+NRO:$2!#TY8I4QP_LJ0.\GO42YY8M>'[JV7:>P%<"/-C#8DSMYTX0, -5!<J
P)^@16Y/.XIE[2"OR;H).M.T%8C78,A>%*L,: .NFJ@S#3DIY>P0KBEA]DU,2(<5\
PRSR\K$QA["K38I3'7O<80<T/A83Q*V=*8H2A*J1AL,@H92YW\Q[(,<%0W? 7&(>-
P<V2WB)0@JX *[N$ G&*CH>14(!NI2><6UZETE2"C@85.L<;EOE(8-0H#K@F2PN,#
P7V+LI!'TUZMYF,E**44B/@N*4':GTF.S#L\\V1KNI@KZNJ;N;+</I!IQ&"PS (_R
P%LVF:'X)LZ#(GZT/4+,# '.4:YC=9VXB[^_]%<!IU:DZ*4IV.Y\1#<5H#6]T?<_V
P4DAD7LHVDM ,'AEUC0A8/UO6?'!'9V><]Z#C^C!KT6OWQOC@ .4CE\#;VTJ/69:.
P?8]=>*/RB;-\HX _NBNY;?2L_7\K T=B^P?K*&(F@IQA=""OAHO@ G:)FU.WVVD]
P"O;2/A^TY.N1_!GCH^_E[I#BTR-%6OT> V%3S$F5!KSKN+[<T0EFK)>(9Q'WZ^3,
P('@8C7>/-%^&3Z2[(O-SW$3X<.J5L8\9U80B?PC"N9W-VY1P< PGS2%E)Q+3T[X5
P;HY04T]$2H,B$.[;&V=9?RTAMR?F08T/_::098OX$J<#C1G(7] ).<ASI)!BQHWP
P_P* T!5O/=='&G576@YJ[/I>[(KW_H(>2I<E07XTL'PMW@+YX\;<NL@.TY#9, ^,
P=G0<\KYXAM-=#+] %6ZO;6TO,5#;E!1DJ6W^_]L$ 2UUJH(5I"R9L=/HJLQI VUX
P_7%,(TL-+MHT<<JB2.X/Y69MU:HX%'RW]A?X:":RB^1%=H/>+>,J@#(R4SK>SZ(:
P;@(V+DT.CA[2=@C7KLX=H:V9%%])V=OO0R/%NW4NR#EO"X$#W\=I7O'!G\Y^?X)5
PBXCYT^"(KB;H2R964*_H7*5:O^(J/_E="BZ?/=NHM]'77H;@VY1&2\K^8?X","1R
PX-3LS _%^D$%<@;8 .EO;=9Q33-UYR0C<,(-M -B&8COZ\:>Y^(&BF<^5%PY-.E?
P8;-NYIPAGJ&^R4:R[APXX</F%._G)J4.WPHR_FKL"I9*+-JXZ_$1$#SZM8;4QA2Q
P5 7L:GGML@609,H&AIM9#J*_K4<,,M'.5RZ>CZRC'LA?.'^CSE!/P^F&; YHU,"O
P)P(RO0JT*:P'D4N$V4C2K-$<C$XG<6667&O\JQ1)]DA1X1W4W @=+-BFC*!6!&/I
P^5D:ZZA4FZGUP]73%?L@.V-4HG-'"N<I1WEOIFNTWN]O#F"K\2&*0," $MTU15$ 
P>%(0ISH%NXN>\9.DPZO_:3\ET(< PA/8]L!.RQ8RI9DKW1F$ FZYR7P-94\9$MM%
P$0,,'.-T*ZSZ_+"43-XY?:E*A&CLT&EQ,1M//8(I;)K\R0":T-NGJ&Q=J&1YF>L^
POX.1&*$G&=@%,0@DL=*!>M=^H0GPOQWR-&+5HJFEQR73<2<!/1<GOI(7;UTX;2"+
P;/&XHB-Y!4<OBOBK+5VVJB)3;:UOMH=!X0@ ,J$X9J+UZ!9"1DAQR5E"*/G%S*^A
PT(,-QBRP)05^HW4*!W[(ZKUHUHU.3/<"\9P('_(9[/J:,L2P*]&'3$*"7%0Z<1K\
P(KIJ3*XF7V-\"UGL*DP%*:W9N$%%.#,QF]M/DA>"0*DD,/XDF-2QG*E!((%WI6';
P^,MVJ<1?#&/9UDXI\G#"TY,[,ZFB'(S*+NYE=F,5QP[P\#E?B<R,#INP0+BWS7H?
PJ=(T:V7:+GNR)A9( MMRH97^MG0WM9(#8G%NH%K)JUR*>.RNX>ST_7AD6T*+)R,9
P+-&(((?DJ,T@V_#F$WP34#2\8\LT6Y^PZ1UZ7-56X[Y*HFJ(YL6Z\=+]/M!LD3S%
PK\S@GWJOW@/J86DF_7'Y16BJ]1^C2-K&UI9G4N39E"/1K37/)T;(U@<$2C=IFX$O
PBW< KRO-EGFBOINBK"IL6Z0U*, LHLU&M3+TP),UI1[O$!2OSPP]ZFPTR#H\12Z0
P;)V:#SP4T.MJP23>M[LHB8J8W/\G.]>H4?F?V<RKF[" K5V!@C;45!L^^>A5#7%N
P_#JBI&^V4.]E0E3>QC%9A+W![%HH*M NMC?)N=? S!/@EFH)3.9!,VFI;&CFT/<&
PU5,JN,CB?2C!W<%=O@HK(6)=D,5DFP87)620'(ZB>/KT+5<@YY5#*L>X1L!@M;D(
PLJ++FNMY==)/GMX+!71%$F^8G\O%)4L0Y;D5'1,:O$\!CE*^5@';B[W0K*$%*Z-;
P^/6Q\!&^=X8E/SD$ST]M#'CQUSL_1\@0^\WV+ZK]AN_^<-.-+P?:]Z9F)3(KJ 1M
P-_#*?N.']B@6QA?T>$!C0'IJ3 DF/V@6TL[XXP:)((UXZ0CJ<J=V5"130 T'"3[4
PO/7UM;N+!AZ1$GIV7VA9A(%QAK0<1\2)I;/6=X9..M2?^^D9U1IIS$XNS>O4--\0
PQ>NDH8#UW^&1HPVGO-,F+SVK\K%D8H=6!AKV8H82!,J\6$>L!DH?'IX\LS>%?KV0
P%?D+[^!*YW*GA=@8N^<.G7BNMQ/FP2^7#1+&KAD&)$TWD;EK +HOWK?BZF$L7ZKY
PAJ(TSTY"^L;4Q(533^J9_C@PMQ*ZSD7-'/HT]@/(276:RTKA'4$B^6^NG#:P+<2*
P=PJL2MGQSF;')?VPKF#?F]#O;[*JV:0Z*+T&2$B[8 6>KJ>#SC)5=3*I>$0:F\65
PU2+^)YZO[Z6J_?%2F:Z\BY6'P #,4J@P>PV?86A!1)8# "< I^P=_JU6LP*28"#6
P!:F*-J*@HRK6:\%-S:>:D0!L*#GDS)M-]!,9* ZW%Y.0?TG4X[-8)US-V<;Z S>K
PJ&0"XK#-TI,0O;]ZZ=8T=W[(^_K%C7P5Y*=P%9598L>X\_]G&+($\TD4$!BE%  S
P\&035PNW>8]('(LJI'IV*1J[G[,GZYKG8I-IC,.I\LI5M1=AQ4C JNX0W6433K8\
P5835_RX38+6H!A_ ]"X+=_4_#PR\R2E^-UA#B39[6B]%NH,/5)CU)#"]W_Q#M/%M
PILF*MLPKI*MTY!X"08*A5+=H1KY'8A8NXG=_?34G0!#/"QWP<RF>X<QF;'Y#(, [
P*$+:TU[0LQ_M:7G46C]T#9%PVG"]/UR_^5&0'U@+<$E6NUA*+$7DE\T.>D:33K@R
P/$<L?R,1SM"TTV;*HN9:8M(_'T3$-_P/VA7+\0O#'SB%H6!1P;\>.P3(X&K>NX&2
P,"K'G93*KR8SSCA55PIT>!O1'XX_E5EFDOMU8O'),Q+J(K'S!>&"@BM?3*7*<SW\
PL0$RN^.!?1/P 5?3O+N2P[W32Z?@K.B9Q/MH[/_+5M09\V%RXK-AK]:^\B 3P9W7
PDZIV09>#>IZ\301>))'G]B$$\Y$+5&.;7*S90.@1SI,8H8(3-X7\9(H_X%.%T#:.
PM(>M>W:S6%EBA K=R-Y,0+*85B"6K[;,BL%!Z+U:]ZW+1>FCJT&P4)>8Z $KLP-4
P9KN-)S2?X4/WY/B&#GRFA-)^@*P>(Q&KYDJA<0!1RDZZ[T!'&R;Y]7[A?*3-EMSR
P>+,S:M.=3EG?+^NT)F*Q..*);ACQHNWEANE$  I$6Q-2RJ/DS^5=G#6MEBSM>$]-
PQ"C*A%V/"8H$Y-%'J]8KO$A*V;HC\DY:.?!AF&=IKN&#-^:[B7_J:O%WWPBYM6@B
P8<#%92">V3P@3C4IGG5 +TN_FK6W=H'> GV#J"(_=W<P_CV.A=^IVW,-P+W8"EU<
P-@-V?D\E_ MQ!+5^B([0G7R$DJY-VT.MS LQ4*FY?LXX'4UMKO#77UXDKSS]#C+W
P-%[T!;A:EH.'!A.7 >L7Y(JA@*ALQ^=(PK*,.EC__]R0%8>XOLABP#E_Q1.-W5=Y
P,FX'>IJ_L7K=A. 32(/>4@:S'IF1O=Z!$ L[QD51.^^A&Q1_&\P[XTV#3K'V>SL(
P&*:#ZP4@:TD0V1FRKDL,2P9B^U-WVP5\HNI^=85XCBM6/E)!=R+M;*YM-NUBH&\L
P.9\\,%BE32*^<1O8VF;3VO7IC_>,MD5!\,,FJF6K-\MU8;2/X'(B%!5W*X=^@?7<
P9JMT6?F;7BZ?:OL!04"2P3/M;93Y_Y*]GSL/Z^2>, T7$5(:RZ[[5F#M&.6.GIV$
PXJ<2=$\^=!4J$P>4:X9'(!FTTO*_:-+3M,Z"#$]\LS5JM=\+4D'!Q^K*\N6=) %H
PDQ>]5VGTI.*;>V_T)_@DT([HZS;;+,>;[?*_]1[<Q6S]_D[R P*SE.\>_E%[FTT>
P8/_[CX[S%KB%ZH*97RMW#F&ZFB=TH6ENB1/7FBV)ZU0PZ#AO$BF7H( TRY/\2#V_
PXN5 H%B=1>7,5]SX%)/\K)56==H0)>#B%3.-R$L,R9=I]H1*,.N!^RQS^CC,RH+[
P#-"*>#4O)3Z&(%\ML7SWW$6FFI.Y0GGE>J'DVQ&?4D]+HS_K_B<J,[A:_1W"2>;,
PR452YF@:^=P!:>3]L'PIV1IM0X3AU-L@ZCPT^%?/MOJ7,&!?K]8%ER6=6<'85Z.C
PJ'T;'J&\B9C6A?EUIJ^E.6K9AZT 295.6Q\TN'8V5MUT\-P6[ 9)];NRTV(GUN ^
P2M@&Q_0$T_0.7IBA#KX]YE&[B.PS*V2O^Y/<K]^Z!-#,67S@2:\8EZ [(Q1>FDCK
P4Y:0MY+GDF!-DAA<8'+EDY $9TRPTV%3:C7BQ1'(>X@,2O#DE]#2&ID]%W>7$Y<\
P)DO9?BI\4LP<];0)N76[<:]4$#>Q=0?-$!:A0!2KAN-UN*<C"T&<N5M6A],0"!S@
PL#;D=R6H]W:GCY:P#QI*Y2KE8W =:O/=Q@.^3MPB7/<Q?F^.R5O#H+'X>B_'9@:Y
PX!;K*I'1C:6E\UJ$*9G[\B\)1Z)MI=^B0V>)[B9-K:9@L=VIU=K.?26I#5PW;B*H
P20G=NM^AYQP$58B18XN&K5B4' K.>.\O0QM=(_!@;,GE^:DL11=[DI$'<?],*F1O
PYT@1#?*>'<R@U)Z.+GMWYUY>IZI]D%JEVW7$;:]EE%51'3^>RQZM@[6 /ZMR_&]5
PLK[QW$'2.],3&3.8]_+Q4'/X;7[XP(:=."B5UBZ :JM99M( %Q>:O3J =V@*H3RK
P^:SS@1%OI;PQ$75-Z-DA1#?T@O3JXX81)!D"J?9$G;ENW>D@T)*3:TAAW 8QLI&P
P8O"];W*,\#91>/AH*N[:;EELX;"4;C0J*;K(*IEA5B8'I_% QZ@LEJQ^OF$C13H&
PGPXT'?,7>H("@H&FMOC_P(\YF8()&& N$5HM +5KS^4.8&J]C]Y; 8]?#0^9=TVO
POVL^[6;&O7I0T[O 'R*Q[<(H3SIVM<,Q<%NNJ9DS*-!.6[957J+/>#C3W<5Q>L?A
PA4K;F[><P4?5I#R00C>=EAO\'9:F31\4^O8)IG DX"RJS 7WT9 3_:) 6.7:''12
PYP=U)(/NT1M&L1UX8>K-+@>N*[7 ?][F<'I)G19L1I,]L"QT?!^Z=,-IQ2EY;H+A
P\:NJI=20BDG!/2T4#EY[OBL#Z.7\,JD"S8MN0Y:-!D&K!MB'#NMX:5BF!--NU.#,
PWYC\^)$/T\ST#[<4(Y#$P:%39<6JHFPDL3O+ES'QG7OWLXYFHB,+E-8KB6GD=;6!
P%T2IL YS.3 \\COE8XO:^+"37P AZA2?JMG@\V5L?>F=P\M0('""7*.BS,8.>?)-
P>HN/T!&Z!7(*"13/[Y&)PRX2U^Y/M&H1IKE><Y^18&7DF2ULLSHM->G20[%MKU@;
P4K]_17MCN*?SB4ZV^ EBQ2=X6I^);2_$1FW11;$H28W)@W2TQT1(V5]HT7CPC2P-
P"#<+6^M U$V%NNSOO;I0< !:L%BCC^G6VP:R3Q\YL>"%8XQ5G_= O3PUMV_XQO.2
P7=D6;05T/EMZY3?GAYP,S^([RYVB2[XJUZPK"!24HR2+X!\6H=2!^>N[I B/:B,J
P_XQ%>-N<4WCRZSAX;& ^=5\IS#E##U32%.RYDY>?%H4;?A3&.9*6[/H1>\'5\I7"
PO#OHW(TP#$?/U)P'-,C'+@_GM1OC-N);4>OLE6JZY'W/<W.6JLBEAJ_L!V.9D-W/
P^*WS?S/"$U\XY783EVFEGH>5(PN6& 0@JAK;L9%MS*A>>0+FHNZQQ_ENDC(KI,?7
P5).[YBIY@N8Y -(; O_1A(J;3[=O6K_A%6[LOU(XPDF,'5E'^"$.O5SZXIV+A3E2
PC;S-I&9S#*5S)IX\R2AGST'SIBI,5@;)AV]H#X$<XXIO>^K!^-IU3B2%9N7ZK%$W
PVV&8O,=AG__;O^Y/%/V\]29H(3P,OO6W8/[1]N>+-][IR4W8%&],I0.W+#,F&!4)
P[N'NBIZ%;0)GWQE<W!EJ.II^$IAUJ'*!A*V(R@AK8ZS6WHP WO#'V0_D0Z4IL7WR
P44ZUP0;N -OB$WZ<A<ZC^"- 4*@*M.G(((4?;NYW25SG=S)UI7PM_(A+0L!]U>&M
P$B6*9B8\/6F.O3E1)$3X0*IL]]:+U. K 'CO9V;C!=<R ?3&$WOG2(K#XLC>]64.
PZ5JR^9K!CN1(,^.N#6%]0\CE?>'AC&Y'^[MRF'TH"4BN+O-.B0*099 M]^E\J.:<
P2PR*3V+<L,!\)CN</'EQDE<1L,1?ZZ0/ 9_+C$,3C $5YB6><_6N]^@QB-X6;0[P
PE".U^<O^77"3,]:4:U$"9MA7A4!"]K(<%;HT:Y=JG\ 6QSG80/ELCEUO0;GH08Y$
P0!%P %<VZ8A*SK]O5\7VGPHV[P 2?S+)()'D"94/+=01?7=B_E?W) 5L3&+^R\V-
P1+,P3&4O2$C9PC9LD?8?0N6FMN8B)+"6<IW=R163G.9[!ZFM^/-VMT-XTVFF",GE
PU)[SD5,^,D=E%>136ME^EAGS?S;+!OUH<&.#@0:;_A-;%,Y8*%N/7%,['G@#L/Z\
PCZ=SD=$T?W3:)/Q:.@3]?J3%,IMZ24-'+PBV#8N\IZ<'SN;720@W:&^4SP+A;9IS
PK@K)?\K,B'L].#J3'B!\\2WZ_M>"V BWK;ZX5,T QT2>OZIW)F'"+O@=@DS:@2[?
PAM>>GFY^]GSR:,D8OBS ++&L]E'I(/C@(>B/D(I#4R_= C2=4!&FH*.#<7P>B<;R
P!-X'Y:;YI:$[D%OC7*L$+-&#IK-Y$&'B3,HW0C1>.+K&U@,6?Q"O$?; /&C7YX2P
P$Q%S:TQKY8VD%Y/('7\ S.@'HP0(HX]L?AYP\/Y5ETE"!9GW[?F*B+<V\["]A3Q@
P@<I]>_F,FB\)E11T"N00)CS'U/T0",,L&2Z!D8XWM$_P$G@S)#77=^S7WO[H(OLE
PQ((@;UP'".5@A1-<W@-"#3'#8$AY_V&=V._2OVO5YC"X'2+#DVUA50M4'13N.1 -
PZ\U7R3DT_0]I7 8H2QLJ(9QDZ.$B1'LJK)5VT;T[G]I2I(I>>FD??0P6+5U#0,['
PZMW1:[F7;8XH3>%=I!@@PQA_9K6TDMDGCGXH/ ^/_/FI376>9Q.6A=W%&W*2ZU\!
PF-J).\.*0I<G^P>DUZ;A ,@ABCZUE.8!-CG,/E:X[Q![1Y($XYJ;GA+LXV0Z._FD
PV1=K(.*D'JQ8D>L7,K0C_F47,S:&ES5X2.?A*=<-*G[[=WO@<%]UC)N((23H&55F
PM=>D&OMB[QD0\I0X/>LG$$?3H#5EGG> @D-*R8S&^N(1U)GUM-F7.JB\$]%#U]!<
PZ2MDUUB-;7C_:-L9'1B3K(K",O-(J5O99BYFY^.3O.&X.\=WZWR<:CJ=,:5,F,.E
P8^3"ET:SHBJ5 C/"H 8$QTF8H3TPF8>(R;-+2_8%2$8,$^+Y+-M^[,"!&Q?,X*C+
P]<N8)\N<LO,WA&B-\C#@F-ND1G7(_(O#'UUJ^A>*X-MX#NB13Y%;F'EP@S[N&@/K
P6O[#XNCW4[I0[,!<"6(/C0N;8NR5'J?7 ? "_@A1#AAM!E'=ICCI]YDK./H(_7Y_
P:J)I<,N22^9?G1R^5:>7=[6A7/$;[1<!0J[!:B>CLB<2/U"MJ_?!>6[U^L(UJ:P[
PX\-[9OCZW4^_O+-+@$!>B8:D&2>NP)J_F4C3=BXX0=BY!P]X/[,7XZ&3EJ)5];JM
P?W/TWZOGNHS3]M^Q@FRY)^N]*CW" :0!"()$KP&=9D^$V59-RJKGMCS#_-JM ]-7
PY<3O85RADAEP@?Q"R_R)/%$A[/11XMV?20B*!![I.>[($M4H7-.R6RD4^Q\)Y8VO
PJNSE9*]229/O&Y"?:ZV:!$AK;0DH#P9 5J\>/?6IY^N<"@,Y)7\O7?ZZ>HL 1,-A
P_>2AX+,=SMD-(2RT : #\,T?+W: <@QBJ:$6],*?=WU)_%*W?#PSA9-OUQT+(#H=
P$R=[;%)QUEL)T","XN3M8>^]$O"UV$L^#4'=>0 #>EX\9V9MUVE='^U>\NRFN1BY
PA%#5-S^\V>9F1\&^F= >$]E&E)CDWQR.@7CLD8/]3@ZN&#;7T+ .G+BU" Q60PJ/
PL#D3<L'3*5H+!=:P*(J%4D[)5WQ;"KL<^)S%!0Q%6EZEU"$B=B43-]\AK<2&6_X(
P\,!KJ2H9/([5_AC\]ZB:H"-F/J<AR318A8CUHJQ(4JKM(<MR2Y-I'[[]QT O)$>D
PW!6%O5R 8$8'XIM:P1O&<:\1QIW!RHLK C]MH7)]=:[YS992Y?JG(;GEEK"R)7@)
P]^'4>K55;)RVRXZ$(AFT_Z\WLK(4]TK87+>^*GAYF1))+U+B0]]C25>];LIZXM*8
P15?%N (A]1?:QW_Z'-;M5-&ALQHC<[ 5X96?-^OG!@--RHDGLZJ ,'$77N2_'Q4N
PJ)0LW")E?)+5!K^?P3F3A66AV - 0J'DA<]6X[&JIRT-<O(]^XEF#4*#O!U%]UO5
PA,3"Y#7I2E;[C/F9$K4:%MS"X;?"BE&U<2N"NJH)D>:Z=KCY2U@,,+9U]JYPQ/3:
PJA$_Y %GJ^0%\XKM-Q^D0QEI9EV-%X:3)IZ.!&]MQ3VC[$_>+L5MS<K3SA23;V(E
PEQR0,)XU@N;KS'+='?S]P;SGX78Y4P(QV(C).\0>MX=;'=3ZM-:_)<" !&1H6!+=
P;=V$5V9-^@A+%ZT7>MT,_@P2"ZYJM\^K9CFN?%]J/EN;LE0Z)T'#]$IYKY6NF$,M
PW_Z;QBG<=E9.[Y[R^"H6BQ_-/GZ3ZP6ND/S0![^W",IG_JL@E5?SXAOT%XF[5-=-
PSYISVDGW6)V%SJYHP8?$4^OU9TROH)%W43[5&$^3^O,4$*]R-?--KRO%\/'R[NET
PZG/7 -4#N/$DMX![7A7IRV; 22_36$0ZGR]Y7'[IH:<GDWRO-L6DMSKIO'L(IH[[
PY)EC)V=V;!"+=OKM<>DJXP)\>>\6?;&5]RC9W!>*?;(>E^PL9 5+[P)*/4>#0E]F
P-_*?0+0_1(X&BY]IEC?YJ%44W,AGBXZ0Q03)T46VGXLD_9_PVZF-PYJX')_GUL-@
PC ):BNM3(&B)A9""BES*Z_"2LB*#1DH#F/=TQ-@]G<8M62X,!3 ;I>%V>7^PS"([
P5+=(P]3PN=PA"$#\*MB3_(PBSUZ.F*$=I[66=7Y=SR:B=& "?7]!%*.3I ]XDA;E
P-\IJG(U<S? "OF$5[U7+S#<T1$QCM/8''&*0(4A'[[["Z5$V)'RSTM_O@+ETI(>P
PI';6DQL!*>J:D2.D.+4BYM*L[7_</(X!"52Q/F3Q><G !%4!2)NWR'XVN;H&@]JF
P:I-Q]?M(*>@TB2NQAR<^%AS!]@Y-'@?3><G:6]<$;'=1&U.2%N6WN'W1'@&.:BU>
PKEWCY6 H%P Q?X_D\<64#UMAT=:;[V"OB]YU<4Q@][7,3!='[X56[L."'$1A^"&9
PE7Q@Z![FA4A<X24S2C1Y'M:6)(HV+2=TI54XQ==%GD.3/J1K-!.$*48LI\FLL)$0
P"OII)(,BWA&F2FSG4G3)F*Z_>K;_>[-;$1"Z)K6IV0!^"7TV)G81,.FVWU8E88^:
P9WU<GYY#Y87$H$V:=DM]5.YX_0%$CIXY=Q'>DXEN]:JP7?V=%T*;?D<>3A4L"DF'
P^?]**[E<5%F4&=1QE5A5+Z"O)X9(4<,I:5. ;):=GN3LKGW2>:<)UE"IL$^PMI#G
PX<V4'DM @S4J-:G6F]B'L5Z;5!\I_3!L>_SY=1<JX"EOM/@>1D;LLZ73\SXAF%;9
PK#NO8XCP(F(0<1<M+DFW&TKU2!=KZC!*EM,^CAH6"&3FWPKE\^0;E&^742]7)9Y7
P_[8.F>S40,0BE3E;:@K6'+L@(N$,UI"GBSC0=\A@0C?W[5B8KVQ3D*J"_*T:B*--
P 1@>,4J072D#Q:E<YC_=<E/61C6B$'J8XE%Q$* -+8Y\K,?+V4/16AEL.H-(&J;@
P0,C0.M9W*E.- HL- O')L?- [I.MPQ_Q/SIMN4]8T+=R84Y-6S2#++99/Y5:5&M(
P?%6E+8?YLXK50DZQK4I+8BP6_>(D\^SOS"@K _E;LY==_[8539!^$)0&M:YQ=>4Q
PQ)WGW_1TS!^,6NI!58J'@F572%2Y5K+XWGD]1$CLVZ:DN7^6$]H06%8@)>OJ5 8G
P,-YR#'"@SZ_AS7#&O.K)I<IT7$<R>C6I'*0F99_YPZ#2U+D7B3 I]+=4AV9)_C:?
P];<'-D+ GU<?@L(NHNEY._ QT&@0P_?I[6/!P3^TM_96DAPJ/*%8@\HW:0YM)J/L
PQ[(A9KK/Q+QU"W;MYT"\O7JBG %ZUU+G/B,N&^R7TPJQ (8N%#2XE<[8U^'A#^<M
P>;@7 UV^J&4;E;Q%4R?LM0L RHU3@L]N)8TI3OF496S9(X$2RB7X*(:HS4=KUY)O
PYG7A I3-\$-!0UZ9&>7DJ@TZ),]X'*I"-39=8*;."S1ZS[XSD%%4DOU/E->-^]CF
PH[R015#.KSW\!?Q*<8T__FR_22"?+,98Q3IUDP$+J%,_Z?8#)HLC&*N5^Q^JTB#I
POEAJ#I+9A(!$'S#.KI@UTA/^S3WSZ74Y<S$-&XJ73,LEO4("Z9<+O>G_Q9B[#];9
PV2#\UDVL($VY9]-F6?(LO87/Y":3,@7C].G^&B3FDNBP2TATF[U<E3R4P@/%GIW-
P+ACG4B3 BY$R>3@#MX?LI'10W*.+31<SBE6 )>[#?D!>ULVK/>3UH\(/+# VQ*2U
P+BMS2RUI[42-MPA:RHQ.>R&W0@:3QRB$1)$38VD3[I2"%:(G9V"Y?2@\K9B=MF&K
PMTG<0#V[UJ!??I :\'SCI5=X%J,"&].5<7$(##:IW0.M)W.&)_"6 $%8M+(T+FNQ
P'_5PH#06-KIC)1([%A]4^Z=X<]UVN1=Y$5 P#X6X2=(%OIKM\4HA7-*Z>LQVO5ZG
PZWE!STQBEP!KDQ& *VV)5)'SH&QLEV<FX2@W[/F?JKLIA0@B&,F0^Y*&-$ =&A#8
P1(D2D55#H !&%)1L;EU^U[>V#Y+=V(LW2$:0.[FCB1A S&LW"Y]YSZ[TZ&W'DLT4
PX\J>2\";R,+*=(R7Z@^>[*2&_,/^YZ/ZA)ACT8,V<Q:S!TI[T9*N1$W%*PX!O$.]
P-.QD++-$]A() %U0'*8?]]42=QK&LJO516U&PR0;41<<P9 [D@_^Q.5/WL8KPJ&)
P$9>!!'=X<D1/%TJ0V5,\W6WXW:PLZI0<QD?7OR,13D3$0MXK^96H0?M;0Z7H7("Z
PURG(JR5V3T*P.HEM9D?X*2QIDA.1-T6N<:4:==U\[^).\'E&9+^!-[V#6@Z18X0+
P4%^8NC>3;?,%(1-.;7J.>I]@EBTAQA<HXEM/)EU#J@E/,$P&NB52TLLF2PI G"[@
PZ744X7T*F#^YP=;Z\Z@Z,I:]H <2L7[ICR5#^23.3QT?>4;=),*!L\>U$LTO=AT 
P*Z5GGNV-ZR8G8^&OT<*QVC)EPQ\8WHY&CVW*TB!>&HMD>V!-(45>02L!9Q-W+#9F
PVV+@L#@R&T,3X5VX4HL'+8^3FHG)EPF,'FR:+S%YAE,K-GG\17Y:0SCR)T__>97H
PA^3OQ@\R(=2_P!398I!I2T@QV2C-QA\?T!H[+5>ZMT;[CW)_K?J\E*-UE-'R6NNO
PF"G/1('W+&!YEKE.L@KFQR(X+NMK5EV8':G#FSNZ5>GK&/^PWMQ[^Z#0CNAYJ*3)
P_N;+8_NB+A>1;<70]I\H\;]\'YL'L99L*=F2^-<J5BUFND_\Z'Z%C7'/OV 6.:"=
PZ90DX=QYL0A-9(!QC YC(K$>9]&O4JUT@^MX#G30EI+L!:A/:>2O*U(+SS<;*L'Z
PLD N:)XZCXD!8%H)YO6]Z!GO^U/@==Y\Z)A,:O?4^H23\D)R6.)\]$(&$T)?@$[W
P 2GW4X3[DXUH 3WPWN43%*[%+_5]DK6,AV-!>"X>%E=_%H(70XAZ4H4U$CGH U!F
P$,U)Q?HPJIZ(:>+UF.!"V&202_9TZ;U->%H0+5'W1G?9?I;K_W6S.+7]9F'DI/[V
P^'R@;# H8>KY*PE36PWTG[%S]=)+PYPP6\</%*QWC)1?D5H +$[,GJN#U9[&""\D
PG\ Q90\J#I1^]CSIE,=^JJ5,;;:+*!K-=CAHV+::[Q6SRXJ2#-2E='VH9G\:T/%7
P151]M^<-%UKP&J)5Y-\JN$Y>;2@(5(/('875TGK,$RN#8CLK]'^JK@4)%?-W&BNR
PY%(^3YX7=\[N%\I5J[1B0R%_FW/=6UML*?8]J!VG^GUQIQ^J2%;Y/.CW,+KI60EC
P$T4L/C:;A ] 6MTL22BR9=YQ3NN@LY4O[) 2)[&<"VN'GJR)IZF(.K^C%<<OY<,9
PSN>EW'U@J"!R-ZLBP]L^D6#]8EG\.QC6WP56)@;U'KQ ?\03<(-)'Z$-;/*WV0DO
P;FT.SX8P9RC[KE>I@32G-1VY]7JW+!-F_R42?/G)"*:01RSI5/V]<TY>NA@3O."W
P/223K:K,"2F=D/@;3YRP<-)+M[YJ#\D8DL'B2*_M3$)^Q7W+;EN8Q[O62A%:?\[=
P3[,;C_Z1SYQV3^[!S\A&?#Q8ZM(-!K=$IZXG2Y<[6 [SY(N=-G4AJY<F*BCR-J@]
P+Q%KIJR!M95%U#L#("Z,>*QY:XB3>[[.O"^_U*<7AXNEE;O3_X8TR,HWB0>A+/A]
PFCN)X>4B_JKK-N9L0QZ6@$(_ 9(%04X>IP74H(S<(SY)+.C3X=H/CW.W'3-?<.6D
P3@*&%J'\=@;WU23OJD>!.KFKR$SOWJ^F/]KL.@U1Y22?-Q;*\C"&JLSV]_2?^J72
PT!^HM[K@U]&D"JR;%LVN7:=P3<+[Y_(OC%0FA4RD*]A8XTHM[)'N^X!>[E+6)#J,
P6?::OXYX RFJ/S$!$Z0Q'O(E;$-BM=KT?%DBMI4WK4O"5*V^.6S'CW7,3.F'MW):
P3Z6#3[7FKL5SVEQ/N3/^_$.3*AG$M("U&A/?W]63.#YY%N_CPKR_,E5GULF.;.:S
P)<SG!O_LY\,,,Z,?Q]8^W6QPLKIO&WUCZ]Y>EIPWB[-Y[#'9TVQ) A@?]R\\W\>@
PPF\"@!]/RU;OS&B/.$XX#$X-:'^4BVLQ$I'[LD,,;Q7FWTBY;[\8)&9FE5'"\8C8
P367Z&1S?>:24 ?&_#'G "*M*M[XP#D_7W]$M+#P;:MPZ?T5NV0T*) A)%#<G,H@;
P7";>?\I<Q"AZ?,@:LUC/;@-8CG,VNS][IU8"$E4$J1=@73<B8@B2!HZ=ZWVQ>3ZM
PJRC>30!?7<?=UNIA1YQ_"9?^#H4V))"*AGTP*1K&XQR(MT@.?=GUM*MUU\@DNKH;
P[4I"P39[5ZXCPDM.@9%$G!]+^!GR=(G31)8;UKOXW/7<C4T7.,@QX"J#S08)$T+:
P.TD47GD-9JW;<S\<(X^?9DTF1;Y\3^3>*0'Y#%L?G6<V^!$VQHLE0\U1,PJ(3O@O
PE]8>P.F31/-*%M::8)B2(KP*5 E/U">"OPG#G]\LF72QJ5TDK'>*J^$21H30ZC'[
P41I2G>OFD<ZRKV7%9D5YS>G6Q%@,F_"ZP$T IRLI;;Y:J^<1R2_>6"@6+"9"O"2$
P& L];K.WL?'KB>0#+8MZNT\G_,TI=%B;U)2WW\,C\'J('DEE5K4OV?YI\WRG,T,T
P,>9[SX/1\2CJ%Y5G19IC9-%=3?I?.B-%N&FXG37W>6;XWE1Z=7R47.N;!8Z-LQUS
P!#4A();DU+S;]54]A7E6O7OO@?-!;[/9'D PNG()V_<$+\KK3A-4LH<^D-M_5T44
PHM_IQW@68[WC=_E]+:@'.S&G5  G7R&X:U"C6L=9_^RY\U2=W=;?A_LC%TP"CN E
PD3!(:BWY3KZNT)6<O8A8"\LCIWFHK^8.C6^G]N:YH&)RD'^Q\A]D>TVY<:;OW:*2
PC^;??\MSLD$1]W_+\L!.CA8'.,)&CLCN?81_BGR.5(A9?5(>"U>N+ M_R.UMMQ7M
P_95@-Z2P-.;-]CMB,B$Z.O";@TUCP3JW4<,?;N)M?F1B( U5KM\Q7L-GC;$NLM18
PH;J5.W:3ZI+2FBQOVL"T<A9WN>X;=?,1I\S+><=4>@S*[F;]PYT-85HL2(B],RF+
PBFZ'9D[ BY"620B+$$I7^^CSA#?7,%DV@<G%LQSFQH3G7'!*^Q(W=9^F^">:#@;Z
P2<'/"1#'TO^47FQ#YF(XF6E1\Y*0H)KA/U^V$D-3E]PK2L]V! -7^%CRB<7%V;#K
P'K9-)8C_%_<]9J#SP6;5ILS;C\(H7QHTOAIU?K]%:G_-4ZRAND9&3H$N-1JC+\/Y
PQW'+)(/X0.^^N;[;&SJ5[TJSS==O[4:XKD*4R!&<$BCC"3TY^MG6V!VSSO;Z\JRQ
PTR4$)RS2Q$)J7O]G5H1Z5YWX@$PIN#XK7?0:TXB<-G5D?FW$HG7H$$)ZNR:CD7V-
P2%ZYTSQB?>?5-F@IPK6+>$ '#^9# \E<^2 S1-R+.5ZFVHJ8@9*\_!1T]RV :YX@
PN__6956^!@_$%S@6[[!A'Z?$$D?UGAILFWR97AP/D$JN+-C7%XYV&@Y\AUTA+\FU
P4V/")GS@I3U<0QR3>M&]R@%#>F\<7_E.JLWW%GY5MJXB-[#C,#K,[3\F<YGR+#I>
P"V4O8:)7#WP<:&EYE1JZ>&D;7#/XI0ZB63)F7(_2CKF'UO%R"^\*>#-@KZ1>29%B
P-L*C>THSP5#;=2K#AHDJ<&:EO]@)6Z8R'J(QO8ZHL5]K?4W7?3KN#)\H.67D0H*W
P3U#V^:6I:>B3T7V]L@LQ)UWLJ;2>S:NSAY(>KTT1C CXR$J0UKZIEZF':O-["P0H
P_LX2D:CW1+;R=/C=1FZ8F_O2.]Y'5M"ED48<BAWT&G-XS.=KU\M)UU6-ON7;(4]#
P>[/M[R$EY13\^7"=&^\EH&#YP#]/R2K>$0K+VYWYX)02O2.=K&#<'A-EU!_=DY<@
PHWUFSB<2KY>58VBIO%+\/8ZT.W_M>29SX(E+N$>F5H/C/6Q9(F-" H(;*O]AO24B
P)&&TA)F[,_GPPDI_0?D:JVP1#3 OL +9MY46XWF9P:-L>ADSQM^&=7P_IT1&#$"R
P4QO_5/[RF=BEH3)-3X)\);0VS5:/\0'3%8M[PRXG9WY9(J@)[6;5+"-_+F[7F&P)
P\RY%^&V&-[0F7/?E^ZT -A^B$?-Q&^YU<RL?9SHM,J&:[T71P]<U*R#4FUW@!V(9
P=&.^L[XYWLC!4_-30-$ '35LG#I1G! YI92>^INTS=@L.T%T@0"Q^NEZ!IE_ZTA 
P%"!OZ=K.#0<EG:9U%B:?POO<@X\/[4T3B1JEO[BZ?C%)&Z1;8F,R)1H&P=842ON)
PFXYDZ,3,O \Z8Q=D<1.C80;F45XH<6,R2 E$5AD H<, "B4,'CA: 3&3VX@Z-E,T
P;F].>(,&EW'[IG&NQY=)E47X-2)!\;FCW)@;W<A5W.QL@+79>GO%_P<P-T_UX<R 
P@*(Q'ILLYM"$-=C;=1B5^MJ8HCC33)#^80=#5T=>B%]K_;()2<HVVU"WO()L?:M[
P,B4?:AJHP )PC5G8S*]RT1WJ5W6J+A!OG3/E &GF73 HK8$0(3HM@P?</N((RA+O
P%3K@2U*9%G81MOVM9WIAH6(2OKO'N@T4RR)L3'42#96L_EL1M:L%/'IMT!V<9A3@
P(1/^@ZZ[8NMU#9'IUAM4XJEHUB"Q#HKL=VXU,*[0S^XY*3:EZXL1GKP7*<#/D0ZG
P(]JBH<A$<A6X(1MM#QU,8%V=WF@*C6V2\,):3!*DD/]7-YHO<A=*#8!-M0SCF@AU
P69ALJ)[N)TM:-O!MA27,MH\JN0Z]]MDY4>XRBL@7 2E1ZLK#(D?@(2Q-J8*!)!Z;
PUGIH9=CMM/3-2S#<@&P7>Q1*F('@B:5,J>:LTI.1^&0U.XFA4!62K2[(YYKH^G/Q
P(%<+5;[U&-S/M6EE;[CH^EF(E^ /,#6671]JPT<"ML+4E\:R?*9M&-C5WM^/;#)2
PM?%@05&"(JX\KT"U0GEU/\WMD()]X-O2<@G2'<?N^+RN('[2BG[;DT(+:TVQP3FQ
PXQ-\?7HKV-$.,9[!V</[EXZX8HL.(Y'!GB1OBRR2ES];L= EQ/TKK]=P4-M"6!JB
PYR*AX=&,Q\4C!BAV1('3%KL0T9CD/MTX[RZV2:7\WU@J>WUOPNDT/ADH:!D\8<4>
PG$;0B;5G!>NYOII:<_+RE<R0:I83D'8@4-9JV@H==-=+9YG9BLY)X ,Y'C#A3Q-_
P%K6N<+/"U)(':T6\J(>XV7=R*'?._PJFN_7/L[AO(2WS#/&QDZ32#Z+"U#;(@(4=
PMX/?3,;,Z2^RQ3K8S:2];FA.>W[,D<'9&C,*+O1Y6^?%?*1/O^*TK1?ZSN#_ZT7G
P(3G3ZNE= 6G2A%8H15K?*=9H38M&P(B^KHK1M.>!#A!H+LS^,]WS5!<@6NS3V98W
P']VU4$/YGP4_U+"]4/$D,\3X!$$=Y_?*N(%,R>0MXJ2>8I3'3;RF'3S]Q_4I$$@%
P,( _ER;N1\E$"^AR='I[%MKHS[G>C"S*(\C9VW4.29-:<+=3ZV::K9MC:G )FP,O
P;3#BE8^)Z*:VE.0F7F8MZ)X-]_@G"%0!/I1GW@]L7O#RU@-1,S*;=B67"6?^H-4N
P>/6J07*-G 69+,<4D]G&/D('AD%>VIM,D@6JDOT?7WWG)P6HFV!LA.^M:([*C;-O
P-1Y<+P<LQHZR_T42/&%\2FQNSVP3T6R+0(UFOC #_\1EA\G5=L%R9T20WS#R#F![
P$@8%+_B8%GSSFUGM-3KI1!>*?T!S0RZL5$P8H(CR>@I 2+I!2N16'\9Q%ZSM86<J
PF_9\]5@21ND:(^D_"/4'!6V[CCZE))4S&%Z#O-'\RUJ'L%UYD^0U8$2!I)PV<NY;
P/@2PPOIP)0#%(N(Q9L.HE^24?B%_THRZD7^1D+T;:444GI>[RKR1]\)<+JQKJGI=
PV'I&F.YT=$/DPWVDVJ^/TSTX=.&84<=R*L@GE&_,2U^ I8MC_@SV03A9'T[,@QRT
P25A)4U[C1$OFGR,P6);96SNKQX/P4N_Y&9+92G*F'R<,:#.6W60:X92?C@S2OO"Z
P.AW0EX^_"T?Z.LMXJ(R+"Q/IZNF#JO"%RYH! )F[5E_077,/_,\5LO>G\C]5A0 &
P&B8PS+.GS( :F6=8JZ^J/F5;C.B!*J*&'N6&E: 5=HHV.O@2RQLLA+A[@1#S&S\]
PR%J?\XR\_83]3P,EHCI<FN0#28/E4@0XPN[ZW(U_W!@VTHWM=MKW<1Z^YAM910NB
P=]_+;=*9BU!>('H6,HP,K5##M2%K?.O2(.@L*R=1J/Z =P1?:(*+.QU?L RPF !+
PW"1-</@*S19*G.FOIRDGJ JWI;2>V&OU@,0MI!,<M-VH".D6GXA%)'OQ:RP6[6"\
P EJ]192 &!&*HL>VTC5#89&0H.1B+<RXVNV]8WJ++CP;DK6KJ_$<1DV'\B@^>/OV
PW(4U!^!I6CA-QLY_,'UVJ_VMLZ\JWA5W:DIG@]-$BF16TBWDUO$X(#,*[.>85M6B
PJM*]$NAGHB8Q*)U-VCZ@PN2U<:EBBDFFU#TEI,3UZ&8QA%#>WQ2S/#48J7#(YD44
P+RS%H*@#G73#/L.V3,"TD3T9FT$ @8+)5V&8$IBX@7C3WSX?,;6U]V>]0V9%JL@T
PCWJP$)TUKKS]+LBJU"K&,:P(BWWT:GCEK'HB,X4A9;&<1V VV!A2MHEFK!^W5Y_%
P\\5EG$KE\P18;7[)1QFLSQWEJ$;!,1:< J:D>1_<)=.K$$29J*C7H%B6D_G5&B8*
P_VO"R9U'W1DXQLXJSB9#M#>B118;KP%BL*LHM3;9W<_QXKH<GA$?6,+'M>*GUO_5
P1BH7/]Y% (=17U$0<RQ]4_YK$^L.+"N%#N>"% SW%\5B\@0\& F^&:D[-8[F+_ZQ
PP^56H&GR<64TR^!E#*BEKN:;$Q;&G]>A*YLU,;&,RG4R;P\6* )A>N9Z@C:S<3Q,
P% + ZRX\6(J^6&<+; \&9E>,4ZP95 :BASC0#1%\2>%NQ'^:Y_QT>-@(<7'B"OKO
P=L(IM<<=7M4,*+PM P978U\QUYMP!TN ?43"(#&783S'4('FM"UH(IVT=K>F!U*P
P3F1']SKKG5%OKXD'IR%8(>R/% )3$)LF PFY-</]A7,;:N9@%Q]),?EM3[.,).=8
P[Q@\JNO,A9DA6[<W?[O0&!-6W2ZYFXB^=WR^QGRE*6($G#0JLCX3A3OOB0[3&_H;
PM$AZF6G NRCZ%].C>.Q)GIZ%IQ4$Z$9R+*5EG'CG;H ZA&07+SG?3 %-B8U:_IQ[
PY-VA^SJN[KBQ+B.S?>_U@"$9KK=1>_.4CLO3XJA4DK>#/1Z(Y2'YF)_[S+5*(X'\
P=CZ)@=1_*0[Y8P3W>)J:UBATJO@AEA!,O9D.\>O[UYG\9"EQ]J+AY\J6:7F3C(@7
P &YRCPYW_)W;116+(E+;ZKRA# D3J^]<K#K41,<33NSV2\BGA=!$5(4JMM=_<\ZG
P0G2;TG^%U)JEGB7Z)1\X&77F" I]B=1U7R_U_!0TL3ZJ,LYK[$[J3UUMI9L_$4GY
PE'%+%C.880!E/3_?YQ >&8DU:#@X)POBG!J0HXQ(;+A]2(\\J&Q[I45(*'SMGR"!
PP5KA[P0(5=F?4&8+@,A%=42E?'LV3;1HG>U]O3IPOS^2[J)/>Z+THJ]RJ<:)/N#P
P >4;4<7V-1:1YNQA'41?;P[Y@"8\*."8 4:5E,<(^NMO.Z:N\+4K\L1>(KA,ND.2
P8AY@</Z&_F[I?V7(&JDH,C!Q,RF\HLYS^TQ':D?FUVY$.8")*)6(!D,)9NW>B(LT
P,G7&0QA&SJM\LF\P3B2,X'!H^KX*TAGH*", DM8Z#A.[4H#ET=/3:/"(RF-%>!^*
P8'Z96\]ZJ]_+APTQV7T_:GZ\%5J0R1JP0[L<B%\67H7]U3K2\H7O,*C4AKLT!D$/
POMQUT>FW(5%!)JJXS%L XL^XL"L82(DU,XV%QB2OFM0%'_*.1=PG&IK%NBV5X$JD
P8AN+#8!1CL(Y4V*CZ?_FM#BU/?00)EPYLEND4LHQ+0I,I#AAVVWT.!^#GW_[98LA
P/(8\S#'Y53!*+OE8H@Z!70*0^/U8!7(!&+<+#$'4P>?C#!)8$",#P'2*]!*["BKP
P;/):QP0YP&J7=N"QEF.K4&F(Q?@T[)C%:ROA,B9!F!.$1/QJ$99(K6#BH&M.82P-
P=)H@%D2SO6EAP>/LB&?5<\]@F3NVK/Z]9WP/XRF$;;<9TH8[ZMBP#388>?L\J:7Q
PS7Q(L-:RTWL#/4K@!6@/P(0C4DTL&0)\PL??=D.,C UG.-]VNW"O3V3V]_#E/S5B
P%B[]UYSKOTNVEP]Y217]PU\R83I$(.WV77\*J[003@M=WQG84WM3-'!PZ@@\MZJK
P4DCE ]"NVH=C*&0*LJH+,BZ2609L\PM7U'Q*9Y>I4,.%:.?M<X\'A?@C@+40&+QW
PFQ]6(6H\RMIGFIHZ:$<1,9O), +2X9,4,/"\QI2$$X7UJ_?I5@2NS)HHN4.7-_:8
P?MOTXKJZY2^:-#%HF@H_[\PI!S8)0Y'5!^$0P@<24?E^^D AJWT0?,+K;$020%:T
P21C*V$I', +*01C@ATR8\9A?E!?:Z KJL(U8;+W!?/)^3OFG/Z2*7CE]80$'ZBP<
P4+#N\C< "32(8Y5E7;XW4_67;-B) C@9A/<8>)<4C1! -[R!57ISN8GU-I+F6$!6
PFDCL#T>)S./?LN+0*,I%^$_P(=%ZM17.@.X=B27?&#(9P&-'%;O$A\NSWSEL,K'L
P&:8?_8E:M#F\NNF7F>E9@:X(M<1ZSQ7+"1*!$+AY_ 3*KSDI&U7W=_#,BRIY;"W\
PAPR*7IO;>[[J$[:QX,\XKD:#N;L!3'W%#?+,N7 ^7B7.B43 OE]MU=# 7U4=[*$U
P@S#%</"XP38%:9;E7,V3PH9O7*LC8 HKWL'E4OE5<D**[EY*-@<5)<PA2WXH4.I+
PKIO.QO,=Z (L50'P3YW4=@[DF2#H?%S:]!=3Z;$ ?.KFUG ;8A=.A8+,W8A?S%D)
PO]\<8 UDV/EZE%G A=BK!T@A$+4[%?''V0'@]CG[<M<G >GY3\'TXZ>:)'F9T^4T
PIT:H\E["@H]LEF2(J.7Q-!+CSA[NH5P)B1BW."]RL;(P,PY(Z.P58B@JUI[=WN $
P.&"Q3.OF4:Y<4=%B<XSZ=(3,L6MDX6^0(PRM//+]S/5#!*9IZ,$3>2:/W$;(3J--
PYAA=P3Z23-*0^9,Q#/8'M)?KX[>E,UOAGU].&%!%T!R9]H2,:F7_P9Z\VW$C4<GX
P/<_:0_RE5_>$\JT:+2;'I=0#C5ZX7TEZPT]!:R$^5;_!J!,E1T1/.J'PL:57B'F,
PM< 7L?WAEK/L3#Y48R1_(18C%G['':NH<>LO%,W07')WS*@W3[$2J4]8ZLJ24V+U
P3LB<M:Z:(UW4PMWMGE/@7 ;C>4\@WC&V<+2O<8!;;Z*V9=G:C07#<QZG4DL&&VKJ
P9&NN6K>3C8;Y/[$78!>],UZWM\N-&@WUKHLY7V>Z)L16(:Z03UO@<V4/XGT$7N#]
PGX4HH$)\>DC.L78@B B<A6@9*)9A6V&%;%%M3IC0>R:ZWW?RO(>*.&?I D:M&[-"
P150OP4(-\HA:+NUI5L,W6]9ZNU-MR4M#7?%)=MEO<I?O74SK+O4^A'CRW,C;5HR@
P1]DB)<GEVT2NJS5)A)T;,I P"L+Q;:V2QI)GTUTL0("2U$M2$ A8>1IETXZW"!NZ
PP#^,"3)-"CJS86P&B:ZZ P@DRG'<%\O+,-^KZ5+T;R=\ N]'2_C)*U8CW"TVDP:G
PPEHC6W@-6G1."AH^Z3*_TG=C)4"]_Z94\->Z-XFFV1-9 4<F[R)6BP+OWEPXO(BH
PO/;7H,X / (>7K42+R)ME'5T"DI>2'3?>&-KQ FB@.PYV&5=49Q,-D A'+) B)^B
PC)*MJ5;U\!R1_AA1*)R%XAYI=@(/65H\=B?(FD9HK;VZF_WEV!!J6R-7FI;/?(#.
PY<B MG2AGS4+^)*XJ)*GDTHQ^L#W5.2YA;#7.QI+1GY^7NOGM)=,L T1D+G ,_TY
PN*0W@LZ@HP=M\)9S5;UJ.5)"VJ'?GU=%IMD>B))\=_G128 !UMP/&#T"5,U'TR?W
PZT#W/ZZ=97/IMSZS71L-[[((^Q0<Y7!0[?P=+W_7N7GF!J?^!'&0689G.@/T^)'9
P>1]';-X+:B?I_?GTYQK$[-;\=5)0Q^>V-Q6K^ "QD5O($V=HP#R4OD, TLPHSWWK
P![RT$X-$ *?UJ11QT-BFP\;_6'3Q]4 &*37HXE(;*H&L#>:#BGKC&OM0S%=?YYB.
P1)7'[)*;?Y6GRD=EHSOGD9,4XU01/(Y<!-[3ZRT*5(E_BQK%F&I6I*S%]6"E$+J[
PQKM+V\T6?6NP'B;.W640@,D\LO S:09\)LGV5FMXQG<]X_[DL7ZIR0(4L+^#\+5B
P%_^UJQ'TQ18 0AXX1-12D'(B.T4TPFCJD$QP[/:0-V/^2.2I36X=HESQ>[1V0-,M
P;,\ER#+Z\)UI#/2=UOII&MTLI"X."YH]@H.DD"<^""RZ%1P$N+=#L=!5IWRQ.\\1
PROD:'"Z5O[!B!9T XG-O,RX<=PH0S+G06H4HG7!6W7V)46><=\Q_^4ZPR%;])6SD
P<:36/=<?L%3;'$%)/J)Y_L%L$EGGL$(^UP\B>"JA5CE,-W"D&I(6_^>$BKPP6"!F
P)DUW"R69SDBL,XDN._@G'"GD$1R]FG4#><9.UA%*"J>LC#N!)H2/=\2BQ B;$-6 
PFM9@G_]\L]VY*$A1D,/MKZV]MAE4L!9B)TDP0V\>^_]%RKEWKH+#;E0:TBNR\&M&
POT.T"VT.T]:%ZQE%(\W\LDZQBD<6G_6=H,ZA0) HR;A_-I<1+VAHY*# .!^BVW\E
PCH3$);>3,<X]0/N!>\88:\>M?4J_D2S83I'O#-O<<IO7,L::NUE2I! ?9TL=&0,<
P$ML\ %XE6'3@F^-_(%BH\::SVB"Z0_C-C$?R^+O":H?,#DKO6XI>MA[=6X?/[W]A
P:RK)1+4MXR!8C1+&@L9!+(=1LD_/Q'5L+$,)16]P3MXVM;6D<7C6'E0'-[*L,1HO
P]\2GN)QY>)BKS?1G:X[2G1DJ'IABB"6CPCK62,N]8-U>,4%6V5>:B<KVI $:&9 N
P"<>-HJ' 2%-(Z;UM%PZF;.Q!;VSU:BKZN4E5+3:0AN(EN:])U9*V*0 ;I&4XU:.]
PWQNEI-4_)HKJ&]QFT[IJ2"*.F]1D8KRQ03./)<:L/[7CO!VKX$,E.XZ'(SAKH-@B
PWI_%3\P->B,[IKP,LQX$[($H;*G\:"SMXE STDP8JE7_:FR/Z4L=L)\OE;2-T[!W
P1F;[(1.=CX9+#=#^O=,GMV?T1.W3(*7N>2W1J/+'_(5.OSO=Z8]"Q"*H>N80Q2>U
P*RZLX/"O6@)*68J_G2%LSQY4:-X[Q/%@)G>395^4?Z"Z!4J)#V(:@-^J:J\-+"XB
P=R*9.KZ7)D;T*\-*NJFS'>3=_\2U8:M:A"-YX/OY[X?U[IES-KP'U^G52,\+[ J/
PE+/$+UY98MJP4@Y:8MH@BUSNZ""+MWW3M/.F$CHYPLD.PR@%*>)-"Z&@Q7JBO %_
P5+#$]"I+#^A.XQ-9"]S)RU'IX[]G>FSAPS'S7AJ7_$T1HY)$_V&*0_'L QQJ^;O+
P2N*-."P:0%KBG'&29ZF)K&7!D-'M;QKYJY7\;!]8;J+%(%:,D[IP3U.XW4>SB3UW
PYD1Y9GA2FT4NTN-V6=Y[:72X%&R45C: ?+,R@N>_'MT=)$S[H.)].&<CAE:AKD!;
P$U;=NSG-3RJ8'M^;(5PT<U>[QW)O-Z+&ESAQ\T^PV*FJ')Q:*3R^C%*"ID1?:TD@
PKU=KO)H_D:O^@LJAFQ/<>^^XF])+3UF5P1 6%GA*LL2 Y63S%O/K",M:O+.(/RD^
P:"T![TX;C*92^5RVI9Y:& "F,6BGM:OUMX3\FV8'TB."])!QL$#QC,7"=6K\129_
P^VV.T WP(5^#VL:PJ&UKR_DJ90P<+_\1U63AN?1J5$#8'[?NB ,N."2H,W)K2C(C
PKLZS)3L^:LN]H<WH>RI!P2@9JYM6W?!SE]%["H2X4F<'JJG<-)J0>.]QJ+'>$&9?
P7KV6]E7G35R\=N!+ K;N4*X1?XQ_F#O1)&$]\(9W?$I.,T:"I+$?S6$/T8^6";R\
P>KX"MB%VVIL!$'C'8?&J?:GC8NG/,&BW.0(!S%/%J/K@8+2+I'V[#E3GAJ&R;MV,
P_WO>#!AEBEELQ&#T+E@PY35WF&H,8Y/P.+24?_KN?:\B:D'G@B;OR.Q-%'1 ]#2=
P_]XCON@[#/M\) <.4.S YG)KF2Q4F?FF_&'I5Z;#1Z:7?8'-W?Q#@S:^V5*!=MVX
PE9D-EWA((;ZT166UHJ[=\ I:\&7DO6#1=$JT"<7+;I\]8426:ITC_.A[/_,#3&&!
P^+$]/>QC63^Z3ES5(E23&;T!VH" L-\>9MA" N>;U7*UL,7BYZWS1F)UK3Z+ /,-
PAT>=HQ(U&VI*J/[V+%<^Z;+MJIKNG@\KH;8Q2\<@MK$@M9"4QXF\5=(S,M?+T5^B
P=?5P=71+ANOATHGN.5W'U<[7TS/^^AS"#3TO,GB9:[H"1 V:7^$G_7L5A)SD5DQ:
P\RXYI+480-'25>QBL>IVXZJ]\G_3(:+K)=^W:A<BY1M!=GV)8\B##$B)9(+=XOA"
PZ3-MD3O Z+3C3F=&SV;&+ D,:,KJ!,X9LO-P?KE_.<K=A.A"HG"H\TT/?HKX&(DQ
PGL-L,)W6@<FX/"_\P"'-$FRQPC2Z=1 TLTN5P"[!.]36^..+J(A*=9NI7<F $T5[
PD^\]3VI &2+VV.'N 8T"]LC%-"E>%;I8?WD&;$_=G8!)ETIP&'=;=MB^W[XS_);_
P2DJ>^IX*5"SP%*^5WQBN'!]YQ5F*7,9+4B<S>FT^^V[! ^K KG*XJ?HJU ,J=5N;
PDYC=NP]HQF6J=OQ1=NL;.\_T-9FU(%VVD0/>)@!D6I;X+^N%N& +:-K@DR. <6F)
PMFW9:4@N^L2)4C^ ,6&733NTB8:Y[TH?\O!'W%=VO#H_:-F );4(_'V )[.0AW_9
P)R E058\@3/.@UR,<9/4@+OB?P%_4A=/JR##N>L@.","?E+F3:=92"ZX_/%J4W&L
PU8''M&"XQ!SG^8H-DX])U0,C^0OI:RH*\,ZJNDD:&G[@AZ=3A29TX&LW?>9'X+8<
P5^VLR[5 D&^%>IPM*GT:%6>R"5<V!?BR-'&W @C6;17=IM\R\5V';1F.MM4:/U!B
P#])65HOH)@+;[,RW[2_!A.0IE+5H9YAD+I7WDM'PZ]RQE7WM:4P6^GE(T3X4?\D?
P\.]O:U T9PJ6HJD1/H[,LX0O4\9*HL6-U;Y,D<@N"Y".4GI.]MU%B)0UB6WU!^4$
P 5];!YRB:^8R^P@3BR\S,F7@,+,5DH5"-M[TB)I.\1=FP_FKO[40DB'%KPS_]U[4
PC9Z ]ZNP*H_?.#.H+LW^\D=NR"<6B%A^DC<4F]QUE7GS7^[. $<^U#MV_I7G,7QS
P9PN6X'-,W[4EF]*>.RUN)'BOP1/0[O\/=2.,9G"8WT64]=?A@"9^'<+52G@9/YV;
PD8C#-$L1W%U7Z6F34\E:"&Q/KR74_0SS^=IBE&$D$'JE%[KQ0QK<=A606H[')PI9
PU\Z.?!M0'R_#@NJ+7<I:*R6OL,/$I2,HFO]T5*L=_"9_K<,XNQ#75P",;==B_[G#
PBD]8[WLL]$E]IGIE][_U<4[4Y&ZHY<):YXM=O)1@P;.6E)1#M!MUG.]D .3L[%4"
P.ZC-G1/BOSD=IH1DN8>OK%8!)N;P9;=DT.L"+/G8'?V;K[BOG:$DOV3ZBR+.6+ML
P/M5,3;GW 'L+\>^I%Q:.II?(P>].J&-U#=D!J[3FEF@+%,D,;3CQ@5T4^[7_]=*J
PG2[AH6NT\D*E$I.3D7Q5N?5G0_[I=^)+4_#T:#.JGECE%380JAR:WM4P8PJ&$F:J
PD>M+E2& 3JPDXFM32U"Y%F;C?)"]%/0327C RD^KX5U=<B .=A#(3NR"(UNJXC%S
P%V5M<N+.4&BB?)WO2=LSF:[C6N@KTOQN#]H+?LSJP M0:SX.S EG,:7XF>(3X6CT
PUYN4Z,'+-LY'W\',V*5S6B@11>U6[;Q(UAE#U3\"TF%:Y6H39SD5M=E!D93'?</(
PQ%)2+7@B5@ 8TE)9N#6TP"^]"R,;GSX-^!PBZ-UW>W?W-L6)FY#2DA:=BT,-F4P:
PL[#/=/PD/YB0!N.W4S /U:G6;>;J.X2'PM<+KB9R7&,G"Y8.PA3-S?OEE$-=HML(
PQZ6.UGJ)"',$M^_ZANS5;] :[FTJ&@JMY5!1!N"-)_"*5K''VULU"%-9!)^VA?5"
P XYU?NJ#HYCEEX]OXX7!ABZ]ORMZ;IM("CR]#5"UL-@987NTF]*;$-8D*9!W(FNV
PK189:3AN+0YM,/%[[-55OND'@Y9Y6;5K@;Q/C4#3JQ0Y#:!?MTW7U%!RP82U356(
P#$ )(9>/HFT 2G1W2#=Y4P&YJGTNW3$#\%3YC]\AAVHATQF^-.P&<$K9%!89F%P>
P()K\-&""(=H%3JI6QAE_>H:..MEYLO9WN_&/C,:QOSPIC=!'1YZ4+P:]G/:VI8,"
PXI<W.V]JRFCL0#JBI3H9O=BB'_7/;<AZD[EJ@V>V%;.LY$/&T.-ZK& L'KL<0WIB
PY4_?Y1Q$>WG:)/T:^,(>Y"JA]-O ?N.'GA9U$)/&T<B_S8HJ/E5/@2#AR( >'*2?
PS J09</./(X7U^0;EGPZ<5(9<CN?&<VPC9/1@(GW?1D-4Q\U-)KD>\H0^@TD+*>6
PE)#6H:\NP<!,4X^OG,J&B-H.MPYL@'B1AU%W7Z;MIVQ_SN%MN@99914D,WY1%QS 
PIQ0>\!1F&>@T7=#HT][W-C65% ,(]BY?^14:"Z3:IMCMN0,^(7]K4XSVU!W5 _&I
PL%S5$K+.;208X.B$?1C/,)X&.8C[2]5U#MY7_:# 5%"PE<XK;G873\A+&71']6V4
P+?45H*0S"2X2$4!@!VXLS,#)X:G1M]C+3&17.!2TG(YGKJ5W\!:5MRD268D+^M)8
P<:E<M%0 .3OH_Q*RX/GX&?![?[5R5D<[[_C(%=)%SDZ<W<Q[]C:#\6W1C7FP!SVY
P!-D@N>&3$,A.A:28.$$O')$%>]$1\(2?KP7V(,#E:/A1[RR^5'C_9G*EV#''[RX#
PXE8L2YHR1JZ+:=Q+[PX??XDWX**2,XN/,+[L0E5H%J*$+#)[8OF_O)@]5CUOEZ_=
P,,VR)2+W9FXY) >8N!('J^ON\M=\H'M%J-94/7W;P"5R=;J %,.D2ET<KK@^BH9&
P8<8S/%2=(*ZQS@L9M_7SFK."Q&QHLE%[3>_H!E#30P%LK>FC]Z&)IG^\L5<0 :E6
P(?R3I'#Q>639?0G;S";24\+_MH*!6IZ$P<C.]AF7<BA=VLNO0X_UNKO1@^+.^GLH
P6[ABM/08,JBP0@NR>BM(:!H9,-D%[,0' ,Y3\8PY$X.1;\LO$,7C'L'&J<DN^CJ^
P62AM.P8W%];<B_6:>BH"K5 ]<+/#.'K\LCV[5%7SX*9<XY$:-(,>)KIV2M&]AW7X
P8GLM4=(Q3&E*OFLC&V5<'V5M^-6:K40U;AV ;*' Z6PS&'%9_OJY-\,F[!&XPT$)
P4#"0)+6H] "\G7H]X:[\D2KA/#^$.0&Y']3U+'*OTXBW93EV]^-85LH-WM"3O-UM
PQ;#X,(/]'5A$CL2]%F"MN(K6.J=S&)&\1X_F6BY ]'NIRFP@U&!)!3X<TPL9W9M&
P=I*Q7DGF8(2-7(,[0]T#J'\/P*6X'4V^>@U&=.8]5@V=FI,*_I>B0U"U_7LF3KKX
PHD@6E--%_QC#W%S12[P*IV.=>9NU.=E&IP2U@UQN;20XD^U0'F"!J=.\23Q][I44
P^;[=+1)*+<Y#.IV]Q%,!<"R@/VW&\B3(GU'B.W.JXKZX)A::<)A@9II>$>=DTFY)
PD#XR*].4%/]0&-_V :K2L^C39$Y@B0N<<'7H.VEAS_M*60=06MHE;\"6'L=RV?)M
PG ^!^==0!@4"HKG'RCM-]4?O&_>YXK:I%@=BS^2IG8H<)LD@[@$?2YPH%@3I$$8^
PA;DJII^,W[),TPM='GJY>AMBTG'(ZPL&Q09<6OE&;KM"VD-K,<#=C)6UK\]1$8+A
PX51U?NM"M;VJYH%1X#IHTRU<CO\7TV_7_9A!"!+1 MA*&]ZKH#KIV'17X<N5'6XA
P\T4DTPH\H] B$O)U(_5;5\G,]_, 45Z<L5TFVPFK^8<$C XC"K)Y[N9;D$19I'-:
P3)\$T &RNZ[O>$@&J^C\,5'M),4<A@-!8K:-"= LE?G-9$'M:<.5(LH!E@OWJCHW
PER5YU,/T2G)'_*[I(OGXW&%8V9%=O5LJUIYS@/]P%PZ)N1431H3;;V:!_7J&,K1]
P!,;[AU:L4)W$?6AJ=+2DUSG8TT *E/<'P?R)]\R$G1]073WN 9G)3?TW@=HTYM6E
PSN&2Q0XM]7YH!MEUSQ48I+:II2(E?4[ESI27@SQ2P^)\]<(<KJ01LTYG)U^A:H78
P=-K?QX/4G:)(3G<NAQ/:;>),E:3Y5EZFL*KZ,.H)[]H)<&SY&ULCA\WP*7Q EW8O
PS?N7:]H*Y-[')5?\V.]#JH9H*,,QQ7 ::K)NP"HRU?UL._&60BE">TH6;:YF6Z<L
PK"I"P J1W+;O:%/-A&<<!Z"0G"T)6DK?*7?UXPS&$&C4M/ [8"&A71&*U@GQ07?[
P[,\J&,5&MB%26Z+1"I\OA;>OZDI'+JS,5,P,Q/M39N#Q$/-T4]BX!Y *@?#QI^D?
PX2EO;NR!XLX"QO'4)PYRYE8_GJ^;K"UI9%+DT#E6UML\]ZO<>$*Q+4AJ,?GJ"UUH
P-+U< LS-P88-.:)[$W_!SA,YE&ZO_8CA?K;L#=X-*A[!"O2;OY!ER/FMR<V#WEWJ
PW*VXL@!J>%?10&=;[_QR(^[%A+!)6&IT'OP&-0Z%8N]$N\YX.YP>L#WM_36M)=FJ
P2T-LJ&_WK"TH'$W8#2\ZM\JRC'C1D[%,5K EZSH:(8OA-EBD+:1RG>C]M9U #T'*
PZ8YWR.J-"YU^LNW1+B*5O,4UK"8M'W;,H3H%C6_J/U+3OS9CVB'6GA1GR!L+2Q5>
P%^9W4V4Y+H*@,E3=6SO.,36ZUC^&"0[\!#.9R\?VVMT05/^.<@O^ '-ZW)LCQ]IX
P;S)4*\P=:X_!@3R57P48?K,_-=4/SI.%L2L$O+LDU?H<RW'.P28^.>&WO]FU0A$L
P)ROUZ)D4J:'M\"=HP-49KN^Q#.\:']/1OKVZ<G6B"6:0C&A++-F@,VMG;1ATWIV@
PX+D1J6HG<6*3![6+R?9+2BFNR+AK2@#OG6;4\\H"()*5F7$LF'OA4]6</M>XCUKX
P?;YGRE(;R[__H=^,ESPKW1/P8!C457?5?[%]C1OL5_#(44[8=&V**Q_-Z+0=KOWL
P#9B\ETCJ6[2)]:&/=62I$/RZ9%UZ&]0'IY#@CRZ]01F=+MK$/1,>YG$55Z73DF\5
PU+5P4%3676KWC:HM,C*["U#@ H"[B/<#'N&#\^NR4""0&),TR?N*N1>;]M"1ZK<+
PMF>ZSJ:'-BB=DGY$Y!OH 82@YR5_4R^@+Z1VW7'T 2]:(&17Z(T0 @B'.4ASS_]0
PA^2'@,L]R( I2B_*/CY/]I>BZN:BE%3SXM]:$T&-FM_[;J1BV!NS*QNGOHB>#)LA
PJ%]Z<"N^O_*)P2_4'F*J!L&M.8X@6O:+0<1\F R1M'O/4;M8(]6N@"KY437GSLGV
PC'!)N86#""I[TD/)K495_.L@K?WG7$4X[BGJ-."<\O>:%;A4OTD1@BWRM%(1E9(^
P&""\-%^\T=)X[X$5_/A-$UI\;<>\!AD]DM48V'S6;9(D3)]2.[;R>1([AN]:1DN(
PES97C*4(Y1@]'D_&HHC0"%VC<^*\/@(O3"4J-^$S#AE'JD ]58+,;A@S5L;T&6^.
P(]7> @';0#B-9!FCMW/>K4"V:]\AWQ?G_Z(JL9,K%I(04Z_M)Y\O\BI+MIW<#DUZ
P27%R<6Z4I=&!Q5!A;>;!^)ONRGAX09):XC4\);Q[G!8/!KB%X[/74 \4T"U4T*;"
P(7[HE<#S)XLM8G\?8,A==?1B>'Z_5EE_RC>,8*_6"^;R1P*6SKS,"C3&9-_8XQ2A
P!VKA1^[7P30EO< O_.K\^N:Q,%<4MM-7>A.O632N!SE@',^H?U$KU%HR8^"@QNN4
PXW-R^<?>DVO]8E& 8=QWC0KWF[PHBF3YYF9+LH&36UQOMO@P;XT4Z(1P9+R7-%_N
PO;Z+M,!EB<5,YT!\7\]D?E=2L-L_HRZ5A781QV(..#F7L=?3=87C+JS)PB?.D="]
P:.+#=G=+0I-I/NK4)V7RY"BV, MJ(GR5!0()3WY^GSC#*:Q]GTD?D,0N3T43SG<K
P:N)=?+!N_=VJ%:LGUMXKL HK-?<F;FWOK$P)?0NE5)'*R\DH@/-2**[6[75$PZO@
P<'%R]\578,G:31V[_KR(*8333)2[]F+@=,UDPGBGZ(_C*2\1(1KYD2AD+MY":?"?
PV(D\^*V^3O='_-P1KR8(B^!/H$K$R@S1!!\>J,U;$7Q&Y&9CDD3,]"Y)./D%+.<'
P262(Z.\B68-L(=RX_K/YQ*MSZ4BF.7>CO" 6G@GS'L.S.W*HQ[S:3V(6+XR-1B[$
PL]_*_Z_K/_3_U4/SXT=1(9W#CQH)(G+EJB.[G8;+98X<V3:([C.YW,I7+? 8A#%^
PKVB+:PHUD POG#4V-F&"CDG>B7YK!$UMVF6Q""L6+W+CH'K\<-0@J?!V"++N%T_;
P/OAY MQV;'L4']CMC@]KT@SK38-RT!Q.A()Z=><:6C2\5W2/Y**W\]S7\F[[8L:Q
PQ9.?[EW#;"C%6[$278@G7AU?CA5(&'OI[=69_NYU*%C]R@S]NGA+PS/)0[2\N\_,
P>TUSLO==40HQCZ67F);(:[M2 16]$.\QR7 N$%<\;V-*!3/+6B,@1 82'NWCY"_$
PT; )HXSD#S!R^AE 105P/,+^TD!N7D"<!;P$ZWD/M(G?4[-"+]4-X?$2/?5_O/$*
P]UC?ZJY"<FSL*,M.N#/X5)B!YH(+%&8H!)@>*NT32I;-14C7O:O1/\O(]M@#2[F6
P(Q'?OCV&(OF;]8Y:K*X7EQ#J]&9IFMWJ#O-7Z2SAE("+?Y^ QU!+WB-%V] &%:=G
P;KB>S=O-+]VGKBY IP=DDHBEVZXMF(#RYR6M'68JM%/45D\+F914WQIKWW=XI6?&
P]?\3QY!@42/;T,ISJ\\2!4;N+/FP=(Y+!JB\R<7;8@6_>$/[*M/$68N-11&R-"D,
PI!/;DQAH;K,YN\!HQS(@'P/1^P?7'N2$OG Y#\++UQ=Z"ZCU#^8=>1T,#1"ZIZZ[
P&1=;9CM#7D.2Y36IV3=_A?<]#'R1.Y_EU6T N);6*HYN=CYFT&V(*C ?; +N@\D.
P._>?/;KQE_/AL65D4UER3??L.V'H30_.HM0MN9A*-0)'?])X ?>UN@D6Q>+&+DSF
P4F@;CFUN&P>H=UQ2H+G^V\J*(D>?B77,C%\#.(6JVF5*;I].&%@ADES$I$;_M*]8
P3-+Q*=>!CX#DY[S:0L,7])'O06DJHV\SQOWE3C560/4*=0QF4E5,HO:$*3"D4 L@
PQGU\?@^Q>E%=.!R72C8=-M#^.1=P M=3$R/IM*V?AQ!1L(ZO$MQ9=8:,C_JS$"NX
P^(ICF4\%#?OE'\LZL$4N(*!R>W="@'6B#$Y.D#![9S.?8*,&7)XY:8M2B#ZU""X@
PRTT7G<U*41XZ8-J<^X1LZL:V?KQ$<[DA-]*/27ZN<4#H4Y6"-?-HN;O'6IV\B:)?
PS#:DXD#D,]!V<B/Z/UVBR89C1X0WG1F5;'Z;*9W^/M,![6YTT3%.\2:S5KUT$7']
P;Z<9GKXKSVS'?I^=W#08BUA-EJH=+.4VF0I?3RKM]Y;&4 0?Z5=?'TW88(<0EH.6
P.-&+E--\/\#%/0Z%<]?.<JGM[VDL^70LDJ/@DL'F'N4S#0HR#7%IR;<4%Y-V8V7?
P$^+@+!#8IK8&\2^JK4BE07E%_6K?#.51 \1Y6Z^<&A'JLMM^/V7SPQG2D<>LJ'=4
P$E_)H!MG/.=>/USJ4')@X2:^O+ F)Y6GA!UB>DIN5(U4HJ8D-LXF-]9V /I@.838
P?7?HIV+$GW@J%O]^5.T)SRR?5KZ=BF?- T:IM2B>3JBL)LCFH#T?LEXQTZEG(5BL
P]-_GSXZ%%8B%G228>PRWN8]1;@NY,:;MB*J<J'2]!*QP!=9AEZ<YW*]? 0,1(\/:
P3FT$,.3EFG"#(?+E"V*N>$GK#S-6"DMP!=M2],*7YO<VL,P%WA?8QF,R5AV[*M4O
P%GN8[V?9W=LWTC_^2#_J.71Q)[\-O&,E!:KTC%NT&M6QBO $K:Y(1F+4>OXB_Z;P
PU"$)>U?K=I2Y<]YB21'T,M5W\]).ZN,0GWMO2CWULAV:S%:JOW,ZG+$5@>QA<Z?6
PE><MTPU.B?X&4<VL@'ZE+!4*H>C_?A5?JJ!2%1[$KPW'F\TXON9YV=P[^E(K_JX)
P3] :L^H.3C89'A!."#ZBCP8.3/FWB44G!-D5])FL_+:Q3\(1 F1$"+2RO\V?J[VT
P^LNDJAL^[,U&%+?Z%FBRYS&[N"Y(XY+S$N6[/4C=H$?$(; =WBXA?N>36'U!H:S6
PA-A  N4 #3ZX?R0!J%C<^!EWX>/U8_%$8OK9*3=4;"$"0HK%QM3J"H:XQ?+1BN'<
P1FA,,Y<ND7TC+3(NK;2%0XME(TO"63#ZX%^P7A7\?<SI6]4O..EG3'@E+3-/+F*>
P% E0^I9ZMY=J>^P%%$%!H&M(IDP#LR)QN2CBR8OP"J]N"2T0$^#JIK9?/N(<P:Y(
PP]RX%2'3F%#=ASE7PH1?Q&M6Q7)P.PQ-[8X&B'1#)TO+.?%67^>#)'J>[_VJ%QM8
P_XABOD29]27!'J]E2/5U"KU$3E;PR+(6#(F7ST,5<C).7C!N:LZ#0(&]#135S_',
PKFEOF6L$W"/5+M@4;/%Y9TXB"C?:+&="]27]*2KCU.^>;R,\P$!O 8UTP@;$;Y#0
P_D$')GR(V:LNM10634C/3%S?DO[[B78M8C-@L_K-X/O0D5TY%07,R3[M\. #.@%<
P_/6DK*=,9GK(_Y]O;3_.O4B6U)!NIDP(\J8D?#90KWZ)JULL)*O/Z6@0#\!K45AF
P1KKH6O!JV!>E(AA$.ZHL='6/NQ3+;OD93&L-8C?L2^#%TCN))J4&#;(IES2"-/*?
P+L'\L4WV]Y%AN)DF?I[<W$;B7"78!NG%@,R+1I<"]:3"B,F\\CZ$B^44I+80LGE-
P$@\.;!%5L)A-KA)H-:#&- 2;QQG0_68XY4D@<FZ7*\:W3,/F!FW%#.!B7;WS<Q#@
PHVUTMJ,[*((<\P#Y+?B+ST!=MLC_O4L:,:G"B@YRIULJ0?\;8@MN^"IRPSGVFHK'
P:+EI+203U+B8[N:%,!YU#N*[.+_*$B]B935O5.68'-E<"0YHX727QT%,5-$,AXCV
PIAX&C>#W&KSG /CO6TJ[DG/ L8-@@]DN)H'+:7M1@X^:FD:6!9+J"'2:YX#5<3K'
PZ!;:0R':MAV:^A&7[";X#GX=R4J&?%IZ/[GPS3E?YGPI0<!5@3G[GAUTKN>J^VY1
PU.^C4= '&/S<)B'*:39G!BA5^\^D+V4JUP//K(BW,7RHLFSF['VO-F9".4"9I2>6
P*\;!T*-6Y#^8=4:),0)QS8<7B7J=)U4*P05S?C\(.XGY%K=KW'Y:@+11<_AG%!:^
PK'S707B-^J<,HFG/YU.T-/!HF7AV<[0*?6)V9X*>A0M)$]OT<+)F4+.S4+; NPI9
P#,XZ)!=E87;$U-JH60.H57],?+F$C^!B8[>^/_I0\H;GI($CX%DHAZ!5.8K3-L27
PKRN7[96F1VD5(]P2W)7]=27*_&G%:3GRU%W6)9SCF_OQYT6.@:_Q(\2F%B*2(W9+
P"$)!QH*A84W<&^+>^"%0]P^C,_ U3?16+TD/RH(.?ZZYQ6",KX2_[0K-U)SL]D4Y
PU[_M<@M)<]@*_(E9U1WNJISGG7A5PRCNUP4:$TA!:&>M.%]Z(A8#U&Z<NUEA8ED@
PF"\]L4WX93\^,E]D-M]>].,YYVZ^M.6+6J!'>BEJ[3PCNHH"J*?(9B4I A</R^ E
P5 @-+@?"I.?V<<9ZEZ['[S'G:FC%\12YO"S[O=P^ (1L$H%J*@Q*'Y!J.8K"=Y5J
PTJ>99O'1\(-!3[[K0.NV_RQF!F0I\U<Z-%PTBU@/AC9Z)LIC+X[X3S44NJ'2]T#'
PF"7XZ:_M6@ZQ2C#]8TA!)_EB.8+YU?"]-;?7^)7M!PZCD,#\YAN,4 @&.N0W6A$5
P>;O "E$$1K,V;$GY,-0ZZD/+Y$SG#MH&IB%*)316K_3\8(^I6R3, 9@VX([FGZ5#
P4_6KZD%PI $V-EFK;#0+N>^G0]IH,_S?()TZ\.E?7TH2'8P@]WB^"96#>+B8KXWA
P/#>PU*/;KN1\9)Q;)W#R0X[F*6S_*0^;1^&*05"88D5AM%B&R7=; ?1'77X7YV!Q
PI:<;,0.C2YXE7\#'VK810/-[+;ID"%%2,RG*7;';^8:D-1Y*SD)EK_4GG.\[R]$\
P2J=^$ZF<R!O1'^X*5DDW^GC:ZKH+WY4ZL%&IDN,\.5_B&T0/B5<5:TI)(Q>O.M:A
P=90"M0 G^J*]0Y=-"W?W]?ZR>14CP^WPC:N;!V*1_WW^SY164,X1$"[@0:$^ BC4
P?*+K<1 L>GY :5;N&_[8%.U6T4[+8_9-RO>MI;(MW'?1&'?RXOM1WUU#Z*[I0:GN
P6CYG22'Z2FD&VG6D-6_&=A306!PQ1, [F*=^9CU0!ETAA$>YKB0Q254(D$^:LQPK
P3\4\KMFZUI1/5!:YT"(;*,C\\482]$F LL@K'(S>>W(75#F*$3L.;-YI> WY;!45
PV@I97 D_LD2MQ0)J9'_?@S30Y? Y*=Q'VSSAJA9G.*]R34%3,)4PI%L$7V2Z]";+
PN)9N\9OB,#C-[GI:M\[F &7::OSD]MC_G^J/K*@&5+.0LA/M!V+$+%7.2L8I?3;6
P-,*#@!$=URN)-*"8$5Z<1 =D(P@X=O8.5-?6'U\W02,$>*ATQH2H+,=?( +)SU3[
PSY(@+&!+^CF,X8'E'TSQ^ME.6%I$S=34$332P_$_K<OK0C$W_SWA@8*ILLE5#*$/
P@!*_?UC_)45)NQ"1>I.DI_:/>!*&X%BM:J\0CV68&HK8HU$C)D_H3%K%$AOA*_C5
PY3+1WEZBFV5Q[^8C1_73GF)>3*,U @0%=M<M:/@D7L>-U@N),9JM$+I:J8!/79\2
PQIUTI/GZYHT*4JG;K?8JO=Y_?@?(@8XE1DHJ&Z&WBX$9+3-IMA0@*F:( MN1?CG"
PSQOQS"TRQ+1@J$M$W\X\DL>H<K][0X:0OP9]O64U\8DUM^#42B#0OZVL3]!I9KRS
P-/35TV$P[IR;'QTWG<5" @2?OXUR<9 :A-=.V95:7=2FO$^Y+F9>3ZFN6%ZZVL:F
PBZ<A"PT'%],.)J^OF&J6K#/3JO3/AHX?9W# "R,1G$Q)8C[N>F#6/RTV@K*BL+"?
PV97U) /.0G,S=;#0S4M^X]<SG%Q4B6/_*6*2*_/RN6[CZAX;Y''5I>9LST0V:K9]
P0ME,S31]%+:7/8BCGV1=UK.@!PP%76:I$7Z^([6&@L[NI08-_'L4C5@)CRC,4]C 
PSU6>RW!,@H*M?U3N_+Q8%=_'']OW\<R],>'N7RX7D>@6P. \'4XEFV?,  -!V*>6
P))R(\(7@D7/U@;<CPQ<Z4YC5Y#W;#C_$AR@F#E;)7?^+ACT,V4,1O_D9_X"L)?@.
P2BD]&R?);D2G;_]]R_X!Y?"6SFQD?:8<N$4 9B!=M?9DG3FVVL >#7H5;$0NOK[U
P69HR';"U_#VZ2^G""QM"60Q('W1X1+!'RO&Y)P-((G#5UGPXF(#T"EJ&MF0FH,>1
PJ F*D\W,83Z:FP- ^V]"V#H0'Z)YON/Z]ATUSA_)6:3HWIVJ\.)N5OZ<#)"=##*7
P"5&3XJN#.WQ%WX!VC<==K;$(X5;U:=)(*M@0[ PVD5TQWX[!B0S0#.)PK#*'XU+Z
PB 0>N5#-V\1%"J-1&4/IW+KH0L>)!5M9TJ70\'KZST*!C^K?&_000T;+RM58I^^_
P*&;M*):*[NGW%J4>2[FHUD/[$'\068AN5;'\(>^%\@ZC\RD'SFW &&>!]PIU'@U_
P6S,]G)?25'8?=WA<+<?'U@?+#AY7E$4L?T\352G)"Y/W?/^Y0<VT2+4,DJCE."-D
PA2^7J"VMO%:!_G3CG#*+@%G= O'\15H:- "EE)K?+%[.F+Y6+7HT"XVT3U]]CA$*
P,Y9XQSZK],>O+E!VFC0@ZD1I^B&I8B99"$$,4.===PI&0SI,2<:A!2/3JEGQ@];V
PF%R0].&4&^QR1L!K&]\+W:=B):GF>U)/5@L(@:@&7=LY4[.@T"2[3H8I8?R->MG\
P=B!<1K;L20+'^"W6Y2W12AH-&^^F:K/F#[>'11(#!XA\H**L=T-+85#(["E?.HL;
P==NB.DO3<>@$<S<KXTU<=8UZ0U=6--L:C#MJ43N&Z>-$7EB3SV_.ODNK4&;GIBMH
P$:X<L"[HKVY=^1."'W!]U-UO*)7_0JHK1UM*O+[*(,/BDA+JIJ_CM( S,T:6+TMW
P=Z:R"89U)<CT<S>8HL;HO/T5K1E,0)%%5Z&M?32Y,;9)+O@\EB>"SZLT89_EZ2=A
P#XQ9L^\_3')9,&<OG3^@M#60P9Z:7YJK(]U<V^?13FS]G[K*/"$XW&BAWL3UQVZ$
PD_H'KRM]+@<Z<A69Y$H(;T]T-N4*$UD05(TGMGI5# Z]XX=<UG,>-W@?$8"=\V_8
P6_YUJMZ4XJOPB)7.-P :DPL1P^J3!]5S@;YRSF'8-#X[W')JJ:Q^5N,?'MH)'>Y%
PM6L+85Q9.=*P?>R>Q2[0USMC^*QL^8HSGY'HIK<8=0Q[<KJIS=># 7<>,A@ _T,I
PIX>ZL51S[YO3!['D<D\TZ=-A*3##S2JF(1<(#*7<SICOTY?$6/Z=+I@GH"ELO8_Y
PD*\[\LE(F\;W\_<<VF&9$!O$0##)&74$=&%*^1)[+^,_./5K\>"[SH5[7!V+:=)$
P\A^<)QY-+>,BU,RR=N$1K1YIQJ5"$04>8!;$#*+2)1Y5)KLSBO.[C,KHQ?-SO,<3
PS%B8UG(>9:Y:EH87\_&"$T+O1.+E ;<F-#QKG_D.[LAQ20=V-OI40#Z%U#>DQ1.&
PT5Q)_WSHY!W4+^5FF*ABF6*40#M/NJY!4%96[VA#'@CGX!V]3DZ"7>0=-<)A:,")
P[7E@GBLB1,,90JXA@3V&<D4C3"K;G2"_/2@!<=GV 4GPO6FKS-BR"KZ,*VS"&X-'
PYD!?8MI&.J/;L)4TLJ]JY=.:,*-6>WA:S"\\CRN1@3741M]3-?9"8L,874:!YE?0
P=9E/<T"2@+0GBCW\/T"(B.GV"N>*".1 :,7Z/TOVYB,6/^KTR6[,Y?<BR=9-]4'-
P8-*C4+,2M*KZ6!>J+MOG72[RGT((X9RNWQ D=!2_83T5F':3H9U_:DA;(^<";,T5
PKWE;=Q[W8E<;>@3]EYI#:=CH!&[95(YQOE^%J*CH7"472.&TZ7_&0Y3!655RJ]!=
PNU'D,9*>MHJ(5KY0 :MA?@M22>6-?O*;O0Y8/YO$ONLZQ'-V$X/?4^C<K,(@#ZHJ
PET30[$]Z&_/X!5:4)X_8:95S8+"/5Z^:O.%&0/< J<<@_8[".E.70<\_&@=>>(9@
P_%,KEC3 EX_7K#3EZ^MX!RB_4RHK[-H)2"; ),4B-<BBPN9 .XHHNUE2L;A5/;WI
P5ZRMTL8]>L2U"^"F9A";X9=!9]\8BY^!PP0R9$T&X;?'+Q]@]5Z(<7\>\_O<H2 V
P4Y/V2ML@[[VL\-A YW_5K7[!-,$E=9FGQ]]]*J%WZ,!U=)]*]64,VZ(R3^<P;4A?
P@M+ 1MJDDF6#DP%4_0+6 EN3*7<F=(K7_O),;+TL$WPGN\/X&C#O05N#2%O=HNK2
P\CQ(^'43<%Y(Z=^_/2JI_R\T6U9OJAB1*2%<+@-Z5>'MX6O;0[#=0591S1EHO -L
PC+&-+"?Q;(+%0MB[XC-XV3X+T6KV/' O=27B@/$@1O$ 5#=G9A]Z1VOG[4H\N#\*
PD1)])JZ'Q5V"2<F;]+OP)Q\JGI:%2.".*"U3H1V4$))[!.\8AA$5(M[NG^N#&4!J
P1F%CGK-W,LN"U_N)Y)FMJ-[[#YTR]UM:L<7%&"./NV1Z?>N4,6-&MYD8B77NY<- 
P[8]<EDH48QQ\/8(<8Q=Q2.C#QR;N3L%XV'I%*=F^\)NSYU\,?SS.(XR4D&B C6QO
PLNV(JG+32L2_@^S<\NK$<(1DD$]B)LK:L9K@B:E/)9ZRY=J<3$/X@SXD;UA]$?,$
PJ?-J,/.D&^G:/T3 OZ#:D.D$L%.XAT9SHF_+GQ;@?U)J#ADDN4XB902U#+NMCH0G
P>B=P]ZW!Y!/.H9'O\Y^6*PV]!BGFP\]%7M3=D>2.G(:QX(D)=;7:9B1C^;41$?0"
P\_?/>OS1>]I%"?[BB*0+_C*K-X:^3,F385EJ-66JG'A,W'<V46ANZF*V?<E%-Y.T
P?(39?>^D]],R9.8\*'1\UDX,Z"61PU38B/N,Y P=?G(!MZ;O'DSSC\G[OHW9-(*O
P@4YA1M?\%OLDH9U*R+E.98=GO8Q?F-7<P (P%:PEH9]:>(Q4WSI)%N$(?;;.9Y<-
P<^W$ \%/?(4,NP^Q@_96)BOQ--M^,=51KA<CA@;Z,7D:[&HN2!# >?0!1-LH1DR9
PHWTKE^I-=G.J_6E=\>^X5#S52D@>+6VX4%F*)U57@K6BO+)F >/]IDAC3+)SXT,Y
P]^KA 2M^9#/&PQD6)9SS'Z?LK=1I[Y)I7T,/RPA.HI5N$W %H7]_,TB[@?4WF^!9
P;"&+\_)Q%Y7X(B SN)!>E&R9R5+&!8&;N"-T4"\?5VQ.1[%0*6G(YF5;>PR4Y2=G
P.A#!;8#Z.\'%$ H<8A@?5U/%%V,ZMDP1**"I_SC,]TX?@!5+]A!)1O]J9H$B\'\4
PPC2H95PB]TI<\/Q;D*<)8*2D5[P5V_AY8KZE)*YI)O,2JI"H0"K,MNR6>J6 &#JR
P.-UU.3W(X44=PR9BIY3BV%/$[*-'N(B@,C&,.\(H6D-"J*R>"PPP;4-E-M."FW2V
PYD]N(,W523Z1VXUYY''9<I?A(FG\+/X;4_)?J5:R\?Q_L A"V2X*-B!=$,J["DBE
P$W_L6O_>4<2>U#$4A2TEB1 +BV7E"0X>^RE&-4N-B*NC$G=*_C^XSPA!%];>%U0]
P!C4KYK"L#4__66<67[^,[QV56,B[?+U2^']#_'N_*0W)P_%Z:5C0<0"?,[2_/0^U
P ETA6_4CCJ9=QII6Q]6T5QS:@!,,(]648+:(F+1=M<FB3>1'Q;<1%5C:E^(,$ O&
P82DBG0_D:)YTYP=#;P$/#?[A_W&5JAX:7M-TJ9!S"6E"F!HPDS/;R!#R4H!7EB2\
PRVZW$IAX$321(MOOD!,^.C?"_IJO)U],N^=SIN#IB#=BRZCW;&R)A+3L.-2+]H,.
P6--"=(,<4K'B2V;@3K/,^PE<.>#GE&>TBH)E?WI<,ZC(H=3M 2(J\<?RP4X@^;3E
P?MU-TL=8V0(!WC^^17S[3@X4U=PXD_*G'E9'K18<66XYUZETMYGC2C-X3G#K4%GT
PQ*#\%WW6T?3%_^PSO6BG4,["U%K-CN14YZ#8)8X?KC$@3WV. _*F% Z(*K SD;2$
P8\^*&5EVBG=11S>Q%LSE(>0L<8B% _60SZU4^Z22H_T=:\#@;*+@& C>(@XO MLT
PZ<B.NW6_9; &HU[2 OQC<7#;C<8K@V_^DKAV33OCD&!+G-\_YN)V0YM<7/FZD1*W
P?%1D3CKGX7&0.*A=/3.@0YH,\<\P;YPDG69YC!W.4-[<2^JFA;:EN5P7#D@>^T$;
P/^/:7)8*,P-'N[@9%*&^:F$<_T;:/4H6VW)G8,!C)H@7@VTM*K%;<-]QGM20I6FF
P7]073 *[HYL=6DY>=1?%$CJMZ,?6T%MD5I(9_B<?\L)EI8>_@KHC0WK/WK::S_BU
P30<PFVG8@H8V)WX?6I3XJ9-B/0 /UFNT3'*IV>%6%;2L2^: H,, 6PP)[D'76Y_O
P*HVA,E&^K'#@T&H;I5 3587.5U1')A"V&]'LQ*",6QNCE<7KDXQY5!)4Y=XU8E@?
P+)Y@9Z:T%]<TS+S5[\0;47AU)4*PET]]:<AOT=IWCI#X9>!VK(&<;;U47W_9435 
P0Y!1\PGA%P\.YRAW<U/&"V"/ %3B/2%HL7&PP:JEPE=ZP/6+WV+"V"$\R5+8F:D)
P%T/9Z,/D*L4K*=SLU?YRY*A MR3[HO9X9L6 @6+>OTK7UI]?$7N:]14-,(3_A$(S
P!><&C)SOS_.6N:5@G@AXG^QB8_ +T^FE9I?.,K)87#I"=:(&[7/H =?H5%7#K>7E
P+;$\*O\E4M0_+\=/_\T9;$@=F\H#FUX!N8V:ZKU;UA4^Y-)4*LB_+WUA42$MK10+
P8U14JK%%ZT X*DK^PGJU8AITL@.IM1Z^.+N8@-)?>.1%G_0!O&[PWU8^N_54PWM?
P]&8?S8('8 8$YB5K2S7> +$!UK-R7^IY\C@:7S;C18U]P/?^-H'[SPC,"?!XZV'8
P"F" =[;+4?^<+T_?>+^-A8.JXTXB&;I"J!$E1J@B2,<DGH^FDMU->/_2_$6H2C.B
P3+N<+YPY  =B'X=UEA!)Z&EJX^RN6^GV;7I5PR+ N8WYO(%EI%>)=CE++\9@?O.D
PJ^Q3+X5\7=VZ\&2XQFC>Y2] D&HB^,=[K_C"SR2P]BX&.R-9YQB_S:T%N#XDL90X
P8'RLO'_36Y[,A;]-SNX@62[CQ7Z^[\\)EJ/%=*:0DK,R)$^R=.T%K5RAR5*<7)\*
PSM(VUN!S17$$&N&N74S10/Z8L.A(9F'W76CLJEG"2Q("/91HJ3H=\OU9*D[B/ JD
P&?+:GESAPBX6<_27&KS-1&TTX"(1SFCAV/<#6;A $SYXF2<6/E:ZZ_,*M-OXG52V
P.[_@$)AV1$#YRJ/K<U5!X;OVO/$&!RN"8%%U\.@^9:ZS,-FP1=-/].5(?EZHCTVB
P'KTNKZG0*BO4=J[5\1P\F$I-@9&-5-J  *\)(RWY2$Z+U*F)?P$;[6UD<=U# RW_
P#7CP(3.;UEH=P_F,==GW[V% [34*J1E7S<SF%(WJ1!'FZ:NE*9K0:65*EG]][.O4
PB/1DV+0W;SN#O'V3CCLY?WG.;U\,?9='Q .>6M0/WK+_""/G'IT]G,)QS1HO-27!
PPF<Z#AP'MLQ:QPM]L=7MF)7FE$#+O3I(B-UK@!2^>J!?V3^-5]"Y<.F"O%Y3='!*
PJA%<X(I?KG]J 6U!?K)9DHNNNS/D<OI74M8B"O\HNK3>0Q5;IN/@0AD:UN=K?=(C
P?7CQ;-HRL< @$_@,\^U^C=E0:T!WPD'QB[(=$QQHR1D-K]**PDX65I**LX+O3>CX
P+\W;6H.L60!NV(0L2RG>U[[.:LTTEV2:$'V))X-["!T%/A_ QGY0L_L=BFXY+U9H
P8)5Z]5^CU:;ZTIY;R%<-)RH3B??+S*R!DI6LTY?/7DX&^+YA\5G;6^MM^'Z3!PC:
P0Z4UG<+.6C"?HJ0<G0"5/SOC3BSR@U"65[M1B8M"(0YHBE[RX41+WZ$;.7Z2O6"'
PDX:F^*8LC5FS'GK2X:TVDZ=OC38-7_H4%=SF9PV:D-,$:1:7-LU+/AGQU7^D5V9L
P<^D^?LET^T49?I0D1;+=%^U:@,%N9@_2EY+D7O$2(ECLB5MMV0NS**Q.\K);>=P7
P+&!I?HU3K4'3?7,6E28 +!)D9>NTY%Z#%T&R=T"5W-K"<A;<! ?-TAKDLT:B\8"/
P927;#AV^@^R0Q&-$$%ZLBL>  "?7AP]E%5PNO<P/1@V6>TS*5C/KE;>L_CA:YQ[Y
P22@('!Z?3D=;.MXF"]H];T%;/^.LD>577],''VS*]GG$*9'4D:F/Q/7/J6%^8,O0
P9[#V,>9;QMBEM=2;)"%O;>@:84Y$[=ICJ9RRX4=99.2;UK%+3N,:POG^;XA'!:A]
PZ6UM&]%W:)%Y^B=@;L.80+N?M.A-O.#K119G^DN]R@$Q_B*\A0$X:&71XWK5O2YC
PLG&9YUV33AB&$QFW;*O!!0XYE,Z[\VP43;5!@^_O'3W/Z3=+J+YQN34CGE("B<+>
PI25XF+,C)99%6TBFMP7!A:RY=S?#)%(12.91M=Z3$'<@2(6?-J#M:6L[1+$\QET8
P,!1>\F09+%#\G,;*8QFE+^-XPHX=[?8GD&@-:N,HC?@JSV0_-;#%8,72$$F:3;<7
P\VP;+H6A2;YX#"JEG2>*5![@@Z*O[=1!*Q+F:!B"?[O1#G^D!O59^0ZJ(M&STI2P
P;/ S"<HW@[UZ![(YJ.(SW5<KKYD:*!619[T7?U4:>%1G[R'2U=3&"E;]N1I)(;=[
PG8BZKB"/O.#$USX;@;D+9-:;#-2QYJJ%?G[V*M<ITU!'; &@14O3^':$=7'51V:)
PQ=BGEKQ@VKA%43V]A;^UZ&$A)7-:FN';2J!0#ZRM&/.I3]^A^%^_,+6(9;:6N8W!
P\$(DPKTY'6QFL5XS,A;\0N$A^\M& !SWP8#ZYW\NC)>):$7^H6[132%Z2CP_E;-&
P'%3L>-4P3]O_:^M*+Y.O2!B!8R 96K=(R/0IU5A"(:%L1"#'PR4E[23-HI17S.]O
P[5M#]\Y< 7SD4$8J.%(3?-D0N!VOX7*?1R\RTN_K9O_K26E96Z9#A=[>&]MT7/UT
P1<?$W@2V\,F;YQA_D_7TE/L<F(=)42@30[2B:<^)&V"W7_QC?U.&]E87B&)*F6/U
P';G&V$32?!4#P\_E0I57Z/,Z!1S2./=@@\']?(N48D?MV&@Q>Y;J)'>&J_*^Y\"=
PU=/&%M()2W?I_40(4_Z V4X4FRR^>3DYC<)[F%+N3.'6_TYH9>@JU(.!MZ*3,1_T
P5\M5S*:L#D$TBG;M7]X4RA(:[Y.2!"@>!ZM(-'1S:$ 9/WFABSXHL:04Z$((4&5Q
P5D<6]?[VW6C)J7]EO'BE(  (CA!#=+NNEE(N!OCI:TQY-KUS[;+FV&)65K%N_7W;
P>B%U2V<L$H1-JJ4O@PXUF1E&JKCU7X*!A1L]9;#'Q.=P*ES%L\C2.''T_3!";QR.
PN,8'D:DF7S)+>E+Q@Z13=M518P6[0QSS??J\9%4JJ&,F)J*M28C=J'P=2&_>I@& 
PA)$+ZS/TDFAMS:/RG$81>UDP#*X!)],;O$61<A:Z^B!4!J*RU=8%+].,BY#%DQ8V
P 40,:$'AC= Z++AY*V=Y,0- 8CHUF[\@>>^4Z3\A4;S;':SIFPA2.Y!'*?#C92\Y
P#L[?AHZ!U9<H,D#?C_-U)GF0AVW%*_I+"[7&/6:#&87UBR1V9;D1XR$",JE3K^<?
P@-3/#%Z6C*LY'+,'>*MST *W35?--E&'(U;B0(1HT%G9@C)9<1\3;O.'4+=#]M &
PFY^F^7><'%'-CN4/+".,FZD!Q',E!UX3]+O8$'*>2"PQ*:NVL4<J4,F)V5=599K+
PD9H(!6=C2DT18FNLY73\D[@<?=@%S9N+>T1RXR/'@Z_=)9T/9U+!F2[EF6]/87]<
PROMU&@-O=.YM2$KV>%M7!@NW#Y#[#*I-]'XN;UIR[+*1Y:-NMB@F!]&>2Q 'D3'Q
PEV;/V.72(L2'1S,=4RU_67M.M8@O(%OZ:2BB'@_?%+'HRZ$P\& J4$\UE1G.>IV(
P691,2C,/KI6X94(5Z&PO(31R=LK"B=P9&' E#A880W;P%8+X57?^5C(= O0XWTMP
P8 29_DQ+I-TC:A@8VL'87:2K/\HA8#,KN1)3+^VTSG*5U1"#<-7/I/2;=GAG*Z H
P,=>9GF,", CD:($VUCZ:7*/F.K',.((7Z?:NIO#23RM*0 VA1O\EV"3;;[NTL^H#
P^507]$ZA/C8M9_ H<"$#+-]:B "\G8F;Z*M<EM_*M/61F=&=%7%K';UK;8"DRC2/
P/C @]\MJ!0KGUM+>=NT_U6*V41)&>;SW*>R_&+%1P25=I,4]K>K7;*B+APG_)?+U
P\7R&* !V.PT"5$:-7/IRYD&++CY>\_RR>'V=UINU!/"7Q (,NV5.0HBOUR.8*/[[
P\JO M0%O7U@)A*0&<(6F]*VX=D6M+=I9+>%I'L7,HBM, ?(*R#T\$:6^0X(M:][1
P#Z0(N QAL?N"]G2-*?5?WXVN<4M]&UD2VT RJCWESK7@*GR2_Y;N+B;= 0Z&V';&
P'//\"F/CGBZR#JT"&AA;E;5Y/[#/KD>2(@RC\:X-^4>1(7MY4 FP4#0A)_Y#_'BT
P/X+.#OB?DF@C""Z@/C$'_!Q^ RY%#$GJ6'X\#IQUQ*^6/?AUDU"_NZ77 WW</+?E
P6N %[(:#+25T7XV<[K]V7Z*O<_/(X;7\Q/K$2/)F&)JW*'1"5#S4LDI)I"D&E ::
P;TY!A)M_G_52R=)P,)XN/IP>#?3MM6X;@0 &+JK('QI);S!"FRCP]>E":HZ*U*R9
P$854^ZA<SY23HKT! PLXL\= E;C6L Y8]OX!'3-Y_,>=:D$&$N^-@D+H*;K9#&2A
PC"CZ,4"QS )-?GR5DA1Q\'  ]:0($CU)/D;'>=I"GQLT$[\B[I\Q)QC<# 3:\50-
PN#&AKI;T:)"5Y(F7SB!O05J*KT%!;V;"FW"9MV'1)U"3N:6*&9'':?6G-#O">2V2
P/*3(8RRB?2-3-L-84?8I@.-Q+5S#=-K=8I."I 34>"D9Z"M_*Q(%?B<GM;C,Q<4^
PZE,,11@5&U*#B/YPJ=_8SX0C>VK'A??"\C08=<%"__3<+[?:18^?9]!654P2JKQ-
P$7V1>L+T1V=5<7!O>%X)K&65+114)7&N=HL0J[,Y@OX4!95B<J_(/1DTEC!4V" 7
PL&]J_\/T)BB%)I!YR8F5&4RN_X!]1%%\W9SP).A%J3(%]HQ7.$!_(,5!S4]F@?T 
PI?)#[7)]PZ:>I0^H>(!DI@&\JRWTJ6PJ8I3BZ&3 &IE%O;LA19^CG+ A'H#ZT_NR
P<%%/BND5-(^M88=^R*HLI.ZN2(3R<DH)5L?IJIY2SYI WD.&P&#%7*TKQ00NPI63
P-CFB]U2G6NA6<'?KC:2_NZVI4W5$2@" 87%\3R6V"%)U0N&(5PL3N>/U$/"^?>07
P)'JW/=(;KJ>1]H7BO1@YBE$8Y*R!#I\ZQ6633&+$ __S=L!*B&;#1TH^3;=LAP:!
P JWC(.BWF- R E89*Y2OCSEML'X^(7J,?#[!?TG4S-@OG&'^.$*7::2T%!)0R?%^
PGFY,A;>+0C< =BJ>?7JD4EJ8QCD$6^:EEK*CIK6;N+0X;DFNH?.]",@9)U("_=*"
PQ)"594;))J8'@6+3L)"<?,<-?M:\S*)JY"PK\.['QZ&,8NNV"(F?=J7/WK(Y2M4/
PF9Q#M51QSYX?IR]3A@[B)KA^ Q9P/H[T+^N<CSFK"\;,T^J@F,_!Y)6M]-D+Q4] 
P'.^(5B=7XODUNMA_N.!F),.8@F6B>Q)O+JC-^E"CHA ]E9P9@[T>BEAU-E-;&4^R
P#<BX%SQ^T8,WQ<YMQILO<0.2%9]S=X>:7\-!RT6JLH0A32;$]]H%6@9CP=6Y'&>G
P;G.-VWV&>:84#"1"-24XGZ#9Y9NMH!3K=]15P>/=R1 ?Z_7#7TCY8UQ:V#K.LNHH
P=$M\E[9]X D#G;=%4Q+ZK FK.\G")V5N0WT$+)%$X![QU.0V0 7&4=+;(^H[=M;?
P?IF9>C0$Y!/K+24$YC6T@WY!$^8!L6)';D0\LMA9DAR#93KCGW)P- CF ,9*1FR-
PAJ&=@?XI1V2K8+6PW L]TU)F%DIU^^H9V_+- T+$2X)1BV? #"]>:[I.JYWTRD:+
P.V6O&8-$C4QQG\QGOR%I$TY+F D:2M@P'@)%R^70.> #_; L-EY/>C1C B%6(?YD
P"W':5O[2D#*G&:G%#[DN6>![5_DP%;EWDC!!-JZ :IT$Q8!%1Z(P%F]_KDE_EUGI
PZN]>_FJB[EIRM0?T'-.NM$M!%E,O0+I:L.%8SWFI.6",3M68^0,?60Y(\?RRU W(
PKH!/[-E! _;[/T7RZ;X6C_E2DWG+D[3%+.FX=:/7]0:OP)U/Z+2O'9:5.)2W[Z?R
P L0XY8F2BG_#R^NGH@DCD6E]E3%^P-=SIY@MAPSZWKP99IN )%D?X&]X/F5-Z&YY
PW'?3C+@PYC^ F1R^?G4P;.<3^C9O,-0=%D,5_J2;#&*$RPL*FEU1+:QXX&VZ$E@J
PK#U5G3NQZ?.4J)O-+,EY$QG.#:+MDU1RJW N[Q!""+K+[X\S^AM;*L;P> (]JLF9
P6CCB&\)S&12&/EUL%1AN#@/T-P!6UE<."U7(2I;]8'B=+935!5'#[L*N=_ Y#T-+
P2DWB/6?\"VGWM]BPN 0WCVF'#<$TJ)3[^PYYGL*S;IHJ$996J/H2O9+YG_Y5@G@[
PC0E9JH54O@Z%<P4?2/#TWPAR.J;WI*^1T:&U;:A$1YZC\:U6ZG+-PT'#CM6KWT7Y
P8A)Y^H'_?)W(].5=$KL=-)G]/*6VL,\_WJ4\T"IG_#>N$+D<U7T*I_HQ\N:2;6=2
P)%*D92N,.I5;T.G,=4?HK?[[^K2W@G:297*!<"<T#^ONP8_0*K1"[>#Q!7!N4["-
PN-].\O1:K9Q[JL4?/*&FI5[B^V[K:&IVXTGO8P6=-8LT/I->)RU?;-Z:AX.,\<SP
P LN(@*1T3Z7Q*9,QG[?E9E<?+2FGCLZ6(S7"IH%V1!V<7"UM-*/VV* LJ&;1L=3;
P>HJR^P_]N7Q7LAYV<B]2O4F=;[G\*Z(-+SU)<)=01LDII3Y!$ W17# +@[\E#&I?
PIL'-+0+CT"=$F$JK)S"](K*&BAQC3!FF:'W$NL\.]*SGD"UVBK?1K/"YN<[9,!E2
P5;BO;[V<U[\ZP34:%$$03Y 0SU*&!_\F@S#+1K#"?10/M_%/=35,W)X:%%'ST5:L
PT*#"-:8S*X:]'XD:53H,JK<O@EPVLAVF+=>XK *AT<'0#X5#2-"6YB>TC]&\ \6A
PK2Q\6+T8.S.&$M1!^M*T+]%(K8 O7=%[TLX?_6^=Z'[E_4#C&[%53\X+ZQJ6NI9 
P\4!'1%AV&AZ!N<$6K/L%7 5J %*45@F!O5CQRS]2@E7VI$B.PN^:G2!Z<>IA^Z$^
PN6OA_@)NO,1+B<H,9[8K9G.?R%?=4WF1"[CPS0TEC84ORI"V,4G^L")N>"SLRICH
P#>H'+("3_M#-#^.0*W)7U[K*-(?:9&[;KAE\G.]+CII%GGSI]]]$SJQD\]53D2(6
P%T<'1:E^S[+OR0V4"R])SPJ03"HP%7<E(-QAL =E* '=&T"+H \>Y2+WAK\-+(4>
P%BS"T?D?*_I=VL[$RV#O<#MGKT8LC?\DGU(_<J^4B%AFI697?4+D57^/4M!>.67$
P=Q5BUQH[&FFS>?4%*MB2P3U&,QL"<2HC!8&]P0N; VH"X%A+O:W+L,"C<\%?GN&^
POG-]-TYZU!L?T712T)=S8K<AR^?K?TFVVHO[>(@^%R(3R%B^T(Y1M5(3LW3T;%T.
P^5'M <:BH=IN_***'7G!3?@7N,VB[EL@DO,<B):I.C':^POL-QMM74O!)C#Y"4D=
PXR7W0VQE"@K:FI#*K P*M\2EH<J$1[$<,O%W>SD=<G%%67%+M3+,I0N27H .4BX[
PHYTF8LTS3/;+NO;.S^@)SNB_%W##F)__3JU=-?PKPC1[M#HC^7?<?0@.&@V419I5
P^D Y]?YKSCPCN0+61-Q$]E2OF%?GI;A+E(DY(A)N33J[<9A'X 7PNLUIII8*8;( 
P-2-+B<!(-R;B!4G'-B88H0NAZ H]0[I[!H]'=,0UUS%*!56JUPU6#UJ73>TG8-IE
P!9?2QI]=DE/YF Q%(TFF4KS04 TP/LR,Z*!*'9?IKLE[/QTQB>+;39EO"2R=&+H@
PN2]T^ALD_OSZL@FR7^KK,H39^4I9:!B9V\M-U"/FXLN^N$HZ _-Q,ZYKJ)?\YO+B
PXMG*Q3\E?VA]SBPG/)7[;NKC3]3%0!;2$)2RBPL4K']]!?[N2N]*@1W$+E$TII5 
P,MJ-C!=J':CH,:?%T^8FWE%FN5)8_EEJ+&\2,=HJ+9<0F-\-(ZCQ8!N67@A<F@0Y
PJV;(LLI=6JI2QTUK3>/@RL\,%;7^UN-)3_6Y;PM(%Q2F^/B7AK0@SQG!C%#A^!C?
PKM2*(*4]3TX*@T2 5WP/A/G'P$#2A!H 4%P:O;IW)/A !53'IM'>DT\*GW:&<O>I
P%&J.]YSM4)(8,7J&[O9BUIAZ>;S2.3MBO:KGM[("&6'=* -67O^;?OC#*+L7@-/5
PW. [BVPQ[;RP2/LZ=(V%A'QA+/2;P714%CK>-%C.Z!\ZBFS]]U^TH+I@1>NMS_<Z
P^:L"MH2FW[.G1<Q*CZ.M<Z<(/8W!@9"O0>P"R?[Z5"EEPW/LMS($'&,!)4H6\"W0
P4&@' (&'#KX(\17TY?-(B4W_@J"^3+YMSAFQ$1^%=!2#.Y:[GHGNP1L-7QNW>#RO
P*-J;U\Y#$A).N9Z[Q+J&$]?P%< $DM>'O%$Q19;?1S3;K<0972QM%'U<W;$M<_#&
PC)$RAXQN>]Q?YWA L.S5WK)5UJ]YSZ*:M#_KKB.U;=$A2?9[ST19@$@?=>L4C!/]
PVL%<()XW;C.EVJ+:QR =R*,JM<I'$'>LR*ZF"(&>I^D9PZUK&\Z>2EB *6<9LRY;
PS*?B69@X5R0\A&YO:1691<@XL \%*WI+//%9E1[^?-"!/31]%.0%;H9CW'6!XOIO
PDKIXY=U0X>QVN08&LCH[0"=6>D)(B1ZU1T:\!N FN/?A8V#CBG3K#0$DH/:9IW#6
P'QI (<L9^AW?'],UB1R-5]90'*\_8*.Z#.)CZVE7JFVC";< 6+DGD.&,1+SH;=2V
PX=O^3(CXPC=+J:]::V&TUJOZ=/QNT6FB\REJ#CK>8!B7:[U>9\B#!"?^A$34B&5\
P;$O1""R\Y;ZG&XR1F@VK#OY;YF?1<XNI%C^PZ[[=C7[H:V,K)V-^(/5?:X>XQX9.
PW 'UR\+!<T;$-L=&96'&3@Q>AS<B*Q@M/](N+T6D:**8N0'04T\WK]_ZER*G#+-=
PB5<1!0<S8PFFMM_=S^8(7Y9S.'=0^W3=Z)$[B9+5%"79DSJ<PX;T,A189_?]QZ$$
PA^QP?6'7D: DDX!4_)2S>%&)]S!8W!(B3$_[#&SX+R%-J0[W8]'.,X/<,\%>9_A+
PM/^,?(%R:F7NG9[AJ7S92^/8C'3?3GHF$4&&UBX>*(A8B6<J;IKS4HD5;7?\MG++
PA-"3DK&-#;U3]"%WKJ)#>B\MC[>G\J(HP1.0<4KX5ZUYEBS2^1&5KN=B#="T=*&R
P\KG#8"8NI7*)N[>;?9RC5'=O=V =UB;Q$BP-[8_^(Z:=-QE, *2*@"/T;<'>D.X*
P?L%96T%5QAR+[?C&^D-Q^[!S'XIAW>#:G%XQ_)_)HYB:^RK$RL[[E+")BP]&89Q%
PK\:MTC$8%5Q-4@4:_V*)!-/P?$1$0.^SYSW%7XHGG8;^C7:<[&<)V?;/3<Q5%UX-
P$[D,'M6!C]@W\4U;,5Z/&6T^8JX''L4S3^\GV8-4@//OYW+G03_#$F)<;D1(M\8_
PN\+>*%,/:<R0;_-N$Z-$&"8H2;<%*+KZ>./[C$5'93%X>_L>.[M:4*@^?"Y0Z!-^
PP4U$! ZQ$8JQL0:YN,">EJ%]*^:3WIS<4, 32J3MV;.7? Z2Z>:5G8BE [QLO5GT
P$B,DF]:NWBS3DM@N52N@$-K!5ZVZD]U0+K=)OH&.R3WJW_$$+R*SU%81PN,6_;P_
PLFYIBZW6#J:1&KR%72C;!S=6H0+I+YB@Q4'3YKT;?)ZV5-H9[:*O083ZDX(1?+"R
PZ/Q@$GMAG5+P+J2@')]F,4"")! O81,TN8[:,EK1Q!TU-2N%WE<:8F(F]:H*O*7^
PA"]L\JWW1\EQ!@0S>*"U7#=!#+"8P"J>1 Y3WR7YZ_9IR&WTW\[O<UE!,+"1!:UR
PF+.A,G*GB4D.3V@%2!M4?68:6:KUXD'Z\;5@^W&4LQ,>'!UX.:"(&<U0*=(3B+H2
P<1_B.0&/N&7-^R@%PCPD!+& O_D?T!A->];847K<^A6:.5$H:!0C, F\O#10VIC7
P1L\93--3:'B/LQ5V\9:"N+ _LT_ED)';EU_]0G5- X<[U[[]: HH?A>%%.="R_9T
P)S&!^J9<X(VDO.[".HUT@QHJ+&T/6DH5 ;V31\+-W/&+JR)5??:C)K;6JPWKE6@H
PCA;SQ27VF&2N:>\_[R^H1>-+21C$7MI]'+-@T_>:P8&D&=H[0-Y.]#&5H_PK#F(K
PR4"UA52+9KM#/WC%9JIBE.'8;OE1I6@5>@:(]B/[GN6!G15'<.K9=RFD$X-*!=R^
P#8P92=;*&^&._5$.<'7P-L0SO%24RM9KS"7)J#HV<.M(XK[#-%\B4D+AQS=ZZZ8-
PT# S.-^[\"90KW$.*J>\KW;#&!J#K_#'3@.)[4ZMY. +^G>&Y[W:[>3%="O!,W/+
PN?ZS<$#'F>6;)V7XB/X?I?N$S(3R&B!&C2%#OTH5\C#-^$;J$>_6-3+AKK(Z,X62
PLZ2'H_V2&0H]B82[0J:,E1'_[ZV7Y@ALX)SJ<2A1]^Q*F$#YP C"T*U?6S%3TQ8>
P-'U)G1F4KRK2>2?1!XQN 3[X7NE:$.8)U[8:J#.@D:LVI HD\.& A(>LX<4S<PS5
PQ5XQ"B@HS2;A*SZZXA3=6PEF/."0YI1M-/6>+YR,<$<G#KA4%J@6#%5^<&V#//VD
P_6R);#M^$?X#59E96M6(6H9*'BD^(;167NQ\8H N_'ICZ40P/@(..W.[(*>4:ZQ(
P3APR\@JHMJ^BYPCX;U6]!;&B&@HU'THD\,V@LZM4I6'$#HW/J5HJ_G8LPF/MA]-5
P[L%73X6/?<XO*I\],"#$9?_.(G+:)>]Z^,=?P$X5 V6=/JD4,O+,TPZEM. *DV'J
P';0[:JR.G@5=R+ ((2/2#LRC9[CT'P8N"#+6L4U1CL MV59V,^)7L!:0$= 42*I6
P@.%&IJA*X4+W7_#>V6LA69+.D!5A3((XLYL>9*:X&Z=@&6F^T[NE7? 5-SU4]A;5
PI5[_HF,F)EEI\19)4X(U3.C-Q;Y)M;)],PHJ C^'6*C3(F<8F@F'/?OZF80^)-44
P1YI%*(B%^HZ6^O(W3*JA#)VNJ*^I>,+CRE&5T*%YQO#,[ZAJM295XA^72GV9N'&Z
P5^66J981!4G!,*A69T)^>!:; 6__D<^0RTSOX]%3K:4;Q%WW:*";C]NQ*+""N\P@
PQQ7;O S, \:C"L%.?8J2#8,ZN%*2<LO7\_BDG\VJS*+AE4\07_13CBS0IQ\T$OR/
P3,@C3LYS34WR \#"?_2 "0S*6'L:B\E5F]FQ'VF.PCE4T/1MILM7<257HD'N?G[Y
PI:"%TQ.WQWRQ"IR@D!$W:#+8ZPRP<U.MB19+/<@MD/T]#R3D/:XLF^[[PG5>^XN(
P,+,<E0VBCC? ' ;%=KDHI5JGA(L6MA]BNDW\\G9H10.;,82@KD&-?>TR*NH,UN#G
PH6AY WG.L&0P3.4Z25DBG%NN!C([DS36UMC DO#D($0*X2?T"#"@E,Y=32A\"&S%
P_!K7A23<5,@??J6)_"Y*I)'#8Q1V/Y/A@N9_-%%HC3J%DH<$8T>Z5%1_].:[Q"'[
PB3VJC X<H"U5!AI6XU%'%FL \9QG[3:KG)RDD4\X%DA_A^O6Y;*SV%V&T0=RF=M(
PR?W:"Z22F_"1=C1C$-TUY^$ARJ IC,ZD2FS.DSU:);%&<[H"OO?YI.#\A[[>>*G 
P(8AGL 'HPRR87?4%K]J3HNM&=OW;))2SZH/%F:-J6>B*9%91?<:+/V>*C)%L"6%(
PK/FT\(=U*9'U)V&!M*#,]8&AVGV*K;;3A!S_U=?\B$V3.CPI/#TI _#HA4!T!)7Q
P%+__$IE>J"-HH>HG9ECOK'#)92JCQ5[V&PDWI=1@DUV_KX"J3=NESF[!EA\8B%*G
PUPB)2 9.5;0F<YNN%DIEJ8 85E6 ',ZR/9'.,L@O/L4("(*M,<C8E&3X/Z6PE5+8
P.ZKP$>26CBEJ;J"/!9I1@(OKX"Y)CIPMQHGO7#B/'O]F&K3=&*IG: @X]R41<LTJ
P)X$0,:I&_E"5G(<#[]1UQY P_6C7?CHIVE!FK(J+)4Z$\)U5=<DYWP#(V!>AXVQ 
P5 _T*;5=%&(M52C#HP K\JJYL/O E$OZ/4@^#5L,^B'$D$?=%:8RF"_U37<\$P3W
P7TXY089?>B>IZ6;6H[46E5UO\RE2?[EAH*HJ]-G$F2IVM-/6A)U1Y'(EF?-(D8_V
P;99T/B$..#0$':'7GW(P;)IF^F)W8QZA>/O1 W%^B(YL3_I\VFZ.8(KK1))&9KC%
P?*<QH-7D7##,JS?:,*-HL&M5VP)0T\SCTNC^D_,SN8PO_W]'4NN)?<KR/*K%(H:C
P.YK80AWU#QNRY5"Q+)YZ*+F<WR*6^\38/]M,AS=(9LR>AU[GX JBZO^MB2CKHCV^
PS/VF%VBJ#AJMR6\03 7. _%EBW@U?K$Y_Q>C4S!='?LKIVO675*.!]W4^+9#O1T1
P&N(WW -J^'*Y_DEN]I.=PX!?PFC! H]$ON?UU 2+TLLC\O[B#X6<+PC3X6!,,\VF
P6DU L-.(:.7X)8,?#"US.BXB8D5O!XF=W+FX"II6*X#&DZY:B? Y@H/RFV>OT/LV
P B<[),>M7U1*7K$YL#+O]3&,%#<_+F!( HDM_X[G@>_F!LD<*LK9GZA?%HUS[M= 
POT&1I:TIZ "BCP_/#>9/1!<#C+JI'O8RM\O_A]1,JK5Y\Z%__?CZTRI$]$CPH\AZ
P[*,<U,<SZ^4!4SVFLB&7GQTE3%R2];IKB"&C1@LL%JCRE^\'\ICRQ/(Z40W=KEWR
PS= MP$"+"F$+\G,,,YW9/D)C2D&$I2!A^+E;,H*ZP90WCW(9&7X_K$0';</49N5S
PELF3HK,BW'XTT*IH/:+INW12-+>RXU"<_:4]C"D/*_O(:)5R^GDFV5_ML+!6?0!2
P+FM^L1G]4[-Q%**:"=[5N7WUHV)CLTB&S^5N^7N4&=R-EEV!Q3N>4CMSDU(\N,I#
P'PQU/*7SEVRV<;J%+N9,MM*;\&7O1)L'*P#B70.D:L,$A6[JJR5O-%M/\,FD6D8\
PN9?M)ZJEG7X8+$5$B*74;Q[K>IM[JF,C^*3M G<DUGYA\!SK&2B:D7\>47W9D/3!
PWR&XKWJ@;,^S=+GO.,5TAGW/AT!^^(O+8KTLE$ZFI7?[:I6(0^?P(5LA6?./*X'*
P=Y(R[L)=6?I_/P_W%H?X,'67#SV%&*6!32.VAY-1[B-H8]D73N:D(QC";WXAFYQD
P?9F]]KE+Y0;!>^I$H->TIG7=O-G(J-:U2:VJ&AWRV2K$1;O5T2H(UJ,[*EBL&555
PQ7>67VWL]'""&C7<U@7KKF7::/JU+#2P1WZ> XJQ2TF+)6)*PISN_!4!U-HS HS)
P;S:J"$>[:]S.J\EJ;FG<4OYP:0D[]VY><+C]4YK$1V\ )IBD&12C]D8GOG#@N)UZ
P4GVSY"U\P1WH.* L7%HV%@C10Y$E<$1=D+UU :I^EO5%2BPC ;D3 ^"73FKYLI,A
P(H7-#<700YY:?^L"Z.>Y,FOE;:S:'R-V^?8Y5V*/5CWP#E_W#B5+>)LXR3>F1O8O
P[*<3IXSXF?M<>A#[GY!N8<)RNH!Q&(:]7R^,(->T_F2:1T8W:+(H/.:R#&.C2US1
P,\!N$]RIP6%IYEOI]H WV&.W09I?R1WQ.Y;JT2.+R>#K!&IB:W9A'6/N_D$UW?H&
P0+/(1C0>22,3WO=8M;\ Z*%XV^8>(U9:;#V(T:(@MX54,4BP7!W^121!G<6[*;%A
P?VYYF]6<_D*\=X$4'K)1LR):],)1O9[O;PF/$C!%R&X6H3H'\BPS0C1E V7,8:$O
PFP./;\.J0CPNP1!E,I37T,G:_/P;Y.>KGIH_F5LR4W@^^&J$7H[?MVW2"D /B+T(
PKFGYOZ1?T3,ZC(PL-3H&<_CLF1%0.%(,-04R_4[%*_GY9? @Z'+6?$N%,:5;^?>6
P.G<\G:>?0Z(^ =,.,;,^>O7A('Z)5SEB4[MKM:G-S9)GG2Z7Q&1A>!7[!7&+JK$3
P\#W@][_)I3'!I)N40\+M>9:N@_+'>@>8*6KX8HN1QK\+L"W=&_Y=J&[665\L9OMT
PR/EJ6M#SX< N]W8FMPOV"*F'@R5GI?C/0!F<6=B@>@'RBKAR]]4B.N;;<!5;0T92
P,':I ;K^GRIUHX(_M]^<"HWGFF7@BQ*E<+]\HW=!SX7/E=O1Z2G IPJ,$L4$UN4S
PUVTB!ZD[ NA'X*(-'G79F*52*/3>^02!&=)$W+BSGS@92%_[4G1UU[R"[MKDEI@(
PP\'M6S>UP&J.::\C'BU5</:)XGLX8\1NV$BXG V^<\CHV4JOYAA=0(H1L##0XVPT
P=A!(C6QNB[6 TCR706"..WV%>-:H%H24O*QTN+HKZ*9_4 N=U>J=8W6<8$ED;4(D
P1#ZQ5A2?1)D,^O%E]WPB/YJDZ8*W+1KL;0*%&U4YJP*;-&]Y]GB7%#E)KNI&CH\L
P_-,2ZD3&7X]N5+TO;S^F7I9=U+ WV)3B3AR4.HQS&K/&U_P*ML#$?!32&[0E5"T#
P3&^5"Y 74P'GO8&;E%3' IU*O2CC)P^W?U_L\O&2U0NJA@^-MJ9/Y]J?7OJX\=Y8
P6[ /TQJM';\:/LGJH:6Q[<V=",U WA!J<V\5YKZ/N_5;*/'KS]G78 <:CW?\D]V*
P<_.#%=E_I"NG<2R2R3$I#X[>7UX-EQ*,$NJG;A%U =9T O.[J\AMP'<2!&@KZ*O3
PC^1NH+T*,YZU!_*@.BI(7B8<-SQ>[=6*H@@1 T6RD1N'TY+%&P&LN21KPSF=., \
P54/&RF<82)AZ03:28#2'-4C_T_^_[7+8,%BCX*,B<QC7&[ETH3MDTUZ/X;<MCX"%
PM?.4>T$#HQ0U'8;5T@*!U[ ;X,JF_J[VM&5:G$@6)?9U7,[\YB&8.:@%]-RLGQ#H
PX$;>)T:9]98Y LQA"UA"[,F2P]4G!L"4JK&P2/ >RZ*35FE!N#:^]29OK6(_D7$T
P1<-=5>CLKZ_BYY^@JW ?*.WV. #NX7#TNE2ZA$*C6$Z;U:"IP)Q5W7Q[XU:U-K9/
PY QF^^A@NN)";R@?[%)N5S#;6@V$P1*4-6K)V0!<)JJ[U66[%?+[1&L23;T0_9/K
P'F:#I8]C@\/)VXA9;.O="P2U!L]S5C) G#LBQ()(2RVZ4VM<-X&WC6@&W->*B3*"
P[SG4$/C4><M1>42FMLL3PY #+%EABE2S?V"['&:1I7H1@2 MC(PYL/%/',V5LU K
P*GG+O>+%E ]&D,=I60EL6?8*F=AMY)CC!S=Z"%7'%*/%12G^(_C/IG1_AYZH(%&]
P+0:@+.;?D="ZY/;>&5N)]I$DV-5O+#O;8C@A-4W$8NK"7MX6E$Y"_HT@9XY4!M2M
P/F;79<_><GF"V.!>6C4E3B4B"3_71=S,1(BB?KIB6!#2$AC0%NUY*P+>[$7+)M>F
PM]E6?>."R(?6,IQ_S:G)"]?W9\-Z\@@9SU-$P9FDLT6N?0&,$"4CU\CQ%1UUV]*%
P)^*2 COGM%Q8UC$+J=$$,/^#?P084?#5,M19):9CE(I3^[!Q<4%5K)WV@S%$7;[^
P'-6F </O/T_^7GR:S4[R?):@S43OA3-I#\=I'<'V '&&A+P:VP_NBF:B,KV2;BBD
P"SA'?W^?2>2WDJ9@_-F=A@!G:DZEJR5$?E63-DK-,ET#)9Q8^IBICN*F.U*I01V#
P0GE_J5 Y2X%*TW_8P5W$B^*6EE>%K0- GQR*^O_*2#!"!,]6W/S9[#Y5BK!<XZNZ
PP:>+EJDG"/U6EA?^)N>]N;0 7LIA00\Y+&60<VY2:B/@K4!0PEP[%Y9E>=_M-U#T
P.@+]0DJS"TQ7)X :8J^];\JUOKGPPF]6,P2/&(@((+$I%N1EN_<DD(,R_7[6S!LQ
P,<AVLY^LQS/>M"'&_38CY+0#3Z$U0MX,J&!YQ:+QWY# ^W_*-TJOE!Q72+_<@6DR
P^_;S^ Y]Y^<@Y(ZQ(F#;VNAG3+=+RQ&+[+3UW;TY*\?>ZPO=8A\(#BP$-ROW$HWB
PP^Y*B!4C(OV_S3)EF^'V\TO,VQ&8^>R:4W4[!,GO+,Z5N ' ]ZX,;C8;SL.YY%=B
P+'Z/I5D<Z,4;M'W Z(H>%QPJ1>]=$10]**2$W>"ED"T6G30!/&^-L]7T*I,:5XX&
PZ"^TW#=$+':JYR$@*'[*%_T$>6?MY=8UW9S#+>F1P;%>P9LR9FCSD/X>"E5(Q.L?
P:+C9>'_*A'2O9I"9%T/.+3+:D12);@E*UAX#AXC&\N8AYBDD%L2\_.VHSP8/Y*MX
PX6 +U+]1NOG/SD^+>-+=!A>[F8(L=#?QXMC2IH\F=VR/>8-'#J."F<N4_^8K=QE\
P<3"'@0P(<=N1$A<%.]U$?D-HD,*XOP7#F@D:]3O1K";BE57]'CNE<P87-7:J9S?5
PX(OO$,#80CO1TD@SM=]"N^^J^ZXY >U6?:=$C5*J9#>.$<W&FIA3>$8Z!,,4^(C2
PB6-&FG/O_19<FFMWUE5F#)8!..)NEM!X-'JG_/!G.)H@$,+R8N $<B+'!5UA/!+\
P]K\+<-BI\B//5 MU/_5[</L(#YK,.C+MZYAI^^6DA[=M5T^__<*'W!<1*XD?TL+W
PBV_W,C8XE5T@YM^BL<M4 2,BV J.A@1;?I1<=ERMW;_99.OBN<64S[O;2![GM,V%
PA<A?,RVJR.=-Y4J$FK:Y!S665R3EYW^PX3'=C#JB@_DR,S O(D6S$N+2!ZU[9&9,
PJ;TU%)C/B,1:T<P8?;E:]T=JS=D0U1*B516CM#-F]C[AS=, NLO;7W;DX!E)1JB0
P3$\6\P[E%.[8U/-*.%XH ]_NB9QCKCT0%;$FLYP+Z(_1_Y$EFZZD_("J")QS2/>K
PM8ZUL-;@T'.!'W"'IBFD1(:2B$I^KFL=M51S"V*?IN6UQLC*SOVH['Q^M7G=*V,&
P.<76+1M=5^XE/CU8EYY..IOG8CC([_(NVC)!(OX$;-62RLUR0\;89?%<,"EZ^"[?
PM!P1)6]9Y'K U4/(E;'G2>>K4VW>YS&1C[/'=6;G5LT96Z3-K6U;4X @$=G89JAR
P!(AJ+(Y?8,VTKOH;3^]]3''K["A%H\%M?S)?=4:,B!7VG9^;Y=,&?*\7AOZC>![^
PK*4X4X\<8^^U-HVR=_3IU//KA&;"&H)3+6ZS*@!#2NHU:!U-;LS>?;-+!.5S#FN^
PN]G HN\4$8Y19^=$OT-M!Q/7IH9>[@%?1/T:*[:0OFUE?V6\!O_T1511#X#NHP^/
PB/.]5B%$[3W^Q:9+#SGIS("['SMX/C%.?]>B[[JJ*733-\5&"NF963L"PZ';LF+#
PSUI@,JS7%]O3)(390HS.<T%1_)!9<HS5-+=NS7Q^(K"LH8T)M3QMB!['OR]&_/.?
P48+=>JZ/.Y.92(1$X17,2XI"FU&GW(K-=GVHE9>'%)](04G4_O:^02&::P(ZB\+H
PE18FY=K?65_[!3TLM=%NH?P7.0_RH[->P+6(*!TW<0+$/!?;GH'+-GX!QG6W5@&;
PG,1_/L.<7,XD!D@X*"#E0E4I"M!6O:Z)!2N1UI*%O2N8VSU8R)1L4 "ULM%9V,98
PT1]&PYC#2"%NM=;15A#W1.76YX$V,H-4:L/-Z7Y6VD!,01BO?;C@^A)CI),2-Y(Z
PL?6; ? "AQZ*1L6K9O2K6+4O$=E)[;0K.3Z\PSF"/QQJPDG:_I<1IQEFQ@4_@J^>
PU:^\E & @G.9-B""Y4[,_X [<B2]N14_4[9TGO+3_2S7A<;:D]7K  G#KP2PF>O9
P$#_(L\R-H9=VB9U%)KVXKGTL/3IZH!$)IN%VQ(?3?!<G/GAK8&*'Z>U%]365B&M@
P/:$J_W1[7CE"M7JX-J.:\:H%/XJF4Z;6=0M?H_C]Z].R/2>]7W5C$ TKSDH XR;<
P%9,MJQ,,#O,O59B!P*/D.W;):WZ<H3 #C>,M&QK8-'#I; X5- 43:76E7N7"%);+
P9TETFRX0M&IF\XB2BA(R979T97F-OT&3T(8+#1/14-P2[(*M#IBMO=5E^^I&^K-Y
PS+YA'HEO$N206CLG[*RG['.^1?_1*Q)3]$#S+)SEY\[/TP]$(9=:0M=2X[!5"95)
P>=+G)9EO_5-*.!=63@C$/_6??BA].!/>AHZ3#*XL^W*P.^0@RW73,O-1K4C)Q_+G
P\?:/YF3"1&WJ5AXD-C7* %O&.5IO256N.9IN<WAO)Z.E8SI#M[*R$@>-TIP.3VFV
P$AA QYS]4A@4>7MUJ4N#J#WY3V_^<POHE N>V7[+WK,XD\;>J! Q5R4M@L*A_9YC
PGC9[KL?ZUKCTM<.JOH0PU_NN-+JB\V1U4K&R-P.;]XI 5$MQNZ/@1#ZE !=K%.3S
P^ O0M=65P.B@!#8OWIP9B9?$M ),3KAL@,"_W)=K@:32$CV3@,7:1L]PN=P"T]6G
P*!G7AB;PQX0DLQ?)USL.1]@T8^^?]4KONMWC9N;X75L(0=H_Z[[M1>7XVOM& \L]
P< 1L^<F'[2!C8D&9#0/4" ,<G&Y<EDFK/%8,$?P["]RM@;QNL>ZN%>8DHB'8:8^_
P_V2N7#%OZ@0(-&YH6QA^6 R1-S@R^R+E$DX,;-NG"(:Y+TD[/ 6RC' JDP?.[0;4
P5-2P[?^9[>+GX#Q58^9JM) X.SA%K>WGHEH*_U7A=1J+0G)(_I3NX10$A0J*QFI-
P1R'J(]\9J^:"U%R_\<)5C 7@<U$87 E_JCS12J*=H%N,#Q8=!&XX+##5\HDPG]IV
P2X"Y[7O\L(RN UCH,230N=[VI553:YJ*/11&NGNL;?,:#, ;H[I[&J_D*JQ-<E2%
PH <4H/I)MB_V2?8WLKG2LI&#849@?)PXEJJNPWOFG0R#F+C'\O_S4K7JR!H5]*+Z
P7^I.H#OBQ\6'3#D_W/@QY8#*5<IDL3P$UU9WSPX(P;QN'ESW]Z61MHZ]C6MWP#R+
PT\,UZB_&JA^UP2>H&4@TD>T-5\WB]4A&.K^1X:\]E0 92)UMY%['!OW+5(99EN0[
P*MY+FK#/#("0( "2HFOIJ92V3)^Y>9,IMK6O5@8*57:.N.$TNN@5^@ULE^("G_#Q
PVI-[B)B//M#16B65=L2L_:L? ?3;A>WPZ0VO-YGU\E&QX>I/GA7J8K%3XJ<D81:P
PKUE;C80.:LVXQ,_I,5/;J/F"VK2PF$)&&"(Y@*LF3LC^':]AO:(H>!-;,@^_WW4U
P+PA"+GV.27:=I+!_T;XW,*%!6B0U;;$R"=9YURKDN&7B)%--:^5B60G,[Z5RO"_3
PML4V)VLK#5!.5#S3;9GK"1YSDFJWI/;=='_ESIYN\3?8UL%E5C6()EYR=5R"??YW
PA 2#J:WKVZIRRP@$+4#*L\L9L(F&O8"/].1W!#B0R" 8?C$\"T,\'HIK63UG !VF
PLRH41?"*<JBJ:H>D^B%$(VPS5B>Z-+V[85+F-CB?]XW8Z-W> CC&T06(T*TSRZPP
P;!.R13N9KI[G%\N:-I]QE<^ 4L>9%1]A-')!'IU+#F^6(' I! <.DP3=FROZSU2$
PB-WD";EB7]@B1BQ+F2XP=?I .UW6:=(B'I SJ@EJ<BUEE6X/AFM+Y1=<R)U30'<W
PQ1=BH9FRBH6Z;RO% L[07C]E\@\7%KW<RF\R6%732MJH^-L[TI\C?D A>LEGN"Y<
P)(IBGS*Q&ZB;G7B8[<+084\^LW2;L%%G\T45G&J+!Q TCTY7C&!IQ*]/;;!\'XOQ
P!,18N8SO1+[NQ@H+I-TP^_WZ5F[$,Z5(*\?7M;M!4?:TK?)Y\-\#E>"%KF9#8PF\
P/\MU[X&$J1Z@"V#;W3S*O-!JAO[H:7^M6%" %)?47FG6!^/I[LW&D^L8"_>*;X2\
PY> S:3-M.5;/GW0/WRNN](G*D$#;=9:O[OHG*;SG>-:D!'F^EX;4U(/Y/ZPCK!C]
P21ZTN;JP4 $^PLFVGKP^'+\KHL9F:^U)%S9)VF\L'[-]O52OOFXYRXS_[91P$F?G
P[*F]QF1MSI2G5.E%T,M<ZJ'.E9FDW8!*1I,6!%HB^67%7HX=5EOM)N3S5-?2<%82
P]3Y*XJ64V*/8Q=)%5K;SFEFS0RW+L=+K'ISN]3U&I:2/'4PG03@S>&AJ(9#**-3W
PJ><U7P;A=#VZH.(EV*\_(GF?13K,N[!>('TL AM^:C+826T A %):T1R\79R$BE+
P;P==3/T6U:L]PM3K!-_%Z\7?L2@1?! -+A_YP2N0")D-!VHBP%I!(!!].V[/&NK+
P:Q@=,>?L7=CQ>BK<#TTAX5M&?2#!TW86QC+0OI\P5LWCZIU$>K861TD!>2R5N#*"
P4=*<]^&Y:8*Y4[M0/@IN9F7E_[8B:2V_Y]MBX8T@F,37NJG2"&QRK##=JT\S_FG.
P5-MWY#.V1"M_IROU3!-2<O!62\(!G+LLIF312@27YSD(:NA*%- VKP-)"@,MH J%
PI!$76(0W$XAY4J2!PM['PRKCO]J_&'UEW,B!$E>,,? H:@0CM]:GX%ESW.9EX1E,
PD'-XTJ24S;#Z-C2>F7^VB;^BT[VDA1IN.'B2.@R;^1=;5!#FX(!"&H4HP;S!^-?H
PC.<L4LG:XQG'^3U*I@/MG78!4@V_KG0!Q_;3F?=>S!*7HJ>_\D(],_L;K4L@:%4:
PGZAE>0^_'5GKS8+KJL/>T7,;,7N/,F2(@>D3T/9E:I>G\X P&C?%?^.MM+0B-OV^
PB2>XE#E0QTC'C2@VL&4--A[-71/$8<V MN"$,:PL0-J>@R8S8OEU5.1Q*3,Z99<^
PV+P9TC74>:D3O/>K)<T[%'F_%MPI'+W6U@P@/85SZ8PCB(X7?4'(;<RC;X$;H_\C
PU\OVNGJJDQ91YL^'%,(,COZ3'=C>UOP++]/Y0V,+^>BILB=.['IC!3/."RR$4:[1
P_I3#\4[>1[W^Y64%%JYS_E$]2#!TQ%"7PTI8K%P5HBC8I&-C;)I1-5X,>D)>]FS 
P^"R[SQVS?#[\(WE3[S3,S%N*"EN:9JOVRD/_Z[G4$<*+P6YRI4EB>"A6# I+#,?H
PA2H1 $WS1J_Z;AO4/;8QTW?JKBNSJKXMS  9G8-ML2N_PE!U->F2J](7.0WN3XUJ
P&[[Y.A%LG2!1[1^(E2J8X!-;0!+I#_<I R-P7OJD+I[D0 960R(JHW4LQ66'X<$,
P<(A )9MBKC16\X<%UU,T.BI& O]WL E$D/:PEVJ?>4K?D)+$7LD_#VG$-!S.D&LM
PX=3=<0C!!=[7'J*NQV[D-T/=),!+.P?&U6K769MA#&0" 3HO)S/%-LXF22@:AA1$
PH_1$.8%[>6!*\90TC"$!V<*7TZ9:? S%9-099&3*AN5 B2WTAO&X4HG>-5RU&#L7
P@$,F3/)!'0IH2?GJZD$90@/RFC7F3>DP.HZ:8([%P6RPNH#+;[ G9JRBA$TV^ [0
PO[L$<H*+=5=&3ZLSC1"W9#!*Z.\^(\A'3WR>8<=#A+MH^09W,@P&A4WCG_HB8?#D
P<J0/F:=T!R1:*TVH*_>-\)P:YP<YHN_47_V(9!;5R?; M'T8ZP"G6 84?+#FH)]G
P(]J2O#KX<1(1\;&-B$0><&2#0'8DJ+>THPG&7V&/?68KZRAPG\/G#^5K98'7)J" 
P?@M7(\@!XW_PDWG2/H7X;X_*X*4WJL]$NG[/=5GM)!./CMD"40\V)SS_M>F]C_:9
PGC"<K-A:G'!:<I.RX)@AB'J?;D>>+I*')8&_0 M_G6;77E#EJ4WFI8 (:@VV#"&D
PD5U^U;!2GL(S0,37%RSCHYS1J3XBJ;/K_R,*U*I#3CF!888)708X&/!"5?312H+G
P]A5]+N$8"BT;[T$M52+EJ.0J(FR#V68OZ#HF%*7G>7-]:17?D\C1.EX'_FH)\X-6
PZYHH,5<7FT>X=H@U[%/+0Q^8H[GD2PMT@?=&$G]SP=E+W%^6AH=%AEAK!^*:'FY0
P,(:[@+6FX7>KL<?;-9A_KO$(6H^#[)@P^CL^T"\S['1@.P]:X?&^YVY!J=MIZG->
P%5Q[)&KQH 2]013X6/DH15-TV0#6Y6?8.\P2'0C,#M6:W_(@[;F#L0;T;_[<R#5D
PBYY_+ZB)6=XT,PL#%X9GPER7/F[,@N/F&0R7A;,@AF(N9B@1T?.L+>OL%?GMHP'D
P[QMRET4MIWU>GB(5)7Q#&>,[$@ST;RV [/YBH>!YTQD@YK8T8P5"1_LZS@^R#CC=
PQ::R9 5$[JJ102OV&I448*I>0^%_:T=3>(Y_$O0:'5J*U5 2?-@#8ZH1:!(@C4 ;
PG&NFX8 T'9=?^(W];3U45HC,&C"^74^TKV>]868 7,[/ETWP2"%QU=F2XHQ%B2BM
PJ&7^=$+X7+?Q;Q[_N>FVLDH14JL6L8YW8852@9/-MAW<7.AH@K%A',44:XOCV*BL
PH+#B7-!;C^H>O0ZT^WB2UEXEO,H7D'S'T+=B8P:?-.T*2Q>SZO@D4;2Q=&;X"7B6
P3")FZ7;O]+Q4'/2]7P /U&JS])8/A#Y@>S;AS^R2I=NS&9PZ@).&'K-V7<]^?:5F
P^NVD[5KH&DHSNX$3!9DZGJ!"CEA;"^0$B+ AEQPZE/@U4^<=?/%U 5V&/J(F)EK4
PT<@(FT.^1ZLR*2H:NT5I? .0VC#,#.QMG9#0#AE-^LEHH&?6:3Y?U8:XO8]+7QY2
PT"::S_#5]Y7P:*JP^I;<_?Q>+N5$]A]EH"\QV+QB2K[[A9X&7B8_+PV9L_N;X3MT
PG:8&+'@)X$2&V[EHGI0FHP]"H.G@#I<#V(.2YGZR*:.=UZ#$H 8:(=ADC<[G?M0P
PXI,6\M=W(\Q9UWP&P%H[!W4$149(8A!"A/SRB$#]"+UQD83)_^\05GI'4<"6 Q1F
P3[EU7ZLZD,?5-K=QG*%A.:U74L#_.^R !Q;)=O+71KQR>K_DM>']I!%P9>GL]O-O
PTW(&RX@=A.W28RMH_']H"89]^'#Y".,D;)&=0/%4OOA^,5>>WQ"+IWK!LP2*K/!M
P8;X_,L05_Y2<CZ^OMJVSBV/S2[UZU@D\X7E%R&*CM?Y/?646HB</R%Y'VB$A$]2*
P"S=+E&<:MX??F*PB+E?;5]X?J_!<^P+NH^6RLP\!8M)E),\2(KF2]4$C!?/@U.U&
P4FW??U8A3L#./_LK"G*R/Q5/3G_C/@?R,/A(B"IM.DM:9#WYS?CGN1RQ&%&1"O"J
P09J1<,]2"_0+]W+QVN5F Q)Z(!R1L)&\>38H"&((B?M5;S&)!%7LV?B:(3'&K^ZX
PDPD.6%6=DO.6<867;^9V0!(Q&E ''=6\]O:\+/-O5DLB@/Y>04D( RNIA-=R+>#.
P!H2K< I#NQ*F!F']57!#7VV,\5I )>=]0B)F>D5S TL#&+MB\:RS?KK'A[#6W]=P
PS]*7^1TY8I+HDF2CA9U;P#=5,)?VP+XIKZ4\-5K*#2@HQ@K:)\@RJ3X#.4E::P;&
P[ODO6PAS1>E>=3J]]V?4%D<> H1<=WCQC8V2-3)VZ%GHMF 2ON9.]!]&P9,'*(] 
P.P6SE3.'SGYUDHTA@:J5=(ET4G@,/-@;;D2V U@]9?U'(RB_& .-*HOX^:PBC?Y;
P6IV"J86Y8D/+T6YZ7Z<94.()3FV,IME_I,AYW-L0,E$R+CF3/92%,IJ)#%==>.S=
P/*VZH-%5228>LJ[]>'F!BE-+SZ#OMYEGY *\3TN&-6\;2 G 0WB%GP1_]/\:=2ZL
P>$'#]A;X05E.9[?G:'HB#3DY2H@OPBTPCOG^Z,0)>"4DV'Y=(Y=D1YG!YR[@Z<.6
P2I6\4J9;$73BL9</ ;!GJA]2]'C0*#$-8V&5I =!$D=0&GLV%B9'TX12+O2J,$?.
PS<-SPQ.(Q*U]>>G1MX\4;:K^#30;YW,*&L3=QK;P\:U]$D+ -7,(YK($U(PB.D-V
PKWIN.,Y[>T>-I\8QFO:ECV:JQ]VP9&F;B>D2*PSX(_^Y&C&*I!JA2:#E:S@S.W&K
PZ!N9%:Q>[QR%Z60F;$.WDK)*5<D!V.^[<"@MJ7&D$_=GH."C#&QF2E=#$J:$=Z_+
P+98=-7>/OYYR^FC.]B9!4[;,&M4X8= O7:R*D*#G=N/ H,2,S$\,")*HD+4K3ZG0
P3O"Y#W(!_+Q-":I,1[W;U5*>'_=ZQ"JXWMGV85_/0Z-]G9L*6:ZU+G1/%;"E;0BV
PRDY)"PXQ;-+@FJV@6WFJ#LHD#L3^G=^,?K<V14B4;4T^QHA0MYH:GT&E:%Y8](S&
PS?;9N,/:!UQ$0&\Z4J/SJ$>0TZN5>=+,#Y\HH42CS5HEG7_Z1YDPRN:T7#+[Z7U6
P,[^JQ?7V3DPW G,J9( C1NKDQW6 ;<M*VAV&0U!!(*5M\X?:E&&*(<7NF8[JZJ5G
P'_BG("!1U)1%AE5P^[6IF=C<&NQ2UC6&6?A_WZ*M'@IV/910I%;/+PQ^V^ SHPZ0
P3[O@.7RP%'^W&;[7<4_)_4>W-! N:ZRU$T6E#F#?93'N_-M(TQJ_%E\7;#;,0]?"
PKX:K \XLX)9]:L[VZB^].+(2P6R7W9FJ#__P;X'":LMECA=/VT RU0@3;%<]14$2
PKP[\E-2$#Z6*#(PR'-L9*A]3-RU.&-,8%!-A#PD2+: R@1&_3:J8XP*+*!I\U1YI
PPU]6\_T)<CK#'D98<KG\I!9RF!-B\(;5<%WT^1_'><#O2"%-"K#7.1%]$4 -=KT8
PG/==:E)$C\-<P$@MJ.VAD"_#*#*2R3U&&\64E#$,L5Q-Z&.<U340FGKIJI8[!F4Q
P $JJVRG-$KM+.+$:";*O:X8;PJ-[* : *C7AV/9VS%9X:,5[7.A\[C8!5Y;!,K-7
P-0) K9D=X#H+3+69& )]XI&*6GFOE,F^\XCYG*>WVK!>*/1NINK[PXMMI1/55ZU[
P+,I\=IIGZRE?<R;G!4/H?+$&\F$$I=03H7J*O5P^6=(H)6^;Z#%K=A'N<6EQNK$I
P6,V4VIJ]DG$%_J/-.EJB_69:PCHA/SO>7-G10C'NX?Q8H15)%9]6<FDOL?G,(L*G
P#)\?C^^EK8?[H<0U5+<"8!O20-)GFE#/L9$23PY(*;BQ3F76I]5YK^JW(84(K6$*
P[ ^>T5]$H]]#KL4[BM-:YS;R$D_1P'NL9)-0#E8'?Y^1R0;3"TX#JC:/"P@30@25
P\PVL17@N!X^!]Z:['27?0%=Y"6B^N+7*$H&A%>A<.&[8\+!AGQP>!N 3\K&?"6BX
PMA>R &6>HU0Q?P:(C%?I:KC@['-Z7O$94'H3:XSH0X.ST<6OV@CBN0GH91E"(%(M
PQ36RK+7.P.JXBW-_^ MEQRI69U)-D+C%X\8FZP[-ZART]F=CW-(XH"&[)MR!>QI^
P\F!RHZO'R/<I8;9X32#@S0##]^W, .@I11K#-X!-(>[J0?VW[W*QR!3GX6U?H5UQ
P_1!GDS>VK>;UIWZUO@FTP\)#&/!SJ% DJTO7R@OYY$JLTKLV085:P+0=*\4'4,$(
PFP/%_?2 ]"*_R\'9N2! 1"1AUU45%W0BT(&VI=U:6^S!K@:25EI[%YB]Q"CZU]&5
P#E8W*1>-\A(29@_:X0U$#_"*>P)]:V"9[01HON#/ =C]X\(F*]7CXM84F;VDZH=%
PV3L<-+-&8L(S[(Y6=8#\!XDCA94G2O63@N\=7]3/<R9]4<P6MH5;P(Z_F^5 &3+R
PW:J5^N.Z_ZQW6":3S#A7S0>[FO*FC?=P S;E6P0K(G;/(9WW&$:?'FW*O&[;UF8N
PX-6Z:3^^KTW*$T!S$""@#>R'8!S7@[!@8<V=?H<9GC7N4>!A0I0U; R_I-LK=!(T
P1'OB5V<,YOE1'!QWR'C@S*Q1ELF)].;A0#10&$@L&O8)I!JAT@;X<@R:1?IYQ>% 
P+7BI'K<E;9#VT8%A<UMN//N%V\QJ)P^SFS%#IQ*#?$3A_Q_G^;8YK"0B)J^@V#K"
P?>LUUN,%XWCR+?[O88"I]\8G;*'; $YK=[]UG%*63J!<?23GZ]H5"]6-$!7))A%X
P17V_HD #**0UO*/DA#ZZYOHK5=2<4<H-&96_-O9-#]6INSU0@,AHWEZJ6P @9"I3
PN=WO]\MNHO;S/9C6B.SA3G+*L787_PUPF84Z-0R&C9X9:.5K\L$4_1?LA[5^1+?:
PRZ5C ]!'AJX%<W?7^+PB5Q/<VD-DDZA<8GQJ:ST1JOSI7G>I[VMTZB)(7?92D;(A
P,^N29AH*.>9'7.;[W/F R*>9:ZTV7S'5]O'7MW!1/&Z$S$H3(C@-[*7V;<KJ[Y&9
P!)P9SE!=;4B1_@4R<4'%%*CJ$H(#\56$[,P]<K!$V9-CY^D3OC)1 -URI0-*P.H6
PQWG70G1EUW1"(S1]@,V]=X2O;\$^?;)=_&S(MV>\AEST)_(!\22&-F8J+#^.A)%E
PF#-PA,_,N "IH'*6S.:>)EPFG3U5C[9Y)<(O][0O;WIG:@N/^[/%;\OEJ5I,B)KF
PI,1[*%KP_-\_ +V>3F^MU?DIIP9H#^$;]2(Y>1FS,DT]$:L10.M*]39CC?9CFB>+
PJUN4QKI;-L(<:T,"%3[Z^$+ROO18;TYY^2W)>N36EV8/<M:_T<-3!T_7/NR;TZ#$
P>QB'2;KH#5W2&I7+^:5WH<;=-J@0J['4G^K8H[XI+FX-Q02E2+A(JE8F1%W7?K'Q
P,S]C1]_3CS>U?A2IBW@F2LJFB] T;=[1BCC"J6,J&^_!XR=.D^-#0&_"_)D%,*M/
PA0@2O\!F'V:AE63&(:]&[JE5\?+5UX^R&R/MA@D:6UY=>P#P4:42@CKW!0N-T4#,
PE2MJK;VMII&%0E;WT0B^M6<HS4&R<8^K77=-7RI8[Z:@#E'.^?E$9M KA&,O&DUX
P@NZUGVV@,!2IY,%+W(A[0;I0DY^<I5CY1H>T%*@@UP>.%[N09;*\-C] /FZ!96H=
PYCL8E*1FE]EBN0)9U%SF32$F>"%$$,$*+W*/ $FIU-VR(37J4*[=\%EHX&L%*?#L
P&J)L3)\76+K])?OTNH43Y<YY/IM2!Z?F+(Q]V_AR$N\Z4Y<-VPHQ-&@"MN%F0,]_
P]O0_<TJ+\/HD:W^$?-3 R3I;>WN3 8VNY[+UJPH$FM72P]7K(Z#/XD Q4+%NF9H"
PG"V&?> ]87G0%*P^E&H0N,!F>ZK_4"JRF9[Q0#[:[6HP&!W-AZ3N8YB/!ZG=*=,.
P[O#C"?D!6*EP9""S%M6;3HW88D8:2@O' A4.3"0']N8J+N3TN)!1$GEDD_X..8:R
P,-HR*Q3*8Z'XE1+O^&T1_!G)[.GM&RV_>] Y06(;=^6#U@:%7H<1\UXN"$S@;GCC
PKU8W;Q<696LWUQ^B9+D@63G>>WTN$;6),N%9=<OZ(N"'_K3W8+5&SS4H4![PLU0W
PZ%7( K1*L/?$Q7TP\!ICIB8</Q21!E[$6Q<K(GKOK@WW30]]$]"KH%FMR<:_O\DD
P0G&ZY+CNF3;"PEAA&O'V>*EH7A!.P,ND\A4WP#&"#A:K9O%M#1]H@YF13&&$6\LZ
P& 66&JHT!HXH5JMIB,R@I/@K VH24@G ;7(PH88X_6A3IJ>@FYF+;)X@$?!N;.,B
PC$AH])'3P\F&F?COG316FS5&-]=TE33EFHYBAIW'K!#^/>". NY=52S#IG2I4_<\
P/A=95#]O)B9GPID#FXP6@-'2>4=\ C=IZWR[6^^^1!$M[K@QE5K'6\(%-"/.B:% 
P^.03Z8!,^MZJ^"%%J?VYM,UHGEZ$JVY<VUCV'-6&&;@65Q+J8":6Y".4ZW7R&R#T
P3RL4?B!/-H\-Z6+>FGM%G/,)8$:DXWV>.K,B60Q ;F&$ .O)IW!]QRQ(]P2ED 7C
P7B$O>0*K\[UAEPHIX9I7\3,H\"FO#^S/?UR]USGK%L]J% -6H,I<H_D,MU)>CGAG
P,LB+,L$"C@^R*1#S-G\!6IYH2;^?B@:).5<^/(4F+^<65J39F=!$U^3AZ'OKT%@)
PMHV/'8IF\8OZM9O\0K5SDKJ7#V[NJ5TFT96"L(#FK(]<^C(/AA4Z!VU[/HTI_+%)
PK5XP5ZPSBQ1'6M3/"N!4#T<X%M8&C5VM-,9D7L8E(,>Q+:9M+67Y%EA6V[W%/(OJ
P.K%!A@.TWDD$44(E*[Q_7G\C!Y@ALL,?W6($_P31$.4FRC5R629_J64L# Q-UGE&
PV>[:Z.7&.-@\]-S,3_]LP[HE!80E6)=WT_; *A2--WB%$O D<Y^G6<XJ#A-"CMS+
P.8ZJ2=7KO9@7E-SF8:MS N[^X6O+..G9335R'''L(VP!U/[\?PF7>3;N<0=4/4OG
P4IM6,;4A*W=XWLD".#BPVA5$\-YK7R#$VN\..YYJ,K4IAA9%L.]D>/9^':GKF?CD
P10_R-F'+@:7J,Y/L<5)'.W^LP;9G.'F[TD<L[EV!T.G2<(@NZ<KL %/U+^U5L66J
P[+O6_+3@1:R3&B[K;KO!@R"UG[YDY<=4RR55>]@29RZ;M'EA?P35(TL7+^9H6/]X
P+11A+@=!C_\--W(".J.>>W?^CX'_6H(+)W=>M(82;J#7*@ $C$])BQ<[_=X&;*+@
P64RFTZR[3X+WR^9<7!0J]QI"N@*GSV#,=@U:""!9<+=JH/5 _<:F^/1ZSK7-6:_A
P /;'2-,6R5TO-#Q[=&%?T*RR.2.=-+981#&._Z9TR2?89B"#4ZOV4:N!I32HK&'Y
P8>CA$SE09H@";W(AZ-2EI8)?ZD+J>&4MISHJ@KUU;T,'A].5MOHE1T!>K%NBH##G
P4V4:9U3N-(>+2%8> 7:^OS&7/N1P0]W".0&6J'A5=P-Q"?U.?-#@)^+RJUEED*S@
PS,-P(#4X/!CN+OG$-)[,YSFE30L']M/.A*/\*K E'V^)JQTY_-WWRL4D_K[O=>],
P@TG\^+'1'><YP^9?,YI*)20 YM"SO^ T#_U<I#;&IL,65#]<_$Z)I])4#L6 5:VK
PB@+M:-F P1*>@HNSB6%\.3X I\Y/!#.*+R<:GB_O#!P_W*[P2DXJ\,<O'PW.Y@0\
PB_LFP>>999>R>:QB. 7;>XH5F0OLV3I*8!UD/&["$HX'KKUP3&ZH5D%=!5L\-\#[
P7IBX#A5PE!:["SR *C>8Z&OI".4^_9D+)*Y*TB19!?-RVK:V1Y( 5HN25)'-1C4X
P4IFD"6R03;, 5^I5M'\12&5>5X.$BH7'G+^%DD>S!T9'W]V>*>X?)??:S^-9>6$2
PC&4WWH9?B[>G^7?XR95]U:V/HFYJV?:D$%=7 T]"VLZ/Q$-1 L>2>YL(5]E82S5B
P#M-R0:4W]XF-B_J5'3GNI<^["G'CP"+-*%$'UAPH+B'Y_BXS'[IPDR*'P[PEVDQY
PX</]X5#OH_D;/N5YV-_7MB,H.+BQ,^<X[($@&AB;K$V0R*%!HCRTSJ"CDY(0T"&T
P6_WFRP"B[YD9,$NY.<]C?@Y-_(GMNJ67KDP);;JX("*>?DED>%XLQZZ%!%6@OW& 
P/7YF[@>+JP.[2,/;QH%#Z0V?HN>$4@VX-^'UTEC44(3,F:DI4,[:/"?YQ143QW C
PKN]9;#JF*034B=DBU_DF2U:&XPM08N6L#1BQ)--7<Q/1FEQ^#,M.E4301$/2]FK/
P'I'8-&>*]B@.B\& G]1\O?\[$].IH$A?81>W&.LD/$EZ+W%CKUF/!?$<8CLL,C "
P'2V!?AOPZKKU!@FEPD0CF$3:N=%+LM9^ZSE8]_2-LUP$WAD6T*K-;+.+ UT]@:VK
PV?V>+QIB#E[E";2KPHA=C/T7)5UX[O$0CO=9F2N6K\(0%P%*W'4'!S<C5.:TXY)/
P)1Y9NH'/NR3.T U_ZA[#-TTF\JQ7E>(K/5(!@%[&^= N?7,I(M+4LJ<IKE/>$NHM
PP'B3?C1E8^T7LQV\7LC-I "&,X[W&KV_:(+85XG?6L>MA4(??><+?QIG+SE7NEU&
PZAZ0"I!Z[K,W0I&8B8QFI,)S52%H^WA5'M&(8-(Z=B\DWJALNS'<^:Q(/'<2FI^D
PPC\/]GPQ1VE&!&4PR_S5H4>ZP:B6C@E.4U7J3UDU^0V\+"24:'A<LNM96*YV5NTG
P&!'R9S#'\V>YHG-7^HW1ZQS[E7+!Q\CL_S,SHV8GJ/J67O !0ZKPMHL\H1C4K <E
P;?KGH%.0(XP6Z*UUY*Z*P:S%U),7"VE7W'BZ*"%,IT,%8*3IM'I7CKG#K$V=4!E_
P.A?6!X*3'S(1NU^^EAM.EJ!!*UL'D?KJZ!.46:64<8VH9%?U_[R1&2#M+$5P-TOF
P-S(^'<A$1;U $2-V)@9Z^84MT 8G]IHFK9EUC:]H6^ OE0@VNX/PQ\H"F:")F!4,
PVH%5]I>:C34L;"O*3F#_4WV"CC2(839+%K[&F\:01KNZ>K17+%F4-(NH>&!^,LT(
P4BGQP$C#AEEAVJ?:$90P,5V1RO#U4-B0Z9!:^1_@M*2+-7<!SB1^8C<^@F".K%';
P-2!!DGV2I[LW([QS[ T7PREMTEH0K8SX]*RJ%EW_3<"!"HVNR#FT*"DCC\'PFB&J
P[FW-<_.P>:^PFIQF=8!\G-D'&BO[_?@ZB@H]N= L82@&8$ Q&S4V0"-<M[D:<K/#
P[S]MS:-8V>.&P"P2OR<K].BVBX=O[,T6P!TD#O6VK@$YRYH-<I9FQG2YO7Q/<)Y$
PP%UZ=]^Y).MS1\%Z9>LGC5PJ)6X>N+JR-O;]Y; [6.G/HX#\_([&&0U<C:3"DW\/
PY>Z6D? O?\YW[B]^D"W,R,;1T,^:?S[SWAN7XQRQ2Q*5L*PT>)\"DYE;;C!NO60=
P1GNX#J]>N!$;'8,+II6/8?Y$(&K\'EB7GY[PA51]-R6JF=U+?J\>?D<:C_ZTMO;J
P@1AU>K;LT?,R04!Y434DWMVT"M6(@K?0QO6\,"<N,I%HN_(=>PFJJ_O)IX62.92U
P3XITDUU5Y_V/_RS>43"C2*86U7R(L^3TJ<H3FBY+9SD*0_Q*:^,@6EP-X"0+N?X'
PF3N+$M$\T]!2=:G&_9)<^WB/?SF3ZQV? "1\S!NL_)#M:0B;GZ]XWA,QO>:_:D"S
P.C]DV![L#>EXB!H6S#H63WGL;])6RT0X$2O 8:3Y.W@1T)#.TIMT> %/,.24EM/5
P[&=G.7KP06+QL<NZ4$(. CC17"J\GR#92'+3XD[6C@UA*!0O7P8V%6IC*<7IO$_W
PT7X#UCG(L*$E#K<Q$H7V/)K;C?7K7L#^><NZD(Z'A.D[ZM;,]B)/@]PFNH937FAM
PC\!YY6\G1B/C3W3)&Q>WR]B'^?M[IR_6%U9KX<_QI>FW,$<@X*IGFRMHE"Y<9^O_
PBA!C >NG]>D/5+] =E )\/Z"SLA9E@G1",@W;8:U!/.4+GF@>(P1B/I86;-_-OL2
PBYYOIM5\>!DG\,%R*U.&I7\7N?*GD&SY0]FYKQ/7"2^0)5,G(^RY(3R>:UFMD]=T
P,A,N&+P1Q5VS#9FQ J5N=UK&;R98AU=Z]F;Q</B1<>GB)@PVIO/C0D2U_DZFG/.3
PEVVE(5JGZBS1$C:S_GC*LDQ!^8S(+IF\.4/3TS2!V6;^8.W\=%"^*069TX6@+40X
P:=<V0_[EPGII*P4B*5LC; SQ_'EP#UG5*QHFBCLUJ7V9/,XIK$4QWJ:Z8P>3!%Y@
P_'TNXJE88"&B62"G- (U+VKT^&>JR5$KJ"@!Q0,5O&QU4Y913T.[E=.SB^(!X(X.
P-,/C-N;J1ZUR<( 5T=8(,_W!Z>U^K!!\TSJ]5(-5_KSA6Z-H$TI9"^*J4OV'KE[:
PZ(.K%U?$3BDI:EI_5CK_2M]C6%P?6^<KWJXA0]F XYJV>1_1A.*:(]$R,2NRBCK.
P!O$RL-7X$5ME;"N>ZT1AQ3X4PN9=:C+VHK-/9 K8D\S/$@A+]_)+-*E)'_E-.)@%
PX*9EW_#C%0D4K1K'% G$UKH#;RKXE6]2@D*L]>378M7,TK)T->' GZ_5P-_B[(- 
PB0.QH[\2$<XM/H(R;IZ@#ND%X-1Z?<!R4S[GI;HG+.L]$IWI4Y2BZ_(=2*9+ASWJ
P%$Z:C:P#==V5)'^.@/FZ-_J*DFQ@; W&!;\^'[!G%FRFG%Z JTG@(\4#KM_:\"0I
P,!WAL85P-4D\6%F=!1QF@@(JK1>C/&2Q2O%;=4W(?2#* ?32?5[(E@WQ-)IAT/0K
P$G9Q=&80G'V3;_OJF;J4P-&;KWG1!H]0C5&#]OW+$-NJ]EDT?6:3= =7ETW&Q);L
PT8"5]!3,FNM6  NQ9\:]%KZ6&S$L&#U/O'CNZ&,WCQF0T9PI28( Q9!^D&L]+2X\
PZ+\BMY3AM3(H<5OJ9Y(L_   K@ABP*5T&X V#"=VU,\^_OKY2]D4K[=9_(B#C-P1
PP?U\T&<#L&T%&XQBQS#0V@+6L21+0[@KQP]9'7[OH3YZR5Y+&RWZ[_O5IQEBBG8I
PV22(0^W ))@F['!Z+,]AOND,2J[8[<71YJ(=VIXAO;8 ! 9]BH'U'NS%6F#L;EEV
P#?GLJVWM\3D<8Q&R/BF*$(,K1V1JP(HKZ-/VW"=DSBM0GS8OU)FAV1('&<M/IT P
P>TET:$?8<0';H3)^).^,EU?.5@).0W:+_P=.?<>TJR9ZJZ6-T=U-1,'%</V+8Z84
PM(G1H:C9\;1?RY'G@%ARZ[*<%,30B'!(5F8E^QD,RTW8<=9L X:Z,F!%!7,'D16L
PN-JJTRHC$P,(("&A,QUVAI[J>;P;#!V\--R&P_9.QX-Z YQ\[;GCOXQ"+%NMW%)D
PM\E (56E-'M7>T =<?JS%P$CF<F=K#%"OH1R_2&H\^O,7,%)Y%'>M -M#@^'RPE9
P=\KYF)=I8-GGFJ3>#X69OW;6K4<<F0_K/6<F:8=9?6-]NZ4[,.-C\*)P!+LY=):Q
P7-GS\GL WVX4S]!OY7%VA<-:UY%.Y<V%&M(7"=>-QQW1ZB8)QLH64X)A#@DICUE-
P;N'?ZJFR9@>%LS-,\JG:UV69ZJS#GNV(_Z.B]4'YL%7IT N^@6R__[_8/8S_;F&]
P?L_ $G4=8\()\H4P3N-(8)K# 2J%)CRR6"8()61I"X@LS*62%<^#2\D>5NE7K);[
P?3U-O?3 JU/1"U,YPF-]QG-5_;LDD0;E$,Q8$-]A$4O^6=Z8I"AXD'$:\<G/,@LD
P!3?+B+D+&!O&T<N94<Z>Q.[IK[" Z%;&;59%;T7?+V D,:!/%8]2I>)KZ)0-+4QF
P5GMUK;%+C2,%V:ST>[%+^)):PU@V/O.RVHS":%X][<MS<*J2%O*<Y6GWZ5&.YD]@
PW!EN/^,X*=B5-_?F=?B-QME/CJ%K>OQ!PHR$_J0UQ4D4RP:"J[(RH_8MY0!)!--9
POL8.](33=(>A^!1X# ]S7  ?"Q92JW.;[0:#)V=C**3\")X&BG#@H$+K&%F#'$FO
P.N7[Y,0>\';O@/.VM<;W/%DT,'HC5T3JRFKK>*!ESZ23C:"?;^DW_O<V@M<14^-0
P.);AN$NT[*-=KRT;$XE9-._EW-@"_'1'/67*(1DKO!XV- SUB]TG:<3G)=HP;)FC
P*KZY7F)^(XL1S,?4M>A_XRM&DC9355-'!W?CHFW]2SURE8B=K?K(1L99D-ELLA<A
PL5AY#YP\AZBUGC LA9 ZLWB=1#K\M8QJ-0^]J%D"GY[PY"#Z(;5Q%KMP!8,T+9EJ
P=VY'K$!C45AJAX:O9Z9,=W69'SXXN54Y4^V"6^.]\ ?&I3DA,\)W=*^*@G2BFH=C
P\(#3+H:%Z?H;[N*@M05,OSTX^JPK2 CE<-YOISC>!4ZLZ?K VZ1>6\">5X .<98O
PR+0$3ONC!&XU9"HT-FFH$VU5+N:'C()_DV)9]P-RP=8RM@S7DA</YE3Q.=#8B>[(
PYVEV^+X[Q<P70:];P"%/F0<Y6KLX?CHEY6R<+92CH-IAYF1(Y@D.Y09,;U?=MIV5
PB6FU=U*K8<!C5!B=;,U;$J\ <CL$52:!6 %%\K9#:3ZL3+<<7Y'O<H[8XE:G!*]Z
PQ:VR].6 2GS*E3!SF\E4,X._]YHGX_"^&]>(DQ7XPL]C ]WX<HE>BQ^-"BNQBH\/
P3/B/< SETW[&+F, S7-LDHI$^N:]/L[>N#"8]BT'L32V'=V=4$));R3&-9WGK;-L
P=MQ4,(G(V-ZF$A!M5N'"R#A7P%0I=Y?*V?3:V4BC<0"=5CXZ5;U2F;!N?6&1X-X]
P_,D-^TEK@,"E8JYOE&66_GDU<T?!<\-Z?D74<CC2U8U+9N$10FK5!?Q?NC(OSJT4
PXJ?/Y3!MY&8&@-MZNTX;[ULJ"T73JG16#9WFYIC7G!C?MTE(_(]ZFLL4D%6?IQUD
P3$0C* @[AU(3CIS;Y9FSDX71-SSM-6SQ,"/QURC8IL=J:#X%YXUXL8["8G3HMO-X
P_DDH&A5-K?< O*(]W:K^I?)=><K)%$[D9JE)3KK/QX_D*<#]A;(B;K/%''1!'-S*
P.&@,U=%W;>1"\M:K5'#Y38.A87"#'CM#H<I4P=H\6T^J88O3T@=C?KA6\M;UI-9]
PSOFR&E(S1&I2\$:75G&VR5UX7]1\QS^%HFIX;.4U ID[Y*^I =0N@6G\0%4TFS,'
PL8VSI_\V>-H',[S\)MN3'Z.ERPC*1_9P8C$M\$<P&R/;G[AN\=R;#C+2ZKS&B8OR
P"P8,D= )?;] # (<>+$^U2+R](_B8,Y"D$RB?(UTJB_D>><\0B8OWE8\;@Q-U!Q 
PP0<+8"HG+I-M1W^:EZ\C'??8C*N/7$0%'%-O=3Y(-7+C!]?3Q^!7)W/VA7/)D'PS
P8,IRM\#CY @BTHS)*WI(F[+U&7F%S\'S.]4>RK0 %0?:C7R2?[:ME=Q>LQU6ZKJK
PF5O]#@N^1. E#]2"=0@F/4PSBU03CU^/RZVS;-)+4?"Q2=/ -$F<Q32&$WW$E:_*
P\P1KQ\#'[A,EQ\9(N+8&4Y7*@=:%36$SN@%<XL'STT1.8,9^LVPG*>V@=MPE..6G
P,$6&PI5*:>CR[Z4S62C.L;*SQ@B#GU?3]O /&P_N8@X<YHU7@C&OPN?G1JT_CWR]
P6&&&,0'[ 9'#JYI@F+6766/^&DGTO'/5-,/QS4Z?CC[$E2K*Q'@2-/>Q\A8"Z44?
PGN8@)1 ,ACHC+E$SBT3$SX(RZM;+?#+!CY)0/#OD,",B@)]Q.BQ_P9XTKFR;%N%0
PLZ3RJDW=1Q<R=2R8.4_)>/6MRE=]0=]7\=?-;V9VE"#?* 0[;!7Z6G8!X&.#=9E0
P,")?^KMU)(JL!,G0TT0W1:CCE3.OV(]<VP++^,!F,:YW0#5WT-'+/VF()TBW058Z
P-]"UIRZ1* &/TFMFESJHYR\(U<*)FR#$6KE,OX;PE2 XT?7YD$G1_?2FVG_:#Y+=
P]F1NUXD/=A*O-ZQTRT%UR'S&P'3ZDC=KJ/ENN)XW"5N:X4TR!N=D+;PMUGA926F?
P=ASA0>_WGZI8#I7>%[JJTQ_' -+P0XV[JNM)+Y3^:$GHN//R]OH>I8?0+MTKZ'Q[
P6%DT_E"7%]$_W(QFI:4Q]^[Z2GN1MV5H'POTW\PCI>P\&[B.-]H8N5>B*!8*R@^C
PYT.389$TP1@[S[K6^E0CH@YJU>M::8,KE\N"@K*P[ 1%:TJ\2^?T434\UB*\64A 
P"$IZ-3"=)(U@DU]].>HG3?!"J:4+.>MM>@[Z@]@-Y]X7=*XG:M8C?% 5',^PFC$X
P/>OD^R-BN^$H+"34\@'/JIW;^/!5G9*6H EG8*FXJ\0/26C'.]^75,%FS4A"RL)N
P%_243UYL@IR$9QO@HPRE8XG I #8^$3LGMLI3-_V76=4 X$8;.$=AVN;M,Q>,EY=
P\Z!RGNR2\I?#V WYOP6OJJ_F\6U[[%S\:36X0O'H^L 8J#JJ2"4J]C/P3KWC10;=
PV</I-O/W$/\.H:Y"O&96L<MPN"P9V("1:^0?FD9&*"U\$2 =6+2V\$M(+*B,&>.8
P-&8QU[Q8EQ=!EKL9U?8A2M^D(;0%VNM-\NMYVM\)2K;?0(/J!(B085I4^PQ67W U
PYS5)8!9>W)<3EM$@ZT = B:QJ1;U++Z'M$E%G#7VEHLWN].A"3@-^PJ$G!92S^_B
P0ZQD5;A$I80K'UHW&8)3;^E5O^-!@P,7DB9P?WM/I&\I\T;)Y81_TIZ/-46<QY V
P+YE\ AE4S[]!C#U:I9:[1M?0,PHXS)T\/:D$G1%G M(O-7BH#!72D2BTQJ$EB;_V
P_%#\L/?KWDVMHHGCJR)+!3]+2S8L<9W($X2_/7$O6[^DW#B-6FE%.\P'NJYX$P[H
P)<;IH$;;Q4"-\64:Z)I?8/V:@P)1$9H DDY]=I$<;6;P%L$^<U!8_>>81^\'PNFA
P$<]@ET<8>6G?#\"?8,R]/0<0Z][D/Y:K@KKB=*\WD/BKW\:/]5IV!/V-/6AGY;G.
P_V&\CA(9U3-M4.RW0-$PI/Q<0I"MLBE*Q0\CH-'GH7Q,'",[LDSIAJ$;8R*!V3[&
P*FEE7 RA12'D[;MU?^E8;C#H:;U[1OXQ-^YVZL4YS.\;5%)34(8!\;=S2ID"0+;6
PN._BU112@N2K*\:/SVB1O;8J-8WF$!6.=@L]%^;-%*"MG;[CP-=@X.4)9[[.1;;W
P]=HQ\$BYTB<SC5Y&O;B)+52R8'#5,:H5'8/OE@W!/?#'DPIK/@93QNE65E8MF+9^
PWY*A8T8VKDW:HG/8Z@;L<M'U+K0R/\+6).5\A?%!I5>?/1;^0(@6ZW-Q:U\+*$B"
PBSV13F-CM"'#)3,K_)75I@(RY?!2(:!@ZR71@G2WH)D3\%8\;RQUF41X7<NS74XB
PR0)-ZE[[]C\U*]1_6.K@ADF3UW-P5U>Z)>*(W*S#0A26JDF#=ZLS"VH!'N<&C'TH
P_%L66H$P^H,V%_)GTD7<FNG7?)V:$O%1?C>,I%<0<O14^$B\P+"\DX8TH-[P6]"5
P2%;))4#FRU4__"I]@]+T"@12'P)8CI0-IZ1![DP BI:S3IW-:,9XSQ;K!M&U:#C-
P3\?<I O 6%_QK&AI[N8N#I"*X/N4(S(JF9RAK!$>6H<4*J>4\0G1F15Z[\'<N$2D
P14;L<Z_4T4FZ/URYRA%'*)&FVO=)O=_]1!6N887CF&-?](_8^=9%0CYO4=$K6$DR
PIC6ABU'>:9Q=E_)=C7>KH"XW%07-TCA[R/MD\'DC&_1,]X*E]N6[U']LEE]+!)M%
P2,76O7$ME@$V>Y^OE]3!X]0E=C@$V)2)(_O;D(UN'5(\7(X!\U8!0TKM_J!KZ"U4
PB??T#.&XXS:G'F4R)V9<%\5YP#WV=;8>S)1E)&4 BXNMZ3HP]DJ A1_GY*:ZRNHR
PS;4P+ T+*03!S*$NH.RWD[,&I3@&++0#<;;SV'4-%&HH+OE$Z"[W&4Z=WR(@M) J
P(NLF!Y16!1H!SQC-)HV:5R.P?GKGWL>3RGO9=1<!6UU_?+5\Y7)_7$T@.)676CHI
P-LOQRTVX@N)?]R0#I>B9_:22+ZY$5$B,,E'3+W<%DP@(L$[BI4_$N#*W%Z4K OP.
PQ!>?Y7TSU6!N-_28K=_@S'UPYNX?IP'7#QXS<?>1%Q#$QLQ:4#72LUFQTJ4\;*1-
P'\[\-C!"QAXAA$OGDK.5=EF/:9J)U8(VTR"76!P9ID5'CR[N6)T :LJ+,]EC)SR(
P$*Y._&-W)-='C]EIM,F3&'6[PK7+E:)= XFLB)82-&YBK$?8^+/(VXK?_(4POEX1
PMP&3:V\-]C+U JA=C.Z\FOE0%+4L'&L;4;*47590A_Z0+O5M4B<?U(OP3LJ6<W]B
PYB<'!(BE[SU+E"QY4(M#$'/7!8.?9)NHQ_?9.I(391$WLA.GFTD:^=C-0%A(BY/K
PS_,)(PI6$2>U]5W9)+RZ&U1HN>[=!R+; ,0%.<ZSLJO5MVW]0\4;+NDM%$+YZ5>H
PY5'(4!.$:1 SLG !@:<HSO%HY\X6/6Y E9)OS190=6I>S.G+ 'N]O:).$_M/UM85
PLO]M&T6"#I>#,QC<>H&245CWH7#_WFC@U<DZW]V] !-;$ :>4 BCN'ZN18NJB<] 
P25C2">AS<BT-T$I'Z$X>YDQ"O97!-9$@?W/71 -@9*GDT$6^8?$$]AJK4$U\%) S
P%#EQ4,>N3:';%-'[\L3F&SEO7JH$!1%SAI#('?KH3MIV'K#')]?C#CM/#W!'.;@)
P:,HP*#\MS.:_L[/U&G_Q\,\TT+4_"!DZ=TG,INKB\;]U9/K+H3$X74TMP\\2BFMS
P'LAOE!S^]"W')^LBP??C<),'C)+*;F0GOP*D&?:T3/U9?R:H/1XA8[UD /O8W5[#
PW#8<Z</V=-!;.CKEHB!*ER'!0^7@9%',3@R;?H?5T<!7/"/]3$Z6U&LAD:MZ2LX/
PQ!;9./-1WUOL?"013DNU9"-+BX;/RG_,>.01K>!+(T23QP]YCR3'@J4L82RRA=5G
PVI *K >D<3EE\34*FO/&[6".3&RUN(&9^V,*RMKL3[;/K5 !":+;19;*X[2M'^',
PDNDLZGT4P_[VC7\!9"PNM=T?CUG##G$4IM8@TQ-%YX2B&68TT-T8+2Q;)CA>X&'^
P LFX.5"(EE$B[+F&,2G@J(U5%&"HQ@^IO(]?#.X=)PT6JU8&N7R=<"(9V=N\ER]%
P##?=<J][)%4SYP9,_A4'Y;TS2'25B6.>$9.6F5:+ 5/36.XOP0P;M.YH:EIHC'6(
PHLE#$>=3>S6GBJB>\XRCP7EYN3MV03,^_]+0&9[U7G+78[G3/OR8*GK"L>S#MC$3
PMORJT<.UG?,?E4$'1 JM9FN51?:@F:7J*Y)25/9(4<7'5U&S"27**I?_81,J4\;X
P-CCGP3[HBK&4G!OYUT% F2"^ 6,OJ!0SRZ?NC18'%I*(8JS]8CP-TOS02&<8W%1\
P0N]&1QFE'+NVT=$/\ #99:FE"G,R)JZ2*:]\FJW36;%3:7)_!3-JR5PEO.JL4Z%^
P5Y/(9!Y[1R$VD&NX\C-TMMI@W;C,UD)J-9'^6D;]I@6S2(.TRT^C\>,ZXQ?$?P#$
PKBP![6WD'JW4&NX")]7I'#)*M5O7O?M1RS"">F&EO@$-IVZ-SR#QGJ)%_C<,.NS7
P\%YAL&#TQFA>KEWUC;C '3?H N+Q+_"LP?BMO_1>Z?%.G2OF*V;L;;]HUR]-<U4S
PRW;:/"_M3V.G_U_[\C6^;>0#? $O^-UA!\/TKKP5T'^9@F\33>1Y,_27, +54WS4
P=IO 3&MN5T77"8\(N"'=.N?3M0X-*T^V'=04G70I)8)9[WFY.D#/^RJUQA7_';01
PT9FZX4;D[*DZ'3H+$Y_A.VQ_9E_FVYJK3@U'P V-D6.RD_'SFX5,NK M%05/_+U=
P@\OTS4J1KF&^UIA1L'Q!I6\OB:_7&8 9Z*B-TMUAVR=U%,I35L#XW[/NA?I9!LY'
P2\%BQ1;N4]_\R;_0YO($G+FZO<Y+W34;- 0:=1U@N(4RO'^"0+(&ZM93UT^4<O#!
PS!I"Z%'Y.[S$C'=[D64ATP6X*[YZEX+3[@NLQ=)*OB_'+?#J[L)(\1-#[M&P!9*M
P@M;34N4KB?03T&6,SL^Z-!Y+,_^M?F8X/JQOX.2>VVCU>1QK1CA["MT*>4JGC.BK
P=MH]]0NW82W8T9AIW2_!/AJ^5S,E=@46E%)/GA7RFTQ>8*<FW*:U%]^>1P4^O^@I
PVQ$/1Y.C1;;K>!Q<W+?E '#WK_&X0?C6>'1ZD%T5)?\,U\]U:1K]QF*<QT?K$7)1
PXW%P3_KYTQ;E#2&D6VHT[!NZ=^PH."1_?%7"P\ENN5G30K'DXRKB4>A70?C$_E&W
PFL2=*T<Y(^H3>>N\Y3<*\UT IU)IH%,UI5CM*7?/;. @/2_[*'AN=I.ZTF[NX;24
PN#HL0%X0"P\_7*T\Y1_BD+^_>2T3!2:\JC&//+'C]6&V3[^*TR<C1=P G JZ@3?0
P,7OB*T_*HKD 64XMK P9A2 0>5\T.0S*@S%6I,7A\]U4*2M"*/2\JRNE DN"XD%>
P)9"&"@R=?O[]#&+2_W#,^[VD#Q$4RK&4E)LL]^!XU'TEGCD6!I:_EK3V!!!!LXR)
P5YZCW, S3"6BL3?Q:T'+#*#?_/><#R;^4%E4'F4/T71WAS*8K.0,U#:!'[]4H+*'
PV9!.GI*V,WK)T\2"/19#<K_M&"\Z<D9T1*I-\+H#^<O)%%U+VLFI/.!#R6E(B'S/
P.U2$TV+5KB-I=97_+K=YV^F'2(E7<?T?JO*3[$? 'M*NRRQ-$%X^A^C7/H(J<B$N
P?778:GS(<*N[R/>M%KUPAH-+RQX9?ZNB(=Q')%%.6*E9!X87U)6!>.6)>N:%D ZA
PU"&D\O7T,5ZY@V",_Z_F]*X)3=='HZP$'<XQUR&'*7^;B %UT!XL!04DDVWO*<>+
P2Q&W4Y8%FWGVY);<M%7R7(:=QU!!?UX@]\7YCF^Z#T_N%,&.PRF%EQA0;_.5DZ.\
PIYP3=ZZQL2)EN1]7C,K\*G$<:>'S8ZTVP?B6X >%,7_H(*[+#GEIVG=)\',EU+9T
P4VND[D>9#'N\UV)V/?V2:[0GU%E@$ VO5OP0H3I"O[")-30>:;U!3_>E.Z&I!9-*
PZ.N,8Y96\ILPV04/&$60Y-*IQI;;NGI\6@K/=LM#_A[9KXYPS,)1H34WXWDW?G]7
PFR%8U:"JIW]XRNH;A#BU($IM0^36;'@N/TMYF1KTTDYGH-!C:2T"C8RWVP95#[CZ
PJTIO/4TCC0\E57$MM/A7'3.ID;W V.X-:;L4G*FLHBI3R'Z*6I9FX#^;&<GD3@TM
PZ)T\K<(LN!_]"?R+ED)9-[]2OL97[TZ&1S%A]J=<A^S<"EVKE%(..)QG3POGZN/E
P\K$FSQ#9-&!6[?+C,0MRG'3*CZ)T79HT9N%:'+W>\4Y";8Q>J!_P]]5SNCA*#J!V
P>(*N[K*N>UHU9RL[6L1!.=XK:HHCNW\,>'Q'9K=% [OU8->87$63+(6W&HB8A1)E
P?JA]T!1:D&:?!/5H[?^]$QU[YU&'L<^!)WL%W#(_?HG6/6IB 5Y9%J)G6XD!>#=B
PUZ6$FRAUJ@]NMVKGRJEGJ;&_2(]SVY;S0*\ ]P?]6+IK_KNS\3,K;%@G+-HV^:LF
PF>',_A>>U0SKQ4Z/;G1.&!IZWI-WLTTP. +734$!(^0DOJ/[+B=T?/>9CVP)<MO3
P0#:.DW_'&; P&JO?J9P=H"!P9^V-Y246>L@Q*^?QC;PRE=F%BVB.$[G"?K6S&OA9
P3-Z,[F^"SI!'%4U;2Z.9$M@?\V)0QJ^R$?/0 B9=C)T4<T&,5^81"7H2+"'\#X @
P3'QM [P),QNROITHJ$ +PS%@>+7J#K"))Y;Y&F3!A\)]#!8K)),<8FMXL17D&S+R
P*5%R3W/2[U VBJK$'K=U/L,06\=:,HG30V+1XH@4VLK?'*6C/[>OWAK1YK]@K[#!
P9_V3U6"-SW=>(N7A%>Y8_,F57GP=]' ):+/(%EN^8AS]D/K# 3W*XSH\3)6[VBZ0
P_$#ULD_JUYJ^0:-B=P+@J<T#W? :]R*]HO)%'25=W@/]2FTFRBMF3 UU .3Z!SA(
P\ZLIV-?M29\_5ZL:<;ZV(T:]V!-I^\Z]UNL?&+OW@![OV)%^$V;O$ORL;8:;[FZ 
P"2K)/NY)CYG-U^A:%:0&I 3V+XQ_./!_';H>J5,YVU\FHZ??M8(E\,.H2@P,"^_1
PL!HT:0BZU-<K,L#3 J/4TZ+=WZ?'#'EM?ZI5]1ILX^Q" VHW4]B.;%4L3[D(HAVD
P'6,%-[O>+5"LY>0-<U5:HJ!#-.D$RFK3ZD*ZN/%QPLQWO@1DX#?#PX%V!O#E8 82
P2O1VR*#F#PC.(,Z<OR!L3UJ5T%;.>AP.(?3_,DX^KQK1:G'&V&&S;P3*<T_:/ I(
PD ;I'Z(N&&5[ 47K!?!+UHHN:%TX>NBW&PQ78=9X<'8/=D\[09D-],5.EN!U+4I<
P;^7$2':\+AUP_1.[BC@T#R''ZF[_> &2G!-B;Y=@'"U0^9H6X$. !GD/Q%-.*/W9
PE=$ 759_D_&(@3 DRHZH*4 >E\V8U:?*GRX#+W257V%XES0C,=:X"="0 (B&/;6;
PWMG*P$7^XV/._,8(_V:5KO!=P .=7OZ=TR&,>Y2-MZ#^60Y=8[+!@+JP&FV5IXT[
P0E#FTQ 'KNHH-6_0,# /DYXOB3$SZ$+ Y>*YZM&:P^$#M=:!Z=& M^CVJHVYV)96
P\1M6;(W>FZNFT.53,S"(Y8^U,Q)E%FZ0-&B?2A 6<I3K4W47\9,3MJL6O[3H4E<Y
PM53HB[3%?$-7#/2-LX&UX6F5+N61&%86XRJ4FY6*1NX>%Y&FQZ4H3L 6H6K;?VC?
P)#DC-2=74'NSEQM? B<8PXW<N4B+Z(.:(41ZWR?;+BDFV)])EZ/9P2U!*GI <._)
PMC='7UZNX6_\YWH#,@8(_[/ SWKH"(8Z,IJ;M7' Z<LK"B-/7D]&^#8C@F&Z]KZ<
P!]4M)HR:=5R%=!8GRQ?V>4T/NAC;\2%KRR.F.WY\"'USJW_$NRQ--@I0/GBBI'1<
P_M[E1_%W-@1B_A3GE[US#:#3DCWJO\?YF]3T!E $Y3WM<(,FA5Q+??VL&5(\= 4W
P <MI--TT'\'R@*23IQ\V$C4OD5:)"(7M4DWPC[B[=74X*OZ5P84L#$S^;/Z,8^XD
P?+QOR60VY$SQNG1M._#L>._]*\@(Z +:+OT-=X:;.;')?I&/!H)1IU<F?!>X)NZ"
P_-0B'9)8F[A,,-+; QXHOJ4FI.DGOOY93PG5@^*Z<D.%JE:[&;<@3!&'>S%&KAO 
PDB]X7%ZUSB19[/9[/=)YJZTFFG.W_!$+&Z+@YZ WY4UU5Z!0QP;0Q36BV OU.)IQ
P1W61B@ @9YU)?@08P.IE@?!C42$07._3EQODH[[RZ:Y_Y0/LL##(])$/ZJ'W,\F<
P\\:IB"[3==>VD:)C[IL79*X:<]P+(Q@0Z^70Q82'K8P-@M&.S\XNU(=S&%TCTFA^
PG$VB8P2E,0F>C? 2<5H<COUY!D#Y:A'#^HHM\@ER@DWRH3GNT']Y]7H!<?D)<H^.
P2NT8V 4UB5_SZ:6_T<T,H_H4;2O0(Z)N,72H!;O=KSNJ(R&&2F*0$+T+%P^1;)L1
PB 3LH+W6(WF-K?8*>95>F!5U@=1X%[$2]QVPBEJI*UX#,D/G#*?.+ ^U0E;MEJ3D
PU;RVO=8..]BZ+&-9F.9(95 _NNH%4!J7J_IF8;G 8[2HTV5LK+-+'_Y)AT 5<?&!
P&X"7PL.%3ZP/5W0R39Y4PNVOCV?+_^)QND(A9*(B7ZJH/77HQ8IP@H,7P2>.8ZQB
PPDC+M,^,-=:.\BR \_"7SPAGPMN?D$_ (JM/8IC97!$/AP#MZYLMF/Y?XM=63U1*
P<'EKC^V:@J(V#]FZ%6\=Q+2O*:ZK=!?_^7Y7,BWG"Z3[DZ\;V6C.6V,RR96^4QK6
P(9E3-(.&< 2"L*7K"^>:@%[..N 6*=X8L$NUUJL1J9ZR^=[]V15R]E"[J):&LR".
PQTKR4-SCU2N:-V@X)3BD*,@TH9^+ #/*P(G=#"IN%+1@8,A8;200LQMMO^&/:KB 
PN\EY.9@&J_/Q-F(DQI'@EVZ9NPZ_EI>DQQ\F:E/\4RKQSGY--R'"Y_]"LF!DYVUX
P*>[!M:D4]SHE-\(UGXX^P4Z29F,9"2^4,T:OC+]987+D.VBFAUD;P3M?#R23?]2?
P.5^/Z>AEBXF_<PP]#[4R:9>B6I-(\6*XPPR G1QDDY[9,M/_?8^64R6KMU3_SE*W
P[ZWV^6(VN:%"OU7T:]25)#P -8NJAS P<HE,2@^G4Y*(,0@XI,5JFT"ZO:/"//KM
PI?@?DGG]1#%0_)YK<S?>'#N:7ZD8]<B_%5#4."AE]P!%!P94@I:=08>UGRER\-OT
P0KR0>.LL%1&IZ$"$I<LQ)T6.@O-$, 41$_SEW<12(UOAFR<E"D&H@"V6AC%VI%TX
PE-+RV[\F.4BK,H,X8P+:R5[#30;17OJB8XL&]A^>YI?R/,W(G^RJ2UM@9ZP-\+GK
PCU/NZ]#P%8F2044%YY'M>;>%UE8 _9<21'GW(4JQ?"UM*'M,E)1#'K: ?1 @L6JE
PVXYJO4!>@1.@_E4FH++];9N%/P:7JL381C^0)"5Q+JMCF08*W-3TB>X>3PL"/7$>
PH-R3.:Z_"Y)!KAHOZFCU; O=M47P%G+O"FJIQC]@H?ZR=&;VXP4B_*(6;X2AF)E(
P5!5-%_@@A@.F;K7"2L5B.SO[S+]\CD*P]M54I)9FZ;(-+UO(BE:O*TAG7W<>9CT1
PA?^+YI&O]_>\Q8CYZNTJ2HP[S0\8N0WJE]<Z_BUGGH_(T;G[M+M.[+F[/K$ZO,Q>
PYA@3<D9XDT++GP7)"P]ZL\:_Q0>.:FD>LA\#>E98L"=$HD^CLN=.Z1"J=T<J["-&
P)Q\VWJX_;=B0KW(!36]]W$;0RN^[359\=0I*5OSV/A4K!CF[U@W4'?$_)G6-.&><
PX?K)(&/VC^9 K_[NF/\V]PEA6QQ[S<B12N41O^#D]33ZP5*)9P0>6(W#.X5KE*L1
P,I1!8@,J\&K@"22@;T8I\CS9*3D9;RB02V;_=9_U AL[$^@CJ Y&N0ZVEWG1W[Z(
PE,J-:/E.3FP[-AC_AY=E!)%1DPS+NHJ#3YVNXDB[:O__UTM,(*Z_WX^"0#*[1ON*
P%!S@-//$_'X^Z]^*$.HK!'IL:RBI;CK[,"LP08#^0R+<M'P^."+WF3H.W-T!K&78
P7!Y\<U9ANWJ[[S="AC[8:5M<*?I''9&F,W"*U6YF7$K8#:L2P15.O0<P.3!#PT>D
P(;A#$9<;UAR?MP69J3WTF53RZ)W$GFB/T(G^W,HR9O$"E%DL OU->,_;EI>#X,KJ
P)-+BI.=[:H)%0#: _-#2)TP!E=HU.V07#C)S$V0M[>I8C?#(0=A8?J%&8$JYTN[G
P#@C>4,\+[=0WXYK8:" C)$?/Z^938-(E:XR=G<8Y$Z_/?+*O:.A356Y2H%+^MU;-
P17=,W )"0A=Z$#2I_!N'I</T>_4^=,#[G9R(.,3,I$EW31C[[4N\<3[NLCK-)ZJ1
PU30.&7A>[^4!VSS+M.Y/_6G#SZ+*,^B^DDN@$:<Q#B1V!1J0U',+554SXR)C*YYU
PC#F:[/)'MX5YUJ@AEI)A-1)E)5BPIJF>HY[(?Q8F3+S&)&@XJ+I"9970E/1GXO_@
PF^! . &Q2//D)LRY\8(! %&G*_F//G *%JFHZY'ZTL$]4UH@!(</?CT=^V&;]'Y=
PN%%.J(HE&)QUF?W74_0%?JO#8\.:BUYRV=LPL#!S:L[G/\SK6IO130&5]W+A]![Z
P$9MA8'FNV8EN')TW"C[?6-#O'X(5]D?'ABX5/M=9LW%F "5LE(J\#,#M=P5#'8?_
P8HEH4#T= ?\\$?X3$X[M8FS(LBO&:3W:6WT5\KS1:&8X74O$%F=(PA<];Q(['9%3
P#=PC,;C?OG\BBR)X$'0_"ENH%:E)^@W%1"S5SBUEC.,USYL:A9MZDJ<U#YH$ 0A@
P27.XV),BIQ_15 P0U !0@&)N<&"-UI*8H!B)2%?A>]KYX'.+6,Q40J<OM)#\#+6(
PR97PS;)M]HD):(VCG_NMKKF!M;P"9/AI$.Z8JM_!6BZ(R?7:ZN585<=?VJ??M/*6
P'YS3P14EHLO\I?J=MJ+32;+X_V3HTWHN^'I1[V9?7FQ9IR\'!QNBX4TGX7-]M<7%
P_3<1/.E)S1?8/C&"M3_3B)38K?&@Q3Z5^YXG%,&!'UW-2CJ3]:8Y9,.(*]G[?T!A
P'^3XE\>!O<E5^5,KJ#W(<.4H57N:EYGW_^L<OJ,#1$@Y\;@ZB@AS]'_Y.!R.YI;Y
PKZ<@&PO;NHN73$_;L47<LQ@*C*+15$W6)&M'?[2U,9NHY-\PYC%2K]C4LF;K-9]^
P2A_Q0.D30: ZIP$^,N?QX%&/C<)8^A',#OZ9?C29+R=S\UT&3NC9SL@:D/4;[0I]
PHA9XMG &G5]C89:DOXXZ!4T!H F&,_V[-MK6:<3&76LSR_&X+.U0$JE+2YAR=W_A
PG5,D+B]?3AQR!<'=8+.G6/P;4E:%O#/SNP]AA1%][Q4X38+M1Q<53XJD31KH$(B5
PR?!XN=&RO@T/3:>-OA+9:]OWB>P(P?S+FUTZTN4Y@#T>*$"C&X)'&4SG>%^:O8RK
P[([A@;_UX!T[J+#-<>&K5[H0Z;31>SM7/;&;H+B \Q2A>IW-%S-.V .I*2LS[1Y'
PV\$//^*JDM8C3_(&%SE0T4%2DMX7FP_QZNANK1[CL\FB>?3$J;C6+")J*AL5#E%^
P?_Z..:17TO)9ZC\<G-0>N<;)VAC2NZ,WF4O5+(.U >K[A7J7,&X!2^SR5:1V]FH[
P30#>0%]<CSS1GDVDG'_P_"GAA[2T6/*N1_RZOAKGWBB($8DQ:I@EG%-I^.6([Q/3
P)D/QL%(\;?(VQZ!=[FA!#$&E<Y)'%+K[>( 8$GVOW2PGJ3H\#:G/^@$J;Q06#<!C
PA+OB1])^#\3:<./3=#"@GX1NY53,M<;_N(F7(TL,IZ@(XA1.VLN5" ^ [<^WSN.D
PFMQO8RBW8B;L,"KY&5N@HJ0%=TVH6% <(9'0Z0GIXHAX(1Z(]SPZ4+R=X9% _47,
PQ^L/@HH)#NU$,2&ZER%J#)@6:X8,E<OD",C#]NZXPW6_R!!Y:SO\HK$HM@8,E6@*
PS5# 5M:0!KR)R$J\.>E4PRZ-ZJ-\JYNBXTU^$H=*,$&^6N+OF8?$.@E3(IG?G?AC
PU%R^'B3!]"HZ.ZF8#WCN6Z*;V!]U\(0'_F.94SH1X4'6EMB#N:@QV_,(-1$;,% D
PEB;S2&16CP[DKN<$10P5?JY/%DO.GY57UA,IQ=.5P)FEG&ZZ6[8ULG*?Q;C:Z$=A
PW<*O9'?.;H,(W^E%'+ONZ7>P'KL7NFESO0W01%T[+?33:[RI!H +Z"C1"B9/A+>-
PO#W'MB8^"*^\Y8O UR5^TMIH7PR#MZH68WLIVX,T=XCC)&RNL(CE/;*$U-7834+@
P+#Y)]M*G'X](W_C!16H]E7/L#%%0\$!T@_;]U0)GU=\::>TL=&=$>(*%X"1D4-BJ
PBVEC6DFNF&C[I*'V;D3P6H<P(R(-E\I#T ,MDJW89/46I]3(W7VRWQQDT'+,.B:0
PZM7F-KW%BI:O-*B@/IW=!MNM%)+*<:B[)B7DD!VF12Q/QB4%3NRB31I!TMC.-MC(
PSU\R0#B"@L$:<=H4%KXCG!H<.B+GH;T\=SG=]!Y95C #:)QU EA@%R_?ID$!9WAW
P%:T%E8#BLL2JW@HTC5J9DEX(K%,K"/7WAFP)C,.MN-(/>,WJ$?/J(B[OH"$@7XZ#
P;8Z?/[, /591#QNOW2FQX)"[-CUZ+FU:3SB++D)@017,CC>/W/";DT?C/NV*TNC+
PJ->YH::DVZ.$Y^OP,<23PY(== TD%_12M$N+V,".D4$?O#X<+J&&E,0:8ZH_F[2"
PYQ,!+0C0SINLE:+ \]I3_.MA+9B_^?@YGE_!(.YQ%X,EC;3S:7^DB$4( !"VH,2_
PP&U>E?P#)JLKOOZFY]'#.E&5:NWY.FQ%J1\@%X^<8*WML^36U\TI8$-2PP=H$H &
P"[SZM'EK^5MWT0$7OMZMD88XM*(8B?Q0"[(0\[UZ9OR3T&0AI'0A')MPN__<GFTI
PBVL8LYWB?B4TX*)U86"L_EQD<\<)P !D*28H.]"FF.326XE9*]G>MA/"F"]1:!'&
P"^Y=$ ZSU77=WO04YL<O6*/Y036'9;[BC,I;D/395_65 @S2".X78_@0L:LST)K5
PDJ!&+J@5:SM=1E;^3L,W"T248P:VV0U'%#38YS51[EJR%S! I)UA]-V?W?<_W7=M
P<7XQ'[FYEH#Z-TII+;@8MJR[_.3IB0*$ZGO/:V]@TBXY!Z,9ZSJY2V9.)KC>4!A$
P@#]=T_H9..DBW=P%D1":BB)RF21A3!.BL7@A]I[&8>!)"F6-[!8=,&#^8<9T;*&!
PLSO<W3HD/,SKM):!$2K%^\[E#PW?+H;(<=XY8%<ZSUZ<W./43T=<SGVI\FDBOIM!
P)X,7X>*0Q$N&EK-I![Q0KF1]AUN 9K,RGKM#KXQ7K#L1T5@:?QDX" .EH#@X[-,X
P4O,H5Q459)U8U?[\ZFOG^Z"5=Y)Z04< GR+F>+-,VIR(.4A&%<%F9UJ#I*?1=PT<
P%=U7]2GX+")%SP!938G9+F52\9&E3\_EG2)PQ%OC.X*[):MM"!QYA-QER[&HR[>@
P$2))E'%R+\K/X8OD.6$!$366TW(S-'QFZ4W;0WZ1]MSKP-@R8D6.$A>W73(<$2 =
P'M]1^\WZ Z\[PCCYM^X4N1^-[#CZW1N.S=XEGT9V]((HWRLW%)JE+7IF>%YJGIL5
PG&M*87(Z)36".NQA_@65\SEO*G]KN43U1 PB(R#"/9W ZX^ZF4N)$>XWHQ_&%VW 
PDMTXTQ.B>3E;]9O7P='0;R(]!M0\9@':\QZ..L/U7S4<#^G1>S<- L! 7]H>G86J
PD?2SMKWUV?=^LT@PL"?X'R4%+@=?S%B&1\8:[^^IU5TP5]$"J!^:T"XXS:G12#DU
P)SH0-<<7(IMU .I-G-.PJ6>^[@ 05V[)R+@:O0F 4,)N_:**^MUAB]VD(M[VE/[G
PBJ4'[25SE0A)(@".68$@%,@44NK6+-"6E9DM( 3-(Y*B&(W/!^ZH-N6&]C+^(?XU
PSTZ0DXD[S*GNXW2\+ T2B[">(?R:%/XP;[$#,\KQ]?WF491",%=&!K]QQ]>Z]/_#
PT':!TEO"!.-"R\^!/*,M4$&I<'G\+^O(HM&S-X_W]S/3D:<RI'J;@1/D"Z+(_3.%
P2H6"3=^I5#/RP7I+,K>PZ5VT@O[7&JS.DQX*.&\=A7[ -HVOSL)EX72+[=NLG-$ 
P:IH?'PCCW$@WLKK38=S[3[9>$=W]4<(C]RMUI?/5\ "*/MK^&.=%Z:HBWA&V@0UK
PR<SYTBLJUG;]5NH/QX@=$']G, 3BF.)8_EG=C1X2HUWU<#(][8D"]LYXV%+#*'TC
PY%Z#PK>CJ1W&-H:;3_L_W%XXM6$#0E)+,'KAVM,K'=G_54Z#/'QJBA[QX-3*<1!>
P(JHU.L-)@\0#2199.9\'[Q'>T*#)<TE9B.];H>">4OW$N\*K]>3>K&[M1*4TT7V^
P.P#R5F4.)0'X56)8+X#S$F)'UFDQ/+<!-7_LPFRL4E4*M!31<$TTI)G ]:!\)OGR
P=!7<>L7ZRJ6&@E4&Y6L,.2=;_'6=?FZSYE"9BX/2LB4A E0N81KH=K=476L<3^K!
P9FA"ZYG\ZQPLO?52P,<ENLI9T$<.;FTA@CF=L83S,<((*',V<10>-)N8L\,JBR&'
PX*I7\4&YHY@9)]D>SBV 9SQ!TQEH58#W4OQ.MQ ?H&D$H^M*Z23AHO[8XK5-I#">
P"CZ**VINY^ 0SJ?ZWZX86\]N?-);[!N^+B-MUXZ3-0<1:S-DCS.1/$]JS1+7SJQ0
P32 2Z9]Q +&GG062KCG,DC):>KJXK./BX&K5#JC$V[(&C%14N$92,!F/EB5+0)KP
PY6+@2VW),H3]6_]WG450?$*V&]&@!5>W@T@S:^#R(2"^_>:EQ&VV>2$8VY;[!@U0
PQMH+_V&<2>,6%Z-T_'/O;0/73!]_HP]@HF<0IC%6!7HJETY2/ICA@_8Z-8!$D*Z+
P2ND+R4QZAY_P>H3.JN5^V0T4Q:^'RE^.-]?8BU?[Z 6M<O*6X#_Z5X0!RX':I,S_
P3' J%" ;4?#1WK2:![1:2DZIB7#:BBID;,[X64X,"VO.%+9[I>.I:J-K3'$'$Q;"
P'#X3.WDZK-XRYY1'&,K,XPV=8Q0T,F/9_E#-DE(33])\-5F.?=?7732)V%NS3'H&
P 9/0/#@G*"7\-6LOWJ=)<1UT!"C?V8P?T1=+R^Z=71Q^]/F2*/2R\<- ]K S'OTH
P$''*[BZ&S/UV<_D.'?])L:^N<K^R)S8OL)\X5QB:*;WU)GRC%/G345A@C +C'.)4
PS2-9 (F>1^<M9$R]B&WW:A]99=39QA0TXP?(!^,#?DVF?0SK37JV[>9:0C44>K_J
PP."-F3E<TES#K_:U."RADU;W][OHLFOP^'1;5!(Y-EPJSV_#%V#$T>^MW2AX7%0X
PA&@R_;>@0BT0(,BDL"%-WM]<2B8)F$%@.0GK%&582^!TB2D8)T'4_[G4PX'EM@^W
PD0?0EYT.O>2LO?K*6G;>=H&$Z!QK^Y(]C'<83I"PY""X5.$$I TK(PW6((.L?1&8
P6]48;]KW^L,JZEY5B?-2$6,84?=H]$\K2?\_90J)<BJ@NY">#_\]AK8PO]QC%_K4
PUYWLGSELJ";(QK52ORVX&RG2&W0].:Q)A6#+J][J?8>0H.+!H]=W9<58K#M5^VD8
P21XQ]9<KDJ<M%7G88^V2PU"8U9XFLFM$#R:Q$Z-FC(HR,*(TH#)*[LCSU-'JCF. 
PFX 5IJ%LTX?7M!9CFA\C;;6&1 Q^512'HH)G99VJSA0XIZH\!%QRON$NMFR8V4@0
P,[DM6[+OM63,98NB&$6*CLP6SQ0?4;[F(E^L]O(#2]12QVF7JF"HFW7 AVM,HT@2
P8XTIM\&B^;Q9\:'A$)2P:>R0B0[K0?%WL[KCSHD+5%F$\J,:<N"PR-$N?M<&2O(C
P"_2#N>/ <\Y+_?=(T@OO.M!XH,4O/8!1(K=9RY2U3=EG5%QS7#(RK/ BEF?"?DOT
P-90:>:FLLP(U\(R/"XD(S0VNA-R@4X7^V5?HLY#/_V]H4*[[W8GCSBF&Y"@6M89S
PMAV]O-92Y"S1##4!^[*+U\2<4@"=Z7B@OEG4M9H=+4*]=C$W4VO"/0SWOH[-.* -
P.9K/#)54]NWNV9121\36VS^R"'4(Y#S7U5GYBO^SS_N>GWHHYO\E%X#P*P./=R!Q
P6>[NWXWI-X#V-U%"@.JR:8=Y2XTJO8?8-M0+ZD6!W=O.>[@9<Q#0V,G2=FYJ,&P?
PBNT?,(;E9?&MY&_[=,5BR!I-R:?(B!=P<V''OBYIT$2),9\LYDX#//.1N2:D70-.
PPRIZW*Z[1C:R@82=GT/NOQE"1$]CP')N]G_-MORT;K#(N0Z&C[T>C7'MAK*%&ZZ\
PD\VW^>7/4(VO(YF<'-6V,Z+%B(J2\O/"[_9X- 9\V]L[DT5\'4-;"K>@)QJ0WG\Q
P!GEC4U@BMG&^,+BT=MLYC8AFQ](?QJ,^>(PGGE]U<L.P-G@G81.];8"<&'ZNQZQ/
PP)G^3 *H*,9W2 +DGL12I^"$-39F'B*LM(B:1@?"R@.TV8BL">4@1[[<6V1[,<%\
P]DXI-W^EF/FAUR2>AQ NB_>&!6=VZN&,-A&6U](6? T21=W)+ E*7FK8 WF2Y&+@
P017NS>X:#]I97;N&5_>W"#<HY-6G;%W._Z5@AB6!T,8/X!V(4(A3<!,>(V=G\=3H
P)WV>XG>%V%)AG'I*0\)%% ,R:#X.ECD.H\K4'>9%+$!01LA!6[378@!AOY:9Y':&
PM1(8K6=W:"?]R(\T>TJY1,XQ#K@)KF*A,TT3N4QT^%9O5E8LL7,)M_7N@!_6?R2O
PVS5MR<AS?'I3 Z293$9.Z+,A+E!^T,H/HW)%;B=3I:J]&N-;B-KC AF\QO72"#0:
P&>^NDS(DND:]R"5K0?47>DC!21Q@X 3RG[/BEZ4]I= J;-J)@PGL);E00#)E*QN;
POB:!^3K0DNW5:$)\0 ]VRV91'%L7,<I87'QGX39D8@6JGXB>N7W:+XCC?W;DGQ0)
PE6/>$Z)/?*RW! O/UTS>!9GJ$2>(]\<("C^M@#/V+IH$O%P)SN\7@;\\4(=*X0[J
PV/D%-6Z&1Q2;/DYE>6\VA4-;468D99@#]<2/\R$*58*[V*2$UGH.GG"MKN5Y<I_Q
PWN9T0: G5<SGG@B2%H@&P!U;;U4.N)M\SHG<3_T;J^;T)SXE'PF C[;#ZX(QFS6:
POG32N7Z(I9 >482E%!^/J^\@1O*H6^\@6"/:1X_U<T70/M6N9XKBB5%V-=VVZS1(
PRVC=::E@[9-@_AD).1)$":.Q[=T*/6BD!1!DH*)43YQABL-F7;-II)=*5Z#ZS .T
PQN)EYHX!QB!DG\[R;*AN=)$22 5&Y/W( %1Q-^D07CZ_+]O8\8^Z#7ZAJ@M?0QG+
PFT>DDV?(6I^K$S")2J!]C?E6KG,74'IN\XUM"8E1X;NWMT\@9890K &BPBZ5-V1_
P^SR%[';0V@'_@0.>9"U/Q<IFC0[?_ L'AO3$/-46LVX&W]9]+/U2^-_E5!CQ@+B+
PANC]U#<.R++]$IZ'R"F(?B\R%W&GR/1BH&)Z_F@4A!2K:[;5$EB!CETY)3"YQUZ!
PFZ<E0_4WCHR&N"B,.<72TT<YI_?8.MM<ZMHG:)IK>:TG6*R33>=U.ZN\5PN)JMBN
P6R&LF^<D,; ND]?<G!:%(I\C"_:-,+L$&,2]/Y"P09LT@=Z+F9&?< UOGR='78#2
PK8>"=%?/%(7:2(?-&8ZTIZIU]M)IPF"YE^4E7DQ+08STW9EP&G6WHLEY#/>SJT'*
POZ0'SQ-)8[=5*6:'F6!=;<]W?-B2/M9#6FB<,JA?L"Y:)H^I+NQMSK:#E6$1?]*!
P3C>5Y48Q;>FA5@]?M6!!O.A8ZBAP7/Z!LM+H)C-7%R@RFQ/\7<3.=HMR7V@&MC6+
P4Y+/:_A^\0OK!%;=?K95PL72?'7O8H_F3<^\QK,W]EH%H0<^GRUU=?)IVJ ;./0=
P6HD<YP[09T"!X:QR?X5'&"<7L_M))"Q:QS??"S^5N3*3$MKN 8V".ZZ[),;2YSQ%
P;O&6O([0JNT1!YF)MDE-&U9E$GP_*K3R+!T9JA[QA7TZW<#\H%+=&%9T@27CSHNM
PRU0G^SI>+.ZXY5(D7T3.PDR/N/'6^H]QD=7@5Z/?:P-=YNAGL=%O,$JN, ZL?M!@
P( @SVSENB0/WCT7#T0^[<8YBI JQ\-@=^I&%,=+L[$KQ<)<*IK@T-[U_96"R_Y(!
P/D'[27MB6'#F*=WK+/3 UB?3PXM-E?]/S2?OY-J\XW^ZOVZ#UQ0-01,-;>=A'!YJ
PEI7] >T#6M[V/$Z&%[>2P 03IWT2GO0A=<V7!3O@EO[O=_;_.) R8&4;D@Q8_;F<
P-LGM6L-7]GHPB6L==SY/GGZO!R<C35!.!=*_VW<A01:]V.B-JYJ3TM<QHGT7P>,!
P;47LAE8YS"*PDP!;?680-J&B$</!HC/8TPI^Q0" OIXI!\&?AHS]>9,[3X'1";O/
P,? 36>6'%M^S""Y0XUG9X1O&.B@$,#)^41G6B>7Q11I 4E^:=G]ZYDTX9>LNC=A1
POQ^=)D$C[X$:RMCB%_%'4<66Z*=])-"K8%$Y9VJPI*+=Q,<FAOV./'$&0-.&%KE6
P]DUX4XGLY; G+1#?@?4MK$( C.=68RD,"FR'Z1$E/W]*OEY;FJ?J8%,2FUOI6#3-
PB*-YM5R]([569*['S.SR< F1H$@G8?.F6>,9>^P>&@AOEU;=WD;^;&W%Y8;DPB <
PKF>NN67L)A\LQS]Z;LDK"EBLZ-Z&;9]X 4IM/O%;L%II ](T\HN[9"Q<M&AT/$3H
PH1RQ+V&6>DKH7%*A5>';Z2BEQ^_S0NNTS8OOS#:)X2?6VEK5^8Y(W6EW/PH8KT&5
PG,J**96#W)@K*)V>ZJ@#XCF3BM8;1KH+]=F7$ZJ%IPY!#Y8,Z/B\9O)ISN@J'OI 
P[DP6R:AF[35X:SY'-LF.5&XFL2F,$;UH(V7'S<*E4BK@=%LDD9[653_21\/'0KQ!
PT ;]RNIW=N#?2;VK=13ZW6#6021[2CLNR-Z(6T8PF=;WMW0KZ>67H(D]J&+?KW>V
P+BNY;G7J^X,X >>N/;&:M+]@0L"#U[)]+R$6Z=GSL@"PE@1L+GKW*@;G$NPH'R'H
P!YY4@B9:=<5*=&@E8%),R-]=5V2EO69_Z]6LT^9K5. O=@2F("AB1Y;N G7FX0[B
P/G2ZK9N6FR*QMCL=^ 6WT2Q +W;7_# >=%Z9G">)(!&U>T=2TY>9+]']^O!+[.6 
POU5C&):/'A$+]C>+VHCQ^^XW1EI9["FX(XL(1X=A<POMA(2OM'G)B10GJZ!\P6FI
P3QL4FII&96YH/A5S+3#\(;&Q")=6FT!_+66DZW=WB8?&[..-ZAJ8!XJJM+O_\DU#
PS\F?D]X A^P$P&QA*7!*<<VG!JRE"(-(X,<EO8'<G='[H4_I )DIW0,O[RQ=WWEG
PKT/UUVE6C@&2#^AGD:+5&</<:>:]NU!(*]HJE5B8,LS3&AEP"?:PR)0!3J.=_'FH
P%?Y(Q[_*^<)>N@N,+'\Z8T3VK+BE4>%AG(H-1\VY@&$,WJJ%(I5,FJ;.J5,%&AF1
PR*&V;RB=YR+([\5[I,_+2\^M/(9*004U-MX94HY'ZQ1=3$Y,9L97H/#7]%%J*DLP
P$!X+TWPA53BNUW,L&$K=F:ZG9D)N0\)CAG\Y2E1,1&IU [/<MM88T5@@-$]9!CD\
PPZS<6A^0@Y^CQ'C3'??RM2T"'$@AB-.^6,E"FGR.JG8%(FZID2MS+WQ"?O?/_(+ 
P(^5-SMR?RVNQ^6H%@W$D@YTCYP]8)GW5G5JC\IOP"$O8QQB#@O;SW/7(TF0XLS\N
PQ"A9 QOX;]E?W1%PQAEX_IT%: YABA=8]#J64DZ[BNI_MQ7S%]EOFT Q+GWFN;%>
P!QU5:J47]]F.N@-PJDIKF_TC#;#<@>+JSN2?-2- O@@D*82\S5M8#8NVP@OD>#[A
PZ@ZFE]_834 D.5<]V*UI0QGXW0_25V^&L98N?W:$@>K\62^?<Q?XY;BT!$S 4^SR
PQB"#-J9HNN^,)=8Y,KHN7%T\OLLF%*WZSV^P/AP=(P5U+:]/JC[J-(O?Q/,>*" ;
P!89%EN=9ZC)N,:X+L!"Q@<G]QWLF#!\!@],@[TA_WDZ;6FF>_*E&%I5M/S!(G7W9
P"@<*ZEQ<:T!3$NMEHUF5F73-TX,)F\">89;4 DHIT*4N &FE=3"\%/FVN1M &/CX
PY#=BN0YU!8[#"]'FZ<R#-47R-GDJ<'OY3E8P+T! ^:F[1]G(DOO(._>A]G84NQ[S
P_L-<\]1GJBM4@-U/7S\9XL@$)'>M'T,O/^]>I9NN>8N6"8G%D2;##PUB1U]NX"&[
PDP3.;JFPI>1'L_4"$;8@4H>G_]$V;OS4ZNSA,G?NT.$MO^QT$^Z25U96#)D+64KY
PKZXQ/^VVF9Y^@\=#]RN^*#Y$&%E:?C>1-,1OO%%G3$,9.WUFWJPP 63$ E,>X- 4
P+NUU5^)@U!% ,_0!-&#R2J&X8(T\ 4^J4'[B)]4/I7F#EQX0WSABW*\^I /"I@M/
P!#(O("E2;+N]-LH=%S#K[,<?SDSN-A0OV4LXP@=V'WEI<#,=>\G5QYBWW1A8AT?1
P?V)7GQ:G^#YJ&D:31',F3?WI<(.H@8>S@!IK,D!TNM;ZLI*"F$;UDEIY/G(64DY>
P(<%H]5<AY8;?Q&E'PLE+8LS[2O2RKH5E#AS\+0-1D8/1'[_6Z)R#W_YEO]'GBO[^
PTM)?H!:)BUYNT=USXU-+J<<@.A<!F97C]W9\)X)ZAL1_FO@@QR$.T>IQL[TIV\*4
PT5DVG^K:AVB!]U"I!>4>%HK\)+)JUB(:28O\[&X^ >JSE7I?YBGMZT?)@Q@NB+T?
PU-2\BN'G6X*2J[G.]W.K4G$P[,"-A$D 5$_2$>H5"#A'2E&?[;O4N[SDE6AA@XI6
PCW-A!F1J?[D#0]Z$W>Y&/P*[N&4789;XWM S$P^2+E1GF0;GL!2R<)%NF4HU36)5
P8H,8D,,!L$6;IU2R<! 8H5MO%.;3=VGG$T1;6@#\?'44Y/773NA[+FB?[QN3><D*
P?["S^($S%+<KI5>]>[ZLNM_ZGH7/@"+O5:8Y",Z$-H]:=V82C&#^N^$/,7J]Z:Y]
P=1YPDE(:2')NT!N\$&TW=H=S+*D=7F/1=<65=HDUV:_D/TRM'FTAA&A]($OK#YC4
P H'GD?S3B(E9U<AQ^-!BXQ\!=#0AE>6S:?(504CJNDC4M#D_ZZ8)],,P#AF_V;XG
PP*L+XM4^RO[2ZR?$%)3VK9=&(WH-EKV\?@L1J93/CP]*RKH^?^SL2Y.9WR?PF80.
P_BL(YA_VR"/6^]M"KV6T[' K(VAA2Q,?4NE:E>;-Q(1.9_5)L/G/LC3D:Q)W(?"G
PPD/1J0D+$H&<.7*=B0=HP%.4*A3(JZG[=%NE.%"'B#,?U!V4+GY-9MB&\*#(=2X%
PU#J,EB#I(*$,VCFNGF3!E&@]G>[?7$E4T>\DM[1?--K?U,7/CK_P#;-]Q"?;"$%J
PLU5IYKQP.@?L(6:&-ODTZC 2*/ [XT\J9+3VR7?<BE2\):WKK71'E^C?Y-"S.2RF
P)PB$H[]8ZF1!4'C1:(G6C([VT.UT"._ZF)A^:$(),_\!;3MXJ&I>V2*.#-P)^KPE
P3W2MK[\:8W8_:Q/<QWR7UN8TX/%>\E [)+R/5#$\A $:I8];<H%:!@XUV2<H.C<P
P!S>CS^R/;UK9O9^GCA'?JL<2=X15Q@),BHT _I*R92KI4G'(2UW";;X/;D8H3!:-
P)LO>.AH[P\J$B!#>\1U_C%9NI!'-NP@H!)B"A1'S$F2Z\%OD#<ZR3).CPM%]5QU#
P_%5_\UN(\01"MM;@/ 7N6.PJ J^A"K4AIR[-"=-E,-3@L7MP'!6QHY26$)WY7<K8
P: K/8@+,GDD<V<8DX;+%>J@I<$0)$^P?B]8F<U\H]N%WCL2OD]0$TWQ@?!)[0:H5
P;VGW?(GA3:J5QLX9-7$_8%/@AFT9Z6,QH06D['F_L="@NSF&&-MKU']::[CQ@\KP
P=TWLQ1_V:-D*';&I=BC2PZ\J.6/!SR#'69-\]SRMC]OZV.S\?'W>PP*!RQL5VUVI
PGUH0;R(.J/Y1"IP@G^G5+FVDYT?9C+RX;54ZON1&+=9Z'X3(\SHG7 )I)L9PEK]/
PKM ?&P??VA,< O* KL&;FX:Z#*-P29RK_N0IJ+>)008Y[[=HLD1U<DLB-5TD>=4.
P-TCQ3SDV"W9]"'9['3<8>_R:D.K!8 $!@BXD\<&3?C+W8!&5 /ECR*8(66] ':LF
PADACKFWR";W5))N_GOOQ%&%,!@8K4]#KU^^N1_<"JYJCM\HMJKA&5< $.#:08W./
P "27=9EEDFHAY>&)#WZF>HCGB3B<-,6[9&A"Y"I/):B8K.1-2^+9^MU$M[IIL.T]
P)9;^B!!X .&]'&#>S8BZNI= ,8<@7ONIT@^5-H:@SNBN,[V[7*48IM=LI@XTRZX?
P\":]3W';SR\$!'8$:M6)W$XB>+@#RR*@]X:(YUBH*0VQK#*MVC?/Q-5ZB98 6#E=
P3:)X.15HM3M#M^6DG;4=ZW$46/>C.F1P.ZR[5A_AD)1U#KKC%D@$RG8ZR&V?#>ZO
PQXK/R$:'*8^R(BAP11DESX#/_(WGAI/S6CGK0R:/%PXOL>OMA3+*,:%8G>+R>^2F
PYJ#F2XE* I,X)NG>J\K[R#U6P_6_MF:V9VI<<TF/+>M=X5PDSGL_XW2OA3BBF0]X
P9*'FI1*_9PN/02<.EM]_87U!*)#F0ZC?B>HVG:GD,DO!#Z6!RT(9\G#J 8P7# I.
P1=20<+9O;0JQ;P4LKG<;'6;IEFG?MO/1K_H@7&C)WW#-WOXA0EFPC(305:%@GZ/]
P.]V;1GL'Y;""F(!'F>/(@..K( =3,N6F:!QLH]T?D(>Y6OLG5P/SI/9_1YPF</>Y
P+A4?UVOU5BVL&>PI^K6YL'\AEU'Q?@KT;(V=NPOPN^B6A_P&7>#ODM-W)<*GAL<-
PA0CY^.T/!LWER LD#32'<[WZ7EBL=S4[@XGL,T&@_XYSE(,IPHQI5DMZG]?LF ;&
PA20BQ54,UE%P+BS7S_>-7:Y72R=+L[S+O3M)?NA8*ODA]Y_"J@%H8$6/[89>+E-#
PCP?C@L$3YG2[3AE*4D-0=X047:TJ-SPMD^LI=F":]1 F=]0%D3)+U#;HB+HR$A-T
P% 6G],HA&.R98K*E'#B^(1))WLQ.X**':+6'Z$\J7L[2ZO.KC!VGG)FIB\W[$KQJ
PM8I?2F\JW] E4[?\]OE<U :\S5-<D\'BYTD:.=Q@;Y'W0V2:6#3SN^ X2LE62B9E
P'ZU()22?>,7O=;+P*T%J%JY+#(8=EXA)5'TD=-<'C6*/2HE/DBH<]@ZG!2/5P,&2
P]SD/!.SV80QCNS^1\5;E\8SML2V#*?N:,-BUZCN,D#Q^-04[<ZM*^(Q6F]#KW;5<
P?%'"D<WE,@]0PIZ0E0>/]T,YU/ZM$.II6E(#9?0;WX,%,I/)D>77Y@EVD?\9KXY!
PZVZ'=W[;^;W6L77T(UMIOZR,F;9(@];*:7=3<X5(R):D1$K06&LT@"J"?56^82V)
P#(BE]]$-^>4B XZ3 'Q4)(Z'VVJ I;8$3)$C58A:TEK\8)1<?\!YE_C@4^NP0+31
P$$/J*JH3QJ#K-X](X!DFEP88C)ZR;KSOIJ$6T\Y^G 8J[^#DVM@008_-I)#= N,P
P(,B'"NHS/VT=[Q_9LJ4(#[T>"!POY*]G8T&;Y'.*9$-?^UK#Z6>\R'76[KB,:H<3
P^DKK+,UZH?1Q(V$C)OX2;4;*PVTH5%%Y[7X53XWNNA_W00$W54;;=VJ(>9>]=1UC
PRL09K];[J=$(8FICP.A42$5.N3#_5!V-LRR@JW@U]9FW0(]@$I$_ !KS+)(Z(A10
P=JB.0K.,R2;FLN(][HT:A+U,-<S3OH[3N%HH^[\SS*7_P5^=]L[SD@<[>0+>EP:=
P%2H1]%$Y,(.GH>7^YASZ1U/!!26-'"@<1)8Y#U!1U6@ XG#,#X_7]6]GKY*PE[?\
PH(N^"Z&JPY=N-:),"'F-JH8X/]$L.%H_6?$#HS!&29]+"=&MK1F"/!L0?R>2>9T:
P9<X$^B%#U44@:G@.'@0]52IQ3FERZ2&41V)V\O'HA<9.:8ENXK4==)H;5NKJ#V>O
POMR@T.!22#>X3WR=N0^$_KXJ&AC"Q]DV5% +N[P%+$07N\YIFF<_3H_O7$%&\D];
P82/ :%'5LHF-;5Q?8H>/KCH>!FI<<K"D:B@'6C=1-G2[9+SNF(D)N*>GHI:BI"2A
PNS\VV1:[FJ1W>[@K2\20822ZD<MK5:*E:H!7L7*'+_(@#PS(]H^P:4B0@(7]AH&W
PB#O)EFAZ4(.MEL 1K'#HI0N-083DA?S7,WSW$!VUQXK /MKZLE%'DF).2H3&3X=:
PJ$Z<7SX;*?N[LNOSW)/76+0H6%NI$^ZGZ=X-0J[?HA5],M:J?9'SL&"SH:*>IPM-
P;CP%Z"%D&RW:-&L;%PWC>"KI\\H\64V%;DQL!T:GJ?DA?O-OB<@P]1:Z]$-3^&JW
PP>SBJ2$U P2#8!$1 P6X5]3[2/=H0:" '!6![VU5!KHT>6L(H1TJF?443J813;=3
PG$N5H(5$V*W;P0;J%T.M>CP6>=](%-=ZH8FF?HSV;!R.=F5AQ>WR8HM^:1,NQ$0&
P7Z*[2B#O]&M3&^35BESO\@CPQ_."CXW0@MPQ&-Y( =6\.XW].<'G=F5SXIX ')Q2
PAUJ[P*'P[1CE>8-0*>6[^B>4-G>OD&_9W=IKLXFO$&,H\#X8[QOP\V/=7@>K9>F$
P3D36_; 6Z>3 @O7U+IT-+"P" ,KH2!Y$C32$"QE>;^31$IX,14>EI*:9<;!ACSGM
PX)!?W=F] /7;6E%C0SPQ*:/,".Y=:V@\1)SNJ,:S:?Z ?\;KS]NOEPJUX*W9]ACZ
P>>*C$WH" S_X=66JGAQN)2\^P&"X1PO*-JJ24[ :+6&6%P*N\9HE4-63Q$WH&6^3
P&);%#"N8J1H)(]ZLVJP=*IQRQ?;$J%/)<7A2\-,^AY+?7<@@.*$/6ET1S"Z1PE\P
P8JQ[=EC\5A?*S);>=QV><SUGIF?+R"'4F:#-K2&OXY#MLC/-C"@N[I[85_ADVJ(@
P*U/FOHT_HA,&?[)O7+@^;#OMR!V7\R,E1&D9TL-#!-:XT'9%=D ,HPH,O.=H8G7?
PLC32J+_VWRF%T\=*J->72+%D+5-\U>3<Y9:M;*IF0H'O"<8&U!7# V=[CQ D1R 8
P<]KAT%-2T*&PN,1G<N=]Y>L"E ^^,(.=S^7%IV_CHDU8"O2S'+ '\4"H5R'M[M@L
P9DB4]6^3ZR+VQ]B0>P/ +D'5[$RCWD=:1Y3Z)DTDB9.SZ6^'%[]6P,(R\"/,%K[F
P5M#W?5^?0.4W1A(% 0 <=6UHV!W8P!_+^'Y<)85"T=E4S:=C?3-@2?9J1,+<KW3_
P MBI7V'7P1"("J,EW9YM;7]HR;'>Y7"-5H+_L)FLF=<#7;MIX\$B8N/#AGIG($A8
P9P(N4#%[](*XDNHG:\=UQ#H-RPNTM6B[SKB6"'-+TO"+^1/F N0I_1</)KCLOGF>
P$4<Z2W0#H%Y=>?7*)TS;!U8+M1XC+&H2K0D 9QD0>-,O7\@*+3+QV<"NG/=Q<W-C
P2.+/:EF%(M/% .?7]-/BBROZ317/36 ,%3<CUDW<='K$\Y@#MJM>\\G^FXQI9V^(
P+KX+BWYD-'>^QT$'3EK<_B[IDZ.+DB+K!CF&RA,]3I09OK$:!- 6[I;QW<?G97-Z
PV=F,APN6<3-BV0ZFPJ-D_4]T,CKZ<3J$\#J1N3 1<?,\UPAC=NJ=R3K[;GT@MWYU
P'YCGVT*_' B0J6S\LXJ'F:"RV\FL]!UA!2NXK;&JKND4&,B@7'DI!&U>X!S4LHQ-
P3H*\!.#79)A_V\,T>EYTO4\A='YM^WDI_:T=X0M)0AHF#]#N<&EZ][G-)*_Q:==&
PDKRWH,=6;_.NLG.(8Q5>'M54^N^CQ)(QFVI37;2GCM/*023G&7"#P1S#55,>SE<6
P.;X._CLHAES7.):C,C?D=MZ-5W%,6WO>%MK.Y*5%2D67(Y^?=F4*J=)&V\V'"D;Q
P/"IS[ *7MT$AQG!2?EBL&9O0J[W$;I:I$0[XO2S7FDAF-E_BPXD][CUPH^'"@"V3
P7/_:W.E&39[?2Z_&@8C2Y.:JJ8N*?QF9:3:3Z_WT;"R7ILJ^1NBY:KY82I3M'2=K
P=M2Y2XNS]?A!EO"LT-C8=DC-50:TEONK-P[(9+@:#$3PJ9C3_2K2WA_TV@N!E)^3
P3HFIR-][/D3X'6]'Y^*1)>GFXU&$?!OZK><! :*9G> $)1B"%$=F\F2>=$NP5)TO
PGEXSE@9JU_MS!PRZP91Z>@]<:55NFSFJ_\L']92SK[ )L]2V&7)"#;%VQ2(^J8JE
P1YG_?,'RT^)&G,[SP(\1;U_5>?,)7M;;)BZFJT>;1O&1T(*^N9O0F$W"-^9_E87M
PGE)8D,(]L\V\>T09[^SX(>!/9RJ-H,@DV]SEX5.D>?5J6,R@;FP0:%4F]MM./;G0
P.M_F0*S%B!8W75I<@O.,M>PV[R)ZG955[CV)N.R]*EN:>P*\K@!7>VCE*5V'+J0P
PW?6%(9N.0NL&(1IOU/]R+BF@Q3P6D; .SEN$4]V)L.^;%$^[:'V7A2^24:"JNE#O
P2[Y5=^&GL[9K378I#?"-.82]@WDIEX8:PXF8-,-%)F=8MMQVP(ZZ5ZI_;Z5.=ER!
P@%K'7F[,BF(@G?(=[XHL/=G/]6]W 2KR^TT^V@D'#?W;:&$YIRQ[+H\<U!X ,H<0
P8V[U2!\7#Y@O"QLB#=PBRI*T3Z<\O_S(I*B"P6=/$ #DI@76CX&![;F09I!MJ*1T
P'_N1MOZM92PUX8C;UF2JT2[H$\^N0J^#\'V=]O6'NBTVZ/F,%LH,3+(>4-;6SFU+
PCS>NT:[?VJ_$5F9T!0PU7_S=916'2H/U0O'C5H2VD,KH>M9^G]MO*>)7_4VPG2\"
P*HLG\=!UJ@A:T;(,!L.A<_'NPS[Q#A[4$P@EXIV)54OE59+PS]J2M>\!AFC%C]=Z
P[SBXV6M38&GD, 3B/XQ8Z BPOO^3@&?^73A%(.I);9U2E8OO4(QL$EK)6=^>Q:+!
PEOT4")^K.-];AKNHR-&2ZW&W>.SAL[#DG/6C:A["4H@HU,#Z$V%K-'O]'W<!.<!S
P(DK2PQ.Z()#8(+,<)L3>LYL6>S;?-^IHY641C99.9W%,O#R&/CQ]4D9KIL65#14<
P#S//UWV%CY<(*!D\0U0L56B9$JT4&#JNVVVY1@[2:,(TM8@<5M^%(A_"0\SL-']?
P;UFQ3&F)+;R>.@&3T>J$\/TI(:G<%5UBOF;*B#]LUSOWWP6%@HHJX=@([SAU#-A^
PFL#;E+>A&2H6R (RHY?@)]%KR3#<[$3O77+ PQ()RU^[PF#4 \/>!I$ZK'VKYWI:
P(*CP\C"\V[C[VQB3W3Y6(BHXR8Z6%9ISH+&I;S9EUIX 7;B/*GXMC:CW09C5U3[@
P_"-==?4[2+]Q=A#S/M_K-M:1QZ'12^O?+7EUE+NI2T^/:,PSF,+5=07DBV?QQUW?
PKSJDYFO<ZNB(+1_HA]AN\,E"<I^ OKH-4H7K/'QHK\B0)3]?SW'@KX]Z;(9/IL$[
P(&H2@DUK^<GC>,UW.YT1U@\?S>$ ).X/!VOT.-;GS>P:*7,/'G^>/(NH9UPXJT)A
P L6W7EE.2@\J%.R9T'.:NP+(Y(WP5O!Q[Z_(9H?N+$!!=N2\&8 69"TU8]$%_9;L
P?5L]%-L$#% 2O4AG=R">42H*FVL79AZ3)I8Q+L.D@I%4'4XQ/<756,QW6\P$87%3
P^*<=1L_><FO.$Y.2+LMC[MDZM'[M'GG3OL4]&#R!:2TZK_X^@LH"W^N1"+_,FL3*
PLU/DUAXT,6+)2 -?=9(H'RJ R@:- TWM#;^.E_5UYKZ?&S$]#.W];L1#_=!U[)R/
PB"P2TS>;<I60B)^DQR O&VC\ M*CH><H.?C,K:_W>WBIF +P///TYZFN],*/87 *
PE"/HXM+V9F(VW](L5BGW11^E6GR]%4&)G.INQ)^ /!NN*E<E4J=0V:.'T\81D\+P
P"E(E]^NKL3$M5M],=;KGT)[;.(YK&AULEB!+1/$,5HB$W7M)$1/F591P8W; 1,R?
P#1F\KS-4"$>5I@2:A+O6^I!>WT%80,*,95.W8_J5HZ9TG%R0$$%CL:E^:CUE2.,5
P(&LKQ0(_>4(STOIO7L*Y61F#OWH4C:E_ <F)#-.;4L+(AO]ZT9NL:A[\2E">Q>H6
P[DZS[>A#!;LT6-/CM;ULS/+L1(1-R9OIFB!J/7+42*H ]>!MM\VS]-B?-+(JD-]8
P3;AH)SIOY)*UD_A:)@@Z1!\K 5=?[0&I2F4PSC3P)/E]EF2IR2M/&_L'L?R>)Q8A
PASOC]"R.'S^3"Q^F#QS:X.'T_SC$DDPPK"*G^?F$K3J.1<TZD>2M[G:/5[,G:UU>
P..XN$7@4QY<<L]I'CV$NGU\YC7!/XU?_D/M2,C]K\3JP2%Q"^#/D)XHR(-Q7ZKD0
P$TL%[[B51_-G)T/@&D,"J_3:MZ$:(.<;$2QK,#*?"8=?3#PHNX84;K[Y&7R$!CA3
P7LT%G.&Y<G^VNP)9#.B+^H(I(^?<;&B3M?! ^ ?U GO%5]O<!FTH-=!<E*P7 2N\
PGFGAL;9FN%R3[KU3%COHVMHDU['6T-BCBOV&C#!/<O"ZEMV4Q$_KM2H'F$FG[?:@
P_[C3EC;*<IQBRU9(Z9@E8J=BK#G\T=.L^\3IS(9-&_)F78_N4?J1%"X_?\L=]-5+
P"'A'D-^4!(SDX0?ZKY.A=5HJ&@31-M)Y^?(3([JQ8;*U/!]:CCG!HJ<_Y,6MS!N:
PPF'5GOJC:?3]_!B;'.1[0?+6_9WH<2=>(3"?UK",0+=*O&)!#&Z+9VCW>QY09[N!
P6^6>7,O:$,: *^-/5";Q(?^6IK$TKNWELED*/WWV_:6 06D?5 #"RVC% EP'!H]0
P@/F $#+%U[%<=M'XFJ(76 3/STA)Q(::N"/2'"'Y8;<TC7:KW+F>F8^$]D3!74\=
PV)XK?@9A_J_W5:-CRO22S!:V0C<$SB5#==N/J#&?>**9?8B/IPMBB+*!5GCSP'^H
PRS6<XE&@D@%7B#R#JN>JB$\/+0)2UO#GQ<TPS5)A<ITC%6@J-6BA/ H[J.46//P%
P[%N,!M.J3S%TDQ*V+4@*22G(*2=V5SPAZE;^A)0Q_/(RYWOGX71%9A/M@^8>D35^
PZT.;$YD\+FE.2#GV#J[U<URUJRM,_+TVGJK5U^U\?XPL/:,00RV0]@MFFQ@G.MT8
PL7[*@6!T0^D]\_N"&[SF 49DQZ:SM0]0&I("0LCK &J/FK"T,!#:\8/X\,Z%_=GB
P\-N* Z0J]8#8\EITH/?Y\9=[A922$C@MLW=C.6C*/L,E+$1X]#OLST@-$<#\!C-)
P-,3MMYTFE;)HE!+!AAL^<.!\"GI5Z7[?=0X?R50:"/Y__HG ERVC#SK?^36(_UZW
POU _H_BP?Q*SEL C@$NH5L>#3"*S I_ AK9]7!L?&4S:(PM?U]R@-'(!LBC Y?;S
P;VOO\LFCP4%>*K_FH\:[;-_CJSRE/2 2FH,KUR4$5#Z&]Q,ZE9]ADRJQ'5?3$WB.
PS[B"AZ>6P'*/0Q@'_Z90WV*\2.H,@OD0F4_[,]#,=.L OB K%GI/.H1W]L<,AI1'
P<O-5L>&[N7R9JSN^_K:M(4":5M] R6!-,_I]$U$]$Q+?+2R^(RS2UQG%"=7'A\'+
PP.\+]!1!85("U3D*.LZPCNZG5GT@C*>!HX2+WSJ&CS3-:YVKDJW3"(U1Y6_L+7_5
P/G5E!=T>3M!GI/N;D K5U:FOJ9-':$LP8YLXM-;E5(@%L7@ZL6C^852UFAHN0=(Y
P NLEV?)[)>.SD=%V"&&'$BJMX!P$3$B/N6=9(HUP@!<LEP"S?PU*+NRU!4;J,!+3
PRM@.!0P&[ [P6@/K3_(J17&F8?")&* "Y4;"RB:S1>> B6R.T7,NB?8^)W_POV%M
PXP<4AK((GJ9C)>@"3;KO]YP5M,)YF$.034W->PX^N$9W1^W',>']RA[('AS76F60
PZ6QFQ6?T$=3/[#7?CF7RB3+#EM$@M>L::57I[8L];+XWM;<C5 M;?(<>X_Q/O_#Z
PS;*1/KL/[:ZR>N?ZLQ7?LH<T>7"3NRZR\F^'*48/SDLG*SG_*7$F<ZDEVC,E(MW[
P"QFUXQR,%,_ JFS6=A1"Z@;UYJ]B##=[$\E&B#*:S)\._=*)D'D=[6EOKE)7&', 
PHO1*HNFK2NP0U/B.63G[#>"17Z5[H_@#QW,(7#'?7FTPT$H>:".U^0VV][@F/R[Z
P>SN=WL6,=[;7E?&Q]PZQ4$B+EG:*B:6%&G1^_EB_05X0:EB"$;#6AR.&A$P: 0E/
PWR(V&+2R6U;1U^1/4&?);QI^%.6;Y3+G?COPGJ0[6-4)KZ2P,#F]A[W>(3]GAA"\
PBBY,\%LQZO<$<O4.WSH)R,24JL[HDS.1#XKRS\@%]]8U?+3SM8=QZD#B+ W4K^1Y
PRQ]+81I78BV=<V6T+>$+XHZ@@"?8.XG961=J01\=3NI9><4W_>0KK\<H<M_/8'@D
P&N!P"* P=\TC_8EO455X)/_\LD'LZV6Y&W5[:O#QDI4DMUZ9PP!=B2?S%@BATG)M
PQ=V^/S MB4U":1C83^ZZO;LU2J;4!+ LQ(#T3;5F9%G;1+33Y&2O $@1,.DXX+&J
PI*?L>;0C 9X/@:S\,+HR.Q9+R=3?ED%JI<AQR/3!3 -6V(2G?;T?BK[N77D&7%:Y
P< #L^R#L %TYT,59TPFCTNU^+JLJX=2;K#EZK^DHTEM+9%^$2)V/H*1S$8KIUJ=X
PR5@8?0-U\5Y18.PU60[NEM.01,+1UTO*0$-ST?, N= ?8-BQ&QQ-P><V\NAJ)&V=
P8!AY-V3:5Y>L0WW3B-TV9>1O-&J@MK5RBXPYET9TZ4YNY5C$%--(L,I&EIT51DA0
PO*NKI[Z*GNYV&5[ 4=KTI'S,4_@9UM'J*5Q;U=C:E&E#WK"<KO7'8I[^EZF.*VLD
P@"RJS3B5T->F0H2U>S QTX?U"P[*_>G=DJV2=YDE6/DMVV[3\L<OF&2/&OTF-J>Y
PKGA2RVJ%'1#%B!X'SCE8]RSXWBA'K80D-YOAIT<H*75FH:@(M88WY8Y3@.]4]NLQ
PH]8A@,R#]7Z2K/TC-"X9MLH4^^X"5P&]"= \G<T<<.\G!>KOD0%7,+'.F[TV,V%E
PG.1W7B#N39J\3D]'_QNF3AVU'POOM77G)U00HH$71[G6$U$4$V<'.-6/9_MU'%69
P;.;X&Z[9A;17XO$S+_WZRX?T_P'1%:WXNQ0BE93D!\%#D+9<&-K\?^V>AC6@Q!3Z
P/5\RG3[+2U5K%D8%M=F$8M1JI U/W?_IL9N8P\CD"3O79X9*CFO#36-#S[2$1@_Z
PF<XN9=HNF3U5_VNC_ENP X/C!,8#YPU0@$,"\$"*NX('2G<H)RQMC M2LIO-C=""
PI<N98^H[A2Z\D"&$*?A1 \#*DY\TO-+?/[+F#C]WH?2S8G*E3"UUC!E&S6TGB'!.
PR"-!82!1PLBV^#@>XXP?$8$L94:Y5X=WI5HDQ>5F-IBX:'Y^H,3,$/\9A%^,I"XV
P86TQT+E^Y27_ KPW'>  )"2]-%K$,C0@0MA]+1 O%&$X$Z[KDC^!Y3[6I$NX1QV0
PD+1MA*-&H=4>$U[D&>C!/)C;Z><XPJC#P.=R)9NKLHVG<^;:RAC:Z'6W7,.[A%G)
PZH,>I&Q)9_[BB\-S297E1VN+;@A3'4Q^61'#)<[WV!^#9KV"<1E;@K<B&PO!#(YT
P7[*F(V8M'3ML.%IDLC\D2H2=&[$=&_5_)1IF!.Y4> V5-M^*7DX0G]/7@:TGZB"V
P0F<NK-(@KN*(Y<"PT!X*R,0QBTXX\*<**X[=ISO7"%FN8[7NT]1,E3@T20?ZDU!U
PVS!1MG%_AS?0<1RFVE.5A\LA[\K05^<5O%*Q2<008:C'5ZO_OVN$=VK/K90JT?<Y
PN [',7VA1NFO/SNE+[*QO;&A&4^<09N2I:F^@7S/O6ZZ]>K:CW,A<6 \?8EL/Z]/
P7I\UST&%)NV OI< 6#C1OU3'R!-.=)<B)LU7;6C.6^ZR8>=A$@'1@/#;78KDGSX<
P;]3VUGMV-2FO&W8%[T^:_"D#T?J#6)C-0F**^:HW I :K)Y=G;D/NV7X@AIP]@_&
P'C_8K3JXJB0L</;=+7_DA5;N@0LI^4S('R@,[ L*AU"X/=@2E[U10TD;#G+Y6*.R
PN)N (O=K% D]H!&&>E8\#MCB"7489X>'XX!,F;>L=NXVOX;OH86TJ.-VH"Q]?9%.
PB188BMKJSH.2!R>%, #4J5ET(_*L(TAI-4C$Z/WE^; K0/ECG1:9TGO7;R0Y3FC"
PU:O-#.)]]Y,^PDS%*[^ 8M<51*?5T,?SP*$ONIX//X3L3+C'$KQOHCY9$0H^KGD]
P#%BI$PU#M:"F2(8;*;7O!HO/85X>=ZE=FD"\F[KJY1=>P0P1698$MOQVE>T=ERH[
PW_Z )[7O5)?8JZJTN$#9M):V77+?4X4"*HP >@%A:G<"/0H38)H0]H-1S)B)48_E
P CT==$ID@>SXMX,4K>VK0,R=-4??_&]JV2^1E+? T-P4(+T$G7]WVM*4DXS\0*(,
P**/V":1(F1YQSSX2EC)#1;I"G<*?<1/+]'P'@<H4;[(8Z%EU<!8/H?7,) 4Y>&Q3
P0PA=C?4ZI$)3P[CLTT\L\L,J<N?K52AG=D4*0+IJT*?I$K0@&X7>=0O#N>36RFM 
P^H@$BW*3,3$K<J2Q6*6SE&Z">4,+:I'(L)_)NMG1''2Z?<?:*BY=_L3,^1$!N WG
P@C@@KE#U9F9VL)VOJ:&+DS:$-JDBF+I9+;1O[NSPN6&%T?R%;$K7\R%"0$KD\39 
P$'*F1G? 7%X^&<ZE9?6;F*2E9+C!6YIO/0BS-8.7"71[0]7F=,ZCGLKFE6U+Z]MQ
P%Q-:;U[OR1)GRI<1U0W-K_ID2E]:\7Y-K#@H,X5Q[6ZRPA+!MQ,Y'\'[GAKH2$J+
PZXY[I6N<AC(Y!M4EHC>/MB6*PS;]+"GU05I#Q]MC?4J;';:IOO,A$3)!EW@_^[XW
P-%X!IIK6GDTX%L?"*$R4%I.TU.URS'+B4]]*-&<F83G9 =F; ^C X<M/1\F]\>KZ
P!%YB4V]6V+R:=>G+LL"R 6E154UPL>48>AB3U)D%221(J"(%W7-!^>QJ) N0*>U2
P>=(?;G,@D9.1.L,2J"%M.<DMDXKA&ERI>-?A7%T5TX_I,""XIT4#]$_9MH0]EO,[
P%C)OQ_P9&B7V HM9))G4IF9(JA, 3AJ18030]E</Q$U^\8I*SW4Q<6*+&ILY>+XS
PM>?;?:VW7EZ<R!MC%B+X>)QEDV(S,J;9)QC'(NO'[\[1]@L9,SH7>0>D>GT%[,'7
P&OKHV H2K9U0M+S "'?1+<!1"J'-Y,3C(^3H_6YVR/LAW)%!$((L;.S_I)7BZ#1-
P-[I40B,6G?7I?4YC!]:8H*F^$),E 4^%?YY(TT6,2XXLWCAI"S,3SN;PH[))1X U
P!8M3LM$#>D$D5ZV?7<4LA1ZWD*L_S8-RGOGGF05M+$ST0)[&:]3AM_R;YO9;N_HY
P>T6H4P>/M&SJ14 !TZ>FMD^KSAB0(^S]&OTMPZ2_B5VOK.]0)_0D;.*!T=[2(L>0
P@55 [U[U@=6:\Q:L;I0^_H]P7:3RZ+VH%:?S@(EOB&1<]P@3(LA5A'0=R*9$SN,;
PD($H0]M?H>0$B&?]GIZL&?OX!*@.E='&3JG(NH1(BP?[UXV-.,)+"Q^*:??P$=7.
P>7:H'3J4Y1KR1?6["K2<Q>?;%&F30=T'L?7*%#S-([W=P[0%D\[SJ/_;B0%6/ -B
P8UR8NUF_P$SCZR'+J:WBE@JTQ@WIQ"!S3,9WQ:BL-XRDJ6 03FEZW2X$-DA#L'F/
P-&3*GOIM\S11D@KI0"C/F:C68 %9OJWTK+4.T$2=[3FM'E!JCS8!4='KM\*UO[)1
PO^U<RR='[-29P.W$ZMA_)%6\ECF+,P4=5^H)'%!1W/P2RW4DTPWG,$2Z;&+\-1@<
P=&@V0'H 7LK>N>=D(9"GP-9P8;LFB=NYST/H+%AH'Q!8BB, ]NI.,.!=)69:&(HC
PR85LR'.Z^DYPP;J9??#;/:RW=\P/IPSY>M)@<$\3)0$<"NUPKAUC7OE",%./@6'(
PF&SV+8^VZ_E<_ "8>H;81V?'U-^+Z3@C_AS5#-%HH?D?0"1@'2VI1>6;,#-&QY !
P\R4(M.F8.P!Y)7R[:5..;G'EYI K9(8;@"Z>I+-]HO%7NIDMXZSR*J!KE+V*J V5
P%!4ZKV5Q?4$-SC[,-N+)5VRU:P=@RIAG3E GQ/3Z'FM,_- @,H!!#@[M!Y7  HZE
PBK@-++-_<]20H0%Y?#V_H/P49J= G;X4'T+%3GARXO??*_F3TP1/D7/_^T>4JK)J
P63CH3Q>19585FX4OK<Q4#)(D8:HE$6H#FY;+BR9-+)*FE!P,2FY1!B$+1@!Q!BL_
P&PVU$Z3GU,3;;&=_<':Q@W#UYN_/8#-F@O?W)OA$^*16W@D 8]6/CJ,E9EK%XID3
P DVJQ?*?Z<P-<;U&'")U'QXC$&,!&J@CZ_D@7+X,)X7>7D_#Q0\L//<AR\GO#J3'
PX%_I3;(L,2L(K408(O35S=N-CPHU.-'U[677?1'!_,88)'&SF"Z\<D GR5@'H8;O
P2]Z@/F,UV3UEY*8,")P*U/>=#P;QNC@#!;LKIHX=VW0>8+9W#8*TQ(7[;#MHY5M:
P"0HSH%,%\K5UF&V(P.&#\:MA<2Y@L4IN'FZ?T^)F$$:C4_(;E&X*['2E0L:IM6U;
P2Q,>EL02/Y)EQ)!2!1D=..KY&4EZBYAB3>=JJXM;99\-E*>PD?<:8W<"5X)=SA76
PI^VVB$0AH@BHZ,E<[>;6A>\H6W?!S02>(3;?Z.@(N7.B(G%^SAL="F(+)?X_ F5F
P;2($4W+$Q.\@_K'7>9KPT=%&R+"JYCHH'_7,KB":%.&MI4US=58P\HM-(;!>.214
P&3K9-:3I75YY,3$XUY[!F)['-XSW\2"$' ^GZ_M$*?^+Q.^[?9U.OBG[:R,C):GL
P:_."N^L9:#AR( +\24+@'DO-C.8VTY6<VU#8XA<YH2A&R0%F!HV9_)BNA&64,(5E
PSG?RA7PFMOG:4]\Q*C!HEV06/GDAJ.X2S*94[N2C[HG=Y:7B>K?0=&@$G@P7RX^'
P7<I9\;/&61$=S?1LLOTP<SW'D)A61^25Q%1 Z5:CY!IFV7O8V?#.@V73YJ7"VWPM
P_N(H13*#@PVTM[RGHMPWB9;8W'PCE>04%=92\EI,@(H-:@^9,%YG2DA4Z@*W?FY/
PH#R*].U0.P3N#O6ZPB[Y#; ^G)6[6L;B-@F4,^4)&A+8'7^$5E).[(%M7RZ8!&)A
P^O>AVJ /&6H&IO+>H)SO)C_*3^UHN!=1L>L]/F0-HL(JS-4U!*P4]OS6&@6'=L)\
PQIX.:LX\_&KM'G=,KXHQ&NV P>OO.>/A.*JSGL^$#,*_*$_"I]<AM=,1B+)Q_X!3
P".CSO"@"K],S>_*&Q,%6"!FI'D[Q\FG9&>:.=3SXC0+RR,.LK-?\,=D?K"!3:5JV
PO"E(O=R2TZ=?@OO!7?P^,&A7Q_)<SC;-?6$RSCQ "+7][CS)8@@-!@C<5L'"=8,*
P*;6_!@M-IE$B_O\J*3=$>Z0<RANY936&/Q6?7\5;G#9#:TN+\GI)7\7</<6:\@,[
P7\"&7%A2; M*"X+B78AOK'0VD7[24"^.;)28;ALMY6Q.<.Y&0-Y[&&C1'('EV1*,
PVW9%1@R=SZ6#F"V"07-)?\9 EZ<-_)"XO@ \B=18#$@D:2"^9L8ZH"EC_',PJP E
P\R-MV)K7H GR4M_!VDE2+2?,<&'?'Z$N]*\#FMO3?ODNA2  T2='.#9Z(+C4 47$
P*JYI*G,W8S>$" RB1.VBK]2'[@9(4LA)C\D?G'<.$<58QT']G@P/R.A3#1YJL=$B
PM>9,7GYQ045**C2;.$E9N8/@*%H>LST3G<AZS%Z$=HY!Y3=JTF.,P.9^E_/!NTL7
P<S'E87<0=NWT54ML3T[]BG!3<\>QLCRO5:+JHW !D&K KY'DJO=W=NI41E>>\#!M
P8T1\7^\$.=890O:/7M]>78ZA/VD!=YO2,.4E'QA9BA5;<%^OEUEXOB51TVF<LUGO
P,<3_D3B 7F'=GV-43H6J#R"AEE*[HFA% KSI;4I0BB>_X59\F.S,!=PD<)R.22+/
PD'+W</F%B !*Q_@/7N/_VNR83?1(<6R^>QN;0S3>@42S_8[MK\<9L3 +AT6Q"7QM
PS]JU]>4BA!$JDE$>3<[=CH-U<4,DV<WFG*L3JX9%HZ,D=#[QC*C$?F02@) ;?/D)
PI'X;@(Q9MR3J!OPZBP2@L'=(".>&[RHAW:5/S*EONN),K]V,MH^$J;<4AI.0!X%C
P9'4.M5P^P!:AG54@CQ4*OT;I0'Z@=..'S<]JI5_OPB[8ZDN/C9QKKA^U@</=70KL
P80$/JJ<A<6.:R(&AK-9[<*[PVXD&F+4R7.TMU"#Z2W<?7%Z.2]W 2VIBVL;BV;2'
P W[AC,\TC/-"*]C/BTREWW8,_3#-\O,EKX)JVX3S(X8$R02=*:'V;U]!]+>6X4B7
PI%E>[;7^C$+"\LG1S*#:? WHX)[.51:1QH"V=IJ2! %E.^ES-Z;.UJL>:?IQ$[SA
PGS2=MR)F6+ARL NQ56&#PW^#GB.RI+%5W*>%7^?GW59U#F7?-'RA^,Y88.RP^5+O
PS95NMJ8E^0T^?)P]?OZ1KF1MU_AB(%5GA6]-CMD@G[ ;FQ#N*C=_.\W5@*;/FY%=
PK^MMBGM1BQ'3A8.EFL[F-D7A.'I__=1#T(+0K\X1V"OADJ"@YQOO5%?Y-;\J=,<]
P17!5 ]DK.:6(RSMO.48SP=5HZ_@H8@WB[:$"1F KH?4^/>>?_)@$,$W^G2<8\<4&
P"3$K'SXW_AA6<^V7'>[^,\V[2>>_+$$1+<!:/-7>5/!_FAI4D?0@+GU:C8CGMPGM
P4\&3<U6;NGK6S\N1+_05?](+24B&@:^MTO)D5="(A",'QG(G(/%*K/6^6Z+E+,J3
P"C)4J")\NLT\[U+0I5N95'^UG@6G_UK':32'(3-HY;^34Y#Z]#K527Z\L="S1R5*
PK<-1@6R/(]7K"12\]07AS@E>]7/OC&(IHD@D1H,DM2HE_B2=T**#"2+G"&6TV%J>
PC1UQ0P#?-PZ0^B-:2[\CE((C8$#JA8BE#^*HJ$>>RP<DOJ%Q2PNAK-_5-:[3VM./
P'>Z&N6@87$\5FZ#M:S#E4P3,XMR_2MO?'>H=E4_I2'J,K_>F^F9,T5/4K9R^E#J 
PSAWOPKNL)Y::>4[V-,X#V E?\"Y1:%$P#C#SW7 DO2">%=H?4*AS'IC@T*U/2RP5
PT;]2I/!Y8%(_DC6@Y3O<\">*Z6^6"WQ#RI5@RZ!14=HOY\!(5BG$H?G1R5]8F]U:
P;U !IB]Q.=+CWK#\['#I<' *LJ6#$[35,W96LU*0C GZVJG=:!9U+0-$+*=?;.WR
P<8ZJ4.LWZ/_$)$K(KD7*J/0@A:E^)@L!+@O'7+O^USQ5NW5;7N;CY'B[B2AMM^XM
P1K2R'E8]!B,#KR_[$N;3^YJI$;R[_=\U=L]+IL$*\"U?Y=N_RF2(>5Z#BKQQFW_G
P$,N^UANJE#S.JHZ$O;6MA_N20%<C^0ZX38AR2[Q2K&8<AAEO!=%_UB-+I9#4_T+W
P_4SFW6ID9UDTJCP=1!\"UF#ZQ_V4#$4]/["ULP)+-@0_T8[!<8-7Y_8$YN?&4E(#
P(E(I*78&_<E-0?A=:YU1G\-H^)M((,2C[E(=2 <N &1=,5BJT0JGVPEU0-@I)/K'
PGCBV+ [<+(T6'I5 I\P7LF"ZC0ZHG02[3_.&_K28PT="PKW1WR_@1" BMI-X6)!A
P'@6H/H[]XKA]><<!*^TY&_?+%\GT[X"8 M*A(\-/S58I8U[W4&#1":$G3_UJEN6Q
P.]KU!57 ?Z5D520B(S-GQT-E-VG2/L*H#[$W5R42_#'&S(VX<5.)\\U),HD<2PEB
P;MRF-TCBITX49(<SC\UXWAF,(O:W +8)K0M_%U> SHY_Z#/.;FT(#^$L0QW[U5(1
P 6?KR=RQM@(#;_I=9I?<+L[ ]D7M6!]TY(J$E]<*_#\0NMC*RF],\,#A$&XVY(7 
P'D)>J,ILX .KVGX62M$".(WMD)@V0_^G(LR@/&73U$.W,NPR$E%%-)A5$E7ET3'1
P^L[QMR%"\X\]8%FQ<QG7-.S+_L+*G],89W00K$,;A\HEK3?9T%JO+N)YX]FITC E
PNK3*)@SM)W]^U72S&GNA+^92NF%2F.JMMF0XN$5!S;$-R(*"R=,C-[:\-7/*!@RH
P*YIL!OP6FP9A<9OMY:OU_]U(QFON^A4R'4,XBEIBXD=!*)*%IU[ %X#?ZQMBM50'
P+\T*/B34[E4)_@> 6YYB^=VN/G-^Y3.48VAIC"&C8M9M+H8ZJ,0K).0_/PXWC/1B
PM/\AL@#=WDP"J ?NLKF@YL"?A>X_=2]:0F)S2:WH02V@<R)4[:^(:0?Z0_@5JN-G
PR$%XS-S]\X!/'!QXQCT0>G832<](A+YIYL&^89MZ).G$C!XYS]-B.&7>*#[.;.C<
P4Z5 O%HVO@-H?(!YH9OJSHZ4JB@TR7:4D4\/I09QE,FY7IJ^*D5$$>])GE%YX*A+
P(N)U=O,/UF=:>D8'-/O00'PD*'"6^FQT&5.*N.N^<^H5FYL)$P%$WW92N&?E*<-:
P N3?P9!0TC3]G'0(0&_;^^Q4FH5)%TJ1_Z1_^J(>)(KRR"W:YF#7,B%G8AUTD%O.
P+]QRQST1%EZ])'QBH7QR2N&K=YXD*Y>G,4<*)@<4P0ZA_?CSJM^()E<$U@9B*VW2
P)W*?O?2?#337%*<@ZZ0*NL #<;RG'CPGUZ>F3:KS<\("4BB^#R'.$23H>313X* ^
P$^%XY,"@3XWOX=&2RG>%"'EAO/)E@LO_(9]?JD/2,FZ=1I=FU:P*<"=WA47];#=C
PUE# UQ1&\&,T5\DDNHV-Z$SG*X@0KFQ&:6P=/\O\++U;^,IU'?[!N)] 1PFD]/H\
PB1QD[)D]2Z 9Y8WE[S_(.M@!5;RWEHHMHU5:)(T@N.'M/E*KX>G__E79CUI*'/4N
PRAZ NS[A2KZ_)R>+/:$M-.:$^TGAN[:GZ?81S=:8MJN/A]X/W!*H]DV5?*Q(+>%6
P[BW3*JLPX]<?B1;SX:=JMY>(CH52$1=+@<&D//_>0IGS!!QL4@*0 !6N;\,.JI> 
P677Q1L_D"<!KB#U3R;='#F0&*J%TG 8\V=3CFXL)MFPSP<!PG_/6>5@_N'\0?J3L
P7[HB4(  1/] J(<F/VOQW\</UHM.DXFJ#/?N"9>6[+++/0F6VU(C!59 -CS=[2O4
P6-[^_5 ]"; #R/)?: O)'B\@XRO@"QMN,'2;CT'G]QI-SVJG?<NH6_N.#2M;!XSV
P ]1D5 U&H2,&Q*D!#50(*D@4+QB;B'LA:SU1@!%3(U[.UN[2[WY+MVFA?U+F> =)
PK[]I:>KV^P:HY(1"FP6R/9^2AVJ,G0O']C?'IO(U_H(M#:)A_IL1<%3/VF5Y)H=L
P84A?N$_9YK;FX;Z(CQR.@+\2-\;/QJG?C\]_[V37G@+DI1#AXAN_8Z;I/?NM53]H
PER6^L$*,-ST%5\#.GD(92JQZ'GJ*7DRX38T UB2;I3[Q=0.=[SVUH_<FR^]V^S&!
PI;!VE8?(&,]<]\ZB.D3D_Q/, -2[DO]2L22B3Y$'AE4@3<.K?"N.1<9V. B'D&JO
P$$(MRXAMEPK81-."B-[H2BII8>VIVL;N[]PO&C?6DWW3:B'C[]Q6?[#UR+?9-!LU
P_T;Z/1*ZVWI\Q^150$\D(\^3;ON5VE5I-%++!Y:R065I24;S*SW$*/K;"1]4(0,#
P59#-OAFC&IRIIB'PK& 1B;XK#PE# )>?8A^$3C<S7\@>HJ)*QE.XA1IZF@/!U%Y)
P567ZR!U67L<-^WI3R0N=%^+T&.NQM18^1.</A>A2_;+$L>N;)&>KRC/H$51KC>2!
P[$_;14>$O-S-C$TSHSY*9!U4Z->M^0'EV*]%3)C ?VX+M%NT&_8P_J\;!1J6/Y/,
P:$#3U7]\0#_474,J:7^WF,)D'8H!G D>X\7/&:UNM?]JWQVT!2\T(NX=%#@SS_J>
PEG#];UFAXWV[[YO;KD>Z+2DWA8[+_Q7'OQS@@K\-4K]HMI9B;@'\8^ZI3])6I:U\
PDN5V5&3X]%/H,J)\H,&*V/F$4P/E[Q]"F#\B5WP-2R'XU\R.KVT4HVCGLT<<2'>4
P]6PAH0'C'$V)I&Z\Z^%GZO^0%'^>;NTJ[+]CP(E8F'5(&ZA^W:4=LAU=9@6/J#$+
P5!==/> SE#V_75O3SVXJ$'^[V$_NE7%6?RW?Q<$3#44;GJ$TNKO.3;U;]_O,Y07X
P[E07+:)Y,%CLE%-XD2]:8%HX;UVR\!MOHAINPKQHODK,+$D12$O1AXQFC>J>&B9;
P$G88R<1JCU0,+C_=B>;<\"C&N1S?4S^;E/(V-,&;)C?ISO7%8Q<41^-2-CDP4J9'
PR406[HE&0,PZB54"41IT!P3!+XH-:1!7=R;1:X/Y;BW#YQ.]]J4K[MI%4=> ?_.^
P?H\64G&%N13TO7%"8\H0=@OJ=GYT#(/XB-%CM3L^/=C?3CX'92<W!-E.VTVF'*>%
P1RONSCUY)<:"1;3\"4NYMGU^$C_P<2GB702/Z[N6,Y D+I?/AL($Y1<-[&W>Z%9/
PK](C_PZ1SW] N^*]Z:F7FCR"NZ48W-N\Q%FUX\<K$K9[Z;#8R!@,([YUKVA1<$/H
PS ;4--27[8?J"/SV7.MR48\6*!5V89?,@2H9!.X/OT5N,Q0Q(YM<9/QPHKIWQ;=G
P:R^\R!#5X<<**"Q\UP@I/XSI/ZK6!J@(TK6!3V 8S%<.3I&OG+(&7A\H9(LKV2()
PYW+CX1A? +FUQHLGFO&^GU8^K _5_?R[ZT9.X].ZAD8>SH0TP IUQDM9Y],SP,LB
PYXI$@LBBALP@B:T@$Y"R*I@'#XNR4A3)Y$ 58T@_>V*.C*-Q!%^T(4$*QMN'RU*9
PW1\ NKF(;^>"__#J*2!TO'N6LP;H/M?X^]?W3!:U)=V2^%H,T3[>0&MW>N[-T6A-
P'1LP;(PW W7159>!4CISC^/''GPK%YGL9ZN^4[SYR57)3/WCGZ3Q;,57/-9P#TQ$
P":XWT OZ6/62 ;)?5$.\-%@O>.X?+Y0 DZ-#&[\!I>!ROXA[6$R$\OX0TSJ].A/ 
P? 5N!99DH2WY@9,&3Q&!Y@9HNI,.G![D#D)F<:49M^%UJ.R$=(FX&1'@"*'^IL G
P#U>G#PM!&QA:LI(-#*F72B(I<%CL1XR;V.4Y,0]!Q8N#H3+4(P(EAZ!%J\U% .D%
PE W'(+DY571).CI]"UXFWZZS?OFGB6SYK*S,J/S>H5VQ!5\G4HS>^]TV(S>..GAJ
P<RV!#="=91\<#[YE1_$W^J9B@U'>^20P@LEN2CE3P7.2Q\'/A;_QB4RU9NV_*(2>
P4 A59OJ3<LLH1-]L/8XZ@802=1Y:G#ST,[EY *ER@_+A]+EG&[.U4H.54]Q;S[<^
P)O50[^R =A[*\DV:J\36FE>(&6TW/+IKA\OK+;%E?D9'L\-BG)YLWE ",S423I,X
P^AKWY.M ;F>U5=B83J6XM"<]U8PB+EF_/G\6?7F9MEFK'? %\Q9TP]11[HT5*3[R
P,HGT=JE60HD7'5?6L:JL2(9OF_QD-VN$;DP*!XPB]<D4@<=EM3B&K?I>Z_Q@BEEK
P/C3T$&HFAG+[LL]LSK$@A7XXS7Z8^'5DF9/\+N3IQP!X;P; ]7FU'*,604<6$I2W
P1*AO@:P(GMLGC9>\CO+O=-&\?)M?MY+!Z#6G1?RQ"O_YCLRUA<-B'*-:50P:S7<X
PB<+Q-<GSSGN5G0U B5L<,AU)L)=N(\F:FFR+7Y^[WTC485(Y*BL")K"SJ9'2QZ[+
PQK-^7DG(3WLX$F(P\T[E5P,S!>"FHP4?2-[MK:1!'(GBP(V')K DJN(+^W!T87C@
PI"7D82>$%$8>8G^&P8618&K&DPTK"1KJP?N"M0BZJRY6[M"%U#3)J-5C[VQ:Q-?R
PT0@'P+L/=N%$ZQ7-XA=94TX!*' "$QY+9>/"J]I$C.]2XKO!!R+N#*E\L?Y S)+Q
P/J,@S4+,V MGG^(-2,U<VP'/6N/'=WN07DTIM41[8H22$,FPZLQNA!> ?F4Y5#FC
PL,=/D7"&YQYQRV"*NX^(5B*L_0>X1+%7N(C^?N/LH%3BJ[JP>K!/O3VCVC2D9SAR
P/SA=U7?'/P74N34*NZ,3KAOEY\6U.M9%LWXR:F1!P+1$.V6_(.FKDK\<'%>@[U@^
P-OM>;;FKHZ;^D8H!Y!%623-=F3IM667V4H2_P3=GS!G,WPKT,R^O7#7'XV?)B-DU
P&6BR+ Q&5T$#.V;S<?C15=P3R%4[D_ER!BU_P-5FL]6UZJ4U#UBZ\*^@T]-R .S'
P8JK\@?0'NE+1;JX=1BIG'$$9QQ0GVQ+D*.:<ZIB9[+?#H<8O,Y;9H[ ]0Y5$A=$2
PB%8]XC>4"/LI_FZ9UI<X0^:[9&Y]]>?<N"-<R>NV>\(PI=F@SP?@\>SILF#X=?J=
P5^^0T2H.I )O*MXVXD(O%H5AN*MR8308[P(5'+@AYI4Z>^/QA _/\L#UC)/2"8(9
PQ#=XCFI"\$(#ST,MK_?0A9W;L(!OO4]XW?C#^]%=^5<U5O-(A&W>QF>6(R<MDELD
P=L^9>C)97H&\ .&E%F :4U!0>GN2<@-D#M=T:WK5AS]$G-A_X1^9##,9G&CK1&_5
P G2)A]3/0#W'!")K@)Z_/NJ]T!;-3S1"'*C&O4'O2ZD,!B7>=UG>.BO[M>WR"= O
PI:7D<Z.VLU6-9C><O5P%#/8Z3\$X_BNPAR4%12M$I6XEDT&N<3 P@6F 2;;2]C.#
P.\&%IMS[70ROX&6WWAS?KSFOA!$O3HH!X>%OQAT27SW 4P8-JZ;<!/&-E?D$>&$Q
P(#M0EFJ?L $^AKWX1SBXWOV@%@ABQ,ECN#)#%UVM6A']-1.TIEVJZ9$.$V:.-R.Z
PKBG&>#)OO3X'!/LB#A0<"X QC-&-E+<K?/ALJH;#E9Q187(J",L/2U]EQIW4/G3V
P&<0JY&I&M&6$9HL#&-_-!94WSF880UEX*T204[02^\<*DT 7N"ZL'KQ(85:AW.#L
PA'W)=_TJ1S]7WXP/ZIC;.)?C7.BAH%\H.RX2#4J9[:Y@FCN_BB^)@J#UF#KLBDK)
P^EVV?0^FKUGE(&% 'K8M8KBWU\!9<TMK)&[(&PMVHM.5O;;0C8@]JF!Y$\2U4JP1
P\>NO6^?-DJ^E9(( [0,*QJV_QOZGGXJ#8A0EAW]P*F C#G?TO?K9Q2AKKP;F*9D7
P-+_\\" 3A6E:[V[6<G =["&!/K JJ7;&57(VC?E79FR10#K&"_M3#4'2<36T)'K2
PLQF08'JPZ=:WS8IMI.AL(SV?H$*H@NN#,</O^1<F27'JBC=*@ZP:J)[OF4=+"\S.
P5?6T^@?3)Z][6"RNCD\D"WPQ#-P/0Z27S'_D@;5[J2FT+T[2_KOFT<?4WN;8:#73
PC<4::UD+/G)9P5D^$XA"KC"Z>5'$NXZV_6V8T6J$9;G:7K\S!UJ8)$RTI%T$4TJ1
PWD(F0]GDTF VC1]/\$5EEB@:TEF)]J.8=P9@=15@SWH\X10XB4AR)?XS;]=9SNFA
PI]3(2WQ).BZ)$,<\;""/P0M9ENA3MW4C/O=RR\Z7@V]>_PS4C5-:17,F97&MSUQ/
P2>8]([_\*1QY$"=^0G:F7"OT#1<R9WU%L^?7 #[[07X:1;MXJIUWX>A4LOFPWD3R
P)_#+FPY]CE;0B%S;.Z\F_2J0/P+7OY.-,H]+SY@0L!>DB?V2R!"F<S<M5CTF(__F
P4@+6C&<@:N"D_TT/G(,"%<&78$JZAI]((IJU!SWC?GWT73\Q00;:.MN<K"<&^2^0
P3FU=307S5Q[$"99/QO")DPG7+H:$@OV!@"83J 0JT@VA;51'3WS@SP!/N0T?,NJ(
PSF(]&Z%+HP>4203!TH?XD=4!Z#BI>X%0%FT3 9^V+7N13;!U["(*H_F)TR'&EVR*
PW(,<#2""I.6_)64SC:=K=Z(S@*%H$J".Z %S+RA4V^AR\M<^OF!%1RG!F^V0_7+3
PK$V(:N,+7^3#KA,-05L?<'@1:0UWS]]!WCEUBD>5MO'W[F022>#9_W':M(,60U"#
PI@I:6I"Y,XL[P21/_+OHUEYTV#24R,V%+)E2PZHTP]9T)6Z@"9G^Z-F,0U;*LHA6
P@ZA2U4]R'H>4XI:UQX3;38%H@)/LP$G>ZI9_37# D$S?E)E8<LI1;V4GT6_#1/*?
PZM=G0SAF^9?>K?\)YN<+$L#9T<I._#<);P>7/1;2Y=]UX7P:>/V#W4V;,"3NE^Z%
P&/P_EY^$.JPC>I]!5!@282$<(+9I]="1#)I3%$O;+K DL5P&?TC(+_GZO>91/!.;
PD>M-R&"_("#T Z?O<1H+VART_#=2,C97]L@<PWT+R#T> ].&Z^ZF36\.L'*D^X]C
PO6*".K:JJ#=#S?472QW=?P<(H PIXI&;X8Z]$T,(^#.617NPM'A<D2$0,H*S7 YQ
PEV+Z)[AH98"/@?&AU@MOKI\%.@?+O$4)F!$@F#KZ0/I27Y7WJ8ZB;0J:%-$N83N%
P73=I!DA70F9.A,=>V_UX..?HG?N[R$#=<2_]/LK&84/O@EU!&6E7=SH\CAE5T)QR
PS*BPJX!LI&MA^)^AVMVXO5*";;9MK)4&C'#%CH)PC=X?AT'.;FLPBJ(-N .,%R3G
P*W$MO%!6%Q-Q%V2%/1=L#]C=0XZF]GK--O.O)-8CCJC&NND3+P-4Q=C'KXKC'$-Y
PKH<%:F-\B9!*9:(L,2[D$2G=T/"LMSXAI*/EAI+NUJ@:(_I<K6B'?0GROPR/Q;_L
P^!=L\S]BON?QX:2KU-(X9I"JYA2^(,M'RUY=, NWMQ;S[&T',^<9?;QMN"\!7$[T
P80OG5I/<STAC@;A#'506U2'\EH"Z_YK74[63:[EXLV=WYR%_LIEJTO5JIN)#J_9!
PHSDD^N/*Z*MRJ3+;QLL])7']6#0-M*0[3T-J4 D['3\JE)M2ZI)T6+@G(:R49?YA
PQ^@<[6U]1(9'E(!3'>S?L37VAP$$5%^7P\5EY861SXJJ([LA$-7%;#,N=LE,IDZ5
P_'/[><JXI."L%&QHQ?[/6"-L6==%R^^4"J_L4NL)#<_2WC?EG89?S%K73YR:"D"4
P8*W9IP46/%7EIG=.$-A8YL]P,->*BN_0'=0A@JN A,A_?9<L[6#>5EWJ.>7,PE5F
P>  5P\X7!D](D.UUK CV+#15;$L7#,L?XWA<H%I68%WP4H@'$:TZJ$:5T?V.UF((
P1J\4 -5BYDD :!3\A^U)@YN1H1()]_!ZL]-'BE&N!>H>/I&W:,C09:2>B2D$-=\[
P_"Q+S./>'6JP$:FC>[ [&C2>ND;*IIY$CV:U0T;JY!S5[ 5[_(>3B*:)?'%;^>?W
PT!/H.G)G3"N92\65GE6#_KP:YM>Z#F5IWBW#[\>K,S'C)GL*(O\YY%9WX/:G@8;$
PW7S34>V!A)<+VS';X@C%3E/I6X+$Y,]>ZTU0BC#"^_PJDG26Q72C<I31)7O;M?MK
P!GM)0H\J(<..'J2DCG?F\?%KV,6WHLH6RSDB$=\8'H _+#!%O#")NLZ+F#89<+K'
PT*:PP-K/_V"WK-S8DBQ4Y)=(RQ.G;:BXMLT?$L E&P/6>IE^,@DRWC '*B.X1$VC
P5ETAP"CV/!,_=WA'7(5C^].D=:I*ZK@@:9J:2DEU,"BO[FP1@\JUZ"[="K(4ICU0
PN8=MX<>BT_MV8M7XW:TZ1;OZE&6!)!* 8)'</2C+[]4(  19F_)>T\J2<4LSE[KL
PN\D&U6L*XVZ"M/&9VK8Z&]WR-_* +J\/4HN%,>Q)>[%>U.DZ[1&:TX-H6M:+N=:\
PFT"VJ^L:+*CZ6MY=\A<WB>Z0A.-@V,C0:0HSJ<)LN@/\1ZQ^$=B-$BW?/5L8)4D5
PP8]J6M(5C6,:*=]OT5GFCBJ5U"J@%.^Y!MT;NE(J< YEB=0Y!3LRX\A%W-4GM*FO
PK^ $&C 6]TMS]7/J+!.N1N%/MSZ7"0M:Y]W4QT:N,L=X92EEP6AHR/B8]R1A"Z[3
P6!#M@;.7TYG;*Q6!,HL<PWY:X8\/)X*Z4.F%IA=(]65"?G523;:LLN+47E*JOA]V
PN"EW0Y+ZTZ(197G;:=OM4F&.WC96LZ:P=->\ N_%-4K+A(@I*'(L4/3*Z!2E->B=
P7SX>:7^-TY'I*J/#"[Y6=>W.F2Q[%H*2VSO/C9'4!;KUW2:29T=CAW5V963FV."F
PC_K(>^I]QH1M2"@IZ*>F*.ZXI/U(1X"@;684^VKA(IIP(2Y-\0+X QI..#$P\T2(
P ?Y\H2/J+&%L)T'$J_4A0IF!8;&3@)C\%(P5Z%?]&D053/@?WV)%;VSO\=&/Z ?$
PA=\D[)9.BP<M7]YVA[XT:JC5>"Z;2DN)8]=S%&P%IVGRCMIOJ>=X0G>PT"TP%8%#
P2[\?9(1#3SR(,]PEK\SM'?.1>I!J,M!<RV")=]I6V5:KWSSLB.GL[O7&R?2#52.C
P,CKN;&^(]M4M.13*%(V)HN%NVS7KQ\2V1R'$C..4;"9[E=31.XV>?67$)1&PS?S:
P2&,E\:T0"CSBH?[#H L\9'QT](GOT@$IEC>OL5:]RO51)N+TO#B:-;<)2V:X* P4
P>.ICXA"H^C,*'-1NAJDP1?QL1(>V>CR[TY..<5S _(1]\.Z\QHM(P"*N-8:2':(H
PEH9-_DAQ@4NS2AVRR;,Q-@>@KBL4>U@%%IECU'Q+CT'_@N?R7"_! 0?$2VIQ)HZR
P/;39W+&:P.&6BIH>03B@@4Z%@\DO"";&TL9\'"7X,'^@@PG9KJI"W.:'80ZSK*&_
P#J5/YI%9<W8$2EJ2+'E#MM7%&:U%IJ!E&:OUL$/3=Y7?I30-HU""0.9G0?*,35>W
P&A:'EDN&7';&J1EHEZWIWU7BM-_51*%^U1FIPO)V\0O&T;Z3MK['BK+J"/2_HA=<
P.#!B[@J,K=>HQ,GQ5B7+68C)X%;M$,4RQQ3]$N\0YBC]YB1F>(=4_.4$2+3.IO6E
PBF'_=\[IF!B>$XS*T!DZ2B(JP-%!A#RO0G@^KXOB^(NM\S2QJ9.-G'Y/<_K17!+'
P$G"M_83 ;"Z.JA2%@A."L?([86"YDWH[Y)='@<;,HMH1G5IRRPD7PNDQW]\!U/R3
P4A")O^&3SJ!/J$?$3UW*X* XP[>+9ATR3YZ;:12KIGK117]/K@KS2-&J6+:BI!. 
PS8BC$F:Z\K:W[WF3/?I2#LFP)NDO.Z#WM$FA>FH3;GDS&485DUD9SJH))+;X+L7/
P\*3.DZSUYMTWC?"9-W44*RJ]2+9]#AP^U&E2/AM7&T7VT*LJA?TDU;WG/5U "N8G
PE&A,P9C7WEJ1DX=KY:C;/X[?1R3;(G7\6QGQ$(O_9TK#R/"0]& )(ZNHNTE>AL.-
PV$>8JTP.FG>>OFSY8W4L6R==U7JJ[SO$L3!@F2?;^5&_FCRC17L&W,%-MSHRH4JL
P8VE%YK^=;?6>8)1==E_!@SI3*/CO90MT+82U1)0,C#S!GL3;/&[;AB+":J>I<%"Z
P,;2S9S[0PMT4*(5/JL?7^$FBAH-8!(]/&)?[2-T!QZ4XK0Q30!MN2 I($4FVK*MB
PY5.T8.F?@*J\LYYA:@Q5:D5,LL8]VUI7@Z>X7WKBG/P&^E(\W5R]P $J.VP\H !M
PM] /B510OJZY!2I$N6*2!DBE9CY=L+MS$,<J><3(/L+G3/>D R:D.7T<L([1\9WP
P@\MP<G_!JAZCF-V.M%-]SLSD:;+B%QF%'5SHERF_5E7F)NGY^WXCN4C%\V-_X%VJ
P'(37[@SB:OIEP7) ZI<-:%J[8YGHCM+?4P$-E4;,O(P C[S[211LP#];SS109D>#
PO6HB)M!A@J1Q-*ZX.<O[>BIW5DN%Q?B0[D<E*R_+@T"["O^)^W#_[ ->A+&Q'!.*
P;;S.P9V1?](]^!S/44=;#"K88LLFDIRM,.OK@&PXS(T,R3/<_DPD&_,_N_#8U@2>
PV[CWJ%.*0Z?1&"">H*)!SO_902P\ICJH-KQW -*BD6XP#C;7!E[$S-D@K=3.KI2\
PS\_>G(RS%W38H85XIR\G^XI[):#F$:&L8A'6H._%-Y'*BC3TNIX'OLT02%)S^Q'0
PASISWXR30IE$(M=R$NI3"&:W/:]F!!PL]26WJ;Z^L3@%!B(.3T#!2]F62'#$$]WS
PE]\(>X#_XM5*>L,ZS&*29Y0VJ[QB[N;.$V5/.5OOLF;()O:?F38,II381%67@3E+
P>*LX#RI0D 8597X[!+Z??.23.. #'=:W9PNX2&V#[FP.I(%:G9.03I9ZK#_]R_MN
P%\&6]%Y'XM/UODXL"$?RH+!(98E#$J8'2+ZEDB_R.-/=:J@:/*NT-!8&<612_&5.
P-F^MG&9ETM<!8$F((8JS"K7]E3?LA#GX?=24"5%'OWGV4=,(Q.SALIO0')BP[Q![
P%&7789@T/>4J[6D\\)&:9FN1%\'=23ZTIKM*;)+'-958T< /Q$GK/OL2$&O'A!9H
P\6J/\L21%=K=&U0(EO$<^5/E(!%OK]6<\ ICF$3+=M['IP%LYS^=/S:>WM-^-,PJ
P34>5Q,@!"ZESP?G$KJ:MC^S0DM> ?ZP !>WZ0B_.E]AWHXS&E;N=*T!D3]GV7VH=
P5+QC9/LJ4WGGYT_Q@T2+@:9$JJK@YWP6^X 8.CQ09@YMG1=/-S.\;/R/4+V^T&8N
P,3=%UIA!9<)\H;RPJ3H!)L"+:=<1[IWT@U,9BR?#]C3%63[=NEJ"=U&KX SC#'XZ
P1#H)DY;LWSI#;M7QT.AMF;PO-3)'E 56>4 [N6V"!>R'HRE14[>RU)Q6 6*,FYNZ
P\UI,QSV#[5TE'1RG+UK;D^(PZ"9\S85$YK?EDQ-_&@]0B'5KA[]%KKUAY"]:?ELC
P@-(4'EBKCZPM3$PN&@>,\B Z>?&16=,QN_&Q-S'*KA+SP 5&[2ZEI68&U.1.)[:Y
PK!/!UV- D$,T[B46!@]">#C:$C=XM$%>^PUQ1P=F6"KIRJ8(0M'2:K2]2JOI_(IH
PU9TIL%)=MP]$V"[LJJ;F>QV8VGR\H98PC-5A[DOG'$W-*!P::G-G")*DL,ZC&^C?
P3;BWJ,Z]A.G-.P]Y&I65K[Y\6@'MXPU4I)\$6%4V@!O8OFDV-)N&=K[H':[C1PK6
P1<RUJ5%1R?TKNJ"VA]X*7BDO&?K8JK9L3MC!)-=?J6\B#.4R*)+_VQF'ESN9=*L=
P@3,ZN60YFK.5!/N\8@]R@R%0L5BQYU ZM<>@6-0\&-(DC45Y9EK#8YB OJK^]?WQ
P,TZ_*X1#289TJOR-J#87<\H_ 6B;26,G@59%#IT#MP/@ $AC,V5S_B.O"_I]KX<&
P)7ORB!P0D >%P..I[@S*MG.E-#GX*VLNIK$/V\T8^6 >2('0W$O2PE.?)L-S4U8H
PS!6FH&HG8/.JQI<6P,9V"\5DT^([*)[Y@V^]@A*])=]00-[\=9;#((2,H</VN8$ 
P108H'UW11YXKK04!WI<@NJSVP?'5$AO])3;$(0G.>0/DV:MAD_"YDJEUO7?H!YB#
PQC!8)F1VY]MA/F,$ZK@*C/MYBR&*O02F(\^,1 5F39T>@H=BXF>I>W8B/0.">$QW
PCQ0[A  O7KKB^H@^+,9;5C^[:%&J<OV@!]2O&N4M46VQG[S2V]]H#&<*F\)BV' )
P?SD_5C.@]):R>8VH![L:OWG?2CE:CQ$,BM9%.]+YK75"\QC]@>91,AM;4,8(4Q#4
P9\_21H!S(\;6KC>SO'OE.G0?$"%\%%A(#D![_1^XSCE+4[/H;'+D*;&&9]#:[=R.
PQU5=^G>V6<'GG(2:PGQARI(6[TZH5YXC0?^=\V_R&&8.'3T,#7CQ3[+1O^_)L1GJ
PN9O>[:H&YNGFR7O*($PQ]U3#F6UOD@$ ,<BPT.8!M_+KZ%8,WJ[ W,LZG)6;B' 0
P:&1E]"2+K;+C[)/@5S]P[)C'EDADJ$^-/Q850NHN][H49.= >='LW;J!4"06-G"F
P6(P1I<)]-[JA/00_Z<5^A /0TKHMLM3^*Y2C^T$\M3ER8JHO6U*%0H#9.'\L2',3
PNU(45=II,^3OVK2Z!M#A2MX(=D@'FGO\FO)_@]HGCH,XB05]RY\]NT1X>U?'!Y<8
P=(<]&01(VE"VVU1Q#7).'^HVRH]6/T??UI3S%!E5%J;#>)+T+,^OZ.TIV:NVOOK[
P1BH;]4;Q;6$CX/FVBVOISJ#OS"N*L<1$"4,RC>NBU1O?M,#-SUC\+@:DDD>RE$F>
PU!T*'K^L+9)>6TB/Z A)F./[F6C$SHL( N8[/@3,;Z:47^6-)+EON.09!?EQE@BY
P1ZQ?Q_ &Y- R-YS8U(RF$H.B9Z/6<'^_A++SP5D#DBFK=8A6O;N.<#Q!"JC+*Q>'
P:MQEXMDP?M8AU.RW,@CQ]K% OY>M"A3R7IVMEW ,N_:03C_+TW$*(8S(1AFFD_N8
PG9SRXY_(_Q)Y*G<K[^.'UF%%%=AL\5QQ"TZ=<I#N  F%;\=-2:H[U<V.'<\3D%Q8
P9U2L]!OJML/IA(34:BV^7 \B@SUG7KR!" 1:'BI0@9QL2JQ#Z'<&#L_,H;L^D^H'
PN]E*R^,-P$/NP$IJ<IB=U8H#@A*-',W)A. U6][6J_#HX81<CP95Q)*_.!KY_DIS
P,;>6G_;\OO$LX..:<HX=Q6;8YSZ93()NY"?. .$J/%:*[VR%P8J6(JUG0*6A(?HW
P\;@9'[7=W/+>A*XU3IG^&F2<7J\K:0.T<;H65RQ3;I(TCZKNJ!%O+0B"2I1Y TL&
P3O\5-R2Q*(=@9P"#^?K-D05D&%SZ?"7F6 SF;Z@V':[/NZ<KY'L:>NCN_N2I_..>
P?NK@HGW2N!T7_,&F;@&BE8('/8S ,G?E.B]E5 VL1A-H6#_R)^L&EPOY+;S/5($L
P0L.Y:&-)ZL6B'3$TCR$(UYT2&?2)O=6'<>C5#KQLUTH174T[A60:\=<DR"@I#)K:
P(/V-=#D_(NR&$#J4\;>T-CRA>8\1;\?Q.0HY<&XT+O%C&S(6[KVG@CO45$P7^VR(
P!W((?_?- ]XP,!(X42NWL?3]P@(<09$6I[@5#XUA!OC-$1ATK95+H0WL?<1 G[E>
P\KM<PU='!7>Z^0'-9_U7*%Z<57%:N[P[ .-^YJJ3VHKM9"5>LZO(ZI%R+SP&>8*^
P7P"J1K!R1L>$J9.=5%C3R)<+""'%7=%MBZ-KSBH5DZ]TVHWQ.R^NMP YC4!"2?6Z
PSA?,,M2\.O4!0F)2NZ=IM4\>8Z"_K5,WC2-1K'3,#A7A3Y+.4U^JVW9HNVHX=7Y!
PK?&4&3.S:!3%3'[_^J:D60<>'4@RC+G"9#SL4&#C0EELV3047HE)&7RUB&AN]?E#
PX5ZU5R4_WZR>],P#2SLBWL!4N(<WY@9B'JP4#"RN@P>2**_HZA@#/\8OQ\8RO;P/
P,]T;ZD)-B8@"C>,]CQ,YJR2OIEW[DKT1N/&'4,_R17UG&IU 8X<$3*^#RPA $S;4
P2LRL@X+;"4,'2Y[VHYO"C+RBH$QTY"ABLX\O( VHX@TF&V&,GR)DKBR9+O39BYV 
P$K$3 X/\%]JGMSY\,KY28,)'OV!M(XLC',M">2,T3"#H!!KMT+'&1";F[R?B9Y&2
P:O[ADV,V>!6+[/-8MM72;C!)>OWF<IA4R 98@LV<$Q) (CA[.MWK@$D']XY]ZNTK
P;*["VZ[$9P_M4]:XO<%;B5T3KZ5-46[D="R0G:1N:1U3Q!Z+-GGA#Z]3AH7I!_5M
PL6L @LGC&8&U"""<E15VYP;T7YC*^SD;*F> R#1VF9L9O6ZFSW>-0N$+NG._[&'!
PJQ_=$:I3'5J.[,.#%K''0N2I7_:GOOVG*6++QCEO9(RO/:(2:Y0#;<YG;\<'Y!1;
PVL1,DK5PAKE#"B8"]LW([+BXQA)F]V=%J-L[ML>/I,I8D'FD$XE$I?M%GWLM0( <
P>+*@[6<4AV^R5=:?Z-.*W22(%=9TN0TE(^ZA!PU17<"W,2L!J^6^9%!M+M1XMED3
P0V$%3 "/2&S@8(_?P01+1":C$_TQ/)@P;\$@"&(3C^,S0;%QSCK<,BX^(BJ*_+J*
PD$I.X.':/1S<?=Z>/\;J"OG?K)F&II"P#)Z9[ZN8\.N@]1Q&V=V36U9HFQ4XY/+?
P&5"*E: +Q#!I6H#BTV IOP[7)WE=K%>IY='6UW%5ZLDWFZIZUCK95>V7J,C$K"/4
P(?+-"1[:@BYF M!H)9<9X*T'_ D$Z^/W_'9  _.T1<1^.ISEL?:^GCAMYU+VLJ<N
P;C=EU<):J99Q3];N=)7 N0K]#"@#.O;QXS;L+;CIBS(;1<Z^3L]S1R1>N>'IP(7Y
PY_8>\&G_H5R53NF0]K/G-P@O%&DC!1-#5IZDMI:":?ZZ\,5PX!T%'S<24$J?TA'.
P4WKIV%LU"6 +)P]/3+ '7-GY'"TR3?1JN3GR#SRTD/_V&+9S+.=*&&(N8;A*;DX9
P^Y=9(<IJM3_L_S1J)8;/]RJ6Y;+:="+.\O\T/$?',.*3Z7WX2E3!Q+*6-LD*1_2:
P#("S+N_V8VDB!V[S8$WKS5W\03#?GT+'/=0X^JY>?-4_',)E+$/_>)DU\MR6"%X=
P *ZB-7IEX4N_1<LAX(/-<99/)(X7PAPM9EG"/UC;>->\F0[H;//2<T%\/4,6/I:D
PW?SW8Q+!$BMUU@UAY/W0\,!M+]6,QD?P!9X0!F'N$V)5.XXG0K&#V;WS_FIX?42O
P=#C;F1CG"Q,NK^SDU-Y%$]=@.6\[6A1Z0/JCK:-(?K[[D^3[D0?1-U0@%L%.%+F3
P&Z=ATD29)..,\0_3(#/X2.Y(;39,':OD]-2*DQX/('COWR_>H?E""EJACJ1&Z:[0
P95<E2+6VAKEKOU8!4 O>E^J%<^ 0(NV67\ =BQ7=C8'T)S^#HY>YH<]DBV"*7!XX
P]O?$D.Q =.0V"0D-Y*GC_OK5L8/=^137IH%[;=-RJE%6@H0%O7HQII9 \Z##C_I\
P8#VU]*C+,DN![S(F-A6@8D<IV5V&IA:;)XV3;B! +X@QF1+,8<G N0P*.:7-Z46V
P/GLK\P+$LO&5<,&HH_/KL5M[^(A?>K%'V>Z%7AR%'K1OPY!#?@(0&B3/08=FUMQB
P-X.-X?)=OUN"4$&7^#;67W9B57H[<-=L#TBPCGO X&6(#I"@"O[14[Z[F=NM(;CR
P:_!)8F]Y@0">D-K=K_(+"]3+*+NBR2%0-L[4UYSS.$RN?O(UM7-"9X?L9AX>.??<
P*2_$I"<U-EX<JWMT.$%C%SI\2D.+^OJF( /M/N50$I!&(!6.6\2ZV<"0'C=2(L*%
P/EL):1UUYH$[\ZWGV%?5NBPK3]"02DUAD:Q4(XH<^=+C;(ENR>FG!^#&).[-T@J0
PEB*!T4(RC"VF*J5[RAG<89 DQY:]W<U_\VH5X\!RI4FWGF/0B6[B^G[-:GN$'<OA
P$(0,4V&9X76K92'=5UJ)YM M+R$"NO5Z6EX%X>72)=8FL>R#TWT<A#C(P)WA0G;O
PFK\'J . PQHI=[++KRPG<E(GY<DGI;2,T^1T'L:SNB5*WN55H[ZIHB\,T2L_#XQC
PA!Z8Y),7Y%L9="5A!LRH%G("ZDS%4$//$4'5[-B1E#@_W+C"^LBJ-.7N1_@2EX5"
PB#<7?L"*3WC9A'Z^*R9S-[Y0E\8S*+H_J134):S&9L6GNJG;3DA[A@8$O=K ;[UF
P;)G40M)5 >.$BH?Y^Q)D"5,W06U"Q%OF!66)\ARZC\_W(6"2"ZBW]^I+OCK?TPOQ
P":&Q+&46HJVLXIE_%Y7(CA7KA[19P5=+=-5XL6_QZP5>&F)(4?; M0R]]^AHM&[,
P07C[LD9O8\=) T;,C3:C1P[RJ+E.HC;64;Y[-K54:2"S.>),#Q>5U14\@GRRG4W%
P@HI'D _?Z\:B1]_ZWIEEQ <UL#J-'9"@MJ5%BOLKE*B5!:V2__[7=_V['_U?."/0
P^=G?)/VMT"Q4%50B^:.ZZ*SK]5RD%S:FRKD^HM?_M>]>HZ^[#^F%'H1#7?Y+<&I6
P\"NU3"33R?T+U92W)/WZT#&1P>RW3@:/CSHRV?ZO.B]6N4S@RB%=5OQEKQGB'Y*[
P@;KK%V4[M$!BC=<'S&#O.XT9[G%4@Z%U' 4_.)^S[I%-1=A@:F&KNY*7KM-)87;Z
P5F.I,/4*-X)'6:\U&0#*(2;9>$%%8H\LUVN7+,]2$;@OY">PMLA,*):9O%-($H=1
P2S"_-<&^<G,)#C&SI4ERSCQY^1(= 8.;E^-]%:>)>@9!UFW/_P[M*P!OKR!3JAU(
PPUS'E 57X$:7<<:(85=PQ,,0)/1W-V,TSD7_"S%=X6WV:+)^D?QRAW;,<"IZ-2D8
P\HQ3::45]+X>JJ^R<G@4 ZCQW(:TT+2]#U7<%6=1G?!"A(YP^)G2%)XB.PA9BIFI
PNSX1[<R$RMUOIMLEO0)6"B?27K/4<?8]KEQ>@D&8ZN^E*">:?4.:$I/YCPX0AJZ"
P<E9_C5(=//AQE-LK6 [W]](5>W $N0>7(DBU5$<P!L[[M5<Y9;.Q+]-+JNS><K U
PMU NT#5#O(!]MI$(>>E4'ULD+RYLN-5,""QUE1QUQL!)B:[PWM32%!CN&4;O;H,;
P&Y?J49'93M^>A<2S[!(A4YQ^7UX;?E!RSW!?VUQX/%/W(;US2<5&DP.@XL;V<#[&
P!6NY+_I?!PB9 -CJ[0;P9I#*9ERDFK;:\R#*@VW[G.=+HVE1+UD!3[E,6BOH3+'X
PZ$U)X5X@ EMAP]O G:3+L$AZ3.SY%B-UVQ(W?L6$ZY&@)9B!YLN(AT.R] [2!!LZ
PQ:SF]N3]U MGN&8+MD>#<5M:AE*_ U4:P:B%K5V8P;EP:&6C,&QF4HUEBJW>7Z1^
PQ+\1\J1MJ=3'P-\!,:0&0+)#_K.-\S9WZR)DR>PC"QK)4P,P.F]>DR\G-H(H!9XT
PG'2ZWQ?^&.#.POE"\D9$2HC/)5T#3&KWWJ2:=K/+19PQ*$<]NMGJW B^@Q]'MD_-
PCP8!%  7KLX:=AO8-PGUD] !Y4G$!6Z#*WNF*B9L542?:Z^J15OD2";AM]?3H=:3
PO9';GIF^GD1(?MW<TXS5H)^*1YBA/_1)Q6BJ# N(=<V&@V8D4#>)1\96E<])8WRZ
PC@=8G!*+L+UT?U0$N%MUK>IPYU^O$.2U=912S"EG6T?XLQ+N5X_G(5?>4"1E7/[S
PG.0,'Z[QM_4YK3%9YA/\?YV_B[=XGE%:5Q]>CR5MV XN;%,XO-Q0);XD>B6\N)UH
P#6B,0O>YWL9Y?QFG">B9 Y51O8VF<\0[]*+S3:MN,D(<V[.ST 3'Q2:/N#JB3G,,
P4$$,$NXU=9!G7A:U8X90.F:J4ZUHG:[_;?19O)84Y\5G476F0=&'9,.>8-A^[IN3
P4%'PY?_$LW;Z\N0=#$KVFQ=L^(0]%-VD\$M2=U.\I6M0Q.T"]Q[C>2<=MW0U$<R]
PZ/PU%38)^QN_!)DY%C\=206-,5$QK<71FWZQ27PRG@:X5[C_$,.@4W@7>+";JJ0L
P:[*@4YY:O:^C&N*&IA89")OS$RK?<^>?>[NGNL=')7P*6Y)INHTCW^$:&?@F1PP[
P98;J,:UG?=:>?=#Y ;.0\PHP7$2(CL+3N[KGAS7G+Z'1A[83DY!T$9PYG>>FB$^&
P[I"X6:^K,\L^XK;!Q"OAD.JMQM\;]A._H^9H M[]1]7EE.A*;$I;Q0YT)1GJ%VP^
P/PY:9$Z@]\L>@:5PUIBS[.>XXW1K.04\5G;[55M5)Y(Z5\I0,")/ ">^*F30)  P
P]*ALHB".&E>EA \5B2"A$V3=,E#+U.B=.1*G(/2J7X^[I"H6Z<[QAVQWTLZJ>?%6
P@=YF>-.J(0-T,+!PR*\F.NM"N$!CJ[@EC[J31L:#M@.3?!FJ45IZC4FVID%R+<A^
PT+",K>59K0 V5'&")>&AN%VQ+FX-F$EKWO@#X?MXW%$Y7'_'E+3..*/Z-DD*.;O[
P'B(L2$<!+[%;,^GU,ZDF=#=$Z"LRC]K.;4X4C,DR(<.T3#0M_^Q\V;TK$3(,#:45
P>F=:.%!"0>%KB_5&9<GA"(ZR^J$T1DT?TK%]LM>NO,0P \@D!CCPI0U*"(^*B_I"
P<_MGV-K._-5"ORAE].)6*3D-$U@R@_:J,UYO5?!(/$,OC0#8^<UMKI50S&%&*!=D
P'5!.DS;;I.5*KER+:W@$0/>628K)JC&PDY><^!&'S+2VQ5J18"L +6;)#2JT!$,L
P$,Z/:'_&[Y[-)N&U:E#@"+C2WT#96E^=I5!<Y334X[I90!?^RD+/,QRVCG>A(?36
P;8G#PY7-C:!X\VJBX'VG'(:A!6J1:_%'FII21B[D>R./CH@!ZMKX;;_"\UQX11Y4
PO'&29(K9"(0"4?76B)HER1U]WT%NX!WFXH(K69L(](LHF;IQFY_SK %D[W$ZD?##
P1_V-E10<['1A!W(I78(8A>IPK&78YO)K9_N\'5WH>KV.:#:KY.CBSM&WJ-8A-QSS
P*@+T6W#A(MP<:MKL;0*A=S,F-]S1O6GU925(U>6W%^-Y98? Z_$\^8+Y22$$5KDM
PGW]9>12SY72V@%D!+TA>IH[;Q'!+[M<B#!M L;>H#=>3 <VM67Z>Q>.0TSH,4&^*
PL:QBZO+9)8R23TCWD(3<L-1=E.K):,H#TU[C90IA?!$:]$XL-39L!.JX2FW_AY2/
PGAZ[J(T0@K0U9Y2,@U:6,FJ;.=!IAPEA#,:Z^Q,:U1A'??H".7)Y?0]0=<FT[]UP
P.^*$N.1ONO](HHNZFCB>A;FBUC3'+O3[UR9SA8*UN5JF9G8+%Q' ]D#J>M=DNVN*
PCB*9V8B5:JOA>SE]$F.="9_.DW0V@%U4+K(Y"1:4CY=#TVG"N#8RM=Y13<8C@"MA
PX5BK):^M(LRQ8_P'9V&2E;*"3)=\9F7P;E@>Z'-L.GQ!<[";-AR.\C?GZ$))9WDZ
P0#ZLEEW@T<4JZ5N3_FTZU>N@,\,87%52%\N>N58GR7SH;@&:;9GSM$[QS!L='B/S
PUJ\_S$9%<7/L8^M(2#EZL_']N_;J]*,0MA-.E$Y,S^%>]&,O9VBWL<NM$"BG\RWG
PI KU0%=3N_6<F/;VZY Q.I!Y+O,8LDN1ES]U5J9C;9U-R!;[-;HQN#Y\4 Q1!-97
P#T@"?5Z_E^WRO)L?=TL2KQ#NN"!]@.N7#A2$?AYAE%P6=:\F0,K1B+'N1#7'G%9=
P.M8]4N[@^9J^N;**Y7+)16YX6Z3[+D"[5.GTI*9O#$["*,7V_(5A!(E&[(H0U^1Z
PDD=*GFALO@6I=&^;IK='9)ZPQ*\JG+3< ;VO;>%,FFK<]_8AVTR<T2%)$?1J4H/O
PO%*X'58W_75XY2?_VP/UEPW/*XG^U?D>QWAN92;-?VH'F </AS=Y1!._7N3MLNK[
PS+)LGRK/=3S=E#OTR\I/7HM]738EWG=3KX UEG]4BI*^;0P_R\D!.6YA(].-R_Z1
P(%5Z%1GJ.UOBO;_$QVF])G/UG!3P$&DOD6OH^ H]00'M2 2P5XAG_J*[Q'PWMP#R
PAVF5F;_\'2>&EB8E8L\(.J(?)FTSLP$-3,7TA.!_F(]^JW_:WD<':@Z< B,ZOGTT
PR@#5!S1O?YQJ'+'>\%63)S0ZLU*XF08&WM1=1[78B\##P%GI[\DOAXJ?98H1K]IZ
PY?U%_PJ&,=NJ7<1QX;46WNK-,A,&T]]HZ*PM:A8,H;%>62<KZM5HNE=:[TI.Q0IH
PA;2/U/(2.2!@,.8L[BKJD]&R^+Y013<:+[QTS!#9,PV*^U-.'+]0JN:M<(M,_49D
P*%<%F^GK?((*81X&;@+YM0W/4,FQNNB%<_]Z]<VFO^T08J-J"3(/9R=TFYB*/(%F
P-4+%6>'&$KD3Y=.9$,G$N4%%Q8-LT5)9IFRF,6IX1&K$R[4QVZ,X# QE<T:TH!(H
P@[)%/<,KU7"8CJ;[V8EXLE7QDSSS 3=394>?BI6\Y=HG:NB&'5IG^+LQU)4/8?R$
P7!J2(%UL);'[29WT.K>%U$6QNCNJ2!.XJ(S,F<<S67MPG)+&=7$1K9-&K$]Z?<--
PO?5TBK[,.,9^U\W4T'&B0C7M7:FY+[./K9]--)XJKEV;U=>^ZN,_&S Y4@ $L97D
P!3\Z>3H\K.^HENX>655/P]$DVR7P<S<T$>"((U$:#5A@@5&(L!>G'8:+VR.:(_9J
PH7E]7ERL8;UI4<F@8O( @_K0UY%@H%AC^!SL\V)$OY?QWR0*RY2=?+C57?(=5U\A
P+O,[SK"R'B3H,UC!VZ2X,(1"\Q( RFE) #!_-H-/N3LU'72JGB(#K/K@4]4KXGL/
PCCE&\3W&(8YZ$S]X&FF>,ZTH&TGQ_U\C]+1=0ETOEKE$"0V/^X0?#+L2^I Q[,<D
P(_=1SKMP_4O /6CG&;9[O">URWDNI1P\B@&;;9_4$Y5_T?,TBFTR'6LR6B7U322#
P%4>P!T,+U-0U$6ZV;4SA^(#?6G:RF4+VQ<EEW,]'>6& 0AG2ME(T^25MUHJC-&^)
P0Y2S@<7I+6FOC0JGJ2=^EI2(U2SV1M=:(-N!=8E!:BR?+/6(=334*P/Z0\0OPAYT
P@2N#/^4".N#,:Z$Z;Q1XCNW&5&Z*WLX"N')G%SY&Q*52F)T"X);# ;+84K^">8P@
PR\?.'.R9)X[R6QNIJQB.^=CH5BM6O%8EVF=W8]CYM"4<$%!2SP5R=#X"4?8LK YN
P++(8.[I2&8*&-@JR.W)/34+>G^%@6:"JO)*- 8J<W3TH/?K.'*Z08YK 1O[L MVY
P)+:A6((Q\JM"C*BQ'<S4)H8,+E(,FUP'EU\^.E3:!)/,&MV^I:;79F+V(K*#WW,5
P5I$X)P)A<=<9<[H(/%TPW.39KD%YX5A]?XXYXM+X(1Z;\];$:WXQM9JD-GI9JWQJ
PZB->LV'\.&,1-MO- 7HFD+!<#K].:A*2 %Y3=C>KT/LVT8VFE@D1(3AUCB]9H']M
PW-IS5RYV,V"U;ZC%9Q!Q+C&2M5)UXQ@?"S;':(46Q\"2!I[X/7VS'OA DW+=>2"=
PY75Y5GEY?<^(6;J ,Y5;YL+INA1-.KN>HUFAFP&D"?NHOOOM"U>T+& GOELJ0:\A
P!Z"OILB;]D2D]])0H[GG]_7"$W"HJ[)PBT:1]:6]4D/(I"R!8']G\S\R%(Q1-C-0
P)/&G]G[\#(0.&E2F$?6'2Y'>VBUN%L!8_D2T:W.0%X7D/\>;+96E&DC+_;OW<G/7
P+H1)'PQL9ZJ5+,Z,@E#"7LIZM>NO>&Y]:\/+9:U'$I/@W_C^@R(1T[<7NEGL8[]F
P@M$UN9)G/8N]6G#&<;.+CLU%<9V2Y >E(??!P^?7*FB]I)'N3U-].K8C;RRLHAO!
P,CF!94%!ARV=TMN4W7X)_(@8O=4BL1)&FNU18LM0R,.H]$68HXP8&Y%<&U*.&CFW
P0"' C[,JA+3(Z:YNTHAZ*<N<G Q&QO,66=RNE1\\+:J33KALE%763^KX,]#LE_JM
P%T8JX7HJKO]G+JHTT**! <UC'/%Q*T3%1--F8F5:OI6?1M<'(.%WH VM=<H_(J+4
P=-EI@W#19#T *0+*!EFA^>'$+AAIFA^YH?YD>X9]</B"N,FT0N51>'P_-DC(AYE=
PX1*+?BG^U P6JH4-.<-LUMEH6OR__ES2V',"KX', 2XJJ.,JUSKRHIPB_5'6&9C^
P1/K?&[]TK"H]THQ'@=PW*U=W:1KL1T>(PG.0L/O,DMWUQO4,L\F># C&EKZS6'$M
P[PA$XZ6SM""Y2*$P\@$5 F$D>I$YX=ADHSAME>%9&AD;_+6W2L%L4\/"#$YW)*J&
P.I%;+0$&;[#TK[QQM"3VLHN)/29 1J6@Q?+(>L'> UO5^CU?-$.N!FA/P.:_\YIP
P(;$Z.G<JQ+6SS<*3\?,)@M!KZF[0T5!>C/@6VL!]26;"G_$W@J)I8:/S4$&XVW5]
P=GV\9;_DIGLQC;K#"/"(JJ[3XWL6D*A-2@M0F]@UX."M?"?*R_$$T+X3/HAP*XL!
P!#UJ'OK=.'%Z@6Y>@KW\C80IP<_'#)_Z2"X9L>)!"2TN-F$T;R,H&<WGSF<UF(S+
P%JX:0R&L(V7.'?&,I]0J;9G \IKI6;'^!+"T4HQ6*7/K\?@.TSY>':L+U\*(W/M-
PCY!]W&UG!AD("Q!4EN.X\U.(=XN7NN<&_'T37#G[!KE&K69B1PCU=^<C'?\%C5:N
P20006E#EH.EDC0:XJF+[HE&:OYS0\=9LM:/0)Y\/Q05+PM[+A-Y!;S$'RT9<'V0/
P6+J5*$+>B,!F7.(]$[S?&4!@I<J<913.!U.7,[KDL'?4T:@>>#>0(K 35%!-+ ]^
PHNR_U7F$H[>B?;D)G4MPL,&"8039/9,C/KNT8$H;0G!:*PO*I!#D$5V*.#DD*4FN
P'7L04?*1B?Z)<[$,&^P4,R;HFQ_ :@WG_2:",.4Z\D#7K!F8!#J1ZV6,@L-GG;V:
P'V&>*"+FJ&L)XZ;X!<MO@[IXPIXL>&+7U%('C9I%:4B70GW.(>R4\FU.72#?_$++
PO];$"\% *M9*I1#<:>5K+'*?+=,1.<CB=U# 52WN@J@YXH79&WUH#B%61H7^2JO9
PHH56BA]D%UD#_,S7D-7_I2>_O"#$C:/-&/D!4!+]I5!PMK0."!!P@-U-_X=6VTC?
PO2W[Z>98%/FERD.-@(8D(A-[/1#)2.[\9+U2'_2#9I P)AVE$%^QXCGT-5B15PZC
P&ZH&6$Q]:J<#0OOQLH48ESD5H7G)YH"CO<7RK)L<C1K7[5_#KK:C,?R$0:$JJ.)'
PI1,[I=[D$AB1")]SG@MR=+O%I0US=E%Y*',P+#4,O<J&?JXJB>J,QJEKO#G__T8>
PYA742]0\4'*+*5/'Q"F=J/17/(NT>WO$LIQ9?\C@GPAY.9&L+MSX_Y%"SI,'4;?T
P <#<*7UU"05CW6R)&0>:N%S]B%?;#:9G8I]#9*%7;G'#5)C@<S7/T0E?_++(-B'8
P!WL3.E<8?SMP2^@'"7C@8?!(#X#Y5B5FC3(5VGG;WWVHH!/7U\'?S6 R2=!1P2[F
P.M,Z_T75;DO;.W;C\;&A+NS$\JR2A?;-^X(_X$IIFV\+V,7B$N4WZ?8;[C+VB=^ 
PQ[S&C0&DM,3"3O*%UZ"QD .4!2PE!X'"#9__.)WO.G5=URRDKR7P]T5;H@5M,([A
PDK)E%J&R*N?L260<*!]LYGLY#>D!+'XW<(+G\Z?6&YJK>XB5\0ZC!_X5\)).OTVN
P>6HW*7_-):Z%[/MY;64MA4R=7H16H'="!9K?.2^6=KCQIA.Y0R\EN1F]??MA$&B]
PJG'WWW!.W0;\OX34,1\11Q"UHV&%Q0@/ Q&X#:ZG!<:1?D"5X:P*^9OA _KJT=N]
P/\1EC,?'I_:AQ\ISA:,[=7A:(N<>Y84.GV#>J4 -XXS&AFR4'U5&)2NI[=>^@> ^
PE1'+"75-TXV14N:(9[3)B^ATHARHB9O"INB37?;719CWR@#Y!\CY_<V096QW\"4Q
PA[>*S!BY\IUI16?+,2LO 3_Q$";2"@C+-;0[,:I''=SJS)32>4BSO>L]6WQ<ZQKZ
P[(HL(%:Z;@"GX2O==IO2 5(VVVB84N2'W93IG"_O0P\F5YI[W7G2E@.^7&;V5MJW
P"O+T3][0 !N@F32 ;R]:F75:2Z+$5A:=X3XA_FB4JI)7FP[@]2\UBYI *34W+DF=
P7%1]0F542_[5-7]XT&%PA:/L+ Y"(2+Z[(K+.*V=38S5A"M G06E%6"4HK70N<[1
P,.U!SZ>"FSY,J1WRZW9"D^XFB%N \BQ%5_Y5M3R0AVKP]^Q4B FS'"6X\RG:N/M0
PJ!_K[?K]WR=LN4TT,]@^-@NOPB5P;\TVUQQ'_JJ+[Y@2DZC6')*>1E,?0/\,%588
P&/:MT'H=R] $7@<WT7%#+1.6]SX#^%85?6[NR$[*^X?QD<Y=A3\Q<0PP[0/['S0>
P[CKAWQ./J+/.S?;ANGK02WP6W(H -3$J-P<A^/1 NLNI%W#:%#O"Z&7&FCU-5((E
P]H_',8GF)LH[JE)"!W@*I5A+R-N_K2BDJ)@6*;/RMD)GA,6K?(&.O8IL-6 <3X?^
P7Q_'4CFF;6BLA\T:H,B1G[$(L4J&E,E]99*3G9>@8![@(QP@\U?.%04O@II]N87!
P6"IF3O9\=ERGQPJA#=C #LOZ1QS9W'KS] X #@Q7*?Z:N-NBVB+$*.8;,.)VN&1W
P?E\(Y#D5RS9&LUZKP2'T1 _N-!CY,PNR--AZTB4^E'VA0D1/WZ>4<NEQ;DG!,?]W
P+:U4S4@!WE^E0FGJMD;FIZE6V><I,X);NJ[L=RDRU8]:3<)\3L._5=;NQ=&)W(HB
P&9W/C*KJ38B?%LIN%_I3/J+YN]&1NW'@X#3T3/R^?F\V.6.LD;K@95M"P+I=X;3B
P9%Q. ,TR[>'2-X6@=-R<TND#)=Q<! FLLGH4V'K@LA$YDP85#FB1;J:F5)1)GE#,
P)[00ED/2%#?2&;/.6H\(H\\WA8%4:1-#=<,GEE$8Z0*CF_ZDJE\H9.+F&UF9$2:8
PH3]$W&OMJ12??KN?0]50JVKETM^CJ!\-(6M=<$#8M'V$)6G.A9ZE?)_R3SKP*T#Q
P-&7_XH#J#X4BM[- T\")6\0$<5I]V+4KBJD$NZ8U7;/4'9DG 1.;Q$HHW]W9#OXA
P*+C/1>0G>'+SJM-US1I6D/09PK]Q1XZ:#"5O5K751;G1WC(1=WBP1JI>EKQ/R7+O
P)URV#PAV,^&QCZ;<I=L9IN9(:N0S2"$_(<#I%[OW%U0!V;5,SY%09#!(>KJ;)]3'
P.1:QPC-89'"&C]"L>]UYB4I+]3;3N4[B)]=]05=,DQ >[X\^5B6]*MU? +FCI8'1
PAUL8O:,"N#"A#YA,CP'_T6%B<#! %-!?IA<X?H8[@U/PV.9''">@U-AG,D_;KW-]
P")6?+@(-46?:[!2("2A%EL%2Z7RAH;_H&[99=6U-TF-XP[D:4?;J]1-$L0SUJODO
PIF"!V*7BNXL0 6G9JX;/Z+(//=IL,40_68@ =C[N>C720><RXR#2,EMIFQG' L*:
PVJ"+$C/3H&LAAN[IG[YV:5FM;QBML="DC9E_H>8P_$M8M\53GU(6S)<U^9I/(3(/
P>YG$;"T-ZD@X+^X.PN,=)P$<.KEG*[UJ\_.[[BQS<<%PM^J_>0N!(TZ2@^*Q>H!5
P5#P_OK+E>+W']P38%U@"E<?E5Z7^'&)546*=75\V>UZ>Z,!7*SK[%3R]!Q#90L4#
PC1B#*[[@81J+>3/$:W<BZ"TE VI4W4&QZ)XQ*/ SKON1*,5A!A9!YHI%U5?+R^(A
P7"!=E>?36#1%;Q8"538>_&.X55C^#';WG410ZU1V&AR>5,[.:7[@V-FEV:ZOGJN9
PR8';*9LLRZ89%=[.%]>CY)JEEG15J-O;'6Y5(AC6$9XCL*0(+%_(R+?GV401SBL4
PZ/Q2H5=0 BSHAH5[* "#'VP,<4[)GMS3B2!RY70E6JZ\3/AT] OFJ GA9/A#1CNT
PZ]#2)J?)V$=BKC,>7=[I^: 6<&5JT1Y<+!6>PE;ZS<3"*W#@(I,9W[ODE<)XI:48
PSK :(BR5J1.%M7Y[/,D9JG+\<G4*P4I#%NN=U#B4NR,YI%T,(5 NF+;E8UK -@1L
P2T*LWT//! 6JRQI?MPL(DHUMA0?9Z3M-)B<NLE./J%0"%$77>-%E\<F@X+2+W<;:
P(!ARAV\%:V:6\W9.XA#CA\7E^!Y:BB&\\4",ZI'8T+EV?D9H$:,/*"%QWQK8ZWBC
P#UMUX?B4:O:/"-6P:VV5U[MTK]H7/NIQ\ENF;H_0@QS'<\# L(8%3PL_8-S]TDS 
PL>DA"-0_YX.?TZ*_VA:!O2]#^<)A-S(E01E\1.LP LV@XJL'\\ AV"&?CK.\R8@)
PX.L2/,3IZX!C5E[W)F4";&_2<1B&K5"IB0BO,K^*%4HBIMG7$5-8:)K$P,0.; 9I
P&:)L";LT#"GWCNSR=8CV;AR*2_$Z6J"AV5F"C#RQ+<&$1U;V.Q6&8>!..#5R-VVI
PH^0_5$A<&*$XMZJ,NTNG'''(I)Q+-.+JSV?9GC)GBZ42!*JNI,VTUN]41NADL6!(
P00#)Z$ OJM=QEUQ.PZ(-=9V\_30TP@)_]#AM3(J1ZU<2>)XK!8U]R#=E;"HWT):A
PTU%[O^]T]":??KT]#E1'>S-JWZFT2>%2ROWNC^B&B-?-QM.VA  DDR"!B *J=32.
P3,3"'N)<-K]R#3Z71"Q]P>$05#A+C4NKKJWI<5_[A6/MVO]=TG"R&S;1R4<@/D-F
PX4O(8"2A!P(#4(JAC[2$Y<FY,B!W4=,NYA=8P/E#ER;[OVKA6?(P==,S-W/9O4'N
PWRCB(Y[B4N6;! 4>1' ?6I#>C'GB&9+/7"KO[2->ZF-.[8Q;4IF:',T>R%BUU&>Y
P]LM\3/[L9%EN^#>WF!/U9/94!L7J4XQNNR*.&0*O#?-D4)MQ:I:K1MC""C(M,DF1
P@HDBFD9P1G-3,2Y#;K485P^Q,<NQD0KOEICF.D%^!6RE@= JDYN3&][LZ8RUUBHR
P#\<N]=XL]L*O1MT7*\MQGDDOE;N&(DW["$=Z,QJ4J;KP65ZSH(S.HUVDJ[,>I#9-
P)>%U%,'PGCW^_ *VZ.T2 U-5H.WC089LGLWH9JI8-I6$B^1NX3=1WE,=,Z,;3^5F
P K>4S-<D!"\?/9D8UK!=A"V)A#DD\4"^P#:-CZMT*^.NZAV'HZX[GI?%+\I-*$GE
P84OV75SW#92NW7*$#0(O3XW]8OV8IS7[E*(S.Y-X?0:G=)QV/4 ;#O$HS#.IC%H$
PA78A?LNW-AL@7(QBN^I395>'F@A,C)4!J1-']K Q$?,7 K9MH\' WS5C>]8*3\C-
P#FYCR0JT320]YW'A^#)- 9F,.JX;BO:E]V\1L]MD;CK38LZL=,A';@$(O-UYX.0V
P*T.#[\PRU$($;+@6!B%7QM(WA-*8FN 1KXO)<5A"),",]P?_RMQQ"SV-6E4IO]OR
PT<)WDE\4KDT75W4SA5&Z0T7*M/R^;Y0QB??A6D66(.F1ST](# !+WM8%QZFZK1J]
PG1]O]%3^J'&S RX?\>#5=LX@<FQXH!<LN+@3CIY";TSJ[V'ONZCZ,56R!$7-TK*I
P)M!$8Q?3]>I8%RD<# P=38O7OT4()(D'LY6PEQ7='1J_;4KJ,M!B;G;?_-YO\V<&
P#@*[P[Q,J6\<J_W/&=&9 2!LE8RMYW'[$U(+^/@@@=^/J3(A)Y.XC2/\W+9"B&1*
PL;& 4_P-[#T;@A725"ZV+ TH I7Q.K:"<FE#!8K5LC00%NJUKN&9[8_ ?HSHZ+SB
P=-^7I.I1IY'YPA+/D/@#MV)H$<?!I?N-X4:+N43#JX+.LL;C>!XAD7%-EF(!*^1,
P_"'P@8I0WE_'^%CNE5O2)-&T=<8RW$X*Y/_EOY'"MF,DN8[B3@$4NZ_[F1G-9S4'
PU__0&_+A<-1P00YYOV6LVQ?Z]WX=\F7LIX?OZSX</V$T7;AQ&G:0_W +3[1O,!+:
P9!1Y)(I!E"ED6:P-E9ADE5\TCU/ZU*@W:S+.Q-V[#DK4]YRGOI-X5'/WH#V;4AK&
PB *9'#?6AEL\UCJ3^G?\$@\<UI3"I%0F'&WV-#XZ]T;^?"B"Z""QSM42^X]0*F@'
PJ94K49OH6)"KOM"12Q DR*9M'%>Q[W?![DLU[>YI$A&UQ0N4,YFM3<Q$T,^+^6Q&
P,R#YGL-5-$.JP<GZM#SRV>Z)=-M>9(6(H%<2LVS1^HU0R*Q8E'_)S>U7SYFILS]F
PU6$ -'51K/X?#%XZ+8F^V@/H3)BA8,E1#+>I4]E B5]$C<8P 3$B9W:+]5 U>,S-
P'FD95OVVQ!.4K;53(T $D<UPFY9N'MR+CA;"A9^.'&46E7GO8%EKLLE2\J7R.6*P
PBD/L\G^YO':Z94W9K6.$QWTJ=YF1.]DLKPX[%X_(^:1!*9.P()E-]LF2-_^I]V[Y
PH,TFA=)S -U6=MO@7EE-;JC4/(=PN..04]^\E2#<WYLV5&MPC@)%IG>>4XB#0:2R
PK5+*Y!.-T3"O(J6W(>3!-KSG>22"9UQ3\:#YZF *K"RE$47LL13\KJ@Z#'SZ!<MD
PIK=B-1V.V3$)YK-GL3V\4''ON:)$7U)GGSC0HZ7D&5D<(Y3HDSG""D_7B) \9M]0
P%$$Y%-J%RYH,>?USL\8"!X!5%E+Z+^HY=CD5N3K?JI2!R^&3.KS:0\&,C%8_689P
P!I+JA=6YBD@$REOC-]D<@CM7(K^QX*Q+LKC/:D;LY'.<>Y4]A^+UKIJ(9 I/E%)I
P3!MD28BHY]OA0'9K+64\<2'#C+'1&,%EIR,N*\6_E Z:[VZLNVPQY5VDBV3#:@UA
P%K_Z*.[L9VZY\8JXEU,7W$'Q7\1;.BAOVR4RR1R33A_W1W'%K>6\[R,N!_U,VY:Y
PLX%%,3L:1M3QD8(73N,\F@W:JUG,QC@%V#ZI@9COOHX^W>Q/%H=YZG9: [ER5#@Q
PANJ=<N76D3Z.H&3[6JKXI>N'CQ2;Y+VQ=.DO//8\!B9R;@(B R+ I$3[4UF<\BP7
PFO$LI(L/*.]$YB^9KKYAI*?"4*SNW<(]5A("0%U3CIAF/HOJFA+8'&OO87A"SDII
P"4R=@"H+;-(=F@G3?TV\^:4X+_56UQ=AM#9;JC6W3<NF?G_Y5=F9$EX-%(4P"U!=
P6^&3PRFWX!*8@&!D\5#66N;TW=B64P$7)XO&-!(3D'-V_?RI=*BS1+-1U4+3P)F,
PR7!Q )?%C\CN[I:G^F%ZND@W)H=ER<E2;(9$5N^= ^^;]RY:7GC&J:52BO%)+F=B
P5!^WZL:&"[7\YR!1IN#&3&BMSVE7>PQL/C3?<*)=4)IH$>L_TU#%P,&4IAJ0V.Q^
P;QT6J2E?-X.!87%:0^MBV;O&D<U04OD9])Q*[#+P>)R^Q/'==1TTP%5"3\$,*FU9
P1&KS&?%?QY#^C^SE*8C= "?6WNT0)8H7M%S_G.I:A-45RB5+@K,)_BLG_U%4KLP4
P\T+T6@X2#M39^;HWP_U[WSW7MC(M1.GBG^2<BP?%%+W>I*Y-:<_A>5%[!:[YE$IJ
P$HCH)!K6P6-V;PKC.Q)M/%-+#$,!:B<TIH/60G/!;*B=A<-'X%.V..DU=%^C28Z^
PXLKW)KU6]@.\@?!KQHG7$_M>N5;LH>E;;5MK:CPH2D-Z,TJ#8K%6[E*'#L]-21HY
P[:R,E_53Y R2W]Z).#MSR8IS,P9-YMI4.D H\GVB)4LRXL9Y$7\6R(LI!IDHRCFO
P)#^]+%+,]$9,%T,V[F(>3/H'2+,MHYF]QM\=XEE$;6DO59[=99J)C]7[J0!"D\5A
PSC-)S]LX%$#&<+&1Y^ "^<.:^=RJ65L]W7"LV$*H%'K7!@8EQW4[NM;9%SEN,XLN
PV4;ZT.HR4'S^N3E'_>U^[4]F%;V@QG+>_V!G2BT@'X)\ISMYD^<O3-W]C8\1F89I
PIDN[<D528#,+*_!2"XE[./=:KUD'*L[D5NG_ZZ*DQ )%U)2.]KS?2;#!6D-YJD%+
P1#[HC[1#WHW^G0BC^B*"]3^Z^=\%VB#_9:$._RSJ2\/\2VBQSD8#^.,Z"\>5#F% 
P9+K:11=TJSDX=KJO$X8>K.N:LE?T8$HF=!<EUT>"W\)<Z!%\*?UXG[+V]$OGWQ]*
P:$U9=-(^JOY)%8A?3W/_X5S]R?V09R=M)+Z\"%'NUYREMW -[_<*TD?KC8-+I#DL
P8;U "PL0F.43J.+0E!^E2J45[+C6CLN\>2<P,QF1:UJ@IP[[@("M1---;F6R;%O3
P-.7/AQ ]'[30]DA%H0GP%0_M$[.:^GL7T1)3XUY/SZ[[]TQ%?=Y%^+U_^P=2/H:-
PK:$.$\"^C9_':ZZ@7M &99:K<)N6^I%XSM=.0JB'QZAC"B^= E/*!W42UPU%/0Z6
PV532:;C5/6 F$5H,N.+F[M<6U;<$?J?I2AB4?ZK0>8L(D*_?F(";"9A?[E7YM:W*
PN+,R]@'G-1[2 AES'UO>,A4\B%#:\[H;G0*8%7V-;"UL:A-OVUC*.Z)_D9;Z,9;-
PD>P,:KEE3B@37^?ENT7A[U\:>;%W!E/N_ 5NV7QI&GU6E/L-3PJ-)$!+THQD6T/1
P,KMF,<\IEX-OM[OL?D1B+N(&S"K"2LMC;GS!80:PNX: V_NF\(F9I\+Q+"(W:+-.
P/D(A[Y(MX6O.[G^BZHD4BHFKDAOM\N)R\,/6G7G'Y64CL<UPC3!4\]'"N'H';SXD
P$@CNQ;YM=DX81K)'L&,;FKD>8DU65BA;AJV(<^"4'AMPJ?5(#-/XMOD>,Y_C)AWZ
P>5S#MOS,%P!:'I%G$%8V!/L =BZUFR@N?RP08@VHT-.A ,8+K8\@N_22S_8_X!E=
PIM^?22F#K@[R'EZ*7F)%A?*7Y?4V>*[:I2@:TWL0JEX+]:[=?<T':!-'-%_ONG]<
PS4)NWH$F.9R])[,Y9\HEEETZ '^55V:(XO9- ))L?!9M085T<@+ZK;99\UF6SS8L
P;*/BIA$:Y9@Y)*R8739*670M? _RU[,V:+O>?9 G[><6-^;/)I>B%(H*JDFV2M=[
P$5H-Z2 (*F!!DE+?;?PJU$<CW>?BW/M8I,JG[E _I_M1(?/0^]OCZN*BQTY<70J9
PQVRW71U_JG$A>EL/O&\2D;LS(B[1A69H:6$U6PF.6P[9J9JFZK1NKL6+G_F %T6(
P"=X58?B#LMVWUI0 #\1CH,G-*L25L@('[##]@Q2A4E712<5JB_L@ <RIIS\ZM0BL
PV<0VK]^J]..E*1A9I<=60@9 )CBXQ[3]K-%@]QKO@KA?2^.OX+Q0[_,>?D/(@$99
P%J)D?+VOVD7V9R'HFW)#\GF3.U<<C6A;;?/4K(R>M6. * 4GO',=Y2<:& 6>[AZ,
P[HHJ_R/OI\B'YN.$N9]Q/BK*>)&CY03R1X1$BV)R; FB@GW>NK'2Q1[S&53^FDXB
PIECD2R[H5Z-Z18Z:OW'B1XK0RQN-LG;6<\QC\R>&/[U;<*$LUKRTOC3176119IU 
PD>@*?$U%2G^5>^$PC"0+@?R-;1/E#$MVPTG#"3'N<NM/%T5#JI4_C%!FZ4\QWY80
PPJD-4*U$85@:RLUA*HT^-R0R*A.W#H];]OX6+EPL8%=I_'P9)"MU"0-<?^8S)U\&
PL!P+OW6SUT-)NEFFF P2@O<,SE_58/E=8P!GM7L@KV>6B6U3NA;Z4TA;:'9U:0%I
PW='@F%66P]A48\UC@='WJ76^3>C*Z<F<D%GNU!<*AH>235$M\6;?IQ/X2OI3)_=7
P2^$ 8K5C,LUW?:/NIM-/6>K+Y%!&X%)8Q._AB#+ZI0++'PAG3('PE" (@IWJ=*JY
P!FH450&AOK[#N<_JXR0L=@=)0ES@TK]<<W*_&3MX.#@<7IH,O@3A_GFSBK$#=\]3
PG%[C-9X,4<JPSI:Z1##-Z^03VU"#&>\OHI(79+03^P1Q,ZR;3J&5R/%/RQN%^]/!
P9N8R_I5<6XL%_D3868&6T)MF+K$T5E'RFSL2Z54'Z.[\\9'9O8YXGK=QZZ6.&/:L
P+*XE>%$<9#?63C56\R;7TH-)>'U-S0Q2NI:3*J%-U$A+@K&1!XZ%$U+-=':0\5B>
P6O,F,WI9B<S CKN2^*$]5A)EV'S)]__=V<];+5'N2=HAP3--?2=R].O]2X-/<=!,
P ?1#C.K"0:/0%N1TT[X]UTD[SB<M.B<JY,'4LM;*]]!5!-$<KPWYHA# *C@3O*<S
P?98G2D@SG7,MO&RK9A,_O8M[U<A2D"X;[U/8 :##J=V_TZW[A2>#"'Q6;VD6'C4E
P(XUH='0&42=K1;@MA,DBUOL\3.. !O_3=)1?#\SNKARE_E'[C.4ASPJ*_OL60F6,
P/ESP"+CX8.AD8MA5?VC[=CL#))Q@_,BROF6W+C5*)NT(RJF16##96_</:G>HL<&H
PI_'X.;$Q2FVL[1X=_ZB:T6,L!YF"*?JO>?SY3,84IF&%K-VU]+=ONX77 9JI)*9B
P%7S<<PZ_K <X_.U!%G!W-<O+ 8S6K=P0[&&+RLV;VVN1CD11L$6TG7F-#2MR][,D
P"O M$(S7<T*=DF*Q@] P-Y0>C!T^IRVVI:<WVWGB\"H]!7L,!0F5JD/7'I^C[?).
P#LU$W8-FOV3IRF]E5SQ_>0Q\,.GP5!!!T4LT2]KV61QF 09-L BV"<O!#7&1T_E7
P)EP5)'(B&#/%/XD U>\W(M=<KZ2<9?M?^S&-%)=!@ZU:*%-*V8TP$$ DP&[G17\6
P/[-N[HA3'SI'4:'5IR+B!?0@,2+HN97M-0IOZ@_1IT^Z,&]D^@0@@SB'PG:9+8>(
P#^17_JQK82Q#_,ZU;I_ME@:7#O\HC-)$,_LG<%N Q=(_+;2EUME ,%WAC6/N&/(O
PDGH#5&V72E %7-LSZM%7"?$PY%1_4J;XW["B\M)_!R9,6>RXI3Z7G]\P8;YL0-C'
P;;R_NNH<](B*C475HL^"$<H7;>UHO-"N']Q6(38U5A$J/>Y!24)T*.TX-7@A3<P\
P1(.T8ID\W2BSY*>[K<\0CQG"F_CP.Y.A_=G]&59S\>!2#8H$IT9I*7A4^C(X,Y][
P([>!&U&7KKJ1H&!O%[*-\!4O,RJO7T73,&Y.#H](^61E_P?L2C3L=QU ('?6705>
P 9!VCSF>'U38]-(XX>[?=_^LI=[&A/%C.*SK^/3CE]]/4K1,N.'^(R);_!?S;L/V
PGD'!  LM'1O\3 27>QP] 5BW/N_54?D!Z\UI 'YZCN&*B,K8)?O!V0XZ38I!]_$=
PE=5 =(ZJ?)DP@Q?^;<R1=]+Z]^O>08V"A%C?/O=N@6B;)R^_S#T%*D.6UKU)#/4!
P[#!HMFBR/O&$N-AA,>)H;/^[\"XP"4 >^;Q-NV[.T;R=9 >[>6=L_,0$GEE%;XS6
P*@ 8R:CK8AH.M&$DI1> #O_P_05#8STNJ5,YHUQ&>A>GNU[R6(64YYN@E8(3<ZK6
P'G'PFMQR(?HN9^(C.E(Z\?M'?U\XPZ?IF6YS)&&4OA;O6A=_^(.S\2N4,VC-A2MC
P:;3(YS/:I=V6S'NC2'#::72MA;IDP:K0X,988EE"P*-Q4/C;P6($/4YWMYE8A<7G
P5WDAL\[7EA[-8@/]?GV!GBF!^53CWF^CR; B&2P5Z;99WRK^3'7QQE'<1?^EY!J:
PH*TBR@@&LR'G@10R[JN+0R,2(8 C88B,&,"&*R\>KK/^^K%98;M,7V_=09 @7P4)
P#N7OWF]M<(8NO3HC?IVAS:OP^?$)-M(EK&M3$/%A1FDCW"//$ ;!)P FLG$4M(=1
PH55E/B.=PW[TG:JE15&4)1,'>^$M#3(V[KL]\T&A18*Q#6BK(M#%0*1OF-M7J8:?
P@W6=('*E/^7@7'A)JX(%PF-]"<016$4T<E@2XK\8_<6Z>@*>42+=>._@T 4CZIGC
P@9-$=X)ZE>[FVL>_E=X!-)'4-S N+I)GN'.C6AXTZ^\M,,8^+LJ8TA?V6U>TOO+<
P((# B/M+5Z#'%:_VX"WSXDE6SM#DE,E?=%]A7U:D>1 Q+Z<@W,$UL=2,">/>8TL0
PBI5(Y\F4H^8E0N;]VK7/^ \6>+";'!6GX"1=_,4I+[+$ZLOW#9P%PL)E'=8L:E?W
PPS)X$SM-<>^&EHBXJ)_F@=LQ( ? ?>-JK<!_462"M8 CK6['=21#V$5,<6RK!SB'
PRM7=MP26AO?W!:];W2S$OU!$SC4&6PY5J.UC*OG="Q0#!> ('RC,Q43L8K"GV6YJ
PQ''7+S&,H.)? _CW.W4ZZX:\(_*4H9!A=D7#V][>$Q5]=>K"7KFZ,9G?7<URB8J/
P;1N1R%T%2WH'2RPW(OS:C76>H8VDJ;U1JIH?4JN>Y,(4X&:XN<[F>&W,_UI"8@7,
P[(JZK'JE31.?FY'7X+K/?<.JM$'Y%D+8[5/_Z((2WN7!BN7,LZUBYT/7P\0\5RVX
PXU?T29D,:MZE2VH][?3Z+;C$A_"JR4JV_\M[^5+2UC\ISJB-,"H,'Q]2!=A_V3+8
P8K@]FZ)](&,\W>AE#J<_E\\H=$.9^G*H-DRB$FI;8$KN[+(YKJ/I.>!1 #(UN(5.
PP0OF!.4 Y@88ZU-=O^=<#W6,8S82U2KWD(NK0Q;$39O9AZ*&B1KZ1*5U!^9DBF*I
PKG_RB97Z5.*C%CCM<'U/BL?:R0*I3[P:D-1)_!:BTA,[(/U*0AX"$/>)]2O-CNA2
PT701P0^#H]C7M<4PC9^SVT?5RQW;%9!2Z12?=BKZ\_ZX-P2&PC-GTCE5#74(0+Z4
P2):@15?3\XME4#[#Z$V9"M6$\]!_H(J-EF1/K'_G8+41DH-0'\H;GZ@F_0LM734#
PC/$U2BLK-$@9ME3D/%% O YI!)L/R,Z=,:1(9)NW3@$93$J]_,+[_H3;0 FM@B! 
PV>YLOVKT>+3/PNZ+$H\]%.)D>UT@,I7@&FHP-S6@]'_E[3^[TBOYQ7GM]Z;\LV<_
P+;>NTXKB>!K49$OS>ZQ'1H3""$?CI[:@PK]K=EH06UO\MHH/\-_5@",G3JB<^1NP
P9)MU]_X+D;E,*3N^Q\&JR@1K-#1G%10X;YE@$_0_]<#4Y9JB.*DH'7V5O%5.K,*7
P< ?@,^2\H4<2U=,EM/F9NE9GFZFG.>YR;:C[!V?$OQ^^9NYF#68\RFE4,"KG-F,,
PY*O_?O2H%V)I2C@:N-5D5@2/C'"O.1%GQM8:O=A3+;;:O*VK"S.K =!&)4[JQ9B)
PU!V#:X_2BR4EK1[J F+B2:2HHVSH"*'O(JI-P@YWJ>E'N/40/ZX<#M< QDEY8NF"
P]YOVVJ9F<*U^EYM"2Y+-+6SM[Z/)6F$HYF:$#%VFL:2/EQF #Z!1[<AYV;MIKJ.7
POZM4Z>:@XQ#J1L40[J7B?44B4_H1 X*S 7(9@'H$I;?3.=I?/&XG)$IC^^LI(J+R
PF7B,U=\KH4ZY#\(IH!8ANS'S.>W![T]VPB9?E8K=XVH!%4R$+,<33+!G!UJ\> K)
P9.^#V.C02,NN_OCN^JX.W2T+UWMS42>,"'NB9<M90!PB1 $LB5XLL&'6H'48YRD<
P'9;#5*L]K+O&_3+/U56<W*4^1S4/Z&2K?CYRAUD%)9&*&3 R7PHTV;X@F7)!B@3W
PE!B@B?HXGW) T4K@_K++AB/@Q*.XO<W\2"SEX!M<BL:H1_^"_U44(+05Q(0%E#,0
P;N-R-2<3^8%!K[!QD[YQDX_3O([3P87:/)?'-0MK4P,-Q7-&3X<R7="=<)OV;Q[!
P<\&7J?K:!5?@:YN,','9D-HCVZP#6M]4GC;\[[%*E3_A'"P1OA=.&['%^X/!V9GG
PH4%3AIH(;A!?CBO#W?_.D68GUS>AYX?0G=J @DD\E*"^( DI;H*T4&(YP3;6C&KK
PHHN^R9[3P!SY3 J"1IH 56.F4F"*2J%?,Y:4O>(.$93O:49LUE<%I-1R7:-A0R\U
P]B;*(A/-H%(';!/"/8@I<&;@R3C7DQJ) @$)?/87RL[!3"*1^ U(F1($ZE/\\ZU5
PS=Y"TQ6<]&TLU@71N[!&9W=>QCTF[<B<-!^AKO3'5ED\BWEM,T,8S[:FI;#<D>9@
P7(EEWU'711,\1$-"@GP4J$[QO-,>M"&B7.<)8B*G(#F9^X*JIX+H3>0+A<X3)A#Q
P@P$%X*SBB-PV"6""OTZA$/ N&L02R3" QK]:23(74)B4I%7!'S<JA*14J_GP]XN<
PT1BJT5!I]CG<$&\"(4[:_;I8$2K#Y4]%BAE.T!4K]Y8[%CO,@IGYP)S.7>4C83A_
PKYGA1D+%Y8"0<HE1^=,SWS+L'A+5#3*^;^; 1LRM_9Z[6ICD8,N?KWNXK>>RW2.+
PZ@54$XTU+[L7!_,7!PSO82NR04:!,#\1PCSW0\<RMF4:2<X?RPUU>[6L=)0N54*+
P?2!'T)L+&1:%D(;W=9RS%)<%9\S*\EXHMZ9V[/6DL'XJX5[@7\B"/[D$ZYBDX7#R
P [>\TF8V$N<P%D%ANN^W#AD:5TZG%C/T:+2Z2#8NB[ +4(SS;_M5@B:!16_HYEL8
PK>5EL*N0RR+(^L2A2D9U<1NN?[(M% GOS3D]1EB[18TZ-+MDRQZ 7;59IWV8QM)O
PAFLEB4CL"]?DA&!%4-E@K/M4H+71NZI&UZ5SGY"*DEOF#FLOP Y0#1"%&:Y14X0O
P?,N68X-6]^]2*;@M.Z%M^=FT+4WEC5&X2@FCNBIP@]NVZ-M6;?/[B6\9(C3;&C46
P5F$CJH0*GMQL\[1O^MTIF-M?2V?DJ@$]I9I (TBR^@GN!#V71)0,K(QH=,S&7?C1
P4T#S9.85!97>H1*QD(0/(^&@^LKZW/V!CB+('I&-1(%@O/JP^AYU[JQJ.U&\[-VD
PL>R_Z\_+Y!4JT^N$1=E\F<\QO*HOW.FZH97IFM)%R1E=>I D4R'<]F+'X) 77T&,
PN>-0HV/LEF%SNB4GSLAR&!J.6.RZJ#O9R=_;(X6TQGB>W:Y9AY;AH?AYG"9NZL@N
P@LJ=+"[&&UX5AJ$]>A%.].!\"VVJ56&7Y[,I0/33^LV5(?:2V1<ODGY)_2&O&7YD
PS30H6M%_%I1'D7/R!;EXMSS#PY'8/K,^%>6-N,]4;M*I8%A)_'Y%J.B<?@*S.O>&
P%&/O:TE(KUT:U 50]J'?L&I 0HB?7&PT+,35K]-VI6$^NBE"HN#)JO3K9AF$]@Z"
P\P56.K<^ZGN?-QY*H@[ SIH?Q_ *%PL8E5 W%,=!!B'I9+.5\+>!BG%G)H&0)SX3
P'AFD@E$;/)7Q\"0Q!1<T1ZZM32)?@I98;'GZQ'^Q<:A+N]?1Z$G$%0]#E/K6^P?\
P5HEII,KX \#BXGJ8J>,8&%&\>I"K/7KB]$R9EKV=U0[-+?DD@H.WXX(]+J:7?$U%
P$3;:])LF2X40X$BQD#OI="!+).[8CSW^97!,=_B7'9<WKH5;' [MKRZ#16MIL Q6
PT+Z7-#S2FYQ)GY_DK:I9VOWF,W-/SXE0[LZ@1P5QNVP'+5Z2A^7"FI9'5UES+;2-
PQ] ./WB;1M#]I:7&<G8B38\OG*!*MEX7KTXRR%B3ST+NK!12WNME<P"0+ 7(ZG5'
PD/I@R*G]H ]?J6J _8_->W+A70V"0[!5=L,G-C0U]YHQ:AV)%G@!U^0="</0#R\0
P24W!P N98&:6U^H@.\8J@3WVU&18C5CN;A;;;8\9=7(6V0FO,Y7FC^6>(2V9?KIG
PJ#B^TN?9C>8$<I_Y%M_"/W+69JSA*W_U:XAI %HB78M,SB_'Q(<L>W^GK]L.<$'P
P?;LUL'@:G'UR!1_-R%%!Q!CE</VDY+MYW];!7(LI<2\8)/X"I#9O<N8CFV9DZV"(
PAVT?L'V5AE(IS)Q:H5AD:,YX1#H9?"+>/W14!V/4,^S=*"S2FR;[%?(O2;)-.CF\
P('CY1FIK$5X>>!JYGVVJ2FL.02"[&<]Q,58?RG1#+3A]W5#Q;3V78Z+8J5^W48/T
P5&1L*IJ:J>_5S5&Z (E&R0R2J;G(CQ3M;*/FX$V5*]QB[*<K)NE@WX^X:$R$7!OX
P::WZ![K%"]*S7O$(="<D/[A;%>!)^=3\NN#[MNU/70.&A9<ETC!.M6 LH*-Z_ZW9
P_*R)!6+LI'@7V:XEQ=OBDIX)H$"Z4S@0\6E/2>-HO(!05AES]3Y !$N^N&#VD-)L
P?/.+M3!'OK8<"49:RLPC\\&EN-O[@_[*%<!*I?5X34[:5LR/=J#O!3;)7M4<@?E!
PZJ\-3I-I#TR$,J'7S&\3^PIX#.T[E>@7^'PBI]DKA(9=4+NW*(P$0GQO3*V=--;K
PKD31^8V/%9S\V2W"###%;T#-SH:7FG_&SHJ!;'_M+\^]%$>22M&D'Z7JM#V(L482
P'YRLO,D+>A+ZN8>?#VGK_ZJC=$NVJ:!HC*1+M897$)TZZ SP24^!!?96T0E( Z!!
P)78W*U&%+YQ4&^4:0_?2$AH.6OO@ R_P2H/31#4G=A%-E?9PWTA/.,4R^6]],V:#
PFLM7X)7;+@X"&&9V.2&D\?8%;S.?,P]Z6#6U'TI@B[$Z9/O;[9 0"WS/S[NH6P^F
PGAX3>GUF87<)',KY=%=WY/54&DZ6S#(\*GPGIA#'N_7)S)J4?B-!_!.G*<V=!R]%
P)(K]*K^N.6_\GST8'&Q?G[_6\0;^WW1O$2N *]8X5K^K@%LE]U:J6;MN;U"_?Q+U
P]P7R>-7QU)* 6IB<Y#/(8H_\P*FA+6>>&;)@UY5+%?FBZX8X4_?,?9B/,9ZU\.4W
P?!^VV]1-IS]%2=PHDAD7Z>J6\3&4\)2A<,X,P0XDW<TYBC-_'Z(H<P2[#-[DKMW/
P$)QR*W=+%/X;82&DO8;*WFE>[5,44/D!CNG), ;=_N:C3X;9& $#C#.!%->Q?E*.
PSA[:ZZC/K_' T(>CQXV@,\=#X&@7+73&"MD7XB@T(^A!,J#6L:']M)76? +6GTH;
PM,LGW#G*' \K]AI^+^S>GV,(=W3N1WQR-+Z'?$AS6*$!Q)R?Q]G[.@S1KN$/U:;\
P7A8R]8+,9*_"#$PHSRH)0PIC*L>FQ@7"F'D&917%I6J*EF#YF@-5J$G6CC\^6)61
P6[R@0P<*9E$.;!9B-!M'BLP 0 [Y4DC+59L'8 J='M/36K=($'/4%D$1'FL5Z)&?
PJ=QI".BE%.4NI"VH_L<?T"/OK:N]U? \AG5N<K/P:?3*[QJ&;F);+9>X_*2<(T2@
PJB]W2S\%3#216R&5#Y]A[UP?Q 87P^*=4H/1\P5;W:0V2!;AQ1$;GUJ%/CM_^!]4
PO<8!=)N/ XTJMJDEG%@:%:^+>+HDO -?<)JL<=<%=)7%1BBMBD)?1ULJM*:)>)FZ
P>Q77-\2FTS)D$UTZ#O<7C0B^E!*]SR>XFB*:"/;Q^WY?)L& DR\4'76>J(\-0)G 
P<]99A?D0S_\58]Z*^H#9UP^R]SLIIF7)Z(PG7CTV/_^=<+N6&EBQ++CE$<_$\#F9
PY.$YG-V*3R0^0C?9?S!<-IN-.XL6D:IGG?_:M3X8".8&XC 6X%V^ Q@K.;_]I3>5
PEL"%(7>UI(;+?F)E)BV]T8F%[@U-=-4ROC7KBPJV#0]5.1Q+0@MT<!YN?C8._;T=
P(M T#[JBM0;NL,1Q:5,+CA519*NM5099$6]2 EWH0W6NT)A3<+4+ZC?[;F6B'LC2
P4WS&UW9N3F7[N!7_TD4W>\LS"V#OW\XX]^[A'J$DM5)7'CU*QE!:V@\Q:SHKH=BG
P1-NQ"+9).'/],5J;NEUU?T;0"61PT9/9YYA)<L^G,ZT^1OE-'B7'&#!QU'%R8QZ_
P:FQS8SK_]?C5BW"M5(_%>R+3\?[W]RF<;,0*--RG/I(M.S]/_MS IC!#8-!/C^G:
P4>V:.V.UK&:)AK('LH_#C:VH\)29P'=\/VKYAPT(X7?J#/9$,9[QFV3(5;!T&/Q5
P[$3I?3T<U!R_L=M51.:E.!0QRNLT)Y:W'K$SU5NXB/^[S9T7.;H#MOYP]IY0%$SR
PR'05,,?Z%FMCUQ'"V.,>7$@Z [1]U]G,RVDJ6%^)9Y&J!YS\/S%A/ DN:!9I\-VR
PO6G4R!37W9_.XQ?CS($EH/J [\6[3A:^(!;XHT"0J/9DA#5L15S<XAV^)F%@_W!@
P695R*+%$*.,S!LR&N<AU\Z@%/A<54M(UNV0S2::P\?M78=N,>+T>A[HX+I!\E(=B
PD/6:ZB[K!,0X>$"T8&.*64R*%!PJ(5=2Z@BP4/C8J2Y_Q,("9<G+/;@'4,T\0GOU
PUI"G%M:.J< IHP;',R@\QAM(6:"F-X'K!AL'PH=_,D D(@D5;+>#<V;83Z;<BI)K
P*_?$3>P^7J1G#1DW^M2>/J9!^)GHHAWID4%#T)64I<#.34]\I4W-0A%GR+XW$>9H
PO@[GGU"Y%B_@FVJ'8L?<6WD&HI;]7X1'JY#SPKPVZE;M.56 (!-]\($94C4" E+Z
PB,HY'I&;T*H+>M;,&_"A[/\.M4VKDM15KZ,]-B<S2XC^M^).G&G4/<%3ZT]2,?HI
P88%GN7U*4X.TA8B]<!8F5;UV$7QM2KOE][@.-Y+AT4V[W\LFW@_1GA)040N*#4@A
P(V#6RQ\?X.V'BG)'W*NVH>99:<(CQ,%.:;8,/9.5;Q$*+_27A!5NQ!N," OV>B#%
P&DCO(J"SOU7UR;MLJ%^'9HHX;2)??_]N&VY;;ZA(8T\FZ%#W=XL^=K%N'0SSRM>E
P6#'-1 'F YBEXW#Q0J2M*//!/_5IA*6=I[NA4?L[N_XDMS? BV$U4G)0?"Z_Q'<N
P6)O;-?FW".BDK5%NX=V3$WMS*2T ZN-U6 L2,36T'Z[:><#6$<U&*<3NIB-+@KU]
P)^*(DCE@_GIZ$HS.*ZRF[ ._G8K#H616&Z9O)=X''SR1&C0DLP.W+@9+R8F)4]'@
PE#_[I/6OM\ @B,DY_DCQ1WFUP^(XZ!1#C,*  ]96KZMO2JW97!>_O4"=1(,'JIBV
P]FS.D/]5?4:M2#3W>,L9;]P"M,NJ%_,<G!)E$\PP37 [O \ >)G=30D=%]J+#[5U
P6OJ#GQW-\\NZT.] (3.XQ=CNL*!UY/&H<4KBH8$K3646'+HN>( HM._6I"B(":DA
PA1'"%$* LND^0]6+<,%"M&@=XG!P2K[7^>=2CW]+>EFZ**7<H&_A03V"7M7;,P1T
P1T 70CFME%*?=$O#!7F$N,P%G\7L6$EPZX*(<4MS= O68$-.3MSZ]*Q&^(GECP#B
PUY*M*F"I=?%><:C&1S%*5.(BE%*/).9(3W[ HF\SCN;J+]P1I3JAV-B<$&\K*JE1
P5^]X:#CWXC"3-&E:3L*HY0&9S.G?2333]]KR;NTDL.09J87N4= L#^20CM246!OS
PPG4&HR:J.*@@YMXXD=>]_I03@M>9;]" FP8%O8MGO;7Z6"/Z%RQGT@43=&:_!WY7
P>:%8V[E-2C^N/]XDDP$(-5F*DXZQ<:CUV7OQ,42B?+%-BMGU/[V7;"*OP\4TQ0?@
PD:EC0A_A'VNBKZ3E,^ODEU@F>M8RYS+QJC353Q2 =GA^I5L9<S'\<_EX'T]F.H2@
PQ95T3[IQ^@1;A)^&S,P$^"O;)[,6'I:>XWP]$86L%!(I2T4],I[B+'9N KWJHA?<
P50$+&&9=/(NI8!P&U1%A]WCLGWQ"RDZ\R5?)4TG1;S3\2-.N15B^B!^]O\QI:L]=
PJSZSD-*H>$*^%H,2)TT\D8XDG[LY/\X^1R-5GQS,-3U!AV#@G[S5^R(@)V&6W][$
P$OCD^S,]KP7%$Q[:)R)>U$#OGX8Q[^$L[7=#&FEO?1/,&L\#@'^A+_RAPZ+ Q6=$
P:8+=V%[7C6OK^J_+G"U3?[FS:%LY$%O/^7@DRIA)\?_6((J:CP&'J-R^OEACEI<\
PSA!D+':P@[6]S_E@\&Z2/V?T+(#$/F,ALSJXOPE$I7_O<)!XGXJ<[LAJ<-.9KWQY
P.#HF"(TM8" \6?'>NR: ,NH(0>FG/+CZ6&:'?NN*RWO'Q=L0N5L)6FB-ZWFDCF6=
P4*V;7:7OR6X88S&>\>H$>TV#^;_]1/-LOSYM&,Q+0KA!+BH?\[E)98A&VW0Z<7K2
P^O[R>P4]P23^'EKZYGDG_7()[NSVM69970\X#;;ZLA,#I/CB<+8V-K^<6DZRQH/I
PA*]_,K(3*:YY3_9UK:L_)]]ZG)/T$%-;(ABO@$HH8HJ+9;Q>]>C\2RCRF(?[5]>S
PHNU4G^"!QYC.17J)A2JB* N&I>\R2[O*\?XNA35] 1#"E>B+6UV:;0:CBN]WZWP)
PRQ9,Z1_77PF,=9UG)L#VM.^6 +F-?FV1<U''V"@@@-4FD'B@KP_392-OS%K9NWN^
P'XM^WH9A]<]9_2.57<:#R:U9.QE[JT+9F+4()Y"9 I1_9C(CGRSIP@1:9#6F]H(?
PDO)2X3G+Q^.<>!PPU5DR# *_%O%C[[ 1 ,*PWWPG ^2W&E!MF4&X>>O4J1<5-O\)
PQOO?V9LW]WO<7SVAA^ %ES5 AQ2H<L=LR[%LY3 X,[#!)3R<<<;E:1:*NS4-E5?0
PR$_EZK(&5_(EKD-0?I)E,5.5OSG.][04KG+?UPT$#2.TFK5 ?+7UTCK]-!$"+@Z9
P>3[P\$I1E&1ZKT/X#!]A35NU*<HHW;N,=)2_@B/)H.71GGQ;LL#50D8OL,U-/UP6
P5O-(C&HF@O3/I$V$9C2E3O %WS@8:GP$F*T:6!$=D\IN#6<J;?@3E/$PRE5(_A5<
P5L;Y&M6 P2G:R,KA$!]H?AR';]4DDEY"6*/-J9.=KULQ12^9:;97L_GKH(QTT4XE
PK $5*O*&SE/C/NL)U:1>\<<+[Y[KPH#^A<O5*AWNV/3> UH)IU:K-A]T[0H3"5$/
P3:*;';/*/Q#A5FZP*1_H9=-S,1BN3,71[MO,8M0._9V?*I*E=7%H2Y3O<BN.EQE;
P."KK@%SK9 6/X3V^JR505%*+3]ZV'_^1=0N"K 7'P3Y\\6PCA$=\E+VI*L''KZA>
PXZ2FPW+AD^.1W#$OGEA3F7:MY]@@E&,9%&/E#\T&7?FN)<N]B(FWX%;&K[Z)52G_
PQR7L>V52F+$Q0EVQ4*,HEDU\VA-L]DN56E.N\DIPBLE8L#$I)HL_OS2U3*0?[^@E
PWK.H'NOB[?!X#]@8!1JBTCYX[94*V X34-2A3_W+%V-Q)8*:9*4"/9OLNJG<A(DY
P,T9+\NS&"?>^8,+(6G$@2R!?]I.F_=/VP9MI(FB'-6:&'(UN<M6(\NR+<PH@:4L$
P<G*@8@+KX=ANO"<Y'Z&YUJ;;X-W[1A Z"V&RDW=4\&Z7&IOK(IMUB<Y96QGKKX!O
PP:!Z2^>,GO3!]]I[K*HE4-<N.YFG;S3!]S$T\_"&9)=.YX2&H[)JXP*/FI\9C:N@
PYIW)<"0MCI)<E@.Y.20IB(%U@(5+OX]"T-;CV&M\2S86>2;!:QU+&RX_L\D EKMX
P@USGHZC"=79PUJTGD*/8T$N+%$SSUF'M(<;P L87+D8H\2!0P1XQ2V=3A#U<J2/8
P7XX\VI"15YSJJ[=*T=I/_9B*Q4 WDV34J$(VRX<)ZG]_$?N.6RN]ZL-DI+Y[KS_R
P.S^!U/3B%G_F^7Y=B^7"8YZ(QW'!I'<68_7Z0+Q,(HCE<#C4R77#6\BI)I,D^V-G
P25_63$[9L>?VTX^#+I'=M3[EML9B,R5B/\:PG9F9/:><&* BUH2IR[+((;V54;81
PD3!7''C,5RQ<XW10;ZQ#1_<1H*C@ OZ'C^J*TW/4M;!N/_AC+MF584MV>U:OXZ+G
PF94G#&(4TM\R9>&42,_>RKMN;CZ#<I@"X0EYW 1"B+^.H,$%U$TO(9X>326TRU\?
PH@ET6&>M@_."6VET/L*7:\N(&VV>A'C_0A/BXRI18%A)6AW/P/I_7P,N\1S)V?;"
PBG!B2/PGQZ9PMOK%=)"KVT1?I0+!0^32^KGKC,SBU&'P%RQXO]I&^UE\)*'68<K4
PU;J5.7Y]<2P#@R<$&Z$-OK;ZS7*L);UNDKY(;DS]ZPC)AB%66OSL&_5DBSPT8,D0
P9>[AS7H4O$BE.$U5$&UQH5)XEA5Q@;E)G;L&E;4,<0A*2ZI;V3M&BT34@\WO*3)8
PC<LQ[OV/+_K"@T\G"%NE^V:AV4 G:\2[QW-ZZ-TQG#[&K1XU^7;=7E%IWT$<=&/=
PI$I,\8$E5_=5Q[O_N!DUS@81 W3]:X#*XKHD9,YL@R-V^W_\_CSM7>*W*ZCZTK+T
P3HW+:8C9@\+CHREM_K2;9=']"53FP!5ZUUZ(:$E*^GH<AX[MNJQ(UN1-"W[TKKB4
P6&>VQ4<H^43\/AYU/"U\D3ZB-I[(^$8(/-]]?C-B6J9!3;,@"UKTQ@H=/RRIZBQ@
P0C&Q&BE!"]%AU6=K>Q)HUB_P^1EM-4=H&E1Z6*#;<Y-OOA@D7Q?6]"UC3H 9XF-'
P+.X("U$^H;@U=/VZ=>]JHD6A9!EDGU"Y_-Z6RRQATV9&FZ&CE;@Z1XH<1\(=RD./
P#AU'[2K7P@R^V6_^#6E<7$19A*M;N\@/&M<X)/*^"&TU1@7YD5UJH+R"EVT13X(5
P^>F@.$IO6; 7N$0-@HDF/,+Q,3PHO';N? M ZW:II,9'8<NS#W!LUB="6L:O/H24
PZ6YMN@L;K-;:31=G:P2#6;EIU:]*2O)QGW$E_!3HO6F;JEW,F\-%H1:I"$I,;[<M
P=0'AT;1+=G;AX-D:>*2-_!4^Z8O4ID"F!Q_JAFE/"9.4/V@OUVQWK8\ED<G/#AA"
P@)L)CO&ANDM;*7;P*1;YSU7Q;1FLL4&5MC+5JK5K;"G8G0!84@A<*:#X!O4'J"]'
P>3_+SU,S@!JL156C=(* ="ERM<1> -VF')M%9$5ON(01;OG7WAC'EEM?>E5E7L"V
P"O&CF! MF\&B^I@;0D/BJT79L;^HE?JJT_3=!\DSV9\!T/G9[#&Y8Y]Y) /[LP?N
PC=NE2>[@[$E28B>!E#5@>_EZX;7U/,"4Z$:^PD_@:4=!_:,\F$Z[58T;%=P=)-D"
P,/X9'J?Y;.>PSSZ)OFPZ 0;S!Q6C)MS- YU#?9+W-6G1['D?KTT+>C?L@V_EYMJ:
P6JX\R$[991($H;&:H%0BG3[C#?!7_P12OKD#V5O7$/^'47$8Q0/@Z#$M6L"/U W?
P!+"(48@BLFZ]M_O,>69IX)#GUN<G*"%G^RI+V*56<H#:Z&EUP"%D]$RNY2$G!@,1
P"MB_][3Y^/_9,4V%+AA$7VF-R!H40\VUR<N1(R)T?T<.0MK# ?P!IJ4GHX3G5)NO
PF]YHDWP>J6AE'Z=5R[Y7G*[9><!X>V8WE)T?[P/$"0?K];(;Z83S+[P7\HI'^(T3
PFYV[E0#OPGI'-+[%5/)&$);ELY#S<WAX9ND[S!8!^V?4/C&6SMA33TB%'X?K6]UK
P+B,]/65 4T[#.WENRK,8MEMX1\FJI>-VLOU[PV )'6G'VP-B=U,.6/"-%@OLFV^T
PS+&Y^X[;8*O[R#Y;O[1'H_9^^4/%;.K[9#F@_J(,II:'>N7JVPU5=5EI^:G8J1<&
P>S!J&.;[E7@H5LMY'5UT&;\9LWG<[#.]%KIR0G^TJ3KE'O14:1/A.'I1:8[REAH"
P2LKY9ACK6 4LFFS.C_ #?F4^1 =WP<_\(6_Z"2@]3DE$1RD,)MX2(/O44N3P>#K[
PP*X*7"[VQQ?V]G,H0EL[HU\BC_PL8IZ6$!2&95#R(/!QQL@54OX"=AE '0<$'$;D
P?:]I!@,Y/NISM,_'#(!T:LDD+'UJ7'L$2VDVQI[9,$>67URBZPOPOLAJ26MZ-<:W
PPPMO$D*QBIF?03LAW(7@<#(+JK4NYD(H7X\OO:6 :>.K5%U2M!L AX/>_Y<LH7XP
P[,P557>[6.':XUMMLPA_&0KM-;P+8DN1WO5.C(]*K?J@"3+[>B<=#Q6*Y =/A!2F
P/;LG\_;U\ <;$D-S1%WM16Z#V.Q*<K/=0 I"8#G*==A^ST, (Z$U?^#7HR3#I:\(
P,A2SQS=&=+Q"*E$G?-/LH"[]QLU_"/C_*>@6.?C))K^7( U9KMJI,[7M'S3$;-_%
PQPT=Q!(T5YJ? XOF$I?@K,G@HW3"Q""[HP\N):>9^T.BYXZUJ _=^T%01*C&.7@^
PX2=:.U;XF#K3)-%J8QA&A)0IM1CKU%8I<JI+:NX=I&M;K#7EVAU!C3_1/H7V:NWQ
P90+Q*>/AW'/:/0=X5 N4CE]T'I05DRJ]"*'-<]L<">< _=5"<Z+SKVRQ:MC5@V<C
PD&@7H*A!,N=1=2IPF4*4.++B+]=[^OI7U2KE7Y ;&XOB6Z+!6.<<G\AF^H_EK+\J
PKH?7BW:IL#]ZX>S%2M><5"?_G:=4V)W/HDL('2@7U=WHCAI7>WY@M9?)P@CLK:A$
P/.*LT2DQ4JK)GZ,W16/<>Y_[)L2K\A>S_6F@=*9@,;#1JO8+SC9@Z^(^Q_V;52O0
PH@BNG@:0(O9"27ZGN_NK-1@W"0Z]UFB@&Q>53DN/S_<T6^11-P6V8>CR33L)5=I>
P+3,A+&B8J;%4^HDK$^S8:.^*::*@<CS,_]KGZUP"W^2M@\" (\$NJ^>+B>N.R^[J
P&P73I16E[6TBXP) 2T@62E?.U<O=C_<WNR9/#&Y@"5&"%W(WJ<]12MDW%R15V2?8
PTO-2I2W10]YCOR1<#74$H)#)8/OQB][4L7;Z46]<TVX2:]=LH-D2]]?#><BOU\F]
P@GYWY&*S&5V"_0NR7-&M?I%0*3EU()D&CBQ+"\T$7JAS%91$L=T6N2' @H==!;P+
PP H5]DP#><N*HR!-.KU SR\\L$H]C(DB=R9_0P4]/'V#]?UWRH]6+K8AR57(GSF5
PL,P:+7>[59S\><X1G;;94#P,OKC'Y@#;DI.X,^*X.+D491<M'&J R@44D2B#3P&J
P^5WKR1P]W75J[51E[OJD2AH?DFH. @)SQ[0S1'G13FMQ:R4>9*<MZ3QD$E-%19,L
PC7/8:6GR2.B#J(*1SVI1G:67(&7N:^UZ#Q+TG/D_O62$KN!;I??X=4V%J,48<8SE
P[[JUBTIH+A")M<P#)ZP"1BE<ZO7HZ">@7/U^'I*5J\J<]7!H0..KZ,0U27M0PT0Y
PK:H^MS;_$/'C,XQ 7ZH+\.YQ6L?Z&0V=)"+0+I_/(2Z65&*J\!K?^[Z+S<6#&^9K
PM:V:X-FIK@?B78-V:";MF!'K;./CE1RH+2'9MZ-LPU@45$HL"%BR,$0OB"SCNI6O
P7NNBE-KA\I@FV^,\(4S^(];>94K1M=\-1IRN8_<,1CU]5D76&A?3%.6P[!.SW_M5
P)9(EPF6RDU\Z0F_/4#ZZZ1(*O='OJ+:,P0W\E%K;?OVM_B0K@_25<33.=#C0G]BH
PU-&11_J"U)<.W_3J@0E^T]+.H633-RV_#4&YP@_;^U]O/TUT$]V3U*K.CZ&X:93!
PIC(]=<P1WD' ^G%4("N/#0[&XR^2Q3 Z?WV7]LXE08ID\$*EO@36S$>OW>M?_JGV
P6^-F>$0*"1A+J'Q1G7FS0N!MW&=1YD%C<]0Z_;A41.M_SX=7?#F=&\=[1/*+-8/L
P.CVJ1FR8#YRUW>J)Z63VWV36(=#OK&18,+J(XS;]%/Y'DS[P9]_>'X/%&0!_/?&]
P2 :+'9"U#"*^7.*<*"6+I=PF"B,O'O>CO)8Y^<J!#B_F$1=>+LQLF"TR[TIEV^EB
P*HH)4I=\FF/R@:T(-+-VS#FXL$+ D;:F2N".UZ8LQ*M9!+P/D]NO(EI (WO--V+G
P0F')_?+%[#+%TIF/+RR2._OC#R1=F5TJLL=-8FD N96'/:Y3K3O+'+RZ]C6-U-HO
PG'X1F.0DX!S]/R]C>=F8XK?M*?/S/.;D.^09>9_=A.\L=MFUX+[B:BF_D>G4@FT 
P&!/3UW7^IXXB!:%8FF!>;[;(I&\ =+%S>WMP<D@&!@;L@9<1'[&"_HL;?&>L)LT:
PBOU+]G?9WT^[J43Z7R+FW"^G+NR9)^T7?1I5B37N2_-<(&Q=P9@6AW(!80.040&&
P"(JP00.Z_@()/=;#TB!GNVGK_L$N^-2[H4#LGI#-RV2K=>49E)Y'D F^0FG/Z93Z
PZ!=@@@*\V:$"2U ,"*&?" X1,ZN!,80R&"_^C\Y%A-M!MG):'#3WZQ#G_)UX)389
PX@T.G<K>TD7<L/8@5D$*<M,H'G'/4#CYM?"@0>4UW?,2P3IK]GF^/42XU:Z2\[UX
PU^[X/:EPNJUB@L2E,8_G(73X!/_31Z;E0@F334LZ5>LUZ^22OF5DS [\S=1OI4Q2
P1DS!WL],7U@SIAZ7EYC1BUL&!1MBFNJ);X)=_HMXS9\[87:N.>PM@'_'\BY=]N.7
P&!@:OV0>K+NLD7 -^-_T_4MD;\\(4X^AA&^A)#YDR[ :!F@PVD?GZB[KH,YT5X=[
P]:QEB(5R5=N'Q6*!H?AC1P5U#VL-F:  #\JT(#"36FJ '@&V.EF8Q]5T6<R"IN6M
P&,.[M.^/ [_-3%:GVK&)KWVT;5R(1W];"??XU*_\F_0O&J&?EQ)B8@]N@)7A#:K\
P3H,5KY[D[UY(L^[T1,HT]E&'ZIN+<1V3'6A82)GW]K]U#EY+F@K]V  NME9'.<V_
P.'Z!MY9]!:,RQ(.;,%5016NXBU"COH7[C5T9M_+]2I3]>C4ZDGR6,+E*ZE'VN$_F
POETG0;IO6<_;!;<S1%2V'(6AB\+_G@BF\P[4E_.ULS.HW.&8I@3)->JD<ATS7RP"
PD97(W"'>NH(Q8%.36\E5Q<*QUS[(Q,<]*_!4$)*.PI4_^IJZL80#W.MYN*IO_ >X
PBH1DEL10CQ)U\-I5O=:$#>-N&!,]JO>*HZ3BP/3 >CR0YX?Y/]Y; L))[@K'G'3Z
P(WLZB;*=?+W$[AJ[-K,JS]CBZOSRVCICPU7SI"55#/W1'E[+K(9)DPJ9^QR;N)_2
P$EN-!["5F<\M4";_@T$_=P%VCC#HZ14UJGU2<2"-U5"\TB:7U;<+\M>^*HLC5^UP
P:F-JK"4W!"&:X*DI[[X-925P[5#G+]!98Y@^KI96N)C;_/R<+N4M+Y(KVCE7W(6>
PC)LE!_JA9/HG^G<NRC1%!;7^ZA*K[7=X0WH)]SGB)FOAJ^(WSUU%96P95J/&/AXG
PW',YI5V'KS\=F>38MG1QGOJ@V)W39SRQZ:#S-; %G;]]4!T9 M0NI"KL#<"]9#)*
PI!1VK==NE1JW]7&WG 99:6]*)THP7B X>"38&,]HD!5X8CWXM Y#'L!AN.4NTD+E
P9?S@VX[J+1?*9 6?"TN]__V8 /'D*K ;?AG@U:17S*:$^&#C)YP1'$-"-4D,O^F!
P['*.)?IGJC.\EIP$9CKY5)8*MI"$%OEDUJ!-:7HM;:8Z=5D;>L"S C9PDW]67@F5
P^;VB.=94(:#,.?+E6=O]A5<XU27'M--X, _[!RQ#IZ\WBS9&M8@[+UW4NGX$JE#;
POSLNWT0*U:]#CEC2":61S+PI4<@S;CW2?OB=0&9,7:(SL2NF2:*JUU,8&J2$PA)P
P3]FHPZ3WRN$?<6?*A4+$5.EZ&E<GKAJ%H2E!=DY5T.F9&_4BDP*ME"/H_"@["1G'
PPN@-U!@=^"85?2SI?6+AYW6^*V= L/NX=QO%Q\Q3YYZ!,.KW#&/BD6CX\)M%]4;@
P]=V.E5I/P[X B<XR%8OV\33_QAW%7%GRK7A^V@<H(@/7FNN#.R=H#Z>#N07,K8*X
P4U^T^N"A"1-/(\?T=H"]D<M_R^@_C?6WC#LRS9]L"8BB8W=N@%1]<(#FVO ; Z=*
P2L!_/!* *_P<4AMS]TQ,L>>^$3'2^'!BA9\RE^#+ #-^HY)5N"XO.&U<)B7+GVI+
PH E@AD'NRY\ANUBDU[B4%+$NGW>_A@H=\UN>LFRY J"C&'_G62HG'U&0*^...M9W
P-C'#*Z^\H_A0B%R]VJI/G*VCZ!HXT]'1Z68&LI3H),[B53M;$OLHG3Z8G\<1,:6$
P*7_QNN#X_2+[+O/7'S"MOQ56*_%>2)ZX*O"8P6OJ["]1!9A([?XPAC2*W7'ODIHL
P".^V)64R(P*Y%+L9Y;GDF M+?[U]5/_8W0@Q0<C3B@Y[4*>*C4<C@)<F)@N$BIFG
PNQ25+K@_$^%<Y^=(B@$WOR#)6Q6L1 3G4Z!))2F=4]/9F<"8)IU_3.)Q' CWC5^%
P\\DL4+\"\',7,I:OO[?I69#8$@ME?R&@,YG](#9<]5#2LFNVF=YD_GLHD-V&J>]W
PMHD?\1&B"W>=IV 0T?+8+XPHS^,%*SHI\=1!A6/Q3L976FJ^.UL6JRP900IC:=]C
P]LY&"QHR$N;SFKSQG%SP[0?/Y*_-[!G#$OW!7@1DM%0U0(5.,#MV_'Q@QP;Y_$J)
P;%^<7DF0#*:55\NE< $J<(6.3:C-Y(2?K)M64P5[WZ>'R<RI\CUMK):)'N1V><.F
P30D;"Y'5? _++0%5>@J)Q%_3*?7]&7-M!6\GJ$;$&%T5=K57FK'?(E3*?.!";YJ'
P"4X; 0N85-L_\P*#0.,9P^+3"VQLDMWCW]F/9$'GR'N!.5@QZOQ^X 7OA9%56@P\
P]5HZ1JE3 VBE+%C;+<IZ=HL=2Z"'\.M^W_<DIB!!]!W6W<%#%BBF=T90(D8T4BD,
P"Z_8N&)U($5XE^ =:S66O$X+/6+I_  N@N;9(_?<OSG+U?_F^#),7+N24<8K'@7W
P_FBG_'="WKNJ1-2WG?!35UA:X;:3*8\&M,@%U[&VT0H86'C[E.6@K))HB;MFV0T@
P1(P$Y=)<M/8B.I*U[HV2[;ZDY)1+U+J&/MX-U[U'PN 3*=ZHF/AI22)FS+@3[U8Y
PU2._8"(]<EXR!W@[V9<S[3@9U)[R!3C)LU#:8]X5V5C]YF W&S.GRH."Q^WVN_55
P<V-<_3#]!!^),_\MV;KK.5/O9I]!V%WA0TW3PH2:M>I"8L?+T2RZ[A5"L4HMQYV)
P%7,?@H+05'XRN:"70HL98[#$6O+8#7&/X&L *1K?4'240HXJW:BXC>ZR6V#,  19
PW7.Q1=3$"ZS*O[_L@0J^+'B_?P40HDBUL0#W<MO<X*OW-B;E7_Z]!;QO6LNMZ*1X
PR,[_RY8GV75G5RE:3@QUOACV$%F:;HH%IU&_J,4[?R.A$L ^(\]6ZQR\NNJ&=I^&
P<'/EZG*^C*\:U]3-?F- %2G3V!G&5.#4^_VZ=>A9TR=%:VN#D^,''\,:M8B]&T3$
PAQ3(B*\62RRA/OP0_9'SES, 1B%1!%_O6:5K5:,LZ+TC$IG><>/<&<GPZ9]>R]U#
P;)I9. GEH&[X] NK&B6,C$P(@8LU*Z& W^$_2P[:,.3/A*68 I2Q!I*'? KYB"5'
P"F0,8H=S(8[W?XT Y="E/4B2V;VF+-UDB=\?9B]3UTM0F0'1$"P1!_J0U/RP1ZFH
P^;GB=YD6@4]-__^6IPH)P>UH;1AU:]D;SO@#I([%&5Y1EZ:3)OZ:J_N-O6ANE'#)
PINO9YBKAK#LN8HSE?)5,1'5',.&_G-E5)K#JC^,A6 91OI%99G<?B],2%G(!S7E/
P31*/"?3/16"-OB_LN-%U!0'?RTIV:#]>Q=9_2]83;(!X@/O:8LQW7V=5R92PA#5L
PN# #U=42H0D(,2H]Y)L8JA?="_'&.>A]=E\!K=?'$NK(?Z4;MCF!;L27=M(.V4$#
PI.7$C 9;]Q4]V G"/'WV0T65%G=.0."J,ZP**IP<G[2>QIR]"\TO0#7W@7^J+*)(
POL20QYB0$X_1F$)K6#RW #EXYB\!CA_>L>W\ =P?Y/(=K[I@Q)@3#K"+-1\$B&6/
P%F&-Z=.Q6!DO[^C;Z6-<!]KX:0%(\:&43]TX@965QM ?*[^+?];Q<.DX( 0%]5A6
PG>WXK'2MJ=H]I:ZI.(,';ESJ<XVVST&/Q-6@*38VRT[]09A"]I=\AZ+;G^>!6VJK
P5NL(523@C.;(>$GL?C,IFK8H@ H($)T.0;GP2/ 8L'8&(PB 03Q..1!E48.!(^5Q
P$669$!%WV\[57@!2A;-B>]846GUP E K$!C'M'Q[-N@BMM]YD!RPR\BDW7];/>0,
PL8^M@1U(#Q> 8V:G1?5\@ O2_\1I2V<.^00!3EWE;48UF6\DQHA0B*(#S4CV0BW*
PEE--,UOO-BQRI,GQP0)Z81U=<6(0L\LQI#'^^XX9078X4 I+NYXPP=(C#F:E)%^I
PFD!&<!2B5)08J08_WL1* "FGAW'S(DJV1M3+#V1F1YAL$%;-L=[*8M2;%-/)R^Q>
PZ2-#J=)^:-3F1B^X><#X\7&;^28O2C*A\XD+PVR_T>KJ)CSZZ%!PB1GS?G#>Y$LY
P@.PWG*>4L'1F-U>^$K?^4_<^DH$.P#R_@<UQ.X7F\* D<4W>X=3X'6H[UUY6:@>(
P#; KEB+N!'J</&;Z0"B##_CX7'^&L6DD;2O1E=_?$BF+B1L3O: H ,18YR]\"<J]
P^Z33Z,MQ"WRS59+L1U1$2>I+_&7N]K+.;]/!IW] 78IFBOOC0W/P"=I6NE\**B;Z
PRE4K(W$)+T[. %P)/8V,B/=I$I-\ 1&J^]9%'^/NM.@N7^N*IG'>!'8Y<9(C@#X(
PJW93'"BE(WWY(XU9$SC0<2R\1D%11ZKL=X]Y._A*GFI+UN<5'K;)%?5L4"%7D$FC
P/>%N'N^9SR$J_N9'VP5Z<U_8L?/V^Z6Z$"3*@.!L,JDBW-"/7J&=8I_L)7S$4;SV
PQ.R1D4F]=2 =$RN:Z2>]#Y*[6(B\N/3!2:8<-@("7(8;>%W*:(SNX&4!H+T\E40 
PY-XO3/+1AHDHE_4:U^K3--4-ZM6O@< <_-8G9!_S01IOF6:3$\<!+CQ[T.K/5E2W
P WI)IE6O:W*[^DFLOUVC@BT5S!JIVHFDV/)Z/3 6@&]=A =%^5YDFP#QL1IILM1G
PRVNL-W 5.SS[I;L<E01Y1L!$%6H26A[DU6!#4U]P%+EE+ KWV64]^B<3>E\T%F',
P:C$U'!"1*3(R<X)]#Q$!(EYFT:3@/%3F;0*(JPAIVTJZ0A7=WHCY-KHKN_T8EZEJ
PSYE#0V^9SG>M"K%YJ5L*8<2@Z;NA/U248W[O_Y:;?M <*O]5;Z'@*<S2+ TGJB)7
P^-J_2ODI0YJ,1AEZ'PO^ IPU6H9)%#X,M&=PP['"9HU]1(+1E<<3'?7:K*R4-#VR
P*_87:;].IO]G-'XF$XFY8<_-Q:&P[S67]Y1.D8R##12G4S[I%SY41%=CI"T;:\<T
PC\VUHP'A/IU%@PTQN%&\T%WVO" ?<WYJA1'7$RE0K'@\9E#P8HO67\ (LS9,IW6U
PB.RSC9.RS#Z-E!W*+MZ4@\)<=AHH[N(^M]7/HAG^TGU .C'S&.VF3BR8@H-F;YEY
P;I?T:_*5/FG4^WRC+AY"@BGQT7+D1 &1D.VT%95BU%P>QW]+L)Y+YMEF/-9U.7.G
P X*N'G$#:OP.D,2<:K9:F&*EO,15 IU2BO53=LM7>?;173<.7L:T&;IJCJ*VO,S\
P[4U5S[QAP!3SD+ -*2?_%U)B,ML#&W!@M_"$J15HJKDI-C04[.[WUZ()(* =%T.M
P=1ZM"]/M/6_NF!RTC?N9W)Y5>K$"9W- _<3+,2D)1U2'[&+KF97*M.GL?AYTJ%%[
P_(7[S^YECL*O%G+^J^A3667 Q\A9E+8;6,YREX9\"QZT"P!=I:^^"V4% RDQZ6AD
P<8R/-M&H[!$8<,SEE^EE6-&BRFZ1S#![IW<U<NM(\$]U#L[YIMRV6MW=7$@!CG]4
PLH-Y[7B6?9$07C'8,#;/5$7YIBO6.V/LT1F9N,\VG-/-.YXX+E_!AW1_?/'AZC1E
P9BI!.)R]A,%U-Q+UW*O4>8"0U.J&+]/FYPDH&UR @[_W3B.);,!/TQIGTZ%6B=Y[
P2D>[Y>@7'%4))#!#[AO@&.GZ0EJTO[.N[_=*5-EN^3V2T82FMA*XB+H%=4D'7[\_
P^T7AM1P:9%B:?M$?2[Q<]\O'#P)EQ5&8EOQ5*UF9^"]DQQT:E93B.67C!<U]4M+V
PM;J'/R%67(=DT\]9UH9>9 !YLP.$ZK)SC(R3R7+$S6%X:BE)?>TOC-I41D%A(C?\
P]\W-Q;X<K,3O*ZE03)2Q,%]&O,WIOALR<L4CU$[ .Q(MCO5VX)7!0HZSZI/J"9%K
P7"A,UUS*)TT9A0^X+L8]0B2J&REM3GJU '(S:*^Z=U\V@)[I^H.= !!B*"E_?24F
PK&-[#I@\UH0$O?2^O>B2,_4&6J E9P(JYB)SEJ]UM!-\+>=G3O)ZPNJ)+H@N7[2[
P3J3SKC73 >K,3-%,\!IZ,BS5%DF,W0\,EG8L@SQFR1*KAXR7W;)!M.9\RI=4CA11
P:2SFI,T>&"X9#"#MMG49* 3V$FXM&;9B#CVB/Y$T431&%P(<)]!'N9V<!<R_<S@/
P7-7:K+K67XZB!VXEQ_(PWBYX&7VBI]%C" >987QF/:S!=9N;2OZM?\FV,D/ (0TE
P[+'=-]*_,2A*(>0W4-[XTX SJ9,42[%^Z-T>([7#% $015^3^F/V)Z@;UQ-!$':V
P"/0G5HV>NQ*@L;O9S!?"\WZN&+'ZH&>F8IV_\5N^I0-9CHR*Q>:?6W[OFN9<H4OY
P4$H$1.E(G;Z^W"Y:XZP.[^5N=E#^L]X+OU3<_BIU2OI\JWE6@IL?PL O?7+73<)'
P72YX"^?.[]KH?4YR_+#3T(:6OLL,K)393^?^Q\.T<?;7>5W%^T3S4SGU^[R108D)
PV\;@J;@UZ?7'2)!H^V.1+%2H"KC8FQJ4G.&QA)0 UDG56+(7<[**;;(OL"EXY8\L
P.2:O3-M9Q7]17J$FR)OB-Z5B7&2!"\Y]?%EUE>E<FA?W@1.=22VLC@AZXCBJ@%2X
PG"]D/I"W3(R1IWH(<%Y*Z ^IT>USLK4N*X0)*34;.7.0\_=MV_!L]3W$9?PKTY3'
P/24)C;3S&T^Y>\FWX+GP@]ZQ3AD  !_YCW*@7P)B4$8@1/_6NN"TP+F*KXVQ0L'X
PMBZZ%05Q;MQCSM\:_4EJW2@B\.U8?9RRN<21K<B;,@$Q]S!'PY05@SPZ1QQ:A;EP
P)A,S;(S':M,?_WF?U<&HY.<U(#LP.QHLQV933I.P"UE@,W6"*<_*7]JL\QM)RU4G
PY1S(CKF;1I_<3$U%KAD*),1>"U:$(L"T2U<':3_WW R9$^Y;OE4R(0W4X&Z"$5Q9
P?_!7')GIDFBGJ-KEL!<5_FKG1K*^1AU/$S!@O5H33[$WW3AO**(H\]4,:7^&$/M9
P/S/XUXW'0GETLJDPUS.X.#WJ-H8<D9QESFZB1[?"3HN25S*;Q52Y+I2TX6#T4 [C
P\ZIGTRUEWV:7+A:S!5P<EZF*QN6"!ER]"N.3L5G&>8S8QWRV"U*\$*HOP&+[V8VI
PM1!1O6N(P0*&'L6F T8&I]";^-N7)+0G\ [5% 2S5$*71T>?;TOO$P*&9Y93X@@Q
P^^9?2:@V'LJG)J=NQ>S_P@#7Z'4AXX]_CD>DS\FX-A]TWUG+S@%S_<W#P;=W&C-/
P%?/#3DEO.7-7UDJV;?D[!!0331BO0<J' X:>"^P$:$(7SR71L9$!O")^#O?R 5GD
PJ%)%%C,A,%]AKN,G*Y:3SHS!5#P;@=& :$4GRE7>!^"5RCQ-0L9+PY?7J^D6W>44
P.V#AJ,WM;C"<'-VO0X]O:01Q\NEQ^WEO]B7DCE*7]N@4NFBD3]-"1W^.JHH\6#M1
PGR[2G,"A)&O*N4J#W>%<VS:T##].M60=+BE#+W#Q'(M,=)=S2TTW"NXGA2+R$J(B
PP8$@WBGC0R=BS!4$'+!%$\)OV_E\."VL*O:_I"G9CN!01HOHC2%)Y"L3M9HVR\:F
PJTY1VM_I&>>Q&&BUP'^DY-,B6 "13MWW=1,6#H27Z;6N#(J/TS1Y0B"?F-Y1XDU=
PBC2\N\'EKJJ)Z:/KMEMA#@MYJJ/FNAE,U(V73[#%D\E3+)P9,)Z%:9%?##X%;\"*
P'5Z=9BOT"9%N<Y!YEARFB&&U5#[-;3A(!W[E/5])U$%(C2F*V$PO4:._/[UC6-6J
P"A1J5434O,I6 -@S=42QPRHW;\)<[DX>-A4D&!R$_<1H)=JD!0[^TL A#Q^4@*/-
P>#;FJT9G\@S:@)!KB/IV238>_/)I5VH]N;BZG=T7E&U2^9(=ML1=_O30/A!;G]UE
PQZX/:I[ 9>$SY.AEL,DKX$ $A;^AU>R> ^0P) U/V<T!@1TU$@:T^M6L*8QRPV_:
P"P RN?DAN/ZNN?,![:[2N!V^D6NQM,=;H:#4*;SVZ80A<].AYA*"_Y4!)V7:EZR?
PK4'\>B7P5"Y&91(5#\/0SXQ+#8D/G6\/]G.+' \+;.TJ1S:,A]A,/]HDBU6OU$F(
P5%VO,!6VV%B--K$9ALZ0,NW\[VC3("[#C94LZ0" N#[D=?O$X]=U_BJ*?7@77OSW
PW<XF4/W)-TS+?/,]G_Q%W,J\/H,N+QDQ(QQ,K9"O7EV_G]SUXTV_FPP<R:1%Z<N[
PJU0+_'U+H<L9+ PH7Z 0"8V@,9,BJ7LE<:7./T)?[A$^Z#:TG8(T+ZAY>RPMLA(F
PJ:.*'Y3+AWN6+.,!/FT!39-I$T:O2]1!@2DBPQ?%UR)(<"=1.E0 (DE0BF@)PPA:
PPD0?&GI5UX"ERY%B_6G$:>4I&F$U6TVF:P.QOMR'^;-#D*COM@:>3_+"QI6A9IG_
P1XXN4L[#6O;-#N8$0,K5>YOBQRS[& .K'BK#T[(8]X=ESSB)IZ4H#^[YJME'?[5X
PDD^KKG&V#G,+G-%D$U5\QHXVO"<#DJ:D7 N1??\31)!< MWH0?NM)]V[40+-C_VO
P-N+W? C<?P>?8M!1A&>8LL^CRC08X6GU/+.0&AZ#DA9 SANX[DP0ZYU44]W29=.[
PKKVL ')V7&8*O6X1 P@)F1I/F#" (&G1%D\.<!23@''EU;5O[]4(*GI/EF3M+20#
PVS7@]M-A_>LR_&TNU-S&SB/03$W!"9@B"Z*3LXFWY@O*/TD%5:V&@B8W99#K59(7
P2P3XNU7>#P@W,<V M]@8$-_?/_)6H@5/\ 5WPZ6I%37YY3/I(YUBOD>LV!<""0$;
PW1$_7/#NW7.9,UD^B8^PM(8^\B]3V8.BKM;4RD;DMB&^YM3$R-[2G'5^R\ZPV"(Y
PYXZYR9\?%$H'3.R0]Y$,#[Z<G01^^K]D/.;@&);(0JS1G_FCSX$-(^*OZ3Z,9[_Z
P4 K@9S_ ^262-#)IGY=0^CNJ1QJ ."T_*)0@+_KO(VU@(IF-.*%>:BAB8'?;=0<T
P^)NB=H!9PI'H=;P$7\?J))V8%2WM^#X=/K>NSC'V1\%019]DN_84AP892= 4I94%
PTBN@M(8'*3(R6 B.^!'J= $Y,U]5HL!<V[%([/>IG!!I0U3;D(A\_Z@\?I6R4^^%
PDCTKUE?53\XWRAMU$H#/;#IP"%62U_ 2VZ^@]TJ ^ I_EX2]KAM;,]7;:QF(5L0U
P=#6%8W'L@!P2+P4OB#N@0<]GWG.XHJ*/9B_RA@D_9F&\O-Y?(*IV0VHJ]66F]TNA
PX,?>_>-OOG>/R"A64(6B(F@._\TDI.0#;":@:]%9U7JT7_<NS"'^YU#8B3S,48/-
PD\9TVW&DBA RG89K[Y/3"7#RK*?QQ,"K"/^&H2%#D#M1 7]$TL?-3]9F)VNTA'.N
P2'#Y6)HU%_!8J%I5V^H:V]-]B.EOIH@9>!@&87Q[$@2$ACLT'4+EZ0M("IK(X%)E
P*?A)V$,7#A'H,C&VLN ^/:6L6DCRC3M"5'I9ZMLV]"8%]V:L/T'T;CTMWGCBVU$T
P%ZR<__9KGA!$\)CQFZ2I 9S<EQG<QGE@B(MP%>B=-"K8V!-<$8"$^]O"'2,X-P8K
P1.7];ZKS8>_DW&"$$HF/UO(@9@\KKF(H,SVX;MMB$97Y!DZG<,Z4DO!IU0MO)M8S
PPN^U3#W^"S68[B2T9$VB_/' LU;O\*0W.6)B ZF,M5F@G2$6[KJRMTP%8TU?8,C%
PE,;4)[!",#Q(UW<.[^20[08Y^=TLH"HE@NT;2L>/7DHU$\[@2G=1 >P:-/+:T7^W
PC<_%LHI>)>HMYTZ'*W4O'=R!CX5G-+')*]MN2/CCCUV,<I$_-.?VZBAN;=,J2ORD
P IAV\VCNLTX!*B+W)GZTFS^UE,0@^HR'FM[A$,(%I>()*-=[X 4>N-]#DVN3,<>F
P4YZM%N+*'G^"&[M[0=^.A2H,PT9TNU_(Q!;DW#-TBPA34NTJT3\UV85EN:9$>1K 
P9PNZ:!K9D$B]B[XG1>0HHLG%3YAR_M$JU=E\_ A]?4>L>Z2[GK%;*(9M 8\XSTT3
P=-$J6TA4_@X+ DT[INVE+21SWI*>&77YXJ+'Y'<QV8)RGFZ8/EGYU3J>:.7#FVMB
PI;*7EIO4G_8DS,_76Y1 1TZOU+%O.'TUK)2/"%@,LL)XN>66H0S2*XKD"4Z5^12>
P=/,_)/>H4E&2_"2^8M.)?Z45 -XP1B=?Y4C'Q[-/+RIQ#_/QIW/CL/QTP*4'E/G=
POJ H(>Y$^2/3#)H0_V,B+=P:&-4">QX-TTTK!9E6:GMP0I,+DJ(_]-7(5C\Q?QMA
P,E0+("8[)(@*5.;<*G)Q>61_Y PM%ER\T@*B"X&HTZD=U<.9Z;1Y"5AWB0$&L&_H
P^*,(IAL24S3E*5N6T?4I\X\C#F^J&,T8C;ZY:[BN$WEI>S;XN(I:]?+UXI_M63D,
PE#>F)F[78!MS'Y2VP<U@$!\!+6ILH]1[86"AA?ZWE'KJ)W4@8LJ0ZA1SK+P]+%1:
PO$:9E'Q?)R"<!,?L3IM*MQ5(9(-?JC9F'+A@W[_)U?>H%&)F$Q%41*+\G8QNR6#J
P0=Q LB=&Z/!X1HO9[6 F_SN3NP"Y6@9CS\T?&!4$Z4 !Y9!(DXK;BM$MP8:.UASA
PF6#/(+'#*[P9!Z<WH*WF//ZI<-0MJ_*+K:QM85&@_85XM#$B V,XO4(EC;-#KXV8
PFP[X8P+1EP:BD!G3E+AJ#VV?N^<> [AF^X%ZPPR*\L*5AQA%V_W<;SZ:#(#IW\7C
PL".68\4'DNJSJ7*:LIW\.Z\7[A3L32^Z;_S-4D2O=%SNML_9R!]S&\JUMJ5/_N.T
P5+97)!<ALS/8+T9?G[.00J&GOF>CCQPA^?6ER-4W;E<76@ ^R;G[.O1#39YFH[K'
P/)=]TS<8_]9#NJU<B:(;*I_'TOE7>T0-P/YQO$LN'/M#0\F>72>0Y.S=E]G&PNF6
PX4U];9/GMZ!E+=F7G\'-SI G5#8_<5W0QJDS4!&$B-PTY>B%+N%$#QD]_5WEO#EW
PW_Y%XG))PX7;3[HF,A(?G6N0<&Z.>5]$S"I0D%?N.V,;Z9T^Q04*QBT.<2"!2-<'
P@P]YS-6CN,VAI87.^28"FXZ G#Z1IW^:$ +1[:M-NRYYKB%DESZ\@N.]P1N,#&H!
P1,**]8MD;#<6!!^V>X)DXI]#Q-3K:MY4".='R)>KGK[/[??F+?LOELM*R29?5?=O
P<M&"XG9'?: VOK9<8^^FK?"MK"!#D!41L# *8'BAEEIC<HEDIW@S,*Y"$)#')4]A
P7&)]3HP3(R?M 4X$#1$6EBK?QL)5^H  H:34)WW@\%;Y]B&@G8#9](+!!5U!&7W*
PU%<9KH?=J\8"0\#9Y1ZQ'AE+/B+B&D'R/&8[QX1>LPQ*-=3>'53\<[R&_Y(Z7GGA
P'[/B7IFI"Y+^;#">9XJA$\EZ%F!16:I9'V^/Q3#9&%'6[[V,=&3."?OQ* :ID_<-
PZMH]KS)>,P1[[_U38I<[E3;MJDG1[9< !8(/FP)L0LT"3MV 2ZP=XXSY$>Q>T30(
P(-I9B9S&PUZ7MX]X"M]#.+ARJ%3F6"#EWB](PM9.7V<!#4[<GKA2)+A)ZB8!+Y"J
PTK6WZPZL5M2N]X]5 8ILMH[*XWWTY:K95-A]O%O^"O+/A%G\\R'FFE3?&\)^T6KH
PM2%HF=% +Q*6,R]F;$#P,N(JJQ^Y1_M$[FI88L'FG:1MSI()X:V;=3_K%(>8X:%0
P.^IYJ,.V1V1ZKL'N_V8^\-"H'3S22K.6*/M!%W,->A5# 2.F6789=.(!FF%O/QVM
P8]GAG!8NH9??0&X$>55'%S@:VG*C4O+&M,/O>X;EH_B"O1&N4>, [EAKV:QQ<PL;
P[9-=2;OVW P0!F(.*PD.B4RNHOD+9PAE+5J?C'HEFKKR*M%VB=5J?A\QOFG70WL3
PCW<:_S643)#M1%7Y=A^ ?\G=N?@83Y,&7W2QD*6D_<TT%2F*+:W?4[Q'FC:Q@%I1
P[MM>>^[+>,AO!J?JN\*55M.[WX6CD_#O,#<:%$(=:;Q !_62]%-!X.V\KJO=RQ!C
P S)/$Z;N*;98B?W&M%7$0_"A$SR*2!T]L+&7'=!);R53K5=4)A>.,9#Y&U[M"+]?
P HIB"<D?2M2/GR3PM!YX]=.[9.?F\B;*V&FO>6"\+"@FEG UNV=PO.Q(%$5***L 
P\:HS<'TEU<8/*V'  @OI!Y Q6#NC!2/2M-;=6CA5P$[:UT<!OAVM%4W0_R6RZ4+1
PY#C*EF2'E6K;+1%H1\CXK'K:*01  >8&W?Z9UIUAZW9@'*%M\N*Q7%49/5<4^XSA
PLMN1U@Q>^UN;<U#IXF/(-5<P$#T"*>];,.=$BN)=_X.-0%7;?#@R>8[AZ!=?80R%
P(L7BOA=WL]LE3BVQ"8N!(N*!Z*$0KWZK)1;]OJY1_VCYL+5B;1)8P@4^TOQ";Z5A
P7%_K4#H!YCU,&#C?$+B]]XO;90GD<TX4N^?8"DZ30>A5BJ_=K0..DKR<&IVI59HO
P,_H./I\NQJIJ*;U1+@HK*1N@8R#AJIX:L84^.)/0:8YWXV^*_)&W/4+6U<,SN3&2
P$P2R'C* 7=*@#".3DR5&; %%NK7T_FCCX6MHU6'PJ9RTRP5O^)(KM,A'^HY:.NQ'
PO"UX)2TN!58B=?C]XA'6JWQ4ZDB>&W_<6G$[+6QZ[L4YW: 8VK6PGS3.-G-);NJ@
PDV9:.GOI$V,FGH54+7)RK7YIMNQG,;YH%C^X46D)U6:+N9@-RX9YF"D@IC?W+Z32
P4B $CQBB+;$&- I(MQ&A7JK8CCZK'0QN;S_DCO>S,P:9]^'7@DEI&'@Q+2')H>*T
PE;41B7?V<&I 9PJ"(CC(3N)DL:3UQ8W@BWF,%Y'534MY _?V3- (W/MH-?=,"?Y2
P]&*?'M\]QVFCW9F^*"S=)J43HU6YG*O'[3M.(:Q/FY"DP .;D%!ZP 8.CC+GZ7R,
P/7.G3V8M+7.F9$L]8.K#-<\18B(LU<P0AQ':ZS?N[+X'^$Y0V0.E)"GBH)219TZ0
PN#75M S*$T3![!5)+<(!1'-*W2:Q/''L^)HFJ6A0^/G.3\L:>E#9:]KJ^/Q6^!1;
P5T!@H9Y\XRGIJ.T 3LV?MEUTR&#JF7P=[2GF<]1Z J"Q(;U]6QJ@)R'&V63@!)6K
P@9A#0<;\#W$W-,VSF:0YD!HO:P3W-)_$MXA@^!8'KKO'EH4];R$&#+8'9G*D7<],
PVR[_WC[2$QQ#@^F;PL8VCQG 9Y(;2>6E'63AVY/ Q'@87$O#22%7OX'2!:(;_T>C
PX'O<S!)(N,NW)[\[KXR:"+4>)O"G,X_M+RM$P5_U3UZ!V'BU/E8:\CIAM_KU 7]Q
P :11+N(.'\W!2'Q'H1\Y*>&3$G_0\M*H("_2Y840),SE];+\AH"0K9._?J#'U#JV
PWW>$_*A2(QH)KW)1J!_E ]?3Z1],M0S)PF\W[J\QN1O;<$G^1C??VZ@3O4PC"A@_
PY2H= (IA>O!SH8&NI@<@B>0P/A=/Z@*]/;&4L-X3L#55>0"BA_197S*GMW'DU]FE
P]8<AKOJ^K"SKT+FMC=&FB"5P\F=[AH+*E-H)L^F:"*9ER?'!,/7E=G,!*@6%44G3
PXJGC/_V9&,'D7&O/=<^[DPQ>A'JBT7G9SRI2'T;VR.!V:7X^$6][E*+M)2$^);4?
PD)'X65BP RNZ)DW/15SA2@S@U$WY51FF4Z,N>A3S/O)Q^2K[5G\D%WC(5<L-(;'-
P.+^9'_(J>'T'96J_S"6AZ$0I@2,(20P^01W?1!^?\-_Z-8ZQ'- K"K\%4U+NT/M8
P]OAB@EYC]+\[.2>D,F1;,U)%R2"&8G=*['ZEE-R#N(;4=CZ>J<"P(& _KW'-LY"!
PC;%^_X?OUT-++ OYP(F ?.(D':;$6?1_,/%,=288$$P-$ [C=W5UT_NW4 ?".*VM
P=SD7'MM6OZT>NH!'@-^_\.JN*/%^6"$T$DO%<T.TP[2HJ-J(QLO]IO"'W-\")Z65
P/O_&3Z^"WL<@KIE9N]/9M)M%R5-H#JX*^Z<VC@#TMHR [_9&4MT (/[_\,3><8Z4
PUM=P;'W,H-\U-8*CTMW\;83?07-E^]6HK/399R>_))CA8N'\L%G2M#UMH);,X"?^
PJ(%(5_5SJ\X>)/9;X+C.EX4-JE!LYO[J>[%N-%"S%2H2,VQ9@+ZHE+U%O6:EK'9<
P-_,F>83"BO1;528 J(8OG1T.+(C4+A*YP"]KF,\' CNF&(:][4"'FD3G6\&[9F3 
P:S*WE?TH!WJ9?L 7M$"HVT\S-F/XCV B7UM4Z=V3=OF&SH?OW[^G4=THB)S:]C!-
P!*YS$:CGE(SNV ;'%$W6:0G%P$VU.!2A<1:9#[>E=+"?L*"=9@PMY+Q64G@2BPL6
P.Q8IX[2A?\WM: F8>-NG,EC\/\3=ZW@#)I]-=+%R[[C"M0UQ4]!L[Y#CZ,<<59Y*
P2K<P,M!XQC<O%YK#Z!(:FTH>CR\)U(NNV!H3S( :NBM]+"Z);'7GM"5N>/I7ET/9
PO]V$]DPJ(DE(ZWT$(U4TD*KC[7B\X_-N:&XYD >V?->.3X[?@_-[4V>; V(^\>E4
P+.,8MH>"EPX61SJD>C8/4C_ ,&Z,,]B@F:W)"HW]E$K =(30C\T"S"[^K2$D#*_[
P+\B#&@L2/B&3#]]>:%+Z*$+->\2';#4TR_S*'65>,_\1^PM,LP68^.UHTV,L8)TO
P89L'VMKQ8B+=DJ4?H0C#L&ZY3JT\GM%PW >5QH74[&$3GS+W%8]4$TJ"_G[M D!*
P<MK0O!:'@W'E#D+LRIIG9E5.W:LH6J,80UZAMO*![B[J11VV$$ZO&B;#Z::$86BR
P"?4;94G[WC#E2G;%YOZ+0ES/70[DXJ/M0=R4@PP<>R>'FWBJ8D,]KE*#["TA.,>C
PQ8*@>P>WK(<=@5M0V"].>3+1?WI.21N2L=U4B\M4AY_U$<R08V\3L[0<V$G/%3U]
P9C)/RI$I[G-<5#-AHJ Y0>DDGJ(T7B.(>:EH(N*ALPY9&>N'VJ.MGYZXG0$2H#Q7
PG1O1#'85G\N!4. ?1=#W_,Y'OO\SR.0WI,1O)(#+EE!3Q+%I@#]8JV-8D6G^^+&%
P3"Q%AU:Y/<X<?I!_*T-#(Y  F$J_%TTSWC55V(B;1YF*(QCO:+MX\Z+@*5KS0!,#
PXH^:TMX=U/_SY_GR-FZ8*8R>3CAOP'M&>.AL]UMT][*QOO;Q&IO<R@U":A3;,G9P
P\7KEP%MHZ=/:(%0KUN[-RXGP/AEZCM.R F(@>N_S<W5I0^O2:R"5GI5;V@DB$7@@
PE,);(Y/!&,YS]OUS'5O(/-,/""%QB-A N%Y38PPV-*Y/ S;+B#1<#W)R!ZC>]NP0
P-L,Q'&FW2DRU$!JM&0V;6M$Z$8R>HJ:-%3+VP=GTYS<1,69!0O&Y_(<?^@A-#?UV
POCJHF_GLJ<;G'/Y5[Y7, EY]Z7V&9SV9+>5JB8_]O3KM_O^\3J^)(!M9WF\UGX,"
PA-\TC5.[I:2KF1R\W6:)2%4P6&P,QK*\!>O!'7M^%)<HL[G0XUZ=OSQD50ZY_4]U
P-H9,R)D-OF&F%"S&+LZ7+[2<.!8!Y&!\R$[6K/FGX,B>7;>L)WME$9P#WK2NN9^T
P(B/Q_Q&$VHXRS=Y@\=%01ZA^#*.CGS"DW=&0QY8&(7Q:^W"//'77<0*<N78\'J C
P/H,],TCP+ERTMJ&HZII)7FQ?O\@>LVZ0[&/'=^ 0_R$[,C=R>S/A20:JA@G[HQCU
PGQR[J]&NDFT.">S2):I#/N[; -U!>A[,7$7%TO$C6DDQ_L6=@#=S@SH-I>4BVU;+
P?>O+& /4&O4K:1&Y,OKY:@D%#BG$_4?%L(G%I\Z*O$0Y3C2>56-5N(+D?1#;8AIA
PS1SG)5139YLWA]5^N%=@;#LC^ MEF@?UVV"K#+.5533_=7MP'JI>8,V 4P#Y_/,M
P:UH.>Y.(#R/8#EV V8RAN5"U:R7H!F9A5]I"4Z^$=IB2_-,_U55M$1JKCQ^YH:C)
P*-*6=OFY*765TD;#E_LB+%LVVQUYQELJ#>G" \Y0D_6#I"&_^1=!<07#3E!H1O97
P*W2FR47V2=_KG@(.1VEJ%2*D!Y@CKH9\HP9Z,FD[[CS3BD?W[HKG 73.<(&P4P(J
PPT@0/UAHAD]/TF_NT_"B#+=>8GZ0SH\+? ,_VFVK0>36+:VPVM+L<="7C(JAFZJO
P^);PVVSZN&TN *_\M0G>.+*)7+V.YNW*:.9P<GY))6RAH)V8-QKCCORY3/1(FV.U
P:#J.+LJP UY=D5S:P!*]YC//1M]X&6!0SI8^K4YWNH[J-TP[QYP"9587XVN;DZF+
P529E^N'6Z8EC\59(!?,?2ST^]+A9LG6=+^RF#O3UV660'<^3ZXD%G<_X+SK=98?P
P'7'@*!<%QPI5B.L&GQ!K#S _ K <*H<@$1B1"+J PT0PPQ+XU-'MSW&WM/=3F(QB
P0F(,)0&JWB(F,(EJ-W&GB6@$6+2\,*TGC-Z@B-WU)$%S5NP:'E=O9(BV=8*M+6\O
P*=UMEJXP-?>(?*87>ZP\A=+5O/#;90BPFTX&5'.A4M"!TYKZ0PUV^-VU4ZY"',L_
PF76J@7'M2D*/D,UD'*!U 5$Z!FNR%=%L3XPIKTD64A.[MA@(SG4@)]C\\Z4CAVY[
P$HSLO@'-Z\T$FWA4I2M%59OF[0^Q!"[+X%CUV<J=+]XVEG?U!RD?PU[+R(##>R=2
P.\]52MGB"2B?"[N.I D>A<P!T#+&S"3##A\U1D5@MW,>M&WH<R8!+J:]/>?N.P]?
P<::%7<K@A'RGI#0P9LO)94SP-Y'"*5U2(85.&HH*!F/A(;ZF3N@4WO"[8$F!!9@N
P'":XN46"24F_K+6;D9S?P*X!M:D%!ZX*0=B;DW0WONM@ $8-((QAP^SP1>SF@9L 
P-#2^?;]5LT3%\VX,W.QMU)GVP3X>*#Q;M!("7.JTEK@%X]P1"PQS?7L2ZO^MC]"Y
PL%.A+:*$(F/^XU\:;ZI/Y 4U\;B\R819]&+\Z;=VK2\@G/-,05Z]E7"=,J0OQ!I3
P>&\YJR0".Z#/$;- LAUH$JZ6_GGUY$GMBC.1 N-M3(*ZR/U:<> I:[\38V%1BNVF
P*GI)"7K3+@.V]1\><XP/![9B41_;<B@V8#K+@T>FR2ASH82!-MY#9^,><=^HQEP&
P_1JS)3T4_$+\]$QX2B*@Z*T4K*G8AJC9!NJC*8.2PB^O6 %X1+CS5MU)O4FQ4\:;
PX^-G"/-B''9VY1=4UQ:SK[>->UCDTVT3ZAO<_77%SUC,AQZ8F#U^3O7M'PQ=2$@K
P+UX9VA+8.AT^D;F';,:@D&U.1W:&T&!(Y*'CJ1LEWV4]#^MO"O.XH;9G9CD$TP&M
P5Y0>^1#Z2>G<,.K;8^_>,<>!=M))O2 &AHB$'"*05T)@:^VZ99D"&]9B$@3R82#N
P,3[AA%+Q8I<BGH6AZ]F@$7YO<T46O>VJ!ZK,2M=VTBGG<0>C2GB0X!Z7+8,[U9.=
P(60%:EEH$'5/U1-#]1(EM&1QOG<5'L,UXEES?_<PD3#V'L.C(GO@4A1P"(LKR0#K
P:SQWJ59#"[Z!0AA. XAS6R7=M=SP2B"M!$ZLR_)[>BW:D/@>TG?5,8)I:VO-TC!R
PB?YB;)',:SKWFBDHS&YJQ0D8^?S]IF4J'23U>\D0S97-T^+&!%3;VE-D$#F0I<*I
PNXM0&O \&J"^&00BU:%).2=!U&V[*4-\-/R#HS&_(L3RZ+KXGFLRL^E0!'3E1$'H
PY&9WRQX"+_:U3H#0F*_A%Q/ 1%7.6_J94<\H$.8P /\F\)7 _:>_WU1_62@5<2F%
P,E]Y:X79CVO]VH++LGDWRSJL_W@AFQE?*4<Y168X0ETX_%!2O\%;),W&)(MER,F\
P,Z /52_%J+XB%MN_L>]U7CC)FG L9S/)ARF+P)CEU_"=]1GNIL#4H!1=<HU3?!03
P5.&1&+&><C/P1TSLR%0KT17<['1XBTVCZ]5H60YT/*!3H3'UQ*#A=><0,:_\!'7N
PL7C01"#JGV.S<S*=.WVD,()H25B8)\['^RE#[&*4CS%9GZOO*^L62/@JJ##@?7>P
PO?AT<YV/&R *);T7:B5?Y1R)\1?K$,&G'.X0HS_D,:\6LC_R]78KNE:3TP<Y0X5=
P+4RD>L*BOT%63E3A>B)YQ\G\$%;"W>7L#S?ELKR]FA0@Y'2_WRC8"YNM"L 9FB)>
P($Y^3P#$]&(N[(BH']Z2_1NO3AQYBT+N<MV0ZXD=/YET@L0QZG#16+K?P8H8<H;U
P+DRR1#L*2/2#&-6+6>/K0HT4B=&>!'-6U7M<;=P")ZS@_%#BCG%GSQ#MNNLAVL,)
P?=B(W<$JRQ'_,Z'<I\>VAB0XN\UD5]L20!Y=I,YO=D[K[NJ Q?0*JUSQ2,)+2!H@
P;YY=JO7M'UTKFZ(G@<7VMM^?HL$N7=[SSU"!/3F/:+V<Q]'H4V$E&RJI.=4C(_XV
PCQ;)3H6L_%]S556LF%^UPV?<C.XX3C"_5'UH@%ZS:HWUR!BUI*HQ.XCY>CCC:&=D
P&_*^M2Z9*:7]?2<K>4N=.XDHJPD_PZ<\=5>%@.;.<YY._:+16K7<)Q*&S+NTWD)4
P@6VR_/T>#86=XMA-\N'._);"V!(U^QX*M!\Y)?83A1\RJ7>XR;$YEO>G5X8X)>7U
P="W0HL<@"$]:Y_3JCX_(#MJLSYO-@+_;:VP??U1,3@X@2/_H[/]<[;:>0%4$PB\$
PNRGHUQ]MN4,%TUWE8U'S36E^0$@NP-"<U/X05++LC32\0>2FA7%TH=7^@H/00W62
PVAIM+)J\M*>LM^N#P#4L*%N"$/6X.VWN.;&6+ELW)=T$OOO"=G*,\8J:ZVL/@=@P
PY&;6FF ;!X8=,DE4 _9D&J!Q-E+)*B#J*//*LT;$S ),CI)_MY3P;(1=RNY I[?*
P$%14+@'?T9A\P;PUT8A0'JE)Q;86?O&:,RA^62QX$9T$)()C'-ETUIIO_:WMWVVY
PB+=9=DI_1E5?@'EE*1@E_]M?LF@UFR7%+1;!L(GG(25A8>,I,AS?<SONK_C#L[:(
P%<WOTL1;0L%,Y#MOL5O:TV9B/&HU)W?'JG9'0FCZ(\:/L\4U\8#;*2I)4W.7UX>_
P39/?74L6P\!FFYQ.F2T0@W[RC2+=!?.Z<.WZ*!D22BE&)XMU3/6+#D5_4$D-+A6"
P:1/_$#_>IIHQA#Q)9^(Q*,K3 P!!Y&::/'AXK*K.0M[Y'2]O#'N%PMX7 NXXXS .
P,XZ^8"7PDG%_B#M3HT?9XY>J+WYZID6GBG1CQJ-P7)F?SF>O/:;( _NXAAXJ28V[
P^TY\&(.,*#C0C!_RM8D(<(#P,R&%G?8(+MF*2EH<=Z>["Q%@0Y6WK]YK"_WNSA>U
P]Q+]!(_%PK:6$^$HL'_U&' %96%VE67+%B@B:V_"QOLE.BIP)PWQ;[S=IZ=D_M!3
P=OAIFQZ/*FKA8B^:/&2*]%P$S\G3A-V;\;UXM%%].M\>O5]HFQL+*I*&C8S9R3-Y
PT=1J]%R8?!_DL?%$]=<D_(Y*#7B\IJX_',KQ%Y6YRV]C0.SB0>Q8^_N"5[%KT</3
P8N"V7>*ZJY9XY ,R?,"5^G-3L9:+_XR;.%DZSWA D(0 2!$+\G+^T>.XIN[O$GP7
PF/:2-6!A!H_<[7 X'N^3+/E ,9%Z&:[X4D+L2QO-3!V'1;/A5L<V0[RT)RO\">]X
P<S6S=O0+!=,A=E7KM?KT%MV_@CX4XWGLSZHJKN- &DD(;>U;97! PN$,A#!5?B%T
P!Z]E.T;[>WE:&S+FH+P114W,:#U<7LP.1^E1O+8^J[;@:ND1AB<UBP 9*+LWIY U
PVVJ9Y=*?Z(_'GI+,Z4@+\7Q4"-DX+V '%OC/+2MJCCZ5R'YS7(0("9=,X9U^K"9L
P,25FNMF1/_)HKM2D!#*_G+*T[AI+/ ,UXJI[*)_B*;  W!FIP"/\\&6A<(JA53QQ
P-,)->A?\\ML6Y'F94+>?1N\X2")_P[/),D'V#H'-\69XI&D-Q&[WH(9+H=5*&HUI
PH&$"V-8[L_RG:F5*04*%7PAMS=Y9"$$>(+];\LRCKZM03,R?@2/"L< ?,&2SU[B-
POY,T+P;/T27=<@X#];OS*>N5 ^+P6( X(MT(DQ\I%HE1^D,V EO?-1(EPGG >.&K
P.?"*W#;1(U/I8[LB8IWQB,OADSS0-!?Q'_/L1AK_O\RYUQ:NA49MLXACGQGOGK<5
P>[A3W08&"G9_O:XEE:J$DXV'[IU\4/57>H5N&D+?T0&FG%.?(%D#94O)S+BYQY \
P(VIG!3/%_1#C&7T("_0MQ74O5"-#COCYLV/&EQ\A+&L^7F$N+97O4+&Y3?JG;(8B
P5INO;3CZ/;BJ W,[92$$A'5^\47'";<*^P";@0X@*6E"/^L<5Q1,PS8]7T?'H' *
P->?*FGDE<N=?J6D%\Y0!8>8"WD[)XW&R_#I'S+ARJD6AAQX1.34 *8:^-P2,FF.=
P\A?3BJXQ8TE=OD4I]F7WH"294<I(9Z!GYV* SR!$DM0MH")(?RML6NUB[('8!YIR
P;L-MKG>0[."Q5R*B&7T$-RXVCP0KK)<*VWPXNPHN\HDW-,UJQAA$@KIF7\->[_;Q
PF+R=OUMI.6A#UWRU=6#DKS.^^K=$ 3R_%3, 0! F@6RPLG"T8C+GH/>[Q9H]*1.S
PB"1L_-HPYO=,+0:BN:XTYB/9N6,@#(RVBL+I=D1JL@!$O%"WD J7PSQZH/4N$TTJ
P_1PUHFQQ);FA-6LT,R3!P'OL7*N\!C4TO_EB% +.U]Y ]'-D=]PWT&9>)N_,T>5D
P:Z2+C;5<2JE<QUP)6&.\>(T-K%,QC:71_)0+C)-3469CH +#"-I%Z*>'>+-FR0DA
P]*;&J+&K:')07L1)J"!HP<!42H.?EF]DG_U7<<68,D/X]F=]++T-K%#]$BZ+CH%T
P8*>!!:1O6AX-B>!0'((HAKZV>VO?]ZB^C_*QK:5J^M *(\YB2OF-JW@J0:P2QGK6
PF.OY<M#:F(.=WL$_'#@B<S"Y$NWKOJ%$;%:13)+BJ0+G14% !VZ2^P)-K6%;[^JT
P*XW?%/;; U:6ND5 N=&HQ4\&"^>V2LG^D,*ZGLVD 7BCZO'Q5W+X"-S:*WD 5&36
P',*2J>N[K(I->4]+*RG<BTBNN?H\+('3E9G2@M"2H-PWZ2PSB"K,M&],?_[V/?@V
PY+ONI<(%Y74"<4TA9E+5E.?445Z1>;OO(7/+Z)O+VJ]%XI9,,V8,'+R5_80L1F&?
P.\\AI<!@.=P2&%":!9(OW$-*QR'MGX+MC66E-03C6I>O ^A,B?)>UA$F2@/V[*^#
P*EN^X%N!$OGB/S]+-,:S%MP$3!81,N% "6%,K$'1<8(BSZ2OJ7/ZY=4;\?M-E'-/
PF!WX9@#A'^B/G33/7B:8$ *TD@*'KSLE,?*:AG&6&]?;++(YE(=+=#VY>IJ?)_KR
PLM<0]1;/H='E:%9]D@K;5\]K/$' E"-4L@BJNE#(WJ(^U2_8H HC>+\--[/:-R^$
P:\W@72$L$#O(+JKRCL)A?&F86:[T[.Q934Y\<[M_X5D9EL3-Z,(_M1N5[C5252=N
P9-M;XXV>BG._&]&B.A<HW1"D/.7WM_2XU/Y0*MJOJVY\591>XRF,(ND98GY!)ZFZ
PAG1ZC@.9]L]"2Y,N\&^$@&]1-;=56-O.)^QUOY?\L NA%9H=^^ 9K(1[_0X&/D_F
P_U^4_:X /:Z]NI/[J78J'@RB]<N.$");B40WE/#FV9P4J; 6-656V1P!OZHHAW[=
PK/XT0R3Z?V%6S2?N4R-FPP)^09HT.]0?9XQWS3*:NC3_G0KO;AM]1U.XO/:-'!F2
P7.A&%:4&UNOV;^:PI60MU#WSU$?QFG2?KG(8[U@CS"P'V_4D+ >/$O?'T;Y$?,'H
PD'$F7_"#?4GBJ5;3]/IC4I@!9BA\1,QB=O;+?Q\R'%28S-"UBWB_Y*[)9<AC TB8
PQ8\Y+HDI#8$400(_'X]0XNN%![,<5#NS"H-2-QY_<K2IMPL?UVS5^2CDK]$_HG*F
P,FK -7:>)Q\H<+WK3W%$ZC*XN4W4#RUF#;&.'$Y!AN_%Y^NOT_K[EB4,G)5GH:UO
P?<N9DKD7I/ISVW$D68NK=S39I>6=W-:*/AB"\\ W*KRUK?MS*94Q[,J7SY\PHAD@
P9<M/^$6W-A%*GZS5NXROV':("AM>EK%$AVI _<P3=$Z"-H_8-R;F/",U5PNA74%[
P4?AZ3I1&J/K->#EFY,@F+OF!2ID\'%=/;.^3R+*OB-X0)@,C>5;X%[+^IS]S@D)N
PV->P7@0U7ZLO_EHM"GQ(-!W9VUBW;A2W724!TI7G+YI;ASIYLVE,V:?$],K;"X2T
P)NKTJ"TA2=@8IF*]F(T;@6@<AC"7LYO!9I22/B,S9?\"3MNHGS:^IU#?"$Q0>K?(
PB3T-/NFI"(H-H4"VU",_2 1P'+(**(^29-2"E"0VVP!@P:KW5WX8!1$3YP',JC*I
PC[1:4>>X']:3<P77?<G"8/2.YC*))6W&5>"55-%)8I"O5GRYRM1WJT$"!%29^M:P
P_YM5/NZ^#!5(G@D8P7.DP+;.\OFS1.2?<6:U?5=L@H0H/*^R="G#AV#E^O5FA++*
P+\V=ZW52/E&1E&$ "+.MK79M&/M519E"7LG!S$&=7QZ$8T([G65,-UWLL4K40ZMS
P0B%A%ZBICR$2-Y\6^P-:G.\HXL"03\?<Q-\?WN%)H6.E$,\;JEJ,%MC8PZYIGYGT
PG1#793JM!V*@(KIB_P&W.JUF;4P_2L1:9KP?%)6\AK6O&'7M9/_2IV?[ Y56 G#<
P@LW5ZL0#5ZRO<A'U==P-G;7@ 0G*=*IC:$G/Z1:5'J>66PH?#O=L[6AC^JD>PR^P
PH%=<$20E5NDVQHFD?+8DJ,D VF[+8(P1C1'\^?'0*B_T@>M$=0(C9D^G!#-9P?0/
PK #02\S\F-AI ?UCL/?1*Y =)LKW,5<HBS@6,*XDJ)BF*&P^%;JAL]33N<XXM<"C
P. ,ROF*FIJPB\A:^($ZV^**MO/I(Y);GC.([X[K!3BK&S%0Z\0DZEV/VE:*6Z4/=
PGPUKR$(IUR]GC[G^&O2WI;9S%%6?(#D*RVXPT(C D^<1=M[D=(,-5:2$L$L8A>KU
P/TXKUV_;UFJP&3>?3SULS&IW]"'I" "S8<F9M2 1E187HC0BF#N]1REQ'?NM3(.K
P,H""8"WGO*QY:AAQFG[[K,_=B BHD^&N2AOLR:W;918</29,@"3,K%N'C%?E-#$/
P<WL!V3@=N($'&RO3%"AN<,EM15<LRB$Y,!SPY*4R%(_C9!6R&9"O.1<C01P;%P08
P8P\ZR$::Y8S9&>Z( \; ;SDT9/P_T<B47Z+8&%--\O/L,56]#!WE!5(30-U5CBW,
P< Y)+GO-4O;_$O)04XIGNMX1KU<K<)S';L5B.(CQ1A7.VL<CZL_#XRU:2/76EE08
PC,-]XNL$MI\@M24AMQ#;I:%@1\"B&?,LN55J">F<T9\_-=>NI[!U >=R:TC(N /W
PYI-M+FM5+A7G5*QAJV>'C:S0)G8K6^WA0OP(>2&2(^G7GW3K[33XTSB@ANN+)S#,
PJKP/(_48R+=><'*Z^DDL4_"E*^VTR0X%#7+8),!UYVCSY^:WI^SIOWYLDI!\Q7$%
P!>L)'?*C@CIG&N.4;0$%#A*]=+_WQ/P_8_8N!SU#+*8-!UUMB#\"+?:B?EXQLL,U
P?"5Q!,:FG1T<&VG0TH 8+92[J__SQ!DF&&&3B@30M$0XW"3M8#YSB0(SI21="XL8
P.-61+C3JG+^:7<%LL[_?93QY+G1$D7O%.)\]4#:18GB$%$!;0B* +=-"]Z;1MV_+
P:($8H [F_LNXT%U^5C+;?%A-.^'"2 #>&<%^'_&+6G<7\$!=_T--R04[ZI3F;C:I
PB!<6%'1#@3SWSU=Q=1^57_[)7KO:2,MCPCD<QBB0!NI(-$&H$"GOJ&)YMKQ#X'EY
P+X,5(4BZC[8"_:&+PNG#Z2_-TS"=[4,5@47#:F4: VQQ4282\G9OJ\WS!,XEP,_6
P$Z-QG5*P_5$5./I8;+O9 2$QF/965ZKDCUOFJ(LYXY?Y[_>/@6$Z.O%5SVM5OB'-
P'3WI2Q;N%K&PFPH,Q3.=0"@2I;:3< 6.4, ZCNN:#MX.K.8_#.?LROON2LQO5DM*
PZB&Z!-9".I.XK;D;+"1;DC>0'@ _[YK.B& MI!/2V,M3#,\3;5&R? )Y6YD 3 *B
P;##'B>4.[';R=1-!SQS#<.P.TBSG%AGZ?;[!A*U=81>W C7)$:<2&HFIQJ]<'ZXX
P1&HV;^BZ=F\6MC5L@;V4GQ,G!0G#E?G._@J@[,$-:@+ //<,0^$]8SI/A?-YK$R8
PRM?\6P]95Y^>"A!F8+/C&(=F_E31Q\/T03:1$62^VP_:J*?T@@)!N&TO#NL78_YV
P#?#(5XM4^27_1"J8I!E8 \K[-?M&K&5VQ43R],3\1B\64DVG.;2&&JG' )FY]3N'
PG[ACMP?."3^(:TH\:NCI5'4 T3Y^&B8[CMCTC+KV!K"O(P KZ%,IB(3/];J6YY='
PE% R&HL$EP/LID5DMX:6O_5\6JV0X=N ?.YB6:_]_CX@CX+WY2B3]:/A/\S(?8G+
PWNQ5L^UC!J$GQ@0([8[[0W)\(.STODN""S8DT[>V*QPMRMNMN&^>8H&!70E2)\-2
P*P ?>8SV=LQ1.?E'<^K3LN[/_U$(JE\-=5/0SY.E;1FET!42+&YW/[OQ+2_I%$)O
P$3B+"DMGM]$=.\?J1^[,NR"<@SQ_PJ7Z&;?H Y?UX- \/B0K'':V:X'0\7I=!;9K
P02790LY_OU>GMP.<#1NF7X2>>D.#CX(9T$*HAQD>3<C]E6\GZB9*@H&!AQ,]F3@%
P.0=BP,@AC:HX4(A\WR7'U"MWA5'0:XAGE[RM@@E\S(J;V>B2R+:"LKL-')5ZU4;4
PD+F3-$[T:IOCN)/]Y($)XA\E@267ZC&A<@/^]T(QH[MU2F4C0[1-4V?/L=*9P"90
P.LQJQI9CB$F&8&S(-WA+Y=O)Q@"F E<K91,F?IS*,:C/%H 4K4! X/J3(?%-TLL&
P=609!L80:$>,VB6&'[/?=R/+(JTE_6"5_A2LTVY&1K/R1!JLZ1#)8G,6L@F%5RH=
P"T;3<6,5K7'6N2_5U!IFR!9#5F*'PJPV^2&"'*XNEMIKMMPL%,E#: <Q<4]X)BTY
PZ!P!W(XZ7P9!3,D,HB8B?X8#36GNNE%]"D4[>"(,V#I8_BW*,^,[QG8&W%E6M0]+
PEZ^?.-+YEZ%E[#U#I55O]SFK-TWG1YR%PJ$T1!F_A3^/NHI#QGJU<HP^T 6)*G,7
PV+KO'T;?BT#8!XJEPH]KK'-A?%#]Y5&)3"WF0ZG1<)) Z- \*@*]O*X#DY5M=W08
PJB[+M*1;4$4=K:8%VM;2NS!C 7AC0X3#[D\R^&L$[\ZR1D8E)KUR28MP+O2QJ-_S
P[MF0\TFY! YCD"N7)9$(,,96! ON(UKE?[WUZF\2.&J;( #E/TE1]LG>:!<7+&6V
P%@807%O[H_$N)P^629B%B7Z\R:M/HG#D@8,NFPBMCHY&.5EK66])N/(QQ87UVMNK
PXIB,JRY5?_:05OZ*OV3S@.(/27EZ]D89QN2RH?Z&J4Z.QB.[ KQF[(5!D6F%A3R#
PMG(+W<G:5DZR*0S^G$HL*?6V7G9'_W-KG/JT^#*R@4O;HT+=7*3 8.%3=,O PM+9
P%M>06,)5;V7V<+W8&QO>];]+OH@R^<+M6GJ3 PC*'@PN^V*V[!M1HJ-RVTBD(:+J
P?^VJE @ELM,&S</>NB%IK3-:'N^;$X4_1EQ7Z9L>9R ="YR98@HRX <1Q8LX(.[%
PS\& ;IRRKXA<DEW8*6*(.GE,ZSPXW@==0'WS28-'NSLWQ2'^0-5'LX!'WA4&/U?B
P,E"IF7%I,4"KJR/S["0GAK;%!GOEDQCV%>TX6O9N&>QP/&XS9G82RXT5T5.J2MPF
P^Q]55.[O44P>=UF[0BC$RK^(N29R+D/!GA(Y@V0 ,!($7*;&H^^"]YEHSCO3V&2Q
PBBI9<!*PC%5SKL)'46,'GMY G%<-)-T0WWM8S;0)3'N>4'ZM=D8<,;R)C.2P6ZS&
P6HA#ERY@=J%$2,SLBJ*#.(AN##C'4O7MS.%K[.'VGAL0=E)=TA+M^=)8S0D\BO@\
P4]2R"@Y0%EA5%CNE/<20ZR9AH N'875QI.!_-.1=$B-L/)#,\087N&/2W&:<4&, 
P@1U_?5<(,S*N^,YJ-9.##>FCVUI3;><DT F"]:JU> ;'TDQJ@(3GHN ?@;^5RT5I
PG0B4T!QB$=51<-@EYC"!$G(L^1)^EJM(\SS_Z#M!<B\\,'WUM-^]H$?YFL-2\OD&
PD'9UB+//_,F$XZD_UXL7@F1:='%^$"3*_*Z_=?;H=Q5E"/ ><;?V[P&A_*M!20LD
PL$VO8H3=<.LP_9;($0CL!R<%D+9E$CU)W+YPZH]N+#889JZXW,A4.#:.P [TU<[*
PDKI>S:,% S*?/ S5/K,K)5B6Q6;^*X0Z25[-;$WAX#Z?RO.=*A>Z/@(V"H#' P71
P@VZ3FJ0JI91;ID[;RS0DZ*-51QL*/.'!V'OM=T(*6(3%OKMOC;1QPQT\0+^1Y'20
PNJ%%"Y#C(O/O^<?MTZTQ_5;X;U'5A$]NBP3<MVHMM<E2"*U#9^Y[Y>&IXJ*[>+>@
PS0WIY;A4%"U[C00Y8)7OS-:[DN_%RD6XNM3)G []SKIVXX61J+5O:1==WSI+E\(@
PBCYJ0QP>Q"\[5/B!(K=Y8./&ML^]=&X5>%GVN[MA_(48I:$D<+\-27:P0(4&8+3;
PIZFV"B!'S"BU\ 0KQ .[8MB:1+^)A6+WN0'9G2$[<*#.7P&A^^SAWO)%&0R:VA\=
P#[G[9O$J*8?AA#[1AQF+C'#>N.PZI(PWT55XD+@@;F&\PN;JJJ.AI.Q$+ P>M.!7
PN!EUJNL0BG;-F@5TPST9W)%GM(!@/^V=GR!).D)Y/QZ)>QG(T)%27/(LLYV'2?U9
P_Z9SP0$:[%JB_[CP:AI2?''V6B""@M==MGSZE#8N#9=_"*XKSWH97RD<X@8Y9TY;
P*((^I-)).W:+!'H^ID5A2Y$F*?$Q8K]ED\O6M!O$'J?7=(R&)BA/3>*M>+4&H?(M
P,%P.9WQ36116G$CN+MKN3+A78>"%0Z(PP6!+]."5MU]J7.QXU;6"1'Q%^YT(SSX+
P#'7*\?474DGO8$Q(:/BM!"=$N.Q2;_^ZUOD44_L#!$5:Z._WJ1Y=N+_J5Y\#ET5>
P,_,(%F*2,'S?IA3-&W7ZTXB>XE$;<S95\9E;M!40WY\],Q"BZ!0G'D38 .2>W2 E
P=^O38TV.I4-6! *"AS=.CDJ"Y!]4"A-C61U#N#+XL),ZI(=!'?_H(>G<\A6D13 <
P*' =A(.*I\0GG>X4A6 /7RA_M?UC4B5M^I20<J7Y(H$#9UY]PNI!K*-6Y>+H</&\
PY%B;<.X<)E+8\CZ=3#DU-:5[: &(0-_%XJEN7]ZGT?5,70<6K"U7D&4*!*@M<](\
P%5?#6,%;[8E7H@<H3U0(7GBG5UQKUP&O3IZ)V:PNRSUE(#E*M2?M$;9HD<LK.F1X
P324 O#A,)KU??]<$D/N*.YA&^]#,/K=?<3I+4GF?<@QG;Z"Z6<K]O2%=6F(5T*C7
P>M\AL8T]45N%!3X!3TG))^&^ OH@%&0:@@P"PW.9XR>/N^:,!W,7*$U\D08^P\=R
PML>]RIDM$HR2%9S?[KD0U;\,[Z_<0-N@>>JNGK%YL(^&@=^#BN,PJ;!VMDR\N:R"
PI"-U#0O>](N @*5[KF?Z]7"%H]CM?(8;6GK;D*.F".RT/"=P:";]1-2^XASMEZ-M
P 4@#D](T4<509 6EBZU<^[&7E?F&QJ"<@X6,NP'7_#3*1EF_PXSZ3WDV=4Q"L=TB
P3%7.E\8*&K,M19_48F]<=0&U"4'PV"@&7L=M47&-!DB7L(QY!_U@K 8USCJ=+2T8
PV(YIP3!;+(<??U7!R:F1EXU.XI8]C.9J=%G4M(S7NPQ4E'0>?:%Y\K"I&P+>BY3I
PH*?Z]Z$@]G"B,@5Z'BJ'42_-^%]87>&KON(GCY36,- VHW^,D-URP<\;+HEUI[%Q
P*$UQGS2D&>/7%?WCJ=@BFT7N'R71CY%U&A!=V*P=>\PP,:3N)=%OYX/2!B2EM79[
PY_=D$S7#I_P/7SX0I1:]]YHU%AO5TX<4B?4D>+?N<8;U/5K8IJ"C.O4N1W@'1K.1
P61<0)B=U!0<B)8O<3J;93J#J:TA2S2S>F)"3% +SS#"Q$F!]D9@=(=>&D^N?>,ZV
P$A5I*;.G:'2VO'FC$TM(7Y\^X(+D& +G,0@S+[/4,801&S=68QN[\>+,=" 0C-U-
PN.KU&P/2S#VRF8(J'N.XJ EDBG?7G>K')U?R3C:$_UJ>G72#EJ,('GDW!,D5H4O,
P^GOQ_$DU,86!)]S)M132B1I>!QG210!QI,8MX@\O%,P4&<"18W2+9WE?$35T<-S.
P@<PD8"IB-$%M-HAZJOWLXV15R^S@]7Q0,;US*MT2340=LMZ_CH6:UQX<;B&U1A]$
P/?Z>S*Y:] Y:M 780AA[T4;ZDC2Z:CIY[Y+ZR\%WL"0RJ)G2']DTP=SG^Q'>_IWM
PQ?PGBTRC@)=V_*^72(]#,^Z+(E"^+>@B/AD#-B/&BF,!]_6U'Y8#7'F=+/8;,&]]
P7K5A^#>BG:#OA572RW*$:0PK</+4SF:H(^N%P#_O&C#$=Q4,(:P\OY?[PZ>J%\M-
P66FU-<5D7]LP7'QE6@967;UTL6YJYEA:" R2W'[M:Z+K0]E6$?ZH#$7">$F/C5)1
PGS^5)<U2^/P48#>HTES4<44&!/9K BN=C?)ND<E0B;R_YHN_1+7&;CI&*<%6Z]1O
P?2KQ<<&[+L'S="RS>#H;Z89<50N%NW&WB^GY[R_J>8+L\X_C: 0YN+[4%MOO;5#=
PV#/$$^?9U"".T]ET".7R)R/R@L7G#%QNZV_<A$!^^#FX+&R%%<%GZJI[NP@;\00,
PHX#V\!2#:X)0;,A]'GZY^& ;_$>D3_RM5*EA-@O]=X:I=!_8\.[>12PIW!-BI1[1
PY[;BUURY;$=&74 OG+'"B@I%EC^GWDG(+3KKRIIO,-].UY6TOIW9NY]=!) J"_;;
PX76KJV#PT>RT3A60K)";A%Q@],^L"731'[P;AZ&S$MOG;$EE^@$??;?1$PL36A  
PK2OO^0J]$M:(;>;IK<>6]*/,O*ARAUB0.&<GE&T#BQ?>#W7$:()E@'Z'X9(MA?WR
P6>IJ&8D2V[G!.^,J<#8]*37)X[CLG3N>)Q SFYE7%IE0AY/M>?=#EZ)4P&'=%#7B
PD<Q:KE )YT]&?U\5N89H?YE\]3[XJ5NH\WGF?1C6:795N*D>)03$)-.&R4-;PK3F
P=1#5)G]MMN&UPMB[_B8BBBA&K<EY8K434B V'5A[)Q"- Z"2_<5Q\-R)?\54@\N>
P&<4.EY]2/ KI3^+?YF)W%)5!YIBM&QFRCV @?J809/\-NCL6I5C^D3\'!=RB/:(4
P;\X\^.#_3[7;P;61).$8/.+')R .-5BMJ1+*\ 7\VU8OO)"CK$TQQ=Z7J(^_A28S
P"-P5HWVIJ.BPXM&%P!4B;6==+[O)EI%T3,QVOMY7=S\O5I;'V!*NZ WKB[[M* RV
P+*.%!@"E:U0BT8"!'&8/EE%75<U#!+&N9($JOQU&Z"P!Z.NI)[L67C!])C!/71L$
PH0D)QN[@6;<F(.[N]K#4G(!<7%/DN3(O_=%/.$1;14+R.T_0PL;V_BT0\"8'@6S_
PW<]WR4PBF4N=G KY=R(_6W =!1!C,$#?8H-Y^3]?JLX(YX.HET4> NQ&C+N;Y3&(
PGX%ZSS%6CBVE3MFP\UFLIJ!0;/)G_^/9--867OT=K@$,;BA#8!TG+5<8-BAQQ[?S
P1=6++-QEX#0M]4 1FK4&"DG,3.\GEOF>:GRMT*KWKN6=C,M=VA[WU'(-)F/;P)%W
P[N" 9W%[C5%*J$EA[,N#M=0#K-769)JMW A4Y8GTM)GX6H^7FJKP4Z@W!RF%Y62O
PL V*2C35SK-#OU"@"JM.:AI*? DX1@E8'G6!P@6/_EJ%UL&3R,^;=:B5URJ,F<5O
P]@%,_#\QO(G<BE%KH"?XHX=W1:[PF#JL^S\@X5HI"5,HV;PUCZ[U=54M8LH?(2<>
P+/$1%_$;YO.]P.8/HZ1R(D)DR=+W<9"3S>O#HOU\V1YW%EXE";?F#W+&:-C WPH9
PD2&930VHP>'D<^GF1DI?6?=<'5??^<[K]39A$-BWN=GC2Y?7!,K1L.MM#A.;U^52
PIK@?:A=3V7@9TJ'1]<@6;,3#+\!]].RU<]@\<D^0%Y:F]NR#US,.-!SZ+$^;IIRB
PU1Z_ON%,,R;I?%(!ZKGUX)9Q_1Z9H9+A_Z-!PMPDT+@_GODB0 CL" MM\;)1NJFG
P'Z$E,MXF@WX?RDZU3TCQXM]CS0'0L[MCVW;; \2GS[8%!01U1VH>&*.K_C=/6%L$
PT@)O"213C<]*J8W=5K9T&I\R'X>OE8*<4C<#FQ6TM',)5,\*X45E!3L8#F14Q =T
P_7%!Z^S>%_!=,WKI03@B:J_Z3"TKTYF34C8#F)J0!-S>IU,S^,U.P*FHX"93;::+
PH1MX0P<>O1N6*^,Q$L4!&*MVP"UVGM/D /%#T5ZFG\CV*8>$O;*2^9&B*\;L[*OA
PL'*+74C\4D*%HVJ6"Q>KHG]N434K+A@-HVIW9X\;[$:;,:=>F]=[]\$( ??:2#N4
PCMZ&6#PZX4$(K:C)\@([(H+SZ8^+*+9^X0>^#BA BE?NX+A47K*PF#C[+",QACCH
PM2#<S2%2TG3NP0+HH?P3JLB_*WP>2\&R50%VEG]3T!]H^69RT:M3K*3H:K,DUG+N
P5KR-8L"5JH#)R'&)XH&\(JK$*]\N-H0P<5:%X-A<D;B@F$E"M532,CF#]P <M56Z
PUW=FTK0N5DO3 '@C1%NW(AH.QAR6Q%59P[K<&W0[5!XD\"B6!:.GF_WZ\U9?2@5_
P6J79335TOY+]$H(D>I';9093++-C[  N)2O.9C"N51L6&5XOH4VGN@IO556ZMKYO
PIXBX!1?,(;VA_9&"O?^K_:=*PQY!':C/&;U#8@Q;$P(2.D_(O &+N !Q8IWO#:1:
PZ'R@2Q_R-(\R/^PF5@@*^Y4+=*?HOL1J?K9U3CU)LKD!6>NE,[X7"FBY^=]T8D^=
P>]"UR:8,0COFTLQ$P#R(H;TM7W.QV&[Q< : 3F"\^'\SQQ?C]-#?1$_B-EGZB^.H
PNL.R))(-.M#/@.J9_>P%.9  0GLSNF0'Y$W _>\>QORH/[>W_GROM93-4=?QS\S"
P>T@P:Q:+%]1/H/<H-3\I*6"BW30<W>X-K;7;,S XEE1A_L-0T6"%K[3.)@]K5D/\
P8@;*:IT+V$!DAX).XK+2& =CFOYVU_:DG2I+I7EX.-"GU"G +$RSP"[B8F+8WP)6
P;Q#'/N98P?,8<M@4#(.7^>X[:.8SBK_$&O)Z@,$X%B,0=-3MBLCBP-'L"30O;T#G
P\IW^64IZ3(EQR(Y()?\1_P@&$(6KHB 2JH%!%44_5I>F&9U=\*3#4U&U8^C4I4W7
P*;5(>D,4.@O[55N-F9#H? V6R0.NH 9&Y^0H78$Z#;A7GGPB:Y[1NZ.V?GNL#-$V
PK-L#:_^EN=@%NAF A(U-?SQGSMXH.N"JA4';\\Z'18)*X== O*IQ+!2ZSPV%,6>7
P7] 66L^>#) >TZLGZ8#M\M/7_5]@>M@ :4XF\[UR=BR;M/PY)@1QD6NRM>;%5N^<
PC<AM$L@Q_@_+#K;,+4^V._F$)^M$XHJ/!:N)'8I;.:[SO>&:86HE"7<0X9%!.G^A
P!F* V4MI-.)UAIR>%+\,/&W9'X14+9$,-F[LW.N#WX52]27<%]88/D.4LE^N6NY/
P#B2JU@AO@)-M$)M^%/%':+#^?Q6YM &QVB!,[D&.]5C@<L2D4#).,3+1)O2B)?>>
P$$JBZ(A+7!3!\@^1>3='F^VE2OFBCO/RAT1>5LQ &?5LRG=A1&DST5B"H#P%]M@0
PA*^&\>==BC[K#)*00VY_<O'_7P).WS=)\ANL&BPT?3#NN4&LIG*AAW>33G%?.O1!
P:8=5+7@W($>;VNDBI).#HA3.)S!RFLY*CUZ>"]DT8H68D\K8/]+I8T,^X6C:^&,"
P,D+S(;\0F<P'%:>+H=REH0VX.OTC[ 4G^0V"]E]9"C:\(8:F8'%L [_K6JR4ARKN
P."/'PQRW^,8OVQRV\]%HL2T9Y^2Z\ )L-#K2O4W@?U"TORA !Z*&3>0"&A,)RH3F
PBWU6 ^>$B_O%?"V$:"$A\>B9L+TY<+L?$3:V'?G:5,\;"O@S(5DE"&64F\>SR\'1
P/@=F=*9/^$B7IZM#QS\AN+'];,X]OMCU]F',G\((,P R$7:)/**\EZE!6$ZT>3SU
P.]@<:T[=EZ2:]RL9S#4+L44.0:WTR"(E/;FZFZY&_7'S)W>]6[8SZA=EOQ6'Z(,I
PS(63)&CK4O>:8N+-<P!OD6DSK=$ZF&)58^9O=[!#!;#\,.(OHT153Y[WT\E)9ERQ
P1]"C)R5QK?)N!9#XVSL*UB6/8(Z3U4*NUB5-(708MBY<F(K&YV_BV=3^[8@;#6\'
P>7WZJ[3UA1.<E@(SJ:[G)O(,)N>"3\S?$L?A?UQZ2O$[Y(=[S"+J*)Y,*8W-:$&$
P]SM7K1$?DK'LMJY]"44572XZCP!:1?A&[S57=U 5A);H6E3^7G=0*E\(3:-K)E-1
PYQY]-'%Y&#0]2-+I#FP4Z9YB83'?7\ZH)%E_"G]%\Z9._&N&0.1MTPH%AI<F5[07
PEQG<XX9O1=&[%ZUA#.6NH<4NCH%GN LA_\'&22=56B(20B"<R!(!5B&;I?04OG("
P3J.V.I.GK'/;IS(F\G.P07(>@*I!Q-1AS94BA(72$8&KR78P7)7"OM)!6Y',[$1H
P5)/<J;C)-JA"83: AB4XI0XISU5)$[N=5[>W/>&R1M_@%H1( W\^*DRL8_76]XJ;
PG",J( ^\/*0E$W*%$8D.L2-(FQ509YN(&RF'*9;ZJSI]JD8S:""+'<;]R@30,4%Q
PBDT6NGW@$#*5Z85A5L/64"/6-Z*0$O(%D_KJKD814"&\H2@QY[_:\;N='IPA(GE?
P5*Z0V$<>[3M4=A2W,Q.T"< U+TQN5O)KCDWINA^8HMBGYJO MM@E-TVV*1JC4/;'
PM@.7Q_4J921I7L\@D/*<S;Q1/\$(>BD3V]C1=F5O?NQO6&:K!+4%>< B.QQ6!801
PA1RP"\H:/=4.UC+#+[<:39CI97:RT+PZ0$%VU&F4WS"L?>EON5_QW1QV35$7,IQ9
PWDFY\@Q3F=: RMVXD5'\O_JV7@3VR=P]IJ]/1#FOJ$Z@^SZ(RX$G_O[:FNL7FVK=
PYX$3-$B1>[R%1NB_M5SG/S)J+.U3,P?.NHWPFK](?K9Y[A[L> H81TTD%KO)$+3@
P7_ 2_4Q7#+6H(Q5XJK<MRM=N53Q+@=S()T_<XFC&G)+(>'O=CG%##2O=TXN4+3@7
P\V6@*-9SM[7^QVAF5[3+.=BDC3D2W@0VDWD;WY8-6[8FDX.K4/[%;I7'Z!89BJB'
P5Z@JHP5[,BK#."RT%:4PY]]TUQ@=#F[7WJQD$#&7';V'&K23C="] W:/) S"O1^>
PENT<8-=P&57]YMA3Q5_@#2)^*\0)SPF-J:H.SED2_!HLH7/@\TZ!^=J4OI5L+'M]
PPO./,9L%4/M+R=IO/,"5SP,Y.K-&WBF/OYRA6EB>)B(R:<(OT7CG!AP:(L0@S5%A
P(+VB[H-M(;WU);,S@=0SBKB$4,,'$PZFK?^DY=]G)1L))4DT*S4F952H8J'VB?@+
P_+/ LIHR&" IAIN\>?8!\V-90L5",C2._37\EVKJ!X,0YK%WJ:VVMD4\%"),G+8^
PUSE'R*,.9P*9(F96V6-,>L9QL=2%*L 7O@_'=-,*#\0\:B-@RUA+TP0N6;:2)@NJ
PD)!Y:/GK&GM>8C!1/&E_(U L^\M^R2VZ9.Z+_?IO690]<^3\I':(VEDE$0%20%U(
P$@KY!V?EQ.J@IK2A[$:0>;,^[B>)3XF3(0V7<AO ,M\^-;"]0?E4R;U*G;UC,T(P
P5A-P,5]JHGID#&B?R28Y)EB*"_<B2.Z%JICK_-RJWD-6CA0 C1@4M%57*>H$D*.C
PL%2UP]@S./U]ARX33M[;;:S 8+5S=LI)P#+=CJNTP'0M\!U)J?#.,6>BR5&$JXC5
P%3_Y?ZW(Q<*GIYKK538"+>5XG_IC)H;*JU72^^NP1:Z1-K4DE+XX6?B4ORH?:&+ 
PL/M%LW"4M$=Y&U(H1=%=":"15OTE;BY%QUOT^\Q%,6^J8-S@]O;&-D]$ _";YTE*
P<CUL"P3)SV=2.XR$W',,)2: #@FR.PG]E406GH)+*W9C]&&>UQP'UZVUI,XGM<X8
P@O1UXGJ?=(2O6;>0JJL6$JE<W,'2W^M/BBQ^\6<KS%6 EX@889(*'&SJ^".#2 !P
P+*>)G0L?A]Y7 =5Z7+99985?Q.8)O>J2D#A!40(([9&??9XENM)!1'QV.A7%JI=7
PX29+0Y%Q-Y-5 _:6<UYC2'HE#)$T*2J.0CWSF2T]J5JZV[Y(MJ^[@-DW"JNZ)9%:
P<>],5< E/("BW_N:3?&'"6>B+2;BAA!Y'YT^4#.X1FW0!()P?&K&Y3$) =P(+B_V
P3'J%$L5S20:M]%5>9.G7XKIACHZ5QP [<UNDUY0^G0/(Z]66T,AO8L]/<'>VF]BE
P;0*PU(OGT'2+-S5;X8Z<(N%K96,%:]M6)9] *Y4@>;DH=UW</R=A2 \7X92N%3#W
P027\4)\RF&IIZ:^_#9- %X7'40>%$0RIS?V.-<Z> G%3XDQ7U(UH4)0W((*[+%P0
P!@-%F 1.^0O76DX4UY.E D+OCU2FR-^WPQ6"",4'RG2Q@;]E"E*46>J('H"F$;%$
P/>ZF$EF+8L]**C*LG4<V@NO,)7&Y&WFK4F\WXD'LC! %.=O&UF-C<C^^4@.(2=6H
PFZF+[-A?=O@!>#K].4!A=Q0+G95NCK4]C\^^F5;0IUFK!_T.'*7*RD*5J V=?6X\
PM8W>L9B"-'%1_5;<QDV:)+_JXN01672B&N;2K6N3F*4@[@3MO'(29!KC2HPOOV!,
PV2"C6,D%-"TI78AA\CW9'-3R(PG@1XAUKK [GIGE(Y^8E&XR#"%][5@:_'1Y:(T1
PFU9/8*E*5CMEB$T9M/_[D#'N1W9"I W5SUU\<OVKK3D,S35 N7.S%)JG94:Y66 Y
PWY$/FD3JVD0L^TL98OCDR^*4X-ML4\(3%$2<%:">:6[&V5,23:NL5E:_]QW0C-(V
PX&_(8ZKJ_G%4O-A?SZ8(B0%^]U]1>L73J!,'#X#CSZ'M4U[S:#1IIB]I84!&AQ;Q
PJ_0/"D3N!(B7EL%,25][@V<!D;ZQ4N@.2# P %Z1V[R=H N'M)$/P^!BURA5GZB@
P7KKI([6]O5M)&[OGU9>E2G)BL:E^^&31S'IS  I(.'Y[Q;T-HQ8D/*([QP@+^G-G
P96E*#E9G8!PUSADY2S9UN\1+09Z=1W%/_H!B4+_E;3>I6N[?%$XDN*1)+J=/FUA=
P+$)0W;RR^BHXV?S(==F'3,\O+'-MD2"@X',T<%5\<"KD\["^VRI<^-H]6\<I<;#A
P_+C"Z8"=89'(4\$Y6%AL=24SY)ZA8=*BACC51^%X  WUSMAM7_S8SIKC@5XX)!9.
PTE6Y@\F5NMV,5C?O(G;\-?KHZ]G)Q(710H 6U]U+^09F?,MC#\HZO_UPNJN1/[94
P$1<+C3TYE?K=;@B K,Q^709]-QT0B8$_6N.:IX:2FJ'B*PY) 3B_=AL$)O&HL"UN
PR1\7QVRT*?->L!'7"0HTG:=1U9.U^;S@Q]F$#=$80>XCSQ)X%FW=G:!]W[,>5,0"
P 4A7P>Q[8/DSB2L:DS7\'E7E5?>I C(4B^F@UG#B*::>$@Z/XRF*[;H(G-H1I!E^
P]M'.#Q$ET#""-P4+<C28JMCXI?I4Q/+10X?:6C]MC%,M_E]:W;B*"5$W M,3L(0/
PDU&<UJT9Z"E_'.ID#9$E^ZG_/HFX"FO<KO5_?@@GF!5LJ#>P:C6ZRR&\=T%L5+-:
P;&6AV"./V][NJVC,2+7B;1/8Y4"W5NAS.QCE,:PG$/U\L%^8]U5SL:Z"5#LYB<HC
P1U3LN'$\+O7G!GY4(%V<$P(>X7U@(Z<E6--E/X7^'65!=#%]HY7O722JD2FRU]IN
P2]Y&T"^SF/VI&7]WQ@FMTS6$0+,PDYHK"1/40SN,T?Z/BEJJ0SJ>IOE]M);R 5AY
PP##$?V"&+O* .[TXP'B9J4N>DZ'I?@V$<"<=V6'2)</EC@95'<XGM3NG03=:MK'&
PKOC6?W;;^,3IT88^0%X*4>/3GE9EUE>I809_Z-YM6'S6FDJP\,]1::,[-33MP[%A
P)PO.=%O_I:B;F,XU'_>4"LQM\KY2+<<H+8_ <-9HP;I[.JLQQUHB29V*=C2$HDH 
PE<-KN5?8RJ1,<-$>3"/XM&@1(U(?;:JC;4QG:QJIV.>ZVV@O:U?5-G%>Z)SK6'^*
P*)1J&"V.[G%W[B]7 G+I;&6*N-)W>V ?G,K]C$VG?(\#')WM*%M'.TR)/WC)O$?*
P/H8RXWGG^QE,.JZBFY5[DE.J#(1K?>\CE7;SWYK#XY>U>A]2,I->S&ELD,=#2L+4
P*3(HD:))^*\%9NKCY=!6U,]$%C>LUG&G<B4SI2ZI FB()*8'U]Y;L<\1UZBD33JI
PYK;M_#[J%'23W[;E@IB%'()']-WU"E",FDA^:_:^1ILK1#%(J9E4Q9N,50R52"HJ
PT0>J+#X1 W5[H0I&QM<)R<EU]TVE*'(SK:?Z@V&Z4'05T>V(50>WPV!FYGV"QA&[
P1.*TRM?%=W-AU:6;]:I :F)'Y;PUW$G*,)3N64]FI^62#7L2[I.TZLE4\QCP5=M<
P.3.6-0LSF,). :7)ZZ'%6I&U:>_)0=PFX2 #"*+0$/YIJBS+LC@=(O4"F9+GIN R
P6P6>A"SXH[S5)4'?$;=37,N3@51:FJ;G#-  3/2GC>8+@+!9,]5H$,&2"DFF/?86
P09>.S>GW7_/MLAB@$PD?R*L*>"R547I@A]"Y%]F"ID$X1F>;;\Q>X"KP3+(H<<I 
PU;_41Y/.AF&LRZ=R(E^Q/7QW:"?2<)+LN3^JN;U"6+-A#DHBF6::_Y+^-H^ZK*N<
P$5=TA)7V+V#2YSA@3M+/Y?&VU[\#";>@XC6H-(SDS%$YQJV#@<D*RWKP ''1/]!M
P+I9CP22(:KEJ:ABB1Z@Q)0/A#;=U/Z9D76K8'/&_EF5T"=UT2GHXP_*/4U_%W 8+
PI*S^(AFM#).7I[/)O5"F5QS>X]..#3T$[]#&$I4_JIYRZ*3084T?4.UG<98!T5,N
PY.-IQ%' [?S)+!Y-CABM;,[63"7='EM1:YE2 Q@37X9)'N< G"?YM.W&SZ"-ZQ7;
P?"BQ)3=^PLRD0.5R1E/P5Z&ZRKH5H>B2@!@).DLA[H-?KI:P"(BL^\P,K 26"*?P
P'H[T](,9%=I,V=_QT&>FN;0)*62!B'X8Z6FBTICR2TM$9&#]SIU]7S8#.I&SDZ/(
P^F@LQSIY.H_BE4&UXHD6#DIR;EC,VN*R,;8\B>8^:5G)0>DDQ_G5D;3/"*Q2>HN,
P:^USJ>6 XA6S79US%?JFR?"4H^\[R?;DMA8";9/S40@7M_R.ZXO=P9QBIPPPXRQG
P;T2FV$;5=7<.(/D,D\N7D_1/9@#"1Z*":)D*,\5[,6FI\WEZ)"A^>(/.2B<Z.O@Q
P,];L-D&;;V,WZ$5W>AT2#Y<-I$B+"5<4H=%7"*5U/MQD3)_,.?H3*&YK<(09(L^O
PK?.UO _;6,[D\3U@U\;7J"#^^R]A)2UT'4T"B_2RJUKZP>3@J"GBF3-N2"F!3ZL=
P2F'?Z!#S 40[4UAR)'O:H\0PU&-5$X88\OGC(59\QQP''\>Z[%OW5'FLDYI=W>I@
P]XXL9<L6UTE#,/FMEX3;%)&0G@9&TDP5U()ZB9#&4SU7JF/(_=_ZAJA;_NZ0D H<
P<K1>%,9S F2KUK>-OH295"2,-P9K.Y:V_-<J/ !5O%G5\VVQPTEOV*>#RWA:S4$X
P^VO@!A[JT8S27WZYRU\"YDX)LJ=G 4XF7PI?-W0JSB ,UUR!^8$+Z[*X7("ZSQ(O
PQFS@,?2K@]H>]%O<P?Y00\V*X>4? )ULYLO>[>*!Z#4I8P E5<=+1NZU6/;__6L'
P0.D)$EJ[LA18X5HEMKSZ'G.:J/<^@K6QH)Y4B(L-\E$YJ2)Q)4'E -B"!P\"[_O)
P'@- @\( >.YD'0 C%8%/8P6O!F5A)JVB#"/=BSU[Y1XC!=MUM\Y&0; /&'TPEXP 
PE;!Q:WQ<[R1@S?3?BH$E.OJLVF<%H]@6O<&68J3!L ):RRJO\;H:6*")FO7G;H+!
P":BUMES-'MR/!9I?C[2JT*?,+0_9J"N(.7RA%IKWK',+*NUSP#$D7CK85=6K*A"T
PNM1;6#L4 \PP7DIG;Y8<?\I$>\<SEM-U^^0[WNIB4 \5381*OZ[@>:[.!%X>;5+,
P1F)%POS48<+).*NW;9(0T^;C#!)<ZFH<RJ8%3D/2_J2<P9V72,!W?&RHP>4*2LKM
P:K"42E(#;+=$Z)"S[22%^5_M6-H6+.5='O; >O<LAA@NMF2!'WZQ[Z[W9JERPP;+
P5<T,9+G[K-UTM\5$= \,]+1>EG+D%W:S+R\S)W)P=UK] SR\(OBHH$6:S.,NGQ# 
P7SM5P6-I6'Z[<>3-.9:V4A7?\A)BAK4&5UA"LRY$]/@:^:0M'J/D8"=, -UKWGH6
P;_J\^2 E)P(KBWJ@?99]5+RL<6PL/NN&=&;LI,>#8E!++?NB@&!(N8;4*:?["2OX
PL'8ZU+*EK5+#=PW^D#5B)-NR,.""H>6+.(.0ZXK1@"X <<_ 05DXQQ:U,AGT[+DJ
PBER>D%Z5NJ!WNCV?L\6&LHP/%#V4$<+<)HH@\$NI:V2Z#KDB[IQ)!T]!$G@VM"0(
P<N)]+_J,U57G\*+FWIAM85KC/M4&;XO,/G4:1*8=AAG/Y!*.J[A?OG#T#(\F0Q?Z
P-_FX5>>4]\K] S1K=!LV+)]1[R>^%/W#:["V.A=1##&OKREUY4!1R$7M IX $V3Z
P1DFO:X("D3_7'J =!1OLQ,]!MM_[/%B)*+1UVP?[YK^1S7DC)Z65FIEP0$HVW@M-
P3KI1UC)3VHD\;R?DC6&.B/H.H24-OT+:TX>@C>A)RI KTF28.J*'^;'PVV#O2RE/
PA/4U12;V]DOA'#/5"JQP['^"Y'+BN=*V@U[P.2N+EP+ZM5,V1+ @"5J/8W>,R)1\
P_ZYSG297>>>V1<+/=QJS,+O\Q@8=IM>)L_@"I^+8Y,=;5YWGY :G=Z'.(>7\&/$@
PI>YGAEC<8B!,+.O);A&)D*X_A((U+MJD<.W3"\XF094I4>*.B9[^>,80Z4=D& *W
P:"AF?C#D^"UP;-3+:?:M2T,>+)E%DP K<"1K=,6\X-[,*#4[CL;-EM;ZAMN$'=3U
P/9'CA<>%0%S]S"G4CUO\1G/>6#1?<L +ODK "DB:QSL9!)>1L@!1D87D/+EJ><MU
P:GH@B>WP>H6&WLQ<J#]7 JV0"Q,7\+P?*@D#DX*PC,@?4L4)2BMR=PFIGO(HE\Y!
POH$HHS=)EE/690N[V;7CZ0 5(\6Q-9?F E_TRS:PJ4T<FOJ^+J L;.C!:]P6-Z\_
P*>'&GW*Y\Q>)S*<HZ!\JG@!T"B'$_6A[5+KEM[&V1:1RL@?(_@/0Y,^)3A9J2$7K
P54LG_J=LWTL %T+09H^3+ ;\CKYLG[C>K$LX23O^R2)_V'9R8B>@!1&1*+YP(20Y
P?/3CWPW8V#0AMK__Y>GD_<"MH(G_NL+[:OKC^H+NL.:<$.^F% D!-8_7!BCOC(F)
P%Q0TOX%N?SZ0S#V"OV)/(D\*<$-<=-FH- \G9')!/T;[EL6$,8:</)_OX!77ELL+
P:<ZT:L5]QK-A;55U!1(LE+%B:;VQ%Z7A$E]7G-%RET.1AZFP:HMN&+&U#HY]T^>.
PP-B6#VS. YNK+?J"&!K$)[/(;?8YW3GI;#&^&$BR)2&>NFU6<\H[GRJY;WAE(SW9
P%$)VVY!I\QWL7E282^&[L554$'+?"?@C!3P])T77@M"D6_CM <E>!=P2^ZRAS2_!
P[(G9VXV'KX].'JP T\@^/@=S!U=(L#P8^HVV^!X,_@#^D\V$S#0-)0>(IU)#"E5-
P"%=OM[9F%1YX>IM"$T]^?4]."B4S_!, )OU7F^*I7<,FX ,)]4]_"]8IULU$#S<!
PY11LF5:@!9'<%<=N-/.<[XE/?.JDX%@=-@T'N]_$WW52(T.05YL!UL?7ZD"IR;Z;
PDC!%(^W//M]W$,X'X87,B6CY .D[VZ(A&*(HYWRR#JM0Z4-K^)/$A<&^J%'I1%:#
PQ4"@'A=YZ[D]$Q=<BP+PVO/WZ\'22LCD*YOGS*-)\TE)_YVWZ4S5M(QGO&HNCXVY
P3\V4<Z5B4"HVF7??IA<3<;O<U>%:1:.D54B#PW"EH%7GD'X&=LQ <$MSK]NY#@8X
PB[^'6B<LIGIPKN7_-HO:$%JX#XG-AS=Y3@UHZ9SNOJ<8:_#.NY547'LJA3ED1I]@
PM8&-3_OE]*YG(FJM&CC>5U@2R$]J%DWIV-I7L$YG8<4RG<8+-O.I(I6T0O:MHH_H
PF/$D;XU-"I$C:E/R*=#K.7O.:-7-IZ$>05!3POZ^G(M;!;[/_*%B/X,C$A6;'R :
P?(Q,3/ I[695M,JI9"9?D+Q15?L89"I%A/K=)-UJ?P:E(ZBB,)T?*YGBR!%J3LWN
PK$1C5#Q_FV_WXMH&=^S_%*IYG_G[^)=<2KLF\(L@_MR0ISG+8/-DS0+JRJW5A5J:
P_2(M^,D4^6;&VA&"@=+"^'(7-Q!V^NN%G5TB'E*:1PHA[U'!I"1KUG894O?6OI)G
P+.(+D.)7[DE'Q+GOXZ0WN\<Y<^$-B@1B-M>O0LKK11W,86RQG[B=-W%RCO7-5K"T
P4RV-C1U5&J*,E\]($@069;#Q5V[:9:["^%K4PM2 LM[W[Y3ZFI/P3 ;9^961%3AU
PL<J=/X!/:0XFJ)^#72)+0Y42-=E2A@YC+JA<A%3G$UKF+$T2H$2HA#Q4PY]VKJA9
P$NJCHN\8K,3EX8QZ0\XXJE(&>( A'R$$J6!/DM4?I>H[B;%#6EW:V^BBW*VIZB,"
PTQC/(E[/@)7W9=^=&^4'W%0+SX\= <5>-4G^29B5LTJ_];4'ZNEKD+-6#N76M0=R
PW\8 RM9N;/*/3E__R;F=_MU. 5K_-1$\_P*^7Q^+,R B;7W[!V\K'[)!$MM_\0.7
P#T7IR315"7?\L;-68,WBD85[L;%_\+<+P[M2T7B!T@G5UN;*9Z?' =_NKSHA"_=5
P?G2[%B^%N06Y%4!P*U504X9_2-!=N2P-)EAPU!5-*%\+%]*L]Z=K%610[2KQ/^)S
PCU7VH$FZPK-/5NI5;4_4KM*HSD4<HG$6Y)2?--ESA+ S21 TC'7<T>[(_BP_);+%
P?TU\T*"M"Y,MU2$P&13J2%%<J7 KMY:9]' YY^G+RQL>?VM' +;.UP\*7P-KG>J+
P?*+ _]8!#(UP%F H5O6HL-;IAHICV5%9@_=-CY[2E07!7^3OJ6B&_B09P'A%W&;5
P)BNA?7I^7T/.0\"=9'RDS'9"67="]7-,ADY)'EWXP3W_FKLQJ^>[1*DR:6B9[AY%
PM(I*7M.ZZ6N%7Z,XR?LL0+PB2!AO*?Z;W\O=X2&S&]-4EEKIL8#,KC*!O"VM#>'K
PY8-WIL92PM;QC!=3<_IK2/5J-EEL[)C0]*$.'SLFLO==7^?&V*@[L"CHCX9+:!F'
P]&UK6!PR;^E#%M88Z><A(HF&8P%*&#4V<<V7C<-AAKNT4NCPFFO.!EK^L8PX.8QV
P!!J;H+?HE)[2U^[53$(.Y*P>'254KSH5-"C)WT#D#X#>U76\EA-SR*;:"S'Z5)6%
P#@R/F/:.HHN:R0-8XDX"_@T[T;5^ODRA>)9V+QX\E730200\,+^[E%Z*@0V#!,/@
P2M0.63<"WZJIJ>!)-\5"SJMF*:5ZU,6/CDVEY,HU%^2Y(FHLP'[=97(1K, [G/XT
P35L \VV8_M8%2L5^;D41^GS_!_7V;ZYP]*F"ZE\Z#<1:-0NHM[Y*C77 :#&UC0+O
PH/3(7S##1)6$<6['N>TRM?$U/'LKBL\<+Y_9/0V+0T9]+<23Z7DTB5/\/O_4SS9(
P_=KKQ>?RGQ35A?&)&LOM!D9JOZ'9A3-7#$8X,;5A)!=Z90N^' DRO%!=B@BL2LK;
P;BL]W0)B&7:@5@C?09?:!JV:9T6I4SI>FM@I!C]=VA8)*UZT;'#3D@6E[%6ZKY$4
P &(_NZ'<[LF<@3-AXK(=1+V=.J!KUU(#X$:3QTKSU$B?G]HS%$.^3A3'%W1Y?M_@
P40K7A\:PM#T1<])@O46:8>T; #:<56-'5KKF$WRYI:U\>:3,[8HZA[#BN5YFCTIV
P!2!:I<6-^E.K6TE5%\&P!=_UM[?6![W(5,# =G8O->.DS<]:KY]7M(7@PR<P+J3*
PR0J<H+'SP[H;@7R)8$149,L6@17[=#GA*#VUYG=GVW<>K:2VGXM""JPV6G-.B1$"
P_>!\C?$CG!O.( J,[8@Y[:3A8)7:1G5KT?9P2OPC!XM0Z=/?W&7UX<(<]SG6KJ1&
P0"7RYMC5?[4'VL_UQ+@ .2(UJ(_*U:+G!??X=8FTN^!6 P^:M9?CAUT:WSS,VRG)
P\1."6%#%&H_H[A\' ,J.W["RIH2C Z.X)^)<A!\>T6W4R%9_9 NBS'/@)CSLIR!F
PZO(/B6M;"?.DYU]6-.:6LT49NM\<+@W%IC=2+G<G1;=??V8 0S3*[Z/.VPTM3-$&
P,4^DZ#4.\I>BH1%J[@3/>=V1X47EU/?#M=."(V2@89&=\I/V5P@ZTOQ8=\'=RKVT
P"_4JKHXV"^G)A'2RT(TTH"ST:[9U>?)^!LA27WQ*_]]9O$![3,"A91K.QR.!_)TW
P)F[1*G&*#DJ/K<96^M(+=]'RN" 7F&LZT55?#42?);#-/N60FYDG<-A (PL3]WK>
P&'2@,NMEK5,$PK/5;5DTTLH=T#=H&@Q=ZY6+BV0E8H],IZ X]8?:9+TS?Z^N,I+G
P?H<V^-OM*>VTUUV;*35)3];VRS0#].+^(%U#O@SNOY$[&Q56RDN5"1MW="9:Z9OW
P1@R:C21'B6B!B:L$74OEA#6^9;VFD'O4>+K32?C*.JH P35O6J%!C,28,T_1=ES;
P]0[([\T!(U;K<5)QHGF4%M5-/ MK5*0Y53*:%Q?W!VU6+-=0C,U;T:AN/##&@*-D
PC9+E,)T>/1>1&3N'^36O]$V6^+ ?EA/[7&6:]]HO4D.7&AYE)_[00U:O9Y1F"[Y#
PI,IDB"L-&OEK98[D/DDE_N_8#3/UCHD;7\_:]N8"JFV>:'9R:+MI7AS\B)=U\90&
P:R6CXEF 4JD2$39&)BH\9T]O,5PWN!EPIZ#20A43=7 %!79U:HKG*Y[-N51/_AAS
P[ _.#71H- MP"9'PL",CG7;)-K9_\Q[<^JG8374/S'#Y.P7,P6,F%R<1WUL'RV*)
PZ^FUU%+EL%22E0?@HUML GFC]P;EQSUD DF>E E(H'YZ^P('FU^$VT1 M7(*K9+:
P-B>B1$H;23_/_Y%45E@RP944RB;#8]MGZRKM,KK/V3ICYVD!UN9 U)+J;C+Q>7O8
PN+E3*4<DS.I/++6@8^4Y@*[#02@F('I/? O.98O&$M*^HVJ8U0AKXDBEZ*@C/2_C
P!;U>B49BM/#%LY-$&='[L.Y3=39.Z_3X?')9:]7=5;W:\4_>2NE1S#Y1D@'94-[L
PAMJ;MY1Y\B]]\?.L.!:P] J&+9,$M2R  ?;QV<XN/9T%X<+D47!"&NM5(E;XI7GS
PO<GM5X[7VE3%'W%W#65&O(* <B@I Q4NN?/ /VP1=_R>O=(K+\V8\K!_O\2YCG!=
P&R,H%1\8IC$C =M0)X@R*NOQ_?#=N2UL<&7)M)6>/?G.&K4FN,8_B4?B @-<T9A8
P8MUH7HW>SN!18_LT#-F!;Y8UAY5RQ-)Q='GK?EPBWZFE%SXBNNP>*Y*IU&F&P67$
P!V6F,IUD],-;L$>B3=N8$(\EE;UXQ/ZYA^HH]RKW:ID@7;K>STJ6Z9:-%5MJ4*>V
P5\M\5L9I3ED,&?_F>)5M*N)'NI*'.-^)&5[JM45AIS<L;LFO4@QW[+Y'\ /9-9AD
PV3W)'XKPD9W.#9U\PUEU\V33+_3[<BP%<D\YPMDR:D^LYPN.(8PV:6=FR\_&"N6T
P_5CX!\$%L02STK 2LH'(6.8 OQN1Y^(@MICXC;,?.7&!)E>%$[23E)+)E$J$DA9R
P4VH-Z&,W\T!RU4)9=(C"APA<@CSDJ'M+T6&0[:?GM.@.Z!6NOF[)ZSCZB0 94]6F
P?:0B9<3WZ@Y\;IYS8@#);Y]-:3>I,RB.6I@F6<V/I7U:YNH?0W4 ],W-!#_W#0$X
P,EL?3OVJ"*/2%$[<_0$QFLUE ';GR?RVA7=\.,4@?D"B-7UBA@JX!:FUZ.PRH=0I
P,O!K4*5GVS4%?QP$BB)I%-D\,; Z.9*0)X">+))E2[SZF"V*0VD/=2&SPC+ +FSF
P)';W0=U (:@(H1M-5GO\F',]L_U_PO+.G8X?<7W6;>M7(]9N4:+-M$F9^+PO0OO)
P%?D+9($RN.YT2'%H(/W>MO<!Q,SKC'Q"H"5+PS\DDDE-T7\'7"%_$?Z$J]V$FY/@
P[%_ K^^FSF*FB6;/?&O9.:XYR<Q9!< [KJL:9-*;\'(=JQV4JKE;TDRGQ-(9V(,!
P"P2:"1 BI202<^O<WF=Q)I&H%_42DQ ]U3$,I> "L1)8[J[RJDI^]KY.-8*FK!Z-
PU'DE5QJ=K=_AYI7%D,X$8-'<*0Q_A*EQ^5:&?T2DZ)>[M(E:I6Q*:8X37J7(B(,Z
P!;*12$I^FQ:3.['2.$USH=$KS]WGL\#SB]VNO/SHE')+V]6QG;;@#/C-G>]$N7\X
PL0%$K1#/P^C@"(&^DR2D\;TB%VEY:2Q.(Q$GUADR'S"(-7CU^.L> #Z&)P:PE//6
PSI>_4UC9MP)4S'?__  'I5_$Z2E;ZZB2SDG:Y')_M9*4CF,S\=,>E&QC^8>L//BP
P,Y<DZKT..O++!J$#C1Z?%[+R6(OBKW"FV_SSCMV0!OR"XDH03IG:E;:T":_0NX<)
P@S8M6$Q0KZ1$$#70:@9FU;V^ 35<>]<[R^4#X>M_\= 0._$_CP+A@\.2Q?Y&<83(
P.KZ&7A-78'0V5W!<X=!^<!0'EH**W NN.*T5/:0QV[.'2@)2IUJ/(IW[>,^2O,Y?
P3G_7ANMYB'%HW)%=J&*H668OA4(#\"["4DH>;D((ON:?1!]G)9AE2'E0S2Q=KS4Z
P5H'PLS3+[5BB.K/'0]3448DG==F6+O"V7CLXV'J;^_/Z #6R\DZ9E.6>>$36G687
P#35/HO3]Y2^:=\CX:(%$34&":,EQ!P?K@EA4!Y?!'K:4_9ITYHBHH3K;N7D&YT.C
P'^?)^2QY:-2S3\R2JE[H,K&89\*/F]]@2%47;F\-]!N)PT8"I'H780<\CE:<O=_X
PE$!?PVS/JSE%:.&AVTMHE_P--UE55K1Z]I(FUD^'#PQ:QAO/2H;T[A'M$DSO;00U
P**_VAA942_ZJ*4:(EW;]>I9"GP9YGX[W$^I"M&E=\T[^0NE^/]RD;SME\,134;_U
P%_:?:69UN.2N/"->4K$BO$LB6#Y>Z)Q8(EHBNKQ'I5J)#<$23JY(O)W2[E#[>3RB
PL/,$OV4"NC2R,Y#SK]D%Z-?EWB!&Q:%.[%ZNKH@8-X!(WW&-9$9)5DRST29O4Y[H
P<^EC-O0$Z !;_)'B=G;A=-U%HI97#/$.\]70ET2ZO896D%0>.*WTO>G)SB)]2'=5
PSD,5H>!-96/!V'60:8A%HB5)UP!#Q#4 PK;D;7;(W';MK!:HSO2ZY +XGJS4/;(*
P\PU>?XGD9JP,%6!C2(=NP'EER!F.Y2H]N9)^)%<="+0*"$/02YSQ1S! 4XF=E@JE
P*N53H5%M_8AN5KJP-D!%]2YXI$X!>/N11EC(SDO,@-LT2S7C58H(=<-0R4)'F&#\
P8B)W)M3I[_G5KM-?AV@:U4QA% 4H.C7-LGM)1.W3SSP8C-X1'4R#N/3Z=#$JV/N"
P['>J]S2=.[&*44-,0Q:X_X.:BXT]\<*<_BA7#Z_&1)940YE8JA5Z2BJ:Z"+=_WT2
P=;*EOG$:QGZ .8A^KTNUT\7M0DX0.5G#5IPV8UQGO_IF1!:<2+<*%'\HC^(-%NNY
PCTI6*5&F1IU;=:3:0?%>')6RR/G?W,_)HFN@\EW"[MI.[2&)V1QCB4B)-\#?;^1;
P'?A7B,W'9EIJC&;0547892G+E /E:I!.N]9IW!K6PG\1$_.\R-TF[B'JLX=XVD(.
P+8Q%Q5$7?[\1]/8G0)[6$1G:QK>8\!FOX4@PF$IA%6D9>*-7O]L1PEZ?K U>*8\!
PG5DK+.Q3']"WT'Q9^2H6.TB \4QWP.QJQ-B<74-]A]J6<5I73 ?.'O7-M>T.)D:E
PYPY*0@J.0,9>62ITR!6[2&A>#+[+E0)G59HLUDS2[WK<N"*.N==Y)*7D*4J9VZ6K
PDB!(L;LK0LT,<%>:?@CN/5SRB J(&T3>EUV410CRZ+A'>.UEQBZ?5ZJ.L6^TS7X9
P .'R]4P)-=YO'CL?N_P%]D5N/=2Z,$4*!Y$I85B8H9+.=BOUV@Q996J=;L0ZN#&+
P/7M'1%$-6\ZR-!!) KWX:K=S3%2DOF4PJ_W"[*@/M<#%^CDGE7X9V!EGF>Q6&($9
P^]X;$4=B6#CJHR#IP1_^5F/F+$HC-N*!*%+:'/SDZ=*%8YV,6=>]YA&Q_B>V66&S
P<;G_]-&9&2P35Y$S]P;"4&'MW$<S7$%/+T> E]0H"H6(MGS;JL%=-B"L,R&'F),4
PY@Z;@(3B-GU7.4+$S4>WL"L]#BAP4*ZF20WN7(\T&HD1>6">00DFP0].))"\[,P;
P38/BK8,(KE)'9"(](C/&(&,^"@&13QONDD*^6>#; S/A[.]!:EX\7&@50KF3T)@1
P?>0HX7"_[N6FI$11_I (VJ9()=:)/G<'Z<P.UC+LE E:O0MD\#G,KQ'S2/(D(32U
P%-]CO%</4&U<NR8]P.3O2 +-;(X_/VI(PS,#H!X\HNKL;S@&'Q*5#,VK%R41&W<X
PG%_:L'"[/<![C#?<Z39J[(S-OQ"#<XC$HX3>5/0H_8?S>@'QK0"E:9G97E2"(;0W
PO?_^FH3LAB0!=,V2#NK9$1#;WA]=P_AO/J*BRXA"%E,M(*U=@CJL]$QR65#=J]X 
P"IBZ#E4J('M@!;" #3;!CF'@G<_;_1[X(6TT$,M'>H]YK4]"=\?4 0,FQ15*["L9
P3!_MNF.WNZ><<9J LL&^_--)9QB6A*&9FK)Q/ !U^.V 501JYL8;L@8ZS@?Z[/8;
P"SMP6<.H,E):C[0>_D&W9')Q4=ULZ4N92;%-!W#F).S[OGC]^/&_M0KK/CHP,#O1
POI*X($;^410#D9$X&9AC'NTE_>"66D#7AQJ:G6VPW;V?<?- ,0<6YE^N902<U"M 
PSUWS6V'9YU[Y 7:=E=)<DJ7Z@C,$3E.N8!+BQ@0/0W+@G42C=_KK<:@>:H\VG(<I
P1;O6$7/<CT?]R:AS?Q;]WGJ\E<ZJ_#N7BBBB(1[5I=*N=@Q&1)I6#,O\=MX48W0/
P?R&0Y>ELZSTNW]/M.W-[5,4IT/FI06;-1$PBJY%0;ZF6M9=(',QZE_D6B9<0RSF?
P+G<K6+N-U*#] IJ%QE<.O&T()MSS[2":(5DT4FKUZ=7"A/8NV8NHK7S<V1I70D_Y
P>N=S3@,T32TLWJ7F6;S9';</(L6R1Q@CRO3BAZ .*-T][6J@@DJ9I9.:YZZ1(^S?
PH_51$+Z/7F#SXKEHYE2;U3/UEY$<[N*-ELXL5H_PD4RJ2\[9#?!;YLH8>#?C/)FG
PINU5*76-Y49EB?5@#MK8DJ-HV>-F^'>K.C,9Q"'%.BW)!:#-QE& $NQYP<IG)-N;
P? QKIQTP$./%\523_/UV\G4U_UU"8XF)4URRDG]C3AFF)AD'<*;M!#[@RS@.DS3[
PY ML69"FP1LZ$Q/SP\=&T2P-\#OOWI)A"-&,12(JA$$;!(@0FC-\KO"=6PJC*A"K
P!6PO)Q]4!B4"^'H-0U?JN06%6C]VCKW6$4M=*V[]J0<:>3TL]"GK@,,/'%*:Y'K=
P)!,_^C<_3[LZP,E(K@#?8*$O/UX<A>C]&UN%=JTP:YS&A1B"FI '7P-TO;* #JH8
P?1*XU=-)[PA6_OO79*L#U$M9HG.<[GG&H8E=G"2VCVNHI(>"^!=<;C*DE?#HPKZ\
P: A$L+G!L'<9,PILDTQ#^'3WTML.5/NK\,2"L>ATQHP,8KM@/J)(. 5&R(Z38E=*
P1X$=>^2M$U[LJ\N&"5#\!F!/^0AY#%E,8 ]GR*L!8A.^^SI;>)N.*,,JE$B;&P/&
P18AVJBWOH6/]+9LH!PR&+\^20"[0R3Y:6*-3J+&U#FG,\FS^. .WC5B0'5X/UH/6
P(T*9'Y4,@YOQ('?QC_J_RE7%ZE85ZW,QHAV]OD@?J9<#;I:6IRM]&!S6D)[]6)A7
PDL/;5[E">YOV1RU^6#UY(.Y)F@!L&?*?H-4RU$@9A7 Z'MV<X/^.XUL*[U,JL?Q@
P+M(ZXGJ.SIKY;7ZQ,1%9$%9F#'@PTZU_WE':Z<B6I,.0XOBB/.7MO5P@(N2K]U1Z
PSS3L\ZTQ *":!!$%_>!9\,\]Z@:U,6*]Y10$)N((4R7T@"<\GL^PUDQ'GT3H09!U
P_33!'"/^+SN:#[&-+0C,8])-_$"HWWDCI56PFHRS 1+U>#2<; ?DU--/UNJMK8[5
P##9?^3/ZV%IA?^SI/RSM<W@7YO3,%J79V8"8&=UNH5"/[X(>)FKV&LU<>SWJFX:0
PW[.GC*=5=$>B]'A,:Y[!!='XYZV7_2*<Y!C%((3_,-:.P7G?ZP0#'KG.#!0#$)GL
PZ#R8#1R@$8C1QR_9VYFAC)FDRVFO.AXNS?I2/OP+PHTS^X9S;;",B1>2;<G-C7OT
PWJ]ZSW\% >*&<9=Y@OR#_Q2]O9GP X0[)*,35<U_A"](.DA+P%P:) H&EW.W^.((
P\-Y#<PA&-\(P(8LOI0S27<B%*:VMRU,)K%!*'V0M@7]QS#S6YE:&Y%GEY"S/=-/9
P6VA/"$Z]\_&LE[H<[^F?B$#6$QW6%'(IW1#1Z0M*HOV#Y1B61ZV/40;O)1).#TI5
P_K;#ZLR@'&WN8YO(:LXSN^-F^$ \DXYQ&%%H03Y!;AH6QP;"VC>ZU^6EW$(832/L
P(/Z5<9XN%ST![=93K/S<V)7"0:0C:P[:#488/L/9V$"EN6X0U23H,\SG.9X:DV\Z
PX"C>R<H!^.98H3 _4"1">BLUFVPNO6._,>_\BJE?CMCQ_FV->Q(S56HH:U=$8#C&
PH)'2MN*Z7J'5YQ.3<<NTFQY2SA+S(1^ 8DIPU87]@+^1@BIRU,T\N03D8QRXK-P0
P;,[6,MJM/;_RK28^ +?E''OQKR!UY&?<S7WJ&[*C$Z\I?U&.BZ!)^4"RK7N V=H 
PJW#(9,)/0A0,"W>XM#=*UU4A@QO#(R<$)<BSH(/MIBM0U!I4/8W"02;UI.[(9RS5
PT[\LO=WO";DG47%V\0PSVQN".6 64^EDJP<QI:>A%JPO-Y9ITOU%?.,XI(1,]ZAL
PJ?K#Z8S=$>K\M@7I4H5K4&*\F5;6H%] ZX/9FJD-[=X\"2QMS649,8Z^ 5PM_*A,
P Y0VD.Y$*/WXIN")I\,.Q5 B("5D8)&A%FM?:]V=RDCZ:=A_:OJ#Z3SZ"$JT^N2]
PGP?U7TSA_8_B:(*UR891.\"Z!NTRTNP9S)1-[+ ('M:J2^I97Q7'>"<>#8@V+VQ-
P&SF_=?2]2)#QPOJY#O@H3'OW-LSY$I/Y(30.*-4JQ3U2O!Y_CC75RBK-?+N(OEI1
P@CT^4SZ82*80DR34RD[<OZK=KWW+5$:&F'8+,8<+]_FPGT%<@"E4P]@";(=YAPM4
P5KQ?LT4S?) PN1,8+;^P568/KEZ9B, 0H!Z:,)'76MX?>*EENB.ZH+PIQI0H6=$B
P8RW?=VTU]@7$O&Z ;5[KCAOT%K%VYB9NH4THYH^ !$#2Q<JV1X5=Y/U9CS]?BL\^
P P<;7B!XO#J34)I\QNS2*CL5D%(6@4CG.!D%2ARM^)T5-0 0K%T3FXF99\E?0%!.
P;AF81[H6GNO6"S4PN&ZD@:>(R/%S-TORJ%8N,,)4E!KU]3!>$Z'EK5>M^3;SEOG*
P,/$"-K5.3@2.+3GCZX3?L?'BI'G.UT9(M/W<> =JIEQ0,C,7!*7Y=YQ,?AQM,IK<
P.Y76[DCZC7!3:VSSDY! ZV<9ZK<REHF%^C P;X"4X;[]MP"=I3>A[PB0]18@:&2F
PO]3A;-!P;AO"ORFI!9F@'7_)&3W*YW14"U_J3VH&YKE4A9?W9OX.>C0K$)K%T9,]
P*%KS8^;28K.9#3$,=[F?1"XQ6SK69$\H#.T)BQQ&_VI%62%^9#$DO+;K<7U(3[XB
PYT<%VEU,]HZ1:9'C/#[RS$SVS&XJVS'?B81[P HON6] >_11&]'+QJHIC+>728UY
P2+H3"<^:<Z<@'1O-&0D"ZN/3\7('.A!?B-H;"6XI.<709!-*;OT2R#)'X#W3(S=B
P8!@%E,MH!&JQ0;A>';AM@P^C*HJ>B*^/]R;&"XHOJ^QEZ>\B\*VF\&!GE?_HKAF2
P@50\K@<V/6)<@8?L"WN;<M[8'R!/: ,])&API6*$%@&NLV%O1#:0!&Z5,'E&2P%8
P\/9B%(AO9MEW1D0;__+R-CJHP W_"NS/4JOMZ 1'50:VP)K(Y:4-@\@,6NY'D/V^
P.')#_.,D77OFDP%NTFY<#QC0!T;2^'D/D-2"UYVD?Z'@X"7#.#J ]BT4/)Z',JR&
P?G$Y]>GFN0V/.40(;__,+/RJG9>+GC369UOG2NTM\H[7V/"XAE/1Q)MDJ**^N:[X
PE.B.F=-!. RSY'''T,2KXNWM2D;C@D_5CI"N.5X[W>0DAH12)3-<]XY6DCZ5G@7?
PLV\%Y*99(/YAT7VE^(5$GM_NY,D8@&7P!^?D]U)E%!V NX&"CTD8XP$((FKWJ5!W
PFBJ5;[")+3A\#C(CW/_<+,>WWLTM_"G+OP6R0@T'50]A;N8C+E5N%D6U3CG\3V+-
PT1%2O.BL WRCO?:<]AA[4PG*D_  X)3,V"04"9ER930VLXIRG5]GI'+.H'XW;SDH
PQ_MFU^6)?=1MG&0D?\R"0O&*QK57:7QPDN$5"!HQ\1Y9I0^P[%9?KNN^G,M@IZ<:
P721RGYXE,X-JN^N((=A$&*B>S>2Y(<H/!X]M&^ICG0/#!@8B#&YCHHL_VSL=^SHK
P6.<PUA3KF8QF^A)I(_D%]0@R-NS=>&CX")"M*UUU#AJ0-*6I6R;AR!VF4'VGQNT#
P:'F98S,,1^]BR)\--5\H#HTEMU G&0.[;D7(@]R4P%[J[RMU7"KTW)(0OW&9OV1[
PR+(T5V>!S.\5MB(K8'#^>Q3[S4=#8BESPJW#!J3K2J.!/>J3]K!D\D9^9K-7,,I 
P3YW$_YXRYS/C2S<D*\_XPHV0+[&C" !?N5;D 1N8J">KXE-C'QK28',5G>&:Y,_@
PV@:9*8?N?BRH6 J6<&/WZ[8OH:G@>->/I$A6)5<'J B\51 "@;WQZ#PIMM0E;P] 
PYP'.6-X-2&6;9_S#W[E"16UB:2RTX),=AMV1JP@_ENA <J)-0<@DO@W)7H=?TQR9
PK;:29Q?\M=%IXJ3PSOJJB!$]JJ96WVT'F1%:AQXW?Z\X[G2>4DW&.DG69;VH\V".
PTA0]8:F!P-ZE8A Y'U8H"4=;C:-X;74S,30ZZ-T5_WH$X_&(O-TL*;(3ZJ4(QLH.
P9D1'#.$=FO7=[/DP7BG$VQ,<M-"ZUU3W'+-5TV][A5@^W;E%"Q.D>,G"EZIG:T#;
P5O1=QPDIUTRIS,4:/*X"IVV1[E$>&5J76G1L-HPIC+R(%5!6CO^2A_0* 4O*:20?
P._)OGZGT29:-J\!]?$0WN.H'9<D2Y)U:*R+^7) !5E_#0ZAQA]YD<+N@Q?]Q 0/(
P*L0D77G8LB(A^@!TSH^[)T9:0:<4X9TVJY1O;2,"<)29VS,:A1ZN/^%;/MAVD$W(
P%L#0WJD"<>,>^34??8!"N (U87IH.N@%F\$;$Q.#)EY@X1Y)DJ*$JYV5SJ/0VVS6
P>G4+M56/K-K?4\I;5W222IPF9WLOIGFT2"VGIZPD5K0$A#;>FH\')1=V%Y^9"SK]
P*QR3FU[0M=!XFG&1-$3C "L@SO8&XY$DX3!&!MY.7WI\ ^RU7"B-/#\"I81F$CUU
P#%(=30D\4(0P@X*O<HUBVT,$S[D3/%W^:OK""<N>DM)-O\1KTHQ?@TID=?%O?IR/
P>O$8XQ#_&/W/C-'C[=FZ,<0/3VZ,*VPA=4:CS;$)\=PY'\X6WA]C+O$]+!!8H=UW
P@67/6M/G!%/?SCXS#Y"@U)E>'/.X<<,>@$\/DMFG7MSH6W1/4U!8[]*/(<HP?7/[
PJ2T@FKDWR'&9WC/147]RE[NV@ KV;355E74#]=G41+"9*#, QCJM*Q;0D,6>F?YJ
PC4X03GD>2V33.7_2I_%%X9@M[YQ=WE&;FHU5D!=2>9WS[,*)DZA[/(8!/LL_ZN_?
P*$@W=_$ATJR9"1+DJLJ '&?%TZ.J VWY#<'W8'/=W;U&K<QNG?:RJ#@,,-&8G(37
PY+W]'?R>:$.B&A#4CYD\?H/"RI0 _$23Y&JV!4V0Z.2!)Y1,^!,"0E19:3=CO1\:
P@G/V%'_CM7G#51@"(CZ22>9,,Q3Q/WA.DFOW5&N0N#/6#9:E^ #ZVG]P9,*4/0R]
PNLS-H[" C35581[=JYMP-E5O7H$BCHRC*/O+]Z]_=_8#CQE_I;(7'DEG)$B-SJJJ
P7J4BN>OH3L"+^I4>A?4-T) O7_37ZH6.V(/JQI]\:LUV;7Z8:MU-^W:\O$!&('5?
P>LJ)Y#M.P\3(9(U.!MVZ*X(P019NA2Z+2M-[:[P9J:F\XS0U6[S+O2*W*E$*IYU&
P_#M=I!N.L:XKRT.?UXYS^:OWZ]V%+RP*(HP3*JN&/1B_)1WB'U )0K*UBO;8+U57
P.;^BX<;&0O&:UN",6]E^&GG AXFW$%B@FO<X9LK#, BA8!?F8WF!/Z_ )K[J8X .
PW;0K=>=7+_U+DH)7S'WFIYK;!B5Z"C(3F82579Y)+F;C)]*: 9&%2PI/+"H4S;&7
P-#*_(R E2ZQ,I8*677F%5F)/?4S5&(S4?>3@5\K3;URV)&^;18]DBJAO9_$I&&:U
P@SOV-D7;%XF-&2@YPBL#1+"LVNHG26(53>SMUZN@-EL,\088%P-$5\'?>,N&]M>D
P6,+D5CEZ.?JV=@Q3R"@Z0!'1WAIH!. FW*%^CI?-L7,7 7WJ5A0@\\<KXC<A'F6<
PF2P9<PQ(6EE4'8H_@N0P/17R0D!?8"8!I$(C]MM%GDN#*#Q/8N8L9 BU0 ::]SVL
P4C 4"\ACS<'+JT "%=1V;]509C>@HB#Z575D3QHZLL*AW^<&M&5V\PT-QDUVUV"G
P $U&HY>A#J[HP*WZ(TK[U.*4?BI<6.6"#7:QEC3CSRCZV[9\O&_U+5M$$];3^OG2
PYD3 F!\EBM7DV/>W7\4]7O$4@4-_H[O*KYE<ES2Z8!3YM(7V(LX]K"-+5CD_+EY,
P%50ZR:'S0]O(-O!<7D(=K:2L6SVTR01P!7KM8Y2T)W5 ,)W;3&0!@5VLM!<W]C13
PUTC+WHXKX?)';CT+!-3O#W8H[R4PW84L;JWGX#U:WIO6TSB)Q%4[@P"RC-FV7Q>?
P-F]<4Q+Z#I%+]YL*K0*>OH>Z?QDO'Y.9FZ**Q-P[$'F>LOSKC-O>;4?.$0N':J*B
P/3(M-2F+9]+.$OY;3R1Z14'QSTBA!0VWB;52D0JQ4^5L*9(B[T/>PVZCUTR3&K/&
P?JO#PDAX[J[3@R:J!_K-UH>O03'NKCG7IN-.P)[,7>>;$T1]FK&5(YNA/&+3\PNP
P!N9$T?Y0ZP!U<F- SK5)+H9T2+^ZQ;H8XS*E,HL>P@8_5M#>[C[@JV):N1?$$,EE
P7!,^DV"'F1P%A9XG(]];MZ>T-IP2RX83,4LJ[DB#\%F^.(0L!M&PGM&6V@VQOY0-
PSV22*9<Z^",8G%\$N9!IG%V(A>N=N6X0,YUAA^)!FN+.(Z@/1:J MB" 5M@-1HN"
P-"]#"-CJ8]LMD&.HWA1TDC"J\CMDCTFS86RW>U$?@-J,YWMM8L#N],02^#7BDD*U
PN#M/1@C)EKX"#XQI[9&VE<MZ-CIK1!1**U1XSKPR7NV%V<H]_6(()KE[H0$OFP4,
P3:W7JMT^N?1N(ZLQ=B_$#1YQ81+@?[MZ$U$R<K=18^BRJ3*ZBSH[C$Y9A":6X/1Q
PO[[4NJN(]VT-S+%'(YOBS&IOE\QE6*35K^U;,*VQTX4G&UX<"V>K*$Z[9J[I.@]<
P.<A,4ZQ_FQW;$J,(Z:.N9B,DA_(@Q2J68/PMVN'>K<N6SQBT5_O7&$>ME.EQ97?J
P *V)7Z8#:)"<"&2(7@F6O.8F\- ^3IE#9TOUH?Y6YF;5%TP:,*=M_K&*#BUZQ-!(
P%N_6V:N>#K_T+,+@EW.OT^!^69L<^,=F=I)Z1#*?&]5GR%TBUZ<EY/.4W&(QF[@N
PY):8?MVT\[W/8F_[#J%)+#&)2-V0UA__??/:[!@Q:)=#_'HA\TS#:?=72D#&R4R5
PFMP&SQG]H]^D>6F!4W[* 0%2RGWO"[D\D8="_4=.>S)ZT%R$CWT6V)<N(>'&JO;U
PE?_GL+0W5A%7&SU"-&\]R8?TSNP1N0D/!J8W6"=+G3<T%??SKR]&;]^XUSE'_#&5
PT3.0@3 5$O?@F-R:$]_XX],*P&G .TIVDF3X%?M1J:TCD-+P3:QC;[E]U0/W(/7Q
P^98R3'\!?TV+20+LLXGHOTI,^J82>EI1$8VX^(!GB&*<V-&]:D5#A)\SGZF(L HW
PW;U;U9#S;#>47<*T)LQ\X7&9ZJQ?:OOE9EE4( "=-\H$Y/\C<M^XN%8TUJ4!O% D
PG>SV:CZ3=@6Y=[FP-\X59[DT^^$'4I9*2%[B,.F=.)6V(?EAUSS45:.430UW4F7Z
P '$7#%0G%/4"&V19#/V_(OL!+'L[4LLBC4Z-2AD)?OE2 ('&%(<Q5D"_(.1MRG[Q
P%A-MTH3J("A#;[Q?_W*]<55>&' !PPG2.NF'H#88@66E&KNWI/Q=;_9<@F JF*(?
P1WS"7R./+$^Y6 :X/1869#R=$.L"XF)A4J::"VNVK(A%$:P\++&Z8G5O:Q;Z#@ZU
P$@+ECH+LE6"M5#91RS"BUUFZKOVQ^#!L#A2(:_K+R%@C'4J&@>0"CY9F5)(&7VXW
P/_J#DY76[5\\2@Z Y$(_8J:0>6#IS:=GZ8:-3BUARGA]MT"!K_=NW;L)%7;$E^5"
PUHQFM%&91:H<+6/U15? Y/+$Z?T.I['/0UKH%5PK5S9[,5>=P1M3="]R@0$88VIK
P[5<"UUZ/#:&B;?0?1E:$W<F:IZBC'D9E7?)@<&ON#S\*]T)QNN-)N_._7&?<[^94
P_^HW)PZ::;O .!^C#XU3-K17RT\\@\Z8L&&<4>U^ZW7M<W%L<FD0.UP1R&&N/].V
P?ZN"G8Q+\)K"/@!C&H-3S- >8]M%QZ;JBTBP6#7]=A#/UABNY3^7JO&A?Z56R6IN
P F5- F[>5JTAO.AJ=WP.LCF U#5/>L*&">]1H'/X^HQGP3QZ<.JM#30$&QN8O@20
P.L9,3PO#PD![3H(34[67(BL3I(E-+RX4D/R/,Z8%[CH=_A;$F./,B,$CDU1'=(:V
PPIWDP_7AQAFGCB.7[&+O+$]5,#P-!8%0KUE\K-V1DUY]!YC$($+0FD::[P6C&*)]
P:$4*:"%,*%UMS^![;6UJ@A=Y((TO"9!5E1>G#+Z*$/7+=J;ZRP5;D]4YDKL,3TXL
P!S#^:DE8KR3DVE/Z7%57FMI]0)YDFV=+0WR]2/SZ)E,-/&,+@X=8.6W_H_,W?,&.
PS028@!1L"H'N9T^#AY&M0W]B_ 3=@G9UATK_-PZ,>NM9[T/V<Q5"A0Z( G6H(%7,
P:S'X?='":2!\++ZVQ)FCIYOXM]/A3RNN:@QWG XK95H,M#7;R P-.ZV\=\2K#($Z
PV[KT[!U*8')"KK_(IM+B#7WPK4Q10<.!68T%EX9-Z5%I;I^XB)Q<GQ@\)&BX4R)"
P2E"X)Z5OJ]W+9WG'2\#>B)3,"X&RICKR:P2M2)([^)P$ST+L"I+6F1!2KK5.2&;A
P/UDX]> > ^.@/43%L$W02]P_;@ZDQ?1#+@P$6Q_BW$7HGAM_U'?"ZC#3=X]J7H6M
P6+:H:-'^9$&D;\MN8"@E*C+^@F@0ZR9'\;>L'IG?B6F;DN^JT>I.)> 0XAS7[,%2
P\L7-H-(O6%G<^X4R^TE1"'30-P,:\PI(=9>K./2\0J]\!KG7XZ(8>*.M^=Z)94'3
P=P=#'0<^GB.]K<ZL^*$!0Z $J-W;SYY7&--3P)L&%;T%=SUCQ14$U6;>U;QNG0E<
P!APV6C;DBPFA%6K<[B^AE1E!@Q_& J]'6JPL<7L?;__']E&@#F?N@\G27I5. D.[
P*906KY^V!QCU@$U((@%T"BIM$A)N&Y\96@[]*T6+UPYG3SU'L/V0L+0NH>GKJD]"
PN@:0(WXN%^4<E9$_)^DRZ.;.18U+;3^&S$?$Q  N;YKTVT$,F(8G()>:F2<P**7M
P_Y!:ED4",-V+MQ"4?/C26%]1KKF^_E#\IUG.A:GLDG8SA>^MKBRZ,_49!9\L>MA]
PQM22X)Z7_G'4E<Z")S=: RKSC7BTS].D\<T:2>41H(6]?*W=%I3DD(IAWH*%>P\K
P\?9-J:D8#XK>X.B18TNZJP"V1A@)2#J<LO8[@^ AUVR:9SC8!I4QPGBMK4S;)-\H
PCPB HA/!A>4^-^D*Q,"XTCF2LSH_/=C*-,*H2ZO#IZL$SU1+2)LCK:9Z(0WK]XM-
P^<-K9OS ")**SHXFA[U3H(_< M#]\F]3*=+I[=)NJS-I!T?(:N9-1D!8^3O!RS]<
P<Y-$$"(]%^&EZ/#GJ1/+1>=O9LT\/.($< 8[OBVUBT<$L4>]9_QR((?DZNY^-)5$
P]_O3=W2#*S/Q-+IGY*'-?P[>.B\]3&H[[3%R28W+$)?Q[%E=SU30Q'.!IRM2BK^>
PM%H!)<FQ B7M=H]KPW2T=NA\.RS4*O$9HEJA;';R7Z+=Y1B9IG761!2S*<@/SBDA
P*O.!1<IN)Y1&N8O*O^R6F/0XJ+;?.JP(W)4O%V5^9+J!A6$&F!JRO41ZBUA3RUOO
PS^5<OT RVOLPIP'VIB@- "R=O]VCJG2L;35[G\#"2==U0ZCT,I]-E#Z;3ZL@J.*X
PV0UBQ768A7NK>43_P_UK07,R5C>**8W7QGW.L -/RE$8%MY<R6<3+#V@C,HBNB7+
P_Y*1U*&!T @]'!/[,C@>![J%;,K'_G)4'JXS;^A$@>@UR/OC*_'PI"-Y?[4[SA>C
P"#L?MF_%_1'UV&F.O;P5K:_AEA3?%C12D$=8SBP8?LA SOAZFB/S1V+^J'%ALGP*
P97*,19RU[#@P7RPG/9Q CVX0KYDB_0!PG[SW ^N+F'%L3?]PC;=V Z^:RQ@GU8%'
PQV.?0F"0E!LQ5RVZN5DH=]UU!9@@X]SYSE@$C*O>POV5=1(#YVS69)1&'!+RV57 
P6[U^*%SFWS-_MS-BZ.RI394S\9-"!50I@X^F?"H-(E;V7< C$K=N>8\>H][E)FTI
PRJ()Q0T](T ECUFW1I>CS]#8M9E\M<6G65<'*<>"A<D9>-MRL (/S 4V-RD9OM 9
P5XGW'W+")&2=I!.?VMT#'BW^7/.<SV6@"5;4!^G*KHP@NQ<H\T@\_&5EE=T_'N_+
P29)SR'X=H\V87 "'RPMLY4H%J2UKR^2C0CV;V/2?0=>P\)N--ST.XXH7Y-=:Q!<W
PYSU9\2<+?]YOP(KC&,7PQ,0&ZG'=ES.8V0*<&W7U)W4S$&OJJ749%UD"P7\M12OK
PH?V5G\R83T/JF0YO(TL3LH>!PX+JQJ'T?.YWA4= R<KK"Z@AISG)A41@!+M#!OQ/
PHK3*+C $-T<P*%-2W/<ZAX %2XNKFRQN0*2W<=8XUN$G1!BA^/#A1D]UL8S3+W3R
P&0.49_+34S3IE%_9DT'KAY9)IZ<6 #"D8&5*2<J++)3&WO0"+@.M\!Z78LM<L.=X
P1+WI9+0Y).O>HX\SCDNRG=-YG-6J,/!F5&FTS5GW5H%W38$L$CV>JLD\MI;1AT7F
P<RMS[KMU.UXM, YC<#&/#]I.%1W3A/).6/)31_'WI9#A(\V@IC+^V*J=*ASYCF6 
P^XZZ7RU* %$ANPK:$CO>[&;G;FUN((I&!G708%BL)$B\P ?G'"79_81Q#"%5'APS
P76SD >2Z4P^>3@4TRP[DO0G[+ST7V2P:H*HG\8$:>?V7T)'V:@(K+0>0!_&P4=%<
P<2HVL-_L NJ%2)!@M:PO*9\]4*][T<LY)X;\G[& 62DLF-'ENJA5T[SGKZ&9PK"D
P PV16R2+IU3[D!.@IO,:*4=TL=X/B]XY&P_E4]P8OD+RO4_Y[:'MH2=$2IB?I@O/
P\#I!/OH1GMJK%\I4%\K!H??G]Q\KJ*S15M45^=2MHV*_K4\M*>93G)E3O98,U7BZ
P)P]IA5Y<V0^[C6TB_Z2X]!O: &, 7RF(],53$4S(>]R>(P7J,)[G$)3H*%%>&O6#
POZHYQJLXNHVPVL'RPU=#!O4;.[L9%__PYE4DTY=LO.L"6JWFF]6FVI&TPQ*K,R;,
PTWNH+RFHR]CLU]R0*KUROT9]R%742$4J*2L(GC=%O$#2?8S_ZE^O$XJ3/A5 ,1V%
P<Z:]U(DX#FUJ1+C1=]0$:[0&^/*=K32!\1"C"S%W[$"6Q/2$C?QV?#;JG=.7$J(N
P88#Z]X-RG**/.&'X^%SF5NG:.OU>OH^-;?+[\[\++&M%J:#CSH$E!&00AHWI)"JM
PWU('T8X[H(DGP$&APX^Z(8!M/Z%4D@*2CL7U;796.;8^Q!HP$)J*$_JA'ZB-8$.J
P4*T!QH&08(&<^1BB6@N%S#DX(LE$K,K3/8-,GHE?:(IIH#66=\@1"Z(29&J :E^;
PP4^[6(Q<?/@;QW"8"#2O+4-(UE?S3M/$!H*MC?J)N>%K8T;K:@?'&1>>(7TX#WVS
PQ?FXW!ROR8P;T2&7!OD;Z,37=Q5"*[FXH<0GQP \_7[^'X5D50H*X]JU7M ?%T*6
PJ?Q&6#?>/1XURBS+!XC7/A U-(OLEMQ*4-!9PSMH$LQE,YNF.S^_S8^*DA2P'WBQ
P1JXCQS3J\'-PS0&2IX-93W,E3V$#]05='&D=4 <M)K.-_16?TIG,BGKOE>%>T@#J
PN:SR 6\KYU?X];$;X?I@P^5/8?L:2W4<&M45#"8['A@'UG-O B!O&_,RXT2267ZY
PK9Z7I-:<]\3"W5GG,)8'ZP6'_ $)+0"[D?UZ+<AWS8J_UWCI0;W:."0'#MRW$M]X
PJY."5_$^PJHQLNZ$EQ*A +_--4%C9,A^0"LT14[8S3(YI>!_U(J*4/"X*M272AI*
PJ=8B-/ 384_==W)N=$<I[1('KG:OWT][VF%JQ_X97)M4$%\.Y-CD+4)TS(WKMS:Y
P^+*O=OV%@#C"Q](7WATHM32@O>S*U!0[T[#[!$G,614?C]Y,3O! NXU.!F8_Q'-.
P?\H@TR,:'[2\B@8O-"B%$[@OKDN_:E=OGAAP*!/^I+8ZXPZMU8E&Z\$I;%HIY=,.
P? D"XI(U61:1 ^NE;D%>$AH;.6_OTEAE0.Z%[*W+(S[S>!:3J0JQ<JH&D%8O5@9>
P*?E 2[ ;3]2NI2[K#S^^J":M)DA]EP6?R1<S91VOP*WGYTCTU%1D?H:X0X3@=D70
P4E=TWEZ+Y3[?8$H)BO!4_Y2779)Y*<Y(W'6RC^:]_4W,+M*7K^1"QG=XQ@NI%M!.
P7Y!*($C!VTUN#(%.*MP$(JW-I2MB0WEN[7HN]PU4($%*WDV$9GW3'ZD3%Q586W*^
PN0YB7)]*R'!53^#9G7A1AK"3*]SR--_,7LA*M,#N4IO<GDBEO%F-4DG;5<S[1IZ+
P9"9K;8ZFSW$1[7*E?9@1UWE N&V4RFM+XW+O?"O \O=Q3*S3M*1K$7>#>\GEW^'J
P[7*KU2L +!G>=8!9F$,@8&(62%4ASXQ80F\\VV8*L<F+I8O^CWWQ5EH*E/?W;.4&
PW8EF'0CD5GE4]!DLN/W2=_HF!7>"/CGU9C*EJ65:,?A*F<G6%U6@81*<Y#!B$<7"
PE] CBB.// 3F<8Y!F#Q-#_^7F.HH:A( &B!U:ER/8(MY?V(06R@G:F["4]G;K&]]
P :YS+R+6SGAL?V"C>5*L9C_Z,/G7/FW>%T<-E*"QF+E3E;PY1UMCB6&;/)-T\<\)
P/,B#=<;EQ;=@O!E]+:90+6[1*)[&FQVDSZ+6?OC_?'9?0ZS538B]QIC\;-RVWTYV
PL!M,_?D,$=!W%2@35(@OM$XGD WUEO^WAM+09J&A(XOR)VA+6Y^<3-H<#V=_'G"O
P8\?$TV?1!W]C5NST6@:+["/S)+Q*P#X$H<'G 21JK<:M.W]%?-K_$7P2FM:7.P&M
PG*/7M/0%P%G+3./.$CRV=%=HMEE_W='WW4/+IFM+,T_:0T[$!8=1J+H-6/'B4).Z
P6[&HP^:.#(@*FBU)_/MF-U7\+L1=?CHI*&SZ!V1[G X7!YMC[,CO@Y\29FPC,#C9
PQA_HL\TN1@'=/^=\(1?A9Z=Q3B2S_G^M!XU9_^(G(RMJ$[^Q)W&IHK3XQH0Y1=$S
P\[^[Q:E_!@_KUCA>A=OT+D;@CZ-+;MAEV@1#1Y&^JGWL#',5(B(X."?$<%O)T6;;
PZ%^$\G:O\.WG"]U)_1YIV33^%5WJ1^*#OO[_XOOE#H_3M"\MM^AHW#T'B(]-XBA\
P9?OB)&8)[F91>"UTZ,<H+>==3#3^VO$5 ;2T#CZ'=WU&&*Z%4O<R?)#QD&9;SPVW
P<$ 2//A^FX010J,>S/(A=XF9D]/5;DH/U<GCZ4&-SZX5W&$P8U=WF^B2@0SS;^J\
P;[ 'Z919>&UP*-;?,I&700/Y8D#;";WDG'C[#I(452358,3N:'?U,5\DO.V^/;MT
PK]_8L(GQ5S8\RIV8FFF"2L7$IXE#]P*L>ZH(C5R%H !H3$#DYJ">%1JL 4ZD[+0V
P=+O4&L0CP1[%F[FO7#8:Q[GQ5U_Q:R)1%!7=_'Y]"8;4N>71K>5D&40Q<@![3@/H
P"I3-V*CBT9O6.ZE-ECG4J&"+[*P(TP"#CL>XGS^,$=AK@&;Q)C&":$:7B3V-_2UA
PFYHEZ\;X2\/@PBB/@U4GX\B^B\%%VV&NGG633]]N S5:RA *E^_7ZI7A"NO84B/6
P [L.0/XR1_7Y<(U2G!!MJPGSXUXMU->%E!(A*=BD,22IW.=0$7B.^DT^,/7G1"9 
PZM1B)Y['/3YN-ST1IBE6\<FV,*8]*)PJL\G!AJ\U)R[H0TY<L-BA!-OIE-3?!'B-
P\E(T-#H;X0/9PY5EH]<V50AM-/?4D/QQY^PWO)I@>URF0\2/E&&]$:^<(W&.0.O[
PZ&E"+;YOUT 3Q*)BS$C1W8LB0.^B1X)E:'*GCSP?I*0HGVO25[-RZ_>JJDB$W0NZ
P:L2UOXJ;7O:BAY1T]L J>E<"M(F)*D-:U\19!"[@L_VARI?\!S^]3']7$3 2.":#
PHT.[E]JYSV=UD-D2L3[LEO.25ER&K2'XQCVG.Z&]V&(0$X#2\'";D3")9:Y=/$/J
P_ 2#MR>GAYGX^JP^^&7TRX.@XQ#^0#\<"[X4D6JJXE6?AG.'HZP2;2"#1ED*9M\I
PSFE/V"2%?-";H#=ZT:AE,B45E8*7"]BA? ]N*0I.DG;%_2*.SSON]<$R<H;S&A$O
P?^RPQITN>%79V1"YF$:V"6GXBR=:_,">CP=7%?UY&I?0XW!H$@.<^Y*Y^"J>961(
P43KJ'?_@+F$#E#C8_/3XKA99Z:AI.F&:2:UH;*S%^#8AF#N.:*D(ZO(OE3WVAR.O
P<JM:W.(V5C'L^&5_A_VJEK$H$YB+P-B?Z8PYY- >(,^Z^7P,]<LFIP[*)HY+Z$A%
P?4M\%36&09^M<NK_MM(=JU(AF/.!)OPP:H,NMU':H6*49,AV#]RE08^)&R&.T0O:
PDI5=.UG.E2C1.0BU+M=^OY![N#";5:'VW)#R]5KX,B+=-Y:X3$VBP6'(@^N= LRZ
P3.#?NN(4M6?S[+OA.?7:--JODI: =8S[E,N9:?F9I)VZV-,#-\>4WOK(&AV;D*Z4
P89S H?TONIAC)H3Q?($\H46O%"18=>!)!U^"CJG&B_/FH8)8Z3G\*/*Z'UZNR<I-
PNZ83->0]AC5,!GZU!S2><F%G9Z2.5(L@^\3B)//:<L+AZ,J,$UF4N?Q9 ,Y><^)+
P<?LUV^<RQF?3#H!WZUFVH&"X10A1V5?/[H&"+<=S*AH.<*B>G:U\P1:C7EVOKD?[
PM<'A+?$B$R!/-L_LQ#9C_:PT8!TLBSUG1AO6OL@$?Z\GO'J/A'R@N\TPX%Z%?V \
P$>?4H<B,&U-] ;%-@FY#3"1Q&D'(6.4HF:X:Z/[.N%4&5!I[N#" FC]9J$>=:]F.
P:>X#RI-+7V.Y:D!N0(>>BDMK53U Y)S16#<'>Y*J KDJZ9HVOX#(1@8P=SPLNA)U
PY4@#,Z>WCD/J+LSQS4F834Z.(PD6-X]OD&*\G=Z_"DN'<M#71Y+"^S.B=@P4E*8_
P,V]]4_#1@*ZUB*(-7KR8A/9;&W/[<5^8>%NS%V29PVB;"_0X5-!/1>'"W7YO-:I9
P5/%?LT_Z5OV"M+!0W>EV,7E?*/#T?EGK!A[T-XRDR\W:U2_F(@LU^/[%R#K&@JI%
P8*E#9)+I6X$9.!/C0(\LX*V#^=J.4694;=8>.\P?B:0]+K@3349%CH;W#_L!%;X;
PFY;.M\#OU&$_E)7F88>A)/:L#A%LJ54!M]M],6\:#?RH2?*[+>'S3]4@;=,D"IWC
P,HI!T];<U30:ZQ$YQM?RS'(WIF@2"0'"G:??K(J#F!(,B.4G5*8A0[;\Y\6Y,.Z4
PJDLU>;*;@$[IZ."7+X%D:O]4DAB[EF%^SO]$:K\DNB:E##XRJ%!W-.XDZ*Y%1< Y
P&(.?I*/ 5 H@V$Z &\LW!6+_(W_IPY=+9)J;GS8498ZPMQYW\&'$Z(%]\I9#0 UX
P2Y: )K\="4EWKPW"](!X9X2[W3084*SI;'B,7-OA1:- (MSZ%S[)QIENOCMJX+=Z
P>&*UU%:$='^:;GP&Q30I?AUS--S-&FH!\Y,M'R<6WMM;_;J7ML+E%4IU 0.0/CAN
P_%YV4Q(%%*0@N8U\O,1*HX.:9HV&->T@(;;T2^"J'A;R;5#:P$K>]MGYD3Q]*L"8
P)]UM:X*[#'/PK*27\Q^WH#D:;F2*Z&0>D9*O@<8@!B5@OS_&ET#1;/7Y!'K5,K3[
PTL>!G"KWG[[#"(!$%]X+*=IY;*T^;/>@QYC07OLGK"]Q9WGBI>Z+'#PL992HVO%O
PO^_A;)%TC6;_:JY[+$EFD;57U8+%QHN_FWQ=J\6P!SQ#U9*]XTLUE[J31?9NH;ET
P&FX";'OD:MF@#JAFRDPP2?@<L<A2FKRX#S-62_RJEE4\8A+LY@'GA8K]ROQWSFZ'
PO:"1R'0<)JZ6: M$?L%.),",HU27L6A^S@>9P4\_D:F,8%MZ O&<;$Z9")#\D1&1
P^"+W?MC7#I,A.<T.B]-Z<GAN:?)L/:IACCX IG)+\VM("P(Y7L$'OD4]BN@D#;3<
P#+8Q/=_?N;LQKU6M:W\</,ZP519(@J_9 H*Y?DYO%R\=N!S"20,=C&<JG]U!8MI\
PV<T]]'S_?T,2ZA>:$W/9F@]+=W2FFU6JW'6OM"3ASK+>-=:4RKP_TA9*Y?^*0H:=
PH\.6O?:8_F-IRI6?Z=PJ^J_VKP @%AXBQKX76R7P=."J5YMW)^60-Y!O(HG*)ZDQ
P:Y8!#Z0!W6!;#!\%..&Q.C, .2Z-P#-Y;:"K!T'M%5\9S."VCCJLO,0/;AJ\<3H&
P\3>0M- QQ<6-)!Y3,^'8T8'1T-6BK:HD;5D2X9K -9R$ UD&G3C"^:K(XJC%)U)K
P.D"2[?0CL7([Y>V,CB;O:M3?/96[J/#V%XE_#OW<+,QH5]L4A5Q9^IU3=E:8(T-9
P1S  )[4 D]>/8Z8%^E8([>R\DN&Z$5!8\:.PKE25]5N O!'!P]0!XK.KR/[@&ZE^
P3WNVG%8, ?!Z],RS:AU9MEK*55,!D=W0B9AY3N]*^>LID&-?15+4F5I;)\+&B2'6
P!5ARRR[A7\M05)WBSY2.#Y$@ )EH4T87_I5+O30#VD;:4;_"TI22*Q<9!V;).R^0
P@7=11G/6)Z0J)G29"S]CF"94'H8)AUR/#!@43>B&XNN[,5?]\($#_I/>+@C,.F=T
P[<#BNJ_%6JD'LA-H"<LB14D.OJ'7MO&K/OQ_\IDK_=,5TD.#43V<HT=K#'431BV0
P$F/-9KQ64M8WLO)&0Y=7AXR6F[2CXG0D/7-=Q=+<9.NX#$K6204P;,-,PM3A%X:;
PR<HC71H=#7-"I1(? "($DSC,V;5+V+\@363YZ\<]GR-E68D.NCF6B0S&:L_P0FLW
P\G=SSA8,#$P*FTT9,\%_DR25&B6 2^6@!'#P,=)U!HWQ<>@7/VW /.E"I?N+*NE(
PD1(0V^]_7[?@+%W8]UK]U'?3TBC:C,,35T!HJ\^7?P(;.9VWPA9P#[\%]MG<:TP\
P5'$OR-V5Q0>+'K];_OQG>'^*45WBYHQ?E?6O7+PAQNV!1"M/]7FL1DT<QD7[0$HS
P(=/%&V2O(#.2J)OVFYF7SMR%CNG6(5,-GNTAL2A@[=0;9!?]4;+08F@,RW/KU4L&
PN"?0,W.R27ZY D[?NNPT-"::*9TTO%WP++8&"WB^RO:!QY85B,(KI$GG-\R*LS1,
PE:^RGU\;!'?A;>!T%ABZJ3PR.13FO-3 RSXE+*;RO&M"SM:KA2QT\9'@8NEPIVXO
PX]-^9TPR0C'AK?=W!@E;F42]']# 5#J#V2Q<HKIW-,US<2%]9<7[6=/. LD]F-<^
PJ[WR)V7QO:8/SH)0$CPPJ@\1PY=O@+L^$E+>U,<A@2DO=O(:NVCYUGH 0$%?\,FR
P6-!,.K']G"8XP(VMP&MWV-<U29]2_FOC__>&..42JVSNGDZCN+C0^VL//:D+]I>>
PL&*ZINS(%PV7APBN,+!W3V]T;007UX6X0Z9=@@,L6YOU7/M3[IGR7M.H),]3]WJG
P("+CEMBI&;+0"%_]VS#?UTE\U;9STF4W:)WYIJ5P!;32'3F)[/:7:.=:8^ERTE@"
P\8](R%'N(9H-1Q$$0*'"^/2,]A=,3_QMN"Q!W6V)5(5V61"DR^EQB% 'E&S:+=;:
PXF^1O7@V'6;5,O]S&&]R\-XS,%AY6%FE"K5RK,JCUGT]BM* +[I]5V"B O9(+P_ 
PCA5]9.B.="I-J-H')MA],W\;+RV)>>;VC*I3YA]+#/ *P@^].NBPRWC*[C&$9K\'
P\O7-JU;#DCC%7RKQKP8K?B,=C"=<D*.Y2^7$D)(DI&;Z4$J&LOKWLQ-=3#;W]L)?
PF$PUM>?DIHFIT-+CGXL)@88TGJS#]6T_%P8[-8M5*H&&W*!^<O_P(.&]8]GWP,E&
P59(31:A;94UXK%4V&!WSH?R5TB%V)HL9ZNAEB4QDR$#%: 2>? ]R7MYGBFI(27!@
PR2&VOL@OL'-!HB[5JT)J20-7U+QM:O7T9YM;9XH;")RS6'TD.N:IIKXSOZ_F[9@>
P>^A]#&NDQK!V6IH')NB0QPWW%OI.UO:()G;H1M;-[/NOB> )KW'95+4ARE<DC;UP
P$T3Y:4PL+\;6CV2'V'J>#\5QK43\.S(M'I0^6!< GM/!0,< )'H^K&DS57&"\20Y
P^B\A%I8)#41>$:'-VHQ-PWWER_3=S@/;YF#94'T&<P^XI1 >UP*[8N!N(.IGSC72
P(FRQO;(V)(L/(4&'B7&L+WJ&ZVD>UGI8?D$6#!0JWF[MNIYO27&!/#&,YE>3V2[*
P\;9*-(^UCO(!^4XM;<. V'O,"SP/WW8'Q]Q"55!ONNT I+U<6-CHZHCY/F] 5DB 
PRN-*S06F:Z3_S)6L(M;"\?G\7%>8_NR# S9.JK6F-E0Q@T1XF!E'N7B%EAB\GO7:
P-@AI0';8^V&7.I\:?^?J'10NK.!BXG_@#68,"\BK3R#UC:7UIIE@1]"$2917]Q /
P$&;J.1_](M^&R=1)/N(7!,UH+A-L*I_(\2.0ZD5*\ (0"ED);9Z0T:R2L#;RIP39
P+VD,\OJEY/SZQS>^X=UTXI&>UO)]3@1._W U5RP8]6DP/3[-Y//C!Z QC@X66WCN
PAMJZNM^TV:L]<JO=<L#.C*8=RGP3DEA#K\.>U\%Y6!]@# -'WP('#?-W>TIZM;2W
P:/:3N=:$MMLC0"1P'L=]+7FSID\,6(%\KH_DP(AAN$M2J0_ 5^Y$VA#T$L;V.UU-
P6*0.ZJ^-DQ&57ZL75 ,*>ZGI90H"D2,W=3;RNSOBZ&0K*VZ5AJ4#@0/R"F.ST=3'
P^V%5]XH1<:YL)L4!)8@38*\QQ2BJC^K:]6_H:2[9/ RV KM5+1UK?0/%^F^^W( W
P81GK;N:#K0AK"[?.%$&=:SKL!&^!7T62D<B4_*P^P4O+[-.I=X2%08< +\)TH@5&
PZDA)L^OP#K$AFXQJVK2[ ! "H=Z[U=11;K^%S^81(5 68JM%:%C&V5UJN%I%/VCY
P0:FLN?>.!-V(*2 1-'YC%,)-14#*DI:,)A]AL#K6U$?>K_YPJPGRE);Q-*#<;=/6
P+KT7567,P&<[-@HG"T/Z6^Q8]*34 4+6VW%\$N^MAI/^425A^'G+@#T%..)G%@'D
PBALH$/Q.8EB 1:[#HDYS0,*)K4NOMD"H\$649]$ V^5\GZP>P:^R<4YA:F,._ [P
PSJ-;=_&E[O%S5JR<@XC"HK_2^N.Y/2ZP]2<CX&CL1Y0*BAC^;T=,R0IQ494I&Q1G
P?Q4QRB,#20#^(S,-Q+I.X_JI^V[ZX$"N(9)>(5Z7R4[85>!J90%%X2C=,)ZO90:Q
P6O$X?":4^F#UM;*-&AEMNG^RR YGX?%^(E \>G)"^&@<=;,7EX$5+-6A8H8)16L&
PAMQ0#L $092F>U&!UQL'P)N!>S[(W?B_C,GYFU:D=K*3OCOGIK6KKHIUW=C+GM'_
PK.,M#+,1 M)/.=\D5\_-#+O%(_BDZ:P&_&_ED0P6O'/:0HO63S?2UUQ/+ 21Y=I[
P,+6A#/G[2I'T\PF3U_<'E.^^I/D#,VN(\DT@*V)*NZ"YPVS[0/,H69_E;?-1ME]-
P#.M3@('42*,IID/B:%L\J(>78 @GE:R> -U%;>^5+'DFJGE\;>B\X?.VU#(7R(*N
PQ8ZR8PC;#5SW,))4 \1/=OGMK5^#<NF8X7O:WR*DI3<9C.L/3_TQ0:"J0GHAX(;H
PO8[8>>Z=^6(.,S#BW:PC5.WB^A(Z^$?W3,E<G3?^@:;-9#U6T?3#"M$"">ISK\_Z
P]7RE,)3\BZG-Q)A1##V#)( +DW!:JW&=7LG-Z";K.>_GM;3:D[3-.\+N)&_CN__F
PE^=  N(76$GWN0?'W_KYA#"-R?XA1U@EKY"C4G8"^LN\N6XNW>>QDMJIWY#2O!7<
P.<)F6_95\C"D&KK2N;-LY<9)'U4%P%3VYYQTX$V@/XFQZ75(EI/B1,H>TB]]GZ-8
P[AB=E (+!<@"E>>\63/W0PWD#\<_%L[(7EV$??<3 G8_Z(">/.86W;49^DA@Y%QZ
POWXEG()MY20T4[ KK0\7-WQ2*F4+WX.7B+H$!0G,5L.N2>PFJ-ILI+DV@Q7DP.@C
P57;FOR^@K+,DRRQ19SQOUL_WVPV)1V4<'L0S^@U: &<*IE44[\F@*_@EWXK+>I52
PE8+1Y-0_G*85!'-D,LI]UC&N/&;=.&G\Y<+8+?@GYUSH[L2T'=?;N_%,B'H%0P@!
P&!ZUQ:A%Z>?RL*>"IV_/$!B@U'SZLU 'HW!$W0BC[B@\9"P(\E_F]",%V)7ZU18$
P=*C-S3Y&G3U%UIJ*T-Y3"_G)DBEUA?RS6$=A?>T427\*10ZN=2^"7L6(0J>>BO8C
P;MS18C.;Y5DR)[)&^T-N"0GPGZT4BSDGP$B(X7@37&EY\)H+#.MN7?[0HK?$*[L6
P&O.K_%&))?*57)N$J!WX0B@T+4&0:;&ZNC*YP;YWM5AP$?#Y HC=_:W\42?>YNCB
P]&'8N2NU.9PH$(F:=]S-:3(1D56!_*_8W4%%6*OP);?A8D^HLMRQ=H%LV/00\:>,
P.\F!F6D..$2S6O,-\*>N2C5XW9=PQ6'][H-8/$YZ2?]#._CA)3K\'Y(LUYSQ10G=
P+ROLML%8 =Y&)X0QR8GAF=E^4@_[1;?!G0D1>,7+T7\GS'4XK7/,(B#[$C(DIG-H
P@@ JO\..=<7GC&G3--M-MWK,;#/<9URGR1WRKN+OM1^D,P'.=IYDD[-]/YH+OV\$
PBKI1R@ZTA**'6W:-:6._.2%(J_G1&+,[#W8P\U;/R-4K6']9[D?X%BG4!IH7"U5G
P*/H:IZE&0URA:$@INK9K<?;9;5UFJ?1]K^19,%3';/C8_H$S,G?:[1 #E<?N]]TC
P]+9> ":#1F@B_Y!QFPOMTC0;>R"16<$3@ZM4>LKOMR.M8TD6S?LE6A]V#@Q";.>Z
PG.JG0+?]<4(F9X*@%[_OT?+!X-D%3>UV3]S!6[F583P(QB <TDWX-H#!9KM?9]J$
P-_6]-'LJG:"Q%62)@7F^%]K%=L;G=KH1GB./_"RU=O2Q/TW?E6*D?E!P[';@,Z1K
P">%HZ"Y*SBDH PA$)08_#TY9" 6?XES+6/4O*"#$;Z1*\T$KLT='/WWP>:=LNS=/
P[2*S/ 787/\V]09M^H+P>D#S#T]S6I@=:?U)5Z^>QPMNJQ#,=B%HBJ$D<+]\'0@8
P)P>(4GE^K795[!/,>F=3<6X*DV<7KPH[6[>#4=F0-HCSRU32G*$,.)8-38UU_3 P
P($ UZTVD8?\K R+,-00G!F)3OKU/3L"FR7*Z+C9=UJEJ3J1D*FFQ2\[1I,FL"1_9
P<[=QD>B!C\8?)IM)27:Q9GJ0/^GTT9Y3X_Z!YF*>E?4EG# 8BWE&8,.T.D=-&H D
PJM[4/$ ;'D6GN>''?4-LA[\"$E=KJO]S:$RE<L7;QY[=AQ@J :>8HVC*Y%G?AB4J
PH/#8HX '$EGTL<7.YW1?Q5 @L_RYJ4%I7V5(BM"1%938.O#YR TAC5]>MKJT6%JL
P$W.&O.DJ>>5=0"QV8]FV8V6+5*/2V(S:1Y8VKH!596DI0T),#8LK>@J)/UKN+M:5
P3E1[Q>Q 9AG,_F(HC]"4YRLKO7B@<QR76@#PKJBR/<X9-BQ]-&2OMQS'$SPBMX8Y
P3_D"BX$XNZ<\^K&E$G*E-?AT(E\_R)W=J4Q4TG@)J,)MU]$U WJG,$1)\[Q'@=5A
PEQTWEN ;OLFT+'@O[&#JR[.GDU#Y,MP;U3I5X.N]08W+)=S!K4V?.$2TC&[7O[7D
P?OH!VFZLE5>#J-Y:-NNP4_%^ZZKTBD,([I%(:Y+GTB(Y]#*$*N3H7>X$_X7-$._5
P?+ZG-0"QE]4?B U7*9S2##= 9^P=_WH@_LDD#Y)- %?"+7/(/TMPP,[,ZJ^SZH,(
P'[-M>K;\*"_E1LR4@#RW][TX%@Z@\T.]N5>XB.?[1(!HUJ2)R$G DR#<BMQFSQ%;
PW%KK>$+#MJ'3JQ!YBP5/DF@!"M0COCENQ=B1IP1PA\EBDUULS(U: [BE9IPC!I;K
P_KQ#8V:]E"_9L[SWDG.WNG79.>@B3^HQEN>VB:UA]0+K.)?SFA%U<8L-O,(DJ!F:
P/KJ84_PW=9TYWXF[H!4N9N*-7UL0P^(%LH.\J2#T'['YK%Q,?8\.X[:8\2C492<>
P<;U* ')402-IT+DXZ:%FZ2*MG5 V5'&QC77TO''3)M<S3,9!3CU[O8MY:IVT;DAC
P;R:I.-KM3[@G<H!J_PS5/?'323W#5(\BW05B!&B6_WH KN<@N9!>D.4S* HFDBO\
PJ$7-PA?.]J6&:^$EI,-5Q[KS\Q!N+H@X+.C5>%I(78"*7QXV1O#:1O]@5?GB"))(
P"W-QCVIR^3LZJMTOHL9/ W,D=:@6;N)CV+0I&0\=[UHQ<;0KO!U6'?+O3,I*7I>3
P=<.4:^TP5^5T>_MM>M9\G.U^)AOR))U/Z!-0EM[)DGY(GZ07[0Y\Z3B4/-EV970Q
P';'2>L=(FSS<=/F'>ML$'#) T\9X=/XI^<2 \P=7@TV>=TT2:!QHWW(Q"X5(7O"<
PHC95J.A6-.7H62"N6GI9I!;G[3MAC B1OI9Z]+F7(AC>5+A'54+CX=9XSM%BR"E8
PFO? @=*5&=2KW%25VKA4.N'.&\E"\PS]:EN!2E0,GH[TETZWT7Y4ZK<3S8"'J;"(
P"O[E\:F7$;Y!(')S(RU_,("QOORA]9G"MA05S#V(V<$X-[^ZD_P5[P>%QX[E&W5*
P6TH)3,9 ^72G_0\-VC.T^W<?D647E(AH6WML^>M*=&+J=;0\F\,)5V,E6WZ,_E@_
PZ0S,W$ !WIPX*19V-S/>L><G8^&.-54I0K=7B /%[B-J*3*KG_+T@HN[/F 'M3-<
P]G(;$-F^5,;$K-!@TMC@ E.]O<J(/8GTK'G6-BX;8Z?CW;S;BP\^C^0P>2]<_)??
P<VA8?+%>(&K?;=MR9627&]J\9OA]$[!2JI$K."C)JBBE.H=R6:J *29%);'1>; O
PY5)?21:RJYEZ!9B-RP9*P8NDP#**6/C9%4^),AUEHA>Q+UJWF5FEK$]_:G]$F5GB
PB&#?DDKFXU&(Y^SVN)FG4Q.JWXDDJF=*SUP$5H7H])K)1D;R7YWWN51OG-#PN"C5
PRCXX C*:,SJZ,SC#!O:D[-A8\3B8!QOE>QT;^-@%D\0U@_FX>D:9='S(T8:;IEXU
P*IQ_$1<EZBULO<A#.=6R)XPN32MQG^8/>> FCS7NXSER 6I."A/,&L[%*)#4#=1F
P1989PB+ZC77JXC6 3U*,"ZROT5V4.*7LT=F/=@*LPMFW2/,4!QBM&;T^#N>!RP9%
PT]05:?V7T[F [>FO6)72*+W) FV:LA28:E=?-'OMR/?_P8B!N\]HE/8.1V]3I&K=
PW);;8G?$K94QJ2$<7R:L;<&WY>Y1FR&H%L/J&YXOWQ0M=KO'7<9^2GQUD4H1'D[R
P .,%LX+_-H4,VRRC=$6W-H.$#0/8@J4&CDEQGWKYCD5EYJMAG#,3%.1N&]$&]^%S
PO%J],96WC.@5:L( 05"2P*W1_>"STV044=23M)5@/ZOZ0UT7XUGM<O1Z%'%?;"[W
PA0P$2!F2)_AO8A(GA-F3U5L*O'G(FH<#BUS?2RNP1L]./OED&J>,'4Z""*-O .",
PY0IR2GH8EI]I C"+BAZN7C*D7_\'6Z&F AL3JE>G?G=2$TVO"OB9O_T&RU1A\1L>
PU+?WS0XQ!VM&!3&.7NV75SD23D?@V%GHJ@SE7$0V(SIH+RH&CT3&00N_53OC(7CW
P;T2%D84 3&)<D4@RQ5-61!H+S#A&16:>)S28,/!2[;[(V@4XZ:;)9*@9G4$1SNJI
P[HOM#8BJB0]S4ZGLM&13P<PHPL^EH^LB+AEI/XEFHX]0N/-I%T=_Z=\WY//FU\PK
P$8958OE!OM .R(AE4-HQFL@.9U';ZEF7;\W@3J#:X"?Q-8@)\00WRD*E=IR[*WME
P(Q/96$?Z#T-GO;#'9B^/*):2WC9^?W?YVY@<H)?AS0MLH/-VT\NQR/Z)&L^JOL-Z
P OU,K=ZDX@K.?WT^U\?<KU5@S1.6V@_O(<6VR)A+S;S@\O<Z/@L')^.+/FQIL+;[
P$M'D?Y7HWHL,P4P@U_B14G= R-71=4@QUZWU>F"EV\F#W9>&J^S#UDPS/!V/0,RD
P#4K-RA$7SP2KP@0G7> UX*2-BH2.JG^Z([+X0,^-0^F5]GP_8HS/Q_F]5SB<FG);
P6>[[=]J,SYJ\-6F=]3"1&_9?T9YB:ZT]L N(#L@*T$DY1G\078B2[U[C>3# 9!DH
PSZQEO:IKHMX XZLO(V_8"A,\TKB/ QN(L1 ^*H3:NAV/W3.XQ/9*REK'% FXA**D
PU3"&;S(F5CX$R_[RIQ*Z/5($X1-M_^-N#H+>3GWX'&^?N"V*B^;90>A3,(TM9*O"
PG(TL5+=9::6X\E"/X1]]&A M5C]K/"TRCESA<JWCGU7CS8L/GPFB91,UU<WE2[=4
P T1&1J"&^AY@>528GC ;E0D-'4;#U*N)\67NPEH;N2J<M;PDT&AXN/(N4K6C0I6?
PMKHJ+3VG#2EQ6JT#D[YG60N$R4-1WD"35%>"KZ:KM,_R52IB*OS)\&U?'&7LEZR=
P'VK[V_V2#KJ-5)!3$4%S12PR7L+LO/ @VP-> TZ]ULRYO/ZG;H?"VY,/.B"^-JS\
P4VG7U78%<>ZHG*( 'F3%:;^)P37?H=JAN 0:AJB0DL.U!($BHK4%H'8$71695Z^>
PP:IT+ U2+_L[U:EO&-;%&_54T]'48?).KUV^ER09\ICZ/T<N+$R_.WWA!N!)F D1
P308\(KLV]\']EL'NLY;GEYD+>KOT$MWZ=82JA:,Z$%GN*'TFAQ F$%AS12$FMI&/
P";>FZ@61&##P?4C@%&"1;Q @K1 JC%C.MT@F]E2#BH_SB#[V\QQ PX8,^,$ \*9$
P';9+Q.D3W!9MHFVXODA2.H,X],GQXJ95C>NEX3^-T!XTI])M;:56 >T1,0;'"7WU
PX+A-L=KO?/MX:"?_>;?53Q$;=FBR4W 9:^B+UT^WE_J8>O:WD?V!X?GDL5T,,7U 
P@&HD/0!UL'L=E7 S&D#RP6_*2S9?V<_%.78)CWVR59_AM6I3>(E:-:=XK$XU#Z\Y
PM+']>\';#KI_9YRQDZ%+A(M!_?G1N&!\/6DBC[2.E]) 3L:]_.N?%3PEG"O3[K[8
P<8 ]$;E-P1ZB:1?4\?&Q/;;>(V&/['7+9AR_MQCA<%']^$CA":[KELJ/ 9Y>!E9F
PC@[$@/8MW!,3-YX818$.2B4;BWUEN_N[B!%^FRQT(XNRHA[CZPQ)[X(##+BLRYPV
P;18;3]MKPT!$"2UD*N;-M:PW/X/IF.,6!^36\-&!WHPH^_BH@!2Y^=2/-7.9HK6 
PHIM1!CPH;PVU2)[M,(N;WF,@^#AOMI*&P4RBUJK%>B226B?)D F3#ML@VU.^:HKK
P:J+Z(R&*?J)A>; GP[NY)S>WN5A;V";Y@9%3E"T]\'Y+S$PV5/=A)YPV2[0S3R:'
P@$J+9PER0@DGS6@CFEF<]ZD&6?F*,C!Q\. ]" &ESP<B ;M/$MIS-5B%V]5B?Y5Y
PIG49T,%=^ES[!YB(%:-AA]O>)8R/MOD"YCR311.9/./"]?&^[]#;%1I%8<_Z/7?/
PF&P,J:13<4THE"L)CA>.>O.29ZNK,A?OR-?QM,*+V.V7\$*)':>'H@:,#<-8XOM8
PYBC=\>_A#&1^7WL;VD4C#G%#ZHB661Z[<\_8*IL?@]2L%,5'?;*B<>ZU460T!4+Y
PQ*BF83W25T;4:LKA&#(:<,B+=ZA 1KZW(S%TWX PP8,W4H(K!?NGG&L!-'T5Z3GN
P W<)JP:@<@>%^[?VBC8EXL8_6GQK_1&<NLO(O'955IK=.1%J8</'77+BLKS-E9=@
P!\J=5 )W),K%?GE%(_J192F3$Q>H4:M!?V/LII'^)/%2:6Q!.HU(<RAW.3/5.Y/!
PYI-BP_8^G<(Z2&C38"%C@>Z$.4)T=9N',+CRZ\LJ  .R^M'0VYK-+VNUB5$GD<N'
P%@[F4+>)*K< ^MO=;/*;[JBPSGFJN$G]!LPXXJHU"N8%[(_W7<P06K8D\GNQPA]4
P$M\?W$N#)>'ZTO&U'0EC(@D(XE[<+=##MKK7@'6%[.1]I*N<M#PIM(3TBWJV1!C=
PNW?K9+(V%*'*:(^84#>>=5)!E& 8)Q@X9:=+^F/0P2JI]2DY$0[/+$T1I#NC2J3I
PA2PRH??HGU!L=*(2UWN 51S/4OATZ$3OZ=VVY\:/A241P<;O##? )K.N*?2&6KWM
P<8L2Z?I.;5PVWLUEL6H*$<O&XE9PQ"-TGU3'&FI1YC5L!]DF/89-Z<^Q)@NA6521
P]\8RFJ=D#L.528F5@IN&J2348\'#QV*M68;&91O;[[3^% RCI^<2 /X*Y!L-5Y;F
P'(OW=M);VN4SN[&!S:%(KSI)%<3FYXPV^BS?DNS;>%'1C2VO4V/@7\- 1T4?]<:S
P-U3R*;^H'Y,);18YD8,46+,XGV8';S$++-HG<@;C?61[#U-?)K)]3&B:23 @YM>8
P7J4JPZ7?'ZIMYT)$:J4&/.?P E[D"64+8=@DNQOF.[$60ZDU<Y-N0(M<QU]V]]X<
P]2 =@4O;X70_/ JK(1H=#N,B%>#4E/YSQM#+IF3J+I"=$9)WZ&[US3WL H(;:J3J
PC3 IZ&&S!^'4,Q=C6I0A?3-6(1;HDP4:F[]A)$8%=7*H&O^$X'1AT?WZ4OY 82E=
PJ@N;>DM^;="O#1\N0XC(?7M_DN49?B\3^ <CRD(MOC81("NP235S@NLN_L*."/<X
PNYP#2+<*W?SJ32XQN$&2^=73!?R6([42>O^EM$BTD5TDAL;K)7=*_N*Q6^9%<>3H
P.9!EUZ0:C,<5,.4+6&T+2Q[(*BH=[C(A&.D"^<>#0,V2,4=+HG&-8.(SZ)"^O8>:
P'L %]C6TL3 1S?^_JY;V,LN&?8#,1QN>IVS5;4!'UD!NCA]BZ)=E])4=(X>C#'JQ
P0=!BMX592 =>'DP(CX-@L>;#&%E56+N9A \HO#%64B<@YR8WT]WN>2G3I38"+Z\+
PS>UA1VL7.$>\[<&]]53 XPT<HR9,9%.J;)XR8+1X";<?8OY360:E:]'2@*AFDQP>
PU7UL;_M>*H4 ^,-R@-[ADPU_&IW5-$'PXR.1+=LW-G9\*0>Y8P_26\BG8MP"VRYT
P5(J.H96:SM\3=99I(E5U-$.<#L"9G3?/ P959]#-. 6%MJD@+;%1M;3\]N[LP-5/
P)%E$L=YVJEQCR9N"E+MV(\UD>I:?2HV2V:]0/T2XN^6RS]'#Y?AOJ51A ::+[0-U
P'"@HTQ$-&< B*0G'8Y.F1DB7.!S.=B%IR!+!P+^$P7ZP;X.>UZ2,H79.GK)=I.H_
PB>$FUDQ048 E>>SSD'-1P14^10 "5W(*%U> -W7NXJX-?PP\T'?F:<:7PS# S);6
P:0$3<8<-R$_B_PN$@9GUGPOPCHA1^0\I8P"48(6G@<;@N%Y<$H;:2]K&&)51C,0>
PVLT:D;I-"C)8*BFUK=!X,]9:-DNO%\BAB!/"DH"#6%?0U"+@V0-QPL^+V;RN$J&"
P]8O@5?(82T=:Q7:$Q.TVY5=SRM43,3&> 7G$N,^0ZRY2#G$%XTU;LB:F7J^+0,TC
P-HY1P+ P14<O$P#;,WQ?! RNV:8.>#D7VE?! %SP@!/@=84'; Y7'LQ[9=8/Y%^B
PDQ/K5UI$9!",R^78'XZMSB_**#TBOC8J[#SG4A! ,/@))$@EN;'W.BA+]Z#)?C45
P;%)U*6HG.OZ3HMUQ)6//?#3UJ'Q5+_>\].O\"H]C86D 7$ <OJ /UN@1-)A.R-P0
PUV2&AG3>W[8AC%CD;M![HU% SJA03[>%E-GDXF-X&AC;D/0?WJY+0.<XO+P*;6\Y
P!SMMF0,S#/^@3OLXL$82TS$/!QE5X7 99Z3]*!$I4'26MZ75?9"W+D_5^#%[2H*D
P:H9K35[]2,^X).#KG_9>,'\Y:(?[T_M>A(U :Y!-(6@K#J%#JFO/\FP4JVI%F))5
PW' ,S=1&PYN)+,#LSB>>V,]<KE&O)X:H/#;UOK QVLEWV5187BTM@WP+X3MK/K9O
PCZL<7VA2UI-%:!\<^'I"&KZ.I?QF)34KA1. E$<82LA;\)%G(;J3COZ?M$+W.1GW
P$PO60B^W&&N>$"AVBMQ?EJ@PZ7TV;HN8=(4]:R6FIZ_5H#>#B;Q"D=J/-8"L*X@W
P93I4]ZPGFX1SHX%-_&$?6<1@E'OZ&X>[GJU,+L3FE0IB97%Z0*N,O^WP;=OITY(9
PA/ %C U9A?.S7K#+3>V2@2\$+0WI;=+7;*+IB_WFYBIOOLOE8+XY+!,;_I; MG4P
P^$&#A<K3[*(@3/- R@+SROG=",7)6H*INN>ZU:>-D+_)/+.)EC;Y;^E9[,U-%!(O
P+&E54,_?>KCF^EL#;U'M^J14" #:FNH?#"O])0E?$LNZHM;=0G;]N)72SSL&Z%A.
PY!QZ7F5?^_%D.?KAN3%HI<XZ%P#3(D*]=Q+D/JADRVIU^\B=!V826@%;1K?)<,3D
P;WW)K;?D62243E4ML67$?MQ#X?*<F#"IL.C'L=%J704.2QGB\SN8M0+9-R%/ET8 
P'M2K9=;U_J6 JC'XR71OV[MS=&R\Y+)"5/=[T(7<6?QHF&8^8I;]H\=T^C+:N)%<
P"6H9H0T+&>^'1%,NX:W2Z6G\= BV"@HC_%2X=D) Q&5&E3EOU>5-!V!A9E_.U?.6
PW<TW]OS6@#6_,2GVV_DR=;?=KXVPR4B]L9M"ZZI7F$P5W4"N#));]&<Y&QU;:"\]
P7ZZR*$I-E=AB:=?-O>P*MVD(YL?OE9AO/+BVN5 A]K'JM;&1H$O)0FDA$T;$XI[ 
PC>;C)';3&3>9!06IM<L)5CB;&LLG^H8F>^<@%"N/-?6]?\#C+2E"N!.I\7FHEW^%
PFF3A6=)H54*RQ#[(GQDP'6[HPQ%B=CW_D9[&Q8A1O(6$N>4G_2CQ<D-GBD9=.'BQ
P;QYJ^O6P&W!@:42*]*;X,/3%KL_"%%M&]7PQ2[C7T_@  GHEC5.LE*O#C*ZYNIPH
P!4LPJQ*[5M2]9=$7E)H-H$2A^.TEJAS'AOJ3_/B].$82SKI7YHZ9F8Z*O.!%Y_37
P-VP5ANN=. L+JQ7CEDE(T%2$OT!XT<Y]9T/W:UY'N421AEZ5K_.I6AJ38$E(M=UV
P.MV^7V( /Z[P^*>_2R,Z9( V2\")Y28O@GPJ6];^'B2+'>TJ"D26\$2:W7$B?9S!
P^>:SZUJ>)+%][",]NJJT09R^NI-K6X8 &'1H+38NKQN/:_5J+(=W"YPP'%^]PLL]
P[_];<9RRKY&+90=;0[5T2_&8="MI?Q'O LPI,,:V7J+#:E[ Z9BRPF5K:V.8K$B.
PJL71E6+3:%UZ[4T9:E&&+ZJ)0:;KM+*,(MHT3&MBBZ7H-Q"0"SJ9; 6PC8 \)VB6
PZ36C*@SUANE_R2V>-)C,+ <6!GB;'%>('W52Z-W=RS!56L0Z7*Y.]3?*G@'.$:_P
PU2;AO/EA4H550STS%0A(@1L8X=JG\&C4G+P7%%\F+FV1@"K^(4^+ *% T6+4,E;4
P0:+Z15 D(+G.+FUN*TL3P76,F>&+\42+TN1"!'M2T;6<0!ZW\,HP])[&E(<\^(N3
P-4.7BB#B\6(C)@/869H/8/# 9< YU#]F< L2%3[=R8I.:-?KFJ_?ADY\I.+^,#J*
PJWE(\&C4T)*QF=;[JUOR8*2]02P*Z^3S/4\H4@T8$ :FY=.D>+RI_:8SW2"94Y_6
P/AU?O1%*+BCQ.,[*!;^NM'',%E2.9>)^>N]!^(N 0%Y!ZT <$H$[=UQ^(I$UX-&'
P,P&\UCH\]78R #U&=5,QFF/793CY73B*%1DDH2@GWNFX#F=M*<^EB\'>-%\'>@95
P8P?]6!_?(5>D=$JPV!A+_:QF.IPKY@\\\^,AKQ?P0X92AV]:9]V.)5ES*![+(XYV
PT\2"< LQ;^\O#C6]G@TS53U ZG*<3JGDGZ[B+EGN'\?^.TB$X/EB]S6N&5D9Y:YT
P-KAU.LJZ)D[AV9=-D.<*2;RM7N\]JW-R(PW1W<ONX'/#J3I(CZ(NM50XRXT1TAV,
PAN(&&8X-*U*Q"!2T&&;2,WGLI!G,H/4<@Q<+>M?TWRH3\&=SH 1CK?D',,5\_]UU
PF0M,3"]+9KG;6TI%+W%FN.2G,;/1NF&9Q*[T2 +5G/+1,RHU8A,MQ!;Y$=$_Z@.B
P%L#/:=305NM%T0)/.K4@953RN9#O@A*W'^QIU(:&ZY@)*)(5KB $CSTH:$M8-H\T
PCF>CF?I$D80EMZ*)AS'YN:H5Z@F98GWP#@Y+XBZ(7<7++V;Q)P0(/&JV$2OAA((;
P,37- =(Z7G2 =]@O+Z1-AE@6E<>HUVQ/J"<V6E\%I+U<07TWJN6ZX4WA/=0JFQAF
P;?>#\4AI-KN\9%>!='PQ"0TBGJF)L (YS'#VEDIS)FP/R-=@/9TEPU 6,ZS-ST8Z
PFAJL3_&ZO*@T!W1A<4<;U_L4,[#NIU LS1ZF4>%!@L]MO&8+!E-6^7NAQ 'Z399@
PH:KF4)B_!\AWO:YJ<EKH>,%P38JT,.402JQ^<6!63"[TNR.VSA82Z?X0LL3Z1\UT
PE8,1Y"O^HJIP6*T0"Y2HMLOOJ$Q4PX;)E+B2$O JU*]+K473Q#LU#3L.QMG9Q49:
P]9?3HM!Y/WELKUB^TG$)4X/1]D! 0-#W=8K9]8Y0C1-TB>O=#+<8<5??T?Z37]_"
PPG*W-?^1_KBY*5;SW:-.99)W6#RE:SK[5,_]]XA2/0Q[B[X0A^9O?TBD-?!1&53=
P7&L._[5%D6]"6H)XPZ:BMNX2+E&F>-*FYB@U>)>CB_>2!+S8TM!PLD[AEA^8%GY,
P99^8??H]T-:GM4[<;?$5]]D9OMX%ALA^2 6Y'F/H)A5C37IRU_:-0D,%F)NC#:6?
P]QD]HZ!B;+6:0%G^#N?$Y@ZK$1&E[RK<]==4\H/ S49T&F51^;3KU_#;XX0*[ OX
P%OH]A4K^KS[V2G"V%!R[$NH4L!^7F_&S!KG)]>T7;:D+'F:2:JTG."0\N[Y?>#D;
P!%'GPC'%.,<VA)\%[:#\Y2Q)F//##<FU\BG4P%2[92$E.E?YQG^LI^C&4EK2W:I$
P)(9DK#Y,\T%JFKEK_UK0Y5=I-$/,)>51,][JP?VY+;JY\BNQZ]W*_+#$H3QAAV>X
PAU\,OF$@$+ZOJ=S>Y(8(EDQ=P5L-[+>-.7='=!^!EJ?(1%@W2'24#5!FQ"B$M+%6
P!L'EXM1,6!?IJF\2^>B2?WT_?H/ON*-65% 7WF6P X2+7+.UC=1=^ N"D8!1^Y$W
PP4#.E2FJB$L<R)E7-'K1;\+4YORS#>:OS/(H+EK"'N7[Y!DZ/5/I%[<2!A@4V'CB
PJ!Z_-<N)UI!&\S<N;82Z TS=(5F'L:@A-Y2<D9HJ!^^[>;BTZ6!_M);^3]SB$1]*
PT.4];1%/LH@<Y>0H@)I#PE\S%*UCG (X[[C&T2I8,UBS1-"//M2DPG6"?)R,96 &
P(TH_[LE57)+"02M\.&FTOIDE2;R40,@8!PX]04O;F47[L?'7IS0*UN\@&6YFKV/7
PMV>SM_F!N 18=ZQA?RSBJ=K'6ZUJ_>9]IZ-*^HP2=</9/H"<VBN@2WH@!&H(.F]+
P5BULQ^93]B)YX(JY(R<^@6%#_&ITOR2<[:+>2;Y-FWW!G8&ZB NQX1IDTXLY!\SU
P1?DIZYG)(1M-XA!4]^;=#M;?_I85BJ;*P*D\TPJ?XMP$;F7L.JN.WH"8(/-E!)?U
P@7BQ"D'5KF"!K'#KUL+$QVV:7I\X0@])1N(1&<:9/>%XU$'CPNQ2W$]US=]1%J'\
P^V*4R\F#RWF+0:JKD=O4S],J7K .)H(O=X@WWPI_9S.QVL\Z21I"A9CD7)N\9GR8
P)P3[O((,9!U0#7ZRN/@!S.W\4X.-"85'S(<C/3'ZFR -L.8H(30:+72+FW['KP6V
PFAI 7.-Q>&4[O JLJLK5QH]\L62(4L/N9I+22T(T%")6]WK^1HQN3OKW.9X.XENZ
P2A7;P0[A^>&C9RARPJ,\ , M2CS%:V ]73@)A[ '):)1P'16*=:XY'(60_'I8I/0
PX2B@^CI[3$7B$=([VOJ T^"B<KG[<G9$P(:P]T;3';]$8/6:+ZZI[)S%K"'_W6/5
P%._)96)T&ULZ46R"2%7ASAVD\>9.T0(YQUJR>097 E$O_=T@-/%Y2ATQ(1H6H5F1
P90CH5NIR%;N*Z2-OO)!14FCR.(QL=V ]-](4Z81HGS?_=W'<6M#72[M1"Q5NS&'W
P0,#_8^$U-DX-;F36KYFY/QPKRK=O'Y('$Y,'9Y^'U>"&#L5YF2V4,Y M\,;LB00W
PH-RC:/4"YL]5@BU\X^XY%V$VE2+,V8S&Y.=,PR'%-$EBU4GV5^(*X535&X1G^R*:
P*>CQ[T\_4W9\G/N6NS9$V2%0?J0/\6KV88S_5WO<C1N*WJR/7HHR!F;?^?">8ML?
P*7*MP>QEP[F]T6/I185OB;EX#)^8H7=40[J !ZF?""K9R5"@3)7=V+<=A]-U;L5F
PW2J X<(B7-V=Q*(SX.Q@]'(WA&]J@6<Y8J F@@W5U)2].#D6]BJ[KEF!*)LH\ATR
P+T?3D;6H=6:K%XN:,B&0 +D-K[W_62@SJ#GGEH%9;BMS;E$#3QRDVD<^4=J9F17%
PAR)[:J>?MGWNQ^8CAZ8MOU4(=4T%K=WK7WB]^!</PG%'ZIQD4IVJ+$,H]A",//*V
PG);6@@1_402:\*V7@A9;X'[V<9JFXY_.D&KC=S"+Z8-9L C.D^F[6E#<>*GYIA;;
P-]!K'I[V=OGC;43ZQP;Y;LAR,#($5;K*:7(/J.CFAK7:5)B\_>2E3Y/'"JLF^Y[5
P;]EBI, MIDG4B(ZMLOF);ODJR0E3BWZC!NU(%(HH)!..7L"!H2N:E'QZ.WD5PB[A
P0,2^TG>!8IT<60EYFL=JZ@P V0%+OL95 K\1/,6O*OQ/_1H&I[PF8WY*! '6!&/N
P-&=&(:3P.8RA#5IF'RSMP^UN)];@P\05%K04QU=G,V+X\/:S2F>??1'T69 >!. "
P>LXB$IU>$EWE=I$DF+BGQ9<:C:;7SK8+.]V'T^6AN]<2XDB=-$).#)M02Y ?_M)$
P#\_+Y\;@VW!<DSO8RKMENIG4S%TB1:M1N3(9DRBA=;)^I^.AFYHB#9!W$MSW%+VM
P.Z8,BU[TYV>U&%9XFK29D2CU$K\D]NS&8;4MUB^Q37$V11@AQE^-GL<"2$'_VF@2
P4@(J$[M'3CDKU,;G[[$#G&_<Q)F'U,-? ;^X[@J\4]$U\2&S%%_ OQH$=_N*V3ZO
PRUY0Q^S)9=60TTMJH^E<41T&2<R.-\^Q^N1A!(=B*'"!*RS>T,"#D&8XE33@]X&C
PC$++NN9-!Q6U(^+F,(@(#_#7G2/PZK&FNQO]6W.6!WKPQG;C^52W,5:#$L&2R>%^
PKBO[ A;\%E2U\EH:7OD=-WG4)^+7/I>S;XR8&W"A-,[J7T[DT#.M: 682;]P(>,]
PJ6LGK,MFDM<,*)VQ[XS2I$]A?_<<^@"P>318EUU5<0("3VP'(K!.09#[:Y=+)Q(7
PGG5GS#GS,C?7E5,RFP;D1BG:U>6B8SS!Z/I0J_>MZ]EZFOB_+_T C[.**APX)M=\
PV<)NJ\%Z<7M%1D<NUNLP'0TM25?U]26Y;0@F[R8]LICNX]\-L;O^!$4V0>N?95<&
P6C5&>()%8GMS!>>B%LYQ3X" GQ=FBK(?8PDBOLO(R_U1MA4R_@@X\9J=L'W&_U)+
PL-])ZK.K,Z2TBQ9\[!9'!\)Y\[-HS/^",JIL6RQ<CQ?;;4E1CMN%U*I>;.>LT.:$
P<WN]$^6J75Q/QBGD7*%7OCK%YK6 B'_,N? 2!HA-F5/IU&&?1<_N4RG[QY"+'@82
POH_9N(%'7 P3;7O-_E#\@Q9A+:/7Q/C*D)/9\TN:"_$S#TRR]UFM",U+/*E,'Z9W
PW8W^9@XJ5P"4A<Q_S,YNWK@?1'Z3'N$;CMVZQ)K8GMY?54"Y@!T06(((Z[).7)S@
P8717,L5Q<:%+QH:0[6D )XOB$^4 %^UC*0ZOHVYM;Y K[LFSY;(C2S\V"@H$^S]H
P_9ZH%22_%$' .X]%/3$(OG&-U8SVPG9[4>4*>I(.KS! ?)--2TOX3;A#ZI9W9>F;
P7[10YY!]JE]"P:<$G_@]%W4X?)7M1=W.WLP@7\ZK]/%Z1C(V&0!=")^V/UD_8<^\
P#"J5DVJ6]^?CH$AIFH9^C@LU>5RH?*J32>U:FD)99E1.S0@/OH^D4O)C)RD& %_%
P_^^20S)TI[% >#7\:$;14;;'9"B2$$:9I)!')\U*O;TIYO41&4+?BVGV(?S%E2[B
P$IU>@>WV-IXWCETO\F@:D'65]HB&+)"W"@V1?]LCXTMN2G1W/="Z7FE9+S_NZ^-V
PTH$% '9N%0.A6\=93558P/F6W@0A?2^^QN2,JLF<UF6=_<,M @WX@\7BB(O@R94 
P([T7D5AS[6S6SGW=O%(I>X9EP%E[N_4Z9D:ZD+WZ[1[3+=;ZC0^K@X@P5D:L-AFK
P\OG1GM1V )B<HR(0IIAG$045QV)/-X 61JSX3UYUGM'&9).*^%X5$%!TXX*5M&IL
P,L;/77@6_'L_8(C#J!&O?WN LM']";I.E^MB$SE763S0R)++[?VW6)VMPYW-H6@P
P"0UH(;KQPYSWBQ*>_-%+=NQH[:>? D,',8UCLM74[_L"C E[XAL&RV_/GQ)MKCLY
PX(A)$J&EI1I$SP.AE+_Y*MTT_'-346-!L-UA**%&KU,,M7#,0^C2MQC@<0;-V3>1
PDV,_=VU9;TIE*_= ,;@>_%!!*DGJP'B69DJO@E7QV0'&MB3QC3%.N 9>W+/O_)K5
PGY7C;&^3N^[LG']6A%VF4/ZR*GC3PLR(85)/HX[,Z-6-[LV9L7"KWF$>PVQD2</L
P"N]+L.AFCY[5T#ICF(+VSVL-<F1AP$.-5.*.@-DRR3RWBKNKW9*9[;( WLPGI!60
P(0S E>& M*WWW/3,$Y%K^5Y86>]UM.2.BT21MKJ,Q/@<QEB-=-?AWWZZ 0-RR#!0
PS0RZ98-P^0C.0?Z1X>X(M$4LX?A4-A$,%='^D7*^J'%P[+G'B+<-)+-S- +/3ZCN
PU)7PW;8. V<D%_QU"<T.DB!U*CX&("*J;] 9[387<+\@=G\Z4!S\]E\(GP0$_U69
P7.6IKRE(8?)>*(JNJ6)3WTF- #D6P*CMX59 X[EH.=S$ZS2CBR: ***O^I;=.I<K
P0#XJH1>HM9"E OE!;Z- 0J.807X(Y)Q[DMS>*331.VRJM):04B<P28G1>QS()%83
P74+%HW0R_ GO%8?:4HXQT U1U7J2C,/=BO%HF=ZUZ5%^??DFLYNYJU<'1II>D4Z3
P;GR-;VO7!J02=W2E!W=+WSX&'O?O?.[&ST%L51WHUAOWA*(9M'34'FD1P='[8^+N
PMU'^/@L)! PP].B6TG $'13@)(AOEAY![RFU"[-B1J5GCL9C[BH9&3>1-%>UWTMP
PO2KE"^[M'7[Z>7Y]57L_>$1*KNGQJ!*G=U8-28-N<)5+%W+8_\XF )Y0EF),TF6X
P/L1N-T[_)O\IQ*61T0+Q7BH6UW!4-8IOI,"!Y[8+APVR<W4<5TOR^"N'38V*O_G#
PZCF!M"1-TE>%'V/_:2;34 HUW:%8]EODH;DJ.;!X3S04&+2A-2Z49%\,<Q6M(- T
P;X99?K# S^%UE,[/$*C/1QG1NKGVW$,_WOH[!J= M&DE\E@GAHF*%M!PW_Y,9!_;
PX@CYOY5OF#X,4_DH#QU8L5=C@$)_>_T[W1F:)",1YM%Q!@</4>*QT5&Z@2HX5G14
PY=$D &W4M#F_=P"0@=-UKP"AI&_=QF8_?"R$DDZYW;PM1<-.H/\LL*)HM VAW*?^
PO(OP69)R]SI[!],:%%/)@TZ3TLQ$Y"7(V=64TSS^>SVFEX8"<@;@Q2Q(8J."L4SM
P\^_[UUVJA3D6P#ZNAO99]6+ L"^_D:+\XIJIC-PFM#H<<$FC]+3-<B,E!#CTU4 5
P=I'A4J"P;9* Q0#K^!@7X&EN/QJ9L@T[/-*"+3T4KD!;<L8]B__>(_YQ -45$%%-
P 4:WZY8M!(4._>WD?L$*\^]1IYK3'D*>'_+6H[YJLN31>2K4WO.!$VN86IJ>P8B]
PY/_)DH0SH*H+AEQ]TOT7 G^)\*3@\$*44-CO)^Q56WG1O<($],'Z9HH1P=(H)^ <
PI?;%J%!*#B$'GU+86WCP:L81&_Q#M=Z12<"34L#RO.5=Z,DYGW^8X;*C+V'K*X25
PK"$%]ODYF2:%?XBKMM=[2V_)!4-.C)5.T*TV$!XD3S-*TB!7/__ZMXB=ZSZ9:U^X
P3-M8V@P__S]!!OBGFEFO$W7$"H'E+.UE?XLQ"(FV<2P,3 !<[A*O;L/W)#N+91T+
PC?($,6+2"$"WG#_BQH3/FD]]44'Q^87LS%8;4Q@DX)7@:O.F20K3 M4;.#M[V2%/
PN0RMOR*ZS(4!!H62((SZ\NW0L9^@/.-@:[HWZYH8A%!Y;]@;#?*K6Q>A-L_7 W<&
P"*%%3U%*P+$]ATP/ M3S/4O\;DK'B) -FG:>4C9_+7I$;WT:_EU&DE"FY@%]]2L=
PXT'=*2L[IGF.>\N];%%VYNY%C#]<S?I?'VUPFS1Q@W>D0("Y1D'(6[YYN-<H$TI0
P*-Q;\6\,EFUH<=B)C"<I%,Q/:5O\'.O*H-),"'2=LL[5\74V,YCV5JI31(I@@+/>
P''1J/PIJ&$M5FGU$VK,YQ2E8>BRPX'C3F;KPH5T9S!!"EH.(/=B+53D'$P_8:^^,
P43/Q#V=H? $.U5Y6KE*_234M[7\XAJ<V$></D.G*Y@:W>15#1?R2HB@I[V1ZB!::
P6V6L Q"SS<P6+O@J/HN X*&<M_((]^.MZ(I;5#"//CT%/, >/.<[X>E8BJN5IA=I
P7U/%+MP+)<+G4NVLDKOH>UX)C/#+<:UR2)1Z+];S(WC58F/TA\/+\KERO!S"CDA4
P?S+WJK-].:UH:&K"+5BEC-+J5K?_*3S4) UGC6&-?\S(#%L%/=XPKH%^XHV/.86B
PTS-L2TMS;T4/QS0IZ8CH_XR<[AGPSB^T+/-6/<H7&7B \K96,(;:/DM!58.AB6O2
PE\N1D,X90873Y$;_%Q1?YX=[7GXH>3%'B_Q"IY$(9DD-#J1Y:A=E2. .0W6J41;N
P2AIU]F%*X/2%:J=_.5FB8["^[MB:3FD6Z2,_$(K(48T,&BFH[A_]B:9',6Q][>F-
P%UJU7I1<#D;]1Z!/#)_O<Y0>TN U0HE]98639H@ZXAXF2='L.A"OTS-$S)S-]O8.
PCG$?[\UI%]+^ A/5=BW@X#?_RF.*#HX9A0@.!)?34E0T(UAIMS?0#Q:W12V]!.2I
P4;J&Q5C0X;"G1B]GK7^CMYE;]DHL%;OFA'!0E*@0'-5M?_+8,@-VT5<[&PFSJ%#'
P!#'7W$@S :X-NU$XR$RX8ZI)?YD<_=G224LU[RX#)GP^9<04TAL& 6EJ-O'W.$;G
P]_Z/GE]F"^SIZO9Y^.!@K(T01,Y<UAVZ%:]<_H5(OMT/K8ZO/[,;)H;Q=B6R>>JI
P+V/V@[OX.=:\G& PC@"N'%(=6SG%<X>Q\2Z44;$T,#?"S:B>Z=O[JTG;C22PY?&V
P9G.;U:_*R0\.L(,EV:0SC;."_C%[6&C(6RVG93*HKH"?IH&%Y:&"O\@^!'H+E/_7
P:::C/URAB4DW>\$[P3=O?%;Y<7I>!)U#2(GGW=PM26>/)"^E/% 'C5!EFZB &+-.
P>O&MO7[?SEK898W1YP#@/ZUTS' :3-CP4\","W+?.<&_':TX;,?AW)VA$*FI]B01
PER]P$8I35M)F(6KV-\,DIE[X?/((_4<0#?9"*MCD]4;%G:3D]]"L5P4S:89A6+TF
P;,>IDHMN3+'T^B;0:.8AWQC6T?'A6,DJ5]E($6=U>-"R!O;IE8RH.\UYJ4^PWLXC
P=YOE;^"R#%N%Q=L,%UX;YR]T=)ZMM![&+[5HG[:1[FT']FSDS!>K-&B,6?]#M<R$
P@^_HN;J^*W^[RR^=9^8HB:OC6^@1DQ>,B[(R[EN@-\-A4_&+$$%GH;O:1=HK5(+7
PP?]Z.UNG:/N(B(W.\U.!X(A'>L-PWQ,=UB0':L?^/9G2ZCSF.)B _MW.6,LIB3PX
P(?G_%:W.&_R%S[S-R9E&5P64/LNV,9)X7O6N_%P:83<:W4(CS=O/%1F%_V>'W@1?
P-X..5;3M+R9HLS+Z*6^@@?ZO?ULOH3(8G#9IA><H(F0$_D+^%VZ%,G1S<J%*9?7A
P$\#OBD1?&W-H$*T70TP.,A>?!*IZ:GJMBJ,3E/J#;U4B1M.DLQOH!8T@Y0.M/&X!
PG3(#:OI"S^?/87AWEH+1V]7B[A>H\$1/ZE**5F&Z.VCQR>"B>$!$?/)WPUSW5_FQ
P>+(-Q9T7KM_KGFL"CN2,2OS8(-TV6Z67#JZ8=,-U%T:#2^43I13.WDWA$^ AJWI7
PB^@SGN#W2/H9?=/CY7E0[7E!MVU98==OX1\^^:G+B7JQ ZK'_FNIXVOF#Z=9 /'I
P\'M,V^Q\OZ8'4?:<[UJLS],VA:ACR[TNGNHR/]-_T6Q<-B>.=R0/AQ.,?(_5F"B0
P81'@"T!FD1@L=P9"+35RC<Z>V##'C!4,R\(OA/D%GZT396].ZC!X ([>RLZBC^0^
P;5HTL:D)-K'@F?2*'$9]?N.0;_!C8E_^P[&>?/V@X,BJ=H)"=:!.KF2%VDNXM$=.
P4]GE^Q10O&N](3K6HOF-ZK,I>2L(O>>TUNZ*85 R/#Z8\0'9'Y&U>ZO?CN)$RCT4
P\K')KI:OVI6^]9#:)?8F</B!D&BC* ':#*ZP=#MP6>RHQI=;.=>R_0%I-6=&I6,(
P'M$\P4%^7_=]+[W9(IZ=I1%=@JMU6AA//KYU[:+=Y%T [@F4K8;\0O]M;"AW+ML^
P&.P^:J6@.;!5I>D06V\T@\3/D?Q[YY)6?="3H+OHV@:5ZL)5QN[,RG4R?OW3E179
PVP)^H3$YK6G^H/(E&_Z0W(OMT\_\QZXKX"T+</H(X*F_BO)![5M297BI<D(4<ZZ-
P:+]XU6/HXU!6"H^3WQLZDJD!=.^#WWP<Q-&*?0OAFPTRV>QX/KXFCP&XE!0(XCUQ
P)"8!4X9)P_0Q( [1&(67FTKZQ8\A;LN?X(D92+9GNQ36-J9ID2I3)4]Y6CTV?',<
P1R+:@#ES$^XHN++=@W@!-.P@4D^G3'XNLQ7$&:2M3T^2,L/-=W@,AM#"YC.WK!<_
PSU;@8TN\0/-<:="W_GSE 1G62M[[V!GS'.^NS]101U;"2>LE/^;]J@?K#4F2IO'N
P2.H[SE63<YNP=1R^$<]KC#SEJ??L(XU,-U]XYJN,IA$M)BK1]4F*]XBZ9G6U'OG)
PF$0,?/G!WQ?:GMC_4\<K#K"&#@B0VL6SBZZ3A$$_<I@LZN^23QR-";TFO9 #[^J4
PTJ\AP\A>3N(^F#SE4QS2QW 0Y=8NT]SWF44(ZIJ9 JY+*N+,'9KC)351]""TBMJW
P"C"31<'5Z4*]<X#(&LD>/WB5!!>JNIM\&00#315#KFAVWIT]']DX3!%R&<]X2L[*
P;[M29404J3$^[A%Q)[R2!A[(7#2Z/935=5;2O3D]1$F)%1'][F+Q,;<DEDBO>72Q
P<!2@E[-XF6N ;&P?+^K2)IN(I ]V'67;S[2F061AH+ 46*;.$_A]Q9L\1=OX['VA
PGW%5HEE4'TC7W;EJ=4<8E:+%(!U[V4E2J%8PF9-S+V%%;C382HY] 915Z"!SP_.B
P@*U&Q(A6]C+M60FB;4<79ID+J%:L%-MKKAL'>WS.0=/DJB&!&\'[^%9A R>4M'O5
PV+_XL20"LO[<T?EG?J-T*^^!1J096Q.C_36Z-/X 7A;K(^4T&B6'I4#93P+GA"W8
P&&NN=Q'1.JN03)OB!=BGR50= =1C3R83M)><*?#-@NK86K@-$F&SU'#$HX5V7K==
PP@+-T 9U+\MT"3B-/(C0%K5 ;D-YI%E/D^5LMHX$4)&+/$5[5T:$D[T7'5F.3!<E
P/ -]F(SYUNESF^H,)6X-JH1AG\O'0TO,'D821DSI]1?BF%K^42NC@@*5G-)Y":1#
P?][*!?Q-D17ZQ8K<>QJNHQ&U_*Q-RO! ,4+C1$@9J3DOVL)9WIH+I)AF082JA#F_
PFHI,4)=($M9B,',$';1,+Z,?^J#H/^"5J#E7)6"?^W@%#B[:'_AIQ<CZ%UQ=0G;8
PZ,ZS>*ZU;DDJ#04^T@=Y]2=H^J!OY(FE.(+/55"%:4[F9EP<2AL3Q.<Y\.YL$Y0Z
PKB;/+1=8<"'A>J_5"\A4E@GE< >A^WH+'_9DI@[9A^^2 Q<25J7YR+,E&_LV0>3M
P=@$F\"96=GQ]>\F%,/I6^DE8HZR3'T"3,=4L:9K3R9Z):D@KQ+FRLR376V3SA[;-
PSU!C+83N-D;E:FG8>^]ZY 0J%^O0_8YH0N0X-E&/X#5V&!2KG$J;+.44?043N$Q"
P(2 $YUCZ8'@6?4:#YQI-&KLN=5."3_=U^)FK$!;P:LZE"<9HXW'R5;BP%PB$T\-\
P.,$S\HK=?C-9)62@.5 /WA?WC(Q0" $QDBS3,/%M=^FZ2Q"+ 0Z^T<:Q9\7,,,Q;
PGE#*_$0A$RN6FW><*-?29OL(G8T FNPV&APL0M(%"/##IR(E_^].YC"-I.UK81'L
P!C$K,H1W@\Z6;ZJ9M<*F<^>/S_/(O'ZGL96RG8:-K9>4*]T<H*AOXB](ET1%P5O$
PD,M96+]R47@)V];:G+.Y!\6RN8/JLVERMQV]YJD%R$S=@&Q;J ![&S'/]& 1<6F?
P<WR?6>!WSYTIRH.=ZJ1\'8"H".S=!/RO*3ERZ$A4OY"#W= *PA63O(.>1%:#N^>Y
P 1Q+.R3$19MC?P,3Q-X*-N7 =RTP]K,FW%U-2!>(_ST+:V/60'QW RP*&<5>B#5H
P4^A%C IT5\=P  IX"5CA"]HHM->1!0>AOTJ;B!5\_0L\LQ%)B\3/ES@NIA7M7PX(
PZ:)4JZ"9>]EAOO&$^#BU_@QF#=WGDF_N%/QEWDC<RQ!^=NP MH[MW69EMI@1Q^9O
P2D"WF0=&UUNN'EWV;UAR%?:4,M.@K0^W?:TW':6-H'+@\6LN-"NKDS0BXT,_?8\]
PJL'UE*59W_*4I:7C15%177:G@[,2UT6-[=&0W'L5]5NM3-KE=HAA2/N!JV#*J=5+
P;G<DBJ;"W&5X:4H6V]3C]A2(UX<HM0)RN]E&\>.7R_PYDNKJ3NZP= FZ'M#G_,_T
P:"1[=6!DJ5NK$1U)HK*_X?Q*>U>?G*/)<04R:N5M+[G7!>H_<NC8YW.T&-7YN11?
P'RTR/*;?$<G 8"A/YN]!$\Q?LNH^G:%#5J\XB,UZCT6?J:25D<>?3FSOV:IJ0HO3
P#*ZHP_*S9!-?H%E?H V4T]A.(%Z/$TM/ '^P"1C&.P"W0Q\G?&H,_.F^*GIL)A^>
PWOBT[+/F;1:16D,=F,(TRNI^2^&XKN2K)QI,S>V#U[%%5UL0V*K>[%VO_!2"J,[H
PU,=^-UTDH4/X1=VR1(W\^MYC4Z=2-+R[-(=L<-C+L*EHB>,-S".-_^$SG3+/?CE"
P@G'@I6>R&VCL<OF!L$-)AUBY*Q(ETXIH.\E!FL6/H2LS4%(0W_+(I@Y9N@P!V]]-
P=(&#JD]^%TQ_36N6)7%&=_HNP]N&=+B-U_ 0<Y#TLT^O+>V*$XM^A)7JE.EH/2IU
PAUH8)>XOS/- OJC4&XAPPO/4*R @'9J>GZI69><B]ON E$@:1SGWR'?D&B%LX\B@
P;?%.[P\5#7;'/NP;717/KV.1N(XYWWO8Y\^'GW)$?2HG<O3\D!PX$Y: &=;CHYVN
P,X5$J C_7<T4A+- .6JP+ F7\D/E;=Y3\R:ENQ<W;W6B#?233'YC3K!9YD)M*HT^
P;70YF,@(>@2C+S\(*:/!7+F-;2/9YEL+0":"YN_S=AILU4SF<$@>Z+ /2^T,+M=L
PB0'XNT(-/SJ;"Z#?@^%#/Y.?DS_S$A\>)LZ+22JO^A2>*&Q<4@!88BL@M9>Q0,8S
PF);<#*6.;D'7H2HJK("$5S.:LRVV!/D4_;>FW&/UR@I#7VW*C,!(W(JDE\(\M(4=
PGK!'$$.1A^=>]?3TO*3X@3.*# (X&KN)0PV_<4C; K)F9#.5BJ;6<OH8 HMZC.%:
PP#:^7UW9Q:MP4W'@?ZSV$4CL[V%1<?+K!RXR'X3C0MRN2M@3*^6]G+VV(M5$9(0B
PC;8F?=_O)]831SQ6H KE1:*->V,Q:JI_IAS'U0F08PY5]RR,RM>)T1OF900!8O.?
P ^!&=_?%D/(Y)F[5Y78M<4AP<'%H-@61D\:9T<;,I%OGB+E=IP"(W-23$?%IBCK4
PM?MQ'_)I5W6<IS7G$7AT7A3D^HH R2N;NPQBPOA#O-79OL K @;3 ?H"0LUQJWB:
P_9($^5!S301F">G$4-&AQ-B6$Z3"\DY,<'MB$_&H_84RA!RE\E&@0](\Q63T_DV 
P^O>! 0(>,!I\T^R:HZ"ZUL&X$ S!4GK<LY42VKN0BIYF&Q#$T5>4&]B,*_='/NZ3
P@.W'(P@4=RF;40[A:!(ZI+,=(\W!-K'C@4PFE4-^T97,:F$)TT5_+)FXHV(7R92K
P+9BG?(/CN\4Z>5Y,1I7'R7EZ_\ 8%\T":B\B/-S\[3YRVD)L+.L^1(Q/H!O/HMLB
P 0PG3N-R4>;4KZ128PTF1-[[; ] 7R8(E+V10-F HBFHRU)5E;4!6GA*Y<JHOF_?
PCGL0PI9>Z4%+I'T+\Z2E" #<]X!SK#86T(?=YY8'4DBT E$\..*A5VY_%BA"M;M0
P%"*M$,P-PNPZE =!!)=3=BLM/B4Z[X IX%[#*2$1[7'FGE&E7ZQ6I=^4TV "*S"U
PQ.F4':\A)J)X/:H]'O1B%#@Y&!6H/+3M+W<^*X"&,"ZX_O=\,%$E#XY+C.3N?43<
P91-5TD0EQOEK6\/O<8=#0-:G1RNP_D6D@(&);EJM"S,/4NPU@V\'(6&LYQE5/5YB
P\(TFM>C2Q09?$ZO8FL?%7PBV0L$6/58U4<KR1H]:Z)("<Z^Y;@4F:!P5]?/^'/1V
P$WUBQSC<Y1D/4X;Z2)-*ANN[+X7;*4">^*#=LW<B%W(5CP7^G5ZZ".+Y0C,U#N#S
P8T+$6RZ#PC#[WD?2M4R6-2AVN;TLC4'C2.80*B0P<^2$'9DZK-5IC&GW*OREY=9Y
PNE>2RD#.0;%64M)\GV [D3]<7)DS7J78EJ)WLP-Q$S?>IW$#-=BH#@HY+4[P;+A[
P0N-7,N7DKX5\YUL%>JN;0QF#0<N,SJ[.;]8PO,]\Z# :%.)9I^?T^V_$#G%1)TU6
PY7X[3)K+-^O<@FP1R&<_0<[!(E2/09QV;"@Z$ENQOKCADH["?CB0:4H?$!N:E4I?
PSO VX9(2/"#P%##YAGJ4-^@/3V(J-IQW4Q"EX4TRT]-5?QVU^#4W4;).F=%#N!!8
P@_O*X7J;E?>OG%B(UAM3+ OG9[%+221T?#1O@_W 8-KZZ@(^!WT'14 1>\\LN^;(
P8V'%>"G\\K^DQ1-A6<0V!G]?I + "O>A>@BTZ8LM@%\C!GZ68OE0_7QWH%FT/V$W
P_<F72!41,58G'3E+?I**V(%MUG@AK8[.H<&N!@5]%?;A,,5&=F \B*H?LB-59_BR
P/_)<"8!?&FM^%*("_@<W1#\<X*3U;0%P>UWA"$776=SKO$U:,N"U'>02QNOH"D^N
PY^+:FK78PC4(=Y&_H4&[/F?FXG@ *-:\WS_U?59RYY[-DJ7&?7L<2$O(P2;44WP#
P\!8>)4DO@IY[%UZ)_7P0F^18.M#/-J6.3.;B'Z7E'Q3<7:'K0Q1_U!3O!9</OSU5
P(UTSU^T:9.QJJ&(U#:CDCZCT83>#;-%1,Z6'"09L\6%13A A^ CE)<TILPK$C]*A
P";Q!-!>B>DG[[L:G1RNZ'O9PRK"BP+C)I0>6NX3^9;-?U!XNZPVC<,9<=_#P:H]R
P\66+VU,C^K:7I-+H@.S=Y_B[322<ZOE++1M1K1Y9Q$E.'=H6.A+ P]VRC?0@M3-4
PWX!$NKM>Q3<:.FSPV=#1"+&K.X6>U9ABC?[J,GR<N=Q('EW_(/^3E-^ZP2\YR'O^
P%,V*=C(\G*4:!OD0\VHH7:B71!K! IU9T8>O82;GR="J*IB,4X\H!P[!KS+]G4[L
P9"X\ @ NQ#_O5&&/UV!K#?%='E4DY+JIA%&561<QY/L-$&@2+_2Z=I7\CW,O(>@H
P"]"[0QO$B6$#?$KH:>)+1[1_T(I@Y:U(>:L)-&*L5M]UZ$QT;V2:*( .5$@A(+F5
P@P\K-@5<6+B@BSD:[UHC VK1+6J39=&7QH>0K$,DZ%.#ON2W34^_7I[_@[:^L?Y2
PR.JUBX$HO;R\I:,+XI[=9JK)UY^4FJB7B(7Y/$XKIS55(MT6W=;>U>?LI#A[!ML9
P_+ZSW.''T-@-V8_[GHFE#_6LL3#)%0=8(R-).9=(*4W,;2D*JI;&5O4[Y%A,BFM.
P.^RI_QR*2W.-+*>\=M Y#;*S,^E3='R.?QP>3?XH&5E*,6@HT!,0'X6%H@"*7+#/
PH/0^2]_!R3YWS$,OV%7?)2L<F8]Q$_1[V_5:@LC\_9WTK\P^&1M^,(P;:Q(TYL])
P+)WAB"^@3RC8_J!]S[/RP?#I4/6E6>_V05AB9U-W(Z6R.6K@<\0E$\S1YN2D^"_E
P[-@=;4B;M1)<R BR# /O,_)%&G4UN..F(\Z8%HL["*"LAKU4L8X58?4E;FS2K\S3
P..IMX;H-,>6D66_X&3?$".0"H,)%Z(E<.8IS.2LO>S(@XXWM+0%??X^D"IF'/(R-
PA?(53I$$U16@L.J@L3#J-B!H9D$[$]^GC$<H.)\1:6?#O949*U%CT%JJ(.TS.V#A
PH)W7)];"!U2'!LS! %?><WV)?C ;J3I(=ZP"GD:0(^"0>?>&N7K G[D%8Z8;ZRY5
P:G5"R/&%5E1(\^:][ $;[M3?V3L)8CT8+KN8A3OD<"H",*I3(#*I;57H34CVG\]1
P+-)_CF9A!2EW@(H!+;#CRC4-6<RV:EM^SL7QO9D<7Q/"MC"A7+&:XE3P]7K:" VS
PH)T!.Z'UL5>*L$J&:.O2"38"MRI>^ZQ1*_)A'*X:00O^>A(YRNG/! 8J25P0Z25#
P"E%N[TJJ<X0S3Z6'8PN?NS@P5\+DA 49ZS4\ $>\8,8M:6UW1[B^72'IX-+Q8'#"
PN7YDF[.E44PQN-TEP6/ZPHX"5@\+FV7./ PEG=<=%^'#M5J5'ZV/G712-5H#CCL:
P:H^GU2UM3&Z/"I"*A^)@/"!(G%D0(;3A,@"D0Z:>5,&C>'SQRY7O%Z3)ETP//X<H
PNX0^0R_/*K.T54FQMNZN8O=X;LF;9@J-B(DTG1S)++ =0Z[&.P;5J%OKFJ$W==5&
P91-JS&07\-:$4E91<JC#O0 8F_H2=J]OO5%G)&*XYS.2Q*A[H8G('F^@ETE"#6VY
PM!C [),ES&*AIF1E-%3 5B)0BO&CIQ] :K&I'5LAIYS$*'QQ1[H$]V44LGW6? !S
P.8#07J]BFMPNKH,E/T'#*2<9]N8RH[&.(['Z27E7V*^&3H*'L8I7EQADBT,UOO$'
P!L66$ -7;-A5XT=2B_J&*KPPC3(6N4X!?#G:T?$R'!.\WD-3<1.'2G 3$L,\:;TH
PT*-LB6BYB -(8/"24%8*D!F^F"U_U$41.7)<@B\'G$+JSN,^202P=)!.\WNNT$IN
P[D,*ZY__,?9=VV(-D2Y2,8WL$*QW IZ3.B?_0 ^'6["TYHO03;W6"%VML5,U)-E%
P+0[W_,]8YZ?*$S>XX]BX!L*#B=MN-R!;>#8C4ZB*S%D!WS2TNN?9RD"9MK@]<PMR
PC)VLV2E5K(K^R7]N^\?!(RG]\)3YJ\]B!8'=S6K6]/PV- &"S)E' ]U@Y]B 7EC+
P.@8C TBS9EC0L]+HY!T_FB3?NC6T%KCU 8@A\4.BV^54D75@:"Y7""4&O<X1A8#^
PEJLGIFJX3?MMK\,07 ;N$PHWMC>H,<5A^3+7<2VA6%K=A D:IKVDJ@*&>>LB#+M!
P#YZ+X^A%[O?DN&V0@LB,/>5KP0SS#BCL]*%0U5(Q B5%&:AC+O('BT2W=%&ZX,\#
PPG2;4_\E**__2^C1B^5D2,"_(9#.0+W6]RZZ35X <AS>:Y.HDA ,2S;:"?-H,<B=
P5NCI:?O\W>$*CSQGKZ!5FP>V]+V/XP=:1)6]L-<LH5D)1A(173Y4"^QI%*"#\H\@
PS%K&;RM/BL(()]CB&/'7-DOI+,5H2_%"J8!Y4MP*/0*.BP4<AV>7_/9LE]<!%ND=
PL7S,3$]N71C=[D:V9NB KQD7XNRKM*B1P#:5G6)L3Q7;88PAZ>TE&]L<#6D11@?I
PMN#+ <I["7<; ./^ 8]A##S)M%C3^'"0(9M:C:SI8'!>\Z,P,:X>.3NIPY E NR4
PI_ \?WQX$ESN;]4'.#:^QD3(GR?&K14D_>S.Q1PIC VMR\T2W2^I=O-EW2K(\;&%
P<"AZ3GRK_D:+!;>@:N+SQY1<:D%>B/_*Y+.9;?2Q.,RI)'*_]?@'F]Z)1.M?<K"(
P/Z6STP<(=PO4&J!^_)Z0'Q=,!Q:>(3"=,0V[<G%0>D?]$4Z$0!"EJRW#&T.K"SPT
P]8@*V/"-.^3:"7293P@?:9KLN.N< I2<Z.!@RXLB#ZHO7OC!@XWRK542LL,/CO-E
PEB9G0*R$<A;%*+>MIG<ZWA@&EER]I#BTQ".=N3ZW@SP#8[;*#+U0=Q]3L?#XV^7N
PHLMT/BI)DT9&Q\^HZ%(VH6**O%X_/T%!PJ"D?1\M^)$WOA7(@ RS-L>"-R]WO^KW
PB/U)7.),T 5"0C37K^._1HI8JV)?MJ0'<LZO+;H::'ZF.<JQO]1+RDJ6 =?K#5P\
P"Y#V=L*7.*F1_:85*S:E"X!SK1(A,]6FLE"DM6F;@2H QZ^&LRU3?"G_MD"0GC7-
PZV?8NMI!A@+21&SI0+!(:#!N:!VY;,F_BIKAO>6+W^%IC#TFO/-":S?9ODEFP"-Z
P0K/7XB_D/TLQTF)I7[Z#VSBEM& K7_\%S8:%)\B>T>+A]-*VLP?P ^O2B\SF%:^U
PFKJY>^\E1FM%!RI06Z:CB##@\'NY'U/EKCG(;Y_LV<.^<+7"H^EV\,]>]4K/1-P]
P.$1K*S73IV*DM2G["W7)"\/) MP%('OT\ VXFZD,%[.F<QTB20LK( 9A#'3\I53L
P!L#6GYB<8&I1&B9T05Z(K)KNDX(H#+US^UXX6DH=YQLX$[?-([T!)N(C+DS[BV+E
P<X%R155/V:M(2BZ\N+O,@!#=%'?D%>+/X4+NWB=*N4=DJ+01LZLFE5CG_9A8BM0#
P).-$HR2IR,N-'H[1@ 3 ^G7.^%++.+#E<;_S1AS%]XGYE_XH>-\0.H8HJQ7S7'71
P]J,O7F5QD_9<TFH$*&9)D\;W-*STSE+IZ5Q2R.:@BVMTT5*9AK=I@E24,D<A:P5!
P6@#0.<Q^U@O4]0M:2@SPE&V5\SU9W\R,<B)8?.VGK)BP RCC<;9H0I6MAD.TI6E(
P>QXRB39V%U4MDY<N:1 %S;(*8A%S>J6*79VR*+\4>.=B,9SV>O@2_; &:%SI$W$'
P1,?G?AO486M0 *6=[C877LQY^G@N;NKJLZ;81J^Z]HCPVKLMTK]1>686 !M\_F>"
P-9[%E_K6TW*HE]'6'-^L?VZ@8.$_D;3B;Q50^>9(C ;:6AK*5;XEH$04)[T.HP80
PRZ<B'51-793!>_IEDY%L&8B@]D50OQE!S*906_4&(#@(%/RA?QJJ<[ 5NE)X:C_-
P1#7+/)V0/>KJJR@."K3U:'!2'=@'>%?=D*B%;F^!\UT$PD-PKYWLPP8'@<N'COXU
P^<_6(@"(B\%(8V>\-&:];DR!<,D_JQWY63(<:$K%?&YE^P+DP5.BD* <^L[?.^!/
PMB8-2-C#N;*@A-8@@G":TD?-Z./(R)BOO(-:5)#BI,P_=-7^VFIVXIJ(ULK?PGW'
PT@$SX)E?VV00E^<(+>34+""7;.<&Y8$ON^JCL'_A![;L!A(%DW].&0Z*(N_;I\;H
P@Z-)4F:1<ETRU2V$NB,D>284@$PA!$9F[(0>@!,*-%JTJP[O/=-\SX/3N*)WV8&A
P3,B _&5"2)^.*PV,CN6#J2V<T:NCT"^UD:]MKM'RP.;P NF$E7ZUE5/Y=_"(M[22
P5N.!"-R]Q^4JJ,,*J5RLNZ4LBRX,_I]$?ME)"65G##2\J9OH#RV] -P IL4A6QW 
PXJD@-C+ZN]O^N+YK9ERD."9"$,I5!D&5!"0)$<_X'7%Z5F9MJ'[UM9_RG&PZGX]K
PF^6M6@R^658@*L5S7NG?I@++;M,?D%A7HJ_UZHN_%(PL]F1R133*4P,2OY?\XV;1
P1BQEL2A'@A[@N\FQYXX *Z/[QS475CX*$0Z&-H/)EK*"2'3S85?U= ^[<IF!)7=T
PFJKBD*IT\/0O 4D%*77P1;2>)P@CC)S -X>3#+=*N$V1YI%GO7^84>IF'N,OKZZ/
P';_#8HHK9*2E>JEZ;I)0_*Z&W*TN7Y16Z7,59%D&%_P L',K-5L.X;M<YD]&H28A
PBC]VMY-/M(6K0=(N:!2(,8WJBF5'.7X._<CL/,J3UW\+'TGJ14;XQ[T%UDWIT-=(
PN6Y+_MSF.5 XFEC10OSC*0I5660X'9 ;?UWU(^;?--JQ*"[J'*R(V7WI3#^&.V:?
P]#QIJF"]88G8V?J+BEXB#*.U[8!,%WFWQF>!P'5S3OS 7XB&8ZC*I*%?$^GO(D:T
PK/T,O^[\C8O $BXG<:P'JT@'ZT.% )2[76+115+I*<(Y%=&S=V,L]HYFOG:RIHHJ
P9V1HC=\JONSPU=9&.::V#7-87@:=B8)#\*ZI5M(-T$O#,;B-!="]#BC-^US,<JZ_
P<T(VJ,[\#1-%^43??M<CLF*$["MXY]&L6D8T:%-@G?KJK/D+R]Y -6).Q$VJ<6$C
PMR_:A,\/2J]=LOHC0V_X0*#S8Z"V_%7OOG5K6P9H8$))R8N43C0CVF[7E;PC(ADF
P93&88+[9RX%I5>-X".4U2H?X(Y.>2]")Y/R0"RUI^DUJWW@G%7H5W<L_<Q3%A]BR
PMQN^W9!Z]VTSTI%?D"YDZ^B,S\F!JW1O5L?&0LJB.&2SH5*:AAC2B&@UF7E+TQP[
P0KL/=#N93Q7)SK-BD;1<$\^A:^KT86$#$^,S>;-4^;X)U:[T;H6*^\)RO&'E/O';
PXUAD1231VAOP]#Z,\WQ$HZGQT? WRI&4UJ_4G=)L;+WC,KJ]M.]FZ_+\+:\U"_A]
P-1LKHX$W8*5QW)J-&ASSU/3);FRD2>0SZV=7)C/?Z3TL.& C:HA38!GMKV/:@A7=
PY",:;]TDLMWP&NTO"-5\ $GQE)%XQ_%:@NGO9PE1!Y5/RDVDD4W$?EK;=5Z0=?+1
P SR]EP2M7MK>US_H2H)-"4J4FC(HZ=Z6K9/2N1RK[@@:R[FO&[_SJ)D)[/2:I7C3
PP:L:DVBD!8\ DM=W7:RUVGA%4@(9I16H%VX(' HD1JD,SAC"AK+*TX':>:0LT_7:
P3,2_#@OEUB,V6\]@D> \/FV^3K0][71-7D>DEB9,; U)''PW[KS'.N6["L4UOM_-
P\-WAE :64\SLK23KE,4U!3@30>2I<J"E[".*WWH4\&K!O'F!Y32#@;]X=>0\/B4C
P+\*]?JV$::A7]MQDC(W"])(#1#K"3</I\@[E*9X]EJZ)RGI.^O50[$^:+%YYZ@Q*
P,)JL//29[CPUM-HO&(9%)JL*E?C.<M:^C61T4,^P1N6=.+<;6G-K/#'C:"S#-=$Z
P#?#RHU=+0U#YFT^3-Y0"O:C1T=7Z+HV)6MNS-ZWZZ>YZ%3QCW6S].ZFM%)J2V>C9
P $)VXJ;JZN(=$SZA4=Y-Z^DK2[AYU4<(X<*4>4-IM,F1XY OO,S'4IIX.@]3'#<B
P3*(@6]=._[F?#&F_+;#_'S*)'AN;-V\$OQ:W&Z,IF^^<22"8H&P"KF+\_XPT+LRH
PAZ^ZL^VZNQ!+\B]TFIV8EO5)JTTY72^M==<VB,VA )E^VO?<5?D@1R==_%%0+-,N
PQ_G%E<#ZNEMZV-09)+4$OZFB:U.@%(G?5W4&#./]#6PP?CQ8;B\((II379WXPP;V
P#(DA*S6I/ KJN$0>WA/!L(A34BWJ.O:%+/=T98;:LXHZC>6XL^M\V<BC479T=-1E
P]C7](53P9"VL@[6I!S5_"5PAJ/*I\3*C)_BD@S\"J&H$68+X'X4QQ6@GE-,*YFAX
PW7J0\E\"-*\.J#&:A("#Q[JN.]S/K6+Q&()=7@!IMAS2<]$F.+!39/EQ2&+*U<E*
P(=S(IXLZJ87Z2!-S/,LP&:QXKI09,4@$Z%B[RJ XVN#<R94GWALKJ ">ZE[^\3JP
P<&L-3"Z12%B.-'7@)N 5IF3KM42'\I-EQ:NR;0B"F</%@!XB"2)6KEGHV-\^?'4W
PBD:@.'4T.K0K0R!$<>2YQS%,21E!8HQ7)EO LRXLWI\VBII""2VQ5<%6WO%"TS%L
P0GLZI9_]>W'J0\9/ZRISI+LVXY)&_V36<+^A&TB"MZ_SJB+N5]^B"K,@J8*.-08'
P@ ;W@1K"(['3#K8RE"1Q3=2F5F$T11@==D;\\;#[)JO5V_[NT5A"^##;W,7_?MYS
P2N>^[QP6E]DKPXT-4G.7V)L-0[D<1ATA]%=OL)_/K I,#NEB,2 Q.5K6G7>0MTX&
P#?$A9@65W*%<Z^%"44EZ(:4-"#>];)B8B'9^X$!'!]2# JCT2'4XLYZ<5_2]77;)
PLXIUK;^!,F%+\)@O .!?9*T_2A#(CS]9K/VN C<T=U$D-\=2AZ.*3OO3GS#N*CUR
P1%Z$W(DAC9)3!C6XE07L78#\D=NF]XP4ZE%K[8W/OGK-R3M;1LQ!Q&Y"$XH#24/W
P%+3A4,(+5"D\M.S1UT>M1X[T#FRSOP)X1OG>)',&LDK>13["0+2:@_C4K^ PJK$(
P;M,%[*KTG$W+37[+G&,:6*8";NXJ149)\RG*(%/Z7@PDD)'5F44/=ER4Y \?TKGA
PH([8Y1700GO]G4FG"_C-IASLM#'L+Q /L+"UW7TZ>&EE.TSB7\)FS4_\9^'UJP7 
PI[H5$<. ,59Z 8B.\'V.JB;8G1_A3?.KM\=@T22935:N4BYV:74Q;WQ#_*ISJ]>X
P[B92H36W;$&FM!!N\EP/X$3!\-ET8@HG&B!N[TPB)>O3XYK,I]  H?@P/2[I\-0&
P/3K_4L/@$E>%KF@^B(:S-<ZDH=P&IO3XWA;K'>Q2RV/QF];U^%WNJ(!UM@UP L%8
P[_38=LSU>TL* +')8,XBWZG/]\XKPQBQKF2LGY*N*;L=C$=BAP4"V3#>H^7;\BV:
P&]S0,+MU^%U8U:M8>ARP%S40#?9]Q(!.O_!NT2$K'$!X<UDB5Z&@3YAP2+X-D</4
P'""^T'/4D6X/S4R?&+T%A<C1Z$/46@I->'TRLVK+<Y5<@-V]-%9G[B8LUUEMH9[F
P%LGFV%4#"%0K@CT>+ -7^U8R+'5( IW\M4!2JT/0B2_L,VR7,(37L$Q2X%Q,(@#\
PNIHCB^')&@Q"O :RU=O<A)?/B .V[RVI9([0@0:"@'F<^6?ST52!L6"HR L#PA>:
PQ3H0#,1S;_.79_.+>B6D\[-(M3KBG@"ZDW!,H5N]\V2?MT4M$DP4>D5Y]H9"[BV/
PEJ$U6S1 +WTM-LQVMQK2&IIX<?F;*%IV[Y7S)-^-#<T980W+<-)T@3[5/UW2_,(G
PJ^N:3,\0;^3 G,;/*GJKM42=BS:A[8<%E.5;W (*;&B-ZGQD^=',>1$9^FUIUY;N
P4]DY#G[B"_Y]"<(*V_5T7B.7B'^^1PNWG$O+EK;C([)^WWM.IX'(6)ZUL#UI)BSQ
P'N$=79-F27-)DVEF'ZIWJ3.K$WH6PMX3C;I++2""=KT%\P&+:\>EBO@T_DP7M5KJ
P@5NHJ"D+.=JBL\9#=JU_N-8^7'V#.9G%NIU(1GII:& )BNZVE7S,)@U=%B ?X ^K
PZGL6%Y P:(YK4) BB\<T^>T'J*"%_-O\>'E\9/OC]1KH'HCH/QL!J+6$^>.6AS;K
P1E/A@W=,U'A=$,>3[N^G Y?%M'E ;]?]D((,IU[6#,@$>3+.6R_#3?GZLJMFZI+)
P2UOD%2?<=**LJ2\1;->@)-,E"6.Y&@/SZ2V//@:%,%%6WX^E>7X>P7][J+-0?7U]
PL5,\2R]\D1M/ ""/3O(HF@$J!KDX]GY@]RU;58KXSU'!#N=JZ9!2N/F%1/H&''SC
P\T1>S$C&62\3D$_[]*$FYSJMN:4W<<W!1$V="]Q(\2$62DW#1=&>LI(6:HH)0?2 
P+/Y=C8GW/0;V8/(%8+AW\@R*"S:<V%5;=KD7_'3>;@67M%1#ZU%^$ @/U<7@4FHY
PLXM4S4>9W45CNEC:S-D=1^;_QHT*ZYR=^7QA&NR)>8P=G1$HW?<P<\CV$S0]9;0S
P*FX4\NG<@B$7?H@AJ_^#T'4])$'$V;3EWS0/8GC%U>@VM":^%_6'X<==<KB$,#Z@
P85W<GC,_5;!_W]\<Z_6N]D3Q^9F^=[#"^68ZK ,?$9>;A2H*5?0WIO)61**3EAP*
PO%K?7=H<+NC'YZSB['ZI59X7'(,MP_@&<WM&K)T)C\4"2^O6G38BV1R^9X4:UYW+
PQ&A+,446O_\X)ZK%F+N/]A864XT=K9G"3?XHO<M)BTN^@'D%7@UJ[Z0N_'$&A=YP
PBU7]!>Z'G(IN+'7E:S%>S46;H.+%C1FT(PRMM?KXSCV>015E3(C*M'ZL[:P>0DZ"
P.2$DB'=BNK8^U@S2YG;3:AZP';8_G27"ANECEDL7)7DI3Y'H]YPIV%O$)ET&A+VE
PXS$)_P:H5X$$[$AV.-F1O#^4<]-F #&80ZG$#>-[/!"0J)I7Y.YH$E;)NT%%W%1U
PHH<WQ'5!R3*WT,^V4&W<(5;M:&;J^2$7*=7,ZSRS7?RH1W)B.0+;<?4OC+I0>^#N
PG'S=NN3?>DFGUF\<N501<TC.5&[6=G&AEDA#3@YRGWONGNA06$J$61R?Z=LP&:3B
P1NI@8X0LK**2W"$I-^@P'[>9&]0313E9$EE>^CO(,6)R.&8:GMT@>CD>JNQS\/!Q
PBJ@-:T"E20C3QTB/DS2 YL.\*@%T<G#'L_IXR* HH6%L%3KT93,M9"B_('2$-1VU
P[-ZK5+!_#8E;KUXK)=8B QEF KA>0&GEO*EG*UXZ3:]J(H-\*%Y':3G+@N//&\"5
P]M4R#$DL;;>(+T&K8TQ<TE=1V'=@Q3":68V8N_D05A1K&1CE3!<;CVZHYF2@=05\
P.M4E 4[4-ADG^LBV1#WZC^.GC5GG28<I;J/8 +/\";^&>7O3SU9*.A>(<Z0.X2YG
P9/:-P.E,<S4[66+WE7.%,C*D CW15Y>(D<XU2)DB*7(B,0+P^"8NT3E'B:M4F"/'
PFH2C 0?)@3EROAS/&#:5EGD"L4'CZ%_=_XWNCZ!UM! 5*#UTZ.! +*A79K ZK*!Z
P5QW6V8VOF^%4^PI>@-!PX\RR+MLD\Y>R:_\L1L_%.$9OL3*YC 1+W/ ]C2$NO$RE
P-#:A0!EF ?DV[P*;MG,K%&E1N)Y_;OZ8<6*56[,PRZI*Y[M'RO$VG&PZ;0$N1"#R
P4/-"\,OFYP13TW-]8J'SRW)[EW^ NB&IGY.?YE68(AU 3JK?W;]NVJ,S^</3FT-!
PJ.18(RF*%&B-2J.[?7EA/=8:@V=J7Q+8=@80M*E3.U..-(J!!Q<F4.W:B)%'Q.QD
PPTE.KX,UV=L"S3 6O.,)\F^[H]=.J.+%&NX4HT,[OG]]4T\<6.0267/Z&[G7!TI:
PEW-<JCU7U[H8\592)HZ/,\+(2:975U9@8/3R<.EB.R8P342;>7U7\]+=FM$IR:62
P52-@J$%@H8ZN3LQY\-XVY:L#!VCQ)@S'6SL#.Q0\,0C+-=-G<:N)S/-$)DO+=7QF
PR8"RL09 N2HZL#^\WNXJ)S?'&E6=-M-HK#=-\UA7Q:'F)FBPI.X$PO!^^]_E8[JX
PS(N7Z+XJ9&3)L:Z'XME.?:O<]/!,,6$%CH\V#.#;1=N(5K]2<DH9?>93P?!2V96>
PBX5,9T8SH)_6D^ZVF#QV]>)/L06-:G;0FE%L9M#>,;I(,HHI']*H!>-"#)&IT.NY
P:")=\W\HYNW[( O>DSL4U_&,S/2[^&3F,XG+;KGC6\:[7LMG V^D'H7<LF:BY-K,
PW])^^DWCXC:ZY,(4]:0A$!H*""QO-9)EGIU6J.L)PE\"*)8$7S33U32<@4:&&V;G
PNFU"$8G#@?%R,$CZ7(X4.M/8@)40D&08)ZI>&]L8541../ <@'A*[P(,&EF-;C;D
P>C&ESLU<_(F81(-.?^URZ8I8C-Y >]]T\SE8N4S<?X:SUT.@K0E1W0I1T6O1+!W'
PM=X=W@%, 8CG,2 [0!G&_M@QW_$-*H4K,ED,#?:3E)W8+<GS(3\T_.#&EA?=I>#T
P9W*V??O^7V%.^^0AD'Z2[R0XIXPD7@:?SYM#&?^I$QC_\SVOV]*K%KL8WG=VA$^N
PE$SQ3;ZVYZ"F/BWR3]E<2A-LL^%(;UB_F^'\1(=P<L_SS>C1[K' GMZ'%!0<6_VX
PWN:QAQ(&JAM5WXLAK: G5:M=_>(?WK(3[.ZH@/LFX0-GRP=8G-0.T4'3[#Z^Z":L
P3 L)ICI\6R3R(?Q3G6<294O>IR7&V'$O];7\\*L$=LBR=,\/<;ZT*(['\*M[QZ).
P=%=A<QGEQ<@VFT2BU:2S5_O>#^Q60H#-_[+XP2K+I!_G8^.S0@;?LRH4@Z4YBFZ5
P#M3"+"N?'-<+E!I/\=XA T=P&AU.SS&!M[:13[%LWK(2XW1TX$=B3-;'UF/T-WLM
PRU<SZ167FJNMP 4S%I>PVF7.'?*$(_HU>@58FX3S,CS7TU7<OE0W;.%V622;V5)K
PC>GVI(43[7&YQW,73 "LY=UK=*&36U41U?71WSQ/_;U'&:U;/7MYM7?@$5 9D>C[
P!(ET,H3DNIB8]=*3PL_1>C@"4NEL%-V#@ZOXHP<N9X,P:Z%F[931SA2AK>'(?/V-
P=9QDL?KP[.]JRX=)#ND&<"H9Y'A';:9[TI-TR#4X^%F(+U+\H-ZRM,KA"Y3,&NOT
P:V'@[IW8$%C)B4PN)I>HA?+5HX178\ZDK89']3,Z8RGF_V^]$(V"8KVGUBY1+,(D
P+NF>KE'KPX."6.M9IL6_T7=Z2K*:>6W$G(QA.18P)*:305=Y'HF:CV7M&\+ JN&C
P9EI.,T//9%E'L-'94+!>,7!6MP1@ZG;!F.V7F[K4JNZ;")\K4.1/,12?:KV9YTTN
P[V*U/Y7A\47BRUS1UJW#3IS:#C<=,*J'*T/+!$L'&D;0UP>:O439\<2U)$H&1I!O
P<IRAHD18GH<3982LNR[4WHPCOS@X^;K\+IWOZFP2=;ZX P]LV7Y3HTD=M!0Z_F/4
P@9D\&*B7H_CP>*4@HD'!1_TM6??\19P)65/OOW(#Z24MW32C72 *L-9-IM03/3U?
P8_% W(\[N^';N1$LW-/C<IS+1(DX(ZWOYL_:8$O!3O=DX%8(U^MQSC$VX!BI!? I
PWF."A+<=P)&S*U#WE.S*E)%SEFH;$ZONEEC\7+4DXX,(,ED9+%#MU:O;,N#,_7E(
P:^M^2A@<U(RQV83<,N+?+3@L?Y=$,R>JN-?_2RB4>A/U,[AFCC]>I<M(K^6)M#4"
PJAP-/9(4ZNY%2*Z[K<79#(PI"_5_/:<*[/6C OI9SP;0BDJ='-]!!Z@"+J9-SD>Z
PKN^YMI2U+V*A!CTT.4P"PVYD30$Q-#A _(3A,:_L0*/1?YB5OD$5$:OZJ2PZF^P1
P;MW&,OE>.L=T!:T4%<O%HK98]BR>G9S/AR> !#'LB9?A(U2E,#R:QF;E1UIY?V+B
PX9B>>9#Z<6*HFRICBX\L4@NKR:IZ_'+$U)V-ZT$9#XH ZPBU"GZ(O!01\AKR;DL;
PB%9"]H)BY,[6]AZCXA&@TSR*-"%  E&NT3HD_-6%=3M1*CR:=E'D:D2P/9-O9^M9
P+4<4J3G7S!!VG0Q,3:Q'*, J/Z@N+/PNQXKNQ9SD@I^R1N@9EH8L06:=W:@O@=J]
PA3U'U956*9C0V%B+<=F[5<OFSV'80DX5P:D@MIT,QHA/]**;5;<+PTZQ3S+DC1\G
PQLPC:=O9Z0HC<I5NX+4[7Y1$5@G3<#B6-I()V>ES0D 7K2]':^=4Q*(W5H$:@@\F
P//LG=.7,(AH/YI'KDE"7*D8:/N@#0 2:1H)TF,XM^:*:52_D;@^X/R0+9EJZ4+@%
PIZ(X)GB>E&5[/A3.&==:S:OR!HJUI1$=MI,6&SKJFJ<TEJ7]K?X+6OT;Z%4BU/^P
PZ9MQ%BNP^[.#"YKM@4F]UFP^9&&5]VF,@!GF2)%6[#$*62UD*\ +OO+2%Y["$1B7
PAVLEG/H(0_MAH52^$>9%2N!;2L5"B@E7F732)A-S:0MQLD;4"[E,S C<3.]]V(A]
P&_PR'V +&@^W.A'=/'U(H3&W:]B/$2I2DAL_C/CV!4XZX]ML@)-;-)^0T86"IUK4
P:!/93XOF5WBYRXE,GP2186C$ INL;"Q!(X6Q:Q?+S$)KSC_)H_Y=2J0(Q9D]E9?)
P/)K]G%+X?34/UTNH[/YI;J4K74V6U.?JK)!G^44O!NX/VN862WILKI/%Z$@&>>!]
P5Y3[ 0%,QY]CQP/N8XEMZ]A"7!M@\CDTG%)C.!)L;<X'F"K'<AB$L?[V( %E(W K
PO]"? \9MP\H0>&GWMO:D'Y(-G^V"%(&*&5*!E4ZB1,EX%O[^P;^  X>-. :9#'.I
P;784(9.#62L#^[ U$"-J)2 1D&70ZX"J7?.!AD]I&X]X8=UY6^>D$/U_+[8DNUE.
PA^SC#.$-.Z&3FJ4$]!DC\00_'IW4Z&@>IXE*NW3._-=:D8J:&,)V^UZ/2O?*;73H
P^'9GP-N9#Y*+K3EKAE'LQ TO875I:'<=:GVV".?F#LGQD]51;/]60.**1ISO)@DG
PW[JQ0!(%Y^CH#!=;)5 '/Y>LG\#3[XJ-(V$EAZGJV=<A(:&P*FTS:,#_UP+9R4!4
P/84$38$_%[XWD6TR,>I*482EJB[4BWUH(,B++UO)>[U0_R<13',^?@OU@\$\I<R=
P?)%%&R?OFK4*WSJ\REO*O5,HB;?Z,$H#6&/R66M3Q#D@9\9$5]M9HZ+2^M*257G[
P//T#1S_$(P> $ =A0X?.>RYH=D_@Y(%#/$[1M'-DSD(U8#X X8_K"_5+]7N=?M:W
P>*O/*XHM(,=.-&5>%3FXJ*?Q\RC&1L:RP-!,!_&_EA-0;8#D^HGO51D/JFV*KC0C
P2&;(2&"Q0R=.V%:]%AV.7I9\V%/G4<E$-"7UC@AU;Y"-"B:P2DXN;CK+=XT-#]!&
PF&D 2]V9ORFV.=AHV6KMT!Y\@D#8DFGF2 XH>-,+F+N&4'&N$X$]>.?RFC'=NYKT
PH)N60'F-UKQTBCJA8&+!Y90?^;A^BC3TF/M/W,=;/X)D".0&<RQ&*-9LBBO2@4N&
P+T& '!^9!L[%+"FJ!0"96EBG< -Y?A3429Z'MF^4-#2S0O8D@ _$OQ6_K.4%3S+8
PU]$B*?@JS\07 0.B<0B@_9.!</\$BUW ?SOCVU24ZQ%/UOG )!(CSVJP]L"X'SA.
PD:U_EG>_ZX9:D:C7=W(Q&+E')4MUGAM?R1"Y#EUWK648B,5OZ\'''M]1]G[C=/H:
P?WZQKTH93/ Y 0R..H]*@87#00>F_$]O2 7O\]4H(&NZQIO[GC=;B+'":^]<&NAE
PA# "Q$U1U5W$MWBT6@NU" FUW4"VRZ /_3S?(O/ )26:.1Q7AV^O]!+H'E580G\M
P:Y,J\!2"AH9E:;-G%!M)WK[!HI8T*:AMEQ\0@C)- ^%%$6Y;![L.+%==9?'S>^0"
P\S!_6SPWJUO<,F#.T2G;/DS2B.F71>.K/+L9 M5/3U3GW*P..2%+"*^K-\+N@5!Q
P^6JBKP'9(K,0D L?,@AL.SVUKMH\0,GO3CB_[ >6[[.(QV']$7=2X@\O44[KF  &
PB)J:O43QK\EKY( +.0MSM-SY5)=++^>1L")LM7V#!QWZHY3OUG_;3AV^L9R($FS;
PE4M57UR*P_@>66]!>G7=SY+W:2Q@QJ\!9Y+\!03-KZ%?*I]R% M*/[+;?QER/3!<
P5BG0D^?XMV; ZMRID,1AN]S$CWE&L;;+.FQ67"MSB1-S#Q NDS)3UY[>(M%4ZW9U
PL,Q=ZHF%#B5QD4_@7[#M<HM+D>E4RPHT/G4OKK?K4#3R2]85Z_4(I,X2^*=MBX8Y
P.';D[WUK#DZ=<II1,#WBWOEFS4/5KVA?M_.SK!Y>,YR57.BL]0AD 5@/2([@\'\K
P''W-C*\-*1<JS?E[MGB]\:]4#9D]6"1A152]+!2V\8V+_L0UO2"0&C+-I#KZ1*T:
P!!6Y.126KI--,C;EI6CR?Z+<R/S1SR240!S:3KT>11!ISSX]9>/&;+4)-$8C&1KH
PT:4;CX&7&TA6XBN@^)L)HI3-!#Q>K 1?RK/E86M:-I@J FOHJ]G!>P73.M7Y1,'#
P>5BF/3=:>"+:)\:83UV>,)5](9RZ]).Y2.D]2_9WP".TB/0SX'DJ["5P$L8D[H\J
P>,CHRD*MK.2$X?>0;-BO#]+;!?>$G^6-[45J144D;F"]JGG9N:C0<)[];4 D;86(
PFCN/ *V;8A!B;Z?798?#UM898O25^=X91^1!G!(TQ'18*>?3?GC)GPW1A#QO;1N0
P#_,TKA6JH&E'\8BIC).-9YCE.(&GKHXB7%+]M74#PC6/>^Y7Q1&Y;\;&R?$TR%Z;
P\ ^T756\9U:0C^@E,$%RN-UDT0:A1$.XF'VRBD(GWD<4I'R7;0.^J*3_*[^1'? Y
PH?;P+QQEUJ.%6-P;"2B0]^P2*\2#R=M6M"FSJ8;>@1Q:4WVVL.&)I._Q0;TIO>1H
PZH>U\ZN'FS1P=@#\U#)G"=47=>;%<40 ]:OEH$/\9-9Y4HQ<4N"),03VWJ(=8V_?
PV<)K\^A?33>>IE_31AGE"PL.5TW49P:"*-2'=\_44$=>EN0(;4@-M5@@NA5VSRD'
P+MJI58&CG#KQ"SDXP*EZ8A@8SBXN;@0=)!^ 9\IQX5A"1=/W!J*U?X=Q86<$3OL?
PIW7"3]>VT+T>[WZR40P8<N]P9JF2CK$S>G3-V+B9'7VH1528K<WL@T17GI[WQ:K&
P>^R;A\!"JP;N+IZ;X\NCB0UKIE2_XV>F:>!:'[1-A%#Z.R-PIE#]T(L;,M>J5P[$
PH9PWHB@5IS=K7[2V.35/6_\4F%V3[H%-LG  901LBX6VO<N@H690@I%'RZZB9&ZI
PYGOZ1Q:N.R$OP)M5;!T%#U<Y:QJ%8=Y*].X(FOG4+1QVCN*:=P-%U&V?(A1'0C&B
PSJZ*=M8J>2NZ$BC*ZJ+J"+I>Y-%/!-P*2&<"@#U@QK6S6XA!TYUQQ R0=.S9,//7
P>,/>[PI(R3]GF940YGVH/98CLCFSE^AAKR?ZOS PX!];/KX!J'+.,6"&CM<71QF!
PG&@I11=+,,*<9.@V+1N6'<I>JR@4<:>4)EPD)(>T& Z-%^]:AGPC!JR;0OJ"&>QL
PF MQJ*$]1(-IQ%'A2 1R'4VZ0H_6JD-VZV8\.[J42<J8BC@SKC&A8C[G&C_^-J$Z
P>-W/0$=3)NWS>*86ANRR#1IZ'#_RB]NA=)42E.CC/QI<'90@&DUVADP:;SK )3,;
P^=IIY*^@\F4 _]-P7)#O=8Z _.0\=#_#M8W9Q?+D+8-*91L_YV'38KO,?=K0E4(6
P@5523R'L/QT\_3]U#^*R/.MMAJH6?MM)\=Y3DQ;6(3]W$ATX>B4E'==LCZW$4O3Z
PUQ(<XG-P<F/X )#SV]SR#-KV=?](%\G!4 D9*WP\GDRD:F(O63%[-X^UX.VSQ6#:
PA/S5<BGV8Q,I6A:4']-A^I:H7G[.Z:XP1TWF^6DE>7&(AH6,(=A\@17-+A_@>6%@
P ;I;8?2R'574L12%?NGAYNJ;:/VT_ O?B97F&U%779P*<HS K0..8'R3)F?)[$/X
P0KTH)O0 E?M& GT8X&;Y0OVK37V9 JLEQ$HQH1_G$I'C:B+/LR6$^U782L]/Z&DI
P@N_-8IU/5T)"A;WL0 [VJ5YMA%81.2O4^&!F!8Z'+:6569Q&=V&*R)T"65 .#V0V
P5< ,645F?[PO\FA14]I&S0,/",+,\I#1#/V^ !C2N.3:;LZ*JA1QS#$WI]GQ/M?8
P)YA(6* "):5FZ)X_[6"7N BSU7N#::]6#U2)5&F#Z?=@+=EV*-";K>A118MUOT@+
P!.[J^XZA\7G5P3348<2X G!N6?1.AOE4D[<F/HO:E119?2E!8M"I>9Q;@3.TEVQN
PMQ@^5^<==$:4[79\,T!NT@\W71^[U\<H9$M;IT,^$@^[R/U!-4:^4(6]7VXP 83#
PA$15HV!#) C8G%:_O]X^@HZCR(I\QEL%@:8;)[KLKF=^U+5ES4W2DM_>WQR>)33;
P68ND**B,_+@)(]:9;G<SX.HG@O+FO,:Z8I3MC(Q_O$VRQQK^L6J$UB91TR@C7,N9
P_N8MEDW Q.LSU0"UK!9DQMUV<!)#0,=:$/FXA53K0.D54%T(QH4I1*23#IEG;EKJ
P^J^9Q5BASIC6F+!#L+2P^[),+A^Y7\<=Y7,@9AM^65_<SAGP[_M3[UIQ9QV<9O@[
P4&6$N=AG5]C/#Y(>.@V;76#K#"'_ZO5KF%.#@'@Y13-1.8+/Y<Y#VUSSN?!,4YA&
PLX:;5T!UFJYH'RJ+'")O0DZC,;&;<?CT=]BIGLH11,OK<4 S]?\OG!NBQ0,Z(@0_
P$Q"F07M: DH)HV,Y3N?N\W2FNU7B]KD3 :5?]_6UKN>P\S^M=N&K$6'\[#M'N8SX
PV7AO[?WSL,>EHIP_K*X?ET%K*L&]LH7J-E]0*\@+&@S#01K]3&5JQURX:*D&RI+C
PF(Y& 4J1K,[,HJ;\CO@PEI73ZZM@W;/D8N^>+%LHM7V:?&&B6\RB]1(H1@[6"F&M
P!/4Y)8ZZ0I-?6W5W31D4:_3-I'T_(^25I+"T);JG'QK[98-)1C&A8/AD[&Y1)$CZ
P; %G+T>P'Z'^%NG"+](7A.LPMFN47^S8 #.$7_W/0?SQ!*F.E.>.Q_IB\[,SB::F
P+0CCFHW<\5<>;W]=;F )GL"?3RR&(BED7'C(XO[@%@Y<*LN,@['!P..?3)D:%,++
PR$3:'99Z7>L=^&9A*0@VZ4Q25PUE_'S'94<I_GH+J^\OL3]3(4'=^,()KOZ#$O%)
P-%-B?^;/3G%W+L=T<%(+YG6-MOY92L'!"#X=!085 IG$!DSDJF1V'=K,:7_QSKII
P4O]%A:! ,A32?;4NV&;Q"%NO7<08PID%0HO_0T%"Q6()@TP$%<L],G/#8VL6Q*]=
P02G]1*TX89D^1-5I&; &7'83(-OP+1L!J&.67NO(H-WITBZM&4:2A\XO2UD/'TN$
P.P#D330EF9NOTR)M@R(=Y"G/+<IDR\T8X=<97*Q03Z3)(:-K>W8,L1 Q..T%'G"2
PJU5S;U\&PEUFL_V=.Q0TGE4N ] F<[;#HG38+R0'\-\4-)[;^#Q(:06I/.U@.>FX
P*'H5RMPN+>S\[:VH91[64U5T202U6#NZ[++_J"%J@<7D\G450L3N#WS0<F_WPJ4M
PA>A]&@3,X,BNN=$DT,4O%E-<1B"5MRWNA? <$ESLU*T*79=SCYSTO(9$%B]5DWEN
P6Z/2S.#2<Q3JB#4RFD%"^O9'"(85<T?Z?#@.E'L )G03F'@@?.[MYHFVS4R>L'L0
P15MW"!+\KUP<Q?0Y962[F =<'<MICT*=C^[#.O^JIZFQT 8:&+>3]24S;.$VN5R$
P5<]$SX*+>E#0X<B5SQZ4@/(;AQCH^(IH-)73#D.<>IN][OCQ=IGTJY33X;'0#>T#
PQ!Q-PQ77Q.FCZW2DRT=+Q2>V2 [1C.A#=)LG>3F.N2%.@ H4>IZN+G:>J2>9B2#K
POM^5D+\8>/0:G8TE\I ^0@O-$Q9<%V/<=:2R9;6:E8R"YJR:+\+(,GW]-L*"Z^N5
P BN$BV*HS!.A-+1MKH5E*@(^5F&T5&0WTK6C/07WF>6YI!^OW&WT6%Q>OW ? 3OX
P>#&K'K%*-B1@V@+7?$.NS1>!8UHQBV(7K@5RM^C^1H&W\?Y](,PULO'JA9@B8^$J
PT^G /V+B#WDNOA/B8-_19R?1?L>X,4CZYVF8G":^8P[ ZT->$5R6U 72+[*F&1:]
PV8=]KNM@W5YX \OLBP;6H[_N.(6!Z\;_"A&0PZI('@77Y+^R=+(9VK[(I*)Z+5'\
P7^_?,N=:0UQN+@@+KUK$3^&C!=WS^#9E .BHWY-YK%*OMLV'&)!B+.LSH5P5VBC5
PDLSR:F4XRP;SXMX[] 5=;SY-[W]ILU]PB-(LU";2M\#+H?[D#1#S3(=0(+CIC,.7
P)<*WJU>Z]/6<1^1_O-EEN.8:)XH018NEVN:DZW^MT PY8 8+/R=G88V](9M.7:3>
PLKF9_EE@<'G@,QY^ME<4,YA/T![%]#[KF%&;83:)MJ]2,I['_,RCQ@8.@ C(?!]A
PTPAOQD%11O@PEHV& ,T!Y0VVT1QEG*MG792Z@>Q3P>Z<*3/8>Q;]5MHM?E[/QHQM
P]R=^$J?"699%-*H3JW2@TP.U>[W^. []IQ2A)2T^]:Z"6)I*CNVJ[XSSD4LMIT__
P6]N^!&H])Y*F4]L_^N)B3DU.5HU$RP==SIX<4I\*DC2>YB)R<UZ]6!,%IS]-6.+@
P4(\\LW^^*[9A]1M;I1G&6R.37\W6,:") VA[U$3%DIMFM/;VXSQ85 <O_JA$R:L[
PF M^["16P>\FB\DI2(!^\#_$!'INJ'(A3C\[5Y\-?UDVX<&M0Q&@K23JISUJ#Y%L
P@8:,JAMHYK.1=OVH_$#W9Y]4X%OUS?\)8;T<&<7E[C(_$7YXM%[]<9C[@!VI-D#%
P+AT$9YO9W'!X:?H0)(+S;"'>@[N\I$\F,E0UO)LR?\PRJ=8P>Z"3G UG=0WUG6<$
P3J92@5,512"<#W1[<Z7S]DT7T'PD,&Q@UW*>*D!^"@3Z!%N]:KPYLT?!QM;-2&BL
PTPOMST0["()<=W<^#T?ST'-1SX__+4G>7MW67&-W<Y\)2Y4<( @'I&[Q^XCP9B$<
PWH[GXPJ.Z@JG%E=_AC9@UQ?-+J'$E*#W#UR$ )%SO+9>SJO8F_BPG=5I?WNFFC-0
PXG;8YI!-#>O5MY\PS+A[8ZY!@VMGR_SH*!6B1#-E8CLA@ W/V\T/TZ#-\[_&[2#5
PV.YQCY(8-?$7MZQS%: 8; B4NQ->@ K6<5M*H@>2MB*\1O.Z,)MCT6=@WA0=_6HW
PH.R];V31SRS>URB&E7-:%A)=R\OO%QX8VN*EXR/UE]C]]ANJHNQ/C'B141X(0PRZ
P_0_K!$RX&4H?@<I9ZZ\9]5.Y5YZ&JUL7SJSH-EE$5:^"%Y) B5)U/IBWKC,>XJH9
PQK?@O+.:8'G/)"5^W\>Q,O45LN(B^_#VX-2:GDGL.-1>H/'OK.4U+RH^_W4)S'13
PA[-I15E*E@#I-L+8RQ!GX4P-\QPE![$;$\3>$(%S9+/4JAG!A?:C52#%92GSHFMA
P0=./525[<8;.O:M"@G<' 0G:6N#;_BT?SV(75[>O?(^L(>99^(=V!W48PLO<J-S]
P36KLX><,KR,=Z['-/;_WU"Z=X<8F@52Z?J2C21&1V?660)A(3M^8T7%\'R&"++ ^
PSQ$2N%\[<4DY*ZJ9D!#'^2"'2L%8".TNL,=[*5J\)R=-90Q(E5^851#GF?OWK)SS
P:-<$>3?&>.PO*$3BR]B4RK1O <G?K#@C0Q)( $F%FUK\#S!1NVX*P)[\!0F4C*H@
P#Y"GC5PRY3"^^.A'?SE.!7=L3D^,Z2QZ]D22 T4@1XBNDS^AEI[=BK^9-WX>HS"B
PPS>U("&_4?5^#QY9N6J1JSWCRY(J6)^$S<-BT[^\;?JM)[3,6*SMX\D5S,B;2@^D
P<MW]79>OA&CLIE0B-8M3:HBI(4O6X<.^O ^:*)[2M):-6G2CH)[%S1.76*+=]F(?
PT.91?WK@',Y&5]BJ_^X F^I+!)-$1;/K:SX8\@W*Z+KD1-\P6_Z]3(.VKH)#19\0
P%6M8]O$G!DR'7H>6:LD"#3:!82UXH;0.,-^,*CA-T%K&)Q<-YM2#.W,%LOM[.$>!
P2#A^0 /DG8UII>%)L?QZ<XI?*$P)-'G9X&)&QS2DB+D#?%;JY\*B,G-8\**%;%1S
P:8^=#+71;HF ,T-'O+@F@8X+=VH/H!8M?7B;FZ3 A8)J$,W)+SV+K=^\JJNYK!_]
PSMLXH!I*@M*TS%TP92),4BS++Q)<C!'_;2>[MI#1*"SY@RPC.@\ DMY<#IOB)RL,
PI2]W%PB_:8 Z>ZD<)M/Q:+H<&.MOFI),A8N(K7Z^Y0P)*:33 5QJSCF&W0+]XXNV
P-M;B%2WBC ]C4#^>J,XWH';]KC(8@T.FQTZ?T>TN2$B4=V(#B<8GH=Q%F[;!0P.4
P'$F7^:_G!5Q'+YZKE,4N F*]A*-VH 5)6FIIL<$:$>E8SG!M.!;^X5L?:BX3G(N0
P^N8%A=T'I#F1VP2^8/(7_MH HE=R2$,!<00@A9H_74A"MX.7#G6N^[UD]8P-8FB 
PAH6'#W:;#X4G:W<J>FB+3 P.W^,EW"K?!5#9CD0CWNWE(MCS [_CW&=Y4J(T*J7;
P9]>HN!64_.4481>!25FPRJ7 $>QM;O*8P*[&YK%,PGR>/5#8;% PO%\X"HDMDG;N
PC4F4]I,)-:^A_P99UD_'F6C+.(OXR)&#R'4RJB,FK&(Q@.H@7$MM-F$.WT%SGML]
P&(@;T6CE":)"1K.3!"P#'YVF^R_JX7]XQID,#IMS%:+F1QH""0?F?/[R\E-B9/43
P'6PKJ1-A5J$E'L*2E*X&K\S%DF&]8"0(;]R?]Y:@#6F8,[K,N8%]=]\Z#X^?RR<^
PN8=43==\9TT"(]#M.Y4A;C9Z._ ?,,+9Q-/HQQDV'\?6AUD5V-0MZ5M:;5?@1\C&
PUZG:SC,@5+4*^4XLKJ8EDZ@,*\FQ9@A*UW16-,TAJYBY4/;K73<@?/0Z(9(7>.*D
P)T=B-F">O9OK1@$C!X<-Q(F1Y;>T3R5Y!!DR(V\*'&]F\3UHT/&,$<?;CC?.O:/1
P(&:@>W^5L%KB?3!$$[X4^5I(;+U/V?CE>*/BC>14O\M)S^1I<#(M$_65KG% 6<ID
PZ5Y[ =81A"P!XVBY07"L?I--^F!W;>T:BM!A:KAS74(7K;%\W <.;(?M02=CR-6Q
P#Z*D0B@).[%<!\"S^>5V6%I,FB4CH;X6[VJ.NRDC!5I@Q119?&@C^9V.V@"1P"=M
PJB>B29VNO/R0NP&OV(/"A/HJ.3BS3GE_#YY!W-TAO4Q9ENB2,O-4 &YN84Z\@$M=
P?\P..L!@5!5D^LM6I=C''W2%\[UL56UM<TY><CS^/+@$I0.L(>),>N?MQAN&=5BK
PCI%A^5+L],J41TV<'>4&C-(5;/I^C^W5&Q8_X<#A4DC$+?:O,P=-6/KUL<[P/[:<
P4!B*2<_)\9$4$)=%A8H:2GBJ%>_H:IDZ4A^/^:Q!EE1Z-O["4WC*2C7#ELXF!)>3
PE.TEF6B=\F\HR7 73/_P]6(XK4*,Q)%8"W7-R\;;;)/2:64^]-'^+)@P@)'(1OH5
PO-W'8VE[[MF>[2^P%@HS<,O ]KKL!?7=,*]L+-F:H$S5X'.@<+#]LH8Z\_Q3.4\[
PT,@K=TNVJU4D,='V:C-Y$@1EO1V>NV,Z*Y+L6(#+VM;[SSK1O+E)8A86DJ,V=;E%
PR4D",Z4-K1Q?^[-S?+GV]]+Q_H-2K@ V98]5-&6KG72=W]@Z+3VAO]W< "6$N:,.
P7V,Y;A&D<M<.U(26/0*(7+&$N(<KS\0+!/U!7WI*L<HB/4DE#QN_\T%;J<IW]95W
P+<KG[7::.@(E- >L+E_5N"C,HTXE],SD_7$T-XVDI[I!A&F-P'%Q=2W _A@%*NW)
P*O/W S1XH[H5&PE#I4*:%]NB"UCLL+"K'?(,U8!*/&NH%/=S2_YTM+!#PG6E6K J
PYE_0<E^!(G7L!MJ(SV5W\OOCJ_9.9'-@ @.S5;7W&K*X(?"O+$L$0[51(;H(L*2I
P5H^8=(;;H33MRRL9IK8Y?=QF&J'3-".1786OF&N5V?Q]'\,0UV>Z ZICD3&K_-:^
PX2L,HCOT][&85"G51Z&I7B?)K3* V)<_4(2"EW[@F[.A(4(C7;I1E0PQ3'DV/YI2
P C1G-1_"--D&DFBC.;J'@NAX;QMMHNUZ.P0Z?5:O-(ED)EJ-4:VX1-!LPF%1-+5N
P#5+[WY/330Y&'1AY +H\LR#4,6G?NZ;!#7%1IL<^ELL('MHZ"96/OJ6:=8YJ^X$I
P5R1 0LKP]].& \E\_%[V[Y8-2P';"?MDSY<D6H1Z:7N*!Y6$O;'+4OVLD3J$>< &
PYE#DJ0=&O'5.[BJ.B66<[*3_<3[!)\'R\V6H\G>]!N>>82'9@/*=*A[AY1] '?QJ
PBR^;G*?8<D+=5G"UG.PH,E0-^3NS)Q3 2FB55E<IRX).FZFT2:2+0NN5#G!>J $>
PF>ZE?B+\B5=#8:2UI0+G#7.1 #W,:A"33K?/K0X0*S&,C0;WD?G _68ZPE#^.MS8
P"<[9MQ<E0=Q4TWK;C#:C8.A'AVIT[,C:F/A'F=*_>2PL@\S9% ""SX&WJ7:T^SVS
PDO*]-__[2W3N ?! JC[YJ>+Y)&H]^L&3I1:BFZST*C,.;4M\[7P%!%$T=8BK>>TI
PFF9^C'#,:C:;9@ZJ(WOC]G,-2@;V:C$LI7LI8<,\J4QI=K X$?R).(F!B]X"(OXF
PZ="28W[[7G'>"B5\%A><0RW^\0$SCEW#AL17ANR?Y0[2\Q7Z1.L2$:0NA-)GNFQM
POYL>#ST^\ X>3TE1- #PGTN";RP>:YO.ZH0@H2PSEV8TB/-8NLXWF7)E^5Y0,AE;
PJ'W"0?<252J.=_!7_[HO"6.FC@XF9%8[5O92:;MF'E^\]Y $0F8"*6\$,'^*Y&2G
P FNZI_$,XUEQRI@M^&YDA8R51KMG4QI\\E7=SA=%OJ6)>6#,7#NZ4DGM[S4_%4^+
P0%.58<G ><O(A?@J,(X6AL2W$2O/60@8GD)H3R/$QN:SXY0D&%,4;V4INYQGV8:H
PM0CVED4S:L%00FN(\Y?*V;U3WZ?D'0'++T*]Q*7(:(]\30C=UAJ>:G183^CNOYU1
P N($S86;>G>&/;B(.#/"+YFG[0@WDP@0HPA+*8%UTD+(1/5?O#8_WC0+ ?'-:]CG
P@W'Y=B1*=Y9_)6XP-<)6EI*33 %!^>'UM[GAV*U8ZE9>##\5SX+^^LO+1DB,(071
P;GHADO#!9P'R@P^K.(;<D#KAW7Y:E)$F,].OGB]V MV1,3%\0(/XJBD-P?08(M/&
PSF'G$\L'#1W83J4*J2<E.Z]MK^^;HB@^)9C;HH3BH3=->0$C5&;Q8@9\ ES9>/>E
PF]+ H-CFK$=%T0;K4;&XLCD-),!*L=W+Y$'<2TR*R:UC;A&\L.O!MG0WG)CALP(Z
PRZA994"B0Q'-.[V&9^_C>SR99)1?_Z>0FTQ57E%6J-8/H ?G%3]VU^&%9AA!\R?6
PW)'/Z'>OXP7A9F&T'3->.""Z2BYF.)/7ZE*BC".@LX%CC/[BQVHO_94 B_#EY5IK
P+5GDKE668^<N#M/VMG_<0'@[>?37BNH8A'W,0B3;N5EI*VZP*Z<=!KG]&6(2!P$E
PJ;O\87,-U[NB\0XD)T64X=/SW# #LI'P43:*$#>>A'5@77B+SE^G=^N-JFF4GXS3
P)B5I9IZ6W::\1IR[QG#_3WQ@L! PAXQJ:_TLNNK/65)W4UC*1RY[/Z&+ JMC7C^]
PO*";^_!_4ZY7#(8'X2V7V+8%V4! Z?J/>&[3THS0JY2=)=F!4-%XH+W\GK[(>>4(
P7N6HK,4BZ0P>D8GMP\2C/$/.+6-V.<K:QZ(6W-<G?R1)F0L%5HW>JA^QPN,O?G*O
PN[6'A6B5$#QQ<+UR0[A@NH8J/.ET%V_-0DM+V!VP&HK24&(+3]:PMJT&>R)! ?5G
PF]\=HC,-:7C.A()%.D9J*"QR0>V QR:FEV0E\PGDKO.7M;B.M_P1DF!/^MNPT]JB
PO73(1FQO8 *9R0TO%4RC!M4-@53[";+;.06)ULV:6W51!^%64^8P]0</^'ZXWC@>
P5$*U,3173W<STP#['5=V:&6BM]<Y!1KP-] EE&R#SO\D3)[!'JH@FHD5BW91(D34
PPH^)+1L[(?>Y?B'P5%<R42OGWW:+'<TRN[STZD3NNNQ7"DOY2WXFJSU6_GN4_T?+
P0VUF/ZRZAD5D*E#O0YH5?4[VFK/2]J0QYQ/I_T(*:=J%'39A?,F[@--E49-O0&3F
PZFX-M7^KY9FV$>)SU^>\CL!SQ6]BT+Y:> "CEFHF 8V_M86ZT)=)X!SL%?_!/_[8
PH=9C)X63&#%1L=05]'EDB;E%N/$;&R$\\I4WZ*HW(C_4J>M/6R*;QH ^"+<FS^Y&
PI2P.YT2E"($M@"WY ?')Z9 U:9-3>13+86E8T^KZH.W:$!@J;G1EGK;O;@K$%M;P
PG1,93*[(D0B=WE6Z>-K7.FM V\@K\/8XA+F6L,-T)B,V+Z7%A5 L$'24)L$*ZBRP
P7--,)GK!W_/MH]LQ$!4"C''UGBJ*X\M+HRXU7=G#&0JOS+E13PXUYAL\6IC*CB+C
P1R7?.[PK?[.4F8@J.8>]J0887''TV@6 X1:/T7&JO9:GHUCUA=MQ>S+.%A3E..EX
PK25*!>!:BCL8#N+6/ZP#8[IQS,CYJ#Z%>XTHYO ;K(7'8A.K78U=E03A^_%*NK0J
P[6Z6!U.[?RC'4?V3&HNNCR1.HL(!;YU@WFVWM,*L2B-PQ/NIBY'3LV,O7%X A>X4
P1Y[OC1HH%W^:;(\@YW3:*MC#TU]9<<'M-]R0&5:8JA>7LXCCQ[C!  68]Q;9YCGE
PE\X5OB_9@S %"$Y.FLSVY21L,K0(/?=1D)6/[HN?2B36XK+)]Y>3<CYX5=#&K:(Q
P)]TC9*-C;H'[AC]N=XHENLEH87_VEXVW<.TER[#)#B;A75 ^<VK7=_20!RE?O@<0
PZIGDS%N<[-8[/9O@R#0(&X, (.4M4Y.(!/;IF*>(VVZJ?YP\M?:^&"GY@4-Y"$%)
P+#/6^441+=\#7&)X'-;;RACC_YQBU=DZY&J1K=4;55X#)?AW*9Y&H0C$5 0R/]+J
PIF!N^BQHWA1U_H2QTB?J9 Y'-=!Q,^EI2#75#N58@+X+8"Y#$:U^YQM5Y!#R;EPT
P\-FE]DXH4E>S)O!SX+ZZ26.UY%Z.O,1[2-@55!S"' #)FZY-A208="274:H?S8HM
P]Q]'UJ8];G\J^PQ0/EREUOB(=H7BOPT>C@W[!3I['@WANDA\U"Z_+MXGZ;*:YMC 
P4Z;8I J.XVA9)V[%5QWC[B3SA<^0M,3R"Q:'DQ%GK31I!=5=S2[RFRKL:GODU<_V
PE+'K]+CUW@;\UG; :.O(X^.9<[ T/@UM,^V0XS''1.@>+L!/0?$AG0LWB-V>.0%=
PAF!(.V!KV[L3&:O![G8_<F8C!;K_K,^#?[;1&H'Y(63<]; ?XNLJEBG[YRUE3\'D
P&O3,0H9YYS-2T(406%D2E3$YW'4JH-[RRDOIF*WL?9%.\V*88L1;B$160%M82BCC
P?)Q8E;WKBO-% $A>02B[L=#N%&0""DU5=S4UE3IA%D$MU?O9"J=TLPPR&M[81-T$
P8J-@_9YF$ND!#]K,RV@+>8B&1WCV#\/M?B3VCX#+'C>(K)KOV<G_0E8G*7P<3&U_
P>AL\%FZ"X:&!MWE-YEB@^R/U6);B(@,Y>\[4J&(4S>6\E'CJ8A\?FEC $5^IZ!;[
P"S.'%^]3OS@HN(:_4AQYE#;.KG/'U-J(K;(%;6+B*@R398?7$(;>P=^7#!F9@$,#
PSN:"3!?;=+"*L9&/<09.=%"559Y$*[=H/MI>5:.)9VVDD;WAW(XXFO>C:XM))M.[
P(5$>"!?J$/WV"O.'I[)+"5:MP16#L<.&DF2T=P\-'L[<F/D2$L$3LD/C_64"]:J"
P+GN["U"LA:TMR22M+-OVE; IE;W; M.+;\UU ;)?5DN5Z^_=<8Y@:K<)0(P+9T>%
PVK( O M^N.<9>=TB--#U04K987L1GXX&!@VF=]>.IQ)4M<DNT;91YJHLNTO\PM\$
P=1%(&>'_B7RI$_"W#IYNU4 :3>D;S*X2J</!&1+7."(>Q A<7H]MH W[(4K7O396
P8S=?4Z^7_8\T=1-M,8PJ?8)#7T5G Q&[!"MX,/;/L5]N',!^P!&F?(BL,ZQR*$<N
P5[C8)CM2$0YEJ<$< M6KU!\UM,,N6:U<*S<(.@N%?\*$%^!AK<=AG46B225X@CXS
P;P/11_Y$CT@N4)(!N*61=(T91@-IJ;EV;K$K[_1!:6B ^OU>2?JTWW$FWF<3D9Y,
PY*V@#X2)(IWZC3!Y+KEW(E;6592KRV FLOW(JI0J8' 5R0";HXGH^OLU\<!23.Q-
P>XK$[U_Z6\!UA2OYU-IS5)PGN[7 S!RR]MP>@@' 6(R"O'I_WRA$F;VHOR=30BC[
PN6\)*XHT=U8&UF9+ZU7RGZ)HM=0%B?UYE>/2M]F>XBWG">R0LC$[05\LG-*_Y.5Q
P +!R'EH&()^JS+SBB@VV*!\PSG:QZ6X7F2YQCY>Q8K/L/C(K7#LQVM&;1A_B0GLK
P\I_/_W*6J\YFD7]I7Y*DEZ7&ZQZ5:NP/&0&.H<I=XY3BJQ7#>+P  $"K]E;NZ5C,
PGN(_T-=E8$X[P+_M!?(>-L A 6J-XQ+!+(L9H<D<>2CVY;$'6RIC> :[E/+E*NPX
P *:+'H2:A5H%R.LQ7#^&1&(_,'A")E8"]YXSO+@?VV3GL#!D?LU@1[;MV#I."@29
P/G_FG*6H/^&:Z0W= $7,>,. WWM(Z$R8KI/L-$P%C;:B_FJ%J@(D[#B?O)\V*6,I
P&;GZC0RT<&P5->-G-YLIC70'_I UD18C5Q;802\K"/(Z,]1:(E\+/$ AZ&5>)3B.
P!?.]P;OKHQBRLFBKI"R#5N=$G#8/ BY@E3W1@1V]$R'"<D3A0)94[VW[G3U\J@I:
P00%IM/ED$PR0X224=4&EI[3>327'&J+3M"%@A/S*7<?'BU7!W#DP49=3PC!3GITJ
P-E&)#B/./ 08DD842\:"]60#$(;$6U#2L52,BKOS6U [GBEFG<,=G>)(V,>OS:B2
P>PBJNT&#-+M*+!+FBQOC:HF>@:2D%5XHGLC2K@<>X]?7VA5J_L3R@Z#S N@2T7@G
PG[=_$95K?Y]]T;FX?:=<@F6'#EM-#!X)=Q>4K>CK^]/B.-9-V9POL/%%B</ H46G
P5)-Y<!>1&1!-.>#0)4XWO4F9^&OL\A\7TY";W*WPO-1.]^W (A[1^4,R,K:J+3[ 
P*-I8X_2DH^H+)!RL.DAHLCKJ*DF1DES7_T\NPBFV"$;N'ALI(>J#T[$[ CA?S  C
P%1,T=F(^:QCZ _?S8>/"1C6RIM 1'$Z.5$<8"AU:\IN.D3=?'U*7\+>.7TBE-"[2
P&:00!Z>:^+R]-C/#K_GW\'H_VRZ2D_91>7 ZGR"ZL1580E!(F4'QZN@DU0;6M0XV
PD9)&.^F^42 ZYE8Z^?B?- 7?N6-O#39E+L.T2I(3N/I'_Z:VAJ$1]7U'(2A^3L"N
P2AHY8DP0'X^=S=&&%=-MRHAN>S*PM6A#-U\#JA(2G]5=!]1K._;T0S>8+'ZYG=M"
P]#]3"=!LG.A36GZGZ"SSMW:I6^1)3O<\4>3K[BK"_4S/DUE98P:/_"@I/$ \21PX
P7/ U1(]:=Q#TCPK^K<>-PK.J'.N-KM@,D++ +8N1<Z>S[X(N"O*"-H.+[SUUL><O
P+9=85"AMK29Z/)-8:P@WV]@BWP26E@"<($0GC)9& $D)ZCH#YL@:3CBAN<MW^)OB
P%=BL<AN1XJCM?0 >P<J/#MM<<]UU7+\ 9JD8902_:K#&M9]F*NM!VX*]X[3UW@>[
PDO=IT]>9X]*Y?ELX7CADYJOAN^'(0F@Y=(,=L1J^EJ+/O=ZE[Y=#7+RA?_8I3F_W
P5DJ)S5^]@N:;]+*U:TMU@XB0KNNU<4)0KDK(!2X@,9F( C+;UN*I.Q5P&KK+'5?7
PEN%]L&$#A;O1R.;MP(NN@&X <4M(*P4D+[9$E;R)8)XFQ"PN!PR]>5P[)2V_^]SZ
PY:GS\^&]/9I/81=J<\TQGOW9S'_>RDE)/')+2J7PD:]%JC'7 ;@@<>+C]VY]6+0T
P_]B$9"CEWWTUZ'W: 6&?VC7-C7/T@(WAM^R,[J0M#X*&3*\]H@M,>/G^#M?GKXL/
PC@3M:-Q4^X?\C*FRM"*HB15=7S+ZK@K@1QM+>=4-A!T=SZD#\<KX #Y,00GHJ4=1
P=,)5U>Y[F2IC6H4[^&+/?-@GM;4W H9YJ5GZT]E+[>O1J I C*G+>RL3G*<ZQ%C9
P'J81_YSU.%A5"UMSL0X2)1+4[Q!/>\/5\$;L^M4N1N_/!D8:G?]?5IZT]E^!LRAX
P+1A(6ULT= L*7B#\+S-'V@U/-@A*SWIS"FAM$;B##NU1'CO2J*H_]QY4^_1S0ZM6
P;LO&0& RB!+VI/81%@)L-AS/7G-)SDJ[HC-'&EPTPVIY/8?F&.M PQ7G)3,[<,ZI
P9"L+XZ>9J[WM[/T\(R9\3+U*,SY>05XK_2OI#1>O_38RG9"MHT1OK@!$)U3SZ2X]
P!8WR%:\T4^F-?T!:0]ZQW-Q.N9\P3=\<%S]E2 \2:8_K3K-5BV2A>"4X.[ B.VSY
P#Z10\#H;02/KQY<.<E5NW-2IG@SNZAA<,8=*-#G3[[6#2#!.0!Z,A(>5_,'J_QK1
P+ZYH%]=S,I Z911R13S-D8"Y?9GJ6QVLFF(;.@#!B8VQ3HB'#ERU4 J^FJ%;!LY\
PH]V=D!CQUU(=QDMS1O)DBW4U^2]T&CII<Y#P1XW 0W7%/OK'R@L^H](I)2PF$R2V
P?8F[R1\DC"@/7#A+KV];"M3JO>$G&OXYXU7C[VA05_[3R RV/!F^>ZI&X-AJ.SN?
PSO\JS<=JG8+FE5U[DY8RX_=NE&JBINM32A%=!G"'85$J6P6;)HN7_(Q8P&H0_QH=
P^%)<_V"RU :E>%"VZF\C2),^OMJXH21&SOS54PYA9R\4GUO/&9%DP&^WCD_4=VR1
PZ8>BYIK^9)ILTE]-1/Q#YG>>(+RD))*_ H*9+B[KPY]45LS"%#A")AM&,0O-. CD
P/ 2:@7AR:WK^;(HH=&YT&$\[$NACIEF&'.WQW8A4W,2Z8JM%H!%W,'NDTG6DLB#N
PI9,%_<Q]_< SW/2HS5Z6)1P^4=0#(=O25B7[;1OA%5LQK4%L**++<[92S^21?= P
P/:MN-A/STC+*W_ .55+ONEL1&4$SY4RW5QV1\<6V$B]CT(1A>\S%76H6&Y&I+G\R
P1BX7.NMDK%SP:YQZ<%"6K<0)6S'PK3>5 0:6(5+C)"6=YOC2Q:B2E ^B1"&>Y7J]
P!R6#;Q?2[:U&>^]"N8<\:*0F)/7'*L6FQMX@?=8(<PS3#'UX+%2D'9#7>4$C'4KE
PIT;5W:[]@);MD37K+MRQ)PW8EFMA,(E!&_M;Q@>@$U&+]"Q>2:5!"TG_$[O+00I<
PJ_^,5-$>A]2^$!:_,2 $LT@66:@7F, O<^ Q4M7ORG;1D6?@EM-U4]A#"@SB0*< 
PM]<-%ZX.I[WCT'4]$L\"RZD*EO_+^'C\@(ZV!FAX:MQ>FS8-K"X5QER:L*J>F^6A
P^0H(=\Z^6Y#J0G,B7K9G0P.(GR.+!XN-D&IIB9_U2*13.'@'>*:N(8 =?H1.0I[%
P@0NTJ!UB;SG!HASM#7IM5+RA>R&0J"TC4=ES<&?X#V0:]6QN6/!_;G9'$B::Q<)I
PM%807-*)4">;F2 SU))<$@S$/*<QV\U\Z%:C/7-% 3:BL(X]M3@AAZO>8K,V;"MZ
PM)5"C:;K/2259!$\4!K,/OU.66+*0V= /G/E6Z8%E/P[C01J#;1;P/<*2-,^L-90
PK$J#7O!PU9"::81[+S39O\ACJSGXA0\9'4M=2[%.I,;M"#FM'95\4R!U^;YDM?"]
P*Z+@F1@4I;8M2"LI^,);\NW]U-3_K<9C^7:=E4?A9E;$)_"+!$A@<E)T0//:CGO2
PU^H2<@"$5*ZEA5 #40*-$FGU,)LI9\U\G8LIY)W &OBZU(>D=['F$?SJPJ,]IK\0
P4'2WM_B3H"8.XVL/JN<>L:0[";X8FP<W%>Y$3HM61\LYFU%9!3'XJ/?(RN=J6"_*
P ISOOCW[O_P94(!RIW7X!<]80*W[%Q%#&+!WS3PP/$9F!X1\N")_V:K+;"1C#)_3
POY]/3M[JJ=P2;4]MZ?HP*!^ZALGKP%R%MY(6CSE1,.\.80[,>M[_[>J_)P*!3Q[^
PP(SI^1/""M\1>(0@GLR/W;;]($?,NZ(?DI%^2"S,?=?.:T?@SR<$N5@7YVG7]A6_
P45^Q7!GZP3BUSVKYC; GSJOYLKLO/CO[UJ@CLWRH2IT+OM)QU52/=X$P^HTM:FND
PY4PM6_36&V.$..GL;![\!DF?4A<P*"M+AG#DG:EQG=;K?$J4HNPK82D]:.=>;:(A
PRRMHMX)AQ))E#_6&2+=%(7IGP0M2#^3B8 >=T(F_I8'S7X!A?K?T(0P:^>Y'R*SF
P@^TJ:P*B)ZP^A:>$?KB[9QQ?U[X[M/:2+RP*/ 0RFQQ*/-CR(%T]SHB[8;S^Y4'X
P+ZL"QZ'BIG-*,S7&<:A6%36LI_ZYO_THUD[]S6Q6DRFB2Q_%+)0^("%BC^&,*D'Z
PV7,[8/=U*Y<L0Y*@(?%UBC;F_+_B;V_]-!3E^Q8EV\G3R(.F7HESY5A).N\F+G !
P3NO@.>%BG1!WAUPEN'7QA]2DT"#$@-G*[!O/:]"MEED0[D.\:8@%9T9_"M=[B%&A
P\[S[$NS%7K35K5MW4$I(:/?N7DZ&\7 *Y15UO,])QJ>"*150V%JU#7=7 #^SW0=!
P]CFH+2AD/^H@__)_PJ/MO!UDO,3J*S>)$Z)8@0[:O::-)PLG/4%SGPA_)$=]D"OK
P_5/61E4G61P$1]M;Z_7IF3J_M/OH96Y3ZD$/VP/59+F)A"AD3+?8EG/V8U,=#V(.
PH2#! S]T/4],*@YB=[:J\<ENQU5C9H&)O5?"N"%)BFI4.GM:,>H YK%1@!C#*[ [
PO=(;] V?QR-SA7A._$31%BAT/LR@"&MHON%B4ZTITAX9(B3L0/VA!W*_M1:MZ/PY
P?RCNGWBG;H/,)FI0N2,O^Z3G<Q/$$UW=PM'VR]3N':ZZAU'R03J96]+-6REHIQ)U
P[M,$C@*^F"?I1 00Q-2U'CTG%U$:'+6%&MT#O<HWX17-0O/ O--BL4+<R<+2)TYV
P;=]T-N!(H+AA_$^+O I166_HN-[7BY\S43N-P<L*4)1F-DQN)E0E]>D!>*; 4M:3
P](+1MO]\=7*M/.69\4,' ';DI$K:N1*6"/1Q\]GUHZ+AK;2OFTRI.X%H1>L'2W&'
PFMDBR[.^O,Q^I299C_9F+AHKT+* L5 ZW)^;B%'2PM![618+07*:J>[;!?\<35[?
PL(QK KBQPK9QF:+CA%0:MG";5)1IQ\^6M:,@<;!V[]4HV%"U\Z*>VM"6,[5'_/$[
P9!?'L R47V+^1:FLY9,TFFR4I]T)%42EO2+7SDRNV)]WU^^730Q85# _BVS7,EY'
P-HKYK\_[@\:4ZBDVNJ&,*></IEHB[668]?RFY::CW*$A<Y%=F&&K!]!UI6N'3CBV
P/K?;FEU;F! E2VV@12%:VX]]DQ*"8"]*U/^:5@;@6?: O(E: UFFE9@PP6P2U(F,
P5N3PXCQ#^=O;W06#'=3H\6D'R6(_@<+@QD:+KK13M"?OW,V.R^4U2^HIV9+)9_'@
P\A%Q&F'%0*^SA/12% L!;0XPJE7[';JJ1/]0'--(;5'4SC/'-[F;?1#66I3?==IU
PVN*0Y,1V]F"^[0D;DQ.X1,Z&$T[=H1(== 45*]0T5M0N&L=8CBCU9DZ_BE@56;ZR
P,FEHJ[?50,XB+H]-+"A=[<*FGK>*F/X_F[Y1(TQ)Q!6\B7$N[OJ# $?A/1*MA_;$
PG0Z8'HJ*D'-Z6L<\TO8&DI<RG8@Z[6D5?[J3<J[ R)I/3%>%*SK?X<BR="_Q@P6^
PY[H7B.0@:@Q%1O"?\4HP.RYG4_\R*/'ZTP_Q\KWF1/&.(,K+.Q]+>#AY#S4OV.0;
PG@;+EPN5.*7R+"O08N^M]WA!/?<O4Q[O[SI_RT.4+>\,+A[_$C:*$>=7D5BC?>W#
POV^@F2#\+(I,6E,V-";6M%S)#FCU:G@R%5+R,!&Z9SE[S(>&L;UT9]'X3)O^JBFB
P<NL%T3I%[8@_)42[/Q%>B^?]J^3M.0RX!Y5VH<#C\/A?^;T(PFGNFA<KATAO)9(9
PZ_0QEQR9W_USI,U6F5X?9&>AETC95FAXMZZ!G%)3YGA^BDA\V%:ZIPO;N 3+UK??
PT3J(*5M4^$QZ0FYITH,=E;A?6HV?1 MLS5ZFM'13,!ZQ58I+&?!O<9;O!]JDR+?5
PYNDW0CV:_/WK?_]*3B)[4TVK1)U$U+4-]'F6M_ D!AW/!)_OSIWM/D^1J1'<XT'6
P]<CX*EA0C;@3!5GTI5$;,2<-)RIJ1DQ:V3E !45AIH$XER"'#>I[.'(!."KH=#5G
P(/!_CML9WROU?0%P#XP8LOX$YS E3I,Z M#PTL&CQ9!B=K8>Y\,2#/X6?.8OI,N-
P;7>[K7*E,M K%B#MKZZAXJCX0BJ0KW7[B%*W3CS*N2@-K3PFWH[:.="^"2J;U,!3
P$#CJIYW#1)2E-!C_>W)TE]@4NI[!EW:?+Z$Q$"-K#%LT5LOL*0Q+D\$AVIU6PW"/
PIJ>CODPA!:QL?]\*EZ! "(PNI !]K@*#:/1KHLA?!6 !ZU)E_XDE)J>+6!O8QY)#
P@ET<+6])0,(\;Y4]Z) 2VKW.RAW+P+EZ:W2/,+$;FLIIL"*RR,AA\"O%.I]4/F<>
P*0OC]6O0M@6;KQ%$VYGP>MIJ*ITL1 @/E;2O7$*BD?$S/C#[3@%+#.?]?XRDN0?=
P$243".[G,@V1]CL=(ZE,$JKP>Y*;'9L.;/=4[+@R3=< S3]$$122G+E]M;_@IAZ\
P0B21(E&A!7P4A;K^D.Y@V[>4USX>"O*D$6TBWCDH<U7\R(L,:6G-!G-429JM,-EC
P':4)0,*D5C>%KD1XB6J&W==9Y&7'9$$4Y.P14PS*3U/3LJXIG,QE+ 3]-W'/U./C
P=]<@]%I%7!(ZP[H</C:7$?W_.B(C#/$-78-VX/QM-9!0W,015R6;1)"W1NK:$=2M
PTZ*VO.?*92,A'WMI+G7[7"MSS#3<AVLGR[33<8DQW7G1W64^-%1--74]*G^2[L9)
P\[(WJ]9&79)Y-\E.W',*MF&+>NQ8RXBVZZ*.:N7O3 HT5G1_U+1<ZJ06'4CG'U+(
PTK%%W@:C^3LB] C][LMY7SB=V1G!:?5)$5OF-#Q%5U"$/G&VEH1ELSS@QI;R1M6]
P3,XK0X==\"@*7*$ X)Y;)LH)&9LVC+N3QR)8]W7FP%I O7^'?R0"6SX=,C+4W"I&
P:]V=^G8Z\CPO>T_!"[P/M";HM#@%Q8SU 5NJ0<[$54I$I&>2>@@%6FL2,PEP6[ZW
P5FM<)_!6Y'0[KN\(?O#X?^GP@EL@)0AJ?<_.=/=E>ZS3JQQ$^T>(0P<ZQ;\["'-=
PU-V(03IN@.(MC!:50*WI"V1,G%.X,3"'&\<\N>F0-<UUBN4<:J46(2ZMRY%R .T%
PY(5:$_*([J:RU'A-_]_T':?YL$)5#\&/O2HGB?Y[]-JTA'A"71(?UYZ45DN32_;2
P$2?$)@,Z6T&(K29RI)D92")-"&5^;O:!ZD? E]Z8\JRHM%P?$3D<E]C@55EOW6;=
PD5+-W=*VC\4F&,/(MS**<O5KN77@9QN(&UN-BZ5)-"PJHOSF[C7(DB'D3GA_-R)\
P%K9+<A\$@?W_2P4A>_W!P.2# G,X@59=\\9ZI#SMO&XK7U<6/!=TI:)O%0:=OSW$
PY&]U)'@Y+.'HY#MRWFH2LQ-"+4860 RJJ'C=5'XY*62!SQ\P^NC;O+]DNH7>''6L
P@*OBD?++!X-0@%29F7.OJZ&_)#*G80=8!(5[_L F?AR0K^4^IXELQZ.J@"Q0HM!.
P_[,<"V_^*1>G)[OJU;%*59KF>MUQ]XM*J*YE^ES-A@DB+%K<[;Q#%?=>L(SM6A\#
P?R$61N##"OZCUO1ALT A+QX+R%?EM0NP2E8),L>+;Z_D$J>8HU7V3@\@!<66 "/N
PU+_!,^,)=0,F9)QS>*\4'$38;4QG$!/NT_D/LP(X&2G3$=O&KM.0*T,<D!W5?9II
PQ$:RV#%9FTRFU99ARK;@ O2=6"#'<&>!PYZ>!PC]3%KM,D,IR:(4-HIZK/ 0]Y=\
P85P^42"M#M1,0'^_T9BH,;=F=#O%%-/ K!(WN3'WV1\M+T YJ+/+)'09,TV!S<U 
PZ7R.9%RX=-+-\V0D_!T\4=U$# 6T<)/)YP;X,,G<C)8"/(,#$33P91@V6TY7ACBM
P:>N52%/[XC<7D38#QMYP32-Q,69XC\)_OML%,@ V6)(1:2H;N]L3.<D871%.KO Z
PE W#+AN4!6C:OT%=G[05X@ QJY< [TSY0BV>/'T^\/QO.-4$\]O,66!F*3WL+RQ[
PSVRN/>XU\FF["I\.,MDQ@HIXPN? (ECGO+0C]_PWL.BPOIIMDK&;>J K.(4+^J.1
P6<8_'.MZ,&>OC!,"J!"QZ\Z;$HHM89#NV45LC<2@[F.<.UD@:(F&,/+L09!X+T<<
PQ%V'#GXUDS[OK@B>YL_^#E30Q9G$Z9Y'%[*'0;;GK2-O?U:(6BF3FIJ5:&'\/6)1
P&'I70P34P41(3+,\Y>6HGT"*:Z9DF?[D#VO3>W<NQ]>G%T0['TN2!>[8'0QFW"O\
P&@W1TI(!^RV(E$$>,VY0F-6("NB-^96_]IN%W''0I4L(O_ZDTVG'T&B-0%ZKEY:3
PT'ZB:EL.1CEI^=YE['&8S*SO&#=GV)O\YT-!6;D([]A4<ZR3/UV9 X\T77R)9]V"
P:\9HEO2HUH[QLBB&@G? ZSUJO@ZWKX.:\>F.OH1F(UF:8S=YX9H8Y^@"B43]X98R
P)-SR[;;6\M>6LT, $CYHM#Q0CQ;CG?OE+O%S>DD'8;9X29:H8WD%UN0$DF'-4\8$
P2"LL+YQ3R>%SSO#%A\^;C#Q,2B'[,G_EXOFW(+W1%A3XP_YRLNNGA98^/<DHT1N4
PG!9R[U"C6+LD'] S!587=%#799&G)?"UK!:=("(;)V "[M10>QE957:!;QD-\9K[
P9(0GEB")J(+NDI;B'2<6@W*PG08OO0V0N(V36)*^3NT=9*.&(X!\=(B$0)UST*E*
PD-V9CQ++.Y@J?MT2RC6]XD)T'&>2^_VD71@"7._Z:3\4)%GUNE%GF;&CDE.S&K![
P_14D#ZE(6CID8>3Y69#OE^KG-G8=E*8#Q1/I3A)1L*Y#W%%GC0%MLA2JKX?:0K30
P[%V;LS 5_JL]M-*L"M=0'&&AJ.E_( [3=_(ZR;&@.JPP1V/A5IDL\T8[^^;/0<T9
P(&&W>&#=E+A-'RU,,^Z(.SVF38D/+OO.D=0!--F@0+<":&4MO1/Y_%!<,.8NPY-:
P ?L2*T#U8(.'[5&84(85N(K]>B*:84(-*CIN2\9]>X64EI3_]X24<TLZ<^0+WZ*&
P0F$2>0)R!_S:5AM 55!CYVZ[H.%'65,\2I3)\[NV'R:](@R"_ALOH@^!_&9P)#L%
P!R%,QE:%_ZSZ1R +J;C#%ZLPN-,I2%XK+[I9)U/F(EQ"9U% 8%#JK(=-!MZ$.AF5
P6+4P*?_(53B& 8*+DQ;QJ&FB #ST3QBSMRTMYUQ;$$/L8,64@*;E"Y,',O<+G&]*
PO%'@ZX5;R%FIE:_*WWZ+Z  [,E# /KG42J\3IM81 RG2-'M+6/5T$8E-UZ6X8I<U
PU_W;F1K@<./2\)7N-.7%SL1L0\J'Y\@9CAA^D?F5&XJQ(L :KZY17NS9ZJGW\--\
P\BS[_'B"4+7)D6'CDMKEVJYYLXMS@:!>O.!\56$7!= QL_OB36#\O!'AP$@'^<&*
PBMHE 7$2)B];U3N14'9)E_ 6K1V,M^Q_SGVM$;87#G;!@,XE'U1L85@6/$+0Q\"7
P"(W'D15_,8OQIYQR%K1FD-VKO[>.->MDO?\SCN$KJ)*8H@#:AIAKLFH$Z5,Q XZS
P9/'LJM%:/3H@;?@*U N9H1;//\(59Q\YZU0W\RRKJ$H2=C:6HHI5PD1 ZLDJ(F-)
P+C@Q?A(&9QP!91*+*/GJSE%>7J-/O-+^I<Y<V[!RLIOZ(D%&,BV46%5B'KDP\_EY
P> V5KI:$&(0M(?[Z21H4ZD^TKSC#YG)<EBS)343<1]W#BG-T8I()>FDL5NK.!YK0
P4_@Q!W\''4,@)'%:2.+/:6?.C))%G?&?*OK)O6M-(X!U]0,@/#]62,*1([(G3=)W
P*-U?8MD$Z?$84T2 IV]1<X2I+5P,T]-;4MFDR$JSK: /$(V#$:S[7=[6X?T4>')C
P1&\0(!5X^/F4@P!%EN3VG+FH[,(.:/R6I(-P>MSRR&@'!&"G8WIOTC1 JH [=J,M
P6$]10_L-9?]@P0C0V<NXJ-K7?6$N:A3UBY9*CFU8K 0X8ZJ\W2.K9UC,[8X *O_@
P, 5ZA:-7MWHK=;+W"\U_2P*/4I=[<!O:(^PW]LJ/=YZ$;L!?/9TF08,&4 7L&Q?9
P9K%6,**M#SM'8A5%PT=*$V-P?&#H Y;"$K8H8+0L;A8 [;+%\8YOST;Y4PPPF733
P3C&187I@9C4&TF9YU"9D9URV$RD)6T5O4FC1@!T' 9-V527]8RI7 87+Y0]96B'.
PW9U"5'5^MVB1N.2[O4>N"C,J*)V^29"O\*0\N*(+#$G+W$]/BH]J&$&&:LRDV;XI
P5-S2Y)81]J/5QURJ)+CY2Y56>6LXTJ,Z@"W<2I4V*$9-&'80E1Q*^T;\'S*QF%"\
PU&9=M.GXJ6DIIO+]0$HH6!BSB9>7M2\CLY?QH69 25'R9Y+;@U KAE3=C%I*BG"(
PGD+$\CH$+7=;>#+?3<FM(5,,(TW%[;T+71D)M<*J_.@.>%K.>L9H3#PK1+OQ=?^*
P%'(X1\S,:OIYVL$M<<!+.(515Y7Z]UU[:&A>>X2.5:(P^:!LE)(#T5 &B:%G1<B:
P@)E.!6>G7^J80&U_:39*RG'>N*)H.0+#WB=8C?></8ZU(!C2V:.\1A,?*_4=*<0N
PG*@HVV79#7V:BV]QNK/2,HLBWN@%^FH.]54CK +(.8/^=E>)<@O'J S\0YVY/):F
P5-,)?J:SDC1J?O@RVW:2_GK=)O6__&+@E!.GN-0,U"4CH/?KSP4-X(Y&Y+(U#1]L
P#DW8^5'&LQR[?&CNBN)9Q3]#_?N@H12E/<UN?HQ[<<QVPGE@15GZQG1 K![?.]W;
PL_7I +GDT[!%(WR5UKBIIS>W>W6O<\^/C4[''3G".+; "AK1U$Y@7W'P#X>AU*R 
PKG>"^/GE$:\9[_3WCVQFB\J\U^>$AM,(X"S_R>?P8U"1-9^O\5D; B&A.(>T.(*!
P=A9-UA^PX8K_LMJ^5N>?5V/+BDG6>M4#=@YUBI2ZWH3W9CL1B(AOMX*)!G&"P9;>
P-^>/=D^V8QB3"!3[/%QX=49%VNN\>)H]@!/9$.5Y&SW&1 :JD6'A+-\JUX@Z-)NX
PIZY1*#EP?92KF"8LE6"S.3*=D&=5^-YF[BWT#BPX_FR5W:VB-DF#=YZ,;G2#:ZL&
P7V&4)GAQ5BE##3(;E/ 0&T]B'68VC)$O?9M.0PASBGSP#I8E43A!FD]J)R,,"+6Y
P%J"?QH,O>DHP'_;7JL3"0PB>2RI$1)R^#+33; M4G7(U,T6T])*>?_E2Y5XPY["#
P9 7LY^>YTJ)B X3LV:]79^87[N!H!8"JCH>TG9S"D'EN(M=F\#V^%8MU FB* S5F
PM?:U0)$G#R*_\AAWIYSB)0D >@8J_3"MP:4KZF6KP7BXZB=0+MX,4.022?%Z<Z/6
P=&R$JU40MLI5=WN)>71O:=]&:9J#BX$EKK<6G5P1M8;4PG6T!!(C3F[J$RRR(YD1
P(*1JD.B%7U5%R3NVJUL)QV3X(U4EG1CDF(A<H G\;0^P9@?W5HA"-Z'_EL ]@N@P
PU"7SK@Q=/UG,QS[JA\^V)92B(Q?H?H9C#_K@6 B_'7Z=H]0K35+ZMXDUS?+T=9E,
P>@_+_PA##J4H*?,P]'GK%A(OO]G<$0,VCN"2)Q$QZHD6R7495#Q[R&-,<^H[4,$R
PN!/FL8S8T^MG<X+K^MDCXPU,AT:JP$3%C,%:2^D/%90B@X+7A(DQ^= $8P3ND@CT
PMV&CJ VT^!I)VSMDEWWC <EKTYO\AYU^"_R7QD:JHU>?H5,7B!%>.Y?NE6?]WG$,
PQI 3+DX<[33:J*6M=[ZYQ?7PNL"@63(^+=>2#(RE\OY(0-119)<)!A)UA2<[/PM)
P.\SAY"<\G9JU_.OYMY9XI.&$0EFH/RT(1WH8VGH@H<^KFNARGOVCJ+YXK:)?"^#5
PQYH'NMZ+/GQYKT+*I75'EYH^RXW+3L66*)94^"9H_2N8J"%QU+G)4_8P'X_XDWA#
PNWKD^+CPFK#Y?Z0 4D%H91W)^.&JNNGHWX*9#Q30U!B@E:I&'J>*J;&+331B5 FI
P*BMBG;ZC_9[!LZ02'+\$R<Y>5OVZ:R3]%1G9L<,[V!&"^CMO^=0;H">.#3XG/VG5
PG+3(@XNSL,Z4A;C,1SR77$!7Y6]# 8YHHJ1?Q@4;%,I42.I>:KM,4P!4G*P"_& I
PLDI>RA7N'^TM^I*!PQCRH)EHPQ'2+S3,)^GUP=HI\R _F]5_ @*.<5<7MTSHHY)N
PI2#, A?@>^(Y0GOA7<^^99 #0$NV<U#R:A-H2GTF(>*AUO1 RH@@N)#0*!\XK-^!
PX=8H]"J0T&\>>JS7>^DR"=S2QS'1Y:XRN7TO9&!)U>"M"C>#R:32S+4>'Q)5ER-Y
P'K-B-O);S9+MU"]#.4_LKOB/[P3<VQAZ*NVQ)V^;(=/^3MR/?=I S="V3F'B1.C<
P$?Y(0L=K,AOQK.&P<QR <S1KCC+I4;I'%3747#$H+R2\(;V2)9;=4$=-:3TIKPD"
P"= B,0J4M?J[^@82VJ&F^1?4\VS--!V)TD+&+"IZ<@H]//T;$&-A.VH"KR=M%F4?
P(XYLWE0ZXN^H%N\=N[X[TZ#U812"X?8H9$<;;]CM2+)R46?C(=2E/ACVC(*3_,JB
P"^QM)8TD='F<5+=,)QY.\>002FYUR#,C:OMV)J@;M\&(0)VI%THO0;.VK=)UF'/R
P\ST9C@J"01J"]W>&D,O=Y-T4;ZJ4/((CF!86RSF*!*EDS=FY'R='2/(0].O5SKE2
P3DG?79+SH$1RC,EI>0?(X;.NWZK?+ _HW,W61&50G,Q%(*-ZES"VI8#+Y/SWR"E3
P9HAQ740:=0?"K]B#(CN*Y1<$_3LA0+@LV$[R GMQW+PM86.M@OCAKA5-\X->2CTY
PZ!<1;U"4<0A+[G!'<Z0W,EPN/MO82ZH4B@]@M-^AS)@2KD:(@_#3;+.&HC(37D4/
P2\^B7)(@"3_2#]=@T30S;"P^_$88KP,/!OK\N/C-2!%V&'-!OB]VX4,?K VYY*,E
P;93+T2W)I#1PWL2\YCTD!2/&)Y"C*91U;J>%"A5(;(]K#0S>%ZU:<ZP:=NFV&,L8
P,2:7U ZX0+&(ZQK%:$KGZZ):]$NQ#)$7 ;^5ZD<7?B+"4)9Y4=UO%6^+XK_Q$5F]
P,NO$R0?\C$G PF?@26A91:M^-2 BB]X\K3HE>H: ;86BQW*F7NWY^D=K5';\IK&3
PY+\[=*.?'R35';Q4!Y\#=E/GBT@Q@.WRCV#+!@ 9XQ%8M=I7J*5QKK!+. ;/(FI+
PH7SNYMHK#PB4&5N?>5'ZC^8PI;-3;WS'RE5SKV#DC\.P2E#^_DZ6]'89?J(7T4PX
P3A0VEL)!8(WY"/(69ND+C*5?>-@4"J5XSF;16'N^8L[+EDX<B#_V_!,<-CW4MDF]
P2EU1O0? 522"TR?QV8]J9RKQI4TF-Y;#U6W@*CC-<V\A-5,UC-$A)U_YE+5YG5T!
PZOJ941@ET@5E7G )HT$0I,+65^32X3FGZ+ &4CP<_NQ>:M:945PXON\A@A8%U?R\
P*78W%G2=#9E+MB#%!0N2";B#J>;]4&IY#(V+'[[)5ZFO2P5="AB2CU(Y P- >U6]
PZ+L\XDS'GK6.6 G:6,%H"XLFZMZ>]-8SO!)38H7>//$IOMI?V"&RQV97B?:@+KSH
P,7_/"*$L6]!VL=AQ%A;6I#CNB&AGZXQX;RU ..5IEADW;Z7X+8[I2_(.9F5X_MOJ
P[A7@[2)8O6_H)7H2_:<*9J/--L_!LM]3L$;M8% [ #P@YN8AY+,Z-)$Q-&H+^P4%
P4L\FJ\O*O*W OK=*C4JZ2O:N2SLWN%2,;N5.X"'.8W93V\!E2FI+:9W6/2_Q0J@C
PP,RFI:3%Q7[W-3)\\NOOW8:(44?3B&2G1>T]]!F-IK%8_: PCO"K1<&KZA^:BFD]
P'+N.M7@G/0)5<.CG?Y%-RZ795*?P:$$Q<47$BQG^63&[<YX 5&K-/[B"&2UQ;:5K
P2JJLD$\^Z5(UF_\OA&[+U*HU3@Y$%DFN;_<X5][ W"X%,A(S-):.Z*4%4'I><_@4
PZ$.0%)2^2U<>R.DWTD9R-57W NTP/1,1[.KGD7 '4HH+G_4L6/Q78(=1FDX=K5E:
P)0)>?^EY1R^$_&J+%.JTT7IQPH1L489]F';]0OO6ZKFQ^.$MLW+F8=J5!YT\5>\"
P1S?'1?3Z*>]O(#;SGM_/:&"+85:%D$OU\S%6$&(P$U PY@?77%X19,D5$1;BO<\.
P&LF(L/#X^;^*O,32--G(P^RF#,_@\N^[N0:Y@4[,6XS^/<-=^9'/P&LR9_C$HE.0
PV3,8WJ-(<%!ON/UG(P3#T)PQY';HU-^76>M_(UR1W?'B;8V41X-3[--NVN44;CTC
PAHY_=IA9]>R%ZGA19OLH3%BDF]X%GL7T&PHG+1$RG:^@\1%_8?N-L0KHZ&_-S1Y 
PHK).IW-*B5/BO#[DHP9F5PC;+]DYYPLD?!%M(;%$&\CY;K9E1S-B#,:*ORFD-B2?
P--OT!^[V[>QKPUU)'O<?3*YO=@RK!WJ&$4)C=OG-YS9]9A;$@4?NN@*)-Y<+!\%(
P8G#"*37\+^J<L\[<<& */ZV*]J9UD.K/,+?Y]3-H?GFDTQ/W]3L512#KJI (H\Y+
PVOL=0.SU2=5  A0%_CPN&AGR</5]<,]1]U$T@+U=49H[N,V7\W=-WD7A$@,R%WW@
P2MWEP%^1)\5&*9VO!:D  R/G@?LB#H-0GURB^856:&@.6[8W+VNP>C&#$OVOB 2"
P< ?5(;KX1\Z .89YV95@C9_%+6,L&0YG1NH19[;?KG1)=J[>@' RI+,XV;6KF C8
P#3C#IDM*2C-4>4980XJ6,>J:F)W2E,EMU7)S) P\QC[M)D\G]\,<1I/Y^UKN][]?
PG.T6.+NT\Y78@":LS0G+,/X4!I\TEV!&# <61RA@$3NI*2RER-05@J1VA<H!\>Q>
PT!F#R?:$9QZ>T;YY](*PLI)!>E6A']VI.!L$ ;_/OR,[&(:-V6"8+KR_ X7=.1?-
P^,\;VL2[?'7HR:#C[V62E,Y/&/.!<VBH;$]=4;XXPLC!_T#P/+ J.J;T[:F, ^D,
P+0WQ=X554WOR8XS.U(A\\+/')!9G=O-F \%F=LCM$V<,.P5%H0TV^-!M6;>T"1+K
P^L-+B'G9^@A/*(M_]0(-7#H!_V/TS?L',X;!3*[*6._0\C>"\DF=>T.K&QYHH-$[
P!WQ-&>-O^!"7 +)L83D/-O/D&,Q-U".Y-']WOG<B.I^D4";B#KR&!P$:E[[OZ 3M
P4RDI7%;QS8TB3G3%,8*AR$@:EKQP#(V.C?AX0RV@=O\A 63 T+,C=@AQT*. 0IS]
P'?@\+O(9<Q]9I*BC K/- " 1)]@J\D;THR/?LL=4_R (!Y2EX9SOSG757VQ&9\2*
P=AS8IWFB_\)!)#6\"]?U;=U#R6ZX]=[ZJZDL5.N/]?FD%QJ/3EOX#(B>H_L-5Z>*
P%+#_:BYQG7F3<I=Y%$,#A8ST!Z?UYP).N;_ ?U\T0+';875PB9/(B<3O0+S+#C.4
P%DSS;QGT/:,O3 J$&(D>KG$E@VMM\Q00B1VPIWA'/U(ZBL3:$FP;:0LC\7/@=SZE
PZB4"C'&1@2]::,$@ZH_6YA\QIO@'@2V B>G)H%*#\7:[Z'.XX99=YXY_FNE<E9G$
PK3J+<C$"<1F(/#R<\T^ +K!TY=Q+;R*)E?@FN#PI<I0/HQ"[6FF"YE7M]>2#+A'_
PGA^)P_GNX:JAQ5;OV\%WUZ08TM)8O.T(41SA(IB!))&6&%WOID.[C5$:(&XA1>C$
P1F2$NECARQ^S#B@1CT]$X;4<;5EM,?:D]V"61=*JP6E%O1AXA^SU8B5D0,WZYL&U
P* UHD=V]N*(CG>C_?[(SVV20'[U)@EG*=0@YT'3K"P2"S^=&^2-&;INKGRPVH"*Z
P3H.[6Z8"]CPLA];&!G,YM^XTW8Z!JV;_*?%OY\YR%\VO1I<8>>(!Z='/;&8;C6EF
P$/H#*UWNJ_'ZN@+^$-*H%"T5-E/??5N;4IYW"X#?#(LA"8A#PD+CDM>ISTK?X7#-
PD%$+B'XA[:6'=&GW.[W599J]$78^7G[F114><^Z^3!YF(BUN[4DY^2K("\TI:^O[
PXGX Q1-5-#JVZQW=9\]F3V891_*+"X#FJ:-G()PT/UVHQ%=(]_HWW+"FA$%=1Y17
P5?_^:R7+&VMRKM8%&8EDB?"W7%CS^H)I$KF_)*4N(!Y&>RT<ZC>Q>KTBBZ[F.$)K
PRF=W/%J'0:4.'Y0,KD. 62P'TT<!G(B&6.#3SP'WY]>/11[5/$MF;@'#1TV[X&;_
P^EG<HF\\GPU\79N9=V9FL''C>[J+ @AQV\8K]MJ%R6"SRQ_6_4NJMM$;:Y=4$(TJ
P^Q#'&4:",XN^2LB*N!M!4$K;%1D.V&) W/OJNSE<+_0&O^1.T-5&6;5%QNL!"P1X
P8S^/(L?D%XMNA;$<L@D*':*RVRQ32H<S4.9+#CX'\NO+%%9=NJT&5*QT'D!O[QP7
PR4IQB];S.=&N:,$>=>W'M:VF^-J[Z3KJA=.H^>--1B9_Y4&07:"MJ6Y%KYGLE_'X
PN?6Y+%/2. <#2:>"UT3"?WW?D7J*/WH5; '>0; @*7#V]Y;JO<G9\5>'T\9WF6Z2
P%%^CG-T\>;A61+4@L@Z[4B!IGM]I0_\CS(OJV732G)#K*![+@KMUU',<>#PF+#-"
P#AG*:YLR9(M^?(_RJ.J NK7 R<.R&D]FFO6KXF/MTB7ZAGI[.LH^#$45T7K]F\!N
P=L.2)_#@,\U=\6- A'?$K5OH9)]W#2S@5BA3O J/1K^?>GQ0@6USH59I',Z39ZA=
P_P#1)6NL$,73O$=6HO-0&C(RK%H:TQ]/K8K&6TT,1CUYC-!YS$755SL9B9X>8;M:
PI?_Y"M+93H8]@@J4D7?8;]!R';G^AV;+ BYNB%@5D?A638'\FJ]!]I%VE-[W1GW5
P+1+7(*_!;JST[7!V=A75 9WV,TZ4#&[R3ZYVS \N!O*$$;+"-OX &4?L)<;J><4R
P>70_M[X7";=DVD%(X^;K2N.@O<#VBBN3RZCDGG==#$%_GA[U.W:F2G;;\*T 222+
PRKI4 KDW,"="!FD)BH:Z* (=LZWAMVY9C:B+*KH_I7%V L"3P7X*T+_NK$PSO['*
PE6/#%YE.A2Z&"R-%L0<\2" %;!=]5+@F,$*X=_MNZ[O1@=^WP8#DV1"81A_;;NS]
P2,EA,39]3'<'B/<'S4<X$UB,Q;B+ ,P\B<@T"Q%KI*?V*UT\N= SJOE"\*04+.FY
P'VM?E_*LJVP/\.O3_C<>1BPT$5P9JGSR4\YDR[THW2./-E>Y$OWJ5/BO<N87VH*,
PJ\T=6I,.\NK-@+B!HL9RB+02D:WSU=):HJ?8:EVI5.0QA$ _NR$D3^EC_SE^E8JG
P]JF%7M3*@"DE,:?BVRY=J;=:A*=&Y'2]%G;=D49@Y[70G"^M;$<+U2WV]"W0IM4)
P*-_E5"/H\Q6)V^<-"%4.H+^)O*-Y'$]E$;+_YG5*C#60]B.5QN?KB('(]+PE2(Y7
PWOGC16A\9DEW(-,D,Z7TUE1NQ6I^8PO]-UM.JM#\2$CS2]=2(@EL0E+Z0D/0 DSS
PY?V3$HZL ZBZ"(*S:XZ/NL0LT++VI59W)]K@H6:.14LZ KUSQI"U,+LD_'H9C[0'
P=P#]WI;R)FD)H&_.S3 F-L?YHXH5ZM,M9>RBL#WOG,\QVYKUFUJ7/_(V]1-%FSS*
PD+]M,0)&G*N3<GY^3M[\!2G]2>(F%2-6TN1+FQ>3J?56-1U1O03+*LUZ,U[?KN"$
P3= H*="$2\L&!OMBFR^O GW:QI'*F!^5)-J>^B5C$%Z! A*D>;S%=&M5]W"8$-:7
P31K*,".B/(5W)GX=C<Z"@],OLC7E02\85IY[>FMP]%P'M3]G?T5P0@=5W.#R^?<?
P+WXP,ID\[+%'G@OP08*+/MZYO'DX9H''.$\A Z[44R/8T9=I^#KM#P!D&P]C/DM)
PPJ),[_1"2&@VRJ4SV#[@+4=+1?AB0P6*%=8'6',G_/*"H) G?I@VTE62/U=Q"/RI
P.T[>[>%;LQ<C6[4[H0A8JMZ*<:GKB548?#,OF+PJY#(E<PC;@7/K4C^1LJP]S('-
PW&58:EOK%[JQ;D85,](V6<F4#L<=O"X4H#NK?2,!!7(2ETR(%2!=M+CV4 IQ_#(V
P(T([@!F8(%R#WZV#$+R0PY2K(?DO-K!&&..DI/LL)9^-LSYZ 45$F,0CIBLGRJ2N
P5'N:/F;3(24+0*_&J"YNSLQH>]$&3Y=?M(F8:.'C/1D1NG74VFW[#;W_=TPG2;$B
PSH=4\]]52N'.7A A'YRT=1X;13[*[:1-+[PW0GI_%!,4HUWJ\N6SF-,,R9,,=I"#
P^'6^C%(O8Z2&F:MU!31(I2$>N)U:+$)U4E737Z.*]A49@.>D>*GOIW>M'R]4AS%*
P/ENK9-%]>%0,$8, >P,ER$1'-]5%=O$"IRO\Q_OS&'$&9:;*QAJN=+;,V2B-;*R@
PIKVI??4R#$P$=?JBU_HTHL\LR%HT7S =&?2QBQ"C1O-#J"0%JV56).8Z_ 9'DYC0
PC!TP16RGA?SZ7Q?Z,$8P:KPZ)CWHF&[^H?\B!/#0R#GB:C,F[:CH@Z)K+(#D:$3U
P5]=VVM9H$F7$8L\6]<J8K*(Q.^;F1;FX"B"[:&/^G;^W^38#B)A,(%MH3:LL#(BH
PE\0Y6@ZFZ3.<^V$,7#-21YQ$_!S8B+]&7-3-@YX%.&, 5[VS/[W.5XG?#GS<0A,#
PF3'H'LHUT#R9UAZS8Z1="L;V=Q!.39+ J:4.,4PE#!CF*7USP(\ON7*L,E1Q\BAC
PDA99DBIA"\Y9HKZ;]YJW:CSD#WLNV3SC=XPF*/?)PF5JJ_GEE?JF5T99@)'!Z=3G
PC3-+*35BE<S?7-TJ2$!38$^1G\+YUV*%\X.V',VJU1S8&)^,6L#L]8.)[+2CN474
P:6:]=MD=6@8!UU0V0#2Z5#A6-C*@\_D_ ;3M'3=_]>U]?^1Y6U]=:)?=&@PY+>I1
P2)S$9WOP5JU@52S.^XR'C757%0W)R[<6H  Z)Z"YYHAU5PGHP"U5+;VEQ"M8)3&!
PL]GLXIU]4JFQWS"\9N8T=%F S'S[7&;D<N^WI$=HJJ*>DJ9D(>PW"!V1B0-7GZW<
P_]G;>'MNO-8IH4+?IA:<TLH[\ F]9Y^LL!C(-VVMC):7.=@51#N<!*A(OYQR24]"
PVT0"(ED8%E1:"X8R5XKUF!U^N3^=AE+V91]QMXWRQIU>P\1G/VR^],=.?'EK=N#3
PTJ.\DL37S333T93.>S?'-*/UME[*G,M591<K@1EMX*O3_+HR5*+V' RO(H:&VAT^
P/?BE(569L'^3A"7O0Z[A(1M[!9EEV)6?8''458]3J[SC"[71@S 31_-E$U@PX+)N
PP)K<0C[$OWP5V16R"]68V'L0[2.!S'!1189MM@EAR.4-^T$"L'_)@)^UPLKD]\[>
PW.L6%U?R""%$&MKX:LDPA+4N.PW+%8S^9;VD!(,N<:2UT.L7Q=)VX[@K"&68=B]Y
P89S$?[2[Q,W-MMI7U19RV;G&GFJ,?M_8UL_K"Z1&^@JE")2V-;F;OV+'<F8>R$%D
PD4)*:I3">WOM<>(?6P_BUP]5 *%:ON'=L?J,6,"I"*)*/\?" []#-BXR-P8#\?[ 
PI74RP CW->5Q8__7- /S]P !\J"RY62#YODX%1C+9@8[X"B'L4X?&,S:6N=6%-XV
PEU.JB%ZAM2LO\#R].\79>8<J@M'FQ$JE+JQK,<R^J2>1AQ1.&@SD![7@JKWR-O6/
P5S.)]D8^F DA6=!D=Y1ZM2X'*VT#%.OB/_.'8\), N]V#DX5!!A;H1[%\C]Z]6GW
PV\K_V]T/WT:!]NCK^6:>QW2VY%/Y\^',2)S07+D;^&S,/ CGID\[V$7O;F'&<\K4
PS0I)0B-QZ\;=31]*E8S!,MRC$:F6%FOG17A'H0FG<:1O3F](,E[IRF$TT[LKG)\I
PCA%BFZO/^U-@6I:.()J +<TPVI/SN7(I5.%'=. ^](D.OH#>697!.927IBSM'07G
P#OMX1P-:+W -=DZKU0L$:\4IP47?^+%&UTUG*H=GOHI;HV&<)IBB^\ODPMFZB_F;
P#S'5(9F20XNX28\*"S&=*Q\=?DS8=0N.1VD%.I:U^6)._!X=X<^)YL5]YXA/[6/P
P%2\ A+K\RF<+]JVN71RMNL42C<"F:*2NNK5$Z?TB#WE@"'D2'2U^GMT*WUCL-'(U
PZO-\)5W'R=BH8IOE'M&E%_T!P+_QTWJY*?Z+C<]S;!!OIU'YSQX*G<$&9NIJ$E_2
P+.CZQ^I\",9^VP2&^1GR4+ >403(5\\I'_HI;BK)Q]LQ*0"6EEB27\$>MU[)9H[)
P(1&RSBH&%5Q;Q;N-RV_'02Q!3J=DB':F\=983.7\]IZS>#IK(ESSO3O+0KYT]>53
P*UIWVT@/NL>'-(H=4I_\*O(HS%VXZ3*;:).K6YE/[,@-22/%@QQG-]U?3Z5R%.Z>
P9ID1WF?;%3(1)ESL((F$X-R+ZL-7%N4ZXH4<QV%EA3L!:CN)KV]5IY3;E*.X:$UU
P1Q+IH\)U:RU28)59A9MXX3.OU43P(\11"!6SLT/@S3XP3A\/.(&-WWZ&M@L"9T\]
P8WXK%OUN#CY+H/Y_,,^=^7T(B] !'B%QE]LY=]W1GJD7T75V/\:0>#('K]/'68\I
PG\%'TLQ&SX3X\"8]S&"-^)O:3."Y(+W8;7Q<9MFZPZ) RB?%_L?/AB,(D*SS'2O0
PM&?.%#R<LN4)9;9Q3H +;_ZH(T3\HCT;WTLR$2OM-_JD GT)K,)UX4A4\15[N./5
P9B@?5\U@V:I-B:L(DB$;ND;0^B.(=S(Z$\([YNA-A_>%?"^$2:;O;LL3B@I1L6B 
PUZ--U>CU] A $ 0W.,8GTXFYPPV8(%I)S_^H><MQ+7VRET7=O"3C+17V%S$AO<Z#
P^!"L G1)6Y]M^;FBPDA:5CK.5GFAQ1PHJ[::[60$OV1MN;2@=S&9J/NC-"-I_ Z!
PV?U%;[QW?TMIQ;_JTLQJ =-/$(E?]5 GY>D>I23-[N.E.81COM?>T(U^/Z"FH V&
P0?&]D$)ETO&)AS)B\SJ2#[?"W9CG;*E"=KW)^_[]#P)V@<>=WOXO+EU0;^KC#LOK
PM60J2C%PL"4E9Q\2.Y<[D]+_B!-%!)U3'7JB%HCR_TF4\&5)N:KN?,E<"VM_:KY$
PK57+.'^L)19?)G$$U2G[!.Q]M9,_T=VWYID3I.TM(L>1D#^DX::K*M1QN?OQS"%[
P83#A!1/F)>L(!74=_7Y]2#DQMD)R35(0LV+9!+SUY GOO H:S0):"]I#0_BS*6:H
PXVG,+PX?H)"[W6%6.%6Z>T0)32]V?*.P<'$\=S(BP,-SM_YM]D6.:RO$1RM:Z+P>
P"EWQ9R%M;Y3_&N9+C'LFV0DPU@.K7VO#1 PYI$Y&%-"X;_Z4IG=4J,&OK!&;=6@N
P[CE@O<]'.8W<K264X+&1#N=#;0O.0RU+R;?X"797CR^;IA+-_^*DB^ITA*.^V/[%
P/@9EN77R!Z0G()8(E4M, 'MCB;*A9=!?G1$O,W00%T-N-X^$N1IR/S:IY^S5L+HG
P:/K8\7$V-K2I#4I7EN?UPY<%SK0+ ZQ?\!>'?K'O;11-A/#5WR'*<:@# &OKRB?;
P:$/M517 X80*IV'*5@^XNP2,)6HR&9M;+7GK1X>FT"V?7 ?LT(5K8A\*)[4< 8E6
PJQ+QJ&3$/]PEAS$C<,RK&G*1R_;Z1V:A7"(HU2FEYQTW3"2=<\ ^_\DU<1VK=];N
P\6=BR@E4=1_]]=UJ-P1/'.U:TZ\<-("YO=@6@'&O#%L^%>/>IP%LF><V97P?]5$M
P,8^L9\ L8RXW2"KK(; XW&K[4^.;%F@"WMX-\XNKD7"$_G 57M [7K5UZVG2 3IB
PK0G$A(COC[U<^Y XMMJ@:-/$)0"$G=I-KGD^SBP-%VQ_^!F1Y!YHIBO5U/U\,#^X
PWP\1=_KG4A =U^"%'-LHO?7^*%8@.JI:IC"Q]KR)C%YE%I1&\5P/Z#Q=45@MF$Q$
P>!EE_OLMZ<^)CVY)91V5JPM!I:L(Y.%?64 KLUUHY$0:W_BMG&_J^0]$C_2/ &77
P/>' +M9P@M<[@CXV"WB5>0PX+:_-0=18K<X\IXMDH>.4$I9A,  A=@&LY-YE$N1+
PS$Q@E&GZ 6U0"U4?\PP :P.EF>7 F\L(1R/I-3=+_=E?T&[=B7X$7NP10;*4#Q3 
PG)C@L-T<A6U5<55S4$]2%^GSET'!1?Q:$;2AQ/_4[?6DA.I+C@1=8S<Y9SNT0R!>
PJU\))1$30"#;,I2:EI+QB*=I9;^F-[#+-P_^P]I3'E]SB0"X\>=AKYGB\P'-:D60
P36)>$");XY@:6K _0MO OG?-J%VO04:?O@DG; CUA)SNO,HK"#674\HD[$<4V*8J
P?BB%.H&P;9&0>!P:GZNN)BNP64SFX/F"&FJ\O$P*QHOU>6X(!6Y"G. (CA?%#]0<
PXJ?&_%$CZHZ-$"# 6U7TIRO(**=,1)U;;@7WH'-**%]N)7L_#)=<<3*,F8Q,;V\/
P48RJ^$QQP=IZWT?89G5D,[-?-PP,@@Y>V%&O1B>.[4>G5IL;BDM,I';:'CTH%M]\
P%3XQ+T$W0%]2C)<&T9R)^!24BRKIIM4X_$8CRHL#?C(J9*K(0GV?MK#2MYD7 @LP
PP!2/@\A^P7 HA'+I+HY[PH^%R>AGN3DPC]>Y-,=#;G2;P1[])%S41&M\>)XT&F*D
PH.MD%%$+3'.GGCL:/#AR011SGT,FY63.MU. *1'./C4F.RP&X<UG3)@D=8"1G\UF
P#8ZC!.?%,6.G\IMI,>U':W]M2&"?3=H/4_\4T7/5YWSU;V%;38SYE#F-7(C%SP[H
PJR/PFS+(^45U&Y9KMS%1#^&X:,*O(!V0,@LW&Z#?T@S\O9(;V.<>#JTAY(UI[9GT
PGQE!$?S/M4M:J(UNW/<4L" 8/M"W3< W47S,&D^Z3 ;I.Z#LLJ?J@-I0['LCZ#UR
PRR(QFM2J3]]5R*YA/W9^2KR FTISI0\WOU2--WP WI32(A/KRBP6-'Z]0U)\[SJ9
PGB7*3U:48E*4I>29MK'W#K52.L>/!U"&[*Z#C =PJ:,=KD)_N)G&47ALP>VM05JC
PJ\64XM8V)<1\O'RQ76;$)1,\?(V5/#.@8=WT$X(6V$UYN(#2U"-ZM*Q5IG IPKOZ
PL*>&, U<F&_ AP;*Q\GG1&@_52/@#> G,0-/6'2Z.P\55+&A1S2#43?G?!=3J&92
PL:N@VC2Y*:(JD[ICYQCMJ49@^)7+B[YHS+D$"(\O.##@V:$<F'0R"4=P:K]&8@WA
PP@IV6=&6416$KBE0\9HLSY\P?Z^<U''MV4X?;^&$GE(")_,H%++-)QT*"!)MJ1JE
P1M^_-\O+9=1*?ZXWJ89F.E)Y3T^)0^NU_\M-[7PZAC3VW+G?NZ50;RVYS.O7*V3"
PE]%Y"7#X'V?Q!H\P>YHM^GM:AX[-3$><HMV_:.6D-J>C043[^-ZHBX?)#39J*!@$
PB(LPPHD %K':9A0F?R]4:,UXGL\YT' /F'F.@BI;,ZO&I+2Z9:>XJ"^)Y'D?!28&
P%%!$9H]60^&EJD<;PO75J]NC'C?-U&@LDFGIV;6R9$B$18'D;J&NPT 2B?HTTF5&
PH+"ERC"]96_ W+4M06Y7+R3R,7JPV9UE9![@>\O*83K,[%R_FU9EV]:^U+H[@%G(
PW0&KGGG8FOQJ0DM\9/E@&&P R5YQPY=E ++V9\T-TSO.\QA@SN5^[W=1]&0:1;X8
P5Z$D1;(HR5&LN? ^?@WX/S"BNIIP,WUI1M,F UUKL-N2R/U7S_F<%\517ZUY2%D-
P;XACJ>LXXI")Z#]'RU<=9W#10$>#R. 7)6Y1>TAH12S/V3:7,22<[MD ;R<G9RA<
PCR"0MUVW7_LV.]!-."F?U<:Z06EOR"657IWU/57**Z@NT2TYPL_#([5@/;7:!Q4$
P.E:DN>N(C\7-NX 1^@,20LXU'F!"XC\ IMP.:GAL):(Q<$X)CF:GF].%@9[ +'1=
PY^,V4U=7W2?L[1H_Z/*TYBD$?1K2*OV1N QO/M,N]%DO>3]@XG_^FS>F2[4EJ$\/
PRYI49%JJ\A1RG8$%SU8;T">+)8>)3;9P/#20ZQ OM<.HUL5>O:QK>$[J#:^C1R]M
P/NK4K+JY**4EJLH6[> >)5M;C"4IW:AN!S.]6#H+J-01EPP!& F8W(#%0Y352D>Y
P*!#:;=90=90MI;8NA=]O@4ZWEOS6UQ03',&+1NU)(-9,QJ7<;@,4)\L74V%#D4CS
PZ_M-7B^.> 8?G0_]8USJ4KA:TS+DZM-S"7D-/B,9]X+IKG$H0TL,5MFI9 \-L-0D
P2440&0_1HE-<8/ER L>ZT&F11QI1]*5_ 8?,UM/4Y_GLD)"Y@LO4;_*641H_E4M(
PGVS.]3 6^JVF_929_#+R01LG0L7#!R)A3=X^$P@R27/38P#8X[/+$EYQ&-F44F]/
P;R(YCLM2\7<KABL5?*&/S@%^>P.I6\O_&CAG]MK7#,Q@>S=V8%!?%D?XBX^C"<UE
P0TE[;#"./XEJ=3'4Y G4:(K:N0*-.DUVKZ13G&A.Q(-JSKK7"__?F7D8A>DEF:3V
PO%@[5GXXTE^+[QYE"76H;;.\I/4][U_:T$8KRQT50'1!_-:;JCEXTO(*A (K1Q1[
P&=Y)1I'QP3LNB"M/V>?$>;-"&F4V8H,>G[*Y@UP4J=NV9B@^PQ8T&SK$?[[12CL2
POAQH,@Q2,3C</4=HXN-OLE,1_>]5OEHF3!&'>X5RDD+%QZ%*8SG?J)X 8)W=9^NV
P<GU8FW=YW\F?; 9&CHLG*T4O$H7!T;H^#/H?YR$4#M'B\5S*3!EZ:+ /YF#JUH 0
PS\K!;"/"8EIVHJ96"[?(4SHK/)\]<7!*\YY=<<H6%<!$_X?X%Q^UC&,V /<NSKXA
P_O<+I,EE0X;(>&!\?3;(BO%@63L<]):T*+.?SV$5E(P^$=G*ZTRX8'=7#,**9#ME
PQ:."1>2)_Q:KKAT1K@\YWAD-7&=K81C^]E9OOVD;Q41!Z3]O_DWNOQ+M5"&1(R'%
P]@W^8 H9+2EK^>#R14R7D"CSO,@GX9TOS(U70<&,0?5:$22A4J,S&FS85PWQ<=)\
P;$3 M)M+.[\T#0H>X43/G-#M/<@_?Q=2_$,S;(?=OM_&F?'P"U2*,;QX/0?KFGCY
P-&YZ+FYK<RM?A$ K$LL[77I?%>,Q>TP'B;:Y^=$E'[Y4T6\P$/$VK<NP\W\M<^W6
P*NCT_:?7X*=XT/?A=:_VU'%A*Y*XW70<HUY,"02]*,$P4GU@MJABC01&LH<!FF^.
PWG'.-Z3(T@$WK;"A7\&\R'#6:H]>TCCV 9%D\C'G;NYERK/D;# U;RG#Y\#=Q'A]
PP]Z.M_Y_:N._X$9L0(7,Q</4W2YFL.\C__AEA@O^6TO62?;CRERS,M9/5O4L0L08
PQ/5JJM'T-"OTSS?/74ZWDI*090'QL;UB" X"&S'H1$GZFM=&.U0:OU\B.ZV=9Q.B
POQTYH@J#;$ZOY'1^"[G-)<]@3WF4FFN30YAG,%>NU3PYE4:#;O!\DH/BBX(D#HQ5
P.C"(WIF*U$.9*LJ2X(8307+^CH%O:!(U3%7526Z<>0KV51177A8F+BPK@'"/6D?<
PH-3NPWV0WZGLOBJ;9MHYM?V\\2]#W%P^'!'!O!8FB'*\JV.:@;3SZB-VX!<T)G&+
P7/=IQ^@TMEA./-^)YB'GG5G]OS55 [3 E0!^9COBWQ/4QI'P\ZA+VL"[^Y<]_TJP
P#W.XSC6->)6/U"\5;EF'>7;+;F\U"A9[_X";G!KZX?JU^>5B% 6?0O:G#&KY@P1R
PAV?',3 C#U5KIW-@>_:E71L545OKC%BNWYWF[F17-)B[+7XX59* %1NW7(S7:E8B
PB;AXD[S(.9Y=\2Z*LMBU_[.R[HT>9]A)@0=5%/\X<JPY5QNO)8?\Z]BVJP^N_% ?
PW4;*6.?_XP&9FRJ\O547C%/"S2N3I_>A55P#\3AGE!NE;.^&C)S!?L-/J4&,@Q]"
P',D3^.3)1Q;&>F*6H3'V^[-/(EX<1'1O2COWSGYD= JV995<Q\V006@;C6-5_JF*
PG;? %R?V$@P*&B'T]_*I_$6R5AORW=F$S[C5.@ .JT6_$U_Y(#*-K=>8O-Q1JIL[
PR80HE"T%:'Y1OY_.P+Y 5/W[(F/,[DU5T;)<Z"ZY&/_B@P]&..7%_O= J9J?#T$T
P-<3%#^ ]ZCZ5BW1N776/+MGWI^N9];!:S6V"-$:O-41'MB\*)FW=S+H0<\F_CS6:
P\\I7:^4N/- X"QX[$+V7<<9][?_M"U2V+1Z9L;$+/KD5-">S"UO!YS,Y!W79N<D6
P]$Z?W:=<&(Z^M_+$V" N2*Q*R8+Y#' H]S'V5UW;4'C5_G55<4'?SN6U^PSX_ ]6
P4\GEM-H4L!1/K9T/P$03\/V]*+'U5D(:+8!\]BO:%(]>J= :$K#3-T5)2 S$[W/T
P,LN>,1@OFBG=?6<-H0\LB-V56>-!_A/M:ABCA>NX1-J919QUW&*4NF\V'V3U#3(/
P@ !RC,D/?L*6/0:.=97$TRT-)/,O]C!P\,!J\"_U%K3R;G$"TL<O0M.O=L4+N!TN
P@&Y8=5/0SU*NBZCPS@^[ A"X5$P4^=];BE]X+IZ&R@T1]U^NH*1BP6^ZMWGD6J]#
P ,F8T2* MU 90:(EN%C9WL?LZ&0QQM!J>?,6.5RM(6;Y4I!4@,6/[+Z+<#NF/Q]/
P C ^?-M*U$EV8F_TLZQX"RT$5Q _,MRP +CWJC#U&'72?*"M#E>'TVUJ'1H>U$PG
P<'W?3/X,F6;%%L;H<FM*=E/'+S)  S!_J,DDX+<N(CDL RS00_4.@Z?>&7(YO\_@
PY*?6N%TT\\+<HI]6I62R6R92O$J5[9@$F&:/%QX^V-##<O,+LBTH:7Z<=@!'3)L.
P_C.SM,=,&6_52=H73GR[=,V2@#&P-_VL8+;F?@7RPVZ!6D@2V.V;2\LPVJ^V7$"T
P8:"D*>'4CD5,J?']M^4C%DB:L!H&) X)V3IS014-\U%USE.F7LW(FBB/&#^L0*(7
P-3#]"M\W^-]YA_)0'\!W\]Q3-9OV L#,X;U@TOQI#=ID1UJ^"0I!5X>*S^-&+ X-
P]\ST[U@9NH<R5'W'Y@,)Y ]\%%2V;M^S"!!KELGP->7? A*FH$_@P[4P-M(_>2KM
P>T6<Z=Q2)9&+?.SC8Y^CC@#>DTI?N(I=@7T^,//SY=I#",\2HS6T)'YMF6FJN"V4
PR'C(FV &U"H$ND,$LFQ^SQ;%PN9V4<Q!.VQ1P)6>;[&>E'+,#K4K1BHI%G<5VF8P
P4%2I3_<3+BMB$@<QA$IGD)P>^+2Y_B]=K7I?@3 ?1::X'AW1VV>JT"SD_69)(Q4P
P2P@?=I'&=<K;(]9S%R!%4M,9$T15*$U]7MK8Y_Q=@N]C^V32+];G_HP2F&?#P+#@
PZIK +UYA3\X11+DP%@I.BO[F58P.F E"H8R.LF%]\G@/8#T_/ .IIGS]0_8C$IEV
PK1%EAO),)3_\K6FY;##PR .=G"+N A^D'X0<;\ BM>B_R\/O3Z'5"N]P"U4/O_VA
P@]XG\GGU^Y^#^:77^82FS2*WJ?F*X-D*#)W\J$T-[8GZ[[>+QE88IH:H-J@+78-H
PES#*9$WT#2,#+2GH_K>R/JQ7=FVNK-\'#'K694*(S/A !@6F<7<ZGVT1 WRNC.NJ
PGF(NHJE3+W1E QC9S0,<_SLW3E=I*M*6-4=IOEU1#74E:H!A6ZQ8YP^.WL0,!T*4
P#[YB!#C,VZ^A4%VR@->QJWA,!>6?+X5%@2XH;\$C>UK-MKIH;VASQILR%H?MBH?T
P2B"^[)COM2E9W[NU?5MO]!H6R23<S"U>,H838MELQ^4-.G8A41OJ1=C5K26O<\67
P/P@.4+G7-%(V?_'H?#!AY*G:5:Q\ST<T[%M<\EER<F#Q3;("RVWPCR-77)U%.'.E
P<DM7J^!AEW[=VJ-"3DN@>GV1$+CI@6;UU?B%I>D*U"'FM)-O22H\DGWZ:!F3+Q(>
PBPH- 9*C&#IS1K&TO:;$@6[OMY(VJ+14M(5,!<BQV'4:C)Y(6S6"ZWD.\(S)5UL"
P:9UQ_#Q@@Q3966S/0TJ58W0G9!NM"0DVT,>FP^3ADL.QV@SJP0I52O5AXT_J+])=
P06V[WP^T!=K9!2T6!_$@P8DH.Y>%)F9:#%[*WTRX_BMC_?([%I'\MBSZI1%;%_HW
PVXXS. LNG+=^#<$=MW."JR9=P/TU5<.^8"&,_O5)\J4GPMS)P:..>],5(C=8!^G1
P9$1^S$E12XJF.5N1]P2:24Y>X"D?1D8PO)4(W8[51J;U[]@WP(OO%PBF!&U,QC=>
P_Y.V!?7W)Y.FC:;/FPA,*]M$F\?MN9DE,*@U\>C@$XBD5D"D Z#MZD?S,VDI =8H
P\Q1Z8E8 $TKHG[OC%1\L1JG[HBD&,J&6RMLW9ZT<T@R  IVW.]3 = -AEB(4U5D1
P9K&T#I-1VE:>=98!-#1^/O'3.9W *V2@L$3J/$2%:*8OH.ZDRL92I(NBR^\ZR;]>
P_P[F(^LGY/_''+P">O:"\/X5VG3F/81%6LK?LPSD#?2I@*6 T.4R]Z_CQ'9&0!WX
PI# \V49/U#PUJW/I?<1B[%$ZS)'73O]]6!]YB>Y94ZO/[;H9:V2KJ,PM5A4A=BHS
PWQWE=,[3RE-*IV#IUY3MHS7)C2Q@;I2)A+H6;U-E$%F"!'R]1W:43%1?J[KKB'5:
P=]7^"^ROU%!5K5NGKLW3C2#!/+ EH73']HV4!66Y+'B6+Q9+W^U"OY@&Q(*9!I*Q
PSG;653!2O#=+A\H_IKZ%\G>!;@#=\9 XS76RU;A1YXQM"L>#]8 /DNLDC@-(S/P_
P;I-J7=K%9SB@5'%,H-BWNNW1R0P[K5B2_%"1-S3C:\^U0Q>0).<]#\;A_IW=(,(?
P*74VOP+02)=G#//#D;*]8\17F'L_)8F[]DC8?QZSSC*/CW9O!D-B%$0]_VX$>9ID
PXHWLN;)86>A-@+K^/(!]4&8JS3 ;@+)9CMH@(RQBQ['UF'QXLJ8UWB_50F_L&.6L
P@,M,J??_/B( Y,!W*&BNGQN]B6FDV^;&8M0IS&J7_KH/OC6U'@Y7%>H6G1(F^>$&
PTZJ0TKR6AX.73GGHSR/HG>J7N77,:^18PBXR3>17O>>ZT9_^3^ML3N\CQ^_\Q(7]
PD*YB:AVS;WR#E7'CF 2RPCCOA)HU4"+LQ8&J>DA=./^IZ1^A)&0?N!GT_;+CXY)X
P"3W%G57N??UE%^/C(C*T_.).'X.C*>E-7K.!RML=3@M0PTOME78HZW[3E$9/J@Q7
PY>+-G5^-X6T<NRF/>G$S+$5TDG;X=V06C9@M"9#%QY"#_!H!7<S6FD_HRNZ8_=BV
P4NEH6@VNKSE=<@\!<8Z@D"SFB^?B5'!5B/!RL.7D:/&T^UQ-JZKZ*TZ U3UC:@FM
PHS#NB77/Y03T"I]MHLZBMGOO<R<PC3LRKT(7ET@]#@I8G;.$_QKR_=Q:NZ[%J+LV
P6\\H1K+QVAL"+;RS,R"N+'C;P6[BP']:^J-@CV="*\:*@_'&-0Z%[RFLH_U +H2>
PL[J"#-SVB<EG,)?%VA2_J0NA.M 8X^B<QC6] C WI=[&D8/$W'Z+"DBXHR?GUZ=X
P+>J8^G %I>(/H-<^,QU\W,0W&AE7WX[<#J7R7NO""%ZZUX49%\DIX345:5;@)6QU
PFQD(X:"78UM);I:I[W<DB-FH2D,C>Z=#5>':7\IP</QZE+S)>E6*NW>9/> 8"P=/
PPVBP"9I0=0G9)^2=\]/Y"I4M3FN2S:C5J[80Q<]D!K>K%?V.([L)Z=QWX")1*@9?
P0.]D\#=\1*!HA8&1)(_2G-L*!:5T&5$:Q9E8=,6HUY#IH(2W*G_G/:>YEH3@LC$<
P=AAUE+6,R-GJ1#N8%LKSP=TT9"JMV=\(]&":.:I$[K!]-WK1:^X=8.)B_#Q 1(F3
P3,RMB=I7M&B3;.CVS^446E'G&F.@ML<O$:: 2F<$3"8-B?(JW, :OR$ "5.TSQ>+
P2.$H@0S5/+3DVKM8*0V?W:IL,JV/I-=<ZULX?!&XV! FMU>ER7&,A43_ZH0IO^1T
P;VH2V*7/)D]R>%0-C>D=M6M+P(CWO<7!WUL*<W[39=5R$H=EQ)DW7,K 2 .LC<T7
P7#][B3H<![)$79O]B(:Y_7.B!<;0LKTLTLS'9QF8_4N<-?G'JH99 D!4OH,52RLR
PMH:/$XWW!#U\VEDEHY93;G4Q,GT#0LF2.[J&0@6Q27C,1\L.WE,2D5,_#OR@AF.F
P*5;ZMDQ4('IC;'C/)7L>!GY%47KV#9U8X"+]*_^I?,?OD>20A56N?7V'NG;D!7A[
P+L#^X>L^I .XM_+ $%9V8-A;J<KO-+TB"V?[^XHWPVVX%@:KS L[Q*;6K$\V&R:$
PT,^Z5&&*_R=K>NW*:%HV75> &2/2UXBA*0@,G3$>X#6OS\*QN6 ^LH_KLCU^(&!&
PC2HI-C[=H-@&"@&M?%Y!<*:\-A^@'9G8RIMW\I"+,M0E*&V.3P92;W_)!"%['7V 
PKVEY$2@,\28'17\;^\_WOAJ &>P,:/Y2MIZ:J6X.[I&;__V<Q&L4O=D'8I12JS3:
P:MAW-I2Z-"\XLC.JG2(\9<%2<,IE24 *A9-%6S.36>'70>5I.I;CR?\LKXK\0RA^
P9)R*:,!L2.^.:T64I=<OI[,7'<I_+KY%_IQP@"^RI],WZ7<>*\6344SEY_DL;'J(
PUTQ(U!K893JWVI+5B<ZU%'P;C?,1KT4>K'R;V1ST#E^*5L5_891")?X,>6@CQG-+
PGDX?XQR2"]VWX-) S!GUT X:)88],?R6/CQ,=E6SZ&^4EJ_];S"WJ,#P7(H@5E. 
P^=FM0N_MC:U!",,16Q0]4#++ZW<^XP#,RQL%8^O>^6(X(IIZ0?%&#%2,,9CNC7!+
PQ8L^W;544#'L^X[XP9QU=[.WTO(!7?XP!0F,?:$;; L$N546/&T5:5=P2:;B+@TM
P49(9P;RW<YEO6DM3K$; '*]CH+SNLVJT!EA1![%(PHB^<,H5*]B[*.C6,)5C-.'+
P+D-L/K1D>_WG'T=:'^_RJW7#TQ'A))/BWZ%T6A,46WLL.H;J<M9H;T00I+GRI$X.
PK?<?&?5S]OD-I=,Y^6K:^DVHHD]@N9^7;R9G3.J3B%[U*'LYX:/?%&S@0D3.5F+G
P^=#'J$;$39E \":"K4NA$;$A+^VNFP_5JNQ;Q;_'0?8[540_X1Z+S&]+L9;N9)>S
PH.2X/@/5:6MD]9='K*F*!7UM71SZ'ZL7!QM1\Z(/6T+>86UEN(D#:=%A2*Z$+4'E
P1<IO9J0YZ;+;=>F,KF0- 2\>&:^+=DCY0<(%^>6?\[1ZPC38D)-<40BHWB-PEL^8
PNJ1;*QT2B% 94[D"W"F-]V79MTPF[CWX^?62T!628&K/#7>8,L0ET6?B=3'>!=4W
P_EPN$(^44A%D38.N2 M3-O&K8[#,%$\>.:@6B_C8#<HG+2J)^4RM2.[VD[4.$+Z.
PY:Z?)Y@M9JIJL*_5L(]#[7V>/?^N_/AKDR$Y4J[F#G7&WO)2PN;NM)"H404ZZ!$+
PD1C9&!$%:W9E-6+&8-I>LYKF:W'V\XL,\&YPJ[R_),'9L;+5:0IJF/;>BZOT%\@W
PZ!7N0U^F,S/!6-#7\]694]>LK)!I$\* 5#HP\]2657DT6'/%9H2LN:?#R\N8L<[W
P<L8.HYK(>%FWJ/9*8ZW?0K$ JVS.)[]:D8.Q?B*NEJN_/'Y?48JNKUBA)\\FCD0@
PAAI;H20U->C!1NCU0)B=/6(=PMLK.!RV*U_8T_^IR@?GT%+:43X2E\]7=Y&GZ!(Y
PF[&B&ZVH5+@J!D&ETWV&$UZN&#F,'N7P7PEI8A;PAL'&I/+L#AS@.7$>"N*5\?T3
P3)R!SN?,(,+1A!E2U%GFBA6S0G._G+B.)+"V]B\:)4CVLN_XYN_=/Z3,GIYZGBW=
P2'R9&''E!+[V?(0]&]2MW^<""V[Y%@#\8V7I9%AQCV3/$SI*I?709RBX_QV%*(DI
P<7E$653QN6IGS._ #F "H]>S[7 _+/&YRL/N(ED[UX?]C6(<.]6]4;.^L]L2!</R
P0F\O(M=BQ*5].)G1_/H&51+/2N''R*@PS\Q.(4?T<CA?4*L\%;) D9Y@,\X'(A#9
P$-]8^I&JG#A6]?E!F%>3:JR0V9.*+[Q5-A6CBMF<77NVI:^4:+:YCST!O^F#!V>8
PXB9RDD(9.&:PX;5ZJ#(URJM !6PPN!'BGWQ%X8Y.0ECP<AXQKT>-WYY+.Y&J=H$Z
P:8IKYI7O(W"4Q)IQW ^F@M=DP31)FF;7U?6PFKW@'R$],.11)J'FKUE ) )8GB*_
P1PP*5*8QH7K#4 0-0+>?3(WCA@5!!,4P@?X+T+R%"TY$R-E%?4Y7=FJV;0MA":KT
P(?LUN>'5O6Y"[&=)/ZSZ28#GW!* /SWN<B];9;KSS6,KVAUQK[_3ZO#8 F4A4F4A
PLC(P"SL4$?&-Q 6JWAH0NN8<\"QK^!JP"ZTWQ\JO?=&V).M#%M<J:L,H\(-<_X&F
PI+E5[61A/?M PD:[9J7 E5XTA^K)V;QE/:F_6/! 9$7$@3(,%.B-C@,""- IT42#
PHQ0,LF!ZN*0=E4UXAIA'2$U:YG=(GN[O3KP\3UH%H.%;8W?H!9N@%&@J> =Q:[:4
P[AW, [!%C/V+?*V'1TV\I@//?[Y=D<UDT$7KW;#+^H@LBJ[8*=SYP&<GS6KNDIU'
P=].S12I)V@/="/!WZR0$.I/AI0(:M=5G@'>L9&[OD>(<>WOI[5;.)W%<6G+"]D_L
PAT>N1P@J)\=A1&/,0!W"->B96EZ3[%=CS01-UI.-%,^H)3,J.<)T9 Q*3:VV@1]R
PD&Q:=Q:CSK[F'9N%""[,=QA?HK.GH@XF W?CA#O/2*J_SD%($Y2=%Y1(%W+Q+CDQ
PBJC=\7$7\C@JY\TUL6:QQM /-X -W"\I(&"V>^]B6DB P/DED?S.;ECHG$6440[B
P;+ZZPK+5@;QJ3#=W]M'X;2PUNRWL',T>AG4)Z#] >7<CBZ.80%*#OZ9=DE.9&F1&
PML]54TC+S1F"9ER%FPJHMRH=TXBAG.!LVA7?%Z>W!5[F#$Y#R5$!Y/%*.K/H-VU6
P=2V3BN#EJ96;7.5Z4&FY-QP?>1%M<X,=<\R28E)0,QVQW(=\-6$9D0O0*KY=A4&R
PY.@0+?4U2R>NRS*#ZRC0 FUUB!O;IY#,"GS(3KKWSBMUF&CMU2@E[.R@(,FD49GR
P72?Y^QFW9T'4!5/S1\+TDO)F1LL@9P\P>SF*%UDOM?O@+;9[+@7M,-%.(3T:@@1U
P>RC[*S>?MZ0D'OX@)WJ^SK;6DLM88-0TP86SB^VX39=^S5 I,&%;[?&U4)I.53Y^
P >0QUQ'4-["7$,!CHXK\6V<+FBMTR47DLM8'SDX">Y[7HP"E.]Q8$[5]])@L',G7
P1L)&:/+GLD;)5;Z%R#''P/S505T"XYVAC= "V7JZ_84-.E#89T7>7LEV1\3$_F&R
P=^%UTI%2[":P.M&&*U--3,E&T@'MF4/KUQR8.Q+-?@^-S"NTD+9]=ZR/\:0K7894
P$V<%?6S. M$#87ZT3;L%\T E,PYL7UP87VMR*%GB#2M*'[_Z>]MKAITL'%O_BQ'O
PR@62(<5'+--!98]"4"[P%'X'$=C.2,8*A>++I'>TO0)'\?'@E82<92"48?*R$]:#
P@F/HB;.O+=00 Y/::860:@]Q<'_M#<7ZN0Q;0T**A7^)H2C&H.]']0?;.O#;?.<:
P!82D)?3[E-\G%_25WW<W?F#;3UW'%,5PT:@<)IA0 DF6$H/(-@:E\KXO#++WAL&R
PU03=XST^KI9*\/E].@Y[0+/<LU^9.38_Z;@3\BX0N?"*KJ 4J;;=*GZ):+"<O6D0
P\6%7M<!'BDA -O1V):E _Z+AYN0A6XZA@51\*@0T/:)]'C2=_@GV66=RK7FLQVRG
P(ZM@55 ;"*EVVIYV+1\:IVD3?4@!]5Q>#;,7Y64OC+V5;.;R[EELH<4J[XT;@:N6
P9P3Z\Y7UW[4M.+/TF7@=]WI,@%KAR%"9 Y*U$QVXXRB>@^'Y$&"?0CU_(RM.D)"Q
P:$1X^XUUBA<;RZH E?DY"G__A:4B\0;$3D*>, JW0T'TVAW'OZWRZ!C+\>6W.6]J
P@$4?@!4RZ^>:0JCJ-@F^'&KNI#5B^+(NV?M<#T+-.C7(P5H+!,5 2B:+NK1'A3RO
P<IX*XQ,'&3/>.1R=;F*(6H4ZZVZNQJ<Z9S%[][)S$<V!RO6T>Z^6_(;1@OQIU F5
PCO5'Y\)1_SG3UF,JPFMP_^R95:B.+)8,HP[TZV%=&/8"W-4&N=>2> 2?3FPH^")P
PF&J6%V=*1U3!"Q_"4)A[U/&ENN%[6M2%_>2;>M10S ^P'9.\>]A!M?$KO3Z=5C:<
P5%UDVV63NM;/ERW@8.C&_Z1Q&D3^Y_,3]A9QWOI0:H+S/1**<GPG$6ZH>P[$FFIN
PP]KA&I!>L8(#BO&3WR $0)+SV[6%%+&=AV8;]Y')A<OC=E]Q8Z1]X.4P,ZT_0AB,
P&89%]MR2@W_."']?5S3%E2&M0%,',G XY"8[C<0KB=*=[?.8W+EL0KL]&AY02J\W
P>2ZQ(9Y^&# 0D](C0,3*:U>_+>]5GZ6(<T!*I(%-H[JJTNS'#GY.0I!<FY&OX"-9
P*@C255M=. _T,=JJ=M;24VW>LVYO# :BQ29OHR<46%GYD^:E+VFJA)!L<98*W"^C
PB"'RLL.I3]S8R2TS9_0XN I[."K-=I?E7;@)QOCVS::IC4W8!$LG>+O#[T21*;YW
PB$7&E,G]-C^DAG>/H@4U.ML_YF,NS2:%_O(6KOSEDWUT@!I@J +RI@Q >Z%C.IU>
PNK,OI:7:_+JZ^=0#%@47:R'E4<=\-4O[ ;1@=>$%J\,K[3=,:M-G-D,4RA88BFO5
PM"PW'C?\FV79(DP+JD+S!&S%'LO.>7L7J8)'*GSE6^(0/B[MG*=;BK[#K2]<(6;+
P76O?]$7SOT#U0=5A,,5WFLD:W*0A-RIOW+/WD!-R-9_>QEJ;_S(KYRM4+@"51< J
PNQ-*ZAE.'\BE;&D9'^4KN'O[BL02$W \X*B-U;,D0369R3N<<9@?OCORV+$TD%71
PBN3Z,$?6/!,0!5%89ZC&^0L]><<(Y_ W&;VG 5'Q52Y/X57<3-DE9Q7Z-R,&_D-Z
PU2< H*XZ]/I?:25A[@&MJ B-*NS9[.CBS>F*'E_-"GK@@^9H[/VCVTL1(1UHO.:_
PY\A\)"\CPD=R:S8UE#R]E.7I8/SE+Z!TWY-=R3=&'X0;![Y"K5FSNZ.("D1=2/F6
P<8-(QHJ*P6N1+G LC5KG*FY\VQ =E6DA-/%^?#Q6]Q0D[*SL2R,V&?$N*U9<)BW+
PK.Y2=05JS6*1%5WQ&X'UAZTB<>? &!0=ULT6=Z_UO7S7,:;*23:_T>3C=K!Y"1U5
PB-,RR1 1-REW,+7SW13'XU?M-I%P^7>9(Y%IM(Z_X7YAEQU,)/Z"/2!_2:YMV1CT
PG<8$=FWT<$Z*ZXAFD?"Q2+84$J+U4U'B6K2=V&&X@FU&;@&88-V?K:JK$,?YNKK+
P=,!?!BE(E_9*;GKIH*\-/P%=T2S:E1FI24%@W6A-8[W";T4DEXG\YX$^FD+<W1#4
P6Q=X;+5U^N4FUE@[ILJXYQ5#EN&+"P$JTGXG=.JFOJN>+[L/T82>1?9YJ3KN8:U<
P6:76[_+I/ $K@A:OM8I6J(*FD\+C"+OFVX/K(GKKM40-4 ?:7 ZPANH#'E-O3U'!
PN9FL>NNICQ8H)M,:(24?1B7+PF$%Z\#(*P(]R_*!I)$XP$FFZ^HUG"MY><+1D_P1
P9?XR[BQ'+Y6\#T[0&T]C2O4)@&%C?^^.G-8:EMO 1HU[MN@L_T\DZAFT+]:CDO(X
P7&DKU[E&@OT7UP@?+P/U21[WX?UN CY]/YX$2#LZ2@V/?<=HSH,;HAC;_QCGH)S&
PUO>M)MO")!:=]=&^OKC-YVRHO4XT*L98Y'N$*TA1QK1D%>Y&M#@K687[<NMDS*<D
P?'D0]@BE=7DQ&N<B_S"U,I&:+GHCLET9HUXMY_'.;*QAVD9QWS'9!/!S35Z8I?S\
PSP.4[!B6//$=U?Q](+3S\"(")!*]2X"5'64+L^;*, *4@_&]U8!NQP'Z'?-6QX=[
PG6T--8/3S5N1S'>8TI@B(#M:C20(-1\ @-R")3(M,7 V.Z1N$#V^4_)#V%I:<?\M
P-QOMTCD49WO+<<:(KO(*4XX/@P%G>=;]OCS"-C(X)-)NVS#->MGA%C/#W83>NG5J
P'6I[E'/F@\23OT]88MX+,0@B3.*W6\SO;F?#,'(E7B6,SCG?R[;/I[+Y0L$>/D%-
PNCOU1B41.M^U:.S-FK[!_*:Q<&D4!$$J3=#FF*;1V"Q- <:6K3=B9-G'ZKQ1T*]4
P)R7P_BZ39=.5GE->LF$]@CT9_V?0T&G^QQ=30TW#UH+AI6;%2FN >J= !.JV]2O-
P*;"CF$76U\E_!V@HW%FJNE2%7\ID""D6[JC7["R"2L/!T:D%S:K7-Z0IB(T(\C'7
PN5)(!*I ;.>&;DXO[]\E+8R,BD$.CL5&!V::CJV1RNIV[RRM@VGFYLN&8(#EZM*I
P"HC\+3XM.<I>+;692Y& .HTH"V=@1E@WY.-_3@+AQE>$^FKDV9<,;N_R4\G/-<^;
PD$C(0W$W= 8$QSHX6P.V]MYMNMKS;K>E>2;0>AU.]-:!IEA4G#W B2X'PQ3I)-C,
P1B*V\5^H0+:]9**D$<H8BZ@1.Z%#:5G$WCYNO?9+8'(>3P0+$&:)*QV77>*@GSZT
PPC5 9M79Q#[-1OL:J'/:)=PS9#/W%L&/F>5[."?X8Z<WC#W%$1'TF+(2JN6QEYDH
P$M3PA<4N$E^RU)Z+4DX__S:2[HDR*"N< -@,CA/"_YKNW)T1K9-TDPKY=K*&SP85
PET(W=ZFAC)UR'2@7!$K=N%GF!5SL]LJ2EGF:WYK;H\!:/%_7$MBTZ)8C*6O%P1K9
PZ&O9-O]2OGOA1VP)G+1HEX.!@E!JQU4/'UW&3ICH^5;<_;M?AXA \N:XM,*01:T.
P ZA2 *I'REISV;&[MP%*M?"W-32)8:%_+?P8!/RU';PD\+J-M)V2#9Y4S!!T1()&
P]D$/7PQ2=T,4I0[@3-/Q]/EM/X:/^HW&4*WYMQ8_C&KJAH&-]2[$BG4\G7?N>/?6
P;(T+Z<#@NZ"IP<2A:!-O-XR6@(KCFW-?D"3??VM[^.<[Q7$HJ9JW<$F"DV[V.SZU
PD,3[D6,UCL3; 13;6A\X;1W?3;RY=9U8AX>S[H2>12+20E<9B;1[7?A;9'!W3/Y=
P.1&@*\S.8/(Q$>;%)Q^&S#WMN(FF#(M5P"/'&](G$0L.6]4GH7",%Y<@<*+*;2D/
PS<3J%R+%-%XD.%_+H.D.]&A12KD9]2E]UXM(0E*DZDRL%T?=X;T9S]4<=VHB5N0X
PN^Z9$"WVMBDKE2C<:'#1KZ>86N82V2&D,A!9XPFVR#58.AN7$4Y]KVI43H3D(P_3
PGK)=H$C+;Q'.PCX7+*9OI04SQXWB8)GE@-E+1LAF\#(4JI5BJSE^WN<0I-M<[:]W
PXUB:I*G=34E]F6&,IW?5=Q63& >YQ40!DL@(.TMM*B)MILN'TF&"E;,9 FH1[QP0
PE]?'KZ>6CQBJ:?.\O2C!.X5R>PWW]K)M.>]P0'5NTZ_V\%L%+8GR'<*%)4=P XQ?
PF*FF5 ITE _VD)4%_7A9=7I1:&\4WX88P"5U(EL]M;5-UZ< *:CD:1?KRBYH2@RU
PC4&P!VS@6(SC7A,L*Z'@W_DZ%"'+D<K:I,HU,//XHU@G8=8Z?0=\Q6_K8&R!Z2TX
P+C:!#2*T4(CL!3;QZ[G:\+8YF..>Q#13R@BBW<^.M2 25:.5$VM<M(1Q87B3B%1S
P=)6&4%M8@I\Z+,>$^]SRDQ3ZP6*?3&3Y\(F!3H3?]70NE["BHUH?"JPI?M^C2F%\
P'@>52Q.(8 Y@Q]A+Z:KKZ'2*2_G;TQ#6:T(..=Q\=/YU9=I:8BO]#SK".Y+61U0F
PKKAKKZX1+7)8Y0N*K;<Z^FF#UO2!(_O! (U\+B8M._>-C9E8'H7)):Z;8-A5);GP
P\3?2KE"X)17ZZX2;V0[WY+IJN'U&1-:WD4*72PADIU6:5::0X@2,/I67GKS"9#A^
PTW]Z&F]*,($GX76JKKS+]J01I5I4G-VKA9C:LX<Y($-YW^4H.^JNT*]D;#\W'74D
P*LT[-Z9*X.ALJA&X#YE24F<\T-$I3\0:M"!=\=)N/BOOV<^.XZ>SM,_Z& R\SDW#
P9)A[K?TG?;G_0 _0*-[@J2]: T1N2T!WM$K ^QXQ,L0M.Q 70*DO'!;*SSXK4K7A
PL@W1G%1#FW>Q2?86F3XE4!B<KBX$TL&BYM]BT.30\&,=3F/NO: G+6;H"!8O$!!!
P!-:#S(&8Y?H<N?U;+S5_@E2BQ3JE0)@8()"M9'_"OZ&E8\MG7X#M*Y<X28@$QZJV
PO8?)'%DP#_W\D\KM0J\4<+G49[S%G.!>PD6U0HUB\Q/!>7N]JN(FW@C GQ6OCC1T
PI(VG^LH>K5<Q0UX+I[Q;P5P8QMJJ"@<'_)1GKOVI'0<*9_V=O=@N?8\5R8@\]@(^
PL-B1=A_97-RPL&1FG4Z!KOBKJ#;<79J&!PGJ)>MP !@=L5+N^)Q$.*U5Y<@5Z/;.
P8+ZEFQ'\J5)@MAPUFPVS@KXT_+669S/$6'L/@^!=A\O"(+TX@$*]T+A7[\13_4:A
PEZNQ4Z%ZO)GOVZ%J+*A.Q.A[),S8G.NOJB5WWZN^[%9X1 T1P=YUUFB^71D23'PM
P13GUPYLG9]+VHUPOK]-M+-+20A$3<^N4"_P4 4M3^= 1ZN@%*+/J!M:/_2EXFT7R
P__*%HAS)I;D*=[C)L3ZNN3CL<69CN/I-[;N 8MH@0!F _]5OW&>G^]N\@@$/=:__
P__=[<'[R1C6A+V!:IH&_:!C-!?]_Q\J/7%CGQ:^1+X(W#Z!C)(_A]CS*)^:I%D\&
PJ:QY?M=,$TZ#)DSLZI2F>F86F>>($N%*B0/]3KVJ0L9+E)1'0U;"T0"J-<5&K0I8
P>V,KP?Y]  HAR79[-]_*Q=2QM\.<])0!4E]$"BXMYM%P$FX,4*5D ,56P6@+2G2*
PX.=4:!!&1<&'8HK["%V:=GDF2R<\8O BK?:PMD*B0QLU/ *"ZM>D7@*?F-BB6"YI
PYAXWR!IJ%U#=\=L*D.Q9$!(L$7R<@G<E3]LGO4N86XP_D?>MM11J!>,>K]#<+#@A
P^^<S&'Z!U3DPKIXQI$!\DJ>-G/I4$2S 1^BH2+@/%"!+L%Y$W#W)RC%JTV\\F+ID
PA4!"P6U"!05#NUK(8#11Y\&@EJN#@N'PRTS4V.&K^;L/1B6.#;:5*<5X4/!FGRYT
P(C3]N/BD(TZ8[_2"TLK,C2'\]K-G!4UT_:3.^M?J_39&<J(I@31^0\^9&U$!'^;W
P(.1&M?.KE)<5EG=<X#14]BP72A+75H<R@-B]6VTEX#+]:I+=Q1:@OBUZHI8$NRWT
P LN%_;I:R]BWQ?A*K-),^K? I,%(60HC*I<<'S;MK!\.^K'AUR WG6Q)!9C[Q8N8
P>09#+0S?O>;FM-YO2PB>N!%R["X[PJEZRV7J(+I^?$J;(V YX<.'#D#Z=2&_F(-Z
P(IL]M_BPXKV*_BF=]YTS]-7X;;'@^0U<E G!_28#%)#X5^_54V_C;_)%9O'0JQN>
PBQ"'LE&B>Q;"+]EEKE7)870GJ.-"!EH/T].[!89TM?DJ=;BC'M?NC"85S^L8W'E,
P==6WV?\8DJVR'$T@DF<JF\3LH:RY;ZF<TB7&O9/XO#*.8XTY- K:H"ZO*U+CUG-/
PY&Z26.1M'&C;:"G;DN)Y+J30V2"BWF40\(M X2"ZH]WYC3044P$@+Q1PT<G&4<?;
PWB=[UB'4&/S7N-D@,#^X,A.#+ \BW GWK\+W_YZ15RVNV?P_%;F- .?AQ/;L#DSC
P-E F:GVKK.A+ODG6<4TJ4Z8=(X"6$+!V@2G_Q&N0AWQC7BG(UOK3XVKA43^EW[VB
PE?@$.P-?#*($5*7WGQ6J=[!PYZKL0WT\%8-UM[RYW8U%CH-]R:M+1=I''UH%@6&K
P+R@T--!]!KR8NG 1.YU"1&X4@Q IKAJ-LEB!1'$:85U1PJ/KXBMB,183'*GJ8.K7
P0MOT:9S@V)S8KF+^TWU6X!!LS8E30I*C4B)C1+Y\K5<%.&\!I#GIN"KJ,9FNN;>0
PBZR6\K@COIJ4/E;6&BLVD=[SC!/C>C_J.I@0:X2<I!9'NMT&5)FM<"<4T:+##Y6I
P:WWOS62Q!Q4X>PPR,63J,YHT8Q8I%)[.G(L[;3A53<X7TG@NV[KZ@K;!/N@,=)PF
PENSC@DU:X(<YY83/ %!O$NJ4KMQ.V7?^_ DU+O.]/4 L3]=B!FZ\;W_W2;51^M#N
P64&,XMW_*[OXS^\P Y\4?BG3XBQHT&24HXG14RA8M\#XRW)V)2P.7UK X'*AQ1#'
PMT3^33@6ZX:?G$"!%X99APS<8QZ5LJ; 8CH924V@Z%YHCU,/1RT0-5[!U"X^W4NU
P&.$3#[VX7,3_I=S'*A>C7_CD[$"NVUTI-[ &&(3;E2'+)5\Y0J7*$D..4I@_@=;'
P.V7!<:538]>R%Z,&:K>&'W<22NRC)Z@K9BXK):)%WY@>+$'] +BH[D[@#%*$BL%)
P!%"JU.E,M0VCGJ,-S!1S^<(!O-]\P,PW; U)[&$C HH[DE-K-;!.1GY;#.34 A94
P[W4U"^J1]39'0!=H\GA,8&KKDM?,)%MSF1H$X/>L?_XKE6XX6RMOE.ESX7;%E^O/
P8P%0J*KT<EQ:X0?!L.J# #1G72O7P)6\)1N-@)&V'M XA<EQ>K/JV^UL1-4L6)UZ
P5GZX_GC6+TNVG.S2_\7ML+\$%#OOU4U.$:$+@^=.P5G D_GAIT=D>UT#[!J%5Q0S
PN5@J7FBT>M!]:>MA;YXE;H8(!&$8"^9NM>SVP?24XBXMJE@IML-V;I^_]^SP$HU3
PYC3-'6B?'>[F-R[+<W[,IV4H8BFK?!JMR8DZ3W?<=!VF4A:T(X:V^7%8 5VT4VG&
P0?M-_316C"ZD$GZ-0WD\[U+QNT"<&!Z?9;C) M5X20][G<9HC:;[8[X"HR[N,+XL
P$T$9)S,+G7H\]@ZTX@RIPQOJ\FN3?"73^/E<AUS#:RU&>D=!T0.$'0\_2[P?S& D
PTH^H!X.M2-)?3KTS1WK(T#A\V9C\:E50@_S<Q[CO9=F*X1VQ761J]H3!N]0P=%FL
P!?4[2*PPM*.&$KUU<5<=5]BWL<7K:VHF"&*-VO +=XB*IR<'SDIO4$N!QP1+&>.I
P@7,VAM??I5,*FT/8XG8 9%@5N][V0@^7_D^V(MA?FFQA[+O2J%C!H+0%/)IY;G2C
P C*@&@K#OPASPEL^1AAN#>/W.,@B;DVB;TB<KUJ'M)])ZK*37SN!.MYMY10+P46M
P?R)8GMJ"#.'U#+\*@)3GH07FWPM@_SU/=P .O0>_F%PPC5%1A5L;053$*+2"C1^G
P]FX0H3P]'A04"! BO\Y73SUJ-/E\:;1/7L=IN';,T.:$;$]WK\CJJER=XM1YURV3
PG$WT&V5&@J:A=$U]0Q/?'ODZO.?Y26;?R_Q2?U&JFL\2VB!E>HDQHQDR7Q.P:%@9
P/= RK27+U[UKLP/6CW*@19?/@#.R,L"@-*B*,%7/F;@FE[\S(4QK9NKJJV<16[J\
PE$<4?5P;:@1[\W\]/6MP*)BJ&0>^YE_8)2PP9F.JJ!CY=_T,!)\Z=[UK/&;'OL5]
PT2BJ@YJ=&XM9H2B?+1]I@>3KY*\7!FK@=@E#($N%Q#W?UE*CTA1A<%U% 9V%/T[@
P$<H'PF9*^E1%Y(_?T-W> U8E^*_5EU>L9L=*W2D1;^N5!49: $1UM,9L'SU?M^+M
PJOD7=J'UJCSQ%I<4R1"=GV5<4[K""W\G*- WP2K6(QJ7LM'QEPF.4B?SFU;FL%VF
P*3=%A7>K<.!BW?7N+@DU!9XJ+D]E(;2A8XGO?\AY1JS'3#@[-=]GWX(D X_HP+=Y
P^4B'&CP@ N.[Q^ A6]_7=8PU(?S-5Z-D,.\T4SHT*R0RFZQSHZQ]$(+#\(!R P4*
PS#(6# ?_KE<&E^=%^35=8WRKD],+'M'TA3N;76R>N@/U:BMKV1IXX6CPRH_2$2PI
P\7#:,D351$.>LKRE \POY<$BS> JVQDQC_*Y]P:(7/I=W])R\J=UV6RU;A;92"8F
PW+[50C,W#Z1HV0-)M?!&%_SY:^FK4: _15:>0@:K5W*6 K/&]6_;;7U-UUD;"V"V
PIO*I:DQZ!ARAG?S[?L<@59,LL4$\?\3K/MKU:1B^S#R8G+^3:>*TC6;E)?1+1MA5
P9"3"6XEXLP0VFO[0GZ(O$XJ604[J53C*ZUU%UH!JHF=QR-("N4L^2"5':!WF'@^H
P&[?<7A(&BS D<NX!C9$(=:O*+[8,N:<H1>&=$^9PTGM0S!RLS3\=*P286/991Z0!
P><,<04U[3I$\ 9N,;[C&^',AD0.;6XSZ*NH'0"%^MQWB#9%.7 '">U.2$2'8ETT=
PRQ\M4^# \_KMF).6:>/] &LB,5K0.X&2;J*XWZJ>]D3!%VPKX)4"F51Z.[@+A'O9
P(!WZZ]]E$;)]=ZG=WPKJF(KF*"NK-FU77D.7KA6Z"V>0VAWN<BLG7+UD17R]VQX)
P#;F3#5(8S@H"CX>;+Q'"["LBA6$FF?]3;J2:YZSZU+N">"MSZZ3THI*X..1@Q%#N
PT>>O0P4WC$!:$C'/UXX.,#<D,'R#>5I<8:Y3E_ ,ON9U>W@XMY XB4-JBHB'O,S@
PQ3$7H@5(AT/>F^A=BN&P1[K>G!J[BA1B@+Q9@PQY,(;254"3.&YE'[ %M&2@J'@R
P,+TP0PH BBJYB,>4LFO5^0S@Q&X/"EI#C 6[;3>?:O;JQGDGC)@N+][.9G>-YN\J
PV//9 (C'6N1LN34:=M*BQ8W.)$"EKGZ]K^04P&B'B=H*XZE)I)&[,E"3YW[N_A#P
PHC].X+LR@#\XT:V\OTR$7$S=&@W$!3%<B +3YGSJ0T[Z5(]N:H3\]L&X+^H.9^6Z
P=E3XX9&O .*,=A*4B>$W(?P+MK$_?P LX")FI)^*&?#A1G8Z@A@<-@BUQ4RC)5^T
PD#4026LE:#*:TX!!>AC]Y)#:W'!>PU.9Y+*"S=Z_?O!=\%WF;M/&!S[T$F?#N3]N
PHQ/I\B/*P7<[%\'4<$G->3TFI[UY(:G[[T]'EPEF#3FQ.DAQC^!_H\IMA_ &1'#>
P7AXZJWXG=B"-7KR&;L<(<T3:PZ^W4:TWMVWO^36[M2(MN13I5@!<MY^%B]DBAZ4]
PO W6S34]Y@@)?!ZUHSAT)IZ%^WC187;]C084+)L%Z!]1%.BC3<O,F/'ZHAF& _?*
P(=$(8Y*8]!!UQYX-/U:0R"TY804O[,WA2O;[CS0G68;GDCXV+T]]>CT(W^AB.UBK
P$VB&0 XN5(L64!=!ZKS+UYS6X1VR(PUM*F-&H!!AEKFS?=9EHAG<&*T?*7 4._K8
PY;D49\7]P< W&FQ\FNA8KC=6&L\$9J^79O"MZT+WPQ9P/SC(;EQ_=);NJ]2!9BVP
PUKDE6CP#2E'1Q4-KTM[VHOOU$AN'S387,WOW=T A9RU<922NHIW0/0= T=/,%"^P
P*8DYX$V/,> &O"46[%1#ZZAXR^H;!5S!YHQ G*O&.["#M VEFB&9YJR^D'3;.1!$
PE>'WT?#,\.D>/N3!63\J\35V=LN_76[(]/7)@=D$%4-\&BQ7HB573E53XP^GS(?H
P0O(O4E4$\N#9B6T5"K:X(@?FM^P+WAOUT5P(B%7=B=<1D38'9\D*&]^-:1V,N !<
PNVWDJJ+R>C@$ P3[/M(;#"V=F%9)V;IOT\EP5.ZW<=4E *>^M]7*=B#>IR,Q=#0.
P?M17SS*E!#0(VWI)+2PH/G9/2]>'0789BTKO@4P11ZDB@D7*C-Y-B%D+XS5CPIS1
P'P=_=>#$I:N:0+R%K;XXG0_N3$([Z S!<JO>047U78.%.-YY.G4/5VO5_7D;AQ&?
PU%_\$3&YK@3'/4"@P<5V3:I],1_=%)4796N[(I]2:.W32ZH&DW.9K%81(X.Q&.S#
P^ 4@>]^X8@II,?<UYQ95J>8*.M0R5A="."NH+.&2/T>*0.D NDE$2E!_$TK:(3@?
P["Y?,556WD7<IK#W^-[N#3G#ABCREP6Y<8&(HZ:"FOP5F%+TF7$@9E-P670WZ -J
P*Z/C'-P731/=VZB9K+?B+]U&5*-WY[$+U(VZ!8CVW*S9X+%O+388]+O@\IX1F6_4
PI*844[O_NGL9U.1\>9XYC ;'F\MAB.AXE8GW^=D"?/0Q>F]<,)FXW$G#S06N<>Q<
P-CQ:==\Q5+4[NQF&?H=0LS%@R"YD_HX(M<Y=$0^E:]%MI2G;WV^BB*Y-BH":@HL?
PN2\]1XFFR#'/BX4+;7";P::D%*8N?,])<WS_EXQF1%->BOZ4<WJB>V;46-YYF5<>
P<W3\TB2[BJ0*J7.2\J:_+-YNE5H5B_Q)I_7?$ Q76PS1^G&O[D'Z$&8RG[, 6C!,
P\V'_M%>/N\'[B2@LNIQ%>L:+#ZWT&YL^H L0^^JKI37[DW&I,/ >3K".:U0+%TD?
P;^-Q'(FM[,X@_$^T AD0X;PX3N$:=J<D#(AH$/^'[?^\JMZ_DPU3WW&=!/A %(?-
P'EMFT8<E)2-&"=ZSQ#X5T5+Y(G+JO#1CU^)@EE-E9I9U5Y#L']I%# Y-H@_E7[RI
P,_<VDFBG&&V!QF!#>4;^<@'*HZIZ**K<I:J(V2.:BV]Q7B3381!R^-" ^Q@6M%&O
P >>1$]G9DU]L)MI=&3"*\.*B>5T\/^D[,74 -_X=W44$OX'KN5V*]SF2)1TX6?.W
PXX$5\;5I/$4PRVN:EYPG:RI0W*J/3)$?WAVQ%^0&8 /-8#L[24E>SCT5/.M/.G4R
P%8P,##I=IVM1G9L4;R2AQWDE>U7:T8O/BY]&/5M"(IU9?)^FJHI!D3?Z2DU,VJV0
PG">'3"TW\XTMQ7B$:,[PP152>IHD*[*\YQ)[;]&!0C]\)F^'?]=UU1MQI?8GKFP<
P<;-19GT+5<'ZV%PI^_5&=Y*=MZ&_+4@5<.1RALWIJ N>-[K)IG1KITS[+O! 4NQ\
P-U$O!_H 1*8NK;Q*VKU&/[4)S?M:6>ZR6ZO JA,?7SK[LM;NRFRBY3N?=,#+"?\[
PP;L2QDD'OKL?%'XZ^!P6S'RLSFLNF6TNZUO):<Z&&)_8L<P;;/<R@%*#=AHD^5ZV
P&/PL[AIWMU;.4J11FSJ4+X1FT#V9:^7E-$A[_%_*21!?MRK@X,> W^N0AZ/,$TG;
P0\63^YI6T/NCF\E_A.<0R4S00]V7WQVXRO6,7'KB<G]W74@P68#X9-SEB?E$^^OM
PPD?*1J'0\ORGO&R6!+ #<"D*14=%$U26L1RMGHXL)O4BWU:5SX1:;K<&JJ!WO8*K
P44 ];/X"%PFO&$5.0Y(;@TP]ATGQCN!R;'VF1^[<F]:I$:BN#'00@BOS2VDRO 0)
P'R@_,_"#P)H8 "Q6D%,.KKG#UDRXE2(+!C.+58Y4SY%#$BUEYE%CT%1$W#6-*.95
P,9W)<0NX,&BFM^E.@=+8@BVA4+JBE31EW9$B*TR#$/W3"/7U""W;F("1(6//SWB&
PW5<>UDHP,O#^!N?ECA=T_ "P2X_<%P O^=+C- &%I.'QP5AC"WF3TW946N44.<'"
PN3ES&Q!;<,"@B[$Y245'3T2 //<.K*>EH\;'9G*0L.@_\$6PB3KYY@,&D7.5?^\5
P,WCFO-5X$<>9>Y4M$$1A/?",W<&@ S".:XCH&T05:I-V*+K+KH7+4>-[6R_LSX$E
P'>%+1]]$\IACD'727E \ [ M!&YAE8O35"MICI7&^. ?.Z)868JNG!M0.CL.(H.I
PG8B9W0EB\I)B"=^E;?U0KJ#,,HIC,:FV]3J<6#8K0AH,P-Z<>0K=%=%NT.&B,V(,
P"8-KN0TQVNGYXRWUSK\ I@!9:0/ &4.EX95W:__R)B,FG,<W\(8[G4T_*K>)2E@:
P02%B8FMK(#=6EMC+K6MXR7UR6#443Q-]M<BP>'I-:7RPPD(E&RLXD#L=0^Z\T!M[
PP6'V &6&]#WT65NO R;@81EDBMH_L!&A=+ P>.Q_42<8E2K[S=3V^M.U1.S&$8VA
P)(_!1'^&UN)LIFK'%C*<>B7M$4/@HPJD<S;I\^4T'OY(687W6PN .%77FS>VS"M"
PE<)?$MR$<?Y3U0.R[.GI!.+V7WIK5;+!<5^CF <K(J!FV@B7>V>%RFK+;$0H,W%8
P^DY7KOQY+;2GO!Z]/T!]< W.$<CL%#$4MK$X7-8ZPR,N;'<5Z-/^OPHQO4^[ V63
P>>:-P$*Q\)IFK?K%&5IN4H'./^E2CRLI"Q09;!=\\@82G=,$,GBJ>%(JG',$[&)G
P/%+#8UN#YY29T"A?@+]9%U1^="MU9>2K]503,>X&J%9!+F<N&0.,&K(T.)7$6.7K
P7B JM"O&["<0XNFZ:+'@G;5SX@[5H0%VCD%.4IRNA&K@B0Y :U$(&C>"X>72WUC6
PMBM@%2R3J_F;\RC\?F>[^,UAY2C3?6X!H94W<TW2XD/O!X3LQ4-U8!>VOF.-M?\]
P]4\2MXA;J"$WY^PXUY+'4Y;V,3FO]2$*IR/OB(3\*R'*J,/R2Q-Y0#S9*3$'3K=2
P<8RU9B+!BR-QX21))1T<H!O\[1:D9W73BAJ+G&'VBX;30<]@FW'LRK:(85P0)29[
PBQ!&*6W&.6H(&1DM-T4#Z YA[(\6M\HK.ELZ,L_29W:<7^^,24BM>+H0 G!&_K:F
P+]Y_<R#B/(+J"^#J7'2,_=P"5;4(/7(KQ>!CFT1FT]#"Q1D%#.1N@8YHWE<+EKQ+
P6["CF G8*L>Q!+JM9CE[-XW-396(,/N<.J(NG#>#+Y:6=!2$/W!;<+B:;*#V5KD,
P$U@L@-5@V3%<E8$%&O,D!5/)$57#(C1?!VO"$V%86&SQ@XF6?S%'N:\VB93B\*==
PUR T99_,J%>FF(LUV\C[W^OGX6'5B42D[N(+:LO)"T&ITI?-3,)?AY#Y ^'[DK#F
P$<:OVAQF3S!V056N&X ; ;\_'3V_K!?O!H5R#\*%) &R%ZZUT;-+FM%<YR.P>1&N
PLXW,3">.T +/OSUY1;'2QDC9.;*L,F!C=*V\)_8:TTSI&"]*N$5G IW90&!F<"K.
PMMG"3X<<5/E)X,3B*S:_7[HR__VKRSMR,6.H*?Y/M.BFQ-V6338F]%^IY<\[J?7W
PH.W5J-)<D<+U ZP<Y-5ADS*5J:>F>(X"_+/RKF@BB?2-[ZRQ,FS5\O$/O#D+Y1/>
P00V>1XR\P1\F27V#3'I.K[.G$*W:LLF@??:4*B1ZE9]#C6/L^K-J6'X;AZ*])"21
PAD4.9"A*\;<(;ADB@'$6IB;Z/@F&ZD5+Y>OGX$[Z/8D:IDCYJT+_S54TUA?E]K$2
PQT>E:/"SEKW>U%,J)'M^X\1-7:4MI 9(3&UX6+)(B[B5%E=:\)3415'7O=RSMT5 
P<'\)KI(Y ?D-OH^3'(?66KM%/'AHR@$':077F7\@QE_N\O_\K0[1,V:,[G>2 1%1
P3,O+*0@2*ZS $9HZ,QO^6J?R1"B(HV?*-AL1$. 6=<8_4L:6<3<*91:(D!C0?MBV
PJ$&0WC[^S'F*A1'_ 'D(\$!>)%4AE(Z4IY=C!\6.[HGG)@Z:_%@$?>U2,-+"C]ZJ
PD8?]!GH2#+NP!K!)=<1F7$>9LV8--T"/0X7?Y_NRQ$6ONPI@[< ,))*QZJ1)7P;Y
P#BF*V V(IH+-Q-!(@/9.@O_C;*>( )*[_J[W6#;[%15E2PU@8#A!/?Z0Q6" _7TX
P6 <&)2X,\\BO<[B;\IQ%/XI4:2Q'WG['1BH0M5E/H3@7L5Z"S<9"2W*"=Z^JZ4_Y
P%6M^C%N3?J!93\L+ K?7?L=IRX'GZ):SNL;B?(M/$!7%4#&"=(A@\CY7C=GN.A<D
PX@MH@6]QC.,TCE.1%K%9\KD;!R'^"@0+Q[F$'W%FUY;SZP3^+$;^+GL&?,6UGF-2
PZO]2/H19X%W"F;2J$R\;(?&6^-_VF"%BO!GM 2Y/]0DJ1] C=.E,,[@'44B&$1 2
P",91FX)75D/@N..:&I\18Z=- 4E]A,Y1E>&+TV8?0>U?#',D*\3@!TO6UDTWAE7.
PQ!07_4F]D_?TZJD03@7?"B%?1OSKZ$,L0SE?/GVY!GVT;4<VII 92H4F4@UAA[@7
PBA^#8<JNJ9W#)Q!9+$I;=N) XO'/J_D!%B.!^TN(&&,& ,'<9*JS89_\@]?6VO]X
PKH1<"9\ 14X4"(J=$$@NVKK?EO[ @^K_E.HHVT9G:=TE5*/2:CC=V6@J$MV?*IG9
P([8#'IP2T-MS$</:^_VF+V09C936YG?*YGP+2*->QTHK\\80A^Y_M69))QUEC?X/
PMB(WW,!3$OU?\H[6JKQ&_H$8&]OQD+K2#'J,MF\Z#&][A_^Q!3BS?!T.V)(5D\5P
PX,1G(LU%KJ_I/X\HB+'%^/?4_!WS'==*:I<E4'2#Z]VGI=.X._-ET;*ET=V4?T=#
PD5ZDY8V:2ZT.-G07-ZB4$K02<>@DIO?U489>JK^)OJQ:IB0#P$)9L*'HJVM$D_/!
PH:[AHZJ8'U3.VW8R-(K/+-I0/7,B*]1W[@/[-A#9"CO7@;$S2;8P ;64]$_*>GC_
PA!E"1&,IG:SK+AB?RO!ZSPM;VJO6OZKC=<+4RXW?[^8*7M'C IE+9*N7K&5Y!>:+
PH,225]+HRV*JGJVQ?):*=>JM:$9&]'"D>_R<OZ'1;-7T8VPH1C>7GHPTCN2)%3?9
P.]5S82T2':7:I*+\H9B-N9T>I%BQ#L7E"IQM>*XD6YK;FCBU1[*>2\"<;'(VP_99
P[]^B=LY,5/A:0A<'P7$B#7K0/>-GD;EL2>EJG&&LUW/99*!0[?O;4DQ3<;.4:6;0
PGD"#L;P)0\<+,Z<'%86W<Q,*;]P<$6##G%Q[WR$"=+E"')!__0U#+)"!-CX!KA/]
PHQW["OFN,-*JW80-=^WZ>_J&:A*2W;TGP-I5J!%V2A(Y9H3-XOLA"V8R]][L=I0L
P.GNAMYI(^E<=6;[7"1?KWNQ=0WRL!U"5< \SOKSX%_Q@^?G8*$A/##O[QKQY*"OU
PV7>OKXW,*!=)\7&K<S_JWAYK ;[KS^,O9&ACJ/ZW@9:;2AG2_(SC!*A#I#1KBA8A
PJS)HQ$1#-/LE&K8.)*;.8D,L6&1'E*PKJ$XTAQG6\15K.PB<N&9_UXI7@UU9W2DQ
P^+,<LY:*R*B[1-NW+? :NU)&^I<9ONFWFMT\5)N8ZQ1,_SQ,M<(3#7"QXG"3_<MN
P)6714R%^K0+T'Z83F*)RZ>@F1E5TZF_(:7928L;&<-"N$@HRQGWFL@R!L-HR.G5)
PA=/L*D=>5(#*0#B^B1MF82[N0G5,F) \)*FX ;D$Q#"KH= ,EVK,<A8+Q_-"?I=5
PH.<@\$0E)KE*'[<$]JXH3AOU&GA&N)R1;#4]I!;-.N9%6^@3Y3/KSEN,]?,?%B]<
P R!?8\D#DYPOZ M2'2Q8ZO6 _=VN"S&?U@B3S\Q0K V=G,$O)< %D=_6HE?@>.Y(
P$)F<"*[&O0VH-1G@;Z_E\!H:+9^'3T05<QB<#'T\U^M#2]9B#\#\B)K8<$^]5J$J
P.;=!C%R]Z-_-/'BY6%9E@1JS-1@6FG3EI <AR!.NH)9A;1+C)==>P[_Q4)!G'Q0.
P[-UMD?TP&_E6'["D4-:[C.ELFW;?DZF[[YR$D(2$;+VE"W/B4.+Z?PKL+ J>)Z/D
PA"V^0W41$"7*IVP*WI>/;1)($W?)2F35R$IXDB:1OWS[''SS7-.V(.W]C&Q%7+8(
P68]#MAHF4!RVTVG"K\C-,T#Q=AIU@_F,_<DR_-N90&Z-S3CQ7=^5;?$$J#Y7:A8 
PR)>F^RX_XZ.YX0Z=9<A#QA@3G7= YI?0DTB$4I5T 3V*I]3W#I(@"91GDNW L[@A
P7X7&/K^3>L<BS"GC0:J"K@.PP<42/E8\^C1*GK4;,$E/HA3V<\$G^8U !OQ,5BCB
P/=OGH]&M=6H6+@FCM.@R-A9HG9!+ 78WN$2@<T#E5G/Y_>$P#G[-.?!5[.^#6$$-
P]IPIR<6*/(PO%GPW 3LCQX>I=]Q9Q7B4UOUJY+,6J&>WI;T9;4?R(QK"B@ ?8"#\
P+1FT,=QAC!^1-::P&P[L FRK$*-&UD>-70Z<JADMN5I$;F3357_WXFE4$6$X!"3'
P.]>9>-_T5**.G8[BEM%Y]E/AG",."[_<L:OJ0YRI"%%,3<40_R-@NC (2%5P$.";
PU9%<\5N6KI?@*C8G+K"E2-=,!GZ763PS0;%2^^32<&-*^O;2Q69/72X@M+M8E\YP
P [JH/>C*/ETT8"RW;[CY@H 9'F4"5=U?$<G'QM]N4\. 8L&&G]]%<6>!YR-R=T2R
P>UJ)DI=*L_\^QX%'S#\6ECPX^:.-QJ]?!?J!1/><"!!?Q7>Q;2STA.7'T$:)0(/E
PK7V'P:.9DPZ4:#HY,YVH6(OV)Q+!AHL\RI_T#72+(:3G)P VVI@%Z7L4YYZL[$G2
PLQQ;_"X[O1X,,T ,_8VI];)$6+:=UW W2M0*NO*4UCV=2GMZC&G^G>]0[5-5B<V=
P<%J5<G;H:QH3#NG=[8/VRKQH$^G"Q7G=&/,)KF;U8I^/Z9+[[-[G D@B1)E'&LU*
PDH6[N?LIN[",I'NW=<)DCEGH3N_18GMC91I6''<HYQ9Q_L'2 J((7TJ/1/FSN=BA
P1GM.=G@LE7+="#S?=>1K85KJ-TAJI;L9 SK ".L=DL2(D,68FW0\**8X9WS-5,$U
P7>H<\<U]Y]E9MD+P">&%[;E;?I@5B'DG9@V,(C*Y,-=:J M4$*;9L*V'>S#:,>"?
P]+"<L5LD716;_[4T9'J>-E(\=*# &4>V!4I=8$YP3_QHKDY@2CTR*"O'-;:XPKIW
P')JF%\*8$SC$R<)&)5+9P-MM'CNE 1&'149A)K,)N-+\36J\PJ;B7$V0R]BOK] 1
P$&3ZKCO9KZ3I2GN#E61$N7K+X(>>"P;3D95;KD:.S%'!QAI:J=N.CFG8W*Z_+SY?
P^-Y4H,AYOX+%_^25U"XWB";<<H1_'HL909@BQP*W'>@E8OM_<MS]G!M7#%G4NU#P
PB4[2A!G)8&X\['=/&L8ASA;O-[?4>[T*/O%VO9%RRB\WDO%:$INKWC$1WQ>)[$E6
PE(#,/3?WC80'DHO4).7P^+T)7<2[,V#X,U.1BB]#]"%AU-' 462Z<.U)#>SN$Y^V
PO(2=36M@EYOB6N832T%=? V.^.MU6R>O]BLA)L;NIQEH$LFY\ 4]W^.  <%%:6X=
P,IKT=AO11V*U791J!L+WA+0'*0'FE<,[WU]"H:,KGA^+92[Z^:L("AG&8^:4*1+*
PS6%@LA' 2G:;;V.UR6Q4MXQS6>ND6+)841;.GAU<QA%%(Y^0$',GMC0DPY/<I16J
P+TIGTKU/<A\: HSE3*!-*/@WL0?F5@%OK$@ [B@\4\#)INLK$#41."H>[ENJK,^<
P&=!AHJ5].A=+\@R/.T^D,0O(J\)0:LH6&>N9(559K6%#/3<4[$B+[2 2L&XLYL_W
P1WXHUZ#8[XG@$_=2$^.V6F'=)8=<UZ/;1[G94\(,XF%Z[+D4]U3\I/N5:/9-L#ZG
PH "]+4)\(]"\8,M,ZUT]$@>FH%Y86$BX#Y^_;&T?3615%LNBX&"539")2%(?U#\W
PE"K=?2S\U:3N>CAXUSV%@C7DL<!&4<0EIB';ZOT8*%H^ =?DO8(@1D=$90BD? DU
P8,<.2+J[0IMTV' 8_:]W0-FDP6^E(*B?5I%W+1SX2NSVEXOC!O?S6NS!(&0XU=VD
PM BV;S=A[]O.WQ* 297:-G4V*NG,7T?OEJIX,+;3GEHA/]DK/8X07E!V*>=0\'R%
P\2QYR^M'T=]/UB2$X.P,L@7=7_,D6OIWAX2(XFEDJ(3>8+A9' -@/'V7%':PB6]>
PC'OIPVTT"1BZBJID#,:-B6J3G?# $,\-!S*+FB]@*_Z0/O_"<C!L^H*2T/,+3J*'
P!8PB>%]P2/"=Z*&U&*KI=>,K_=I>'@,["80TG 50L -+FEA<)-3W/)=SR@A0P*LT
P(<(=?2(PVP5#CGTAP7,IRLAN!%/H)7Q H^-Y5TB!*>EL$JVUD((Q42J4VK[,%="'
PK#7B7[TT'A_+UI*09JAL:GQ'\*O2 RV#]L("I#NE8];K_O9'1P_-2KL'3)?-3FGX
P1>V9<+:X*R*CI0ZF\Y3-'#JP:E[>"#%X&+;DOPF&IZ.18343FS4JI6VPZ,?YF)RV
P.R:DF=1(%>7?LVWJL4)_%0?<6;V;1KB\=OY$!U:FM0WEO<_5HJ2V8T4(-T@M/ XA
PUY5G0W2&HV(#MF'%EWFF7Y*_=L0,NC0B20,S\E4YE0/ 8W*TRN(%$6/_=/'MZ0K[
PW&)VI%GH33"^]W+@EZ^XWS?%A2.FB[?H]<@'.0A'Y6J2]]N9E I$N1<[V@A,H,J+
PW[WLR_-?<B8G6+N?PEK1(M7G]J?(6$'T$#U:_2_L1]W:[%YB]>8DU GN5')[L;42
PI1+.7?]PB_<@?<_&.ZI0)F-H0I%T+>3K)C-4-!$TK2*FP'V,?EF9%GL1D"[]8?]Z
P*MI*MM1UX91?6G5EN8NK G=1?BNDJY?3H3K^,?^"0UK(;+7Z>>64"M/S.+496'*I
P@3(S+6E%Z5]3,TI%8/9QN1V"EJ0L>T$]4D>FD,^-)4=U2MJCS*Z/OR+ND.PJ2CFG
PZN0?@E:<30$VHD775Z87GNG1O'RL<_3@JEG:^\;-Z8F("^C]^T@RYA9T"76O#(.%
PQWF8$CV:S&Q&MT[UQ5"G7:RWGI1<82WCVO6O)TT&AMI@WZ&3WF1VGK6<A<MXV!F=
P_4.S<A46EDCLT]5:-*5$M6MOMA'JB1"6DZ;P3,=<$%PCTRP=%KFMW5X8/[NRI40D
PZAUP92!_U$5_O?9_&@%09KB)!\(3+@9\QU.[]&N]9#EA>>[@!_K-#H;3Q%](\^SW
P5<[3=0M>-V\DCL>^G&H,^</+VQ[RY_Q'5PM0;)DY;.OIWJXO+/.V+T8 OU7QY#ZE
P@"A I^3JCM6O8A(*PQ"HF;9UH[HEJEOE']Q!MUX.;$EIOSG^65O0 @AJ,<-*#KY1
P8GY/2@U^\&L12#/^@$=+KVDQN8!)2+._(!#!)71HBD:-.%?7QK,I9<]$Y-2X-\':
PW#]B2UC%G[]PO7'(PDQ;LM!5R;3:[*_1\^1HDZ,FAPX2XLC8W>L=54.]4AT^)B#>
P\54F>S'8()BGG[>XMT&)M^(]+;#4ZMW1BNO\B'-7,8_[8-+UDL&NE+3$8TJI )8G
P75YO3' L9:?G<,T5="HRN) 9CC2ABH793>1X.'F<MIYJ:'L2AK5G?EQ$P*YW(Z&V
P25'Y&U&K4VVP#\78F24XM&OWE"$>:R4@3ZD0_9B[>'P':'3W"E@"KYU=S#N22WSQ
P/ FENZQSH>!:QO[TF2/':!\AYM(KTA,2X!:>/=]_T-X=\N7:P.A8(QE5;74' ;/E
PO0VF<YB+>6SM_*-$@?7?T6N_UEGTA6-Z=:$6WJ3OWU:K9P,(3&#;$L,G)O0P"[>:
PNG8MB;-B %:C I%GL-E\J7P><<F1\-OVPMUL0;R9_>IH&JW8.,>D9NH7,5,S^+?W
PN_!B&!].JK#.'FDE/>KA\IAL/9^H(Z*/OFN3K[KEJ^S?TKVCPAB<))\Y"25;9WH[
PVU<9OPEV#!JM\,?AF,"2-G('D.HOUTJHB'$;F DI!DEUPF/#;.S20GKV)P)UX]Q"
P/ONR)R7C@"Q";Q\'1.S6[Z^U.HUJ3V1F1PU:9_#!5T(4#+[A&FI)23.J+@)A?7?-
PE1M).),$?K_')*Y#@W<?;,>V)Z,0U#L'JH#T%Z,[B44M7@P!#39T&GV>H8Y 7M51
P1$:HA:!?O*+"L2SH<;Q)3[D>/T XP4I/J7H]B?H'$-/ZNMW9[6\K5V,O\O-UH)9R
P3L1JF"H&LQ8.1VWD:R.@D+$@DHM!2P^^'',2\0BXH1G1J/_X1/',6P97:5)&P#T]
P>&D2<R@,VB5GK$\MCA*H#%%VXU3C.IB<@2R+G,=I3M1=$\3\LBV;$BX@)BN8&$TV
PL$=+%U)^SSSJ&^_8Z8**.+N_VFP12> (%$T.!@HL\^>UZ_1J.]-Q;]LBL73/7Z/D
P<Y(@7MUVF-[E,78U&*;2PQ0DKQYJRUOUBFHE>C"0'Y:HOE.Z(V0-B=,%=O5MT7]R
PA"4V8T%E8/TA5 45 2$U],<?:!<&0 _J+NJD%)E[AULQSFR]^&TXPX)*-GIS;_UK
PZZL^\VO@#%!-->3,7^0KQ J4YG#]J;.>^K?+)P%JE!KER%]*4?\?9P 1M/$B<4,N
P*G"W=')8H(^42UK6*NQLA ].!.@&8":]@AD3'  -EYN=P"2EJLJ)/75NY7 2X9XH
PU*/9-__%FH"1W931<Z\0:<?]_!*A0[JXQ1/RBE];@(ER5<+"!QDZ9?#,EB?W,J8V
P224^C!DM<DKT*&330XO?6L.)]<0@LNO)T&3U 1(Y%9:\R(EKMT,%M$B%>\8G>F(1
PI^Q8-0ME^?U-E@9PY%L^QC1],%M0\F[BBP5F>!JPUKYLX:.DPD4P/Z''FH$=FVOL
PZ9BULE.8P?-9+,]A>RU#EPZ[L)<"(FJUVJPN]0T]=GU"4+H9Y%M*"=9U.M;VR:;I
P7WXZG69_)!!F!BJ\L[]B?<%9,%"6?QT7(-,]Y)CKDF9#$V%Q;RH2M)*$] [$+3PZ
PZA.4'@R+K]6RG)V:*!PN%7,^)UL7C@E;J_6)1/'5U9]LJWX>+XC>%,Q":1-]:$S$
PH&D>SD&T<-L'VFFS5>O2*LMC<\A):Q2_/NJZS\!';SX4 7C=OA+.F"!4O.:ZXW>L
P/\FS5Z9T&<?>ST 7W2^FC4]Y(L%4F**.=_]6M5OV.3U<HO,NU&1BZ[ZX[_%MC!5$
PS6&S-U@N('ZS/3(:"PH.1I00$,L2\J[9++\/10M<OM?:W]%DEVIR$AS>%F1#+J%8
P]_BNDS?=2%:CVCL9R=( 6S#XVHYNCYGR;[)J:,Y?5N1.)>BB-/@'--"ISY5SEC I
P3*C('1O7N0)6#;;/J+<'HU*,F=7P<CA7;,)H];@\_@B?+#N&'8&HRS43^$*+@<Q9
P.GJ!JJ>4=AD=PN<QYY_G4^JH9>.\?LA"]=V?,$#3E?VU-T@]%L?V^?6."-_WI-"4
P30QZWVK #]):JU<C>PV1U@.8GQ<W FN4C^"T\U64["KFAR:C%>!:,SNL+AE"Y'JG
P)V@F5<@P2RK0T8F:-PM^ 3*Z)]$$+?17VED$6+&K!H Q6E4YWCP@!H#OR?LP: 5%
PLF],[W93<&>M4+H%N&!$R($<69*.T !"&W#R;79I66XMF'TS5TE<OV5?=P"@7$6E
P&:)4)#5)F]48!>?V+TQ=;"22FX))WW74\*P&;T!QA>/Z;XVDKDM%F?A(H'N2<:JX
P",89$"WC?E// _[3M@H.J.]9SZECGK+*SF3KV9&/1544MN(3: S/P8,VP_<O[=$\
PSP*UZH)0%#V9DJ@1,V];P6@B"< VXKJL[%\^[WZ"OPO%.4J0H,/J*:SZTXM;B_ F
PE2L&-0'--V#906NX=5%Z .E[K7F>;YCNDE6''QJRK+LGWX]Q/GA&ZP"]3*0_<()U
PC9<"RQW83[6/NGZ4\2I:'G^W/P"0(* JMS6ULGBJBJ*!GBWV+I+S&,/TN.,A_*%(
P4!G(";.K)HLE$4@. )""X.ZD.C,S"0ET0IL3:M<GJ3*3+N#K5WKNKP.W.CY;;L\B
P1R![@79QK@Q.D%GUL(IS3L0A'1^1908^]K;WZ;@_L^7&'8+N9*CSWV %@L),I0>'
PG6@J:UVU(KQH&]#L:%3VACDOX2KT3BV*<*(K^AIW3]!]4SC41(,&RQ>-<Y;"0F9U
PH^T9W$U[8&H BFCB=<C<H;]F)E<X5/$7-U<F7C=D6XFRL1[/8C@.(P^\0OT%-14Y
PS)P-X:Y>MMGY6\571N?@%+BC0T+9(G"AV,LZ2P"92#!BW+IS^3V>)G(/TL(9W+DJ
P_9Q,L,L:ZXF2DVNFYIT9 28>_5W[FP!M%![&P'GQNI10GK/*R8J,3"?[E]DZ4U;"
P +X*BN8LTR)G VCLB)V%)*0+7J VJWG:L '$4/*T]7?+<& ]_922;I72WD;A4L0M
PLV<:DUGSFJ-V0X8@_:7TX^]PQ_L&I>'EJ .]R&[?6+Q FR_^+\?Z+@?DG2FD.#X^
P0NZ7*>-C@W=R/*/TR1K'IR%<7:J/SU[-#YT\E"<;)Z>^W3US.O4(9+I=\=-F_BI#
PC"FR[:5F81 .P-.I&_%6/3,?>5X/,Y<H2KO6HR"\9OUDR*RPIL3EZ25YPC'$V%*(
P:M."@_."W*HOJ >'\]F[4+]EG.NMR!FIAU160*15#+Y +_O'T*9/@_@%IOX7S\9M
PHY#(Z0%+U0. ^$^$[):7\,([QL[$:T0H<ZFI_UM:RGW_)/\,K1<=.D7?1/!>HFD;
P*LJKG6OT"JA() !(YO9&5B2_L68>%=1%2SJ0PH6G>A^+:M?N[J_J@"@](F4@O?DM
PH>MJ&JNY,['UAIC'4WC>T9!6E,(='7>R&,@:=KMQJ4O* ;VBN2^>V>2(;T\$PN(6
P^\[%2-Q_8@@^1S5>7^\@OX"_ULW/^:)R$_\$TD&\NW7/WY1TX4?W344F2;+5:*?(
PY E':,[X%4*@M^OV0A)(Y/_<[AZ_D+/V//M%,(RB18'#6!N_?_(]$TDJ#":$]^MV
P,6'S1C5)VRUBCFQPT^#*V2($"KS[W->4BCGT':[=(BBQ4$)_HH+^6.QZ--XI9JEG
P66&"-H,YPY"N#*V+K6)1!OK;S6SNI(?0.*LSP"H/Z&=_HV#?V6"A7! ^\@#\-**1
PSF>L\X^?!2HG_4D_]/"@$>WVV\HD4LH$24G_J)Y07STKPB[=YYLM1T&$ #BM?HLM
P )8(3>7MFV[ 8E- ZTDMW,>!L:$_LVQ@TTZG\EIV_RNF]/_NIQGT9LZ:.[=C04=%
PUX*#S=M+R*+$NJ(2$Z&24\EGRFP<0'>B0\)F9U \J@5^ .F?^!6 U+=:;<U3"0\*
P?J)A04#Z*I(C*;;?R.BCQ(EV;\(IF'(<-_4O1E3A'[Q+A.VG+_0B!,+G:X-/%5M,
P"]Y/=I_9RLYL'9#S#C4H@A=J*3<5*G8,.XJ!>3=+VC,"!L=SR8(.?D;'OK[*ZF?S
PH%1:;U,57_>_SIFGDY(?_XCLGRN+:R2/<>LO75J=71U/;-T]YQ#OD2] !.<<"O%\
P8>TYB3$E8 <16>""BWO@PF:(=BAGN,.%4P@Q4B?5R(\E-&9SQDN?] =>):AXW8RC
PU*PS1#VJSM:Z6707'B)O:U8P/A'D80Q!$RK)V+,H:#(R4'7-*\_X&DU*77*S7#A5
PC)Y]\,?L4_]"(G_6!\,I8J5IT\:7SI8<9:?Y;CA593(26\@C[TRX;F^WZKS74_@)
PV&NMA 3OR_U$\9YZSZ'#VHNT *4I]Q:SFD@MGC7U1RO1)I/KI+)Y5=1G.#T64%#A
PXAU>,;CJRW'DB+N#9%943SZ!.U&R7.L"0)6D?40D"!/"(E"\H=XS<."]1@^07'Z6
P&I L2&:N0H)0\D67Q1+6-1I]4;6E+F5 _ L\*+L/E$5\\W018^WA7T^_FV+W._\6
PD+-FW?\KIK;:'LK_)P5B!I64QV<>30(]Z[>D0%Q@_>N&9H%&+GD);64*6:[T$OBF
PA@/1,@&+AP_,RE:V^B[C-M]_+3XWY5V^671)M3M'R0]RLJ__'.VE1VIHHJ3 "X/M
PB4D/90!&$W\8K\A<C!O?;0K#QH88/,53TFW' ]#XT)7WJ0F(K/!HT4SR@G$O$ZXH
P635-;MNLP<2T%P#8"!1:Z7M1@J;QIYX\;4QLK-R%O-PH7*P=2A%A9DN?\F---GY7
P>K)C)P-(,II9^<@WX8KV0\,P_;7 7@V[3@<N2-=.2/G,I2Y'WJ/X*=,FCD>+2\0Y
PBH4#<6;])>C9)-X\LSY69?UVSXD+:FCS+/FX4,SDB '(R@54BURN ZD(@*B+UDH$
P'$\./Y*G/_:2K9,[;$#[M!3VA@P;#UEA6P1%!RU,B(S_:=7.2Y/E#-CPT" )YK81
P@[@^Q_8.'K&$#O=JQEN;RN3 WI_3'G;KD&HK99KJ]VP%B$^U*G>@FVE*L(D]<L8=
P]-*R#;X&Y_.9^SW8(:X:'(1Q%>^'/V<0-&UPADW: 5$> <Y$ZD.E#A]".$VJB9&_
P)FZ>#>O2SBJ%M%ZXQC'@.Y^#<+8 H%QA@<27H;C\[7[>G)=E,KP5?T?1'X47)E.!
P.-;DV=&P[77L?2C2%NX,C'V(&^4>KBF0/BBI'LE RRM%Y]7R,?'*Z[\BAO:*QX L
P'O;H1]6.9K$)'! _HZ,H[H?/6AEU<)<R*(2F%H"T<QT:6-B^UI6.*<1B,1'SI#BF
PNSGW27\QBTAE->+C&Y<<ANYWO %@LGG\,Z2D$EFO^N1JWD$<XI>,:I:[N"&@7PK@
PE/R.!-8 .861M@ET#-/ZA!%C3&(Y0[9/[0UV"@2P=P\0W'@1AC8\A<?GP$/N<_HL
P0(A-S<3+8+L]ZU61.HU [?940\?)Y\QZHE8K*'E#X=UOBCUL 6UMA/PWYS+QG($?
P%IF6GCG!"Q#(E6E%R&*[D(>%3LR35]5A84A2$>U[6F<JDI>4IS(!H_WSFANITL8C
PFL=1C/<$"GJ,^P+],O8<$+KW9P\*4*R9WGK=*;4]^210CY4[LS'>K =__=3#5L,P
PI1W>+M)V8]JJF'R>PDX4!:>"A-KX,J(4)R6#A+?MTH^_R;7\XQ;V/ >-RCUNP)A"
PWY.LP#WJKF(DCBLQP.R?QV=LPYQ4QF./XN.D':"!!^37"6\=D 6:T0^=X^YL%F<H
P;*/BOJ_3W-98F94"40WJ)E8_G=:^09HE <ZGRM&(,ZPQP[IT^Z;X0__G\1E$2 P-
P2 6*T.P[8:&IH22\MUDM[8^:\1@A-BVCZO@ S(@";TY63YCIF<.KGC07(YX\V"H>
PMPJ/GZ0I?&LK7 JP4A/!99'+ JUOD"EXA5-".-7.<!!9=#5%R Y4MVX06*?^]+R2
P\X"TV)F :0WFAY*)8V+%_.]6Y'UN%:7LUS;4LW#XS+$JY?%)PMK/3(AIPNU-//16
PAQ(A%93=&HT@B[(L.3!.VX.F7*\T_6T:\2S4EO2?+<P]T>6NOTO@2%I^*7F;PZ)C
PL]_R1%_P@QU+]%24MBB7S<I%Q-/@G#;P?5=X2(KG@:,E;(LL+T <D@LC8R=^P@L6
PSR'OY^ VRX%LYRC5HN3[+?;4OKB>,<"H4.(3A90XFF7!"CG*\H%BIQ2-+#VF,UOT
P+^I=D/^4528F^XF;C^3!0K>JVFM*AY]8;^0 -WZ53! 76R/<#;X^]311&*:VL/NA
P<YF2<$/T,FS$6193; YVXK51O%,JG30H2^+O[D>$C$8"'+69C8"J\O'*>$98ZGGY
P2O>71-G:6:5AP.<LEM 8VJODV#2O5X7K5'.1IE3*%F 2 ':JNF%0*7D6_5-XP'0(
P)%A6EZH+N\#5 K#G_T? N!H3MGG>VC)]?JH.2<)'[D;U@!-J/C/W8 T+ D$D%86I
P1$8+G'-2!R0RX[7TKMSGF\U:Y0/$F!8!'HVV]^_#.V;8_YD!K<^+;.X*1C?\1U[#
PI=I6WFX2DS+X*;;PR5.NUM=O=[4Z53YF!%<(50D$-6J!$>N^MF)NSX-W+.6_*:ML
PSI"AM#3IFP/B>Q(#0S$7O2>#SS5=7A^-E"HY^-'#"O!I6'.NR04F2:@A^S+N?I )
PD#0I&WSY!XDH][+]2/L1/K2E:4E'H!I@&%8[)&.V!QKSZVE0/]P!#=S070YE##>I
PN<'810^5J59-SCT?5XMFEPMTRK6B32%'PLDXY-+57K@WE PI.KZ/"I-#Q+=L\T1,
PZ_.5P)MW6FS&.XAN@WQ@-IW-F]VY707L<$#4=2/?HQ[&'6[^>[AH>_GV.O$086%K
P+5>'QM&0K.9G;.HR-WZDN($5WW("F0DZ@8)!+AZ)5S2FXM+-X)K7L)L6WW=\<DB'
PB*Q%*GI8DM>_V1\O?-Z;7CD.8:FY)>?/X\V2)4PT))6S[.7N\@TR IC&75$CKD6:
PC;G;#E7 ^39Y?'K[XE+41*K25&4^:>!ZO5@>PS-)?U!QS[. R=!K>Y2.7U(ZN&M#
P:MJI,5PQY*TB2B^3_)0#QE'EFELZR4G\?#?[9"+5-'IM,E\^2R1,;KM521VX%2-#
PJ\"N1=4:R[XE)RB,4'OJMOHA%R3P:B:IVV/S]#0ZXR!LK"U^6@,N6G*D[IWL67(;
P3ACOZ"*SEF R>H\WFP0+8OKS(]H+.HY%<EB"497] 6* B,;+2I_!\8;>T7_O;:1/
P:8.L=CC+$#8704=0I^P1_Z76/EAYI=Z7M:?HT@+,/F1COVY)'@\2S#A7/=!CM3)F
PCL+&7=++]_*AZYT>:RAK(-PC]&Z KWC7+9IK9EC?V'!].T@+?8$G"_V,#.[UMC($
P##<6YA5OAUH$[;J:,I[G,#C<&Q0(CK/P]&0,O4JP0ULK9=.E,.R7"%X$I#Z5MWP7
P\T>\+8;7B' R]9$":AB:?0]>MWN;O_;+Y'0@4_'GP]RNSA4/H>^> U($+5GRZY8$
P0$;2*-4]]?!/'Z50%+R#1IEU&M02,D#HPHX$:J?=7_P5K0M==?! 5PSUC9W71^@!
P0<\]2ZL"HXROGO_0=;$KSEI8QU,,8^O ?6):[MNY/ (WT,K!;]VT'0[_B&;22X2$
P?8=TGP)S9) =*-41SY9NKWX,![<&4\MFCW*OS@%WN*@RQ5N,4*O,73OW9JG26<N]
PIRS)0GSG7=.BV(+OLYWDNMQHMBRK*5\\CV^TT1V>C ? )'\R??X^A//3ME5@_;:!
PP^SDO=1*&^>K=(IDK /].^947DXR#\O8,[/MHR&).J1XU.!&5NKI_DEXTT++")>1
P+D%U3^$4U'_V.B !Q4Q)9>AWMO)+.81Q37>+H/]-4PH^8OK]9P<T.+37ZYP/,2""
PAFY4H_:&)^9#?X:F$?>&WM*JE"M=(<QZ9:,^:U-T<I48^7G>+(%RH&+2%69V6S$9
PZ93' X!$7+'_@QD4E\DM7M1Y=:NK5I-CK%8=*:GL/77]0+SW_\F[ @0.VQ&4=70S
P:>"ID8U"-RO4=__+C.6(( A\\MV1Z_4K]*B4U7)L:NI.('HB+\7/A$57\ZO1-F$J
P653*H[B(5TU$LA'P+;(D4PG2KV M]%:9U>XCNC_J'9'\*C5N16!GW\\4M$^I9EK3
P?_JXZ>;SE*)9YA(A\+3'O2?*\$EW^08>XC6&#91IE^2$ULZ(WLGVT]+PJ*L^%(DB
P;L7<!H829EBJ49SS("K[J%+;.\%R*BZ:.FO=.$=YV04A[<6#]V)Q 7LV%M?UH QY
PQWQ57E[7@!=7F'K!0Q4OQ@[1 ,=ZWK2#G&HE>;HH%92X<_5L20H;;%?U@+F$'B@R
P$)1),<9LB16CS(/HG-(FS%'=84T)AL"6X )!O894F@]V_'VO&"N,/"(>OT;.-V]I
PZE*V=7T(/$[&B4:2V_3;8AE.'P3EXWDX'A>.6<H&Q%@^C9 =,LJ9;^I@HA?;>%60
P#EYH",> [7>>ZY#N9QZB??_SWS'>3SKJ90V!T\Q&V,^%/M^DF=L)4UZL'T^+5VTZ
P4;_K\U-9H8P\[^@I]FSRYHW-R0L785Y+1<$@&]$%FK&K*)L8ZDWLU*9I.2J&^]W3
PWK+Q@''\2W:J=R+$"9VGCJ2"O%G'@EJ[PJB?:U#&,,CI54Q)[UH\%TA>4(N<E+1A
PQC8S"7%)GFHH<VPK0![.;!&$DJCW]YJO=@OG@UGW))26TGH)M%]",>ZV-@T:6,TI
PX+],NL$QS8>.=D37D[I\5.ZI<*&,BC;22)0GQI2>V</D7*:B,=6:56#R420@%UTI
PXC=B.O2:.*^E$AC%7Y(!OO[K17,!:\;5(8-QJ.E<.+X0^71>;0F!*I='4_-F&[&)
PS6UK=P-Z2M!],?93\+(UN'"D9&\8=B,$>8T=7"/-T&H$6^,[,<=? 4/^SLOU[\U>
P<<Z/B)7YRX<^2IY7]Y>%+=  32@KSUJQF4)-DK^&5T$UTQQPCN7PX?$:=3CI10TD
PO@DQ.51#@@>NG+=5P +6;O07 *Z>!X-<A[C%1&K"CYF<3A>"HE.ER@?7X9$FZ>FL
PS;WPV-G7X=2.*KP:12+D6PR$XM[+^JDUTBE]X%GJ9JC^\46YEX#L+;J>$L L6GIX
PP4 XT3P!'VFW=*LNJF=W&@@@OQ=?JBW R&K(54T'/_/"/7)8V1AX9)C :PY ONQ>
P+>+"80R/+ET^U0Q^,KD6E*K*'QZC,Y^9[]_((0AK$H<MC# =*A<8I$F*0SNCGJ7]
P@/=;3!-:;ER;0-2)VGR2U1175C7<B1G%]R^FD1M/E!91H@H5C,9[F$1$QIG/E7[.
P_-VIU@RT_!:]$G-.W0G;&KS2\K<L\#8ZJ4_4XE@\9(?M/&EG[6#\#N:%<-5QUF7X
P^<B>H)J&C=IZ+<_-/'608\%\0>E%QN(H@PM&6)8E2&=!=5CMFQ 9\S\.4:6WZV^Y
P[")=V$E!D@V3%>RADGKUZMGB$RS%C)U4AEN;;B3@!XA*%0>5DZ%Y]B03M?-(O# /
P]C.(MGR IIPN#)]L,;"17G/_AFN0^RB=7?[^N5VE7K0%<+WF=M"!D]?18?967#=#
PQBO2<N-@'$%D/531A=9%_FH.4/LVU\'LWW*J'4'CB4^1:5FS[(/$Q>K5LR&^NPV/
P*'9#=@G))+[)H#F2[VOUE6E76(F+$A*E^AP7!0$^9VJ0,IP:E_3@%QAARG>P>K[V
P18WN7>D%)R'P6KS7#"X&(VRQD>!$>@B3<OTGK6V+AH+)RKC :5M!T3,QB2U]9F!5
P!-IL[@5]E\F(26O](ASC&)UUMUG%A9#4*5_!YY0^>O=KT<.T-M6ZY]1B,1&VY2^"
P2OKDV$2(==4UB!X1*G3&]ZLR<I;@RTFYY(+%'\B>>I67ET1Z1&&N9)$!;K9WV6X^
P+)A"H\\)D!^.5J2PTBTD,4N=I-H-/K!#8F&/+N@NX6V5'<U;*$Y C665>\;+2AG@
P@3;^7D<'51* B-D>4^E13:P=\KJ9/PBRUA0)-0280W.#@Z[ZL#OX>Q66P?OM$2+L
PE:B%,!-PH5$:D$E5JRE)B" 6U1VYG4.9NB1N^U 8">4S%E$L9?47$>WGZ6#S1W0_
P]?FFK!7G>V1"8D9+Y^-A_ZP9= QQ]U@Q<6K9T)>_^,KZ.2!D\8<_K6U:OF@F:00=
P+8>1'N=L2A<=2S:&C0R=A2FPU@_B(I@A(USO+ I(37)BP HMV# =]Y_QOD29ZT:O
P\_14V_2_"F^S7'GY<ES"4U6<\OF>+(0G]X^:_O-K* <62C+)JCS>O3V%LCO_=2#"
PI:X_$,0$!O-LUT(AL-W^6@1#H:$+==;+=,F0Z>C%&H"Y#?NY@C1P6,G,\8^0KA_*
PL2D#Q^]#A<$'H2A@U,39*Z#J71JKFWB2MSF@'*.9PCFH+LL>7KC!"8>G4'%(=E !
PC4YL_+XVGU:TJ[=&R/VGO,:KE#" 39 %I7$;74&E\M&N=-9X29NKED?^LP'I5!Y;
P5A^,K4^5]HT-SS?Z$5M2$?M/2DDXVX+V3C3Q2J4'HEE,9T(+C(Q^-A6I-J629KS=
PNE,3$F[W>!\%!,1EA&*>(U2"!.O6;^8A/CF<<L A;WU.%&J9D+KL<_\Z_=3]=J\4
PK8J*(P'JT,8TE'&?)>*^B[75 ".1@NK(JDQDN^+,,:YRR=1\_$L&!12B[.B[I?:<
P)$DR!9+3691S?B!)IC-Y6&P(-9;9L]:*W-V]QUU9]#SR!1Q+<<D,GXIVYKS0N)!7
PT1U:(X8S*8KBCM'='(56'RFRR[OM0]%%H985NVJ^TVUJ"OW]X9J7OQGW2Q!-9//4
PJ/41D?Z0VPCLD6$&15.ANBDFB  ^RO#= +PXO1],(J72KC!.&CV9(53C12"\\*#N
PSUN"=P^BZ)HX'2--#"URG-_U^# O:_-!"[VB@&I%VQY4G-SGQ7V1DU!<'-4Q5E_K
PE  / )WQ0]*X3!E^$"U%>S/:8(R1V.M++2"/_J*L$@Q<0_IVEAXGY+8X-,H8F7([
PVJIQ'7:KNB"HZ':^5@/+]A8CU-:YD:Q[$=,BN]!J_V58*((CHS(9(RCMSP*P6W.2
P,]_8+2,8)8'3GS&'(N EP-'P0%W/.X.KU#JVJJKT=>&NAE#=^7N]1(_:IT--6,D1
PZ@]8A$Y\:.-'"EUQ\T#"5[,ODF;*?3S[8_J=_B%Q& 4:3LPP!GD"+:@D!OP%J$EU
PX336Q8B+CLK;'UI;MAO^@M_?(=5ISSZC&//F]TA*Q4,MJ=S>_=[T;FNKX*_;G2%T
P[3@I_CON.W,FPN"/T^CT^K^$Z5JC;TXN8M'O*GK3TU3PCMOUG9D6E8M'H#D5LMJ9
PC8\T6!W5!OU4O*5AMT&JV1SC=]MF&RBHW3EVT*GZ"G>R.NA;G?'808;3;7%;%]1Q
P#54?\(1/I3!V[)-"MZ=VONH<$;!Z!PE=Q8^V^A>.[:/&!U-CCLG;>1A -:)%%#HE
P1=:XD)%G57B4,&TEP<P&O\_$PS&G: 'MJ-J:79JJ&[E%93I'O4T="O/A:C/:FA,S
PO+FHI.;+YU9.[:0LEVTSQ:QO9A1"1B<9M:P.H'<1Z59S.6&#;R/O+YPEV5LQ?[X\
P&(UYD;</KLW?3$U<,/\Y0:0X3TT<>".R@V7A00]T60_P29R$8M/19 ) 4->GY(4V
PSZG>W@O*:,G6Z0, =F([ "\A6W-_6+Z46!3=G-I!.B^2$,\T;?: 271[)^9I=PK[
PAN>%7L@7\'4AEU&4[FX3^597,31T^9"JA!+S=>_:V8Q=9$ROB5ZCGT3AO?^XIVHV
P;J49VA*(%?)O<H[NK"N[,%"5S,6S&D4! /Q]%T "\2^?:-$P*2P4!A428NI'-_#+
P%E6!'IT.?<@S=*$3H9@"%L$MST\X];TLW 2X?YMC2PZS\3]Y-_[8"U"431^,.:I+
P9_A<!XQN_?;+W!NX#P3-G*&3Y*];NVE;.?41[-EQ5W20Z..FR65_P)!)%JZ4#.UT
P4;):MMP]C&2#%D@@!T;W[8,%\A64O;11O<.0*P[$;A/<O[GB(]D,_HUH-$R^_*SU
P,HM9Z&1K1XXI%D6.;"#S]]&PDVL^MF]EL/ZLM$46WG#?6A3<AN%[6PDNY](L7+*:
P NLI.=-T9_"#&'0Y]L=-7@[8PG]'<Q ]$D\M+^WFBZ-R0,9I&JKIC(^&]B(!Z $L
PE.ZH"WT0 $(N+:TQ/@RS!>,SOA>^)%]Q!455US":9_W^;U3V6_G"Z6U:,OMXDC\,
P=9(5C!EU=JK5BJ*(+(:T##)&0''MP_(6LY@[(:03!:">,B3D<%S5.)+)H<Y2Q]4N
PY(4M?OM=>GV3Z_,E!#@%T9@^H:P\!B1'  %E>SX!&S4A\2 P?,WEEEA;M:A1"(2_
P,=^(M&=R7Z;'R(MFM"P*QNPB3I8V@?0**.M@843"7:&G!B*4,'L)1[9XNZ9DVTIA
P.$Q/Z#"$C4<IV2G*O4=ZPA@'B/!-ABEF=[T;DP:!\X-)CPJ,C-GSJ_G[ 524+"L=
P>JQ(I9/3*6?T1MHGV5"MHKCC'"5%^INJ&^D1CH$-"^LB-2FK@AOU@,+L7:3M.-!/
P9+"Y+MGQ1Z0ZX:Y?38+ ><@W"*E1K8A%4CF]B&[9/Z2_"&*PUDV<]GR:T;Z/4R[C
PNI=]D@)F.YP:Q@*WPVH))1YKLJAE$_8LW1#,9XWZ_4Q&R@O$"PRN1(KD:="EF""N
PF4Z#HFGP.$7Y EEC\B,"TA E!'LR!"^S]QK>^^"^<I#"2(J%EX8A>O C=I ]0G[(
P(7;_-+769@CBC9H@'?V*@84.F/"1HDA8C0,7[8?9;A?*^EDR>*^G4X1[3<3;C[GZ
PJAK2BR_#:%8)!M=WGQ51W+4R,=K.N-M4O7WX9L$P8@#3SO>T%QU*:__]ZC BLI14
P!5:>*W*D=#5D>EY7+7!"8;VEQXPR$#K,OI]_KX4K)3.0,E&G^M!HL8!X6\+SBSMS
P)R[H$" IQB6-+899@4A!1\,RF#L"]#/^XE?<NTC1>PDUE9Z)@2UU83[:1OB&ET:=
PW?P?@TQ]+(4U'D@7C2YE-ZX4[F_<6QV5W??-M/KP)3?0]T]*=PRX<PL;Q\-+&:ZY
P"ZJK\:Z]]X.OD\DB)MC0V^=E'V!)6'45U&>$$?P'&GOUV+2(S9H]I]O!$84M;B_*
P!88ND*L/=H=!&R\"&E0+QJU&$C])CTOI.?G]S\9$@/CJ.Q2D27)&G&C3- /+P!6O
PM"C18"9=G#EO?5'GELS4<<Y=$#"6U6.&#/%)FW1(<G[P4_59I@1\FTA<V':JMH,5
P8SP0K%;FVSBIIU;>_[G+[1UTOQKG_T8-#]DAH)$YB'&"6XZC.0/8!UK?IIQ8CP2:
PR,U.W)T1&WJCN 7#\]3Y]&4SE]!E6&M2&%X=H%4%Q&&FR"?T:T'1K@:C0'?%%-")
PK_RW5*9Q9=^JK\[VT4WVQC7#O[A&E.+NJ!DGME(/Q?1(!'\Z :9HA5$DEJ"> R?7
P12Y#WO4 %94"6R./VAB;3!;_'*-D8/_M3!,2[,R:#LIR.QZMR&IWX^0MZ;TF)]%_
PS(YR\OIA;%38H./7EL "GVR'.5M]P-NY# V$@/ *N8^9&_W+)?WC-8(!6!I;C"2R
P;B^@O[F>.(*B/G,8HV+#FYHQ8?8HW_6 AKYR1RYG14<3+NFC"YJ.S(]KR'=%$Z@X
P#]_K'"]7AV\6=Y?8GT0RT T]GNT\\]CRTBIJ/BL;16U8IL6 Z3H^^8^W:)N. U.[
P?+BF0C/FAIS6N:)'14RWCU XK$%@[L5TK$RK0^99+('$I/*6'X77$%1R+R\E[2U#
P"'E9/KG=5$7ESL$=GV"WXT[W$<$]]V<"[ER"4 O.7>&]>^EK+-'7^30@F.?MF3NF
P[A,+Q?OUO_:V>/EMU T<!_SL(3F:7D+HD4' AOYJ]S_4<3XG_M7JSJOG5'H3E- !
P\8L$RB8[Y?1-ZBL'E%P\[-^:X&%*%F8F)<V,V$A2GWW_>+NIU]_=55^>;OD,69]Q
PM?/(@7LMCMSV>I5?3^#">B0)#-<]"*/:'1'ID<A">Z/4@7!"T-JQ'-(>[TM.P)Z.
P]@N20NP:0X?VYQL',P\Q&W#UFA*)5[]U>RWY!17Z6NTMHT&JK4*-^V(Q$YL9$71Z
PD[GY\/]27YZ!9IOW;_=G$'WE2)/,0E^;-,9)#/&R^:BRT9&##U/C,Z03^D\7.=6C
PM3RHC(E3CO3A>S0[[#$+0,:>48Z9*F]42[U?Q;GGTI6MZ9<F9K)G@G@"BN:IY3I;
P$^"]\P_V?)F:N_D$FM3R" Z2)$A\7K&+Q/14D?QZK7>ABEL5/^2R;R$PN)9&,)L:
P5E),*>!S)_#]8R#9G'!^6AN65P]P<X5G:$K RG=,KXPE!G$V7FO804#:(]]L.DC<
PD:\84KZOZ&K.;D)DC*;7\M>)&E@VEKN1ZTW(RAC6L#,,6_IY7PR!D5II^>'V8_\N
P^"T"X/I"3TT$I=<6";_A^]3M0[YN7L)=09AAFB'@UX[CK"5+GM,Z,G\G W:\GU5'
PX&SY[W0<%\2$S:)]^71^>#3[@0BFA7Y4L*T* FK*')%8\H;\K(PL'D%4SA#A\<AU
PC]O;E3F^.]?%23,6W/7NX\+B1SRS719,(YVB\R+2N)6D9E+&=5B2PIYGC/J5ZG;8
P>P$N S6P8_]CL=.FBEB\B25QL ,-F5Y<C.D;'5+_%%^9]#M0LT@/Y'6N62M4]Z'\
P(^0YBCR"PHP/4L:?>A7R1!I2E%7&]5]^D"NBQOS2  3QHTLHDHM6TG> *O0V2W:K
P#2/[2Q'*D=>D" _-7Y\O,@C&BB]8]/ P&>.,6L8-$K'"T](+61[BU/I-T0HJRMN_
PZ>NZIG]>$^4.>.&$GTT0#-!()Q!X'>"8<O[0%#JEF'4G7WH_R3<F_C*JA(*IW]JA
P ZI< ( $05A,KLI&E;^M[*=8+(TD0S V/5 O,I<\=S0&OU5JQ#;*JD%G_]0S'G;'
P5071_<>UG/BJ?S=H]^SN-\0N3NGZ=)2S8SKO[-2GOMP.X?=?Q[].[8=>42Y7'ADP
P)_@<NRTGMH3(,6&6SU@2="YEY*I1^:8$":4XB^<E<@>RV??"&Z@,\3%0S[7@*.7>
P?H^+03\*Z'N59&&3ULI*#$;&WL1TGC#]=WW?T((OUJ[O2&M-^P.0"))JPA/Z;BNR
P4U=X7X<64NAQ'9L.N<ZOWJ^=>+7P$M,X)$F&6<WCRAGMJYWE*S_+3U5B"H*,KMNM
PAI))GX>VUVWJN/CHR71/'3\8<6,PT2WYK<D<8+(C4$8+-(PA_T&I:@G=)<#O[=>:
P2_@=)#F.%L:5=:%);N<GHB3:@5CQ>7Y(! AQK*> _CV5\%WXWJ4?D=4,#'8H,3R"
PB2QU#"=YZ01[C>6,RV.PTXQ'24! 4:GPQ:^4U'*;&AIV_4VG]6'S$=/(AW1A<2[$
P(#!,3WUY3JS-#\A0RW.W^#SP=F=$ JF;R"VEFM_'G""?Q/[C'-!DEWZIQ<ZZ5")@
P1S)5LMMT<Q H*XB';-]C=ZLZ=ULXV\EH3%(I+NM<$ZFF,3"%R;0 'MX-_RI/3<B.
P,%:T%]X>B0AM!?ZGK(<R(\Y)S5X-PO\7OJ A\(Q6CX7HL:V?(9B;3]9.>1]<;3#0
PDNS8C*H0F$(&L=F?@CM%U-2V1!6>9J^:S@YN)V.;5G/[P=+BWM!XO&_<W-\[;(B]
P@QT='F/B*:")1X[\ D=K+%5W\MC3_&%YWZC"WP@F.G*/IW(CMF;@/TY0DM 'RK;9
P9.2N!O8>GE5=9&7<;[6C1'*_7?&RH[">K!50PGK[J<0:D=IL,K6_U(:[5(P;CQ:!
P=']8&?1Y9:Z4-\Y3Q4M?,R6V#[/)_G2/%2=]KD4:(JMZ1<C3FK.PS2<>4Z,U@Z8_
P4"Y_>RRE&=NCXPN_6/4<K$R3,C: <J"_1A'! :6@G7+;MJR>8  /4(6]@BGU\9,L
PA=15U!XK<=[7>6;XA!&:W, '5<KV!4#+1&UZ1$9<LG<B?2=Z:;<5'K)3W!$AQO(+
PSYV]3LHH-%U1T$'[. "CSNP)L&Q:BA <\&+CK,)YT"FE]4E*DJ[VGV8 O/AEP)&9
P7:.V\Q0]3 $=DT? #%$6F,JUI6\RM!EKQ-=&[0O(C+JYM435)IRM6\*OIE>Y.9C-
P4%QRWD*T57IF5.4%<H+907IVMVD-M.+&BG=EU?-T.7J=-@*3#_03P]^_P[ )OV8'
P!^/.:(Q@HSA%=$D4.,Z2(4J.C(B!4_XS6:&X,<G@(&/I//_*6@Q@TKQK;IAIJZQ?
PDQ>!7J?"C]0[AM!"18>1>,<#V5C@4"J_&0O;"KYJ6O,#K1X> C.2$M=)]"=/?TT3
PAJ";_]L3U63$^#?^BAFV=%"7@(^.IZNWJ="-)RHXF5RE%A4$CZME7I(U0>6"-XH4
P4O[96_N3%H8X&#]"ZB2.Q<[YI9QNJ<)!E.O,;^4I:Q'X#J<S&DOP;PB$(AE04R=3
PE2OTE+Q^8B*T_AEA]N2A.E%/H9Z#F19P>Y5#Q HO'9E-K6&Q/"DY[%G';QKE!:,0
P[LSC]#W?[3WSEU2^9S'BHE84][;#K1G<6[NXU#C*0X8KH9 A4@0(J]=^;T"6HZO(
PW9,CZV!KML2<@NF"--#P)<!C^,![]NHB+;_')-,88\Q-W.IJX[%-,RCSI-&=) D;
P%&#^CM &V5OG6BYML06.:5'_5]%-GY&U2$MP41NH<XKV'AH&C=_?LN(A4@*9D>SC
PS;?II&IMP)W+!SHQD6=:(=#Z2XQD$Y"U! *#>$AO9*@;+[^!(FKC[KP^9E_(98AH
P\%S2P4"A^!;15UCJ O?Y"_U]_^/CVX%&T .,QC8Y%!*?71@>&5"M+X7M\Y>UE"S<
PO:N+/I^1+9_3_Q8VSC=!![FO'HY8W(K;HY"W5R)^SWS6E("9>'Q0,:23C-MN$YL=
PPE^DL1+WRS#17.AF +3S8-1K]I^]JT.AR0@1N'N8)6=P+>5P''"ERIR\?&NJ!F2_
P]+_N8XH@6MP% .*9#"GR<#+=L@EG(7MO>D=/S$0+LKK;'O8[RX8Z/"MA_].>K^JB
P6NHSL-H' ER.\Q.X,C)SEO%4.'/P,.9T0,[LR!F=Z_"M:)SMIU!0###_H/]]# D=
P([C$I"B6#GADN*YN"#J>>QVK$U(8MX5N>*:D'VU\(T1/7;0Q34B>%'[P>E0:L$K2
P*%7H07J$,,O46=5$&Z@[N,)WBM-RC62!7^\D(;.Z@'IPFZM(_(N=L%'Y$@J+I6V&
PBK-CLT3YIQ,FVZCQEL*IC0@6]^F@Z:K2PP#WTTB0=Q\,\ZL>UC=@"4Y ;/WW%L"G
P>V0-4CZ89AV;0*$-%F3*+XBS  6O)X][WRCU8%+SP MXPKD&/HQ@W:@J6EO-(3[[
PMW^REA*_*3/XEY8;*?I38382-,,VJD>,?Q7==D6>DT<\ORKM17+=IV[2$7,\MQN3
P7D##L:-5<'[>"PMW^,V#9O%^4 83V6R:^(5D:>,44UH=6Q >V]2,J$9)B=5T1>JI
P:L[RCMCK0F%-^>P_T6< _0_/)2<:^ U#]WB6IL;J*@D^Y/MRRB@>F#K4,W;Q*;C&
P7+*?D -I[_(FW0_%,R4:>F (/=NBXR70?;D=^UO#8??FZZE9?HFB"K :,:"SA-]_
PG5S74<-3S. J,@[TQEG/^[<]XF*>G7#3B4G_EA"E-\]F[<8?4&>!?-PP.5UAC2D;
P<OYM6=3CP1=J9;[$C>-ZE$*?,.GT6F[Y$4*BLG[?J1FM[TRWT;S&D>]>>,S/B:G&
P]4*K;0;\;VX UZ_$2T/2-#T,O0F\&>M5P7J6'$Q%6T4[P3(0G.DV4#+(0$4DI7/F
P)$]6M'+@[;F?MY4C.3E4,5'F@SBQ&[],NS&. ;B^V,M@;&1XF65L@UX"%5SYP%L;
P_5WX:LHAV1B4[H;^QY^M]*GB,D".7WGJ$S/[$-G'V$^SWD";IQ0<B0)MYEX+4+4Z
PX996PX+<%@$B"VFB,H&\?'>Z/V8KX6];F3A#D&$RAUZAVV[2.HC9 9PU0E%IRZ6-
PQ!YX:*!"86HB9.<+@X:)#?A(?F)>IH5@I7 LNL DC7  432,IF/Y+WPU:+3CG^S8
P=$&;(M)7*NU9\I[_[H#E%A)9@2RQY-[*I4R,[GD;G1"6I@BXM3NHMEL8 N%?X+^I
P!59-TZU)N75^F^@XV:'P9[&957P6JV3X4><SLSO>PB@H63A=VTP3WEGF]X-%UC:-
PI$ .60GS#DCD#U$#^[B>FG7/ME"5UU>9\8#C?JWXSZ".#^>\*.2PX9.GGA3'B@HS
P+Z7SV$JEU8.8+EW.QQQ- 59RFV(FOI]D[5U?YB)H8.N3L>3Y*6'&&R.4L7K14<0;
P''07;+H[LCFA<?JD8K_%7KO1KL/A>-^D*0EDY]'-,'XPY%N+@=9*Q] TYO"/MII1
P,S+SU:+RM:Z<)8;DJ=0N>$=FI20/,,T'B)#^BBH=K">MRV'^H]HCF5-CO0<^)M+ 
P7Z@"0S*HQT]U#G3%Z32;;\@Q-*_/4Y2!,! +77MJKBF">7GAS<C:7)6*AO/P1D].
PZD&7FF7YB?:MM_C/F5+#0[3IE6>_>E81K(6Y.&*9'7'33D80&3&,G+05G[*L+;L"
PN@XXV40*<YA,;+]ZBY4ZVIL)_>O%/VVLE3JZ_#XUD(7^Z+4GX)=^&VY."=SK9/ S
P)S>61%UYPU&_J\\2&-$,U>W&X@YE*$LVJ$SLF1V>NAU[ZUUX1OU(<G^WBB_'"#/"
PVP@8/WX=,UH3QBZ)X/GRWJSJLLL2.Q3:+P1);:'E"F;<$*[;-N8/ZO9I,<6NMVY;
PRML/=@2_FC2CH*&?)SF$G7N7(,:?7$\?F1< WVI@X=2>!=_];-^<W"<>?5*GSQ@I
PS-/Y& ?RV@K< DO^Y@7O(Y+!+1A%15V1\L<0>48]+6U[NM9I26K'<!/"*1SUR^XH
P;8O&Y9!&0&U=@#+XXZY05FYKF %ZSM7IA$'T%Z[3I'KAKNU?/UCVU8ZT73U<O F=
P#/L%J<FZS? R''4?!1YW"^:D?IE1JZR/U^;9=+1D5=>!(^WSN* 11"H30]]AIV& 
PP>(--S>\$F[V%.D\^_^]I^'K2,G2+9\+N89UO4?HW$Z<G]0](8#8:?/ L2=B4\^(
P)..(UF-+,UFPR]D+>R80M198+!_W(P:.+U-L:W @&X-4,\S/"@X,R+=R4!/:(2(L
P^C'5E[YU!E%*TV2@3!:(4PUQ;$@<1]<Z1:!UT,)V].^=ULH_4,8S%)JR3KZUJWK+
P_./B)44SRQ&?9G]7B1^B_^W\"4*J>Y5$9J"--IR8R-#&K;FO'+B.\T1H%?S3M#&;
P=L<LU^QM<<;05$W=4+)^YHF+%<'5(!?'_N$DK3)@TDZ@"1D9[>,<#"L>J("CUZG1
P=K9XO*76]AB1[4(Y'M*3!N*JRX$G\LZ>A=T60Q6)DM8S4G ,ZI"7;(:NH/P<T]#I
P2"'I_P#^L/OY4J2H<+I1;#205&?1@=UO\=>(DE[8Z5^8V9<Y-.BG%VW)K,D;*D^T
P2'EPO/09*@3,"Y';PUYQ;:^='97NR0.;Y0N4 -J931 MN$8<U[NPQ@T5M )QTVG,
P=W<' Y9Z,5<]%B/'B6Z<HM()+[ UYO0T5.69NI1B5)[_Z5F?>*DH?@;,&>Z]D/[D
P'@29KC.U2VL$:8"N<-A)'T1J$'Q#NX'?VH"+4SZ@>H.?A^D2[1=V'((KH[I&*KZR
P5[>$V-#NZDM]E&:1YJL19NMMNH+.WF W#_^,N[CA8U!;R0E)-NVX"X_#5(3:H;WS
PYT 0E]$Z3*YCYN:5"_>2H<R&=:G'N=W?<OWIN6=+*Z*Q,8@(3'LP[^@S@[<DR;*5
P+DA?A!B<JCT6 M- +GKPFLZS7HL7OUYUG>F[2_K2X WC$V.M1#XVTDBBN=KZ%O5_
P7TGD7K.PRX.^DRQ@1#U:U,#4U86T*U#UG^/B.)!W^XEB<'+ )F$9$.*-Z&+_GVK*
P_?Z5$WP? %KQHX$(W4S$),;F2*?<RQY WKB8@[FP.XL I&05!4I59R8T["L8.$N\
P.4/6=*O@'SAE7NH<V**+Y>ZR^!'8V7TI@DSAR75W2&F&F^+Y]X0:2-=6CW%O^FS1
P0P8@'O3B("W]+0&)6[5_J9.M5(*%:[#;[S!,'''7A5@>N6S ROB,"<^R84:QU;D_
PQ4.VU$Q2I<J$((LY7=KT]AN)7N*$2A,N:$3M&E$Z[/@$^F&&PQLO$0-+*=U\@'"D
PW Q)MJ"J)234!W3JQ(69>$!:&]^J5N4R_?*@UNAAURK4H"IA<4^=+FY]2 PE[ >;
P(G:/I/WQ&A$1:?0CP8"M%I>FWLL'>CG'WBC%T=ZJK]Q'06@R(IN65[[%)QI7(LR:
PE35ZK2O\!^O?D/C)EL_6Z(-U"L*6E@2"8#,BWY\A'0T55  ;W=R_2M$$$!6D%%6V
PU  BPW?*/FMJ9!B7Y2& H%,^#P:56,(*(C((8.XE%$G^#-_P]@8VE__Z44A/*Q=-
P\_^RJ%PHV$<1;KIC];,DY>'Z6=W9XT. ?P[:_VEKF#H(A/+O-TH+CNIFW.9:2Y$'
PU^ ;%E5#*^<U*%%_A+Q@-V&5T)0%0WQ%J&#V&13[% A8*CS#BP[@#=YU_JA_Q._"
P5CFA;&<#SNB';>FABSB1*6=0B4KA7V, T.Z^>S<5.JLA62\M46;ZAV^B$GTJ@SK8
P?1OJ"%I 7VR,/P#5[:[-X_72;895+R\E9"8"LISON[M<VWT,)M#%/5-<^_ZA,K-?
P 'W+.].L5IGAB8\K6EOZ;>#4J)OV=?&_Z*+2B-Q]42CFB@11QHZ"CG,V*SE1A;-P
P92LO7?X=E[%I+;3\KPXS$;T)4[=\&]R21_4XD'K<@=&Q;9I<Q?J4;/$8CWE_O%W-
P6HB74C>V:K6?M\T[^A*& !J[&6&JM!(=J_03V!=?8MIZZ&U"3K3&-%]*;&M?H_@6
P!'B1<GEZ4-=T%2,Y&QAWL S8##A'8D2H6,  %AY\Y"L:?%YG7JII'NC>/#,(4_==
P2>OFT1YU8G?U;R4$$*8#6VV(>@G .VCW&.ZAOO^R9CQ:2PY3-;6LUQ-D89X6?I3B
PB6.%[=;^PX/8';G#PJ*9I?"6\UT:8KJ_N0K"E\L7K2(F 7;0:X5]I3HSJ6RRZT]N
PZ&"R2]_/@'5]0[ $484$CYK<,72P[6LFP'>["CM.1[(E=7[=R(@P2\]MRT7H:9<9
P.RR18+^W '_)WL#:2(*.Z#4,D7(.<2V'J';(7$(T7: *-V<NN]N,4IG+(C<-=HA=
P[DP%JW>&T&#'RH\\HMZ&Y-\./V;<)V$Q/>4W-(:Z29.C)6%(!CY2$WJF.=(-8]J0
P7M?NMWO^V.-IL8!C@V'4X\'&Q+QE,Q;S]/DMK;6J\_YA=; VPOT3MT$9I<(NY;0Q
PRO"FL_5<K?H8Y][&!DR0H/)'+!@EOV<TEF?SU(ZEL6+JDI[H,W7=5B2BIE;,^"O#
PA5GU:%U?#(Z11_.XY'\YI]F;_#S1F&\EK1=3?4P#'PY@W'A^!";JBCAS-0"YU0*[
P*&O2A &/YT'6I[LX-.*3:6L61$[M;/<7QZ:<$N>0JEJM.(MB]3_U(FFC A2RX\P 
P>SVRN2(8G/O$_VSOT.E*:I;3'LF0+I7"C*L..VCW0241,KI-QP#\$E?DCR4!KD3E
P69YQ_,%^(&*#TK&\LYZ&0P[PHPU>=8"@8D];M:)2N&Y1==1E=EPA*2"%;7_"9?!4
PZUHQ05%[G=^,3>_7_,(='[U^D;P88Q[*BZVII&#TIN/YC1[AAD]D90ZTP8\W=\IC
P,:)!E.^UL8C/N[YRY_L@Q:V6;C.1L%&C!TKD9V4D& H0S>C3M %X24NZ*Q8H*8+F
P@^KT0*247PP>'2H_5;_>!"'LS@B^V&A=]]2++T1>6Z-=:@F2I=I4)HIW19'_!@H)
PH.V2]*3ML_(0T>.=$=ASC&'1CC";,1J9ZF#X)KT]*)/K($(,!ZZHS"FSJC?EG^""
PN.18NX,5?K$F<:G8; D=;A1JXR?G B!-X;#%6)]>1GNT-N==YFTXN$%Y?II+Q[  
PJQ=:L<4-QP*KOH5WN/A()CK2GB,\JT[^,!&)@E#/FCX<6 1<,M\9:*_7OL_]>+!D
P._ZQ1$]M[/!ZBQWJ+>B 1GEDXR7;$JT6$,'A-5VS@*;#EWP-5R9</TE3B0^4I1@%
P\>2G2?N*\9RG!0O>5<6IRY[T:!FX#BQO=6%.*;1/RK(+U/?8 _0(3[BAAN()'[41
P? &-Z-7+N8 =IWFJ"5YZLF6O_< 1%\IU#38CVOI[^T?6]:Z;:2M>M!I::R/R)=18
PI&VH'L8M+O5OS#92S NG1"KII+2Q+Z;H5(!MF;P .>=/PB-$$\\ =TEB>PXVMBG7
P'B^N*(JW28 GN:^:HJ?!!L+=^N,H67HWA#HL[9H4O)SVB!Z)X*8LYV+M5'I"J(%M
P'-QU3Q!BNJQS"F&ELYXP@S*[CU#\>Z)_MG)8FHC7I4P\N+V/40OVZZT,;HV@#JUD
P^>'C<C$>=Q\2DN;Z1HS[G09&*K4MKJ#&V FQPXE<. YC(TOU'8[4_7G+Z0MH2%R)
P]8QIS&;;H**^MIGADK2EM?\S%1U'HM!:L ,CR'P>H:6[*_M8C3;YRO].D3UT2P63
PF8WL+JGX1IB&?G#)=U^V@AK]"XQGXE?TFK/8[!HEDL#?:B:J3^$TCE<-WH>;T:WA
P_'%5VY54N*S)+5\<;"V[E0GD=W=!1"[/V?:)G^_>";*O]K@YP)87G+RD9HR,Q9!-
PM7=69G5[>LQJ-"!B&1AF% ;Y<=HRU$!1CWO::K6#AK5:_;2A&_=WS!"X^PVZG'>T
P>1BQD2?I(<4*_]"&[T:6N#>H?DE3M"1/M@K+OFJKC-E;+!S";1:Y9QCP6P(!0T?5
P7QWY4H'B)6]S:EK9_](1_8WB\[3*4I"9>^_L=L_YOY[\[?DAP$2S)EA7"$ZZNJXF
P/I<)EH_%=XX]6;NHU#<S=GG4?4,.\Z3SO_KM9:U&T%:#1;#ZJBK 0!2TX[R/6\Q"
P'7'>+FG!&IWDV5CR@#)</>.&"!'S&<J+]NT\.36UO29)^P'=Y\N;:55\,Q8$S&;U
P-I46,,/50 J:HED-%G^HY@3J,@RR:1@750(*%$'R)MQ@4/].;4\I@IXC3+USWOA+
P?IX$1BKG'DY4#Y7WRQ#D0'=K,F?0L1M%N?)91BYE8>!*C'(H(?/DZ9FZ?!2W>M4?
PH'Y;>"#_+RJ_!&VR[OK]VPYGYWJ/%"S L(50GSUWV5:,W>!@^LE19IQ9E5]2;4>M
PS8PXB4+(KY:*.G,)&Z9;J-ES!CE< 9R %G4$IKE4F7$Y'OX_6VX'9JYDV426ZJ)X
P!:4!3I@E^5)'BH#_:XIP2)(;U>T[:A^P_9XG65:R0;.;0F:T3>SUJ5JR<':I#Y>0
PJ>)A;\NV^H*'I"*R9@ WF>9_!B$'=Y)&9^327B!;)$1!V1=.!.\@F 4]7*ETWEQ5
PHC;7X"I #C95_Z.<@;8==\MC>A(7LL#6&%^C9B9&9]K^S-#Z=QP]DB]'P?5)EIA-
PYY035FB=]GT+T_,5*C'93P,M;?]]^+NZ3]/ZIN-=J C<E6L8$P3;LDZ8B"6FN!)I
PT0:7Y4NV)8GR,YD^*_I I+P/5Q'F2-.4AT@!E2N+.6U*"9O1F=_?T?<K([F_$U;8
P%G%P6K7JK6ZJ,.KP"IJN(^(4 :&6USJ][??V[8<)P[O$I9&V.:>JC.=2\V X)JYD
PO,,H86R0D>T_'%@1XW2G"%\L8Y(QI-Q5OTQJ:("7"U:SD=!X+$0B7YIVQ_X;_2*C
P*75@>%O$X^+L.>GDQ*3BIJYPQ?H9I&*A^B,6#DDH ":>$M-52)*%1T,!D$2@0N ;
PTM[87X.51[[+;/U![]J9\Y8 7FG]_@$57>WKD*1E\QN;D_']^%+</O"MG\9U8[N7
P3A!GF3*]HH2'%!1-MT<U!5V3PSWRK:9V[] FY9@:]G!/P3D./!=8/3D@?F)+964X
PS<3C,PL%-E(UY/6#H)9OL#>*H\M(E2UAXJ#J3T!0(=4.!Z!-B$$OH[J%S0T :BU5
PK6Y4P?<Q6[@9R1R:#Q^3#S%_:.=$;M0D2+R/-?8!OWCQ7V['W2'@$XQ0T-5@O[Z0
PJBN@%WR2=EZ) P:G6>*B;97.H,=\"HT)4VWN, %X%OR=C7L)8RM[S!FC4RN@WDMB
P$%"@3+FCFQL$!KB!-N8V_$;2HDWFFGE+IT:?YCP&ZLW8D02]GD&X4-:6\,$TDUY4
P7 ?(?!YMM[P6XJ2 ,D^U<3D5G+4TTH5Z56<!UB?W%'KJ&A[^D3EBK ^*"B:3!F#?
P!6$T'N_[(@E"HR5Z2&<O8RU!.8%(*E!W?WT-T.[]+M7 #>7$^)Z98T@ZU4#-QZ[A
P]+8V+@S5ZTWJ:\"KP2YZ](?X/-@%4Q244 \<,?,&O_5N$WU%*E3!7Q!M?K<04;]"
PYLV1OZI!&G(NRE_&S]NZJ> VV:(3KK3]W;C""R\&@\1:U52<& 1'JSGZX8A=@F*D
P-[-MV]>3%'3G&^DO/= *=IIP4=;A.LF7/A;;W*V%@9).)R$$,E[HZKO]UC ':8A;
P<'.U;S]>DN#;R"D0=<_5=YC[8%)TS3QT+_])7CQ+=*S2J7(E:GO7\!C(G39UJH_R
PXX\G+1"8B) %F>N=-=A_2;VJY=?QN*P(U-G,8ICOA+T\1-"B3S>C.VR!%Q*"$</U
PF1-Z-U56F K;02BQ8>KH#L>'R,_E3$GD-X&5 E##XI,*NL3QIFAL23^!Y%TKI, N
P[H&!%9S">5A%+R7&O%X;D_4R:WMA;7AHU V;[)G;8ZG#)?SC!^DXFN$<*--.H7Z^
P 6^W@>-N[_3?9)-7U0\[.^59W7?G-794C5OC>#"6&VHS<$:TNQ!R<21,ZDVXQ\3J
P!APV6AKXZQ7M!I3.E#H9[A]T8V0CC!/]&0L;9%I%^'G"R&@;;%NQZA@8%HK%:U4,
P/\A!4</-&6EELTJ5)N%I<C2S#;JYF\^!X<2DD+O-O9P4Z#@\H RLR>J$<^SM_J-&
P,OF99FYYR%B?2ZN<G2,$P]F01M@-RU;U)Z7GDZ]>#,OW3QQ0\'!*JCR.OXM6GW$H
P4Y/,5'W*5NRE*,E-/  CA)U?[,?C3@1(T7KPLKI_J&:0I/27B2/^R^]'" (J,X&B
PR>M<G6FWPH_'RG8AZ\ O2FVHP0/22S[QUB0I=FA'<MGZP1J=5+MM.(EX""N0 CSR
P/8<I2-FR;@WWZU3\[,P+*1)SAL^D3$==U5W4D["FOI$>R%D6_@.0)\;1;1H>P<1F
PHLNI2GM9LSDO&!9=BVR;_W#3!2D))UIMG?3XY+][+C*YI JK(H3LK>P7J2XHR59Z
P2>:OYZ^-=SUXZW^]]*>W'RVZLNDQIT:ZZD@UD;],HKH]=9O5'#,P+@SP/B/1H31[
P+6I_^]"%_I@NIK(U#5@W&&"$DJ_W^21IW4Q4@YU3F;F1KC64I"TYV[<,C8V"RD4R
P++./V5#?H".^;$AR ^P^D03RE!A'3A3%\>#L:CGBH"GIZ,T)Z#A)ZNCX"9UV&7N3
P4%BFNW[2:OB<5,D=:49E-,R_Y>CB*/R/F(G_K\,M<$TD+6LY5%8AZUL<.^VG5]VI
PBB//$(I ?<_IS=^SV2D=2IO]> +-95054QGJZ=LE$8:8!6E^-_W4H7M*J$Q,,X:C
PM([#R0 P&I\*6\B%2QE#/V?^TS9[-M;$T#LD[-5%/#JN6SXC6[B7CH):AM;DD$K<
PEC)Z3\4PPQQ+8#9^+>,=;6.N3F)PGL!0,2J:Z-.IUDYK'71$F]YJHZJB(=.,0KVB
P@*C>R":R=C=#;96AH6$WQ3)@969YQ<%B(""+,IL(7%Y6RE8C"V/D':<B &-8YVR*
P:#'*8_; [*9:T"X8:'DT!'IL^'EL]#G[!N6OC&8'<TFJA'D$.22+?:NNP(X"[)[B
PQ3$IL6+7N*5.GSB_6C[_%5.[T-W+#$VW6ZZ"Z"/11JL&WS+$"'D?>]8-NH1U@FE:
PGD<K&R0G9C5D#KJUS4I+9$[Y!"/8%F/NL: #LZEQ84-$T0>*M:DI4J'9Z.38SFT(
P)Y+TF*$89-"_G%;&B&';,[&DAIZ#DJ>P:@23H(C(0&B1N]0\O"N636-!H_L05#ZM
PR=#/6NM,V12BRA(16Z+?]$[.Z+PN%7&UYPM=OC4;]#H^7KP_6GG& &OO',I+72WZ
P2Q15F6 ;/6.'QUB\@&#D\M<M2%P.?-!ZO&.$RJ:';@GLE%X.G!P1''1'*'=^3:9)
PI4@-$R%\:BZJ'ESLG#SP2;<S?"C:V9XBZ3!K+:^/B0*2C2JY<Q*2Q][@\Y]Q[N@/
P$#(I5O[-GD^S&Z*FSNFN07)I?X/C0W1U]S?F&U$.=E6_KAFMXMENGW-F;7#70TA=
P%]:%A*<-J*%V2W^HTG@JUDCA%!'FY__JT+^.M1L&WXNM\_^*4HI'U(3A$5B%Q5"[
PYY2S?P >9T-WLSL7RM:\J";M^(88KE:*:Q-+9$E V?W">,(NCKM<=W;Q5LMSW +^
POQA:OJ+7%.;NEG)>N0+1\I3T(\E) Z*2 WX;^VUW0R!K?L(H\FHT6(19^;X*]0E'
P%? 1B_MT2YAZ"7LUVOD:W[20&"QOTDO9]K9F&9F0U*U7FVTMN;8B3IS?R;=%(WD-
PS[$B[HO(!;0*@N+)8KUOY@;7;C/VRM3F)2W QI$[</:7SL2*H9Z*G,CK2'S !RIQ
P=P7LS0ROOH%7T1:?2PCI<'74PR.1P(:MNUN=V<T/I_((#T1/S\14W>P#>/ZB-P-P
P'U?576HM:)ID=YP 8J+"6\&FP.27C= *:&.?6$RVNY1M6!-2<E/K!($O>)&QI;.R
P;0>F^YF',VE$GSG;6:L\WBK$ <VZ25_$Q]SQ\>JX:UW!ZD"V?LH+86;JE]:=0.RC
P0G'S6Q<5/\Y"?,P*]?'LD%^';ZXP!&^Q?*.'9O,__&I!2VJ!+Z#11!/C@D4C*L<-
P5<&<*+SYD"2^ _\&7I,4=DC1Y_0QHK$NY2#/M2RM6Q[",QD?#S:<'.[._:%WR!QX
P>QS]^$7YODU&A*P: 41R2W"::M@9(L2DPZ3ZOIH>_PPE5%JE".USJ;94/5\??>R.
PL_,ZN&R+-7PH57;%K+-L$7!) ..=M!CP!,;_C)Z<KR$5TO1^FK%@[(%8OZWV,=)?
P'[;7:;&BKAB>O)?D+XCC/3/Z!^YKP3D<CSXC=3O6I1A"%J=%\74(^1T(F@(:EOLR
PN73Y>A#%U(!_P_CQ'K[[-ZP9=LPG4=U!/DB*';\6OYB=0)LK$/$[GP1H%XI?*ZJZ
PK/;B2FQWK/;7%M@3"Q#&6Y#-8/Q".J0W9U 05@D#%'I&48L9@JO%VZ:B&5 M6VWS
PJ6MNX:SYD.=J<IM_%9D2P.XO:X+Q+FSD:AC3)5,>6II>7:V'>OD*^2SQ]N/KVH+8
PZ9T&A5+ ;099"RAGHT5@JBR@;7)? 1>$+;EOA54!$8FK#M?81XC_L&F,M_"O(640
P5#=,\>P&:05P?,U2^^?/S'@M.4#%7&,6'!TW. GKD_>^E<)J5O2G&PX,M5D6W!GJ
P_1.'XFOJD,2C;6-HG38:*48Q\Q^&C@&_)?^)$S]?[I;:J7TZE7[%!),']WT@SZ-3
P>!']\,=IDXOGA&S];%.;R<4/0>Y9.&"I1+*;).@HZZ?KQH"]*O>#5,D5$><6.0:N
PR6B71_^4AXK(&]4C_]Q(+KHO+=3OOGHD.<OLJU:A]E4%*L<')5"@8&K8%&4\CMVO
P8=/$U&7\O)51AYJ49&["@.!"0Y/)V^83I9D>,ZO^'DSOD#BB?JQCZY5$)QOJ80FV
P?N=4I2!W>8@+A/A[L!VE;'<:7 U A*@H#O_K3\KK*BFY_?9'TQ>O95N! <EPJ!"4
P%\4QM67HCH2.8;*I3%).9OQ\EE. A[Y-8KSRQO(,^!L[L6^KQ=7-KK?'HBT2H[QR
PKQ"/:.GZV5+!^1_&8&_G9V7-C7-36M5ADU@T;^ZV,2N\OF0O-BWWJ/EL\0^/KAU_
PQCSR^_;&%"U4YGWH[;U2E&DF41"N162'M"24?4V5]9X\D&.RCJ'"03'94X)9I1^Z
P0W&3^-XX$1.^-P-8Z^F2*,+EYS<=$,2)$174ES4&O HH+HNS@,#8GK#XKU,X5G)N
P%[<],Z/NZ'SL$'E3GK!V1>21/@,ZXQN,;*A'1WAB/_@L72P<5/]&4S335Q"C.Y;H
P!7NL"SPF7M[CSIIR:+D2:&A;KY]XP W6I!1LR\VRRI_&#-[N49_E:'-_85D'K.<;
P^V#!(;N$OO26&F2)]]4B4Q!QX@PQ=$:/Y!!R<=QD ]HN#" 1>JZJR-\%@O61(6_4
PVQXH8J#I>/J(,O%.0DFY>'W&1B6F<V@B\=_A')'I(GU<YG<W52%UM<<=S$8 L:>'
P9U7#<J6\T'", <.;]H/S:(4!_4F+'=7!LJ]DNDMOBQ6P^_JR%W?W;8A04F&0CN+?
P*J#69]\'LU$IFE_J.K:[+4[O0",V<>S\VSF9361X#SWJ)EJ;UDO DK8-^:(2F!)&
P?=]9KM1/*@"GCJ>TLL"U/B6<_D*8*EYA&W.$>X+3*O0(R,5068GYT/(JQ'O'/8P.
P.C>EJP"M^^69;O(ZP&C6VNB+&-6X%5.&C0+WXK O=:RT[)#.>\I*5V!LT)G+JTF/
PW%M1W5.H,ISX_@2(\J1Y)=9YL)!(\D'%3*-LSBJ<2XL);9\YIA6VI 9Q$U0<_GSY
PV/SAEA^%097X/F^ .C!3#HD*\;!$@D5-.;U"-)Y!]BJ6Q><0H]YCP0<T="3E[4\P
P2M0F0LS&$E7!#_ W/B&4T@L16Z_5C)V<L[( J]'A)CK[=W0BN$QKA[R^4^5A2/&9
P-/8B"'3R/YXK%-XZ3U*C.>* _FVJQ22SO/C66.03GM T/2+>A\-?WTQPQWSI@H)1
P::C*\:_[@=[N@E2N%>[!/4DJ [?UO*F=OZY+JMEBL%.A)B2<UP %RMGK=_HC?%@R
P1DVV0D3;DD3=2MHR%CM$A6>OY[TK33IFOJ<P>0@^@;#/ODP>HH\>#I*@WT\4P5U@
PRVJKB:J9M^2 Q%!R<Y2_>!XE->_(R#F_,KPHRX=2R/Q&25IY[:*K?61F"/X32_QZ
P-G5_]JBWGBVSHN'S5,=Z1@#.7IS.4S!(2#*Q#34QJ^-R]&*WZ!'I#7<0+E1+GCO&
P5:&PP:G6!V3@%XZGO-I<0DO-((LOB>=:UXTR(OJ&A]644->:&XZ&;?6 $6SD:-GR
P@<]#N#").]])#^5M6(^ML)Q%2GL(.!0"XM"?T8-DB$73A1Z(>KV3W'W $XTG+A0@
P:XA:I.(^=5"@=G><A"?,1!^5=36+[N-<%$O#K+<ZE"G,C(9P%Z<+?P=BKSMZ8)Z+
PH*96T=T/+H>TG2<R1@MNV-[;YI1(C:$Z.E&Z5_>)J5J9F"PXY 3]RJ7;X14_*%4[
P1!7)5WSV$7@]6+#"_ TP73#E7*3.N*;B$FU_K+:S7+[[IR+4AI:7XA8T,[%UD#Q4
P8N?3:Q[D%R%I4I(@Z57GF!G_SWH46];N"YF=K&)OD0"97II ]:$VQD?OWN?,F*X%
P<V 6(K2&9,((@_U&USPD'&]!J$=V;L.RK .L\FZVM2MA;PR\< F+1BNX1<X!2S[$
P?C>23'5BH  V;I1GHA//:J56;!B2J=X9BZL6[CY/@Q17-O-"8'S%+A-J5GOU23\R
PL[7O7%2+)2-Z$B5^ZF!5<I-GI0!.V5F%[!M_W/UJAE,6S8)'+G7""FVF@0NE+ PA
PVW.U4D.WA"5DB,!^Q[%NZO,NFVH!:O!>1@Q>(WI!^]9PA_E:0;>":N?F3EVBL=4E
P;"*+Y1K$:E>4/NOA4R;' 4J6))X!)1A/I(Q>(9IQ#,_9X:.WH^Z>\X3IZ8]/A:B1
PDCY6,V%&D$XD/"H42M8=@+;6DB5T+BCU<6H;DD2A9]*F6U3I-'2M^O<;20.'"XO+
P^<R@E>M/J[Z1R!++N9"L8,U8OJ#F;<X)M259AJ'K,'I[E-3!A0H/!YG;7U\;_\=>
P2+I8RY YAQ.*-RJU+0UA>K.G"0NF[<_]&P1? 3N\H9!KK=M2EH%?$UVB][=OCPGE
P2Z4BS?^TLW3Z;B@J/+1NP2=IQW+%W!1V=>_3H ("4DFB4*G=FB?0R0/D;OVL/IIN
P0^_9N4<T(8%DZVLH)!/;I]$A03R-)+[.L]A*CA<-_Q33$4U_:%MRY>*\]GP?SEK>
PSRC_:2(C1D%I!$?)+W ![R M\O"156_7R$F"Y<6[PU^=<<S@K:\UOXMQ_JY48GX1
P#U>D,![?^O(X\\C.Z>C7<PC&--0"(9*4)C^^"9J$Y2.+R]Z5&ZJ4DRJ@ 419^Z^*
P?^A?,O(840)H\L$2@@B+PY>]?_NAO%0'U>Y3>LAG!X^C_%0#HYI8M%IW7T&!1YMK
P#&3/I<O.^^X#5@>"<[Q*L6&*QYW%O=)F-G4<TY^1V?PXT?I>W O/5QS]L #Z&0%I
P_8BO(K',P<MLE%ES%+ 4&Q2\J,BFJ:/<IK*7XP>4H2")\O0UQB_/Z:SJJJ2:,*YC
P-'YCNBCA.RBVL]WJ(P6QX$HD-KM@B,4P[39Y!GB[Q.:;NZ_'?6GR 91B"Z@=PE9&
P).<5*DEF/,R4>T;U.(V[9X(E0PL7P!I_,IA6=M>K -&WG*EYZ9P?#?VBKWTWX]!8
P2<:U'5]#<3-JED%\:]KA7]MZ&POD,&ZM9,$]&TLIR"\M>%J4R*L^0"%/*]$RNPTA
P:7ST]KF!.(#%.TX\97R2O;YJ=!]IJFC!U[AW]'=]0.0S&:4Z0D@H)BT*OG82?:8(
P[OW@FW6\5=FBXH3GH9NQWP;4G"[?EIA(HFE@3R.T')V\3JR8HBY[ <*3VY#_&IX<
P$18+T2"O;'ASB)>FTWZ$ J'7^R-<LPHGO-CF 2<BG'O[(^XE8B,M7NGJ"@FZ;5,^
PT(%%X@XI\)\2O%)(.U(EUM*,0NIOFLPVK'DVQ\E/*U^N7S"S.1?R4QLNW$\9X+DV
PJJ;:Y?^@60+U4AF]90;<-_H3H7*9JSO/O'(44?"T8-YS!@W)@U-(CF"ZO@1"3K0:
PJ^F&L8")[-Q\$;D^0FBLN:[>8+X9CDQ.(W,,<DU%:WT]JVYJL)U%I+[;??BO .)Y
PQG0,3),]UJ +W\GLV.B\J\?B*4XG=ST)1M3$L+);NRX3OW@'-N@+K9L9LHPYQ[#L
P R&[H=+.CTK7)-8"JEFN3WR2)6?$K2##QC;26@9PHNM<K>R>3 W&(!.BH.U7GG!X
PH/308]J@=+U05DMC3TBT]ZZ6MB>AP?($'9PVK#7[_CF8=D4.A[4)R^Y]280/_>5B
P+9'59D .NF9;#9=)NF';)NJ>2Y\?[9$?F)P@*,7^^%V&R4LL*_-,<3*4&TEUY^?$
PTZMF&_[@S?W@'DH(@))Y;-4+"6H?2M\W?U\O0+Z?R? N$F?GTZ#A>^S^.9"'3)J]
PZ_8]G@)LLRN+]]Z+)+K#F.>PI(N*V*#"!+WB V<<<'5_EXE?1<)=X-(,GP43,U:B
P+..6V%SRI]!37&S)\X=N'NV9V:S(JYFN[AX:B+!H-)5[J!TLC7(H3?JM:P'$D0WR
P19BX&BB/_*X3@B%:V(.])0"I0C%%4#BR].9_%]3MS!#[*K;\SD/G/4K/'HLBEDTA
P=&>_WD/LE?M\[Z8RK20EIM5O<K[Y='U2]$6"QQ_J_/J-:I1=5*W%-5BG&\WT8B9G
P50]W-!Z0PT<YQ5?)MZ<M6+9^!'"G#\T\]LG8!7HMD5*/F@9T"!L57M\-NY&+(TW2
PR&C1W1E]_;9,=T_F(O15O\#FYBM4)=Z%2Q5+FX Z2,M+\0739DM4))L2PL[?3H?2
PE*W"6XLFX4'$18C6V7T 8O.*'=E+2<T</WTJ&:26CHA[NAE__(Q\:O-7N!+CJ1XZ
PDLCM*!GK=N?K,H[X%V>J"-(N,O7%VEJV,D1$<UB#(/?%5]? >R9!I3GK6H4DJ/ZQ
PZ$'WK'%02@;(56/,5?'20,!=5^B;.*R\@5"?0I>#-=:1)@+ECI%&G/4[,KS\EOPM
PC7])V#,"/[&=RR,OWJX;R;DS6'2-VY9[J9O&-6IQXMV@Y"4> O*.\5-=_KS6JI"R
PD>><26QQ__ Q5#=]GI&+*.+]?(^-Z8^D";9]+7H4XE=C#SUBLN/-<8'J\A@W12R?
P+R4=Z=J_HP&D6<)=L]V@.4"$A#&3&>NC)B<0??WSJPR&$^(8"YZGZDF@9I QX_I,
PVCH5T,5K72Q].<;[IJ><#F\KC0FP_8)ROS7:3&TC2(#O_Y/S!J=4,OZ_<(&$$S#2
P#@:FW*$%V8\==AS[>2S$%);H[(]$ZGC)-4*I+*5,/S/F4GC=%C;H1/2$AZJ[.4',
PBNC[2>8,=X\25=;F^[RN\*N9,<=YUF'ML[[\XV3#Z"GTT>+[%-!7V_X//^#L9X+#
P!P_^*28<9 (_OM!F1C0"Y]3VGYK%D*;[Y*C&6=WZI'RK+)X@)L5+!H]H]1*SE?N8
P2DEVR2WPH^DD0 NS>*B>0WGZH$="S4AZI/ZMH][$'F(//+)=UGI"?Q=4*_7HTS5I
PD5PU@Z1/FU8PA=-EZICNCM*"5'\1/6M1+3]%^[Y%CQJ0N])(Z#^SS9HMGL64S!%[
PG;+^4*8%!GRYF53G,.&>]+:7S*K:(NAL0O&Z[4BQ[''Y5:^3C(P5(QO132#*L6[W
P"35B>;ZB^^DM2S&=3L@=H=I'HJ0Y\XCH?8BAY'1F4;$U?-2VCKN'IG_9;LP!T'.$
P3==%#3(=5P@=(M9!W[\((P#IT&N_-"?2M,+/F^0Y--R3^G<,&!Q=;SRP05C/+,QX
PSZ,%1(<O*TR/^V6R-9M%>SI&*!=[>.^7F>HF5OD1()5M2[-^7JC$&QBJHV R5QZ 
P3X[$NH0"8M-T/0'N$#W"@>6.7-9+^.]Z5(N*G4I]QQK#6U6^)]4+&27-2&..3L^H
PXT#X$%!(@!P./2K]:OPPY-[AK18-8&Y>+CLZ[GN[Y WP+GU&J]^B_5LR^+%3<QOO
P AY[:;="4@7WAJ7WOU(U%S=4^HPMZ^ZI,G\1H5F7<^_=7G(1B/HMG++RX'O-3F\9
PV-0_2,?7SM"$3M<B2&4A)_B^3IS)^E\-*N(.+"=D-DFQ;WRDI#+M;'MP$\!V#=Q(
PC?@5]G$W+P163'@'F0Z[)2&0_,D1,BQ*=L@$<A\;TE_P,X1^=R"D-R\$E=<XYI:?
P=ZVSI!5-:N6 HS8'OP!.C:@N6LJ5-HD#">\@TJ*!OPN"/;P1-CQYRIZHT\]I\!TQ
P;\':E2.M(5 K[.9WT7 HEXM>,8IPWS.0^L+%OJC%M6XD@12>4A@P2UE52N>\R\I,
PZ3K<K)B">@#SHK]JJ[>1AT#'=)!Y49>"2+P;WG<B\'JER13;N7_9_E_P=7M(-2X=
PNAAGX3 :Y7/5"%! 5?P)#5*TFTF%?!-SG#6&YTYP4Y^5:-'3>7;%S]Z7'6>_SY_;
P=_#PG0"2S+V09^:\!,>'AW2SSI=A\IT.%(O2+[99NQ7/;K7(M8[C[$3J-HCO$L7.
PY(0X/-^=OR=N^]44HZHI,X@>^:C*\M'\^<'L-]IGX(+5LI=RY(2&3["Z9G1=Q/@;
PT@FW%89'E!NCP>J1%4E2W\X@1+2DXSZQY I01AKOE\;I322!%?&:=[R$5DL4?5-G
PT\WEW+5U'%I,(,]49]1_&MV\9WQW,H<U<,:>[OZ:>!7+\*7XRTM6/S]>@A)B@A+ 
PK:8.\S510@&/F0,(6&@^BQN' 6;,9FI"=7EK&-\I-_! UMP-^P*S>CET&)4MZG?N
P#]IX9>2+D[TT>C<0L%U6==;:&5PJM]#M/.>V="(&]QT3*>VM'L5-T) YV1#4-T,]
PS1Q8'CL$2'-@Q4N:3$I<<>Z#B?&NHU98S\,\,VBCX^_U))3QYHTS1*?%[][NL.ON
P O9^^1G$6Z#,&%DU:AL]:&@E?_NL#^.7'^$*?R3N>DWF=Z45IM&OJR>3:]U(<7^>
PQML4UIL;@U0+W<$0N"J&:B*R?X"Y6=47L$ ENC5G_PX%T1=SK<1]BF]@?6],U',2
P8GP*889QFT4>!QTSFB:IF:W(T+IP&A#M49P_7\H-AV9D33+&B?Z["PB /&5KO1I)
PU[D"O9V:7Z!7^5?9]8]?(0B65/>7! ID_\/0@\=6%3BP=\]3RS]A-[#-+(V8Y<*?
P"((Y? 09UUEU]@7*^$*.^U#T<S:8'D1RQ#HQ[TEA=]('5D0",%*I(SIX!D%%JKCM
P[V1)0[H7Q%,BP?.#:=H8<<4A/-#S,-_)I=BCX%[_@](W.))]#M;;0!5C,M9W,:8-
PU%-<9:_R]&O:YFY%QV@V\$AR%!""/R=I*%3<ON=.Q?2:OO\'1Y3$&O"7V?LD7OMU
PVY$HZ@00G3'P6X =I0X+&6WA.:;1]K\TA8!2,:ZK6,>8DK(7,QG8JH$VY%[1 ^;/
PREVXOJVO60HQ7K.;,J>,+5>#:MV@G]4$GTK@,JW.G?CE/ -3F!1GPRJ T%?R+!5B
PQ@BB/TZ&AX.<,IJY:2,H).HV[FKZU9O9I("::\3;D5<CU\\'))JX82'30'WA%&1&
P?+G#@A<V=Y^54HD!L<8>4YBJ;RSV*LESM>Q^6O5LN8\:#E)8/MU8:%6&-[=3_:++
P4@Y^S++?8U?[I9!P/-:QM]4.U[%EGSGCJD+8<%A)]=F^CS<'+9TT0]P1QJ[==0.:
P%48K64F/A*?MU>[#)2_<AC7-+N#/B.ZI?6S" P/0P)(ZG6F1M0<]*[;;I0("LF'"
PE0)63JO4Q6$Y^&X&BWA)W$VT+;0CQNN2LD: F8L<@:>"#I1&$Z- =$7=KG*> K@7
P7\VK?^<#H030'*X\=<1 *!HJ -[=4PJ\_P3.,166T16%8R1 >'WD8<C\[$+?_,1^
P;.TJMQ"F*.L504RA0GI^<K^Y;\4O5VT\HU:/\!>XX]UH\[F6>L8])@*B:I>?Y#_]
P7CCA_-YU60@T\-R9 Y<FMSP3R9_.'*UVY993%XXRBCH.=9CS?+2P"N>S[\!%%PHA
P?$2EJ4<65Z0JF-1HMIU TG_]D> L\!BU/#EC00#5R9AZZ3.( CI?R%\1E A>LN 3
P4.W>TVFRC E,]H3%:JA1IW 6],CO20[58*5PV/D9W>T%#:LH9#\2(GDDC2%!R@X!
P6E=W]E[E#PB ])'(\N%66ERT BYMS>SR;"LOKJ\1NE/"'U6\UD@>]XSTWJ.E^(2O
P*/+/%];83[&S[F>??-S:9,%O+QK=D6%( _+5P^RMOMB")D05.[/1XD)VO*_WB$QI
P:-OMM$ZXA<+?A+&"B^Q?S_]6F)$/%:\'RCVU)4)F9DXSNI=9@0*!VC2U_*(9-)!9
PNYV3A[BJ5PG?MQVW+'0/IZBKQ?I#ZMDQ9["&O#+\?%,!82OYO^&[W[;W)3->T._"
P<P5PA'GO0OV94)['AA4C#0BI6S5%&M7D.W!Q-K P-D<_!  NZ""D;3OY;!JAO0YQ
PI+OD+"43;&GC*?N!4;WM!$"5O;LF]J_>P,[0>]&>Y:IZU0AZW]=<%:0SE.^_,!^;
P%"_>@M!<YN_;3@!LI TD<?(&U54A[P/4YA=;V46YI1"/"'"TO#Q+Q&_E)>=;-)FF
PTW:QF#! H=I;EE$:G^2$1O44APY^)5"I?D-EM)-LD""XN:?7.6O0[: ]<Y(-_FS'
P&>C5M%.&-JG]$?-&F;<[#-DIN34/2G10G\+$ RT/M0UPEX[]AU+^I43!8=%=9"Y0
PEAW9*$?SC^%#!UE;YSZ%943X]C#$=TM,"C31'>%.2TET1R>AWDX!%U)\AVIPJN]5
P$J7B&5U#&\+4!4M#@=,[!YN+<@]V*"%!2 J>BHTT%>"]R/&/\S&]P&(+.*^&]8K5
PS8G-V,;?C+IM03N99W>2+FH$;]?IX83_V9B"X.$)/%/,B1J%K6.H.C^?$8&&)X+8
P%-9?J;/U-Z4(IWOXR.:O)+4X#[3#0_*26*P2_/Z 1;ACT98.WC\,$A:&%$.=FO"[
PVA&!Y%LUH]#16#A _Q..A9CXRP7J";,74=^Q%F-+<-7=(+"<L:?N:4)3#D>)YQ?-
PBDU:' 9.\LEOOF57O3LW<.6\$,Y>5L!YKTRDI9?ZII*6'IZ7L;4E]E<5PD2ML# =
PJ$H+EIE_6$1?P%VK>5/G913O[#:_IGZJ@N$@OYGNJA@8@;)&\D?PG\L<]"Y%(@,.
P0C[<-Q]MN 29V\H,'>:@E^!EA3F%/Z'JRD?":EC![8Y@NUVA*AZ;S@4J*.R>)3UQ
PP=SKE0;FYO!;<CGS0XQ!J"=E@ZPKELX <')F\HDMN?^YD1;(*'FN0D$=_(:J*K:K
P^05YRGG'7NLU"C+[P RZO]DPM9:#ISNJP-;[?QCD'"TQ7#^RJ\]VB5@R'N:6%N;'
P)7QF5<C[U[*B+NKA<&J0&S.:^<Z@OD3?37A4?31:-[_*U0'%5)&*)X,)<;O2_5P\
PK9-Y--OJN*_A;Z)Z*XN\ SY]!G%JR<@Z&!/-.N+\3UO/QT?Z+(3L=7Y;W7>E0)P2
P/;X)\WC\T22\3UC&]F-@%DO"'OY\[<@U4B'S@[MQ<,!4LBH4Y^#TI4W]S]N$'R.F
P)*:P^9O^8=,P K'O\ZT,'DY6T#[5<_5C<'QJ"0L)4,K5A_")X:C?M>:LAAN7U9V]
P7,.@O]JQ)>QI+>Y":_K]]\\CCGQ"ILEA/>V<L[UTIOAVF R72\]^-"&7AD>LRQ$9
P\VU0XWL$N>LORQI[<HEEQC9W\: MI)_T[G)1KKCPS*3 &[JSX>(_R:<RN*_'CKZD
P)IO\N7?N_R:>;^8+)O.LU;_#6L(1&(.$L\N7;2*A?W_<3?6C@&64<)6>/(Q:D1#V
P\%+8/-=<*YN_R9S$Z? [S2(P?89_73838_FVZI:^?77:# X\'Q#2GHXX6;'BV/P[
P/\*K$?[9EK'>OX8?I+D<;>B:V"D7G#F]G.O(*_\R?EG['W;VB08\K8, )@?1PT[[
P<WCOF/0WKXYS[2?EKZH3I$3FX7%G<L ."T"\;SB#0Z/9X+9SC6,<)UNB!0R-BSY-
PGG(-9P\=YF#5H#!RM#WS="Q1:D9P$#MA"!IB2S'M>L5DE]/SG\&X(JLR[8IU5J1D
P.IQ&08F=[H0Z/&WD'O'K-M9NRR9V#J@OQ9,$,X2E_4]9*8E[CHR*FY_[^LKL3M)"
PF?M-NC6AJ(^-!1N4A@WJD'W!8=0+T8#VX4=9YNPO7IM#N2;6P/!P\U5TRJAU* 96
P]S# G#*>)+;\,5*F<$.9@+Q43C'C^-0:!K8=[/AC)UJ?J_?S"<@Y\G]27^C$RA;P
PW:;!A])[,CVLOIWJ&;\\<%B*.33A_G@AV$<%2;%B##P+&'YM!WKUF]G.5+0/0R\?
PBFX%SM-]]><+4DFYCHG"K)1MP&15O\/B&JCJ99:3;I3HT[[TO8Q)O]A2(1DZ/:GS
P?+E)<G@L#=*;:&=1MRD<0X&N$MSR1#)_ZR08+"&A3>\)+4*&I[93%0;!O&ER3UWK
PZ.TH,HA.!'+\U0M7G+#EHS'!?B%KI__L@?FD*$S6F_3[>5_U+*5]_ 9G\;<*\'W[
P).5+_9+$\!ZRAV+FQ)(0*.8I'4=H,Z*M?@"TKU[;']>@[E@A-\'2#0/YE:-,5KWC
P M<O#2 9>/!D.Y\J/]%YS,@=L@\XV&T9YQD&NY76?D&XXP*GNNRO:6%7R.7=FYP6
P3?V<SEH0M6)H(#GC<?@5_+BXXI:WCH GH*0E#ACV8\P@+&"&T+'Q1S&O![@'T#@Q
PXY+?C,]2'.8F-:/7VW4O=*%F=0BE1RP_EY3<7+YRV0S!<FC8LQ*I#KUN"5N[8.*8
P5?>&@1=$L<4:*[3$(TRE8W)/!Z@ORB?&O<)A!V6BVC6?^V<%+R"T%N#2D"\;!Y7?
P/&,T?B/P8U"!%4X-WS)JR9V'X0# <3 ECSR4=\:S.4""452/^(/^PBE7QRQ^*Y4+
P5_)!^9GLD>V ]X!<1>$5^Z =.FGC(A)*COUMK(1AISNPS1AS[VJ0>W=-4=Z,S3'&
PT+J64>923>JZXVSI]$.^MFR4PU!V-VPXC,/' P?X0>*_^@M:SUA0\_%*?Q+)OC$/
P$N;@P].>QTWL%_)3+K0Y1%N2!P;];OKB[8"%1G!0%'8CB3CB^>HON"%Y@76.CZ/C
PV5$0*^1.ZHG%EUZ_Q--5D"CQ0P7K5,VNT#JBX?-O&G_ODGOGKU:M?8/[:RS*[2'N
PJ%PWD_"T :HQY*Q1@!7RTPF2=)QO-D6 1UPJ%+MP?H13J/_L!S.F+%.M'4$Y,,\^
P)%L"<62/8!GGG]."8AR'N$3$VE6]^ FG7"#=*,3V)3D:YP::ED![IW($D36O5"JK
PKP$SF>WLO6H/59X3)FZ'Y[XUS^-8:(:^[2:C$%R<A42<V3/AZ[Q_:RJAH/0BHJ[*
P# ' @:,)#/_B]M;E=(ZOV2^)2&!H)25A#"AM8CJPUACH\O+? JIC4T:*U!TTD],^
P2CNEIZ6D%H%,([5Y/)9RMRG7)T!C@AJ]V9S8VV&$OL)-T<XE*TLC]5O1@Q;?@9-0
P74V ;VIX2QY8\'>WF>E683+.!XH$(5H/'G]K]O?>4MNT"1*-%$9__HZLBAW]UEQA
PI 9.7W3D]= 2YBO+XO"P%!V4K"^%+Y15:93I_,Q/@PS!;=?6NHP*IA?9\@LO-O00
P+=/KC[]H5+B-SGL2A\'J2%!S]S=Y3:>LZ@]X/A:RNK)WX>85MJ]G8T*9.EB$/]YL
PYLG_@?8\LL+#2T-^_#8N, 'H&.6ZZQR]^Q%/BI-#T=1-57""!1=A1&COK.9C]]E3
P5/Y8($>"O)HS%+BG23<#.:V+[+UESH-"=MG,8[S)CDNTV)R$:=;L7/]U^(3J%?^D
P1"A^D?LHOKQ6%^+E&.H]%.G<;):SZ"^:?028-!6;3*K<WWAN[7_AIJ[*35).3'_!
PL_#O1C"SLS!ZE=3U>N*AT#IQC.F#25\KX1<[<I5:'S&2[R'[O9^JTQ7Y+0]_%2*Z
PP&8( ?F;L_DM$;C?!^4?+M&2!/$/, TN2@TN)(RJLYH1"R7"/%-)&'PK)!72Y]:9
P36F3-:>YD9XEJZ)U]D,4^T5PV%BD".1+-E(B#FP"NO;FO+G%<S/#'O-2=4?U+P"=
PI7,8-THT[7S6(9L$FVD(U;;$&%6M^;%W"?S2[;D@5)Q]TMK1F&C]UCU!A7EWX?<O
P27Z19,NQKE2JG%#=K_=!)\MN\TCKD+IF+<H6P6HO2+EMS3V(X^YQ#&AC%!2#N)3M
P+*B'XHF<75@=[VUL< -EN;HJ0Q/H$N5IIT%;*/6HZ\[2Z/K< @),)$6[-K!%&):]
PV[NH"7,/Y3V^%8^CIU]-[4&OO%C1&^[4!C+5L'V19 W17_N-0V1'Z.E.82K<,G-U
P[Q>RTTL$9#)&?"6VET)(=P5R-^Q6,=K9S(1C_CLF '8FSE:HA^6%+"2/TUA]GE>9
P8./"8XCW+T[KDI6$0+A)VK;T*9.30;KP0B2#]%51G;K14.PRLJ%35U;V428-WJE 
P<_.*$7+<WNU%VN_@IK.?VXD09'$*!]T@5!5WHT%2;R@&O8>2U5QE0KY A-7E5"TH
P*WR$/X(F9Z C!U1ABP.#;TYVWTC2^\E/6B]$GNN]G1D6OJ"LM+\0'XBIKGLO[1?I
P >TU3B.]8?1($&MMZJ/HC''U6:C:]":?B+;:I"569M*?$VMAW+2CE\9X^^:&4FO6
P6 U'$K6V?Z"+A:C!]"5EI**^!_EZ:K9I0_S!"8L0?8/014EG)3AR-,6FBZO9G5VA
P<J=LM-L($3.CQ,=8Q$<8"-D9)CN(:)/=:/("JAY,&/PV#SZU*>5-O<TZJ 4ZEL.E
PX>["Z'U/+W<HI?>=-2R6H/$4RT0'V2#6PI_M+KW")U['E[!QNJ?F[3;QD,\$P;X(
P.N<[@M0#\UD7]CPM$;3GU?E2]ZCE&<&3&YXV#>)AZH!FJOM1NRRT!.:5S/\++37N
PLB@8>W^16[[P@Z9B]7]-CLPU.M'TM+58PDZ<_]5V?USQK#;SQPR5LZQO/I^94<'M
P34W1\.]Z/]<=?YMZX[P#U2<6NQC3<3E*FF2^FR$@6%)0ZQ%];\YWH<RK17?E\\6]
P8/KT]W7"Q)WE(.L2!T>D/+1#K4)^_#KHP-S^-4I$7T68W-3D$/ZEHB!R=<X77P?G
P7?AI.19XOJC0;RUH0#[A]QHS5(^'PZ*$<-\:68 <09F9:>K*_/.D^>O&@9B76*WU
P%N&H*^C3DLBT.L,GLA43+,9[JL<9I7AC/N0Z[^=)N"6B4OUQLB2"T3!;6@K0YOK8
P&1B/Q<W$RS$IR65S=:$TA I^^1>R=0-ZWR@3V*3Z?*TZ6UKBR+ BE%%%:$:Q9VX%
PTG9+D;@DZ4(#=7-_*NEG"\.!^^A>V;JZP?)#2N7=I!@BD^$_Q@?SNI\I6^^H\7NQ
PM + 322Z=(/#>FC+[<,^7;CO^5&CQ(^",CX=+?H);&V;'L*NNAC&S!;6,W&-^FHA
PX",??E<\SJG=P+)N1]K,D[#K:\_G:1HG #E?L<Z'1Y*Y CPCZHXZ<;B!+CSDU&EB
P %1G,N8*4 8CLA'F4>U@A3X@#&F6DBPIRY9EA?>)NHR%U)T[37JMVMWF@ABC:RC]
P]*;8'F&HH3DQ3-L08!4CE!$&O<%Q["8?8..711]VD1F:'.)_0T#N%CR?/D#K!>;:
P ;W74'SH_ZVOP.V;WX!#&LLM4\,/I9R1-G2[FMD2=NT;\]DWQ[#8:;X#KVFW:2^X
P-;4KA$90KN%->,#TYLPRJCT]W#Y%IX#K E9&-A27=VJ_(QJ?G&4ZU8SQ'R,QRH/#
POOE#TS;@<4.B^T\$=DJR"'OAHZM!!<?*3.UZ.#6VS\_VJK=(T9FG$T@=A(%-&MD2
P>]G%7F^)1*0+EBQ2V\U]/5-.KTS+5E-1['4%(0\("-@BIRQ.KI$-@TKT<;)O2ZGG
PVFA+/V._B"0(3'Q^NZ_C[Y=DM2=LN3K[M1J3<\^;9F6GPP6M^S8,EP2:; .Q62,P
P971K1EE'DG_NBDT!]SO[_K2@!,B-VK-Q,82LF%P7++UQ $1?A]L1/P[WTU%I)BP)
PJ'11^3SD['XW"%$!< BE#-&CFRFD11YD,F?4"PNA,+1X!Z1W?V@H.3;KFB>??>R_
P*+FV\ >WL%FA;K0#H3KCS7QMZ@&,"T)_AUZM3BPQR'4P$O]PGE0+;%ZC6FCG7:JG
P.>KMS>BVP,W"/2)T,UM3-^,$>/3M[C4Q*W]CHMN4TN513]-U\L2RL53#(2W*BA#>
P>Y7L)5+&0L&'N_A 0)5DP;1J2,Q.SPE?4V7%]S0U]W=4-5QC32D#YZ&A2RP<TWYM
PI+1R/@K;SIG7<7&^C.W)"K0]ZJJV%JQ&$D!Q';/TG$T8"FX9BEP1)50Z.:(Y3>NU
P^2Y$-IDWA>6\5T^CN69%E&Z%+LZ/S9::&Z\@"TB-F%UZ!(B@ )(7Y]&4S)81EFFR
PKD'Q,<;_Y-[$_IAD#)K6&O* ;6GE-5P8HYBVJ^:YC#I?)+12+ULA?@EX%:2ZA.H-
P!>O*J/@F=:[GR#;=#L1@D_-1]T=**,7Y)I5Z&BG":^V-=[4-"8+;FC28N#\UL0,=
P^SE'"Q)<"&3I(ISJ%=YZM1N)I6H^WN)%U,VT6'CURV&6G@S^UEK9W1_MB0C_UG4<
PME/BI5KHH9@3]I9C%=Z"4]6MM.'6C!G'TZ7Q#+%]D59%$HU]"X%_(PF5SUKHOR#A
P *V?H LOF01V!]O'H!UGD $%*I7*3F]2 6T4.K1S*'0+%(RV:\#UW>XDY!!R<WQ(
PK,=N7"3XN/D-HV=[PD9'4&K::=@\<N0OM)&&</+Q*5:O=$4[W<]2>@HC5THGSN6P
P/QM+K#HV@U[V!*="0;B^-W:^CW3^2(-Z!"-E^B4AA=;N;\9OI^GM4A8<%PC4IQ\7
P2%E,HIW-*.YN:?IM)SV2]J'+6KX9#8<XW4OR-X6P?($O&!B2I=Z7+DQ2JL16//*8
PU#VM,BG*FR[E4K7$^FDH*:?S'>[) Z<_U4F99^'."$2YR:C.^9JDPU9)J2)$U77_
P0D,LGRE<<?6-#POX)'#F .]P5-HVO^$.49(CRKZMZPM8"Z&?%]"Y7\?H1LUX)'<+
PVU'[4)+>PG:(.L1^%$0.RG/ XS/(;-:;=U+<)1#8U!;L]DK2*1!!-_@<A:P'VRW&
P'SVE3)A3H!Q$H;Y'MB6 B!B!9 $ <%&BA_3!: Y-M?C$ZS?9:A*IB=.AW\"ZQK4(
P]NGR+^1>&%_:&*>SJ![+!\T7[Y7,OAO_#CZV;G1LPB-=E2LA_I/4'5%HI,9;\ZIW
P>CTT:!ED,NHH*B$X?9\2P')-XO*F5T"!YN'?/H:SM.YKF<(/6D\^V@$JS$0AGG$>
PH.\ @-3Z>=9MG'+U=?H&C;0I"<G%:7P5;QC=J=^8[[192R9V*X<QL4&8BJF%:;AV
P%N8^&%R=O8Z(C>JHU@7?YIO*LWE@P](.5JS,YPO ^LH.4SE2_[(;$X@/^W55CR%W
PN[-P\'O0<G&-W[HU):U0YZJO?$&86>80<G7<?4NZ[(*KM#O'J:()=Z!Z7Y3?Y(%=
PFX(9A$V$\KI_J_D2<?R/QL.L8'AN6AS1,.6U>I%\0YQM@#'^)#]-Q[MV>RY4-=L\
P:'V^O@_+TO]&JCE@I(/@SS<C2TOLCC\IT/!)-+G99C;T_S&$(IJEV\:."B=TI/TY
P/F@$Y.!E#>!;3GVZ8F@/P?_= 4RG_$S&F1'R1L5V4.:H+SR(7S03#A"EK)WR7(=O
P\W64+!D""91M:JP0E"%\AK*ORT.-LKLR]9D?MX!FIW.N0$,^\6RV I,I38 ;?V 7
PB2>83#:C;\Q%=+ZS3K$B!(10-())E:Z 3<I/DV9TH\X(#Q,PUQUF!.2U'QKAI'(^
P:NU'PMNIVE-NZ84>LE(+$LHNC6$ZM0K2>(GZF(8H/<>!7Y_'GNI9T?ZBJS4=*DXV
PHJ[W>2VYL<$XCY5?H=S=7W"MB4MW=N90VT-W"%%)D2H99D&H/TCE^HEQ:%K[!+UR
PJUWS <#AI^AM;--?(!WC&/FR+[_20,;7 +N15(\ =!4P8%'3&?2]M#VTB79!!&]/
PPKQ3TF<+\R74+U5E[Z&\I/IKVWZ?%W4"$@!;"1H0\T$H<G5G4<*WMJ5 2'5&C6N,
P[0Q:/@9PY"<\<5:ZWTY[V/M4 '2(C-$H,,\T%LX0>&HN#;)$D^ IC56O-^NJ_*KR
P7N0H_I\H+J5'G#X>\4R703+-/FL7N *':8KRM\;X5A] 4K$G[E6(JD8%%1L\6^ED
P]?'CC@^M;ILV)B#4S"]5A]/."I,8S<'0=Z)A1V!(O5 E:=U9'*()=&2#DI6>;A]!
POQ<MBI*8GTDU )1GI[O*UCXAD2(#NW865JM!8Z;YYP12($F[L:N%'?0785$.GG)Q
PC33H 8!I492V$M^+),9&\.H<P^3$YCP,I[G\?_7^8M2AH?/_Q H;! +LA_H$?.I7
P"ZC9,MF<=WOC**3.+%50.\+-\ Q'#R1! "?Y\OPC.>&N29'OCR*U8?\([BUDETMM
P6!,C%*042I<G&L?S<G0F<LZP]"<+;@4'/(&CIQC.:21':$_FVRU 5T&;3ZS=..'M
PI=^YJT="K[%]6\W8Z\Y'4W>L"7Q;:ZJV$1 NXE[ +\SG[%CP95 +C9).[;#BI.I!
P(/=DK"K,1^J7(Q@[AHAR(G?ZAJ-O6'?6(4X<-OFWM^C[,RW?2H'8;"FC&HELI7B5
P![U!%6OS0ZM0_&;B<VSF.7).8--MA!]V$UQ1Y9U]#P-^=/&]_7)BS?=?:Z!C/^_]
PT]P@V[8H&6UISI\G]VS[O!RF+[EL]A4CO3P1X&2>Q0E\0B),KZ5(\&3/4[JP6EZD
PT 1I^>,A\D^&3CY$_OESJ(#+>BO,@"I<[2>^/$A.OG*Z?MG4_KD]\$;,SK8I'+&%
PD098A_J84[UXD\>!N6E#P *VZB_J]#51L7_,"H7XJAE&S1KY4.4(22G1M1!7+ER 
P'=)D7K%+[2,OBWQ0P5KIW8@ +%5GGND?D,?;=&2.JNIHHCH8&_M<[S/# _G:O_-[
P%_>OW];(D]P 3GV2$AMT,K'J6K3'2A/XJYI/C GO^6G0I_BZ+&F5+,P067=30#V 
P37B/I2N>P;.3;'[K\+2>U;M?/-#E^!JR Q"1-).XZ;U>"%[4;>0-3R@ '9K9^0AN
P1!R,/B_SR$30>,:H:=T6V:Y%J9_@.H X:AQ=@_Q.(XT4RE+\Z;XB;I"5M/MP%*-_
PY<?[\PO) A+#^2(WUD>D2BJ.CL&<UN _(DF0#9(]S>PQQ7<:OBB;%LG+(TG8[M5=
P/6%&E&EIE&_<D>73 ;G5-@H[0NK_P(X#XXKAR7?PG0+7A M#YX^V7953V>Y;D^MS
P[M&<?32?=EFE@MC>R&,C<&5\P3$?J?ZDT1V=TEP)/F#C!_K:CHQ\KIZC.4% _VVH
P=TA1>(U(?F6Q##I[^"D27Q*M)FI#Z$X=<)&Q@?^('C[[#M;IU??PL(3B1&PIP#.>
P)4-  ?M"C8&!2_&PR+U<BZ"RTCF=B^V+H?.H3EH!R]+A+:0OU?HF987!OLCFG6\_
PGPK_ W4]/'%6HUVWXD'$IL25;5^Z9N@T+'B18A6L-8L'&EPBJF18SX(,$JDVI]Y>
P0-085AYZ#T>Q!NM>\)\]HM''9HD*'>W,: )1**T$E#G/+YP,4.A,P^DF:Y:S:P/%
P[8(F29O4#A?&',,;;95-%KF-N(C(8^$D5K5A26E_:'4Z?";; 0:+\Z>GCYH+0?2/
P PCFJTQ.KEH9YJHUS!W-GR9^ [>I\;'(4FF?CPAT<YUP_VGMB/OH$W!7B&IPJGM9
P]N52[]N'LV8C[P$\*F3Q8#IKVWL-!M-8,KG!L!H76-3N/Z ?FZV*J3&'C#<[V@);
PO*6E8+C*BY3GS!(A)2H&CF9]C(MSR#&[Y7FXY^U/JK[#2:^?-_U%C4*:.663\!V 
PE_'%S.X?D!N,5Z6N-_'VAB-\6JM.-$V9^HI5V-@.R%)!\Y1[6[]V2X7[%[4^3-H1
P?/E^8V(!  ]8(BN+&^"+,M\&*&8B%%2M@ZZ9VDMIF\@KNVF-</;#OLCAJ*88J>1P
P\:59Q#EILMK]S3BV:LN+^JR*VSJ'?Q*>-T8 D1KL5''C0KIJ)#'3@7P6TIY5VZXJ
PMOYMN7ENB!.UJ63<]Z>4N5]MKD?O%,WZ!VO-^CZI,S:DE!2)_UX'LM6QK.V\8F'1
PSY[,Z9H=[MH34[Y\@NYBWDG$GK'%UZBYC-#A?T""&JVK?!<OMOL;CX=-CD2(F+^3
PS#L+60C1LY/![E83-BO?+]\REB73/XT\>4?9Y'KJA:LGW%@21=(7S(+<F28QA:^6
PX$C9OEZRA<EJ,LM2SD1.!'=H]359%?/- N2W9%WZ8S2I,=5%E3ZQV!2^5>L_W*2,
PL -D6S9#Q^>TX:C@F#3=2)M*15M/#"Z.#6'57[DN6.08!I!8@&(E94<,SC8/>I9_
PS,D($\J%U/T+X-P4].*18##%5)Y$2X?-QA./MLLSKV]7+@&4+<!QD<5>WN2/BZF(
PSF_#Y.:_WAU++"ZR:+>[H!O5SM871W2]Y'A=%5L:G:,!H+EYJ2C7(3G2GQS)\AZX
P]-8<T,.23R2!_49CWZ+*WXHC_</*"Z14*R<>-# JIN67$JX]&-*7-IQ< ]&F>I(4
P!JERF$3#WW!AT%W<V\ES[P)A(G)#A<9(&:X$(,)UCX.LR+D]=[M3?SJTGW 90&IY
P+%O WJ+W(X&,#S_\#-R_(;/"9P@6[]?)B42F@]E&Z1WCX87@C.UT4YU]5;XDCFVR
PIO[E'U,?HX/K50/6/$RX5XX<296T#^I^9!I!MCEMB/A_@C+B,1Q\/5S#@##BDK1\
PHS <YH2))L^^RIHA)E4&\/:?/B^6M_L;AZHEM(N-F?@/1W9'Z]/SG*UO0&,67[@V
P>(S9!19N4P\<&.0 P@;C,5>7L@F%^["N0MV3V[#NO_?L1O0@O1JI52(C4Z* U(F(
PZ=DX,PM.=$M@[FFD%=E*Z0)3X&&?!8%U)"K/RG)H,I+<V'_5!0<T2#%A=-,WS$I+
P7<RF064C?)B0_OB3I41NRH69Z<195?MFZ\L >N_=^$G+T*H;\YNRXWA5<4ZMY!9'
P7]?!Y.".+JCY\?? CELV ]:R8@"6@^(Y^WP<4 LZB]Z\G"=.P?B>TC>FOZ ;V)OM
P6=#?ZVK1M!.N7C; T\F26-X&[DU=Q4*[XG;$UYX"(IM:I[V;<P%"<7E?"[HTJ4<R
P:6!/"=3ZG\DCME/#+;UI]\,'%'=$*6%B;_5V\SAN9K5B]YJ?74'[NJ%B8.%V4$6J
P@)!V=+9D,]TAK?TJ<!W<+NWE4JK\']12AL7.<#*SM4['7)8-Z5A!03G[+\-29EB7
P8>B0\O^MH)+3BY>,EEJ[\R&%Q18UP,R&ORM[09^4C^[O \D\R[?</J!G*U%*0_(-
P6W O,RN<SQXA AV892 TJCPOS(<WAS-?<.GANFD,7\V.?XH@,SA$F*B).(AWV*UU
P1HE(@T[J$21L@32(O&K5\'E_,(1W&D0=C><3R:/IHR-6B;N&\Y3TS42YJ5JMS$3K
P@,R%+4!O],YI3,-^!VF1TM">X<XG*O[L]5?MM4;>HF2+BL:$JE_->[,AI.?N3=8Q
PXZ2VUC:]'7/5Y24>#DZJ9,+D.L,8<V27DB*[U.E_HD3C*EZQC1^QU<Y8RW7$@-G_
PB%AX.1,"\S%=<Z<<O%*1%&\9V3R)K5@PR1;5^R+)^KF) MD>^2S;_&=IZ=(.O? 5
P)!<^\+3&F[4<62*H8CK>^67IF8B&+:/(^&(D1!,R^,5\!&0L0!TFW!OKC3L&E* (
P]']O:HQ@O^L.D+%-8)@@F+!R3IU<"IJ0'RPQY[B"5QK,W8BXX9U>U[B21(']'YT_
POC4HBNX:3=ZG<1T=<D_WDAPH9UZ839@/HIUBD\A'W?B$F&=#>X6'S9UJKE!Q_E]M
P:@HJ%5^GU[SZD+RY&/O>C<XI]P2/F$$^B_@+41;-)ZMV,4[&T4\G V.T%EZN&%UP
P#Z^C@_E2"<)*<JQ4:^8L!#,HY(<HVKRW(IVJ7H[RX+\H@]S+1+T1Y /$F=39<V$E
P[,:3-Y<OI=[MN]X\$LN=Q3R/5+/##&!@BA.2K#GX>9)C 96\0,$1XDL\1U(#^2-%
PDC'D[P=$PGRMXK16-JIH'C-6&$?5G&*%O>B%W3G?P-)Z(E:'AE%@@_)]8E8\*L =
PJH%A<5_/%O2X UQ@4+N9#G, 470U= <0GY\?G'75L>;UTIJI,N_!Z<P*4UJL%++-
PO]ULYFL]:EI>P,E70O3D;-9R..R]?B\1)8YF5V5_V!S- =VEY_/QD8OT%;)ZD\@_
P'8 HO:0^A+>WP#\5Y2+JL57<26M!J[RN^?)3W\"DL=$F==K)L-U6DQS([V[WCTDX
PH"ZN+TZ11W^?:<CT4"/4_A:FVLC>_ !+GL-A3G0Q6-TJNKW]:[4BS4(?_MZ4HN9+
PU:#:1IVS@$\ ^HZK"6@<\E"7^GDC@,EP]!H%XR/\ LXL(2M;G0)GP7#7NE^Q/CB0
PO@X]D9C*^_>[CA/#2A(YN@<L!C6*[ZJW]?Z0+Z:I/2_TZT;3E^T(1]4'=(U0>& I
PE?&4PGP;,3$E3^U91KNN5CS)9A:%1]N(_]/J4&TB?RU#NZE&_]G?%>X TX/CZD=$
P*DG!? R;W1QRQ#UC3CH)QS!IU6PS'<-!E)X4/6ZFUOAQ I_AMNSQ%22N\S'&](1F
P 'M*RRGW\C=D)$.$Z<H7:W):H$29JT6YC(HSG"(;UXTZ$S#-41@!V7[EQ6_)B^:0
P)9.I M-^^=Q;-M[2ZILWK*Q7ZWDQD[!(^FDR:JG%L/V#;X>]49A<[YZCBECEQ&XJ
P@6MEXDHGT(JSHJ7T,BYB:)4A5AU&R$#3M1"2(K9I:GI&YQ8POEA^@4^A0*KZ8D3C
P,4IOO_6:YJYOG!AM(BM]FEL6]K%8 ?0W%9GTV@:Y;^J63YB'K(!-2>+P8Y,=,.Y3
P1WL=!W7WAKUE?R7<?I!.>FS22:Z8#0#B3._(S"A]+T,N$B1%S+FIXC@81$\7G@6U
P2I+0ME8E[/_DAU9$>0I%[7@>TMF.<-.\7&B)7FV=5'JZ4H6'TD]%=."L).+CTL?P
PV7YRM55#-DK\>KXMVS(R/== .Z10+7A71.+A;F-(&EAYTO@U;[)UQ-W%C;Z9KUH8
P894E,BS/ ,H/.X(V:1H!N^>7MTU>+>T12922Z&$(1SQS,\.W$KNZST #;&#2'_]0
P9KC"$-<:>0GDOT#(EG;N_ U?,?#:;=MH-3T;T6@KS==*7)!^[5M^=/L$4XK)/DX#
P9[U.]3H(L)^R$LK)8;LOR:[5'K;-=UK0K5L)B"K/H3[+,R!4U"Y*!(.5=/R'[@O4
P#,WX4H".R<O%A]R6'IBF3_]\1+S;>P=!&\U?2%ZB!^EL@[E*!-YSW\6>< 161Y7Z
P:?\6<]BO"$:6+-_>E<1VF1+C&A^A+^9+M%[H'0"C%V!4.4!<*L*)I=7*FLJZRYLY
P!+P(8NY]'PWR&I$(IXC7E;/TL_M.9:!]/AHFP$A%@,=4ARB^79#J*QI.!MH=?MK)
PT"U8NG>E*RA?[72'-++%^WJ5#/%Q0OF2KQ9.$,E]' ]'>VKD&SY4Q;]RL W' Y3>
P_PR;L.D@RI$YA3Q\%;03-,L&'X6"SCC=*Y6V3AHUSYQETP,U='H%T1+Z4#C3?@6&
P4)V-\&0@7;_]I0&@VB,H.\P]#G'N_9AW.C4-#DD27;8!<5=Q)F.>%=/BVL='9%0^
P8AH]/=RL4" +2\9D#XI-GGAV>3[:&%.!**#>H>B2@;F(%O@PD;SY??E 86IT8A^L
PKF73S>2"E_[IZP93KP$Z=N9H3-N'_CY;Z6)=86 Y_&E(!^E ^W32BH#-0AE&'_AZ
PQZ"%5J9_@TI=K,XU1RXG'BEM4PO)@M+(2*^;9-"9:RT,[G=<$$G)Z&8&<^]Y..,,
P$-DLPP(K[FX'FU4F[%OOS%,":A27[KMF'JL*W1ZHLTN%<P\3'8"&Q^3P9WG.*AG3
P+N:!7R?GXF:).!IX;\.*I0759@"R+ Q.^UBJ;25^;A0HSA UT#@;:]?>R8OF<?H$
PE QJX R.FR<,*$KR<)_)0M ?XM#/U\/_-,X1(X4318-5R&>.4)*$,-$FT.X(?# H
P#$_EYE5R+_MHH>,H 0J*4"D>Y.RH5BB "U#514][HVOV2,\%Z=_<AJA)]]-W?ASO
P:.38JOFC\9/VP1 SAV]\O$ @]S'+-D\G_S0 J KTI7VA*451!\Q'DV'E(+(5!A# 
P[#R:IL2)B?_\XN<5/92B/)-U 9)VJ6)[7^!&&VAO[7<S/:553;UZHO%J=41=G+H'
P=X-H.)#?APTO>H"1=-DN@-; 1A]<)G72?\7A#TE<V4('[2/N^07M(7LA^%+O-+4N
PVJ%Q<NYJU#0$XY+U2C_.25\!#M%*:K33_4UVV^R&0AO?.F73Y>)M?\RR)*@FX1'0
PIH1;S<_0A@G0#VUP?IL[0L)0U93Z@JU04):TPK7M CT/CFC7YH(]]J%-M4(Q\E@Z
P)P1DK*>B=CR$.HA7Q4K?%-8H?58X?J9S2*9M_Q(Q&FQS3WXWSQ7?;E?:Y'8V+)QB
P?K"/_HJR(?=(FR&R] 0<DRGC*,1_#$+#G6L;1_MF2EMQ6,W,AP(2<0[!U\/M)#)!
PX85V,S9UFFET:CUYTE@IG"(:I,9VWU(BQ]GI^#WZ_$DLZV[F[@$/0EE_/V,F"'4L
P+ CWHJ<F'CD=\8F 74 BQ$V<=TCSI&++#[^^)S@C3X560[&A;:PO-K.?VEVV2V3H
PF>G<TXH^C[6(8J=P1=L;*?&><"4_V WB91:6K"O."05<L[32<*EBY[U)/5>>5V"'
P0%30XZU>O/1+VZP'6V$V JZY81WY<AJ2K1;#M2K>2!J.R%7 M>NCD.A61,+S2J:M
P2+"<Y&I#]3AI:_4D?D'B/3/^1IVW^:06OZI!^Q;$=]9_=#HT]6%[D]TB=?HWDP(V
PZ+WVT3C**_5.,Q@02O&[/\0\,ENQBO1(O#5=;#;$E@._?Q%$N044U4=R"FB*#-_9
P4[G!Z5G46YX X7/QXG>WRHVVA-W_"BEEU =%*@L3C*"PWE$=260,KO,"BWJNV]-V
P&]4PF6^EJ\;L*UEE:+KSGFOI(.$\%G4\F11--#3<Y:0RCBTR:#" K.,'Q T23M^*
P*R\$T%35\#ZG6[-Z3UMJKRUR1+'6@YKWVPL&+/64H+OK-3%ZON6JC(FTS%K S63I
PV7^&+[Q#M+F%Y//1'*,2A27SDRFOB2G8SK$WH58OX)7RYZM#X$!+QQL3#ZH[IU =
P7)J%)F 8I45E*NMAW[9GV\.+2/KIV*>-\S>^CYVW^O267;I#^HT8W:%>-0L_7F_M
P("IE%?RR" [,+8_7JWS80'?30,?<_P-U_!>]P-W:DX9G$7,O(>^U=!J6:;*E#T_%
PVCT$>3,1'KAR"VT1C;'()V!E1ROZ7K7'#S>+MQRU$/PG<!/@YO;XG4C;C>#ER_@0
PBC<X5&!(]&AK0\\EO=:39.?1P55J&R\3F[(VUG8 @=T!Z"N1@IJ:])NY7%;656?D
PEFTNZ6\]7JW$[JUD6<YUK0G32[S"C$?(%%S2 :P.;N-@[FAK_]5OGPLFLLCUQ:O[
P>KE!IG"S/M+!!8:(!DA<F-""*(8H0J?"E>,K^<^T7X,B.IQD<4J PF?#>"1)/9G#
P'*=,O0NH6-LP8A@Y.WM*JU[32&-_0VTA^&TTG!]L"E>]08'SEY''HNB%*[%^:T@V
PQ; 3SK]8P3\-^V??@TV'</[0?T5.)<%:^@M!6B^*XXUHFYY%/#H:W)VR&!^L)0ID
P5]3<9:]&R(3E'60N2N"/>SU3@4G]W082+]5P>G1.O+OW^Z@%6RU@' A"F8:AX#(%
P1U)F#)>/5%[\T_F<IR44OJ>#Y:5Y2F0.^MH=*C0R*]STO:K#?$!FBV<[6+&8GK13
PFYN6S/MTQO*D*MC]]M$GUQ<1Y(%0Z#Q')31J5:J@!BK ]I#W1YZ5(YJ[G:52T^:O
P4>]1D3JG2ZX"Z,OALUG.?[^/>,9&D%V[-Q20W5)B__9MC5LM9?@U.N*+1V8YRG#=
P5-)[QQ60NXSRHE9L<X37EBN;P[G<U#Q^I(!EEMU$#:.:FQ7&?'S[C:;-X;&:3>M/
P',(64]5IG;I6;E?0;C\>Z /XJ5CA$G+\(]I-86R"E,)-8")R:"@IC3VA[OYA_K9#
P5^Q33N'OF-+C]6%ET7__J?R!.VNZUA[NAM>#^9AWW#IC"%YC$M"VJOCJ$!X@&MDH
PZU[>\+;NP+/$$+Y]<H0[23C6B\@3YN1,ERQT\Y]KZ8CK2I5Y,R!-8<E(<7%6PKMA
P/A=06TW"/CS2/KR-6JA9Q0]3%3O]KP>H;AF5AB5@&#[2G(HY88P&P3Y5)ST$G\KJ
P=4Y+E$#"<;:D\$):I7!V$+KHU4!4T8RFH$'?90ULXW)[-%7C/["V2EX:E&W=69%B
P3[0_)N+J=2D3 !6E4M3X+Y4PT11@'&2G-CN*=-;>RB==5,R1 H()MEYVCN(,AK9"
P-D3^FS!_%_M67EE)<,8+B<]'R6WI3.DN3""OWYB51^+6$\<K+Z..KO-.T$K8&6_Y
P,E7&L2IO'6[;7X/8H=G0,A$9_A15_17%?'$_?9T0P'OF]4Q;&.C#L0S\GB;/>Y0=
PUKBG_H[!?/@5ZR)(!XPY.3Y7:VA"<1CRZ80*</4ZA9*(&JL7K2,MSC$SQ?NV.[;"
PV&J[G\((8.Q4&PU;AKN9AV-/<E[62O% )]&,(3'D9+FEPJEU<Z'8RR?%5L 80?ZZ
P-2QTSM:T3LW5(B*4N6OJ.0ECX"^EYO_W3KSXB>[\+8MJ(L%[Z:JGP[8+0)0)'Q=;
PA_>6=!%<W$Q!\YB*<6V2N_*)*G+[X;__DC\JLET <J)-R2+EW=RDIQ3?(>Y38#2;
P'BQ>IN"#%M+8QC$8B-54YTTC$:TR[!1U_VE9C1[KON>'/Z?V-/Z^J0PTLDMKN1^&
P5VIMSP/:452@G4..OHJNB64P?_45[]UX'OJNOJ8/#658:I2&QGV?8U(0&\M0M.KD
P8S+0QA#M ? /+<\(),>NL='B]99^0B(TXO^?CZ=T]]A'*X;[WQ:.C7>%HV.\56,_
PC]O@!E;L2S$=B=&6/S+1ZZGY&/==G(F TAD,K#9D"I]. 8]%8]OPZB7W@]Q[UO1V
PI(/"A">K/(O\K[&K:SO$UK0)[0+52_G9'.I:0UI!*$QF4>J$GY#?8U[I@I=?"&O<
P/3ARK='UOXB/5DP+G"[,1)*$ZZS3X]^=&9-L:=7S0[QJVDI;48_;;#]]'!5WR#>1
P(\, 7-6W.<4\_=Q@OK2!<#9[0(!3>6-O58NRKM@8K8TX!LBC5&FMS^>3N2.[%DX_
P<#9G^]R'^!59EJ>,X1@<2J1@_F!$EPK(\!R1M@Y63$@%6LQ-V3JX!$'PT@?MLWVK
P7;VSC]M_A278RZ;<91R[AA./!$OUFAZCZZ6T.A+\CY6A3&57:VXVX2'1E>@E'467
P0_>HTT^L<0%D_BWT_283KA,O-N_7<TK0#[R^>B/T%/'^6D.9X4.I6+D[<IS'"O'X
P2X4&8H'I*HNEY3T+'$IVY/6$HS*-2)DX]4XW@:A(9Z"'U/0U4W7FK>HVIYYK9GH(
P>C$P/D"+10:[.@0V;\G]J.MXV%BAI#GHK0.I9Q5@6U77#@Y@[:ZY5#-1ZMOO(:QI
PLAM!P.Q&?'(D3U'!EF:%X_0)%%6.SHV/D3UXI.W6DJ)4W;\1BLUQ-!?U-2T&^I).
P4O>5!B60WD3K*42"^]DQL_>T%+K&FKO.7'8GU?E7C.Q5D+1I;Z"AQJXER3?F<<Y?
P#A[A\M6DZ_3PG7G:=$HR?CR'6"HQE+'6SL'#W*\MKFM#7 ?&WT@PB("\R/P<0R=S
P51;04LZW1G3&#^[3>(N_+PL=U9^"%WALQ7_0?0REKH8<(3-\AWCW07D+:Y!F^H$"
P7*M#IM/<RN?&TY8MP/<OC_D@34_9Z0<Z/0V]^2$DB3#D9"/0 )W^*7UBWBO1T$S*
PB =G:4Q"9_ EY5B[#I!@'+3B!;,=P5RK9^.KG6@M!SE'J.L3T2KC94I)'WML99A*
P)-/H[B:S;12.V4":%F("1),E"\6C"4Q%^-U"79Y6Y8&_>J5"%1!YTHT62FOBVO\3
P[G[N)7?A52?R96_L$E[RV>9W,[QWNZB&?([1;)>H#V% A)'7BKR3!+2O@['M;?[H
P4V,Y*I+434YII,M3B(I,\.($"=[Q6L/D4S[N%\*?W(-9*^*:4.D56E28AM4F8;&4
PK-BE[^C.X)X\Z>9X,+/,C75[8Y5_$$\(5V[40/.M1>6?5A9I-JQUF?%$R*'Z<%O8
P45K(ZCCW=P7_-O X4B*:_BBD;AUJX=R#M[R>_6"R<@2A2QQ>?("RE$0YU88ATH_N
P)63>@D\\M*LG8;C%K_-?TNU;]2^P>%$R3LIJA65\D" :35R"2*)X;(7@>>3+A1[:
P[W(7=M@:'(W-MN;MSN9R_J 2Q2.Z@V:7;:U053)5:%SQGL7@VHX4:*6/+4V+?CMF
P>E?I0)?&C5P54L#HG>Z#)UMTW[=$&Q&-_NR^3WF[N0[.=&))#Z$#7+>,\V(+I;OI
P\$</X$&7$2.(\PW(CZ0,^52E5&N>EJJ-P9DM:5+C5TQI3Q2#&GSJ!;7]#C[3"BT\
P9PV,9-08A^8=N8/*R;>F;VNGOS3/-?]U=M)5G'%V('1*\4,2+2M)/ ,[&2_@V*_4
P]1B#AEA[=&HX]L?NX;U;AQFX "DFQ3-^=8N01: '8-05EWF]@E^ZSSO2Z/A>IPN[
P6W&"<76IS()+2>KX;.'PGQ&Z!ZA#\(C6NY[W_0X [DEF]^+@,P[16T+O0ZILEC=:
P: O NC@<;E:WEJ)0I TY:4W7Y*=\5+B?TP--D-&SK#3Y\>J)^QRA?UKF?JCO#7.#
P^SEIN:P;6/2D\D:O^2R1A[0N%3Q].7O9I3YN8180L58P7 R, 54E"RLLF=Q#0\\ 
P137W'"8C>EUA(;%A@/5?S((Z!?>L$<?/!9O3>4]H-?V *2"(%E%/S4J.\+5[F&BK
P/^$F.!MA0:HEV+T:*-Q;[U]6_^?),XC5AE,:O-R'0;VSJVZ!(UXJ8ZYE"1LL!3'K
PEZ2U+ CR=!)PX<Y+C:]WBKCC%/O LF3F,QGH7^?^336'5_!4$;"OX[URO>+;X&>@
PIV3ILEZ"?Z>@Q6I685Z9X=:ILP54Z:CV9?@(!;#N;:;8< X/<XMF&VZ*RKD<Q%DD
PJA_)<.@:TY =J^#_F>&2(@IX#^1$0I$R^$JB2J7U2#;F[>&P+TSDAXC)"H__Z#]*
PL/]RQXPELDO?#_#(R.=9I:[1(2"@OG<Z<<SUGPZ)"PL1 X>L<T8=?Y"(+2HUAJE\
P!NK5:5574WH_SX!KJO=*P^P]$G%O95>G_$*1PTF.='N\)*ISV%5D52L:VZI=5;-A
PYD9!>(=T H%&I9;]3WR54UT9]4-CFC,392?&]1#+$<.M?Q9C^3)Z*XCP$NY%T<SV
P6[H6;')<5*H*P*50<CW0:-V8GG6:%$A>7-GH7>KOD%*.JW-%-O:!-8C1E>Y8T;EK
PG#KJ$?A.GJ95QYP%&4,-H]ET%U*%N.GZ? Q23.0EP*QU$&(#20E85G?6:JN':/C%
P:9"-9MG=J*P!6J- =.J^(5,T!=79I&;6P,\)/R)1/"&I5CW4-DE>G!1Z+6 8W5#$
P9%5\/A0$R'?1VP[KP+D=$O;?MG7.Y G/GO@2RA&.T'VW)(?3,]B]Y_VTO\[%;D[=
P^8!P=08-K\DJ<<RV'8/W^L0->/9J6#C'@JBZ^_9^3XDZ3P)Z+%F)9+T]N"X,!C[K
P&##[AM(C:UZE2E165R*^_\Y$U:JUOS>4PC@D:I* M91NT,^&>N\U&S1= 7!OB:6=
P(H:-6XS(9NLA*3Z816*)*MP[5 ^S8W I?:ZSS0#<$EZPG/9C!<87C=)K(FU$/7XY
P7G4J[.L!:YBUE-)SU5<@@K=[9',66I7[88?>:!XUI&I:;)OP4?W?-V!%<_$(0Q\*
P1=B9Y/^S%M[P"]2_V(2_,+$%URP9(Y&D<B]"M+BQ#3N>SJ0.:-P6%:30\8I/S#R%
P;C.**AO3W*![$*^+D94>JD"UMFF$_0<>514!UV I.6"]"?S^LF'&331P/#34=>G6
PUZ9;!UJ[J_$> S8QG:D$((:^/E6>50PE3;"X<]_*A7K7]@RWV3HP4-XAYB7(TRRE
P$^[*K84_H'YR&D4N&*6[K//<83BP3$M\7(K_ WS.C4H#F%]'Y8F]WM4S:#ID_-[_
PZ[/W=G>I\:%R.JQ[@'47$=2&>1>6F BYJX?^')L;D6Q%:57^LN(D>4[#C*@5C\V9
P:C!@??D>8Z3/G9PQB'Z\EJ>!NH<_29C.\G6'!ES?5T[X5$TT&??&W'-,>LW(^@5$
PUN?8D,+'7FK/A__]C[BZG$\-3M@:,KJ5(*?[[P65]/S, F7)!8E34KW@%R6EY@:C
PF?6S4R)$L(RW.E.O F'D.K9@X*6/.K^"4"95<C_WOR3 &%^L6$!PY,U@E.$*(G-E
P\)8PULUS 5Z8:7N/U&-J;,O**:"WLGXB], ;CD)_\ZHE) ZEQT1=( -0E.-:KO7C
PBH=&X)$;T)\L0:9?/L^'@2K?&++Y8=F[&65R:KT;WQ7O@;#J#9M#,)$0' ]M:.8@
PE!NHT:,V02_*&VAM5XX^-UY^9G-NI&8ZM$K4._65N,K85"+MS;ND5\_&-TAH)$($
P'MP#YS&O5MW^P"1[A;$_=]JZI! 4I"U<:N<@/Y;#)7S<PXJG \\/B+53G7[:ET 4
P*B;KB?TG=,06ZP?</@B3VIS6:_,47!<(^]T:E"/QD45X+-+W,'/KT$LO^1-6:Y(M
P?4FM6!,1?[)X^RO"0RGZ;TP9B<AI0"K&))YA&]G!T, E.GX)C+HG3!ZUCOPBJ\UF
PV_K%L!;7;8@H^W^LF^<;S>%%O:)_Q(EMP?2B^8MV<<6J)=]=T_$D7G:#ZL'_L$(M
PQ *\9$%S"NOI@?%<>^1]V5FM^USA<[.TB0#SN7B]*N!5D#/R7QBM*#2?_.[I"X-*
PT3&T2EX3A+G?7_L,U8U6/I2 $Q=%#,7@$C8.[CB&!0-8LOI$3.UY%82:06'N3234
P!(X$!Y3.Q*:MDPY [UT]W"Y%:4[V44NG6HZ^N5ZBJ@_0]_D,5O<0I_;\CD60K!:6
P?)!$^([ZJ?,>0:$ 4]E!2'XO5Y[]D^5IL3Y1B",4EBM/?^Q__8N"S UOQG)ETSJP
P/2)(%B!L]PN!I]<D*>5V\CB$V,*[9B&>9!$!J]>)UF(?="M!@6.CYSLQZE-@9;V&
PAC [7 BS=9D-%RECL3TEBH%=D6 #I[@9&.'XS#9^S);O-6DR%GJX&*4MJS!1K-3Y
PV7KY'\11L'&SYR--GZ16+KAVTG8QBLPB O"5T?>GYG=Y3#C.G1Y@=K</08-0S9\L
P3S%[1AK-09ZIYTGO'#4N)L-)5@R<0@JM*@0@@6 CJ7&=L 7#IM"'R:=3%M4&O1"[
P3K9VM_(RRE+5#^KFUE91)L!-@O <#/(D3!J1>/<Z7"#2]J"L5F[G\Z(R*IR3J_0Y
P4^A<A3DY%BU[G*8.T=^6'P:Y>1RO&M3SRXXBE%PI!^IV9[0_<LG.7S=33+6!V:!^
PAI3B/78&UQ)0OCZ79VB6DOR3I]G\-2TR.K7O"\N;&9()N?&=V:2?I]-=YLPG3S98
P=RW$4_9?#OJ0DEGU*&_I5;I8O%9$:@(.UF;6@1=8@Z4"*8F'K?B2!GK-5AU>-.GN
P5@'1?YIRMV)HF[+D.VB)A[?+8N:ES)K$%9+ZGDOYLF>GUL!PYM/6F5$\_4?)-3:%
P(XOJ7<$LCF":[)?_@L:M*\YJ>GZ5#3N]T' FV3JY5)W?G8IAURDZ-#YVTFX%R_7V
P!<Y ]U=_PE2:8G/EW15SN>%?MH L8VW9.<FN5QN1.&!#1,EPXOGFHM&VX(H/**0*
PXJ=9,2_H>5 '4QI7$SM+Z  '_X?N[5J(I910,3V%.TI48JW'K3_.H2 (& W/#7@Q
PF-H373IA+9P :U(Z&$>N,TA/P0FB$_EB:6QTSO#XRWZ@>RR?  ,O[N>R.)X[^Y-/
P'B H>%C(*G-\?=822SJ> 1+#GE@;F,O,*+ZY'O(SW4OM(1.FNQ>I6+".RMHX  QG
PXT65MTT>4)JD57;ZV[OJ;&;+;+B&-O^8J%1@^LD,;%!>&EL:-VRR]96-,3WK@B"Z
PJE@<\3'%NC(>C*=J9HK6")BN853OW+<+(M</-/C*&-&U5]I.SQJU[AQ[!GA_P$I0
P!3WK4Q.>G8\<!1RAY;>\)%HWPE1178.,EQTF/C..) 8(.,I-W<7!LM2=AIG_*4 '
PRST+V8?3*!(#/NCEZJ8U/^)N*9"XTT[G]POC]Q$$3T6,KPU^;?>XZTL#,9/)^K:8
P?;7OY,H@5H.].--;(\2O(>B="(T0BC7(,Z0CXJ/2W Z(D70\C48_:85+9>#Y:>O"
P2*)L3+QN+;/O^B,0V$P[$UQ9U9&=>9D@U\N^; ;;?KUW1]#JUM>S5E @N_10F>IA
PP?8Y6T::<>5=W?^$)M_'4SDI8EZ/R+2;"T3S^J#F[CGB2VKF;BPY#YQ K1C[YKV;
P434M>TVC[[%1K[<A HKN"P['9,*)=H']H-$H4 U N_\-Y-O=OR;="WK'[,?X*S6[
P]H-(###OFS=QVQAUB@:;^_,X?MC-#(2BE<06X:F84,A/@ M'^ND4M":B6 5.D![_
PLIN6C*4,ZR)05)_V?(NT!79'E2S[ T[MO\.?GJ:1RV[0[D9YU\YOPQ1'B>EN@@#_
PZ:I;I5QRF0I7V8F^%J:$) BE E4,*2C>G$CVC)7>K(G@9;^\]3[/"X9F>8H%!MJ;
PGI,@^,&F/#K-JKRASEU7:VV=PY[<1U,9&*V_%'CNA0$K7R7WZ?(ZL:6@+JM.3MV/
PUU$MA!1G78Y%--4AFZ8:A6?=(+2^R$4KG(DJDBF-U('66(K+@'IS-0?2M1FOIG)W
P+K'+R^F=175<;"XAP!JZ5 0>MP(!;K%=6P#L?3RQ$8S27C"'\#!S3)T3!KHFN+L"
PJVG/QY[L&-NB7ML=?2"9&,PD.U.&4N,=4PDUF <6+B6'!X.Q:PB>8JZ0$3=XE3?.
P_6HL' _SAUB/@].U%!#/$MT?*E-$E?_0\!HY,&NAIPC9#'(%$-""@H*Z;:O-)=4S
PG!MDTA NI;"HL[&_AD\$+R.15<VX3LCT'(0"ZF _V"&*LFNGA%%A@KQF_04O?D'3
P2U96OZK@PLEYY%?5!;/+:0EB?#+D(Y[+1+_PO5KB@+ \M()Q'<BP;%ZK%P%E&/O,
PU%7]KRP04B(!^.TFQI\8.!7;IR8Z5MN#/ )C!]!4C)J, &F)-THD4X+.Q2203K0D
P_;UFGP<*C;3]#8>[L/S>[P=P"PO&EN+:+K<Z  9M&_J]]X8F2X @2?1UF_^CJ#"F
P)Y[J$?RIKD:KANS@U?A>+DE0?*(:]7T7O35Y#&*K3==)_<D-1_'HV<*/O)JA,PP@
P(X]"F>AMW\;@?9!09*=:6(DGQMU3G\!KK<*?^%DX9(2HS3S7]C ^\#>WC6I,$)1N
P(7PP83 6:^<@()<FP G"]%[N,0&BN_+_,^,\\ Q"YP,()^[5\,@IN:=\,S!:'80#
P\,GQY*IHG>KU0FHJ%;N@]5A+84,,=ZPM:&J@303B>6+FP%;NBK9*A'B7 !Q:EHWQ
P:3U+8:Y!P"$5?#YA!/HSGW(T^OZV<X,76U,SKIR,[^K%[QM<SH>SF9)-"3=6BA6L
PWOOZBDE*CN$XJ[A6PY3>PW_D]X.5<S1@+XPHD3,=*H'\O>&+5G[OIV+3>8M=<B8:
P?7/["84  =<_T7O0KSQL8+6F;^9*;XLW1ES7>Q5MHM RC3:GKC#(!F\<ODM,Q<S]
PD3LDM\T]5:@ H(KOK*OFEIBRXUN^VZZB\\ R8(_8LAY^*YU0[]#-:\8EQ[,3I@3,
P%X4"_* >FNU'05.W7&'"HU9KC)HN-8B_L"_,7P<$DJP70<-7"LQPF,3K+_EZ1C17
P>XELJ8M@ZG/VC1.* MI0_/KZAFDK<RCJP9!2DT)YOU59/LYX2^"+K(Q-B=:Z8&_>
P ?V67MZ;B@U5 :^F.43GV\&RI7S QL+I(1/<N4 -[!!T8^N 7K:P$]/^Z[NP ^V5
P#W >)K28'O3D&N)1%>)JBXK_4MF5WQJN)[6G$TOFT?T(*"7E$?9W"PZ&&0PD$5>1
PD]?!9(W,=C&N9YY+5")M)I(<^C1.>C@Y4@MRFDTO_0=R3?#CRK_>[[0S+RD&Y-$P
PZ:$H64-_.!K:Y6MFN6'*"E'R@Y+(,.VI U>#T;^NB8IDWY+G?T!=)&^ZBPG;1QL?
P6]QV(;8JP&_42.].L4DN#)G8<WXDW ":NKZ15JJD6@3& OC(EKV5YU/(7^\^=.JZ
P.XXJ:23PFMB[5U<+IS8[2(A;*3CG6!3/]5*#*?-_VBEC7.VOS_3PZ(<DO*CBR,-U
P&WG?>61G90J9Z)M1" B^>:"/Q]C>Y4^.[GS&(:%9P?:/*@7AD#]BUWPC8BI.I#T>
PT WBS+$68FX3#.(NG&9GM)G4A0&S<R(=MI5VG6&C4"1Z)4WP^G3JMR':<B\MK:E3
PEK+&5,^4@.HV6Q86QK0_?Q>R/76,JN?T$I,G5,UCQ(D?1(42B2&2<U,I],$Z2=T\
P[CUA$*VN36 ![PC<^T69)9/\F V@E[:7S-@J0:-^:00,;%.L@577C(_8O#X6(E2M
PNRV=,N#(2C$5*O$ %XIG/F6D@#U(H6SOZ00D*R/<U,TK3H/U94JNY7:4> -%)$4[
PO_\N'D[[2&S!&+%KY^%I1DFU'PZ0PTB=G&8RV+M6JP2LU-APHCC+!LLW$NMFAZMJ
P8)%H4SP-H#)3FDE>]M:S&J<0CW T5?5&\WJE<"F+8Z\HDK@"L-[?F/7!I)JG]>I?
PT%M5_YS>K S5BWG)\ \Q0EXK%D9!D/V3=JWQ8AUE''_E%?R@4(32!%DQY<- ZYV 
P)"_9];M648[_? .O4YMDY%"BEXH&%-,LFN)GK%8E.ZV2T$PYL'&M%/($Y:J.VRVO
PQ9[=/[CE?E^YZNVW>6>@*N&. <2)Y51K$32IH4)B$MESLDY(@XL5X@^KQ4+R7 GI
PFU:#NJ=8 MT"];%I$@/"6UW3L7DP+]*&6B)UXCYL2*X7*%$([1%>ADF6;_"D>WT 
PQ&9$1>;6UK< 5\U+)MK/L/.SCO!2P*2)<_L> CP1SVFO[W5P>= [GN:YMUF,1[_O
PJJ69"L-"QTV'2W9JLYG:OA/;\&$V&34G+:$="6 _[2*ERY?0RI>>1#" :*EU_5N_
P,.6K$1;R0EE#D+IQC*MH*,=-6/;Q:"9%R"X)'8BZ-G#]NY3F:.D2>/-_?($OI,^Z
P&Q:M#Y G$Y+[\8X[)-8\.JALMKE 5\AZ2M:F_$H\%<C[?:/I66,70J,L@5Y(T-_@
P]]0^2_5&S'\2-N-0=CHO&]GN>W[_TF>H!)@>X*)_JT<90/P1&^9)^W__N:NI91.0
P_!E7\W4+==2<B*5Z<^-*BV8RPO0E=F;_/U]"8[M22$ X9_O'3<N(T+>AJ#I50,[>
PY4-6U RC&].^^.RF)SE-$F,HG$O YY!^K\\VA^LHB-1D5#2O:6PZT40F<-/:*E9S
P;ED).XSV_#,#N"(%3QYL=/G P0VZ,W0<96J^F>O_U%J]WXH#0*/[AHHLIO3Z'/5;
P&.<5&4OV(#XKVQR@41>R:#^'/;\5>".V;/=6HW+AA 7MP]L^U B':!53.=>NEZ2F
PV!;-7P,"?<VVF'7!-S0V$(/L@ZTP/FD+KI[R7W)U4$M=^660SP/<_F8"_IER+3];
P?%:T^=$16Y$E[?V/E*[6H#(0$="RXP<Y-IC<#MLC>9UPMNW[%G@;U\O P8M=6D>9
P#"?.K[9?8N)OZY8<2NO%!V/)C#X,;\F^P[Q+NJV9VU68^#B&1M>"'S.T&X>_\F%)
P9Z![K0'>KW+0"GQ@K#*V"3H]]-KX@[L,>@[RM>7236:2?3V9#9O,'8J]OS.0%A+N
P3+PNZ=4X;C\20HP3O^!6K>5#JS-]%R_A;\8P1&*751E$/6=<_2&V?'^! EL^=5=P
PDH,4ACA)CX(/VF[3'"O_T;) OD !_>AN5;J/L^G0;G*B75& P'!^C@&>]J)I%*A,
P$-Q.U(J*RR)U,D?N4C^P";I'SB4A^L/=*Y-&^(,]3D=(4@JN43-SFQNNIF0;/04-
P$8Z!6& '-F<-Z[<,\D)NC,8GIZ8\5TZVNWW/E-T>KL28,X64K/.HHUIO?RQ>[NB?
P#Y%55-E<_Y,R*-*UA3S+W9DN1/,=#-5<R= )#>A))/BZ^__%XO'.NI-+!)Y>T;7)
P[8E1:DHP+XFFZV&%=[YS]O,@>ON4$CIR%/HHFP\4B'A6%P/N Q<.71N%W\F!C2V7
P#]T]M46$^S)>'%2D-X3<K?^8WDRLFSDX< (T4:AFBZQ$Y'#M"V7(-,MX!S=Q?^%5
P.Z_U!O3C5DX=5#]X<*?LF_EEZQC=)S'QR:+?'^6L-JYL/)_^01Z*$XUU71_.V]>S
P]2S9Y0@L/:)EHI5)NX_;;60YC@IA?Y,3[(5(/0U_9W=^#8'@+JM=)11":C CMW%O
PF1?G ;)UYV4P_$1VM/3ZP.RV50*Q*B&7/=,%1(P@\YI6SS<I=B$!RE(TR'>73')#
PY^%Q*[YYXWD"&P>IG8*;&$X:,,L,^'A;>ZEQ]E6WV[::[@S.&ATLGN4K\3B@9TAG
P)5LU!M75'E*2X?7#7%G-5D!LDF\'-*OZZ?HP<:3]4><03:"AU6U .%IB7/^Y_N0E
PZ#R((<'ZMLRG&G:XSJ>624;MP5@ KOTW\I_#:JHVE5F(50CYY .I2B"^U\3-7LUN
PU\7IA8;:!G6W?9+:>PU$TS#EO1X_%9@66$^BKMUG:,*.RMQO>*PF@'"N3.:.8$AW
P!=3,LC8.T)JPG5,3JHZ%^67SI5A)J*-@-NKD.!Y_W)(\G'0*?%%/*EV?58'^QOOA
P@9/P<:R2W6NC^6VG%M4'J_HQ2HZ:X?K?@5'0IB$/Y!)SQV4!$#IN&YD'%VO*P_H-
P1L6_%WA%--92WUIL^NA#[;[!0J+<L(]9;DYIJBI0[^D:_8[GO]Z9PL0(E*%+[/,$
P&:9-;SI&6(4T3,IE9ZHS#64M_9JVB@58:HN&Y^K!%!\WP($MJ="154VQAD'=I,24
P3"W3&1G^*4L&[HA]8V!T4^':SZ1#'S+&!$IOCT1BK2QT+@V]ZDDP0]9.0I86;=_%
P7IH4L.-R$3L5O),GC&H2Y2=)O+>L-"(&)N92AJNU<D&+\$G<UX7JELYKYY5/A[%Z
PS=X]LNE+N?92S:-?W8GKYBRI'B D@O5#C_QZ8#8ZR$X:('K9A&4TQUO_L9*D"B5X
PCF+C>@*M?.FYD9U._(_G_(U3P/26,<C/LQR4:$ZL^DCF!_X@H/G[),J8YG,6B;B 
P>"E.83&E+>9B#'C\H,74Y$/(73*V[[Y)G,C<TCL E=D4S[(DC5=*H+^5O4AHLYIZ
PU?NO@CA-2Z4<" =OHNO-8L:@A _F*EWWCJ#2!H?T[@VZ[Y#.ZME07VNT.R;+!PLB
P6C>Q-:H2*/V'QP-!RV3B0YGE JI;ZNA#DL""& K1Y<@FSN]VL_$J&$%JR M?:ND5
P\,684[,"@)A8M:EH4]4<9R@#^PZF15T4)=-G@3B\VYTE^*B9=)-!7[K)"O*:W")%
PJ-P)T%!<ALZSL_VT:O!^ZSQL>E126[>6'-YR]2]'J%),?T%;7VBR][J'=;QQ</'Q
P0KU:L&^3474A:4 %#XR$T ">G?2R6J<*OTQN\Z.1\00?4A9T=_CO7LP/@<9>K&[?
PVS*?#[S')4H%4Y=<1*J'XS7>BN!:>?8$(O 8^/E+/ 8-\,,Q],5#.J5X^Q_G6 T\
PV=7G6@SIES]G_NU;U)%8@"0V^>VCCOL$MD@Q2TS[RZB(11R6BF#YQDB*?E7+'$4F
P'_M7TG K76C@>0XSNZZ6")1QK&)-,>2D92,*#+C6H/9.OEI%8LVW@$$*A:<;$2\C
P[YQF>+YR-2-<FO950I$V"Y$0A8#33I034TE[EKZH,@\1GE;?\.7C&[K;T?Y<BE<X
P^^VCO\.&1Y8'B'Z<;U'3^4* _R"7QS?VJ-,?Y%T12.,2'%SV;>@55YGU)<5X=5R>
P>\SD55ID,3':$>52%@%]"L"M);;-D(U3 %1GGSY=':.S6":/9*J<Z52.YAA4,+:F
PQ+MIFV+O?]0:&V^X>1Y7AM'VIT@:X;U(TWS;8"":&O1#+?MD5<>^:1MU1D>RLY?;
P3LQQ34R(,;!_$.-!F^SGT(FZXECQYQ]DY0(_O9S]&]T7RK#YO5=3T48T3,Q?*W>8
PU%Y\O2@!@2FK5OO+ $- REX5#4P2EZ3IG"-I^Q71C0-1;I*L6_2YENP=&I,,Z+#>
PIOKH0W<2;TV$HF;HF2_E*TA#@H$^6>+V,Q2&>(>Q0O1!.<6UZI&: LE^]HVO]2!V
P#1UH@SK5^7G_P>X-^OA,ZP4XTY?D0JR,B[CW$'32[_W+'C! ;H: ?!$^]4,HJS7I
P RT(VXVJ&3 R0!&M:##(IR2#O.]_/.$G!!IH5Q2(W#,#CQ+:J:0A\-W'I?,<46-C
P$2@%@33A&]8F" =9I%:.XM_J&[6U7P+LFK5:2;9H<C$TJ"4 &+612$W0IB_K#'[Y
P-5\X*PH=37ZT)&MP7J;]-_D)/MO+:7G.!G4"'UXI5#E/7>HY8-L65IZRI\\\8D\4
P%8%\D#2AM+,O"K!ZA%XVEX5;Y.*:./U;U;#SBO&/)O3FJTO;RH@#VFC)F1GT,5;3
PTDIJ:D'N)5MO?+7_F1,FN?WFD&J,W/]8N1XT'RY]FW[+*<1Q&8)B7B8I_^1:U3&-
P\'YOJ$)?H>)+RL""L]29Z,)XQ>%4$*?8PJQB,-7AM(,B[$N1RQ)PV3:>9%!HL*.=
P1C&$4$27JZ"Y$^><)/]M\#3:1*CUFSX1T&+Q[!6'%;U-#PHXKT75O>I1UYSG.J^$
PH;7A6[JS>S?%RQD:*B6.;Q[2]A%0'&L4ZA9T)8*4&BI+?ZM5TB_2P3B*O=#IE!!O
P!<D4829'3L(-#/"R?UA937$YT6 X^BQ1\E7C5):.Z[2O@V/#L&$R&=^RJ!P8?K)Z
P@QH$'Z?T;:%_F]TW2 UY9)-!/HJS^0*$=G4!QZ,,,6E=^U]0\Z6&(X0LL]@&X_8Q
P!(+V8IKA2*@!)2=[O*\[9V*7]54D7(BU^,Y=YC._1MP#HP^(++_K/@^@/7GH/8O$
P<FELF\AL]2 RR@X;99_=CKN]F?F>%R)X9A/!_1*7F';;[?KPP$.8W9X1(M1XP&/O
P[Y%Q&O^C-BMOU]<4D8D2)@;ST4(N*HR>6^+!'N3G?H[YB"TA\MFJ4-9::^"B: ^0
PT]UXF-0?UM%*D;-HN+J/XE<;ZXDRY*HS!X?;'OU5/VUX%HW^J:+ ]#* <\>R/[D'
PJ2W'SS-#GTJ5_>P:NN ?;^$*15*KRYN5\45QV_E/?F0KN G>B[E620<ET=4F$[\Y
PDJR5DA3^=EHG9V.]F0G[+1Y0=HL47J1ZU=MC=.ADV1)#S:=C,G9_<$AZ41YT3;U>
PL#(ZTL2:#O1&07RAG#^27$+IWHMBU#"%FLUYPZ"T(=C)&QVL\;]>/@^7XIEYK###
P/#,K8VG\!-SEQ<[N#[(B=*..Z;OPVRT)#%^PU(Y</O:"Q305,(,\]$2XBY/]8N7U
PA<S)P"Q \(V+442D(\6*^:4<J6 P]D3563WNU'4'?5L3$>4#ZW@'K^BV==:LJ;T\
PGO:'_XOJ'M9#+(&\HJ3+)F6]S#BRB!2Q*K.IP;D.9*P313^BCW[GX+-,%N<$VS<8
P*\YK>(9FM#^KP4F\3]UMN4?C[(YF;C&3 +BEBET[DY8?<([;_K\#C:,BS./*(!Z'
PG5I0LS._!7 _8VYJW)X+-D"40C>TA?)X!["S*8%EJ%\:\P"VI383XP8U5, L)<@W
PO0J59M[QQN:M'0(YN# _&BO[.G3(NIW-VZS(!@ M]._-U6B1LS&L@-@P/ NJ$6?\
PL4H&&&+\JG"/Y9XA4RTCS6T#ZB8! PH?O-7(N$#UXH75XPERRHVO_FJ7"!WHY^%^
P7&-7A/I4L-4OE:7RU2W9U5\#.MCC.DA@6J0&5/+IC3\;HB:U4[^$.0)JMNKV>''K
P^":6.C4YR\A55QR5'#/HP]6N5IK@GWZJ?Y[@<:LHTFNQU#PPA%4YCMH#'*E*&C",
PJT"GT%74XWP7"1*;1)8*B$"&!8"&"C%9J#I\-EHR9P2F^8O=;-W+@EAO M63ZLOJ
P;]4X>+G*Z(U&:>GC+&O(.&&J]#4B0+TA<(YK)4E2^3WS0%@MQ08.2T8&H$XRY<!Y
P]GWX9=;$X:VY<E\/(EN,ITX3_RK+OL[E;"+[75!O964?#16V);U+85%R+7[D[P.5
PA<\P<#RQJ@L:R VG6V@)[VWFY:-?G2> M+9-)"WBQ6&TF+WR6.H#7\AY?3)35/SW
PMYG<\[6^&;!3BN=H;OGRE,P0 -$YWTAPS=RX\%+>Z>63KZ+913T,[1T>5G95&D:>
P$)>?CT34$MV_W,%M9D [()D+:R(+DQ5 J1^5!N" %A0!..3^LP^E^?/ZF#P+EGS[
P+06<[I)4CC*]0%G'?#8A5SC1%U><()H#XXZ)X,((9&D<.C_>DK3IZ"B &KK'MQK.
P-[?>AVJ[@=VQB*4X\#\H/;&]XSO]?RB8&T&,U>[J+$'0(%V^C.&(]$Y@V/BWR=\R
PWT("W/$VS;G&].I3ZMYR[!T.P [N6J620>3M)Z_0M^T($U5YH;]'5GKY[+A]_%3'
P!XG[LN/?&!0]L'!@1R[61#1B@;2S)VR6>$=XTR]H4,$LGDX<0='G5M3J)1>3?<T@
P[)B8ND5TM]R*3E%K+3*=+.EEVZA-#$%PSQ'U".3C[1[RL?.-8\DD<)<R"",1%QD\
PMZ4P2/W\K5CP?DBV0M261L4U 3:Q-IA,HURV]7) "W;/?!NRCQ)T@E2^!>6?$>+@
PS5+:JYG#%DX&1JUO,I/KJJW>[7G2;T5#>M9[! '^CZ_VL[A9SD<=?IUHV.21JEK5
P;+*5-)II'=83,*"IO7C2GJ=ZYV(??]$05J6$A%P77(%%HD85M)P>/<;*7V;@[<Z'
P1D)>&'P+>F<[_VX36&]1?L:C3 [Y<[0F0/MMBTFX=%YS%?]#<Z]/&XUN"\E<'-S"
P6/.6?+^E%Y["$,OK>S@F/BM?O-V;&RSM[J/PV<:HFN$S?D\!H\&S+!:!+*)9XNP<
PYO+<XTL5##S3;UOW7C <8WT*&GCZ> X]8SCR=%8FB#7L%R>$R2'D[*]ZU@Z85R4E
P"P%S<EU#/Z0U^4G0EWRU;,&610&XGU #H4BX>XNJJ:D%GCO[.3) <C@7BX5D(RUP
PPVJEJ,(Y6FKACHN0TP[%7K/\R2(UO+JZ):NIO<JR5I+4+!WI!K5BVYR<."\ST'Z[
P?YI0Q= '/U>C>!(CMN#+#5UDK=&&M:\&.X<F<;_^)69+O03Z]<"WBZM#:'Z)F05_
PJPZ!09I^*CH=']8A[Q'$H=GL;Z5Y,OPJ#BDYUK5:I"H6^^[;/8$S$0ZO!,,H_PDR
P=V[P:E..N9^EA2EAQV[+N6S[7VY^ZV0UQ?+XC*6VUCG?Q>,GY:=5JU,ZD['T%M!_
PN4?64; =.4(<Q(9OWE?)3G'N*-XMP3!V53&'.._VKY,V%,AH'=%+=PNB51%N.%4^
P/)G]6Q><"9-,8KK%9C).W+I(YI6GYG]O%FG^@KX9!G"*'X4&WE>_G^M2(<>XU:@0
P]5S2EN 8>$I]K&RV\(I+ZTN1,E"[LR05H%JY_+.]=-=EV]*#!%8J.AYW5 ,3_Q% 
P)' PYN WR90'6H&R)(JB$\KJ9<&B 6J<F:_9!8T02-(XXM+2T]M86#C=MO9E,A= 
P]K"F@YJ=??>O9,'*UIOZYK]C/MH!+SOO70\=SD481!#J:SSU7"$;UF8OG0.IFY<R
PYOF\-'S1$JP_[A"5=5@(="*TPDX1-JEN]*8<K"286&2(G>KV>@^]I6H2CWM>8LS/
P"7/Q?XQK"R&0(PG:,KN*-D!@7"!)-]:^_9#<-:N$ 2DB1D66SO<T*6P0D>@Y!LSS
P6P3]E5R&Q6SX7U/LH+V1.3:@,@.*59RNV/"_[RE^.T<GV(+P8T<TX?!+5'85^QB1
P7,DU45K8 <;G)($WE[PRU+6-DL6Q8Q\U*RK>PIE!,$(YCQ6MVNX?=W<<4A7(AFP.
P-S?A"IW##2R7W\IGN-P@ W0;B0C$1$K#0\@<=J(O8.2^DXL2>6W]14R03Y$C6D2(
P/'3C-TH^3:*'S+\Z#/<[.H2ZK1*]?>^\,T[>7T41&(U0Y0,*E>*^.-XF3V_X2]D_
PS OEZ[K /3L1@*H=;CL\6_6@%BY[41-GB%I>E@2>Y!;=O5B^I4^/([^JQXH=^^P3
P/)1T=N$J_CCS<M!! @UN"%.F:="1G$S8;LJ_[@9VGRDDI-?*6KG>-%O[69P1*G6G
P^8I\Q_"T3\<%Q7O-L7'&L0]$*''2J/&^:K&?&L<'^+R5!PX\8%MS7\,MQ)^$ZW?3
P%$R^_^+6=7IX)M>VDJ*,\?8BBL BXTCZL*?6Y/GO99&4ZUZCFY:=U0R[D,0,.G>R
P?*MM&")+:2$S^NXZ\*B,Y2SW/-Q RDL+)1./ 7Q1L7TZ.Q4&JZ!Z9,?9\ SBJ>Y,
P5.2QQ0$(JGLT?2!.[>6*DU51GUTTD0]*0NWX'2XSCD:5JWU4BI2T.4XJMK[*-$(9
PU5IL2F*K@ZV,-'WC'(T1$C9\AP#XIDCN0K[13"%H=2%PKEDQWW;;9A@U#X73N5:!
PU2L>F\AM'H$>=<M*3_F$2+FQK7^XM]7F<<V G%$U#$%QU:0;RK@.&[4.\7%U?XEB
P5A:<(TZ0X^[K3 \6P?)=U/0^44JJF1#Q_=)XP[U%T8=<.FH.%>14DK"O)@N%1=^0
PZY<AS&L.Z^(,*&+:9.WYZ6\0A"5ASN"1<KR5EW?P*K<ZHBY^^<;YTKY'%&BI"P@L
PS<*%5L7/T=K3"-\M5C' \)7/+\:'ZR[S$8(A6QJ_KI5)R9<A)8PT@Q'T5:%V*>ET
PO]56+A6H2>LFLFY[&O5=)) .R/J6VP>EA"S\ R^@=F,7B-U*0(M9=[0@(QK"S R;
P9!WH9R"-5 FNAGLKNX0@I5'-?_Z#JV:O($[\5^C8S5F?BO#TX0K\P0ADX".5V?D2
P3Y4/TR'IX5!UX]>^R0M,I1$ZPUW3-I"!V)G<^I,#&&,/Q8.G83(:F;@0$3M-#2ZI
PRT>R.4*;^(Z452>\<=[\OQ0[C$@RN!C>6/=Z8G-^LA\3=*;V\^/K4;DYF"JN)V@Y
P.R$WZ)8O/AW<;<5M.-\E\0,48*QI%C*I(USM[-A5$PCP$[<][(>2DN1S:^!FHR1<
P40) !ZB9);E<.3?E>=C3QNU8CUV==P81K6@XDP[:IU.%9 Y%B]O$OC-+\16Z;>]F
P2W'3 -8F-H3LHV7(UN*?"I'8F@ZY?\P--#X/JEIS<)1:GN$HV9OJBIRB"1T%R(/3
PN-28)1<! 4I@I>\SAC"8_YR#.X".N52>&(ES;'0Y(_-2%]7J7^\K9.AC0NNLB76$
P<RA52)K>)2@M9?C9$SJ"SAQDII$]&@>2P;PI=#^,"1),,889(TGM*0,&A6K&92G9
PMT3&\5E '#C_GY-DJI9]Q#*T\L)@KA=]:7F1VB?S\Y#N3-('9?5U]$N/YK<]Z]_/
PLTN/?A5.Q-OJQ-,0/YE##67?\XQ]C,XBAD E8WUC]@-1D9)R4+P:00J.U1I0S8H<
P775=-57?%7 CA\(MG4=&\2Y$[M<B@V7G%F,>XU*84N;L0'8*#97X#8+EH(G2VP2#
PE+]+D;62E37_IU[/R6%&??P(,)(:'8F$+0 ^Y:U2D6H'G]Y2VPV5\<=@#0-XNS^=
P#QNSB-DO[)"$ O:D""4:68,YG"+;5%*./,41IUR$^G@TO^%%$EGS6)$ 1G"N F1M
P4NM6GLP+Z[;8M&:QC_+L-L*&HM3BV<K/3%ULZG.%T[,G>M;31DCI;UHW&+3:(,3P
P81+FC49U^Y0&YE,?P" XZJR]:JM6_QT5+U$)J?L>K"_SN8C$J@<6:FL4]2P>^T7E
P[:@KI8\[&^O"&5<)80O 3'HST!#+[C!/4KBK@37"3"M:]C*1:8XE;K;KI("[)SL$
P<6Q2>^A#FJL1DYRN,D M(IH;?1<M1(?FU<E@=)QY&(=U"BE%6KE<IIN@-MH,$4(D
P=\T9,Q+-J*,,/K0&[2J>I\F69@#D"U#J,)XRV.R*U*L!SSAT3?-,<6QT(L4:'8,A
P9F^\VA@C60T&?.#*C+?ADU+A3#/],!IL.(VOS7V.*?B6EO:NT4Q'\Z"!<V=\?RI[
PS?9#%E]W \(3R57\6-NL36*SGW&'7\1P6RH9^JEYLA9\WGH7W=\@V<FK/A\%,<D9
P7F.J!;JM!?4),I[;=1&=/1"$C.0?)+YP1!-FG&0: 'U(9,30^5/2ZB7A"R,L(^,6
P[X6>]@*U(AV9B,'C"OY X63G[QTR7,,XO8BU<!.ON'9!L"MKJZP?:!9XS\8K]K90
PH?5L2)&P9Q6C5Q>FP[:>16$2V_60D(0DY6?'?/T$IJG(@\)RTOD5SA,6H<@B*VP=
P0ZGHC:I"@(A!'/"&463264,QF X:?@^& IPHS.DXR!X13=W$M"\$2-W*#*0ZH,; 
P,#Y),W.]T7"O4J/-4']A$, 4%-HL@G9I;*U@Z'@O93/#$:.?",?C9^"O&GXSA^FH
P1H^I8E"T<O5Q*I!0T8NVPLT,_6JBAW_Y^D0PI8&.AQ Z4!N5OBNAENT3;RL1,_"M
PSD%$B":E1,7OA+N]-CCD+0!%#OY)O)M 53C'5,%L)."L'A-DQHYYHS?7%'6%+@RA
P(PG&XRAM,34AE2GI^LDC2Q^3 LH,M3@V5M47:7*G0%5V1]<AX0@H2W,U""DH1"W[
P6=%W%=N#7L_U0>L7P#66H8VA:[:)A1&YF1%?U%#*@U28.5C48K=&/XY5VL1^'$9S
PXM43RY5<! >Q!PR.<=:4-A._X:B89K%8_DOS(()NV#;Q6X2'84ZG6@(X"G6+*O-D
P46E;<L4D]+D0XQQ4.9R3V5R<B0;G8NWP,G-T-KN;_F-EIVJST6G/,W6R0:;GB-3H
PA<3VW&.%WB[L;./GC0?D78W\!TDO6#0:M%QA3I[^^=-*EI@<,+<)9/"#]6T:'U8U
P\;.T4+7'/G)<-]7<"C?81]>."HF!0+\W_5",R).N<8)( ,WIG]Z/R,!J-2^QDQQ2
P7"[UXHB"[G\Y%M'HZ_<[IVNALC7B )S.GSKOYJB.LB-E9%IKH/_C5>1.E8&'9/TT
P7R;L=^F/C)WQ8T6Z&/L?+P>K5CJKZ\I3K;85A^\]W+@D3D$GTG1MS=8Y#*>>7H9K
P?O,2+YA-DE;9>@_8C>%,80:1*/9V@C)O9HU_0>S<K9[<[\."I #KH +]AO&'N!-[
PV@O>&=/@'&(\0F7E G710%TY[?$M-'^R7?&91]1K(?Z^T,<XLS^;YEYUF=YJL[>O
PO@Y>:*M@=J6AOS3]!W* B0/[ACA,C#CU/.4BC:?.A%,"TN<8M9]/!M3)OX[[0T#"
PN+L0K8!/;PRU$Q7U1H4EU&D2(95U,=,*+Y3V'\]8R6R_<?KGKLM<,H\,P74]9S]M
PB]0VZ  <W+/"J5>U;CRRLWH!X= 8#3;XO$3:BLFB8;2B8G]1$+V'B>RS1Z<L"E=/
PX;D33>V5ZB>)+:U@BI_0E3?#NW@G^)4L+V^#R>7?$^A&*/$CF7IX2W4RC;>1#VPA
P<34#<^M]!SO9:#:RK"CSAWZ-U#=L::M.7B[<UCY.;<$@6(V#T"70!\/BK'(U.$?Y
P^D]@&I;$K%20(,4XKY5J-/JK$O#_OX<(! NJ1O7*/B$^5%DMEDV>DW&&=O"3 SL'
P+=1DKN- /:OAA^? N7Q+3(&Z=:YX\*3_%5,C/7%-V;1W^)"#ETTW\>?CG'^Q325[
P&_LL]LTNX9OHT=[(JLW4A Y.BB^AC$6/9E=6TJI8' ZP3I1?X#?L2]IY=GBJS'AS
P3?J$T7MRV7BT_*_TFX7K(XYR(VI&?!'.5B%ZUW-ULG <?R;!/B1'B##\E^B[#^F\
P#I9^.M+/@MLTF,OXU2F:Z?G9W</9$&7J*^2'_<")+%^L:WS;T.>]#?[-[Y2E65[C
PQ]9\P6E7;(UL&;C@#T-T=]@?*<*3(-(N[_$A0@>HV=C>H52]*S->CBW-*I.K./9O
P:E2LG/-+WSJ;A%DHVRZL#(@1S:/YL),V5\49M5@<+Y06B((V%=-%:,8F\!NV[0D<
PYWZ]6BM/=+,-:K%5TC(A,N]65')GMK#N$S4HWKPGVO!SR5PK'$GLWI=I2::5B(:%
P?YC4\3=V!XNA']0(!5]G@HJ"C"X\H,\DL:6<.\IT6Q\Z2,8D5\+\O \)]K1BZY;K
P;.^7.X)L)SZUWLN+@$NT$.?'5*S(AMKB*WVGDSY=JL;Q+G%86">USPGC7$ 7:"@'
P;5V;[BX[4( [;/5;Y1%;2.W:CG<=/=A9D<X-5I7TG2R14ESJ;;3S3H;VD)#XK=X 
P(C]]T!RB];QT^CV4/JQ=$QU\LU(=&[[_>KR189P6/S;L'@1.1QE*Y=8J2;[NE!UG
P*:>"-\1,6^.JY%4,^K3L]IY2(60EH%0'R!^</LV"(O3%4(]*<X$6%M^F3($"*7;4
P><[LT48[[0VO9)B(SZ!-1K3*"'4M&H*S^(?6O'(C$6"8O:N@Q<\HU'N5,2-H8Z'D
PIG)!*IY3"DO_"M3H _<4C3J5<(]<NOBC0QC(A)C3L(8S!/9\AT')6C2G$9*L!-A,
P+4!N@D(QMN%3+T'2R-QHY;75>\;_Z81%CCXUQZ>B#FICK4XI0,RP8-=!AKJD6[DO
PCT24QJ'7.K.V WJHHW H\YVB/3Q0:BB4PAZK@/>@64J*-ZU#$Y.ZX;]+A&MCV*+4
P&VDJQC/'F/'+;O<X&Q8O;\YM# \]L5]V>F$B,2J=WTHR?('?N_</<,W,6OD(^%)B
PY(R%K25F%V%G\[WR?[S)L/#91W/QH"QT+=8"PUSPMBQX1!ZL%A/D,C 1JR:HIK7X
P;EU5'PN#/F#5TU"]HV-IT<B;*C&_@UK891G]$,P,(U_[-],'BY?Q-1,%9=+'<:RG
PWJ;"5K*(0$BNU#FL*\KAH!;,1.G+V.=F7=:ZH[):457'I3(VMC5\U#ARX>\Q.>[H
P71PYYC=PTSO6,Y_,.55:0I_;6W&Z4K0[T76-%./4#!.-EP+3_*^7YS$LG_&IA[4-
P1W)&F4<CA'4(3:-K.B)@J\5?<O1N36AG^MGCEV%EF%6C=]$WF'X\"-P_E^F:O!=V
P1F(R0&B5$ ]G=AE5/G?&",:&D@C?/*M!+HP<?9/=N(S<>^C.(H5$%9 ?%X?M$8\4
PLF/28\%SWGP6O[>+695,;JZ_A1\@VCQ2;<H+S#X55Z7XY)DV+C6 \_1[KO3WG@V(
P*%,RP<J7V"F M/IP!_MBM.'9$6??+['P!DK8F VET_OK*[0&67F6T-VRB[YI2[&B
PM8U+9\][>O66>-ZI[>%OMPI41?'XR["/;D2 "/T;<6ETXI"VY695<S9LGMJ69BDZ
PB?:-3:/^BY+)8/M8OMX\=,_=@U0]KN;L19F4%'<1M5^E:!7#J]I+:RB:DE-SFNL*
P+S]0[S1SO2WHE#7H#J.0=<I]/.5E@ C:V0#@GBF!?Y%2S42ZLAUOV:U"_3\8"4<Z
P!T@Y8O P;%B-OM#'%P]!LJ DITB\2A5UGV\H)=ER.B>QXOD5NVI?RKZZB5D&YK^U
P0YQRPC[' LB]T4] [A4^)SCP>I6<.$C_G^.A+R/'BV9HC:NVRQN!7O4OX%'X<#R-
P1VFD<+PM,.6K_NVA-P>"M2H7Z."-D0(O)QZC'AK3 [[7!2BBA'+$>1<5KTB>_ Q4
P3]=68K8>GP,E(A'6.<G&MYXS^N7B,PW^N_,%G_UV@^#?G1)Y*&!"M?83GN?YGLT=
PS+?AWJ^6\,8(R3\/E((42X^Y.U$5:^/5Q*9,WP<'24VNX%=O]TD"$>0^?.9W<26.
P  N XJ68.4,N)!H>^V$I1RF#Q%R7XI'-I6(,%QDA;09*N8"N5VG=WZVZ<'",:V"*
P#<=QVX"FV+41!9#AWC\]#K;\MHA-TUJ)(FJC)%_8C<T\X5OT UN+]=D01MD#:"HN
P.3/%CQ0(YX1+(?/+]J2D8?:6??H#4H,;U<CRI\U])7*0Y<HU0EX7.X*E%*'X":SO
P/-A,0""''C&_!WN 'NR#B!TPW1BR6LF^IQ IV M"/UBU&Q72M?R*P;2'%O'>3&H0
P%:F/6Y' )6!25V,1'Y4S7/1JR<VQ:^U?5A$JL/&<FE<=*MNSS26N ,\U)2W-I2K3
P;6_RB4O)I3$R+U)+SS)S+/0T]0K:E&% <LG[SGXE;-K33=!1)$L6M?.+>IZ.OO2-
P#76OUC646EF;(T@GKY04W16A::@>7T!(K//I,)<#L<N(Y/;F>(BE?@"T($"W!P!@
P" _K_^R)^>+#T8'2;D*$IZ)#20E ^.GA**Z8.'@D*X5H= #UO@[\;SCB5CBAVM1J
PJNN^+YJPSMH?*R\>9[+Z68M6.P8(KW^#T[3@V6*1A.;\J )T6L A#%L1<W 23RJ*
P7Y9^+;'X-)V"C_,1E U7$B,K:Z+,F0#F1!9BSX[_&,I#!!9_3@O?0:C>89[U$L 1
PQSNJE,,Y7O<?0_[U L((>1T1G9^-(/YM2''Q>A\76A,%(OA](RFH#ZN2WX^1F[Q.
PH@@FN*(:0-?_%Y0/R'<@4QX?(U[$."H6/Q[%Y'$R02G--5V1,!3?-VIJZ3BSQQOQ
P-U__"8RC7/?FUZ-O$ZH=$=YT"[=<+Y9K*C$*]6UFSZ3%H;J8"3&@  .-K-QXD#.[
PHC0]**;0;B])'!DD=$A/0$$<"V_?H3MI=)C;/\O$*=",=W>,-H<'Q5QY/Q%8&7PA
P_&>O0^S2/D*C^!U;&@(4Q\ 1,?P+PMH'$AT$WP[2KO]1+Z'SMOS)HB)G&EA=?1\P
PL2O?$KY=E;6>*G4?\$6N%W"$:C?FI&33]PXFR.\(A\G!F]^E"?C^PC]EB$.O^DUD
PD6I?RWO)/SN.\^]B4W$E,<:*<!57?&:5[^5Z)<1Z/@9"SJ=%J\3[>D1"0%",VG(\
PIV[$G$WB_3;1_X1NV-?O/>"XGV+S.MD *]EQ>7^M*VKXH4+UF 49LP8Q*_S0E\%W
P6 O8VH@$<,J6W3O$J(,_0D^&@D9Z53CX!W2=+@: _LQ\76#].G^PC-]6ZX<:5IK/
P@TULKQT!;*SI@("=J3.78JO!.^=C3C-Y"H",($+]OEF$5;AYR!92N[G*-"FT >QM
P^YX\]QW7$*/ @VYV%C$_D)M^[00$VD=$^#[,^YR^T%"9XO1=$1B2L]I9!"&$:2?*
P-D$\-M9 %!*??%EJN.LEL"GFL&M'>5B**P)1)42'+)A4M0'Q/F3,J6Q+CIR5TT0[
P\,W8>_-=K'J>R=N*2$58@0T.HFG5>S"\1;> 'EH<K2^* TYN5+IU?E#<WB!\I%:5
PFFSK,^4-F91YZ9X-O/:;CRP#O:5'*L3=WC4!O=]?^Q<; 4@U)W#X1IN#'[UIWGY=
PWN%4M%<O8;P$V<RPBO#6"8))?<GI$CQ!,G?.L]#":%XP%/+GU8L.4B <JCL\89UL
P._BWB9]NI*I"6.!ZX>=D/AED%T'O$888K3TE]%2CTY.7!]+AO/(LGVT$S^THX$_C
P*?C1,8<6/HS%\LYL![]+*6M-)_YLI,%SZ+"2,DUF(D++_E!K?@/PC7V@TNJ,K@:A
PC05A)=,UE-\4)P2;TTQ8X;MOZ8<P-T&G-(+%8^$/((O?IH,[(*T_''XT$"3D03T:
PPEP >B>XSM\%.2*Q-FR _+T+6.;HVZ+C-6BQ+<PZ&XC%5!A=C@<ZFDT*=%00D,PI
PIEUH46 VIB3U>IR8 XKX<'')S.+O9,0^O-'?3W4O#N4N-BD]>S<[PXH:XBF.U%S+
P9NE65%M562GEZ]FC$YG4N+ SN.N#!"@C&$$ MA1F)*XJ[O10(5.*KC\@#Y<GON74
PRE#DI?%9TCG?02?,@7]O9]KUSUM09;55UIB?]!0JO30&34GW,4$^Z 1/JQ!F<B4_
P ("BA*NHL=&RM0-_ )Q<3@SQ /@6I7%"H%9RK'H%7U<IU"5XDL5S5+DD*Z,G]X%Y
P;?B"%-[G8+9K:UCG'0Y"X&:-,]DYIQ2F)ZW/%O!GA6^/R596PX+A9E?!)LM4'EN!
P*/D,L;G2^RL?#W@GJBR@%*\87M43ST?'..0B(;&V/PF+=;4[AZT?I^$H/AHSJ.K*
P3#*U(O?J"2%H+U*SRG[Z$@J3@H6::<PBP=GQ5Q[M)-MZ(RVFXE8IVJL<)9RB)<!T
P@"1,-U1(9VWB=OD4$+1;2GUTWS:'1S B_/%NNO)?=VKV1]/:C3  2VR4H=3H&43H
PK5&:5S6)!=^/X5?K)M#DE!4O5@O09=XNA-T?RTX2:'5):@U<#ZONJH>I2S1K.7C-
PM&NH%N2B$>H2JF%GVF)S6+/2:I'K3H%%;,(V!6H3$@_QZ-M44!W8S=!SSL;D_'+'
P "U4O6FT'PX)0:SKPF(5S&%WV.S83?.-6J$,HIJ>20"TGM\28FS3R4)/:&]N"SR8
P'K>=W6XS;67HU68*J/ ![L#0'UZ^\PULRK309C4O70#!1>U;I?$VH4DNGLE)M5L4
P<:3L-;K/VBS@Y8"5J"KTPER%X\LD0[A1#=)&, 7ILRL-4MV#KN$F?#1(A;IH8F"H
PH;5M/#*,5 WE91O=PG\7DSX8)->A%)*!65]8)<4B!MB3Y,!'K=#_XX7=(G<X H U
P#MHG7__,5I0&3/ TX,-'/=.(D<;RH(U(A#)S7/UTDAZK=Y,01/A2 ;;M27QGT,]N
P49 O!!"2XI\_*^J3-<9 7AGGZ((K5AV-3\0?36]8,O&4F(,G/.1#4E;; I8--#()
PID\.4WF_[B &U(CTW!W\B;)8G4!3\&>'UJGLLJ]PS_628Y2IO'%C"HW">$/^D4MC
PEECZWD/.T>3K6)P]GN^TR-\UCI_V"I[H=2@\:+?9HFA'$85_4R4Z 2),?>IX7]JU
P\[NJ%WTA)4Q-UH]>$F=V=.5 YQ8(P_*:2*/V." 6+S[V:G"A*#,%'N.W2E[FRQL4
PTBAE,"ADN(/U^[PH(>,X_Q;(B)8 4W%OTBQ+E\E(T*Z2WVRD. F^[@9V9%YH16,@
PQPV L6N(&L9LC4+J5N&ZH5P@H#E)><]P[@WD*%CI#=^#8<<^]39Q.0(-Z9=1DSX[
PWN$6/+/99@B_ _R@X(\W(ESJI1IA(BU P(,Q1/"DME?#QIQ37$%84:)/M/,T\QP4
P<XVFY9N;Q7+DCN^0U0M\%1<]0Q6/E,-O)Z,NR&5;;#UEQ$>KRQLK!N5-,-A)2W98
P[$EAYP:5>H(\1-, (#(KW!8.U0YDW N(WYI8OX]5%GFB I@*U-->Y$_0(9T,4YK'
P<9XBV,(SS9(T13\%4-^2^@VEL:UM[0W@@?\KF".@JKEC2>6P +K%<NT>)1JS,RM2
P_5+.C+T2#,/9%X_L=,28J5H>G,S^G@[B;TRLW;,&Y,--WT7<R-F_4VG^\W)\L=&W
PM;1,[W+!&/>H79U4+GWG4JEAM$) L9!53,%/689NGKT]Y63UZ7&\)1P5]SNT$7WI
PF#40%PGJS/ESBGUU#=3DN'(5[^+C@)W![H)SH>3QI%QD*&IDNPQS?!F>)K+*2O'O
POHR9, 54Z,!J#,;BG&0:^U(P]//:(*(TU*J*.BD%C6,W^?2R&5Z)L01&J\I;9NS>
P<8:6ZP\JL^6;LFT:53O-(5:-<Y5A1&US6!XEM(\2"6'),=:\G\9K[GL4#EQR'YS+
PNCBM)?-%"E @0-Y!PV,&D!\?5#T:"ODU=R4W#*'N@3[$XN@\,*W:%]]-WD!\/J=?
P@O(<G +DZI1W9Q\XIRCOKB=!NIBB)CGS1@UV/\9%WL"VQP_+B6SY^A9^2JK'/C:M
PT'!E2KL5SKH.RV"]P4?^9H(H=7+P0$B]42MO"4%,=.E[L)5Z*S,N;)_X<$];MF?U
PO7*4JQ-@M=YWDDFD[5LBV.R$YJ*W-LI _*PV<V,(9@?FF<USRJ]WV]2[P023-8I"
P%M%9[OMP4;P<:'+?S+Z!Q,89,Y'+)MH*/J.,[G<_^Q4&<C%PX!^]_/?W=%X\YX\,
P?ID+A#16\=UNU&J75+4LI0W6;RA622>&&"EZ:.5 TXH-_&]5Y8%4M&;6BDL9V? 1
P')!=8ETX"OLF/7Z05=*,FU(P1?I!Q\F-G2&!TJW&/XO/-JU6E+7Z(<5H:[RX5?]V
P_ $_768G?9"3S0M@1_'.(-$C<O)O)E1C9,A7*:-&XW8//H!EL-*^1>T6 ^35YDR3
PB++\ZFD^$R0RJ&@-FGXF&MH!U(U_OB92S3V-Y 4Y7U$H+%L-O<&.N* _1F1ZF!S3
P$F;([N:.@^8>"SIBH.L=QK'0?$S?8Q>1>$O .:[O#@NSE *"/5Q,[*R'X@*:FDO\
PJ';,FJ')^4+ZG/A"-Y%]GR#]2\T>"=0MTL?"(Y-_M9MV4%>-G2]_QGV.*H4]7,H<
P$'4E<F:?B!QR\EA.7O"^(H3::NZ_4?;PXMAH(NIZ+O:N02_^NK)8O%X;T)!INIY9
PYRCC5AJZRC*?M4R],.%WM4=_+ILP8-;0*^YLCU3O /6O=Y6))Z+ ^G''JLS/!S08
P_P@G1EW/8P[3KYPE\Y/8FF>U?]/9V)NKH%Y[9L;'09-L)KUK'LXF, *B#BS/48>J
P;2!TU%/F3%)$R3M,^#OY^PU>!14^M1++)7<X*"'G48VH[Y-F# G]ZR\$B>^U;IV!
P,$#/$7=6#HQH8.TC0PIJESM>LXPC=>&G.BX-M^V&M^AWC@QJAE*P<K-FT)A._,3O
PN""4P';^G*Z-PF!7EA/9\XB_?'INH!6=% $,,<O6 W4(S)E=P-%U$#>L_O71.D,'
PBY2Y,\+?^>KH] 4GQX)(TK[(XZ;?D3AGZ]=$?$S14"AS6D?F^DM<!J!HN58\2NO@
PZJ(0+I-.S=6\#HDD99M_.-=;",L8$ZE!Y-,-5BD%<=UL@&0Q.H<JM?IQ8[T)XJBG
P#,WD)[B3D,\AC7D>F1QF$@BHU5]W+H\V5W>6L?ZA*\3><B# &;$42$TE1LV5%FSR
PP]T)O5[)3T6 '$C4L* A"?4;5NXM+%97@+>#KJ_2C0A*@N^WA$$@$%)81::<6[ \
P)TAW1-6UGEW($(H8*GB&O!G5NFM8]#((07(R)D+WU07'#XL_?9V@,;?'&4!'0YQ%
P2CV,%L&6']/6E1Y6/1B#1!).,+?0,H4\N$ ^:W(\6S:<@35/7E%T@&;#RW]DXX+Q
PL\XN\K*1=[6T)C0:-_KQ*UE1\<(QY?R$%=7\VP^&Z&]9I%?0,)]/<YF!*9SV'7O"
P,<UA=LE%@-9,IJ4TFRO\\H$6#0$AT%MC!/74U# B>+OLA/'G-QLPL+/)$>)A98T*
PBMRS_?'T4C$)3>Y2*[ 1XR+7 'I-EMO=64'!37,!] P=55M?S''O>!&1G$;>/1XW
PS7O4!I,?-\2@ 0/ 92KO'1^M9+:1&3/#(C[KLJ-DQ@4(??PN4+W@>&;*'T0WOH26
P$QW'KCZ$#M,'A"Y+R[ZL=B7>O$AJ[O.0JY;F+60X1O_0!8<P-DF['D$U&U:E;(I>
P8/N?'(/4!\\VKDF7[VT;ZZK3^Y&1T:806.]2]PTCR\^8'])E/<"=="2OX"'YL=5Z
PX6PRO4 BKZ3E64FZ+M!&*E:0T2+&E;-TO$-/YPU) HZTQN;T]>N3$"WLY:+*$5(S
PU(>]+J.<TK0H_)7%RU'.?,X A2OV9P'GS-=]7WA?\\^EB&HW^Z&C!*X;!-S6U+8 
P\5RRGK%C#$6ZG\/-?T2@7Y(9EFHK?^';!IR"@0GS#F$_H<05N*UT[6XGBD4D(KX<
P_%^<V "$.TOF4_0NLY'V1=\T]_I!/[XFUE>PJPEN>\]Y<$D_2@]YV1RPC;3.C%".
PZVSNS+?9P?95!UU!;5QXVS$:?LF@).&4^7D-#U"V+>:S0""%%"FD\>'/YBF6<-%J
P1SE.^M<45";*>Q.177M,NP@P,[0JMMIJAU3"FN%$F"8Q OVG;IT4C?O@%BV1T25:
P0F$/Z H.D':5D$/_\;".N417" =OZ6^9@\51@;T1^3U.>:/73M&.32\L)%#.2WB1
PI?42LT+>SQ<,]8>%VTP#?JMAW;T^6LV2"H(IVK(;.'W_<S3(P7>"*0%0VL\)1"S 
P>"^,VY-<4F163ZN\;6Z@D-OF&+4"2+&-2O 9_FF]+[?L30)Y)3YE#C'Y]/8^@)5\
PS&P76YD-(Z? LJ:\N.A&NVR=R3PKZ9%/'&I[I@&?4IKIH+(B1):;Q;>,62@0NMER
PTZWO_ ?EL(F-9N&J_SF88#G,-*&8WDOK+$)4F!",BX+#O)%VS#?8X5%V,_O.,EQ)
PW&1$ M%H(MU!G \;DT9=OQ*72?GEX\8S!02HE@A@%NWD95HQ"Z$AG>-?6=RU\"U]
P_FW_6L;][7#K^MGZ>>8UJV';71FGH@!'B3V1&OL?*]C@29]85-BCH,3)VIK(TSU4
P#_2#36SZ97EQO8"B>NL2='I+CZ:=+\Q+<-1@GS?"^)8YP1 *[RS^?D0.+J[W\>4K
PEH/K.]W*9?"5T;$()X)0L<PG1G*26C;P#,$R\(96.O&N>>&]I%M^=R6^-LJ^.DD:
P4Y*C(KDI7/:Q"7D -.8.2BEV<\;#K>%_7A5%BK7TMAE6T//<;@'UTO<N 6563L_.
P=DIP S:]WTQSP6#K$\8'1446>K$M<PAN_4;*QR^I ?MIA0)1%K?K8+^ID8(]#SN7
PRJ1\H4KI''\LTK,>"5?[8"G5.HG&[N^?VJ":+3!-TGSK%!P?(W!Y'("+ZTIA^6ET
PJ3QE%Y-K2K$QTQD52!>!QP=L[LZ2H%&ZGS/>3E5H.%:&]_S)52S$=5R]I)2#06A 
PZE0Z#H["+X?B:Z)Q+*,O?NMSJ;%N!ACZ/IL<UC!%!)\:C*'?&%:%EF/^_U#B1Y,)
P#P#D:XEJZB&%IV.XCXV-T[M9J-4]&_Y6,PI(G45ZY/TO3]ND.:9W-#,1DD41/PLI
PO=OB[B=["/G *',QI)>$E<!UZ0HLXV*NL("-"6A+WP$LUTW$:F2Y-18)T^W()XV8
P.6,R09R16M<CD!3Q)+?7JZ"@7O'&4JIZ%UKBMF4NCNLES/[.%QKH30 TOWTV:M3G
P=JH*<2O+_3V@T7:AXG_RYDH?H_ ZNG7QG&+')^W(Z,E)\YR-!<>TZ?]>?8$7";D&
P4;HF$S%=(&]:0)/(]HC(L.>(PK#(G9I:7RIC#;8 2&5G2,BIXP .],C($DHGCE_"
PQG."-$%JNJ.:-B,4S1(T]O<KYD!N-EE@@2NRYL6"H%#:=\R=:#RF@>D?&_Y*K@V?
P3BDVQVPDZW(Y/=VV9E6FR3<6-?+;F"6[IRC/=3I.,M\+\<A/:(%GPJLHEX>O%6<B
P?>LJQ87OACJH5YVIXMS],=_='7AW_9T@EHILY[OPG1W >=GJ%C0F@V)3NFUC &2G
PE(=7GCY9D8DJUI ; W_66XQO$NM)QF^!,C-M&W=6)3#4D!YEI(#%$P)CK;U 2'S-
PV)WUZ@#A@G4I.0U1U'>6*,H0_[;]C["3TLT2(D<66P8$3I_KJK9&%73?']@T)PF1
P63;3M^3M'7UD:C30HGJKNJ.P]1RP6>,A:(G-'G98>:&93=(_ "@@88VTZA0: B@^
PH^^H"Y*"PTS>@TW@1IK>E1=5PCACS=C)OHLL(HA>H[9)OMEKO3V5FZ!@=6D9M%EP
P8G.S\2IBVHO;P[I5A)44N[& MTFF(LZ[BT#G+870T!5AY=\GE&/)D=<K\-:KW7S;
PY2->69_;^]D)<233S5 /X:,*^$78NK@I$,T%7<RV3A3RWU8,[#9?= V=KT=*^%6W
PI4$_'KVSW,T6S6 @_'W/$"S>NS+3A*J19;8?EOCI?H':C*&?5V!T8S##S*';U  M
PMGWJ'Q=K/YD=8)]<:-TB3VG<"T=[RW,SHH&7EXF6Y(IS>OR]Z^;ZB5 9?;5S-PN6
PP1S[!0B\8JE)26\]C"4_ ^I9N8^C4^/'+9$XM&%N@ZK;[A-;ZTVQGEK79 E$Q"!#
P#-2FW7B+770A5/IG&CXLYCHD*N=J1=O:UF)_4/'VW66<;T:*KWL[MER1T*4%H#8/
P1T=FRHME,5WKCU D\Q+DQ'OF8D%RL>+>$.?FU52 Q(YE(ZM320KZO:#NJ,*'S2QD
P3 57P?@6 +(BF.($!<,O0D(;"=CVAA(P"XD[V;.80)"OQ?ZQVL:FY:'F(:4G^V7C
P&$'KOM/;M#=,GXN"F<$P+QT'/5@2 \O'.BV 6/6,$V3[!67>:&C)N2=H^<$*S).1
PI38\;I>56/!^.,6%PWQH_R:+PN5Z"C? A/O PG).MOCCI_M'$R16)[^=V&S2>U2[
P3[[:^>H'^86B&Y^;9G$TK-4<8L&S'=P]^('ZOXG$&VXG9&^9!AL1A%/:30-3Z$DL
PU2)7XSO_5M&Q)6);3FR'':&8Z5/(PT-C2^._TW+:'><>>6'L_.^NP@R=YJ:S*L^#
PH+JS0,U*SK1AAQFW]ZU,^H.YO)Q2^2AG@ -E$\!Y25+&*(C*DDKM4-%0!L#9&2SN
P86%_B'%[QM9RH9GK$W&%DM@:Q*@BV$([H%M(U\.WCQ)(F(G)/8VR(HOR 7LX!4\W
P-3TX<5VET:/B=^NJ(32/QRGJ HZW&T<UP?K*GR3F>+A><GF-_Z@<:"$2:L%;/=PM
P<])/]?00*:6VGNX(J85;E69P5/EZB_]4M0N1.L7H&")^.K2.?*/WDK(^5-KM.=HH
POSLGB"I.5)4?!<JA_HV0%[[UYFWJ,[9WQ])P_/ \,X?X0)?E\%8:1A?U>\;U5ZL=
P%!J</.\+!41[DD$=_O%9H< ,%]62,:X=1@J6$+RM3)ZMLMF=I5*X_:6TEI4)&/[O
P3D4+3X8:O[VBN(V#$EW9@]_K_"0#5!K'+E#M=B--"4FH :XAD1$U;*G[</^Q&09R
P_I0EEDZG7**=-X>+OT0]\QR:P@G]B789AT46]:>R3TOE3S\53K1EBGK#U)([0TA'
P.F<A[8X'B*LCJ!3MD&6";T[#=Y_W8G8:'P)?'<+*\L.39>^'B4YOESKU,TU);F++
PQ+[%231?[\L69![F_H8(Y?,ZJBW4Q"-!91UT\UFSG1M,8'2':_;W;,9OPYG[ 4LQ
P!$WFEMS@3<)60D[)*Z- 0/Y+<$8:LPI1\+FY+Z2G(+]0;2W=P^TKBW\9L*_@W1#O
P9_D#:KX,4Q>L;V(T$"(1^_N,EK*' 1[T%^]X?Y."(!#;^\^3;+&'&=,99?+&U)T?
PR_!K6;2O-5U> \?"">_-+G&(^%.W>U2R;R?:0\C_DH1?\H. PWX>47&&^YOF(XAS
PD 3'-[@3/J<?6MC(^^0YE".47?CC?4\11%$>5E[M4B= 6Z-+7 R!_8O%?%#Z2M[0
P<05>([I#7_A3T$8> ]?"X1:UZA&A8;),%J>]/O\-_SP[J-V6QKXXX.!!,9/,W&5H
P&;'?*6]R/I?!R15^(F:+QXC!JHZ.KVZ@E5JU9E;!1J$^W-ZSG:T5W0%^<#'C#]"B
PV[NAED&K021+5@<'YPB:OM+H74C%MXY!S>@B&/(N495/D/BR)?F.?$Y-K4QV-B\P
P?4 >\'L'@MX%TGQ8_UAMG5V,4$ZNY8.)%YG.3D>"[S#D;%VH2_NK.FT'ES&JN+/1
P"/5JBY]Y-$B+UJ8R5NK"\O#3D<H&687Y-1<! !8\B>'[&-R\=.*A4$J]?E6&6@;$
P+G)=2"*0)II9(RZIK4]Q./G-[,-G-7J?]S"\;+I9OF20/S!<\LYLVE%VK#LQO2RM
PR.>(?2J4+<7F?V1=]"$NCB&BR"QR#%=)1K*N$*/*ODM$(G2Q1T-5=*E3$=7,S,G0
PC+-8>QO!_$)U))6*_6=!)[;V?H#VR'[WV-U#L+(13I(A(MR2<OE,>23Z,(K[SC9R
P&PW^K(+A]B39QT4P"8<3EW0&]HF.P8CIC2TS=ZR"4%IAB5,OZ *8"&789^QFK2H!
P0MG$Y]Q8(*3ETR]U0KU7^B^OFK^@/WF(9RU.+PHHK1 O]?CJC8[>0SKO_4^0PP;!
P-EGAI[O@&LG*['^/K=EM&8/FUM<WA+TC-WL;:]IAU?7!UF^5*E1-; !9)_-RWKL,
PSWMMBA0,S >:*BDTN4LM+BV]VZ]D=0C^O>#IIH1Q?RP=#&G^ZMOP0:_.<MYV*>8J
P:1F;BQ;U1;L$UJC(&5&2%NB-R \ORWU+K\"-"*L(/H1X'F0< .Q )D"&M)+ZCQ70
P9K*L$O;0%;XM5].2D+?]P;,>$[HKB '3,:#E%.J&&:?:';ZK1'RSJLW,[P';Z*T=
P:)6*DF3HL5WR'ND70AM>N3]=H/0S*\EL4GZX$$.;P]7F:?QLP#_MB?J@M3&O0FX8
PCY ,_[N*3&UI1YMGQ#0WTT;)WU:M19EZ,^O;/+ZBY2D&?".5#NC!>LA!4:3)'-M/
PAKO^DHRNL$[&:* S<SBO/UZ3.+1$CO&?=@*]VNHV^S%TJ-S&##F_--Y\VX%#!G:6
P7]%P;FV$KB(6Q%_T?/$D+[DTU&'5:($@+5_XLF1:XR06[ FE<IU?3<C=6/\I7O&?
P(;=Y,2KQ91\N!:-B!(AWZ&Z631N6H"$8UZ -UTP4F#KEJBN:/X/E,!NWGH_^'!<(
P!:S+$I0;E>*=ITZ4*#0Z2@?GJ3\MO&S?@L2#(C3(F^L"W,2-L^?N$O>+H34N+46V
PC[$7_JELL+FEZ^AT5D?.F.+<":.V@V6/KGT__J[W,#(?.3 U=C6+K+GI<(7])@C*
P]-#ASTX_WV4Y%/U$[DMI:_K'QJ5\I,JPR(1]D1M3!F"=;^\$V8 *4&F28WLB.+O&
PWF 2J1H+K0%/95T:J@OH*[EGL;)>]#/YCX;1><S/G.]%2V0T<$9;,)UM)(>SS.P@
P>M")3D/; ?\ T:PI&\7HZ^Q@/8\363-JQ)<RS&2EDCW:KD;HB2QEN4[W=BX::O06
P@V:-M_\C$PA+KD\HF$MLV2JA-F5J)O; $+&MN?FC7GP[,YXL?[E^VUG4;7TR8!)T
PA_@%;$L=[;&Q^&F0U; EXD9I<KR(NL%**9@&Z<@>G')RQB]84 H,PA%]"'G'K75]
P4:*3</SFAR(?=ZV"*@[K8,8-.YX6O46<K]#"SW K$(@!EH[DYPM6?!;:6FQOEIM>
P1"V&>@?E;K9P''6FL9:A_<F^B)@4?8\3A FQ]GH%13V:B,51VE>N[$0M04[B;[;K
P>$<+G"#@X%>V O13]^Q&JCU3O7]E89_(].OLWOB)S0-+.*__&]1DC-R]A7VNP?D=
P,W!+GO!-'2 9]FF<(QQ5;Z LQI=>4C1IU*GO5588S#YM.ANRR3C-E?,PU< L?#2&
PS<'4@?1M:ZRL3"BW/8=G@_P5\0RV3/42FF0=?HRG(MLEM!8*49C3>'ZR.\BED5^2
PB>6LR4L1#W=&<?8.#H8R@9Q^^2ER+2&1?J+!S4=%>PJ;"2XF^3V. (C[[2O/#4QY
P[U>#L)6']3-4%:PVIS*8C3D(/(+^E_D$)=1)4MC!EM,T@]1"1^=IQ.S@!=$^,%?0
PM-EVTQ8K0XM-:RR&:FSV)Q&\?S2)]K\>M*^4]I9U!!.Z2-Y2EY,L$K20"IE3PLUV
PAF< Z2*NCZ[52A6F'/1_ZI<07D(TXAY3Z^$R[]'#N'7OZG*2;C+3I04T8C]^,%?2
P 3YS'&_[K\!AA[@8"/'05&52?^LB\MAE"QUUZ/+UEF/VSOF=>=*[L /?[1M[%E8^
PIWQ@AJT]=QC'QZ["T1;R-Q&)?UYDRAOD???FNGK>Q-6!]]HE!PH V?:T'3<,\D9K
P"UY2IJ&M)72P5NHV,V9)/2]EXM:G,9)/^T%('WLHJYU14$#I7ML4R:4%X5I8R^?Z
P (GKA4>_(1A4#23OCH-G&(YOL]6Z+SG&JR%L%6+;TJO27[!Y03F-"(*4A\.8-'5P
P(*_,)DC^9&_O"FET%O,]M;\VN:\GYS;Z>WFJUIF-'C0DRL5@Z2VF'*KQC\?X(-'I
P(W3]B7TP+#G5U^<<>NH)&RFB?X4Y]NR.I6TO\RU%W\(N+KER,K<IJEHFL;],@K=*
PTVH %Q:5,^R;6B#A;E?FI_:SP7E8<$# O;,7&0_V]X,)J##.&ZJQS.I-&CR#PK-8
P*&@7!"#NND#5QQ(SQ:4[9ZT5#%; .(N\1MVCE%&I_CS#V=BF?#.LGPT]>([5*:&N
P,MX?BXS!:DQ2G;%D(8J+2K=[]<1'K5SJ&$2=RC>>:,IC;LFO2)@'%AS)C]VL7Y>0
P<!!;X[IOAN!E!17 =!(#UL=?+(;2AQ<!S>Z:2DICPBO7F7"/C/.6F0[[>JH?/&,$
P*#L5F4?""']H3H,RA 23X">;H3IJ I$+_L0%GCT2R"(C49>4&G5,7JQ]-UA:V*)B
P3SN" I-Y7#A<QD>]QT?EPWJ#0PFLI7B3)^L9<N>L=.&U=E,&L>';LQ^S!P+[@E4>
P_F-<"D1:FU.\E*5=LQDYIW8](2AW %S+. L_I *A;8Q:MC"Q'-897X[[FT<X&F]M
PLOI26ETD+4]ZC_:B#K/,*:[C"[Z(AWG(QRI"L_>:IO :C7_Q RE<-$*>WS/TS@KS
P605]5TT-*<<]0VH4X+2\@5+VOEY)<7VPW!JQ,9X@IU);BY@(D,?(GN8V//"KC%N>
P"FR=RH5)D\:.>D?*@:3*[:3\SM"N>2D_*/7J4XC1\72*%8;TJX4_F&+UB7WA[QMG
PZ"1+NJXJ;4+FC=FQ5Y^IMF0(647/<09P@4$# BH5SJ'2HMHCEDT=J_.+-IH&7WTG
P?.X7\S(2KKSEVQC8?KZL/ST&Z(&H38$ _(PZ(3WW)-:WD&>.8=L%@))(K1&Z$F]P
PN10=O;07#NDU180-\=0\QG3G=>)W8D'2!\#,A?T0:=P;7]C:CDT(KQYX6B=AVY\1
P'"GW6;(6:-UH5X4<2=<8"YDSW&#M^X&_01C?M[=,?X7?[R]:TL9.[X/[#0WO.%R+
PE(I<U[?U_,I@0DAUA\7@R2.-$)O-0>/1_DRML?>7G%LIOS)XK984_V]E6%S$39\]
P4"FF]_JL5*K^\Q=!8/(0(@ K(YR0(B<]TM.VS'2W#2K&Y=_%;VDR1H=/:$KFG/:M
PM9D_'90'ZCA;1[Y;.>R%BE.#&^O;=@1C*5NKYUDZ<!X%<=;RL\$:)87?@%,N_(_S
P>6*.+Q)#PJ[MC<C"T"URZA2(<BUT+C3EP*%I9BR?C)&U(S< #!:0*6GC6(\.N"$<
P;MKQ/?:=+OPI[J6)&Q97U^6;^$\--GH%@DD#<B/!>D*4U9WBAZ4]!0A.R2SQ 3M;
P<D7@2$P%TYZ'0=LS/G:<OK5OV'689:\<!8A>\M26]+$5_!40!&0+RHY[4(PSM[/=
P:MZ**Y?1"@E?M1V']LO^20V'CLU5H65.:UU4L3(3'=\TYPSZX=V0S/6,J[Y58<VR
P=SF*;=CVSO?L>7HF2?/(FOEQ(00&:.N8 EC-2*<[^*MZG^BR8W];K-$P<"V\Z&+U
PO'!D%I,9SS<C4*$&LY=:-W,+U$=CQ=^)=Z:M>$@#,@?9,*7G(EMW]@&;;>A;=\\3
PS[N(-7@UE,+:AR &V'W5XT&]PK<2(I6-3SNU<"X6CM-^GU5O)P0I!QTGN/7XZ7/.
PURR,N *AD(7BGO,)#0F^F/S+07M)B+;_(U#H<?A7.@FC&08.J8W8.:=3!=%.JM53
P8WQF[9%H4*QYR6+O N?L.H:2X21%/%*M%C UV]";C J]/X_T>T*6IYKM.48S"%O(
P1=D_U?B;,T-*@3% E.W^Y+:A# IM\<QG?_LCB$<K><E\\]/P@5=*U3IQZ-/Y(!RG
P@X6GIDT8:52DXR+I7B%N;AO"MI[)SM/;PQ7?#-'BF$4B+6#LK L7& S"]>M'4"CY
P.?]NYFR)EQ.H'4T00(X'H<F><I/>I87Y5_>A/U,<EE?<[6JV!M=Q*^X4QW/(Z-K4
P]U:O,#/&6.^*/*@ZPA5.4 ]>RA.1YY('UD4HOW1#$6P%V5WHBH>1[L OW?D8*(UB
P"DW0!",2(#9(-TV;BG;B59.SJ3NK4:2J/;OE1W!3?B*XE<.FX00SU5U,., 8M2#I
P>SMO3A-^YLRXKNF\=9A[-AJ)O,"@!,-FKZ=7GWSK4^E2.):G5;ALX^F9T,]N^! ;
P(1/R,;F:K0TD,_!P>,F1E,XXGW7Q&[P!W/N6UU5[,8]DL=J3YMNTOZ2^AX9R%DZV
PX+@&"6SC<P3KZE[1:W;2!T$;@2K%69-Y(>&P;HM1$Y//>^9^04P1L3+3TU&3H,27
PD DYRA-4X-8\O%0T.LD8?IXY<A 8 B%OI@#*PN#H;K^1O89O'[XG"1ENL=P#'WT#
PBFM%IJV6&,Z/.K(E%'A=\"3P/]3&"7Q&>3.X';%$X6$Q%%O$NQD1XQ=*@&:'#<#]
P?PG QA4[\/UUS5?%D?/W,%:6ADW2H>4UBE>B$26;;DJ0O0BXOYR'ZP+Y+ 04I6 4
P9LJE1X4L7+XL<7[/FD@PH%CK028BO7U>"\Q4\&-R*^E9FG/,@KP<U%A@X7-)]7D1
P]]'G:_;YFN'-L\E-6R8MZC=N:.]8=24%R_B/H<*@:O;GE4M<Y-B1T9.Y_[AI\T_D
PZ35@ZCD6,80;0[LNK[YXI6Q *E+H=P@9R^M;BH7D<0JS7SQ0>]''<H+HASQWH QP
PSF>556C4Y(*)3([O&09YT/"&?U0([ ^69Z!W2NEZ923U,R\.1T/[[AD :*OI7=-S
P]_OQ9C][H;Q\CD4I'=6O,1!*V#Z#JG#K*KKG(N8/4RB\=@;HE!]+A+E55SC3YL+F
PUCEI[TNX3M2709=$H?Q8Y9(P?S=>TCBW6\Z1I,ZQX_1.A/GIS;XT/\ ]2!@&;B68
PD-"_69'(]^\ V/]/[(FE&#JR7HT+,CFZ;53^ENBMD$!YG]76O4WH6)_Y'XSO_0E4
PA.LG9H__CZ_D0)IOI3/ )-Z;DF\""EV^(AS=>=T.=]9^&"^3)1_/C,J#^=$ 5-S8
P4K/5X,M6&29&<AYA?]\[5BSUZ2C2X9U]_M@+NP5 4Z,<I%;5VJJ4<[Y/K^=$S8L<
PF+2I%074ST HA\DU%5C2:TDLZRK5BVI!<WD K>DL$@?2PFN;!0J)5?::K3=O9.$<
PQPZ-.*:4T>PIB^^HF<P;TG9PEU5WN .U9W)/!\8<>57'%4GFHZ/C?N4.88"$YA1Z
PB[F8KH*V9WF;#XTN=".UB7 L3<%U+3YA6#((R4#LI&81+I;6AH 0*+YJ00# &H1!
P0K89$V>"?QFJ6'FSP?]&-W;SJ_G%%,.%16R(U/M#VP=;R%'ITY:+E)K9MIN'QKA9
P,=6U*Q!5UJE_$EX8@=_/,#P-J O!85C@C_*=OT]WH+-,=2^LH8%A(MI"I LA)I;6
PKDJD%!4LSN;-G@+HQ-%%(PG0VKR%"/KI&]HVYY,P*76J,U,4!H\J];@W\O\&,-[P
P)XRC,246&$<JG#.0BAE$:?!X+B1_;/@#+%;:H.>803D9P.2_::%LA]4(XYMG+H9]
P>)_@Q+G3Q3PAV82W^W4('+V9N$LU(.RW90SPQ1/RT3=\?8AS#[9ZABFKZV%CP3[9
PL=8QXV4)XB6)F%#</H:RN</5!_/:OV/?D@[% %)H)A''?9KLT/A]V$U.X#1)SBZ6
P!"O[B;\#$&!G5>OD6M234\<4VG?;1&U'IZNB.'* 7Q/PX2 P* S%:VC19CZA6RD,
P<4$>^S(0-&$?+S#L*'GO;I. =1N]T+1P^B+R%__D085TX$63W,&T9*6\PC$7W_[=
P(O:#_M%HS?_%1-$<O>V('@('NYW5P[.P=I(@!YH*_EZ@-+8I$]I@S"$T7]#+7;H^
P)NC%H.,LIG^#?%:NH:#B)^R'.A!'7R</";#;\844!&C$.@04.&A!'7[&WJ8/BUW-
PP>UM\.NW)<5)N05\/=@M[YX$-2EK"]X06'GT8B- '1:L16P99@=5+9[29SI3&:$;
P0J:'+")#=MC)NG.FJ H_U#<5-,3"Z$8ZH)'[)9<BS;A.&>5,-Y2KYGYGFC)]*TPF
P<9IBKF#!T$TFSL['O0\?SJZT!\7@*\(%];Y:2MTJW45G F@UAK>HH+?]*1(NC/XF
P^D,&%;/068( (2<RQ)GVNB-'PBRC_0WQ3'LKO>SW; X<97BGE9N2)GE?.'N7>,.P
PM@$7JE4>J/[\N'BCI UQK"4 93@(D_3/!CRNJ5<0LDS_^2P@\0.&K1N)3[O'@T-B
P1_N>YONE>/?D,P9X@5DZ&]ZH%!VA GD3ZE:B"L;]T@>%BJW+&,Z RPM\I,&4?LP]
PP9L2344=:K<5P_M6B,M+%P;R>+_(6VL 1'SSL&>N'HI2(DPW(3@KTD6$];:PI#CS
P;2D!OS&9L,/CY__XYWAWP=#VP4UQBKU>2-28-GQ8J.3P:/N2&3M'G3W Y2JI5+/=
P5EXJ2YP-@W(EWBMN )2NF!"BT+<&O2\XC2-SO^A(+>:T%.WW^PTC7>R ;\NF'.81
P.YSUE@7*S*T !#-8;0IT!+8H:0H,!K;#4KZ+J_;XN=U>'\DF^Q1&Y(A;*G7=B_- 
P"L 'A%6Q4&AW!OK[M<$Q5Y"MQ/B!AB%.>MJQ']2I7&MFQ"#F%*&]E!* 4U*)>3&_
P,*P<1<D" 8 I0HZ&%1YWY\ZOB,5 VESC3;BM8O_V"](7=K].G 2+76[L$=-05KPB
P_+"B#:9\GYAIU+:?N)ZKW!P_['$Q-)\C."-><#BDY22D'5&^M+%G> +/1_RS4%TP
P.3#GARBCH!UV))[A^CA_#*7L9<X[_AS8TL+G?3-X _]"&F=:36B1XQY9J<VWW\27
P]]/)YX$<!J_0UC#-\57CQ]1=A@6'OK./3945 YM;V Q%F><N[:ASV>UOHPZ"\R@L
PTV@^Y77F",!^[3KY/JPFW(6" JVS=L)/(KSJPALAP^B1]1 0U ?9.< [IUL=Z>;6
P9QCZ4( -F12Z]Z^QSNSK-XV3Z4,NP>2Y>U$TWP%-MC)[B8WWAZ[2_$"_Z07*P+P;
P9T6_;$4./A<1DAY"2QKHTA:(0KU\?23=?IH!(>2*EI4YV5QXC3>,D^_=>O:2]OZT
P:@$N$5P.#8/='W%8IK6*RF#WHNZ/(0:3^S,#V:_0B(3 &52L5=]N"^/'T(@N9VW0
PV809?VP3^<J0S:ER;J27!3>+Q-\\\:_E].8*R^J++WI2LUL">E.N6L[]=8/:!3B.
P W,7RZ[";'RJRXXWI8US_^_JPZN8C>K0^SZ<&["O=<T;S?DLT..Y#7<5$)%Z9D15
PM7JRY*G<@0%OZ0^% 3\UPNZQ)E)=B^=6Y-X2</RMS[P*1G7*5T6I<N-5(15TA,GP
PP65((_4O9I.6XUR]/\&H_P70@M*5QVOMB:F6:?5/"Z9&Y)Q?@SK#]L*U/P#=C,XM
PA$KI4M&=<E'AJ#3S5.B'%9P BNM;4#JNWS[;.&&6Z!733K^76HZ72/]=Z)MDVC9&
P(]/_6!?;KQGV'.>S\W5+!(F8^@SPAW-,WB'7""$4A-Z"YY,9QL)R85_H%0$-%@'R
PR<Y_>( H>:W>M^!S:I*/_;B^!K*=1+R?M9+V-2?AB3$>AQM[^D1"X%#R;CF&$!V&
P>3?P,G9'@G]9YIH,F,?&6YU%,)<1RW:N927YQ5K8YIVZ((W_L66M31)NT8(-9EQX
PN:Q"S#O3!MN&3@;>24X)36=/=Y$\:$U/'+SU>+Z]F<' L,R0_"?+(15VDE2"&M4&
P>AB =3AL8$;!?LE.OM(%-IHTENBJ6AB]IKEI!?E?G!<]YB@!ZCI!OI&!!361DQ$ 
PKA&X#0D?N6;@:[)_U+/'4 RY0UU"=0"LX8%/AB)*L,JTF&KI;,5AADV4WWOW:0F!
PC:N(ADW(@^D;06$4)S#ZTKDQ?X@)9I)K/S<$CR@HZ^C&.M2QKN6+VQ]&7KS,\4M3
PH^G;Q^C>1]R &6@+U7D/L\L;'9 7$I([.U_3J$&FBL^%7ZI^Q+M,5,<+_Z^7$X0-
P:JEC8\BX2,EQ]*5'1#V9GWI\S^ D1^_&+@+\LN\IDIS8-^79Z>"A3GT9NZ:LO\10
PV<;NP;VK0.:1<AY8 F$3^B#_A"1@&([2\@PA$^#R1LM.WY*DC(&AG@KI:S?4L%JM
P4_=CWLP,46[KL3TN>GAO9 ?IGFT 2+,#B'ZM<TKO_B-CC@=\GK0WRD,E.GV0@>,;
PV6@>?K(W-O\,66Z^L4/<BI,<9C%^+PE0HI%'L+S$ AIN+)A]&$CN[<B2@ ,)PR  
P'B#P3>7RG!R6O'W;TIK"QPQ1B<_H9IT\UJLKTA-E^B'O0E/*'M!OMOIA_).\J0,_
P3IE#Z$W<_,?3WUW2%4,3,N,EWMGFYU!VV,42@>,!WS@/B*TX<0I#<2ZFY3!0N#IU
PMQ)H6^UZAJUEDC[P;-\,HM!5B@'::50N>^O 42RQI!L9FXO93#TU_BX@"@O%'8Q$
P*PE&(F FQR]Q)!IF/BC5+ +9L""*86 WO,;1X/$\EG@*D'SGT!![F1(3&82&1CI 
P<:NK"X"AO,&O<;%H:H,[I:=H.Q7JA?J'V%RF_NNT)A6-:&=M9B@+C,?IXDOZ)"$W
P71-34PPLAV!GR0,#LJI%IZ=KDWE/90#PS0(I#SX+AZ[YW3V%[MIP=@ WQ=Q!X7Q?
PTSLB70EDF*)@"=KF'42G/T=AF6KE]POYN?NBPLC#%]70SFK->"'HU%<1RYT0J#9X
P>N35735^L^M\;O?<\*=S8?XMY&1WS/V9-K3(OQQO1(_$Y!92QRXGG(H0P4X/RWV#
PG_LM/J6FMV_L9U,SQAU]EMG<@[&@+]"%E[T&O;RLE O<-PDMC?P3JI6HRA(;;4SH
P='_RG7'8Y&PJ93SIL@N!'%6;&-?PL:&<6)/R[MP<&FQQ),*MP(?N:[DS4:'!S (Q
P'F-=>V]L]-Z(Y_W2HJ(E %[Z2+LX"1<X.),*H)G 64 T-BDU/4*(/5=&M^,L$".\
P!'^6T \FD).'\VM%1&,0,S,"=2$BDWVT7*5_B-P!F> 8>$^E*T_=H--:=3M6>KV3
PK!*"77%MZ'(U>'R<S_!V@3\T)ARJAT0.R;M3)G%146RT78/<%W;'@L^[*Y?FA[?1
P>G^#ITRHMD?7H71V" ]:APB9-IF95/ G35UT2#]N29PTOK[V2:4:;J:][M^T-!J@
P*J>THN!SFDE?N:7BST ;%[&\&A^=X]:K14BKP.?9<+8&Q0_Z;Z>/&.7B!6[X345C
PIK#_;",WT9;4./=5Q%LAED;Y<@[E^RL:3&.\D3/XGU)8>IHD^GD>7&9 Z1UDA;LK
PU/<F5,PQE(0?32EP4=N>&?NJG<1) 1RF&<S+A86SC$9:WFP]SS#BKJ)NV_/PDSAW
PRXXW(FY6"W=I(<A*.%L^[MAW!?9.<*"#BFCUVR"YW[:H:.OR-#RE./TVR\.XG!1"
P![:YR\"_/MU[<3I$MZCJ?U23BJ40^/,"3#.%K>5F3>.= ^,-]5>[A!H= PX\]VH 
PGX/G@:"9C]X.WF?MP6A0[^G4<CRGKC1ZC)T!%XY3G%/QDL ^^@:>$(.!_:\7FF0?
PK- ]4>[!"C_]\%3*R4Z<7ZVW+Z)B_=4JN,MKG7AD1:'A:< =B'T\M0VWW"ND&MD$
P%9.8CV>EO9I+1).JX\V,9$P&Q *-*O@7 &MYIK/4U\8_NR[\[)J47/DZ#-P44Y2#
P%KE(64W,++>B,\8+OXJP2.Y7Y)E5E3"=?.BN$!(&HAJ,EZ>)_[A4")\Q.3U/<#.T
PJ]KYCFPYF=9.Z4/9%;V!7L\;OCJR^Z9L659\>NVCR0D9[=1,=K5RH;$G/>:2OF-C
P'0O[48)7M$<4*C6,9&MAO07X J@16A/7J*L_:YKD*"[K6"S^U6@:9@4B]QN!,/KT
P.FUR'WIL/EKI*4# RJ$7"=89O&,:"HGS3:/2'..4R)Z*>C'N,M-L1/JAX85?"LQO
PG[56< $!#YMN98J\*3<U$NS-WC8E#G[^%88A^:8F"2-3WCC?RE3<-U![W(8(^>KO
P79KDIZ.-AC0RA$S8='^CWHCZ6'G\$5^(^$-;+N*[C?Q>Q)Z-XWEN-'#O/VMLN3V#
P1N_#H^+;\76 -<M*2K.R- JVFC#B?#\LS\9(J:NP4U#@I75:G\6KKGM9UQ?:Q5<9
P&X%#4M"(B"FMX48_-)ECVA4"OW#4AD-M13?5LN%V$7K_:IE_-A&:D@HU>7>"-AKU
P@"E1Y)L[H.KL1*ZY<Y0^D[=NOH?"MBQ3#KT39&H=KOO";&-#W<B+YL66#EU=6R" 
PDVQ2NMLLD<)KK!/:LTS+G[5ZS5*F >Y?,L=I62^8@-7N1,'N^EOG= N5A'L)+&)7
PH\6 #@2!,,ZN-YDL.5UD30R8U<?-/)IW</WYYKW$F%K]K4:G[?E[+$-)T4^"]K:W
PV\F# Q3@RM+(H&29Q(<HT@<AV1+_\BU3-D;P6I.Y.X.EIQ/L37<1:!B$!9E3QN).
P.:]6:,:+W\;*Q/D@A86F/M?"G[,EK]8$%[QRE=\.Z8=+*>%R[V'^C_4.T3L$RI2M
P)),K(6&#DNF>HWT=.X8Y2"6%#YR',2;>XZ(JVQ/*]L+"MI>J7L3>1"CU&ENQXGV[
P+2XF]%^J;%+(F(N(E&M+R<]Z!A0B/N?!];J&V"WG,>=_9^2E-R?%D:*MX'(#'H)J
P2RG4-,1"GOI'8T;4E:;R!0N^<NADMEGZ <_T44J&Y[E/BY%38<PRT3/_C0_%U%3+
P'6@_CTOCQ*$+ Z7#I_B=>M#:2:6.2%C;*Q>:U-D@+DGO3Q2;]5S*4$%:KIL3/- 9
PM1NV\I9@2NXZ;3RV>R-]'OO:63Z%5\->9E*$53I(?\S),DZ9R.Q"Z?@\V.=+C&?-
P1TBUF<7*+V$O?>E<JX!#J*;1!8)3AH9[;=,UH-XSG?.^#)>FM UJ4[=F"O[#_';J
P>5A&Q4\Z !HW>P@@P3F#GNH< :_Q>*.&8/R;R+]:._A\4(].^YZ"0Q'F1FD[6+'.
P,_/TR#H,P3[]BN$+UXU8IQKY.;\3EBJ1AT+?K,$IY@:GJ$5E-"[>70>(WI /=<(Q
P:&'^A-JHU<\T??O7CA#HYR;J-(.#<%A3L]KK78^S$$%NAPU >X@IR_-S/RO(IA\K
PWRO)_" W?,9#%4EID8([ J&=64OR.G[E6;*!LM_'G3\XGY8-^$'QDZJVUB!#;(EN
P/S&7U"%1*R0_9ZX4-<=+(DCVGTGOI WI/',\<([LAM*D(I% "!DB$G=ION?@M(.3
PEZ(CQ<TXJ<W,,[9UA;]MHZ_"/YR7R15@)Y$LA]JAR&=N5:,N?9)J<".%Z*N+.8Z"
PW<C]3$WC(6TVAOB=1OK*B:V.D50'<]** 9?9,9!DOQF]#& (EZ0.D/5^6^GG!]L?
P;KKO!8L,%_4S'46-CY@N>\'?N-]*7911 X'"'B%77H?B'!D"88/%R-W4V.*/=I/V
PT-]HD/B0VSA^4L"#97U>USKX/09&G6,%,KTS*93$9"C2$]-^+*&LL'*:;<Q*'[_\
POYLX_93ZY,]5R6#U6S8]<A20L<_FZKSZ@3-UR1TUP0]6>RF@2FXE@7<&['I?$V7Y
PV3F7D8N(#5A95C;GO@ZKJS7+U95*U>NC?#VW-J"/+(7<KI](5[&BKJC>JCJ&I4'B
P8IQ3T9&IHD5B_'ZA.#R_:>*T5!TUB'A0VR*%'N[%4T08D\2Y$9A"E2>)R-H^,!.A
PXY$TC4Z.6YD)2BAO*.>.J@0B3G<$J,P+T</?9M_+6%0W:1STLA<#0')4^' 4+17]
PH2'G+O48K;2DP-N"X:&"Q(<36#5'KQ/ @>(7ISWBV&V(G9CAW?JW7N=EIC.NOON9
P4HPDG8H8G'6M<J13I=NN5S\R:718%*5V NLQJEUN3OSJD<K/18_B@_\ O^%A@MU+
P168,A-S5)Z#_/*M'!D?%+DA9T)'^HTX+KJH9*V+.O=QU;CSBQ__>T@F:#Z ><=1)
P.3CU\[>RG@D>^Z7148(<6[%3WR]R^A)!*AJ 52U*:WS0E0%+]3/HO(-KNKY\2N=^
`endprotected128
`include "ddr3_parameters.vh"
`protected128
P4V[.70) ,).1O @97-VI4_[',2FN*E>SI&7 :QI<CU%-#(C8BI#3B[%D_V_T-=P"
PPRXK(&>+YC$MJ(YAO7.9<:K,L*7.6.Z"<X*F->KD[=;DX\H"O#T)#^-VE"/V UE-
P!C\31&95K N:Q@IAMTD* YWW5C>&:)V3HYBHUC-VS]<7/?'8S>E"68*T6+H."0:_
P[0&JO;N)7$4V9QA_M%D+<[[+J"O?:UCUY(M,W^:,'(J."J! 0$Q)!5!8'4@27>PE
PH'Q831_02+3U>2\2I59Z:"%>]1J%M L2=V8>,_)6#8+"2X<5J@%9+#<8)3@OW_Z:
P:"GW0CCI=J:P8_H2_/!F7X0A:>",5=*Y/"BZ8&\2T0$$?Z$[RXHIP'?X?2?ADB:%
P<_C.(*PTIR- EDZ$:,.63TF(66;E&1P^E'DRP55-^U#69M.?^;M>WN=((-W*//[\
PX/4!\10<!8@^A:!!5QNTZ24K07#3(7,Q5<%<0G5B-"&GW 0M)DP /3B<=(QCFO;D
PE#\W']+7@^K,_JMJ45"7#%&)T'&T0E+YZXX2YOL&N/XQUX02$FU&AITB%J[L8;K)
P.QJ )M3UR[D5BH$ G$FXOE=H,'.W#*'B:6.L3JR28KTR.*WV"%H-GX ]1NK:>%++
P;=U\O#+C<_8R"A*>B^>:9 *DB1@10@PI9*J?_.="F=[11%(R9';[  S&]F6459N,
P3<^N:+!]DS$TRQOJ("J,O16AGUAY\\2X&O07L:8EM5QMF61;NJ;*0TT\#2DW5TVR
P^PLJ_2DQ&QTNJ'5PS(IAL3,#@J8-#E:\4E?2@N:2J<= RW^L6TN[NU@UQZ=9S9=_
P^:]XBL?^K%9X-:R+2(%P\#L)Y.EJ!CJ4 =3/V>IP&+R^U3"HBSDUHLF/$B."IV>.
P2KSMBTCELXJ^FLKCB_5 )VB7RL/@]Q^][ZV^=&2KD=X'F,#%_P-2JQ9=+V37D-IN
PG<\LAUA*-%8O*/LT"NFX&J 9@6Y)P@@!YSW]I>^4F;!>ER(;/6O\JW?U27Z,(.N@
P74"V:4LZ[C^0\#'N_[_T(K\0S00Q*X%^^#)2?)R;9"^7PQ#D+.],3;:GQT8?LJG9
P'9G_D1O/F[N,-@F,,\ZL(7@\6LN^HF?5U[W)@^49!:H.&)OK?7"G:*C_D (-SD5+
P>1#9B#&$/B*-#[8'<97>E?=GK([(-CI8<K'NEX>*'ED"K1)$K44:TIQH NUOX1=0
P^-MH51:G&7X17"13\F208'# J;P,)'4GA<BN. )'@"K+XU#R&O?!U0:N-'Z+;K:D
PCY]]FW9BIY)J"]F/G4IKIJ@U@+-82*:^OJ&5VZIH+%]6POQ9-GH2D-C"VK+M&O=\
P\9FCM, +P%7'S-B\#[$:DBJ*-&-B@5W3NJVM+S.881^&;&#\"TLWZ35.Q8C>E8*>
P2+#R59*>7[JJZ&POQT)5^?PI W(S1.!&;]0)(:SPO*Z"[C'6;Y$,NGO<J#I>U[UB
P)GNEQ),8*KZ1U_R?>9[P=_\Q),45\5^9"%L^ _>O^XB_2$Y(]@B_$Z,=J$H:<&SO
P5;89G>[GK\?V5R2,H\"++5YT,Z;_ _/'_U4*L.<EV^2T'MM$4J4O;S.C,>"S"K- 
PPOZ0(B-]TJ9GEX>.FLW(<ID6BK/L[_\:!<ZO27\Y6FV?%4,>Q?NJKGNN]6GV.%(U
PI.B7>I4UOK]4F\D=LQ8K6OL.2G="B)(^*R^E?W_[PPYJPGDVD?M#)0=W+Q"X"* _
PUN%1BACV6X@AXXW>9ZJD;!J_T4 %DKF$79*;DCYQ;93\GJ9M!$ *GT><4IK>7974
P<WA)%WIZ.F8%FZ#SJ2VU0]US+'E^7&K[E9ET-S<W>1YQ_3E;5*^80O4/0E-4\F39
P3$4WL>.("$#-G>.B:I0>J6B[XLW^R&7^A:9Y0?5RDK2?#\*YC@D9A5W['JJ^/^,Z
PV;5$;E]VKV5-2)"H)(%9S,JOT[,4FD5%>ZO?PII;+>)HGZ_6=J>%<:DOYJ7OG:Q;
P3,F;8V.1=BV$$0#*IB'%/AN7K9LRQ?+]:^8/S4CT\0?] <(?U,U2ZNE,6V,5R2J+
P#:*8*Y'08[5-^(O:8*80@M$\*12#.4Z(<6)0'AU&#-+"5,A1Y%C@9!4A<$6<@CW]
POTABT^ 7XGQF"Q 50CB.K#;_ P9C)I^)>.XC'NJ'A8AAX"E>T=\N>J(Q"Y8@3X5G
PDW QNK 37NB"(AV-F=4C"!4V^-JG36U?BF*N/3T01H$0F]?U@27O,8G'JV+CJ>YO
P<EL:CH26_]0S]3.HL(:-$_Q7O] M-E%?W@OW(#O7%H3+9XA4U^5!#XB\)3D<>&$F
P&!Z(Y3LTIE(3KV+0QKQ(D"YQK4GG);G(%@OP,E9F(PY1R8GAW%1#+$!V5/-"/IJ=
PS,X 4UMR]I.[_#F#<0-,.&Z_^T+6-R3)@.C^0 ?8'AU.?6"$@BHC?XUO7[^(9MT:
P2%%(V'-A3$_BS09?8$2C:^V":)):GC376-K<Z0>=U$JO_<O*B[/I26(Q_.ZOM!I&
PH8E.SI7"M4:*FF30!97\=7['M'/PT*M?BVTX[*WBI1<J/8^(=7WBA G4:\M/'/,9
P,]AY7+2>Z9//ML."MT,*4$:G\ZS2:WP9BU."3M7RLBLYH2SD8,HF&%/K]J)<TDEI
P(Y_\<8IXC1.(A&TL<'(_'&2,B0LP6^\1TEA'&'KGC6+K[?@Q6Y5//]G!DYS[O#B&
P1VZ 0QL>Y0SCD&/M9NU+<C/=P';0H<I(Q,.9KQ<D,CA=+_Y14YN0AT<\.H=RWX <
P;5T=_1.HYTA'1)SILI66UECX61Y.$3P3%V1*>CGS::XKLIV;>/Q09XV2ZI(3]G:>
P>(M[7]R!FA0CA,X\[7C9V5/G8JTTN<_N8]J@E(W5V]"43:G*ZBMY.)(/X=%V_%N/
PN;"1'TQXG"82Z;",@#>3)204-+I+ZW&U11/_0<;%\ )=$96N5!W/Y4K2KZ>+!$8F
PS90==Y6]DMVKML5_G':2#;QE'5?WI66\0@LBEDGZ;U:S#L!619Q+>CJ<*5*X1HHC
P+OZF*'D3^5>$/'3DEIU5+]-B)0Q,RSTW^1E;.J<NK[[]$[>U_Z\4JRHQ^LT.PM/^
PN.-6@%JR*734&[&.@(['N!*W1Y+UP]C2\+@]-*?]/"IM[FXOV$7YF<,O@+0NGC8\
P_=^]$]MD==6>%QE5!H@QG[,0Z@F\>0'O?C*QL\]'7HD/3AU-@MGC.7YX%IB_8[QC
P$F?ZF@+9TVZ,<NIY:.27,H"K@+3L.9>DV-@-<S?J]C HP\"X0JE\OT6KOB(_U<O:
PD3K3AB]>2)6=J=N55#GVH';IH>V7$"C961$VU$R#N,0T<2,5TL/\J2(0A%%D&6G 
PBFLA6K6*$BWKV:/PAKZZ8>GY;I$@"/%5T(<%7T<,+%)&BU-*V*T5+@TO#IU6C +T
PL=$ H*KCTG6244%=GY7/Z(T(+_S*?JO9FNF!I.SEKO\\B>A\8\#+^%J\(&N ";8V
PEITC=M>J3H)%)?BKP7;267O=M-/Q%SUR%HX'7:Z]=O\U(;C_FBD=%>V2BD06/"M%
P<?530Z%KS%3^AY'7?EPZU;'8]=9MF Z @#3:FZ2ZC%:^&[+P]LO.&1X-S>]HHB8]
P33DLTLJ(@ENH)F)?)=6'!+&(R>LK=<,Z?5B7I<$U&\FP7<<W?%2WOACE[1= )GR#
PLF%G6^O/TFITW1WR<*"D>]J[25 7IP6VJ7&__@^0H=1(\\E#%PK=&_CGC>U1Q<)-
PUO]C3/U8KQ!W3LF0^0#W%OBMKS2$CXNI^DJM=N+N1-Z43$G=FGI4A ")@_96$2?B
PV'0/P[*1Q]%,DSHP&OO>O9V$65 $:U%5O'/R1-'(8M)7K9L]3 S_6X$^29LTNU!Q
P6E;O;!F+W1; \4[8#.@H@2-W5%,Y(X%D^FR 1ZM:6]:-+ ;[8GTN-B8U_]M4%[[8
PXQ-(,$$UC<]:D]DP:O/J)#;*^#%W<&0)B"QC#NQ.UK5)BD!(/Y(K4[&\M=V &VHA
P6KZX%A\IX";_>NQ1VXI$<BP1_D$O:"C\*U%VXM-5(,E"EG;Q@&8CX1R8". ,1\5C
PAAD/BJ_G.=EZ0[7B*;DOAR;+OJI[Z9L\8W=%C^&@2(%W+4Y6_T42K%]QZ7GLW1:!
P&A"U_<_61P&1B[K$]5OXK=SCCPGS(#2+0<Y;64%MWVG6(#IQ+1A,4?\FRR:PF?TV
P%(8_U3^+[(Q#6 PR[7=&ET<:J[S_&:[SUHZ.T$5-QQNV"1\9RW[>]%J]ON0^-I@C
PTGLQ57\FZI:%)."$C!BCWU26+@30"DY[4[GEF3U93VI+3K%>3)2W,3L FH(ST@[O
P^T^<;W8E]$CJ0+D+]9M8@U].;=;X[S]607(%1H<D_Y\/O&2P*=G^\QM:COILW1CP
P_^D>P4A^]6,=EC]"8XGDXW8FBHE3+AM3.*.0M",];1^'7BMG03"4"IY.K4'NMP<6
P#?)#MP1J2AI?/Q."#_-T9C$<//UN-2[.R5$;(7&I@I.6KPV.."]0Q)CS^$?_V8;T
PIH/PGU(>;3 H:^):7A:Z;01U2DRTQC"$P')VMP88W+/6_DH^S=($*4?!MH^EOUV.
P[]Q.T)]6U>NE)S:0V"42AG[P1=1B(<Y02\^"%<IHFU<J$O6_E(;<HCZXT<O<*D@\
PDQ%V?=LS6[-W"?Q^ R(XI7R;*V<6%871*@N#^Q>[,U%-,,<A0TZ>Y!#E6#N;C),Q
PK.QV?2 97-EMA:<2'SIRNE[S9!+=(28=P+C>D=^WKC6L6CG5]Y:EI'-'E^='^V@=
PM*1:FB%20+F__ISL\,F48(5;-0JE%_*#<JC S9,+_779XUT];F]Q<5TY)732E>B\
PI_WM!/O4J<*!V:Y2%&#^:U=;R.(?;/]O:H@<7C&R^AWDES[Z[-V.;)Q!\4\4.!A/
P9_\\T:2*5&!@8+0%E4Z-?56 D.CKLUN.Y7*_W?L@A/X#EQ(")F1O\E?WKY*.8*I?
PLAJC'[=\,[M)$&9%43GQ)HQBHBDKN_QVPS_" ZDS;2X@[R>UZ6<?H1R2P_8M8ZZ:
PM[(4[X7$7ME%I8U5DD-LZA.PX^NP$:BUI2,^)/<DF)(;W U99 %%(A7EI^=H5CC\
PEND>FT/P/]T$LW;^V@%_],H6/%S\LZ4[IB"P+<-4R!5@'00]TBM  Y1#_+92ON..
P$FB_AXPP?/ZI?TE+KHM0.(RWRKI%47%F#F:4S<Z_43'.T@G;"73.$EZ09=:,Q%%D
PPR/\+5]L8#UR!R1@_&^$03+AY$]R*OS3=_[T=BD0BQ3QGDP)(7:^Z\DE9J9EZIDI
P_&NT1_6PD5IA=CKD!H%%Y+<N6-E$0L+WDVTC\^]11D)ODE5ER908;<D3-6_6D6HI
P#PE_IM$(=8F1Z9!RC]W,>U4R] N.G2#7;!7.0%96_>C^W>,_,BQ3V)*V=]RRD-/!
P@S703S_+V4YFXX:QAT)@""GSIG+'F/JIPJSR[+^!F*]ORC,[XQ-W91+GKJPXEQR6
PVO_)22C'2UQ@_O=PQ!MZ9OT\,B2]J.I*$*A^(FM08E9@,..SX# .Z<)XGB:X@U>C
PL>1,;NX"BSS15\*MR77\:,CA".M)=_BP'?E^:+TS/NF4)Q/5HIET7)U-A<S(\ K,
P+L6D7CO (%.(,<G,@9:Y<2JB" ?CDV_SQ*X+#,=(P%MVU@I\%VTG5V1H"[FG:;?'
P!:F61UCUZ^N)UHY&F42W0>U6XH91 S:8W;7WU^AYN;OZ#*2D_CU(+E^G.4PQ)0^Q
P2\,(II5$ZV<]!CVX+#747)2CWIJGN=,W\ N$ 4OM'A>G;](/LKUY_9HI]V]5WPQK
PB]UN;;6*T9N-+U8901[K4+D(ML6Q"XO _(9@N*GIX$?;2B&[!!>;*4E+&G[1_4+O
P\I(L:83;,Q\LH=&>29\T#ACW&B3CO.WP=!-JB;)WPN2'6  AZUB,V]]M$NM5FZT>
PJ4!*B3[)=)R2!  W&^W*3R=WVRFU&U20SD"PM= @*7/<O8_Q_EDX)[U8 04 08Q9
P8,T*L]P*N[A_X4-7-_S74F]>=5,6J.Z+0T_S/7 D@=ACZB?#F=^1WC!'Z+#50X2Q
P<*F=6^4Y6+L 5[+(*NMTOX)$17 +HD%3;BYP^O&)]V_=\9^R_24L1B]'Y^I6_B^G
P+#M1 ",8[Z9 B#0XG5UQ&0= 2JYV-:Q;P>;4@Z&WV2H;E]T,_N )5+\/(O]=/N,2
P1=J,2C3ZYT5B(8?=.G0&NJIE'L,0>>>\[PR"W@/$.DDS)9[;9N8%\)O)8D^3(?Y%
P: KH=1&5, DD:I0%9Z%M.6]?RD[A?6'-GQ3IR/$P6[5M"FQ)=CZ@-?FQBE3=C4QO
P[X2QB*3PG!,13RRBHXJ#+S@B8R?@9F7\M4]Y<KO>_'>N9"]GLST9:,H[+7*@.Z)M
P(^'53PRQV^J6WY^5=E>J*?I DJ$9JI.8QY2A;3V<+NY@RK6S]0J9BH'\UQ#&J5J 
PM@B%#0^^>!3^)2:,?8J74W5PY^TKWZ/,ZIA+=TPQ>X%U %_*3KW(N%--$,#=.<76
PJ/<5KI>X+\(/[:K\?<_F;RS.0X=>!@;@!=])?1?-CB-5Z+7GA#V-:=H,-5)\O:U!
PKBP4!D%>Q%5>8/R_S(7TR6B4(\IK]2S)0/HQ(UV+!!PT7NKRK'D2UXHH-*"\K(PX
P-=W;M%X.!_3BJW6%&XY0.F^TEZ!(.Y4"%$FOE%$O;8]L0&2$+#4HTF1D"^;..N@N
PXWD:,]NVE+=8J'MI"M()9 W(.J(N#_>'??@$[^[GONIS9XIKM:B,_L$U:Y/7]]ON
P',ZY0J %PM9RBX$9&1MUR3X.G.EOTH(CL:M()%L;AQW-"AFTY$^V"/LN,Q)O4_;A
P<@SK?MKK_62_BG%-#_V<4'57V!"JX_9886O5[MI3G5?>*XY-'G_1-&=AY*/,'^ &
P>E&#Q:G2I>JA KMUA&, ]QD8C(J?2."M[,DDZ^^DS9K3!)GM@L$_%<R-X?X9:<WL
PRBR6R#;"7V)\J=6V^).PC%/J5;J-*JEP A&Y(F(^^[TK-%HN18Y'3)&R*O^[.B1=
PG_*.!9U/<I@U!-O0V#)M'1:26+A<>[V:!P=4$24!C@AM"/[>>0'(KN9=2?!"PT+F
PXBA=$85:&2YJ@\WVDH[.%4V/$O"CDFV*1C]>1'(PZ%O)P&L&T+^8#C(,5!5P71PB
P<C)#)_]KS??0KS*%9]U+!VP_6@Z&)5U78\00GA.L!>B(0>ZMB/> (9<''L"8OQKC
PM;>LI,KXKU)W\M&@]DW[."I1N/6CC?!;(HV'YK#*2.<:67UC?\R16P"^E 81?GOB
P(?\P3*47U@G6@=##=#&3R?Y7Z&%>(\N@ZIR.:'6&<T1,W=N?+*M#3MVBR=AR5C1B
P,>Y*'=*9=JU#Q!TGU;:.633ZIU[&:,W.F$GLN+^EZWI_#F5X\2,RXY9),.^MT!AL
PTFDEME@^:46EI4SL<T>)TW&A6F!@SUIU]:H;1SP):IE[KQO-4D>@CA]_JC'1LSUP
P3M&HL8OP1AW3L@G8BPMH)P*S7!^EH*'I&W+*/JAR[SJ3:\Q6;.EJCE,7,SA=TS_[
PB6#HG0<1,7P&I^-@T &-<REGA[!"9WQK"8JHNAZF2O%V/TS64W+*KKU%'$LI(=$@
PDW(_:?:2@YZQ).[*/PO:-)SVF?](Q[+;"E;:+2=.0)-VO!,GK4"@>W=:X$I?Y;V@
PS>^-(^1P<DPB0@]!L7!;G*@M7N\M)3K/^<_Y)^PP!C(DD*WD!YGY9'Z0WQ2<-L(U
P_=9"P'K*H(UT8&S>+!NM4QQ9.ZRR@)"R][A2#[!>=(-<9QLY5"$?%\0747HK^%\.
P5^SVP0A[J,] C$H2VMS#C0PV(<8.FQ[B%M_^ A HY 0*7SF[9NZOG<CH8=CHQI K
P^1XP#Q*=AFKYG%11.FMDT4BC.WR62HRUR9&Y%7-->/V.*#C=F6DU%AVQA%P<IWFD
PT?.-]$6I,OCU0 U_XD-TRE\.VKP."DB__0AC(4QS5;9@>U(1\O!Z;%4V\[!DIE$C
P2DS*Q$*A9Y+HFZE-9SE" F=++Y]2NBJSY!;.7OZ5'7@S_EUJ-GBPI&]R3S(HXK\(
PCC8A3 CW?V,_]P+3?<;P5>X5Q7L[GLJ9G8;SJ],_3D?$$U+TLF73?B/IIN<EF;PL
P0=&ZBP@+-@  O/)#[0<+7[-?TJV;"?@N\VNQUNT*HX&G&Y<[A&AL!+H$S=%M&'D 
P./S<1_Y8DY.0AR.(^>(CKS:6*D0 2IZ2X<4OSJQTBX#1 ^:RY68@.VD\QM:N2QWR
PUE/]_Z1_L$DN>*VVG>HR*"7P\!9)R(^.V#'WIRA_&-P/['_O6RQ(@Q'EZ"NV5PV0
P,.KH#CCH("V1B*KK@*P:?#X;N9PE'HS@,-.).;.=M8@DA.V[O/QD?NL!?X7J#MA:
P=4/;ILB@&+T(B36U .Z$]$."%,4Q;H,C#*#[8_\4S 2%/5EGCTW!]_78>93 3940
P15R%#5,69W4?/<H%KL2T&9ME :52IC9D"V6) >A0Y?IQ'X5@![ATM^9O,'1)P>1C
PV4?FCMII#NI6)#Z D0GVR5T/26#VNC3)JHKMNP5];%/ELCXA>IN>3Z[V2=?B;6$*
PJ;O82E7%1'FY0[B5GEWZ!"-A'44 UN3] F=526<I;UM\<,S,>;0#9M#_'!%+VI]>
P!(\AT!?2^B$0RI%W,[DQ@/DQ&_-@5]5BQ^/@LNP8 8N4$C/$QIV_1^1 ARF%:?5B
P3D]^%]X-"JD1X<YL;CAP+F+-N(8>TQ:# Z=GEK#5'?M[D.!.6J3GW4BD_B" \.&W
PK]_D-#A!D'\/U<I\Z 1-]4LQGI2=CDMCTF<M7EQ%;K>.&#0M*J#D)N/Z9YSAP!K+
PMOBNLI^0J@D;X2AI(Y9/NW+%AA\5S"">>:OJD-.>AB+:^^+M []9'HZDQS?X,^0W
PQ--3V.$6-/O.**G63?BIE]1ORD]14=K4J9.Y867DI O4W8*^>(M.)2N'!GZ)Q!M+
PKC^"<IX+?['BVZ0A\IYWGH #%1[IT5Z7@258K4V+,^]('(??9G*&.8D,62SN;-/?
P'<Y<,IZ) (7G$*V JE!IAPY@NO0_NW/Z 9Y;#Q9QH&-:[+I*O4RT6NG)>'?S.4LB
P^?:1;-,A!K>FK"PQ)PUIBRFKWR"%  *^MH:X8'>4VF?] BI%7;/X.[R#2O $&@+Y
PWJOS%V=TMX;.38RNU".9XU:W.R0>++5T\:,X ?=JQ?BY)28F"A3O#ZE9/H+ACJ/C
PQTYW"GUOG$,X'MP>HJ$*/2<%AO1CCOTBQLX33QD;9Z9!WJJ5E31/1FU*!F5C6,F7
P4>@."2N[KN"&_^VJ5N=W=^A7Q,S;*HC!I[S?O=.9%7Q\,G#R@370PAZ>58 I_:43
PCE$V53&+[;WO:S9-4_\]86/C18W=#BPR!C)>>5B*4U9=(C"4LFNY"8CB37%Q?H3.
PD"D-*FI@HSO2[=.L(_2M+LJC/T[^-_TM7I4W[#:M7&(A)E;S2ZUF7X\^+;U9^T$7
P$O.-H'5C.HK$6DW/FY<X%8.^;R23'>8N<YKF04(CMW\[7PZ0%S[/F99;Z#0R+IU$
P50X>W8PY;T]0( 7Z) 6\G&Z0.H;.-^98W+3D29,/Q>%)D_""4+R=$@SW^H\8*'N+
P L'+/DM;)8&--1#S\]U.GZXUY:>9$6M@A)8I&E$%]OK_Z/\++[R>7W,A@S+]=G!5
P&2V5VT7QF:5I#K03_@)'0SQN4IQH&R>(&&D.Z]'F][\*5[3,"@PQC%O]P&FO= F!
P23G11.@P%!CFW$G' %"("2*L*QE(-))JI599;=5!BMN%J,?0VBL9H=U'AV.8Y$\U
P1,:A131O/AK_5S739F<+V<,YX\ ^.LGAE2^F'6Z>:V<V<Z#\RSHKM0H1[E3^1*=J
PQ5&J\3UROY@=FH&'@YDNZ#=@Z&'^E[6W*.DCTFQ^Q&! QI_R+U4AQ_7+?#S2MEW>
PK2;HJ(ZT!?+HM2&*(F@GBILC@X<S@IRZHB$WD/@I)HL^Y0@ X_E<(^V"/E^./U=A
PD<]\F86_AKQQS29$)CU \HM4(^]E6.;^.9"S+1!REUDE_E5SV*=QJ!PK$(/([1;]
P:LA]@#A4J]0?;95?.?"KP_;F35FM[X B9H<',EW>:;-#=[ (Y#[GQB>'G S#6-/U
PT4+')G)%P,I@929I<\0&EE7.-Q Y_-Y1> UP<*REU'LR;2-FOOMQFJE/-%5=:7]-
P'51B=E!A3R[=A9K8=7ZX1OC#/QZ1C_?Q[Y&(3@3Z:<^W/9\;RNI'4QL4[LMT?5IP
P@+== ;"VL=]KDM2Y+PX*/2AH:+V7MIHG'NC/@.TL!U4;Y6FJ#/6I64,\\7D&*$EK
P;;S<CFPC%'\A.]T\L>I 'Q! 'L2WV_R)2>!H*L$>DO@KL9E[O<-LGP_T5P U'4]%
PD2>P26\,$SM4*D! ?5M)C]A%=_[Q93Z1YPQ&11U2$><!(7)ZPPUM5]BZ"S?SJ8KF
PRT<%@-E*OC$O1_-,:#6<O![VL5$Q[+=L!2XUMY=3=L.\F9_2Z/9]$=92\02*C6,\
P"';Q>GQ_'3KY>I!?L<QR\S__*.Q;ILRTD/2 7N0OIXC(J"[?3!QLSS!2%RY_]R,-
P6F(9KUA3]H1U ^O0:9'0338"YY4UOGEM^&?!BO"XHS>!MU6,%7#;HMI;"2XXVV#F
P-= 0_SL[G"*S;X=*%ZRC#E2=%4WXM55>(G*]+88SIF,?"J.%M)/8=X4=ZYUYS]0-
PFX<IS-ON<)^GFP*-PU76_2'KG4'[.,[@/MTA*P3"E#SQ_7@0M%(M=G339,<IV7,_
PS0O($ 5B"'CC^(8;GS?;DLXA"P2ZQ/U6M. G*VP4'Y1JS3/%LR)E3I('R9VA2XZ^
PKQ-C=,2J0>#["XJ^.'[JH-0,S^?!=1R'F&T0@U(SNBK 8>!9";%I<B!DL2?8].Y;
P\&?UTRA0*!LO^+W"C!+C>2:NEZX*OUBUN]TLC2YX+8@#J2*LK;ZTX03.WVL]?;O6
P0"K.YN2,9>*W@M5^[ T?EQQ>F1YH!6Z^-QQ4'?I:IH\[K)RZ,]9>Z_&"./DE6VTK
P>]ZL><C?E(Q30@B,,N.=\AO#G^R8K:IH9=Q3_TZ-/.<;EU)X&3/Q=&#$/M*@8:W.
P)]U520E\&')3X*$4:T>!O[3-36J<=$N6RM\5/6.&@-ET6(Y"#'DX($X#,A?R@*QW
P#=H[&219W'>AMT$2E34[RVF&J1TLK*&V.0;(>M[<%VUE.204&53N9A'33/>9J.2E
P\ @.D(I8&<=ZF49-3G(([]<_V;G'$ULF@FNEW#)5R6Z(+GP$/ID!O.I"5G]P'E12
PQ\@*-S&JV ]R ,U+)#;L9P<I_#97%/>G7D)RY%:,A(RIYKC9E7 &P^D[&P=RZSW;
PRC&'[R;G<B[*P?J0#": 97")YFO:]R")=N"QB7XO>/U-S$I1AN;4CSCXVL9*>8C0
P-4;S4(ZOV.&>1P/4"/&CEWTI;"<&QQ".'! U)N:T9O/>>7.W14^U@"2/8:&K"-OE
PV&+#*. @ >D#H':C9D)\BYI1/?*E#K.;[\^S3K.$#1('TG)Z<Z=69R,GV<19J$P*
PH$LYB>R,6-E']+C56Q^7?@%[LXC*W!<N CNCE)K,#6<8MP*PUG1K;!*D?X%\WY^D
P0R*WL>)36R?6MOJ%]3%1]41/47ED\$3#,[HT<*^F&WPK MG[<?,*NT&^E7/C%&2V
P-XXMVMN-+65(VZ&)<B^OA%E0-?G):%#PS-#3V 3]:L3,356#(P-V[= M\?PSPNR<
P8[I%GXF1N;>X\P8>#A;IX.M5S'T?HAN]N'*$5+S, <)2R[G*F2B ]7%, ^ :7. :
PZ__>%.9(\V3^BOEFMPL (A_304MC8Y[6-?-![GO\3Q+30H#!OS"]ZO89'^F=[E67
P!E76D^6MHVJBO'T%_#NTFXTZ9.=N-!;_<3UT?3F:1ADKXNSXVW_G2;@EQ#0YAW]M
P88D1!ZW/T!C5-0=M-_5F806J=G'-J%ZJ*S^".Z1+)[=Z+GS<$-%0#;G!A'K%1,LV
P' \2%JJ=O&\]=Y4XHWHV\\SRZKS3-6'&Y/\TJ9?2ZEB,%]'8W_ &8Y.0NQ=+\YT\
P$B3+DPVM0^7RY*;7HOX0;@TS,[PVRT]O:Q3T5)0RI+LK0@=>SCDURR$WV &A.)<J
PT<[X=)QER9H,E+(Z<NC6U#TOF2%>A-FL69B>"^'J3_<R81@HP_H0X7[TZ0-H*AL+
PI0K>,YS'1_T-*CE7!^4MHJ/K%7<4 0+6'^;Z>S<G$KJ[;UAX*?X]^* B@!)/-ZHQ
PM,;;.LPZ?H9R/M?_(9LC]7317C"5C6?K;W=E(?Z*OBUZ<V0M02XE%H:C+?5XW#CL
PJ4_/D '5*DN%&C+UOYF2X:;Q-\@G/=>.I0LKHGF;U43(#'6"!C[SUI5@'GHNQ?ZG
P.I9,5_P[!90%2D=FD@ G9K8K9>*=*KTJA8#"RX9_<+Y.]^0#[UM/K'3T*/56%2@V
P6CI#W<<(C%LLFP'SIEB)K:CG"N[IU0]:7.VN-XM,RF7J 3^5=R$0J\/XY-G[;5*9
P3PG$CB?!2-S?+"$D7AD #SR["DC WIF#C*T',&'ZIV3;D,)RY]@&#&1?9$1=_'&\
P03-Q/L+7N2NQ"64JDY9LEP WT]1M#4Q@Z,#=&-BC=598#&!<(2_^"9M;#47&/KTE
P7$OXV1)F3!0%N#ETX-,NZ4+-/RU7J[A!X]NJ.!87Q1=>=%0&9WE#EU$F0X(%9D8Y
P 9D$U4/>DJ4JX*I6ILKH*DHK%SYH#YCGYZ_U$55HLN)T8KE0MG$TO!)/Z-2V\'($
P; 1GG6 4Y.QA4@WOY_^TB>2B(]0[08)^^EI/_"':=[)Q@WZ4BPK'B3F^L716=]3Z
P<)@_XB%>4_O<*"Y2B!&'U$?46U9*PL\17)O*1PXVVV.%>6R;$+^IXIX)NL!5Q[CJ
PG]O\^+?J<YVT1->":!Q(>''RN .D^-1]AUN:L)%_*%]_!(%7NX%.WTOGEHMS=^:N
PL7$Y?OMDJN>['C@HZ ]%-IU()RZ6*.-V)-+ITX7L&22KH[9L[3X%NZ:DM:TE94]D
P##IB>%W#A&DR?+]WWEV)7-C&*.JHF1>OBGEF&*BSS(]:DZX*PA2&*%3GQI=W$Y95
PM:5.&'*.4_,;=U*#)!IDK/B>]6OU 8C+2?M#W5<V0,G# +F_8:\P[P4#.K,QA]N8
P)*J?;C4^CE]Z5:P^F>[37C"@IV'5-F6S+JIJA9]9P#7$#DERE.SW]$\[)9/>J(K/
P,K<D]Y:'+-2V-NB+A7A\SCH2=$\?;F$@B*A?X%"YX9#5Z/9KVQUXD<OUI;5))DTE
P#YR*O7*74^Z$U@/SFP/-7?B698730D$8,J:MJWMC:$P"SU"<U@=7<%T?M"14IQB5
PF#9_U@>5-C4%>6E-\ITGS%:\H71;V.RG[S3<&?%\T7W)*6X[HP1$ %H*Z]]E\=?=
P4(:S99=4YNY:_3GY7HWNT5Y.$!6C<;=7+ R-U)[.XWC9.QBS+[D^<%3HR+M!%0\1
P+]=R319*5DQ:[YL3H[0D>KM@:L7*Z6B LV0\2GN-1[(4*YCU2;-Y5E; 7@&=D91B
P]@=A/!]IBG0*3P2YM*V'LV\YMD@<P]"A XPZ;V'\.#EGUZ1@Z=3K?GC=4&W,F:JX
P1HL4O^M^1#!E=8%ZD9=JJKBT/6\H_[$*!T*04Q'A+\/>A[)76PI(10J&^OT$W39U
P$NP[IBY!P\PTHQKU6^W3([-72CAZ43#'^A/&>3>.#QHDKWA4VBP2SX^B)9B(5P%3
PBJ[DUF7F->SLRX%JL'#\=3WFX^C=[TI?TQOU".?>:2^'>#E3.DP$M2?J@';!<0YA
P:2V(O998]$]AC';U3VFVQGSE<0*ZG1IH\>EE!/JE9M]9W'SY:=M7&LJ:B#SRR6EW
PT1U/@+E82)C4+(WF$Z'LI+;FXEX^1H7A(_4\,_6$#!6\U (]LQ@J37O78>->"AS'
PQL/,+Z7DH9!5V:#E#W$,]HG].R>P6YHD@/C-4CS&.A#!*<*3[ WWN71!.FN[K)YH
P;07?M5MGGV<U5(I:@FV2WW/-&28@$Z(Q^=(%+%<"CN8^;%YUGO>YX;G@ <DN0+"2
PMM>C/TGI<6GU:S#Z^_^C,8<L&E^G6:W_S(H9U]_XQPGS^JKM>)*42 _J-OD?4KSB
PZ-)XUD_7*".H@L_O_D.$&APEF=S$B:)$N8K/!UJD_2-+FJT*7HM"R./6+*T-;39K
PL-_GG.,&(LB+C&<9^-58@/L$K<I%\$C"!]/NFQ]3D!6WU7&D:OY3;>N&]Y:D&=Y!
P/Y53CX.>[A7+XR5PT'8%L%.?"H#5"'[#VD)RM9*Q3I+@1.&,I,E3>%AI[C&[ZQT6
P82J_7B.)^W!2L6*'<; 3>6K]")-HF55MQ3+WAZGM[F!2]ZM7/S_.3S6$6F2.O08=
P7<WUD^6[-&)WD>^/&<B#ML8FUF]RKK7N,C),V'I)BI;BT4F143G:U7;[/CCJU=5W
P)%4:<LS&!2VG1:6@'Z_>R5Y%^)5]U5E(^:GNM!3&T]F#N-]N N .">=(81PH\N+9
P7T106#:86VP7^%28W>3GFL.KD18',@;A#>=O0=?XJ0A65Q4R5N)P]&*%!Q&YRCO[
P.IR6V(<<A1N9!9X N7M"J'+8,0A@TX$NN<$[/6%C(F%ZHR=KF7E(QM&UO#?JRW +
P+,.WW(/+DMO,2 >'K(-/B?W8PS"7TO1(V?QA*?E@Y'";,DN 6]>#&F(36)<20MGE
PM?@\=Z=;/)US-L5*KKU0VVDL^'_[$BI)N68:(SS:9A'\^+0;;$GJ_4YL.@JEI'_R
PCZ+4:YO0M@U1M]WVTYHL Y=%(&MJPCAPP88!9@]%S.UO[.NP4F6[>PE!IZ4B0C#S
P8G//,=83>R6"73^_I(HW^MO41*2>S9%;!J-4$Q0*:GK^.]MQ6))CC!3_SR1F<5C,
PQNA560= S=O:\QS+8$9+^'VQ*PT;E5G*6/Z?X)#B2.NLK1RF!KOL/>QG<*AJ*E[=
P':4.@NW/6FHKD_Q-A?HQ0QP*S=[0AJ=:[F@<:R?K8_L3&J9%_C43$!ZX2$JJ@Z]#
P(5R[:S%\0QD<[H>+<D%\2?]Q(M;@/8B%G7?;S#!L_V>]1.-I'+,A4Z*@5F7OGED0
P5#*HQQ^P?!!<<0H(2A?D;QCDXP]M<F(KV$>>;/<:@XHX)]R.7K>_#J6 ZHO)Y 3D
PX]%CFZ%43*^^'!/@2%;J8[/M>Y,@XP2$R.G7AG$*&U=_=B=X!(4#A--(U)X,+HSZ
P]1?2A0@=-K1$;K[:6[@O?B7AV86U32C\[=#&!:63BY'$A12+1U*:"B=[V8.2.LN!
PK9NNC>&&%ZH6NQUA&)6OR7\-W'%DY#(D9 N@"B;EQKZK4J>-#7 1HL IW[A]BR*D
P7U)^+56F+W?T_/_/(1#F9YY+:8HE"><.X0?^V4!.Y<M:#QM4(V AGH?O8I+]L&Y:
P$TFDM?YTZ@'$CD6WC#$K"QJ+%)PC(4$SB\H_E3^!S_Q %Z&D[T**.WAKA-MBO^ '
P4H;J;7:_1#>#"E>:;LCQ&%@&53.4S=X%LX NE5#7JO>0G!DIZK0IY\*Y!+D<*"S[
PY4?X>7PSH29AC3 COQ#%81O/56RANI6XE:.]/H]VNUC&^$JY'W"T^W2,Q_@(N\UD
PIJM7R)3.75ZGJ+4'SMR&DJ92R^_LAG>XS)+'F4;W/V=\8SZE+H7V:U\;6'&^S]V>
P'U-N6XZ4V1S5M;#@A?^&<FG#J=&N]F%\+<J-Q3"Y!X"<4?[<SB('O-\I7T?\:"J-
PD2VCS0*%G<&]/;50>A(@S"F:AGR%NBZ:1E@AHZ<AIZ@\SCK9M:V*9;4F&'DY:>I$
P C)U&D%C!B]\_2YWUZG[ID#F%>[B\-#S>M1*GK7C5BTL>_.B^GUL6P[T:K-"9[DS
P13M99R]V!A/>-&AHW0 W2')_(V4 .'\F+/VS+(<#HPPVXU(%)CH]<Z?J:'#^7WWT
P? KU)!-4NQA&06)$KT_TC79!5,-1_H_,U8CB8D5],LF;GXV3F-=MWQ;.0NJ'ZX<A
PTH!,>6ON*>7<HB"C^\'I7TY4D'UEH]"\%"EPJUI75]U, !%C/TH@9X*YZU: %&0+
PZF,_EBR43=%UV@@ME.Z;L(T<=?M2A56<V6O/G/ -B@EZBU.%X %(V?B,K4V4HZCW
P>IQ3  J[-\Z<Y!U! 4B?]I.V$41[N[UZ\+B]6!O@I(TFW+-Y,&6-M.,@>GO1( W0
PJ>FKEIV+V4N&5OH4O7/"_QGM<!OEI[YJNS_#5U%5R$-1'Q+@YWGE)+,4<,7LNGV6
P>"NF0X*-.%'%GW].__BA=L((/8?8O%=(E7<?CK61!#D'RB)53+J R_!9]T>-XJJW
PU 8E:.E&-U<Z$8:S&5L[&;N!-=-V\#N>730W)BIDRZ$/ZE'3ST%&F&L?N1#)KV-)
PP<YF]BW^XI-4+R2@N,1[L I#^"D;85*W<HZOP5$^SU1<:V\\O%9&+.%3F$8W2;QH
PTU'GGJX'H57'/TC%D_;^@&,HREF(\S.PYLA\;<%P6:M5#@>'T37"4O4LO4;$AV],
P_PUR.^/BAK'W&O7?\OUM-)B.EN%<CVYK@\UNB^X!\T3Z$NT9->,11FH1!/"^,CJ4
P'411 -:T\%,(^C1F[3$ #0J\XOIIJ/L:<L+O.=)%"&^$/^*KU7#W(\K8_:TUZ>N&
P+%4PQMN!TFFC207X8(#^J-OFX%!76NQ$H[CB@Y=JV#4CV;)991PV_],-#AT\3T,X
P3"PH:/5KV<C4TA\5TS@4;OYF@\_? 8R/P1WE_Y*:GS^ORGS/D@;_MN\7G4F]9%"\
PHFE[B;)FX;6SR 3(\17D'</DW-> (KH]7/+K9C[-_6U3ZY.1+0.1?E3]--WOAUI[
PE!7+ <,Y'XR9#Y(N5%"9>5WD!=ZBTYYZ[SOYF-#/Z/KP> =3]?Z-"6,!<IVI'%/V
P?$=0AJU X"Q3!\:[S J\80/36MH/W'X9!R[>]LL#ZI85PG!%:HD34^#P'7.J'?$1
PQ$M@)&@E"M/,3HZLX,UI-!-X5/;IMQY*L)P:U1?]&-KF\;=+,WL"30BGYHZB')$C
P($//QX#/#!%\;OLRUZF/RL<K,)&;IOI'S6>P?[-4X 0A%=LFQ=2Q7]<3M[%P50OA
P\,58.E!HJK.F0MD:@C%*#E1IQE:U4.F1=V>Z0FJSHK/196N-$F=&/KD(OJ<>M^M9
PHZVAIYF/O /2/'1P6^ \";-]!$\:#K>!,[\?0<*ZD$_8;-0#6QF$@[?SJ@EX!K )
PZ^W/@/L)7[HF> "ID###>.O^E(NT?YDEV,I M09 %KK^M[D>M)1"=JL=SL(D2MJE
P M3O"PIB]Z8W="-\9W3XW=3U&@'?GR;ZJ+U&,;DC7I*XQ]RXPH[?%N*8W8%:LHO7
P&$0,<_V3+NE\P[F.HP#J:CF=[3%'URJ41<7[Y*@+6_[R(/I*P0O$88_-!"( ,!B.
P75W.+&#2/=05/'^T98R\O#D3&-;LF:\+5[P1IEV4]&?XER5C8X=BFE&^3+,%&,Y=
PU.=<2&*N/\/52T8.,UT?-6H[%N5[D\_UV@&OL%?IW.;.YG.4H73WXI&Z?4DG/IEC
P(B^JZ_<H;ESTY<SU$-IBU)L@/T?"4'=;XJIF@1>7L\V*AW&J^#/C3@QTS9FM36(W
PWMF$DU\)NNI3.866+X>@^DTD&N%KR8&&RG0C;ME;@:2%6Y58WO.?4)!6+9!D>CCY
PN,#9'-XITUM0[YOPRO CC<49 0@/]LO@4-MIR]B4D!YL;/F;0]"]I,?&,%#Q5T;P
PN]17EWKZDU&-F6F3<E_-<P("5=8T-G>K+6_*%PSRAU6U:DX7ZFM1[(7%.L1J"C#B
P,>_?)=7!-(NK#KTA5#TUW!BL_B&(D%E^W%:+;KAKAE.ETE"3=LA)++A-:^QSPJFX
P30C"W!H@8OK'64-^./5AA'J0X)&4M!L?S*F.2 ^,)^A7GEA\<F3Z('Y-),=X"5_L
PWW=^.W)K>S:N+"KPW#B>#BJU3JG\GGD2+:9ODK)5HJ^$]N!B%,$MO_4L1U=/803M
P?9_&>"$W8--A+,M06X>K2"D*Z_JS[DB(3709M' $XA?#?#P>Q>%[&N-QIYI![I?:
P!L5%$?R-S=$AHZ?.A^N=0M 59L)O\X"F'57A"&/^SZ/]'2WN]7=!E2DJDM]&TF((
P59#HCVRGO/@R> *.GU'HA_B'Z(8KEB%X#H85+J',!%_O>1A#_4BK>J_+3E9TIJ8K
P@7@!M#9__80GT9,$]JQ;'\^HLFQ0)D:[DZ&SM]7/^"&X*CG9*\B1. +"'H%_Q'DD
P[_6^47)D0I2%<DN3V3:C9Q43V0UB949DTV3NPC06Q9FX<[JZ1=Z9Z5Q>Q&6JC?3^
P@_S;+18+"=SG?_"[CNJ8#__:%@[(,']]_[/*#OM)HVP0-\T/)4^#7ZXABF7W_2L]
PI$[68^U<'P)YUDT8SRN>&U/_.,8Z_X4<[Q@7I%7\*/TXFP14VV)?H16(*Y_1),(H
P.O#I*FJ51J;9+6M+'8W2&FT]"0M_Z- ? -\OB=P,:#)8,O]?'=$AWBF_2([3E4'0
PMNN@.EB@+YL":N9)4?^A);$C#CENRGOT7!=6 A[.>K'AG6U,X#!([DCYZ^5LAZ6Z
P8JGHH OD6;X^G'.!";??G3YD%PNI\JHM50)AT#TY3)2)I(O:E%G-"2/MB"Y9,M(J
P=Q<AYPV@7(78]TV@W_.5XI)+[@XYM"OO/ ?MPA15U+SUVIY'/E?K5(89JQ+N_-.M
PGOX57F6F'=Y:@MIM) \*SYNEU^U\,BK.I_=.Y"X_K@YYGU*=<)G&K"9FT([M>T= 
P_W*\^:A!2P]SA_FC,/$8RY0:^=+L0\UWGC'_5G(PX]$*+<],25[R5?CV3ML.66ZG
P.Y3*UDO([F3"'TM24(S:^AJ4J)E0WV%Q&.#X_/#U51U,Y>M9W#556.8>IG;:+'F2
P%2/5]"Y1'*)]?.[#&>3T/:C#0 ;UEBT6UW1!JZ:55*704ZQ0=I&8QKLADEOYSW;7
P(*5Q!<PHWZF?A[Q11>"!X'S[N,[0-V6=EQ],0C_L$;RJ:"7K,+L>U"DHI;!# (K#
PS"JFK,].93+L=&W1BM[D2@;W LD))TC)E%XO_I3.V9AZKP-$^E$40U43]6DC:N)D
P$-8\3YWS;UQIK[Q> 4,93MI1+/WEC,2)06^?%T#GTE0A&S%*^)&D2A(%H:DI%>3?
P2>D%,0,MY:>=RK]F(T<_0.CW@^@$Z7+K)#\.Q;?B @EG5S)N01\T5 ^+'27F>]XG
P<!%$QVQ#< T0]UR'U%!S;(SN8HLT%D7;FT,D+64 ]N7;9J*K5*^;V=243;A/57#&
P>X#,/"V?).*#_S_<KZ=@"#2JV@9<M'DH5&ENBD$99P<:,JJ$6W56'V$*C1,*SDN%
P$<PVO+S:M@2I@MLT,V2=A(WXE(R]#PQ!R+T<V[-R:7>Y[[P7?B>U3T<]LT>'N#"^
P-3NM^$9Q#I@7E)+(YT"MN_O_*%6<K^>KH#0E^E^""O?@ONP1Q!0(=5+?98+!#+E?
PPRA+%,%$YUA0S74]%.X;1,^A:K*6W_%.UE=0<\5^O^9&<6:%.7IV/<7&EFP%?13V
P$GS&O*O!*=H@KQ]ISL7$(C-B[5N26L!OF_P?K\="Q%WP*HH\LXFCZX-N]-#DJ1T-
P5)-K-0W4H<6F'B;]/)*-Y7!^F,ZC</@VOR>!V-*L@6KH(=FA#HL[Q:@)E$>LW0*?
P3H)V^6+;<;5HN[HWR0EK+4_X35W%7(GWEFZ.ZVNC7+L'GO 8C!#[?7OG@@\'1A,.
P<N^T'*#-KTPL5-Y)P]A[G4\E7-WR5'7LN,_?I>3(#%9%JIX8YO<)!+'#(%JQ[BD@
PP9%)PG)92AO'5G;9HWIZ@6CCVJ'7PB]6V,)&.>2>3_ EK6 ;.3S&#:UV^J'2[8K&
P1U-0.4U$0]R8I0I?!?5N*;7&L'0BS34O6EU8!Z08DW#$M*>>E^D<3HVH\#GQ!(RH
P53IHG2<SQ\&V&P*]N8LO*9HI1''.T-4.(JG+L/D$&H,3OO1CN;[/>674S-W8L"4J
PH/E%(U/6+HEQYJ;R^I*$)<<7+H39KUV=HYY:XVW]@#AH@LUQ4#!0?'Q@"5BL1FHG
P^(;HBDAZB[C=S8H+#B%>VT/QVDQ7=+OB)J[L+3B;Z[="8]C&MTZ:5%FR-)4!>S>G
P1DF]S5*[VIX)\XD^TF&UB:D"2-_G7N]LI'7YK+U!Y.&6-#;3YZ-.G=D'F*2_0Z[7
P=HQ<DX0H0DB*SF1YI-@8E<6=RNL#<X(D5R3\C=/IL9S3]&PE ,8W#39+-K1F@J%A
P2(=;WE[$&(.8_HYUF]ES]S8+K#I1I46;[K8$">9D FDL]W2"F<NL4OBK5EDA.4@N
P_OI&Z.S<3,@!3)R=N(-98<UV05^,JGVFJ4#JH<2O)^+N)1/D/K+F)W2>[^IVIU7>
PUJS,0N+_&H#E8OV/?PIA)!GXJ/]R3@C,0I-*O=GSQ>/SO)SIL>79]/;H.BI=R9&K
PA.'^X,?Z+51+T3=KKSS(;PGLACW&2LXJA54.XNOF+O[EQNN&E/;=>"J _9K1\O<4
PV4\RBL6_M!OF)_--^HII=GO2%!F@B/BU 9K^K"+I;\CD$MDG-I:>5K;9ZT[LU_3P
P^'6HH#L(__J_3SPM I#;ATYI5']/=P"J."PM:'BVV28Q#]PCT(NVA 4HI@G.N1\>
P-3$3&43 0$,N7'Y"<@:S\)4R5"5C5#4CU^:#*5$^&@'F7YU-<N/SNFK^.12)F]ZD
PLE!I2\!Z4L;_'1,3Y+_(_GA)#\ $,X*!5']6Z(TG"17Z%60IH4=]<#M>3]>5M\6O
P.M<VG_%E ]D  G$(Z) I=:U4H=O =1@S"WMC<>1XW8%W83@?]1%#\=[Y,7Z0G*XL
P'LR/?QZ0RZ7J97 <GN>1;?_=V]MN*V4'"0=MEF-6D8+YR_[BZ4U1BS&]9VYI$@T#
P";>SK2M)&(R2VA%+YB.XYT:=XINJ@08-;_9(XQG'\R<0TP.9.*SO$']1;JR7+ZC@
P@X_XZDRO5!:194!-Y@&ZK-3N<W@&*K5\_UHWM$Q)402_.E\T:I&'0U);\4RS%ZF[
P0*K_1Y,<-XI>^F_2E%<_.R-%OSKN_&ZX>T=(T3_BV!9G*BC^.PW:/'_H-KX(7<%\
P;SU= L^V5UI3H4M11VM@(N8Q',U":%*4.$],GGF0!CGH_(JM!]0F9,\!KO!B=,\E
PW9;2R7JMKE$A+LX^\W/%O(10Q_!A[_(S=3!$0&T7T9?=JI.;R]+HQEV$J15JGL^9
P'R\YL-28E=GNI#%"E1:)ONSL$(XSM\2E$0=N+I,T:S]CGB"_"V17W=6C+.EYODR2
P=P_YO7A%R;'I I"$ 2LX1C#E\R*X=4#_@\+A[3:D[<(VFK?)?WXNDKS,1*+AY<U<
P@$2E.VJT\;_4C4[9E>FOF[1'N.&4,QAL#36<$9 ZX_\7ZT\(S./CI'<K&9%^:[SJ
PL"PYU95@N_<23K!"GO!!7=X8&%A8L%@6K @?RU_57;J=^IY$2I?&%6DI3-/"]_UO
P98&]!.CW:%R=[KD&UQ=Z6R4OP!.%*+\+*>P!6#A]"2ZLN2>7(0\P[(!W2QB9>5O<
P KG]MRR.)XUEC1VPTP"69>[\/$KDS[BYE [HM$ZGG#/3F78^OFZ-NJ7XAPYJ!B(D
PJ[J5C<QE#SEBPZRB16HY1=*>X.^8:V6PIFON33+X?#?1=T?,>=(MK_Z9CTT04R E
PG7-Z:_'<E+165F+52[N2;ZHB%,E+%LN4W_1&(%4#7_QD'+#(Q"+1-SU#HHZ8DC!M
PNF)NPQ4KAKS+0:?R) %'%Q-76.&EDC17"'/P,"!TQG#$O7WU)F\5?%%K2"?FE_-&
P 8T/N!5_(-YKR3)P?0EF.)4\8G AT&#4"(>/UQ K!5^\0;/BW^<B<L)7<?(*?7P1
PLH4I+R/Z%-PM:"FS8S[)D['Y^?=5S[#*797[0&3=JLF28?+8K:?*0"R.1<-;[%XM
PK(!GG^]\9E@%,:^0OV.J?PF+?6T;'UVV1A*8@SL0: H;Y+$M6!.0I.S>& ;<XK75
PN*7MBL!UHJ[^N&L7O!@A/[MS<N\JT03H:4-\(9M 736JA71,;HC*?%-_ E!&U]**
P(>278G)BYOV7-,FG"N:3"4#[$W6=0L73V&V_R$+6V]TA6/J0;;IHB+T"G^R_K1NT
P$I_0K#TJPN+GR,*-EM6D$F!<8A1AK4:N6H'UG,M5 R6: ]?0B.Z-"3,*M1L4& \?
PSS\EZB_[.UVNL?Y3I02W6*X_/4:WL8!-U-S&MKB^/S54)V^M"3)'UN&I /S'QDMA
PMW&-0K_I\$5_6I][- S3,J'(\H!+M[3HCD$JIFV'1R!HFY]BY["SMX0J=B.J,A0D
P-SV>84P@ !Z_/D31#0UZF[%GJC!4L2"G',CS!%L 5HZ.K!0"L-'5P79B\5U&0Y(P
P!IT9ND]B/PGKK+"B,^5NB[ HT '7DH!T^E538<"DW6G7.C'B\SE<<JG)KUL<VGP>
P;#K^0H(@<+"\Q \)-][?8>?K_ZLB9,/>8H?)0OK;D\?*R&6.!8/=P7\+-AG4@1/R
P?WX;<V -B5!2+,6Z97Q4>)N;X;O&=-EG7XV..V8&!J_0?\Y5G&KR;E[.*=:AR53E
P5_#'Y![]SVS^0U*.BJA^P-UL6KGY,>[C^1!LE4KAG8E$:RCYGA<PGL.R-2H1S#0G
P9_FF<^=<PU%EJ]Z,D::.(M]LI-SK)4*:\48RD+Y@X30'*B"R MVOZLE*9"<+1]+\
P3H> LU3F@K!!/.1;:B'=H;IIR&,['W$2@K!!1LY\M]1K@<8#K+,@V^?VF>M(:['>
P#UI?V!D![G@&5^3G5V>"#FU 4#^*'H>5$;XM8Q-&%P.EU.D9;R-:LPM96'W,G./J
P)MN2!2A08-/)K.1F8 _Y&J1^$"':PF*@"<P$?C=Q7'A_>/KW^+!_@7:MZC.\(=R-
P?,.@&IIL)O>('.7( +GN$F,;$@V^&?GG\R$NF(2VVNF9TZ$2TAY&L.S S.O_VRV+
PD)Z1G+;V:2Q1*+B&,5[V\":D+(5OT<^)*S'9OO]^M<)=_7CT42VY;B^AP'GC$#:G
PF5W(IY\5R^J/I(L4KY=?'G(TB5=0T[3#$KS@# S&$(F\$E<^U%@_U9]2LN["FW#M
P;BE]D\9C1^<75T\"H>_]RBLR/*OQL:5.2?!*!F%LT'J\=@'.LF7 E.O,.VWB(A"&
PTHW7HU,09(00_>00) ^&1Q9RH$\*8T 1* +4DEDGV*J$,;,'Z=K6E-FQ,#HL ]MF
P=&O6#I"(BL/G'2N9KU]J<'K1&S15F8Z<'K^8*5EV;]MISH]H2!,T,LENEC[KC=A9
PU:+S,^+LHV*F!\&C&:21_^9/[7J7UJ8JC6P.F6&!1W(/ZW4XN)BJ\H[WR[Q9 B.^
P9*\[%4:RT28L%$SS^#"URC->Q/Z.<-$$KU. FVF=]VN\.24@GGN1[6Y8/8LCC;!C
PQ@-\K.=:L(+XU9R7<ZHQ1CH+W2XRAL9GMY;2+((>9W"I"H60]FNB1F@*B5]W9C6B
PZ0ND:'VN^+BW=D47%RHFM=J)G,R:9G2E=%+ZI.^FQ6\BW?UE(Q0U8?D_=@*Y" T'
P5-LA=3$#%3*&VK9]F8KK>3=+?",ZV4?3 :0))X*SEP,A(#LM@:8Y1Y/O@2C@LZ[)
P3<@8#4&@QLRH?1OF+L=/H:_)?#_-X&,UOX%(0E4+>Y@A1#)5)4;:^S6?I:>98GUJ
P^GH6%I&_F]N94JGD"O1?;:_(-Z,>9B\$Q<[ -6O>I[PCG3R'0/,:]1KMS0,#9=22
PI1#K]BGUBXPG!&P]2#"-Q=W,PN3U+-H].[LI*7&@*A$QDM7N--#OABM3'PM^/E3<
P^(BW=$X3'!>IPBJ^AG=*<-EWW>$'B\)+ NW*.WH_@'O&B=U L)Y_+[7NBEUS$G?P
PGRX>8E7P:4WHS@]"GB0H)O#?WJ6O$.]8'$]?J9+Z4%"/D34H!N/_7E%A_>N4)X ;
PB/LM3#&E],)V0RX[P'P(;RRX%8P^8]R\AOFY<%.O(\]8OYZEN$Z<F9KQZ05.7I'3
P><(5K :BRD:^.WT*KCB>*'U_S80#!L"CKD1J+_P>M;MM6H_(RB);L^9?4* \DNPS
PF[WXTRP](S>Z$\%QGET>-%)"GN*P9\H&IJ!:[(,J &W_>1H*_,P&&/NH;X[VY/A2
P',Y(93_[6CNOQG(3L_]&&//6")<#(ZH?3(2_(JN)8&PLO.O-#NFY(#+=K W5*[<\
P<6"O5<DY"#9'E;Z;)=%9_X""3P ?.E Z(*VU?@]%J1T+[@W"R7STAE:.6&4,G=1%
P!7X5P?=W=:\X;*M6;M4,Z1Z_LD1IH#E?67_CC[MQ-2];;-[NKU4&#R.I,G@%\LI7
PP77$U#:"$%87IN60<]EP!^(F6DXLY9K>K<'W\*Y+1-'N-M+^%TWL 1G'D.@#[0-[
PZASR4ZAOK=I]X=B:U0&07VY.@[@,S:^'4A%?HD<AGU:*$>"L^L/L<5@6B)1/Y(/5
PN.G#@&1C_-=N9@I*/W.Q+XO[[3= \@M!*/K^3QZ1E>CLC&H+O@2C4"@0Q<P6N840
PG37#MU8^%)W7W1?41CU><%\P4+*9'<3UMG._2\YW1_4]W=(JZF]P$=I\W]M.."UR
P2OT(\4UI7TX-^*G'7!EHQ!7ASYN3,>*903RG5U9=!$;Y<A^K)I<+!Q#*(],=#D=6
P,F4#CD*7V9!M$S3=)7P@MH69&( _HU@_2]7R(4E#SG4?I36G-+>\4:E.'U8-EFM6
P3A)^SU:+S9'*+4 2)AXDRU!T.^Z3A_V]JOSSY\X9XCC(;L?%\@EAJ_=)S&_,UD*+
PT<E?<NM( T$+45?E]OCVAH$@(1Q2K7:RJ/PQP::?-;4;P ZNN7ILPM1.5)W$&<@Q
P/^Z@1-'K&J4K$C2+6Q?FO#(P\C"<S%&(BE:).#W<=7_2=$-'=^F/,B(*!I:/CG"H
PF)PC<Y7^N>\I!^91T9![K.@T8IH$/5GB5PSV"%:&P"LP(*PY[S/%\6WZK4DD9=+?
P?ENEAT /K0:"3="[]G3!^%+OL\=+*,FJ-%[B2S")!K@V8^-Y2N%;9?4I!%M\D(@7
P?WM1XRS[QDE$BL,PW^ 7\7- >UM'"486J!S$)Z7M0R#(,DH"A+K!R> CC0])_=^%
PYTK<F.MOT/"]QT](N1E6,]28%]>2&>V\&I3+8U*QL^0)DZ<>-BRT]:3 &X%>FLUI
P'I92(36+W&<A&\K20&NC/($_81N;Q].".SLVG\Y1Y*2]]>)";5MR7?5SZG/%IV'+
P+(1*DR2K;FYG>=59RY?A=8ALH'A'#(MUKB,P7/E !TJ T1KRBIJ8#+:-"[MY5-[/
P_U?^%(!* R[)FZ3?QW6"?W-K!&;4KM)E@_X8#[U>;0CV.SY!LP"CO>.)3-V .?]L
P/E]_>U!'3##Y*N7:XM.*C<](8IA2[0L[AI_U!E:)L_TM!K"Q)7HYD_<G%_2$EN2W
PUD:FJ:L'#L[2$Q!FW&UK(EDR + 7#O/+US%M;M+#_&X6O.>'ZB<7+A2E\=09<NV2
PCY/40D4[Y2.>U[W<U,<3VPM:XG9#?-=KW,MGR?"R4O*\I>2X2^2;0/6M1W^HT#$7
P=C]S7*Y29 +J\J#:V![T"I,:^_=,,M9ND&,"H5F[&$Y"8K AR^5*TC39?=WY,E?Y
P\[(/%/_J,W#\/%"!D?8^F< IT'TN*(E\+U@<5(\ILT'WY>%$X!6A'GCX?_%624*D
P7^^ \]89+/0A*[^0.0*<URX>Q\ZC;)'5&*]WMF#_)#AXT,5TU)S6RM_1X$;&B7+'
P:DT!4Z*RP&]1AXOEU&X-W7SU):612BAY'?L(29P,K4^:GT[IR!0);X=(F]]]/P<U
P]IQS2;@^6V;0>_'I>>ICQA6G_E3N(6/95]0BSS/N]H+*&K('200]N.&RB(&Q;](.
PH9&S0A2*$:^5VL.V"2>N+E;8Z&76JXDZ7Z"EFA-T_L'PS>/JD1?L81')-'S5_WG:
P[*:\=:SL@+$R>'E;V?^WQI#_(4=IN-N@>-9OFGAJ,;B!K[W#@9,%[]V;, KK_/6J
P$_"6 $ILK^.T%E%Q<9Z+#3W=\_<"[2->Z0I\?RL^[DLRJ)"CG%O6/^_6/Q<C=2 /
PS0[4]6VNE0NQ!/AEK_-!"XF(&QL,00XE ]27F_R>M2-9S8\,49H$;NF/+UI:SLN"
P$^TIJCRK56BG,@ #-$R%4N!BT&&]QZ=U)J9B-IWLH\Z*:HGHS2@.4.M_\3W?8&S]
PT3[G95,:^=-.>7G)!.F#6#''WYMI!5M &SE+@+!TU')D0H3*WQ;_[M"IA9O!!<N/
PR:%28$.*2G^T2_$K[&B9\(2@*F<&2VTU[UF9X3ADB\UW(T J=QQKE]?_>K(>V9%)
PG$S]_[V=^S"?V.B?[:+(89#(>N./]I)$;]?^=RDD1 63Y)I_\O)QG:7DEB23WHJ^
P.\GVVL3F*K-,H&+M]$8,$/ CU:$9EV+2$FD,X$E<+"@B!O5^1SD6NRKFS*QB)#AI
P3)QW?@^>*I;A9=,%X>VP?X;+<F*U?89.Y3DQ[8Q?.:6[E[R$S?KUJ?%F5PTUS!?;
P28(9T .?*MB+V=Z:/W8QL9NL>9XDBVUIQNGX^GXJI",7^WY^_H3*ZMA&'I4_K7 /
P0IC6KY-.3!37A+>LH=[#(?,49?H=1F;\%RKR.)]:D4Z=^A!8B?1XN$N\6MB"TI_G
P2 (3**H59OJ5@\?&(]^+<_?N)WH3B)_78(/V[_%PM8G"SPA#PM(V&=GXW^-M_8A:
PD)8[C_4!V4LFRV;TH[4:%-H(X9)Q%?J!GKFF(T8LX#%:T_?T%O#2:'KN_*B<^6E*
PMT33C7T;59!(-A+^.KHX_-&'UX:=*-*E(?64K8P4FVDH;?_@L_1+_FA*GI",+%&%
PZ7CY*GO>]_;<X7NNN#+-MS8'2XRDWV9))1=%]CV2"Z]9O]+SV3%?RR2I]SB<-0G)
P&+L_,<6#AS;*.#76:W+7VL:80<IF4!MTY<@$D.KF^])$\ZB%#HDSDGWX;WD,;2,?
P;%0DLM^(4U@ (X)&V>.DDN%(S7_/DVF+WNGUE]Z7QA?20</$Z8/+>3'$-L"1='CH
P;59@?)T8EME-*'H>A.2WI0,UT.IP8**YC45V 6J=2X")<R2V(4HJV*A6GB,VOR=T
P#YX%W,VCA@^BRHES@<3=]+T3*!X4I4BDF1^AJ 4E^X@$;;O1ZVGEL(Z,'N*F)F.B
P(X?K_!A@-./(0"2S]_I09LY-+A=^WB.$^TP\_;#R+8XA'B(JGWQ;J!6VN _P.3';
PM@;I$,N3QY%;&2'Y7()\\0AH5"\#Q7(*D-VNG]6LCT4Q^UC;F,(31REG\K4;UA4?
P/FHVF8*U@U D/LR3='4.[LNE=%-NT4IX05]SJH[L[*N<J;?63-\JA;2%%!98V5, 
PA>1>W;5<T2C<W5?+26:M%2C2734.AO,*WY9[DQR,EWM_,/)P3#O_W6:H-M@2X).'
P^W!0(Q[]+,1YN(2/,U)C'1CS2_L'WM2>K60GX;;M"T:*7Q@=PE UN,,TL.<?60\V
PX <KW05HM$,:@(8.JIBT"LWZ?5E6=O_F%1X?6ZZVA62B;2M5"#92 75BAQ(8FM2Y
PK75 ZE,M7LE?E^86&\R1K=U1:QT=[#6;E[Y@IB+Q[$QIT 3!F>4T,7"^G-86+'W9
PZ:S<5SF.K(O%5[Q0;<CC*3M.51SO"UVKAB"XQ5GPE#&7.V$TT>A=+[M_8. %3BR<
PEV.JJ9@P_/AH)4R4H9,TVQHC[@Q&%Z'5)'9QXL42U8Q*B7(G/^)D\XS0B;S)SMFR
PK_%'TLMG\RGCZUX4CX E6)HP#.NTLCRT;E;ZX8J7(]D'D.3I$OQ%OG87H\2F.99I
P:ZF2.EUSGQ2,UIAW=6-VOC%R\UND"6/&<J5#_"CL*W3X%[,J)%C.?*PP$-I(3W\L
PS[;1GUM9$]!L\#R;1!5R^19Q,N7(T5*= N >>Q7HC98%]<<=6[<F5RXM_9Q)RGDD
P.CE06;/N_7*Q5>%6 T+F2"?@(#.A&FL\*\>";N,)!(/P7X(:QA,0+8T!%EYWWV6,
P"K@IZ))$T%] [X)L1(*(*!_+]DFVXO_)K((&2>7O%X#?HOB2.9ZBS23%6/8?<_E;
PN>(&Z- A3?>U9(]X??M#APW/."(CO.-.?P.8%:-.JOGI*&K?@G3#%1:?TIZ,N:9(
PX@<PY_J"GW:Z!:O (HQV)"2SF?ZFN<*O++;Y9>44!/9K2AG#SP$UMJ:D[#K]PFBN
P@%H2S0<L"+?X]#H,K78GIF9M?;=7TEK[ 1?PEVP[D\C_5O,6E$$@<F>L9Q05^^:]
P 35H$4 BS+W1*Y' R>7>%>*)#_,%D402?*.7*MCG"=%X62I2O9Y;'C\^8$UO\+Y&
PGST'YW*VY)Y38<BP;KU%NAMM@T<W0JB9!CDHZP[A0[:&IQ!BJ=G8]VW'-,^IE,Y>
P8?+?2:%<QMXZU<7Q%FG\</R>H_]^M/2Q7!N1FDWXQ?:GIN-[G$[>=I#^,L,H[-,D
PN@L#6#SL*Q$YXCM=D<QU+G;9<T!#EX TQ!E><:%FFJ8@>X#>A+^YH\0L3!%TPZ#O
P#)M^JT.D,^W[E??A,\X3R\,A_H7#MP'_;6E9M4.8H)+?A^WKTE7+A.&Z6^BF)VO2
P-]O\6;R<F89)X^2M7I]0@..T!9>J77B*-/\</:57J3?L'!(:T).?U8@<D3CX:I'?
P/)_/KR8%,1NQDHA"TB147AS/M\@W5 3]4G*,_<]8CVHE\G-O*.I,GJU;UDR]?(7$
P&U1/IA+!U$5@&8,?=CE_QCJ!_D\PS.0/U^QB>')<)DJ7B@Z;5_()2&[C1H 9?U%.
PN4?7H##&"X3F095&=!YE<*G7^?-U.#1\10[N42?WCNP$S@EI57(D%285?R+NL\-=
P)A4S*8S[L@G=/85 X1;'@.)XG[95V<?ZTX/$NFT.EZ6L;VKW\@N1.^QON CA,#+,
PN.8#QZ\/_JKVO,*E_GQ$LK'."X'E85WG0!,L\<+;9@Z,_'"9.8C 7/.AWNIV?PF(
P:3WX#^FYJ]+4^,L%>P,U3J U7O]XE]N$'CK(OUA!2.+QP@V.H,OZ-(KB:O5=*Y' 
P!)-6,S[%22Z[A3C02#W;S[K'UIJ!_T]]RB,W<#-19^S-F *<#K9*XN<A2=1^A2(]
PXHL+%4GK]4=W.3!+8D:=#KG<5.NNZ1)2+8TI"3NL<DY2;W:L-P7 0@XXSE7J304$
PV_73A-+Q$J_H;W]^^F\S;E9XW3Z3QITT=CK0D\VZ9VH]8,TB]]=)"@Z!\D.UH<FS
P90Z_Q65WQ#QXM_-2";4V=PE(VBQ9VP?*4PSG_>OK/*C@R?L-?YBN%GZGD:XFJ,]H
P:=0&3$ DS_/[GYQQIGUC>&X#A_?"G#0]^ 4> PNZ53";CSH8AMD_7N_5C MWQ\0K
PII@B4TK!N%(=,6,X@J/0H6"@&1F].-6FS_DUN5O0Q*0?%TX?(<#4H<'J]Z]!=3 ]
PZPK5$>K'RODG5/]W2C#FG7I[ \.K!:EWSXKZF:&5,'II[!G3I%V)9H"$B;?$UR/-
P8NK#:&5BK9%&W=8*ABQ.;:<A0(<ZUJ@-@S<5R?9YGSA/!_;-.D7IH2EARG$FZ4Y;
P\+O*(?\R9OWU">7S0?Z\N'XKB';)3;+*N;V^DJQ5DWA"IP\ANJ(9DFV@CLEAT?"=
P<OGN<MAB+7QOSZ6A.N4G1^X- @C18(T-!X:TRDY(X!DIE*E,7$:U*QE."5">27*Y
P2TO3P.*?W.0H/*^$+O?<UC=+V0C0X30SFBL\)F<.]BX8!KH@P"#EW1>+>?<JX6M6
P%,L!N\H2)TK-C]OO.C"X_J"5OU&47.)$#K3S\P!=N>8&4+!\2)W2/?)8EW2.EZ]V
PI;%0!-%A).3@LC^_G*LM"J9RKB9K76?!4$4(U4OS/)5V\6@P5O0Z<VIR5@0V<A_"
P$!>PJ$36J@VY>Y(6I4]X[;M?_A#@:NAJ]L+FUH7,T4X D&OD/@YW6L_BC<B .X_J
P'BMH%^", PF24X'U%K7G0G"H3>P(RV2_$D$XM?M.+<&0TM2EKN;HW4/Y6XP6^6 P
P*-;EE8)@G_?&AXW\TAZ5GO5T8\5Q&LY:F^O.-J,JIR&2(O>H4"6Q\IV=)_+7S&Y?
PD).G/Q.]HRN@XY#5)'!N"_?U *MZK:6WA;"24'@)7W\%J,\5G)47F<<UH43OO7\C
PG @]"3M$53X^/R?JS@,&?7= A]R&ZL>^/^5,Z8^2!HK]: 9L>?:0*(WP#D0$8(4*
PWYFP):9A):-HI7KDCDP*J%#HFD.+8N_9#[3Q(J@,#77QTL%NJ4ZJ)5W\,6N@66O5
PNS>ZN>T#YP%.4+OI51$)LUDU_'P2P!M')\.BFJX7P<0_&D>)6SZ('%3S7+$:)/Z"
POY-+]7;S644P0/QQ+N[;3_Y^4"&W5Q&8'C"X;MCX_^BJ5$!<#P0!=,> FS_]8Q6F
PM@..:UL^CC..X*&UN@'G9R-(K BIM")EH[J6:,_'7V8H8N%XNG?$/ U=),25Q9'L
PDCRA7H,/!>@L5>75_&TY-N<G43OB<ZY:JF+&;JW9J)W\"(7=*OS\;G)3+>1@<A43
P.1>V?4>#6!(1A0G!Y*_4ZUK :\R[+T*W//$5*9E\&/D=/33^5'GKRPD*%@HNS!OS
P/QTOO+!D:&ZCG]?>1S5M[%7B]F'HI9$="IHP#@"T5*+.MS%Y6;(L4P"@0;UH 8,K
PDR-<,[8:!NHRZA%-HYZ.F$OU;000CC'W]ZD]'UD!GU&1Q(W@84';19T"W4_;_7JP
P[<X<AM=I8.M$JW8D_77,AK*(K68[R<4, AX*#:. I-C68]\-'&(<=VKJBV-Z8E[6
PN25HST30P*65>2*@7K8_]4I90U9^;A*Y.@E_>TJ8\*#CDK?B(77?&N/9OJHL#O.]
PDJC]TBNKGKS]CT8O<P,TPVLX",G=CNF)LQ<P=CBE[I\&D>G(CK4@2^OK- ,;T,8W
PE?)W$+! Y%O@&WI)4F]E+>RY%O][SZ,F064;4/D\/!>Y>KUVD42>(?NGH:?XW203
PYA(31B> "0E2:VWQ!UE1,?4N65GZVO/4Z^:/@&9;J>9) ^\Q+4FV^V(T44N%R)0-
PNE1J*:FSP&TK(/I$^QQSBHZ-L5^/RW@W0^0S+!U5X1[L0[IQF U]FT#\* W<1=9^
P.VCM^=C:^N@0H>X!WH_LTCTQ;6<DF-C^[*CYKZTE>8=X%^2^.O#OU'R:A)P':<8W
P6MF(WJ'82J6]U> /[0O4(TC#FSP,00LZHVDONI;G=1,_H\]R&>-]&;U#(;U!(J.!
P2ZQ;W7%>\4+^/GPH*M.4EYO\).\TW<I9G:S*F8V8_NR.3N;4>+ENZ>9+3>6B0(/4
P-AXDKFVZR&V];<\@2^&2A^UM(XJ^97C*TPHR3^C\$DXA"_^LT]1DP:I ?9H]$$1?
PG9&K#MNE=IY>Y6R5"HP^55;DK!\N3V4QD0AD2#&^9',L*K#N!H+'4DS& 5 VE;W^
P04J7MV)=TE$5EX/;/D/#3065 5)$;>N#N)V9>+'M?7=XN@9&FWU,/5.^CB0D=?2,
PF9&-K2DA:F@H(>WVJ!F2F^+&T>-FY1H^13E1'5ZA-V/K[E"6<TK02'0[06/#(LJ.
PJ(:OY4=?%,6F5Z;4 CA.T2J4%KWC8<[7].P.]EH"^6BE@%<_8VA?CSBXT(?09OV(
P)AB P1M=O+S!X+QL)"GW/[XMRQ)"B%V7=##;L]TJ^S/%U2WMO]_B,;#(F3$V:6B'
P&^ 9X)5."Y97[5W 5B&+*R$7A/NH82KG?;F;<1 ;[5[Y_=2%.;S23ZB)<(=XU7D!
P4P.2DULI57(3\NBR:R[3H"."2[YZ<@Y\*6V*@%^)IU8KP>1&^+ 0E$%5IZ7YJS.&
P#UOM0SERJU[U%R8U8S"5<TKG+75'$N3UWXMBS5:;BBRT39Z,SEH,Y@XJB4U/]Z&!
P_3DEJO2'G8) VN&H>@X*0/Q'M&9*[*X_T@H%V8'5%L,B6)O_DJX\4.TL-CUD0,E^
P5X3Y'5+;#G$U_*TW'<;2:XU<M'[[,K^)$*E%>T[8_3>6?@4A1RI#-4T?48KB?*E[
PS,HF,G/JUAH,KA>4MU&@&P%%SQ.=K(7,=C.T^6R&$.UM=++]"/'U/R(/L1SR4J"R
P!W: %&(*VKOL,5^&J5WC[(^<\>89X%MC^CN:CI+>TP>A!XH95LX<@\M*,2F=&(P#
P:'#?J/Y]@BJCIBOS_E/.Y3)KD];]9)-P-2QYNKF4:CE08%YD-!FB91,HDAZ-7M;(
P:5Q['V5N XL&$%NS/!\'2B##1L"E6STDK!"?S8(*8<XI^Y13PRUSMB0*QGD BSWS
PXN[*AK",\9K6 WL.Q)6\Y(8.N)I=&E]9P 5NXRT:#D 00M<X/MA21N!_(:+ 2%N=
P8-TK4 "4<.\8,)%"\E4"H"LT7<2^\".K#/$J>S,+E: >109!%<+*C0S;O"#+WM=D
PP*)D8EHO_*W[.6[%'P3CGGM1L%&D>JQP*__N[@P0@ &P[1VQRT<T.$U\HYF2(ZMI
P)*2#JF"2GJ'>SK\U/KTI^6E$L]C)HXPCH%^GV[7].IB-"YS%5&/)M9T_+Z"\AVO%
PRZ\[T^,&'F[7]V7&)(OOT?S-]0*SCMD+'JG61E3.OKY<LIO:1:'0Q?;:R4T['R2O
P]5?W%(R754;5!*&F7K0XH)R$KWE<0+[B/R3-YUO3%@*9"KS%L%2TN\-TR:M@==T3
PL%]AE@&A8'0-H'>!PV4"B6-+E41.,8S=>UOO9 @?81\$F@1Q*H/NODM>O]TM1S(T
P?"6K'BBX]#Z(K_GZG5!/\SZ6(\ML(009#@(/GQ.N.NP#$_V;&B/(*H,B3_#Z<WL1
PSHN.PJ,)Z*]T/>,>WLD""RKH=U_FV:W2 OQK/?75CN:MSU<[V)AZ"[7M5_^G$5S<
PT^>$Z;.$W\?'Y<BRQ^(ZM!L1 &;+EU9HJ<Y) B"'?CD,]._&!CT1C,B 8EG,I:K^
P[-9+(*,@NU/*,N4RBW"($$]5>?V.I\6(;GK+(F!Q J**"OMLE- 8%4U9]24Z2191
P=XXZHKHT'[?JLEBD=&R:'MY;(+ZA?\*^5*.ZK 9(:D!NQ'K5=-]-BW%Y0<P!!^O^
P]^DOG6CE)* !?X.U:?+$T#W<+0FBO97"!/R#"P_F1/UIV)A"RCOQI5]^,A?!.HM@
PC>RK?O^%2"LZ?TE\7W!?(Z(NH^P<DS!"R[-N<>:,#HNU<ID-^C,YOS4!F7T[!D7$
P32>]0N_AC->$O5PB(BKF"F>^<866'U2.X5TH AUV+.C-@XP;(AQ -</5.NFI?*XR
PK('MEY7#N82(I#1WEG&3> 5R1V8&' 9&*NCIP+8,6_Y:%"9\8\00>/[>N$SPA-<Q
PK 1P$2C(&J?:KM_#$0F I^BF-!C"2HU7*NZINTND63<?5^Z2N)V"IL1XEAX0VB[=
P/7<,X(06Z#TD@8)'K>4E:WR\#+XYM\7S$(\V?=MFVO-_'7NBR)HRC 5*S\3HV,*L
P""VL%R5HMU&A[)D;,OO3 9NG-2!%;A/P_6OL\/$IQJNURY4A]'QK?XD,8\A[P>?I
P+]PV.-1- RF12')95@J6U&LG_TJ82-P!0CF2+31A$O9I?X8MT>5Y&\W'<[P*& O9
P60'( 1,?#1*O0E:!SFB=,D!,X.[O,NL @8$+-'VE*-Z-"CIFAFE>!,3I*%*U,FN6
P%!7H(X93H5S<I\SB'L5VA#F=F=0+Y5 GJ*DL=$_M6LV[PAGT8<MC/,K4.<J<Q'Z/
P53I .0=!<0LL]IOU/E6F5'1X"M4G/!E7'D$S2ME&[A=?$;D2#C\C18O$"UH>^/@M
P'K')%#.^!PQ4J&OL'%O9;=*9X+L>$XI?@]Q SE"IB#>8<<6U-99DSPNIA^1V/S)0
PQ-US(!T"$S<0,,G@XPPJ?]W9)B#I]*R.]I,:=Q;P\DX!<Q_=9JL&)CNU/A^]*F?(
P4NV9$K6\PKBH/>KMR)3(VQ9NUGJY!EL&=>LSRTL:"PP8BY*M,O](,7HW'>BT/&IS
P":X6,^ISD#1-RE*!_W-XS+1_UHBZ/Z]$/0H*A9Z#>"3(&8;27VQS10 699ID]+"Y
P0-X^P8F>]RL&Y\<?,/PSJ_8I'ZL]&B*BSJGDC4)?;)J$$"WF6%$^;=S1BS#Q 'D,
P'.G[*B-H25'Z?V862O!Q]AFE5<9.W@B:UO7 !+*@DY3Z.Y6\GO&=60#Y16E[Z5&W
P1_:-MB,8B22,B^>WH3H8X\/W->4_.Q11B4&2D(N7Q@AF]_\QY?L?+;]69:/Y6R>P
P^H%2ML.F,%S@]N%'GL\M4&DGFFE^!JOB5-YXJM>"W.9%OOR&HRAU4A@[;O"?N2;S
PC9.,9I0C"LDW-=^[ F88FH^^[]>OC6YT9L1/^(W!P^(ATT859D.=PES]CK>QZP]Z
PY3+9]WN\5>#EEI@@\\G5_HRU08SZ!,49*SU^"]XD"NXH,?RR1=7[Y,9I%5[Q!K^)
P"P 0EOM>OYCD-KBBRSXWSNYCL-0&7_S+6AL7CBS\A914=AK*Q!)C1>5/)J' V>@#
P!*'G["\\P_%:Q3[E/ %TV0DG\ IR6Y,EQ>$FP252;-U^H$"&C]URX ;/"328=PQX
P?^/V*#V?9(;CQ 2+W.3>\JA[S>JN$$6KFL>,%G]B&IK(U"_2$2YW2\$O9,OM;_CX
P&SZ2?]KG@,H6(Y.G8J3[O9FVYBVRH4O"O'8-;!8*\D3#++Q_Z;<?P2EIZOJK6JS/
P)[PD(MF<X.^[912BO;,CO0SE!@V]'DKG(Y]E)1X)(X+M.6%D%%K[&C3QPT_7%2I.
P9NGI3 /0'#W N/W0@#%:;.N2RU+[(LDJ;%1MO0=W4#=*^)L:BG?R ;A[6 D2>PVR
PIR^5F,XO D4 $TW:-T@LI:WIFM2HZ2VQ26K ,)&FS9\[\>$G1B= B1MOQ7ILQAE=
P5U$K^<B.L+Z0$>:[2^'8:-RZ>0AO<^]R>PU*!3NEC)$',$O2,-&A*?+#MJ)S<B1O
P57J9J;CC5TFI11Y#_,4YE.3IW4I9[T:K@&Z*H8ESM<  8#2VE_KN_#[-JCSUW.*3
P'OSV>O%@CIHXZPLH3$V.ZX&/T+]LIS+DPFTBO?W<I9\00T710L+3F'KS*55>[M2!
P8:BU0F[<XX"T_F)OX\O\K=13%OSD@>ZTI 903@I%N38G4^VR92 7Z/Y)9S9\XVK#
P.?6E$"+)<5V"<U^[VR78VG4-/H/)X>M*%WW)@DH/)FO"C#B/GW$B\0D2_K!5B 'B
PX2)$AS*A!"F-G827\3!YTV+=;&N+$T,F+H1@PS3-@21SJ>+4"ZG5E23FFFH5T&0I
P($V\_&TMK?25";<.88=R\&?Z(W4V5#+,5:>&?;MKLJ64+L!PW4;N$&65GI"2>O.@
P<IFJ0]WI?\8^$/5"V?_>@1'3T"<.]3#5!QZ\.,C"Q48HCM:"RSC2>L<P-M[!A3A^
PM\<FFNU- ?9#_K]OG0D-[-Q!D:J,D)&9BTQXN3'%M029%GS2+"\D4X[*$NZ-L>#4
P*VZY)5*/YZP@-F#1FVUD(8# ,K<MC!*JE-75V("Q#3:/[@879/2_?6X2Z!9ZTBPY
PR_>K=#AVW<C?UVF@TUUZ*N868+Y4F ?O\,QQZ"9>Y;;_9=TPFYQA6<2V;%,@4YNP
PK(RTQF0ZG6<R.@\C,)ZL&- R:W".+2UVS\3*FABLF:JV-V5@-;]-2 '\J&#HY0E;
P^DP=9MXOJ 5RD7>0B[2J+M>5%$-0T1870U8V6@:"1ZF.92Y#?:$6X_5+T2$G_D"!
P8%)L;NT XNU^NG_'[!RY\:UT/U/4D7YU)HMFG2>TKPBOBV3C)M<V!N.3L#GL70E%
PP "&(RV?BE&Y^.K63H.BXAVPLC#:+V48E!*+,L9N4,WB(GN\IJR].JSINEA239I[
P]=?QRU7UD%WL\R%$_&Q)O7=4U8S,$&'P2;$M\DVJ2/*E*\*P96S;48]A:(<,BJPO
P,]P,?",ZVV;MKF5615=53Z4V/D#'Y&*:"YG.A+<=9.>UC&B3AB[*Y& U];92I_& 
P7W/=IB:Y\;HFJ4R;45>LL0NN<6OTCF:F5GP_>CK8*<D>:![?U[P>NE$?=M61;,P\
PR0;MYP\FY#R.2&P.;4(PS%G:5"!6TK?@GWON^8'](7  G EC:S^BZO* <^_V9QK0
PS7JX#.+ O O53O] @9((U6<4P\5.*(**(>,2]#L9FJ'!I;S>]+RS8VMR6&:3))SP
P8WS^IOTXU@R-%NFF;J*N%_EAEG?:O)13933[[-MTO#W;@CA>M2/9<?^X<Q]T2Y]"
PP*^YXE[KY\@032+B)4MV8MD'PQ^BGPI_UG<0J@=BL'PG@"Q#5%J9P_(7TM0XK@+"
PH_$^\IZFR9>= ((HQCE4;8<_ORP^ET8Z/QY <I\L9"[DFC[IA)1DO39PA$**.=28
PDGX@;(#L,A-\VOZ[?GI0@(;(ZXKV+(/MKO@(&3A'YW4O&&5@YD\&0W;+KD(JBW'\
P6=F&6V% '^V,?0/H#T'V+4&_>R^V^%+% !NL9+ GGBZ72]#-R9 [-9EBD&HVKEAQ
PFPWI2A8_:8^;D_](\P:&BM?.^R2N?BFA I4WM4T?6WV&' -4BN&//#;<4%*8)7CW
PXW@;1 3J_1FFF*B5*5A84%GNJ+"ZFS6"5=NNYJ8A7T@T.Q[(]VP<;1F0ETOH,D'U
P>UPJN5;Q'M$GM3Z"M+2X9,>=YD[(HA=ENHSJH#FG?_7-NG:'0,K/THATQ]_:BE[Y
PY6!"IPV;@!R/EV922#%LU50ARH3 :"^\G*V7Y5G ,'_6]L (A;).T=(*!N5\D(06
PK>T*;6.9/V7+#M3M#0_"VL_)=N>ABXE)I(8JIF&8[H9)RP /KC(X5@A9-@G02S6"
P:5;XHQN*8&!Z6F?NDU* O:XNJ0>+ZUF"M!A44):C@XZ)F=Z'-<\8:1H@==A*SR$%
P[^:(UAP5"&$45; Z9FZK\,H&09&N5H6D>[>8#N0\X3S+/%Y:PA,*-1H001Q[>+A^
P?_Y=;X&=(C]@$K)U483O/7MYZ.@GQL,1@BR>N?F]YTNUGK$+U-IUCQNJ]U%@PC:D
P\J;..OK<(TNQ%?802D==P_Y5B^_[T]_/$1&AC5)=QU4$H3N!N K;F3*1@3T.$WVA
P8^VXQ!G3^"25+?52K-^!TZ=5O?J4JE*]X;_S7MC3"U.V!'M79#)5\EMG>=:YHYP-
PDFK,+!]28DNZ^HH]C$,13!=<KT]PD_3P]%94[ J5?X:33T*\2AS=^I;.R,$T&X@I
P^YO*487:M'H?A<$,[F?IY)K]5S6+X8#($C'R>=<S.G3SS97M!P9GP'^F)@L*_PK)
PMW>OT@?#@T#<[5%L1U]^(T0'/I>P+[!,*/FEFB#4G_L-YSO_=Z4^);FO0'?H:QI?
P2TJKTBVZO2\[).1 %ATBLX#<A3F1-*#[AYT81\(E:#)14=&,&&K3J]A:TE?7W3I;
PC?U_^T%!\W*;])\@F1A)=3@XJEU/.J8V-\?L@P%R24LXPYOO G.*:9VDLFXYH ';
PLJ<NR0@N=/#.(]U+Y&X1EF_H7T\Z_5OUZHQ8U.%8EWI5$-=5WA*];HOG*OGU'-Z>
P-D)=81^V!="3#?]VPOW3NC;9,"19HP\&R$0(B^4CD*.'CACO5M+W_2VN*45LJ^5"
P@P40UY\<1B21:/G%G>N;0M3"/=)2]R*%S/\-I(!KDW(=,G6%)7>]Q+908X+?%.!Q
P/-6Z?-!+9T#O;;<CQ(=_G&K(:K(C94NC85/T'L)@RVT&YO0GX%)FDT<ZKN]<83;?
P?>AJ,N4N3!\(3%;FQ: [_U%](#C=AQQ[@?A%OR( >_6=PTAV-T8FJ[%]KA@U_S5O
P/DFI-RL4B+H.#?,PF9_PJH%I!<M-EQ.P43'I">QZZTEL":%>HMP(ZQCB\2RDVS.:
PENKY=XN41_\.%_%PNX/^$H\_Z+N.3U<]='[S>VC(+NJ,'^?Y"#&M8GSQ>.P_:09(
P:X-QGL1!R?( C)C26\KB(JY:S 7)O'/J<_44"9GQV>\,0F32IF\-7ZA9>B)GB4BB
P$\*&*DNXO(^ 4K6T:.G\@RC4:5UKN=R/='0-=$WHX<P!*I]I*<KP+;!^45#'80CE
P>"7-'4Z6>W?[]9+?R2?S7:QI-TQJKUFL054"A[EZFU@)<Y$Y_-2\Y'[09V9WO+2_
P ]8_^>/;@XU9RJDPTZ8>Y%R[0-]LRUJ)G858+''6X?JND(HK[LJOOY^Z\&^W.)IV
PU[J?6K(Z[7W6Y(#$>R#_4"+Y@< /?$6.JA2O;[%(LS)N?& N"V'QCH$WRAL:OY=N
PQU=<9HQ(9:!GT$X1@D7?G@AL4V+/)/QN'=9U9D\B"MH<O"4 A&,J%2HGM-0S@=/<
PNA!W.8*EDGSO J!NUCV#R)ZPF"D2+)$F]EG#X4GC,SXFIRH*0:D\+"-MNL;;2T34
P*A"8H7#A5S!K=)!FN;AS4@N-DYC#>(L\GM(]GJ=+ES8Z_;J9:.O$GOIXC',O4(0D
PSE6&Y7>(LS?EAH/*E%"-'[9 +^T&8^+#-0T"=$$O$FE00-)>N:"^YCHT.DCA\B(Q
PV]KJAB\K.5_=PN\S^J,/Q9LH)]B#X92P'OD#T$S[DNV34T&$[54@?3!\&SBX5BY.
P?(Y5T@D:9H.=(03H(2>!>??TNS'AEJ:&70MSN VS%-K'0!G-A?]K;<=2K)EZ<[SN
P4?Y@JC*4]90&H<SD!B"B0RT->9L@^$T6I& UJN';?XYML/5O)(=MJX5)\A5JPO]Z
PK\C"<)WL]V #]*QNFJ9X_/C]#@Z0Y1SCWBO_Y@4E18[IK'ZZM U073+SV:V\4SEJ
P4I9FG]EK %M62&U.')R=4=3.>W>01E)NXS%".%-JCHJ00L'W'458Z;)S&XTI+H\2
PLXU@<*'UTD'N'X-^2JK^9G+%)<X7NFPI6 N"< XZL;KW?C*C0;^#K)G8ZVYI(@N8
P6RU;=.@RH#Q3E*_QJ^3?FHQFUA:W4X$K2V$4@Y)O**_E$\+6Y=RGHY.72X5CGQHG
P^/9*+H5<SH5B!'(9^,$"LD#$FWKBJY6D$[6^[CI2*0TF_I'I'#(*"^OM?@#2:M7(
P\55B36+V^HK0I62=="+K376?\V]3,+%=ZS/6;7=?ZPJ=!Z4G'01S8/FL&P4>. OW
P0 +3>GO$>>(2]*H;E*7<L[EX413=,=9D#QE:W[LJG>:8_&)X%$0F>YG#AL=*8!:5
PZ?6\(6/4R0PBV(*ESU$I2AN/=X%K:9UG!-M24*[73*JSZ<+V2]N%E*M"GM"T_M2F
PU,AZUDP@$7ILG/YDO[.R>>Q0(RW3/L@DXK2[V0UW=8)4A&&N407XVVC>GR#@'G'>
P;G+ XF[C64D0VCJ\5S\<Y(2?S<!?KC1,4<57T5H)Y'R;JB?EP@]WP]2\%/#3=7-<
P&F'I\>6"[=U%QWG@7ELGB=HM%Y?H&-@$8;?:VK_?OG]K&:!RC=^W:3=2F--G,&>*
PN*=<:]5.\1E1()3O\.1O:JI-S]1YRLJ?CL9X(21P%TF/F7G@*!+%JM(B27IST,D4
P5Q?,/GFU=H%%]1/*&;32QGDS<!ZTU>C:V!IO!,\Z0QY)M#%UA#'?);;$N0AFX\(F
P:R9.K(KO%VS<$EL-X<[F2X5U%?-,7]PJF=\B;D#9Z93O(-%"E9.<J>BF:"(>!5!R
PB]P%J\?CN$FULQ.&>3K#HU#<0?W;/9Q;[)'IG_R3\U'J+!QGA*T["6.!-:;WR8-T
P %+$S2AV-+E$_N2J GC1P%5&Y2,3ZXUT$9:G*=")V$T'.U/@BP;8AT<^;G]F&'*B
P@=_Q_[._.*FA!C.$$?[[-84TX!^2LO-H<F5X+ST,:MC!=Q9/"J+9%O+ )/>R%-V$
PX5"#YE(\BIZ?;NV -Z;=D"L;_SZS!79T'=_W^YL?KP2S!^N _04)5Y0;G8C?%&(B
PK%>!%PA\)L?$2QVI0/H;[A]]/!AD1.RG2S$O%Z^?0#IEH$VYCWF(W<(%850K=^-X
P@O$"X81&__8!HZ*W3?A 4E!P7A,9C&C/RI(G,GHXO1Z?RGM68%7GT>'C/U83EU5$
P/'_H- T&QC1J6!8E@;A_0/,W:P<Z_<G-)R64)U?"!60_ERV^FA=!&J8VW!&>X4=#
P<3)A5Y6!2#K@LV5<=U6_\]?2\?)D+"&2_G@Y0 ,6.[:L"C8]&*\Y/;E0/8Q L+CF
PM;K@22),GT:A7D-"/?:-+] WC*>MX!^1K-8%'.&S91X*V<N7V;&/:V6W%B78,-\Z
P].J]W/!I""G;-,T,D7KSG$[>#R3[J<QC+.EQI70@^2H*% " *1,N)2YVK DZUM-H
PCBE1X_:PDRB2\$#-MO%&D"31*K&!1&C#=JMG4;!,/GNDB?(OT&K*EH4>S@^2;;4W
P0$Z<9IX ^IT,H8-Y]Q'0P"/INNM3,L!_:F2$V[%DH]*-!3)'F8*$%@-D/&O;R<UC
PE_UCM6>-U<.%'845F=H8<"2>9PJ^&M-6^7Z3?&*%'WS94EYG=)A*4#R$Q]ONODY 
P5L%*YEE8:I_!JP+"W"_2X\)2:&R/:X=,UN?B%\82Z7H.^K8BXVYD_=&<N@Y&,@)\
P,WP(3W,#;5M>#3ATW49_*@W'OYSF:*S)J#G8P#? XZCPH\5:G^I+FUF=59QT+L=%
P1=TJ8>5']_^:X.@F/U,-Y&(1 F=-F+'$: 6I^C&$[-T(SWR=?#%HK,O@XT>;!IV*
P2 J%^JM;G%6ZPF31:"/8)8]EG']@/ L)[*5DOY4;B!)V?GK)0N%D.K]E_G0YFH"3
P'.57^N4&%X:_)2 ]1],I8K"W <:+&H1\FYGK=47%S V0U.X+2;Z_1!!630V4_N1>
POHL;IQZ! L<%A21%)7?()H+U$2WI^%T4<)#4Z&T+9;;$=*I=73[X6A*YH$-PHA]F
P.<@^95S<DY1)7?/:^F2;(<X* )Z\^OHV>=17FI^+R2T3PJ0#,69XOJ.<580E.-[&
P3>$PQD0O(<Y_@-C:ODTM%J)H8 B8\@#G 1\-YX__]^$@P!P<0!*Q([./=0H"B,*"
PT$WXJ R YW&)5HI\\7T[*TV%A:J88#5QW#HOK/>-6FXR\C"T.SY5+2T,Q$37D#[J
P) ("%,D%.*U_8"B77Y1;O8F4U^)29J3W\+N:JDJ7LO&!,OPLUR!:_W"GE6DUU,]*
PPP'0,TIU?[KB>#*N<L=5A!B%N-FT6%_P%2.D^KQF[<DUPOCP<-(_C<5ZB+0*_"$]
P?&OU1]!^7W39834=U-P?,&FAB:XP/H@CTP.U>=OJ!!;F+W>#3N8 /O &ECW7F"<1
PG+]X\JYA9)OF4,3@3DA$\CMK!9W U!9^[*J1_9E)N:<C'QDJSA[3).+/,UI?-'3M
P7JYU>76<_:I6UY.:,M;*H2I,"<H9O-,B*#P Q* 0"RD5H!^T*+ZB&A,VPZW9$OU=
PC$<3&=XM8+QAIFAZ-+ %7 ]@7[XYU65(0/?+1WAK]EOXJ6</<H51:IMS8ZVNVX9>
P9 'Q74^88]DP7-S*3Q4-%BQ](=YM+-;U42]\"G^8';^@JEA?VK86NQ(P1AUT/O/ 
PBYQ#[&YF^T GO.0@UPIV;!7(L'*Q"(\\!9M**Q4B>[XDZ6PV90'UY+SD95"LFP-?
POUA!FT$D6Q:UO?[H6!2HG64L/C]7RME6Z B"#/J7\(@<96?;=FJM'9 1"-;IXA!2
P8'U<6[3&X(JJ1LG"/01U,NB^^_TC(*%B4A)$OLU]>ZX=>&=:$+&EUYK_4CF&^,BT
P$F32$L"JV_4VMNFILDLH<(-LS^$E<0H'?K\4U]DHTZ.R])#8R"WM[8RY/MMY0P@Y
PU!KS# ;6+=0)_/",7<""IR/TL+/-23DP 5^/B<#BA761_H,@E:?P74NG2\6(LV<2
P9 _0''-L E&X) X\:QKN6<8'Y%DR*G2,^KYR9:3,?8"!L+N.0X=FS2_$/S[,"WU8
P6*RE<'@]OQMQEQ*<&W7I5H"^(>?/QUE]5"RTMO(5C795J#2:HUDA4 YQS]TU@2?Q
P?78<UOBN6FA[$1!'GHS'WE#?!Z+2(X_OUI$8A>&R3JQ0S:#=S4/#]GE/ TO((5D<
P#]1(Q':V:;*JCX0>4Q2ZQ<?P:MPR96[]^FCZ^B4N35\\UL5P7<3@@:ZW@1],\/(7
PB33!9V-N7@RN9//411WV.GI_>EPCDA*9,#4&DTG13V0P!?>K''LNZWSU1KVTNM"8
PX_9]FC&? =UPN"#_V0 0Z<L4_/\_:O&FXA%WPZ]YQHXB"!B,8YF9[G0C:PN[8B"_
PT0IFMKWV3O^.%*O-J1>9X8]X/^5.WC%B#CY'#.6ZL%XXU,I;GK]_ZCGFE6Q5\$"T
P0"\: ]LT1SHBU)0(E(HT@#!(QO?O=_9.-Q^>^BL_W'P/BJ<'S$P *,>SB"O>[&C=
PK+?R/D:0?D\=BZE ER_]:T(G+E>O3.9-W*BFF]K6S<BHHF,>N9"!_OWQ"R LXB'I
P@(-4]*I<"4^*S'$B1G$1+P$([OB>H@] "F[(!RXUL;$\'"RTKNW_\);1]TI_'FI_
P&9X6#^ D"$/%-9>0P%-.(U%BI]]ZN3^%2KEY1XI_N^!$N5PT@R_LL '"]88<S> G
PE@G&KH:>( H+M-)"84Z'B,:,_7/_DUPMK?QZB?^X\>:0')(V["!RVD,XOZ'U2DO^
P2H_UR]9$;U<(+0WL,'3OLG+P/)&GT4F:DD_Z5O0)4/8PC<U^A45)M6AS%C^XQ2JV
P#"TBX5J9FTS,GX[IW:^A?VP'*;V-F]"@L23DP;#:!A"B+_57:NU%2>_#,**.FYL1
P*X^.VR:+20"L/+KI"O2E\%3#AXF/O"34V_"GKIG.=[<KY/-4P)%XGCOB*-URD/9Z
PRVN,C123"^1%&$I^EFD_UDF1X>WY-FR1R?3[BU,G(6W4ZZMI'1A?(4RV9XYC$<7/
P;T2A;FC+^'N N\KBCBV\&FZ)'C6?T/8"52'T0PF7E_5QKH0=)/*M"/<UN5M-[R8J
PH0AKX%/Z(4=M%1\3G+<I-XZM^O%RS4.!<DF^\F]VJ^K@,]512%NP+338*S5WFF!R
P>EMKHR;FM=8CQH4CV(L5?U;/S+==<=&P'))9),*HHC(<DY#JIZ__DB(S_T?4  \+
P!OXY:5A)1[IX:;8V.YP>YE2#4X?^TV@(O"N<[4E(410'OJ4ZE)#!^^4[SF38WS'[
P0B:CN&3/4X%)+EFJX)'03B)PRG)_ND:;L[>(J#!6A =,?9N'IE3Q>9E#K&]-?]@_
P+73STFHC)U1OI#AN=\U3S_@,:QWB( &-QA[>S> 94')$;)*I8(>I6@2K@O>_8HFW
PLT72?@"V\IU-HFJ7>Z)B-/*T >N<E%0U=N4@TS2#M<0ZM"<V+-FO=?E%C:6\N;9'
P3HG"_OWOAA0+O_ QL2[>YJ8B!1HN0JY61RPI/!"+$ON]G+\@JYTM<C.<41S-_0&K
P-UUA"F]:AMGH+_C>XQQ70'\:0,U&[M'\@2YZF #T1F7ZA=%)Z,.--8H2AQ_*BM%\
P!4@^JJ@8X2BE.)J@<X/)M&'=5YH<B_2" A.(],<(6M\:WL$#DS^XZ&_AII@/B4#!
PRD6CTN!?2,JW+M(@_$F<Z(UK;)M#*I?W!!4]RU$3ZJZVK'#1("_Q<A(0(.HC.!$0
PN$XY$F2@+\&'VN.1VW\2]C6];Y?[DNC^X'H&?]7T<M5$'1AFZKIQAI_P+#I;OG1X
PL0P;Z8/NU"F+@P7T2^ 8-'%L^IY4%/\DVW9=F(O)@/ZE]%#3L?.#2TY/<I7, WJG
P"6J*4E)=J3M[:.I"M80AIEOB$;GS9[ #4[?FG2**==FR_>+1Y#>ZH7?LLI3KS2_$
P7<C*$1V@]PKQAQ:)B\"!"\G4K,0T"$!&B, 0ODZ 9 %N^]?R=M +-W Q#R?PKHF&
P4;JSXS>T!]=TK2.9!?^\S"1'>]2Y4B-_Y1UH8_;;UZ #06^!M/<51Q-OCE'BV@,Q
P;49^8E?W3E*/#Y$8!!-;"$IH2Y"#G>\#0;B]J3!U2W6+46-WCVC$=$G+\^MF@5 0
P0D]-:Y0 &R\GZTMC4*J=#V7XFT@[G%N^SLSO\0B824S^6^WE]W1&\NEY>V<W62I=
P9E&X!=,NY(QUILQ/&?+Q7AXP['_9)ED%$+?O"%ZPKWCMH)#8*=_I$F* YL??),H3
P6:MUCL':<%_F7Z9O^[\_#0VEOE-NT/SP<17)^B9TPW,XUN6:S.BRM^S0%-BSK2E 
PMW!]-J&.(?>3R$XKCPF?V-WVC* T3"O5'@K/M<,#'IB"!.6"H6^<M2@V,;3Y"H22
PQ4$4<ZOV9+0%WD=[[[1Z@WO\C/"E)"5SO9*NF.Q>[3!K^7>KGE)U+2)= 8_0)) Q
PM$D1QIYPRS$VXEYQ2.Y5#3WCG[UYQ<:&M88-4&N*J=R1WU6YWU.3W,IHEOCIT&X,
PG4$@XX(,?[?KT8 )(7!W^S?!SZH JN--)GZF/8*4GVA%7O/.D.27W96KVA\V"!F+
P(,UL*V.'P;2?RRV,?3<&I@/WNCX;;CK7A*R_H6? !AQ"4N^%JO-_^0ZKI, ^CAUO
PTY[O4I8%_JQQJBU^Y0.'3^*&!+5,^#QPOEOOVUQN-H$4.R-S?:'ES0*="4PPF3_=
PNXF85'U^:,C>P/D++MYD+R.%^2(6!;I0!#/74MG,3E% +GF@T24"4*R:>V\03-/7
P11PS&0#/Q91)9,Q&7TDW;&@A^_3-T1=&\X;UU<K3\T\ +$E=]B0DQ$$G/%_%(Z$S
P!JA? ]>E+EOV3\M+.B>SB]$#;*EO3WF/38%1HL83MQ"'!&U!( CS=[L537;Z2+J%
PB:^+1G*UP%X"GH<3"&_);4W&>C''$:Z'Z]-FFV"C8L.P/0\P_,[]CLO?'<1AH=$E
PALH0O#987\Y'3K$^,8YYZ^NQ24_$L67X61Z*H%G>%ZJL&6*BF/9D5QR:&5ZDQ&_+
P7D+1]K]D=H)=V:88*6^MK1(C:?A="P&US]*=PZ*^>Z^V,F!:HDM)1V>XL/=('O9G
PD4 =,7\LOG,8N'K8O]6J<9@!)[$QF_7AZ+$6KU,JJR:\KF!-57HY7X.+?YNS!XSY
P)/YK/SM<*C]9*&6_NITP<)^#:KJ%A]+=!#)_4I)XX3W':V>Z@^0@/85!M'NL*-=R
P1,)K']QLSX:5[[&T!E/ID^00A9G4J'MQZ#2!)?ZFV(9WUR?K7<JN'$=I!EV3F[S2
P^=>:'5C-U!ULA@3NOF&B=H.=><Z*;59+14N20R IKD0'3%)1),^VPS#6.F]O7O0(
P@8HB! &)F /I:C/FF;UDE/E+,("R>G4P7=;C;PCB,*D]/U;(NL,GEY6EF%W3_M2\
P%#\3JXJ/-)F3X2[SZ'P-KY@D+ZSX0T3!QG:XN 2"*NP*PR<36!N T5,;DLDW'E'_
P 4S@LT]@Q'A:+D)*5L(9' [KJ+=D+=NJO= 09_?O:K3GC&HL@ S1YAS,C*97A&$-
P:Z&-WO/3.=4%.H(%0:UM^!.!F?+7J<$O>&XM@NR499AMU]?!WB=X1S^7X]TT0*<1
P)'TX,YN:) UAVO(M@, [EY9\25M738+<Z:$65,-JU5EHABWT<1 BY!Z 4!1)[X:X
PYL&73%&SH8G6/)-^6.R25V,4Y\':/QENRQ@:!11ANU_P/TBU5M%(BX)(TL[VU F/
P@95#MQK UGVE1VK_([N<_P[RR0AECGW3)2*L"A>70K:VB@D1LU^29K-1QI83[E1C
PF6D4G23A 6_ )F/9MQA=5R%W+9[W]?_9+)M7J:'3#6\C^C7)E:]^OHA]'O(0 7G-
P(<LX)U0,@\ETY#(V@%OXJA%%78 =5*IB\V?5*/OJP8Z00$'TKP+C_]*1'7CO87A!
PYHQ$O::VR<O%57XD^"W9./L;\Z9=3 )H=MKNY&RDO;^YSZF95D-L$2!-$X,!F>C$
P]_4C3@J>]\-::<SS'7EQB)S/ 0_15&:I>*97HT'V@$Y-5("^$VZ<4L)V9\H @(&-
PL#HZ\[6ST4WR6'>47V4U?@%PQ9>P^]Y<&3QG)0&DSD0HQ"10J09+M65==.P/;(*^
P"U#4>_%JJTF>2H_C0=Z+E/0C+Z>S^BS:HNY-.KN,,SD"=7A#1YU[-@JUI^TT86;Q
P>RB/ N"@[$J%G)+'Y:R&DGI+@3G_\&:"BS%I_U)IZ%75#*[6T4;<N(^G?#]]*%V;
P/3<J7)I%;1=$R8;B U'CDRO_7,22B=%?-2=EA6/X7O:1\A_A6D1_ ]W%[5YF8P0F
P-#?=GP.3R\^)EMVSW50G-1)>@A*,-==.A1GE?[S^?:$[B3+.Y;Z;Q-#YX8!54*,8
P C!$)NOY-J>)]8)_C/'ZD4!MX , /);2X'*@3[88Q7+>B2Z04Z_T:)*U 82ZQAG3
PQ;'Z0 CQ54'\^FZ6GA>1A&A))7_%R(\.U3TTCD2?3O>,\ 747<+]189:DBBV&/*B
P56>"RQ4WY_[0%4O^RQF7;0^2<-."!_&WDIRH6P*=J?VLDJBT/C%;NB?6WE$6KJEJ
P)13!1!LU$7; HVVW%D^GK<=O"B2*5I1J:E]08'U;EY\])$<3!CE \Z\X8K1PY?M.
P-M.W)4%F%.$L;G& 7/VKKXV89A '>I4^#BV5YIU!XK>76MZ6>Z8)\[<-WRA74/7;
PF@_?E=R'6(WTS_7.8;XO! 09@+_(8.T]/I65;D5O5.7!V$^O6,9@=W-J:"P&W)-(
P%FOAJZ</>H^^ $3#/OJ?@86N%GYGY@P7$SAIMART/&8<-D=^'LT!C$*YPQ=*"UO7
PZ"E*V''4;<'_W#P\+L,363Q"3W+5[67)"30N#]37DWIZP+9!;AB[FL+%Q&(V4HC[
PX67800Z!@U@8#V24[;6=JO2XS$,PS#?=[^@/;%]Z,F[,EP%D]7N+45"?0Y'0+*Y 
P))M_8D;([;K-OW#HX4IX2V0JX7NH7US'%W_"H$1RJBTU&Q?#O0D @SS!;B=C#N%I
P;;1X-"#QQ1S,C:&#_&I+Z.HL[P+N?/B1:D*612Z)70".:2;0F+"2\<T)$R JNP0P
PF$#<P,3BRQX(ZYE$8A.$>R[XIXJZTFFWFYRO*-4>#@F<6[IT^2[\URE.XYXGF!H?
PXE!%_9C\-" ?:NQ  PX>#7Q;57CD:"P2SP2;MD:/\(C*W[B6>"4H)0&5PG!12W5E
P1-D,7HXA.?PDC5[,S[D'P-\5ALE!K1HMWZ0]FNOR#QX+[5%K!PU^'3^Z:E_]N\&&
PY\E+4CT3S"3;W]8K_AN&EC<UJZ?4H8_X$"-!5)$!*^9-(=B2C$&R,6B,DOYWQC2,
P9(GVVJLO5>C558>%E;SK9K[)':[?4!!*"=4:VF1H7&KOX![('ZI['Q=>4))OXZ8:
P+T>W'XS+[9FH6;:L[1.;3"^_?2Q-:Q(N?$?:;$'N^M?YT9*MC(%9<"61U#0S/:EA
P4RT;,KF6&22#)PVT.P$XW!BBD ?OMO'-+,QU:8N==)>IL/1N?NJ(7[,IA<G]'<U1
PA&*DY)Y;9'W/?H^M7HS*$^29<)1)C3!Z2OKCP=7"%BP"GFS;+>X, VM<V/S)BAE@
P(A*J-UUI2ED7RQSXN)*\\D >,>S=1YF..C2!9+T$=XZL2=7.K)X2CE\H"@CL'%7]
PW:_5TQ[0N!39F^H5D16QG%U]*2607DI[M$,/<]Z.NB@J0\04 Y*I3 P3J&3[)Y5Q
P[5/?+)"AKJ\4\6[QP+/;J>KG>!G8N%GX^!!/&*X3A"4;-J#L]K_VL;%9F4L#="T)
PAU05]5]PP-<0<;F[+D%GG]K2;\.6%3?<TNT33^;3_YE$S)QVW6#Y21*"I$ANQBV7
P;622.Z;;/Q [*Q#0''F#JKP.(H1=].H>VLH)^1K&E_2D$@84PC/ /*GEJ9/*S+[6
P6)$_\)*9!WM[SV8>%4O^RC+J1]N<JV&.QJ_AQJK>1%XF!CRX][TS)I]VT2X2<D_@
PD?(*K+\,&R5R@[\OPB;3[SQDC%UPSC"]GA"E6?I)-.@R[QPN,/_'VG(//VV]6<T'
P@Z3F%(%",X+A#G[25GXZ+>%F*=!>G_.O21ZY4#UA$E3Y/J_SH<M<UB+G0J FC0'T
P_;RP_.K(Y;+=.^[4TQPH,3B+!.Y?%4L)9"?\5=<L" Z6GX;U>FVL^XJ60/SV1!+:
P-_/V20KO[=!YP7>98B[WM?Y!3= 65G,<86O8]]5*DZEZ%X42UZ+E;TIRYWO-24H<
P)./@[MZ*RJ@B'FZG]Y2BFV[HEX6ORH<8K/U!WI,J8]!R,B_QXU\P=&')-='WLN:B
P*-$R+_$L/J86&<DE+WC&U(_(V6HQA8F W':W%*U<#%&/><KZBP\5QT3EPX746U!^
P;.3-E?"^_H%L5N#E@@<5K>X52ZP,=]]?AS9:QU'6MS"9NKK\<JRN3*Q8&-;^DBPC
PRZC8@ %W3L2KQZN4H3"1Y"C/-R&&3_N1:.)3O*58%(4I$LAL?3<J!(SG<XJ6%Q3T
P*C6!^GU*1RR%"78R/0Q_&SZCHI\B_4TDA.8W*;:4?SRM+\?[AO&%Q9^3^RD]+!.%
PY%XAGIRV0@QN;JOU::_R%KD+9>ZM&&AJL0PBW6#IZD52QD 8+_PR[)T '\K"H$):
P_I\XY5&F[R,H% F(2('C=5'1FKBC8LK<<BQV9GO^J=3H=CDH.R^BF_'/WX7TH4:#
P2W)'ISF[PG2>FM.1U;/QID/RRDF'HF+6_T1K1:K9T61YP-G:^QN7/,_7J1EF U?K
P5/\*L@3#"_+!$KG#0YY*#+Q?V<#WI KO#/;$_/'B$$C;8!^6-L6BNM0Q^^N[;>F]
PC0)=07PR?T2^E.H;=,*[VZDM]>,<\EB%:L).!>1V#W-MFYM>MX%!K8]B(TK:W&KQ
P,B]7SY<U)BN78;Q97YA,FU(BU@ZI:'/%G8=J&K#2WX/MU03+C8051$<( [YH9*6N
PAVA5E%5!$ ?JV\$^34-LB4:'^3-9)%<")X412Q\<6\I2N\U]?)-HC&-O TC<(]+)
P03"<]RH^JKM>TP+:N2)7IK2]FX_JX#ZT8,'\\<^FW3'4NHI;FTV*Y *0^I";J,$F
P1UHCO"$(%"7:M:T_B;5'WS$>)_? 1#NJH&MIF)LWF#@Z0*!5"8ZE"^C<V, TQPT.
PMH8&S.8C1H^U*L2/HX-M<7-.HJ1M1A1FS6F\MK!Q8&7O'FEX6A&]>)VS:;T!:R^-
PJ"=_VNFLBRRNZXFBA3J<@$$NK$C8=)U64M.=LC Y.1E[[&;3$"C/1K>W,0/D/DD=
PA@-NU2.8RW4V,# D%'CW_3LCM(.7E2UYD@HB0LYXT4'R*5:J5@D@U?,J&LI+MQ6J
PO5#HI:[.YH%K!81FT+B+#-)$KD/[=(<Q85)^="X'Y>&$NB])A&P?VDM@!$>B0*H<
PG_1Y$T(,\DWHE<W2,_ICUTD93G;8P4L&*7_,5M 'U'8._\>5[@;%A9P;5J*Z2[JT
PMO.%"%RP[%^@\N? =\L\7_/6.K7K#&#N(GW4HUY*""B+5>43J@2QOV4BJMA!C@<[
P30!>[\.<Y4EQ[B^3QW!38S<Y32L G=PDF[1;>V5D?U!=K,F&(BQTL]?-#ZG2S4CD
P.&*.L+&'S:O.G$3T#UM..%S\>7MNQUZM2H.@H:T>0L#N>\H;"K8()'W-2;QKNB')
P*_=(/3W'%0#(=4/=A-T3T/4UV:F4D^NVVWF4J"UW)K\HC5"8EOJ%K>.M<HA#3_.5
PY2!.J9BV*8&*U;HH+=Z^@5C'$%K^.SC?/]3\V27M$H*K'VDF!M0%5Z-0"XS)2<(G
PGM(PBAQVN99_AQZTGHVOH: U3S8\OK[H*Z("TSK@CODU\Y3+,QFM31<4E16 M6,(
P8;OMSD/<WAW3Z09Q;XC\PLC\V>/=8$%$.$]F>\]=POEI-WVK %3 ;2;_ X:P\Z^S
PM5S6]VN3<.3QL F 5_T0=/ HC*-DEI?#L8T5"BR83D(/.?)2%GPN.'MKAG(P.EJ;
P[_^0-HH;HH#27S:9'K\TVBTT72:C1X="A2& 8D;J:Z(^>[4XOZ0[CI1<T/$4DLK$
P.2<)ST34TF"M*]+6FFPNNI9! 4&= J>T8WT[& UG\J+A* %-6R([KF&/&(].%'0L
P:.Y?7#OY'BI29<7>4:-;M_2CB/2--%_$@#R86<OTX@G&[G"[I_)2^=-J33@S$])/
PM7$X4**^;<YL)@BC1?JBYIFZ85_PZ[V@U4;(ITBK-S=1RS(_Q+]/?[9-#6NKV?V<
P7>JC7&I6?I[]??&V46[X$Z-@Y2"_S75%F&5MF<KB5:@#*"@,(D*#5>H!YI A25+X
P06F/4VM+_17\".F2M364W(CZ%IK&/"N2L4 N5_Q*71-L;P=KVMRY*7--J-CT6%R*
PXOTMVP\W.(I#[V=NF^11P;%LZ<RTL3+2^0T^J54$"U65_P%MP]E;ZXGZ>SJT-J7U
PYY^.H#D8&) >PTQ\!\G4^ZONGGT162\&97TR/&[ISQ>A]/L,T-CM*=AW;"#\KXC\
PL]NT-WHAJ-L?JY= /4@'.6MN(=XTZH">88"6XB9@SF>DR,\E:'E&Z.Z8M&%,N#H"
PYOKS4&:I?>[!Y=X52BV-YTI@,&BL\AK').]&&B:HNPY%@-N)0"5<F8%]#46A]7@U
P7AJ.49?C<I\4W2GF$<)(5*0<3PV!4!+8++Y1KN?'*'2IA99 :/C'_V5,D.RJ*"BL
P_^K0,G$823((F_3V2\("4VYH!@?CDNZ(MM#Z?*#6<;ICU<E?*BU<'.QQ@.OL&B;;
PC>?)NXJEW4V3RJR:*O#YI9?('D1CXBJ_;)0$)IOD0#(XQ&&>E)FPI)XL!\:9\#[ 
P&?CD&05L'Y3&=#2LCQT>%O/A2\O=$)Q&E;;A'F.:NKN$6YS-\3[+ ^[2RE9DF\G$
PHC$7IIEKZ2U6F6X:D88Z%&K<G53UA=^9 1;T8C?"4,?8H_SL2DL-UO9'I_.?((=(
P$3YP=IAML5\P R8A81T"Y+Q2V(($ A"ESSF5 OXJ-'MTT=AQ&_1305.E=-5%]<K<
PP1]VR&006I*Z654!/Z\FN(^MW7J%,GK_+X*!_!M2W8BW>V^;"31V:Q7#"UY4J,"E
PQ<#R&NR5CRCOZ4Y5 N&5\@12)3#FZP*,$, ;QFD=+NBX>B9]75G0)67.I6#YI+%"
PQOB;X=RN%A:S"Q93]W%7GG7Q#/OG^80K:?;L7\:9MU4G@6;,\-D=L[HQQ<< BHZ[
PDG=4JK1*S("Z*6^ 8AVQ]QG<%M!IN<3<R@G%^]S(292[P$H=W'._5@Z*12$=X"[Z
PBG_I .>R[(PIH "B<"(.DI"*J7UFY*/]<O,_,!)T0I3HTK$XFYRW@>(C?3 B["#:
P:$^79AGW<3&:QB-YPZ55(.W_8X"Y@!W\1,*#X'1,&%ANEU8^87&]+/@V=!*] ]^:
PH9/O>=F>)GP\A*+&R@NFM\KS&0_SZ-W_QHI5(8(./'!(0.DX>J-S9YQ,B:)6(V4G
P)> P!I,\\!2EM#%PY:P"Z7A)KC)U#FF^Z/1C=4!\(!Q2.JA#-;R&WF)DXK9GN?2"
P(FMZHGFK6!ZI..Q1>H],9SGO%E^-0LFB53:\S-O[Q"HKU]8$LPZ#H,41,@ICD1/2
P@_[&%0F>2H*2!8I1UP?UX\IW5L@S_&8YX%Z5UC; =+0HI'6$/E.^AZ!=#!<KJL4S
PD+;MD+R>"CU_:'XOSMO'K9[Q(KW8HX!CE[F@F:VE3C.*86@$N;(D8P8*@6MB]:9>
P'BO;B>R-8HN94L+*M.-:@R"=/QP,MPD%36*4A(P9<9K/$W$O&=3%%T;UIP',KQ3'
P%V),F)KH:<KTB:TA9I(24$%#7Z*-76BY$$I,Z1ST8N$>2)Q2:#]I_+\8\CY5<F5;
PYJI',++1UA E2RU&]9I3D"C0=KS&,VL$I(DH@^L,4?PV9[]%=3)^VKD!F7I*/**@
PNO()NEF\;K]3,1XEB164#.SU:]%G%"*0E"R)NYE@\LA0K!Y75Y?Y/&%W* )8( N?
PH,/UU"FD&E8YXAX(IY>@$SS@=]@.VC?!\_>.<P>5CREXQKQBYRH2%\ND%NB;\5DU
P13W5.K=Z,^<.6N,NL$L0;?R@FP2.Z)1R0 VY[ML]*__'JAJD_48-TG H=;K9W&'T
P<)ON">*96V#CB1455C1>^RH PSD4+1%U.A*;<R!FFO-D[2\/7D1<S*1M>6,46#I)
P3.HP@YC)^HFR5'1A_:L-LEC\7WV9/V(7)J"-I-A^H-/^1-!O8*]6D/L,X./^H07@
P-![E+KG0T-%#-Y8*XAOU"^L%_1*)C3"ZI5U4'LG%;Y5H@$[01_9T--FXG"#*4GP;
P B)Q(*5!NQ"096Z,:Q+#<0L;L[PLHZG;?70)%NB>$3&CS(9"^$BA1?/ \@FD8W[(
P8H(8T]+8<E60>)A\&J@&S:Z0U,C=(,&+:)!Z LCYS8/C_)"YY"!W.I%/,\JZY$2?
PG.+SLD1;E9CG=*W6]PC^)D/_,<&6^5-O#DNC?V5&;*\8LAR# +?W*<=)!4$@Z]:&
P[_Z?+XC[0K*#?KHYCO/>A#Z%R#E(6NJ3"6(&8>7]5D(W(E/U4W<]?YN#0@(JMW)&
PG/#X"5OR#UU+YJ^-WD<,':N(<(+Y]^I>QIX$?5[P6";-!AZ/..VA[<^7+RB&I\WN
P6G9IN"(FV%\]F]S*T$U% %-)S1392M<V3<$^/@@.%KA7].%U1[:,GP O0)F7Q5[V
P>>5IHE,]JBB),@BN- V0+)SG_JLHK(6^E.R]*-XF]K8*5Y1:! ^3?S4!$ VNA+XN
P/NHV3KC7X2D6I=*$"WO'<7%"!<>OFOB#WQU/+-NVE5C^I:A?$!&>^U=O6]QUV5H=
PWY]%?YIO!I]:Q3!XHS^NKR%,4H1B/M&/;RAA/2;8="0LKL @+4Q%\WTD*(O[REE:
PD>HUTO4 7X6!OL1:.#6)[7?(BYF42*O 5FN7('LGG"I@4.[CV4>O,-<H8Q>)>;4:
PAF2OH^PW7:BS0/?!2=9/#H&G#/=!#D#W9+7UY(*3(TG/@B@6A3%=?[9\.?,LW>W)
P0^H-\GV\[Q/*+7??-S=I_2GASS<[A>4:1YL+='=/;H/%ZLCWCF9<?+IM8\T-J@<?
P,<VUL04P2T_4'6&O.<)6@-+X1F]N;U-EMEJ*K3IF(3D)XI-C=6F6.C5GR]^QR;2U
PKU$1E[LP#4@%&C3\J-2'BN377VK):UCS\.YX-@Z!ZD*A>)+R%8&/( JJ/RD64'+ 
PLO>TMO.?';V0/7_:8/Y.AU>4E6LO=5[F#ZD*F%&9YIL/??U+;1Y]^QS*:04?61=C
P1W,P8%_ !.K)Q%,0K1<3@A.#6H-"M3% %.3ZR1VG^D)C?4XO@73%99G!-]L8C#*B
PW>Z4?T\($J!1_=(*M(ZDCM(L/U1_^O,HYD%"22N< M%/-11[KEU\>MNS),A3L[^Z
P/T'^5YOI5@[+RF&U:<W3@=? 1$IS*:JK$ME^]^LNO)K>U_SB=]EPNUXI?I -QU0,
P[#E7PA70:Z?WFUGKR(HRO\6QGV1-7.0G ZDNC1R<MCYE[J*Q/SY9(W'1S4PU5\3(
PNB=.]<$BQJ8NU9TL^WZ8DOZ4TI&R+UEY:D;Z]5!KV%0:81Z43)D\$L_<2'G#.^7U
PBJ"/LW#2:MQ\:+.U0DL?1A^3RZ,XSWOSM<O.*N9#L9?C2!VT#I4[67%'FW1-]O$4
P#^ON%%MJW$)P_8 ;WR=Q?-MBXTS%(%K0'U^' ]\0!=Q!"QR7P'V=MUK \LXR]"]/
P"DWZ42?3Y;KP80RAOXQ8H'%3QGGWBCNT$;R-O"X&8?P$6^JB(H(7Q]773LW<B(YF
P=S +H=JY)ZYODEM/<&[?3]((KG!<X3",H>T@;(E!TUL"^4_):07 R,16@!R1Z%WC
PICNSFZ=-@3I9&T0L3>WQ9]IC&TKL= )7ZM\$PI$Z0;P\RBPK4N!DMRE&$\5FKE>?
P)LQ:_EYZIBO:.U_G,]AP+4WL?=IT32)F^<)_X+F,,K<MS =BZCC@M]6H0C_QB]*O
PGF+]'+>I*8H(FZ$/Q_> 9YS>\" /,8HKAL=DY#/\!F<6K>XG2]8>2-NR/T':%$ C
P><2+G08\HR AP='B:!NV132L^$LN>OF.!5E$27SS#4 &IZ_I3&W3XOAWU/Z6)Y?V
P(1T$*VK._"R"B+BKB-85&=T79&2C8];?Q>BSSO36CB1 ,%E2.89,Y9<X'7=VQ:2V
P/*^FM(@_+,LO9]3&YRO8273#MSB[(SXW(TL8C1KNZ160$35HY*QN,4YGW\4>OOZ\
P0#D>+HV6U\<!+R"364(664RB)-]#I'K<^?1.ZX75'R-!>(#Y@/_'*],-%VY#3S7\
PE8U,ZA:@+P:6MVM00=8:%+OM)9SR*B]:1MSU]LVU-NDAE_D36LS<+8XXUH]'2[PL
PX2\Z1;-P T#DW]V3?/FJ1:SA?OWA#:_%6'"J5[R.]GZ#Y:ET?LY_,)I@I\9@WYVK
POJSEW1*_N\T RRJ2CXA%=1FEB-(T #SP+AJ*W4NHJZQ#&,O$^&1_VD8N;2+X GKX
P-@28S[CZTT\NQ&NB$(]"*Y3O8'?8(D N@=F[DYR_=6+K-'1$!L\;J(,I90FR!M;^
P'\E"5MGRK:Q"@W$AD1&V,47.^U+>-1?$#LNFR2_QW;T/%B9BSEZ:*>DG?,PP4]VR
PHW*%^&\%]%=OX?>Q)67)ITO\X>Y4)REX$1EXEIYG/%^B>O:RSU)SE5F#P6;QG#7(
PDI_X=5=ZK:\29R*+?.['V*E%YI!->'D7%JX0S#U1_J]IWFFZW2 ;SPV5'BF+<<8!
PV&1-K&TB1*8$NWWP27XH_&II[E=O,50A$"/K$-\[@L(*I;\<P6_!"1M^$6=UBC$F
PC!O]\5]G(B$_D4"!71D?$^J2X45: /X-@>P;MQ$E)"*8,B_0>D>.[7(^P2)RO@GV
P $"@K1GZ= !]8R,O?)U?W:##EXJHB0]>N:\M3K?HF#3<U61">UCWY$,:4\PD+1?O
P+812076H7^=X&5':3,+^JIUVU,-,:P_+H[QRE7C U-KK;IBGU^<==Z1^^- 0Q4H-
P/C6IQJ=@R+:*BL:6!;F7A<FJD,#MR/OJX6J]?B>C(;^ZJ'W\?#0PLP2^O*Y8/I@4
P$8ZNB6S7L.MH"H2OW>._V<:)SU"B 6F'!U(*ME"0I<PL)>*='- ^9BQMWLG!QYQO
P=LS>2)+7&,,Q*C6Q1%=\=AF@G.OAZGD8(/),8[@N0L+_B-!/0XG?Y4KYI*M667(!
PGNNJDNAN04?G>5<98X>WW4I3-H+GY@!%BSTZ"Y*>)_(YP@JL#_GTN']H4FY0"-Z!
PL?P[:.D/X-N=S*I<-,N ^]@V;_%T<]S$7A7C!SK< =?RS""<SJZ ,*F4*.JEQ(T)
P]8*C:J=[WV:E_/=UQY_EK+WYFFY$^HR&]8T"-0 V,7=QCYT VKYD+DR6>'DNB:8W
PI<)G%'IQ(-U1I&*_:8!FO?5S;SC==+A8&&-242=,;BT^(9)P-,6R5>>@-$Z_S1U?
P&CW@%^E[.)A 7/>SDN=-!"^<_IVYUTP#KP IW;,9;K50_Q!6%G<DN&VBQ#%#E-FR
P#<L*+6@/D=WX!<2SLTZ?]2TL=GY@S&PT5FAA?ZTS^[%K.YJ6[L_.AC8>#G]2 :ON
P5[KYS51".PZ+,5-.C!0^/P@ZR^NBP*_8\F,+"7F0&=@._,/,Y/*9J"#-K(&[1S0!
PJ_*AB\\2\&_&S(+7Q^/H00:/5U:.$LAN$PWIA#6Y[6P5 9)3':59S4$B?Q_6<G*&
P@ UM*T@E6U8)^L#0IX5LH8$WYV7]%3\M VY,501^AV.(,(E72/+M.UIG6RC?-D[[
PSAI&VKR>DB<!B9<+^CH 'YQ$R3RB0%GW\)+_*MXYLU'("H8]RQ,B*4\-:/6230QG
P!;<!DEQ >9J8FJ&5#*U216Q?_]@I?3H>83^UN<2N1,$)7C@R]JY&;;3,N#$W=+^2
PLE^OGZS.TCO[2UB,\F1@;Z)B\'50W(MD6=,;]]O#O#?K7923[WJ)987!N(N,V%4%
P2<P?COGY-F'C9 XK@4^$#=6$^#J9M4RIP>L:'8/NUGP2.[ %++)O4D'_]VUX62,'
PD*@4MC6F+#OE)=TX;#YZ\4_FF?R?H'O<=$/N=6TA\@,TC7^N/4[7HY?A@X3"2VX?
P2K[@+8V>1VBSWE_1L-)K/!O,\4I*ZJ=:,9>+]/R"/\PIWN+KZ#%_;ULM6/8A*2B3
P[=Z]#75YL.&06^RP!^;7C^=<U3)XIMT%NH73))2"\-HOW2,N7SF?''6#'(CGDN5F
P'<JZ3?8*^:BLNC"3Y"Q2=LY+?52?Z-[VD+M45 8:+6T>1#6,B4F^!G;#[LCG]QS3
P_Y%G8-Y;/#7"@TGD(N?$QY&U+\EN%)Y5%&Y5[\EY1NTEBP%U]<3#F/Y,<?,F;;';
PHL&S G9E#)0-=R"BWC"[&749]Y*)Y\A]^2\++63<]#MG55=1@EG4;.")JM*JTVAF
P<0=@:>^SCM4!.,4BQY$WSDNOJ7PQA<"5E3YIEI<!PZDZR+?/E#I90IUA ,9JGGF,
PO7J0>@%SX%].=<FHD4@T)?#%"N0)<.G9_T&C'U8X;WY%^)@@E,></,N'=]<_ K G
PJP3=F]VUK%QEKA. "0NGJ&(TZY?X=3W6T->OA&F'.F8:9/N@+'(^R-7J&(\_:OW%
P"E>-V$E=#7K:OGOQF\4_RN(0RN5DTZ9=).A)%'OLX=[ %F;)TRMXMQ/RVMU^2>M3
P@3HC#E[>.9,7*&#_[&D:.")8+]:#^"C0]T_ 2KBRC6:L+VY[=76Q_5Z+RG>H([<C
PM*\I *)/O53T4LF;RG\J F84RI,O^C&%(L,>;H"%VD]X^%!YL2-UL)9IVLC3\O(%
P!IS<<I3C$I+ K[21>2SLYFJ\4!:Y,3E@6#?'::> %<7"J?XX S?$50^HUV^TT-&F
PD9+9VC Q*9HV_@-PB%"XIA(0T<%3]*6C=I;W:Y._*(=K:RLMWG?FTF9ZTL5 #L]M
PJ5*V/1"<<)[AI\SR>.$BS7EQ^I3+L 'I*]S7U2SYO")?P:JJ"6UT=>ACPJ2#/V."
PK'P4\#)H[TW9:E\8(]Q^/YXM0<#A"Z;W254U)I8XB @[/J6BLMU6!'!V(*1RBPIQ
PNVX8-^R&QPRE?]@$ /K60:(PY"M1F%'(>L>.:P,ACJYN_>](L5 %='<*-E^/]D+6
PE,4IRP@6A?*/+YKF#C1_@[UAG?FZ_VV3HIN1R"$#6Y>F0$;QPWX&\ "6SLGQOXP-
P:5GGUE&;=W6:U:.?'#=Z_7^K:Y0C@CSJ=2$Q^JE"C2I5Y"Y>K%D+-*QY'+RPDO]I
PSJ&-,.G\EJ[B^(G1ZF=SM7V3C-DP%I(Y\D',.K$T; 4 P" W59RI,M]=WO;0^-+G
PDYO*J!&34 .,8D'E3R&#N=]KW(52$LRAG.M3<),585'9@@D7IJIG3+UI!6HBP_A^
P8K0&%7?H1CI$>J#] ^S4O7LZK4UADF#W'O)T!036=@NP^).+6G.7(;_?0=J$W=2(
P:)Y6G X4N<*)$'XHBSZ1&"VG(X1\7AH[I2L&F5TO<OQ5=D':UU-T_"%,9YFK07''
P>TA+4EY+/FRU"[^_ [^IA3.3FTDFS7I"E:PJE<CGJ',2Y9,K<SG3E,^<WY:]))]T
PF"$P5I](KWK$XWTB8TE*#RMG] <+.91N(MG;^3^21.^ER(#,_RZ?X-T@V^'\8BMK
PD;<%%UD X91$(RW5;EQ#;".F*8+S.><^+AAZVEUBK3Z1FF-6715Q:8Y$E4UK"5D"
PT!3Y9,OC6&%U="*1-<.L?N;0.ZV?A<$+LL)\1:O^F-95CN%YY 4HW?A\BP*-S1FG
PJW$?FQZ,]94%?#SS:-.Y(#UBES)^#%TU<R!W9R4*. /OB\QXLKK6R85F?B]RG)Z2
P"U@'D23ZI#CXO<EG9ZDC)TYHW\Z;A\NS=N3DZOM= 81"OQ0O='?KH0[J\]1<[5@?
PAHH\HN3V#.\'-VPKLDR9D@/62E)0?<0O[[?8.SJJ\>$%C&"O;1/%6*\C>?]%4JH"
P=!Y@_1W6!G"/QI\PFDL,B0N$R3&-\A,@6ZU+SZCP-(MJ+[!P>;D92E-(@T3RC\AA
P/'"H<2'Y)G6Z-.9%RV11;=2@>8/P5\K-JH+!C1Z%_?WPZC*K\=9NN6F49,.%=IK-
P<0H7GN U/JXU">(]P >*[)G_'5__.59H])L._*^)>K4KO;R?.O71)O)!\KVTRK?F
P$CAWH<V3X^S3"T60X_"&]$B)K2H>)W7.P^D+59(=&;WX"%A$EFMI.GJSE-)*'+PD
PO%770'-N;ZSRTT%&O,UOIE)#&> !<&+@/8Y0$M%? *1A>A-8K":=!SI=QD*S(!04
P'E9A6[(JB#GF 4'2/T1JX/)R$=[#/WW##)%=52Z4I?OJD?C"Z67@,B&PF&=@ES4#
P-&L*CY^%(U[M]R>.''>^QQGY39JO%&XL"<(\L Q>5OGB<NIXXKR?F)(8!'&<<S\C
P!@0##O/TEV:&G2?#AFJH2'%MW8X"'U';VFA/$/.,X!EJ*\9J D'RYQ*=AD]B&EB<
P7-J_E>ZC$%=4UAW;@\1&PH2.='8=U/!SYR2 WBY6S &-0M6]\, "BM9]>K/P$NNX
PXD=&5;51T;M!7A[+/+8A_Q,LQY@(]3/;I9 "N+PXZ*N7)+\4T E&)Y2>C99@E6#1
PMKE/$&$<?_%% *."P8_6#GA"RC'C0MARDK\4OBNO!F0B=W7-FBEF]7$;=N3YIW,O
P$X))BC7.P OMX\;"R_S#3AMPO,*M?J&:<G1DX0:RLYQWA:=?H)@2H7\U/0(A7'J0
PS3B2 12KA_V"(I4R7X?B^#OT(T?QJ<(_(;++EB8"NDMM<(8?QZ+2W*\RM]=P&K W
PK.O\=^CP8W.K**P(*A;6+'[%D7@!RA/+"K5Q+TF ()-56<3&M4MS2CSV_C),6N%T
P/  _,TGNJKB]MXO40[-OR*4]USO+ZU4&R5WE,.&2GBQ25; X7MX@34O&#>UBW1#<
P\ ^L-'/AM&O?\L)5I4.T:=W1#.J"?\>NAKRA!)IN2C<<S&?-\%HW%_$IZ ?K_UT)
P,W]6.6!(H\"56.YT,*L6[TQ]<CE^2]4G"#C :5'-I/ )9NNKA3VZ#)L)\HH+S-U.
PO?IIF[NL:@=-=_YV-FXZY\,V%8MNQ/O47;+*=)P"B27V)B!A.361JI%RN5$C (=7
P*[WG$/\?[XWK96,O)2K_<*: JF)HW=JJPE47&/WLZ9[Y'>6U@2HHX'95]L_EZ[.8
PYCN+^@C=;TIY=1^-:JWEO>(_$)IY =(\48SW@W5H;QFR<5QYWZ.D1BD([0E7@N@0
P)\%RM?NH%0<I>FO9 /W&>H.@ @H]YG,1+$L_>%,"4LSFP%=<%C="8];QOJ(_=#FK
P4.H\:0A\K5@?KV=P46G(V#LX.'W/.>R5LYFV@GK]$"J"ES2VU5'ON]BG0;->QGV0
PFO+MC#9=[/#&5LO76P;O#OH5: U\N.!?[L[XI5ZU=S>I)]WQ;<<)GOR3GZ2WX.,0
P:+324"D$$[G;NXRH!4R\^L]Q836M)-5WL.#S6O.14HO+6SQMGC-"$C)(J7!M1FIA
P=1G7K4#2PLVE+UL@Q>948W):IM?NDU6^EH.7S3 #76^0D@E3>F^[/3+DK 7<>#& 
PZ ;8L;FD9>@7+!>%#%9]EN+5FD^!=DWO$3C(7H(I69,9WT 3$N;6.D)R_43X9Z;7
PU/E7+O*P:$A8!CU?/S6*LWF>RW^$GB?8*/[QZU8H:WPD/* ['W,0$4DJM3E._^PA
P-YU<O&,TM(<<K:R(>*SF>VAJZ#'=)6DT+P >\Z?R77X<M0V/U 0F3)4734:2.T\Z
PF:2&DQ CV\X>+4+VJ.TK6JZKVG3AN$6'9<_SQ6QU WV.SR@/A#=J6#PKVAK>>>(\
P, 1'V OAZSR20QKP:6UR5CPW/DD3H95LDJ(T=Z=]S$N(>,$&\'2%XO(*"5\6)8DB
PT4(TA.W'55:=QD* 556V0Q^'$0%YLKQF/0Z2H1Y=+H05)F_I!K85N%0-X6;N/C-W
P&_,J'RHE[60CU\ PT#<3O-#4//!=  &Y;P\64(T#*S713;)RC KUZYU][=A(CLW-
PZ+2DYJ9!3&E!$@B#RM&9*B#C^%ZT_>X@@;K+-<9H>LHT_94+=W9![\@)'92*$F%\
P4$5#S5NKM&ART-N*OQX.)K0U6,Y8P+RJQ"Y\,DU6G+)#5K;; RBUX+=>2A440=S2
P>TG=+7/=90IWJN].5VXTWL^LEL<F)CX]S3@H:5_LE/R#-@P,'2WSJIO &8"_79Q^
PJNQVTQ]7?T="2@[I%_/:"RY/2<"$S>+4MN3]D=WYO8"@&'K$#T#&,T&'3([C/^ZT
P+*T[4KS5L;*F[DNY._72MQU)F([IKGJC\D:F8)'@1$B&H@MVB*<^&L+$H866NGCU
P:GS[V5;ECU\!XMXV?.T[?T99X,XPI361JHITANPF$=*(8,!BX.%_GX&MOJBFZ(L_
PKBW6YQTW2DX&;8C4[LJ/U969=^KW'M0RZB/<*EAS=#]H@B)[JMW,UCV[?(]%GWUN
P.87$ 6G1:??1W3:/B@+:':;_D?FW%Y9159-.=O/;_T':&[/,(XE/3F4?N9$$XQ(+
P&V^L6Q#L=@+<%7C/;.47@&^/9(B.9/H4F&"")(IWL)/A(*7Q!,4I'P<FVX25HQ:G
P;AV1R_[#Y%,7G2,2GF]MV:CSHZQ(!&S#)PKKQK<+CHY+,/43X,]>%^5Q(1? %1S0
P"IF(0?8[ O_-@+OH-^JPM^Q)%GL4R (2A]?SV9+0+C2" /6N%NDK%;'\A;S2ZE3E
PNGE1:6(='<I\)5-(!-<E#V)!G!U[=O$R#RX-MOI(IJE;Z/1Z55^9;&!BV+3-9[X)
P^(6A)-7U8SFVXRK',Q.F2E9]7>;?;S5<DW[).X[@3* .M62C5%J"S<Q^XB"923$4
P]"[T!$W3]&ZV5DRY^8<U(D#ZXXO^V,<WI4.<"NE08T8DHART1W-$GR9W !,:88A 
P$"WNEO2&%6_42-UUG2;1GO/Q2N'L<ZY$'M!G>"I'S[]@.<Y* F;R,B7 VZ^;Q[QM
P[ST'*&6CE0;2T0WM8D"E_Q6YJ5G/*7EVW7N65+!UPCX(AI/8JG:%20FOL./X HQ4
P]F27<(T8*L20\A9OH4?PR"!MEKD;J<G*LQJA',XB]YL6)@"5<_:>3:VK _?\5)PT
P]7V/NN63) N>?,Y=[RP2.2U&V-3N1>\&Z+UQOC2"4HIT<A9>VM_.@)1C'&_(0* E
PV2U=Q@L_3NO!21W<IW/RJ!XQ@D);J?'+4Y,/MK)X]&S@MEM@M[BV<&&F-!Q2J3RS
P%ZIO?)TA-#/\VC*>I+.J.GQ$]) ZQ\A!/40URB15EOEEN7ZCVD8>7]=!S$^47"SO
PDOJH*&H".8S.0_.A#22G_IO#0K7AT"SN!KS!L&+#&R06HKVPYV)@Q"(*B )+)UM>
P170EQS]^]%QY*#DAV9[^+_S#2:YT71NR22HBK! 966=$E(Q$7J*ZK@$4XUQ4IF2T
P8]W;7(3T<#/W&:*(\3-H,(AKTC_R2, :KU59(:[":=1[9OIN"9@_;NYRINT. EV9
P@J1UEQEE%0/L.Y&9=:S<C3M!GA2K+AI-%1YH<\1+=MK&)KWA^=_R90S(1RR!0E*/
P=^N;6:=A7X&)+<2T*#HZ(R0A_FY-\FZ9F, _L)%<AW[Z@\<&MHN+9&S<VV634.1S
PRG$8U^VLJ>U!6]@D:[V2O>;> :]I-MR>P]5 TZ8$A*QH81%U)XT]NIE$5;\>+?\$
PI9UK)H66/^8-;HNAB;8)-*1Q..G0J6#8E-Z,:+P=]:IZ 5@"/J"#=P>A;ILFQ9-P
P.]SL2=!A_K,U\LN"6JEAQ130H/MC#:$;/1ZLR6I_R5JB)EUXFJQE\MA;'C- ]M8X
P -KKUC.SJ(0AQD72*:2BA.)WQ <3;G&O_PJC-#M1BAH.CJ:M&Q*O_@RSFCPJJ% "
P%F&G[3-1!C0L:,5_XQS^ELR-72 K\')!57 VY/.;:WT*ZV$#JU^%@1.F-=M6J/KK
P'7& *$A3E]:=ZBY>LY$QR*UAS1*<R#N'@%G,RU2:67ZK\>;7 )O[(G.=HB">R5*U
P$I.@0#)*N!+;:N8-<#U?S/ZY?8(\R"$B7@U4=B$15;("Y;4/E+0>!T%(CJ\,ES+G
P)I#8VX6$#4>PQ@_G9B2"OV.3JK>C-P$X%GZXBOQ2!Y+\/C.$>Q<'IT:0'(RU -G>
P&@\1M^IF4#%J8>6I:3@>9((80%Y>RDOKKN.!3<VOM77U:F4=!%>-9?#Y$PV)KB,9
P0:+#[K^ZTM7J=S/UB<UG<2:R@^3'A(:S*>O"0,ME55#H]15[^8,,NH[9N,"Y26.<
P(LF\^E*N\U&"X8I04(JG\CKG<U?797;ADM#!5+H8'+3JW_>W]_.4:Q5H3?%3Y*9]
P?2,W4MZ]IBIEOJH7&NR8? 05TB2#K"5OZN<3F0"09J?[_S<[ I4D1?38ZR=CIJ*J
P-;-6D\TRVQ_;92$W17[80,J9D2VWVUI);*DN>Z0.Z1, L5OK=8->;V16]L_\MY*U
P;CL3M8M?[@*+"EWS$VW$&-O4.O?:/QY@::_8B,,_$5'*)FW<+@+;=.$8H\@,_["_
P-NF>[Y*U1=:BB#=$)O>9[H)$EEA2"4DP W;C[D$()#'D:_DGP(+_WPQ$[S*9HJW<
P?JXD;$L=Z'I.6?_+_T;CC\-%!"6RS3F5 _0@AS]F +E:A]9U[S_<[LL<6CFL6QI/
P5<[_0#O^6\YPW#=@"\H"7K<9]:<!6X]='\S7K@/P% /$?B?H_*TS&)L#1;004J7J
PYI'XQ2[Q:A\M^V;'M:%&]+P[!5HZKDE C0:X#RW<0[:'[3BD6X[+Z?B"NE;P\:K;
PX=;-N6V(>G?ZDF[-BHGKPSW(ML)A*8,*1+(^;V?$4LEPF*0>*[57=-00\((O_*JQ
P%Z'Q17O+9!*FC"0X@'P^GQI@KUVX@I2VC+\>'X2<H98PR:"6_A[YLRU(<MWXVXH=
P%!).(T7  (F5M(ZYR_$I8-JD)'ZJ6.\Z^?U<[05HPR4YSL+\1?%X[Z[:UN&EON2)
P[*V]ELWK,BTL_']XV%K?(SW!"3(2U *K/?_9^X_96XO:>KQ9Y5HFW^E:>,869^W;
PM/"B!)^'2CER_JQ_]M"_H#4R_V:VK&CXHA9J,?.LIKT6GYIJ00$H44=<<LVD7YZH
PY7\@%^OPR9\><I,+3!"@!#BCC?+@WWKW%/R-V8W3[6@VG70.P&;J^SY%&QM\/L+D
P&6\"R"H!."NK4A,"PUL*,N;ZH2X:.@Z*KMM"E?"5]?PMT[WHISDZ62-7]T6O'.(Y
P:V:QY/O)NU]LYM[$20:K$_[._+:E9MS9/EZL1[([G'5V^MU?T5MP%<7%) +H31HL
P36TE+LZ4+5P"J5K&^I[Y[/]QEC'H4JUA)H[SPV_P]28T!$I(/=L1M8WF6_W3=(0:
P0]O[ P%% FA9PWNQ SDZ$\U$%MCNDJB@T&<V+2%BB]5RAI)CB;D^8^9E"ECI>?#(
P[H YSDAY<S5'8UE-QN(<_'626\88$ ,?V7=TKMLTK\P%2M$TILE>#S:<]#.P0:23
PZ2"><+"VQD"6N(WNNKKWC>0SZ+IWX( EV?6%:ORI^+U'^#RY#D4_>V>L4:(8OVDE
PSBM$B4@_D[/MC">VW@I*-=<>PM,]L) E@ :.4S-!98$GXFBI#2,1S_'IJV)4CAQR
P:@V*.$/E00(X$$:82M$CCVQR%]-7:R^MU1B75:BU>6KI ZN$F$M_:14Z4-$;D%!%
P>HKPJ2J-\ )SA3=@.&3R@R4<K;,4H#A\GD_(2.$E)FVA4J6BG"%2C4_!&^7GNE%N
PCX[@>--[_26D?[.+HO>TE4V-'U=2/:4'M\\78FL0#9@]?%-XC"6)1V8YE*<6BY,Z
PK K@HR;,0OA.>@LW5.U(5#0,2$/WQ P)\?C8>*9SQFI!*IZA8&F, !ENQ!Q\LPDD
P#)4*3FQ3HLY%0$K@%HA+WNNMD7PLE![K.Y(/2]<&%&^V$FD.L9;R!X#:TBIEXB?(
PC0C53:/D(+C ;QOIY8W3>@HZ!8HQ$%+A?;NU?YZOO-8T(:<BQTK)1NS5SPZY#C$[
PW)S_>H5F'X"7D^%JQK>KGH2Y"F'-V;F0P)9QQDTF"V#2DUQ<*MDE7EH%@/'_O-,U
P/XB"MUS7^:;3WVY<C)+'L%81RY)0X%>^V]@ YX#5]3$>,\C,RC:DN'E"-2!6[O!Q
PN[<C1RCJZ*.3(<2%',%?79.ID0SO7 H8T'T*T]T9\_9OX?NF,<C*RFV3IQH:(F1U
P#;<Z9.1!Q>"52^ <IQ-CI?)#J#)O&2(N4L(AGNB<@H0[+WDZ7MT#U2BN,T\'7JJ4
P4^'C&6(7QG<#7&XQDX7NX _+ASYHTA@U3F0TU*5/7@273+U<4*P#S))4B-D?J"3M
P^7HMJ25F2IZU(B9LE*4UZNGB.69KRH1:"4] 0U%=9-PB=R^H,VSAU&\7M?JOS:]'
P>QA7T+O?KE-%&T7X&1O'_B$O4@\8UV7-_S^K]/%BL@,7V1P7]$=1 @%ABNX-,66%
P 7G?$ *2"D,'L4X*0TL?#HA+VQ"+[9+3\_*62X*K@')1$>V^M,RD403E=X<D-M68
P"-<JL"M"(\QF\$,Z1,;F\7VVV3G1F/X,3!7"<A*V&O!81QOB9KV /B#I2 &_B6*.
PP+4;?!\FM!E\V,=F1YI0M(AV:7J3;E-'DQ"1+O:8SA\0(>]^RIQYXG(*9GV]^$73
PL;_0 1:1G3"X@@,?GU8KE/,T1BI6C\?KO-<V_@D7H!A(0YNX^_KS\X=.](A*7Q@,
PJBBB>Q</G#M5+'=H&QFX'Y)%YE"' M5E%*$LZH@=>P$0&K7";R2 &VT]S-7UN2=J
PA+M]X)@1KH&4K1C Z+]*&6ATA3"TJ?#''%-T:=F.Y5]M\'//G<^^N\W0H.1XZB5\
P-G\Z2Y8)@L.KH@VG[IZK,Q6[N?M4NR>#S=$=V5!(8Z4^>R,]NC',-,SIM]I/](4 
P@TGS=$E5PJH-_-%H.X?OW65ZV]CVPX[P1,=(L_N6\E7O#$@#+<;/YBA1Y[B KVO,
P^PG?0H&,ANDX;!GOM* UZ>M_RLYRN^(=&AX"5F1<]C$,*\L2UG#H5M_MI1BED&00
PY]6E)"9ATM@BJ;(5\,:D>273QUVS'"^KQ>2":)*B'H98 VBY+Y5ARI,+ 3^LL9^ 
PV"Q!6C8:)QE]ZRZ3T4 B4VC*@@6S63A8(]V#$M5-X-YRWHKY:F%-;0+N*5;0<79F
P'\XW7_:I^F(P<>P3TJ6W&JU:=@OZ!KN>)9 $:?UVXJ1:=ANQO^!8A 0R$&.4[.43
P]K>5C:2Y&DKSG>%HHM3AHLO"?XTW/)&'>'[$-19(998;!!J%-BJ)2II1.\EBC?I/
PDM2-AYSXO\>86H $FT&S\&DDK:@;0Z2>0!L-M']HI,DI:EH_9QS(,$]P=.L('ZQ'
PB%3CDOYY9KO9W1"FGD4$R8'\T,W0 /UDS9;&F_N-;<+/!.1[-7/AD _?_,*3\!]1
P5>FJ+.JY/#N$?'#U, <88/K@<3TN/M4/U$ #;G_::?ZZ2#XTRCM L"X6N<(O,"XN
P8U!.P!)S*KQXHH.ZNIHG7=16*I&.>D/%VT2]7+7;;/-V7GA74W5N']#.1 :%/=:5
PE5HGX)0!511SW0JQ;0C'+;4YW:^LB*/;3*W'4)>9B*-5-7.V[@6=]\(K')$M9R-O
P_T+%LU$6MPP8QIIP%56TR3*.5/5-]^.;\X_: =R#W("3_H/\H>8%"K!$5KU#_T/=
P'F8^&B7O$7N^R5T1[?;C9C?Y:<H-H0RO:MTR3>*_NF+G#@)NZ==TIVB^@11O[PJB
P\B)<@7YF.FV/NP$ZFW(18%$Z3?OG:7.=$ITN@T<_S_B,LW% *TE-6"M:X^B=.&*^
P/ AF?6/[,%253E1VVB!$\(;SRP^9;%3![$=GK;78,>?GP!D\(/V\<,?S"_@M^2M<
P?!B-+]*U J< 5OO"8PU*V";22ALIJO]@$=8-HM?W61\7TH[PT.HI/,W9]V0!:#=%
P+1]-B?N7DLXB9-TD_\@\O(MSEKHFVN:@5;!V3+VSV)U6> 3C64\4&I!3'!Z]]H8V
P_C2OJ&VEIP#]KLR6A0=,_\I8^HP_3\3&<XLF(P7OR+=N(1V_GOGAVS,'>7A8<=(/
PCS-ZK+&R?":->#,(4-(YO76A97- @JE N-5RL\P4+4/EV382-7D)$H=-"F/UO+#[
P..$3XTY U,1>1CKV3QG>-]S5JK"!_!>3,VFM'N>+&_O4)IDOCSRP_[(,&,8;@OW]
P$G""DDK3= &"E9LP?O=PZ6E[-$(OE^\90JRIX,9Z*_NW?C!:\P<+"9&W*/1S\Q>-
P9A&8L\?R=EEL4GQ%4(._%J^P:ZOS$ZG\A^EPD*&N!9>6<Z6S!3Y0[9FFOP]D4^_]
PR>B5Z,<-P!X%RT-B4P#Q);:Z?T7"YZA_E((I!G7=B'9&6T9836KVNU?1(*,81VG$
PK_+O-(JQ*PG* &0DZNW&.^'ENC4B*?J5CF,+NQ5MB^'-D^FB(Y@;%MQ;4E_DVU\Z
P<A2%OI.WU.<#:H W^D&YC5_J50^0&K)'&YE9"<',"(GP@D"-QN9#;6N=X99XNY.I
P3HR.(UX'J.)CF"P.X!&0-UCP+0!<8?Z=W9G;#W7>EWOO8I?MRC,WW-YS80>O8BM9
PCWN/@?]]P#2@U9HS>MI"=DY-!!3D^8L 5@M\M8I%R6UFG3X1#"SE0;"R*'.LI*-H
P#!+518>\;$8W(P/M/VA73MI8>S2$[%=KH,*1!]U9@^S43H">7B(]!:JKZ0IOI3ZZ
P5[N?[PT/SD]KA:>+B0HLD.=&-]U1E-T(^K5[V^LI-=TO]UB"*D?MU0S73[1/W/SQ
PE#1Z95D6"(#ZLR9F.Q?7L@E5PDL=><!(ZTYVX EQ+2U&^2K1>QO%&6ASO2)- /;"
PC=*4C15 .(=H0T'4)R^?HTW_J+FI-)!CD0<O  *%$>[]#6LR;321LVN'WHP_G&)6
P'4.],3J66"@H".FC_LT4ZE(;X^U6'GA7YWEZ(OCU^*>6-!4,KH,RW?) RXU01_U8
P-\*GR0CN=1R1_)\;BA=B(HA')@N9_HANX5G;.*VA><LY @WWL-HD'*0 GB[QATSE
PS8<28>2ZR:3T$<)WV="[5IJG"I-@[953S!)X%(638!+#EGN$L\*//7O#$R]*[)GV
P3AB2J@Q7<[B$!E>E7,Q=;E[B $2O 85NMG(P0!O"RNMQ@^;OZ;A&B]M*T[+L"NO"
PKR]'Y3^@EGF\N[Y_!^S<<,_7=&[3&54L1UW.AO4VQWI(52L=3QVD/&VL6T$JSJG2
PW-%K88G:N:E-C!5Y0\N['E4D0(/]K)8V2!;':7EP;7R('Y=82@5;B<DB^_(6U7L@
PBYAHY<MMY0,.=;HV<K%ZM<N0NOG4937=F"\H(I5R18*>,^&CFRNSM,9',F!UO01H
P&$U?J09A$)LR:3M8[/P;L+3")6,0'IK:WU;'@NZ!L=YR16G>(F35"(+WZFJ8FC] 
P%<S]$^3&L8SH(>R3.^-96T4LRUQ"?(A00AF"RBGB$8A +O[..,"-%+$KA19%$%N3
PH@QQGY!AM,&,OFO6L:'G]$T1(<=4V( JU@8\6V@<"*3[IU&2H3[UG/_6=%1$G\ZL
P%\KZIR=Y 05)&4"BPPUQPAQ:_IE)Y9?D81_KOV[N=]BC+T;0AAS2C^#L.'()OOE<
P7D@I5/VS./:'OP:'WZ2*+K%M$WYH;_H(M+3,6O%U]K!9Y6VDPD]"\*)+7C>_K[H6
PP,0)%C 9'H-0O&S^#.]G4E\XG[A:U!46;.MJM9X'-F#.VJ-1 !G9,!!>4ES\NF!&
P_DQ'U!,V( AP0N$9OK2V8[>STG\+WH,?[$UN^MD$JC%O:C@(94\Z!VY=>J#0+=?*
PQ+0**_:H@1<H61AB/C?<_V(?$**-ER2W,>3-L-YXZF.\ =GS*;;PD9DL7L+X3"++
PLX"YB-HB@D(EBB&?N='"K7H2J,"'/AR<M^ G-LM/LY4;=5#RC\W'L6G0A0W6%K<(
P 3UAV$(E_I\ D6"X,%ZP[>X+>H*5R4YM;*+&8<"SY S*)X5HIG]B?"&P-:D"A!@)
P ;[&U\'A2 QVCC,F(9HX0 !4@4>0G/\M.!<3L8HA-/F$26E=%3,P8T>:"F5J(#*J
PG@V9)@)LX:Q<_8X*L[G<V^AQ6_]B2ZD%F,=; H\1^O)R_E=0S%:ZO5M=\)4"-E'B
PE"][]CC^H4F!2-&U2RZ5T@][#KY5B<M;/P 9FUF0\4S8>H[RGU%N",TV,2&B&WT^
P,!WQHAJ3O_;#!V_/CF=@"B2G^5;@NF=$,YEPSMW.XR)I2.N5@7Y#'Z\-@BNHF'J&
PP+333!H>61A6B!:[M;!L5)V)K2+'P7^"V55J72KPB]EXJ"5WTLR1 N(?$6)'-9+"
P^.37/3*%]Z&H-\F6$@RGV#<Z*>[Q;THPJ;HI/<AQ=D:IFU#'FNZ+QZ31X%V7-^_<
PWQZ)V!0#6;RVLB 3UYB+?NH@RZV(![XL9#FPJ?PJV8O)7L>.AW#]ZX3&O;]*>4G(
P DG#P9L3HE!ETZLU[Y&1A3O5D^?=2HMFC0;(.H2P>;C:SFN(F?D[G=V@&>4SA$VU
P-D>50_,TA=S9N>&@WK-07%S$<<\B9O43:*XQUWQ.RUC.OA:BY/-/D5&&P'IS=.9I
P,!?P"<;1W@>)60HE9-Y;XZ^A[I]JA@.?-5WS;Y8KP#^\!YG$EIW?-VJAT9[K73Y>
PV:1!,(WG.Y8B )?H"^SU?!6D=EGE\W.W=P1%D]-;IX,GW>HEB:(=(H<*R.>WTSBI
P?!FM"FS@114-\J"6Q8=<+T#"OZ:7FER5SL(R"[F-!)]77LU$ZD<G]W"*3+18%ST;
PWC5S1X[+Z^YR10:XMK$WUO'O]@UTK:&;V*=7Q,&=JIO\01C\]30.8@R*/84^,V T
PVQ;BCMHJY*S#KQ 74@!@457.P%0L2E_0S]XQCBUT)0%N5"P"#S$^+< E(V2<ON5H
PZF!RXP-=]RN<!7\-/DO1BAAL('RJA$1U#P"!2DN)R19L0_7HE> 2) OJ"(U"WWYZ
P25T?THXP]-3E4JW45484"1XL<9'X'.N0:8#]M:GSF*@:29F$GSN$G\AT;8+(*<_&
P:E\D\Z%A.,A/_"$^;.V<;&#-8*C7L'O>,^7V[@ *3S*$ ,XO^Q92$YFQ\OUUF/G 
P*!0E4,]%LDPB&7G^7H=IY9UD1U>RAB>+;5[FF'+E:T+E[@P,G!TC?S_1588@Y-IL
P[PWA!UI(,FD,__MDXI"]>Z]!O-LD-+V;NFY7S=PP9:D+:!A?3X\W^DNY3D%61N!$
PHBF-\3>%5USA)![^CAKEO?@7<@8&V>C9"NWM9#"M.-(PZGQ:\XCTP>4B3"6/LSX\
PO/AU0A%]W?W;/3KJM!Z-\NM;'IQE7F(#<[%R&R4FGKZ0&[B^NV>M-Y^"TE9S2W*"
PS:RA":A_\5!VD=F\*='W^+P"EVEMY9)Z05*Y\-LSV3FXH4XCP ;NAA\.@>2ISQPN
P U5D+LU>,U_[D: :7!/D&)+> (<4[!#^T5=/D.\HA.>,L\^PHI%51([&GYT)\(LI
PEVESO8^;5&R--LPA_M:VY5KOG%\J \R7DCOH\E&IH5"EIZ3N4>] "^ADP ZT,.G"
PNP#_NO0-N2D1?F[(S?3W19-Y$%(L-TO9#KJ?M8/F=$/?>\L-Y4+JG#^GC8+/FZS3
PAG1K/3I3ZUOLC[K!%Q[UC^KP\J9F9Q=FI@5.L)%L%9M:HZWJ,!%$F'8V'A\ TGD=
PF?BM;/1>\C_77NI($ETSWBX7T(M='!,Q_+ <9DDZ0N%8J8.C'N!K"Z02>UJB9!V)
PA18RWH,5W9;6G8ANJFL"&:)RV2M,%P@^U0R;6<<"5];FHDT;PK^2IK&%[Y;]SBQL
P"5(]6C6#:XU[5LOGM<I)UJ0D<S=J&C/._O SED[#V3PE\R9(_2"%\G:ZUU_VGKDC
PJ-TYHP:2]M[M/\?4/IZ#?Y:*"]T0Q9,YX*X@$X&@43H>Z[.W["6M'Y.&UO5"B<I+
PH4@2]4UM=](\$"9TCU(D1^:H90O\$X;@_<IYZK&;Z'S[9^H[@70Q+.X4\(3\?]^/
PY^LNIUMM?4M23-E8Y=V#_[I)S&NT<Q-)"NDU6%YU;D]9^UE&?KB,>=<L0N)PQ<&,
P2TUF(GN,#,]%Y*2!7\="AWP:6MW$A%E1?*#1G?B0?U1XX:S-SB_!07B+/O0MDIBH
P>DYVAX)UZ)A(4OGR) 1D6JA79#/+54*ASZ:1)BYS@Z6>"IGG*UG/B,\.GEV+M(9G
P&@H[XFT-W=>$ME@H)3Y"4*Y3O;=OQY*Z/OI4[K4/1#Q/*=@BV8TEJ>TV\I26S6X[
P+7[T'-:"]-\:^]*(?@B4 !DN(0XFFQ1?;%%G7E^RKWCL)/>/6WE1XX#)!5 ,@\ K
PL>KV/@D+L,H2@8.J-!GB43NC/[%'\4S&\T1^N'T(OT4XA@&N$#SZ?HP47L:%06II
P86@]'\+N*I]C-%$K9NB=<O$S7(&FU&9P8V,CQ*6O?/]VZ!M>J(A_5ZU':3IW; X&
P/Z#XM"+YZ79W<^LWY-P?/27\WU^Z9K;SI"XA&;/P?(BPSU;1;!S0483-^(5!(X.A
P SSFB8PZ_@UUNFL:\WV4W6B$%2G>3XM).63))TN_>*8]%E/IVVG((66R7&069G;_
PP2.-VC)QUT@V.[O'M3QM>*P1TYJW$VW?*<9$+OW64IB]<_*#X/5UC; =*9,&]MPI
PK :=MN?_I2AN>):2DERY.5C(Y7YXW0J%>^OQTU7]+ L#X#8"&QQDZDU58M_D!-=N
PK'#_>4%S+->_7)6HV7EN@.T./'\Y< N>J5PM-$5H11"D16F"'YS>3QN=,Y-S%N3@
PUUBPO&H>7;/7W&V_Z%*UCJSH%U2MKDQ-9,.T&6;(/C%(*V^4DCZ<1O]"2#CGE2L$
PIUDZ)KR9,TA !^F=DW>V:;"!-G,:U(Y)E@BWGG79H[N;[F<1W.6[/Z]>$S&/O8*Q
PS[<-8BOTU,9J/]5=DL=*C=/*KI 3&2S72W-!6JUO8*#8(.%RK@98S XF8IR7NU;)
PN7DY*%ZSY]1H3OKU(&RYV^F*.S_S#)2:BA\O3=N9;+RE,M)1T)1A_>?;[.]><E^2
PPD@K1-FV;[;)Q=R0NW5S6-497A5P:X3X<W74LFP1I2I4TNZU/VD@HY/9O5WTU'*P
PA;XO@?6CJ_V&HZ/^X:Z4*M HZ$FEJ%^^+1I U&0U)V-Z]NFK&VKII>Z,6M:3%E_I
PS!^]5[>%N\A+N/@\HK^59ZDT)F P[IS,OPMQ@IE%MAK<+JI(MAM_0NO)0U F\,67
P[7,)_]%12[VC.2(I(SPQ9KP[ C%(_TNP'F"HVL\;KU;2YTA[P]''HP1#IO2D#[K3
P$R+J=6\?&8RP\2BAQQ0C\9MFE*7](6H"!0;!A[A)-Q)YV?-ALD\BNV^+!6Z2</'I
P<B-RL*FHIZJ48Q%K#>PK6LL'^]_""%-0A7V$%FB6H8'@8\GB#9/>%IS(=M2F3GBN
P<?1P-=XN@K],55!#M&"1KVBQC6750WAZ>L7F?^;=2[0:!E#ZMPCA27>5R._R:I<H
P--8G7P#E*9D<>L1_?SZ<;H]&7TQCN3(A_3XYL2J.78:XQ+<L#)7"KKXMRN+4*'+"
PI5HV],[3^U:YTV"#\(3CV* L%1+*]';L574<($] SKQB-TCJ\+%25>GO>&R>QO""
PT0AB8]GKAZ^P,VG2IE?WHH:*^I:-16 G]OV3@_-QQ5WF]2D1)F-69WV$Z57$#@%7
P/8&OCJ*N&^)#Y$SK-R]A'9?/#2$Q'.$_W]8/A_!!(9=1W/\<O[C9Y@2CPSH"*[<O
P.\4"K%M%2KD%B+<KT*(/"KINO8\40,=3]" RA.E/9N_5KS[WDJ>/]7%_OGZZIL&.
P=,B_?/N+3=@"-<QDABH]D0E043EO_UWFW<VX2T8W8AX[7';/$DU->2,2DAV76Y$V
P(Q02U[%8/UK3R3$H]G_A@*K:!:IIPU>\JZ8RW5NQY:J=9Q"Y%^L%Y*TO5S /7#'7
PXG5 N-+E+$^DE(9^N!S-H-DXK7)PSY%C/QC&[;[3.VG9UPX24RU,[!GY--),IH.Z
P,=(' 5^CIU["0\4FOK8+-C3WM\5_FK=+G16(O8$X!_JV#VQ>RMQTOJB"&NQ^)8E\
PR/4N)MFA]?BV@ R-(!FSE,_=42,:\@-[U2921<.'ZU7B*@4B1N=:;768>V(W"8DU
PB>I.?+^0.T^I\ B2]FKE>2,+] L&.N4N*JQ7CFO!L\_[9 ,/B]/%C6A"@,)>@YX2
P1_Q'J=F').C-'T[B*E$M$GSJ; ;),J 7T0I:.WR6.^'1,]WYP) /EI&)@*=Y?8VX
P4/':/ FP3A[3<2Y"+6&[R:AD:U$-7(GY9%M?5@./"1%DR%Z(Y6JW2U/,QWS/[4:*
P<V.B7^X8N\%ZW!D-FI$^8L'MDG9SA:W+4[!H( ;BU8>H:U=_7$%^4GR"9=R_KG,I
P(C1Z@H%2M#Q-8GS"]'"9IYK'A5:3P;79^^&FX8*[UN-XQ@<4^;P/4![>^=[L!V0/
P#V80JQ\ ^-!/-]\I&:Y"LV14?E$&[ 14F?70A&^\4T-1[H%7^,F\]G=1J)#7E=+!
P4EDD1&BV!CN(?_4EF.8=3Y7=)YTMG0F>VJ@@846<Z$W_!"0MWT[51%%3ML@96Y63
P1BP.O?L_R0D!'S74 LSR1Z$&62%*HV^!EA:S(:=Z(G%136 25U! "ME4>W=>L"TT
PM1T()1GCEW":S=+/+X2T.V<'>A $_W3>C19$8 <F'-^@D_0)X6;<RKZ<SWSLG-,Y
P1>TM<,04W".$>6#W.>9]-/0<3W4WY<.@O+W8=1>2".7^K'QH_H2SF/1/WL9W7TST
PKIOJN*[9L_@S(T:._I?T+QN:=]]R]/M6;&.IOAO+<MZX%6P?M<9EA>Z;J/%/MY G
P;Q(F%GI"QD(?)C\L]C HRD_)]#_IGD?%P>>B.K.[E4@^P)2X@80\  @4BD1C?AKM
P/(PSV/]1UTE*.J4<?0^7W]O%L51]V_"WJG8K[+U=U6.\*K=V#]_3X#K\;**:)A]R
PKL)GR)"520ST?=LS,39R34\N:,BV6 Y+S(0M,.$M[A%^7X7<4"N>\]I0!)HZ[QJ*
P$<G4H)R/T;HF7@:8"I' AL?+^_XMC(H,)U_9I]_5W0AU__+O#-64?]&DHP(25;M9
PWV4KU-@/K=U;H-=*/%EMB%)EJ0^QU].GUK+6N'>ZT]EP/:F"%>,3$\C3KGMC$IH'
PM,;>4#NJ#K'Q*=/) RA(WU:5:]!Y_PVM'&>?!/\3*$@C=Z3N^.$94IJ&]_($IM*V
P ^J9?,C3XCQ874SV0P/R9: V^4D+K*F5/M8_G_XXTLP>1>Y7W&UJ\[.M*,27X2$:
P#NL-U>?^^8,^B/NV4C_,3%B#FN;@L;3]2[:;0UQ"%S.L1MY=IB#MU29AWI]P/M ;
PY7:"GI\N$X+Y;2<R*D?R495B3O_1A,TMW]I94DW1.-7:[_2#>/[1R6E;AMXBNNF6
P$,9 KK<TF"& @U/P9U,WGNZ;(U@Y5I*2DUDP+H^>"$"WC&1,+*!879TBY,.?_\ES
P]G/Q"4P5%W0UZ]]>\3$U<!>XSUL)/X,B9OK9X$7UKY-ZS-@*^ >UUJQ>\QSJ>$PP
P=FQ1(H2Y1:=Y8UOW93\5D3R</V+%&"N&'-JMB=Y$+3'KF8B;[TLB)./(924=N"ZC
P=7I.N @<S9A7!2NO<83#;;8CNDQ)(@6XADQFY(CHW &:5#+#'$(7!DU8J5S1*:W#
PN^E<\!W.>+9!]FN LK=Z,U.3F*'K#0UFI '[56B;U8(._VJ H?C@1P8L<_"0*7NG
P:&K3=JBIMW24"@\^)G&3;IIXT%YG'5O>/.+;AMHE%I;X-XL[EPXV_WY8-TSUA1/_
P>YXHV-]H:)P%+RG31JBDPGBPR=1%%E9UV!AHS-H?&+;N6OR6,4.]TYM\F&L@F\D+
PI+*:RHADPY</U!TA>N3L0&LUCVHQ4F4]!?GKHL1A^8-*^@=[)M? DML[A:^"75MA
P\R0_QA(SUQ'./UM#&2;]T'A.IEFFOL%VN+6Q5]@C0OQ 2^C;&25PH/ JUXD!WQ9=
P3KLPI5@_8@!0MY3!6S&P<ICEFEH0K%T4JIL(C!1SMI^O;#6]TEAY&^7O=:0MZ#$*
P&T.9%%)R8[45 ]8B#[\2!?+>TXXL1XD=C^49E-^V6R*G4"*@"KTC^?4L56Y>:P:1
PF?L^0!&?3%$!P<9-I/AE!"<=T+/<3H,!H=:IF4BL9+&G>&^\DIDJ^E<KF:HZFQB@
PW.XX!<4)=-3C QBEZ A<>]J@(<5+:YC[FJL_", -(E %5-A\68H@CZN^0=K)S4AL
P>)TF:G;<<"0=&]LV9KC_7K-<ZQ'8AO":1[:.L\YWU6Z:Y4VKJ!WS#Z3\)@Z!DI@[
P+$T%"<H'WL(&B$6^93S%8P%4BD&#EDA_!RLC/UY*#Y_5K/*G846WHG1(5-8L59%]
PW!8:(/UVLSNK^D#HM_7T]<^3BN9Q^IIL25\U$S8!)T3SBW*U0ASO#Z>E5#'_,M6O
PEF7Z!2T]V.1N;'C'C\AK;E:%6E)<..4G;M%G7YK'"S\7_MU:#P"\O!S\[YZV,J$G
P%D:=DG-#::_XT$AL!V%)\X"%V9!U'G$;+.?^=]!)'=]11+0_,L//X[ =E&;Q/8%)
P"KW1! -@XE1GG-BP*HBZY>610QT?57_QA^KM*7&EGE$2_?8UT-1#!:JWI/.'B/EA
PAB63=_J^'\E$CKT#R"L^X#LD*3TD!2'%2/N!K+HMBN(\@'"_';&/B%D*+#<^RBGK
PZ^:F"R;%SG88C[S?.GY.)460R'!]@#</<5/Y=/&C[^ISTR6[8J]AWZA'SVL^F"P6
P&SB8+8!D5XC.)Y<C523M]$:]C)U&R9/0[!R>>S-_\.7>^T>;RIRV9Z>;X^K%;KK 
PH P[J4[%XZIB=.S@<RX$*,4G---J-X6L1(7/4]=X11S'(_3:HBA4L+"YOVK?3%WZ
P-&ND84,\3S'I6%JXO5R%8VI"K+]BIHC[,X ?MEL.I,*/:)Z>NVA,C7)[:YRL[A,I
P^Z9>+^4+% NR1=:<KJRQ2!FM-1L!A[/OSO.32ZQ;Z[IQ:'S+IY,D_0BK9TF7M3JA
P><1,X<$!5"UVX]R_I_3Z&J\RZ-+(]#?M_ZAC% 88BYS!(0720"+O>/9)6C0%(_\"
PB$-]>G#=,802L[ZQ_QA@X(6#UH"=7M(JG0=7(+-?6#\D[ID<GQQR*#^H,EXM$I\-
P:E\Z0'3:K=+F&NCFDNQPUV[7N#"5:/*V+.T!PWF?=6CS8*(L;R*ZX;_AA'(<$^!.
P<?).]&0LK+#"R5H@S.4X$R9#U5;@A,<FB'J?O>959J#=[C8$4=V::2FF)-7)0>_"
P#><&*H3HG[8<B_GT7!N0D5,,6)+LHL#TY#E'V1)7/F9*G6;4<TF]K^IJ'$2+^D42
P6BC3?EVPQ66DGBK_[,2!S-:R/;A>76]L]#>J4_MQH<(B"=KA,$&?ITL)2QGSM-W/
PC:@V6020/TKNM>(%#+I620\#]EZ7+RN*0Y=P.D;[INBWCNAB/UKD[>/G18L6U'30
P%\\F>^4MU<6;<1.D6"SVJTM>(8]^@_9'DZ,OV*0I?-#>MNA)WHW9J(V'J8ZZ/ L*
P2?LN",K,>K;5_*?P+6F4'!?]'0ZWF[K,1.$M\[4.;RS'YJ6K.CJ!$'Y<)'.(9,#%
P'PUSPN\XL75,?H4HS=OX,::P@ =OV6UHRBCMU_M:CMYC $MM0>\!5%=RC^[FI[(I
P*-C)QUD*1_*W/(/-_FVC3KGWQO%E\:]2?%7638![,*DRKM=V78L1PWQ?(+]^5 ZL
P4)&CU/&6#&]35=0T4"%=,^[C/8XM)\@ ]Q1ECQFV(FT<'6(78"Q$Z8+\3!A;M:EF
P50U'9H_O,M719\-XCDHMD>QIH\J570";Q9X"SA0Y,=BO>S9'T<+PD8GF>%ZI$4>Y
PC'BFC,#9W;F>,ZJ,^>L%7VQO^L04G6N;&Y-J<>/_]Z)1:HRAX+SAQ./7EY1TA4_U
PL[I/*OR$]G0#X(3I3-&B)6(_X;YT@@*1N$!*G9]\67,470Z;N$]5H1;ZUJ2.)*8!
P1'/UH=L<C@G<Y#NO*.4_(3\A]3QS&.BP%4;G6HVJ^J."*Z^>Y-=2*;C?.%A1#&C.
PQ*'D.E^4,XF1?U-ZS=H7"^17*K7$Y;ZK[[.9(1:B5)P2^)IQ(K0T%<Q(DH WLM&1
PMU#03&<Q'YA_)ADZ0"$D$?M/Y[#A N&;7Y6RG73583B6,WN$NQH@5 ".)BV1AFDT
P?ZP%1'?M0"P@R%"VIO<F>(CZ##0,^LL?OBB0GA&/:\ZUH":[VO'Y/3:[:9X%9ZGX
P?VZGNP;(-?J_25.)A+Z6N0-S?8EW4-79?4,4*5Q<,GY6;%NWNC52ZUC5?IBIY]$S
P%F5@XE?KDC@C29R2O8^9II*%$$1'=-74>8"\0L_QBE,KTTX\FI5=TZC)IOYOE0@"
P/>)+DHV:K7>#D]#9>G=@</>6FK5K/.0M2Z/CGP#"Q,/=+V0^V4B=^6$&_/G+$5'8
POHP!Z,A\XY71.<LDMLYA^K#G%P!WK.0I6B!SX7B1@""@=/VGMF-$&#"=6^=WGEZ1
PHY&8LJVXX,!8IO%Z#M\XH>5Z&T)!5INZ(/XO6=4J>ZQ;@ZV]1J)I4 O'1Z^HUU&Y
P7"SMUR]\BO0+ES4N)!\;:I$" HQ\#:U>MCJJ#O4$7TG^KW0GX7>#05"R36.8,@9M
PEI7M.(4J6=V3*+?Z:Y.EMACLLP*;#D4.$4B,:MW)R< KB: H@W.%G $>IEL6]U9H
P8S11!YHP;K^\5D,=D8DNM-8<U\OFLW(#[9R4BV$<>C4$+&C&%/V!WO$'(2&*Y'$L
P\_X3QBZ_PARH1_I$#E 03? #%H/K2@^P8UT1RB_L">Z)6].WXV[>LQ)$U-/3EQ%J
P0D'=TE"W6E+T_NJVF%73HLPW9S*$OA'K_VI8M<R$8AUL4_$:RB2./#'/)>C3ZSHQ
PD<08JN\B4$QM8<DF<?4?Z,WG3'>A #1W\!H(0$* _M,>7 O>0<W\? (2^$A%Y976
P.<X?LS*1*YL^].H2KTPQRBH('*TH%K)6/M'JL<\_%\7Y&<:T_!=2NIE!:<RDREI7
PNW=+X11@OL,)\N;MG6SW%$%6,O]%NJX[(!Z(DZG6"L9=!N&.Z;D_/=9G#4/C-A6N
PIY6GS2!<;5(9P8>0Z8&AGUEK\N5-_%(H:>4Z1)0R)T1(9)00Y/1YRU0#?PVV<H=A
P)O"55AZ><M6*O+ZY".*5D.*#$4%E;<JY+YYUC<)&.9::T$G%3PZ=2E@AXGWIMN-=
P$WIOG>UKONHU;</6\FDI"H3->MGF5"&9)QQ:_:U#Q.EI$0!6&:"P$ >=V^7%/>(\
P7N#3*^V85$*#),.9S*;#!\7O"-HMV3IA#FJVA2R;(;/K#X]?"$\4)'>1CQ+KFX-N
PVLR\Z4;F2G568C=I9Q1FX*(.1>!]]1Z Y-KX2+;]',8/W0)\-^4A'&#>".&;5@?F
PD 2)N]/U2<!]AZ9'2_Z@]:J._,S--J>I#$E"A\1KAV?_L"P)C<R W49U"M-CI8KM
PK!78AWK7B6<\;DU (AA3#(OY9+.RC_\[!L_3F"QKO;*/[8<3+K>[!-_)SI%[!H$[
P[/)J3BB1&^OFC&H1.IQ'F),1JZ_DEYE1MDKVE;)//M:AV'_*[-5H>\*-)T!G0Z8T
PT57X!#FJ*L[K5)=U>>KK(P" \+V*Q$G?^=7WS^/@',P :QM3V4GM2W6Y*N6/CEZN
P*WI/0'[IUVM4,ZB;&?&I"79#\IA&R&^Z%?+H(!0D6,1K-UN!N)OT$-$\E3<^(\9W
P^,X)[VT03AW6U%P:T_1G)1W4Z1"41)<4?V:K8A*/W^,X=3L2I)R, <9H'J^FULD:
PVE_914M <(062SA0D>KB KO&K\0EK1@?H_N3W)E>*PHGA%*[L$(B9MAI]*V^,JCR
PQPVQ)YHA@.+IAT+Z<I<(LZ8Q@R=#13/R.;H,C1H=^@V4>$JF1!EQ*JDW@#$O$K(:
P&SQ ?+?1H7D\KYD&N=!,\8R3\PL)H7I.NFU @Y6@/]?FA]"2HN_9F9ISM_S?E@3@
PC F<*U\Q6>>Y,$$J&HA4'V&2,'A&S(CNX.DJ6<([W2U^PQ&0QFY)ZC= N^%;F[.%
P 1O&R_#VBIMM_[3C,M 7!A507"#IY.8"RL(VJ:1UA]#+VD#_645.J<1J\*,])JJK
P8@(1'LB%<.M]E8**.7$2@8$#(1T02>H 0U&U<@*I_54/;D;NZ *<_!@>*5GQ]N#;
P!BBPY(C?$K 7^([BX"C"01"B6W$\%[2K6ZQ$\-'B4>]+.=S:NP$2]9"5B9+*574>
PO&.Z&4A)1U>9:3>?,I#0M/.(G+)CM4'*K0R%[WC2L6+ )"CXM^RI?A/WF,$MY8B1
P#)$&\NS:3NR_P8_AC!"XD]2CN1@5B@$2_\PDI4"'PPA%()Y[9!<;'PIW.)3N"J)N
P04B='3Z=;",#P47'-7X"^?B0BH=FU"B6>;M0/>2(*NE%[Z/,>& X:BVL+M3CV[BP
PU&H6+HIM31)7I+E=Z.10S:4'P'JZVQ;84> 2[Y0R2U,S2$7M4=G^7^!D<'V2*R'(
P =\(+R9D/4T^Z,.%,K+7>#3+)QW@: @VD81HQ4XM@\$,-!*DCCRS_#N*&I_IN)O_
P';X0_28+DKK[U8ZBFT"><LU^O5,7;0^K,B@(" "'HKSD*HI,KB<NBJX;0/!*J2J1
PVWM#!'A3S =3).-0]J4 4;&HAR/_30!Q>K I+!),X.FZ0"'NX:/2P'/IASGK#)[Q
P;9DG$CI]<QEU>K;]NYZ_:S%R>Z$^*Z A=/;7%UJ= JW1?5Y\AX/ZB282QS 34\\S
P$H\K1>EG9=5P(W,!KC^U8L/ D[*N/O&Y.KUH2UF1<ZXW[[HU@>B8$M2,G?=@?5%$
PP&#<]K%:"M^5W<M;DV,6^]]Y4[9JEU_HY1G\NU>ZD^E5!WQ+>^^PE#">-_07-_E5
PU3E"/IFZ+'*=7&=-]1NK4X2\H!5,-&G:YB3#*_>$=^SH?8-G)K&0Y?20P%UV[;39
PWLQN1_BK1R'"]R+J!*)8O:C2]&M1.E_P]+H;'^RSQB2!-?ZBPM4^?%VJFF;]&<4_
P&"P!OMEBP+X-UQET"%?^N5@L75'(N.;%GG2:C$:A=G, J;_@[DQ00X.8I=$@'$Q=
P4)1C>,8M2.\*R'K=^@>FR]61)W7*Y%QVZ\6*XV5+8)"Y^3QF57\M]#]_J@#;6ZR!
P.W,-2M$G*'^(+VB+S'K="-D@Y@_^_L8U1XL7WMN@>Y)K9@9:Z,FDA"@\XT;!)![&
PV/?3%'ZWWQ:6R O?_D-3/AD\&5U83UV0!H^\"ZM0!20N@<%IG!B>3_*8@>$FEU^2
P275DOGS_>"XPQGVB8'O.DV=I_#E]WAGG-&9,@G*GB#OA;G%&\V]6HD=CY88R'W<C
PVJ[,'46%50EJ59GAS;4>]BZ2#2KK5V[*J3\J((>%++_S'\TR\%NV5&K]Z1@U,!?P
P ^?#VH65F&7MA2T9Q=>0T".N;#HD.3Y$.E</QKMALX=!M\!BQWYV-?]FW->O'J=0
P_163B\J\NL8<J*H:IDL;(:^?*M[<2CW6>3E(\R-I4=2Y<'(.H1*=W39KK!SSC1N^
PMM?*#L]I_Y1TN0:%;I'R.CFO4-Y\) FL2Q+0(O9TM?*F[LUKL9G\T_AA.Z\A\@)O
P(SA)\,F&Z.%ZJN/J05V0AUSI=@X]]!HH*+UA^X)># :9#.0W!U?8F+(!ZT47T;__
PHKX\XK&-]5^_#UI'Z.)4<+-"\IB/JAOTRQ<AEH/"=@<-,%YQ::+)\SE#P=ZJBQ$"
P8!F(UNA0*.<1\E2E^XJ$AU< W);;W-Y%E-%(DU-;D0OYP +*XA! NF;X?W2]^R^I
P*F#J37+?Z,4Q*YM!UX#(VGL-O:OR[O>)$$==_M'-%,,TPAFRWKBZATW:P6< RRX0
PJEJ@>'8E79G4T.Z%->'@@(*B*;ZGR8Q:T47+_Y-/]%1*6<,5?B%"A&_<=K[.H T^
P["S$AM%.C%![E#/O>3:D77S%;==TFM4/>SK<BIVJA&16(C*&A3<SBY9<++JC"ATF
P_?'"%KOB@ U?;E+;J30#73A#438?6*H! .*1FJT7F7,>Z81;^3UZ."B@ /OIW)7@
P 8^0@;D@0$D1N":Y??J$Q<\&XHU,U:O42PDOJ-%OG\LZ<,H;"X37.+%[7_$MIQ&C
PP<?D^.D)?_G)@4YHQMZ(>,=?7@0*3-"._$,59;-4Y$))WFNIY$R=<'JU[3D0&C>Q
PB:'5J:7[D"O5/_3/CAC<+/X63NE]N?P*W[=%F/XIS5A]@M+99<QSX4T*DL+J5<5%
P(@CWCO 1Y3S6T0Z!??#RA(*5$EJ&M.%G##/>$V6AP#/Y>>X6/)1;5-9<3&>;'\'?
P^OW1QQ7"LRV2(MF'!(:0YC-'&>3^ +'7/]@ZFT:;$7,. $788>;0&&ZDU8I?K5S=
P>/=$+RV^K5P[:O=Q/^*"HN8))TN\AU])(280)"\:/W:->-=RVP<I@>&>Q#4LE$MN
PR6^$:\>M3<0_'$!!#4-O1% LEUQPC5&+F*GQDA2.X=/"A@B4X)GX8E-,,-<G-4UF
P-B\A:)_OI$-*U<5!O$55A55>YGH0C'CS%[8__WANJGRL[$RVVKRX'=&H[&U.H\1N
P(2N^M2$J*@.C+4>22KE] 186%?:>VV^"E#*:W$E8@5'WK)JS'OD?0@N8#S2<6M)W
P82F6Q:S(&:-(C'32I:TN:X]DD90H]0>G$V:T?7#;0$9K_5"C4;I#?55E]4YOZY7=
P7"_2"A6[_N[$JAG@E]^.N"Q2(:A<Q7\]<F)&6EZ3RG%/=*2)N[*<+(H?)E]HUR_M
P#\N,7TZV._1?C J_RFL[F9#'.3ZVTJ96/#0;./'BP+>UUDTM6!<*3FA,SWX::E3+
PU"XS$V0Q: S>)YW<JN!)/^Y^6_<:V\ +Y8@MYZ==$^B'\:3:)(,?.6Z]V#QH%AKQ
P+-$E/ &?^Z_U+?ZO)KGZH-043[O4@I2SD*&>>-O+N>(/KF2>..%2W[OTN7/6+=K;
P-4*HN+>)W*K_I=^P]J;6VR=6[H!_6Q7P2%,D'@ HI_:5.\.SW'<SZ$8B_:EG@ZDX
P!+^@]FJ8&)NM)@*Y!X@A+TMRJ;)&2@=OY#)D![CU-?92L&#X5$#/TQ/>OG%!%FL&
P IR6 L ^NBAL:@RN\CE\[L*N>AAX9HLN!F.WPA1.OQ=]Q2NE)-'6*N11+@M8A>UC
PL=VF$O^IF XTJ0]Z)6N4+S_]2=:ZR<)G:@F)J)5--4<S==A;JS*.RF(UKP'5*NE 
P#S^JJE [O.8&NUW6)WK1.GR49%"85!45[847N_N>@]"%R*S'RAV%CC['@:R/?VF[
PX]W_5P#"]4<Z8"@^\&=O'F0S"3!]54$P?O@<!=QC%2(@]-K]3V.>(OW-T,\^1A4.
PT2;-.3^2X#YI?XC;"Q!G#PM8MQ^5,6(L^\'*A) $K7FU]Z$BS]MI@9])PL\S/]+J
P>_2^]((@7&H8)// CEU?Q;71KAKRWFKZ4?W])YIHPN(+S-$B$ESD'%M.QH5[B8L<
PO\;UF"&45.YOLH%=< -Y)R7O_W67X(K=@*,EA UFS4%#>];\2IYEQQZ^[9.:".FJ
P%O@5=E';7MVI[>+QS3&*^$7"0ZSAWWG&YOK#1(MR735.$3FE-\2309= 7 &?FOZ+
PQ"*$X,&D_UQ)6Z-!"XA^@!SSOU/ /-6\HIX0:)-7%5/4]AW24MR8-L0U $'UB85%
PO[W[40XGZLJ>XI8?ZGP3"NF01,C5CMT9"P TCU?SW6K%8]P-3^RXI#J1P'%!P/UX
P72!=)\ 61#G/V6"N'-P*8D<7#:=LJJY_W<Z'YS*,Q- W8Q'D$:809P9"&V9RD].,
P"]<5JD4:F(2A-+WJ!8+!9G/2B]M7BEIE)Z@SXV"PJ8#-+95?BO6I/%FQ <TO,8P<
PS$E!>^-8>51G*!F_,2$&6I)6J%MN.02GDNG?L@-"60G+X383:ETUWU1+RM=!,:2+
PH %ZJ?D5MQ;%V^07)3!/L[S_5@GC7%W;(R8CV/\-\OR/(,U&F]%V / IA#D:61OB
P47(A@J(-#X&!\H\1XU"-K7;L/\N#86V21AY_\%OZ_[E\F\F+R31.4=+[F!\%;$@H
PXI1AES<MY_(]#X=^@5+NHE=QWU@J,/5*;G3?2ZEKO-3PM$K^0_I-(F'EB#;:P[$@
PRM6-OA&=L]$*I4:%;%I,TX1."X,S8<<XR+D)%[8X49''\)W>"TI'JN=+:AFM0#*4
PC*+7MFVI+7^ <"2)Y1BXAO[C&NI>T[ZMSXKB\14(M8',,K;ZCR9SKS(#_0#XXAD;
P.0,A8+8V8"2A;DZ2,NN(XOXK&B(-- R.M\UHF< R_>-4=[:&K39S=Z@FXKJ.^.<L
PM+3C3$3[I:=L?V)=W%LF^)KW>#"7?L[+,/Y"B_-)3>#^1&Q0^BYFT,_FNE-3 5(I
PY,:#&^VR33-#N?]1"B+4CMG14EUO7!D?SMKLCLTZ>30<V]Q T]Z21T^R(0A+9B<:
PI3<Q8_I)]]"9O$'&*O*8IU>Z]%9D$:V_@BB_R!#:LL);)$#;H0J)K+>[U+O9,Q9)
P+MF<7S&\R 1]88@&2Y#O#HKI%&S(0;>FN.2]0K'P*K9:7_JQ3\ R+JC9K>VXW8@O
PF6/\$&?E95O3V898I\N:A04]\KXDOWHKGC5=S1^TF35NL+W* (;R) R!W%>;K@AH
PI'*K M;UO,'89B6[/><J;H@#5WE& G/C_W# T/*RA9Z+'C$>\J3:QJH'*R5!L2_;
P!IQ.D%AB"O!P).9::0Z6K&IV/_&[F01?GMN1L#S^L;D-69Y.JR!^L0*T)[7*,[.<
PY@0;Y VI!ZW&'/D_ZWRCT-494#2NB;E\><M3&]I:4C)G ^#=%H*NYXV8HM [%&)>
PHR-MCZ,2O)THJV6Y?#O%CYL<NV4+^] *JB_/**ZY[\AM!7?/U;\%M>MH_0,.AB%F
P@+YR.')]RX$HF\$KTP%)HAW*!*5L0#GK]\F6[]3]!UV9UFU4R_7_5EL $#I)27<4
PBL=>9;N,VT$)JW;L\MJ4!?=TB&@BU+7I;&"M=Z7%%O;HCL4=R1X?B+$-=T/4LNP&
P$<O"!F&^%>L_^BEG(EA.=$U5-'3\N=G6>:QV@FWS15!:+ A#+EO/!1&)B_^B\CQ&
P$>EP'H,N+Y%RWTWPO9<(7YP.\%.X?E9KY@H'.I<>FH^0OH^PS$V*\+TF[;]D%D(;
P<12_O&LG"$?0UWVQ=5@<J*1^Q![5>"K#T3FST\]0-0783@A?1&<S6NE4?#B5E ,,
P @/#^S+:/K8<-IG:J[++,H!T5S)?A<7R_V)\!,JP$TQGPM</)G*Y<P@HG=L''Z08
P=CW#)*Z24/9%EYT\#,]K@%@>%'(%Y.+F'V8@_#!G SI2_E'-?> GZ9KE0)(XS#@.
P/A&$FVHE.]&^>H;F^/L."-/TE%4ICGF]PT!1I$C$YC[\%D^O:9I3[5+=]%4)FLI*
P6AAU2>F\63X#&-LL:,.Q7(OC1\:+*?ZCF>CLL$T!S#0<-W9M3_/+S$OL>4U<LE )
PRNY94H F&Q$S??[39G;10^*E\1*!F.Q%QA_))&'#<K 9*<Y6P]$5(8A'AG)^NIK-
P()DN:N-K.^_ TJ/O78[<A7VX4?B'V;QRW:3>A[!$N)^/E-ZT:(LCKF)4=T@])Y70
P)JVF+RGM3=QXSH_!<CPS7&C<G;<8"W/P)NF,O;T $K24O\.L7_:I1_H-B:H'J[(1
PZ\0I"FP(Y E@3;*]]6Q9:L$_$;JFJK<?!,"^ZY231G\!V0J<)=#BTZ'TQFI'HOH5
PHI?@""AORJ.-I0^6M7-YTX(2W2,\-06&3_#(%+-E.T0'4O@(N7;HIZ1-*\X9HN%7
P(5[$6 J_4:&_5@8^(CD[EO76P"PLH"0AE;WQH;B^9]0^?@:4\VJ4_?[]!8$\QQ/L
P4!/SW.SC'AS1DMW6_<]BV8T"_P1?RF#_#)QE5L=7CR6K@67-OQ]UU23YP.[.AH5-
PH%E__K4@@CEZB+[76VW4$H41K""6:I*!#?#G;X#E,#9$ !W2M[^@OR4NNBQG;HY5
P,:*]BJP ^1 >>FQ8)[*=%#)4RDR:KJKQ6+$1DLZGP5K[1+#F"A!T\_C%M8&*)5](
P2E2NQ2-[<?@5&ZB<T>#R0)XMGY?>  MEJ&/+[,,,_]Y<.D@*1">H,*>'K[=6+@7:
PT=CBS'-;2M@IC*@=,1,C1L'J(7];]*;0)4QP^[NP>F>\RQ'MD%!.C9:P\BZQS*!J
P+667=+P3.&-CG%;6)E*HW_#VS\98P/-2&LF$G\IU)Q&6(#0 4RQL4><Z&V("I\;*
P^DE7W^7-1)6D99S\\@Y+$3[,+]/O $U6_P(U_^D/DT?T6,KB9-"L^:BI-GID;K/F
P8$J"X3ZP6]&7N)TV@#=NOH+H55M+&\N%=I-,>].%6P+,T%YFXX* #5JE&T&A-J0H
P\TZCYLQ'SU<CQN0F85?6;1KE.J'>CCJTJ7];5:PS'5N'V_M=YNK]&P1TN6#"5<&8
PRO@^HU. Z42=?\GI792!X9\,[11 NYO3^GH+!2+6XQU0^+&,.%FPPIZN3(F:4R* 
PLS<',?+RD-64\4T)TM;4-#1*,92=6@4[/]WL>QQ'E[I4/1'_,SC%N>BQ8@@GZEWF
P"GH,9+)]/9N_1-!Z8\E^<Q).8%\TFQ+IF_P&G:G\<<[VH=M=$:M]MJD8PQ*M45]I
P'KM_Q_J[(R0,_P;OJQTG&1(T[84^>,OT!^ZX+B+G\5<R"&E0ZR-&(L!],L=ES^Z7
PY95DII<\N:G0[MD!,A>IJA/%)9EN<NKL?4V[I*Q,B.ZI)M5@E3Z47[CT!:7("*]-
P8J8':\*1C;M6/3*GFU&T!TO?U@9BX7:,YBB;R_A9:6<-,*3I:XF\R_;&T>;4ET*Z
PEMLXEZTFHC_L+PF&0-B&MT)[7T#JG()NG$RG2D73IK(C&\,9:02';F$T\?'CI&(8
P/<K)*2VN]IEY)*1?MJ,VT+.>P2($2SK\WK+%P))O?6\D>0B(O<.T8J/GB4S@=2=2
PW)8%3%;G?<TNMB&XGUC_%3G?M2$6F1I4A5"_UKK RYX&;\3771ABL. $1=0*L9#N
P!HKV[+1:[72[*&K*(1R$C)PU\'\:LJN-3Y4)BXH8_\I6\R\!T#"FPDZ"(I2WH[,[
PR%>PL-Y\DN!!E9N94^&TBRINNU!6H%=;3/D. ]POQ594P+*X'-;?D'3CP<'E5F,A
P1&O48K\?>SP3=-R@67[!VWI3D;B/'41VU"NR!]621KE8"J^B1JA9?#^-][;[Y/MT
PHE_J["#"E\2\=08(9C,'EJRO7JY43LAJBL,U7>%X10!CNEDUX%"&EH5%@J+:K[-X
P/G?;.1>)KG@(G;..>2)AN>(B\2P,O.#*GF[M+O@*73V>JRX]VERJ;ILWTBMMJ-P?
P*ARIN->I'A]19^G6*))_*^(F 'Y+PX7XL-7ZS#QNKM]O 8TGPN6:X^WAGKFE^IE^
P+JS[>W74 =3AK/C(EQ1=3Z0Y%!9>]DZ1"WYJYG2IMEW8IE\A6FD,D*Z[D\4L;?%S
P.WTW\)Q.!1D*P=VQ1;MKB0#KPW0Y\C'AI[CBY'G%+RM@$$LX#I&8CZ(2V&K*NJ<X
PD3Z2PT30X+0ACR=T1,'Y9%.\6'JW1,'Q4DHYARX-(*'C0*/3CB$\GN5B=E]8CDD7
P)3?%-\S^]DC/YIOH77UM#Y-7T".BZ&^4 JB,TTB^CVAS4NZJ/YAB$4W4%Z(&)@60
P4>PRKL!M5F\&SC8,HJ<P2U";*K>E3VH<J]#]4 !66T-!?B6:AWI#9R1XQ-;_/Q= 
P\^\@.@Y<N]C342?),GD8/\7=5V.#2^=]J;+!3@Y@?0-"D2)S35[ :E'"Y6UZWQ7F
P*]OHK<"3*W@P?FL4YA;6F1/A&(I[.&2[^ -GX6#\^!K((O?8>]D1,%(@;^4@*[WV
PU]%'#?')B(D''^W&/LYU4'3!,>AJ@)OKW(W9!(#I#Q3O'T+!O!]TW;*>8:2_T\S_
PU=7)OE-VU^-SB<?W1>QC+RK'W:V.)>?VZCU[<S09X4U,W67BQHE@KQ.@6P.<U@TJ
PQ]_*5.#6#<%<SS:QG$)&)#(]O!:S_%L1Z@#?1+_M''/GR;!<'LL:40CMN(UX)%#@
PB'G] X:N7:W]J"OM!> LK,3<L88)$5!^O!E0""_Z!/,8#FWZW)$Y!YZ"8S$(21UF
P/)7C3KY#3<:**3^==+5\PG!=*Y3A@NM@S(NX^ISG^7U-(:3 NK@SM_QI1=_)RR>G
P5TF2[6 W<Z"@(Q9.LHQ_Y'GZ'B.,X#JI5L9-8EFF@5F_!K=_0.>&@:</T!@P@V'.
P:1QJTV/!K(%U)6964SMV%*>XJRWKII;0* Z,%I'85J64$E>BDT0P/90A7VK=(&O9
PU!U'DWI@KX5J[-7'8B1KK0.M:GGV][810_)4E_,U/FV@ASH[IU1#.HU:H9/D?]+1
PV=L>S5)W$-&Q,QE9?ELGRTZ%T2&<7N(@_(&*J_,>TQ(SJ[ (FX#_HC45]0GOA*9M
P]2RQ9R_.H7 F]IKK3UX,J-PS)WT9(-Z/T8[TI2VRZ>WZ@D9 *(/]+W?C@Y=@P@"O
PGV[+<L)")RC$-/O:H\C0"P!>$]OFQE4V7[(ZTL\CQ-7G%9&J,L?/BGS0ITZ_-WR1
P $O"F328T_=1!C*_UKR2H*<)J+4GD^V I+R'38 _FQ:$(1BI[@QZ)Y#K,R_J/@KE
PKHQ394Z]7-8[M9R:=R:K!Z<D4)>XJSK!5.3]J<\66+9JN:!DR) R_M]:.LQ1X<CT
PHPW+_K%ZJ?!](#*X5FY'J>)U_8 UL3..])9,LJ[-881+!?J29R^HF:6^4:7/AF05
P&S%^S(0CEXM;BL.2G =V,Z&F!;R-W5$NE;E)OB9OXP'US6>-CW*A?L$W4+7TAF.X
P?ZZ[J2M3)-#^(6I&Y:E!=,,=7X!$/%X8DL=_L -=M%M'0P0:")RM7SO^FBF;DCPS
P1XLK.$D]MF=VUMZ0RT?_6( ^GZ:[19+/TN[!"9;1LTO;J,N.$&@=V5%YI-,D,AV:
PA?>6A] *-5Z)JN_M [$FX( YE(5DXB19XA&PVF3Y%[T2FK?(;5[K,UV$?P! P"=[
PW:^\<79-B2.)LCAKU]XT2;_$M<O0FUYB)T"3U@#/&6$$5(O'2VB72>@1J2Y>D#*(
P0>I,^>PS:XSE1Z[19]%GJNE[6!:WS_6"Z0UV:66D#D*<::['=NK_8E(H6="Y\._+
PBKN\?]Z0W-Y1N3<*A9:F1]],/8]7>:6'9(W_AT%T3BOOF#CH\(0N'9%J'$QP>\(E
PV3:EQ@[;:-M58T>L85JC4&;G N954P-3UQNU;+H5RW1/O5/5".IF&W,3Q ,#;WX.
PFGLMTX.G\Y@-IW^]1?&K]3 ]>>"\_SZ%6WRLWG_HK1_PS*@O?;>H)9SWEN39"FA^
P&?^46&C_)D!]7U('<_39OA1C%+J>LD74O8E9_\@)R_I UIMXF) TJ7X8\$RL/Z%5
P-3??VI@9=PRTE6G)Q0755/%%-BU#Z,QI/33'K&A=4'OVGJN4E/*UU-LSDF7(W1GO
PR?E<94MW9UJ'TP#L6T^$6^E2;E$%FZTXM,\6QE*! H:\\S,];#+ZM[.0$$B]M=YR
PP-_?18=B_@Z#6"D;"X1\. $Z]V74C(S*--UYLI3:Q(V2/&7=R4BNN-P8N.D>/"K\
PQD)<I)("_'XXFZ(S]P+R@YSV-7*!?L//YDWATQ1W.AY']@M"1KO$58,@7<"\(R/C
P!;(D5O=9< +_@42@I?]ZR,KQ6.4SGR,:/ -4AF5F>.@X<V!K0@)2\B8(+WQX[^F7
P<6',.U]I=7E^4<2;R1!D4#$R2)\YBEX[[Y6]$XIIOC3 "#+P-N&5"L-]LP7X D R
P%+J,9&,&->C7Y,2FHP,$0V@MG+Z.*:+L>TO:F=FUC#!C"(!S$0RH-_CL:P_BU=:?
PC1JEZGU1<C<QP>4PIF[-J5W3FK -AG:B3V*P"\">$QF1/-HM&!5/4;ZZBV7/H/2H
P4EY.3&51%^U3EZ,/;;A%1OE0(G^-+_ ;L6=EM,,3ITJDU\=FIO. W#IU^62O>8B"
P)YSK;[DVOR;?^^FS\4/<8IT>;-;6SI3\'J-W"B8:@1 <_J- 2T"C.C1,7F&'B% N
P\WZ].)1?EIP-!\$ACN3$CM@VHFM>+15/EU3A[EH'A0]7)M:,$.>1"ZE$ML[M_;9Z
P3DJAV$&/BJE,G/8XCV89;YJ=R@0NYSM_#=7.*_]$9];-Q*D'0J1*B5IW6R(.J;B?
PFUKMAOP)A3'HN)%AO0XY]X%P;'6T:-JXVQ-MNQ5+85'0U2XU/5<K//% $NIK!RE:
PZU5@R-T$=(;;,->F&;)@9 M3;N9;!044K^]QM3K$,ES"GC97+@>GMZW\QSPP,E( 
PRT*]YN4'>Z&W+GG7<<*0:2&'@71$,V/#UR7Y[M/F8"#^PE>'K1K]],I8V\]A9H7O
PHCKA2DJ*WWPK;=[ K$#D&/@7WXU5D$AQA[0LCB?@F"%X-P5;A<$K-@01F)<LNO[-
P=M"8O)YNNQRE$LE],+F/X^,S)^OCL+5HJODZ 0]I^GX8JV/M&<-H^?XC\6RB-L)Q
P&'PJ"Q6ANZ9>O'>3,&*KOBL1W0U"./E.^G_"H4JQ2KGG*C<K\%P"KX"XO7#3(I4%
PU"6U2P;%DN[%7S:@477X[P-'=V$2_)EM915+LG1)W*;SUY3'J"=L8GF@_A)98$Y4
PGO+B4<64B@1C9#D[%69D*(]@5*/E3&B)$=3QLEAFYPF(3:C/IYRPJ8IE&>@'1P-I
P2/+MMFS5<#=Z7?3]< R>=(KV>J'\B$1*7827WNC,).T-(#IP>]@LZ6\I[FU=0H4X
P;D0(0HBV(-TI*$&I%_F'YA6<F_A+N:3!M&W,_I!6S,HF<5Z@52%>K$9(6.Q$@&FU
PN1$FY3+2>INDFK:A'V]1\E\PHR>V99$PY_GPM#?HU(]0@*J4/,''^!Z X/#,D<SU
P>"!.T@6YW]7!Z]7DKVZY0H^,]TWZQ)\!KW%WG5H?"!9PAT=, (AO^D=_X H3\TAQ
P[OG/AGK;;%)N_Q[.V WEY)F@:)J#ME!@"G?/,&.'K_N]BYUOB_$OYM(9I7N'+#! 
P%&M1BYZ.4%%]5DJN?GX/]"OUT#&0$1XL/5[CZ544D9352,A?(X#1%RELUX0@%EFT
P#QGLW.X580<=BF[] 9J9D*):LZ[T9*]C[5?"/E*#(NOO_+E&:.$HH]QB'_>)CK&7
PMTWOHC=A'N6NG%YZH-<Q^]7ILZ\^I!6FZM]!6;B6 86(D"<8JLP"+..'W+SOV4R+
P=2$!>V=O\7L6S(%GIA]+0#,5X-\=YA/?S+H/LJD)OG#2RQ.G7%O%;D'\_#C+8#D4
P0)@MYR236$U]@96E4KV$[-I+G>= C_]#_3 3.6Y\J\L6DT--6%B:<7 KA1B!1W+[
P7I*DFK>6^E/)2>E'?=]W_:_*A+ 5:\#158-H,LE5>%X1,>P_=+S'K$6,>+S7-M\9
P"2$E#MU^4 P(T,6PTM^-4:I\H<[_/OIK)_M6P(\)_<J72"VL^'^T*2!W:$@3[5J_
P6WMPE$M'LN]?HCT3/D1@0MO99?#+VKE\3V],.7_8_LQ.-#"<W[:!"<"6"^%JR,!+
P<[>EN5X9 =PV*19P2!&W[_RISIVZVOR !]&F:F.N&F(,KWL0E-:=$RK! H,L'PZQ
P=9F=QI-4S\UWFH]31+@VQ?]BJWPVXZ6"3IA!E+7*<G2,HRE6XE4V@D>M&:$/86/%
PFR#;^R<'MG.J339D:$HX';XU"=59%K"B1!=3Y96$G@NI5X*#+=0T%3<C%V5OO0RO
PYVIBO'1],79H1MOHSZP:T165@R.O[$61/RJ: I2!13A#6(OQ+$JL[QB.5VH*ZY4E
P6F/<CYO)313J4?+Q3FL.H<;ZR,+OWNE=WVTERM\FR"2#HCVJ&):&31OQO@DD+]!Q
P+AN'W2UNAW<\OAV#&=__D(>!+XA2")K[(+JSNJ0JQPS<.^B[Q:6AEU0R5AJ9(19^
P6*;9&A/0O<>'74N.3F#USVY&'7"GDY4FYY\08?S'#M@UQ*%.[(_M8Z"PX(WD.]"-
P;FTCYM!E QM8R<=.@S%S/R174M580B&VY?'/V:!^\!I%NTS973PW^"+WV!V4ZO>0
P28C%'*GE+"=+00A*Q#N8*^ZE+&@T):>3(7OUY.7[(%IJTHQS')S;&+4Y01KU!4,*
PS&$U8V0-795^RT6GH-O&BLJT4U%%\SXKOV.*X>"02BZ1G\;F ,3Z%9$:\SLFFV.Y
PH*VK'O*W7DIRB>]:;$8YDB5+9 ?F0*(E>Y9-Y<Y-X*\IRW8"H<A7IG$MR:)QL@."
PP0V!P[*?I.>H9#(A\X/6H;JMXAJ+3_B+BOOGG)?S4KG^)B-RN&<S&XYIF[)ME?$>
P5F 5=!WF*(.!ET!V_(I7S=\V^5@0X;#_"Y+/BX.T\')KL'3BVNITY\3["U_%;II[
P#X 1PU#"UJ?BM9#NFG9.P;HY7/45.F8E""7Q]M&HFI%9?KC+#PY^!,1-Y$/.MR5A
P^LIET_A@:.:CK.RHC!%A'&[A$II^";\UFEK88NGV4B1&BJY.(_K^QMR+Z9&L@]PZ
P?20%G3-\J-2Q?P48]=?@EO#0MR>-L50W:^CHDP0W(!EJ#D.C!DMM&?- Z-/A.BW.
P UR4>OS2P@S\=0HT3G\M,C86\EV7W)&^+A"1-HV<YULKPALY>GLDB'U\ZI- >V)4
PU!@,&H[;RCDTUN>_9K-EE?/X._)XB;>NHN85!-PI+T7-!E=NB5()$OTLEK8S'.7U
P!'QZ82&;CR G(W,GY$#>G,P@?(-/+XY4W* )(K=%)N*)B]AO*8 N59;82@>^E&!)
PL>:UDN1ONMYA?!&L9QZCU?-+3]T$<W]<B)^P"QVW1$#'$)^-/%9.IP*R=?"K*ZFI
P;(Z<\"KUG;\L5?\ 6KOQ\B83PU0,^XIFAR+5(0VB<A#6)'6,"M%5X!]WHD.9!!X7
P:1$@BM%;1.^]4\AA/ S-VF$7?F!MLN>-3]SVI5++^@>_,8V=DKCV)?D86YDQ2_;%
PK(U*T6W5LES6UMR9%D0,:$P5")LAHUB5NK;OP(D_MB+D1P^>S(K,(-,D?$F^8N!G
P<X/P0!%'HC&YL]P@-24T1.IEF M,"- ;>D@@DW D^G^[K^6)VR;F)WZY=AVKB0#2
PA,Z,8&^T43A1Z*_?Q\FD4C>>=[K,<:)0_'%!)6(PH_KC6J"/C/<LZ24!3!<JQ@D*
P3NZEBQ)!N4^$%.1MM3EB:"O<E[FQF,X,D$(?TWX!,]T8"R7"[<^P)J*TT'R20Y'7
P*,+0ANKF_K_8QGX^W^92*H7"3?DH1R.HM=>1&79^OT9\723GN:X%]F/85DL,Z[%A
P!!!D"$7A@GP]B925%VP^/"0S+/_C3"=OJ\Z:'_P7T9VZG$T3N3-.#%N@M,9ZX13!
P*[V/ '0W<3#RS9)C^[K&U+9)\+=U&?/OJ+<JVQM+(WG]% R@9_6FBV:E9X46)?6E
PPHF,>11?P&1'C/0A>X[(J%'$LJ,QRW->9@IS:14^;.)\3D+ GU5/$TM--[<@F-%2
P\W2(RYUS2[AL+#'(7>9(:JG K?MCCCX@"OGO14;HP@#<0WG-;\/OI'S1CP2H>2HU
P5:^QC)X@R7Q1YAS-40C6M$*C5 V$SP-M("D2-"&H-C4AZ7?",O2.+0#+/<JD?<7;
P?PEZP55<QLS>SFDW,,!A3]DW>WUG:H(DBSH#UU[$)AEZ;4TOUJMMH)B"/1V+P;:2
P5I$C#;N]ATH+WM[\<U5"IHJ(\@8^65>]#68$WF(N<,";?#)_XS#T7;"UE-$^TTT5
P'#^&/\;UM4BYZ L#+J\7(SA>*?OL7>HBD0GI]WD2195.U6UDP)<;^CI&#)D)X[89
P[49QC>@9D(T< 7H;=MQT-@E8_Q_E@P?2^\_OPMR857KU8<*;] V;'*['$!P^&)\%
P^4A<%W6FRT!SYXCB=).*GNN6=RL4O[RC%X9XX]L?_+]3$(<8K3F(PR'E!_6E/@-Q
P@X(=TGER(WDW0O[9BGN7[<!5F]2WX%BY,*AC(C(DW>,4],+;Z-PE)36]"-S_F M^
P)0QA:G[K#RW.;FUEII_J[(!P'*-7P+BO6PACKC J<#1#ZEA^OV1_I^-9NN &J%B>
PV7TKFX^YY&NP%1A!L1GQFX!<7GZ/H8)!3):RH7#M$C!H9H^S&.9]P8WXMZHPC97=
PQ2NS[R<*:J.7C"O^E;(,[R4R:S$ URA K(T;U02^:53#TVF]Z&54,^+JMR=A7&U5
PU/Z@<0%GMP=G,9<S1PR)PIAN%)F.2;&F,:'U<_-XZL*D=KWSC%V=Y7@12'>Q)YLU
PBZ X9IHS*6DDEZ2B(RVA5)1CVJ<V=Y33/A9?K'-VB[E@B?S#P2Z1%L/:4 (-OV/+
P+TJ[ O%"JL%8UH(]#!1PA@IVXN<'TY8+F84^KZ,-%:,YAG)J'*:+"Z:$%Z1XW>0S
P2X;#"'98"45F!51= 3#P_JNUK=8^>SAYSQ\Z> B5AJT+F7A0)J?=*C/G<\[36I)R
P#Q3,A^'DR!-B#&?@<VS!J5 ''-0\F-1'R=Z,BV-("1!MNH7B[OX:2J+!O=.-XF0[
P!N6Z5J*CTKVH=E:\6_W_-Y>:_/,>*W!XF)/3)5?[@:Y0%R Z_O^'E64!X-H.?V7\
PT55FKH;^WQ1QWNX_34K4L 0BNE.[H.]/YC>5R%))"GK<#'.#]F&_5.':+]UXJLCA
P[8F@82-T2MM@.X BF=SBUM&#-AE_,X;OKLB_9P9P#MY4FVDPC:G$RD6=<6TR #JW
P[)_MWMC%DH;5![[S@//C<-+\TRB(0EK_4?=']ZFWH!6=K?2F[F3(&8]DAIOII2:3
P1%.ABCE"=:I%>:6N;<PY'N7;]%'"I5+^T$$\(OB$.T DA@+X40PFLEHX@#9D;SI=
P.V:@)<'>D/G(0$Q"X+W@/)OQIWDYWYP>WX 7H/W,U.X9TH)(B#T9BK5W(\GI4OV_
P4C!:<!MF=X4[/(YV5GN'XQX9"0KW^45_2AO*:V)-:$'KSWSXL30/N8NA5D!9'VS%
P\3?K0^7#>?_] G,^E)78IZP8&QO9QUPG5^VOS?(N)_VVNJ\$LCT)J'4@N]]=QWD9
PH!@U*=32MO%UZFLF*[]-42V)TW]$79W[)\B$O; :N )LE)&O(MQF\L-IP)BSP.Y5
PCAW%M$[.:FO)<(5#!I*"<&*U17AZ1@<R/=W^'"?#D&J)L W1626:#[H6%0<.0DUI
PE9[[EKQL#)JU&(U(WXP.QE "5;I&8]B>J4L;MI?%OIN'$&Z]'F>D<9,R[(VE1^2#
P9JYD#9U:->5E;13R%*2"G(24F\#?SAYAZ_QR5:B&:Y>?HTVX.+V&7J7/P:<-.<@H
P>7O^-D@F7U8_(/!TT55B3<"T+VE0W:MS8GO!<G0ZXIZ7PJOH9K6J^278GAEBB@&G
P2[U;1>L((_UL+?EB&,M! A<MLK[*:UN5^GS*!9?%"0J#V'G<5D"!^^ONEH=J\&JR
PH\/=GQVU<@SJT5OF(A@"105<DGC?QC?GB*&1I<A-,<T/.GJ[BA9T-!U[L3O'[=V@
PR;!4Y &C"50L3S7+:HL$4RZXI\KM_)<+[9"O G4?13N\?RN-OM-XX._Z6AJDNY0F
P5N2-J)(E_S6'P5=?2]55#;M&=5RH?)U],S].P$K\OE7X&5JML!*_N(;^[$OO#<Z@
P;!T#;87]Y572V9B!0,);,M)#6A&UUA?O4N<%O!5I&@NRQ ;I?WT.3<<"*VP"LFT,
PI/VA!&IMTWCR12(+D(XO-S%J5#N@5! ZL)@:,#1G(4?Z8Q8]:?-NLSQ8H.4.!55'
P?E0^'\P+A[L5=DNM@P%7#CO;I(#WCF?MRRYQJR:'%W[:DE@.L0C_&@N\.;N@5X\Y
P?(:":.MVU\8#,06J3DIZ!&-,MW8"GV\6(0XL/045O)\4!B4_(F)X%M3M10U&8%8S
POI+.<_N6*-Z^,RL!</CZ<,@^2.V=4J+0'0%2 M ;/YMMP%D)2?,NYB/(XG]' RK$
PPW!1H#)M@I=I*AK?B)/??D)3KI!0UP /8E<<+<H#=TNJ%/C2#0?&<_*Z'4K7^?S<
P+9P^;C>+PV^#>$>6.UJR\;VZ[>D886'-)I?1G2$EE2L0REGY6L'W0N_0"NA=6=*?
PKK.9GME/O6WU287!-4L)L@J0$R"!\&,2<7Z'N?CEB/&L?;0X+-KMWGD=$VXVAG=.
PE]=5^31!O]"82GU%PC[(+! /AA)S,Y%DD->YXX1&"8NI.)'H#V+;#EWJRZN[G6-4
P=23AS?E"ZFHP;E"\]-5*'##R-3NB7TJ^^"&2BW)"N($CT?O%DR_Y($[Z";7FGE\"
P'@&8[S)6!H+!AP+_V 2X&:\</GDN4BCR*<45P!XORSNV3=TN;JMOK]*L$@H0N;T"
P!8M13FA"(H7> ZN^MFXF3H0T[CH[SF$ F9K$DDFC1FE7;3I1R-Z!D9^5>O1_)1?L
P"JQ=Z(S?-$3+L(79[][0>JGE-/[RH7K!#E['N?.ZM<DJ8GYF+, VB72>]<7)6@)(
PED>"JT"A704AS1TF23]H,$B#3?>XVIQ71_%#6*'!$ JW?<]*O\])$WQ5>W"W(1'8
P03CF0_]:_)#=)!40X/L$Q&S\RB61!BW FD0$PY-XK"<B=1S^Y.0C:*?CUQ(X4E&%
P]N2"_B7O*0NHBZ303RV?4/KHD139; QIR6[5R3ZTD(!W2\-YJV3/Q@SNZ1$J;DO'
P[LEZ1!G81:%?Z^C7+M@Z5HB *LXR+8,4I*C.4#)1?N5M?!9.*Z>0VE-0/UFH#9*#
PM98*VLKOFZ4K&&#KH##!/4"G,@P"S:(-,C]4$ ;L0*>?-3.$:BP+($$YGJ GT_,!
P:!0"7[7F3B ELKE0NNX<T*YFI)-Z?!]'HZ;$9&QY3"BVG'4S!FZL_+(16[\:]V/V
P)T=^\X%[*;0E"D/B'@TXQ1EI?&?L',Y+&/CA1M$(!W)U(I8R*R$?K'DUR?R^E,$S
P$^7TGTF.SVCMG/G<=8@A[+$%:ZTJ<K.B0BWJ.3FK]<J?L:Y$DP=9F8!!\SX)'U4G
PK1#B"' >12XW,MJF%8VT5?/OO/P^BK8+.5SY@\)U+P A!7P!UD@J0RQM#@K7.GK7
PJUA]S2_GAP".,U'/V43<SZO]')$^K;8H!)@&)P4D*2PX9@UWH=JZ1@D/Q5;=*.OA
P^P<NQ -[)M;FF[9!R%]M#[6MI[$\-I]]X4(,(-\>SQ(U#O+X[$IYLM^CA<UC%4&+
PZ 5+C3:I/F]T;^C&HXA%O!HC:#"\P03N&XVZ@@"CMEQ0L[A^\'%R2QSELY39G7W^
PVDC](F271TVN3XF4!]$ZOM20[I?$G24XI!R:-K;]P+5DY?'F#F_!C,$!;!7L)PSV
P$N@>^ ^\6T9M?6GJ,Y=4T-XE29?Z;5Y(?,"HQ$$K0*"(<QE$_5_5*UYLGIAT%S=,
PZX\=_,])NL<=/@HW ?R=Z3;@Z4SE9FD$0IQZ'/&E8-<<TJ-39D9X0<]B:NXKCI<\
P&+!2;\;C "0@)3/8+@U1CW_-H(LIBU)$_%03$"V-JVO5,H026E^Q_#S3@%*WN4LL
P2S<>D@7N"/4BG26 &[9A^C(QR"PMC'0N*-4>_)GV#^G\+I9>MIV3_DVC!R3Q'\^3
PD8+2%**EV[S3QH6%Y_B/9G\XCT_L?1V_,,!6< _OMKD K57V<0](-VW6N4>MN;8'
P>ZZD-D,:EP;9E"Y%,^!$P.L(U%ARD1@/Z1+3+SIX8B7K4=X(W-!XU;=27MLQ+ &_
PVF'SGHP4PL?+3PO\ >#_M5,=H0#,HD?0_.PMM0D9H)[Y9'(9TX6">N/AK6#G>]HS
PMVVD!BDVY%8?NS\]BK++1L5G3FC ', 78M 6Q5L+H)8@V'18 I>SFSU[&U@6SY]$
P%@]S)A?;,C8N)(57H&S%YE3F"@38H^RJ#4\L4<EU/C:CQHI<[WN?3@RM11C+I,<<
PNIB[))V7G2@$%5U0ZV"LW$0$IXA_C1WE[U:L5^?&^ <1Y!.=Q=[(V=U43 H KC*_
P[FL/"A?>>8" Y'L[P70F]71Y&?3M-6@$9U_1UH:%;A89/"/]U--BB8R@2H F^&AE
PA;OOSV+P@0:)39,@Z+%AT)#>H:A&><3H2CM;G3]K*"+%OB;LG"CSAZ:VZV#$'QX-
PB*2.E*[(ZXJK.$@G&B92 "3W@NCZS.PC=^""OV)XX)C?7WS^<;T"NF+V9W[&_:PW
P2@F_ G )U3]1DG;D@VJ2>8'1R1[*Q?WU/%DX)H=SJJK6+G6$3TX<+ECMNSS3?V;/
PRHC[]6<;VC8)E22FDM&%ZL+E>Z \I[_(EE] U@H+E+*C8*((&BE.';["D&5IBM2Y
PN@"A(N01#<DLWTW>J!_@56)S-")V0SQ]?*K.O.GEF1%C(V**AY25V_EEN7< T L_
PEDQPAJ3>2* DFZ/IZ6%(H&?B,O^9YC(D)/F!TW0?U!*:I)%H<+J:[."),[:<=3G9
PIU/[9L>Y;8WGKP!MXSHO2H]N7F4WN=6>F5\Y2[YJAZK_H&!TFZ@1"G>B2;6_ W7!
PR,( H!_6,Q#$OH1>#3E%?_%OZ%1E?8MKVGV--.CF\)&4*$ ]K-::O^92Q,1OO.18
P_D1P*8FS&]]]*/\4+1ZEOB+DV>436W&&&B4R&H=;."<C 5O9/K6PO^5H"YG:NJ7I
P-(0Q,8]2ZGZSLM\N!W"+JMP0;;A;[G0<>\RI\!PXL"$>A%W3-?8(^"2YU<2D>IK;
PL9IGRW"0_(A<YU(=N;?.NRQ:.T^C[_;*WLA[./CA=?2_L#A/AI( U/*$K;"G ;_+
P<^Z!&)+/H2 /A*(8NWVIRL=YH&M2384F#)A@#G+[WEB\AU0\R02I$SXM>FZBC%O[
PAWL+;L'DV+*./QRH28*/ %PQZI$1TAA9DNJ9?4*1?<)K,DM:;_$*BLK)X8$S2;1+
PO!6"L2%0)5EE%-&!\A^E",T5K 4LWQ5A+"/$)+19.WL)W?C>N&]E,(A>'R=M/Z7P
P#?.AXK,''$A-LCC'$TOTJ*-88;OC;/\VH]DR.8B6F5?E^I 9BRQ6W3E@@]50+W<0
PW]M+,D4^9:&B2+XML%@MWX&V\GI(4LGBA_-B$PIQ@1%V+LE&>]]AW"R7'IC.[/3\
P-1M9C:T"K<I?_'Y&S:<*K</D$346=_>2<&78V>?.'@\JTG69Z$=_D*' CRL=8>&F
P3.97./VBQ2WTPK'&1'7]=&F@ EII(IGT*471-8A_\&9LJ\&LXMOD2]?,&0U9;_@"
PR 3KPADV_WSYG[HC?0NE'G@LA-Z,3+SM;Y#ID=DRR(N@23V7+$EKADQ!.YC^E/>,
P:*5>B:'Y-3-_<=?P]'J2+"HA:++[]'E.3Q-Q,RXBE/ZJ3K3Z%AH<=-9S<Y6 4]U>
PR*I)8<NF*[:@'@R?#:'?B)9@"X7T6%]D<!!<_Y")_O#;0RPX->)3U[@+87M+(,$(
P^>S@O1>O\#AK'*\F?^/CI_9Y@\5UE7=L$%5$\T")W![_-1T4(DYJ#?_Z1URF2UO&
P)UM?LNO![5W9Y#7W+$;/W4^:8D7&+#^KAG-# JJX97N/7^N9M?66^0!XOLL#[LPK
PP5'S2-9G;4%3WF67W2QXD4N!MX$%3S+7$_8Z7,6H0N%[/>=S;&P_@R@E$3S>;>4-
P4K6 .#U*>'1*,AO>@/B6V8#UR2"31.?'L@<"%T-BI_D#F3KJ;>H?O2&A)'6:Q?L\
PT!^2#B84RT?3R='#X95_AP_WNJ53J:;[JSU$(2FG%+'0S"P71(1< *CH":FJV>/3
P3<4X93/H-]EW&3;.FUU8H:?:L*X$G]W'I =#XG<LO"M-03="(W9L<G-P:].-X#17
P%9K"+[H$?@_'JUK=B=-DR=/4^1^*H1:Z1>P=72T>D5^6%/YI1O@4*,D=!85,E-*#
PHQ$*KUZ(RV(_2.;ZIKBS&\D2KL0-J)BS8Q--VDO@!93.\AO%I"MKOPPW:^I[2P3!
P1^KL+.'@'#VJA34NH_,G4'R^/>6X]H%H<+R2 #J]*;,LGNT(VVG@DE7$G?G2(4I"
P[Q/Z<E4\M>Q!Z,D%8C S7\2Y1\G= =@SG_;U6?Z$Y9MF7>9A?,LUK<.7PE-('&94
PV3"0< "!0#SY*>$&'.S?#JFT$#9W:A\6Y /'*5+$@A[CLK)\O=4T(/,9U<5,1(<_
P61%'N!$=1=F]:IFS0C):3ETD5IRFM61G?RII:$2=9V%Y9>K#)3=49P*GX)8"+QTX
P$0,KV.M_M0=E3#T-D1@O72O^D@K8[^K=,0&32R29^7VVN :]-)&P@>-J(*+;3[1]
PJ-. ]9&GL!2C,W3Y1^LMK/39/O+,<Q4M-A3*Z;]L'OWG%$GN0->_(G%6YAH!>\:U
P/()^"X@+$KJZP_YI[) =[/&1YC4L'<Q;JP"<LE!3F[A"EI6VFC(L!_E' R326G9Z
P NBROPEEVW3N['!/2!A>QJYY:$>9MH9]83DP7 DLN>6 4@'2@A63'?8=,QN&.P<H
P'=54;BBT;A@"CO*/]-F]ZW97##=M\&.SIR\*4>-]89(E[RO;])#DZ3]_?S4+,[2/
PZ0W2;ZP**@K!2[&G7$K+N*2\&-,<Y!DX4R@+*VFNC*2H_>7OK*UO'$=6WHFV\ F+
PLLC*"PNFZNV,6$=F#:615@(H=J#9D#WO^O.E0;$/697\#7MA!'9=WS/'MRG2296R
PNG,26?]J!(3-7@M[_^<+.8;@9SOX?DCQ1A9:?=81X!2-85<[9I0)DA6;>;!=#N*?
P?AN?AVH@_W*U+NTV1["NV$[,=;+/%+'U]C;LL<G H/C..PVCMN-N7))#S91:3YTK
PMT;RL;[&X;H!US/>JB<JZ*P7M9 KC! V/CK=K$-;!^/"^7F<D"*LFW@ PO\4U;K[
P.T2)Y.D"-!_'/3=1%[Q?40#RR$QT*<3[*Z']E+$7GL^K7?>\U-J%='_C'X\/E-L!
PY@7 4!1V:>:- ?(C#8>1IQN3@_/$@]TBS6JLSN"&^7<WHR3QF57IX6E>TWLA*Z=G
P<\GDQ!ABYY+RKWX+I2QZ,Z"&& %:C?BY[J3&>*R:NHP\0[=A$^0%8*AV/(F@TPIN
P.\WQU0FU)@8 0@X28]F,GU2#]%^]I"C0C8-<L#@HX_8M3I; >JDYULZ]\6%+E3W!
P%)U^)JL0:D]"D#PE\7--SNIY2*\]CIQQ6%W?0-YA4EL(U<B^,G\%J;L@817:7S(Y
P<6806N[09'Q!X1)=7!Q7>/H[R=>@JC^8I$8M_=JI?P(BEG!YT307$QUHIE1"PS5/
P,\PC;FZ.T#P10/J\,X4=B!4/L1V3G2%(,PN!5NPS-\S>LKDFD7.>R3_8]C(@AOT,
P&Y#1"@3 ^FM3UQE8ZV1"E,L$Y=_+8/[_GBSVP&W'?EP>=C1@?!L78LE'/%>EZT*;
P01>HFFIJ22"+@VJ)VHR9C1M5Y<N\$(_([_1C4M=)[=Y6/)5&[Q4LBGI8:<+]B&10
P[5'W2-R)H!\&U=#4L,FM9M?>]:)JO>4Y-D ?;OH&31*2R0$.A_JC)+KYUV2+D"-N
P.GYXS&$46FTE6)-B()PA!X1B[*1ON;)2CCKQ?/TJS#&TOX0^\U>-T-0B##Q-D^2D
P>F/&\X[;HJ$ =(?"RDN?_,2DUXV(YCNK(/@Z[IBYQ&2<M\,D@"ML4*=6!YNJ[-&=
P? A(7_GMU+%2^6Q*@LX)C=Y^9:1"-74=/H4\BA@U(]'1YS:^>)J*L4GZL]_>4<X4
P_-O5;/VK76\A_8!"(8BD7N>I:!G;L"8KNXG+DSO"P70'QTX/X6]^0ES.,V!^HY2U
P#\HVQ]KXC]U'?%&*%6BJSAF>86LV?Z(VKJ.L?X'+@2*!J#I>#J2K(IIN"$/M^PPO
P__6AA*$Y63;Y=D?,9EC_3O_/QD@OD/M.O[&^7]_Z"J08],9E/KC^^HOO(DY!&D*V
PZY%VO\A/VW_S8G)//@NY>Q(^FOD*T&S!'#T!I8*XD@@U]79)U0;YW=55#L+>L#$;
P*K$UM)*6&Z-'$#RY @9*X][2#<M4^TR[ZB<W@>.0Q/X+U"=M,3<C+VKQUBJ#6Y1<
PS@.+?65\%C",_DK(%<6!V*X)N1HPY15#N/A_4=A!_L]E>YGS9".DA7@NEQO%H6Y<
P@.<.0&](.!"CV='\DJWW[< T'9BQ9O6J?F+P[?[+FB<UCDI0W)AJ_KS*83@PI:PH
PWRH2:$PZ*/W:).NTV+ Q[X&WKTDTAV"S1YRL6:7)GP@N<0O[%/S]_GB!0F)+$N%4
P\HQ'#3Z1=N7(H>; 5RSVK<5A.ACA(^H9:X@X%KR\;:P[=+5!FK6L:!?2#)AI';9W
PZ0/0SX:87FECZ2#2[:Q$*VC_5A1MYY[2].K!*F&;L9E1I56;R $&<!P$1]HF:X^4
PBJ/'EL5ZYRFX>2C&8SPH6CDD*MVBD"F.;-;'J1N\N]VS74NZD%"C)UUS/4K:H L2
PB?^.%8E=[,#NCJ1DCC=Y!P6#]4_8O=4'-A,6_26%N>:P'^3*$/M34'+R=E@8C.)G
P:!(;:;B]G3^1!IB--277LB6,1![L 6R]BO?8F^7(KQ@USPE-+@3T],77>B$VA)[.
P+D03U\Z\,GE=@XTI5@VJ'!&-&7>]B![+;5[YF65->X8&&F<>8IXQ?^QKM][95-R*
P6A_5:5#&\^S<9 C\H9"1!F/?I-#WHO0HU2?%0GP-R;KFTX7B[-6(A+CS4%YD=NU-
P[LW0IPLPF(IME#+&SE(Z54OKX$YU.&49A9S3W >MF9K##M_W$^.AQ<'J+>. GP]F
P<)6HOF#/-=^&@)V\DYL\9[."3A]UQLV>Z#N7HCY4/(1P">%NPV1ZSLXX&5@\!9:\
P4;WN4*#6-3D*HZA(E)*HQ-#0!1LD!>X2@P) FN>U6]&TF!I.]?GL M\S+,A/8XSB
P.I"VT<0N5&P0)+:U(VZ;BDWJZ%=V&#O;'^*R+ZNNV2SEOB:.>';=.,Z6!D+O0Y%2
P4$M]\Z?.^_J&!:E9<9-3Z*KWIM$UCW;>K'W=PAP5/".@ ##^YZ@/[L[;B:$GG_4Q
PZ[3_9%1KFVJL]ML&.9>TN<ML<G%>+D?4>74*;6P$5R"_N_[,Z%55:2#9J8"XAHUG
PRIX"6PF&Y<]0: [,12* 5^EB^JTYY5ZHV$=8#D[.<;S??@/M@15G6YX9T$5E#)XI
P"\T]V]CQ+XM5S.E^#KY"K')RTAEB1[5(L'IP-/2).]-XHLB)H[H-'AG4#/L;FO!=
P'S/^H/U,KD*3 ]&Q(9Z+'[Y5H#RV]/*[@Q;M*5 [UB\V"\>*VTUUE8IB]$&,$])V
P+A*WU9Q5GD:6YJU6/=LK!_1/Z2R0MGF_6W^&<VKXCC/)E1M\Z)<C$SFGVT-5M PH
P#8D.61(M574V\[FZ1=KLY%N(-:'N8Q)!4P&,^=W +/.6A.^ \.WMI[<F)%]X4*<>
P#BGS2608C+*JZ?A(,QX@T/[EB06>$?!/1"*8#-W.09P95 ]MR'%9#"I?$2N*:",7
PQ;KQCXG:OU=C)&(W73<][/BILBH,93U?B$8<=P1['^WQ+UU00N6-B,JR</S[;L4I
PD$(M0#1 \WBJ,_)J!U"QC.4]5;PV+5BUTWC<!.FV( L_ACUG<VG/%L1P#:52&F,!
PT>VVX"@5*'55.0 UQ<1FTJ&0QNVRFZ!! A)U82))/(-9VQ,VZ5;&#3^]D-LKG^OK
P)7@.^'FUL1WES6;Z^B_0.CU/HP (HHX8/\P&*P0AV-L9K=7-=VH[5JZ2#_.]K?CA
PR_!YHT!FK]7#)1W(P(\>/TS+W8#8W_J L7^N$&S3B+ J-*VL]3"&I:/%45-YA0+9
PNG.^*D/NJ\ZG'7@CPJ\UL(%D(S*\40^KV?/M:C?).PK6-D[ ;8U#\JZ$K122H;WN
P?38?J<_NX6R?CA&V6TI[/CVS^Q$HG/!_\RN&3U=&$2*,"!- ;6.W_+VT&H;9);!8
P92!SUDU$;\PBX1 2((E3JG;O^]I8_&3TEOB_$Q/I=Z6+PB?XPMR2=:^JR])LWNVU
P57_GB'%"ZA1=OTXO#\"2IE;S7#W#"W1*GOC=)1Q=XXG\ .OK6J$T[J:F&07K:[KO
PSMW[5IT5G2-0EJ>_E*M5/O,Z;)9P!^:H>)^'-</FEJ1\($MLKUT,,?%96Q,0^]KH
PQ:*G@HP Q#WLB-[ZX)PV1#XM_A.:9_VG7-V*MKVJ0+":AB@O#9OR81 &#1T8S7TU
P*W%W'ZC8/0'&.:L+:.2[+Z<<UBHB2VN0OY"_M:9E$9^,T8S?(_,QQB5Y*-+M66-X
PO]+JT2$'H<")"C3<7SU;R;%O.SD8GRM2[0N6T6TLC&9,Y;HK5BZ&U3YK7X8#ZCR_
PO3+ZD]S>N6&AY(>_T2MSP(/1EVIGSUN!T="'S43,_[I[_*]H4UF//(!IJYBE.R.>
PQ.$>SL WB[^_0Q=8:X]$6+L(L8"J=O)!]JQ<5996N8#(-.0?FO'X2EA%5/U2L&Y 
P8<P4;'9-KMOW2B$%92K2E 07%-;R?."D]'M'Z4;I!/R*CO\C#949@6QR(=DRI_5U
P319/()QU&Q"E?F/7&T#AIE1=H[\"_\?T.*D&2SG]U<8Q%3G^%)$WG^T)R] 0&FF4
PE&C65T$$_5M37WQ(GKO+^-N5;JK44!I!&N)*YS2VX8S)FFWSU<K@[CW2=K^R>!OR
PNX05\Q?VEWDM6J=XC8U.?A"9E,"'<4\4+O^*6M#)F,IP$OL?C@1?$@8KOJD*H$RE
P$*;'0792L+--(=6QL1%S&)QZ<M;4UH=@3-F20:'FL1*YM^PA3MAA:E3G &AK?[4A
PHQ,=,^/Y7(C&/U1S))J1HZF9>0FR2F:@17'BN"L=6.*!9>I-<[X;YR+3'XT;X4,8
P-2'@9JYL/U"0(=X+ZZE+[CYDUE$!G!;FGH]I(1XFQLIBE@['=*R8$[ K*D;+R[,(
P!X>IDA0J*Q> PE>9_A3YEFW.#2%\[:_0*W)?DDV0Y]PXD_XY:]AB(\8.P,(UA=E<
P(*U&U>0?] VC7HKXBDE] +ZL11BA0;N]]NH/X,JRXRIO9^]01VCEW+^\JOMKATC 
P/]$!O9TI,@1.0H0<]'TI/+)11^@ ?9S)Q#V]VHE3G&MN+ZZ8&D2OLAOSKRE0%,\-
PFRA%%,EB++AOMB8#A\)IWZ8;+#X +D 4XL%?X5%MB-")>F5M\14EHAW.5#IV91O3
P8I1GMI!D<NQLY/A^Z02R"(<*@3/!(5[/>_@_Q+8!F BMQYVM!3=.M&$T)?6 \#WH
P_-Z8@M']!TJHQ#ZAANI1GXZ.+R3= .JG^36<Y8\!:^18$'1]ZP* 8&UMC>\>FZ]^
P=RKVHI@24DSY5(1BKH-+4;R8)'!'1/!S@*KXI\'Y[V,9W]:R@_-CG2;:/R!'"(GT
P[7?H>+)![WPH._VBYU%@)J%$>=A47156RW \-X:UAU*$-BPQW@/[H=MD'D3;3 7D
PQ-(G<GL*J];[ 5R,Q5%:2H(CH&I557;^;2H.;7?EZR*US\0$D(7AM),ZD\=M.6\E
PC2+[I>+]AC#V@$LN:X& 2R'63]K#1[\H,13N>:;ZGUBSQIOQ8:V7/3U9'-#,0WEV
PYXKI6S,GS9H1,JZ$<IHQF /W)MY'SFH:M61K\C@_\P"$5\B\B!W<AC$(K8(0[0 [
PQI>9S+PQ>:EDH=A-0?05V?-I$!EYOV\4<K3TZF/4L.7%/() [IW%G"_XWIT8C X+
P7U=5/#AUI#F'.^L*4HWN<I4%>O)Z^T#5AC5:T?AJVPG14%(0?FHE64*@'UW'^2$E
P/9&2ZSM#B=ECP__<-W")@F1,?0MS7,BL0:LQJT_W/87PW@;N.9(@Z*L.STYS .0<
PS]3VWR4T'KF9"_QP+M$,;;OV\ K (DM5_=,GN!W!)SE%.5DLK7-X($^J3 N3,38M
P!QZ->'P&C:FP?)<@$A69]*'82/GDJ[D&&R!'<:#_^J('>V\?,O!,@Q.:\4K=4MY-
P0!4];?8\OAS>01-4=# &4$ATXP'?9HEJ\%]WH U^FNNY2":@N?YM,F'HNWJ^HC,C
PX!-4GX'G<->.>5U:9NJ%7:FZMWWO[<AX,*O5E$K&>%?)/XO4@RQ<API7-O:)< WE
PM,8*"NX<R[52(^C=R]R66<SU.<C]L,^;9M!GKH52@ %N@6"U:"' 1NVSL >82==M
PM@:M(%WZG_T.,11S,&JD<,9*<=6Y2^:WRPMJ&3[] -?.DEK(& B,^NJQ9\U$ES7T
PDC4PRXQ)[.;-PY9!P&@P03BE]9#6>(NA?"V][,"H-IDY68?M,5P(4"EY47CHI-^?
PB6J.L2\2=PZN,6".5%>[;(?N4:,N[PMTV0H] 1V>IF7 %]B)1@UC>;QC)/2=#?9 
P3.H^L4]U#NSL-14WN<':!$7[27R6<.LSHAEBUU1BC[+.K=%<." 7>CD,2$28OAG#
P:"/N7];6JO/6&CQ6+$-1-FTN91C:-_G1'ZDR.K/1B. :C%\<P<JI-(&G@R<M[P*>
P2DD\<!()FC^$**%TP8\,1]-X6H58 S=OC5RD"/HK3@\+^R6-=OJ )^5P2K2*8X^B
PQ8DDGE342;1PUWY](HJ]^=]^O6*$P/10IS06.-5)SE!L])RJ<EF;O!;8&X31\ 5B
P;DTP?CY*A:'&:T7E=.,,ZO7N'QD ?1W4; ;>&SO9M)U6@BR<F)P$M^/'J<NCSE+K
P+CQB#D'J+\?+;3[T-S$]0"Y;UTM_MI23.7S"(7[BN!<-W7[M]L_=U#(S) J<S,_1
P<PL3XD'WJU-[-?;94@K<C3O)&L;-01>"(^I*K;RW,"S %3W9'Y(45XC%E\@2MWG7
P^L[<N7U-F(G>BO-<^LBX8=8[G;O:T3BO56HF%8RSQI6QNV!. MS -2F"T);!*F"T
PFO//I9%*J_1(>NY$D5W-WEVI^S3A?F%*--=:BP>>:PGICNW\;\_8[%<"QTFI=8<$
P">D([YV1 '(ZT.OMI@J=<EC@XGWIYR+56U2=X]Z1G'>,5<PO2(:(D]ZF7%OF>?(H
P3J)GW"XJVT*]6.ZNLHMSN$_\M+Z :3R69)+J*IYNTREE$M>F^,6)ZR--97B/G-$X
P9_1&/^".+368KU%67OS>"I!B@41GK4T]*<.U>]@Z0&Y0PY[W&VKU!THH<%#C45L[
PR7 UU$-9YHW_@/B9#1_X6.#WQO"_ ']W&,RR247APU0D(/!/*5O4P2N^U2'W2K#8
PKLT5_*O@&_'C0:_-*($M3V+")."^J$)/VX9\\C]403J@@8Y[)#\Q92L%S%)?W'\%
P\W_YC)>+<6ZL+SO?S5/IL0=M>%RMR<R(I; 4(U H^2H)#RC?0QR#_7#@=5<?;EU'
PN;!S2":5+!^5.]>*[N9@Y<"\")9ARN/(F.2-"NJ5FA#1R"&,L+#92\ ]MZO$LO$8
P30)WW9 +E?FUYWG&D*85^\VT1)C5;-)!P#_X*15C0)<%NYC5-2:XL)>.L.VG8Z+(
P]-YD@JE6S&(-&@I%X\I%*KW?\M:#]'"'"+-U[*=C@2D-S#@Q2$> $:K""48DKE_I
P15IP3,/WID!HL$"<X0V=[V6#50:T@KL0PD,V=2UAYZY\;BT K;U"V-),091S>,6/
P4.)L!^5[ K9U4EDOMD89F^,YHF,\[CS*R W.=@/_@-429,F1B);\OU"]#'\9O2'C
PF%1E'2HT'<QVL8B)K[2>)@"/(5V\-9JS0=>3.\&9HJ\3'L'3F&D&DR8=ER>;,(U!
P4^WU7H ZI;"$B%A>X4N?"8/]ML]Z[YS@/99]$T@__@EHO0R*>)G>8YLE0)1%,^V^
P":ZB9RM1R36-*\G(C&SM= MVO#A4^CF;K9@)BF:?\9/?/J<$;,[>Q;W6A1V$71;A
PHE!:(/=L8GKJ3#]$>K- K/5I([XNE)MV2D7'^27@@!%D*3/(!)D.,1!Y92U$939!
P:T'O0^8:B),.%LE4_KO >ADK3SB$VP_G%DM(Y16A[_$&AP%)2YV^4#)K/FL@+-Q0
P3D+=W@A_R('KOZ'P#B]12@/G,R.^JC4:($@.DK^Q?FI+%7"DP BQ%GDT!SDGX@(D
PJ>LO$!,;D&&VSYL# O<(,>J=P*?BD\2625A06&+_9 :G^G4:[H2=A55JP(2U]B7R
P;\IR4%"O22P5;R-=@A'8P7WWAMW#++WPOA%UM(9QPQMV<-$0^C$8O :8_(9H.&"7
PS 7>2TK/LKDFZ\JEV?/W83\N5L4:72&Z@8M3G1,)YHVI_O[CG2@*!\ZW><):Q&W6
P:#I@R2/)'&D&-R8 !7[4]#=T!T[H6BXK)M:26V1*/U)RE-BL;S9#@"00:+:E'%&+
P^/?&#+3PJ2V@.U3GN2.6<KQ:9XF(QNG=T]C@W8"Z-.J"?!@L%8\C M#\/\VHHB<(
P%\5 RI^5@UWKBF?RQ;1U$\+0<9683.*E.H<1K".@QJOL7.[?'6SF4&&+=Y2@37PJ
PET\TCT/I%FURT0]'_T>6,"M+ML52>U_W^MNYU ;"8A&/@=K>5XKQS&*3AUOP)A/D
PIC_NC[V=57X-BL+#.SYY@U6-N7/_-T(0#W(9*?^_*N#*E F(=].!6)-KOP -:%U:
PW4I-'ROH>1G-UZ8IU0E:).$KV*54U^\'VP46(6H%2.2["WIK(.:DR)JON/4?DHSX
P_4F3LOR/]BA+TU=637YZ%"';4M9V9/I)LO*Y<8Y;LB-I+=(-B)B87<0M(PXL2Y<<
PIOR>V/IK#B!L5PVNRY8(W60$ **$Y^O/&5  9&\GE-!NKC_#UZ?VK@A**07621V(
PUR$-F]UBV/*G<19WTIYA67+RRN)^RXEECQ1<#[FY&_TK4,3)?8W7$K .Y8]WL9G2
P[C5NX&9N2OTL<^ELL['L IB&1F]06#XGF;MUX_V5=@Z6$HD-VYT,<Z6N0W294#6?
P\ZP,8/R) #V60%KT+D#(W@2%9YK&')0Q<CNPZ/FDH"N@*=JG#9-6O_KFSXG;T.GT
PG7]C;$-:H)BHACDH=I<=F*0Z7X<;C,=52]PW&/CB ;:KF"> 7W7\BW/6KR9R\EM"
PH:MWKBL4-@O@_8>BV/6FL_'8QC=9F3  3J47A_>0C1B;'1TEC!V(V8H@;.Z6A)/E
PZ$ !_)(MHS"<[/58$;/CC!KO)_H_:Q&P04==C-YNGJK/7=W%&Y8U1CD;"PNM*ZU)
P)3]R.7Z%T4\>2I(@1MGS,JX5XX^_Y+)<<4P@7!,;#-IC3UZEU,78" HE,N>B+Q3E
PV1PQR,<\>WU*R"QE\6V-ON%2/R<[)>R*";TY!,5B]$.EPR)$+3D7 (\EQAC',\BR
P+>G%+M([XB;L5T)*K9_ C_)J^/D>X/"47]O1)N*5<JYIXW3;#DU@@X"7-MW^P:UF
PR$LRG05D\NQMAZIU.3VY7[#9VND@GBN484XB?_>14%^E),M]2!I(P77GT4'Q/1WA
P34_OV"@7W(QPL"%3+O"^15[M!N!_;+ 5$#V[DZ%8-0\Q$O'OO-A&%_+RHER=%J=*
P)Y5*;FLB(B_6)P(<(/8*3-=R-.+/2'_5=A#70/D>5).A4=M6(W:I;C;^3PE-9).O
P-&6Q:L.KFHC:XV%UUD[ \F>>[I1+WN.9T?+]S%2*S[J?7UQ$55(]D7L?;JS,E%/D
PH.$H>Z6>T 0Z87S]FC@BL\[*#1BG: HU/J/Y9"*:@W\O :\U-.3KM0PI ]8RY""/
P?%\X':J6TT>NM#NF@0[O+%R1F-O)0S)AV%!:OP'#8]=)VW6:#HH[/X.W2)I@JQJS
P;TK!YDU:MXXSQ69=F\'[8>278/]5/Z?E+>Y\+26-?>$V;#:4_R49(@#@<MZ?_GK!
P4WGJJCZ]^_VIT09^L2+VNTK1%T2%*R"^>-X&6O.IZ#-V;=(L#E+A *+B]O%"N84^
PMH1<,OR70I#_?&$]; I;_ZZ)FIS D$3-G"#HZ4+DTM+,#GC1P?RMI$% S(S1SMH/
PVD'RB=_SQ-=,O1MHB6@N>.&H)9-]*^6$(51;P-IV7;40&[TR9EAQ:/D>ZL[S8=^8
P+VM"';J#;ZEN\( _]3N.U'@G_H.(AFH.)+I]I1;49A>K;2OUXI>BXUK?A>PO?W&;
P4T&6ZL^:M_H^Q0@?UJSKT]!#6X'RB.XZW<HXW*;3U "0WJX(2X57+$]\J]A(I#K*
P=75/F^<YV.HM]##AU\_3#,NTB@#5XCI4)DN[7!L?,[+0<1'84-,:JVA'(\!D_DMZ
P5K?]1GQ14"$[)M9]:N9,4/+#L=1@-ELSGD"UB!XNR[WG-HL?@7%FY0;[?WZJ!@SM
P4[/\B#@D[-2NR'V(?05-(^\L'Z^YK!KI"'IVAROA?-U^Y4OX9G,-<MCQH&<ZYXXH
P"X2^>NYI(QQR3:J*2!+:7=N?-:K<A?,\@$8<'MM\\WW3D;AYOP6;H[?1&G[,.XCW
P2FH)MI80#=XQ08D 4K =X[]#L:D 1?\MWN$%7XZUO=.4QZTF@/BKI9EX,RD)4&^J
PG;M%_H6MUAYTX]V*[S!KN8M0.M[.Q''9<>],EADA.T(%ZVP9<P"YM'TE7"M[RJ=(
PA7YC,[#8F$G1)N/DJX*;@A9O*_T!(@X3F7?JS_/L)MWBB.!'%S!RQ9N08L?Z785U
P'UB0!4;),;:+SC8Y*QRPMFK^(^H5;_^8U=L&CA0V"X0")U+U71^64\^_[/]4'[3O
P<>977I[5M#/;4T[V6LW5 P<FQB4$!#H@/X=])U%0[P?HMT;-M&W\ARA_EH#N3<K0
P3XJ>GWVQ'D:D[H2!<6B<E574>5?O_,N66AF#A$QB4L-[07>^<^@T2$:#/]:G/^W$
P MVX11!Y,3(5ZR5"%9;7?G8.H;YW " 4[L:4J;987/UY^TL()%N0M'N7/*CUC%]0
P[/Y4%Z&%IYC;K]OWC^[?4=,CN7%(IFLPOSU3DN6%&L7J273H4E6V44.^ "QD5KB7
P]A5U485C" ;6BQLE]R_2 B4%Y&*5 J/#&\9?AX!QJM[';D,0>8H/]2R!4QG?*.K4
P:B_"\"1)*D# SQ"RKIL^-1X>!]UMGO+DD72?WEI$*'88$5#41-[JD2^!%L+D!SFS
PJG)0^JH%Q=3Z;"R=5$B]P7S%F7&W]!_\G89X_[QS'AVBJIH9&]('Q :VG->2U;4/
PI929-[XA^Y):;-&RH.I?EG 7^%2Y%G84 ^6XEK_E*\9CSF"$6!F*K6,\3>7!-)<O
P7NW+VU:ID?RX%S<SS5O5E>!MEO+;0\ $/YP^58%=SFI\UX"4#:F3,KUZ0T_*4\.!
P7>5WA$)S.<5264[EMJNO #D1EI1-:L1,VC8,0G#"^G=(+UR_6+JU1.;9YZ&>NECI
PMF! :G*IW8*?>OW* =6KI0. 1P*L/BZQ.WEOM6;H6[_L:)^\(Y_IX6Z?"H7$]:&D
P"9\/@OJ.S+K&;$#X6-'H6/IE$^*OS8QI)G#KF8B_U@,4![V44RR\U\M4Y_C82F3M
PG3Z05NB]R -%:/L4JY<P' .)*>%$)P4'BXG_*^#C08V#A@51L?&^<LN</0$_J(U!
P3KS=.GPX4+N7Q;H:Z[Z_*2A7"@M@_BJW8<:X>(&LCA6E%ZNV(R'P3B!MO<<PB=@:
P;?3XF6.3#KD0[T??RH.A_5S4:TSP]MB358/E!=R<U-;1S>RPI 2Q56;N[\\XOHIB
P(IB!3FLZ22JDZ2#1%UH3VIDYR5]'W:KM0F,ZA^JL?X6W<>O>V XO9!J"!+OW"U6'
PBW\G*$N\"8?"2=T1:T;-[!$P1;V5OW&D9"$U24VMZVZJY*0/@,>O,([41VJ]EII4
P@_^A;5QQAS%BN1+/SRB17>4)>Z3X=YF;S2$4+2>N=8H%(JM?B7W>ZYRN\^T"_U*!
PS SOJ8%"!B%I4K.Z'F%S.D-5L53%P,:6<<!:K.D_N\@'%E>='B/"% ^ _K-VM4DW
P/](D.-J%UM66&:E6[_XDHCB@IADQ-L_!HEL3G%=^!75>HV!P^I-TG=XJ6&A'B*!;
P"+%6_&Q31'$'HB$F@[XE>@8%J:0>\^=+%IGZN!\+[J$DPJS+=N1V%8"/H7NP."4)
PJ<[_'1FX85FX3EW,AY_@4C=HQI&I)3<W0J.#5+%P Z;MG:,_^HJ1=.+)<;LH> UA
P^.2@.YV1_T^:MVDF8@+%UGHKF:=.UX&-H#K2<(?=2_4(Z<A>/C&IZ<YJLMMJD"'O
PQ*>"ICM:0"ED;>IG4:.;BEANYJW2(0-D?__%<>G'Z8T)'>O:V;Y(&4DK>-6J\"O.
PR_I1,=>:5S#AL^K&N,E[7H)2,_Q!\?UQ]&M73@(7&ZZ(!/X'P'%$N1^=&$@.,HR#
PT'-EGKSD5A]*336'"?IR&NF"5*$OG.HYY Z85M#E?9#\D_>L.\]BN#"Z$<PV$L4[
P!I5,7 '":^M-XX96\J$=]X9DTL;5%7I4\9A,+'D$]2BJ/:C+6W:FXZN@N*G%6XT$
PEVTRC G"\.T;J$,I1(T'9+/RIE;1T=M^Q<D_"_B"NHUS(!3B=@WJ>[%#1"C[O^)*
P7R/FH=W7=@:Q?8G$IX9\5L[\+?=&7JRKGTFH@KO#&G=;I%438LAME@J("'UM5#6Q
P]D0H!;&CG:-Q"9FG=@5'@=5*(2.2Q1^]E\#MR!+_Y:5K;0M^:FB!KFLVJR'"<E8?
P"PMRCOA)?2$S;? 1.7&L+4X&/_N/X1!%D;2(4::=MP6>A48SVLE 0.RPOD=Y?!H:
PY;0'82TH#A=[7^4,!=S%8&*#4.;B,G@&)W+;=::Z$$[\-PD.0.YM]%\!T6A<;C[R
PDV%\C6CW/<"QMP]48$(0$G;>FR,@I'[XY"0:0K>Q0-_0_WFF3D4]UCX/#($E%O*>
P7Q,CN&+A!F_JQ&&K9-1O7X.T,7WAT,T&%Y]^8+X$[[S+%C(V3S:+C$CXL_P+>_SZ
P%^#]29KF=@>8*SC?R^(V8!D>6(G;O(O;ZS++_Q1DTT_.@=+Q=T=(!+U>:%^?TP>5
PNALYGW?7_(08W6*\SD"R=R<85 Q='1--S0K^UF=#WREDV195OD*(</=H]'-]Q@/4
P;V:C"&L.#*/BCQMY(C0^H]3-2R6-T#Y'. !%HA]3>5LE[=!6AH/%H#H&!W3\-]YF
P/>4PS,733DD9\1?S<Q\T0"08EXQX(XU(A !)WEG[3<D.Z)8\5FF\H8O&@,1K6+>9
P]G]I#>RX(NMJ<:DK-1*S]Z)^DP,5 :<#/2=.?E?7>;CDR!<0;2MM]7I-D;W^X4<)
P\#33=S77-.H$@9;IVNL\:H9]1]<>"?");=YP2TAT*RX8@;YLEQY<Y=\S#0>'PO.I
P7"7&L"Y-(K7&X+O#H.5$E)LE;$Y*)!_UAZPM,MIM#M%ODD0C@'^PN];V:I#:UBE;
P4F>U*/\5QJK70+1(QVVHG448;8ZIK[_UY)X2AXB?,Y2!S676TI]#AX:X3Z84QW&^
PI#% =Z8BDF$_AFY8<]LGDP)"R69=4/A(F<IC+W]J!OM9]BB"-U(YF'O2'"'3C;M[
P6OYU/*VP8?R$WZ]^M!,Z &> 75!))[ 45*FMP?O?W*"WC<MN_<$13]D+JT]1%;N=
P\QHVV'5X:2!, N,8P9K);A;ZBBI''A"Y'P22QX[;_WTX9RE-&NIZ39@I)>IG*%Z,
P"+'4Y$%[<!C]U73^7?0N_-'G%V W%N9K@C*K=5@J6/1WS)=0]NBFRL^'_6HUCL0.
P>B*D_)D%@EO4G]8T]PS!E\_;I'P:]OF%27\ES]#UF1B8_27WU(VV-YUJ>8,2^B[4
P3/O:LGJ-9EF1P6Z9&NV@6 M@U!3A<SRN8FC^2('#O=>:[GMWT=)7DFL<08C9I,(T
PQ+@VL$3Q%4/3CAZL!Y_IU[YBD7?"=K&Z,FKE;8?W5P_86)\+:XE9ML@_52Z;[T_.
P8 8TOWW6B(A6)< JKC:63,8AY@]>+S<H*2-S%(%R:KO4VJ@]9SG"XT>7KW!W<%J,
PO?)$>*!N\5<34PLY,7XOA[MB[([4$#,=DH,UB\-"<!CSF<U+9^VSAIT<O9+Y<-.P
P/;?#S2%$?^27,#0PK1A0 %A\$+&;3?J/XE_IZ3$"I-'N[T.J),4)<9?'PEFRPH^9
P@X0+ "JW\JWY19BNVHO (Z-XK'^A]T580\]1F7*3!&:YRC#-K9@*)-"0KS&@U''>
P(-,E@>\/2FG6-;Y@]]X",!8)&XPKR9%#2\))F=\2L&=;VMW?E)'V+84ZU6O(*(CF
P%*__8".0(]"QD](-R<0P'1"6U0_FHJ-#\=F)":B,7K(,=%,40Q3844)LQ! #(AQ$
PI2)0XSAKO^KZW0*3"^90"EX?HEH:9FLVX\!#I@O$I(N%^#V^"@0IP\P_$3;Y"MB3
PM[EW@[\L0';[A.IV^)*!MU=VG)V,_DQNR\01.)N-\:X7S.-S*XJWS!LFS[@5I N+
PT4.F-4%.+7M#5-^^[6-1&D&,=]5#*(^:?@D7&1E>F1 ;UX_A$\I(YZ022UI7))+F
P-NQE*3B,P4+ "O)1DSA,9(AR3R%/(IC'5%+FS+:,3:N[X%]/]>_^M37E/%2A49D<
P((!C#ZXQZ2JJ2##M@VT1G?\RMQH3GDGFFBH##-6X*X*KLL1:D[@8QY$I$Q7V<"?W
PK%"2HB*]UWFX-^B_$1[(O?_S/ B3&:&* SP!T_"6^#*'( %G4 RS6YD^RE:#'3Q&
PH #R5U-IQG?#"V-[>O@%KM]F+%RP#+=,;2=>:9XS_*3,%K_!KKP2Q9_$:"SMG4=/
P3T):*F147?M"%][OM?SM_*HD!OYNM:#@Q<45\CS[L<#1$,.7"9[RQNEP(=+9H\RQ
P[F9VIF:)G]$,7N^,D%ZZN?;T]*_173J0<::_F.0XE'3]Y\$]V69C(C7<NOY!@V"+
P!7UXJM64G15-"U;4LC"6G&1 [#G5#M,(.3R5H6 ^TR+PXIK?@8T_+QG@]-#5(\BN
PK""T[84;E_$V).8"/D+3.O%^])G(:!+6VA ']]WK^-L&.*C$]T<_P_:O^P3J!AN(
P'[5-U+DXB1F$)IX4SFJ88#1.1^-+4R/%0>OJ*H5%(HWZ8+[4](]YCYQ46DK*A;85
P5LX.^$,NB_-]<XZ.C^]Q1L+B)*?>&9GP"HJ00/WG=AHYZ,LC04;OD-%G#<,7L R\
PRT(*+GF3M@$0+NN-$&U-9U8?]QG1YJ3NS,.\[=BG,P_/FV7K._E-Z3%2&F)&_M'&
P0(NY_$3QZZ\BQ(*9K@5#D<G^=CY8$$>324<U*IY1.N\_J1\TH9^^^[L2SC=\%CWI
PC$U'=3:0,6K]DGH5,/Q3$?V_?AB'L%NT^^2E#_(N5A5GK2_\;'!0 RTLXJ3\%"#-
P6)KY?3?#!!8%VN,;J=GQQ_?)XPN<B4"3E27D+ U]1.0?=8&+Q\G\H(DL'4\Q<J%6
PKU#+4QX\0A/B$6=SB5,EQJ2U]SK0,41KJ/D .KAB;]!#G&/?Y>DS/91>G2#F3/]R
P!,F6JP5,@4L][RW)RT:.\(JWXT_N'J\9^@0$ABB$@<!;MH0!U+X5;]MJCH\2CT<A
P%5CBU5PYI<MA_\1H.]L*U&_)E^#*4?H"GW=S\<RK$X/H9A[3*&SX30SQ&PWQ3N%.
PQ3+4&[B%J9;E0*$1\(ZT00/W[*UDKOQG#Y*;6%&?O70N(6Y\5ON+B(6M&RS7D<9/
P7]C=OTU18'R<0I;N_YQ3(W]..Z=4M[OR[BK!S5Y6]2W6'=@/9ZS4Q>'3DIKV84@ 
P4A^I0["U5^Z9&6\7EZ7\,QP18;<3T8M&'Y&41$]U%<*'2NT.9BY;.6W'>W](IF7Z
P<O<IR&*'^UYD\.]JU&Q+$%"I=#YKR'6RD"G"_FC7U5:T]@]=,RSMA.^X6T?N6GVP
P<[8A6J!\T?^,LT$,)):["\LZ-EQG79W32@O'55HU=Y#A!W(2CQ)BL>.Z^5H7,_Y]
PW9W2^4_&(**]E$/_A[TRX7?WD">I:W71>23FB[+30DO(WZACU>G&Y>7/(3T%S[TN
PL\,/5I*&16_F#.@LC^#)\0Y;85%Q/6L7^?'#A0[R7NN-="A.7&OPLW#Q0]+M>SE\
PC\QEN/ I#>Q+PNJ.B(T^J%K9'$]#ZO>)+T(LRD*9<B<CPNG5 H"*G+O!R_Y04M'V
P>B?:@IU,*!>ZOA+I\8ILC6H;BI,\6/%+\!.&EBPU\,\T(6PX:AL U;I8S74@SO4-
P[=M._"_SYYW(#IZAY?:ZA=6&0>80T!O6R%FP#XZO3ZA7U\.OM-[H^XQ@Q7$/5(?;
P,#GPM[Y:9MNZ#O<?)?$#A-3.!![^MK?>7Y>S==R]EZ( T)4#>4L"F)-6_[E?>/XC
P/0,E$BPV.HRI^Q!:H02>H@O)8M%=!-FI0("3]@_?TGQ<Z1*Q@-('T'U6$<Q_&:(R
P0X&.2K$'^LM"A*;UOB\=FP%P=L^G0Y":%G)MXTC!6R<_LB<%E4$:Y;4WE&L"C."W
PA2N-7H-,"-X3];9*W!$:0*4#O.BRUEF"G,NW]%0[P'4V-M06/2BA9^=TFD@>I@U!
PW7;!?&YKU<$#%37XY8'=,:<\H.N&NB_: W/2MFC?Z.B+11O<E,Q.$V7>O*R_5[^8
P8RN*O@2BI JW;0#=VW4TJC8+Z>20;\'_'5<_K?#%ZH/*F=;M#@&=,5E_!P<8-;>"
P6\,56_<[O::B,>KYZ[]Y1G79SHBT6()(0;=_49H':XIL(TL5=+TAX9&E<##ZSV)S
P&5;(VG[82Q'@K?'=\]1J89])]_4LFC<N4K96T$/DNJ-68(=[8_?"@&PIE;J8%8.3
P"-H.\)$E1P=^8J1%XUX:I&=/;/8:,\8Z[/QQ'4%_/'U#&X.K=\GD?CS+@/YBG8QR
PB&:_B- %^ 1WEVW.8ALY*YTT$U=OS>^/#T=26Q6J,=A$#:\?==:1P\2M3N-Z(X?Q
PO9V3 B1HNL+-=\ <E\BRKS83<6>ZIX/EXG"X+,T4F!>C[%9OW2V$*@"\P6FM2O)3
PKJ0@^.9ZWA38G]HC8\D-.LC-* @-VQITO!'$(M86.OTP>2NQ76)!9W;>^Z4[ABN\
P) !^+M7QJK<H%\+MF#J!V$1>#6FC.8TI7PP6>^_\-H;*O8B\0DD<RGDL&"58]:F@
PK2<%/W-82)S*PZ)E9H](PE)':&PFG"/D4I ZF^TH="/P&O#;?)FO?CV )7D,&&70
PK TCL64P#L*ZA'']ZG]KTIA<JYGE>46)7&7('W5;6$Y:J".;DE,PR+_P_8$A"6)[
PG/YZU$'!0 B(_*XJ_0Z0#6C57"#F-%VG3HW3='[9)$YS(]@_'J>P]!K$$(4,-NM$
PMHQUOGVKV3J/?=&>ZJ-]3;8GAC=%.:X\E]1@&TNX/6[-E1T8IDY@PM!U?\>C/V(&
P+N-:9C'!G&2MI:G,<4+!"!)^T+<-FX1Y&216U13\4;*6//K5=!W%8I"C#MW4F,\%
P):A47>X?RR1LH%P.AO<!;51A$HC+VUW7GM]E4MI"8<P![=V8)EHKLV7UE?GD& QU
PLO"CB0CIE1S_?];N+O<<B6UGV&L<Q<8QZN&/5I$3M4$DJYS*Y[$1-B>+6AX[43!L
P&A-YY/;1H;I<9/DY"=N_G'@!6;&B..HPUS)>01Q5>YOICMIRFY8?#:K57LW/H9C5
P=ZBNJMS>*?T@9WA/E^EL_ND&%J1]WAJNSS ;9SMB_'5H&T,4%(YU=,<ABFWM$8_D
P2A;8-_X"(7P>PT (_4Z\>5&2]X];-I/*WP+T4VU/FPK2O[?T60B\[*%\4SJ-2(_B
P2.3%[0SFZTG[1]YZ::,M<2\%\4\84U"E5=%YI;H#?C]$1^I3D25AZ6W'3-E:NH.]
PV1GPR04IZO]0NW0^HK#0C!- BQUN?2[):FC" @TD244M/OO]Z6<K"X'D5YGMMGQJ
P!4&UAQ&GIWH?-8KF:.1B^4[B\K8FB5>C7VG8<%VVQ K(,*JGX -P,%.<"[/>9)6#
P)TU!?K!/!-B'6]3I#?H=3CII%_ YWQ&5-"$2V'E>BG*[#-,V0WIK!=,9:"_#X>L!
P *.068,3C_G-T* RQ6&<W(+?UFWJGLQ<_1($ 3A1)#EYTP(G:ZNOCI_P:B.H2U[;
P5]\2FY4L(1JKCTVU3Q"Q'B#/5IHH '=2>JJWG=7+=3%SL=XA*$HLH.&ZI>!=C:O&
P)KYZJ*<=J#$OF5]P>S"E34,"1!@X_;2-2-EZPHIQ5IW !3Z]1CV<)KR?,E/NL7]=
P$A9XJHAF6-\P ./ ]^Q?NMQ:ET5?A#V;R3PCO7VE.+*#U-%_U3VIF1MA"R"9W@M"
P"':*Q9Q&_#0KB\G<]6ZSG(8:YDPC^\HGMZC_P0)+EE;S.GL@@)[[:,YY=&5&>;9O
P93_)!5 R8= X.A?G'W\IW+7;;\UN6TO9&H?/K@V-4BWPP:^76653X$E#YV=&3^ &
PA*9S#XCH8&C-IJP$3DCUH[]*G%\K1G GT$*.W ^VT!)^Q!T_(ZKM59+B]\UZ0@0T
P8TX4XU=#-1N]ZU.&7W;!3L 8MELY^'*C5-4Q;BEIX0<(IQQ@KUCXG,8]J..D":L_
PN0>CD055TFAGYO\L'J _G:BT-CA $?#OWAX4Y+/87P3*#.SR@5;T=G^^H*6_,KH$
P@"7)^=)8S9FKZ[]L# U$V*I/K! Q"+^X"_]'#:5O<RB3/[-?EX,O0;0S.YJO9C)'
P]>M%J-6= [ VW^=>PW4LB/OG4/2+\WDF30.IF>LRCOAE<KHY)+3!(*!N<=H)0S3#
P-KODYCGT9WZ/Q8A2-U^[.;@L:K7EGA :%:B%A=><1?ZM:F^&#]]7>W8$^AD 5X:"
P)*#3_=^SJG\:EL\**(!:5(L+/P3-3/Y,L]>QA0NWYKL;BL3?Z0_8N)'-> GZ:]Q0
PR)H*=I:8R2!,=+1B*</):T*,5Y_C%BHAU$<(NSA>"3Z0?2O[FV"B?YXX8)Q(%1K-
P/U8I<IB&QTQIHVGW,!B$ILY>65N-"O&"K?2#ZD >2^K,UGKILS9Y<"6L\H*AT%/N
PNUE?BMCW] 059S[":G/ND@.A1VP,B+V[<@XT@T\^)SW8.&8"G.B>(F#+H8_,9_#'
PI*# J=^XA?"$<^(04;#"[;4QZDQ)3/*3S741=/.S$S/X>'+6W'CO4:1WK8R&YX?9
PS#YA&#R?</1Q$,'"IU(:!CT.ZN([B].%@N(,J%#\X(7X)8I5:H+K+@^1()5-KX(<
P!,SF#/:"0N3+^]^\Y@52<-'K&?-=K_ N(32[5\"Q#R=NU?'N(@D.M11K\(#](URO
PT30O;0K6M^^%U]_'4-W>[HU[=BK)>LP+N8BNQ&S(J;7.O,'B[6QV#I'JA<%&$P'7
P7>RV/.?/(&@_XD 9)^0$>=[3 R_:>'3HF+)6.W&>*)]UF%=78H\S6S<  2+5^]@N
P#V]3,<0E>Z_%CN+WCJ,I=G"B3!&='I#?W0.6X$X+B46U!+79KM2P@ ]M>WPET4[>
P)O6IRYP"D6D+]XZ!T<8?GGZ8:5]=?]"AX/?O<]@5-:\M>U?A;)PZP,AZ0LX=SAI&
P41+?:\"E>#W*)50</9/YD-2$"$T(X_[NW'R5(S>[*>KT!+?,.EM![I'32>8+!:%,
P33@5L9<)Q^Y]7K>RO#'WT'RF&A(<[\8'J; OW[YOZ:Y">EA.\6@VZL3S\J2I^_HR
PSQ52T=!AA--(>9-&FV)<<]:2A^.R7?%EB=/ZFN$G5<F#3.4\_#O^L$_K/1B27M3I
PW_X-11]B,*VMA=4?PZJ.F\"E11 T>UV086 3'C4M'=Q. V$1[#HC16/5'<^IK$&(
PHNJKUP\I9GS[QT-:TJ9*V=F:^L&+4I1@-H"^J"W:'53J_:^P?+Y84;"$ E@F8Z<3
P@O':P'/M5P&*[SI(P!_G2UKWR@0;?[R'# ;QFCI)"W_>&R\#W?%S_'HR;F@JN%T^
P]!-;"0^NU$1LJ)XS?)^7"B(1GJWWW8L#^QJ$***RSD(L&PW(=#14WH&UI,U-QA2T
P1,9-:U&A8=X9JA*PK[U 9YRG-G\[TA)R"9,_L$B9@-8MX8I[,78*1$B3 'WTX$G/
P)LY)1YV4JXCD./A,Z2P%$+KYQDUPI78NJ:&N%^O;S"B^Y8)#=JQB*Q_=E^[4_&3T
PS8@E9G,8B<5L* I;GNE]C$E8$Y;,&'>D!4E3P+@U5B]IQC)0D0S1I\P:H3BT(J#)
P'7!T]EJT!&JK_5AF7<COYA;I1V]%L*PPCR %I/B"DT6NFG#=&Q5ONV?E5.=G2O2J
P]D%625BE%D[R+XZQ?AFST;8?,A_/_=_FTJ%.QX$1IM*$&B(BM03MK),R1?"R9J75
PM)%'BVI^MG[,6+P\*4[ :/[?(JE;]Y3A4$27K%@H]<BS?*E<>:6%'9$P:NRRERYM
P;QS:\?]QH^!^"K,C^6)0QN"6].HE# 1OI$J'(:G;]&-?,BIVB@0^6QP>&<P>G??6
P(@),-.(@>:6Q:[]:/21+9,4(GU2#6HA<:UK#3?\J0?X- Q\S9,3H%7.8>MR&CN4H
P!V)H<-SXX@F(T[Z^XV$L580BNM+1EIB]^S16&*3NDJ0H>7O1=34U2)#\N* P1]Z>
PP@)*YJ;^[-.4KF)"]X%#]7!I0; Q0<N'00Q'Q*@EGLR#=I?]A)4/W9&!S)]K+/,,
PK":U1CLZ0<Z\L[%EMZ8X^5PH,WH)@@.OGW>IAK JD6O#X]U)'#B -_QNT#JW$C30
P]R*RG^&[@5ENL(:WHYW?)IJDN+?)=AL^L@]W_H EX'^930QJC/:>'N"G]K^TZ&VX
P#2RW00N?WOD?RD+^@I"<2$B5TC3DSC4/-)[5Q0X3OHXAI.=7;LDFZ"87=AADE.&#
P"LQW#G,='6'J*;^*X93!$H0D]^^OP)V<'-<T#P2,_W^B!5Z[#AQI@L;>Z:K\V$ R
PJUV,=<C':FX"HP85Q%E+Q?(LCM@";HXI5UY;_84\E?V?K;TM#Y_Y\5N\-'IJ #8=
P>:4-0I$FL'./0N%7M\6,FMOE8[*E:N8U>QD-C[<7AYJ"0EW'/E(9_S%*$BO*)! 7
PFN+?EG.*LZVWGPQ:+#)J$ 4_*LB@'S-M9+"ZJ^]E0<GK-ME)PO=D.#28\K$P\7DD
P";IT0^$1:-[L%(# _"GD&[$=O0&BG9B2(HKS]_^!\RJ",ONTV/RQI><NGJZ;<2"7
P*+Y:AI0U?>NC(L0NE;4D@%8A*FN\DD^#UN8N(;TD- NKJGD9)T@K&%S*ZU."L8XM
P+1&<^15%G@88] 0)VJ@"]N+"D!8H.FK%("RR3G1D4X&2[2H]4/@+9$'HP2@^K6A,
P!\E\#B03BK[4S(NC\<*?#H]635_0G7-5QMU-J5)D-KC#M]+.ZPJG,-7#1.NCZ$\O
P^<*!$["2+_XU]?M:CHH^^BKSW[CO;M]0W%B$3O".D1/]5Q\2\8KI7WISA&^D#/(9
P.@C6+@]QF- QI[Q*;"0:32>$-1#D)Y'RV6K/",IG9E1$@71:Z8]8NH+B #.&-U#5
P5M,S#M!^.)>D!97(]\#V X4IJ0CLCCU% +A&%))\4LZH7#E.;I#%7U/>YD%JT>8C
PPGR/ &+[72X,MGH_W]>E#2[NR+W,V3;L\2^7V_[AE+K:/F:+C@$Y78JMU];"Y.!#
P1DH@0+N:I)F%Q9O7O'HM) Z5P-%FJ:/V'R-VX%0D_$2YMNF[;[J-0BE]-0RTOP $
PEF3\YB"(^WNO8B$5%99MG'A:QL'<20.6,[W\HH&(QE7IUWA%0JN8*X&@P=T#%JOI
PRO5_&I,%L<.(^O@E^OWR[=:7.?0ZZ"_3;@TT(^>TCX+I;]8['60;S9_/S7>I->,U
PFCMZG=I;F;[TL!KI!6WE8P3#$TN"3:16<W#N"FS&7L3D[[.W'9&F<A*35QKHK_?C
PV5ST19LU- NHNUH8_:]J(<><MU1[GU%:(7N/,Q'=:AM4BOYQTFY;%QMT"F8,U"O^
P=^\HW<6J8(T*-I<N#+Q]@OZ;80B?\D.@ [YEW[ + _@(<?(SD,?%7VM5[/3;"6EP
P"MNQ518J=^S9>K76.R7G1#$I$2XVWP0=8L4)0>FK4]WW%I$>,J)7IWX4ZB2,7-7>
P4')\8E?TVOXAL5T*08<Y:P/24O0MAZ"D=C9HZ:8#3MW]U8DV;\K296;+<S&#'JK(
P4BQQ#0.R;RL+K;A=4-#3^ ZK0V=D6EXKP!,4B-IYFE#,FG)"C<<?Y#O!(XL--<TT
P]VF2X[F3O&AY$I?G!JP3<3ZBW^!#'=?:CZNA<+0.!B/B,3W99U^D2TB)>%94,'PB
P\K$"S*=<?ZGR>"SMA402LZI$1DP2:,DX*NP1&>J10-:=@-(03L<3'$ X^S]@4@H)
P0U\W-3138HZLJ@U==,XKJU-1 K<4I 5OFX*=-^OTZ(7\?_ /Q]^8FK(<) (JQ^M 
PM\]44[TV0.4R^9DF&=D]12^T%EQQZXL@R*_/-"0\B%(+<>DBLW9SH8;S("P82@S$
PTEQPEKUP+\^2PQBEG;O,5@HB\_&IP8&%'$ZFS/ZXRD BV5,AU:'^5.3S^==?C;-P
PU9BV$WP7&RT=L+>4T^@L'Y4R?*F^?$SC,=EH&/J/G$4QMIC_2_;*8[#JA-[WW'AA
P<+MZW./ "E@\&8!%8(,6@UNUG5D%>NE?4FLX#*?>'?-#C--VLM -P,\'2COI+A%!
P)*=8)P>:,RDHHE >8J7R7-8QU[#"@ $A!_.=Z_L\#A#(?-V91.%MY0&GCC"J$6JG
P-*1JOI?FI[XZY/<+=GLM/O;"38QU3#*D\] KU!)>C0E/!5[KVQO7$0[>+^VJ>V,$
PF>[SAS=8+KV3OQLN0'$Y@+1B4Q 7$NO6V-;AK6H]-" HZ)_ 1W7 @RYY''%RS2S0
P*&^3^V\>=TM5.[ -1<IH1PVG 0Q4!=QT[%Q>W8G8^AW=G/L6Y' *1<D?V$FZ7>'0
PML*O>/L[[><\#W.\]+;9F+JM1 ^E>#YKNO:*"<Q<F^QW2&ME:XJ+LT0W5OBHT0ZF
P>?7<J[EL==G: *17];:T2"[<S-*-<1U[]<<A%U'!%BV=S%%L\N]D\"\+J;4XG.[W
PF25W"$[>W8N% O2+K3%4SG-^339#W"U5WGIE4!@46AND?;ZEKN@*F$Y_D@!;-1H+
P7P-:@4DU'K[R+Z=_,J1"A=5R#P^LQ(DNJ00-LG=')'?;T)*()592LG/ 7RKIX?KD
PI A1?$DK_O._]AM^/9]BXJ:5S=KXGC(96LSC(Q?Z_/V-'VLNIS?]9UR"0:@^?*GE
PM:F3Z&&5%.F38F" +628;00![*X58RDI:"KC2B3FA-!H;FPAKA@_>4< ?M)]JY'0
PE.0<U;-U*O?]<S]2E4QBJ1(1O73$*^57M15J#VL]Y%W%R<;?[V,TA9RFH6+N>)CP
PZGLR$1%'1"(^9"-UG5__JYPV4U0)J/XY<O7--M@Y\*],9T3"K3>Z<8-VK19%96 !
PF@W0[W@+0[-*:!1EXER+8^@32T8-&7?RTG+'"_8RI]^&:,UTL?^)"GOJXN_<%:6L
P3PN-1X*'61!,'Q'>RM9GDUS_L^G\L588U5QF"K5H>S>:DWK6L+,(">YE[A="7V8]
P%"U--TNFA.[$1G6?W&H+>*&0C(3X%A8 I8$8=E3-2&)&VBE)(GGK8N&YRP+?PV1J
P]&6?9#A5?RC"?!_)BB!;0?NTP0/]ROK"XT_%UL8^5?IXT9''C.'FN$@*AQ$%+UEI
PQ&9W-K ^ &\446(;S*ME/WM2!(%.[/]^$)J5/8<9T]M\4[G2G4>?BFC!,\^[<DD+
P5OS/[XIRZY]N/85/V^ SG!V!4[@OCJZWZ0*2]:-^B #'1IH_(43ADLNF+J]YSKY$
P/,!H^1(SV/Z7W<BC:-&?%1#;$7Q39#ID",://;R]<6P\+2_PH/P)[+\YJY8?OV+@
PJ1_^V?')=@? :+C"%#./ZF9RREVPJ%2Y)AP3.<$QN3R[Q70W>X%=9H01#==WW!]4
P1>K!HRNODXD"\VMC/ES5/I)0!RK*3B>(?.MFH*OP7R)EY@CB)]5A&@PLP(:P.DQ[
PB>Q:)I%NXO#I'"(%_-G8842Y4!5DGD;2.2(=:1TL *YO69KRR*C5KEL)QBE& -G\
P<$7I_9R1(AC.LZ+%JI4$,D:PA41CJBOZ[] H,CCOJV\\U1<O^@V)%N\XT3F5Y^_X
P_;SN4BS,5H^K=E.$,W,K2!\1:]I^J3KEHGL %R%Z8 -2]P2K;J0BMG^>3W==&@6P
PME!P5*"42_4WNYC.UH3=GZNRJ55S:ED?5/83DF\<G.E.JFS7[>\*EV\SR\';WS%1
PF;)N/!/P?3>=J\U1W-)$/BXIJXJ>U/O*.E8?TH['?!WDAFZ@4P^WXMSXM/.L7#L!
PMQST/[R2$2YUM4P6$&D3U5/Y =P/'+T2\63,="E.UF-)5G>J3+8H*"5HA;QF0M>J
P]"&NX1UGO=<B8?P::.DL@Y=!WB@65+V(#DF*X*$CE&JJ2;UK#_:ZO#?W6;I>O(W6
P?XGZ,I0)B:#4+<XZ_N;R*&]R(\'TC^S3=[![@:I45ZB=Y]2A [4@OJ/MR+(@N$[K
PW<C@EG=""3EC3/A'2@N2E%CLI]KE$&ZS57TKFG;K1N*#2C_*$$/,.@X<PS>/O%*V
P7+J,67VG\]*P13:"HFG%+0$5^H-!8GYR'/S"N/+/;)X'#9QAEN9ND<H9'SEF8>E\
PIX]\F% NB-S;,GRFX"JWQ.L[HF30 VH0&(FI&SP%=.699ZPH;?EX>\2E2AFMT$ P
P,)^D$D1' ZW1^L>P>^RG40+/I6A;EJQZ-!\[;T7AG$#<AW#*Y&5PI9 Z:6=8$[R"
P@BI/,Y9G";A:!(\,\?$W1EK<Y=0K1#6:'J+$I_7EW!DR5S;5U[\UQ)FYZ(8MCX]S
P2(R_K<_\W.9'U4757??76Q?E%.U+-^"JEHP%0(NK3KBXCX*JV6X[0G$DT-*I;TBT
P19XB] =O"B(/[$*Z6U^]MQ8N+MW>?]U&K%:E,6TRX>E7^948K^<^L+U$?/+<M)X6
P)I9E+\'*U0H3E"(U?[C\@1TL5-DW<,YE&P//YUW2"M>\@+3$B]MLJ"I^:M^AANHU
PNEK;B<3YFV,V0U<,&&/11P;_BMD:L$?&9P])I1..K:EI@U%K8B0D/B7<672/,P+]
PGD(Z0WJCVO4?'?N2QQ1C3MG?!*KT*SU@$Z1%5I2Q>+8Q/GF1=K&.<!Q(/E%5UB:6
P7ARV\'6]5E0D*8TP/C"#<X -J>K:D;UJGT]9YT9KV$J*E,= @)-7<SS"D;\46^V"
P"VQH9CZ6"B^X@V8LA>,V["Q^4+(Q EIA!I ]EE++/$('U6[E?>;:XM]K)18O5HZJ
PJ$,(>]@HW>HSE[171X+ KC[[MU:"U8HD>]:J]@78]JNBT%TZS3 A^%O;,HI$U/CB
P8A7:FUPS5W/:F6\6MM=CG>^][4;'8$+CT<D06/.J&)[[GJ<[[BVVI1.YTU+PK\A6
P-AC!=>Q_ '_PGE4^U]A$)N3 !(<3R"LU().6RZBW5O5W7RNF2B3/(,9C52U$3%<:
PB' QMS,$"TN>=^&P5;1*T5X-ZW1@7YV@?,.YNDO\?#M80P!ZD.0^FKL,X!OOE[=F
PZX),1I"9AMCD3>!QXS CL)<;83:1:8K3K< 5XK!=<^D21?JV6MX+T_B*<'!2TM<A
PM:\<.],UF+3<+M4V5X[%$#LYO_ZXB^CN:%2%09XBKEB_$T-"=,<'0:#BC53RY8H&
PPGT!33L#0*T/F2W:932>4%T<AZ0YW#,LT]$\<Q:^@4:C3T!1=U^Y\OQ53=;K% 7Y
P8REMJH"G@O8@';GA9G=W'<L>F;4$0^!\=2H.V/<E'F-H]CG-0T0LH6X9H(K6>?2!
P,W^^MM:;,)@7L8:LUH<T,[:BSX&GT%]H9Z>#^^$(PDJ]CP\N=#YD&LE$E[$FB+N3
PO]2X]G;K3H+;?F<GB@9\'M**M*MLK5I98+\4@_2FMKN$UP?F42K+>("G2/'/0%#D
P*Y/C0J()8MSM# 4?2QGGW$A/P'244AWQ,9H9W\?EG$LYZ4*&!HR&$YJ 2!7>92I@
P']:Y+8^R+61G4%P/ELY$04,EHN?!H#*C=)OZY.5$BP0)=X?!!"UY;%].)\Y->CD1
P:I%P^.K,X2/V2X7,!^+?!&':QZJW$WY3@2*#V,J(B<XU\$@9PP$"VTN=65M@)%]!
PM+F*:=/,,#@V@:, XU6?7O&PN_FKOU47%*3[@=*+]4@QJBR&'4%T-Q4\&BMJ4UE1
P'V*&27R*E\EX&FS0X8W.HT'43,$= OC$>YZ%:]9W'Z%\<-%_Q^(Z37@'(WOR'SAW
P?\]30&%FTN#FQE4Q?=02UQ[P1 Q,0A]Q.U03TD:^DH4AOQ"K=BS1$,G/#U1J=4^A
PQK*>'#02E\UZ%_#*/\K%XN\/VU,TOWIIYR7WMNGF!Y>,TP0.0JVEW(JE/H$2Q=JX
P[Z%@].#J$-R/97[20-[) !OK;#S$,QZ,G9-3V6X*Y3M9M]<GRDA%&-G>6\2K-# Y
PG:/VXK5'%M.=/Y:TZ 38*:A%D-U+("BFPKZ7EOK=>7JVBQ85ND#L^PX<ZPUSJ8-/
P^VTP-/$X*Z"38=0T>/52W70\BL\D1Q>O9' >6)I<!C7G:1:?S+%3O>:\^Z)Q'1K"
P<NKD6"&Y;4W[#^JM)KUTO:CQ#YW'JAU+95NRD:XYX8-K(X]3OZ5CF!IU]4&-6C2,
PQ<,RK6Z51-6P(.;S.MVT)G4=!1K ^W1?M!?*=O*G01!0[J+_)7HFA![R/Y65EA,8
PWA^.=-0G*ZLHMII__:08F#.Z#$[,)?#)HAT&@NB)>GYPD$ ZZ "<J3CTYKF*\FC;
P6HXEF1X*C6/3ZOO:Q8-$IUTY7JL@DWS'\&"/"]H6+0]?F3^'IQU ;%*5$* V;+AF
PD 57H'<9:"^X(7BKO7'5E0UV]D'QW?;MWYK;72*4WWUYHR53OIR/5@.&B9;4IKPA
P%BD)W_8-A="\Q7)ZLO3/^@IZI.'UE;==\$8?X?1W0UYV22VMBJLA,ULG=#P'[;\V
PU"*]I]32*<V5@/UHG^@NX8*24G#FML.:7"<65^L6!U\%C@6$SOYG+=/\TBVKQZP%
PC;%\S+S/KG^.Z\MS#!^BM]$2@L)35\54AE\^)B\9ZI?Q@13$"PG.^(7*#3$X>QJ;
PU1XN^\*+<BLY5>D'1)6'K7V6=U_"J5]_/LW6B(KS@A**VV@[N+F/TGD2A1#UI@!H
P4"T"K A--N!\=I(?8@F3XHN7I/BCERGMJAW!*?HE7_-47^V*1P:E#/_T3Q'(AY14
PYNG=>>1(&!0%_#8%9>#_J^[2.+);EL]8L&8E[UY(F7 @I/EQ\K*"_#X;:<H_/X<@
PH-_ZCYA].%)"0B]J7.?Z )B\!H=P[1Q<S:>_;&0\WV6S/NC0YS8M>R$X5*G@1K\<
P^EK6'LT2X:4R.\6])PUR]Q;_3^B$ZCUCVR1H^:@MPD!,<(*YZY'T@Y*62SBJVZJ-
PB_S'\5:=CO*!!<OR,2Q"7L4.#T#.,IIN0V28^^2:Y$GGY?L^(6[GK5ZU.\3M5K>1
PZ;J9[099\T;8.1D[^RO[M<?5(U.@!":?2-1Y";O(5(P*$5'&OD;1=CQB%-E@OZ,S
P#[]JYGF5<G>O5>ANSF/(4PVE+LKYU?9BQ2C"*J>F&$-FO5D3IPN=-!T&NI$$ZL\#
P;+18OA/ZCC);'/*\ !8'ZY#B_)V(:H"=+<>RWXSN\X3*S0X>+QVN'V]+&HU^>S'F
PJR'(/\Q7'HB'EUGMIA_2CW/:=<3Q8Q8&@=^3Q,33=,+?('MZ<5D+U\%?SD1+*=;_
PHGSCQJ'R+<&'\Z7RURSKB6^@/A<;3LD$RP&]'=0UT0VZP6^O]RGO5^PG33\D7XXA
PUFXA\6%M$2V@_=A7(,3X& $U:XN3(0I"%MUX3WLN3U:J[8Q=\'U. [RV(@0KGRDP
P69KW^< DH@_;# O<1Q:M1?@"J=*$UP8Z0)8#(P+GX%L-@7QU*+-.@3NEO4ZD7B\0
P!.7;QQ778-!-$@PYQWFK>:V812=N)Q''4V$+[/#*DY;P/()2>\K5I8RB)SX LKS'
P )H/>56]Z_?69XO#0!0[FHM+#*G\28:SG C3B7N6G<YTSX T^SJ2*(T("O3+X+.,
PD K&4$A:/Y\!ZFRYVWCHH2KU\53AVE 6@KBGW0X%:;3:+I]/3%N#IL#-G4Z*Q1F4
P1E=QN^M_KC'I__(,E!S?#YJ,0$?][0FX.%%5_.V',UYZY-]Q[B.1<QX6^?#E'OM 
P/!Y5V]01)S?0TJ>^+"2<U0<2GIO<X!\59:57:X6Z3HSC(Q9* +?T(IM?+DI:L7QN
P:ZQY![$*?KBJ>?!3SO+9)K]F"2)]$Z;=F:2- )PPHD& GHC-5J8(7A1".7''%_7I
PGUP5?D.C0E5&6>1A)_[)U),R 0&A3Q77;7A19N4#J009J29?+5?8W=O-(R_B*7G,
P*O_' 3D,B-=:0!,\<2>],YBN)@CKZ:@;!QIE"X4>]PBQ\73M&0R,1F8[<FT&-Y _
P;CY8E";;68M,B]U6 8OC9FLJ?+L2SSYEAT,8FP3G>PCA-[E9AJ5+T:\^(9UH<+VN
P+W!VB$#VG]<NRMN,]PZA3ZRW<CEJ1SX/"KS/[7T1=C3[7WFITAR^#[U2VW=(IU>O
PXZ8V"[+Y06=RU6Z%T0P:'&XWUQ46->.K"\4%\[=)5O#5?BIK G1+F=T8V).OPWYO
P@F+IX9RO5EQA89[']*?DT""4(%?Z60B/RQG4/1'>X;J.#X\1U9'!$]:7A=V-HV)^
P )7^G_!_8'%NYAD#A.4(&L2#_[S['FBG$/6^^X3'R)3!LO^B%K8EUT5=@9WO!U9-
P-0&(PSH9P<Z4X%*J;/OK4Z7%ZZ-+^B (7!V 'KMFV)*R !>>B3^E?NE<4>>:N+(8
PDZ%QLAF\6NEB75'X]419F)C)QUH%PZ_A-VJL28X6RF:$ZV,J/O043>*]_V: K?J3
PK8\M&YY&?#.#^^HG!A'8J]2I]'V:O19#N+;S/QCM[U]A@^+"]$K(D$9+]Y;]+A6<
P6^NLR0CDTO:+VH\P(<="V\#6XZ4\)-DOJ9[K^O8IAJIT2<EM,6R21%$(&'HVO[D!
P6%5@\"]&6V;^/Z/@8?N&?I")^%MW("8X"0"/XB0?XG5!&:'Q(&,R;)HOF;!2833R
PN'8CC%P7E0$W9%H<!4$]M_-K](BQ5RLKKHWR)U-EUZZ]&M5H=;WSCDI03Y>/R<M'
P"2"[,<DP8CDXZMU-9XLTI'*N$9,I<U&(8NGSM(N/N& _55#[)85>ZGP4;[Q>5*W;
P<>-"/.EW+(G!ZKRX<%ZBD@I(I?3(XV2'[>[VV 5Q"Q(%F?38%ZGS50D#")AN:<,(
P<>Q*$X^"8LN#&M(9%:",L8B&MCZRIN!4 ^!-D:#07DX=%R'O(EI-I7GTJ>>8G<CP
P6>AYYLTT.:@AG)^:!?X:=G5N_9E7S<35(K[,;ELPF'6'2*T6UP92NDGYRL=MG9-L
PC>7SR9*7@>3( ?#H?FZ+"F"QQ="_S5&Q0@QCIW@XK*>= @!XQ,9_UXY3?WO;0E(I
PG=3J0IT^/KNE9@Z4[50^1=9GD!HQ-GS*1-3^*:](XZ$ZH""_A?<_S[X/H6*<_JYQ
PMX8>>D=G-,G%# L 8B5*#I>5'+2;])O.4]XNW&L88)NQY%1^21\:SDXBDKZ.H<"O
PPF6QSR^F^3 B_AI?[&:Q<&W8MJ,09E&G:"B=A%;!5Q?/4=8JX,F-S90.J#PY]@3F
P1]H[3UQ='R=9&)F:,2HSX] B_X\,%411/OF?_;P#R,LDU=*CC"!45T; G9:_'NJ?
P)?(+ND63)N[C-)R]%/I7)6M^#0+62-.AG?D>X<W@I9 5AI-;+:0;*PO#_(>*>%UY
PE<C_,X^YKO:6T]HN&(CI&!1%O@(H?MAS?'N[*6.PO?I5$:%:;U%\IH4\NQ1\R^X%
PGLT5;=S_ ,I4=.&F267AB!G/$S.FHYAK;)12[J?BZA<V*W=&C!:$;O7D5@#D/'_7
PF@Z&0IX[INIYCGNO;J1;6,ET*Z >M_KI[+#18&;)\F"2W1/$N]?5GVB46Q3IJ?MX
PH$L]07"G90281>1TOI$4K"I<=Z7'33MG.0BIQ;B!Z=9Y&':<-_\"<ST&-#L\4.(H
PD!6 R(E<S@'@27"AJ&D3JVHCJ?E>"4GO\K>%NY%&39(VC7C(+:**/(<$,PSL\(P*
PH,AB)B[%!VLRFEDF7S.=2;:^,NA(@LUP+M";P;D2UZA]@.5#T&'*XJQMQ;;2'ET3
PI:P\S2HTN0*2QPH&V\_T-.K5]2A<V4G?55/@0CY&@?Z+;U$\?G\>PSE_*G#Z1X7 
PH>18MT3R"C(_[02S;%VU+#.Y!CK2$AT1_$!$-W\/852TY#\YR=%"![5 PTCX=&:>
P/.0FRY> S=VI2X:,.!B25D&4<O\'^S'I[B%82W#KL#J<3M0$YL5ETHV H=5N^CN:
P=;,@ICW"2B!YW.#$V_C]A[_MXA1V Z+E#Z*, O+/0S"!&)29I>^UWK,+^.[@4"%Q
PWFL=3S;DJG%KO",DU26Q0A<I5W?QQ?R;+=FU\6!](E5:^CJXA9I(@ ';08N[)3F;
PC*/QN)M(Z :SKVL1_ ]S 5W^EOG:T2&5S@U/M]+))"XJOH@(XO_'LZ$9P[VBRQS*
P9@R-U#7S^)"J]5*(&SU!,TJ*:LL_AK5CL4H/!YGR/]DKOG)!X[^'N,Q4&DZG,W@:
PXV3L@025A\@'01+F1J6H/F-I^=3>9E^<8Z<(_:%?JU8HX -O!C8(4*#"-[/?PR2>
P*H:MTMJ<F+(V$]D?M#@Z(&5T%;"[-#::F,Z,D2LUQ-!>F!H$R\%ARH,,+@ ;JJJ+
P$(+N5;))Q%W5EM=CPHX +?:?PP1O:&11>"#GX3_?RK99-?3W$GS613.R1.0EB\WU
P3R=!TM2=HCLSN=4[&&5?_=B-2!',LA;>0J.0MD+\ A6?TY)683*Q<>3>/F6[RRZZ
P8J4;0$8-]7"_6AC^JEX\HQ9CSY\K]H,H(*&!6^]LHZHE)03+^ER%K=8#@989C)F%
PE#1/HJA.&P ??-F:;"XF\T-3W*?KCQ;G^%<Q\PX.F1-2=[)(;D,6R"MV1#0C$$[[
P3FR2PZ8-2"W[M3'!;TV94,H,7\C6</%8/P4_-NLSO_8@@*;3!20T1\!$RF&E<;XQ
P%5&M:ILK=KVI6NBMNS;T;02RD "1[YC.A0@+B2MNH(!KXCDPN^4>B0>J2K;*7?6F
P).#S)YGFGQ0&UH=,3LVH5AC[D05!EU%Z6*OZ!Y9X,?QN&X ITKIR\;&XEG)&?.)&
PW7NF YP4[]/VG94(4-VB< C"L'.F)P$K::JRT;A6H 0.X:Y_$MC>?5T$&E:^5%@0
PI5+1-*.7"<%N=2K^FE^%33)JD&/R=U@VYHN/!YTAIMZM[(G0\W,*/9;[G'D1#;3O
P0)0?G-\J$.T\_.:]:Z#"RBB3BNU<?Y,*4@@_Z>'F,:^>/_I8":#%.-_X9#X3=[A/
P&S<P7-BALG(6Y24%UM%PG>M/SOY3Z:0C;1A9)L6]O\EA%=[^E/N&T^Y.JYK>N602
PE)<P8"R8\H3@W)UV(%'#4&%@T>=<3=4C$_=E26TW< Y*__+*2#U"D1?$^+43:LT@
PRNJ*_GT,5A4;O3PL;%%GA/ILC6I*=[M9RR>O!&8PD7GAW)"PB<4+L:A:UE Q ]$L
P_O";#F)4M.72=R(@#X+P2"F-L'>K94A2;D9O79^/\2UT6R[Q;?W^$XL&L.<)*<L>
P;+C($6'5-H)3-E/F<%&EW6#I1Q60)=V?>435 RDQ[(*Q#=._YMGN6AK5:%@^--LX
PUP?)3V&B*$K:XYU^[UV:EG][J)-9J@(M6>*W'U6A4T4SB!8;%W*WGQ2>]LX(","F
PKTY0.@P@!07%#9*'S[,30%(8";M)R=?-ORN3<[VBB Q5/[90F])NBLZ0EU/R']DV
P; PJ52MBT-W$NQC&-D1<D_;QZ;=Q!V_',&XV)#53.68L,)1\ZK9FD?!*60F?YO02
PZX8X-%W]IQD8'-N2<^,,0=&[YK=.HM/E_Y6/;][U5\9#W%]:9_O+>/[$J!)^W16)
P6H^5_B]L3UZ/;NM:;%1F&_-X/ZY_C8<"%$^Z0:.7G'_%,WW7'&_P%1"R>JI5]Y8K
P;3_O'()GD3.<DH;O\?>EO3.[9_5>[?"UCT;CU#+-Q@S,!%F/QJ1D395LL_48BS);
PQAPZK_K+#WSH/NIJFTY\,5-KC'4'TC&EK/O'I>XWU61LWI]^\VN/R^+ 9H.,-Q3.
PRN<\12?RM ;+"'KJ,=8#OV]"_ 5_F]SGU_SNGX@33YH=EFC;[T\4QQW$HH4YC^_B
P6^E1/[$ 7$9-6E(!XD"3DE[T)"%K6.0ZKBO1[15G_V ?6;_R9OE\T#6X6X>B-/D1
P@-RE.[=;^GD_' 0DP1PA(B/D4E!J@0G7DV.;8 CA5V99N?K<5@D&>H1*3:H)XEC&
P0Y^_C=7F19 R@7,A2F'G#!^#;OHC1% 0<SG%@Z3F@I2,='HM9U3^'YWQR_V6C(X5
P@M&;OY%=Q24\%8_-<W7+74P:@LON1-_ICB//N$GY*0H&?)9,\8@^\-^<+=R((SFF
PM19RL1>AF88@L$))&VG&A7W Q<*8&'X<*J3A@-Y\%U=Y*F%\87W)]8#YE.[7R<6/
P!V1W":QLBH5@ZK.NBIOC<83?5PM,+0VE9;:^=P( $,1<4Y=.:^S[R/MP_!*>.4;O
PYAGV#$HK+-TK G3MZE2Q %'0:8L1V-0[]TQ#K4))9D>"X\!AVC^K[\'E>>, HE)'
P>-.JI[@N!R5,6UBL*_ 5C_R7/=EMM'R.? :0UGC/UQ1OR#E*V#*XW=,V4'&Y]%[V
P,T<@GI]'[9!#MT6%DP%HNT1;_HJR>6UF(,G?1%ST&Y&:GUN_,:*(5/ZN7N_?X)(K
PY.'&I'ZE!A@P]\/@*MV.+J)3\C5*<4RR]1S8%9GZ8"1M\>/%#<FYA8C)JE'VY1YN
PA@'RFU<5D427B@0$K47 ^F+,TR1Z!*PQ&SO>SAH)0TM;,+#JE 9(@Z6ABBYN>7^:
PH2U?9G'L04A1:2@[THEZ)MN[.N ;PSSOX!"Z)?$T][=JTAU]UXM#, ;W[HZ8?C?6
P2>:NWL<7+4IIUYTS\,[""=!%_A+/L\+*3;N7S<=P")F!S9O!N?Q/>-%D6F'W)33/
P  -I!\.+PG!:C1=*T38A:X)@,40JG.W;RU\ S4V3UQ-!&HU^G<+MGQ#YD[9]WU#U
P2'P>3\7U=]W&RDU7K)=[2<V%9F?"?J1 UY*9O^(Q=#_TV&,&+2:\D<J,^%0-@&Y"
P#HOP ,T>FI/;0NX50>BTB>:9<IW<8()_P.;"_;9^E&6HE0HAQ4ECT&9SM(0T]%3T
PCH[1".ZHA6(5,C,O5M6\T$<EQF0LBU_VO,Q]%V-C-'&VY@IDI#E)G$G'GBP5C2!^
PUW:Z2TLE]D] P@O7R<71T1Z<@N0HT9W\!)\^Q(9AK8#I^'>N+& )A8C:EU?7K8 >
P8_L*U3(MV.*1XG22!![EXJ&Y;I6,W"5T: O]@M E^\;>F3'%RMY!Y3)EAF.]O]!B
P^_8GX6 7V%CS9*<#%.;]O$=]@-8%E1Z;D3*(>MF,DKNT8&J[@$G7UV>?H7L/UNN;
PQ>O16MEMA:(Z?@<?E^>,EULC\: _GLZM\%ITM:S@\C>5XC500,LY>;BZ@0W"W_U$
P:4)W1"1&.)M2BV>(D8-!K1^/"R+895LR&.B4QD[A7LA-*"M8GK?&@YL L,E/_/ZX
PQZWLR%*[]HGBZ"JJ,?]KMKF%%;W!@"S<WG6DNL.GD*D+9">M+5\47X6M:Q]C.?&:
P+"FAZ5@6K\&28.&^/,9T2)#5X1=C_Q\#ULIJ?G+686BJ$!OUZZHS6';T?=%#1C+!
PG=!BU-(YX==S^L7Q\[P[C<'YD7-I8N_9R:E=2F>"=+I#DVW0@.:#0OZO4:7)]]O6
P.L^1X3^]@###^@TYKCD"@2]M3JB2JR;)LVF85W<-GPP67J*7K)5N6FY$VS*UC?)"
PPT<RRQY[I7TSNHFV@_[-:%JT"%I?A:X,'!DF6M["U*_%7!"S.Z$?9");[@ACJ7U2
PA?L(C38 %6<:&X#]$LBB91GN SW]$OTD&;4^WR,CC=NA!AT"W8SJ./3Q\UWE;OER
PW@TY3*^7=4EJH!5_8GW)5JKMB\^P:I I![+W!<F4$5*S;.L3,0Q^0QU(D0LE:#7M
PP8$"',*+T"O<&SA,?K0B=>L%D>NJM3?%!@2^93#+QX;\(?I&QWN*R(#IY-Q51C0P
PRH3E_SQ;9AG/S1CQ&BJC*_E<''0[^D(2MAU!9G0._W*N5%!)J<Z&F8$VZ;^$OHM,
P(-:P<3S'5L=FQB[Z#;A>+KD/)1 $*2]\;1[I5SAND"DQ.)]I'$3Z/, &&V$+BKRD
PU2IE\T3:SX$(>TK4HFRH:F%)\[:-[@MJ!I!X1#C$)?+=Y5;RW,]V!(QE-_%#H18I
PB2'M?RP-_PC<SX42XT GW!X?MQ?)IG/S_YV:LH+YM;_B++>;6\Y[9^_(PIF8XAON
P =4K37%.FC^4;M.FT@Z/[1D3[9SOSMP;;5X;7*(5%P;1AM":;7)'+9Q^\)S[Z"I;
PL@Y5<\=:2*=)^I:6C7^+Q.E!6?BD>\7I2"!+RDQOKE"U?%>XSI[_EU@C3 %?CT:3
P,S?.<;JIK[U,;!%,\'H\<L0&?L?#V1^-*#[ &8VRJB0MI'E,TK&^5IUS&SZ^G6$K
P]WAOFBWLJ<P*#]T?[%4AQK48*"@75@)P1YNP*#<,S6P'PX[3G=( 7V8<']6?9]"P
PZUT?KS $VJ'2IGH@;L+](L1ZV<Z.>P&\7("\3ECP?F<BW5G-P#&8ZH^92R(8T1.H
P*"YU1H02OQ[^Q-F,<FKE.%EE>XHY.*FN,XD=,G.83<E!HD_K\,#CM'8Q373HI1,M
P5[H",*&W0]DXO>C]1PI'R8KPP131:="8$?+!P[EZ+$;+)]YN4<?I>G::M7"42X1)
P(_4SBG>1"U K*+]S]U$M<K6COUGDK11OOFAW(B35@=_*"PAF6U>+U6ZV"O8VLW^O
PE,GE=VVXV;(@WVY7MK"@A20/:CGXA4\LVCTE?8NXV3&"O827*][S=E*PGJH/L,&O
PSRVCI;7+$H(K#\[VZ1W"=0;^%,0SP =A8I-[4-\2J[59,<%42SB<3MM1 ?LM;A#Y
P5QXK+'!(\D_VR"#(_E0"FW=R%HZ#W]?Q%WNIF[#D)A,?=,\D]#3[99)C#3#)VIYU
P"S2OSN:_#5\GJW#]GW:-PI^^OE.R=XX#<O%U$VVH,.+5Z; D?56?JGF&3P0#K*36
P'*]+A,T?^_*C1Z8BF_K&>2!5!'OU(:--> %TNBQ>?>0 4@/GG#/5E4TU0SDK:L*%
PH87SWB U>B7SG;.+\V(:_HVI\8X!_%(KQE,U]]G4SS)[>:1,Y-W6+Q P0$#ZLJ#D
PFLH?A8P5'2N:0C"9TFN@'ZTYJ" D>O8YS>[F15R]JI(ECI7"E*=]C&  JI!F@9.+
POW(^;GJ2^O>M4/K K*A4<27Z#,.'@XJZ+1LG?3[9R_NA^!\Y0[S;U<H]Q<L,ORKR
P4(=;OYD8+#0PKPZ%!WJHUL]Z/DME0J810J?B9%_TA/HM!9&W+D+.I?PAA6<''V,<
P@MF%)99.\<U[NJ]&T)2A0&J%S9UBCOQ:!LW[-M4B?%B9F8OH1TL7ZR(X1"A=3?=K
P:-<#/5-C\H[;2L:HX3)$.*'F -R$F:#,\E6&>2!DKJBNI$M%V-*91'XQPH]CF%LU
PCF=C7C]4^?6#6Q\#6-_*'Y,S@\_\J+VH7XR8MD*N"I\=1T< YA)(0MTAT/8<FM@B
PE[QW 6[%7PC.Q%\(2+*N]I52IF&(J57TV*H70.L[;W]5!5$7IETAY\B.R0%MS'EO
P/7'>+PL(.HQ?P,6)@7'(<>;!\GW=^;3OC'5IUE)T.5B%6L&BIQ1K&9T/ 2C]89=)
P#)M;Y[O'<H)%OJZ6;(@!V$C,DW"?P8-7-B[Q#WFO,>0KU&,$3P,O4$=M?%QP6:7T
P'V263,@66'\LF2U@4LYZ417;I@SXW*<2R.OQA6[#LW@$J*RB<VFJ&=840X?WX@>>
P>-;2>![H:E32C%/Q57SB_%7X7WU&W,;Y,EG8N67RS]R][VU\+9QT"F]CUCUND>9U
PW:\EU=LC2;?</GP@+B!&OR2*O5Z2,+"\C!W@=O'R;T,,' ZD-J-\"4A#!%T'?:Y\
P38Q!@*XX%B^8?(15$9BUTXWYJ0T)>V5,15N1&!U$^0VAYN)R^9R?LAP(QXTRD^*T
P;@>53JZKFCG()8PG( K>XKP#RU?+$>1\BUP-KFWB6G"2/=*PYWT[D&0_4D@C,,22
P_>!0&_L%TW$^FP/T*=_*VEQ)7!YX1M#M2B[8EANS$(/"BQRQ-%0#FIAB!MF\P&76
P1R9+]Q;/(BV<._A,_2IL4NQ$0.&%.(Y.!WB2=^>_>7W_84AU?Z[;=KP2F FO/_H5
PBP^R_18BP0<#)9X)$]N)2Z')9MZZ0]?@TY[-O=QY8)F<"832DEZ6IMK!<ML &UJC
PW[^BTGRAKPNVQ@/VDY2LGW*AN.":@90Q"97)]D$M.J0JCAKF,-?!(U2*<)#=<SU>
P1[1KS496'PF_"-N@=_C0KR ,<3+L-2'^VFWEEW)+"\HF>\%>FBU8"BLH \MDH*Y=
PB:G6 ]WMUV]2!-'[UNG-.5/\)N<V1V;C'WN8/]U*$K7]TTZYW8/A!_SYK*:DM%FS
P&O]'DOSIJ-T-2?S&$O<2/3DG'9OP%.6I)N\L8";](84N3]0YO5O_1R!H&.&_/ 'Z
P_-#(LL[$U]<U26@_P6 2(BH]V'>?**/;F 7<W_6Z!<5S ,GA'N^&Q:@4(Z8-$:ZT
P<3<?W)3JP6R/--74-^&;PH>Q\5!.M?N>%NE"*-S1L*>:81(9K@U,!SBGW1FGK(G<
P:+8DX'>>SIS18G$.%<@5:9"-PX!?NHM0#O4XNV0N(]E PJQG4/QF!]F+,^W576!O
PZATAGB9J,JNXXG"_SJ,33?^U'F$,4^QL9CK:&[O%F^ T6"0K)!44;TD]':'6ZB03
PSCBPL^GI!GW23_1,\ZS #7$+V.&&NI)BH9G$W$00(6AO&&A=^43 7(5(YFXDT0PA
PY2DQ_Y$[GY>%^ZNMH$\> /X+!;[%0]I%GBK#CR-QW\H&M3[0-#.%AFD^0W5Z_Q K
PC+Z#R9$[S::9D3,<^KA[*G;/QMN]"/A'&-MYKQ;5QQ@/T!Q*#(0X/YOC>$*M:&=^
P13K4<'QA(DPP??A6RM6\A$4C.DY._0G2(N&VGY_0(ULG0!S+BQUAQCR*6^.6NG, 
P0(Q9VH(+/%#6BSD 6MY6,0;,3(2/T:S2T1O-2NA( -JDW0&$/=C)61+X G0-G/)R
P7A[]/YT,A'#ZE7%X:I73DJ:'C>J_GU$=*>:4N@ZD!;&:G(/U"<C'<WL<4-95K-NK
PA[9-A_H*))Y'5!:IJ#2)Z886*,,ZL<=I#=0P=-,(8>\[)M&.L>1@.*[9S-D6#(&3
P@JW=&69V7T_%Z@$M>6<PD*KGH/'LG&3GRY7_[^9KK^Q2V)=1 Q4D70 8$SMKG<GS
PJQ]JX2)N#C'Y,"34HW!^>D/U;OT<?-O-8M$;)'KRB=*!/\@"^:K6_Y!8.CN.6W<G
P'(L!1;?<*>+*QW&.0.6(-L S65>C92SU"!\2,;ET:"?X.=X\!D!H\8V8-$EJ#I[E
PLRAC;ARDO*P(7ZZGX!#92:HJ)*N*Y!C,N.G">=OMK"+ 06UVF6YAKP6BL20OL@Z-
P=]I^^Y4HM\Z6=)1^T#:%C@:'GA1X6*FQ[CY+L*Y!*'JI5]]\=Q=<NIKEGR66(?GU
P6D]QU)EI668H8;U,/N)&\OO?%%Z4GKWC49E%\?2K/D:?@ A\;O5EA=Y2CG95*M!C
PR,S([OF 3G2>>SCI<8C"W-O6;N?KDKLT1]\6J28? APU+$:AX6B-A<*^I8?(")>-
P!=+ICOWH+? ][QGM;6ROOOB0]P"PU,OJRE/)^,W$K.^0G34"ZU:PC@D31$3'Y][H
PNK4(HA/KHL$!5!*-N#J_%WKM6%F5'(B' @"'*B^_$$VV397^RW167G42_.L"9:LJ
P<71L=6L6E8Q1B4'4>>?)_LP5T 4R&N\8(T48YD[@7!%P37QH'TWRC4/0_U PZ*%L
P!;W:56WUO-)F2+A U"PA&*<>#%O<SPW'5@KF@=1YNB JQ,G?)YQ71 DN-,VAR'#<
PD/S':'/\X1ASI2W(\C2%[S'(6]?GBJ[[:$8+3#*0: ,_."!B>0CHX/%NCCXZ_%L\
P\?JDE6*.I V.L U"B%U&3FP,+.0N^L$N.!SOD,+^VU'Y?L]0%QDJ!%;?4,@F7#+)
P%Q<&2/5]7^EH:/-.$N,.2X<\&ZB)3^[+IE  -(@?'[HQ ZJ>8?+6)'\KR&+;YN(]
PN+J-BE+LN&G%H+H)#XG!C"'>M\T]"FP7EPPN[X5"PX"PM)KA;:?EJ)B#GF]W*8C?
P]M$8-6)PBV5>Q>43-DDI$^,?+GAE;-&V<W@W(_1)&!.T5L.2T'FTZ[GWMEHN]G;R
P]1K:_ [1_#4@T\A6RR3*FB7 4K?6)F867Q&I HLB+.5LZH)B 8%P6-"&?KZJ]NT7
PN."B/75!&DYJ1,@V@R 9%TCW2/5<6Z5$V0LC]Q1A5F_KL+S&G2@$<DC=K?,*S:4^
P(8GZ<4=S[$-6!F$$#SR((43 3:5(_%$HX1D?^#MQ\QX)9#LV.-'9JTQ;MA2_W"&!
P#(@-^3(F]E6@;SU'Y7TOGBOD GC80F[$2/W.KV^OIX-^#ZX\4F5AP>U-[?QK:>0X
P"_TDQ;/TJ7$#)+=G.<&QUTYS#!2Y9;I0()P$'&>,=V0_^74V6FC^K!9;#_WH+'( 
P*'RJ(5ES(2N?;TC] _S&A-[)EU^=6X%"CDANL*Z!#E*H F'S<BMRH1]OEYQ1#)E,
PD%&H0H3W_M4AP+4!<)!)F&? !DJKW6F^2>__B2+6V_%#4S%T(H$IAG8<!186X71Y
P3ETI:]EH>%+M;GN>^OJL1F\KR5W<S'>G9"&2LD&<Q"<7BXD(*>Y\1@OKUOTXB.G#
PF@_&M'^8E._1.^<XK_,*^DG+,6)I:8"*?X9C?6?- XS'I&\38J!F7+BH8EN7N1Y'
P&M94%\.EQ3,V<U&837J^=6$9Y/U!-\JCYRY9=$%JZE[MP4[A.XO8K!5/H?/3&]9\
PR;^%X/7[#I%U)P^E@QQH%C<K%9@T;F7V*S-$%5_[8$J7.@PM[QAG0S)G-@AE$;%6
P*1Z^]G"C!-W<TAQC8SP4$>$,Y0VP:%B]1'],TN3S%ZBO -'A%,5RADLVWH5E"/ET
P;1D(-TETK%P/U\^FZP.M>'%BTV]%::#D2N:NR.2;"I/RW%.G=0.&.[4D!M>P3!9S
P'WUPL\\\%NI/*AJDDISM&S!FV_H2L)-*=B2=;(9J<HSS"#$2GVTH(8JA3'(ERTIH
P2\6Q$)D/Q47,M='TKU+(L8I.,.:$%6'<H.^3<Y#,F@(U4!];D6AH\/5@;99&^^)#
P+UR>=2:J+1N>%.O+%X0F)\0AX'UOA<!"?*WQ]W<R6YY9.JW] !#1#"<P#JOR&>Z-
P9 [(,)U9PBACDT9=T__*N.#C>4.=.L-E3."8=DD' F*+1VM-M'!A)G/*@4M&UDXZ
PKC2[BM-9K=2-0=2/OWQ71.U1_^=Z]/P8X^Y]Q.Z"*G.7/'S/==>X,R2Q,6,GIQ!9
P1G0N\"'Z6/;L\$8?3Q6P1;C"FMG^3[F!]+ZU4BY8>6_+Z^@(?N+LWLUI3=(S!F=%
P  [7.N6Q2D99^^2#Q[%.G*CSD^KMY+7X K0*-87B?SV+9]J,@VQ[8[FA8ZZJF]E0
PE/YJCU\OT,/;Y'R4<C"UL.X\K!1_P)?\U07(W":SP%'L;O)74S%:,*T+$<2(,&"&
PB-,%F"3*,V2FE&F,WWUFCI_80]/6T!2D$;6?83SU?1'^EP+99*'Z9<BC;G4^2S2\
P:9B9GHV0IIEXT6R#TRN\#O0/ZO49+2$^?N87JRS6K9"RNM5\5856Y^F=@T@AIMMM
P+P=7AKLT6(JT<>A:)CM\L6;D:[)V:EEK9JL[O3;T,&20$^P>4;=N>,JV8[%]/JDV
P1P-/B"8+"992(\_<ON1X;Y-)GS&),>@R:OP2O&Q+3O4\N-[=>6.%AR!&#/*T-CKB
P)U?TK J_@ZNX)T-4"?[[ W' SIA_6M#6ED819F#&)=F!C]=],397%#/>^U%E4;["
P+A9 '"H.DXM\(!5U^\O:6U("[<LH7T"8//1\:3*C_J(NE,I.3%2#!KOW)9:2QK;Q
P&LLP_D1 C^P=^P28 \Z!"@9!:)PB:@HE>(JVM185$#D*[/X0^4T<EXZQO=0IT\G/
P5]!ND N6E:N3B;\-2&L&E <>N2S/W.7ZX9?*N*L,]KP8*/^]J91^DI,56?O^[[5)
P,74$E5N(IV62"JO6C3!,@NE80](H$O4C?1U/+AB5R!.[PQ=FG'NT7FW2+TQJ'0MT
PPE7H"+:6+15D').<:2<F1Q")= -[JIG$KJ$ZT>XMS=#"7+B4;F,4%5+$Q/_5>U5D
P$Z)ZD+61F'!YO'Y(#Y.2$IAZI/2@/O&4_R*5-\(9ZX,:UR[FCT_,=O>&2//A?W/V
P4LMT@9<O>12NDP%61#P(:7%!>^56@W/#%1=9I893Q9]38PT$A-FH)DU+8AW6><IT
P<Y &J[@VN%L8T63OZ\08%F/ 2UF1N0-3M+='C2E5. /F1SVY;D=M)<J !PDJ&.I1
P-QP#7)%8'M!;\\AE%;R\!6T6''J_3M'E[@LGX(GBW+]4S0F8.,BC34P=?=_GN7(R
P["C;KZ.\N,"3/NSGJO6%J!5#_UTU5&) :WM,J 3XPBR+&O4M"T4@6*_-!<P,=%K'
PQKM76Z+6AFL/P&MJ]GL("*FO$ L7N\,(!'H9:NT&?A84BNMOH0+/UL;-D=>;'A:F
P2D;6\BG<(RV.E^BV3J:K'_ $"@NM;UF#BAW(D"\*VE^GT=-"H)CI ->#WI]/P(Z#
P@52A'  V"1AB'N[Y0D.B&S%7H7L'L'"/C/67HB;R,CQ)\N]$*[:)ZL//E"/OJL$0
PJZ3^@'!ZYI/4@!'1*9\"2NT*A-6OVVXY%!U;7?R&@=:9(C3!VFM85?H=N;;*3;1#
PA=K0BFH2L\WBA9K=T\?=_ :SZH6RY:;@%&S0S'7%E<S<F+B.Y(DZ(R)6.?24\J?6
P"L=L?F4;BGH><RG #DO7PMF_5:V:!"+AB-\!R)8OG.Q9JW%%\H-V?=JT&>H3DA3Y
PW&(]?HV3<M@P=P4&,1Z""EIF.(. G3:6HX\)8]#*G 3XW3-[M2&8?A+LY>A);)'Y
P8#Y\>!+"U@E[N!]=U0L!>JN2;-)SSF$?1!"+LSSA*F7\E3:383!K>P; I+&RAXMB
PCLW,.$^153$%[#=N(]/9KIS3R_EX"HH"]Z1#63HJ/T1LJ1NFE-?7UCPIPA7P]3V1
PT6G:&5HWT3.PNK7F9H?NLAP@'OA1C,K5SL[V9"#7W"\#5\&W\F0P!D/KN<MCX11(
P6?5L>GJ/5N^8+/OU+\PCC(9\9PJI3!.^$&<\C3[E@B0<R0@Z;!+?6^R*#$Q7@3H(
P<K/L),*F&2JO>!%NV*,CHBM_IL;]-1A;0+I93"Z-@<C]TTCU.<T8&?J0 ,QQ5U4X
PO%EF8/S!L5W8S75_"Z[IX$Q!?0H$SWM>.+'95M)RZ1/H^T-3T3(:TZ&LWT,4[6E0
PTKX(J13H/JGJ9IP^^K,6K4]N$E[?]\6$ :$F3^([.<< BF[YE_2:A%KX3ZSE:X@8
P0.W_ EFCYHR%ZGU7!(U\M05.QR]G\*$T;8]:0-_8Z&.]=N#EUU  )W&N3JHR;?U-
P9OL"IV@<T#?RV@THYMGL"^#+KH.N]2NZR1J+L@XJ-?WQ+:]EL _\7.CEL-7_1>^W
PR 5'T'2--(#.Q%"C$.P6:PU"B54&3NV)%705JT43^2@+0CL611I@B]M@F&4OOOE,
P7Y1K\P3[.?=YE@5+""([8VQ)_0**3R@;D2=]$@YY%R_G+)5Z7Z*$%_D(N74E' %D
P%2Z5 HKW $'G[5#U0(HLG^,V3ERDH.F")&/+(+*)[RJ@Z01.*CCKP?/^$+)WR%] 
P=,V\2U2(73KIQ^N1<LQ<L+%[VCP3GF\0!Y/9U@91H35/WO=7K=Z@[S+<^ JYGRAY
P9<\R.KNS'%ZIX=@(Y9W;/U\>0&\73&%!T-%W2@O^;>(S3^G80I5[<*?$<Q'1Z<*&
P80#'$5*I[JA;7(#!]S9/.4%%.M+>'['#SR4,S$.1;_%X'7U")&[/M!(GF7EZ)[9$
P64!M,IPW^F;S>=%JKRJG7%Y"S3LA9D+!SSQ;_7DMC*U9?>MIN_M<1^;5%=0SJ1Q^
PD&4#[7ZK,-+LV#VJ-21S9L+5NE%HOS#$R6=S<;SD89-O5ZJ4,/D:K=T@$E.6L$*H
P@7KU [,!/]!)E7U\?[KRWY>>IG"Z0%2FXV'V"NY<:5Q*6)YV]R&AUG0G<?Q?]3;A
P- IO=M^N<%*M)PP=HH,N8/K8@BE7W)[SX(*\/?3*KD!3$_;PGJ62%FF[]KNYN@&+
P]_CR>:BJ2^P!<Q%DT Z>%S6IY5AFMI<1E64@WFE6RA*O8K<3TGI8Z$H-2S/OQE^)
P]78JM2>GMJ]4PBNEEL("C"XBVP7P$#EG_[L[$0N6C^C"+@4!;.=[8.J^''D8N'8E
PG)B6 GU9/] BEFWG:3Y4;U:"4&EJ ]+AG[=5!=B'$^E:IFWR?Y8=O8! 4KL$%JO(
P1(!1J:EQ]3A[U(4I4#0DUQ@Q# W.*6\V<EX+FZ:MY#PXW+9%$7X&:-I.[30R'[D3
P;(8J^1;5[:)_$PG:H. M6[)NRO&-4F?+FEU@MY/-*%8'ODE]+@")R#.H"#G:BD66
P'<!<A2]MYU 'V0)(ISIEVKMY8(]=T\#]W@V4W(\_BA@?<4@*@19NSG8!4VI<?&$<
P[<O-MF)@SW> (E"&YT;-5DE)>-=][RKX]XRQ\>X49P-4Y#.Q&AH1F"T(V)8961U<
PY)E;BRV$8(V=21CKZ=@JD?$GT?(!L8@Z"$^3,WQ0IL_0*= *#EEQRD4^/&CE<@X\
PV'_C[6VG\K*;936%R0!PK_\_0"Z9^\2$XFTMPH&&E,XO)9 WIKLPPVT.1Q)\)W*'
PI\\M7$ [/3"522NJN.HL+:PDP@GRLX^BRQ7:G,\1(>KP9YT7G>])^*@+EP[I75!@
PO?-%M^=\B_L,899IQG#*HL=A;*F20]18U^:2 _5C/EE1?%P 54CUF6D@SI](NG#A
PJWS0U(C.WHXD4 -5XADTS![>M3R<5WD,6*\-?);=D#*X^U1BH?@;JC J$56OA_C6
P]DCKT9!5CN1:'O]'1#^(.]V[TT":AFI]63&&?@H\ /J6+X#^7W-%#KWB8860/(N;
P8,7=4M5NWZ3V)\M">7A,Q:DI D_A0%;'RU>PBYX.8)IZD\HDW:=B+TXP6KTS%L.T
PG'X@!U_9@^MC4-WI6$[4&B04'9WN4.PMO[Y!>H(BSH:E3J:_00P5["M!Q(&J?I+-
PB,O4UW>I)*O+A-&0>2JU='W>['YAAF#09?^*.;^>#D\.<$K!%D?A8.7T2GP<91M,
P^>QF_T+,O0/3 \&*I9=U]T.W6>@T+J/8% -W1'9ERPT@=:K3A^0J1T#Z'Q9\ZPBL
PM5'W$@](UX5W L07N2U@5[NO9I*Q.-29!$;CX]JWCB1".F.*=-5,/JL+2=")#I3!
P]]@G4;Y(JG3?(A+T*I( # ]AY20F_YI]L<LX8T0Y*IZ47E\[W89#^92A^M(> "/0
P>(74@IR<:\?Y!GVPK@($ JR$$_(B=3$O0U^+2WQOMFQRW7=-0:>>\G1R_ZW;M6%C
P9KTA"L'R*>E0?!B;@<%U.!\TN:*^A#[/<96?"LL'>[Y0WJ"-"57\TJ,G+HP**:5H
P/!#JNX-85)&OC4D;Y>2'Y:]9?1-GEI?\)RIA[-9>YS(#TS6?EN<^=+RPMNS<&Y >
PR!1 Z1R_QKD-'^;^X]-12*L56P:!?5Q(Z2MK6_KVGZ9GKJS8"7$R?QF0WJKVS3)L
P8#9P(&E# S7* 6M[C[S HU_L,Q(A+=<V180 V7T3Q )/&<QB7%<&[RT;*VC%V]]9
P;,;Z;TA*82_W^"!A*LH;Q"N$ 85!.1"^O(5>0Q=[_5SJZP<#-NCC3_^K:I<30@A=
P*K8SX#)IS((K?=22<VWU^@7%-1,7Y$G!ZT<FHG0J(9QYF1D55::/;+O1E=<?MK(.
P(PQKLM'TH(C<P,*8%1( -9 *S7;R5B^!9&ZU$N]M@?V0UQ/@#Q&EOOJ>2H7Z1@-M
PE^;X>90;CKBUE/<3*(!F"$U9&<NQOS:_M%;>C2UCJ8A(KOG'T;=.K9WSIF>4/E_ 
PS ?#MM9_./XTVC W=5<C5D(+A%G3&$!;KO?-"*4JTV*P?VX@I8H@^^3C5CG&XN5[
P":&N9V%YF\!6LDPA)M:@[743V'=2%7M9D-R*YL<"]KG[?3(?EP')X599>9>F',G'
P!$'(LS$ NP$8TN^*%YP!@P'G</&Y/P 4&SF&5,I'.OV?%ZFN2Y+*K0B[:@"+"<P"
PAATP=!W.-B;LIWP?3 >?.73$/0JRI\'2U&B0AEJT?+03 MF5-N_3O,I]H*XOA31S
P_>Y=H)E"\_].")GXUNRB4H.@SE74#NR=J]T9#02+0%ELYTJ;)S&Q-M.+^H\-)#4G
P$>0PRN]O&4F0I@E]X&7%>[>K+!X4MD'DU>K'H?Z=BRJOV^VZ\H='-BDLT(%%^S.%
P_T@7Q(-G.C?C)/,);D%P?9J20#_M5^8D\[R%ZU2&+C<91J-SY<79Y5)M QCVJU[Z
PW^50Q=$3? 9@0);4?"?.(F"DB5,"(I[,!7MY%X,;2UXU3)^_C>MU'!2M=BX3C6W3
P@MZCNN<5"%.00]%#T:R1&9W_\!?L0YPPBJ95SEX17\<Q(_/*;1>V/WQ@C*Q>-;R!
P0Q_U>M.D[& ,7BC+C(E>4DIE2QX*-QYA1[V0"+"_7:>+]CN#P5^0B+Y@'"!6L!37
P=+9(,AMZ2+OH>"%_X(*L SZG(VK\(?W9G([K,6;QT9/ZQ@; [I6Z-P"YDB>T'FF\
P>F\$B'2-]8SR<^M#Q%,:-LBR9#[,0BEVTGZ']0X3!)!S?IVDWC4 ZHQ.'!I1K=OE
PS&'X1:OF."B5\@7D0L$'[*?H*D(JDFC9.I"S3R'/LEV5D$\\!:Q2?UZ!E;K6K%%'
P5_(7?7R,)>,<_*=P(.W,/.IMJ0A<7+X2+&1"9-P( >Z #Y*EA1^(>NF>*H3R7.Z,
PMV[%;VY*,J8190H,3%_5,NW3[OE0YQN.C*OUKEH]ZH5!LM(GH6G"BP6WTLCQX6L8
P'AVC\M@%4[C)_WL+/:UYM>A7%U@I/R+7H.[61".(0J'@IK"5S.RQX8>-(AL69R'S
P).'YU.> =;$3??=O"C4AIJ@X,KW6"HA#+5U)%H=XL2-&C#0Z1TG PUAH*V[,.S3P
PG0A+E!8:9+2<5D> ;"H)1H_@HRE?\W'O!KW33,QG!MANMZ!SY>&_JLO@'(_AFY>V
P@GELB3.EF_8$^I[,C2&Y5;2KV;QDU1U(&EY.Q\/<<YQJ2T###/UP1\T][/\/NLNL
PET9JB="5H> \-T4$7R'$3(<O#@VXFM!%L'MPMPSW.Z+2J>"/2A'TL@R_"6EV/G8Q
P?ICQ"Z$OTBQ1P8<!<6'WX[JV *#X/;= @P1ZSBU]N:_$;][SK</>)+WR50+KZ)"2
P>WB+V^[AMLL@0'^#2:CSO#"V62R'%7EOMXE0VLB39AMLTB),_B/:@GQ#!_7>"8,)
PI1PS>,%0/OHU[O@6Q/[!AU+C,6FZ[)3$)H1SYM!/CN^A-1G"OWD<7WHQ6[\M]:UJ
P!M80E T \%'-"6KW"5)<B-7V"\7&MS)2F\YQ&64;WN$*VS\7T^Z,>G ;ITY/F_<9
P9.(OWO46CNP,Y40INZ?WJEAL;J]RLL;?M5&&?U2<X0P[E+_T+*BC?);M36C^:QS5
P6V.;Z>!A:%>]6?%[I^YF<]=<J,:E4*13D2DY")9\PV$^\RM9;MH*XM86A[M//Y4I
PAZ?H(\9SZ7\F!_8 [SJ"926O*+Q;^W[+%3FVG7DG7=;'@ZT4D_) WB,V#T0B>N:/
P42<PSX,6>Z! LR[0(CF,]L02"1Y_,(]R:'B!&N@U<>1U<8(5(&=XIS.AOG$?=;^M
PJD,Z!PAK^%J_9%GY!H(,0TI^%?0'+1]&&S.,[V&NXLXM,D+;S8M70$="$#*L5]2;
P\0$FY?[49>:EXKKMACR6Z1D('P*;&\G .>%!H-&\\PU#2,.&BKNK>@0^C0 K8EJ*
P;J5I>*>_$%IJCR"V!D^L6J].-T(W++P)R\!=C>$);,*Z %A?FBNU=O>^R;Y>T0B6
P$!S/5-&(]MY0L:*]EHFN/M)9F?\WYDQ&[N8D<=NQ)SV/<$^\,W D*;#PM->.)KZ8
P=U76#-&'8+_22RW#*SU!U5 )I!BV %:-=J3L1/EXN6B->>".?-*QM>*%DE:T[6&M
P+%*%'T ^*%(8$^A-2WY]%8D2&1V_D9OD G>,(SM]SJ5S]./PCNPJ-<%"\NDC6\1)
P9U=4>2PAG7^ #WPRG@H=GW_:*[H<]:_X#NCQW.L9FC](%Q1?@]/&#['",2!L#78C
PM4;[ 6T]MOC,]N+;WO:8>1J?L&T5R= L&I;;CJ8.9MU;V9B"N1U<!;@^;P;$9FU!
PR.C?'CSS3M>!D;S]@(39&L\#"-FFVILW,MBAZZNR<3_X#T;8 =59/=:CV/>*GO'A
P60H23E.7(.'440^TD/*BY'69EY\;D]D'!O0O'-E2*VN$B@_B?)!N!GBVNQ Q0\Q\
PEQ'M88GTIAHV]!.=R\7[6655,G.,! ]-[[]O/%["?HF@\.!Z,_KENQZ07^H<;(X$
P%G,&%H'4 !+?D#3)J=_NTE,-ZQ1J<W]PD'-73B2BSI]*Q)RNNB'8VF&D2>_:RMQ!
PC67:85WY 0CZ^WDS*4$;;(41E(]=>O;=O'6F4>FO>CR_F!*7L@K"U)FV9AB[4"KR
PA'+^U"/:NBTU6$9_KI119?P<\]!4J$&_LP^N)GGV<V@E+_>4(KPAGI $+;8C5K:8
PZY=$;8:0TP&$>_)SK'NGN!$J-O$#1[1$0>GYER[#/SQ;XDQ'9$VZ;05*8S9'S[,D
P(: G58.VOK#6YVEMTX.E'M._U,M26&R5#6EVZZ/Q)H%* 0-Z,V:L.K&M4WD5RZIP
P0-E,4""OI@&X13I4+$#D<<*<MW-D8ZA@>2*KHY&LU]@+,"X\$"*+Z?3Y*P+^_ H3
PGZG-2-W(C2;55CNVZOD\U*LA2/8PG\!JK @H$)?_HR#*0I#/'%E)=UXO.[3L3=9K
P^<6>UZ,XR9QF#_A=!^I4(-J&T1^/)%;<>$2<G]:U\1>4)D\A]4,<'.>>[QIC.3OU
P]J_7W9=V+TCZ?);]S<$^&9!K\!MIQJ<ZQHQXK;JW\N10[B68>X*\^T!U\3Z1^WV-
P_B=F8T& I/21*[I>44([@T^V?8"=5^A1[&9QW#2>#LJ3-SC$XBV1$>LAVU=1LH,X
P>4#E?Z-$>*WN,P>GWWF4C^.]#I:' MBED@FP[<,0K(Q%62=?GK;K"<O4]3ZH%>Y0
P106YZ->3F3[IH<(@=*!MI2B*;@CE->R1/G;=EO-JM4'$/3KP$UD7J!>R2M^^I8K:
PO.U)OX9L<2ZI,2!7@,A@P+[!PWZ0W=K=55V?/>=CJGJ"M+Z'>;Z!L^YF0*$K;Z:$
P?0WFE2K-:DDV$?OJ281[:'.+04P:SW>8#H@P5B''&)$[(.%'D6QQH).!1.G<E6N%
PI=9 UZ#$3RMV8 I'KC:)(X/C1']H\%-"=\^+W@YG,.G^Q$]H MI,;M-_K',R)]Q*
PC3=T_15S"$+I:F@H9-8JDJ7/#[U)L:VDI33N7/"'E-F^..%MXQUAS'$W\2\DD_JY
P52!I ?"4'=J'LT&BXBO+/3@,AS*O;-U.DJNG@:RX)GE)V?5-CWG[2HWDEP\4=QPU
P.2N_:*-U=HN$)R;DL/-S+"#]SY$ZU3_LE&9+;<W],_$E6S#;)RDX-_S_4_5PI1.;
P7%L%8E"4_2*')NU.<=#:$NE6^9X^Y1R0B2&%JT+U'Q^QTF$2YX&Z2H!YV37Z3Y"N
PH!P'8?64*O #VZ:*H0+S@,?ZV0TQWM"9U)9:@&K[,/[,]?(821&=8%@[ZL2$)#.%
PD?/6Y3\HH[,G102)Y#([F8H%ZP=&O/NZ(03^BO-;M*7P[_D9V1[H^!1E0(JD3E>)
P\P9[1QGVJ<0?,#FWF*SSM'*8FE.$<Y;*B@P>12NU<TZ>TKPW7@U%UJW9TR\ 6R:@
PNC'Q:3MI_99ES'24"6&4"G!*_52&,S&MF[W_<PCY\4_,UR!D*6Y\QEKC;[TI66@+
P?GBAOE6QW<++1&U5+:?C];AYQZF(*U\D\BGJD+A#:!,1LOX#&4*U;U/E9D?QE0?&
PGOS:TK%0VQDL\A6@M0Q*D5Y_3ITJ92R"P</B%PG%35M,A;TE'8%\!2!0+XL9P\ZT
PF<)>+R #:V@5TSP*).^YZ[L2$R91Q[*>??ZO7VLC3!I_:+J*EAG3_@R9E@@O%.J9
P2A%LX5QV#G1RCL=&S$R76[NQ*$O!PB9;3K%4&)R#+!M@A+<CU9$1*7[&"!*.SE(P
PW8Y$A-<?=^!HMMF6VBWF;*)0H-1[@3R\\<;>G<%XH$"7:'ICAXGJ>HR_>/9D1@]'
P=H6P0W#"TQ""[<"SJD17_*$-0(1#S(W9)/>>*^JE@GY1!F"],O!A-_+ZGE!JY%:(
PRJ^P;#8@%3)#_H!R4YL@":, 9.L]D-[,[5_U]4P*5V<)R9V,W!N'W?NIB_#=M*&=
P_/R2TQ-2TTGG('^=J.1J:%35#E< /8Q?YVIUA$Z[38<O 5KROH^0(+89[HK(6R/D
PFYW@FY_@\@A7*^@Z22RBA(^#D"&5=0"N&67A/7=.P_+'C[!CR/64+:*UL=^[(]JU
PR$FEV1/?UUD3=\QO@&M102$ID9'L. >U[NR7OIG^AQ"RSHA/YTZ800HQ$S\)M0ID
PS>YRIH=;U?-O8SF5UROA?A.6[[LAJQ%1H*E94KQ#CB(%N'??H96CP>#/A3IZ,A=7
PB3=N1)]8%]S Z*4?<TL0?.#,H5/+B!24CP]=(Q430&50.(N/%3E[$U8F&$@6TW]=
P[<U)K(BHHH[Y!2-IH:A -"N^<?<?)KP=WR8K,NG<H@CU#"#?&JFWHE, M>[I%1S:
P;<!/RSVW686X-]:RD)UYXC$$,I6+S_:YA6HKC?C^W-%\RQ^SWGI.3&H.LSBQS%%7
PT)P:$DD\T50--U,_;\LTZO4UBR4*L3!':N5*4IR:P\/L)X?K*38+YOC5A<^UYC!A
P.R1/=^RQ!%#,U'U5XRJ6^I&A4Y6.E #4EO%?!&0VQQ4W=NH8XA2K,D<>E7W]NB//
PLI>TAN]2)P6Z<6<;NQ_AM[[<$X\FC']M+C>OFXV<C56TL$F [95@7(^XM^G'ELB'
PV0MXHK(4 SAGH(_=;LD#F/PQ6J(7X/LM8^^CWID^S5JSB.^<)^Z?8%L,KSU<@GV=
PF,._IYH-B=R+R/*ROR6C]'J%_,5D8=&.P60&F+5<K(<&F7?6\<R'4Q !!V03TFKJ
P^JRR;SO!''KCERA_C39IE^J)X\=D-_P6 .G#(:NN*!#8I(!-Z.JTU\/!K#5?I'O&
P1>E\W!8W7)/D%FO[<FX%-4@S<FJ#KOU^Y/_BUW4$-I!99="WTF6/W6JOOYPM%! ]
PVG,C/KHUO/!.'\6X=,P(]GL3A4"NVRZ@6/MG6)DYTLRZL/:!0G-;-4UL7P$UAN)X
P>W&P[WK(DZ9AV2O&U?VV]".Y7(I)&5';57F4U:&CAEE8G]HG_Q'3#Z*,.T%0)%W6
PKEA:!13:/%&AGD>_^3OG4$C6:2N:)N92Q!4"QMO&RYPZ/=,%,B?@=BG8O35VUO^;
P!1J LA9&;3:F+%.>[WX 7D8=W[9VC/TDF,I?:JB I8,;Q*_6)+RUQM0QH0#I^#N;
PUC@ABDGTY.%Y;Y$#JOU7D=,OP&GQ+25KXZ/: X?TM4I\,M<99T80:9E0P2!U3&[:
P]9BS3!HLAPBI9'^)J$K;X[LU,:::V))988$VP\4?77*_])6/HKX<A,)(01%&X<$U
P6BG410]# $[!O>SA86>!&ZY<F1$W X[DV2@4Q2'HVP+*=&!L[.&X%<]0GSZ+P63(
P1;V)8$&-J"X=UI=G4&#K0J)>]( 23RATH397:^RQG,TW34_CVOOA^OM?MCA7/9;F
P2N2OF[@$=+?"Q<. CP=M?MR>I)UI7<XVC,6&5G=^-@/5]4>#, @]&DDBIQY-WN.P
P-D"F6ZF6,7$]K$(P5_I,?<+#T-.'> IL*5J K;0<DZ090A%"[A2=.Q$Q,E2OO]XO
P'GS4(I@N3B3%^K@-JIXR@K>H=/I@9/JI>T_F"L8!A;<S7E!4?,58^<FHIS%AJQ+J
PL5YM/?P;-4]QG@3[DHMO\MS3JQ AS,?D#-DG0MC_^U"6*Y]\X0W#%+/2-(;DB61=
P17=N^V S^@.@/&R+R$5;FY[;9UP#"0G@&F..A=%[JUDVSSM21LTJH?2OADD16*:-
P[41;(T!;'[G=PV"A>C:/QI63=[5'RV_HX.>?1ICE:_+ZBM#A1[E^C*8M(7I4U8@;
P3EP""Z!+=T0%=D$>0H6Q&SW^ZN+XS&'&6)TBY\,*#F^78M$D>:#OY!K($@%6EK2#
P6&-$(1;%7;80AAM7NQQJC+VV>%FP "VQA(0.5DEGO_3#'!F2JJ+'G2B)' *3;'(I
PXBQWF(&>#0X),7NH"Z[5#5ZI;VZ6*=H9O!^* 3RX=QD<$'V-9B6S?+:J6YP]NVDC
P?*:/LFTSEH.7$SD\($$::6;2#H"BY[LX<?YX%&L(YHA3(E29-3./ZR@N> K;D7L-
P@@0]T]%%@5IN'H?P57:[E;<!2DOD*TG.<8<7@69P9#JPZ15V.TB/P&RIHMK*M&]R
P<"%0\S,,4-E;VAQ9+#!6;93IK1XVD5?^K>(C64AYV,Z#C(._<D]"BJI>2C#E<:D^
PG/WB6\!2$PVF&WJH61^#N70!V4<Y1N:>B[KSJUL,BM.)8>"O@SH'7+O3EM*^--!I
P\ U17?J.4MMU0'Z#0I7%V>Z=)IC^EL1(GE;N5Q^Y#Y@D('MV&E] :%N_R5.WL5;0
P4/'U1%7[#AEX]6E;SSA=LS%3I2QK)A055;:1J*A!PW$MJ'Y.T]\QB,OSB+O\@V0X
PBZFOB[D((ZPA ED?#-].=R!KE(-R"-&XXI>3Y:$-G4N9(U1/@W63/MA ?7IED1:0
PZL*AS0&8$T2BU]GA_!4[0'H3OM1,28(0-*;P+E+Z_$40O4EYSE=:9]_0#<YZ@-H2
P$+W10'14F[TYW8_JBE5#EU#C$!FI<K=R16I]FK[OZ/IQC-5^'RU3"E5]'>H'=($A
PO"L7TG.5+(BJX">*R!TD93QQ_.O#[<FG[Y<7VP7V/H0AP6C'Y4?L3]3I^U=70<Q(
P5.*SK\*"()8#Y<PXVP5Q;>DY/#.]'@F#3);7ZR#[4LL^;0)8ILX20R<;$QJIC(SV
PP.[B3YOSB040 0E6994J\R(5UQ:W#14"O<[&'T18.(@T9>'<4+UW>&YV>,(Z/8>$
P$]Q#$U>IC83B1MM\H)[_O4.!Z:-4#H$-HZC<2(TU<'DXQFN":O'4B73CF-X9 %RF
P58'>/I&(^];"R)H?E,\LB4K &; ?_] Z@//2L4YAUWOTMG".(.F?I3P4[M1_SM:N
P/ED01 +(N"Y,3 6N>@(Y.%)R$9D.O^D&:1M(7NK9M98"=#C:["0UF_.W(%S;$>.Y
P0A<_1/L[!/B"I"J ,Y)85WJB:6,Y=C!V>:U)K20Z^KV*P'7LX7C@.:7F>#.&SB_3
P%^NW$J1.0:-+G01QYS%NA_&KN[IB^.G#84#CJ]'?T<LV4NL7JOUZ&8/6QMP,1/X9
P<AR 1)1Z_]X>E0F]!9U9)WUM8X*I=)I#BIZ!\(_UI4A?$X77'%8)W9F<A&+60?4D
P*"$*LP@BKK_H%>!JB_/AVHZ_/%?M32YEA<13?6".][MIX3XW[M?^+'1,_@YA9ASG
P,'8W0 Y+4*8NL?[>;V&R/@*9YOQQ(&W"5=&G*7V@>9\T9GP.?;SF@7]%=L_]O-I9
PXQ-/*)6J-1Z#SH)1H.#AWS2TZ=PV89_/_(939$3F</D,;8 [D64EX0Z+6P41J+S9
P>DRPXK5-TH4((3EOH3QW]A C6Z*3[[3LM@8(@H=>T]1]5G\?ABYA_%AI(:@-A.)H
P<N_[(1@F+86-7_L;%!/NRZ[TX.NWW=]-K[Q1\'T4D8C"B,+586>%S#&K&;?AW%AC
PG\P8J9L;T@)9.+_;1DE"DCYL?<T7SWF*U-FAIM^]N6 9D..8+*<E0YEE ^L"J-17
PF&YBBJV5[,$YN#A62XF'R;N1O4BA.S_O%XMA.A$)+NN(#\+OD-4OIJ%5BZW.J4]R
P]O2Q;F+YJ=T>_MREIJE6-&CIO><8ZKD+&P6'*.[()Z050"M[,SK!"9J_#V.1UR!W
P[1](Y'>!P.6227+[%HE0ITW"$$[\\V]E6N,/CK5_;@8&Z#V![KH3B$MT!>IXOP&;
P**. S:I(.C94W$7P$4AT(@M43.D27D!7Y$>Y,25Y4'59._[MH(I 6L.!;@F#.0L-
PA-@'>.(=Q\FK<>Z5ZZ-W-X]7$P?[]>_U^-9IK/3*)A=@:+MQG*%QO#?4P>@4I+;N
P.!43X.(9&-?J2\X=AY9^?/D6VUD;^O8+'\;)A*H&GW#.EPJ]YT)O/WV/HT^<FB5C
P :3$2AX"$-&.K6M,SG":NH(<H7WFI81G$&XQV\X SH-"M0.W7RLG># BJD3']A8'
PM) Q/X]IF9)_ UH$TAQ7N7/M#'%Q[!W7;GXJ[*H^W+<C"<C:YYQ6ZVL2Q_#^("&8
PC -=H(Y&-RKC38K &X+<^C -NLY3&/T3-<?LFMCE?93B<B-*H[F7EK:WC/+[<%_!
PW?6HSH@CN$"B_,YU%$W'0'.-2Y<?"8<@[]J=E$/O3F7JD86H+YT:%C0.!NV(7QPA
PM)N7%"K4%/\>".*C'1:%);)X_D:0C62MO+QBGM_K#!(5 \;M)_;F+UV\&*_TR(?1
P:XA;#$31(S0W,X3[6%@%X38U"]W=V..X>;AV8L?&)7W59YJKZ[ Y]]2RPE4_;!J?
P;K<ITG#3TU^%O8\T'8 O&"D/#64MC&I!+/3\;H2<J([A/SJ6IC'^7\PN;<OI&L:T
P@Q8)"__'K7WC-C=N?'+O"QHCTLWL"B0:F=Y.86\RM5:5IW^52MK,?;_C,]%ZSCM8
PA4X:OQ/1!]]Z^(#7G#GSP/F>;:%<_[DQ1S<L0K]K^0I(H/=_>Y5H<!M%74N\F'GE
PP]ON+_1;F9'AK@?,4VFZV+A4]V"$+$$?2(L%V<'P*X/U(/IF9>+4#/'_VQ$YI# "
P?,FGF!YIFOM=+E)5ZRP$WF.[UHE.N7?[KQTK/*3,*7+6>O^UR@">A@*T<P#417?5
PQ_E@:5A'W^* >=OZC1KR?J>0*]RB(OZ7:TZ5^F1B'046>'WVE7UC](/2I=[C#__"
P>6Z<4_&_'@6T_TXH$L<,]^GM_OO])VWK@1AW9(V*-;E7:36PW<V4#LW;N>0$A"!V
P9O8*X+W,\S@*;"B [G]BO7C6K!WCQ@:+T?U'=':AYL4^$SDN T!P:Y]'=.MN@CII
P(6!U:;#<(5A#5G G"N<&$0!Q]"K6>O]]0:].)-<T+&X3-Z,)J]Y+AO:JM7^9\.,,
PH#VGDVVY45',1H.IV[Q:KP48'PL8,M&.D&N\]>$6Y3-78+*<%IW<6#_7,74D! 7'
P/16E(SI%*CK!.!Q8:DFM21E!N%T$6]TV)X_>2T"_5]+#<;3Q#P&]\8$PO?F8Q)+?
P4&NM&*N61]<25 3 !B6=0F"IBM2C9UWPV3/#C#QAV<]"V%][[2OAW8D?UK^_:!G,
P9V,8_<V3D$9?3IF!7ND!^$"]>EO:IMEX\<&3\=1+>K$(BLV,PO<I/#E=4E^V8!.=
P./D]JXLN^8RZCXDEV50]N4P]'B]0O.)#7M_K\E$OUZN9\%*QE*;>/X/W!0/3Z%>M
P_PGU3VJB*P*:PY'29[/@I7TP;)),[2AU*8:NF 944>!=(?3G'PD11).(TB?%,6^-
PY+ZD$ZWRNT,S?ILPZ,BZ:"UO\I;3*CS/&,H:ZF\:<MJ=^SA6(0==1L&T(PO(&$,]
PFKSZ:]/FAOK>#LW;3M<Q,$<-*DBIU1H#'+^R'#4#&XL1S-F35*&?X\8Z'5_C:=! 
P-X!Q+OFX5JAI++^!^^@@WPCT-Z1ZET(&BAS^DLHB)ER<FDL<;29^G@Y?U%XLZA*)
P4">3X\Y^SH7\3[EH=A%9(49QNOO0.;@<7+29-X5JK@H&<T<^8>%#G:RT7+_CPA;]
P[C<,^WBK$*UWCS5^LA'"5O'!7Z*X.B5!9 >) DZM]>D<#"4([HG0J>"5H8R>:40K
P:'RM]Z6 )#N/&OQV#,=Q:[OY-I23A]R8_G%Z7GY["8U9D9M)[-I/]*Q'MW%,3YM5
P=+.01CKIFEVX?F#_W86))=GM#CU)SSP('(<43/24%4 IACVY #KOY\W"^HSO)"44
P.ZI5H>3#18T;\K2C[.8ZIS]YSDF/T$J#$/BP_S%?E=K*]WRY-B>/70C%_UHF)%"P
P7]%WS![@(=2/4KC_.EP^K,&3^HOS9X[" JA--TFU+SWWGM:@P;L:@H*!;?T8W-I*
P<^)>UN]N;07E$49^D>@# J:\RD*I8K G;WE>3:!+)+0Q]2I4-)Y4?.IY+VT)JP@1
P\(DXTT*;-PDYQB "BP (K_41,S1 B]2-M=*NZ^Z71SQ6V;R? 8(X<BCZUOJH?C15
P>[P1MR;(O C<$2XWUV,^DO*VN]RSB?@8[Z0$M-7_?E[RJOJLT'22MO!-Z%?Y9AS@
P*<B+&).-R7[JI4$-2B8%RY2$6"OSNA+#D;=_3 -?J^$7VS U:-?U#9CQQYK5-KI!
P&T=0[Y[4V&A_?'@RPU+''V.0,FE,1(L]9R>$T7$XGE4[,JDT.%@Z00"IO9[AJ5<T
P)WJA$#ZGY[_UR3JHHTJH+F[V"1M)'89(4,O=Y(TXJF['^);-E4.U:X&FKAM]EE>K
P!12' H*+KP[/+N$3!HT6S8$3K>9&'I<\ 6!"]'KXCMA@UQ6W]HC,:DA[<YT)OM^/
P(W ;;6=I';E6BMJN0= 8O\ *)8W3!%^512+0B:G>9C9@(9ZT##UYO+GTU/T>L0NT
PXT_Q438?-!VWEO*\/2IS8OSX:%"JQ(.F%JW'@P^>6DFI5)['TZ:YG8A%S'%\W9DD
P59GG2021ES.=FS44UN9H$[,PALU/O%AD<@4D23<#U2CG&I!BTMAVIXPTPGU*G=_N
PNRV(ZJ8_.GT/QCZC<_&[KJ9!*INFDZ25J/B9BA_?52WSA]0^S"IN>^F7>[#/*%&6
P>_W^O)<'=]^WIRA6=6]MWY7+4D_5?YLE"N[S1L=Y8\$UYSVI%C:_XEFEK([M,9QA
P 7_6C]+>G9^A]2]?HC2$:)(X$4EP5?F<EO3N2AK];-R(FP@F6E+_?<3&%W4\"&#G
P 6,.'&>WVO3^.R#B=.G:#VQ>==DKXM.-3%$?AO3LQ6HV6X (JD3_B'TS39E[")!7
PLN;X)?R9.KU [#7,EADAO+&MLL,3S)#IK*1</^Q.0")L<CSP?B?]\]C5OMXX4.K3
PT'_Z$U6(.I26<7O.&\AD[?*0^"AX',*+>;YB/RP"+!_@-A[OM*VD66U981.+TQSY
P/).ZKNM@N,@KUKI/?Q%2]3M=.;B4L]L[)(HNG_>SRHG%TT\H]@[7>1I!'&2: \>$
PD4H]OUKDDI(5<6=3+M!O;^OKT6&6NW_Z.J1 15>@D,6K.O0%A(.4..I)P/-HBO1:
PA9?W26OZ'=';0HW;;0#5,6%P4Z+ I?;F7W*G;$X84 DVI94U(93Y ]NCD;7!%;TI
PBK\:6E-0HL]QQEE? 7C3!K3B8DSUJ=;+@OASZV/+;!6;_LQR!":\S>]LGT0FF$=+
P>[' =\4P/&I>,8O>5//:]",WEQ/__'G]U)!U*CL= 1((LRHLW^/Q\ZJ\(Q6%/ILY
P$%&8%N+%=O;1U#1RHC9F>=!U2[4"JC5%G.@@@!M9N@87BMFOF>%L U4!SGSMSZU'
PNA^$X"YIP)%2A\X!:C7(1@-/-$91-1Z-@X9\?HI 9JS>,B@.Q,]BAQ3?"T*]>=[D
P[.,H/K5VS7PI0EKG(@*K-%[%ARK1 M,W4HY-RS+>Y2+W:D.K-[S?6M#2@:NS#R$!
PY/36'_5*9T5^*Q#XMS7=AA16MZU/N9AD'Q//OP&SCYHRF1EL)Q\"32U.!0S<L78A
PHA@>4PL?H->)TP;^^9CRA1K<-B)/SMH SQ=XQL;(S-*8!PGMZ1<LB"#65[ 8BS9H
P/LUONT1%J6=J?\VH#ER=M38*$PZM47TB&&$6L#S?DRZXPO[0R%1E\+>V6'7.F3NN
PQ-6K=6*S+L+%D4YF 24-EB%U))>Q;31Z<[/#]$=;MU!PRRZ )F+FG2P/@HY)WO]W
PROOP^4L!1?O6)6IA^GCPFL)4(=8XK+[-B$#O= 'X0HUX8"2K/U![643]$\O8PBVB
PA/PJ(*?\N(<T^;#S,%T7/?R\OHO;KO]5<]**H1+4YIR-G+I-$*0F) XZ,R*/&/^,
PC8DXKO$ODER"JB>GB&@!?(Z?.6#=@%=6Q5YDG^PF0?S_*I,&FWFDR8-!"B:5<;Y@
P@;NZ56Z;8(5KMN^!U0 D7DC8[)/--O[7#L?>;53L/*@DF\S\7.=W3GL9QA8RVJ;6
PL^?Y?>7*^_7AB6:%_:B+2CD6?JN!A<W_QIXR_+%@=L8(?F)&F4M/**N3@38Z6CVI
P3JNMW),^M@/0UT]G=9%6IB&Q[4-^@0-P&"CEIZ)];0#UD'@\AWLUY[RZNNFP+,(G
PR8QP &HJLRM4B5ZIW]"<?_5F)CX?Z%)Y=((AN-$/_9?(8TAJ%H2[XF$L_2SB8-'T
PAJ@2B=NRROUW>)5WR_E=Q@*F*V]R%K0'A8+$_H=H"WY%)S:?3EJ,(?,GPXA2Y[;:
P_AN9L+ ZH#);R"3E.*48*9S(.$AQ: $Z#NOV\!VHV;<CJHWB>^A2\2AP.A"R_>/I
P)QBR2PD%;\SSAK2>ZXJ:MO?C;]&O/655\F<Y##C#LHJ'1 ,U!%@V9_\>A/N/LKXU
P-Y4C, B+F[?$8&"8'DAR4&=:J08>-;;S9_Z5X"',ZPH3(65);:8[4S:Z0E,K6+._
P(<EGGH:K;I<>8,A-J6,]IRF0!23Q]]D=[J]7N+WP0XH!2D(>GK?AH#.=KL0FE4/Z
PN07S)&,+58BG2$?;43S\XS.O9+6"1MM:JA(1M@40!PF"%/#A!4=AJ1S9L*/)/('9
P_2_C4:A(E;@T+D]WA9"5DA4$]DQ,L_)M-PR#BOQ7+$&;HF'+AR\W:A&\SC#C0VS[
PV7>HI1?SX9RGPZE>F9,46H#(; 3+PG3;"+ID(LXA1PL4(YW!+0J<NX*?9Z*I<HQR
P*SZ+;9MX(AJXW6I7/%5J3 \+EU;%FVQJ*Z[1N\-M.L7^ESZ.$A%*LG3]?*_FH#1_
P+%+9BWFI$%(B/JFT/P;Z]]FED<SCIO4MB@DOJW=L)O0]"^D)[OS#EA*CFWB(*@P;
P7HY9FC*'M%V9JA*FA*XH._D8!-W8$-0OU7WQ[?(WZS=/TKAHO7+0G_@YDQ[ 5]]E
P!HN*\W2-#K]HN^:HYX$]Z4%(3U$56ZNR+7#S1G=IH2_5@XNJ*H33Y:KX43A?ZU] 
PLC":+P5&2H3PMLG#:DVRZH#57@[M:Y>#7==+7G5?L,9!?M\8D-.7@WK%!5 Z+MPL
P--!ZO1V)"_67[$S4H >9,7B]US^+ *I$X2C/;HB41P7:YA%=+Q>WIE^^!&2GPR_N
PX])L,%ZJ-<VY[ Q[(F<%C(&W.H"$ZK >^83\)\OYVUGJMW,D!!F8YU_1N7_F?/LU
PA$ FIF0*RDH7M)T;G;@[M)#\E-7&D;.#F[H]1_'K_J)HSE)".XC+XVU+VD6"N98M
PWM-6Y)5/0NA]T:3R83G#VCN*DC]GB<RUJ2AU4&"'(=QG1+70<AQW7<1S&W!G""W,
P/0^%"U9QZYPPD0G&==NVRF:D;$$!$VW;B8A6\I/&?LX%-_XF".OJ>!GX5>*0:+8\
PB-T<;NH^U,D[S-MH^JIV4OLTE8I6*G]X#&\91UIU:K6X<,V(S8RGH"PO,8F__".<
PK9$&"/S_;LCI%18(SYS20O**LQS\U^Y5>'S=M@N!']^RA"^56ZV/>-@]\A&N9:!J
PODK_&:R9X4S$^^#64QWLT^+A,7=\Z<9%5/J!CPOJP*N1KEM\*<@"3VZ16P7%' (/
PWQA>CK#C0=^!I]85D#A>PQ>F6Y[+"=4-NK>'S>/2;DHW[1=F">M[PP1YM,T1D.B3
P&:2U\@F['8(@*-@2)BB- XR ,LZR90X-Z9#C1^A"VQ8]6EK!4Y^(CKSKFX6F+#%^
PC?;#C=3#]H%[!4('"#I?7TH*:>2EA*^IN5\I*I+ZZE2*.*QW#\T&P@;8(S=U)MXB
PM-!"O-1M[QH\+MQP=*!V@M3415RW#WG:R"%/9 >0596"M:L@9^B7QG_]Y:K.T8[I
PN5Y_U91F6&/=A5NWXJN MF2QF,-@'[B714@!&E#YW<@[L700<3%LU=IJ8).(#^=^
PH 34IS:8%3\==4<(.O^ON]%[6J"2"% D7>_ES*!SHSRS1>9&$.'_KZBJO%\?O7T2
PV[JSR(:SE'WKA@V.? =D/O,ZN%8* /=\!+CL:LF6G!LJL"Y54DPV$E!'EEZ[E/1+
P67P#!VEGN?+<NR[)4J-@0/Q5O\YHO-(!NR5>V^9V$C?R+[F%Y%&M,R-)W]Z@,:OB
P'1+:][X+E  +Y? %'O,]QF61B.A1+;$:X;J;]?*^0JVZ5VD2KY8=< PBJ,!F@N28
P,*>7#GN]HH*Y)H(<K--=98P6\/4@&9AP!*:?]R]L$VXMUMW\9 *6W[^%,+<OHZMC
P@D<DW#2K&_G2"!M988X]3DY*F7+%680M_;3([$#'?*P5BG3-\C8)=HP.M7@,'2#S
P$[LG/"7,/58Y=3031(^51\6<WA8D.T4%)LDW"HA]:CZ"QRT7 Z2=E +73P,8U1L+
PN/WF*2C=FQA/ (W,P%A1]5]SN'O2V6I/:YPPJSF]RE?L=@!F4TM%81&$[.T7>L $
P3@E%R'@HU*&K<ZU&48R9LA4P8H7-4:S\T$9CUH4Z;^(H%31X*(W%&^J#]^=8C=TS
P!'R>=&W*AAUOP$V$2J<!CQNRE3.TJ5]?!1>U@JY%KSRJ7%V@\&151EO51OCMYM&)
P;[&5,?> U603&%S.6QR]NPI,P"4&*Z@>5MW?#P2=<>,VXB[5  ZS9P,+Y/E%_]QH
P8!'1S@N+% 49^M-4ZIZYR[=MM6+6GK79H$=[ DDP1,JX&N(^RH*D[<3 U17?L9>2
PE\M#X@A'#.R?23\\6(0N%!KGF39E6R]1F(/*]14$&B3,*P/E,SGHLXB+1&@YM:[,
PZ6AP_+C$5OX":(L)+2QUKAL7)L::/?S<'V3,!^HQ&)L7%%50(FK(^JQH+ !,D6:\
PA%;U/_F4[T]F_<)_Z'ZRY)]@6EBK'*O36NK#OV_RW?H?K4UI3LE6"]<:YBGO<JXI
PESOIC^9/@.;E^M,JN]\H DCXD!5T#%E;)Y&OK6CA %[],WP"!=KO#_[G]:LN^KW&
P]_N/R7H8F-X#9L,&60@CP&6G"[?S]%GPAZC^,5#IIF^!4ZR_^#QK7-B)(L_?W"QM
PH]4<U>$$,?F%_7@6#O#7?Y8!5R/H;1L_D-K$$" POOD.U%&S\M1[;4X+/Z1Y54N\
POA9[J0$GE/8[6/NGK$^46U^!MY[\X\V8;0 E>2A2KA&OE=)H[8X;*4Y7'ZHSXKVD
P).BL]N9UC"JMG:P<(J2JD%&QF1,![P]#V2(MA%= /NM R:X(<I]BZ7ZCI6V\D/3O
P=U7(%&-?\(&>BS(C#3RD5%!#;UCO3?05UR!8)"++2)XK 44$^)._*4E*P)[_-8='
PQ-M9,\,:W:E$2:^?-3%XNP\'UGA,GN/9Q'>WM,%A'O1B[AG!,PZVP)*1@T@TII@S
PZA3/4TZT04 "=/#)C+@5O%M(&,P>F4G;+0B'0ZQS_5B>\ 9,'M(_!R%$.>QE/U0B
P=M MT5&N.U7RB'U$NX"I-^(S]L*0EG,VX&"X]HET=6__TX0,ZJ/KD6<M 1F@US%C
PVY@365D"AZ1L9<\%77?GM].8GX<(;8\^)O.\%@=*DG7#*ER 7CWW4T_\)2M*QV2P
PS#*/WH2,N B/#(!VWIC.#5$T% ^5OLS(&J)I:30DD"Y!W7O(UE!D@HD(/ H>#)$N
P#/%L&7P;BW2STU=43Q8'.F74,^,OOD6!*C.*7>=A\QYZ X?)+R4B\7D1L&Z 5JW;
PG8L\1N51-"3*/"/P"<L07[332VV<%%K7N>%HI7-J/AL(?!85A"JE2F1&@!Q2O)!C
PE^]WL8NE%%%R503NBSC^8O4/N_U#L>5_B4B:C1"H3\8(>2( T([O18#C-4437TW[
P";O9;D>%57(+N56P*2Y)WJ0 YY(0^(PEFD-A'V(3^CY7%=N$6+I)F51X:!A$ 5>O
PC_J8JUWE]SH4@N2(;[-K2 7]"=8SH5#P\[G\H<>\D&P#^C5M*I"$OJ\%3/(%>7S?
P;8!"P*&YX=*C;%WZM"K@B?-7"8>9M^5RH/_ QM0$++0MF?;D'N'"-P1$?5[7SAI(
PO^%!>?HB#R[KL0T[R%5EVI?FITD^>K:@ZMA@""!CJ>AFZQ^=%5-G*7CL'T.\ 19%
POVAHG3 W+>)S((/TC44/BD.27Y?(S@5L_  58Z5_-KAL+(D Q'G6!NI5;GDC 6$S
P*^'P^" Y+M:5;F8;+>H?*SE2VMW[I%USK<EWM1=XQ3I5PUXS.WX\#/QS5V7LO@)3
P@T6DRFN/"4SH6J]BG6FC_F^-;VL:Q&6WE79@@\).Y2P()) Z=RXTFXA\ODU7FG<Q
PV_0X?-P3NZV3XS$#$-ET!Y1)UYXF:;MY:TWI4KT>XEII9863^GJ*[>,61%/S+GM+
P5)!.BNPD\8;\=Z2(=A<;5L)< T>?^'L29N;$!'';/#VS%1:;\G\7G(WTJB1VK@J3
PK0*"S)C*"\Z[DXFB:\1QQS$DR4%(\-?V=<64CR:X+5;3=+9"S_.2\@>/H%U!;B*)
P@/L(J@-BPJ>L9KA]-NMPH-+=X9LZ%#U:^0W[,I!>&X,7VP4F@KLUL;7W0S[DLB8.
PS9\S]/3^BW+(U3%8FZS[<P2_DHY#.XLG/""/[OV HQ8"+.LP[0AT"]11B LJ::%-
PK3$7F'ABS-.4D-RFX/#<_"@P9A_L"KKDX&BJ#?T3X?H,VE/>X*'&N82%6Z]FH@4<
P1<#PMS0_]8'HZG68CWMU$C#A]TJJ8:+">:?D$2J"@8>.R$F@2;4-AE+8O47)(CL)
PV _7@SMC.FQNQELK6)-JV-[?CK^SJCS,Y^9<X2Y23G,48ID>Q2CS7MM,W94OYM=5
P\]DH*W959@,5U(6EL!W;H0*EIM2G.;5AJV%O\(7)I8G-C4![L#*>EX>I.JJ6 $',
PUHHXAO)I;#[%NN6N>366#R_@2='4554)O_B3]X1VHZSA\.%3CVZFD*V[V4AV?*&6
P<#R--8YD=%^Y4L4Z_)Q-GO+S!\LK7(?&[.NO@B#A !X9E]3)"^8 W1 H'4Z>%06U
PMAZRF1H*Z2M#=?,=P>QFWXS,!4+T(E!E(2F8N=/Q$ZKS/O.-6R23!U';0I_/4;@L
P':A83FFES9EETYW@CRWD?FBT3P:1[HV)1#9,S2NC(+5.[YV=TFXI"</U@4>!J^J&
P<"5P5W0M!*B^W$#K'003;"N8<F;CL,C4C:G246-?-:^3I['#0I3B+\UW&5^"%@ND
P";\,JY]HBGGGWFS>F9R->]NJ<('F !N8"PR87SQ]"%\Q( ^@2JB<,(*4[=G:M?8]
PBKU2UZ"@M*SYHR!QH:I'+7H(6(W8PKE4 T*]W,3A5QY&TFM^2.A.*%%%DQ(KH[.W
P'(_PH36,3WV?RFS-B&#?O19(?W1 ([AL7]Y!4GY5%@&+[WV<[M1,EO_$<4Q"DNS4
PO<."+2=]$:FM%&YY#Z05OCA,,[\&NBPH]5*)A\L&H)E[V5YY:B71M_NL:LHQW<-_
PN/92;I<B@<I<7I%GAC%]6ARI*0;QU%3J6M1_R+A!T_J*-6":3<'<R&CU3$>>DE30
PW_INYFS((Q0>4I3"*/YO1\+&[$!!FVS_?YJ<.F\5&Z>_!:@F\8GU,IB(I#M6B^.O
PF;SS%R[J?WL>\OS$<-:;-I_JQ%8@@A([.JF8+B!5STC'II Q$B?G0#4DA &[W>W>
PIX6BV[J9#3D2V(9M#F@W]'%S&('U-Y_?V<'[$ISZ:(ZX)(,?I<+&/J:?%L !SCXY
PA_@6;GJ7_!ES+W\&)5(PI3$5/T'NJ4EY/*&8E-DI-&P57--*AC\_;\6YK!3T(]Z-
P4M[+8./)LN/!^G;8\#]:.OS<??VL7<ZF2<*^]>-HX'C*&F=O$X]$Y /@R\+A\#EA
P36"D4<B6F4%MQ<?K]N#!FXR3A]64S*@G5Z,,V-XT3P3&A *./(;J(8S(L:8K07^8
PJH#32Z?F_QUNIJ"C+DRLB)^BTV-V/-(J*V:;>!$MR^S \2"0;&TBAUK89(]3AQ-U
P*7,,G^OHHTF6&JL/0QHYBAU E:D6QS$P/+Y]XAAP?W&,MK&X]0*R<B%83%>KV&'W
PE";%X2+MMU#]>A#-[S#2"G(*WI8 Q!.9E:"B^]*-3:6B!]999QJT8&87IMLOU6_!
P]QAU*%P\^!\MSU@K#7\-\A-382.9Q)'43Q'6 M>6T85<?_["I.@ANCLBO0#HQ?8@
PE:-T1U4#,AW<&Z,5#%]7"8'"<.R$,6#+]Z'R]CAA='Y,N=JQ#D*QY;L$OC'R6-\"
P *4FBQRYT 8/P>R0R"ASYT&95,]F07>W3#GR=LBS3$-04K:?[0.WM[;/%U(%^!!^
P"9D BFD$1HMC)B;UO.XR($,)@@L]BHNOT $;CZ>K!T1K6L<F/F=<@^U9,!@MG(**
P] 0JRSR?X6<P)A0>".-#FXJ'*^ETFV$1\7+?ZF-"%%@,QN?.I@W0_Q+?<@9)6><?
P<PB))V[C/4*0+OP<),. *4?;)CP%,*YD[@O PU)OY^2]^*=/>A:](+ 9=!TI0J8&
PHD!_=;D[OBF#/$Q4G2M2)1\M/*V+2HF"X[9/4$,IC@5Y80*U4C3(]M/%79D>.@F^
PGF,/8YL9KKZW&_M&;0&J2?3W((GFSYEPJ+,>ISR8L'&,26/U._]DY@C&3><"^3?G
PWQ085C()B,R:7KWU8B^OE^*U'JTNN,9[@F]&SE"^$<TQDIK8#+;KON*J3DS7)Y(T
PCXX\\<\4X4\^/J G%M4\>,=T[K&"]'UKI#VQ)@+2>_(;&73JMVML8BPIJ,[5UT<8
P]EC*Y,$>!K0U%U  '.Y9;KZ:3IDLZ*+N8(+[=)U>4D<#Q_E60B3YG<,.0RJ2_\SI
P*RNTX:NJ( 27/^C'0A'*9^TL2#^1@58@L8(4W&<ZF+QU_U[M-SK0) 6%%TY\V?R[
P U@^D2TFEQ:2@8$Q&QS5M]Z5R7WE]E ^7$P_;WYRC]8%[5AEFR^4AU5P9H&XTQ4Y
P0_MXVCHJ/#IZ;AVHU]&V)U@ V"M^B;-)-=;&.-E8,FI1K%2R/=4\&;B9H]H;[W'\
P,04&Z05L!)\_P@;2K.*;.8]5_CL%.]W==?D-@Y9PL"G8(E#/G0N@27?(F\<%D *)
P]&@!R8L?3D6ZV;TU=X,6TQ14"[/%0>%NBU@%BRT[Y\03X81I *?G?K"!N&O\<6O_
P7A*#-M12<IC>4IX\V$PDI('.8MJZ*Y=GL\5[ASDT$6=E.A-,KC5S?WM@?GWL).Y)
P**TF/DHS7Z7GW1P!:+TE%^)""O"LI!@$6TIYID[P4%\W\='5W6/*=VD A-!UD\D_
P2)']83C;"/3[2=PUQY>9X9T9GV>Y4:25Q83YMDVC#Q#A5U*0 3Z^_X.^X)YR+CJ&
PK=#*8RG;DT;D)(\@6"-AKB,DK5#*YYR\NU'+V7O"?=(,I< _Q! *5&:=I$S@]1.T
PK]MJ>^5><VSE*VU<C/;E*4D9H7!9T(BM4L]'ND5H!6CK=.*42]<5/[\B8'B#T>E>
P_C,O5?2"!).(_YD5YQP>\NQ(3@:9C6]1O/<LQX!S=OQ#"A&J0>6-;;N]DM08<=5)
PG[K858B?+JN==#BCK:/+[6KZYR2BRRA!2"'^=UJ=/93K>?\ PGDL+$.I'7>PL;G4
P%S%N^KR'^!U>$99&3$I(##VSLM,_].,3T8?2VJ3VZ\;AXPB&U1X;F6=D[8HC#Y4S
PA'Z>V9LS J?^D!0&*<;'_S].F0E<-IA9-G*LR&#&8\Y(F$<X"J_MZD';I:$G DIL
P0=)1G-"IW]+XO&@1*A94=8Q-O*F&R7P:J*?K05VS]I$+_DIBR:S9&"Q4:?<63)/Y
P4=]"]+4FC3N=O!;TD(&'?;G>G*+HQ2#W@4# P4W4@H&AW9=SD$+: %+KUO=DA9<9
P$-N4P706J0<>)(P[*B(*S*BG5-*KJE ZJ$TET:Z:^K&4%!>5T*5('5)#01@$_1GJ
PVPR\FH4F*AY5)E;F7U<LJ)44R6$;9S&T#$?^"#2Z#&G3$3N%?E]HU/&1S PQI,T 
PX!=G6:GH018(7&"6GT-83)CS^3F*FXH9("&72/1-U X%!/'?!Y97EZ^OA.D8GGH#
P;GZ*23:8V&2/F9I!4XJ>'3JEQ,[.Y<(6KSZ&T.I3&<.@)CL!AM2I&3PS'%M?!M'W
PG=X$-^:NG/GS-@DCW#0W5()(D@*M^*2>)0_T%F"Y8 ,NC6("UZ"L"K]CZ@ZRAO"Y
P/\G]O;5&&U$.*04*,WS2#',_MC+RO \?'$;9#-*YQFY[XBJ-)X[O/*QB[D0S<LX=
P"&.HX-:KHH,.+R%3UU0L%#A]C^,\.08G%+XR]5\%T?<A8L,$P![2O9<B3TGCO[+3
P4I!89&G1[/MAFA2\=N%J9F"4PQ@A0M@0A]T7* %DU9/HL--MH OHD(+\&0PD+<+>
PY3G0YQOI<V?O0FVO>YFYVV\X9+?DRE'H- P=[C#6O5^97N++[G&Y]Q_B6=*"=(<U
PC#'?\MXO]%8&'U><FQL!BR2J:%0BA5AQALJJP .1LSE-C4AUM@$R-4)+U'I:%!(D
PPI7L/=4#Z@P;&=ATYIHRMY=V6!US _%?"!NH;C46*\@/N<CXX Z2.KZHQB:#N2B)
P\#>%.T'R@KG@__JJG*_0VS7'H0?(>J"6:JRU#'T]I/T8YM"Y]Y19X/Z(=CX<3*<X
P18N\@%F=7PX5B_^/OA8X!%+/?PS+1="X;E\9=.APMX:Y2V4>V7@KPTH:A-7;UV)X
PO!_0%Q$-FPW\$GPDN7IX?L8)[\S;0FFA5P@1=Q99O,.LIM 2%(26BOI3/2LE*O:Z
P@X/OE4S:G5;/M'!TH=K1R%8I/((88Y ,'$E*KZG%+;<X)URSB,WGJ/M*'.PB,126
PMGPBK^)&T$YZMVI>0GE2ENVS**51UMX?8/^ZI+W K _*IF2FIRD%9@C\40Q_K7Z%
P'SF6YP<I[$Y!5T1S&D4<&%9([X"QDQ^U-2,'6R2(7?:264X4H.^_@Y,KQ^^A8 8*
P?'0-U+):.[.]MG7&@M?7!:U\Q2,A?ZBE"LX4G>04>)[?%FPEE,CU"*/I6CYY)G9.
P!W#/05[6P9) \SC)3IZR.05%JP:XV>>A#W5I=\S1&TNL,@V5-<'-*#I8S.>@MX:/
P#)8(M<K#6GENQ<<&@3Q,%Z1(^,=VN0SA)(T*396-J7\4ON()Q%(C.8&%R4;;UV?@
P3T*&=S$8U]N=D^C5!+]>5["^BJ%(>2\G0'N@%(E6,72/.VX[:5,Y#.M71I\F;ZFA
PE_':$F9=]ZP #LATVT=,V.%67>?!K-C4& LS3.A XA05857AP66"V.MA5UI>?&-;
PM9T)W;>]<=O_O"6895.6#LL.<J!@,/#N.H2P4!1XA6*']:2I@KOI:6+RII\C^XO_
PW=I/Q;S0,KM 'Q ;R,U$-O&.ESTVHQ;)_(<B5PI2:\3B+.6XZR7S$FST9 +)>TXW
P7C^BVF^5D70EXS@-XW2 J%;T>JM^^1:;+(1;VT%;1+]35?MNX*JAY5@TO-H&9"L&
P+$%GW/@Q2XF'+#I\B"\Z;0E8^4]Q1=B:EO95"CU3HI$8-2U9_T4;\$WOT@YO^;;V
PT8Q4=E8\AH@LC,M4' ,YA5_CD7\_J9UIH/S'Y'Q5 WB("H[,CEVW4LO ['RF'[Z9
P#(K(C)'$4__^?G\PL_36Q]%$WZQ)!M^EANV*E-HS\5_"^Z-=3:[L"&//*M:/#OCW
P5="N:]T:_4>PS<[JFJ'_VZ1PV@_;E5, 4$)L,>CJC<Q"FHP MU/%>=;^Y[NZK8KX
P^9^C(K-.#"8[V!!P$!*]L)G/>/(!&8$ENJUO%^&A'1 &Y;D'?/#F8F40V"J6J%C+
P"V@/2Q20=PHPW0D4*!LS+: X8HMKRTOW)+A' [ME('%J2^'P+*P622G-6!^<C Z:
P+F6]!O1 9,[3J&\)'^PM#F8UG3[S9U\+@*&>0:;L(P&-)4SLJJ/;\NQ?/!O&I"L9
PWI79K6NB0S>/AU6\J2F&O:@MO1=[BF_$.G^4[.V4R832A"9V:.$*%K?,>\Y[(>/S
PYM,'4ADBA7E(_Y4<2P\=D:'DHP;\9$ P,7@L>PGFRB<=E>,!P#;LEF);>KIIGV[C
PJ(WY6 XF"(V'M72\E^RE&X*9CWKBSW[ FGVPJIJ.:(R9:P8AUECJI!Z=ASEH<A=3
PJ,8%X#7N!$*98[0QO==$_@C,-H'_G%)_O@MA ZPHS]"D[?;XSO+ [*U+5Y2W<#86
PGI,6I2Y&MDN&GN9OO42.0R<>@6'% E91L.Y 5R_T:(_)S +7?7!Q"6D\1GA2F2\(
P& L(&44'+^:(=P6]",@6['GN->ILV$O[VZA9H#+*ZX4"O1##0>V?3?9GN84T% C<
PY1PVMN@:-8Q5\.H_/=J !U$3*/TZE8RE+^7$6*AV4T)YW!RR=?%XD5K,9<;CJX?&
P2_:"L80+?P[;H%-Q!F_S!F1XW:".*-6!0R!5^.^S9_,F#&S4$X&0UX>\7F+1 H_'
P_DJ88?A!4AH2!._!TL-RH^)QC1SC.&6E;?6",,]6)W&V8%9;NY*D0WTGD#\#-D0#
PY0,[**#>&'8%.84>D0/U1EYK< W)V.?WNU<4XQKFK P5!YQI#+V.U$H6'H=2ELF6
P"7.9?(=0SGXUF3-4#0@'Y?_:>_@J5$:R&N$)'2BW,]QH$^'=HP$V.2:_"'MKU;N6
PU0V[)]_P3<FQ14RA>_-YB!H]PCD@&R"^<[MJ3(=[4S<YES4$N(]QW0IBH@D7NY3'
P9T/X8*8%OL_/;NX!T=9_:H..5CK'R 2-!\IHP?'VD7B7MQ3N1*#E,E?EJ)UX4C.+
P?Y!&Z)M<"536/X8U$F KIJK@5V)2$K[RSXPLSB;;4%C908/6@LO=S_LA;RCU6. )
P%Y7&=]/1_/=5XA3U4OYK"\3/25>Y0RTKNH Z6.: DLF<76<5I]P>_A[>+/<1'<,:
P:[[Z$E39Y3^.<@XF%'0!U;[DPUC#SFTH[M7]4#'G2%%6I-@&14%XHIM5FS+5$J18
P+,:S=[;P]%*8LGR0 #_8[5L9B@S(7 N ')-$ M/UAJ<JJ\AP)SL:-A/U23KI"X#S
P44I1\V(A(C;W91DHS]>F#TDNBYN],[562KU++2>-,L),)3H\WWW),NL34@!>B0GL
PK(??BE54W+QX'H%/]"ID0_TMNM A8VGZBPNZ(Q'0*W:,QQ=VK(/<>:Z-["X.(RL4
PD=J6;BX(P,\T>%PHDED-@DHU"T;]\#/\)D M 4A^@*+-!-&.'^*C2-#8+XX\NG)O
P(O<\5X'8@%DITV*KTVL3OXS!RKN:D#G@QH=[YQ)638IB4R[;N5IW<_IC[N!:YSDQ
P -1\XOAQ6A ?T(,211@)-]NGG(32&KYM-375M\!O16#6T*]1X*-\P)=&R^ E&G9 
P/X("A^5$?\I0\/S'@7@"+.4&U>N9V%-/GQY>"9:&-:(_Y&U=:[PN)?:_ZK4<[NN;
PF2[0<Q4WJQ&5:>#?83T*P9"#!-3?Q:!HGB3)R).;=V:%I%I9Y+AE5H1^"65][D\)
P#+M_G-:/ I1N^<M45 /I);YNKL9"'0..I*WS."4/ AT)?F$R435D*OEQF89@@TG%
P3 #LRXX>#95\--1.DVOG:7&Y>;V,W+RNPI#G5>"G20XQ?G4L38]D^-(HY#W:AT47
P)B'YH<!,K4SN+*5D3G2D5/($B "^<F/Q?IU"9TX?>.HA_1)I/]9-K\ -V#]A,8Q<
PUEMD8J6!U3]*JVVL!O;E:=*^(Q#?]5LN<;EXSK(<L*B>GGG2*[.SP)R3*#&JU]:.
PE?2L+9T"\U$01U>6>"0"NT2S(==N%EI'E@%.;!4THUL5BK"X^^*>] /"SMVA91V^
PJFA&282Q1*>?RE02!!:YKY -H\:)-#/#TJU3;-XX?[#<W']+(0G%6-M=+%L[3=?C
PY@]OVP7)ZYU3BX6UV(__P2<Z2R 1;CZ^+1S<$S1/#Y:<^2'_82VII#[AQKUF@5 $
P0>ZP=R*$N5;)?.Z=#T[COG* D*"KYWI!<.=A-KX&1W3BB,5"+".[C6;C @Q$?,V;
P5OQOF G1,K^]*#[,[KLSUVNN8ZLZ ]?4&1.%V=IW@FJ2Y@N+R&JF4@"-!S%GL4D[
P__W%P,AJZR'L;[1R0@:YOQ%GV*XP5/96_\E\?S\VLZQFO/Q;*6PNN)J/?9\K@@OU
PTP:Q(:(?18=\.Q*6VIH$ <>>2 _ &ZC/9N#M\S05X#(G9@NID3,B3^'![T@E;4]*
P?O]QJSTN%4=7\=*0[3@XHVC;H-BP2F?%Y)L;>9]^A)QI!)=W4F["+2S0S%$PV[:+
PQ[3N>&QK\UL]P+XX2@V,1[UC-9/-"Y4K<8!HR.LH'#=#4?&*E$-)EU,SI__[C1&'
P0>80>1@&=JII/-2KV[5F>9-O!<LE>_F-$!5\5O:Z*=R@*:80[&P@=OA37*/^\ IL
PX"FS&/^E<OZFTJ C_UNN7I>=P)G&&P%K+0&E>5I$7L-\E;8L8+NCG0;*"O3M8 4I
P[^)^5AUHK1*62:1>F.X,M&7\J"&9RR&6SR:!"5Y-6VB9I<X8A">JS3A<#AO/*Z;%
PLAHQ!<B(\[J6*W7YVR,5Z=VJO<,N!GQ@J@Q9>X!$PW@W^C;].J=)#O/NBAY-@@7"
PDCJEI"%=NUCL3"@JLJ+CA)DD&T5XFB8)M<L-8N)-U-PLN@ZMP89SR2,8Z!&,^E7-
P7HH)'7A'#04_AW8];I&F;Q#Q@)TAOS5L#Z)I3]9=[GH7WNJ'(;<$'0)\)6$=;MTN
PYE(_-\L+1\T0IS+"X=144HG<8(9_2^(T"T:OQ$,M8XB"&]2<HU#CSQAH0W0.-D7_
PXZ2-;$SJYFHEKXI5G@K[>%J)Y4JM8S,U:L<F.!KGOYK!JUJD4:[AQX:H<VRNV?#P
PG^,Y'Y@^R(+4H*QIBS!7[ZR70D6@EB\.SF<Y:O[\NF>Z**&1Y(P,)]11H,7^M5G!
P%%7)_ ")2>4NNN- !#T^L53@>R 4IRMZ+(-"F?$OG,A/CQ@D887;U/,K I?W;J]=
P192T1@)B\6D^K*Y1OC2':88,TJC@B(>V'Q%0JR1O3[C<>H:T<-7?,>WJRG$W-V63
P.7E: MWLA1:NN EO@ZS","R%R9^7RQBPV#O-NSG--Z-4"MQ-<Z@\4&9Y\V%>$<UI
PN3JT6<Q+8VE#9;+^\ER0M.'WC='_^Y@3A^8HOXU"U8R/N[6XATQN%OY>E7]]TDP,
P7&"9SE$V9?, <8.[\%OZ/!">X5L:2[KO0C*/5[XJG-N:."2]-Z? .?9]%:A670'R
P^88D&-X#!&Y;&.@S>IR>EZB8J[)L_7?K>MK0QIH<PYN=ZG8HPE()'V)&;_:RI5A]
PJ(6@U$8^AS D"*BDB[/[HI. 1+Y2T?>=:P"= MRM-)+F8(Q/MLWC.72F/FS9'76E
PE,<V7G0Q#AW_V:R:EJW+!UGN:R\#U5ZL8_8E4"O4BX*N8T'5@,)!HP"U0'&$W^C'
PL)R1:G=02;4S$@*S"[Q0Z\_V:LTX(+/O4=8B#6'U&ES2-/A =<# ,+,C_,@E>21%
P=YDJ-I@4RGG<"G9JB2PEK_R-TL3H:]'NAQIDQ-*SA7?>Q *ZC"907;KB5P=R,SVF
PD[4%?VD4XX>=VH^(_TY*7V,GT<MD=R%<:=8\7"K#_@TPQ126_8[G-\%7-N/)5:H.
P$:WG/EI_G"?82(%5*H9E+_3]OVD"DBX<&,P*(Y0H6VQC?!A+F+V40F%:,)-Z<\IZ
P;<.SW()4KKH-I38-.!_W+Q\FNL)5&%;(O(CK%J8E?TGNDD1G[WVT6ERM#*$5GG]3
PL?=RO'TQ<6RI*,W;@1:6=>\""0B'.]\JU6[V,7?'L@LDTBSG:(9&LX\47I-NBJ*#
P'F;XFB3HV$SH86K5>5.B "-G(((PK"#FHW/@[,2I[0;+-KH:3P^Y>>()?(W!2/$U
PN>"TB8+W;R[%W1L>W3R%_@Y=$04I%<CR^^<U+F\[ =!-NJ3<@'A1Z.7J='5?=GG3
P7OK^9QK0@1WR= SU%-("_BR8Z4560[1LGSPL9]K1*'[X)[3XX/HAME[XQM:=M'G!
P[38.,W(A)E3IY)/P@ VZ*Z>>764)6,X@)2.$ &>90I]^_T/Y^@D9$J3*5IDP-H71
P[QLU2:ONX%SCL2D1$*J7:0*+QR; 4>D)2?>5=S\NJCU@%'^YDC%89[Z+,?K!;SO=
P&1):?GB-797,I%/=K;PSZ=ST&IH/I&+=1711_#;$@SV@(-F4Y+WFGT++'I5^DC%+
PW.57%&#;?_OB@P>L,%$5FO[43G&R:TO4G7X79O7^"A^Z<@?DJAQ!5G/!U+F+!'6(
PC*D)G><M*KHRB]!( F92KL-1%@YSPNY?U+$NY[EB.6*<C'K$4,&Q@:"DB-'*9P*(
P +JH;4!D>0?16 ?_8G+CI'6'(HS\NT55*")4#+]1D-[@JA'@#AT<*=7QNS567S&:
PL)MF:7(6QZ)'LM%'Q+6@F"BDG6O1C\=B\)KKFPX?NHW3#$O)])BQDYK\YJ?N1Y [
P!\76AO[I0$T*8G\4!]4TL9G#&[I7_1+16(3MFX1NQ9L%" ?S_;?QV/'7FEIL4^C]
PHQ<6V(KO]UZ,M=GG+#UQJT>XO%(?HSND/\V8TD%9#8R#+17H,45_&.ACZ)=99#(J
P.:>11A,\UW9WY&'S\4WX2)DE8_Z2T",-H$01!?\0&*8JY0/8MBT&_D1IC"Z\R:NO
P@/^C?'HFHP1ZECBW\DG^M.IE-'9OMGN!"MHUCE0L ]"7!(R8I./M%.NO'L;XP](!
P<<JQ%/)BZT9&[0_)#:F4U-VD(^T-2 DMJ'D3-!#OO;_@7R]OD\V2E&T+*1XN@MUS
P)ITFS0I4:7@(-HZP9*FV&51L<9[.Z(>'NZ6T]U>XP@@8%C -#EZC!F/W? -[9H2D
P[LY0 <W-I'4?KCKAW![805JLLK2M+>0B@P=6&U:@WHM%VK?A Z_KPQ*BJ!I(NGXC
P59NI+.J(@/BL^"*F)]@!"S7T/YI)3)K\M4@TL7ZRQSS+0U9,#H)3FO<\?PXJDRV7
PL0Y"ZFU6M+1RQ[+B/ZTO(.-07@,B&>3OD(IKTO=&X0&QAROALFW@3*_ 8KT"A IV
P$R\!JQZ3E]H@" *1WG\3/P3,KK%1K^T5CLE5P&L\G8A/<I<7\$O;@JJ\9!VR.(_L
P8!8H<@)?!< ,80XR+4G1S?FHOQ./F?; D%;>!GD2Q''R#>JRZE3H&#S@ZPR5UX%+
P"L.FX)4.6\R+TQ@Q L,G+LFP!,+U7+0TNKSU)CQX>FBNX[8QN)9+V'15^](/8GF\
P@+^;7 FB]*7B9AOVPG [TJ:4$F%ZS]&Y=E(RPR:F?[0^I,U]R&.A P<CSNR,^6G>
P%BELOEN_E6\BZ^)- 0<6IPN**56^]UE]?N9%=@V#7GB6)]-J'*BEM6[*^2'@'H=S
P+ERE$?_F*0#7*\H#4BQ<66D:7;7* E/_?(!1;?B\E; 4C<"PH#A?-_1<-&8)3R+D
PRBLOV#5SY@4@EQP!]I74%\C^\K02;B8A.MCP]884GJAY[B;7(;=*\(B>Q(O=GS? 
PB.]C)J$AWYC?MM]&#Y51ZC:]"X7KJ0 I\#958PVLCP_*\5^PN]F?@<H"$REO/"Y>
PEK+,%6=>.$'43X!9!Z-Z8+,LM[0E9? U17%"&9A?C55+6W1 G$<8<A^1.^-Y.'25
P0#98*"/1-[[4P,,>%ZL=CHE=V1"!QE'=&8H/R;U$3A%8'MT6G]QITUW?/'WYR5N,
P--*W@K:8A4V*0TGG1V(]<A-=<4;EK;15J[1(,*2B>0T\W?]I?L=O!"S"=IL/]#O(
P! %P>U536" 3JLP\%KE5/( CSM)@72FJ\<T#+*!XX92A78V 6O^<5:%I\"P!G#YO
PU'"E]R(/$\#M&S-$ 4= 5JP1)T#=[KNO40)'6^GM(*)84#3DYY9K@:6Q<)U%?LEG
P/BJ)*-G/'%P='-5BLV85G$)MM0ZIN@QGN!EUE+,E]C]#,/Z((!2&^*&K.*RT(FF!
PZ-2ZEY $\255B2SP]Y\&%,._I3\0&@7,1:+NXKV(O!7!RT7*%T:T\H(WS'0<2:L,
P]=YY*=U4U[>:6EWD(P,>]D)B"0"]XG3HB<@#\NW,S+ [X?(4G,N,EBR5&U[B!C90
PM&1MRUEU*# DFR;P^Q> 98&6@ZL;9=I=,7IH_@V3T2.9R"1IM+9\=<E_2CPFIAJ,
PB5J/+6.L<WP"[=T)QN^9M2C@ <0OL+LA,\4L=RF@8SDKKM?4OI@LOF[JSNH<LFU.
P69'Z4'2Y5&^7]',T=K3\Y,]2L:VC TY_M*+ K1!GXR,?@X=30DCL NPO04AO7LZ$
PD.\E8@[=EX[@7^Y00L9F@1',0LMB<N[QLC?I(^V3\<KT/R_EI+I/!!42:Q-:%E9U
PEUO("!)$:;O@NW0!?N^W<\L=< 9V?L-_Z$>W;MB,N^,T/E.#I_<,EC%^_1\RWZ$[
P).SPH13)J0]_BKG<.$FVM)A:=FN 60M"JR+:[B2H:LO0!@\O_NW:FOGYC,W6A9:#
POF)<:S"GX5:D"P O,*M=3RL@#"=<#+E  [^8SS_E?" 6')^MR=,WCPWE0AIM5S!J
P6)("8FO6T?IQ$EFJO#1>"]@4AIR;P9G[$PEB6?HM-RU8XU>F 8T113NG76N D+&<
PEF%6Z%ZW;<H$=-$[EG[+&2P-=18U9E)A32<&<7@L=Q*Z(5P$'- 15*1K*T;M:0EO
PH::Q@K<P#8_,E!5X)LF67AX7PKA?#;0WDW^U"AL&C6/>:2\-)?M#GZEYT4G'\4]M
P^?DX$3TRB]3@PG9:D^]K=-=R)(505?TMM,F0&#2Q33C 0AS8!]6T,T]6,W%<N/4Y
PGF0A<EE<\8K %+XVM-=_^^LB&*1E@&DNOO)JDZ/)A:)6,<3R7U-L1__<6=2YP^^N
P915U9YM5;UF</4OG2@ E*>:O[\[B05#J/AC4&"RGW2T07S3T8:.UC.K_&R'7+&:7
P5DN*7N=I!/JH8#KPV1R+-I']3_LKY=*<QK7QS;,7@6G)Q+UP6S?M@;O?R/+M2>=J
PV,I:E'$-MG)=-+I&;W,P*+I27!=<;874_*[6HA=:$*$"VI:M$>^28)F#V$,P\K9]
P3J@0Y+,_%T5*%WXI9,]@@7%3C((%X.G,X#&2_[TMD$_ 5,$!U*U70\!>YQ1OAT10
P'-&+D0:JNJ<F6G8=HO9_ H 8TZY1N*Q;<(_%/$B14D11R[AYT$NWH4M6Z[_A;%DD
P%DY;EA;HB;J>W58[)#.Z=J(5:5-5_&1%R9GX#1_/$DME(=ZUPEPA-- (-;Y'8#X9
P86SQ<N8-T5&N=S86JM*5M6<1HB%97'NR;J?%(/^B-_3]*C#]Q'](#8!L,ETJ7"V'
P,B1G"P$!E,(,@J:U.+/YGW76)=P.(=)NP:GQ&[[8X3_C-4VJ+_=Y")I)HH\CSYA5
PRPXFW#,O+EZ2??H#S1)2U5^Q]A5&GQ=..^3&2$:% ^J8\<KOR<MT,0[!Q\-M"'U,
P@N<:5/6WMEEZ-X+3@E;I)^Q:0M]<$D&OIR 84H+YJS</]H+CM'PAMT!]U$T\MG;>
P"+I8N(6;!X#K".0 #CAI$-=#D[^)90 N"^,7[R8(!5/@O).\SB*B?!2Y[VIJJMYE
P,%/>)(QO"H;;JS;=!V&S=.\MJF9I_3FW\=QC>%"2L5 GT\W/:C3*3'P2RIAD2P@M
P#"%*W/]6QD],(4)>OY4@1[2=5YE$5-$N4 8F[O^B.H/>4.L\\[:)V)"1E]CKZ%:8
PTFU=^RT>)-WDU/%O0]Y*O;%%C(FCQ&%Y3^%9DM@V&QP^:NQ9P7YUM.A8YQKI87&S
PZA3ED2&.F7QNUXU')M?!ZQ3V<?Z_0^NMC%>@/K0MHSM=-75<1 F TTRTZ%ZY68$;
P$=6^GFRM*O"42%?#MK_K\I,P'B]7:<F1IW_IPTD@/N)RR4VP\5U:4,=:X#9S-]NM
P"N(WCYJ&+P,3 DRN)N='?D?]NZ=]\ .648$PY2R8<%4HO?W(+/%+!,<"H+ V;DS8
P8C,8EG)Y,16N*0NWB)>N\*G(]*#A*"\0^F.-2^_86D>&*)5A+KM+4X=*Y;6X=!C*
P$(KV?G><8W.HN^X4>O>"/,/]7@E-\_/!\TU!]H@5-L]Q^@Z)UF,9K4L P^$+1[9I
P:Z+7J8*3B7:R7#_X=P) 04>IK;%$4F.P^08\:/BGRTG;+N0ZLI5RL,SW(KP"-Q<$
PF8 :2$?HM+MDD*:X RJ93)8:TN+P?\_T[;BC92*5-6U#*FT<QL'<V8Z,1<;NA>AZ
P 'Q>@H5=&&K,0#M=HK&A!B717TW$.O/@B*HOD3)^<'-S%H890AT'5MHZ3%WT-'%:
P=K<ZI/X;/-E1!JRDGZL!+A[\A%1RA*B?/A4GM< U)O397#+M5*6 M2_H<]$!.]/8
P=TW _NLO'P]1K<4>F*K53YRZ1N@0<67^A3R8&L'6N=I?9 1E. B$2FB/>P:F[F4]
P;YT;6[#)1)&A^/<AH@2W0M"FB&RO _"M,.B/%5"_BEWW&UA8M'GBZ7%07LJYJJZ5
P'M\9Q_I5A5H39=6",<%GZX V+.O$\;3]FBCYG;*4*"AOO-O*;+DNNAF]T]W<,_*#
PZU\S,JW\[AU2U\<YRT X^1@[*NE165_2_4R:M/O<^T'<S9B8)(K?2XLBH-1UJ"B1
P'@X<W.^T[:#^K*3[=:#_,AB5)_/9Z.9&T4/3IH,@%@-$ZL'C_'F?$4V%9H-;@AOZ
P_0ME8/+"A6B/?1T_5KL#L]U3OGW_@!_1',<@TTMLS^-RD(;$B$#'#Z*[T)FKJ[:0
P.Z#2MG>OB,2H??._Z@$(YVSY?IY7PT_JGC:M)6VL"T6ZUB:%\A^#21( 79& LU"L
PBN(EE"%?'QL,8!+78QK#G!7;I[@J*(32P?1J"$=,C^H1Z%J)IV,Z>(G8S:,)ULR5
P#D[Y7#S&Y^'BIG"F'X/SNM*Y+?;@UL4QR,S9LH<-JA69+0W!X@N""?"*K]]_3(/(
P+0=(ZB&:_ D]NG$+)G1Y6WY*_336JQQ0<;P/M&)K\II]+27UC>A0_,0Y0U(H\_2&
PXN[QEYTBTW-^0+^.$A/%%&S,5^:[C RND=Y[YA*/QY@'W>^BT3?B8;+_NX9NNY+H
P'!108:,&T$E#Y/<7_-_YRPZVH3P5TA$,KY><11X0$ZJ4&W *"LMJ.ZU/KT31-N(Z
P;H6<J9 JXPS7]7JE*B*%2^N6:,M[[S>,5< _$Z[K2O_Q1K370)C91J$AV'C7G(='
PJ=9SYVHW^\!-[IQAK%#TP#V7225\=&@SZ/X78MIB@M<R>F)WRF6KWE#)5^PA>^.H
PL*$#_@_JJF36ML^+>BP&_MK!*O+_>[>[>L\CQX04OG2T";;'#&%@-(JP@2 R-U&H
PKP'( W/L9HY!DYB.MEPPB6VP2#3)=X.J)4>V/?\"\),7=*RA]%)AUQT'4:?L2/9Z
P6*XGNH91)P<E]XNS:Q'<LS6S0=?AB6OVE\JQUFDG<G5DF1:\:]YQ-8WC]1[>P,/V
P-]N!P$K0.<ANK.ZZ_DX -  V/MU7GO=#3"Q:-&U9J#P0)U6P\\*?$W*!!K#($4ND
P.%XS*BY"M?DJ&MK!_K5Z%:$P/E .^0+8'QXF)KF[ ?KM48_F'X*L'755NZ:Q_6JK
PCZ*Z M'V!@".MJ%!%'E'Z,YAJYX]$&N4<=)=EHH#(_W>,XM"/7%.^>^40:I_^X,M
P+[.\U.L#XB\3TN31/Y7"R_RTF&#'MGTW&.L3GZP9BQG):SK1>Q:L,(B[5,%%(G((
P]6H.,Q.VQ \7^X>GGQP>"BW,N2=$W==TFK#"I->G25J:R 'N;8"Q'2HG&<921Z 4
P2/9#]"$(Q=IRKP9="*MFR4# 0%';4P T _'4H;-^Z5-N-@GE6Q+R=)!YUMFY)"#N
PH":7V*Q1>;?!<$HD\#)NH1F8+\ /Y.^DN@=-AJ>,U_'R[,(I1YDRTGUZ'!\*PUHM
PX%CX:KS3Z.#3"+1L]YP+$U!3-Y,%$!+(NUL\"2#@TN:X0C\GK;<AMJ#DJ&"9:P,_
PMR!*4JQR^V2$<D\U7M%(,\;CBS[D$8GPONN4<C0>D1XWID><P;=F8:WZ/K>?F-X-
P*3!2?R;4PE2,\)JDAZY$JIF#?M+0-0J;U*.G(JKHSWWO]P\<?V'R&WHG2HME]>@1
P\-W_WV1=*=\F(E%<H 6:^:??^3W]P[92+FY\77ZZ\W@7WM/\\##ZC!"Q C_83\Y#
P*06S;:%[Y.9O OFY;#:.969E=HUPXF2M?C_GRY!=)Q4"+RZ;4RG10+HV#16UKZ"7
PR:?T:./A'_MC"X^48"F;)#99&>V\DE@L<Y"M%"@^L6+ S?C8T_%@;6_4'0@IX%D'
PADA<KJZ6((D"!T?>4G(CMYKOQ:3LF0YG8:=#@.O9ZQ3A[UR+18A'K;3!A>-N'@PW
P^!QU1!+L0/.E&O(?1Z0;@V'K!11WD3IU;9L9@  33+H36(2<$,K@]:CQ*%.!$PB_
PR&?O")3+7)LA%9BD#037[;,OR,U1H DBN*\6J#\-8.9;K'/ OFLW S;:$27H?\M6
PW>:IO$$=7Z*J.C#EU"J/]_NEM^C@PPRRL&A"N-). ^#OJ^2- Y+)7PR.QL,/R(W%
PRE>QJSJ,K&AA!W66DI"H;[2@>^2T(7XK;H2ZM!RB\N3_.2_IO\D%_0WB:BD#J4]B
PWN\M!2E2(+)&-]\1<HB^*#NU)K],!FIDB_TD']PXH_ !67C;[I.X9ZK'<D]XZ%E=
PS,=ADS!44.O-A6T1P@*6:ZR/<B(-K-@6_:JBQ% P6%IQ-X3P^>(\(,%C\5/-4[&T
P9)D"_QQ<GXCS& Q%^M'9WZ]%3W]ODUW_4IK2]\_R M86"A5!-;LNT,$6@R&T-^9P
PCDMGZPM</UKQ4.)MD67&7Y15M3179$+B^G$0/5E*(HLX#/YI,9KV6+ ]6SE9#OF)
P9D;2<>>&2\Q(G+=/X;[CN>W/FC7X_&6CJ C2+)*5<NSR1+%W&T)AH]]">4+@Y-7I
P?<]^2.2&K8TS#SEDE"DW3"UGU^V _^#=][3]?F>QS-)OIM -#DH0=5,+1#1P_@@R
P2H)QC)*V,-#NCMM$L5<00JNLCD> BFXF$L2S_ACD7C*$;Q \+$CYL8VXX)%=BL3D
P7$MEV,N738W@[86?8J>+VVM.^G_=('6 Y6HG%9+R"?I3+,HPT'@]U$VXBLH?Z=J3
P+[Z Q,>_9HU0UQ3$PZE PJZ3!(L5V;2)NWHUVY<O,H!1L]"47A\A9Z@2*;Q9^UJU
PR)C^G,Y/FWT<E#:L"TYD2^%' QIJZN,\-C+,,!$_%3)Z;!>#QS9H/H0#W,K4A' J
PV)B"RP$)2U+SN2R!0H0?2/2"IRCA"R&9RKZ (FY._=X(PV"T+=NT))_(/[DN:H==
PA%I_L4>6KQYR$J?3G67F9]\@T^"Q&\C[?GH-[&$-AI,7\LHHAPQN'XC^)0<C1J[O
PQUF$*\U])X#LH.A\K4C)1W*X:\4N3>O:/'\CV.61@3L:73M^V4C[\>G6CGQE<-C+
PK<E6UINM33LOR:X4K]JQ(8'6?G-]@!,J<\LX]*.O93DFPV><7;=Y@33QI61YXGJ9
P3"OB6]#S(3HRT"X)HDYQ3\PML<Z5#L'BD67/\ $^1+UQFT&T-"YY*=4VZ"2/[X$'
PT( L!H4$+U%<P=G/W3<3RR[Y 52617*YSU7R0*LCK*NK=X3AS:;8.;U_%9QU][-Y
PSN0G)\]6!?<U+4C_?R )XF'E7T!<(NT2BXN.F^[N3HT14 B.\F-9BW,8U=]RSK.%
P:C#:_T'N%?Q!QKE@%HF.&)O9^$6QR%)".C8E7(2[S%JL.V4MK&\6;NHO)5TH(,.%
P&8:^LJJB'J<QQEK;21&S1OUFOB:C4-7RVYD-Z$6_R%\8]J4$ZTL)W3\3[HPVW"%1
P&!QD-)&]MG!-)L5BAKA)@+^,1I()_^L?;?0*?"7=*JN6XR&U/9RB(^&'AI[9^R:;
P5^OI%N;X[N+X03DBQ:O+-#.4?VI-._APJKO"E5O%^:]V%GQJKU3I=WT2T;N4F$F=
PVS^?@O8LTM_:-R;,,7$Z!Z8DBQ+5*']TV\M3)O)6'<-HG <$?7;&6A.,"I*)GC[?
P_=-6 0FJ+K3P;S'=-]W0% ]CE$=:-O< IZ'#Z#2_\^<=2MMM/YC=T1Q:1G8%KBN-
PY9Q%3F]<OI]E;E:O]U2]^<E ++EZ*!+]*&A="WN^5$@2Y.J1S?X.T7F]HXY9F6<S
P)SR'SS:;OW35MO!5MQ?.#1+Z.1\/T!?&&30#PLSW5+\<6]' =/5)58;XCD3CIV 8
P5*KGN&FG6=T$22 OZ83)=A@0!Z*U.OGN$;=P*V31N'[DIW<\PV:^5+%PF*61G$VO
PK[MJ8;*< =<^.[.NN.+@5AC:FBBYET+TZ99'0YGK9YQJYR,Z3W0O7%@F6[4AI+^T
P[QI4[Y;>E=L3JH2P[8XT\">M$-QQW/ A:WF%>$JK>.\,8F!\+CM9<QYH^[.GO9/J
P\H!N:SH"=4 NL[@H2_ \CATIQAKHA_U=WR<T]5!$J!<OHR&8S5H' +1"AK^WYB>W
P,CK#_,8H!FB[H2\RJZ;&1J2()/R)"SH ^43N L$NLAC%?%6S'(ZXK]0T>>0V_]<H
P9JS.6C&O#TJV$]NOF#=K:]!XI< 8S6JWYM1=D=8M[HXB;G8& "C<EY?_FW.P[PW(
P?P]0L&[U:$O4A)YQW$?@W"W)Y@$_>P(Q?Z>*XQ\YUP!NTH,>JWI==#0A8-Z<"-U[
P':.BXLSIIPW-*#6DAI&<^CU$V1Q=XP WJ&?3^67I?<*6@W3R(%WLC&Q!=<J%24B!
P"KY=WE\B_J1_3LSB2TF@/T7URGG_5-H3%"'ZB_N;F.B4+P>ZS?[P2XN,6&)7U_KS
P%Z03^3PY2Z(B@'[C>"^;BWV.@# .$JG T%N&V>:3Z$_7[#<":U]!,8:SK6*?OMB-
PHA0]1$OBCQ/!(KS3LT@6&!9I7:SK0*BUS&O[^!D<2#1W);)LI2]M'/^7>2;<0\%)
P63AZ:[?Q]&F]1ED4X_!&]#]X0LGU_A20D[TG6?P"1/V4=7QZ"^$$7^ ?,(QT>-E>
PCN!/>W5<S$QN:C1,'^Z9"YIOB ;08<&=+SJI-J 5?=OSS8EA#';E^TGDM;BQK.IQ
PE2E<+RY-F,O5HB.6K Z'$1!"@W+0M%,]U[_WVHB._^H)\B$VI97'B*J V8#TF,IC
P(_8JJ5^Y>TXBE.5>4!K;K+/ATF#6RZ>DQ.I(AI$F[(=VON$7?TT,3$1!J5.C "%,
P;@.A;0&7(!&\/N=Z#W5_5%'"77HK]=[YV"$R;?E<W0JZ$U(8;A98@^)*J[.WY$5U
P2(O40S]FM54/BFY52@:N&_/3[C<1.)L4/"XTN$7ASB)HK!^]XN\\+/5M\QM (779
P81EQ&LG29X,:<ER'=4>0:9Y0S:7B/'M%X%G"_1P"^=G/;PDHP8F6[GW13G/R*<DI
PX>U4$PZ6XTV>:&H60N*@!;M6*8%"9:C*^W[L)C?'3'N'_HI5C&0K<3](?35HS'E&
P*]1CX"V><9CG9=7/_B]F_T]_W!7^PK<8%3NE/O/*R!L8@@HAHEML44>,AIKV*S0R
P%T-M-<M7K]GU7UMT59.F!#7V4XDXTYL:*V#@_.7$RW1.' 'U2Z)N',"^2H'F[1OR
PD/<IVH!58AX](SXXU?NT0E5=BM;:!6ICY)XPU#F]$,*N><0/+>&OR+)+XK-*T9TY
PX%<0F. $BV[D82:9S]X!5*W!9Y.:F?Y_WI1GW#2OAVG,G3!^=-,TEZL17ADAG1><
P=-D:\>R_X[C$7JI6!>^7Y- EK.H<B ^)ER]LP>J/_VG< 8Y]7>ZXEG#O,55&D/TH
P41KZ3.@/%,"TU@%\_JCM"KRPHJ-NM1K_',;P*;_:>V6=2%"OSY^K!1+&0:^')>@G
PVLG$SGYFZ%U@5;G^R=HVR#D:BC:=":$OA6-?=UEB,HWX0IGH_KJ1QBFP@A5]=FV)
P)YVMSF(R84?.1^ 'S4/3AVY?/[O&[+TVPOZO5L&8"V"H*+P!VEE+9 DUO F_]B0%
P]N#$.!5]MJ).U>UEC2@Y+ID%<R)!)/M4*0RB<O4+I_"(K5SU(*8VW!.^09,_#Z@M
P3R W'MPYC!.4KR4C!@\EMXM:M]OZ:4IGMO>!RMT4'T%9UV"AHUQILJZ;K.'Q6"S 
P18#W -WT 2.D'B+%9^I?N[./_MXQ#0_<7KC?B/MD;39H#332;V.U2^[;V 2P'JQ/
P)R'A?696LSMF7Z.FIF9 L+)-J!@+8*6!8XX6#CLV'/6L T:.T9$X3 UW@5#[*#/H
PCJ,&&'J5TM31"#/ _;%:+J-I!"6710_&7R_QS(L6$K,G8.\XQUI%&AK[+_E*G T9
P/[61LX+T]HV#212%A5R!$VE>.Q6(H>*/RA#B14AR9"&*6C6+B(.W':T$DU#O21C5
P(2&"$IH+*KK"PAM@-LHZ$PIZI1?)XKW=EEO:87*5;'IF897-.42]U8/H"<>5-Y =
P%L[Q_>H6$]OI_8</U"[^^#Y4)E L:O*-S4:.WS]5!IAK$<(4B6EEL6WF):RW#D5\
P# L%U1B%\V,#_-YIQ.A-?<T[^*VK9)NK;D(%[T!VTX49._"C$?ZW%F%,%YJI([T$
PZ6&+.'IM&@^^FT$RF;=9VGF!^[6#[4CI7C@T+:Z-OBBME+$1-83BL20.K%-C:]-P
PU,S5J&D$T-.4B0((S";"HHB)8E8[JL?)(T:E*%6'[N0NZ*91>YW+ZHL"(XP"=!$F
P]NT'_!<YF'MB^1*H:X<IA\$9X1X6</$*?R'^F51! JP%U.ULZE!],?E&_\-/JQ\%
P&Q/()GGXG\HQ.8J#';.[_+6M5*;EL6P^FWH*5;/FW*??B6[14-00:3 >?=,9B&4,
P5=6?Y+XHV$LQYXE4]\$79P/S6 L('FUY<EU(9+("^"K!OI6<-!])0((B]>HM'V[2
P&(D=!]WS39.#7<3S^>5,J@?(1ET_I$(I/\@Z*4FAX'#0EW5?,;H)!@UF,#H4%<<"
PL$X<#1! RK8\P))3E(Q:1/'?8S%N6^%CY&WL'D,L?!,RLUV)Y"_?+O$A'A#JI7*'
PF):^#2F4$E#.9V]SNB)\UU=#/#7U&S$F#74Q;4*AJA^CYDS+1D-%-8DZYO+;Z#(3
P?'*DIA8].+8*<^GAK[_;WQS9*E?9=\".4<8)?0JM&<P^H%X1#RY2B^V^#9)9?!=F
PS0%9)^+Z4K_P]PPC'P,E[R:#\D!?2T=!Q4/$IPY\'41042L:MEFHRO6!\^#(HO4^
PD+'8-0K^VA"5L582^2P]O6UJE ,THYSV:N>,ANK:4E&S!!RG^<E.@;8P;A&7K))[
P%A&TUM D:(I7+Y_/A M:^@UM2]_3JWAH 0& !_G,+1X&_$7]%G74V.L];H'N9_\"
PUV[<K#OO("A(>^'T7O#YO=<6/K<&',%TOPJM>7C-ZNYKB^R!7L5_1]J&I<\34$:8
P*$34C">4M28$'4,=G C<5-4XA8#T@,A4/WU]ZU!Q4,]V'7Y+%667NP%!4,RMS67J
P]XU9I7@8%"H/X'Y-Q[<2JY=6_)1?Y:'Y%Q/5!E+CEW5H/ABX>>9 OHD^BM1]VEUD
PKB W#<GM;.\R8/7^,NL$K'BG5\7#2O(-6MLW"S&7TD70J7H\Q)IP&SBYL#-#S02\
PQ;J:WL@&/+?W1=Y*]1_TVJGRASD\=E6I$Y3>N,=B(W3O3*QL7#MT"0P+CO6?U:IT
PJ*X<L0Z-_<<(4XE^#LRLI8<W7P?["E#1_#CY7IY:G"KI^:(_3Q$DUKF^%S+S )$C
P3>B=1_?%8IMX:(#C=0;QU]4X5RD8V3K!0G!SVA#0&<>"%FI@:@X-WAD0Q( W&-#Y
P-6)7LOTN-)8Y9)H:UNI $Z?@C]F^GD;0%7ZH198WC@N.,(3GG26 A()I/A/?D>C$
P9O&;/.NZ+Q 0HI;J2-=)"V*+FW#P[2S(; =R=EB(K=31K>+!PH3MS-M,@F\N"CH!
P24:V0MUC9RRZ@*M_HYJ%D*3:M6(&+#D2%C)WO=0R @I9GXIP4^M=0C[+2E!E.#/ 
PA-SQ\@%&U*4),7!4O$AGI$M'V: B8K;-\W,2&@:Y!&?SX6*>>"-AV@LS?J::<^>P
P-QY+LK1@0A'!K/E'9)SG$%2)#J Y0%3P:+7(QR@T!<;J+XL,*CONRE-BOL[>OGS<
P<+:TEF?T?*VH@];A0%&AR^1VUG\58<VHD309L(9XNAMQ++U-078EX4($ .I]+C@>
P,0GW/AB(*$L7F7_&;I+%6_\:&O'@,#AJ',7&9+:V?ZP#F/*/%BGXW@N]D.:^M0F$
PCD;UG<O_IN\NPG0 V>R?:RBN.5L!DF!/*N:F7NI*"R>]8%S'R!P1PP@V^'#E:(X7
PS:X_-EM;]Z2U[.8F7T5R22#"+N'3-$,4!^"17.CMYC5C?+IX">0\2_V1824WK:DT
POO(WM\7Y+%0V(+)-!7"3 ['4H-H&Q4?\S12)QLV6>[4UYFWT@<3VDH9ND""=QOEL
PK]K^<5W7$-^L6S$<H_QOD O/R-ZIAC>!07=Z]LU<>&R(YG?<COE0;>?(QS/E.19V
PQS=)X)B$BI47E4>^U6H]R$SA92'^(6$,;*.VT7A#OF;8!='*LIJ!-A3'&(985TD 
PY0DC6".D%<PT:BB%E^),E)!NJ%; !N1B9A$U1A;RXQ] ;C;U(!\VK;9]G$R_U0:1
P8+YTD2N(V9-?RQ54IH'%G0T+8)N&<]A^VOG8IY2,']?E4!GWR_J@C)<\@I>8_36+
P78;BCA:T;3)OIV#?$NL&>"(VETU72=5AE)5]N7%IC<X< *7X_0P9:7DPL&)7@])X
P'4=XA:?/WJL'"4 DX4@2[3I)J00-\<2Q]]APQYNXGIM34>_KI<VGI#U,8F,H'YHC
PWA> #2 L0-N1SGIR"U(I7)\Y=-DBNXPON@P^RF7K]N]\>)HMUP753_B=0OS<2#/V
P.@<9^$)**#[7VGB(,-K.?X4XQQ\8=XWPL<NT!C_F,1XO'M+UD+&*CWCF\$$(M"Q*
P-.]?! XN5E5_)F7]@,>P7O54J3=KBRK:^V+!@[9-[:%1\?RQDK$Y[R7K?21'PE?R
P0QSP3+QDN\]M1V^8(X3HJTMB!FA'8DUA)P7M;8+UO;>8OA/L68-\0\ /6+%I3J&X
PG+H*[]U[8,Q>[/=2'RK@$NURGCS+00'X<DKVL\*J<47[#+H&Z/A$!ORQX7J&8/1[
P\__D0 &\I16\,M$G&:F3)?29)CF'(K)"T?T+@<P?$1*T\[Q+$Q#.+AD;H7RTJ&KW
P9&&H5^FW#[M3OH.I<+R7%#OMG306>S6!(?:L@D+\FYF.4JX".U A>O]O3P!'^E8V
P_^SL^\BI$GMG( $[5%3/ P5=OCG]!-2'MW7G+0!_?JZ(ZTF)942LN=V#[P>"NRTD
P->.;>9&6-@Y5MMBM>A#G;T0,(L+:\!_6 D?AQCB81I3;TQ<7)QXJV<^PX<;YWF\>
P=Y,$6EOT4@1D[>8'[GD%BW[L]S'75RYJXS_! ?S:FD?'+P0[4O3+YG.<)+!8ZS<M
P4%^L&"<C:=<%QM[]4#1"W(*3H-XA++X3=MW,7\$VSZLG8PF#B1"$5@*F5ID*P]&@
PO?^-E;E-6I?8!TA4]@P4SUR'\]#:H*C)6!PJC<"+L!&'K#"!P/]':@.V_\ID,GA4
P2<#ZT<+:'U5C#E+YQ#]GDIX27O1E1K*_Z25FXC^W4:&A.@\M?\^*'-6,N70W!)(Q
P]3ET_AH27-NAD'*#ZE?J?#XPC!#CHFC#>9GO2TNIUZ6 )+=JZ\[GE$&HS $G.7?[
P3(TMX]MKMA-RXVP56V4).#- [QN/;#';$JS9N4V$08;.SHUJS+B6.9<^\)U,OG\>
PF&,0/J<;3F=6Z?TY/[LT<^KL4ZU?.^QP?9K*^^B?_M'$?:*B<;IRW3""GPJ[WVL 
PUJ<@Z!A\V>  7L_$))\24E.3:OKNQ5T_M$R0POK=G[I?VM[BYWPW,.$5%B=<AS(@
P$_&G)?S2CFZ:/GK7];&.N.&W:QGF8F&-Q=D.$E"-[7V9+_T6^ZA.6X3F-P/HV9:5
P+YD:?PT?.[+A=F>Z)DS2EL2=UW8L%2H>Q/<$-%@DL !:$!1-05(\6]J\WK=80**!
PWQT8KX>HQK3@DH=YH^3R3@XJP]K40YA5$.O)A6%)R#F1N(J;,+_\3 J8/7_DH*BC
PJ4;*@8*JAM->K2> J4LX&^&44&]H.TK39-6(*;6TCQP$,SKWQ;,]1%X=3'GHN29A
P']S"6C(SC,Q_!H'\IBF>CJ$+7P[&,UKZ ;7%=FI?W[LT^]=2)VIIKTBGBF>^&KD:
P.LK+]AA6:OB&:HZ-NXY1?5:GWPW^+C0Y-F)GM!=21._8[I'*@PP9>6<K+FNJL?I=
P%$K4>2O[(_?#PE&R%[MOUKA[\Y6)S<:,94CY.QQZ &K:!M@*=.;IC=DICDP><?11
PDH#$[.+;.=/]*JF1 ZRW>RWQEY?1Y];8R1RJ_4])X-!0RO_2Z?1Q3G9?25VE/7X_
P"<7!B@Y'WL'2_<@TZ[/GNOI0S4<PW, (M*5SP4_7_38,JWJ(J<2'-'4),E-<L[ZB
P$<YIR0D4+?,6E*C?O:9[1;LPX?PLB710V]@C9YOC+9F*DLB94/ZQE,8Y'B)/+;U,
PGV<0[>,*W#QF9-OK_SQ$YL5$9"N!PY"0!B_!Q]=1>E3 *NL-\1^ELY?!I?-?\1=V
PT[XT-4)+6)E-H)-.G%:A)SFLCC4 6_VV'F (H+[8)$$&3EE!E[7I^]"^PYTYUTRC
P^Q-O'ATI!LZN@:,M1#9&M=]VH)^QK0<=KYO/0ED1HM*G)'LI.8<=(U#_S_^8M^7Z
PKUCP/"KF$@:(]HO+7;IW\)7G>^MO??6?S.- X2J=<>Q3$!^(Q(5T:4T-\W-2DK_H
P9Y\CWMC'Y?G'9H$.4@NI!B1>]7+2K'!KP_@+.W5J\Y(2(&#0A*\048F!=I,J"#+H
PE+N1G^XF;\A/4AR> U4O^Y]T)%(K@O!5M='6_7(UB[KDR)*NH.#R*[CG+B=\^W'&
P:I]D&&'O9>EJIJ/8(>^6B%GLQG/'GOQK35<)_9V;<*RLK\BE\+/%^9 (9&.@GT[/
P0_OOX">?,#_S_%:TN+M2/.8WW?USO;Y@43'V!'&XGI5A>S-U8D-6"ULE971RS!U4
PZ_(6.3.*CRN<@13"Z[1W,7J&*W"6V2'*%U\Z$ 5?0)X1Z^KO>5$6VB.99U!)EZ/*
P,9+E\<'C#>[Z.+;T9_&@7W#9!^V'7ES.!W$< 6E[=MM%%B+J=I;86!]\VG9*2S2V
P!HI4H]8Y?[_=,*-]$<I"/;>T<Q^K4>+3489W"@YNT]U]A%9>->2_$(*OD^BKHURN
PO9H/=1!X1Q:WGOP4<T(,N,;3N_@G M6E$D;5$U;H[MA/%Y"_NFJ/O7110ANU=_\_
P&'7V#QIZ(J("%]EV-GPLRHBR0<]<N6K13Z=8?RB^R/)ZU#NM@8@))QPXH;K(K'1*
PN#JMV'7W/9M"()O7;VB2ND?I/;Y<F8L/<H?"_AG*96 DO=#^$I[;*0T?^Y19C/*P
P78)+^5(2QV+U3NZ34>".A^1'M,<[)#"G3]C-8H]U;BEG%2TVQW$P#MG=KO['K:1I
PJY8]W]:N !/EF4"W8&\X:W,0IA9TU=]_MGD<?AL%)TG6C1W;V\'B*!^PM=2V4D(4
PRRV(;WG6[(+^M" $9"E609GX<A[!JV(939SRGS0=W$0%2+!7@OPN 4F$I>06:@&?
P G?>[3.M!F]JH4 ;[\Q8\[J_VLT<O954'^U- C9Y06_@=T-\W@,@-YGMK5RJ8&DI
PI\UP=FU7AE4PWJL"_QPQ5X)IY3<)T"4ON9N\BW3G?C9[YQE7BKZ\7YVDQ[*[:=3.
P\W4LKX". =*R]B&I/@28K-E4L?*Q(6+>S*"M-9 I0$#%KYC0$T C*058,$$$,)0+
PLUTWU8,>R5F<S)HT$^(B>J3IW[62,SD-$EA28'<9T_/G+HX!ZOQQ1Z?B&1H*'L;G
PT'QP'=@M54NQ#W0L18U9A5 0-U=RT>49?ABKT^GI]ERC' ;X2$+)Z#U7S4D/3)H$
P'MU2(:NJY]SM:S]X?T_:/>LK8I8%SK6U"8UI7:?UW&HCG!&^NB^E-50:>SW>41\C
P-J[?*(X5%E?_FOIME!YVO'4REFH2@"D71=D)M:48@I0'_KM/<T'Q1GZ1Q*+%XQ!8
P^C<<Z*78D=E:O F]35B]GTM#,0E$0R;6.<V5GJY)VG/_;/?39@HFYKA*M<7\I%.2
P&3;\N!_(DF'HX7_;O'\  4!'\*A1!LNC@RG" Y6:?NV'/,*?8!:$(CAW#S?@'NW]
P;W?%:L9/V.L#^WRD19YLD@1\?)ENASBD1.'LBL)/T_->]HWD-$P"@<I?H;C]N$)*
PFA/LEW5TR3F*D.*LS"QYN^@ZKN2V U45>4(K7/_6'VZN-)>?'FW_ZKI0;GN><,N,
PNWMGH9"O,_!1G116\6.&.)S)ALE57(W!O9_+G4#"9D@FFV2+LZI['!<56;KW(PB>
P[4XRJI/>V8UUH%^0$7WK<6:Z:T9T1RGCATQ-R G:$ E$SNO14>NA6"PG;K'0,.-0
PWH4K>$53\BTXG!R+D-6E7H\;AC1'=Y&OMPWX L1B_A2))#.'['D*SI _P)V!:57D
PMF %BT$M@JQCBC[^N)P0J'MYDS%?:I5!XK:>FI=6\[\*H8A9"A=([ 4CPZW157Z)
P[(A"F#; [L8=6S-].P&XO*VTN726>;D9 >06X-J,GJ$W'\$Z3$ NR#9,B$K\;$^2
PC*08*2]QGI:E!+6XVMJV+L+U'37GSK0HT]D=!^7DL[ZO:QLHIWO>9WI>7F)[0RE6
P7KON4Q24_&_MZ5K#!IVEK>,F5E:3HP/AI@RKLQ+#KO04IHRZI/HI2"9@]5<'&VNR
PF$J;P3*Z&9T>'$]#FQ;&C#4?<]%XM[@PI8U4#[(*OA64[9>SKD[23R<YEG!="%4@
P.'VTR?A\K5;C/5^^ T[>;[8 V)U!ZLG;PS(]1@,S7C.0&_F;LLBN;0**4:ZOXL*:
P7+2,!+.56FJP5WHAMB*09%RAB^].I>2/3 ,I3@+7805G?%]XJZT=_ZT,@0[T 'UA
PX"M1KL5,M!1+ 24((?;_V%PA>8V#0:.L($HPI1(\U6GQ)GZX-LB.H\\]%2UA#.U$
PX%SDSJ,8U%W8:V#(N(N&_269JX;?F3@?$-3O1Q2!"B'VRN!Q1VK#?'H8%TF/YK7O
PSK^Q'D1M\E+?DA^=8O!\$Z!N(WB0- ;3-]0M%=N\NVM>KYI:N@3&6@2PE?L6Q&@[
P24ZNOOQC"?+F]LJ><%I*3_ KE7!'S:K&SRJ)9N\E55UH[8]]7^M%E(3EA[DHKU<P
PM!';U_9\ZO1ZKQ>DA7<06 40.;\.UG BY:@ ^$=RXY-17+N=36V#>KVYUQ)/1^ZF
PIK:*G:>HV7&_DJ\A]RSR'\\O*_M2!IA:;NV>-%[CAO+@MSD%^C"%QE=P,56%'\W7
PX??S+IM]$(:<\0.N@2?ZU.6E_AKL$KK31(.8RT3/'.&LQ!S9T^%+-J*;Z$9KF)VN
P]R.-6@U&)EG WY8PIR3YL%^'YZAYFYU7C5/'N)F([12%8>7F=%H!B VRTN?*D]4P
P2-9'>KR^WLL8&J0'I5U.&#AA2T7 \TK@OKA]!LUY!4F8(*HXE%8L^(=:MFWBL4DP
PF"%TZX^XRD%2>8+<3]&"[)#S2R7S3/I,;XV)!P&U@:0$4FO\S]SH_OSUF-F10(#D
P[ST^KK D=S#\XU^^V&V**:5?GDIEX722EJ%)T*"B%BP* I$UV M3AZ$FP6/[")= 
PR$QLC?Z.S,@'\.>%:GS5=-MKQ90Q=J.;>)<$GW+W;@?LDLGP>8NNKE$/02GW^ M/
P,O6:72AT/)?S8RTC.#&5R<=$[-WXW&AQMS(Q"9H!:4^*L4'XO1H) <P)%S9->%29
PVYY=NETX3R!DDE:,PNS->U_QBMSM!;M_C#R_R6"^=O[\G+H-[00/MQ7;N9!C4DS=
PFU['/ 1X(;;]=]3;NE9X9J$4EF.O+/L+4&(B?:"98*R6O'!1*IV.X^>,+]&;J%U<
P:,7P4.PR6H'K8'?=VT+R!7GO=+/YC)W4.B6[A':YJR?&4R?\OI46 ^\$GJ-:QY=R
PAU4L=H^)&'VO_P_/?UIBH@"ZSU]C&?I;MW&_1P:\,>D0S=9<7N?T-CL0G'H*B+SV
PX;SV]%45)1E0UY6%XSD/*5Y6=R2[\H#2P@_/; 0%2PMI1N*\B_K LPAYF3F73=$L
P$/@(V.*;J5CX[ EP[W/T'2Q[#)]W@4VR1L7CB'"JF:-AZ!H)^Z=(C)MY,ZD!PQTC
PV*.?DDAYHJL]$*E<H,.-J9:T*I7+P.Z]94CDD1'CF-3N 9;\.5HD@M%!1BS*.H,3
PXY@ (B$>&\]/%$$%=@;5/E;1/9)!3I=G(5=<9LB=KPJH7'! K-1K[&"B"-W7YIIC
P3'\-6K0FN_U)%5%43)QYTIOA4@ J.VH8]P83.!!"6&W1X;@4FE_;O#U+RX_%)=TX
PKRIK26W=ASB?T\B9F'A:&MO7824&+"2&T'1*1<- O3U31W\=YLL"IK*%P-O.(7[Y
PA9+(@QU427_0;RR%)*E^NS8P1OO\,IU;LB3!=7])+P%U]?/L]5X<DR_W@*9EI+*+
P8F%')5$9=6\*R99:'C>IY<OP/A=-.E5Z8WM\;[6TZ>0;_X#L2'.) CL8YU;L%?6D
POYA'2[9&4'OV<6_L)&&7E+T;"7X[VZ]"2\_J 1K[7+C DA3L8743P0(XKO+2M L7
PY>F*]JZ0GM(J%/#=JXO ]/*39^O2\(P$.1SQ[D"JPXGX'5TZK6\BAP,D)U"GH+KC
P7,;' ,,;Y[J]BTG?=DLY4\0[?Z'^I$P+]%V*9=L)+3Z05K1D-M207DW%RMQHO+ J
P?9(H;RXN0 QE#(-#W6&1#E_1_3_X\5KG9T &I6B5XQ BH[8Y0L^# 4+ T7&0H0C#
P\RTP<Q3SFYLL*=:&U0PL#N_D=%$,YGVQ$9Q,@G#TI>,"/CQL@P+56/-UYWR'/SYH
P[_H5V#;YWRQ>9')[:0A #RT1NA8;N6AF\2G:T[ZGU7U 00BT,O+_>[GY<VPZ_P%Y
P(=/3&8AM1_NI!_I&G!X.D(1;]^DE5_/M&*&1R0B^2_,6+R!D .I\=[.S,@0 E$;^
P?X9PU%S!@XQRD4+A!XHG7X6ASOZG \DH4<C0-<-2&B W'(ZT-'?,3R;XO&!D7IG[
PS*KJS@$=5@*[2JF'JJ5C2D0KM^[;>$,E+F)Y-!EGY-$->V,XO&\*<P+_'2HQD(U-
P#A'42.--Z44AO5.I)<>X"2ZC7"57F=H3VB6>ZK([*W/=KA27)M>:Z*5.MMJ#FNXS
P(\WCC<LR/9"N71O4FB1.&75[T=8B.,,5^LVM1/WL]&:IA$:>I+:!2[<M^G"!\POT
PSFF"Q^-#%*"6RL5/J\W91X"V"3&@0&_EIYK#QOXHVGD[">8^?[X5?U\#UW:2AHOP
P%6339.:>@6LVMG6W-JI4(9O8XMIQFT3+:KA?J3ZP[#W#L"3E!RI1Z.,5^Y:^Z!2_
P&YE.4[4\&GEHE4-.@LE2]8(I_8=>M>V!@=+]CM,.2?Q(K.9 \P9YAI"B4CS9F5WY
PKUZ0@C1]H;2KAUU-;(]B$"HH2>+<.K5N0;G\8+A<*9PC]ES:;[D8X7+^4)3#EO ^
P1K<GYMKM_QK;7PV4L1:".$6CE@)"Y\&?.9XA'+]R%;!9EP4=%K=&ME\,"SCFK$7,
P-*W2S@SQP8K#"@6Z&?B9C#%EC*U='F)^B_$4GE# 5A$95 HJ+6RAR,7=\N6Z)P=T
PS1WY'86(ZCE_4+)?KQ"X9P&<4553UL1,/##;B3=ZW8H;<H^T_8*?QN*\]?CT:YB2
PF&+MD60IV.(IQ::Q7-.7J AXP-[55U.4A,]WKXD073RY2 :2SF3"44=RZ1A%'/D+
P$]?O^Q:,]_=927I0..)BE6 :W6^*=E(T8/J>JK4+;E'MS'<'KX_,5SWW(YX9CO'-
PJZEQP%QS+&^TR;\2>L7UY*U)'Y E[4RI<1'4'I4MU&\DWW,3WM5\Z!WD#FUR-4DE
P:<]#%";QZOFLVEP"M;M[K%'.TG+-$(?)4-#G5F4F<:16G*U8>6<[=B%H$=K-2\?.
PSEJ@5G2:--6D(@+G^R:Q4(P"1R_$<G9YA?K?K'1U\&@(L*?7K<%(R&_9_>^OM")@
P*#-OA M%RE6GHPHCOL8/).ME\4*+:#"OJ3*3X+>Y&">5[)Z(=&CG/\ATJ"UAW_-%
P#6]U2:CODCERHQ_*A2%;KVW7\:]9:K8=D1NY'A+[VT:VU0]D,#G6'7/R','V&6P8
PWP/L:4H)T)L(_G+,$7:#@=]"2NYP+R>0.OZ'BPMJ$28(\D8HI=?]F60I#8.*C'.]
P@CN\7 E#&^%4FU=@ZQ[-<\U@V$T\L$*VZ3418FC!P$L+EI&50R+"==:W"@X,DYB[
P.B:(IAWBZ)Z2&S-M.<Q4B6XHR3(B=42RV&3U1UU+&AMZ;]I-;]4_I];T&)(1G%P3
PYW;=^T;$L9:E2*;>A74-[EQ0'KAT&N^K0?CKWLA?IT,(X^[8Q+S5>FBEX)9%L4PN
P/4W[-EX>CRM)H#A&(DD7\,80/"=?:>L")42%BHV+&TGISG,8!R*65#KS2NNDZV3.
PFS\>RJ5$*H#WVH73R;>^-40>O#0M\6%5?::I_%3-YKGA&:3]HZ^\Y$B7O].A[-LS
P\4ZL1XF5'^RW[@(U -Z>W?PT4$UB@5ITZW([O=A_UG8$DBZ$.:?,$8V'>=@8TJ<4
P!15"^O_?>[(F28_['1D1*S@\A,K-M[S16"D8KVG2CHFW(RX:"7"&7(-O#9(^I&9C
PNBL@Z0"J!6;-7Z'I%?R=JC6%X<1_@C(W%YS5!P*B]_4:@WYDK .0UL'@20R30=K1
P_/;*U;,06-B,0_'*,6;%F.#U!:,W*9&BN3)@2W _0U#75")<J$;RKUDU[U9OK_HA
P "WH-B=XW%D@4IAG=[Q8#1L(L!D9Y8RPS/2FA!2R&&Y,/'8#XP>/J]NS%B'!84O6
PL#%$XHJH?<$>.ZD1:.),P5/#$SWH_V@I>B] '@2FV;FZ%=V<.-F$M(6CW TH)8 F
PLH()*V*!Z@-\UJOMDFXL]06=:%2C$[99R^TKT[&JC*V7[59UR+G*-GVU<-CN/;EK
P!&,!6H;I&\RW,&I7>ZM/!:VS([$*YVDN-N21_(G'0=P>NL IWI8+2!4JF_'@=/X1
P].90*E1I\R372BBL"D7S?Y1Z3F8!_'XWW<D@^XZK4&:#DTI9SZ+F-YOCT#[.YT&,
P](L[$%\1!^:63$'EJB7?^H<(X =+]-I%9B$EHB!>! [:I\9<^PKSN>*C[G2809$J
PF??,<)_,/Q,%_"&U0G7CIEA 7,4!\<Y!?V_[12I;]RP5<:@"7XJA7I@I8SO6YU.%
P-J&8F:!?J%_3F\I4L8#]*0026/<0XF&BSV&?L)199"F=0,DP3O4N"W]K<>OQ$<MS
PA0A#E)GW8-7Y&KDRP_SM_DM7)4?JOCA3#>:]O4)5YXW<PE:%",I@I)+A$],$)OZW
PS6Q_2RCZ# ([*[**#"?A 8HQ$,Q%,EZ:+=?0JNGC?-/JFIUWA^WI8>H=)RC^L]&6
P"CAH!+<]=.5U_PR&;G7K.2(:,X'G8BL1%OD^>$%JTD?+1!)1N8+E(V];[1;C0AV<
P]3O8))UIKL,BU!U=4J%#TU",<NBH.:)7%,[PN/[,-R0\OH-L"EC[2:,/\OML5RWW
P;3+GI3RBW,I%?1_ *MKO;H!:1X#.%$GNPP8Q4' :.1\#S52+9M,5BS88#WT/.GGU
P+])E97X.#:935BL%](3U(,8XS8$^=+#3712Y9>\=]GG4!^-]VZRS0H%S6E>EP1T<
PFL+,(725,4Q[?M'M1I-Y5\TU,-9W@G,=J>."H#NCFZ/(_"[40B&4[/O'.<$MJ!F6
P S]"R44%NVS27EYG/_^BE5ZE,E(L,-_Q;>NT6&O0'E!M(@U0\-&1MX,<F1%TN!J4
P10PN?\F/VN'X/E$AAF7^+G^CT.C_;]+PG ;F\3V]NWRC1YHN@0THD#1T[M^#=F3C
PYF'K0HY?N-A<M EUE;))&D_]+BJO0DKV=L6U)-?EEJO'7.SJ]M04EUPF ;??'??W
P8^B[E\,RNOO<- +Y"M+01Z0#'MP32Y:N:5M-0#(G3=@E )Y_O4N,B%IJT?=<200/
PA&L;<S[2124X[L2].6$71ELNSKQ38]Y@?L-Y7AC9O:LA.;Q9;DTGN<HTK<YWV"#R
P?HSC9OE7I";6WG9H=J//\K5YS\7];Y3WQ&$JN(=.V3*'/3)M;9SZDW7HAB#8#94_
PAU-$+Q/4%4-'4N+#:6-GY([VAYGZUUGG&0*^EN*-V^]U!"3H''(OTF+N SF[L1K)
P9J8D;KU!*VO#ZS6NI4)X]OCM]_II>2>]$X0&J>N7@YUF-T^AQAICG==C?817U=BL
PU#W:>VW!X?O?EUXRY'+"9WR?0I!9"H!(%(OPQ1G:#Q?A8T5JO.__2)<(\/B+(>#R
P=:=<@U*!?6O5=?36!Z'%7DGQT)I7J%_:E+N2'#914G\Q^%)^F@',QA!2;G(='IU?
P\9Y>P-<$2>\*<BV4X'2<I]K>0@7#8KN:/U'V,:.'Q'$&I$LJ-!)Y-]68?)FPP>QT
PEGUNC!5>"J]EK<9US3GB<G =^Y)-^"%7=41*8"7K5Y23)"ZFYKZ*R@YZ[_RG'AY'
PX[^4]L)+SF+;<KKA>AXI:&!0N&;7*>O"*DY81^8 @DD?6PR 7'(H:;JYL9;U'5GW
P1T),DXG"]>A]_\I A4T!,]]#::# MI0Z)G(+P0\RXXL"UU5ROAVM!2<NN&WQYP]H
PM]S)@)[U&V"\Q\I!^@ZZ;L&U;-\$ \O^F[*7RU8M2_7N(+!3 %Y1AN@&_KI+X%/A
PL93:<)"$?.Z[3\T4NK[@.7,@_$BBG=C-CYZIR>%*3NKDC<Z !(=S92U O4C^\DVE
P@BJ=$M>]<G1C""V:$2Z/BNFMK$5Z2-NI6@6'G(O'H#R&Y2PHG>]7E9#&.EH@<1NB
P%8_:?.457(11PN",ROO8#<S(^RD3K8K)#&/ZL0O,7[O8MM-1:)R@Q57RL*;H/32<
P$8$N7#*ALFT'&9L0MB!4-B6)Z>(6#ER_T2!P<F3U!9C>RU23\>.#VN A=+CA[@:U
PCENFXLW(9NB-<_H;^Q/XC*_>A9Y_P/N+B%O#H2Q>U>3QRP-03$A3^%*%Z(1;7"6-
P]7Z3-!Z)_K4WIUCB,RF%(E/\./]$$%QW-D6/,)CGO$.F[7.^01"VAC@ ':(RT*+#
PM_5#A8*+J;_@)MM'BPF\;DZ>Y<=X^9$V9%')@4H"7M8X5#\7G)DW+^5I" S>W_ H
P#8%LW)9C=37FFSKMST?00S3Z4HR G[([H/>\]#)?M^AP6VZJL@=*VJ;I_+G=EZ^T
P7_#H9ES9TD1]J"[01"20:5<JR*I!:V0[!<ELQ.,>.8M^_2/X)T:-C>;IC[NZY/O*
P)L%VSL7$#8 A@Q2%9*PC6&;JQ^->"" @ZAOOD>WX@YY540@X*"_[,_:@E $HTQT!
P#Q(DED3G9)RX) O.=WSU0F;@, &*Y'6?DZZ[^N*)L@D<+$4^Q%',5YMH?OT77 ?=
PG.[K *]-<0E%_I[H8WMFTA:\=G9F[^4,1J7H4L4:PY^AC_B:=THT=PEO-P0BLDB6
PI6K\<XP<T$"4 ,$6Z-;_[V2O1Y#+"8&=_^J$@5: RH_8:;.FV*$X0:M>!B,G%KN>
P?LT#F08QJ"-^O>-"<IQ0GP0X!Q"8*KSLFGAO\HW?#>O5UI 0^I+]8V"N>M890U"/
P6^E:,.*%BY:%@3Z"F,;9]8L%<"FC:4FWU+K]]]22*RW5;<*]<@._F:C]L,US>F A
P]9(OG"OONAGE4[HN5>:W1P>Q"07,ME&%B52/6GAT=,9_ JZQ%^=>2CVY;)4"SA\)
PFY!JM] *H)]N+&/Y<ZJMG%Y (*UE6:@C&"5F,P.8AO8&>\6)R8E3&LEP6VC5HQC5
P-43U$B> R&%@4 $-RJ\@)(]'_QB$"V!7Z[T'X((O=BJ W!XJHR&'88^4F"023C0'
P%_5^HC/,6511"QVJ9RA:&?^Q2E1(HZ)LO#CF9??,3I]/=>Y#A<IL[]\43*[^4?.[
PH8XM:)5<K7#LF<M"(#(#QVGT #FH@!$SE5#F]L-(7QD&=;;83)SK)BWHB5\.&NFC
PFT<BDHS42U[>"3B 582<&V]TY_)\ Q"NR$[V]/&SDF$&%Q]!3CZPE7YA1+[J@P'O
P;!AIWF'$2"O]<J]OEAX5M8/WM'?.7S. OM@I^O!S2_?;%S68IIJ9Y!4Q[%(N Z!J
P/.+5L"VU8/XQ6?\CU<^41GF?TI#W_IDCC@[A;6>) 1@&L_,8QKPXG2+=YX?%&IMQ
P 5: U :C%,CHTJM8M;<COH$_'VL,@@*^I- JC@2[+OMM(5]<@D=XR2F2[]XOL^NT
PA$N",T-)&5E0[*\U6\FQ^-B=#3% WA9ZS^/HF,<.=.4<H!G8.>.EJ@+?_FJ\^-Z>
PJ3:M16SDJ;E=AA@?-YCSH7:/N):5P;6Y>?WB]V'>[UDUDGH79A%[U#H8%)_:2^4?
PP4C 9I[%6EI>D8P;JAGL-O*!^*;4XV+C>UQP@N[$P4XKPG*/C<0P. ]ZIW*K(5^B
PRF:K8I=:S#.*"M,](O@&]%EYHV#>2+\9WT?>)VVABU,-<U^;0RXJ7HUX )[8N5,\
PGV[UY.^:5_=%0_.% R$Z8!C/XE:,P>[%KRV+]>SL:R-"NEBI9T'Z#\ [?YDH$^;5
P?L'N.75N? FQOLCEB2Q:T?BB>W]R"\FVIVLUWB"W0;:;HP_4T9ZR<[".=IH_C5H8
PG&4HS43+I>%DSELN[JIZZ4V##&(>A8G.=JGQ&FXBDEFYAN>H25;/^>XK*RZ%UPGY
POO 'B3PQ$A$MSM@X&9V<>TMK(\0^T;\3X//F7Q6L#I]$2]'!Q)1.\N:Q\X*R5OI4
P!3T*M3I@-O(ZJH:@XF7A"^?TOF0T%H)5A5TI:C@K:*'DP0&H!6K^X#IA()]I-KP0
POT)HI8'Z@Q"36MIS<8*E &C\H1U;%$?,<X')Y"Y_X@%S0\SY4^EX_\Q49U]>;47+
P]Q9&6>(YIJJ/J5EW@I7 0,_[PCD-P&Y3J,>?[H]"*->-*B0G9#8JG55*N*&W"3/'
P !+3@K-3M L E[$4_0L_O'F7<IZ.?_;L?^GUH4+5T\B4]X9'=>-:N!H$)6+.EJ-<
PAWA$?P[MLE17J#MT/B9T#3 <!X+'G0(M(*2XDS>_1Z[G55'DC+O_EK*PFODF#S5R
P+TBR:TPL7X_6R]_-#3\9ESZS]VC,Q6+&1"[?O&V:4.MN-F !DJ_FY<68K7<5(JE'
P2*- /VSWGM*M1H7J^BSTCFMWK:YA>FC>>;#I76@'JK:X.QX,_NL$8UQ1YC?Z$?#D
PL3K-H7X $K7BS:>DV500R0PCV2_&%U#4%REA[/F1R)(-.L8?\+6:,!8^'!DH!<B#
P=W^(#@RO\OU.P0>-GO*<_=V+J'4Y=HO$5995P/7Q_\WBFQ'J"FY%,:[6+-T9NHZI
P!M5?L <OOETH,SI#+YB8FW*N-/<&?_[,R.D79L(H-'^;!@5>!==H%YD-[9V+E?2%
P '5""]5!"&J48I<R$D6Y2I# 31.,M Q%9'!I&W\SE(SFV@+Y^[C ,]_F$)ECV#M@
P5A8,4'T7D53,@Z99'*9+0;1*G*@,N4-S3N[A]-[IKOP5T%,;&@TNV:C]^'75(B2K
P=O:Z)C+'@,QLF.+;.ZGF+T_$]U?*"Y'QW-_7_)Q-K1?R%3BN#1PYMG($DN+RCJ9;
PF8!F)-DL2#"8R@&1@E]XM@K -9J'HJ7_L3Z>UY '610A0^>/W2$*7RVP<&5S+Z$;
P:HP;AY9JU,N/PZ2WK.%J,YI?XW4:\D%%PEX;.'DO@#S>U0:W9%OHW5Z[!$S>$6N'
PM'S6* G-4HPF 7<08WU=049%C@\O3WL]?" F7Y)<Y*UGNV:U-=N+BTT]FON8N-+&
P[E="')AZ_76 >FZ13/[#YET^+L/ZX%VLQ.<^):0%A]%JB)!#'G(U_DP* V*J@1!,
P,J329R'9V^.1@GB$_)G#\_*-/A;T0'U];](W\!%HQ6(ZA6B,;9#NL^\>]X?Z[>:-
P,I/!)5E\^3QEXH[D@G#]=*4T*(_9<;M@,]-K>!KU[.1$ CDD$\FR/(X2A*<7$U]L
PG!$MKY)\?_KXW35,+7\K2X>G-6]F4.L$Y)2Z-J-BI@,CKM)O,D%Y.A&H\X6ND<"D
P=/P/A@-V2W#N<+0?\A3I4%S0WWW&J\:VMKV6"U]@P34Z,GBOZIUSWL.(5:8F+MT6
P7*^BC"X$49\ %TP#VJ]:Y<NF1XJ/:<=]3WW;!&].NV((>[FU06+:XN#)C!M?@1/3
P[+=:EB'# 2MRVC[_#D1\)NLL!S%N UENS*DD934<KFDBD^0B4'4?J;-9?I+6E1)0
PN'Y>R+WX_$!/-='3ZTT(8-RJ1_@\V,H,]."^>P_RSHI6Z$AW$)(VNE/Q",DG!+FZ
PE_XLQ_;_X%\O_A69*&56_/A?4KNF9F*&-NSR^^1T'TW(>6__EK\05G_]BY"88*^_
POC]D^@#Q=Y=Z+N66HV81*O[#@$X#KQO0J#N9A%D/>?=X4%Q9ZX$]6?0;%2FP\:Z9
PI3LX(SW$4O66A?J5BU7[76SXU$64BB-/0J'$>W3S@&QM-:N]-G".<WM.!^)GP3J/
PIXMH_2@QB'MW[ 9L# !#_+SG<6G#$E2M*@XSSF>.0>$X:LH2#73;312P:JYZLKA 
PEQ1D#S*7DUBA5 C^A4IS;["64+5<I6,@1(VRURCF5_\2\:,0'# OS!0U,L1^R7IX
P%%\J<+9CYVDYL@%#5'S04;S$X"HH-?'W-47]A8/AYZ^3_D)R00,3QP 7P9CV8YJS
P:OXHS4]@UNJHTN1FDY+B@=V7JDYS(+3M>#<$YC&H[7S,FOM5LG6T.T=XHN4ATK,M
P9O*2!0(&:^;"21$V;P]]Y19FQ7+:'G*RA4@@P*)O;/*S0&.SXED]@D';92?4H65!
PHJ*;W,.LL"8WT2MV](J;,_7.)2)C.KY!E5?C^PNA(;(#PEWJ^1!F6%;^%(G?7"+R
P<LSJXJ&R%D%:)6"8YXO61O8UO R^NP1GO:Z7P/@YN_90P4>_?^VDG4;R9Z$LRRL1
P_6Z&,9':0!V@)_L LU=E@Y&C8U_&*^E(_(FF)#?9.'*3409)X]W)9'_3"QKSVLMZ
PPLN6F6WF; 3+3A1&I;:^HRBHI*O?V)3KS:&*L7DP8Y*P;N7_:-"4U):[,M?DM870
P>Y]]FHH[Y_%?&@0!U_#U\[Y0B1N4%:V:C^A^>9X<7A4\.@"_W:C(W7;-N1\BP#>$
PC?WK(ZW 7Z56@"MP*5KKE!]H@8UL0*_^[A[)G96(:+H+")%V2(IR\Z/1!](*Q 0=
PE^IXQ;[6Z!^7I11[BB8J8$_M=GML2=ZW1!IS6GF^OKAC:OQTQ?18=0^;H,2XXZ/T
P@H)2+(GCS.6(3973F]R+!E;HOIE@?-369JH'^4M<N7+C?0K-K=8X?A"0P^0E"5Q>
PI!@;)P.QD^V;!X\;<,L%\H4W.MC%?;-5U;V*9D@#[VW?/*T?>F^'0$&_ "J2'%&_
PPBLB63LQD\W4G<7"%-%>) VE$1N LIJ_N( #XNK6!V5@%T$P"ZXVEW2V'NAF;:T]
PI-EU/(1S,.VUNY[+G$J)D#-LY]B)(M?*[78<OA:9_7-3\UCOZL40J5BS\DA\,=J=
PZ+KVWXVJ;#0>M]FY%=RP)0IKU)B'5*Z&O;!X=T-"S$X12E:&*D.*LEJ+_@LP::4K
PI5ZQ>38; 2>.)V$4AU +@-^K>RLO(N%JG0'.,A*#6K@(XH&V-A[Q/O.S7#9T-RAY
P0:!AE:RWUWW7K@4O6*6_+-B4XBL4"D#HJF<0@_R.Z["F)CE:P!/-LE)_(SXF2<NT
PTF1IIO^5T]U87U@F[OZS! ^[NN FDMQ^9QBHWCC&<A1J)0'UX%6<O1QOPQQ2] F^
P+O$Y';JE9Q4V60W))+NK4#W(3;V*55'8MFF@P+-L2:4[ 4MH+ZH3 "V_;,.[<OSN
P$>[2K@IVN_;R0Z:L9,.7*6?H_8 6!H,Q=%-@E%TQ^/YZF2"(E#5-EGB.U8E$UN$?
P.3'>H<5\-\P_U"1N>/((V/;?W_%D)H@3*KT^_:E^?UB \AB9EA'H[IQNGVV3E&]+
P9.E<I1&#5L<I[$.BC^2ZI:Y30#SL1ATT)(C,-/_1+H;PD[X*T_'-#A.B&Q_+C:&,
PJ4E(-W(>;*T]P<0>F5:\ PM\%.T40T=ZJ2MF9,$/CRI'IMO959F!\$#]FPC5DJ?:
PK=G_#^$9G/6/.9.A=B-O;#4_UBB:+R]%'6[\"33<OW^:\;GP45LT(D(?]](QLLH\
P$OZ2T@VL!O45FM5G$M*(XB!9"^;T%2B$1/Y;[!(N.K5 L4=CZ2(%^2[XR)9PF\_@
PQ6S+TX!G\\Z$BPP,;F&O[,*=M*NJR!JG G)5/#J.:\F:=]X>.^M;V<;!W@E) "QS
PPWIA\]T>:"X82T&7TN. _N&,$TJT=5MLTF&$OR3"GV-.0W6?4O<(&G5H72+,\:"0
PY0-7 0E#;[M>%J =M$3_FUT)6&+X#,IYT3"T5LTR.M%,7)$. /6$H41JJ;+HA-VM
P: 8Y.'P["!Y'->G59'=;(HKW]Q$WDOH?$<:80;SSFGK$OG"T!8127"^54*Q+;S$M
P__+]*_@A[W%<IC/^[X$QM.NT5OCP+(SSE<VNI!^+ >0NB9U'*A$I5N8?AR^>FTUV
P!+/*DF^9KF4.C=J\G5(@TPL)^VFO;CI1?<5"EW'G@>QF>JF[GQ4D90+"$>DA:#P4
PRC*&&M4*OCG*<_--LB/@U/)IU1=/8+1%):)C@56)Z6KFKA2#<_8%49YMA!'^&1FD
P9<KK'[R5/O+144S$F9 &)PHOBIXVU!*V+6X^IG)0C%:-YV&71!CFB96I"OTFS\"G
PEFQ-B@WO;Q%:[L>WY3)7@0<GF3^Z<$YI?&?O0FN0?G:,N29+VQJ/-[U&]/*S"D7G
P8"(L^F_7)L9%+@-X6L]0<NL>3R/ZXW\H>[AI$@RKQ0>C*GNWXF5AAS>\H;^^J<6/
PWDIR8ARCXOU9U;8>;2LB5=JG)X-$<HSN637#JCY9MQ@I.W+:\K(4)R<%6ABP[YJ)
PTK%FGVK9NPZP7#UE521:NK9Y7<L*MQ,,G9!.<V)^_/>QW[0L_GF,[(B]TRY7^C!!
PP"PN?$\\$.#E4XG+TJDL_UFI^Z7L-ZYBT5CK&R Q9258/0CC*8>A%8@8@0U:.UV/
PVVY:JIP(.,!<YM][.%"E!JZ@F="[33I.CTZ)IPZYC'-&,?TG?K;-CH&6?7,Z9FA_
P6G8ZG<81,U@>=0Q-94C<GM[WQ$/UM1QX?H=:MS.XJ.KV)^0?Q!LGOZ^R&];VB#QN
P-27NC;<<'&52S_KDS"OE.>,D19MN$C_K0K0LQJ-+7I]+:-.6Q';PFV<0 ZY/?&]7
P;VE7WL'WC$?6AS<EAZ9#4YJF)=6\4^_L53*D^4AR%\M':Z3JF=BQ1#N:\YH8HQ3]
P>C*)QU'5WL9>C[+TF%=6?K5.!IX_#N@Q*Y"N;Q;N_.V$=BS;X>NBM=(K0G_W'51Y
P")?Z%+>M56+IP?.#BGDN<]PPE8I4BB$ZTH%YN!Z2.MFWFH$L[V*2TDNZ(M'22&6P
PQUED" .Z^$I<*Y\VH/9E0<8?$M=#V-KW(6LBV#1O7+PP]Z K3S5C!A8$")JXS0S_
PST'15K]8I9V9>"+LK-MN@L^,#G7>S"Z7R.+KY&$&.4@#T3<E(W2([,QA5*Z"8 V$
PE,O%.'BD#?KXT(/.>_+I7PL)-C<><@YH(M=H$^4]+@?NVXO#!7IUEFD<MK?JM08-
P&^(JLNBWZCS#*O+!HO;/!*%7H& %+_W>)Y:B;_&@^305D$VG/[=[?X6[J6DH)*(5
PO7\J/Y;WU\RV])\OU6=N67&S#1>4F;W+F5*2F:4^+B&P*H/!N[ %Q:(A^UN\;3%Q
P:X3%57&UYVIF/9=4>Y#]%%T<5"6CKK;82&\B-K:H:-T@BQ72?;1(?-]/)3+8BT*,
P01FLK-*I_X'OQ2HTCCVZ%PNJ$)CPIP:Q.GD2;S'4D=YN='9EOUNO]K&*KD^KVLB#
P\K7VR4KI3$Q+02E-\F)?6X>]T1:(S5H:U\L&RUK]8S\#SQW)F<9H0_]NWD>" %0_
P@I$R%ZR<E#TLN( &6-*C#0&,MIS*/-M4\;NQAEI7A%K/K[7.84"'WB7V=Q#68-ZB
P4>U#<X-K*P1/ ^KS(\0\&YY3ET6I"OX:#L>##-ECGMZ9<"+_78&EY6TW 09.&4^J
PNA]X1+"8EOA8%TK7/]U)E $T0:<N?(0T\KEMO1#GW#%7.''#[@JCM*]XBOH?M8JI
PY%I,;L^J]D1OU P:4M[9O. 3B:9M.&.4\2:JHF0 ]/KF_CX+=V(O"3D?Y4L@QCL#
P<%JY!QHY%I)?WD:#UJ9 +JLSUFG? /@=-Q"64V&U>/ OR@1?_^IM-1K,>[!KLX^%
P?S> &HV61!4]9,HB0)AU6KD%&+5UIWK$D2<4TZSUT;>JR"#SI71,:.=H0.^Y?D6I
P:G%YO6^=NGHF59M&'V;3YCZRQQJ8Q&BH'>DY!9W^TSAA(\KS;NOF:Q0<X^4&]Z S
P0W&>VP=.J)(I+E"P$6; #&$X0)-668*W6&.6HW_5+\"UQ"42R_"RFDV4L#]T8;IX
PRM+0C/[YE2U?[Z[/>7XO<="7=;HV [K-TUJ,N/Y:$6C^4^W=&UJG-HD%@]*RRYWF
PJ$O!UY6N(9$<KO<$M6?0PEP&%>9$WK&?7&0+3-17;F5W>!*[:NE>*ECZ>M5$#0$V
PS?\J)2&TU&P$O:@!'?E*:#>D8^Q]G<6.P+X[!EZ@')EE%AMQ:F )2P&?%+#5O9%!
P.&',71)GX"M[+&II>6!P'WARZI%_;&U]XC)G!K&Q"OE]PLDC @I2:9(B/QYS_L#S
PO.&+8A?3OS-\Q 1Z;&#[P\FMXL$<R:]/C[OGMSS6]F4'+\,[U/V-@3>"0O?Q/Y9K
PV,-!/(,8IZW:U[YMXP,+%=\I2-0&(M.WFF)+>\C0/YCJ-.1_P?=KJ1L^0-V)ACO.
P3*5)P-80.#0W1L&QCZE-FD7-S6^C.)?"KU%C/Q%>QV[?IF(LEEKZS"</)>)5:HD!
P81V5IIGA9:(29(:*R/S<E\C,_E6W3>>+UU]H, 3"EOGM^,;Z_ 77=\(=OV_;$4^^
P="6A6&5^%P"OQ..N9(5-[.A<F-RS3G92!Z@Y3)3+GTM.)K<:U(+<71M)LM*+H H*
P6,/V >C8G\2WI()6S,$CT<=2V5NS&__H?SJ,\WR,;@+GZ@U)1RWLA9I':-&9$JX,
P* S_$*K,"=?: ]@]B21+)KOZ_I%*&9*^=GJN.Q30&;6ZA?8L45(]#5V92 6C#^D&
PGO/]RBB-(<<!RA']I ^I09N3IE!@A^O/0!W&>/7 18?F![N12FIMH=OL4Q1YV5SB
P:-4QK0YJ-E?-O FB:E!LO=F@CR".DCN$N_AIM;+;%*K_'_=Q2CYC.,J6@E-VD'R6
P@#,#&,4^/31QUSEDD8"(Z.8E=<!?U SF3,:P$II5J'9"M#6T#N[$="R(012M\GII
P]\_4DN(<;:U,9%,#+6OB'<6?3;JH'NRHVP0/B[_$>S%M;1Y].-Z3=:H*:>GQS;FQ
PJ6LAK' (,RPG_S\[,=$VE3 SH4C!)I?A"Y]Y\;*:%2[<[Q)F4_RD)R*;3G&%]04$
PNW&<\FLG?PKKNW;O)1.*N2&C:_(6(F1=UN!\=46T1MJNQY4[@K28R(.D8-N8BC9)
P,%&?76/^W;X8;?P#I];*"V@+5I@'YQCO15#8)^4<7SEF6;U?-%9(L4%)7R>-+Y($
P:+!3Y'_+ZGI+&;Z#/"CG"6\Z?[5%+ID\OS%K$/H'-9X$GQWK P@J(D,2^RCL)LT%
P;^#:;QV7ZUNM/?J!R%$Y2]WIOW1+6&88F<((* ^7%X)(Z6PR#-=Y'Y:Y:3:@.Z$V
P'/@K:E+;^GD0S!*@0I%U3FY+G/A6C+Y'MQ%)_G? %Y9#$?=^T=.^M!3NL@)(NQ-H
PVJ?3N1?%N#5I*-\$8P,P+IX1= K T=TM?/COF')2>TQOV 6D+5) JK''4FOY0,UK
P$,,XA7YE3]"W:YXSBH'R!,BHK*82?, =?+.&/B-7A&5F+&C#IR%SH<MT*Y%C\,I1
PJ,DI)[S6=@MZ/BV12#^S3.TS+>D@K=7;?E33EH(*\<7-ZBR-67+?BJ%M2 G87BW'
P/O'/ DD[$\CVZQ<* % 1L&;0^%HJ=W6M# P_'#"5D6./AMU^^%@ET);#>8.V1WU<
P=[/PMV'9=8AX'VK?L2RFSG\#^ZTL?=OR\CK-2*8[]X&8 /'MB!EZQ\X L0*7*WBT
PT7!%IG+S,\S#1N>_8IC9F:!:/]R"B]@31&9"FMO(]U;EGCY,..WW(IP>3(!-CE=%
P")GS7A(YINV,*26=_ZK35X EIFROA8]5O[_P+2^1R@,;W&16TQ)RQ'<P"'.FKS:)
P0'"RHZSPPOHB"L]&KK3D8'X:L^FQ@#2=*Y>S%T1;@?%&L0BMEA_J3MSTX;531BWH
PFM?7%JHKSY;6^T(=4"AVFU8N)I_PR25^UE4#*%<&#L.<5^$3K.7D]@ 2XEY"=C-/
P((-<K@SG[6^GLPWZ0',*X+1IF*_*T%8\QYJ99J?*,Z42>Y(P;=B8"U]FKBSE.(64
P/R<]2*CE23C3R>:+8#"KDO*]D;)0.;"QE9&5=N$GCGM%[5?7C)UO+OJ;2/@ZBELA
P@)$6"Q-4,&&F3KH&?'4],;_[7E?12],G2?H#LL8\'B#%P13:64!#'WY?MOQ=)/*P
PJ[;7V])X)L3\8YHK.><0[-DY!"''+@8!K^ZXJ.-6#U9H;HB:/.E.^/VP=AHCJ;[P
PX< BG18,H\%D [%ST1RTX'=>T)[:@]:=:#&4F8H-JKJ:XB.QR,2FV[<=<<9X"T^+
P@Y78Y90*H,BF GJ]\/1L,$*)5"@.%DB2T^,V(L,=J+MA9=:IR6*"O"C*"3#TVA@:
P';/_(HNAZY,')!YX__-B<E50(#[E:WW?B-?0\9?I=Z[SU#9!O2)[Q]:DD6\Q[<>8
PW^*=*;%_$^PK?'OI_J";"S<']UJ]VP5+KAP&/V]:DJ?D^> N> _T)MZ]T3>T[>@E
P)466!W-DPU5]#U/A0@+R8Q Z!C8+>JTZ3H!:,,>=X.\U*8L]PXF(HRSJ@@-O=%#W
P:D]1*LN9DBB +W^82S*H ^.+X]S5Z+@OCKPJ;<#V5"A*\,!2Y@B2%52BGYDT6'R$
P38TG(Y2UJ<>$,B4NNGWOH+M#CZ (BQ?]=EM-W!/1<'+N5(U$?JL@$1*;;E)5;K?F
P\@8<6F"M;8DSTY?JL_ 3LE@J&]G>[H#3-N'E]$ZX^A_F&0) /&^M*>6V/IS"DJR!
P2%\#>AB7WEQ<_I.HHL'=DYTWXIU">F8<C;0NY])IG(K@!-Q=3*T(_B[?C3G/#N!J
PYR0E^J&2/"C52"_%-'8X\@0NL/2 \R!C480)N>_V(_EIOZ,$--/RI>N*!89!$@I\
PQX&5L DH8\25IH*$F[BP(/Y4;LG#35%8-MH?#833DR8AA[863Y(:S['2;UH^\?\5
P.F4ISS+X=\23XO:2/5 I9OUH/@RQ'^OY/>BKPP8]?6Q_7NDA0%Y1U@>TBOC&+WW:
P)EW$DOEZ9,(3#&![*$?0E[6B;^=X\K6[@OU=XIK(F,E@C00S\?&+TO<>9>Z\DY%"
PL-[/?1JK(I99V6$ #LN$9V11KH5N6Q43R%,PHQ08GBA=40S+. $#@NAM0+<3TTGW
PFRZ=+?WQ>$<T1UW@X]J&W%%>0X-FT)B&61P\S'$4VAG,CH_FE]^;X"R%8#B7J$7 
P=LM]QT1XK]&M#!JG>=@CW<B+/8U7J]QB_%4 A!C*V[N!@L)UO?I6F8MHF(" 4_G[
P7\DQ3&?W9?JD&;G-'"YT1EV-HD"ENHM<(MF(\>2_#KCE.16 M;\[,$RI[WJPG3!&
PK(>$LK[+!#M^'8LU\IWA3Z:G,2_1D_>>L76Z>W,BI*P\)OD,#=R;.?-C=<+3J97$
PH[C_C/3$ERY"A6L=.V!AJ@8;+J=WP9&]I6I4'.R,AZ(OA:F-.-?1HEI*&"@__A(J
PJ#L(Z5L4+& B+T?&?H3PP#FHXP7>ID[+OS.&AGI &NF^:!)\^Y#98I3$N:;0]P[ 
P@.?>F6\U?<YIN;TCU>C22]_[EEM)*^:5A\$VAT,]QC2N#RUN>!Q \42D7&\"U W?
PTG/X_>S!>RQWF0I 8.D#(6^XDR0]1L- !X:X,0E21&"Y8H\!02=)?WUO^=+ 1VM#
PN1>(/6<X\)2B@&-U"<209&IG<RWMOKNV5R#WM8"<@%%F>1*HD*J/,^:8V:R= N^#
P/_L8BI(I.)#&JW32KYV(TB2HUM#Y&Y0MJ/7P)O-NMCG4;]:.)BRD%W-M+ O^P]!X
P$B];4M)"M,K6>!YLWW1#A2O=QRJLG9V8!F18?FMXIYJ5_#![Q6-%O8">0IN9[[]8
P(F594K52R;"5I:)+4OL*"P#M[@D:H$:OD2W4QF<_@K@0,PN-VC6>TLBPGN%D_X',
PG3>K:7L9K61]Q*VDRH;6=CO! $AJ(W3G @J7NL>4C\6U>?6/OA#G<Y<D=2\,"6)3
P2HNBVT,W9;2%'>A7X]Z.15O^<#56<-3(('WGW& G)/?:":!ML0IA&[>)V.O-QQN8
P<M1)@?J87+1O)I%T6"1V!<A(?T(1EW]$$6@6&B#QR:[*^G\S MM'P >('4P@52_8
PQ5 +^:/Q<6>[K.;(G%QRB 2I<H1%> F:#SO#)K"*XCYKXMJVJ^74%]!(G$@^O^+-
PIZ&5GS533@KY@5PY<%W_LZ.RIL!H<100\VL>Q=J/I^_M_S-YU=KVQ'[7&+XTPUEQ
P^/$0];<FN ,'Q!%O1<WZ/0D' JTZI#'P:I)[#:F5[X<5S[UXB8OE&D0KYU/OQ&4>
PCN1'3OH^ 7$: 6-IK&9%=4B )4']=LQ!0+]L[!*U!J[^AJYKP?V#[.UJ$"L>W^FS
P(P1+!(JYPUK)N(0&WP?@!@51CYZ;)?D;1P9@P<VDD:UQ/U*DQ(H7 S''$IQ.2P#$
P7N<B 3RA:EC(Y]R+C8.D#%+IMRK '*Q^]X(0H_=A1_UDF]+D+*N3K 0?H3G=Q>:;
PNR)<L"?8X($E;!.B6Y]8&E\.C#2X[+78:^-K75!>L!"%9LX5% 1Z (<Z?[S[/^# 
PO[7/[,G"R!.\[<#+T(@T6%D;JGG?TG!+^<Z_&E":(/<&R+5F3J@'AD,1]+_.K]A.
P9UY36,E24[-C)X#&6N05+#S>%+.LQ\TA2W44G5]/*%P6Q &W HY'J]L\'1HO%9B&
P*(HP!UC.4IL; J?\D\[3*8[(M0SENDRR^<*C$6S<S:';?4/6V6'[GO*?K<.Y^H82
P;B5WZFHMQ-VCL%76E-?<+-/1=VF<=S@\U=NE2?(:R(T=]L+_3H"$.H*]#0GGT3K6
P4_FOG@PH4'82&RE+[J\9T"K0B,?.Y\6^;'4L>?_,M33=://$@T,U'9*+P1E IHX3
P,$LR%3+6KST+1RI*,7PH>%=!R8^Z3E-#+*G#OP$<4I_,;Q9,3O27^8.TI&39^.&M
P80Y( '45;8"\BJ.:#CL"L-PX5.^TT@V72\?J7ZR"M#X5T5'V_*[>5C?;*PU8!E.K
PV@HPL6$EW"+>I-VD=[0[= Z+QZ&!$5(!_F-B'W'1W^91CC;CN6(K>_G'7:GS.&;/
PA':K*GP5$ZEYBV5'P@DV(WL./1*Y!'KKA!UP]IT%[ .A<HNA.39Y)R_L78'.:/8>
P7:%W6'[>:@O*M^5^X+1 HXU .T "US'XFKCY/U@\9\3M>NHXBG?I^E>'Y@8U;SE0
P/,ER$;]BO9JOMK(6V"@)VV;TM)R1;NC1-6;?\AX"MN09Y44>@'Q"3E3G;B-Q %KA
P1W.E9.S\ D$&?^2WF$V<IOP^["E1?-6D/P!&LZTGWYGM78<&SNK?9QOZ 03G"3A*
PAK&A#\"N<MD<NO=ZKYRZEV@)EM5@Q;H@]T^YQVL3B6UI:5_KI/V@">OCW%8: <*=
PVV<V+YRD3E\4G;-%I&C'N:EFO5FJS-M/6 .QXH2.M"3Q1N9]TW'D$..M[Q"R^X[S
PD128:I"ZDI%37)W84!Q1J@C<,<UN]BYZ^!Y;*I4KZ("%PYCT-U9A$\7N3;'+E-RD
PA6FG50R62H=W+H7LR^Q6UVC9W^IT1'SM*7@TF"J2F;X-4N:;6H?XXV+YM)&B$7DL
P45J[JA-+3K%<4D;P0@M8#O1JM='^_$_MIP*R8#?%V\,.$$2SM2&PY;P*X(B@O:F!
P&,6LA/9^'6;$T(C.4(Z=K9P'(EOJ.V (GE+\>3$B2]OPKDG*_.C2" ZE]$]%*%)S
P(JZ:J<3F[W&W/)N=4.,UK-[:@,O#0RF]T)Y7 =_AFJ;%(O,EG[(5/@K\M,@T%%GX
PV#%Q$U7YUQY\ZKG,KI$)>ITK8H)?+"0"P 8)MH)<A-D]0FI3T)X ')4JTNZ=_9Q&
PX^FK2E/@_9Z47GM M0PJQ=.I?Q&[I8D&/K\OH>"JGBYTC!_Q!DV[#,#Y6J/)'0/X
PJ *I5FRM=&<O&;N)5].XT5,+KKC+:$3%)L2O@*?"AV[\QDS EKP,Y?#UKX[*AHE?
P%P(XKD?MF##Z]N\>,9<\X3HJRI9J^R5-,*A)@2 %P(6<^K[TJ1Y_?/>8_,OQ7D2<
PSAJK3+()#U:/V;&[,[YI'#K=AB33 %/*T@G 2VDU%^DETUVLZIWYFAVM\QK'S<(T
P6I#!FM6]*WY_TXE2/E)+<%4.0<(VSR)5?[VXC;J\[-U_5^-OH#F>,W("ZC^1R=SF
P]6.A#=03J]XIZCD?9H#_LN.MOF3H*VJR5BG?CH^0FUUGIP+][+I,1;NK1U99&EA9
P56#!]JF.1KU*22.-Q5_-V3=P$G.;/.!Y0O$]Z#JYK3$Y-7OA;\%%>Y#> 5+3$$FY
PMO5/V[<#@7DUH\"A:^C$1%YB[M17JZ7!I,]/#:%DCS3IGRLH7/M[PS! V,PAA\[^
PB2[:X@)BXT713_^>O7#-JGJ'!/_@:X!H\H;QCQ9?L4D4&E.K*188GMU."OO$(W=1
P$#T!(%^[N5\:4DNC*0*Y(%!S"]8F #H=(^WEL.)&:C&#(;.?$&,PSJ#Z.6[L;\1?
PP!W%H?P@8D><A>O2X 2KF0(8Z-=#UNE.<5SVZ "(EM[C>>U?&]'9 29QO]-%:?^\
PJ[<7%(3.\2T#*$^P73![KZ/(DGAM6"KAWIN$(]N=WOR<J0>ALJT+9N1P8)N+JGO)
P5A-&UX IQW@O'(LO[,[E%L"%$^"BR)=DC:Q)&AA65&7\C,99T32(N^%X(WB<P#83
P/=R^3"4YJ=%C )C \<J!J\L\82ZY; 6%)/W!02BC MXG5R@M+G."3[FB&EDA%^F;
P56\)>IS,P:3X1T3!.-@9P_F=XWQ/&FLS*S[_SRK<61WLYU:=)49HJB34,Z&L5?9-
PN=2$X7^&B%]>NLAM# 8[*8^"O0^"_R#K"R4(%].X:;/S*&%"1WN:0%F5MO/[>G3\
PV&QSMU27'*3SF>&MSW+AOK!5$Y7&+4,+ J(-N:[#@25"]YP<).=^'$Q('_PO9"JB
P;J<Y7KW)10&!/%N4Q1A;_.)G<2<UUA1Z&AVN'F]#'_ZT;L8#_BK8XD;:R'K!O[ &
P9Q+@XC\Y ST(L7EH&$/#,"PJJUD@EGO+K@:B@9MK+Q%FSVZ/A]T?FHV3NJH7(!'R
P=!>5,P Y1,$$1JY1#%;[TGF_"9=@Q^7%#KI;$G&5J;$6%8W!VX%4^(<YG')(/AI/
P]B7QRC904B8#KIH6AJV@&S!8T.,@V(.IF%([@2C<,K\Z7GA2@,.'UWR^/N?GNNO$
P.)@I_:!>AB%%C/,52^S7"FU;=J)(E.([@MLS $2G3?'C8L(+1_0Y(L+ 6,[3VYP/
PNJA11CLA=PB3E.]^JA,?;#=,:*^\ATGRNC<.J:\AV=%^C=>&@'WYN*32$$@L6WP?
P6DEVMK414ZU&AHL#LH\U<Q'0<R[8J>Y"HZT615VLDKP>4AI]M8'I-#7.TW=>-:F@
P\CG,/%6HR5QYA+JA0&X'-2,];5!3_&J):? MDM \0PWD (E:!K0V\%;JMXH_ JS7
PNA>OM+UOT*'ZPD##]GALX#F'PA(E&,01=OE]IX<J5JC<;G:%WVBCHEQDT 9J\^FV
PHZ\5%N$L.P(4DC;<$5@H]1<43,BN5T%].LIE<ULS0&[1<'HELA-?(\G-MXL248T_
P'[/#>]X;.XW46%;E&= B"$J8S-6>T4'SD85RVA1/XL;)169M/Z[B[*(.RA:S/*["
P@,2BZ(IN[_MI?V&05HO5D7B+ZK15PV[=*(Z]6TT;B3D9,'8=[1B/J4VU)+]':P;L
P,MF(_$MS#Q!*(!QLK#L8C"H:,VE+MZ%^IHG-YH^<E&7^OGE>%BF!N+\(IN=4"QR%
P-[-Y.,E?Q*^!;+!M;6B]?(7%_>A3_S6K*=71@W10BX*L2K)Q[67>HR9L7%"DQC8_
PDK/[_2,K)-)X_+$<:ZFPKUB> 6D\G4H,D>R;!%GJ/J[#+8I>UUD(U4^%9V-1E@E5
P(!MONOL:JSC^R ;RZS"+Y[764>D/[18+M2^L2450/:@DWK'Y4;E;>]U^:449PS6"
P] .?T,@S1-D(7EPF,C*<;2D_1ZKH^Q52-_Q*+=O[*7P*MGSBC9-CC)0J8(]S,Q5(
PS='I01(P.J!^M!_23='22K0:R7 W\G*'C*4HX4$ITC+-O@-^2PJ<0_^2QX!LN_X 
P_[C,KRI40#V"I)6"Z!]4=R"'0P%5>=$Y&W_IN8T35WXD-F;.^E!N69%%P?:\=7/T
PDU1>)YJ9?A+R">2HWOJ[GT+W[;D,]V7Z>0E]"<>(+\/VG&+1C474P<&37&J_R1EI
PY1N/J+F:QGETJA0R6!.I?#\:NA!+I)B*(8ADX<$B<K]E$]:G./P06BJVX <2GK\W
P$OH,Z?P' 0'9>"'%[<=%L42Z?$[_"\C3A "1.R*+N_R%;5B*P6NF6EH@-SQPNNB$
P,9"T]-0&"%%NX2DZ IZ0_AEHX8.MV2-2D@Q-+I+:19%XD;#K&;3*"@S_[Z G5H]9
P=HR_LIT2*1B^>\*M8*7+#\6O=>7>.C*53P?TX3>6Z2>XV#FO9\BYB/KW0&+&2K'@
P_.4-JO$@(:AU42:^Y+>8B#BFB/#5C_T 48XQKX>WCV?,[7=/X(QO0%"2EJ!4>W(P
P<G[]Z-\FKGL!/^)F!+-&O7CB]^Y?\R1G+^:H=DSP':FM?Y[=R2J8^*WY3R ]E/2,
P<JSD;,,06B-="]Z%9='\M4[QH(/F;!125.T9,DP $LUX<WAM(3U]XA#F*S9X9WP*
P]7/O>VAHPI+JM<OR*+7^066M=2D7=1[DC@90R;K;ISS[@]I0G$VJ/FDXOVLGK-]"
PWSV9BRWPDX2;U8*.!G2#EY:VL&5>*A1$[0M7C%+9[(?GG>):@ZAB19TF :=L4Z,J
P#0Z#R <ETL1 R-4K3,5&=+2<$N^G.4;KQ(569"->/.V"Y@Y5>G)/0;&+](;*<"-/
PQ#7%"WK4B?OOQ;4O5UJ'AK9%ZO)@^![X0][+.X?(O]W43XXAG*^@!FFQ2K&%<1$S
PMI,'[SSVR/[^S+ ;!!75L UJXTJ<9NX#^>GWGL=K_-WSD@*Z:4-D_; 9%=Z0J57P
PW^[M2>&G3C)-N]SM@=]M-"T YW8Y"RG)P68'-S X#AOT X\@Y['MIDV2W84A?H0!
PHLG2^T!67 Y-\NT!-)A<>J]@(<C87*.D&J3'RQ^S< 0^ D /TZZ)LP+;<&S9_&D'
P[CWGQ07$]$;VJ3C> L(N#%%I#!N13Y7_>T%81##;DVTLBJIO1F-SU+FT)QBYUA;H
P?ODB[8T Q)\_!;KKHB&=/V&SK_Z\OM3#, J(]28#?^M;N]&PLL;7;B#9:2PH,"T+
P;_9Z:1BS;MG4%L J[5Z0$1$( 0D--.ULL'-A]*SPM64ZUI-Q,]S_'9IWE1R$",T]
P +U9@_H:.E.K.4!KS\"6<A)E_+V@*;3$W+YB6>" _MO:6=X=5*^DLV_9V:C/*KAY
PF656I(K4V>RK+%23XI*04%EU46&FSP3D\(J(I\J]<33-J16X@:7HG/E(,<:EPQ=B
PG<T]IQ(CZWEM/:2\8 R&SB51V6#N*00W!?76D6B0T>G)XC=L[R7X%0RZA0Q91X(,
P;?&=(_&!0T>384&KNV (8[&HX[VNHI]RG3@8S(! DM['J_<.1MM I&53'@TN:Q 0
`endprotected128


